// Benchmark "usb_funct" written by ABC on Thu Oct  8 22:04:27 2020

module usb_funct ( clock, 
    clk_i, rst_i, wb_we_i, wb_stb_i, wb_cyc_i, resume_req_i, phy_clk_pad_i,
    TxReady_pad_i, RxValid_pad_i, RxActive_pad_i, RxError_pad_i,
    usb_vbus_pad_i, \wb_addr_i[0] , \wb_addr_i[1] , \wb_addr_i[2] ,
    \wb_addr_i[3] , \wb_addr_i[4] , \wb_addr_i[5] , \wb_addr_i[6] ,
    \wb_addr_i[7] , \wb_addr_i[8] , \wb_addr_i[9] , \wb_addr_i[10] ,
    \wb_addr_i[11] , \wb_addr_i[12] , \wb_addr_i[13] , \wb_addr_i[14] ,
    \wb_addr_i[15] , \wb_addr_i[16] , \wb_addr_i[17] , \wb_data_i[0] ,
    \wb_data_i[1] , \wb_data_i[2] , \wb_data_i[3] , \wb_data_i[4] ,
    \wb_data_i[5] , \wb_data_i[6] , \wb_data_i[7] , \wb_data_i[8] ,
    \wb_data_i[9] , \wb_data_i[10] , \wb_data_i[11] , \wb_data_i[12] ,
    \wb_data_i[13] , \wb_data_i[14] , \wb_data_i[15] , \wb_data_i[16] ,
    \wb_data_i[17] , \wb_data_i[18] , \wb_data_i[19] , \wb_data_i[20] ,
    \wb_data_i[21] , \wb_data_i[22] , \wb_data_i[23] , \wb_data_i[24] ,
    \wb_data_i[25] , \wb_data_i[26] , \wb_data_i[27] , \wb_data_i[28] ,
    \wb_data_i[29] , \wb_data_i[30] , \wb_data_i[31] , \sram_data_i[0] ,
    \sram_data_i[1] , \sram_data_i[2] , \sram_data_i[3] , \sram_data_i[4] ,
    \sram_data_i[5] , \sram_data_i[6] , \sram_data_i[7] , \sram_data_i[8] ,
    \sram_data_i[9] , \sram_data_i[10] , \sram_data_i[11] ,
    \sram_data_i[12] , \sram_data_i[13] , \sram_data_i[14] ,
    \sram_data_i[15] , \sram_data_i[16] , \sram_data_i[17] ,
    \sram_data_i[18] , \sram_data_i[19] , \sram_data_i[20] ,
    \sram_data_i[21] , \sram_data_i[22] , \sram_data_i[23] ,
    \sram_data_i[24] , \sram_data_i[25] , \sram_data_i[26] ,
    \sram_data_i[27] , \sram_data_i[28] , \sram_data_i[29] ,
    \sram_data_i[30] , \sram_data_i[31] , \dma_ack_i[0] , \dma_ack_i[1] ,
    \dma_ack_i[2] , \dma_ack_i[3] , \dma_ack_i[4] , \dma_ack_i[5] ,
    \dma_ack_i[6] , \dma_ack_i[7] , \dma_ack_i[8] , \dma_ack_i[9] ,
    \dma_ack_i[10] , \dma_ack_i[11] , \dma_ack_i[12] , \dma_ack_i[13] ,
    \dma_ack_i[14] , \dma_ack_i[15] , \DataIn_pad_i[0] , \DataIn_pad_i[1] ,
    \DataIn_pad_i[2] , \DataIn_pad_i[3] , \DataIn_pad_i[4] ,
    \DataIn_pad_i[5] , \DataIn_pad_i[6] , \DataIn_pad_i[7] ,
    \VStatus_pad_i[0] , \VStatus_pad_i[1] , \VStatus_pad_i[2] ,
    \VStatus_pad_i[3] , \VStatus_pad_i[4] , \VStatus_pad_i[5] ,
    \VStatus_pad_i[6] , \VStatus_pad_i[7] , \LineState_pad_i[0] ,
    \LineState_pad_i[1] ,
    \wb_data_o[0] , \wb_data_o[1] , \wb_data_o[2] , \wb_data_o[3] ,
    \wb_data_o[4] , \wb_data_o[5] , \wb_data_o[6] , \wb_data_o[7] ,
    \wb_data_o[8] , \wb_data_o[9] , \wb_data_o[10] , \wb_data_o[11] ,
    \wb_data_o[12] , \wb_data_o[13] , \wb_data_o[14] , \wb_data_o[15] ,
    \wb_data_o[16] , \wb_data_o[17] , \wb_data_o[18] , \wb_data_o[19] ,
    \wb_data_o[20] , \wb_data_o[21] , \wb_data_o[22] , \wb_data_o[23] ,
    \wb_data_o[24] , \wb_data_o[25] , \wb_data_o[26] , \wb_data_o[27] ,
    \wb_data_o[28] , \wb_data_o[29] , \wb_data_o[30] , \wb_data_o[31] ,
    \sram_data_o[0] , \sram_data_o[1] , \sram_data_o[2] , \sram_data_o[3] ,
    \sram_data_o[4] , \sram_data_o[5] , \sram_data_o[6] , \sram_data_o[7] ,
    \sram_data_o[8] , \sram_data_o[9] , \sram_data_o[10] ,
    \sram_data_o[11] , \sram_data_o[12] , \sram_data_o[13] ,
    \sram_data_o[14] , \sram_data_o[15] , \sram_data_o[16] ,
    \sram_data_o[17] , \sram_data_o[18] , \sram_data_o[19] ,
    \sram_data_o[20] , \sram_data_o[21] , \sram_data_o[22] ,
    \sram_data_o[23] , \sram_data_o[24] , \sram_data_o[25] ,
    \sram_data_o[26] , \sram_data_o[27] , \sram_data_o[28] ,
    \sram_data_o[29] , \sram_data_o[30] , \sram_data_o[31] , wb_ack_o,
    inta_o, intb_o, susp_o, phy_rst_pad_o, TxValid_pad_o, XcvSelect_pad_o,
    TermSel_pad_o, SuspendM_pad_o, VControl_Load_pad_o, sram_re_o,
    sram_we_o, \dma_req_o[0] , \dma_req_o[1] , \dma_req_o[2] ,
    \dma_req_o[3] , \dma_req_o[4] , \dma_req_o[5] , \dma_req_o[6] ,
    \dma_req_o[7] , \dma_req_o[8] , \dma_req_o[9] , \dma_req_o[10] ,
    \dma_req_o[11] , \dma_req_o[12] , \dma_req_o[13] , \dma_req_o[14] ,
    \dma_req_o[15] , \DataOut_pad_o[0] , \DataOut_pad_o[1] ,
    \DataOut_pad_o[2] , \DataOut_pad_o[3] , \DataOut_pad_o[4] ,
    \DataOut_pad_o[5] , \DataOut_pad_o[6] , \DataOut_pad_o[7] ,
    \OpMode_pad_o[0] , \OpMode_pad_o[1] , \VControl_pad_o[0] ,
    \VControl_pad_o[1] , \VControl_pad_o[2] , \VControl_pad_o[3] ,
    \sram_adr_o[0] , \sram_adr_o[1] , \sram_adr_o[2] , \sram_adr_o[3] ,
    \sram_adr_o[4] , \sram_adr_o[5] , \sram_adr_o[6] , \sram_adr_o[7] ,
    \sram_adr_o[8] , \sram_adr_o[9] , \sram_adr_o[10] , \sram_adr_o[11] ,
    \sram_adr_o[12] , \sram_adr_o[13] , \sram_adr_o[14]   );
  input  clock;
  input  clk_i, rst_i, wb_we_i, wb_stb_i, wb_cyc_i, resume_req_i,
    phy_clk_pad_i, TxReady_pad_i, RxValid_pad_i, RxActive_pad_i,
    RxError_pad_i, usb_vbus_pad_i, \wb_addr_i[0] , \wb_addr_i[1] ,
    \wb_addr_i[2] , \wb_addr_i[3] , \wb_addr_i[4] , \wb_addr_i[5] ,
    \wb_addr_i[6] , \wb_addr_i[7] , \wb_addr_i[8] , \wb_addr_i[9] ,
    \wb_addr_i[10] , \wb_addr_i[11] , \wb_addr_i[12] , \wb_addr_i[13] ,
    \wb_addr_i[14] , \wb_addr_i[15] , \wb_addr_i[16] , \wb_addr_i[17] ,
    \wb_data_i[0] , \wb_data_i[1] , \wb_data_i[2] , \wb_data_i[3] ,
    \wb_data_i[4] , \wb_data_i[5] , \wb_data_i[6] , \wb_data_i[7] ,
    \wb_data_i[8] , \wb_data_i[9] , \wb_data_i[10] , \wb_data_i[11] ,
    \wb_data_i[12] , \wb_data_i[13] , \wb_data_i[14] , \wb_data_i[15] ,
    \wb_data_i[16] , \wb_data_i[17] , \wb_data_i[18] , \wb_data_i[19] ,
    \wb_data_i[20] , \wb_data_i[21] , \wb_data_i[22] , \wb_data_i[23] ,
    \wb_data_i[24] , \wb_data_i[25] , \wb_data_i[26] , \wb_data_i[27] ,
    \wb_data_i[28] , \wb_data_i[29] , \wb_data_i[30] , \wb_data_i[31] ,
    \sram_data_i[0] , \sram_data_i[1] , \sram_data_i[2] , \sram_data_i[3] ,
    \sram_data_i[4] , \sram_data_i[5] , \sram_data_i[6] , \sram_data_i[7] ,
    \sram_data_i[8] , \sram_data_i[9] , \sram_data_i[10] ,
    \sram_data_i[11] , \sram_data_i[12] , \sram_data_i[13] ,
    \sram_data_i[14] , \sram_data_i[15] , \sram_data_i[16] ,
    \sram_data_i[17] , \sram_data_i[18] , \sram_data_i[19] ,
    \sram_data_i[20] , \sram_data_i[21] , \sram_data_i[22] ,
    \sram_data_i[23] , \sram_data_i[24] , \sram_data_i[25] ,
    \sram_data_i[26] , \sram_data_i[27] , \sram_data_i[28] ,
    \sram_data_i[29] , \sram_data_i[30] , \sram_data_i[31] ,
    \dma_ack_i[0] , \dma_ack_i[1] , \dma_ack_i[2] , \dma_ack_i[3] ,
    \dma_ack_i[4] , \dma_ack_i[5] , \dma_ack_i[6] , \dma_ack_i[7] ,
    \dma_ack_i[8] , \dma_ack_i[9] , \dma_ack_i[10] , \dma_ack_i[11] ,
    \dma_ack_i[12] , \dma_ack_i[13] , \dma_ack_i[14] , \dma_ack_i[15] ,
    \DataIn_pad_i[0] , \DataIn_pad_i[1] , \DataIn_pad_i[2] ,
    \DataIn_pad_i[3] , \DataIn_pad_i[4] , \DataIn_pad_i[5] ,
    \DataIn_pad_i[6] , \DataIn_pad_i[7] , \VStatus_pad_i[0] ,
    \VStatus_pad_i[1] , \VStatus_pad_i[2] , \VStatus_pad_i[3] ,
    \VStatus_pad_i[4] , \VStatus_pad_i[5] , \VStatus_pad_i[6] ,
    \VStatus_pad_i[7] , \LineState_pad_i[0] , \LineState_pad_i[1] ;
  output \wb_data_o[0] , \wb_data_o[1] , \wb_data_o[2] , \wb_data_o[3] ,
    \wb_data_o[4] , \wb_data_o[5] , \wb_data_o[6] , \wb_data_o[7] ,
    \wb_data_o[8] , \wb_data_o[9] , \wb_data_o[10] , \wb_data_o[11] ,
    \wb_data_o[12] , \wb_data_o[13] , \wb_data_o[14] , \wb_data_o[15] ,
    \wb_data_o[16] , \wb_data_o[17] , \wb_data_o[18] , \wb_data_o[19] ,
    \wb_data_o[20] , \wb_data_o[21] , \wb_data_o[22] , \wb_data_o[23] ,
    \wb_data_o[24] , \wb_data_o[25] , \wb_data_o[26] , \wb_data_o[27] ,
    \wb_data_o[28] , \wb_data_o[29] , \wb_data_o[30] , \wb_data_o[31] ,
    \sram_data_o[0] , \sram_data_o[1] , \sram_data_o[2] , \sram_data_o[3] ,
    \sram_data_o[4] , \sram_data_o[5] , \sram_data_o[6] , \sram_data_o[7] ,
    \sram_data_o[8] , \sram_data_o[9] , \sram_data_o[10] ,
    \sram_data_o[11] , \sram_data_o[12] , \sram_data_o[13] ,
    \sram_data_o[14] , \sram_data_o[15] , \sram_data_o[16] ,
    \sram_data_o[17] , \sram_data_o[18] , \sram_data_o[19] ,
    \sram_data_o[20] , \sram_data_o[21] , \sram_data_o[22] ,
    \sram_data_o[23] , \sram_data_o[24] , \sram_data_o[25] ,
    \sram_data_o[26] , \sram_data_o[27] , \sram_data_o[28] ,
    \sram_data_o[29] , \sram_data_o[30] , \sram_data_o[31] , wb_ack_o,
    inta_o, intb_o, susp_o, phy_rst_pad_o, TxValid_pad_o, XcvSelect_pad_o,
    TermSel_pad_o, SuspendM_pad_o, VControl_Load_pad_o, sram_re_o,
    sram_we_o, \dma_req_o[0] , \dma_req_o[1] , \dma_req_o[2] ,
    \dma_req_o[3] , \dma_req_o[4] , \dma_req_o[5] , \dma_req_o[6] ,
    \dma_req_o[7] , \dma_req_o[8] , \dma_req_o[9] , \dma_req_o[10] ,
    \dma_req_o[11] , \dma_req_o[12] , \dma_req_o[13] , \dma_req_o[14] ,
    \dma_req_o[15] , \DataOut_pad_o[0] , \DataOut_pad_o[1] ,
    \DataOut_pad_o[2] , \DataOut_pad_o[3] , \DataOut_pad_o[4] ,
    \DataOut_pad_o[5] , \DataOut_pad_o[6] , \DataOut_pad_o[7] ,
    \OpMode_pad_o[0] , \OpMode_pad_o[1] , \VControl_pad_o[0] ,
    \VControl_pad_o[1] , \VControl_pad_o[2] , \VControl_pad_o[3] ,
    \sram_adr_o[0] , \sram_adr_o[1] , \sram_adr_o[2] , \sram_adr_o[3] ,
    \sram_adr_o[4] , \sram_adr_o[5] , \sram_adr_o[6] , \sram_adr_o[7] ,
    \sram_adr_o[8] , \sram_adr_o[9] , \sram_adr_o[10] , \sram_adr_o[11] ,
    \sram_adr_o[12] , \sram_adr_o[13] , \sram_adr_o[14] ;
  reg \\u0_DataOut_reg[3] , \\u0_DataOut_reg[7] , \\u0_DataOut_reg[2] ,
    \\u0_DataOut_reg[6] , \\u1_u3_token_pid_sel_reg[0] ,
    \\u1_u3_token_pid_sel_reg[1] , u1_u3_no_bufs0_reg,
    \\u1_u3_idin_reg[13] , u1_u3_no_bufs1_reg, \\u1_u1_crc16_reg[15] ,
    \\u1_u1_crc16_reg[1] , \\u1_u3_idin_reg[14] , u1_u3_buffer_done_reg,
    \\u1_u1_crc16_reg[0] , \\u1_u3_idin_reg[12] , \\u1_u3_idin_reg[16] ,
    \\u1_u3_idin_reg[10] , \\u0_DataOut_reg[4] , \\u1_u3_idin_reg[15] ,
    \\u1_u3_idin_reg[11] , \\u0_DataOut_reg[1] , \\u0_DataOut_reg[0] ,
    \\u1_u3_idin_reg[9] , \\u1_u3_idin_reg[6] , u1_u3_buffer_full_reg,
    \\u1_u1_crc16_reg[8] , \\u0_DataOut_reg[5] , \\u1_u3_idin_reg[8] ,
    \\u1_u3_idin_reg[5] , u1_u3_buffer_empty_reg, \\u1_u3_idin_reg[7] ,
    \\u1_u2_adr_cw_reg[11] , \\u1_u2_adr_cw_reg[13] ,
    \\u1_u2_adr_cw_reg[14] , \\u1_u2_adr_cw_reg[5] ,
    \\u1_u2_adr_cw_reg[6] , \\u1_u2_adr_cw_reg[7] , \\u1_u2_adr_cw_reg[8] ,
    \\u1_u2_adr_cw_reg[0] , \\u1_u2_adr_cw_reg[3] , \\u1_u2_adr_cw_reg[2] ,
    \\u1_u2_adr_cw_reg[4] , \\u1_u2_adr_cw_reg[10] ,
    \\u1_u2_adr_cw_reg[12] , \\u1_u2_adr_cw_reg[1] ,
    \\u1_u2_adr_cw_reg[9] , \\u1_u3_idin_reg[4] , u0_TxValid_reg,
    \\u1_u1_crc16_reg[6] , \\u1_u3_idin_reg[3] , \\u1_u1_crc16_reg[2] ,
    \\u1_u1_crc16_reg[3] , \\u1_u1_crc16_reg[4] , \\u1_u1_crc16_reg[7] ,
    \\u1_u1_crc16_reg[9] , \\u1_u1_state_reg[1] , \\u1_u3_idin_reg[2] ,
    \\u1_u3_idin_reg[1] , u1_u1_tx_valid_r_reg, \\u1_u1_state_reg[0] ,
    \\u1_u1_crc16_reg[5] , \\u1_u1_state_reg[4] , u1_u1_tx_valid_r1_reg,
    \\u1_u3_idin_reg[30] , \\u1_u3_idin_reg[0] , u1_u1_send_token_r_reg,
    u1_u1_zero_length_r_reg, \\u1_u3_state_reg[0] , u1_u1_tx_first_r_reg,
    \\u1_u2_sizd_c_reg[10] , \\u1_u2_sizd_c_reg[12] ,
    \\u1_u2_sizd_c_reg[4] , u4_u1_dma_req_r_reg, \\u1_u2_sizd_c_reg[0] ,
    \\u1_u2_sizd_c_reg[11] , \\u1_u2_sizd_c_reg[13] ,
    \\u1_u2_sizd_c_reg[1] , \\u1_u2_sizd_c_reg[2] , \\u1_u2_sizd_c_reg[3] ,
    \\u1_u2_sizd_c_reg[5] , \\u1_u2_sizd_c_reg[6] , \\u1_u2_sizd_c_reg[7] ,
    \\u1_u2_sizd_c_reg[8] , \\u1_u2_sizd_c_reg[9] , u4_u2_dma_req_r_reg,
    u4_u0_dma_req_r_reg, \\u1_u3_new_size_reg[13] , u4_u3_dma_req_r_reg,
    \\u1_u3_state_reg[1] , \\u1_u3_state_reg[4] ,
    \\u1_u2_last_buf_adr_reg[13] , \\u1_u2_last_buf_adr_reg[14] ,
    \\u1_u3_state_reg[2] , u1_u3_send_token_reg,
    u1_u1_send_zero_length_r_reg, \\u1_u3_state_reg[8] ,
    u1_u2_send_zero_length_r_reg, u1_u2_rx_dma_en_r_reg,
    \\u1_u3_new_sizeb_reg[6] , \\u1_u3_new_sizeb_reg[7] ,
    \\u1_u3_new_sizeb_reg[8] , \\u1_u3_new_sizeb_reg[9] ,
    \\u1_u2_last_buf_adr_reg[10] , \\u1_u3_new_sizeb_reg[0] ,
    \\u1_u3_new_sizeb_reg[1] , \\u1_u3_new_sizeb_reg[2] ,
    \\u1_u3_new_sizeb_reg[3] , \\u1_u3_new_sizeb_reg[5] ,
    \\u1_u3_state_reg[3] , \\u1_u3_state_reg[5] , \\u1_u3_state_reg[6] ,
    \\u1_u3_state_reg[7] , \\u1_u3_state_reg[9] ,
    \\u1_u2_last_buf_adr_reg[12] , \\u4_u2_int_stat_reg[2] ,
    \\u4_u3_int_stat_reg[2] , \\u4_u0_int_stat_reg[2] ,
    \\u1_u3_new_sizeb_reg[4] , \\u4_u1_int_stat_reg[2] ,
    \\u1_u3_new_sizeb_reg[10] , \\u1_u2_last_buf_adr_reg[9] ,
    u1_u2_tx_dma_en_r_reg, \\u1_u2_last_buf_adr_reg[11] ,
    \\u1_u3_new_sizeb_reg[13] , \\u1_u3_idin_reg[27] ,
    u4_dma_out_buf_avail_reg, \\u1_u3_new_sizeb_reg[11] ,
    \\u1_u3_new_sizeb_reg[12] , \\u4_u2_int_stat_reg[5] ,
    \\u4_u3_int_stat_reg[5] , \\u4_u0_int_stat_reg[5] ,
    \\u4_u1_int_stat_reg[5] , \\u1_u3_size_next_r_reg[7] ,
    \\u1_u3_size_next_r_reg[6] , \\u1_u3_size_next_r_reg[8] ,
    \\u1_u3_size_next_r_reg[9] , \\u4_int_srcb_reg[2] ,
    u4_u1_dma_req_in_hold2_reg, u1_u3_abort_reg,
    \\u1_u2_last_buf_adr_reg[8] , \\u1_u2_last_buf_adr_reg[6] ,
    \\u1_u2_dout_r_reg[30] , u4_u2_dma_req_in_hold2_reg,
    u4_u0_dma_req_in_hold2_reg, \\u1_u2_dout_r_reg[5] ,
    \\u1_u2_dout_r_reg[27] , \\u1_u2_dout_r_reg[1] ,
    \\u1_u2_dout_r_reg[16] , \\u1_u3_size_next_r_reg[1] ,
    \\u1_u3_size_next_r_reg[3] , \\u1_u3_size_next_r_reg[2] ,
    \\u1_u3_size_next_r_reg[5] , \\u1_u2_adr_cb_reg[0] ,
    \\u1_mfm_cnt_reg[1] , \\u1_u3_idin_reg[25] , \\u1_u3_idin_reg[26] ,
    \\u1_u2_dout_r_reg[0] , \\u1_u2_dout_r_reg[10] ,
    \\u1_u2_dout_r_reg[12] , \\u1_u2_dout_r_reg[11] ,
    \\u1_u2_dout_r_reg[13] , \\u1_u2_dout_r_reg[14] ,
    \\u1_u2_dout_r_reg[15] , \\u1_u2_dout_r_reg[17] ,
    \\u1_u2_dout_r_reg[18] , \\u1_u2_dout_r_reg[19] ,
    \\u1_u2_dout_r_reg[20] , \\u1_u2_dout_r_reg[21] ,
    \\u1_u2_dout_r_reg[22] , \\u1_u2_dout_r_reg[23] ,
    \\u1_u2_dout_r_reg[24] , \\u1_u2_dout_r_reg[25] ,
    \\u1_u2_dout_r_reg[26] , \\u1_u2_dout_r_reg[28] ,
    \\u1_u2_dout_r_reg[29] , \\u1_u2_dout_r_reg[2] ,
    \\u1_u2_dout_r_reg[31] , \\u1_u2_dout_r_reg[3] ,
    \\u1_u2_dout_r_reg[4] , \\u1_u2_dout_r_reg[6] , \\u1_u2_dout_r_reg[7] ,
    \\u1_u2_dout_r_reg[8] , \\u1_u2_dout_r_reg[9] ,
    u0_u0_me_cnt_100_ms_reg, u4_u3_dma_req_in_hold2_reg,
    \\u1_mfm_cnt_reg[3] , \\u1_mfm_cnt_reg[0] ,
    \\u1_u3_size_next_r_reg[0] , \\u1_u3_size_next_r_reg[4] ,
    \\u1_u3_size_next_r_reg[10] , \\u1_u3_size_next_r_reg[11] ,
    \\u1_u3_size_next_r_reg[12] , \\u1_u3_size_next_r_reg[13] ,
    \\u1_u2_adr_cb_reg[2] , \\u1_u3_idin_reg[29] , \\u1_mfm_cnt_reg[2] ,
    u1_u2_word_done_r_reg, \\u1_u2_dtmp_r_reg[12] , u1_u3_int_upid_set_reg,
    \\u1_u2_adr_cb_reg[1] , \\u1_u3_new_size_reg[11] ,
    \\u1_u2_dtmp_r_reg[10] , \\u1_u2_dtmp_r_reg[11] ,
    \\u1_u2_dtmp_r_reg[13] , \\u1_u2_dtmp_r_reg[14] ,
    \\u1_u2_dtmp_r_reg[15] , \\u1_u2_dtmp_r_reg[17] ,
    \\u1_u2_dtmp_r_reg[23] , \\u1_u2_dtmp_r_reg[25] ,
    \\u1_u2_dtmp_r_reg[24] , \\u1_u2_dtmp_r_reg[26] ,
    \\u1_u2_dtmp_r_reg[27] , \\u1_u2_dtmp_r_reg[29] ,
    \\u1_u2_dtmp_r_reg[30] , \\u1_u2_dtmp_r_reg[31] ,
    \\u1_u2_last_buf_adr_reg[4] , \\u1_u2_last_buf_adr_reg[5] ,
    \\u1_u2_dtmp_r_reg[28] , \\u1_u3_new_size_reg[10] ,
    \\u1_u2_dtmp_r_reg[19] , \\u1_u2_dtmp_r_reg[16] ,
    \\u1_u2_sizu_c_reg[5] , u4_nse_err_r_reg, \\u1_u3_idin_reg[24] ,
    \\u1_u2_sizu_c_reg[8] , \\u1_u2_dtmp_r_reg[18] ,
    \\u1_u2_dtmp_r_reg[20] , \\u1_u2_dtmp_r_reg[21] ,
    \\u1_u2_dtmp_r_reg[9] , \\u1_u2_dtmp_r_reg[0] , \\u1_u2_dtmp_r_reg[1] ,
    \\u1_u2_dtmp_r_reg[4] , \\u1_u2_dtmp_r_reg[5] , \\u1_u2_dtmp_r_reg[6] ,
    \\u1_u2_dtmp_r_reg[7] , \\u1_u2_dtmp_r_reg[3] ,
    \\u1_u2_sizu_c_reg[10] , \\u1_u2_sizu_c_reg[1] ,
    \\u1_u2_sizu_c_reg[2] , \\u1_u2_sizu_c_reg[3] , \\u1_u2_sizu_c_reg[4] ,
    \\u1_u2_sizu_c_reg[6] , \\u1_u2_sizu_c_reg[7] , \\u1_u2_sizu_c_reg[9] ,
    u1_u3_buffer_overflow_reg, \\u1_u2_last_buf_adr_reg[7] ,
    \\u1_u2_dtmp_r_reg[22] , \\u1_u2_dtmp_r_reg[2] ,
    \\u1_u2_dtmp_r_reg[8] , u4_u1_dma_out_buf_avail_reg,
    \\u1_frame_no_r_reg[10] , \\u1_frame_no_r_reg[4] ,
    \\u1_frame_no_r_reg[7] , \\u1_frame_no_r_reg[8] ,
    \\u1_u3_idin_reg[23] , \\u1_frame_no_r_reg[9] , u5_wb_ack_o_reg,
    \\u1_u2_sizu_c_reg[0] , u1_u2_wr_last_reg, u1_u3_int_seqerr_set_reg,
    \\u1_u2_last_buf_adr_reg[2] , u1_u2_word_done_reg, u0_u0_T2_wakeup_reg,
    \\u1_frame_no_r_reg[5] , u4_u0_dma_out_buf_avail_reg,
    u4_u2_dma_out_buf_avail_reg, u4_u3_dma_out_buf_avail_reg,
    u1_u3_nse_err_reg, \\u1_hms_cnt_reg[1] , \\u1_frame_no_r_reg[0] ,
    \\u1_frame_no_r_reg[3] , \\u1_frame_no_r_reg[1] ,
    \\u1_frame_no_r_reg[2] , \\u1_frame_no_r_reg[6] , \\u1_hms_cnt_reg[2] ,
    \\u1_hms_cnt_reg[3] , u0_u0_T2_gt_100_uS_reg, u0_u0_T2_gt_1_0_mS_reg,
    u0_u0_T2_gt_1_2_mS_reg, \\u0_u0_me_ps_reg[1] ,
    \\u1_u3_new_size_reg[9] , \\u1_u3_new_size_reg[12] ,
    \\u1_u2_last_buf_adr_reg[3] , \\u0_u0_me_ps2_reg[5] ,
    \\u0_u0_me_cnt_reg[4] , \\u1_hms_cnt_reg[4] , \\u1_u3_idin_reg[21] ,
    \\u0_u0_me_ps2_reg[0] , \\u0_u0_me_ps2_reg[1] , \\u0_u0_me_ps2_reg[2] ,
    \\u0_u0_me_ps2_reg[3] , \\u0_u0_me_ps2_reg[4] , \\u0_u0_me_ps2_reg[6] ,
    \\u0_u0_me_ps2_reg[7] , \\u0_u0_me_ps_reg[0] , \\u0_u0_me_ps_reg[2] ,
    \\u0_u0_me_ps_reg[4] , \\u0_u0_me_ps_reg[5] , \\u0_u0_me_ps_reg[6] ,
    \\u1_u3_idin_reg[20] , \\u0_u0_me_cnt_reg[0] , \\u0_u0_me_cnt_reg[1] ,
    \\u0_u0_me_cnt_reg[2] , \\u0_u0_me_cnt_reg[3] , \\u0_u0_me_cnt_reg[6] ,
    \\u0_u0_me_cnt_reg[7] , \\u0_u0_me_cnt_reg[5] , \\u0_u0_me_ps_reg[3] ,
    \\u0_u0_me_ps_reg[7] , \\u1_u2_state_reg[0] , \\u1_u3_idin_reg[18] ,
    \\u4_u0_buf0_reg[28] , \\u4_u0_buf0_reg[31] , \\u4_u0_buf0_reg[9] ,
    \\u4_u0_buf0_reg[27] , \\u4_u0_buf0_reg[14] , \\u4_u0_buf0_reg[10] ,
    \\u4_u0_buf0_reg[13] , \\u4_u0_buf1_reg[14] , \\u4_u0_buf0_reg[11] ,
    \\u4_u0_buf0_reg[15] , \\u4_u0_buf0_reg[6] , \\u4_u0_buf1_reg[10] ,
    \\u4_u0_buf1_reg[13] , \\u4_u0_buf0_reg[7] , \\u4_u0_buf1_reg[11] ,
    \\u4_u0_buf1_reg[15] , \\u4_u0_buf1_reg[6] , \\u4_u0_buf1_reg[4] ,
    \\u4_u0_buf1_reg[5] , \\u4_u0_buf1_reg[7] , \\u1_hms_cnt_reg[0] ,
    \\u1_u3_idin_reg[19] , \\u1_u3_new_size_reg[5] , \\u4_u0_buf1_reg[28] ,
    \\u4_u0_buf1_reg[31] , \\u1_u2_state_reg[3] , \\u4_u0_buf0_reg[0] ,
    \\u4_u0_buf0_reg[18] , \\u4_u0_buf0_reg[19] , \\u4_u0_buf0_reg[1] ,
    \\u4_u0_buf0_reg[20] , \\u4_u0_buf0_reg[21] , \\u4_u0_buf0_reg[23] ,
    \\u4_u0_buf0_reg[24] , \\u4_u0_buf0_reg[25] , \\u4_u0_buf0_reg[26] ,
    \\u4_u0_buf0_reg[30] , \\u4_u0_buf0_reg[3] , \\u4_u0_buf0_reg[8] ,
    \\u4_u1_buf0_reg[28] , \\u4_u1_buf0_reg[31] , u1_u3_match_r_reg,
    \\u1_u3_new_size_reg[8] , u5_wb_ack_s2_reg, \\u1_u3_new_size_reg[7] ,
    \\u4_u1_buf0_reg[8] , \\u4_u1_buf1_reg[6] , \\u4_u2_dma_in_cnt_reg[9] ,
    \\u4_u3_dma_in_cnt_reg[9] , \\u4_u0_buf1_reg[3] ,
    \\u1_u2_last_buf_adr_reg[1] , \\u4_u1_buf0_reg[6] ,
    \\u4_u1_buf0_reg[14] , \\u4_u1_buf0_reg[10] , \\u4_u1_buf0_reg[13] ,
    \\u4_u1_buf1_reg[14] , \\u4_u1_buf0_reg[11] , \\u4_u1_buf0_reg[15] ,
    \\u4_u1_buf1_reg[10] , \\u4_u1_buf1_reg[13] , \\u4_u1_buf0_reg[7] ,
    \\u4_u1_buf1_reg[11] , \\u4_u1_buf1_reg[15] , \\u4_u1_buf1_reg[4] ,
    \\u4_u1_buf1_reg[7] , \\u4_u1_buf1_reg[5] , \\u4_u0_buf1_reg[29] ,
    \\u4_u0_buf1_reg[21] , \\u4_u0_dma_in_cnt_reg[9] ,
    \\u4_u1_dma_in_cnt_reg[9] , \\u4_u0_dma_in_cnt_reg[11] ,
    \\u1_u0_state_reg[2] , \\u4_u0_dma_out_cnt_reg[11] ,
    \\u4_u0_dma_out_cnt_reg[9] , u4_dma_in_buf_sz1_reg,
    \\u4_u0_dma_in_cnt_reg[7] , \\u4_u0_dma_in_cnt_reg[6] ,
    \\u4_u0_dma_out_cnt_reg[6] , \\u4_u0_buf1_reg[0] ,
    \\u4_u0_buf1_reg[12] , \\u4_u0_buf1_reg[16] , \\u4_u0_buf1_reg[17] ,
    \\u4_u0_buf1_reg[19] , \\u4_u0_buf1_reg[1] , \\u4_u0_buf1_reg[20] ,
    \\u4_u0_buf1_reg[22] , \\u4_u0_buf1_reg[24] , \\u4_u0_buf1_reg[25] ,
    \\u4_u0_buf1_reg[23] , \\u4_u0_buf1_reg[27] , \\u4_u0_buf1_reg[26] ,
    \\u4_u0_buf1_reg[2] , \\u4_u0_buf1_reg[30] , \\u4_u0_buf1_reg[8] ,
    \\u4_u0_buf1_reg[9] , \\u4_u1_buf1_reg[28] , \\u4_u1_buf1_reg[31] ,
    \\u4_u0_dma_in_cnt_reg[0] , \\u1_u2_state_reg[4] ,
    \\u4_u0_dma_out_cnt_reg[0] , \\u4_u0_dma_out_cnt_reg[1] ,
    \\u4_u0_dma_out_cnt_reg[2] , \\u4_u0_dma_out_cnt_reg[3] ,
    \\u4_u1_buf0_reg[16] , \\u4_u1_buf0_reg[18] , \\u4_u1_buf0_reg[19] ,
    \\u4_u1_buf0_reg[1] , \\u4_u1_buf0_reg[20] , \\u4_u1_buf0_reg[21] ,
    \\u4_u1_buf0_reg[23] , \\u4_u1_buf0_reg[24] , \\u4_u1_buf0_reg[25] ,
    \\u4_u1_buf0_reg[27] , \\u4_u1_buf0_reg[30] , \\u4_u1_buf0_reg[3] ,
    \\u4_u1_buf0_reg[9] , \\u4_u2_buf0_reg[28] , \\u4_u2_buf0_reg[31] ,
    u1_frame_no_same_reg, \\u4_u0_buf1_reg[18] , \\u1_u3_new_size_reg[6] ,
    \\u4_u1_buf0_reg[26] , \\u1_sof_time_reg[2] , u5_wb_ack_s1a_reg,
    \\u4_u0_buf0_reg[2] , \\u4_u2_buf0_reg[8] , \\u4_u3_buf0_reg[31] ,
    \\u4_u0_buf0_reg[22] , \\u4_u2_buf0_reg[12] , \\u4_u1_buf1_reg[1] ,
    \\u4_u0_dma_out_cnt_reg[8] , \\u4_u0_dma_out_cnt_reg[4] ,
    \\u4_u1_buf1_reg[9] , \\u4_u2_buf0_reg[19] , \\u4_u1_buf1_reg[27] ,
    \\u4_u1_buf1_reg[23] , \\u4_u0_buf0_reg[5] , \\u1_sof_time_reg[6] ,
    \\u4_u2_buf0_reg[6] , \\u4_u2_buf0_reg[11] , \\u4_u2_buf0_reg[10] ,
    \\u4_u2_buf0_reg[14] , \\u4_u2_buf0_reg[13] , \\u4_u2_buf1_reg[14] ,
    \\u4_u2_buf0_reg[15] , \\u4_u2_buf1_reg[10] , \\u4_u2_buf1_reg[13] ,
    \\u4_u0_buf0_reg[4] , \\u4_u2_buf0_reg[7] , \\u4_u2_buf1_reg[11] ,
    \\u4_u2_buf1_reg[6] , \\u4_u2_buf1_reg[4] , \\u4_u2_buf1_reg[5] ,
    \\u4_u2_buf1_reg[7] , \\u1_sof_time_reg[11] ,
    \\u4_u0_dma_in_cnt_reg[8] , \\u1_sof_time_reg[7] ,
    \\u4_u1_dma_in_cnt_reg[11] , \\u1_sof_time_reg[0] ,
    \\u4_u0_dma_in_cnt_reg[10] , \\u4_u1_dma_out_cnt_reg[11] ,
    \\u4_u1_dma_out_cnt_reg[9] , \\u1_sof_time_reg[10] ,
    \\u1_sof_time_reg[1] , \\u1_sof_time_reg[3] , \\u1_sof_time_reg[4] ,
    \\u1_sof_time_reg[5] , \\u1_sof_time_reg[9] , \\u1_sof_time_reg[8] ,
    \\u4_u0_dma_in_cnt_reg[5] , \\u4_u0_dma_out_cnt_reg[10] ,
    \\u4_u0_dma_out_cnt_reg[7] , \\u4_u1_dma_in_cnt_reg[7] ,
    \\u4_u0_dma_in_cnt_reg[4] , \\u4_u1_dma_in_cnt_reg[6] ,
    \\u4_u1_dma_out_cnt_reg[6] , \\u4_u1_buf1_reg[0] ,
    \\u4_u1_buf1_reg[12] , \\u4_u1_buf1_reg[16] , \\u4_u1_buf1_reg[17] ,
    \\u4_u1_buf1_reg[18] , \\u4_u1_buf1_reg[19] , \\u4_u1_buf1_reg[20] ,
    \\u4_u1_buf1_reg[21] , \\u4_u1_buf1_reg[22] , \\u4_u1_buf1_reg[24] ,
    \\u4_u1_buf1_reg[25] , \\u4_u1_buf1_reg[26] , \\u4_u1_buf1_reg[2] ,
    \\u4_u1_buf1_reg[30] , \\u4_u1_buf1_reg[29] , \\u4_u1_buf1_reg[3] ,
    \\u4_u1_buf1_reg[8] , \\u4_u2_buf1_reg[28] , \\u4_u2_buf1_reg[31] ,
    \\u4_u1_dma_in_cnt_reg[0] , \\u4_u0_dma_in_cnt_reg[1] ,
    \\u4_u0_dma_in_cnt_reg[2] , \\u4_u0_dma_in_cnt_reg[3] ,
    \\u4_u0_dma_out_cnt_reg[5] , \\u4_u1_dma_out_cnt_reg[0] ,
    \\u4_u1_dma_out_cnt_reg[1] , \\u4_u1_dma_out_cnt_reg[2] ,
    \\u4_u1_dma_out_cnt_reg[3] , \\u4_u3_buf0_reg[28] ,
    \\u4_u0_buf0_reg[12] , \\u4_u0_buf0_reg[16] , \\u4_u0_buf0_reg[17] ,
    \\u4_u0_buf0_reg[29] , \\u4_u2_buf0_reg[0] , \\u4_u2_buf0_reg[16] ,
    \\u4_u2_buf0_reg[17] , \\u4_u2_buf0_reg[18] , \\u4_u2_buf0_reg[20] ,
    \\u4_u2_buf0_reg[22] , \\u4_u2_buf0_reg[24] , \\u4_u2_buf0_reg[25] ,
    \\u4_u2_buf0_reg[29] , \\u4_u2_buf0_reg[1] , \\u4_u2_buf0_reg[30] ,
    \\u4_u2_buf0_reg[3] , \\u4_u2_buf1_reg[15] ,
    \\u4_u1_dma_in_cnt_reg[8] , \\u4_u1_buf0_reg[2] ,
    \\u4_u3_int_stat_reg[0] , \\u4_u1_buf0_reg[22] , \\u4_u2_buf1_reg[3] ,
    \\u4_u2_buf1_reg[20] , \\u4_u2_buf1_reg[27] , \\u4_u2_buf1_reg[24] ,
    \\u4_u1_dma_out_cnt_reg[4] , \\u4_u3_buf0_reg[29] ,
    \\u4_u2_buf1_reg[17] , \\u4_u3_buf0_reg[25] , \\u1_u3_new_size_reg[3] ,
    \\u4_u3_buf0_reg[21] , \\u4_u3_buf0_reg[5] , \\u4_u1_buf0_reg[5] ,
    \\u4_u1_dma_in_cnt_reg[5] , \\u4_u3_buf0_reg[6] ,
    \\u4_u3_buf0_reg[10] , \\u4_u2_dma_out_cnt_reg[9] ,
    \\u4_u3_buf0_reg[14] , \\u4_u3_buf0_reg[13] , \\u4_u3_buf0_reg[11] ,
    \\u4_u3_buf0_reg[15] , \\u4_u3_buf0_reg[4] , \\u4_u3_buf0_reg[7] ,
    \\u4_u1_buf0_reg[4] , \\u4_u1_dma_out_cnt_reg[8] ,
    \\u5_wb_data_o_reg[1] , \\u4_u1_dma_in_cnt_reg[10] ,
    \\u4_u2_dma_out_cnt_reg[11] , \\u4_u1_dma_out_cnt_reg[10] ,
    \\u4_u1_dma_out_cnt_reg[7] , \\u4_u2_dma_in_cnt_reg[7] ,
    \\u4_u1_dma_in_cnt_reg[4] , \\u4_u2_dma_out_cnt_reg[6] ,
    \\u4_u2_dma_in_cnt_reg[6] , \\u4_u2_buf1_reg[0] ,
    \\u4_u2_buf1_reg[12] , \\u4_u2_buf1_reg[16] , \\u4_u2_buf1_reg[18] ,
    \\u4_u2_buf1_reg[19] , \\u4_u2_buf1_reg[1] , \\u4_u2_buf1_reg[22] ,
    \\u4_u2_buf1_reg[23] , \\u4_u2_buf1_reg[21] , \\u4_u2_buf1_reg[26] ,
    \\u4_u2_buf1_reg[25] , \\u4_u2_buf1_reg[29] , \\u4_u2_buf1_reg[2] ,
    \\u4_u2_buf1_reg[30] , \\u4_u2_buf1_reg[8] , \\u4_u2_buf1_reg[9] ,
    \\u4_u2_dma_in_cnt_reg[0] , \\u4_u1_dma_in_cnt_reg[2] ,
    \\u4_u1_dma_out_cnt_reg[5] , \\u4_u2_dma_out_cnt_reg[1] ,
    \\u4_u2_dma_out_cnt_reg[2] , \\u4_u2_dma_out_cnt_reg[3] ,
    \\u4_u2_int_stat_reg[0] , \\u4_u3_buf0_reg[0] ,
    \\u4_u2_dma_out_cnt_reg[0] , \\u4_u3_buf0_reg[16] ,
    \\u4_u3_buf0_reg[17] , \\u4_u3_buf0_reg[18] , \\u4_u3_buf0_reg[19] ,
    \\u4_u3_buf0_reg[1] , \\u4_u3_buf0_reg[20] , \\u4_u3_buf0_reg[12] ,
    \\u4_u3_buf0_reg[23] , \\u4_u3_buf0_reg[24] , \\u4_u3_buf0_reg[22] ,
    \\u4_u3_buf0_reg[27] , \\u4_u3_buf0_reg[26] , \\u4_u3_buf0_reg[2] ,
    \\u4_u3_buf0_reg[30] , \\u4_u3_buf0_reg[3] , \\u4_u3_buf0_reg[8] ,
    \\u4_u3_buf0_reg[9] , \\u4_u1_buf0_reg[0] , \\u4_u1_buf0_reg[12] ,
    \\u4_u1_buf0_reg[17] , \\u4_u0_int_stat_reg[0] , \\u4_u1_buf0_reg[29] ,
    \\u4_u1_int_stat_reg[0] , \\u4_u1_dma_in_cnt_reg[1] ,
    \\u5_state_reg[0] , \\u1_u3_new_size_reg[4] ,
    \\u4_u2_dma_in_cnt_reg[11] , \\u4_u1_dma_in_cnt_reg[3] ,
    \\u4_u2_dma_in_cnt_reg[8] , \\u4_u3_buf1_reg[7] ,
    u1_u3_pid_seq_err_reg, \\u4_u2_buf0_reg[2] ,
    \\u4_u2_dma_out_cnt_reg[4] , \\u4_u3_buf1_reg[5] ,
    \\u4_u2_buf0_reg[26] , u5_wb_ack_s1_reg, \\u4_u2_dma_out_cnt_reg[7] ,
    \\u4_u2_buf0_reg[4] , \\u4_u3_buf1_reg[6] , \\u5_state_reg[5] ,
    \\u4_u3_buf1_reg[14] , \\u4_u3_buf1_reg[10] , \\u4_u3_buf1_reg[13] ,
    \\u4_u3_buf1_reg[11] , \\u4_u3_buf1_reg[15] , \\u4_u2_buf0_reg[5] ,
    \\u4_u3_buf1_reg[4] , \\u4_u2_dma_out_cnt_reg[8] ,
    \\u5_wb_data_o_reg[3] , \\u4_int_srcb_reg[0] ,
    \\u4_u2_dma_in_cnt_reg[10] , u2_wack_r_reg, \\u1_u0_state_reg[3] ,
    \\u4_u2_dma_in_cnt_reg[5] , \\u4_u2_dma_out_cnt_reg[10] ,
    \\u4_u2_dma_in_cnt_reg[4] , \\u4_u3_buf1_reg[28] ,
    \\u4_u3_buf1_reg[31] , \\u4_u2_dma_in_cnt_reg[2] ,
    \\u4_u2_dma_in_cnt_reg[3] , \\u4_u2_dma_out_cnt_reg[5] ,
    \\u4_u2_buf0_reg[21] , \\u4_u2_buf0_reg[23] , \\u4_u2_buf0_reg[27] ,
    \\u4_u2_buf0_reg[9] , \\u1_u2_state_reg[2] , \\u5_wb_data_o_reg[0] ,
    \\u4_u2_dma_in_cnt_reg[1] , \\u4_u3_dma_out_cnt_reg[9] ,
    \\u4_u3_dma_in_cnt_reg[10] , \\u4_u3_dma_in_cnt_reg[11] ,
    \\u5_wb_data_o_reg[2] , \\u4_u3_buf1_reg[25] , \\u4_u3_buf1_reg[21] ,
    \\u4_u3_dma_out_cnt_reg[3] , \\u4_u3_buf1_reg[0] ,
    \\u4_u3_buf1_reg[18] , u1_u3_buf1_st_max_reg, \\u1_u3_new_size_reg[2] ,
    \\u4_u3_dma_out_cnt_reg[11] , \\u4_u3_dma_in_cnt_reg[7] , u4_u0_r1_reg,
    \\u5_state_reg[4] , \\u4_u3_dma_in_cnt_reg[6] ,
    \\u4_u3_dma_out_cnt_reg[6] , \\u4_u3_buf1_reg[12] ,
    \\u4_u3_buf1_reg[16] , \\u4_u3_buf1_reg[17] , \\u4_u3_buf1_reg[19] ,
    \\u4_u3_buf1_reg[1] , \\u4_u3_buf1_reg[20] , \\u4_u3_buf1_reg[22] ,
    \\u4_u3_buf1_reg[23] , \\u4_u3_buf1_reg[24] , \\u4_u3_buf1_reg[27] ,
    \\u4_u3_buf1_reg[26] , \\u4_u3_buf1_reg[30] , \\u4_u3_buf1_reg[2] ,
    \\u4_u3_buf1_reg[9] , \\u4_u3_buf1_reg[8] , \\u1_u0_state_reg[0] ,
    \\u1_u0_state_reg[1] , \\u4_u3_dma_in_cnt_reg[0] ,
    \\u4_u3_dma_out_cnt_reg[1] , \\u4_u3_dma_out_cnt_reg[2] ,
    \\u4_u3_dma_out_cnt_reg[0] , \\u1_u2_last_buf_adr_reg[0] ,
    \\u5_state_reg[1] , \\u4_u3_buf1_reg[3] , \\u4_u3_buf1_reg[29] ,
    u1_clr_sof_time_reg, u1_frame_no_we_r_reg, \\u4_u3_dma_out_cnt_reg[5] ,
    \\u4_u3_dma_in_cnt_reg[3] , \\u4_u3_dma_out_cnt_reg[8] ,
    \\u4_u3_dma_out_cnt_reg[4] , u4_u1_r1_reg, \\u4_u3_dma_in_cnt_reg[8] ,
    u4_u2_r1_reg, \\u4_u3_dma_in_cnt_reg[5] , \\u4_u3_dma_out_cnt_reg[10] ,
    \\u5_state_reg[2] , \\u4_u3_dma_in_cnt_reg[4] ,
    \\u4_u3_dma_in_cnt_reg[1] , \\u4_u3_dma_in_cnt_reg[2] ,
    \\u4_u3_dma_out_cnt_reg[7] , u4_u3_r1_reg, \\u1_u0_crc16_sum_reg[1] ,
    \\u1_u0_crc16_sum_reg[11] , u0_u0_T1_gt_2_5_uS_reg, u1_u3_to_large_reg,
    \\u1_u3_new_size_reg[1] , \\u1_u0_crc16_sum_reg[15] ,
    \\u4_int_srcb_reg[6] , \\u1_u0_crc16_sum_reg[0] ,
    \\u1_u0_crc16_sum_reg[10] , \\u1_u0_crc16_sum_reg[12] ,
    \\u1_u0_crc16_sum_reg[14] , \\u1_u0_crc16_sum_reg[3] ,
    \\u1_u0_crc16_sum_reg[4] , \\u1_u0_crc16_sum_reg[5] ,
    \\u1_u0_crc16_sum_reg[7] , \\u1_u0_crc16_sum_reg[8] ,
    \\u1_u0_crc16_sum_reg[9] , \\u1_u3_adr_r_reg[10] ,
    \\u1_u3_adr_r_reg[13] , \\u1_u3_adr_r_reg[3] , \\u1_u3_adr_r_reg[4] ,
    u1_u3_to_small_reg, \\u1_u0_crc16_sum_reg[13] ,
    \\u1_u0_crc16_sum_reg[6] , \\u1_u0_crc16_sum_reg[2] ,
    \\u1_u1_crc16_reg[14] , \\u4_buf1_reg[25] , \\u4_buf1_reg[29] ,
    \\u4_csr_reg[1] , \\u4_buf1_reg[21] , \\u4_buf1_reg[14] ,
    \\u4_dout_reg[1] , \\u4_buf1_reg[18] , \\u4_csr_reg[5] ,
    \\u4_buf0_reg[3] , \\u4_buf0_reg[7] , \\u4_buf1_reg[10] ,
    \\u4_csr_reg[9] , \\u0_u0_state_reg[13] , \\u0_u0_idle_cnt1_reg[1] ,
    \\u4_buf0_reg[29] , \\u0_u0_ps_cnt_reg[2] , \\u0_u0_idle_cnt1_reg[4] ,
    \\u0_u0_idle_cnt1_reg[6] , \\u0_u0_idle_cnt1_reg[7] ,
    \\u4_csr_reg[30] , \\u4_buf0_reg[30] , \\u5_wb_data_o_reg[23] ,
    \\u4_buf0_reg[21] , \\u4_csr_reg[27] , \\u4_buf0_reg[25] ,
    \\u0_u0_state_reg[11] , \\u1_u3_adr_r_reg[12] , \\u1_u3_adr_r_reg[16] ,
    u1_u3_buf0_st_max_reg, \\u1_u1_crc16_reg[10] , \\u1_u1_crc16_reg[13] ,
    \\u1_u1_crc16_reg[12] , \\u4_csr_reg[23] , \\u5_wb_data_o_reg[22] ,
    \\u5_wb_data_o_reg[7] , \\u0_u0_idle_cnt1_reg[3] ,
    \\u5_wb_data_o_reg[8] , u0_u0_T1_gt_3_0_mS_reg, \\u4_int_srcb_reg[3] ,
    \\u0_u0_idle_cnt1_reg[0] , \\u0_u0_idle_cnt1_reg[2] , u1_u0_rxv2_reg,
    \\u0_u0_idle_cnt1_reg[5] , \\u0_u0_ps_cnt_reg[0] ,
    \\u0_u0_ps_cnt_reg[1] , \\u0_u0_ps_cnt_reg[3] , resume_req_r_reg,
    \\u4_csr_reg[12] , \\u4_csr_reg[15] , \\u4_csr_reg[17] ,
    \\u4_csr_reg[22] , \\u4_csr_reg[24] , \\u4_csr_reg[25] ,
    \\u4_csr_reg[26] , \\u4_csr_reg[28] , \\u4_csr_reg[29] ,
    \\u4_csr_reg[2] , \\u4_csr_reg[31] , \\u4_csr_reg[3] ,
    \\u4_csr_reg[4] , \\u4_csr_reg[6] , \\u4_csr_reg[7] , \\u4_csr_reg[8] ,
    \\u4_buf0_reg[0] , \\u4_buf0_reg[10] , \\u4_buf0_reg[11] ,
    \\u4_buf0_reg[12] , \\u4_buf0_reg[13] , \\u4_buf0_reg[15] ,
    \\u4_buf0_reg[16] , \\u4_buf0_reg[17] , \\u4_buf0_reg[19] ,
    \\u4_buf0_reg[1] , \\u4_buf0_reg[20] , \\u4_buf0_reg[22] ,
    \\u4_buf0_reg[23] , \\u4_buf0_reg[24] , \\u4_buf0_reg[26] ,
    \\u4_buf0_reg[27] , \\u4_buf0_reg[28] , \\u4_buf0_reg[2] ,
    \\u4_buf0_reg[31] , \\u4_buf0_reg[4] , \\u4_buf0_reg[5] ,
    \\u4_buf0_reg[6] , \\u4_buf0_reg[8] , \\u4_buf0_reg[9] ,
    \\u4_buf1_reg[0] , \\u4_buf1_reg[11] , \\u4_buf1_reg[12] ,
    \\u4_buf1_reg[13] , \\u4_buf1_reg[15] , \\u4_buf1_reg[16] ,
    \\u4_buf1_reg[17] , \\u4_buf1_reg[19] , \\u4_buf1_reg[1] ,
    \\u4_buf1_reg[20] , \\u4_buf1_reg[22] , \\u4_buf1_reg[23] ,
    \\u4_buf1_reg[24] , \\u4_buf1_reg[26] , \\u4_buf1_reg[27] ,
    \\u4_buf1_reg[28] , \\u4_buf1_reg[2] , \\u4_buf1_reg[30] ,
    \\u4_buf1_reg[31] , \\u4_buf1_reg[4] , \\u4_buf1_reg[5] ,
    \\u4_buf1_reg[6] , \\u4_buf1_reg[8] , \\u4_buf1_reg[9] ,
    \\u4_csr_reg[0] , \\u4_csr_reg[11] , \\u4_u0_uc_bsel_reg[0] ,
    \\u4_u0_uc_bsel_reg[1] , \\u4_u0_uc_dpd_reg[0] ,
    \\u1_u3_adr_r_reg[11] , \\u1_u3_adr_r_reg[14] , \\u1_u3_adr_r_reg[15] ,
    \\u1_u3_adr_r_reg[6] , \\u1_u3_adr_r_reg[7] , \\u1_u3_adr_r_reg[8] ,
    \\u4_buf0_reg[14] , \\u4_buf0_reg[18] , u0_u0_T1_gt_5_0_mS_reg,
    \\u4_csr_reg[16] , u1_u2_rx_data_valid_r_reg, \\u1_u3_adr_r_reg[9] ,
    \\u4_u0_uc_dpd_reg[1] , \\u4_csr_reg[10] , \\u1_u1_crc16_reg[11] ,
    \\u4_buf1_reg[7] , \\u4_buf1_reg[3] , \\u1_u0_d1_reg[0] ,
    \\u5_wb_data_o_reg[25] , \\u4_dout_reg[0] , \\u1_u0_d1_reg[4] ,
    \\u4_dout_reg[2] , \\u4_dout_reg[3] , \\u1_u0_d0_reg[4] ,
    \\u5_wb_data_o_reg[26] , \\u1_u0_d0_reg[1] , \\u1_u0_d0_reg[3] ,
    \\u4_u1_int_stat_reg[4] , \\u4_u3_int_stat_reg[4] , u4_crc5_err_r_reg,
    \\u1_u3_next_dpid_reg[0] , \\u1_u3_adr_r_reg[0] ,
    u4_u1_dma_in_buf_sz1_reg, u4_u0_dma_in_buf_sz1_reg,
    u4_u3_dma_in_buf_sz1_reg, u4_u2_dma_in_buf_sz1_reg, u0_u0_TermSel_reg,
    \\u4_int_srcb_reg[5] , \\u5_wb_data_o_reg[4] ,
    \\u4_u2_int_stat_reg[4] , \\u4_u0_int_stat_reg[4] ,
    \\u5_wb_data_o_reg[16] , \\u5_wb_data_o_reg[24] ,
    \\u5_wb_data_o_reg[28] , \\u5_wb_data_o_reg[21] ,
    \\u5_wb_data_o_reg[20] , \\u5_wb_data_o_reg[19] ,
    \\u5_wb_data_o_reg[6] , \\u5_wb_data_o_reg[5] ,
    \\u5_wb_data_o_reg[18] , \\u5_wb_data_o_reg[17] ,
    \\u4_int_srcb_reg[4] , \\u0_u0_state_reg[1] , u1_u0_rxv1_reg,
    \\u1_u0_d0_reg[0] , \\u0_u0_chirp_cnt_reg[1] , \\u1_u0_d0_reg[2] ,
    \\u0_u0_chirp_cnt_reg[2] , \\u1_u0_d0_reg[5] , \\u1_u0_d0_reg[6] ,
    \\u1_u0_d0_reg[7] , \\u1_u0_d1_reg[1] , \\u1_u0_d1_reg[2] ,
    \\u1_u0_d1_reg[3] , \\u1_u0_d1_reg[5] , \\u1_u0_d1_reg[6] ,
    \\u1_u0_d1_reg[7] , \\u1_u0_d2_reg[1] , \\u1_u0_d2_reg[2] ,
    \\u1_u0_d2_reg[3] , \\u1_u0_d2_reg[5] , \\u1_u0_d2_reg[6] ,
    \\u1_u0_d2_reg[7] , \\u0_u0_state_reg[12] , \\u4_u1_uc_bsel_reg[0] ,
    \\u4_u1_uc_dpd_reg[0] , \\u1_u3_adr_r_reg[2] , \\u4_u1_uc_bsel_reg[1] ,
    \\u4_u1_uc_dpd_reg[1] , \\u1_u0_d2_reg[0] , \\u1_u0_d2_reg[4] ,
    \\u1_u3_adr_r_reg[5] , \\u1_u3_adr_r_reg[1] ,
    \\u4_u3_dma_out_left_reg[10] , \\u4_u0_dma_out_left_reg[10] ,
    \\u4_u1_dma_out_left_reg[10] , \\u4_u2_dma_out_left_reg[10] ,
    \\u5_wb_data_o_reg[30] , \\u5_wb_data_o_reg[31] ,
    \\u1_u3_idin_reg[17] , \\u0_u0_state_reg[9] , \\u5_wb_data_o_reg[27] ,
    \\u5_wb_data_o_reg[29] , \\u4_u3_int_stat_reg[3] ,
    \\u4_u0_int_stat_reg[3] , \\u4_u1_int_stat_reg[3] ,
    u0_u0_T1_st_3_0_mS_reg, \\u5_wb_data_o_reg[11] ,
    \\u5_wb_data_o_reg[9] , \\u0_u0_chirp_cnt_reg[0] ,
    \\u5_wb_data_o_reg[12] , \\u4_u0_int_stat_reg[6] ,
    \\u0_u0_state_reg[4] , \\u4_u2_uc_bsel_reg[0] ,
    \\u4_u2_uc_bsel_reg[1] , \\u4_u2_uc_dpd_reg[0] ,
    \\u4_u2_int_stat_reg[3] , \\u0_u0_state_reg[3] ,
    \\u5_wb_data_o_reg[10] , \\u4_u2_uc_dpd_reg[1] , u1_u0_data_valid0_reg,
    u0_u0_XcvSelect_reg, \\u0_u0_OpMode_reg[1] , \\u4_int_srcb_reg[8] ,
    \\u4_u3_dma_out_left_reg[9] , \\u4_u0_dma_out_left_reg[9] ,
    \\u4_u1_dma_out_left_reg[9] , \\u4_u2_dma_out_left_reg[9] ,
    \\u1_u3_this_dpid_reg[0] , \\u1_u3_next_dpid_reg[1] ,
    \\u0_u0_state_reg[10] , \\u0_u0_OpMode_reg[0] , \\u4_int_srcb_reg[7] ,
    \\u4_int_srcb_reg[1] , \\u5_wb_data_o_reg[13] ,
    \\u5_wb_data_o_reg[15] , \\u4_u1_int_stat_reg[6] ,
    \\u4_u0_int_stat_reg[1] , \\u4_u3_uc_bsel_reg[0] ,
    \\u4_u3_uc_bsel_reg[1] , \\u4_u3_uc_dpd_reg[0] , \\u0_u0_state_reg[6] ,
    u1_u3_buf1_set_reg, \\u1_u3_adr_reg[0] , \\u1_u3_adr_reg[1] ,
    \\u1_u3_adr_reg[2] , \\u1_u3_adr_reg[12] , \\u1_u3_adr_reg[13] ,
    \\u1_u3_adr_reg[14] , \\u1_u3_adr_reg[15] , \\u1_u3_adr_reg[16] ,
    \\u1_u3_adr_reg[3] , \\u1_u3_adr_reg[4] , \\u1_u3_adr_reg[5] ,
    \\u1_u3_adr_reg[6] , \\u1_u3_adr_reg[7] , \\u1_u3_adr_reg[8] ,
    \\u1_u3_adr_reg[9] , \\u1_u3_adr_reg[10] , \\u1_u3_adr_reg[11] ,
    \\u4_u3_uc_dpd_reg[1] , u4_intb_reg, \\u1_u3_this_dpid_reg[1] ,
    \\u1_u0_token0_reg[6] , u1_u2_send_data_r_reg, \\u0_u0_state_reg[5] ,
    u4_inta_reg, \\u0_u0_state_reg[14] , \\u4_u0_csr0_reg[2] ,
    \\u4_u0_csr0_reg[4] , \\u4_u0_csr1_reg[1] , \\u4_u0_csr1_reg[2] ,
    \\u4_u0_csr1_reg[3] , \\u4_u1_csr0_reg[2] , \\u4_u1_csr0_reg[5] ,
    \\u4_u1_csr0_reg[9] , \\u4_u1_csr1_reg[10] , \\u4_u2_csr0_reg[0] ,
    \\u4_u2_csr0_reg[2] , \\u4_u2_csr0_reg[6] , \\u4_u2_csr0_reg[9] ,
    \\u4_u2_int_stat_reg[1] , \\u4_u1_buf0_orig_reg[30] ,
    \\u4_u1_int_stat_reg[1] , u0_u0_usb_suspend_reg,
    \\u1_u0_token0_reg[0] , \\u1_u0_token0_reg[1] , \\u1_u0_token0_reg[3] ,
    \\u1_u0_token0_reg[4] , \\u1_u0_token0_reg[5] , \\u1_u0_token0_reg[7] ,
    \\u0_u0_state_reg[7] , \\u0_u0_state_reg[2] , u1_u3_buf0_set_reg,
    \\u4_u2_int_stat_reg[6] , \\u1_u0_token0_reg[2] ,
    \\u0_u0_state_reg[8] , \\u4_u3_csr1_reg[2] , u4_u3_ots_stop_reg,
    \\u4_u0_buf0_orig_reg[7] , \\u4_u1_csr1_reg[3] ,
    \\u4_u0_buf0_orig_reg[8] , \\u4_u2_buf0_orig_reg[27] ,
    \\u4_u2_buf0_orig_reg[28] , \\u1_u0_pid_reg[6] , \\u4_dout_reg[22] ,
    \\u4_dout_reg[23] , \\u4_dout_reg[7] , \\u4_u2_buf0_orig_reg[14] ,
    \\u4_u1_buf0_orig_reg[13] , \\u4_u2_buf0_orig_reg[1] ,
    \\u4_u1_buf0_orig_reg[0] , \\u4_u2_buf0_orig_reg[23] ,
    \\u4_u0_buf0_orig_reg[4] , \\u4_funct_adr_reg[5] ,
    \\u4_funct_adr_reg[3] , \\u4_u3_csr1_reg[6] ,
    \\u4_u2_buf0_orig_reg[16] , \\u4_dout_reg[8] ,
    \\u4_u0_buf0_orig_reg[6] , \\u4_u3_csr1_reg[10] ,
    \\u4_u0_buf0_orig_reg[31] , \\u4_u1_csr0_reg[8] ,
    \\u4_u0_buf0_orig_reg[20] , \\u4_u1_csr1_reg[1] , \\u1_u0_pid_reg[7] ,
    \\u4_u1_csr1_reg[11] , \\u4_u3_csr0_reg[7] ,
    \\u4_u0_buf0_orig_reg[28] , \\u4_u1_csr0_reg[6] ,
    \\u4_u1_csr0_reg[12] , \\u4_u2_buf0_orig_reg[10] ,
    \\u4_u2_buf0_orig_reg[12] , \\u4_u0_buf0_orig_reg[22] ,
    \\u1_u2_state_reg[6] , \\u4_u0_buf0_orig_reg[26] ,
    \\u1_u2_state_reg[1] , \\u1_u2_state_reg[5] , \\u4_u1_csr0_reg[1] ,
    \\u4_u0_buf0_orig_reg[24] , \\u4_funct_adr_reg[0] ,
    \\u4_funct_adr_reg[1] , \\u4_funct_adr_reg[2] , \\u4_funct_adr_reg[4] ,
    \\u4_funct_adr_reg[6] , u1_u3_out_to_small_r_reg, u4_u2_ots_stop_reg,
    u1_u2_mack_r_reg, \\u4_u3_csr0_reg[10] , \\u4_u3_csr0_reg[12] ,
    \\u4_u3_csr0_reg[1] , \\u4_u3_csr0_reg[2] , \\u4_u3_csr0_reg[4] ,
    \\u4_u3_csr0_reg[5] , \\u4_u3_csr0_reg[6] , \\u4_u3_csr0_reg[8] ,
    \\u4_u3_csr0_reg[9] , \\u4_u3_csr1_reg[0] , \\u4_u3_csr1_reg[11] ,
    \\u4_u3_csr1_reg[12] , \\u4_u3_csr1_reg[1] , \\u4_u3_csr1_reg[3] ,
    \\u4_u3_csr1_reg[4] , \\u4_u3_csr1_reg[5] , \\u4_u3_csr1_reg[9] ,
    \\u4_u0_csr0_reg[10] , \\u4_u0_csr0_reg[12] , \\u4_u0_csr0_reg[6] ,
    \\u4_u0_csr1_reg[0] , \\u4_u0_csr1_reg[5] , \\u4_u0_csr1_reg[9] ,
    u4_u0_ots_stop_reg, \\u4_u1_csr0_reg[0] , \\u4_u1_csr0_reg[10] ,
    \\u4_u1_csr0_reg[11] , \\u4_u1_csr0_reg[4] , \\u4_u1_csr0_reg[7] ,
    \\u4_u1_csr1_reg[0] , \\u4_u1_csr1_reg[12] , \\u4_u1_csr1_reg[2] ,
    \\u4_u1_csr1_reg[4] , \\u4_u1_csr1_reg[5] , \\u4_u1_csr1_reg[6] ,
    \\u4_u1_csr1_reg[9] , u4_u1_ots_stop_reg, \\u4_u2_csr0_reg[10] ,
    \\u4_u2_csr0_reg[12] , \\u4_u2_csr0_reg[4] , \\u4_u2_csr0_reg[7] ,
    \\u4_u2_csr1_reg[0] , \\u4_u2_csr1_reg[11] , \\u4_u2_csr1_reg[1] ,
    \\u4_u2_csr1_reg[3] , \\u4_u2_csr1_reg[6] , \\u4_u2_csr1_reg[5] ,
    \\u4_u3_buf0_orig_reg[0] , \\u4_u3_buf0_orig_reg[12] ,
    \\u4_u3_buf0_orig_reg[14] , \\u4_u3_buf0_orig_reg[15] ,
    \\u4_u3_buf0_orig_reg[16] , \\u4_u3_buf0_orig_reg[21] ,
    \\u4_u3_buf0_orig_reg[22] , \\u4_u3_buf0_orig_reg[23] ,
    \\u4_u3_buf0_orig_reg[24] , \\u4_u3_buf0_orig_reg[26] ,
    \\u4_u3_buf0_orig_reg[28] , \\u4_u3_buf0_orig_reg[30] ,
    \\u4_u3_buf0_orig_reg[31] , \\u4_u3_buf0_orig_reg[5] ,
    \\u4_u3_buf0_orig_reg[8] , \\u4_u3_csr1_reg[8] ,
    \\u4_u3_int_stat_reg[1] , \\u4_u0_buf0_orig_reg[10] ,
    \\u4_u0_buf0_orig_reg[11] , \\u4_u0_buf0_orig_reg[12] ,
    \\u4_u0_buf0_orig_reg[14] , \\u4_u0_buf0_orig_reg[16] ,
    \\u4_u0_buf0_orig_reg[18] , \\u4_u0_buf0_orig_reg[1] ,
    \\u4_u0_buf0_orig_reg[21] , \\u4_u0_buf0_orig_reg[23] ,
    \\u4_u0_buf0_orig_reg[25] , \\u4_u0_buf0_orig_reg[27] ,
    \\u4_u0_buf0_orig_reg[29] , \\u4_u0_buf0_orig_reg[2] ,
    \\u4_u0_buf0_orig_reg[30] , \\u4_u0_buf0_orig_reg[3] ,
    \\u4_u0_buf0_orig_reg[5] , \\u4_u0_buf0_orig_reg[9] ,
    \\u4_u3_buf0_orig_reg[9] , \\u4_u0_csr1_reg[8] ,
    \\u4_u1_buf0_orig_reg[10] , \\u4_u1_buf0_orig_reg[11] ,
    \\u4_u1_buf0_orig_reg[12] , \\u4_u1_buf0_orig_reg[14] ,
    \\u4_u1_buf0_orig_reg[15] , \\u4_u1_buf0_orig_reg[16] ,
    \\u4_u1_buf0_orig_reg[18] , \\u4_u1_buf0_orig_reg[19] ,
    \\u4_u1_buf0_orig_reg[1] , \\u4_u1_buf0_orig_reg[21] ,
    \\u4_u1_buf0_orig_reg[22] , \\u4_u1_buf0_orig_reg[23] ,
    \\u4_u1_buf0_orig_reg[25] , \\u4_u1_buf0_orig_reg[26] ,
    \\u4_u1_buf0_orig_reg[27] , \\u4_u1_buf0_orig_reg[2] ,
    \\u4_u1_buf0_orig_reg[29] , \\u4_u1_buf0_orig_reg[3] ,
    \\u4_u1_buf0_orig_reg[4] , \\u4_u1_buf0_orig_reg[5] ,
    \\u4_u1_buf0_orig_reg[7] , \\u4_u1_csr1_reg[8] ,
    \\u4_u2_buf0_orig_reg[0] , \\u4_u2_buf0_orig_reg[11] ,
    \\u4_u2_buf0_orig_reg[13] , \\u4_u2_buf0_orig_reg[15] ,
    \\u4_u2_buf0_orig_reg[17] , \\u4_u2_buf0_orig_reg[18] ,
    \\u4_u2_buf0_orig_reg[19] , \\u4_u2_buf0_orig_reg[20] ,
    \\u4_u2_buf0_orig_reg[21] , \\u4_u2_buf0_orig_reg[22] ,
    \\u4_u2_buf0_orig_reg[24] , \\u4_u2_buf0_orig_reg[25] ,
    \\u4_u2_buf0_orig_reg[26] , \\u4_u2_buf0_orig_reg[2] ,
    \\u4_u2_buf0_orig_reg[31] , \\u4_u2_buf0_orig_reg[4] ,
    \\u4_u2_buf0_orig_reg[7] , \\u4_u2_buf0_orig_reg[9] ,
    \\u4_u2_csr1_reg[8] , \\u5_wb_data_o_reg[14] , \\u1_u0_pid_reg[0] ,
    \\u1_u0_pid_reg[1] , \\u1_u0_pid_reg[2] , \\u1_u0_pid_reg[4] ,
    \\u1_u0_pid_reg[5] , \\u4_u2_buf0_orig_reg[29] ,
    u1_u0_token_valid_str1_reg, u4_match_r1_reg, \\u4_u0_csr0_reg[0] ,
    \\u1_u0_pid_reg[3] , \\u4_u3_csr0_reg[0] , \\u4_u1_buf0_orig_reg[31] ,
    \\u4_u0_buf0_orig_reg[13] , \\u4_u1_buf0_orig_reg[9] ,
    \\u4_u0_buf0_orig_reg[19] , \\u4_u2_csr1_reg[9] ,
    \\u4_u3_csr0_reg[11] , \\u4_u1_buf0_orig_reg[6] ,
    \\u4_u1_buf0_orig_reg[8] , \\u4_u0_buf0_orig_reg[15] ,
    \\u4_u0_buf0_orig_reg[17] , \\u4_u1_buf0_orig_reg[17] ,
    \\u4_u1_buf0_orig_reg[28] , u1_u2_wr_done_reg, u1_u2_idma_done_reg,
    \\u4_u0_csr1_reg[10] , \\u4_u2_csr1_reg[4] , \\u4_u0_buf0_orig_reg[0] ,
    \\u4_u2_csr1_reg[2] , \\u4_u0_csr1_reg[11] , \\u4_u0_csr1_reg[12] ,
    \\u4_u2_csr0_reg[5] , \\u4_u2_csr1_reg[12] , \\u4_u0_csr1_reg[4] ,
    \\u4_u2_csr1_reg[10] , \\u4_u0_csr1_reg[6] , \\u4_u3_buf0_orig_reg[3] ,
    \\u4_u1_buf0_orig_reg[24] , \\u4_u2_csr0_reg[8] ,
    \\u4_u2_buf0_orig_reg[30] , \\u4_u0_csr0_reg[9] ,
    \\u4_u0_csr0_reg[11] , \\u4_u3_buf0_orig_reg[29] ,
    \\u4_u0_csr0_reg[8] , \\u4_u2_csr0_reg[1] , \\u4_u0_csr0_reg[5] ,
    \\u4_u2_csr0_reg[11] , \\u4_u0_csr0_reg[7] ,
    \\u4_u3_buf0_orig_reg[25] , \\u4_u1_buf0_orig_reg[20] ,
    \\u4_u0_csr0_reg[3] , \\u4_u2_buf0_orig_reg[6] ,
    \\u4_u2_buf0_orig_reg[8] , \\u4_u0_csr0_reg[1] ,
    \\u4_u2_buf0_orig_reg[5] , \\u4_u2_buf0_orig_reg[3] ,
    \\u4_u3_buf0_orig_reg[20] , \\u4_u3_buf0_orig_reg[18] ,
    \\u1_u0_token1_reg[6] , \\u4_dout_reg[4] , \\u4_inta_msk_reg[8] ,
    \\u4_intb_msk_reg[3] , \\u4_inta_msk_reg[2] , \\u4_inta_msk_reg[4] ,
    \\u4_inta_msk_reg[0] , \\u4_u3_buf0_orig_reg[1] , \\u4_dout_reg[20] ,
    \\u4_dout_reg[16] , \\u4_dout_reg[17] , \\u4_dout_reg[18] ,
    \\u4_dout_reg[19] , \\u4_dout_reg[21] , \\u4_dout_reg[24] ,
    \\u4_dout_reg[25] , \\u4_dout_reg[26] , \\u4_dout_reg[28] ,
    \\u4_dout_reg[5] , \\u4_dout_reg[6] , \\u4_u3_buf0_orig_reg[17] ,
    \\u4_u3_dma_out_left_reg[8] , \\u4_u0_dma_out_left_reg[8] ,
    \\u4_u1_dma_out_left_reg[8] , \\u4_u2_dma_out_left_reg[8] ,
    \\u4_u1_csr0_reg[3] , \\u4_u3_buf0_orig_reg[11] ,
    \\u4_u3_buf0_orig_reg[13] , \\u1_u0_token1_reg[0] ,
    \\u4_u3_int_stat_reg[6] , suspend_clr_wr_reg,
    \\u4_u3_buf0_orig_reg[10] , \\u1_u0_token1_reg[1] ,
    \\u1_u0_token1_reg[2] , \\u4_inta_msk_reg[1] , \\u4_inta_msk_reg[3] ,
    \\u4_inta_msk_reg[5] , \\u4_inta_msk_reg[6] , \\u4_inta_msk_reg[7] ,
    \\u4_intb_msk_reg[0] , \\u4_intb_msk_reg[1] , \\u4_intb_msk_reg[2] ,
    \\u4_intb_msk_reg[4] , \\u4_intb_msk_reg[5] , \\u4_intb_msk_reg[6] ,
    \\u4_intb_msk_reg[8] , \\u4_u3_buf0_orig_reg[19] ,
    \\u4_u3_buf0_orig_reg[4] , \\u4_u3_buf0_orig_reg[7] ,
    \\u1_u0_token1_reg[3] , \\u1_u0_token1_reg[4] , \\u1_u0_token1_reg[5] ,
    \\u1_u0_token1_reg[7] , \\u4_u3_csr0_reg[3] , \\u4_intb_msk_reg[7] ,
    \\u4_u0_dma_out_left_reg[11] , \\u4_u1_dma_out_left_reg[11] ,
    \\u4_u2_csr0_reg[3] , \\u4_u3_buf0_orig_reg[6] ,
    \\u4_u3_buf0_orig_reg[2] , u0_u0_idle_long_reg,
    \\u4_u3_buf0_orig_reg[27] , \\u4_u3_ienb_reg[5] , \\u4_u3_iena_reg[3] ,
    \\u4_u1_iena_reg[4] , \\u4_u3_ienb_reg[2] , \\u4_u3_ienb_reg[4] ,
    \\u4_u1_iena_reg[5] , \\u4_u3_iena_reg[4] , \\u4_u3_ienb_reg[3] ,
    \\u4_u3_ienb_reg[1] , \\u4_u3_iena_reg[5] , \\u4_u3_ienb_reg[0] ,
    \\u1_u3_new_size_reg[0] , \\u4_u1_iena_reg[0] , \\u4_u0_csr1_reg[7] ,
    \\u4_u3_csr1_reg[7] , \\u4_u1_iena_reg[1] , \\u4_u3_iena_reg[1] ,
    \\u4_u1_iena_reg[3] , \\u4_dout_reg[29] , \\u4_dout_reg[30] ,
    \\u4_dout_reg[31] , \\u4_dout_reg[27] , \\u4_u1_csr1_reg[7] ,
    \\u1_u2_state_reg[7] , \\u4_dout_reg[10] , \\u4_dout_reg[11] ,
    \\u4_dout_reg[9] , \\u4_u2_iena_reg[1] , \\u4_u2_iena_reg[3] ,
    \\u4_u2_iena_reg[5] , \\u4_u2_ienb_reg[0] , \\u4_u2_ienb_reg[1] ,
    \\u4_u2_ienb_reg[4] , \\u4_u2_ienb_reg[3] , \\u4_u3_iena_reg[0] ,
    \\u4_u3_iena_reg[2] , \\u4_u0_iena_reg[1] , \\u4_u0_iena_reg[2] ,
    \\u4_u0_iena_reg[3] , \\u4_u0_iena_reg[5] , \\u4_u0_ienb_reg[1] ,
    \\u4_u0_ienb_reg[4] , \\u4_u0_ienb_reg[3] , \\u4_u1_iena_reg[2] ,
    \\u4_u1_ienb_reg[4] , \\u4_dout_reg[12] , \\u4_u0_ienb_reg[5] ,
    \\u4_u1_ienb_reg[0] , \\u4_u0_ienb_reg[2] , \\u4_u0_iena_reg[4] ,
    \\u4_u0_ienb_reg[0] , \\u4_u3_dma_out_left_reg[11] ,
    \\u4_u2_dma_out_left_reg[11] , \\u4_u2_iena_reg[0] ,
    \\u5_state_reg[3] , \\u4_u1_ienb_reg[1] , \\u4_u2_ienb_reg[5] ,
    \\u4_u0_iena_reg[0] , \\u4_u2_ienb_reg[2] , \\u4_u2_iena_reg[2] ,
    \\u4_u2_iena_reg[4] , \\u4_u1_ienb_reg[2] , u1_u2_rx_data_done_r2_reg,
    u1_u2_wr_done_r_reg, \\u4_u1_ienb_reg[3] , \\u4_u1_ienb_reg[5] ,
    \\u4_u2_csr1_reg[7] , \\u4_dout_reg[13] , \\u4_dout_reg[15] ,
    u1_u3_tx_data_to_reg, u1_u3_rx_ack_to_reg, u1_u2_rx_data_done_r_reg,
    \\u4_utmi_vend_ctrl_r_reg[2] , \\u4_u1_dma_out_left_reg[7] ,
    \\u4_u1_buf0_orig_m3_reg[11] , \\u1_u1_state_reg[2] ,
    \\u4_utmi_vend_ctrl_r_reg[1] , u4_int_src_re_reg,
    \\u4_utmi_vend_ctrl_r_reg[0] , \\u4_utmi_vend_ctrl_r_reg[3] ,
    u1_u0_token_valid_r1_reg, u4_utmi_vend_wr_r_reg, \\u1_u1_state_reg[3] ,
    u4_u0_ep_match_r_reg, \\u4_u3_dma_out_left_reg[7] ,
    \\u4_u0_dma_out_left_reg[7] , \\u4_u2_dma_out_left_reg[7] ,
    \\u4_u0_buf0_orig_m3_reg[11] , \\u4_u0_buf0_orig_m3_reg[9] ,
    \\u4_u2_buf0_orig_m3_reg[9] , u4_u1_int_re_reg,
    \\u4_u0_buf0_orig_m3_reg[10] , u4_u2_int_re_reg, u4_u0_int_re_reg,
    \\u4_u2_buf0_orig_m3_reg[10] , \\u4_u3_dma_out_left_reg[6] ,
    \\u4_u0_dma_out_left_reg[6] , \\u4_u1_dma_out_left_reg[6] ,
    \\u4_dout_reg[14] , \\u4_u2_dma_out_left_reg[6] , u4_u1_ep_match_r_reg,
    \\u4_u3_buf0_orig_m3_reg[11] , \\u4_u2_buf0_orig_m3_reg[11] ,
    \\u4_u0_dma_out_left_reg[5] , \\u4_u3_dma_out_left_reg[5] ,
    \\u4_u1_dma_out_left_reg[5] , \\u4_u2_dma_out_left_reg[5] ,
    \\u4_u1_buf0_orig_m3_reg[7] , \\u4_u1_buf0_orig_m3_reg[8] ,
    \\u4_u1_buf0_orig_m3_reg[10] , u0_u0_usb_attached_reg,
    u1_u3_in_token_reg, u4_u2_ep_match_r_reg,
    \\u1_u3_tx_data_to_cnt_reg[4] , \\u4_u0_buf0_orig_m3_reg[7] ,
    \\u4_u0_buf0_orig_m3_reg[8] , \\u1_u3_tx_data_to_cnt_reg[6] ,
    \\u1_u3_tx_data_to_cnt_reg[2] , \\u1_u3_tx_data_to_cnt_reg[1] ,
    \\u1_u3_tx_data_to_cnt_reg[0] , \\u4_u3_buf0_orig_m3_reg[9] ,
    \\u4_u1_buf0_orig_m3_reg[9] , \\u4_u3_buf0_orig_m3_reg[10] ,
    u1_u3_buf0_na_reg, u1_u3_buf1_na_reg, \\u1_u3_tx_data_to_cnt_reg[3] ,
    u4_u3_int_re_reg, \\u4_u0_buf0_orig_m3_reg[6] ,
    \\u4_u2_buf0_orig_m3_reg[6] , \\u1_u3_tx_data_to_cnt_reg[7] ,
    u4_u0_dma_req_in_hold_reg, \\u1_u3_tx_data_to_cnt_reg[5] ,
    u0_u0_mode_hs_reg, u4_u3_ep_match_r_reg, \\u1_u3_idin_reg[22] ,
    \\u4_u1_buf0_orig_m3_reg[3] , \\u4_u3_buf0_orig_m3_reg[7] ,
    \\u4_u2_buf0_orig_m3_reg[7] , \\u4_u3_buf0_orig_m3_reg[8] ,
    \\u4_u2_buf0_orig_m3_reg[8] , \\u4_int_srca_reg[1] ,
    \\u4_u1_buf0_orig_m3_reg[4] , \\u4_u1_buf0_orig_m3_reg[2] ,
    \\u4_u1_buf0_orig_m3_reg[6] , u4_u2_dma_req_in_hold_reg,
    u4_u1_dma_req_in_hold_reg, u1_u3_out_token_reg, u1_u3_setup_token_reg,
    u0_u0_ls_idle_r_reg, u1_u0_rx_active_r_reg,
    \\u4_u0_buf0_orig_m3_reg[3] , \\u4_u3_dma_out_left_reg[4] ,
    \\u4_u0_dma_out_left_reg[4] , \\u4_u1_dma_out_left_reg[4] ,
    \\u4_u2_dma_out_left_reg[4] , \\u1_u3_rx_ack_to_cnt_reg[4] ,
    \\u4_int_srca_reg[0] , \\u4_int_srca_reg[3] , \\u4_int_srca_reg[2] ,
    \\u1_u3_rx_ack_to_cnt_reg[3] , \\u4_u0_buf0_orig_m3_reg[4] ,
    \\u1_u3_rx_ack_to_cnt_reg[2] , \\u4_u0_buf0_orig_m3_reg[2] ,
    u1_u3_buf1_not_aloc_reg, u1_u3_buf0_not_aloc_reg,
    \\u4_u0_buf0_orig_m3_reg[5] , \\u4_u1_buf0_orig_m3_reg[5] ,
    \\u4_u3_buf0_orig_m3_reg[6] , \\u4_u2_buf0_orig_m3_reg[5] ,
    \\u1_u3_rx_ack_to_cnt_reg[6] , \\u1_u3_rx_ack_to_cnt_reg[0] ,
    \\u1_u3_rx_ack_to_cnt_reg[1] , \\u1_u3_rx_ack_to_cnt_reg[7] ,
    u4_u3_dma_req_in_hold_reg, \\u1_u3_rx_ack_to_cnt_reg[5] ,
    \\u0_u0_idle_cnt1_next_reg[7] , u4_pid_cs_err_r_reg,
    \\u4_u3_buf0_orig_m3_reg[3] , \\u4_u2_buf0_orig_m3_reg[3] ,
    u1_u3_buf0_rl_reg, \\u0_u0_idle_cnt1_next_reg[6] ,
    \\u4_u3_dma_out_left_reg[3] , \\u4_u0_dma_out_left_reg[3] ,
    \\u4_u1_dma_out_left_reg[3] , \\u4_u2_dma_out_left_reg[3] ,
    \\u0_u0_idle_cnt1_next_reg[4] , \\u4_u3_buf0_orig_m3_reg[4] ,
    u0_u0_me_ps2_0_5_ms_reg, \\u4_u2_buf0_orig_m3_reg[4] ,
    \\u4_u2_buf0_orig_m3_reg[2] , \\u4_u3_buf0_orig_m3_reg[5] ,
    u4_u2_dma_req_out_hold_reg, u4_u3_dma_req_out_hold_reg,
    u4_u0_dma_req_out_hold_reg, u4_u1_dma_req_out_hold_reg,
    u1_u1_send_data_r2_reg, u4_usb_reset_r_reg, u0_u0_idle_cnt1_clr_reg,
    \\u4_u3_buf0_orig_m3_reg[2] , \\u0_u0_idle_cnt1_next_reg[5] ,
    u1_u2_sizd_is_zero_reg, u4_rx_err_r_reg, u0_drive_k_r_reg,
    \\u0_u0_idle_cnt1_next_reg[3] , u4_u2_dma_ack_wr1_reg,
    \\u4_u1_dma_out_left_reg[2] , \\u4_u0_dma_out_left_reg[2] ,
    \\u4_u3_dma_out_left_reg[2] , \\u4_u2_dma_out_left_reg[2] ,
    u4_u1_dma_ack_wr1_reg, \\u4_u2_dma_out_left_reg[1] ,
    \\u4_u1_dma_out_left_reg[1] , \\u4_u0_dma_out_left_reg[1] ,
    \\u4_u3_dma_out_left_reg[1] , u4_u0_dma_ack_wr1_reg,
    u4_u3_dma_ack_wr1_reg, \\u1_u2_rd_buf1_reg[19] ,
    \\u1_u2_rd_buf1_reg[1] , \\u4_u0_buf0_orig_m3_reg[1] ,
    \\u4_u3_buf0_orig_m3_reg[1] , \\u4_u2_buf0_orig_m3_reg[1] ,
    u1_u3_pid_OUT_r_reg, u4_u2_set_r_reg, u1_u3_pid_IN_r_reg,
    u4_u0_set_r_reg, u4_u1_set_r_reg, \\u1_u2_rd_buf1_reg[31] ,
    \\u1_u2_rd_buf1_reg[30] , \\u1_u2_rd_buf1_reg[7] ,
    \\u1_u2_rd_buf1_reg[24] , \\u1_u2_rd_buf1_reg[21] ,
    u0_u0_usb_reset_reg, u1_u2_dtmp_sel_r_reg, u1_u3_pid_SETUP_r_reg,
    u1_u3_rx_ack_to_clr_reg, u1_u3_pid_PING_r_reg, u4_u2_r2_reg,
    \\u1_u2_rd_buf1_reg[26] , \\u1_u2_rd_buf1_reg[27] ,
    \\u1_u2_rd_buf1_reg[3] , \\u1_u2_rd_buf1_reg[0] ,
    \\u1_u2_rd_buf1_reg[12] , \\u1_u2_rd_buf1_reg[2] ,
    \\u1_u2_rd_buf1_reg[8] , \\u1_u2_rd_buf1_reg[18] ,
    \\u1_u2_rd_buf1_reg[28] , \\u1_u2_rd_buf1_reg[14] , u4_u3_set_r_reg,
    \\u1_u2_rd_buf1_reg[6] , \\u1_u2_rd_buf1_reg[5] ,
    \\u1_u2_rd_buf1_reg[9] , \\u1_u2_rd_buf1_reg[20] ,
    \\u1_u2_rd_buf1_reg[22] , \\u1_u2_rd_buf1_reg[15] ,
    \\u1_u2_rd_buf1_reg[23] , \\u1_u2_rd_buf1_reg[25] ,
    \\u1_u2_rd_buf1_reg[17] , u4_u3_r2_reg, \\u1_u2_rd_buf1_reg[16] ,
    \\u1_u2_rd_buf1_reg[4] , u4_u0_r2_reg, u4_u1_r2_reg,
    \\u1_u2_rd_buf1_reg[29] , \\u1_u2_rd_buf1_reg[10] , u4_u1_intb_reg,
    u4_u2_intb_reg, u4_u0_intb_reg, \\u1_u2_rd_buf1_reg[11] ,
    \\u1_u2_rd_buf1_reg[13] , u4_u0_inta_reg, u4_u1_inta_reg,
    u4_u2_inta_reg, u4_u3_inta_reg, u4_u3_intb_reg, u0_u0_me_ps_2_5_us_reg,
    \\u4_u3_dma_out_left_reg[0] , \\u4_u2_dma_out_left_reg[0] ,
    \\u4_u0_dma_out_left_reg[0] , u1_u1_send_data_r_reg, u0_rx_active_reg,
    u0_rx_err_reg, u0_rx_valid_reg, u0_u0_ls_se0_r_reg,
    \\u4_u1_dma_out_left_reg[0] , \\u0_u0_idle_cnt1_next_reg[2] ,
    \\u1_u2_rd_buf0_reg[2] , \\u1_u2_rd_buf0_reg[31] ,
    \\u1_u2_rd_buf0_reg[28] , \\u1_u2_rd_buf0_reg[6] ,
    \\u1_u2_rd_buf0_reg[23] , \\u4_u1_buf0_orig_m3_reg[1] ,
    \\u1_u2_rd_buf0_reg[19] , \\u1_u2_rd_buf0_reg[24] ,
    \\u1_u2_rd_buf0_reg[18] , \\u1_u2_rd_buf0_reg[10] ,
    \\u1_u2_rd_buf0_reg[4] , \\u1_u2_rd_buf0_reg[30] ,
    \\u1_u2_rd_buf0_reg[27] , \\u1_u2_rd_buf0_reg[3] ,
    \\u1_u2_rd_buf0_reg[5] , \\u1_u2_rd_buf0_reg[8] ,
    \\u1_u2_rd_buf0_reg[26] , \\u1_u2_rd_buf0_reg[14] ,
    \\u1_u2_rd_buf0_reg[0] , \\u1_u2_rd_buf0_reg[1] ,
    \\u1_u2_rd_buf0_reg[29] , \\u1_u2_rd_buf0_reg[9] ,
    \\u1_u2_rd_buf0_reg[21] , \\u1_u2_rd_buf0_reg[20] ,
    \\u1_u2_rd_buf0_reg[16] , \\u1_u2_rd_buf0_reg[17] ,
    \\u1_u2_rd_buf0_reg[7] , \\u1_u2_rd_buf0_reg[22] ,
    \\u1_u2_rd_buf0_reg[13] , \\u1_u2_rd_buf0_reg[25] ,
    \\u1_u2_rd_buf0_reg[12] , \\u1_u2_rd_buf0_reg[15] ,
    \\u1_u2_rd_buf0_reg[11] , u0_u0_ps_cnt_clr_reg, \\u1_u3_idin_reg[31] ,
    u0_u0_drive_k_reg, u0_u0_ls_j_r_reg, u1_u2_mwe_reg,
    u0_u0_chirp_cnt_is_6_reg, u1_hms_clk_reg, \\u1_u3_idin_reg[28] ,
    \\u0_u0_idle_cnt1_next_reg[1] , u0_u0_ls_k_r_reg, u4_suspend_r1_reg,
    u4_attach_r1_reg, \\u0_u0_state_reg[0] , \\u4_u1_buf0_orig_m3_reg[0] ,
    u4_u1_r5_reg, u4_suspend_r_reg, \\u4_utmi_vend_stat_r_reg[5] ,
    \\u4_utmi_vend_stat_r_reg[2] , u0_u0_resume_req_s_reg,
    \\u4_utmi_vend_stat_r_reg[1] , \\u4_utmi_vend_stat_r_reg[7] ,
    \\u4_utmi_vend_stat_r_reg[4] , \\u4_utmi_vend_stat_r_reg[0] ,
    u5_wb_req_s1_reg, u4_u1_dma_ack_clr1_reg, u4_u0_r5_reg,
    u4_u0_dma_ack_clr1_reg, u0_tx_ready_reg, \\u4_utmi_vend_stat_r_reg[6] ,
    u4_u2_dma_ack_clr1_reg, u1_u3_uc_dpd_set_reg, u4_u3_dma_ack_clr1_reg,
    u4_u2_r5_reg, u1_u3_uc_bsel_set_reg, u4_u3_r5_reg,
    \\u4_utmi_vend_stat_r_reg[3] , susp_o_reg,
    \\u4_u0_buf0_orig_m3_reg[0] , \\u4_u2_buf0_orig_m3_reg[0] ,
    \\u4_u3_buf0_orig_m3_reg[0] , \\u0_u0_idle_cnt1_next_reg[0] ,
    \\u4_utmi_vend_ctrl_reg[3] , u4_utmi_vend_wr_reg,
    \\u4_utmi_vend_ctrl_reg[0] , \\u1_u2_rx_data_st_r_reg[4] ,
    \\u4_utmi_vend_ctrl_reg[2] , \\u1_u2_rx_data_st_r_reg[7] ,
    \\u1_u2_rx_data_st_r_reg[0] , \\u1_u2_rx_data_st_r_reg[2] ,
    \\u1_u2_rx_data_st_r_reg[3] , \\u4_utmi_vend_ctrl_reg[1] ,
    \\u1_u2_rx_data_st_r_reg[1] , \\u1_u2_rx_data_st_r_reg[5] ,
    \\u1_u2_rx_data_st_r_reg[6] , \\VStatus_r_reg[5] , \\VStatus_r_reg[1] ,
    \\VStatus_r_reg[3] , \\u0_rx_data_reg[2] , \\VStatus_r_reg[2] ,
    u0_u0_resume_req_s1_reg, \\u0_rx_data_reg[7] , u4_attach_r_reg,
    \\u0_rx_data_reg[3] , u4_u3_r4_reg, u1_u3_out_to_small_reg,
    u4_u1_r4_reg, \\LineState_r_reg[0] , \\VStatus_r_reg[4] ,
    \\u0_rx_data_reg[0] , u4_u0_r4_reg, \\u0_rx_data_reg[5] ,
    \\VStatus_r_reg[7] , \\u0_u0_line_state_r_reg[1] ,
    \\u0_rx_data_reg[6] , \\u0_u0_line_state_r_reg[0] ,
    \\u0_rx_data_reg[4] , \\u0_rx_data_reg[1] , \\LineState_r_reg[1] ,
    u4_u2_r4_reg, \\VStatus_r_reg[6] , \\VStatus_r_reg[0] ;
  wire \new_[1995]_ , \new_[1996]_ , \new_[2014]_ , \new_[2015]_ ,
    \new_[2018]_ , \new_[2021]_ , \new_[2022]_ , \new_[2023]_ ,
    \new_[2024]_ , \new_[2025]_ , \new_[2027]_ , \new_[2029]_ ,
    \new_[2030]_ , \new_[2031]_ , \new_[2032]_ , \new_[2033]_ ,
    \new_[2034]_ , \new_[2036]_ , \new_[2038]_ , \new_[2039]_ ,
    \new_[2040]_ , \new_[2042]_ , \new_[2043]_ , \new_[2046]_ ,
    \new_[2047]_ , \new_[2048]_ , \new_[2049]_ , \new_[2052]_ ,
    \new_[2053]_ , \new_[2054]_ , \new_[2056]_ , \new_[2062]_ ,
    \new_[2064]_ , \new_[2065]_ , \new_[2066]_ , \new_[2070]_ ,
    \new_[2072]_ , \new_[2073]_ , \new_[2075]_ , \new_[2076]_ ,
    \new_[2079]_ , \new_[2080]_ , \new_[2081]_ , \new_[2082]_ ,
    \new_[2083]_ , \new_[2084]_ , \new_[2085]_ , \new_[2086]_ ,
    \new_[2087]_ , \new_[2088]_ , \new_[2089]_ , \new_[2090]_ ,
    \new_[2091]_ , \new_[2092]_ , \new_[2093]_ , \new_[2094]_ ,
    \new_[2095]_ , \new_[2096]_ , \new_[2097]_ , \new_[2099]_ ,
    \new_[2100]_ , \new_[2101]_ , \new_[2102]_ , \new_[2103]_ ,
    \new_[2106]_ , \new_[2109]_ , \new_[2111]_ , \new_[2112]_ ,
    \new_[2113]_ , \new_[2114]_ , \new_[2117]_ , \new_[2134]_ ,
    \new_[2135]_ , \new_[2136]_ , \new_[2137]_ , \new_[2138]_ ,
    \new_[2139]_ , \new_[2140]_ , \new_[2141]_ , \new_[2142]_ ,
    \new_[2143]_ , \new_[2144]_ , \new_[2145]_ , \new_[2146]_ ,
    \new_[2147]_ , \new_[2148]_ , \new_[2149]_ , \new_[2150]_ ,
    \new_[2151]_ , \new_[2152]_ , \new_[2153]_ , \new_[2154]_ ,
    \new_[2155]_ , \new_[2156]_ , \new_[2157]_ , \new_[2158]_ ,
    \new_[2159]_ , \new_[2160]_ , \new_[2161]_ , \new_[2162]_ ,
    \new_[2164]_ , \new_[2165]_ , \new_[2166]_ , \new_[2168]_ ,
    \new_[2169]_ , \new_[2170]_ , \new_[2171]_ , \new_[2172]_ ,
    \new_[2173]_ , \new_[2174]_ , \new_[2175]_ , \new_[2176]_ ,
    \new_[2177]_ , \new_[2178]_ , \new_[2180]_ , \new_[2181]_ ,
    \new_[2183]_ , \new_[2184]_ , \new_[2185]_ , \new_[2186]_ ,
    \new_[2187]_ , \new_[2188]_ , \new_[2189]_ , \new_[2190]_ ,
    \new_[2191]_ , \new_[2192]_ , \new_[2193]_ , \new_[2194]_ ,
    \new_[2195]_ , \new_[2196]_ , \new_[2197]_ , \new_[2198]_ ,
    \new_[2199]_ , \new_[2200]_ , \new_[2201]_ , \new_[2202]_ ,
    \new_[2203]_ , \new_[2204]_ , \new_[2205]_ , \new_[2206]_ ,
    \new_[2207]_ , \new_[2208]_ , \new_[2209]_ , \new_[2210]_ ,
    \new_[2218]_ , \new_[2220]_ , \new_[2221]_ , \new_[2223]_ ,
    \new_[2224]_ , \new_[2225]_ , \new_[2226]_ , \new_[2227]_ ,
    \new_[2228]_ , \new_[2229]_ , \new_[2230]_ , \new_[2231]_ ,
    \new_[2232]_ , \new_[2233]_ , \new_[2234]_ , \new_[2236]_ ,
    \new_[2237]_ , \new_[2238]_ , \new_[2239]_ , \new_[2240]_ ,
    \new_[2242]_ , \new_[2243]_ , \new_[2244]_ , \new_[2245]_ ,
    \new_[2246]_ , \new_[2247]_ , \new_[2248]_ , \new_[2249]_ ,
    \new_[2250]_ , \new_[2251]_ , \new_[2252]_ , \new_[2254]_ ,
    \new_[2255]_ , \new_[2256]_ , \new_[2257]_ , \new_[2258]_ ,
    \new_[2260]_ , \new_[2261]_ , \new_[2262]_ , \new_[2263]_ ,
    \new_[2264]_ , \new_[2265]_ , \new_[2266]_ , \new_[2267]_ ,
    \new_[2268]_ , \new_[2269]_ , \new_[2270]_ , \new_[2271]_ ,
    \new_[2272]_ , \new_[2273]_ , \new_[2274]_ , \new_[2275]_ ,
    \new_[2276]_ , \new_[2277]_ , \new_[2278]_ , \new_[2279]_ ,
    \new_[2280]_ , \new_[2282]_ , \new_[2283]_ , \new_[2284]_ ,
    \new_[2285]_ , \new_[2287]_ , \new_[2288]_ , \new_[2289]_ ,
    \new_[2290]_ , \new_[2291]_ , \new_[2292]_ , \new_[2293]_ ,
    \new_[2294]_ , \new_[2295]_ , \new_[2296]_ , \new_[2297]_ ,
    \new_[2298]_ , \new_[2299]_ , \new_[2300]_ , \new_[2301]_ ,
    \new_[2302]_ , \new_[2305]_ , \new_[2306]_ , \new_[2307]_ ,
    \new_[2308]_ , \new_[2309]_ , \new_[2310]_ , \new_[2311]_ ,
    \new_[2312]_ , \new_[2313]_ , \new_[2314]_ , \new_[2315]_ ,
    \new_[2316]_ , \new_[2317]_ , \new_[2318]_ , \new_[2320]_ ,
    \new_[2322]_ , \new_[2323]_ , \new_[2324]_ , \new_[2325]_ ,
    \new_[2326]_ , \new_[2327]_ , \new_[2328]_ , \new_[2329]_ ,
    \new_[2330]_ , \new_[2331]_ , \new_[2332]_ , \new_[2333]_ ,
    \new_[2334]_ , \new_[2335]_ , \new_[2336]_ , \new_[2337]_ ,
    \new_[2338]_ , \new_[2339]_ , \new_[2340]_ , \new_[2341]_ ,
    \new_[2342]_ , \new_[2343]_ , \new_[2344]_ , \new_[2345]_ ,
    \new_[2346]_ , \new_[2347]_ , \new_[2348]_ , \new_[2349]_ ,
    \new_[2352]_ , \new_[2353]_ , \new_[2354]_ , \new_[2355]_ ,
    \new_[2357]_ , \new_[2358]_ , \new_[2359]_ , \new_[2360]_ ,
    \new_[2361]_ , \new_[2362]_ , \new_[2363]_ , \new_[2364]_ ,
    \new_[2365]_ , \new_[2366]_ , \new_[2367]_ , \new_[2368]_ ,
    \new_[2369]_ , \new_[2370]_ , \new_[2372]_ , \new_[2373]_ ,
    \new_[2375]_ , \new_[2379]_ , \new_[2380]_ , \new_[2381]_ ,
    \new_[2382]_ , \new_[2383]_ , \new_[2384]_ , \new_[2385]_ ,
    \new_[2386]_ , \new_[2387]_ , \new_[2388]_ , \new_[2389]_ ,
    \new_[2390]_ , \new_[2391]_ , \new_[2392]_ , \new_[2406]_ ,
    \new_[2407]_ , \new_[2408]_ , \new_[2409]_ , \new_[2410]_ ,
    \new_[2411]_ , \new_[2414]_ , \new_[2415]_ , \new_[2416]_ ,
    \new_[2417]_ , \new_[2418]_ , \new_[2419]_ , \new_[2420]_ ,
    \new_[2421]_ , \new_[2422]_ , \new_[2423]_ , \new_[2425]_ ,
    \new_[2426]_ , \new_[2427]_ , \new_[2428]_ , \new_[2430]_ ,
    \new_[2431]_ , \new_[2432]_ , \new_[2433]_ , \new_[2434]_ ,
    \new_[2435]_ , \new_[2436]_ , \new_[2437]_ , \new_[2438]_ ,
    \new_[2439]_ , \new_[2440]_ , \new_[2441]_ , \new_[2442]_ ,
    \new_[2443]_ , \new_[2444]_ , \new_[2446]_ , \new_[2447]_ ,
    \new_[2448]_ , \new_[2449]_ , \new_[2451]_ , \new_[2452]_ ,
    \new_[2453]_ , \new_[2454]_ , \new_[2455]_ , \new_[2456]_ ,
    \new_[2457]_ , \new_[2458]_ , \new_[2459]_ , \new_[2460]_ ,
    \new_[2461]_ , \new_[2462]_ , \new_[2463]_ , \new_[2464]_ ,
    \new_[2466]_ , \new_[2467]_ , \new_[2468]_ , \new_[2469]_ ,
    \new_[2470]_ , \new_[2471]_ , \new_[2472]_ , \new_[2473]_ ,
    \new_[2474]_ , \new_[2475]_ , \new_[2476]_ , \new_[2477]_ ,
    \new_[2478]_ , \new_[2479]_ , \new_[2481]_ , \new_[2482]_ ,
    \new_[2483]_ , \new_[2484]_ , \new_[2485]_ , \new_[2487]_ ,
    \new_[2488]_ , \new_[2489]_ , \new_[2496]_ , \new_[2497]_ ,
    \new_[2498]_ , \new_[2499]_ , \new_[2500]_ , \new_[2501]_ ,
    \new_[2502]_ , \new_[2503]_ , \new_[2504]_ , \new_[2505]_ ,
    \new_[2506]_ , \new_[2507]_ , \new_[2508]_ , \new_[2514]_ ,
    \new_[2515]_ , \new_[2521]_ , \new_[2522]_ , \new_[2523]_ ,
    \new_[2524]_ , \new_[2525]_ , \new_[2526]_ , \new_[2527]_ ,
    \new_[2528]_ , \new_[2530]_ , \new_[2531]_ , \new_[2532]_ ,
    \new_[2539]_ , \new_[2540]_ , \new_[2541]_ , \new_[2542]_ ,
    \new_[2543]_ , \new_[2544]_ , \new_[2545]_ , \new_[2546]_ ,
    \new_[2547]_ , \new_[2548]_ , \new_[2549]_ , \new_[2550]_ ,
    \new_[2551]_ , \new_[2552]_ , \new_[2553]_ , \new_[2554]_ ,
    \new_[2556]_ , \new_[2557]_ , \new_[2558]_ , \new_[2559]_ ,
    \new_[2560]_ , \new_[2561]_ , \new_[2562]_ , \new_[2563]_ ,
    \new_[2564]_ , \new_[2565]_ , \new_[2566]_ , \new_[2567]_ ,
    \new_[2568]_ , \new_[2569]_ , \new_[2570]_ , \new_[2571]_ ,
    \new_[2572]_ , \new_[2573]_ , \new_[2576]_ , \new_[2577]_ ,
    \new_[2578]_ , \new_[2579]_ , \new_[2580]_ , \new_[2581]_ ,
    \new_[2582]_ , \new_[2583]_ , \new_[2585]_ , \new_[2586]_ ,
    \new_[2587]_ , \new_[2588]_ , \new_[2589]_ , \new_[2590]_ ,
    \new_[2591]_ , \new_[2592]_ , \new_[2593]_ , \new_[2594]_ ,
    \new_[2595]_ , \new_[2596]_ , \new_[2600]_ , \new_[2601]_ ,
    \new_[2602]_ , \new_[2603]_ , \new_[2604]_ , \new_[2607]_ ,
    \new_[2610]_ , \new_[2611]_ , \new_[2612]_ , \new_[2613]_ ,
    \new_[2614]_ , \new_[2615]_ , \new_[2616]_ , \new_[2617]_ ,
    \new_[2619]_ , \new_[2620]_ , \new_[2621]_ , \new_[2622]_ ,
    \new_[2623]_ , \new_[2624]_ , \new_[2625]_ , \new_[2627]_ ,
    \new_[2628]_ , \new_[2629]_ , \new_[2630]_ , \new_[2631]_ ,
    \new_[2632]_ , \new_[2633]_ , \new_[2634]_ , \new_[2635]_ ,
    \new_[2636]_ , \new_[2637]_ , \new_[2638]_ , \new_[2639]_ ,
    \new_[2643]_ , \new_[2644]_ , \new_[2645]_ , \new_[2646]_ ,
    \new_[2647]_ , \new_[2648]_ , \new_[2649]_ , \new_[2650]_ ,
    \new_[2651]_ , \new_[2652]_ , \new_[2653]_ , \new_[2654]_ ,
    \new_[2655]_ , \new_[2656]_ , \new_[2657]_ , \new_[2658]_ ,
    \new_[2659]_ , \new_[2660]_ , \new_[2661]_ , \new_[2662]_ ,
    \new_[2663]_ , \new_[2664]_ , \new_[2665]_ , \new_[2666]_ ,
    \new_[2667]_ , \new_[2668]_ , \new_[2669]_ , \new_[2671]_ ,
    \new_[2672]_ , \new_[2673]_ , \new_[2674]_ , \new_[2676]_ ,
    \new_[2677]_ , \new_[2678]_ , \new_[2679]_ , \new_[2680]_ ,
    \new_[2681]_ , \new_[2682]_ , \new_[2683]_ , \new_[2684]_ ,
    \new_[2685]_ , \new_[2686]_ , \new_[2687]_ , \new_[2688]_ ,
    \new_[2689]_ , \new_[2690]_ , \new_[2691]_ , \new_[2692]_ ,
    \new_[2693]_ , \new_[2694]_ , \new_[2695]_ , \new_[2696]_ ,
    \new_[2697]_ , \new_[2698]_ , \new_[2699]_ , \new_[2700]_ ,
    \new_[2701]_ , \new_[2702]_ , \new_[2703]_ , \new_[2704]_ ,
    \new_[2705]_ , \new_[2706]_ , \new_[2707]_ , \new_[2708]_ ,
    \new_[2709]_ , \new_[2710]_ , \new_[2711]_ , \new_[2712]_ ,
    \new_[2713]_ , \new_[2714]_ , \new_[2715]_ , \new_[2716]_ ,
    \new_[2717]_ , \new_[2718]_ , \new_[2719]_ , \new_[2720]_ ,
    \new_[2721]_ , \new_[2722]_ , \new_[2724]_ , \new_[2725]_ ,
    \new_[2726]_ , \new_[2727]_ , \new_[2728]_ , \new_[2729]_ ,
    \new_[2730]_ , \new_[2731]_ , \new_[2732]_ , \new_[2733]_ ,
    \new_[2734]_ , \new_[2735]_ , \new_[2736]_ , \new_[2737]_ ,
    \new_[2738]_ , \new_[2739]_ , \new_[2740]_ , \new_[2741]_ ,
    \new_[2742]_ , \new_[2743]_ , \new_[2744]_ , \new_[2745]_ ,
    \new_[2746]_ , \new_[2747]_ , \new_[2748]_ , \new_[2749]_ ,
    \new_[2752]_ , \new_[2753]_ , \new_[2754]_ , \new_[2755]_ ,
    \new_[2788]_ , \new_[2792]_ , \new_[2793]_ , \new_[2794]_ ,
    \new_[2795]_ , \new_[2797]_ , \new_[2798]_ , \new_[2800]_ ,
    \new_[2801]_ , \new_[2802]_ , \new_[2804]_ , \new_[2805]_ ,
    \new_[2806]_ , \new_[2807]_ , \new_[2808]_ , \new_[2809]_ ,
    \new_[2810]_ , \new_[2811]_ , \new_[2812]_ , \new_[2813]_ ,
    \new_[2814]_ , \new_[2815]_ , \new_[2816]_ , \new_[2817]_ ,
    \new_[2818]_ , \new_[2819]_ , \new_[2820]_ , \new_[2821]_ ,
    \new_[2824]_ , \new_[2825]_ , \new_[2826]_ , \new_[2827]_ ,
    \new_[2828]_ , \new_[2829]_ , \new_[2830]_ , \new_[2831]_ ,
    \new_[2833]_ , \new_[2836]_ , \new_[2837]_ , \new_[2838]_ ,
    \new_[2839]_ , \new_[2840]_ , \new_[2841]_ , \new_[2842]_ ,
    \new_[2843]_ , \new_[2844]_ , \new_[2845]_ , \new_[2846]_ ,
    \new_[2847]_ , \new_[2848]_ , \new_[2852]_ , \new_[2856]_ ,
    \new_[2857]_ , \new_[2858]_ , \new_[2859]_ , \new_[2860]_ ,
    \new_[2861]_ , \new_[2862]_ , \new_[2863]_ , \new_[2864]_ ,
    \new_[2865]_ , \new_[2866]_ , \new_[2867]_ , \new_[2868]_ ,
    \new_[2869]_ , \new_[2870]_ , \new_[2871]_ , \new_[2872]_ ,
    \new_[2873]_ , \new_[2874]_ , \new_[2875]_ , \new_[2876]_ ,
    \new_[2878]_ , \new_[2881]_ , \new_[2882]_ , \new_[2883]_ ,
    \new_[2884]_ , \new_[2886]_ , \new_[2887]_ , \new_[2888]_ ,
    \new_[2889]_ , \new_[2890]_ , \new_[2892]_ , \new_[2893]_ ,
    \new_[2894]_ , \new_[2895]_ , \new_[2896]_ , \new_[2899]_ ,
    \new_[2917]_ , \new_[2918]_ , \new_[2919]_ , \new_[2920]_ ,
    \new_[2921]_ , \new_[2923]_ , \new_[2924]_ , \new_[2925]_ ,
    \new_[2926]_ , \new_[2927]_ , \new_[2928]_ , \new_[2929]_ ,
    \new_[2931]_ , \new_[2932]_ , \new_[2933]_ , \new_[2934]_ ,
    \new_[2935]_ , \new_[2936]_ , \new_[2938]_ , \new_[2939]_ ,
    \new_[2942]_ , \new_[2960]_ , \new_[2961]_ , \new_[2962]_ ,
    \new_[2963]_ , \new_[2971]_ , \new_[2973]_ , \new_[2974]_ ,
    \new_[2975]_ , \new_[2976]_ , \new_[2977]_ , \new_[2978]_ ,
    \new_[2980]_ , \new_[2981]_ , \new_[2982]_ , \new_[2983]_ ,
    \new_[2984]_ , \new_[2985]_ , \new_[2986]_ , \new_[2987]_ ,
    \new_[2988]_ , \new_[2989]_ , \new_[2990]_ , \new_[2991]_ ,
    \new_[2992]_ , \new_[2993]_ , \new_[2994]_ , \new_[2995]_ ,
    \new_[2996]_ , \new_[2998]_ , \new_[2999]_ , \new_[3000]_ ,
    \new_[3001]_ , \new_[3002]_ , \new_[3003]_ , \new_[3005]_ ,
    \new_[3007]_ , \new_[3008]_ , \new_[3009]_ , \new_[3010]_ ,
    \new_[3011]_ , \new_[3012]_ , \new_[3013]_ , \new_[3015]_ ,
    \new_[3016]_ , \new_[3017]_ , \new_[3020]_ , \new_[3021]_ ,
    \new_[3022]_ , \new_[3023]_ , \new_[3024]_ , \new_[3025]_ ,
    \new_[3026]_ , \new_[3027]_ , \new_[3028]_ , \new_[3029]_ ,
    \new_[3030]_ , \new_[3031]_ , \new_[3032]_ , \new_[3033]_ ,
    \new_[3034]_ , \new_[3035]_ , \new_[3036]_ , \new_[3037]_ ,
    \new_[3038]_ , \new_[3039]_ , \new_[3040]_ , \new_[3041]_ ,
    \new_[3042]_ , \new_[3044]_ , \new_[3045]_ , \new_[3046]_ ,
    \new_[3047]_ , \new_[3048]_ , \new_[3049]_ , \new_[3050]_ ,
    \new_[3058]_ , \new_[3059]_ , \new_[3061]_ , \new_[3062]_ ,
    \new_[3063]_ , \new_[3064]_ , \new_[3065]_ , \new_[3066]_ ,
    \new_[3067]_ , \new_[3068]_ , \new_[3070]_ , \new_[3071]_ ,
    \new_[3072]_ , \new_[3077]_ , \new_[3078]_ , \new_[3079]_ ,
    \new_[3080]_ , \new_[3081]_ , \new_[3082]_ , \new_[3083]_ ,
    \new_[3084]_ , \new_[3085]_ , \new_[3086]_ , \new_[3087]_ ,
    \new_[3088]_ , \new_[3089]_ , \new_[3090]_ , \new_[3091]_ ,
    \new_[3092]_ , \new_[3093]_ , \new_[3094]_ , \new_[3095]_ ,
    \new_[3096]_ , \new_[3097]_ , \new_[3098]_ , \new_[3099]_ ,
    \new_[3100]_ , \new_[3101]_ , \new_[3102]_ , \new_[3103]_ ,
    \new_[3104]_ , \new_[3105]_ , \new_[3107]_ , \new_[3108]_ ,
    \new_[3112]_ , \new_[3113]_ , \new_[3120]_ , \new_[3124]_ ,
    \new_[3126]_ , \new_[3129]_ , \new_[3131]_ , \new_[3132]_ ,
    \new_[3133]_ , \new_[3134]_ , \new_[3136]_ , \new_[3137]_ ,
    \new_[3138]_ , \new_[3139]_ , \new_[3140]_ , \new_[3141]_ ,
    \new_[3142]_ , \new_[3143]_ , \new_[3144]_ , \new_[3145]_ ,
    \new_[3146]_ , \new_[3147]_ , \new_[3148]_ , \new_[3149]_ ,
    \new_[3150]_ , \new_[3151]_ , \new_[3152]_ , \new_[3153]_ ,
    \new_[3154]_ , \new_[3155]_ , \new_[3156]_ , \new_[3157]_ ,
    \new_[3158]_ , \new_[3159]_ , \new_[3160]_ , \new_[3161]_ ,
    \new_[3162]_ , \new_[3163]_ , \new_[3164]_ , \new_[3165]_ ,
    \new_[3166]_ , \new_[3167]_ , \new_[3168]_ , \new_[3169]_ ,
    \new_[3170]_ , \new_[3171]_ , \new_[3172]_ , \new_[3173]_ ,
    \new_[3174]_ , \new_[3175]_ , \new_[3176]_ , \new_[3177]_ ,
    \new_[3178]_ , \new_[3179]_ , \new_[3180]_ , \new_[3181]_ ,
    \new_[3182]_ , \new_[3183]_ , \new_[3184]_ , \new_[3185]_ ,
    \new_[3186]_ , \new_[3187]_ , \new_[3188]_ , \new_[3189]_ ,
    \new_[3190]_ , \new_[3191]_ , \new_[3192]_ , \new_[3193]_ ,
    \new_[3194]_ , \new_[3242]_ , \new_[3243]_ , \new_[3244]_ ,
    \new_[3245]_ , \new_[3248]_ , \new_[3253]_ , \new_[3265]_ ,
    \new_[3266]_ , \new_[3267]_ , \new_[3276]_ , \new_[3277]_ ,
    \new_[3278]_ , \new_[3279]_ , \new_[3280]_ , \new_[3281]_ ,
    \new_[3282]_ , \new_[3283]_ , \new_[3285]_ , \new_[3286]_ ,
    \new_[3288]_ , \new_[3289]_ , \new_[3290]_ , \new_[3291]_ ,
    \new_[3292]_ , \new_[3293]_ , \new_[3294]_ , \new_[3295]_ ,
    \new_[3296]_ , \new_[3297]_ , \new_[3298]_ , \new_[3299]_ ,
    \new_[3300]_ , \new_[3301]_ , \new_[3302]_ , \new_[3303]_ ,
    \new_[3304]_ , \new_[3305]_ , \new_[3306]_ , \new_[3307]_ ,
    \new_[3308]_ , \new_[3309]_ , \new_[3310]_ , \new_[3311]_ ,
    \new_[3312]_ , \new_[3313]_ , \new_[3314]_ , \new_[3315]_ ,
    \new_[3316]_ , \new_[3317]_ , \new_[3318]_ , \new_[3319]_ ,
    \new_[3320]_ , \new_[3321]_ , \new_[3322]_ , \new_[3323]_ ,
    \new_[3324]_ , \new_[3325]_ , \new_[3326]_ , \new_[3327]_ ,
    \new_[3328]_ , \new_[3329]_ , \new_[3330]_ , \new_[3331]_ ,
    \new_[3332]_ , \new_[3333]_ , \new_[3334]_ , \new_[3335]_ ,
    \new_[3336]_ , \new_[3337]_ , \new_[3338]_ , \new_[3339]_ ,
    \new_[3340]_ , \new_[3341]_ , \new_[3342]_ , \new_[3343]_ ,
    \new_[3344]_ , \new_[3345]_ , \new_[3346]_ , \new_[3347]_ ,
    \new_[3348]_ , \new_[3349]_ , \new_[3350]_ , \new_[3351]_ ,
    \new_[3352]_ , \new_[3353]_ , \new_[3354]_ , \new_[3355]_ ,
    \new_[3356]_ , \new_[3357]_ , \new_[3358]_ , \new_[3359]_ ,
    \new_[3360]_ , \new_[3361]_ , \new_[3362]_ , \new_[3363]_ ,
    \new_[3364]_ , \new_[3365]_ , \new_[3366]_ , \new_[3367]_ ,
    \new_[3370]_ , \new_[3371]_ , \new_[3372]_ , \new_[3373]_ ,
    \new_[3374]_ , \new_[3375]_ , \new_[3376]_ , \new_[3377]_ ,
    \new_[3378]_ , \new_[3379]_ , \new_[3380]_ , \new_[3381]_ ,
    \new_[3382]_ , \new_[3383]_ , \new_[3384]_ , \new_[3385]_ ,
    \new_[3386]_ , \new_[3387]_ , \new_[3388]_ , \new_[3389]_ ,
    \new_[3390]_ , \new_[3391]_ , \new_[3392]_ , \new_[3393]_ ,
    \new_[3394]_ , \new_[3395]_ , \new_[3396]_ , \new_[3397]_ ,
    \new_[3398]_ , \new_[3399]_ , \new_[3400]_ , \new_[3401]_ ,
    \new_[3402]_ , \new_[3403]_ , \new_[3404]_ , \new_[3405]_ ,
    \new_[3406]_ , \new_[3407]_ , \new_[3408]_ , \new_[3410]_ ,
    \new_[3413]_ , \new_[3414]_ , \new_[3416]_ , \new_[3420]_ ,
    \new_[3421]_ , \new_[3422]_ , \new_[3423]_ , \new_[3424]_ ,
    \new_[3425]_ , \new_[3428]_ , \new_[3429]_ , \new_[3430]_ ,
    \new_[3431]_ , \new_[3432]_ , \new_[3433]_ , \new_[3434]_ ,
    \new_[3435]_ , \new_[3439]_ , \new_[3440]_ , \new_[3442]_ ,
    \new_[3444]_ , \new_[3447]_ , \new_[3448]_ , \new_[3449]_ ,
    \new_[3450]_ , \new_[3451]_ , \new_[3452]_ , \new_[3453]_ ,
    \new_[3454]_ , \new_[3455]_ , \new_[3456]_ , \new_[3457]_ ,
    \new_[3458]_ , \new_[3459]_ , \new_[3460]_ , \new_[3461]_ ,
    \new_[3462]_ , \new_[3463]_ , \new_[3464]_ , \new_[3465]_ ,
    \new_[3466]_ , \new_[3467]_ , \new_[3468]_ , \new_[3469]_ ,
    \new_[3470]_ , \new_[3471]_ , \new_[3472]_ , \new_[3473]_ ,
    \new_[3474]_ , \new_[3475]_ , \new_[3476]_ , \new_[3477]_ ,
    \new_[3478]_ , \new_[3479]_ , \new_[3480]_ , \new_[3481]_ ,
    \new_[3482]_ , \new_[3483]_ , \new_[3484]_ , \new_[3485]_ ,
    \new_[3486]_ , \new_[3487]_ , \new_[3488]_ , \new_[3489]_ ,
    \new_[3490]_ , \new_[3491]_ , \new_[3492]_ , \new_[3493]_ ,
    \new_[3494]_ , \new_[3495]_ , \new_[3496]_ , \new_[3497]_ ,
    \new_[3498]_ , \new_[3499]_ , \new_[3500]_ , \new_[3501]_ ,
    \new_[3502]_ , \new_[3503]_ , \new_[3504]_ , \new_[3505]_ ,
    \new_[3506]_ , \new_[3507]_ , \new_[3508]_ , \new_[3509]_ ,
    \new_[3510]_ , \new_[3511]_ , \new_[3512]_ , \new_[3513]_ ,
    \new_[3514]_ , \new_[3515]_ , \new_[3516]_ , \new_[3517]_ ,
    \new_[3518]_ , \new_[3519]_ , \new_[3520]_ , \new_[3521]_ ,
    \new_[3522]_ , \new_[3523]_ , \new_[3524]_ , \new_[3525]_ ,
    \new_[3526]_ , \new_[3527]_ , \new_[3531]_ , \new_[3545]_ ,
    \new_[3546]_ , \new_[3547]_ , \new_[3548]_ , \new_[3549]_ ,
    \new_[3550]_ , \new_[3551]_ , \new_[3552]_ , \new_[3553]_ ,
    \new_[3554]_ , \new_[3555]_ , \new_[3556]_ , \new_[3563]_ ,
    \new_[3564]_ , \new_[3566]_ , \new_[3571]_ , \new_[3572]_ ,
    \new_[3573]_ , \new_[3574]_ , \new_[3575]_ , \new_[3576]_ ,
    \new_[3577]_ , \new_[3578]_ , \new_[3579]_ , \new_[3580]_ ,
    \new_[3581]_ , \new_[3582]_ , \new_[3583]_ , \new_[3584]_ ,
    \new_[3585]_ , \new_[3586]_ , \new_[3587]_ , \new_[3588]_ ,
    \new_[3589]_ , \new_[3590]_ , \new_[3591]_ , \new_[3592]_ ,
    \new_[3594]_ , \new_[3595]_ , \new_[3596]_ , \new_[3597]_ ,
    \new_[3598]_ , \new_[3599]_ , \new_[3600]_ , \new_[3601]_ ,
    \new_[3602]_ , \new_[3603]_ , \new_[3604]_ , \new_[3605]_ ,
    \new_[3606]_ , \new_[3607]_ , \new_[3608]_ , \new_[3609]_ ,
    \new_[3610]_ , \new_[3611]_ , \new_[3612]_ , \new_[3613]_ ,
    \new_[3614]_ , \new_[3615]_ , \new_[3616]_ , \new_[3617]_ ,
    \new_[3618]_ , \new_[3621]_ , \new_[3622]_ , \new_[3624]_ ,
    \new_[3626]_ , \new_[3628]_ , \new_[3629]_ , \new_[3630]_ ,
    \new_[3631]_ , \new_[3632]_ , \new_[3633]_ , \new_[3634]_ ,
    \new_[3636]_ , \new_[3638]_ , \new_[3639]_ , \new_[3659]_ ,
    \new_[3671]_ , \new_[3672]_ , \new_[3676]_ , \new_[3677]_ ,
    \new_[3679]_ , \new_[3680]_ , \new_[3681]_ , \new_[3682]_ ,
    \new_[3683]_ , \new_[3684]_ , \new_[3686]_ , \new_[3687]_ ,
    \new_[3688]_ , \new_[3689]_ , \new_[3690]_ , \new_[3691]_ ,
    \new_[3692]_ , \new_[3693]_ , \new_[3694]_ , \new_[3695]_ ,
    \new_[3696]_ , \new_[3697]_ , \new_[3698]_ , \new_[3699]_ ,
    \new_[3700]_ , \new_[3701]_ , \new_[3702]_ , \new_[3703]_ ,
    \new_[3704]_ , \new_[3705]_ , \new_[3706]_ , \new_[3707]_ ,
    \new_[3708]_ , \new_[3709]_ , \new_[3710]_ , \new_[3711]_ ,
    \new_[3712]_ , \new_[3713]_ , \new_[3714]_ , \new_[3715]_ ,
    \new_[3716]_ , \new_[3717]_ , \new_[3718]_ , \new_[3719]_ ,
    \new_[3720]_ , \new_[3721]_ , \new_[3722]_ , \new_[3723]_ ,
    \new_[3724]_ , \new_[3725]_ , \new_[3726]_ , \new_[3727]_ ,
    \new_[3728]_ , \new_[3729]_ , \new_[3730]_ , \new_[3731]_ ,
    \new_[3732]_ , \new_[3733]_ , \new_[3734]_ , \new_[3735]_ ,
    \new_[3736]_ , \new_[3737]_ , \new_[3738]_ , \new_[3739]_ ,
    \new_[3740]_ , \new_[3741]_ , \new_[3742]_ , \new_[3743]_ ,
    \new_[3744]_ , \new_[3763]_ , \new_[3764]_ , \new_[3765]_ ,
    \new_[3775]_ , \new_[3776]_ , \new_[3777]_ , \new_[3781]_ ,
    \new_[3782]_ , \new_[3787]_ , \new_[3788]_ , \new_[3790]_ ,
    \new_[3791]_ , \new_[3794]_ , \new_[3797]_ , \new_[3798]_ ,
    \new_[3799]_ , \new_[3800]_ , \new_[3801]_ , \new_[3802]_ ,
    \new_[3803]_ , \new_[3804]_ , \new_[3805]_ , \new_[3806]_ ,
    \new_[3807]_ , \new_[3808]_ , \new_[3815]_ , \new_[3816]_ ,
    \new_[3818]_ , \new_[3822]_ , \new_[3824]_ , \new_[3829]_ ,
    \new_[3830]_ , \new_[3831]_ , \new_[3832]_ , \new_[3859]_ ,
    \new_[3860]_ , \new_[3862]_ , \new_[3864]_ , \new_[3865]_ ,
    \new_[3866]_ , \new_[3867]_ , \new_[3868]_ , \new_[3869]_ ,
    \new_[3870]_ , \new_[3875]_ , \new_[3878]_ , \new_[3879]_ ,
    \new_[3880]_ , \new_[3881]_ , \new_[3882]_ , \new_[3883]_ ,
    \new_[3884]_ , \new_[3886]_ , \new_[3887]_ , \new_[3888]_ ,
    \new_[3889]_ , \new_[3890]_ , \new_[3891]_ , \new_[3892]_ ,
    \new_[3893]_ , \new_[3894]_ , \new_[3895]_ , \new_[3920]_ ,
    \new_[3921]_ , \new_[3924]_ , \new_[3929]_ , \new_[3930]_ ,
    \new_[3932]_ , \new_[3934]_ , \new_[3935]_ , \new_[3936]_ ,
    \new_[3937]_ , \new_[3938]_ , \new_[3940]_ , \new_[3944]_ ,
    \new_[3958]_ , \new_[3959]_ , \new_[3960]_ , \new_[3961]_ ,
    \new_[3962]_ , \new_[3967]_ , \new_[3968]_ , \new_[3970]_ ,
    \new_[3971]_ , \new_[3972]_ , \new_[3974]_ , \new_[3975]_ ,
    \new_[3977]_ , \new_[3978]_ , \new_[3979]_ , \new_[3980]_ ,
    \new_[3981]_ , \new_[3982]_ , \new_[3983]_ , \new_[3984]_ ,
    \new_[3985]_ , \new_[3986]_ , \new_[3987]_ , \new_[3988]_ ,
    \new_[3989]_ , \new_[3990]_ , \new_[3991]_ , \new_[3992]_ ,
    \new_[3993]_ , \new_[3994]_ , \new_[3995]_ , \new_[3996]_ ,
    \new_[3997]_ , \new_[3998]_ , \new_[4000]_ , \new_[4001]_ ,
    \new_[4003]_ , \new_[4006]_ , \new_[4007]_ , \new_[4008]_ ,
    \new_[4011]_ , \new_[4013]_ , \new_[4017]_ , \new_[4020]_ ,
    \new_[4024]_ , \new_[4029]_ , \new_[4030]_ , \new_[4031]_ ,
    \new_[4032]_ , \new_[4033]_ , \new_[4034]_ , \new_[4035]_ ,
    \new_[4057]_ , \new_[4058]_ , \new_[4059]_ , \new_[4060]_ ,
    \new_[4062]_ , \new_[4063]_ , \new_[4069]_ , \new_[4070]_ ,
    \new_[4071]_ , \new_[4072]_ , \new_[4073]_ , \new_[4074]_ ,
    \new_[4075]_ , \new_[4076]_ , \new_[4077]_ , \new_[4078]_ ,
    \new_[4079]_ , \new_[4080]_ , \new_[4081]_ , \new_[4082]_ ,
    \new_[4083]_ , \new_[4085]_ , \new_[4086]_ , \new_[4087]_ ,
    \new_[4088]_ , \new_[4089]_ , \new_[4090]_ , \new_[4091]_ ,
    \new_[4092]_ , \new_[4095]_ , \new_[4096]_ , \new_[4097]_ ,
    \new_[4098]_ , \new_[4124]_ , \new_[4125]_ , \new_[4126]_ ,
    \new_[4127]_ , \new_[4128]_ , \new_[4129]_ , \new_[4130]_ ,
    \new_[4131]_ , \new_[4132]_ , \new_[4133]_ , \new_[4134]_ ,
    \new_[4135]_ , \new_[4136]_ , \new_[4137]_ , \new_[4138]_ ,
    \new_[4139]_ , \new_[4140]_ , \new_[4141]_ , \new_[4142]_ ,
    \new_[4143]_ , \new_[4144]_ , \new_[4145]_ , \new_[4146]_ ,
    \new_[4147]_ , \new_[4148]_ , \new_[4149]_ , \new_[4150]_ ,
    \new_[4151]_ , \new_[4152]_ , \new_[4153]_ , \new_[4154]_ ,
    \new_[4156]_ , \new_[4157]_ , \new_[4159]_ , \new_[4161]_ ,
    \new_[4162]_ , \new_[4163]_ , \new_[4164]_ , \new_[4165]_ ,
    \new_[4166]_ , \new_[4167]_ , \new_[4168]_ , \new_[4170]_ ,
    \new_[4171]_ , \new_[4172]_ , \new_[4173]_ , \new_[4174]_ ,
    \new_[4175]_ , \new_[4176]_ , \new_[4181]_ , \new_[4182]_ ,
    \new_[4184]_ , \new_[4185]_ , \new_[4186]_ , \new_[4187]_ ,
    \new_[4188]_ , \new_[4189]_ , \new_[4190]_ , \new_[4191]_ ,
    \new_[4192]_ , \new_[4197]_ , \new_[4199]_ , \new_[4201]_ ,
    \new_[4202]_ , \new_[4203]_ , \new_[4204]_ , \new_[4205]_ ,
    \new_[4206]_ , \new_[4207]_ , \new_[4208]_ , \new_[4209]_ ,
    \new_[4210]_ , \new_[4211]_ , \new_[4212]_ , \new_[4213]_ ,
    \new_[4214]_ , \new_[4215]_ , \new_[4216]_ , \new_[4217]_ ,
    \new_[4218]_ , \new_[4219]_ , \new_[4220]_ , \new_[4221]_ ,
    \new_[4222]_ , \new_[4224]_ , \new_[4225]_ , \new_[4227]_ ,
    \new_[4228]_ , \new_[4229]_ , \new_[4230]_ , \new_[4231]_ ,
    \new_[4232]_ , \new_[4233]_ , \new_[4236]_ , \new_[4237]_ ,
    \new_[4238]_ , \new_[4242]_ , \new_[4243]_ , \new_[4245]_ ,
    \new_[4246]_ , \new_[4248]_ , \new_[4249]_ , \new_[4251]_ ,
    \new_[4252]_ , \new_[4253]_ , \new_[4254]_ , \new_[4259]_ ,
    \new_[4260]_ , \new_[4261]_ , \new_[4262]_ , \new_[4263]_ ,
    \new_[4264]_ , \new_[4265]_ , \new_[4266]_ , \new_[4267]_ ,
    \new_[4268]_ , \new_[4269]_ , \new_[4270]_ , \new_[4271]_ ,
    \new_[4272]_ , \new_[4273]_ , \new_[4274]_ , \new_[4275]_ ,
    \new_[4276]_ , \new_[4278]_ , \new_[4279]_ , \new_[4280]_ ,
    \new_[4281]_ , \new_[4282]_ , \new_[4283]_ , \new_[4284]_ ,
    \new_[4285]_ , \new_[4286]_ , \new_[4287]_ , \new_[4288]_ ,
    \new_[4289]_ , \new_[4290]_ , \new_[4291]_ , \new_[4292]_ ,
    \new_[4293]_ , \new_[4300]_ , \new_[4301]_ , \new_[4302]_ ,
    \new_[4305]_ , \new_[4306]_ , \new_[4309]_ , \new_[4310]_ ,
    \new_[4311]_ , \new_[4312]_ , \new_[4313]_ , \new_[4314]_ ,
    \new_[4315]_ , \new_[4316]_ , \new_[4317]_ , \new_[4318]_ ,
    \new_[4319]_ , \new_[4320]_ , \new_[4321]_ , \new_[4322]_ ,
    \new_[4323]_ , \new_[4324]_ , \new_[4325]_ , \new_[4326]_ ,
    \new_[4327]_ , \new_[4328]_ , \new_[4329]_ , \new_[4330]_ ,
    \new_[4331]_ , \new_[4332]_ , \new_[4333]_ , \new_[4334]_ ,
    \new_[4335]_ , \new_[4336]_ , \new_[4337]_ , \new_[4338]_ ,
    \new_[4339]_ , \new_[4340]_ , \new_[4341]_ , \new_[4345]_ ,
    \new_[4346]_ , \new_[4347]_ , \new_[4352]_ , \new_[4353]_ ,
    \new_[4354]_ , \new_[4355]_ , \new_[4356]_ , \new_[4357]_ ,
    \new_[4358]_ , \new_[4360]_ , \new_[4361]_ , \new_[4362]_ ,
    \new_[4366]_ , \new_[4369]_ , \new_[4370]_ , \new_[4371]_ ,
    \new_[4372]_ , \new_[4373]_ , \new_[4374]_ , \new_[4375]_ ,
    \new_[4376]_ , \new_[4377]_ , \new_[4378]_ , \new_[4379]_ ,
    \new_[4380]_ , \new_[4381]_ , \new_[4382]_ , \new_[4383]_ ,
    \new_[4384]_ , \new_[4385]_ , \new_[4386]_ , \new_[4387]_ ,
    \new_[4388]_ , \new_[4389]_ , \new_[4390]_ , \new_[4391]_ ,
    \new_[4392]_ , \new_[4393]_ , \new_[4394]_ , \new_[4395]_ ,
    \new_[4396]_ , \new_[4397]_ , \new_[4398]_ , \new_[4399]_ ,
    \new_[4400]_ , \new_[4401]_ , \new_[4402]_ , \new_[4403]_ ,
    \new_[4404]_ , \new_[4405]_ , \new_[4406]_ , \new_[4407]_ ,
    \new_[4408]_ , \new_[4409]_ , \new_[4410]_ , \new_[4411]_ ,
    \new_[4412]_ , \new_[4413]_ , \new_[4414]_ , \new_[4415]_ ,
    \new_[4418]_ , \new_[4420]_ , \new_[4421]_ , \new_[4422]_ ,
    \new_[4423]_ , \new_[4424]_ , \new_[4425]_ , \new_[4428]_ ,
    \new_[4451]_ , \new_[4453]_ , \new_[4454]_ , \new_[4455]_ ,
    \new_[4456]_ , \new_[4457]_ , \new_[4458]_ , \new_[4459]_ ,
    \new_[4460]_ , \new_[4463]_ , \new_[4464]_ , \new_[4465]_ ,
    \new_[4466]_ , \new_[4467]_ , \new_[4468]_ , \new_[4469]_ ,
    \new_[4470]_ , \new_[4471]_ , \new_[4472]_ , \new_[4473]_ ,
    \new_[4474]_ , \new_[4475]_ , \new_[4476]_ , \new_[4477]_ ,
    \new_[4478]_ , \new_[4479]_ , \new_[4480]_ , \new_[4481]_ ,
    \new_[4482]_ , \new_[4483]_ , \new_[4484]_ , \new_[4485]_ ,
    \new_[4486]_ , \new_[4487]_ , \new_[4489]_ , \new_[4490]_ ,
    \new_[4491]_ , \new_[4492]_ , \new_[4494]_ , \new_[4499]_ ,
    \new_[4500]_ , \new_[4501]_ , \new_[4502]_ , \new_[4503]_ ,
    \new_[4504]_ , \new_[4505]_ , \new_[4506]_ , \new_[4507]_ ,
    \new_[4508]_ , \new_[4509]_ , \new_[4510]_ , \new_[4511]_ ,
    \new_[4512]_ , \new_[4513]_ , \new_[4514]_ , \new_[4515]_ ,
    \new_[4516]_ , \new_[4517]_ , \new_[4518]_ , \new_[4519]_ ,
    \new_[4520]_ , \new_[4521]_ , \new_[4522]_ , \new_[4523]_ ,
    \new_[4524]_ , \new_[4525]_ , \new_[4526]_ , \new_[4527]_ ,
    \new_[4528]_ , \new_[4529]_ , \new_[4530]_ , \new_[4531]_ ,
    \new_[4532]_ , \new_[4533]_ , \new_[4534]_ , \new_[4535]_ ,
    \new_[4536]_ , \new_[4537]_ , \new_[4538]_ , \new_[4539]_ ,
    \new_[4540]_ , \new_[4541]_ , \new_[4542]_ , \new_[4543]_ ,
    \new_[4544]_ , \new_[4545]_ , \new_[4546]_ , \new_[4547]_ ,
    \new_[4548]_ , \new_[4549]_ , \new_[4550]_ , \new_[4551]_ ,
    \new_[4552]_ , \new_[4553]_ , \new_[4554]_ , \new_[4555]_ ,
    \new_[4556]_ , \new_[4557]_ , \new_[4558]_ , \new_[4559]_ ,
    \new_[4560]_ , \new_[4561]_ , \new_[4562]_ , \new_[4563]_ ,
    \new_[4564]_ , \new_[4565]_ , \new_[4566]_ , \new_[4567]_ ,
    \new_[4568]_ , \new_[4569]_ , \new_[4570]_ , \new_[4571]_ ,
    \new_[4572]_ , \new_[4573]_ , \new_[4574]_ , \new_[4575]_ ,
    \new_[4576]_ , \new_[4577]_ , \new_[4578]_ , \new_[4579]_ ,
    \new_[4580]_ , \new_[4581]_ , \new_[4582]_ , \new_[4583]_ ,
    \new_[4584]_ , \new_[4585]_ , \new_[4586]_ , \new_[4587]_ ,
    \new_[4588]_ , \new_[4589]_ , \new_[4590]_ , \new_[4591]_ ,
    \new_[4592]_ , \new_[4594]_ , \new_[4595]_ , \new_[4596]_ ,
    \new_[4597]_ , \new_[4598]_ , \new_[4599]_ , \new_[4600]_ ,
    \new_[4601]_ , \new_[4602]_ , \new_[4603]_ , \new_[4604]_ ,
    \new_[4606]_ , \new_[4607]_ , \new_[4608]_ , \new_[4609]_ ,
    \new_[4610]_ , \new_[4611]_ , \new_[4612]_ , \new_[4613]_ ,
    \new_[4614]_ , \new_[4615]_ , \new_[4616]_ , \new_[4617]_ ,
    \new_[4618]_ , \new_[4619]_ , \new_[4620]_ , \new_[4621]_ ,
    \new_[4624]_ , \new_[4625]_ , \new_[4626]_ , \new_[4627]_ ,
    \new_[4628]_ , \new_[4629]_ , \new_[4630]_ , \new_[4631]_ ,
    \new_[4632]_ , \new_[4633]_ , \new_[4634]_ , \new_[4635]_ ,
    \new_[4636]_ , \new_[4637]_ , \new_[4638]_ , \new_[4639]_ ,
    \new_[4640]_ , \new_[4641]_ , \new_[4642]_ , \new_[4643]_ ,
    \new_[4644]_ , \new_[4645]_ , \new_[4646]_ , \new_[4647]_ ,
    \new_[4648]_ , \new_[4649]_ , \new_[4650]_ , \new_[4651]_ ,
    \new_[4652]_ , \new_[4653]_ , \new_[4654]_ , \new_[4655]_ ,
    \new_[4656]_ , \new_[4657]_ , \new_[4658]_ , \new_[4659]_ ,
    \new_[4660]_ , \new_[4661]_ , \new_[4662]_ , \new_[4663]_ ,
    \new_[4664]_ , \new_[4665]_ , \new_[4666]_ , \new_[4667]_ ,
    \new_[4668]_ , \new_[4669]_ , \new_[4670]_ , \new_[4671]_ ,
    \new_[4672]_ , \new_[4673]_ , \new_[4674]_ , \new_[4675]_ ,
    \new_[4676]_ , \new_[4677]_ , \new_[4678]_ , \new_[4679]_ ,
    \new_[4683]_ , \new_[4685]_ , \new_[4686]_ , \new_[4689]_ ,
    \new_[4690]_ , \new_[4691]_ , \new_[4693]_ , \new_[4694]_ ,
    \new_[4695]_ , \new_[4696]_ , \new_[4697]_ , \new_[4698]_ ,
    \new_[4699]_ , \new_[4700]_ , \new_[4701]_ , \new_[4702]_ ,
    \new_[4703]_ , \new_[4705]_ , \new_[4706]_ , \new_[4707]_ ,
    \new_[4709]_ , \new_[4710]_ , \new_[4711]_ , \new_[4712]_ ,
    \new_[4714]_ , \new_[4715]_ , \new_[4716]_ , \new_[4717]_ ,
    \new_[4718]_ , \new_[4719]_ , \new_[4720]_ , \new_[4721]_ ,
    \new_[4722]_ , \new_[4723]_ , \new_[4724]_ , \new_[4725]_ ,
    \new_[4726]_ , \new_[4727]_ , \new_[4728]_ , \new_[4729]_ ,
    \new_[4730]_ , \new_[4731]_ , \new_[4732]_ , \new_[4733]_ ,
    \new_[4734]_ , \new_[4735]_ , \new_[4736]_ , \new_[4737]_ ,
    \new_[4738]_ , \new_[4739]_ , \new_[4740]_ , \new_[4741]_ ,
    \new_[4742]_ , \new_[4743]_ , \new_[4744]_ , \new_[4745]_ ,
    \new_[4746]_ , \new_[4747]_ , \new_[4748]_ , \new_[4749]_ ,
    \new_[4750]_ , \new_[4751]_ , \new_[4752]_ , \new_[4753]_ ,
    \new_[4754]_ , \new_[4755]_ , \new_[4756]_ , \new_[4757]_ ,
    \new_[4758]_ , \new_[4759]_ , \new_[4760]_ , \new_[4761]_ ,
    \new_[4762]_ , \new_[4763]_ , \new_[4764]_ , \new_[4765]_ ,
    \new_[4766]_ , \new_[4767]_ , \new_[4768]_ , \new_[4772]_ ,
    \new_[4774]_ , \new_[4775]_ , \new_[4777]_ , \new_[4778]_ ,
    \new_[4779]_ , \new_[4780]_ , \new_[4781]_ , \new_[4782]_ ,
    \new_[4783]_ , \new_[4784]_ , \new_[4785]_ , \new_[4787]_ ,
    \new_[4788]_ , \new_[4789]_ , \new_[4790]_ , \new_[4791]_ ,
    \new_[4792]_ , \new_[4793]_ , \new_[4794]_ , \new_[4795]_ ,
    \new_[4796]_ , \new_[4797]_ , \new_[4798]_ , \new_[4799]_ ,
    \new_[4800]_ , \new_[4801]_ , \new_[4802]_ , \new_[4803]_ ,
    \new_[4804]_ , \new_[4805]_ , \new_[4806]_ , \new_[4807]_ ,
    \new_[4808]_ , \new_[4809]_ , \new_[4810]_ , \new_[4811]_ ,
    \new_[4812]_ , \new_[4813]_ , \new_[4814]_ , \new_[4815]_ ,
    \new_[4816]_ , \new_[4817]_ , \new_[4818]_ , \new_[4819]_ ,
    \new_[4820]_ , \new_[4821]_ , \new_[4822]_ , \new_[4823]_ ,
    \new_[4824]_ , \new_[4825]_ , \new_[4826]_ , \new_[4827]_ ,
    \new_[4828]_ , \new_[4829]_ , \new_[4830]_ , \new_[4831]_ ,
    \new_[4832]_ , \new_[4833]_ , \new_[4834]_ , \new_[4835]_ ,
    \new_[4836]_ , \new_[4837]_ , \new_[4838]_ , \new_[4839]_ ,
    \new_[4840]_ , \new_[4841]_ , \new_[4842]_ , \new_[4843]_ ,
    \new_[4844]_ , \new_[4845]_ , \new_[4846]_ , \new_[4847]_ ,
    \new_[4848]_ , \new_[4849]_ , \new_[4850]_ , \new_[4851]_ ,
    \new_[4852]_ , \new_[4853]_ , \new_[4854]_ , \new_[4855]_ ,
    \new_[4856]_ , \new_[4857]_ , \new_[4858]_ , \new_[4859]_ ,
    \new_[4860]_ , \new_[4861]_ , \new_[4862]_ , \new_[4863]_ ,
    \new_[4864]_ , \new_[4865]_ , \new_[4866]_ , \new_[4867]_ ,
    \new_[4868]_ , \new_[4869]_ , \new_[4870]_ , \new_[4871]_ ,
    \new_[4872]_ , \new_[4873]_ , \new_[4874]_ , \new_[4875]_ ,
    \new_[4876]_ , \new_[4877]_ , \new_[4878]_ , \new_[4879]_ ,
    \new_[4880]_ , \new_[4881]_ , \new_[4882]_ , \new_[4883]_ ,
    \new_[4884]_ , \new_[4885]_ , \new_[4886]_ , \new_[4887]_ ,
    \new_[4888]_ , \new_[4890]_ , \new_[4891]_ , \new_[4893]_ ,
    \new_[4894]_ , \new_[4895]_ , \new_[4896]_ , \new_[4897]_ ,
    \new_[4898]_ , \new_[4899]_ , \new_[4900]_ , \new_[4901]_ ,
    \new_[4902]_ , \new_[4903]_ , \new_[4904]_ , \new_[4905]_ ,
    \new_[4906]_ , \new_[4907]_ , \new_[4908]_ , \new_[4909]_ ,
    \new_[4910]_ , \new_[4911]_ , \new_[4912]_ , \new_[4913]_ ,
    \new_[4914]_ , \new_[4915]_ , \new_[4916]_ , \new_[4917]_ ,
    \new_[4918]_ , \new_[4920]_ , \new_[4921]_ , \new_[4922]_ ,
    \new_[4923]_ , \new_[4924]_ , \new_[4925]_ , \new_[4926]_ ,
    \new_[4927]_ , \new_[4928]_ , \new_[4929]_ , \new_[4930]_ ,
    \new_[4931]_ , \new_[4932]_ , \new_[4933]_ , \new_[4934]_ ,
    \new_[4935]_ , \new_[4936]_ , \new_[4937]_ , \new_[4938]_ ,
    \new_[4939]_ , \new_[4940]_ , \new_[4941]_ , \new_[4942]_ ,
    \new_[4943]_ , \new_[4945]_ , \new_[4947]_ , \new_[4948]_ ,
    \new_[4949]_ , \new_[4950]_ , \new_[4952]_ , \new_[4953]_ ,
    \new_[4954]_ , \new_[4955]_ , \new_[4956]_ , \new_[4958]_ ,
    \new_[4959]_ , \new_[4960]_ , \new_[4961]_ , \new_[4962]_ ,
    \new_[4963]_ , \new_[4964]_ , \new_[4965]_ , \new_[4966]_ ,
    \new_[4967]_ , \new_[4968]_ , \new_[4969]_ , \new_[4970]_ ,
    \new_[4971]_ , \new_[4972]_ , \new_[4973]_ , \new_[4974]_ ,
    \new_[4975]_ , \new_[4976]_ , \new_[4977]_ , \new_[4978]_ ,
    \new_[4979]_ , \new_[4980]_ , \new_[4981]_ , \new_[4982]_ ,
    \new_[4983]_ , \new_[4984]_ , \new_[4985]_ , \new_[4986]_ ,
    \new_[4987]_ , \new_[4988]_ , \new_[4989]_ , \new_[4990]_ ,
    \new_[4991]_ , \new_[4992]_ , \new_[4993]_ , \new_[4994]_ ,
    \new_[4995]_ , \new_[4996]_ , \new_[4997]_ , \new_[4998]_ ,
    \new_[4999]_ , \new_[5000]_ , \new_[5001]_ , \new_[5002]_ ,
    \new_[5003]_ , \new_[5004]_ , \new_[5005]_ , \new_[5006]_ ,
    \new_[5007]_ , \new_[5008]_ , \new_[5009]_ , \new_[5010]_ ,
    \new_[5011]_ , \new_[5012]_ , \new_[5013]_ , \new_[5014]_ ,
    \new_[5015]_ , \new_[5016]_ , \new_[5017]_ , \new_[5018]_ ,
    \new_[5019]_ , \new_[5020]_ , \new_[5021]_ , \new_[5022]_ ,
    \new_[5023]_ , \new_[5024]_ , \new_[5025]_ , \new_[5026]_ ,
    \new_[5027]_ , \new_[5028]_ , \new_[5029]_ , \new_[5030]_ ,
    \new_[5031]_ , \new_[5032]_ , \new_[5033]_ , \new_[5034]_ ,
    \new_[5035]_ , \new_[5036]_ , \new_[5039]_ , \new_[5040]_ ,
    \new_[5041]_ , \new_[5042]_ , \new_[5043]_ , \new_[5044]_ ,
    \new_[5045]_ , \new_[5046]_ , \new_[5047]_ , \new_[5048]_ ,
    \new_[5049]_ , \new_[5050]_ , \new_[5051]_ , \new_[5052]_ ,
    \new_[5053]_ , \new_[5054]_ , \new_[5055]_ , \new_[5056]_ ,
    \new_[5057]_ , \new_[5058]_ , \new_[5059]_ , \new_[5060]_ ,
    \new_[5061]_ , \new_[5062]_ , \new_[5063]_ , \new_[5064]_ ,
    \new_[5065]_ , \new_[5066]_ , \new_[5067]_ , \new_[5068]_ ,
    \new_[5069]_ , \new_[5070]_ , \new_[5071]_ , \new_[5072]_ ,
    \new_[5073]_ , \new_[5074]_ , \new_[5075]_ , \new_[5076]_ ,
    \new_[5077]_ , \new_[5078]_ , \new_[5079]_ , \new_[5080]_ ,
    \new_[5081]_ , \new_[5082]_ , \new_[5083]_ , \new_[5084]_ ,
    \new_[5085]_ , \new_[5086]_ , \new_[5087]_ , \new_[5088]_ ,
    \new_[5089]_ , \new_[5090]_ , \new_[5091]_ , \new_[5092]_ ,
    \new_[5093]_ , \new_[5094]_ , \new_[5095]_ , \new_[5096]_ ,
    \new_[5097]_ , \new_[5098]_ , \new_[5099]_ , \new_[5100]_ ,
    \new_[5101]_ , \new_[5102]_ , \new_[5103]_ , \new_[5104]_ ,
    \new_[5105]_ , \new_[5106]_ , \new_[5107]_ , \new_[5109]_ ,
    \new_[5111]_ , \new_[5112]_ , \new_[5123]_ , \new_[5124]_ ,
    \new_[5125]_ , \new_[5126]_ , \new_[5127]_ , \new_[5128]_ ,
    \new_[5129]_ , \new_[5130]_ , \new_[5131]_ , \new_[5132]_ ,
    \new_[5133]_ , \new_[5134]_ , \new_[5135]_ , \new_[5136]_ ,
    \new_[5137]_ , \new_[5138]_ , \new_[5139]_ , \new_[5140]_ ,
    \new_[5141]_ , \new_[5142]_ , \new_[5143]_ , \new_[5144]_ ,
    \new_[5145]_ , \new_[5146]_ , \new_[5147]_ , \new_[5148]_ ,
    \new_[5149]_ , \new_[5150]_ , \new_[5151]_ , \new_[5152]_ ,
    \new_[5153]_ , \new_[5154]_ , \new_[5155]_ , \new_[5156]_ ,
    \new_[5158]_ , \new_[5159]_ , \new_[5160]_ , \new_[5161]_ ,
    \new_[5162]_ , \new_[5163]_ , \new_[5164]_ , \new_[5165]_ ,
    \new_[5166]_ , \new_[5167]_ , \new_[5168]_ , \new_[5169]_ ,
    \new_[5170]_ , \new_[5171]_ , \new_[5172]_ , \new_[5173]_ ,
    \new_[5174]_ , \new_[5175]_ , \new_[5176]_ , \new_[5177]_ ,
    \new_[5178]_ , \new_[5179]_ , \new_[5180]_ , \new_[5181]_ ,
    \new_[5182]_ , \new_[5183]_ , \new_[5184]_ , \new_[5185]_ ,
    \new_[5186]_ , \new_[5187]_ , \new_[5189]_ , \new_[5190]_ ,
    \new_[5191]_ , \new_[5192]_ , \new_[5193]_ , \new_[5194]_ ,
    \new_[5195]_ , \new_[5196]_ , \new_[5197]_ , \new_[5198]_ ,
    \new_[5199]_ , \new_[5200]_ , \new_[5201]_ , \new_[5202]_ ,
    \new_[5203]_ , \new_[5204]_ , \new_[5205]_ , \new_[5206]_ ,
    \new_[5207]_ , \new_[5208]_ , \new_[5209]_ , \new_[5210]_ ,
    \new_[5211]_ , \new_[5212]_ , \new_[5213]_ , \new_[5214]_ ,
    \new_[5224]_ , \new_[5230]_ , \new_[5231]_ , \new_[5232]_ ,
    \new_[5233]_ , \new_[5234]_ , \new_[5235]_ , \new_[5236]_ ,
    \new_[5237]_ , \new_[5238]_ , \new_[5239]_ , \new_[5240]_ ,
    \new_[5241]_ , \new_[5242]_ , \new_[5243]_ , \new_[5244]_ ,
    \new_[5245]_ , \new_[5246]_ , \new_[5248]_ , \new_[5249]_ ,
    \new_[5250]_ , \new_[5251]_ , \new_[5260]_ , \new_[5289]_ ,
    \new_[5318]_ , \new_[5320]_ , \new_[5322]_ , \new_[5342]_ ,
    \new_[5348]_ , \new_[5349]_ , \new_[5351]_ , \new_[5352]_ ,
    \new_[5354]_ , \new_[5355]_ , \new_[5356]_ , \new_[5357]_ ,
    \new_[5358]_ , \new_[5359]_ , \new_[5360]_ , \new_[5361]_ ,
    \new_[5362]_ , \new_[5365]_ , \new_[5366]_ , \new_[5367]_ ,
    \new_[5368]_ , \new_[5369]_ , \new_[5370]_ , \new_[5371]_ ,
    \new_[5372]_ , \new_[5373]_ , \new_[5374]_ , \new_[5375]_ ,
    \new_[5376]_ , \new_[5377]_ , \new_[5378]_ , \new_[5379]_ ,
    \new_[5380]_ , \new_[5381]_ , \new_[5382]_ , \new_[5383]_ ,
    \new_[5384]_ , \new_[5385]_ , \new_[5386]_ , \new_[5387]_ ,
    \new_[5388]_ , \new_[5389]_ , \new_[5390]_ , \new_[5391]_ ,
    \new_[5392]_ , \new_[5393]_ , \new_[5394]_ , \new_[5395]_ ,
    \new_[5396]_ , \new_[5397]_ , \new_[5398]_ , \new_[5399]_ ,
    \new_[5400]_ , \new_[5402]_ , \new_[5403]_ , \new_[5404]_ ,
    \new_[5405]_ , \new_[5406]_ , \new_[5407]_ , \new_[5409]_ ,
    \new_[5410]_ , \new_[5411]_ , \new_[5412]_ , \new_[5413]_ ,
    \new_[5414]_ , \new_[5415]_ , \new_[5416]_ , \new_[5417]_ ,
    \new_[5418]_ , \new_[5419]_ , \new_[5420]_ , \new_[5421]_ ,
    \new_[5422]_ , \new_[5423]_ , \new_[5425]_ , \new_[5427]_ ,
    \new_[5428]_ , \new_[5429]_ , \new_[5430]_ , \new_[5431]_ ,
    \new_[5432]_ , \new_[5433]_ , \new_[5434]_ , \new_[5435]_ ,
    \new_[5436]_ , \new_[5437]_ , \new_[5438]_ , \new_[5439]_ ,
    \new_[5440]_ , \new_[5441]_ , \new_[5442]_ , \new_[5443]_ ,
    \new_[5444]_ , \new_[5445]_ , \new_[5446]_ , \new_[5447]_ ,
    \new_[5448]_ , \new_[5449]_ , \new_[5450]_ , \new_[5451]_ ,
    \new_[5452]_ , \new_[5453]_ , \new_[5454]_ , \new_[5455]_ ,
    \new_[5456]_ , \new_[5457]_ , \new_[5458]_ , \new_[5459]_ ,
    \new_[5460]_ , \new_[5461]_ , \new_[5462]_ , \new_[5463]_ ,
    \new_[5464]_ , \new_[5465]_ , \new_[5466]_ , \new_[5467]_ ,
    \new_[5468]_ , \new_[5469]_ , \new_[5470]_ , \new_[5471]_ ,
    \new_[5472]_ , \new_[5473]_ , \new_[5474]_ , \new_[5475]_ ,
    \new_[5478]_ , \new_[5481]_ , \new_[5482]_ , \new_[5483]_ ,
    \new_[5484]_ , \new_[5485]_ , \new_[5486]_ , \new_[5489]_ ,
    \new_[5490]_ , \new_[5491]_ , \new_[5492]_ , \new_[5495]_ ,
    \new_[5496]_ , \new_[5497]_ , \new_[5499]_ , \new_[5500]_ ,
    \new_[5501]_ , \new_[5502]_ , \new_[5503]_ , \new_[5504]_ ,
    \new_[5506]_ , \new_[5507]_ , \new_[5508]_ , \new_[5509]_ ,
    \new_[5510]_ , \new_[5511]_ , \new_[5512]_ , \new_[5514]_ ,
    \new_[5518]_ , \new_[5519]_ , \new_[5520]_ , \new_[5525]_ ,
    \new_[5527]_ , \new_[5528]_ , \new_[5529]_ , \new_[5530]_ ,
    \new_[5531]_ , \new_[5532]_ , \new_[5533]_ , \new_[5534]_ ,
    \new_[5538]_ , \new_[5539]_ , \new_[5540]_ , \new_[5541]_ ,
    \new_[5542]_ , \new_[5543]_ , \new_[5544]_ , \new_[5545]_ ,
    \new_[5546]_ , \new_[5547]_ , \new_[5548]_ , \new_[5549]_ ,
    \new_[5550]_ , \new_[5551]_ , \new_[5552]_ , \new_[5553]_ ,
    \new_[5554]_ , \new_[5555]_ , \new_[5556]_ , \new_[5557]_ ,
    \new_[5558]_ , \new_[5559]_ , \new_[5560]_ , \new_[5562]_ ,
    \new_[5563]_ , \new_[5564]_ , \new_[5565]_ , \new_[5567]_ ,
    \new_[5568]_ , \new_[5575]_ , \new_[5576]_ , \new_[5581]_ ,
    \new_[5582]_ , \new_[5583]_ , \new_[5585]_ , \new_[5586]_ ,
    \new_[5588]_ , \new_[5589]_ , \new_[5590]_ , \new_[5591]_ ,
    \new_[5592]_ , \new_[5599]_ , \new_[5601]_ , \new_[5602]_ ,
    \new_[5603]_ , \new_[5604]_ , \new_[5605]_ , \new_[5607]_ ,
    \new_[5612]_ , \new_[5613]_ , \new_[5614]_ , \new_[5616]_ ,
    \new_[5617]_ , \new_[5618]_ , \new_[5619]_ , \new_[5620]_ ,
    \new_[5621]_ , \new_[5622]_ , \new_[5623]_ , \new_[5624]_ ,
    \new_[5625]_ , \new_[5626]_ , \new_[5627]_ , \new_[5628]_ ,
    \new_[5629]_ , \new_[5630]_ , \new_[5631]_ , \new_[5632]_ ,
    \new_[5633]_ , \new_[5634]_ , \new_[5635]_ , \new_[5636]_ ,
    \new_[5637]_ , \new_[5638]_ , \new_[5639]_ , \new_[5640]_ ,
    \new_[5641]_ , \new_[5642]_ , \new_[5643]_ , \new_[5644]_ ,
    \new_[5645]_ , \new_[5646]_ , \new_[5647]_ , \new_[5672]_ ,
    \new_[5673]_ , \new_[5674]_ , \new_[5675]_ , \new_[5676]_ ,
    \new_[5677]_ , \new_[5678]_ , \new_[5679]_ , \new_[5680]_ ,
    \new_[5681]_ , \new_[5682]_ , \new_[5683]_ , \new_[5684]_ ,
    \new_[5685]_ , \new_[5686]_ , \new_[5687]_ , \new_[5688]_ ,
    \new_[5689]_ , \new_[5690]_ , \new_[5691]_ , \new_[5692]_ ,
    \new_[5693]_ , \new_[5694]_ , \new_[5698]_ , \new_[5699]_ ,
    \new_[5700]_ , \new_[5701]_ , \new_[5702]_ , \new_[5703]_ ,
    \new_[5704]_ , \new_[5705]_ , \new_[5706]_ , \new_[5707]_ ,
    \new_[5708]_ , \new_[5709]_ , \new_[5710]_ , \new_[5711]_ ,
    \new_[5712]_ , \new_[5713]_ , \new_[5715]_ , \new_[5716]_ ,
    \new_[5717]_ , \new_[5718]_ , \new_[5719]_ , \new_[5720]_ ,
    \new_[5721]_ , \new_[5722]_ , \new_[5723]_ , \new_[5725]_ ,
    \new_[5726]_ , \new_[5727]_ , \new_[5728]_ , \new_[5729]_ ,
    \new_[5730]_ , \new_[5731]_ , \new_[5732]_ , \new_[5733]_ ,
    \new_[5734]_ , \new_[5735]_ , \new_[5736]_ , \new_[5737]_ ,
    \new_[5738]_ , \new_[5739]_ , \new_[5740]_ , \new_[5741]_ ,
    \new_[5742]_ , \new_[5743]_ , \new_[5744]_ , \new_[5745]_ ,
    \new_[5746]_ , \new_[5747]_ , \new_[5748]_ , \new_[5753]_ ,
    \new_[5754]_ , \new_[5756]_ , \new_[5757]_ , \new_[5760]_ ,
    \new_[5761]_ , \new_[5762]_ , \new_[5763]_ , \new_[5764]_ ,
    \new_[5765]_ , \new_[5766]_ , \new_[5767]_ , \new_[5768]_ ,
    \new_[5769]_ , \new_[5770]_ , \new_[5774]_ , \new_[5776]_ ,
    \new_[5777]_ , \new_[5778]_ , \new_[5782]_ , \new_[5783]_ ,
    \new_[5784]_ , \new_[5785]_ , \new_[5787]_ , \new_[5788]_ ,
    \new_[5789]_ , \new_[5791]_ , \new_[5793]_ , \new_[5796]_ ,
    \new_[5797]_ , \new_[5798]_ , \new_[5799]_ , \new_[5800]_ ,
    \new_[5801]_ , \new_[5802]_ , \new_[5803]_ , \new_[5804]_ ,
    \new_[5805]_ , \new_[5806]_ , \new_[5807]_ , \new_[5808]_ ,
    \new_[5809]_ , \new_[5810]_ , \new_[5811]_ , \new_[5812]_ ,
    \new_[5813]_ , \new_[5814]_ , \new_[5815]_ , \new_[5816]_ ,
    \new_[5817]_ , \new_[5818]_ , \new_[5819]_ , \new_[5820]_ ,
    \new_[5821]_ , \new_[5822]_ , \new_[5823]_ , \new_[5824]_ ,
    \new_[5825]_ , \new_[5826]_ , \new_[5827]_ , \new_[5828]_ ,
    \new_[5829]_ , \new_[5830]_ , \new_[5831]_ , \new_[5832]_ ,
    \new_[5833]_ , \new_[5834]_ , \new_[5835]_ , \new_[5836]_ ,
    \new_[5837]_ , \new_[5838]_ , \new_[5839]_ , \new_[5840]_ ,
    \new_[5841]_ , \new_[5842]_ , \new_[5843]_ , \new_[5844]_ ,
    \new_[5845]_ , \new_[5847]_ , \new_[5848]_ , \new_[5849]_ ,
    \new_[5850]_ , \new_[5851]_ , \new_[5852]_ , \new_[5853]_ ,
    \new_[5855]_ , \new_[5856]_ , \new_[5857]_ , \new_[5858]_ ,
    \new_[5859]_ , \new_[5860]_ , \new_[5881]_ , \new_[5882]_ ,
    \new_[5883]_ , \new_[5884]_ , \new_[5885]_ , \new_[5886]_ ,
    \new_[5888]_ , \new_[5889]_ , \new_[5890]_ , \new_[5891]_ ,
    \new_[5892]_ , \new_[5894]_ , \new_[5895]_ , \new_[5896]_ ,
    \new_[5897]_ , \new_[5898]_ , \new_[5899]_ , \new_[5900]_ ,
    \new_[5902]_ , \new_[5903]_ , \new_[5905]_ , \new_[5906]_ ,
    \new_[5907]_ , \new_[5908]_ , \new_[5912]_ , \new_[5913]_ ,
    \new_[5914]_ , \new_[5915]_ , \new_[5916]_ , \new_[5917]_ ,
    \new_[5918]_ , \new_[5919]_ , \new_[5920]_ , \new_[5921]_ ,
    \new_[5922]_ , \new_[5923]_ , \new_[5924]_ , \new_[5925]_ ,
    \new_[5926]_ , \new_[5927]_ , \new_[5928]_ , \new_[5929]_ ,
    \new_[5930]_ , \new_[5931]_ , \new_[5932]_ , \new_[5937]_ ,
    \new_[5938]_ , \new_[5939]_ , \new_[5941]_ , \new_[5942]_ ,
    \new_[5943]_ , \new_[5944]_ , \new_[5945]_ , \new_[5947]_ ,
    \new_[5948]_ , \new_[5949]_ , \new_[5950]_ , \new_[5951]_ ,
    \new_[5952]_ , \new_[5953]_ , \new_[5954]_ , \new_[5955]_ ,
    \new_[5956]_ , \new_[5957]_ , \new_[5959]_ , \new_[5960]_ ,
    \new_[5961]_ , \new_[5962]_ , \new_[5964]_ , \new_[5965]_ ,
    \new_[5966]_ , \new_[5967]_ , \new_[5968]_ , \new_[5969]_ ,
    \new_[5970]_ , \new_[5971]_ , \new_[5972]_ , \new_[5973]_ ,
    \new_[5976]_ , \new_[5978]_ , \new_[5980]_ , \new_[5981]_ ,
    \new_[5982]_ , \new_[5983]_ , \new_[5984]_ , \new_[5985]_ ,
    \new_[5986]_ , \new_[5987]_ , \new_[5988]_ , \new_[5989]_ ,
    \new_[5990]_ , \new_[5991]_ , \new_[5992]_ , \new_[5993]_ ,
    \new_[5994]_ , \new_[5996]_ , \new_[5997]_ , \new_[5998]_ ,
    \new_[5999]_ , \new_[6000]_ , \new_[6001]_ , \new_[6002]_ ,
    \new_[6003]_ , \new_[6004]_ , \new_[6005]_ , \new_[6006]_ ,
    \new_[6007]_ , \new_[6008]_ , \new_[6009]_ , \new_[6010]_ ,
    \new_[6011]_ , \new_[6012]_ , \new_[6013]_ , \new_[6015]_ ,
    \new_[6016]_ , \new_[6017]_ , \new_[6018]_ , \new_[6019]_ ,
    \new_[6020]_ , \new_[6021]_ , \new_[6022]_ , \new_[6023]_ ,
    \new_[6024]_ , \new_[6025]_ , \new_[6026]_ , \new_[6027]_ ,
    \new_[6028]_ , \new_[6029]_ , \new_[6031]_ , \new_[6032]_ ,
    \new_[6033]_ , \new_[6034]_ , \new_[6035]_ , \new_[6036]_ ,
    \new_[6037]_ , \new_[6038]_ , \new_[6039]_ , \new_[6040]_ ,
    \new_[6041]_ , \new_[6042]_ , \new_[6043]_ , \new_[6044]_ ,
    \new_[6045]_ , \new_[6046]_ , \new_[6047]_ , \new_[6048]_ ,
    \new_[6049]_ , \new_[6050]_ , \new_[6051]_ , \new_[6052]_ ,
    \new_[6053]_ , \new_[6054]_ , \new_[6055]_ , \new_[6056]_ ,
    \new_[6057]_ , \new_[6058]_ , \new_[6059]_ , \new_[6061]_ ,
    \new_[6063]_ , \new_[6064]_ , \new_[6065]_ , \new_[6067]_ ,
    \new_[6068]_ , \new_[6070]_ , \new_[6071]_ , \new_[6072]_ ,
    \new_[6073]_ , \new_[6075]_ , \new_[6080]_ , \new_[6081]_ ,
    \new_[6082]_ , \new_[6083]_ , \new_[6084]_ , \new_[6085]_ ,
    \new_[6086]_ , \new_[6087]_ , \new_[6088]_ , \new_[6089]_ ,
    \new_[6090]_ , \new_[6091]_ , \new_[6092]_ , \new_[6093]_ ,
    \new_[6094]_ , \new_[6095]_ , \new_[6096]_ , \new_[6097]_ ,
    \new_[6098]_ , \new_[6099]_ , \new_[6100]_ , \new_[6101]_ ,
    \new_[6102]_ , \new_[6103]_ , \new_[6104]_ , \new_[6105]_ ,
    \new_[6106]_ , \new_[6107]_ , \new_[6108]_ , \new_[6109]_ ,
    \new_[6110]_ , \new_[6111]_ , \new_[6112]_ , \new_[6113]_ ,
    \new_[6114]_ , \new_[6115]_ , \new_[6116]_ , \new_[6117]_ ,
    \new_[6118]_ , \new_[6119]_ , \new_[6120]_ , \new_[6121]_ ,
    \new_[6122]_ , \new_[6126]_ , \new_[6127]_ , \new_[6128]_ ,
    \new_[6129]_ , \new_[6130]_ , \new_[6131]_ , \new_[6132]_ ,
    \new_[6133]_ , \new_[6134]_ , \new_[6135]_ , \new_[6136]_ ,
    \new_[6137]_ , \new_[6138]_ , \new_[6139]_ , \new_[6140]_ ,
    \new_[6141]_ , \new_[6142]_ , \new_[6143]_ , \new_[6144]_ ,
    \new_[6145]_ , \new_[6146]_ , \new_[6147]_ , \new_[6148]_ ,
    \new_[6149]_ , \new_[6150]_ , \new_[6151]_ , \new_[6152]_ ,
    \new_[6153]_ , \new_[6154]_ , \new_[6155]_ , \new_[6156]_ ,
    \new_[6157]_ , \new_[6158]_ , \new_[6159]_ , \new_[6160]_ ,
    \new_[6161]_ , \new_[6162]_ , \new_[6163]_ , \new_[6164]_ ,
    \new_[6165]_ , \new_[6166]_ , \new_[6168]_ , \new_[6169]_ ,
    \new_[6170]_ , \new_[6171]_ , \new_[6172]_ , \new_[6173]_ ,
    \new_[6174]_ , \new_[6175]_ , \new_[6176]_ , \new_[6177]_ ,
    \new_[6178]_ , \new_[6179]_ , \new_[6180]_ , \new_[6182]_ ,
    \new_[6183]_ , \new_[6184]_ , \new_[6185]_ , \new_[6186]_ ,
    \new_[6189]_ , \new_[6190]_ , \new_[6191]_ , \new_[6192]_ ,
    \new_[6193]_ , \new_[6194]_ , \new_[6195]_ , \new_[6196]_ ,
    \new_[6197]_ , \new_[6198]_ , \new_[6199]_ , \new_[6200]_ ,
    \new_[6202]_ , \new_[6203]_ , \new_[6204]_ , \new_[6205]_ ,
    \new_[6206]_ , \new_[6207]_ , \new_[6208]_ , \new_[6209]_ ,
    \new_[6210]_ , \new_[6211]_ , \new_[6212]_ , \new_[6216]_ ,
    \new_[6217]_ , \new_[6219]_ , \new_[6220]_ , \new_[6221]_ ,
    \new_[6222]_ , \new_[6223]_ , \new_[6224]_ , \new_[6225]_ ,
    \new_[6226]_ , \new_[6227]_ , \new_[6228]_ , \new_[6229]_ ,
    \new_[6230]_ , \new_[6231]_ , \new_[6232]_ , \new_[6233]_ ,
    \new_[6234]_ , \new_[6235]_ , \new_[6236]_ , \new_[6237]_ ,
    \new_[6238]_ , \new_[6239]_ , \new_[6240]_ , \new_[6241]_ ,
    \new_[6242]_ , \new_[6243]_ , \new_[6245]_ , \new_[6246]_ ,
    \new_[6247]_ , \new_[6248]_ , \new_[6249]_ , \new_[6250]_ ,
    \new_[6251]_ , \new_[6252]_ , \new_[6253]_ , \new_[6254]_ ,
    \new_[6255]_ , \new_[6256]_ , \new_[6257]_ , \new_[6258]_ ,
    \new_[6259]_ , \new_[6260]_ , \new_[6261]_ , \new_[6262]_ ,
    \new_[6263]_ , \new_[6264]_ , \new_[6265]_ , \new_[6266]_ ,
    \new_[6267]_ , \new_[6268]_ , \new_[6269]_ , \new_[6270]_ ,
    \new_[6271]_ , \new_[6272]_ , \new_[6273]_ , \new_[6274]_ ,
    \new_[6275]_ , \new_[6276]_ , \new_[6277]_ , \new_[6278]_ ,
    \new_[6279]_ , \new_[6280]_ , \new_[6281]_ , \new_[6282]_ ,
    \new_[6283]_ , \new_[6284]_ , \new_[6285]_ , \new_[6286]_ ,
    \new_[6287]_ , \new_[6288]_ , \new_[6289]_ , \new_[6290]_ ,
    \new_[6291]_ , \new_[6292]_ , \new_[6293]_ , \new_[6294]_ ,
    \new_[6295]_ , \new_[6296]_ , \new_[6297]_ , \new_[6298]_ ,
    \new_[6299]_ , \new_[6300]_ , \new_[6301]_ , \new_[6302]_ ,
    \new_[6303]_ , \new_[6304]_ , \new_[6305]_ , \new_[6306]_ ,
    \new_[6307]_ , \new_[6308]_ , \new_[6309]_ , \new_[6310]_ ,
    \new_[6311]_ , \new_[6312]_ , \new_[6313]_ , \new_[6314]_ ,
    \new_[6315]_ , \new_[6316]_ , \new_[6317]_ , \new_[6318]_ ,
    \new_[6319]_ , \new_[6320]_ , \new_[6321]_ , \new_[6322]_ ,
    \new_[6323]_ , \new_[6324]_ , \new_[6325]_ , \new_[6326]_ ,
    \new_[6327]_ , \new_[6328]_ , \new_[6329]_ , \new_[6330]_ ,
    \new_[6331]_ , \new_[6332]_ , \new_[6333]_ , \new_[6334]_ ,
    \new_[6335]_ , \new_[6336]_ , \new_[6337]_ , \new_[6338]_ ,
    \new_[6339]_ , \new_[6340]_ , \new_[6341]_ , \new_[6342]_ ,
    \new_[6343]_ , \new_[6344]_ , \new_[6345]_ , \new_[6346]_ ,
    \new_[6347]_ , \new_[6348]_ , \new_[6349]_ , \new_[6350]_ ,
    \new_[6351]_ , \new_[6352]_ , \new_[6353]_ , \new_[6354]_ ,
    \new_[6355]_ , \new_[6356]_ , \new_[6357]_ , \new_[6358]_ ,
    \new_[6359]_ , \new_[6360]_ , \new_[6361]_ , \new_[6362]_ ,
    \new_[6363]_ , \new_[6364]_ , \new_[6365]_ , \new_[6366]_ ,
    \new_[6367]_ , \new_[6368]_ , \new_[6369]_ , \new_[6370]_ ,
    \new_[6371]_ , \new_[6372]_ , \new_[6373]_ , \new_[6374]_ ,
    \new_[6375]_ , \new_[6376]_ , \new_[6377]_ , \new_[6378]_ ,
    \new_[6379]_ , \new_[6381]_ , \new_[6382]_ , \new_[6383]_ ,
    \new_[6384]_ , \new_[6385]_ , \new_[6386]_ , \new_[6387]_ ,
    \new_[6388]_ , \new_[6389]_ , \new_[6390]_ , \new_[6391]_ ,
    \new_[6392]_ , \new_[6393]_ , \new_[6394]_ , \new_[6395]_ ,
    \new_[6396]_ , \new_[6397]_ , \new_[6398]_ , \new_[6399]_ ,
    \new_[6400]_ , \new_[6401]_ , \new_[6402]_ , \new_[6403]_ ,
    \new_[6404]_ , \new_[6405]_ , \new_[6406]_ , \new_[6407]_ ,
    \new_[6408]_ , \new_[6409]_ , \new_[6410]_ , \new_[6411]_ ,
    \new_[6412]_ , \new_[6413]_ , \new_[6414]_ , \new_[6415]_ ,
    \new_[6416]_ , \new_[6417]_ , \new_[6418]_ , \new_[6419]_ ,
    \new_[6420]_ , \new_[6421]_ , \new_[6422]_ , \new_[6423]_ ,
    \new_[6424]_ , \new_[6425]_ , \new_[6426]_ , \new_[6427]_ ,
    \new_[6428]_ , \new_[6429]_ , \new_[6430]_ , \new_[6431]_ ,
    \new_[6432]_ , \new_[6433]_ , \new_[6434]_ , \new_[6435]_ ,
    \new_[6436]_ , \new_[6437]_ , \new_[6438]_ , \new_[6439]_ ,
    \new_[6440]_ , \new_[6441]_ , \new_[6442]_ , \new_[6443]_ ,
    \new_[6444]_ , \new_[6445]_ , \new_[6446]_ , \new_[6447]_ ,
    \new_[6448]_ , \new_[6449]_ , \new_[6450]_ , \new_[6451]_ ,
    \new_[6452]_ , \new_[6453]_ , \new_[6454]_ , \new_[6455]_ ,
    \new_[6456]_ , \new_[6457]_ , \new_[6458]_ , \new_[6459]_ ,
    \new_[6460]_ , \new_[6461]_ , \new_[6462]_ , \new_[6463]_ ,
    \new_[6464]_ , \new_[6465]_ , \new_[6466]_ , \new_[6467]_ ,
    \new_[6468]_ , \new_[6469]_ , \new_[6470]_ , \new_[6475]_ ,
    \new_[6476]_ , \new_[6477]_ , \new_[6478]_ , \new_[6480]_ ,
    \new_[6481]_ , \new_[6482]_ , \new_[6483]_ , \new_[6484]_ ,
    \new_[6485]_ , \new_[6486]_ , \new_[6487]_ , \new_[6488]_ ,
    \new_[6489]_ , \new_[6490]_ , \new_[6491]_ , \new_[6492]_ ,
    \new_[6493]_ , \new_[6494]_ , \new_[6495]_ , \new_[6496]_ ,
    \new_[6497]_ , \new_[6498]_ , \new_[6499]_ , \new_[6500]_ ,
    \new_[6501]_ , \new_[6502]_ , \new_[6503]_ , \new_[6504]_ ,
    \new_[6505]_ , \new_[6506]_ , \new_[6507]_ , \new_[6508]_ ,
    \new_[6509]_ , \new_[6510]_ , \new_[6511]_ , \new_[6512]_ ,
    \new_[6513]_ , \new_[6514]_ , \new_[6515]_ , \new_[6516]_ ,
    \new_[6517]_ , \new_[6518]_ , \new_[6519]_ , \new_[6520]_ ,
    \new_[6521]_ , \new_[6522]_ , \new_[6523]_ , \new_[6524]_ ,
    \new_[6525]_ , \new_[6526]_ , \new_[6527]_ , \new_[6528]_ ,
    \new_[6529]_ , \new_[6531]_ , \new_[6532]_ , \new_[6534]_ ,
    \new_[6535]_ , \new_[6536]_ , \new_[6538]_ , \new_[6539]_ ,
    \new_[6540]_ , \new_[6541]_ , \new_[6542]_ , \new_[6543]_ ,
    \new_[6544]_ , \new_[6545]_ , \new_[6546]_ , \new_[6547]_ ,
    \new_[6548]_ , \new_[6549]_ , \new_[6550]_ , \new_[6551]_ ,
    \new_[6552]_ , \new_[6555]_ , \new_[6556]_ , \new_[6557]_ ,
    \new_[6558]_ , \new_[6559]_ , \new_[6560]_ , \new_[6561]_ ,
    \new_[6562]_ , \new_[6563]_ , \new_[6564]_ , \new_[6565]_ ,
    \new_[6566]_ , \new_[6567]_ , \new_[6575]_ , \new_[6586]_ ,
    \new_[6587]_ , \new_[6588]_ , \new_[6589]_ , \new_[6590]_ ,
    \new_[6591]_ , \new_[6592]_ , \new_[6593]_ , \new_[6594]_ ,
    \new_[6596]_ , \new_[6597]_ , \new_[6598]_ , \new_[6599]_ ,
    \new_[6600]_ , \new_[6601]_ , \new_[6602]_ , \new_[6603]_ ,
    \new_[6604]_ , \new_[6605]_ , \new_[6606]_ , \new_[6607]_ ,
    \new_[6608]_ , \new_[6609]_ , \new_[6610]_ , \new_[6611]_ ,
    \new_[6612]_ , \new_[6613]_ , \new_[6614]_ , \new_[6615]_ ,
    \new_[6616]_ , \new_[6617]_ , \new_[6618]_ , \new_[6619]_ ,
    \new_[6620]_ , \new_[6621]_ , \new_[6622]_ , \new_[6623]_ ,
    \new_[6624]_ , \new_[6625]_ , \new_[6626]_ , \new_[6627]_ ,
    \new_[6628]_ , \new_[6629]_ , \new_[6630]_ , \new_[6631]_ ,
    \new_[6632]_ , \new_[6633]_ , \new_[6634]_ , \new_[6635]_ ,
    \new_[6636]_ , \new_[6637]_ , \new_[6638]_ , \new_[6639]_ ,
    \new_[6640]_ , \new_[6641]_ , \new_[6642]_ , \new_[6643]_ ,
    \new_[6644]_ , \new_[6645]_ , \new_[6646]_ , \new_[6647]_ ,
    \new_[6648]_ , \new_[6649]_ , \new_[6651]_ , \new_[6652]_ ,
    \new_[6653]_ , \new_[6654]_ , \new_[6660]_ , \new_[6661]_ ,
    \new_[6662]_ , \new_[6663]_ , \new_[6666]_ , \new_[6671]_ ,
    \new_[6672]_ , \new_[6673]_ , \new_[6674]_ , \new_[6680]_ ,
    \new_[6681]_ , \new_[6683]_ , \new_[6684]_ , \new_[6687]_ ,
    \new_[6688]_ , \new_[6689]_ , \new_[6690]_ , \new_[6691]_ ,
    \new_[6692]_ , \new_[6693]_ , \new_[6694]_ , \new_[6695]_ ,
    \new_[6696]_ , \new_[6697]_ , \new_[6698]_ , \new_[6699]_ ,
    \new_[6700]_ , \new_[6701]_ , \new_[6702]_ , \new_[6703]_ ,
    \new_[6704]_ , \new_[6705]_ , \new_[6706]_ , \new_[6707]_ ,
    \new_[6708]_ , \new_[6710]_ , \new_[6716]_ , \new_[6717]_ ,
    \new_[6718]_ , \new_[6719]_ , \new_[6721]_ , \new_[6722]_ ,
    \new_[6723]_ , \new_[6724]_ , \new_[6725]_ , \new_[6726]_ ,
    \new_[6727]_ , \new_[6728]_ , \new_[6729]_ , \new_[6730]_ ,
    \new_[6731]_ , \new_[6732]_ , \new_[6733]_ , \new_[6734]_ ,
    \new_[6735]_ , \new_[6736]_ , \new_[6737]_ , \new_[6738]_ ,
    \new_[6739]_ , \new_[6740]_ , \new_[6741]_ , \new_[6742]_ ,
    \new_[6743]_ , \new_[6752]_ , \new_[6753]_ , \new_[6754]_ ,
    \new_[6755]_ , \new_[6756]_ , \new_[6757]_ , \new_[6758]_ ,
    \new_[6759]_ , \new_[6760]_ , \new_[6761]_ , \new_[6762]_ ,
    \new_[6763]_ , \new_[6764]_ , \new_[6765]_ , \new_[6766]_ ,
    \new_[6767]_ , \new_[6768]_ , \new_[6769]_ , \new_[6770]_ ,
    \new_[6771]_ , \new_[6772]_ , \new_[6773]_ , \new_[6774]_ ,
    \new_[6775]_ , \new_[6776]_ , \new_[6777]_ , \new_[6778]_ ,
    \new_[6779]_ , \new_[6780]_ , \new_[6781]_ , \new_[6782]_ ,
    \new_[6783]_ , \new_[6784]_ , \new_[6785]_ , \new_[6786]_ ,
    \new_[6787]_ , \new_[6788]_ , \new_[6789]_ , \new_[6790]_ ,
    \new_[6791]_ , \new_[6792]_ , \new_[6793]_ , \new_[6794]_ ,
    \new_[6795]_ , \new_[6796]_ , \new_[6797]_ , \new_[6798]_ ,
    \new_[6799]_ , \new_[6800]_ , \new_[6801]_ , \new_[6802]_ ,
    \new_[6803]_ , \new_[6804]_ , \new_[6805]_ , \new_[6806]_ ,
    \new_[6807]_ , \new_[6808]_ , \new_[6809]_ , \new_[6810]_ ,
    \new_[6811]_ , \new_[6812]_ , \new_[6813]_ , \new_[6814]_ ,
    \new_[6815]_ , \new_[6816]_ , \new_[6817]_ , \new_[6818]_ ,
    \new_[6819]_ , \new_[6820]_ , \new_[6821]_ , \new_[6822]_ ,
    \new_[6823]_ , \new_[6824]_ , \new_[6825]_ , \new_[6826]_ ,
    \new_[6827]_ , \new_[6828]_ , \new_[6829]_ , \new_[6830]_ ,
    \new_[6831]_ , \new_[6832]_ , \new_[6833]_ , \new_[6834]_ ,
    \new_[6835]_ , \new_[6836]_ , \new_[6837]_ , \new_[6838]_ ,
    \new_[6839]_ , \new_[6840]_ , \new_[6841]_ , \new_[6842]_ ,
    \new_[6843]_ , \new_[6844]_ , \new_[6845]_ , \new_[6846]_ ,
    \new_[6847]_ , \new_[6848]_ , \new_[6849]_ , \new_[6850]_ ,
    \new_[6851]_ , \new_[6852]_ , \new_[6853]_ , \new_[6854]_ ,
    \new_[6855]_ , \new_[6856]_ , \new_[6857]_ , \new_[6858]_ ,
    \new_[6860]_ , \new_[6861]_ , \new_[6862]_ , \new_[6863]_ ,
    \new_[6864]_ , \new_[6865]_ , \new_[6866]_ , \new_[6867]_ ,
    \new_[6868]_ , \new_[6869]_ , \new_[6870]_ , \new_[6871]_ ,
    \new_[6872]_ , \new_[6873]_ , \new_[6874]_ , \new_[6875]_ ,
    \new_[6876]_ , \new_[6877]_ , \new_[6878]_ , \new_[6879]_ ,
    \new_[6880]_ , \new_[6881]_ , \new_[6882]_ , \new_[6883]_ ,
    \new_[6884]_ , \new_[6894]_ , \new_[6895]_ , \new_[6896]_ ,
    \new_[6897]_ , \new_[6898]_ , \new_[6899]_ , \new_[6900]_ ,
    \new_[6901]_ , \new_[6902]_ , \new_[6903]_ , \new_[6904]_ ,
    \new_[6905]_ , \new_[6906]_ , \new_[6907]_ , \new_[6908]_ ,
    \new_[6909]_ , \new_[6910]_ , \new_[6911]_ , \new_[6912]_ ,
    \new_[6934]_ , \new_[6956]_ , \new_[6959]_ , \new_[6963]_ ,
    \new_[7016]_ , \new_[7070]_ , \new_[7071]_ , \new_[7123]_ ,
    \new_[7125]_ , \new_[7130]_ , \new_[7131]_ , \new_[7132]_ ,
    \new_[7133]_ , \new_[7134]_ , \new_[7136]_ , \new_[7137]_ ,
    \new_[7138]_ , \new_[7139]_ , \new_[7141]_ , \new_[7142]_ ,
    \new_[7143]_ , \new_[7144]_ , \new_[7145]_ , \new_[7146]_ ,
    \new_[7147]_ , \new_[7148]_ , \new_[7149]_ , \new_[7150]_ ,
    \new_[7151]_ , \new_[7152]_ , \new_[7153]_ , \new_[7154]_ ,
    \new_[7155]_ , \new_[7156]_ , \new_[7157]_ , \new_[7158]_ ,
    \new_[7159]_ , \new_[7160]_ , \new_[7161]_ , \new_[7162]_ ,
    \new_[7163]_ , \new_[7164]_ , \new_[7166]_ , \new_[7167]_ ,
    \new_[7168]_ , \new_[7169]_ , \new_[7170]_ , \new_[7171]_ ,
    \new_[7172]_ , \new_[7173]_ , \new_[7174]_ , \new_[7175]_ ,
    \new_[7176]_ , \new_[7177]_ , \new_[7178]_ , \new_[7179]_ ,
    \new_[7180]_ , \new_[7181]_ , \new_[7182]_ , \new_[7183]_ ,
    \new_[7184]_ , \new_[7185]_ , \new_[7186]_ , \new_[7187]_ ,
    \new_[7188]_ , \new_[7189]_ , \new_[7190]_ , \new_[7191]_ ,
    \new_[7192]_ , \new_[7193]_ , \new_[7194]_ , \new_[7195]_ ,
    \new_[7196]_ , \new_[7197]_ , \new_[7198]_ , \new_[7199]_ ,
    \new_[7200]_ , \new_[7201]_ , \new_[7202]_ , \new_[7203]_ ,
    \new_[7204]_ , \new_[7205]_ , \new_[7206]_ , \new_[7207]_ ,
    \new_[7208]_ , \new_[7209]_ , \new_[7210]_ , \new_[7211]_ ,
    \new_[7212]_ , \new_[7213]_ , \new_[7214]_ , \new_[7215]_ ,
    \new_[7216]_ , \new_[7217]_ , \new_[7218]_ , \new_[7219]_ ,
    \new_[7220]_ , \new_[7221]_ , \new_[7222]_ , \new_[7223]_ ,
    \new_[7224]_ , \new_[7225]_ , \new_[7226]_ , \new_[7227]_ ,
    \new_[7228]_ , \new_[7229]_ , \new_[7230]_ , \new_[7231]_ ,
    \new_[7232]_ , \new_[7233]_ , \new_[7234]_ , \new_[7235]_ ,
    \new_[7236]_ , \new_[7237]_ , \new_[7238]_ , \new_[7239]_ ,
    \new_[7240]_ , \new_[7241]_ , \new_[7242]_ , \new_[7243]_ ,
    \new_[7244]_ , \new_[7245]_ , \new_[7246]_ , \new_[7247]_ ,
    \new_[7248]_ , \new_[7249]_ , \new_[7250]_ , \new_[7251]_ ,
    \new_[7252]_ , \new_[7253]_ , \new_[7254]_ , \new_[7255]_ ,
    \new_[7256]_ , \new_[7257]_ , \new_[7258]_ , \new_[7263]_ ,
    \new_[7264]_ , \new_[7265]_ , \new_[7266]_ , \new_[7267]_ ,
    \new_[7268]_ , \new_[7269]_ , \new_[7275]_ , \new_[7276]_ ,
    \new_[7277]_ , \new_[7278]_ , \new_[7279]_ , \new_[7280]_ ,
    \new_[7281]_ , \new_[7282]_ , \new_[7283]_ , \new_[7284]_ ,
    \new_[7285]_ , \new_[7286]_ , \new_[7287]_ , \new_[7288]_ ,
    \new_[7289]_ , \new_[7290]_ , \new_[7291]_ , \new_[7292]_ ,
    \new_[7293]_ , \new_[7294]_ , \new_[7295]_ , \new_[7296]_ ,
    \new_[7297]_ , \new_[7298]_ , \new_[7299]_ , \new_[7301]_ ,
    \new_[7302]_ , \new_[7303]_ , \new_[7304]_ , \new_[7305]_ ,
    \new_[7306]_ , \new_[7307]_ , \new_[7308]_ , \new_[7309]_ ,
    \new_[7310]_ , \new_[7311]_ , \new_[7313]_ , \new_[7314]_ ,
    \new_[7315]_ , \new_[7316]_ , \new_[7317]_ , \new_[7318]_ ,
    \new_[7319]_ , \new_[7320]_ , \new_[7321]_ , \new_[7322]_ ,
    \new_[7323]_ , \new_[7344]_ , \new_[7345]_ , \new_[7346]_ ,
    \new_[7347]_ , \new_[7348]_ , \new_[7350]_ , \new_[7352]_ ,
    \new_[7353]_ , \new_[7354]_ , \new_[7355]_ , \new_[7356]_ ,
    \new_[7357]_ , \new_[7358]_ , \new_[7359]_ , \new_[7361]_ ,
    \new_[7365]_ , \new_[7366]_ , \new_[7367]_ , \new_[7368]_ ,
    \new_[7369]_ , \new_[7370]_ , \new_[7379]_ , \new_[7386]_ ,
    \new_[7388]_ , \new_[7389]_ , \new_[7390]_ , \new_[7391]_ ,
    \new_[7394]_ , \new_[7396]_ , \new_[7397]_ , \new_[7398]_ ,
    \new_[7400]_ , \new_[7401]_ , \new_[7402]_ , \new_[7403]_ ,
    \new_[7404]_ , \new_[7405]_ , \new_[7406]_ , \new_[7408]_ ,
    \new_[7409]_ , \new_[7410]_ , \new_[7411]_ , \new_[7412]_ ,
    \new_[7413]_ , \new_[7414]_ , \new_[7415]_ , \new_[7416]_ ,
    \new_[7417]_ , \new_[7418]_ , \new_[7419]_ , \new_[7420]_ ,
    \new_[7423]_ , \new_[7424]_ , \new_[7425]_ , \new_[7426]_ ,
    \new_[7427]_ , \new_[7428]_ , \new_[7429]_ , \new_[7430]_ ,
    \new_[7431]_ , \new_[7432]_ , \new_[7433]_ , \new_[7434]_ ,
    \new_[7435]_ , \new_[7436]_ , \new_[7437]_ , \new_[7438]_ ,
    \new_[7439]_ , \new_[7440]_ , \new_[7441]_ , \new_[7442]_ ,
    \new_[7443]_ , \new_[7444]_ , \new_[7445]_ , \new_[7446]_ ,
    \new_[7447]_ , \new_[7448]_ , \new_[7449]_ , \new_[7450]_ ,
    \new_[7452]_ , \new_[7453]_ , \new_[7454]_ , \new_[7455]_ ,
    \new_[7456]_ , \new_[7458]_ , \new_[7460]_ , \new_[7462]_ ,
    \new_[7464]_ , \new_[7465]_ , \new_[7466]_ , \new_[7467]_ ,
    \new_[7468]_ , \new_[7469]_ , \new_[7470]_ , \new_[7471]_ ,
    \new_[7472]_ , \new_[7473]_ , \new_[7474]_ , \new_[7475]_ ,
    \new_[7476]_ , \new_[7477]_ , \new_[7478]_ , \new_[7479]_ ,
    \new_[7480]_ , \new_[7481]_ , \new_[7482]_ , \new_[7483]_ ,
    \new_[7484]_ , \new_[7485]_ , \new_[7486]_ , \new_[7487]_ ,
    \new_[7488]_ , \new_[7489]_ , \new_[7490]_ , \new_[7491]_ ,
    \new_[7492]_ , \new_[7493]_ , \new_[7494]_ , \new_[7495]_ ,
    \new_[7496]_ , \new_[7497]_ , \new_[7498]_ , \new_[7499]_ ,
    \new_[7500]_ , \new_[7501]_ , \new_[7502]_ , \new_[7503]_ ,
    \new_[7504]_ , \new_[7505]_ , \new_[7506]_ , \new_[7507]_ ,
    \new_[7508]_ , \new_[7509]_ , \new_[7510]_ , \new_[7511]_ ,
    \new_[7512]_ , \new_[7513]_ , \new_[7514]_ , \new_[7515]_ ,
    \new_[7516]_ , \new_[7517]_ , \new_[7518]_ , \new_[7519]_ ,
    \new_[7520]_ , \new_[7521]_ , \new_[7522]_ , \new_[7523]_ ,
    \new_[7524]_ , \new_[7525]_ , \new_[7526]_ , \new_[7527]_ ,
    \new_[7528]_ , \new_[7529]_ , \new_[7538]_ , \new_[7540]_ ,
    \new_[7541]_ , \new_[7542]_ , \new_[7544]_ , \new_[7545]_ ,
    \new_[7546]_ , \new_[7548]_ , \new_[7549]_ , \new_[7550]_ ,
    \new_[7551]_ , \new_[7552]_ , \new_[7553]_ , \new_[7554]_ ,
    \new_[7555]_ , \new_[7556]_ , \new_[7557]_ , \new_[7558]_ ,
    \new_[7559]_ , \new_[7560]_ , \new_[7561]_ , \new_[7562]_ ,
    \new_[7563]_ , \new_[7564]_ , \new_[7565]_ , \new_[7566]_ ,
    \new_[7567]_ , \new_[7568]_ , \new_[7569]_ , \new_[7570]_ ,
    \new_[7572]_ , \new_[7573]_ , \new_[7574]_ , \new_[7575]_ ,
    \new_[7576]_ , \new_[7577]_ , \new_[7578]_ , \new_[7579]_ ,
    \new_[7580]_ , \new_[7581]_ , \new_[7582]_ , \new_[7583]_ ,
    \new_[7584]_ , \new_[7585]_ , \new_[7586]_ , \new_[7587]_ ,
    \new_[7588]_ , \new_[7589]_ , \new_[7590]_ , \new_[7591]_ ,
    \new_[7592]_ , \new_[7593]_ , \new_[7594]_ , \new_[7595]_ ,
    \new_[7596]_ , \new_[7599]_ , \new_[7600]_ , \new_[7601]_ ,
    \new_[7602]_ , \new_[7603]_ , \new_[7604]_ , \new_[7605]_ ,
    \new_[7606]_ , \new_[7619]_ , \new_[7620]_ , \new_[7621]_ ,
    \new_[7622]_ , \new_[7623]_ , \new_[7636]_ , \new_[7637]_ ,
    \new_[7638]_ , \new_[7639]_ , \new_[7640]_ , \new_[7653]_ ,
    \new_[7654]_ , \new_[7655]_ , \new_[7656]_ , \new_[7669]_ ,
    \new_[7670]_ , \new_[7671]_ , \new_[7672]_ , \new_[7673]_ ,
    \new_[7674]_ , \new_[7675]_ , \new_[7676]_ , \new_[7677]_ ,
    \new_[7678]_ , \new_[7680]_ , \new_[7684]_ , \new_[7685]_ ,
    \new_[7686]_ , \new_[7687]_ , \new_[7688]_ , \new_[7689]_ ,
    \new_[7690]_ , \new_[7691]_ , \new_[7692]_ , \new_[7693]_ ,
    \new_[7694]_ , \new_[7695]_ , \new_[7696]_ , \new_[7698]_ ,
    \new_[7699]_ , \new_[7700]_ , \new_[7701]_ , \new_[7702]_ ,
    \new_[7703]_ , \new_[7704]_ , \new_[7705]_ , \new_[7706]_ ,
    \new_[7710]_ , \new_[7712]_ , \new_[7714]_ , \new_[7715]_ ,
    \new_[7716]_ , \new_[7717]_ , \new_[7718]_ , \new_[7719]_ ,
    \new_[7720]_ , \new_[7722]_ , \new_[7723]_ , \new_[7724]_ ,
    \new_[7725]_ , \new_[7726]_ , \new_[7727]_ , \new_[7728]_ ,
    \new_[7729]_ , \new_[7730]_ , \new_[7731]_ , \new_[7732]_ ,
    \new_[7733]_ , \new_[7734]_ , \new_[7735]_ , \new_[7736]_ ,
    \new_[7737]_ , \new_[7738]_ , \new_[7739]_ , \new_[7740]_ ,
    \new_[7741]_ , \new_[7742]_ , \new_[7743]_ , \new_[7744]_ ,
    \new_[7745]_ , \new_[7746]_ , \new_[7747]_ , \new_[7750]_ ,
    \new_[7752]_ , \new_[7753]_ , \new_[7754]_ , \new_[7755]_ ,
    \new_[7756]_ , \new_[7757]_ , \new_[7758]_ , \new_[7759]_ ,
    \new_[7760]_ , \new_[7761]_ , \new_[7762]_ , \new_[7763]_ ,
    \new_[7764]_ , \new_[7765]_ , \new_[7766]_ , \new_[7768]_ ,
    \new_[7769]_ , \new_[7770]_ , \new_[7771]_ , \new_[7772]_ ,
    \new_[7773]_ , \new_[7774]_ , \new_[7775]_ , \new_[7776]_ ,
    \new_[7777]_ , \new_[7778]_ , \new_[7779]_ , \new_[7780]_ ,
    \new_[7781]_ , \new_[7782]_ , \new_[7783]_ , \new_[7785]_ ,
    \new_[7786]_ , \new_[7787]_ , \new_[7788]_ , \new_[7789]_ ,
    \new_[7790]_ , \new_[7791]_ , \new_[7792]_ , \new_[7793]_ ,
    \new_[7794]_ , \new_[7795]_ , \new_[7796]_ , \new_[7797]_ ,
    \new_[7798]_ , \new_[7799]_ , \new_[7800]_ , \new_[7801]_ ,
    \new_[7802]_ , \new_[7803]_ , \new_[7804]_ , \new_[7805]_ ,
    \new_[7806]_ , \new_[7807]_ , \new_[7808]_ , \new_[7809]_ ,
    \new_[7810]_ , \new_[7811]_ , \new_[7812]_ , \new_[7813]_ ,
    \new_[7814]_ , \new_[7815]_ , \new_[7816]_ , \new_[7817]_ ,
    \new_[7818]_ , \new_[7819]_ , \new_[7820]_ , \new_[7821]_ ,
    \new_[7822]_ , \new_[7823]_ , \new_[7824]_ , \new_[7825]_ ,
    \new_[7826]_ , \new_[7827]_ , \new_[7828]_ , \new_[7829]_ ,
    \new_[7830]_ , \new_[7831]_ , \new_[7832]_ , \new_[7833]_ ,
    \new_[7834]_ , \new_[7835]_ , \new_[7836]_ , \new_[7837]_ ,
    \new_[7838]_ , \new_[7839]_ , \new_[7840]_ , \new_[7841]_ ,
    \new_[7842]_ , \new_[7843]_ , \new_[7844]_ , \new_[7845]_ ,
    \new_[7846]_ , \new_[7847]_ , \new_[7848]_ , \new_[7849]_ ,
    \new_[7850]_ , \new_[7851]_ , \new_[7852]_ , \new_[7853]_ ,
    \new_[7854]_ , \new_[7855]_ , \new_[7856]_ , \new_[7857]_ ,
    \new_[7858]_ , \new_[7859]_ , \new_[7860]_ , \new_[7861]_ ,
    \new_[7862]_ , \new_[7863]_ , \new_[7864]_ , \new_[7865]_ ,
    \new_[7866]_ , \new_[7867]_ , \new_[7868]_ , \new_[7869]_ ,
    \new_[7870]_ , \new_[7871]_ , \new_[7872]_ , \new_[7873]_ ,
    \new_[7874]_ , \new_[7875]_ , \new_[7876]_ , \new_[7877]_ ,
    \new_[7878]_ , \new_[7879]_ , \new_[7880]_ , \new_[7881]_ ,
    \new_[7882]_ , \new_[7883]_ , \new_[7884]_ , \new_[7885]_ ,
    \new_[7886]_ , \new_[7887]_ , \new_[7888]_ , \new_[7889]_ ,
    \new_[7890]_ , \new_[7891]_ , \new_[7892]_ , \new_[7893]_ ,
    \new_[7894]_ , \new_[7895]_ , \new_[7896]_ , \new_[7897]_ ,
    \new_[7898]_ , \new_[7899]_ , \new_[7900]_ , \new_[7901]_ ,
    \new_[7902]_ , \new_[7903]_ , \new_[7904]_ , \new_[7905]_ ,
    \new_[7906]_ , \new_[7907]_ , \new_[7908]_ , \new_[7909]_ ,
    \new_[7910]_ , \new_[7911]_ , \new_[7912]_ , \new_[7913]_ ,
    \new_[7914]_ , \new_[7915]_ , \new_[7916]_ , \new_[7917]_ ,
    \new_[7918]_ , \new_[7919]_ , \new_[7920]_ , \new_[7921]_ ,
    \new_[7922]_ , \new_[7923]_ , \new_[7924]_ , \new_[7925]_ ,
    \new_[7926]_ , \new_[7927]_ , \new_[7928]_ , \new_[7929]_ ,
    \new_[7930]_ , \new_[7931]_ , \new_[7932]_ , \new_[7933]_ ,
    \new_[7934]_ , \new_[7935]_ , \new_[7936]_ , \new_[7937]_ ,
    \new_[7938]_ , \new_[7939]_ , \new_[7940]_ , \new_[7941]_ ,
    \new_[7942]_ , \new_[7943]_ , \new_[7944]_ , \new_[7945]_ ,
    \new_[7946]_ , \new_[7947]_ , \new_[7948]_ , \new_[7949]_ ,
    \new_[7950]_ , \new_[7951]_ , \new_[7952]_ , \new_[7953]_ ,
    \new_[7954]_ , \new_[7955]_ , \new_[7956]_ , \new_[7957]_ ,
    \new_[7958]_ , \new_[7959]_ , \new_[7960]_ , \new_[7961]_ ,
    \new_[7962]_ , \new_[7963]_ , \new_[7964]_ , \new_[7965]_ ,
    \new_[7966]_ , \new_[7967]_ , \new_[7968]_ , \new_[7969]_ ,
    \new_[7970]_ , \new_[7971]_ , \new_[7972]_ , \new_[7973]_ ,
    \new_[7974]_ , \new_[7975]_ , \new_[7976]_ , \new_[7977]_ ,
    \new_[7978]_ , \new_[7979]_ , \new_[7980]_ , \new_[7981]_ ,
    \new_[7982]_ , \new_[7983]_ , \new_[7984]_ , \new_[7985]_ ,
    \new_[7986]_ , \new_[7987]_ , \new_[7988]_ , \new_[7989]_ ,
    \new_[7990]_ , \new_[7991]_ , \new_[7992]_ , \new_[7993]_ ,
    \new_[7994]_ , \new_[7995]_ , \new_[7996]_ , \new_[7997]_ ,
    \new_[7998]_ , \new_[7999]_ , \new_[8000]_ , \new_[8001]_ ,
    \new_[8002]_ , \new_[8003]_ , \new_[8004]_ , \new_[8005]_ ,
    \new_[8006]_ , \new_[8007]_ , \new_[8008]_ , \new_[8009]_ ,
    \new_[8010]_ , \new_[8011]_ , \new_[8012]_ , \new_[8013]_ ,
    \new_[8014]_ , \new_[8015]_ , \new_[8016]_ , \new_[8017]_ ,
    \new_[8018]_ , \new_[8019]_ , \new_[8020]_ , \new_[8021]_ ,
    \new_[8022]_ , \new_[8023]_ , \new_[8024]_ , \new_[8025]_ ,
    \new_[8026]_ , \new_[8027]_ , \new_[8028]_ , \new_[8029]_ ,
    \new_[8030]_ , \new_[8031]_ , \new_[8032]_ , \new_[8033]_ ,
    \new_[8034]_ , \new_[8035]_ , \new_[8036]_ , \new_[8037]_ ,
    \new_[8038]_ , \new_[8039]_ , \new_[8040]_ , \new_[8041]_ ,
    \new_[8042]_ , \new_[8043]_ , \new_[8044]_ , \new_[8045]_ ,
    \new_[8046]_ , \new_[8047]_ , \new_[8048]_ , \new_[8049]_ ,
    \new_[8050]_ , \new_[8051]_ , \new_[8052]_ , \new_[8053]_ ,
    \new_[8054]_ , \new_[8055]_ , \new_[8056]_ , \new_[8057]_ ,
    \new_[8058]_ , \new_[8059]_ , \new_[8060]_ , \new_[8061]_ ,
    \new_[8062]_ , \new_[8063]_ , \new_[8064]_ , \new_[8065]_ ,
    \new_[8066]_ , \new_[8067]_ , \new_[8068]_ , \new_[8069]_ ,
    \new_[8070]_ , \new_[8071]_ , \new_[8072]_ , \new_[8073]_ ,
    \new_[8074]_ , \new_[8075]_ , \new_[8076]_ , \new_[8077]_ ,
    \new_[8078]_ , \new_[8079]_ , \new_[8080]_ , \new_[8081]_ ,
    \new_[8082]_ , \new_[8083]_ , \new_[8084]_ , \new_[8085]_ ,
    \new_[8086]_ , \new_[8087]_ , \new_[8088]_ , \new_[8089]_ ,
    \new_[8090]_ , \new_[8091]_ , \new_[8092]_ , \new_[8093]_ ,
    \new_[8094]_ , \new_[8095]_ , \new_[8096]_ , \new_[8097]_ ,
    \new_[8098]_ , \new_[8099]_ , \new_[8100]_ , \new_[8101]_ ,
    \new_[8102]_ , \new_[8103]_ , \new_[8104]_ , \new_[8105]_ ,
    \new_[8106]_ , \new_[8107]_ , \new_[8108]_ , \new_[8109]_ ,
    \new_[8110]_ , \new_[8111]_ , \new_[8112]_ , \new_[8113]_ ,
    \new_[8114]_ , \new_[8115]_ , \new_[8116]_ , \new_[8117]_ ,
    \new_[8118]_ , \new_[8119]_ , \new_[8120]_ , \new_[8121]_ ,
    \new_[8122]_ , \new_[8123]_ , \new_[8124]_ , \new_[8125]_ ,
    \new_[8126]_ , \new_[8127]_ , \new_[8128]_ , \new_[8129]_ ,
    \new_[8130]_ , \new_[8131]_ , \new_[8132]_ , \new_[8133]_ ,
    \new_[8134]_ , \new_[8135]_ , \new_[8136]_ , \new_[8137]_ ,
    \new_[8138]_ , \new_[8139]_ , \new_[8140]_ , \new_[8141]_ ,
    \new_[8142]_ , \new_[8143]_ , \new_[8144]_ , \new_[8145]_ ,
    \new_[8146]_ , \new_[8147]_ , \new_[8148]_ , \new_[8149]_ ,
    \new_[8150]_ , \new_[8151]_ , \new_[8152]_ , \new_[8153]_ ,
    \new_[8154]_ , \new_[8155]_ , \new_[8156]_ , \new_[8157]_ ,
    \new_[8158]_ , \new_[8159]_ , \new_[8160]_ , \new_[8161]_ ,
    \new_[8162]_ , \new_[8163]_ , \new_[8164]_ , \new_[8165]_ ,
    \new_[8166]_ , \new_[8167]_ , \new_[8168]_ , \new_[8169]_ ,
    \new_[8170]_ , \new_[8171]_ , \new_[8172]_ , \new_[8173]_ ,
    \new_[8174]_ , \new_[8175]_ , \new_[8176]_ , \new_[8177]_ ,
    \new_[8178]_ , \new_[8179]_ , \new_[8180]_ , \new_[8181]_ ,
    \new_[8182]_ , \new_[8183]_ , \new_[8184]_ , \new_[8185]_ ,
    \new_[8186]_ , \new_[8187]_ , \new_[8188]_ , \new_[8189]_ ,
    \new_[8190]_ , \new_[8191]_ , \new_[8192]_ , \new_[8193]_ ,
    \new_[8194]_ , \new_[8195]_ , \new_[8196]_ , \new_[8197]_ ,
    \new_[8198]_ , \new_[8199]_ , \new_[8200]_ , \new_[8201]_ ,
    \new_[8202]_ , \new_[8203]_ , \new_[8204]_ , \new_[8205]_ ,
    \new_[8206]_ , \new_[8207]_ , \new_[8208]_ , \new_[8209]_ ,
    \new_[8210]_ , \new_[8211]_ , \new_[8214]_ , \new_[8215]_ ,
    \new_[8216]_ , \new_[8217]_ , \new_[8218]_ , \new_[8219]_ ,
    \new_[8220]_ , \new_[8221]_ , \new_[8222]_ , \new_[8223]_ ,
    \new_[8224]_ , \new_[8225]_ , \new_[8226]_ , \new_[8229]_ ,
    \new_[8230]_ , \new_[8231]_ , \new_[8232]_ , \new_[8233]_ ,
    \new_[8234]_ , \new_[8235]_ , \new_[8236]_ , \new_[8237]_ ,
    \new_[8238]_ , \new_[8239]_ , \new_[8240]_ , \new_[8241]_ ,
    \new_[8242]_ , \new_[8243]_ , \new_[8244]_ , \new_[8245]_ ,
    \new_[8246]_ , \new_[8247]_ , \new_[8248]_ , \new_[8249]_ ,
    \new_[8250]_ , \new_[8251]_ , \new_[8252]_ , \new_[8253]_ ,
    \new_[8254]_ , \new_[8255]_ , \new_[8257]_ , \new_[8258]_ ,
    \new_[8259]_ , \new_[8260]_ , \new_[8261]_ , \new_[8262]_ ,
    \new_[8263]_ , \new_[8264]_ , \new_[8265]_ , \new_[8266]_ ,
    \new_[8267]_ , \new_[8268]_ , \new_[8269]_ , \new_[8270]_ ,
    \new_[8271]_ , \new_[8272]_ , \new_[8273]_ , \new_[8274]_ ,
    \new_[8275]_ , \new_[8276]_ , \new_[8277]_ , \new_[8278]_ ,
    \new_[8279]_ , \new_[8280]_ , \new_[8281]_ , \new_[8282]_ ,
    \new_[8283]_ , \new_[8284]_ , \new_[8285]_ , \new_[8286]_ ,
    \new_[8287]_ , \new_[8288]_ , \new_[8289]_ , \new_[8290]_ ,
    \new_[8291]_ , \new_[8292]_ , \new_[8293]_ , \new_[8294]_ ,
    \new_[8295]_ , \new_[8296]_ , \new_[8297]_ , \new_[8298]_ ,
    \new_[8299]_ , \new_[8300]_ , \new_[8301]_ , \new_[8303]_ ,
    \new_[8304]_ , \new_[8305]_ , \new_[8306]_ , \new_[8307]_ ,
    \new_[8308]_ , \new_[8309]_ , \new_[8310]_ , \new_[8311]_ ,
    \new_[8312]_ , \new_[8313]_ , \new_[8314]_ , \new_[8319]_ ,
    \new_[8321]_ , \new_[8322]_ , \new_[8323]_ , \new_[8325]_ ,
    \new_[8326]_ , \new_[8327]_ , \new_[8328]_ , \new_[8329]_ ,
    \new_[8330]_ , \new_[8331]_ , \new_[8332]_ , \new_[8333]_ ,
    \new_[8334]_ , \new_[8335]_ , \new_[8336]_ , \new_[8337]_ ,
    \new_[8338]_ , \new_[8339]_ , \new_[8340]_ , \new_[8341]_ ,
    \new_[8342]_ , \new_[8343]_ , \new_[8344]_ , \new_[8345]_ ,
    \new_[8346]_ , \new_[8347]_ , \new_[8348]_ , \new_[8349]_ ,
    \new_[8350]_ , \new_[8351]_ , \new_[8352]_ , \new_[8353]_ ,
    \new_[8354]_ , \new_[8355]_ , \new_[8356]_ , \new_[8357]_ ,
    \new_[8358]_ , \new_[8359]_ , \new_[8360]_ , \new_[8361]_ ,
    \new_[8362]_ , \new_[8363]_ , \new_[8364]_ , \new_[8365]_ ,
    \new_[8366]_ , \new_[8367]_ , \new_[8368]_ , \new_[8369]_ ,
    \new_[8370]_ , \new_[8371]_ , \new_[8372]_ , \new_[8373]_ ,
    \new_[8374]_ , \new_[8375]_ , \new_[8376]_ , \new_[8377]_ ,
    \new_[8378]_ , \new_[8379]_ , \new_[8380]_ , \new_[8381]_ ,
    \new_[8382]_ , \new_[8383]_ , \new_[8384]_ , \new_[8385]_ ,
    \new_[8386]_ , \new_[8387]_ , \new_[8388]_ , \new_[8389]_ ,
    \new_[8390]_ , \new_[8391]_ , \new_[8392]_ , \new_[8393]_ ,
    \new_[8394]_ , \new_[8395]_ , \new_[8396]_ , \new_[8397]_ ,
    \new_[8398]_ , \new_[8399]_ , \new_[8400]_ , \new_[8401]_ ,
    \new_[8402]_ , \new_[8403]_ , \new_[8404]_ , \new_[8405]_ ,
    \new_[8406]_ , \new_[8407]_ , \new_[8408]_ , \new_[8409]_ ,
    \new_[8410]_ , \new_[8411]_ , \new_[8412]_ , \new_[8413]_ ,
    \new_[8414]_ , \new_[8415]_ , \new_[8416]_ , \new_[8417]_ ,
    \new_[8418]_ , \new_[8419]_ , \new_[8420]_ , \new_[8421]_ ,
    \new_[8422]_ , \new_[8423]_ , \new_[8424]_ , \new_[8425]_ ,
    \new_[8426]_ , \new_[8427]_ , \new_[8428]_ , \new_[8429]_ ,
    \new_[8430]_ , \new_[8431]_ , \new_[8432]_ , \new_[8433]_ ,
    \new_[8434]_ , \new_[8435]_ , \new_[8436]_ , \new_[8437]_ ,
    \new_[8438]_ , \new_[8439]_ , \new_[8440]_ , \new_[8441]_ ,
    \new_[8442]_ , \new_[8443]_ , \new_[8444]_ , \new_[8445]_ ,
    \new_[8446]_ , \new_[8447]_ , \new_[8448]_ , \new_[8449]_ ,
    \new_[8450]_ , \new_[8451]_ , \new_[8452]_ , \new_[8453]_ ,
    \new_[8454]_ , \new_[8455]_ , \new_[8456]_ , \new_[8457]_ ,
    \new_[8458]_ , \new_[8459]_ , \new_[8460]_ , \new_[8461]_ ,
    \new_[8462]_ , \new_[8463]_ , \new_[8464]_ , \new_[8465]_ ,
    \new_[8466]_ , \new_[8467]_ , \new_[8468]_ , \new_[8469]_ ,
    \new_[8470]_ , \new_[8471]_ , \new_[8472]_ , \new_[8473]_ ,
    \new_[8474]_ , \new_[8475]_ , \new_[8476]_ , \new_[8477]_ ,
    \new_[8478]_ , \new_[8479]_ , \new_[8480]_ , \new_[8481]_ ,
    \new_[8482]_ , \new_[8483]_ , \new_[8484]_ , \new_[8485]_ ,
    \new_[8486]_ , \new_[8487]_ , \new_[8488]_ , \new_[8489]_ ,
    \new_[8490]_ , \new_[8491]_ , \new_[8492]_ , \new_[8493]_ ,
    \new_[8494]_ , \new_[8495]_ , \new_[8496]_ , \new_[8497]_ ,
    \new_[8498]_ , \new_[8499]_ , \new_[8500]_ , \new_[8501]_ ,
    \new_[8502]_ , \new_[8503]_ , \new_[8504]_ , \new_[8505]_ ,
    \new_[8507]_ , \new_[8508]_ , \new_[8509]_ , \new_[8510]_ ,
    \new_[8511]_ , \new_[8512]_ , \new_[8513]_ , \new_[8514]_ ,
    \new_[8515]_ , \new_[8516]_ , \new_[8517]_ , \new_[8518]_ ,
    \new_[8519]_ , \new_[8520]_ , \new_[8521]_ , \new_[8522]_ ,
    \new_[8523]_ , \new_[8524]_ , \new_[8525]_ , \new_[8526]_ ,
    \new_[8527]_ , \new_[8528]_ , \new_[8529]_ , \new_[8530]_ ,
    \new_[8531]_ , \new_[8532]_ , \new_[8533]_ , \new_[8534]_ ,
    \new_[8535]_ , \new_[8536]_ , \new_[8537]_ , \new_[8538]_ ,
    \new_[8539]_ , \new_[8540]_ , \new_[8541]_ , \new_[8542]_ ,
    \new_[8543]_ , \new_[8544]_ , \new_[8545]_ , \new_[8546]_ ,
    \new_[8547]_ , \new_[8548]_ , \new_[8549]_ , \new_[8550]_ ,
    \new_[8552]_ , \new_[8553]_ , \new_[8554]_ , \new_[8555]_ ,
    \new_[8556]_ , \new_[8557]_ , \new_[8558]_ , \new_[8559]_ ,
    \new_[8560]_ , \new_[8562]_ , \new_[8563]_ , \new_[8564]_ ,
    \new_[8565]_ , \new_[8566]_ , \new_[8567]_ , \new_[8568]_ ,
    \new_[8569]_ , \new_[8570]_ , \new_[8571]_ , \new_[8572]_ ,
    \new_[8573]_ , \new_[8574]_ , \new_[8575]_ , \new_[8576]_ ,
    \new_[8577]_ , \new_[8578]_ , \new_[8579]_ , \new_[8580]_ ,
    \new_[8581]_ , \new_[8582]_ , \new_[8583]_ , \new_[8584]_ ,
    \new_[8585]_ , \new_[8586]_ , \new_[8587]_ , \new_[8588]_ ,
    \new_[8589]_ , \new_[8590]_ , \new_[8591]_ , \new_[8592]_ ,
    \new_[8593]_ , \new_[8594]_ , \new_[8595]_ , \new_[8596]_ ,
    \new_[8597]_ , \new_[8598]_ , \new_[8599]_ , \new_[8600]_ ,
    \new_[8601]_ , \new_[8602]_ , \new_[8603]_ , \new_[8604]_ ,
    \new_[8605]_ , \new_[8606]_ , \new_[8607]_ , \new_[8608]_ ,
    \new_[8609]_ , \new_[8610]_ , \new_[8611]_ , \new_[8612]_ ,
    \new_[8613]_ , \new_[8614]_ , \new_[8615]_ , \new_[8616]_ ,
    \new_[8618]_ , \new_[8619]_ , \new_[8620]_ , \new_[8621]_ ,
    \new_[8622]_ , \new_[8623]_ , \new_[8624]_ , \new_[8625]_ ,
    \new_[8626]_ , \new_[8627]_ , \new_[8628]_ , \new_[8629]_ ,
    \new_[8630]_ , \new_[8631]_ , \new_[8632]_ , \new_[8633]_ ,
    \new_[8634]_ , \new_[8635]_ , \new_[8636]_ , \new_[8637]_ ,
    \new_[8638]_ , \new_[8639]_ , \new_[8640]_ , \new_[8641]_ ,
    \new_[8642]_ , \new_[8643]_ , \new_[8644]_ , \new_[8645]_ ,
    \new_[8646]_ , \new_[8647]_ , \new_[8648]_ , \new_[8649]_ ,
    \new_[8650]_ , \new_[8651]_ , \new_[8652]_ , \new_[8653]_ ,
    \new_[8654]_ , \new_[8655]_ , \new_[8656]_ , \new_[8657]_ ,
    \new_[8658]_ , \new_[8659]_ , \new_[8660]_ , \new_[8661]_ ,
    \new_[8662]_ , \new_[8663]_ , \new_[8664]_ , \new_[8665]_ ,
    \new_[8666]_ , \new_[8667]_ , \new_[8668]_ , \new_[8671]_ ,
    \new_[8672]_ , \new_[8675]_ , \new_[8676]_ , \new_[8677]_ ,
    \new_[8678]_ , \new_[8679]_ , \new_[8680]_ , \new_[8681]_ ,
    \new_[8682]_ , \new_[8683]_ , \new_[8684]_ , \new_[8685]_ ,
    \new_[8686]_ , \new_[8687]_ , \new_[8688]_ , \new_[8689]_ ,
    \new_[8690]_ , \new_[8691]_ , \new_[8692]_ , \new_[8693]_ ,
    \new_[8694]_ , \new_[8695]_ , \new_[8696]_ , \new_[8697]_ ,
    \new_[8698]_ , \new_[8699]_ , \new_[8700]_ , \new_[8701]_ ,
    \new_[8702]_ , \new_[8703]_ , \new_[8705]_ , \new_[8706]_ ,
    \new_[8707]_ , \new_[8709]_ , \new_[8710]_ , \new_[8711]_ ,
    \new_[8712]_ , \new_[8714]_ , \new_[8715]_ , \new_[8716]_ ,
    \new_[8717]_ , \new_[8718]_ , \new_[8719]_ , \new_[8720]_ ,
    \new_[8721]_ , \new_[8722]_ , \new_[8723]_ , \new_[8724]_ ,
    \new_[8725]_ , \new_[8726]_ , \new_[8727]_ , \new_[8728]_ ,
    \new_[8729]_ , \new_[8730]_ , \new_[8731]_ , \new_[8732]_ ,
    \new_[8733]_ , \new_[8734]_ , \new_[8735]_ , \new_[8736]_ ,
    \new_[8737]_ , \new_[8738]_ , \new_[8739]_ , \new_[8740]_ ,
    \new_[8741]_ , \new_[8742]_ , \new_[8743]_ , \new_[8744]_ ,
    \new_[8745]_ , \new_[8746]_ , \new_[8747]_ , \new_[8748]_ ,
    \new_[8749]_ , \new_[8750]_ , \new_[8751]_ , \new_[8752]_ ,
    \new_[8753]_ , \new_[8754]_ , \new_[8755]_ , \new_[8756]_ ,
    \new_[8757]_ , \new_[8758]_ , \new_[8759]_ , \new_[8760]_ ,
    \new_[8761]_ , \new_[8762]_ , \new_[8763]_ , \new_[8764]_ ,
    \new_[8765]_ , \new_[8766]_ , \new_[8767]_ , \new_[8768]_ ,
    \new_[8769]_ , \new_[8770]_ , \new_[8771]_ , \new_[8772]_ ,
    \new_[8773]_ , \new_[8774]_ , \new_[8775]_ , \new_[8776]_ ,
    \new_[8777]_ , \new_[8778]_ , \new_[8779]_ , \new_[8780]_ ,
    \new_[8781]_ , \new_[8782]_ , \new_[8783]_ , \new_[8784]_ ,
    \new_[8785]_ , \new_[8786]_ , \new_[8787]_ , \new_[8788]_ ,
    \new_[8789]_ , \new_[8790]_ , \new_[8791]_ , \new_[8792]_ ,
    \new_[8793]_ , \new_[8794]_ , \new_[8795]_ , \new_[8796]_ ,
    \new_[8797]_ , \new_[8798]_ , \new_[8799]_ , \new_[8800]_ ,
    \new_[8801]_ , \new_[8802]_ , \new_[8803]_ , \new_[8804]_ ,
    \new_[8805]_ , \new_[8806]_ , \new_[8807]_ , \new_[8808]_ ,
    \new_[8809]_ , \new_[8810]_ , \new_[8811]_ , \new_[8812]_ ,
    \new_[8813]_ , \new_[8814]_ , \new_[8815]_ , \new_[8816]_ ,
    \new_[8817]_ , \new_[8818]_ , \new_[8819]_ , \new_[8820]_ ,
    \new_[8821]_ , \new_[8822]_ , \new_[8823]_ , \new_[8824]_ ,
    \new_[8825]_ , \new_[8826]_ , \new_[8827]_ , \new_[8828]_ ,
    \new_[8829]_ , \new_[8830]_ , \new_[8831]_ , \new_[8832]_ ,
    \new_[8833]_ , \new_[8834]_ , \new_[8835]_ , \new_[8836]_ ,
    \new_[8837]_ , \new_[8838]_ , \new_[8839]_ , \new_[8840]_ ,
    \new_[8841]_ , \new_[8843]_ , \new_[8844]_ , \new_[8845]_ ,
    \new_[8846]_ , \new_[8847]_ , \new_[8848]_ , \new_[8849]_ ,
    \new_[8850]_ , \new_[8851]_ , \new_[8852]_ , \new_[8853]_ ,
    \new_[8854]_ , \new_[8855]_ , \new_[8856]_ , \new_[8857]_ ,
    \new_[8858]_ , \new_[8859]_ , \new_[8860]_ , \new_[8861]_ ,
    \new_[8862]_ , \new_[8863]_ , \new_[8864]_ , \new_[8865]_ ,
    \new_[8866]_ , \new_[8867]_ , \new_[8868]_ , \new_[8869]_ ,
    \new_[8870]_ , \new_[8871]_ , \new_[8872]_ , \new_[8873]_ ,
    \new_[8874]_ , \new_[8875]_ , \new_[8876]_ , \new_[8877]_ ,
    \new_[8878]_ , \new_[8879]_ , \new_[8880]_ , \new_[8881]_ ,
    \new_[8882]_ , \new_[8884]_ , \new_[8885]_ , \new_[8886]_ ,
    \new_[8888]_ , \new_[8889]_ , \new_[8890]_ , \new_[8891]_ ,
    \new_[8892]_ , \new_[8893]_ , \new_[8894]_ , \new_[8895]_ ,
    \new_[8896]_ , \new_[8897]_ , \new_[8898]_ , \new_[8899]_ ,
    \new_[8900]_ , \new_[8901]_ , \new_[8903]_ , \new_[8904]_ ,
    \new_[8905]_ , \new_[8906]_ , \new_[8907]_ , \new_[8908]_ ,
    \new_[8909]_ , \new_[8910]_ , \new_[8911]_ , \new_[8912]_ ,
    \new_[8913]_ , \new_[8914]_ , \new_[8915]_ , \new_[8916]_ ,
    \new_[8918]_ , \new_[8919]_ , \new_[8921]_ , \new_[8922]_ ,
    \new_[8923]_ , \new_[8924]_ , \new_[8927]_ , \new_[8928]_ ,
    \new_[8929]_ , \new_[8930]_ , \new_[8931]_ , \new_[8932]_ ,
    \new_[8933]_ , \new_[8934]_ , \new_[8935]_ , \new_[8936]_ ,
    \new_[8937]_ , \new_[8938]_ , \new_[8939]_ , \new_[8940]_ ,
    \new_[8941]_ , \new_[8942]_ , \new_[8943]_ , \new_[8944]_ ,
    \new_[8945]_ , \new_[8946]_ , \new_[8947]_ , \new_[8948]_ ,
    \new_[8949]_ , \new_[8950]_ , \new_[8951]_ , \new_[8952]_ ,
    \new_[8953]_ , \new_[8954]_ , \new_[8955]_ , \new_[8956]_ ,
    \new_[8957]_ , \new_[8958]_ , \new_[8959]_ , \new_[8960]_ ,
    \new_[8961]_ , \new_[8963]_ , \new_[8964]_ , \new_[8965]_ ,
    \new_[8966]_ , \new_[8967]_ , \new_[8968]_ , \new_[8969]_ ,
    \new_[8970]_ , \new_[8971]_ , \new_[8972]_ , \new_[8973]_ ,
    \new_[8974]_ , \new_[8975]_ , \new_[8976]_ , \new_[8977]_ ,
    \new_[8978]_ , \new_[8979]_ , \new_[8980]_ , \new_[8981]_ ,
    \new_[8982]_ , \new_[8983]_ , \new_[8984]_ , \new_[8985]_ ,
    \new_[8986]_ , \new_[8987]_ , \new_[8988]_ , \new_[8989]_ ,
    \new_[8990]_ , \new_[8991]_ , \new_[8992]_ , \new_[8993]_ ,
    \new_[8994]_ , \new_[8995]_ , \new_[8996]_ , \new_[8997]_ ,
    \new_[8998]_ , \new_[8999]_ , \new_[9000]_ , \new_[9001]_ ,
    \new_[9002]_ , \new_[9003]_ , \new_[9004]_ , \new_[9005]_ ,
    \new_[9006]_ , \new_[9007]_ , \new_[9008]_ , \new_[9009]_ ,
    \new_[9010]_ , \new_[9011]_ , \new_[9012]_ , \new_[9013]_ ,
    \new_[9014]_ , \new_[9015]_ , \new_[9016]_ , \new_[9017]_ ,
    \new_[9018]_ , \new_[9019]_ , \new_[9020]_ , \new_[9021]_ ,
    \new_[9022]_ , \new_[9023]_ , \new_[9024]_ , \new_[9025]_ ,
    \new_[9026]_ , \new_[9027]_ , \new_[9028]_ , \new_[9029]_ ,
    \new_[9030]_ , \new_[9031]_ , \new_[9032]_ , \new_[9033]_ ,
    \new_[9034]_ , \new_[9035]_ , \new_[9036]_ , \new_[9037]_ ,
    \new_[9038]_ , \new_[9039]_ , \new_[9040]_ , \new_[9041]_ ,
    \new_[9042]_ , \new_[9043]_ , \new_[9044]_ , \new_[9045]_ ,
    \new_[9046]_ , \new_[9047]_ , \new_[9048]_ , \new_[9049]_ ,
    \new_[9050]_ , \new_[9051]_ , \new_[9052]_ , \new_[9053]_ ,
    \new_[9054]_ , \new_[9055]_ , \new_[9056]_ , \new_[9057]_ ,
    \new_[9059]_ , \new_[9060]_ , \new_[9061]_ , \new_[9062]_ ,
    \new_[9063]_ , \new_[9064]_ , \new_[9065]_ , \new_[9066]_ ,
    \new_[9067]_ , \new_[9068]_ , \new_[9069]_ , \new_[9070]_ ,
    \new_[9071]_ , \new_[9072]_ , \new_[9073]_ , \new_[9074]_ ,
    \new_[9075]_ , \new_[9076]_ , \new_[9077]_ , \new_[9078]_ ,
    \new_[9079]_ , \new_[9080]_ , \new_[9081]_ , \new_[9082]_ ,
    \new_[9083]_ , \new_[9084]_ , \new_[9085]_ , \new_[9086]_ ,
    \new_[9087]_ , \new_[9088]_ , \new_[9089]_ , \new_[9090]_ ,
    \new_[9091]_ , \new_[9092]_ , \new_[9093]_ , \new_[9094]_ ,
    \new_[9095]_ , \new_[9096]_ , \new_[9097]_ , \new_[9099]_ ,
    \new_[9101]_ , \new_[9102]_ , \new_[9103]_ , \new_[9104]_ ,
    \new_[9105]_ , \new_[9106]_ , \new_[9107]_ , \new_[9108]_ ,
    \new_[9109]_ , \new_[9110]_ , \new_[9111]_ , \new_[9112]_ ,
    \new_[9114]_ , \new_[9116]_ , \new_[9119]_ , \new_[9120]_ ,
    \new_[9121]_ , \new_[9122]_ , \new_[9123]_ , \new_[9124]_ ,
    \new_[9125]_ , \new_[9126]_ , \new_[9127]_ , \new_[9128]_ ,
    \new_[9129]_ , \new_[9130]_ , \new_[9131]_ , \new_[9132]_ ,
    \new_[9133]_ , \new_[9134]_ , \new_[9135]_ , \new_[9136]_ ,
    \new_[9137]_ , \new_[9138]_ , \new_[9139]_ , \new_[9140]_ ,
    \new_[9141]_ , \new_[9142]_ , \new_[9143]_ , \new_[9144]_ ,
    \new_[9145]_ , \new_[9146]_ , \new_[9147]_ , \new_[9148]_ ,
    \new_[9149]_ , \new_[9150]_ , \new_[9151]_ , \new_[9152]_ ,
    \new_[9153]_ , \new_[9154]_ , \new_[9155]_ , \new_[9156]_ ,
    \new_[9157]_ , \new_[9158]_ , \new_[9159]_ , \new_[9160]_ ,
    \new_[9161]_ , \new_[9162]_ , \new_[9163]_ , \new_[9164]_ ,
    \new_[9165]_ , \new_[9166]_ , \new_[9167]_ , \new_[9168]_ ,
    \new_[9169]_ , \new_[9170]_ , \new_[9171]_ , \new_[9172]_ ,
    \new_[9173]_ , \new_[9174]_ , \new_[9175]_ , \new_[9178]_ ,
    \new_[9179]_ , \new_[9183]_ , \new_[9184]_ , \new_[9185]_ ,
    \new_[9186]_ , \new_[9187]_ , \new_[9188]_ , \new_[9189]_ ,
    \new_[9190]_ , \new_[9191]_ , \new_[9192]_ , \new_[9193]_ ,
    \new_[9194]_ , \new_[9195]_ , \new_[9196]_ , \new_[9197]_ ,
    \new_[9198]_ , \new_[9199]_ , \new_[9200]_ , \new_[9201]_ ,
    \new_[9202]_ , \new_[9203]_ , \new_[9204]_ , \new_[9205]_ ,
    \new_[9206]_ , \new_[9207]_ , \new_[9208]_ , \new_[9211]_ ,
    \new_[9213]_ , \new_[9214]_ , \new_[9215]_ , \new_[9216]_ ,
    \new_[9217]_ , \new_[9218]_ , \new_[9219]_ , \new_[9220]_ ,
    \new_[9221]_ , \new_[9222]_ , \new_[9223]_ , \new_[9224]_ ,
    \new_[9225]_ , \new_[9226]_ , \new_[9227]_ , \new_[9228]_ ,
    \new_[9229]_ , \new_[9230]_ , \new_[9231]_ , \new_[9232]_ ,
    \new_[9233]_ , \new_[9234]_ , \new_[9235]_ , \new_[9236]_ ,
    \new_[9237]_ , \new_[9238]_ , \new_[9239]_ , \new_[9240]_ ,
    \new_[9241]_ , \new_[9242]_ , \new_[9243]_ , \new_[9244]_ ,
    \new_[9245]_ , \new_[9246]_ , \new_[9247]_ , \new_[9248]_ ,
    \new_[9249]_ , \new_[9250]_ , \new_[9251]_ , \new_[9252]_ ,
    \new_[9253]_ , \new_[9254]_ , \new_[9255]_ , \new_[9256]_ ,
    \new_[9257]_ , \new_[9258]_ , \new_[9259]_ , \new_[9260]_ ,
    \new_[9261]_ , \new_[9262]_ , \new_[9263]_ , \new_[9264]_ ,
    \new_[9265]_ , \new_[9266]_ , \new_[9267]_ , \new_[9268]_ ,
    \new_[9269]_ , \new_[9270]_ , \new_[9271]_ , \new_[9272]_ ,
    \new_[9273]_ , \new_[9274]_ , \new_[9275]_ , \new_[9276]_ ,
    \new_[9277]_ , \new_[9278]_ , \new_[9279]_ , \new_[9280]_ ,
    \new_[9281]_ , \new_[9282]_ , \new_[9283]_ , \new_[9284]_ ,
    \new_[9285]_ , \new_[9286]_ , \new_[9287]_ , \new_[9288]_ ,
    \new_[9289]_ , \new_[9290]_ , \new_[9291]_ , \new_[9292]_ ,
    \new_[9294]_ , \new_[9295]_ , \new_[9296]_ , \new_[9297]_ ,
    \new_[9298]_ , \new_[9299]_ , \new_[9300]_ , \new_[9301]_ ,
    \new_[9302]_ , \new_[9303]_ , \new_[9304]_ , \new_[9305]_ ,
    \new_[9306]_ , \new_[9307]_ , \new_[9308]_ , \new_[9309]_ ,
    \new_[9310]_ , \new_[9311]_ , \new_[9312]_ , \new_[9313]_ ,
    \new_[9314]_ , \new_[9315]_ , \new_[9316]_ , \new_[9317]_ ,
    \new_[9319]_ , \new_[9320]_ , \new_[9321]_ , \new_[9322]_ ,
    \new_[9323]_ , \new_[9324]_ , \new_[9325]_ , \new_[9326]_ ,
    \new_[9327]_ , \new_[9329]_ , \new_[9330]_ , \new_[9331]_ ,
    \new_[9332]_ , \new_[9333]_ , \new_[9334]_ , \new_[9335]_ ,
    \new_[9336]_ , \new_[9337]_ , \new_[9338]_ , \new_[9339]_ ,
    \new_[9340]_ , \new_[9341]_ , \new_[9342]_ , \new_[9343]_ ,
    \new_[9344]_ , \new_[9345]_ , \new_[9346]_ , \new_[9347]_ ,
    \new_[9348]_ , \new_[9349]_ , \new_[9350]_ , \new_[9351]_ ,
    \new_[9352]_ , \new_[9353]_ , \new_[9354]_ , \new_[9356]_ ,
    \new_[9357]_ , \new_[9358]_ , \new_[9359]_ , \new_[9360]_ ,
    \new_[9361]_ , \new_[9363]_ , \new_[9364]_ , \new_[9365]_ ,
    \new_[9366]_ , \new_[9367]_ , \new_[9368]_ , \new_[9369]_ ,
    \new_[9370]_ , \new_[9371]_ , \new_[9372]_ , \new_[9373]_ ,
    \new_[9375]_ , \new_[9376]_ , \new_[9377]_ , \new_[9378]_ ,
    \new_[9379]_ , \new_[9380]_ , \new_[9381]_ , \new_[9382]_ ,
    \new_[9383]_ , \new_[9384]_ , \new_[9385]_ , \new_[9386]_ ,
    \new_[9387]_ , \new_[9388]_ , \new_[9389]_ , \new_[9390]_ ,
    \new_[9391]_ , \new_[9392]_ , \new_[9393]_ , \new_[9394]_ ,
    \new_[9395]_ , \new_[9396]_ , \new_[9397]_ , \new_[9400]_ ,
    \new_[9401]_ , \new_[9402]_ , \new_[9403]_ , \new_[9404]_ ,
    \new_[9405]_ , \new_[9406]_ , \new_[9407]_ , \new_[9408]_ ,
    \new_[9409]_ , \new_[9410]_ , \new_[9411]_ , \new_[9412]_ ,
    \new_[9413]_ , \new_[9414]_ , \new_[9415]_ , \new_[9416]_ ,
    \new_[9417]_ , \new_[9418]_ , \new_[9419]_ , \new_[9420]_ ,
    \new_[9421]_ , \new_[9422]_ , \new_[9424]_ , \new_[9425]_ ,
    \new_[9426]_ , \new_[9427]_ , \new_[9428]_ , \new_[9429]_ ,
    \new_[9430]_ , \new_[9431]_ , \new_[9432]_ , \new_[9433]_ ,
    \new_[9434]_ , \new_[9436]_ , \new_[9437]_ , \new_[9440]_ ,
    \new_[9441]_ , \new_[9442]_ , \new_[9443]_ , \new_[9444]_ ,
    \new_[9445]_ , \new_[9446]_ , \new_[9447]_ , \new_[9448]_ ,
    \new_[9449]_ , \new_[9450]_ , \new_[9451]_ , \new_[9452]_ ,
    \new_[9453]_ , \new_[9456]_ , \new_[9457]_ , \new_[9458]_ ,
    \new_[9460]_ , \new_[9462]_ , \new_[9463]_ , \new_[9464]_ ,
    \new_[9465]_ , \new_[9466]_ , \new_[9467]_ , \new_[9468]_ ,
    \new_[9469]_ , \new_[9471]_ , \new_[9472]_ , \new_[9473]_ ,
    \new_[9474]_ , \new_[9475]_ , \new_[9476]_ , \new_[9477]_ ,
    \new_[9478]_ , \new_[9479]_ , \new_[9480]_ , \new_[9481]_ ,
    \new_[9482]_ , \new_[9483]_ , \new_[9484]_ , \new_[9485]_ ,
    \new_[9486]_ , \new_[9488]_ , \new_[9489]_ , \new_[9490]_ ,
    \new_[9491]_ , \new_[9492]_ , \new_[9493]_ , \new_[9494]_ ,
    \new_[9497]_ , \new_[9499]_ , \new_[9500]_ , \new_[9501]_ ,
    \new_[9502]_ , \new_[9503]_ , \new_[9504]_ , \new_[9505]_ ,
    \new_[9506]_ , \new_[9507]_ , \new_[9508]_ , \new_[9509]_ ,
    \new_[9510]_ , \new_[9511]_ , \new_[9512]_ , \new_[9513]_ ,
    \new_[9514]_ , \new_[9515]_ , \new_[9516]_ , \new_[9517]_ ,
    \new_[9518]_ , \new_[9519]_ , \new_[9520]_ , \new_[9521]_ ,
    \new_[9522]_ , \new_[9523]_ , \new_[9524]_ , \new_[9526]_ ,
    \new_[9528]_ , \new_[9529]_ , \new_[9530]_ , \new_[9531]_ ,
    \new_[9532]_ , \new_[9533]_ , \new_[9534]_ , \new_[9535]_ ,
    \new_[9536]_ , \new_[9537]_ , \new_[9538]_ , \new_[9539]_ ,
    \new_[9540]_ , \new_[9541]_ , \new_[9542]_ , \new_[9543]_ ,
    \new_[9544]_ , \new_[9545]_ , \new_[9546]_ , \new_[9547]_ ,
    \new_[9548]_ , \new_[9549]_ , \new_[9550]_ , \new_[9551]_ ,
    \new_[9552]_ , \new_[9553]_ , \new_[9554]_ , \new_[9555]_ ,
    \new_[9556]_ , \new_[9557]_ , \new_[9558]_ , \new_[9559]_ ,
    \new_[9560]_ , \new_[9561]_ , \new_[9562]_ , \new_[9563]_ ,
    \new_[9564]_ , \new_[9565]_ , \new_[9566]_ , \new_[9567]_ ,
    \new_[9568]_ , \new_[9570]_ , \new_[9571]_ , \new_[9572]_ ,
    \new_[9573]_ , \new_[9574]_ , \new_[9575]_ , \new_[9576]_ ,
    \new_[9578]_ , \new_[9579]_ , \new_[9580]_ , \new_[9581]_ ,
    \new_[9582]_ , \new_[9583]_ , \new_[9584]_ , \new_[9585]_ ,
    \new_[9586]_ , \new_[9587]_ , \new_[9588]_ , \new_[9589]_ ,
    \new_[9590]_ , \new_[9591]_ , \new_[9592]_ , \new_[9593]_ ,
    \new_[9594]_ , \new_[9595]_ , \new_[9596]_ , \new_[9597]_ ,
    \new_[9598]_ , \new_[9599]_ , \new_[9600]_ , \new_[9601]_ ,
    \new_[9602]_ , \new_[9603]_ , \new_[9605]_ , \new_[9607]_ ,
    \new_[9608]_ , \new_[9609]_ , \new_[9610]_ , \new_[9611]_ ,
    \new_[9612]_ , \new_[9613]_ , \new_[9614]_ , \new_[9615]_ ,
    \new_[9616]_ , \new_[9617]_ , \new_[9618]_ , \new_[9619]_ ,
    \new_[9620]_ , \new_[9621]_ , \new_[9622]_ , \new_[9623]_ ,
    \new_[9624]_ , \new_[9625]_ , \new_[9627]_ , \new_[9628]_ ,
    \new_[9629]_ , \new_[9630]_ , \new_[9631]_ , \new_[9632]_ ,
    \new_[9633]_ , \new_[9634]_ , \new_[9635]_ , \new_[9637]_ ,
    \new_[9638]_ , \new_[9639]_ , \new_[9640]_ , \new_[9641]_ ,
    \new_[9642]_ , \new_[9643]_ , \new_[9644]_ , \new_[9645]_ ,
    \new_[9646]_ , \new_[9647]_ , \new_[9648]_ , \new_[9649]_ ,
    \new_[9650]_ , \new_[9651]_ , \new_[9652]_ , \new_[9653]_ ,
    \new_[9654]_ , \new_[9655]_ , \new_[9656]_ , \new_[9657]_ ,
    \new_[9658]_ , \new_[9659]_ , \new_[9660]_ , \new_[9661]_ ,
    \new_[9662]_ , \new_[9663]_ , \new_[9664]_ , \new_[9665]_ ,
    \new_[9666]_ , \new_[9667]_ , \new_[9668]_ , \new_[9669]_ ,
    \new_[9670]_ , \new_[9671]_ , \new_[9672]_ , \new_[9673]_ ,
    \new_[9674]_ , \new_[9675]_ , \new_[9676]_ , \new_[9677]_ ,
    \new_[9678]_ , \new_[9679]_ , \new_[9680]_ , \new_[9681]_ ,
    \new_[9682]_ , \new_[9683]_ , \new_[9684]_ , \new_[9685]_ ,
    \new_[9687]_ , \new_[9688]_ , \new_[9689]_ , \new_[9690]_ ,
    \new_[9691]_ , \new_[9692]_ , \new_[9693]_ , \new_[9694]_ ,
    \new_[9695]_ , \new_[9696]_ , \new_[9697]_ , \new_[9698]_ ,
    \new_[9699]_ , \new_[9700]_ , \new_[9701]_ , \new_[9702]_ ,
    \new_[9703]_ , \new_[9704]_ , \new_[9705]_ , \new_[9707]_ ,
    \new_[9708]_ , \new_[9709]_ , \new_[9710]_ , \new_[9711]_ ,
    \new_[9712]_ , \new_[9714]_ , \new_[9715]_ , \new_[9716]_ ,
    \new_[9717]_ , \new_[9718]_ , \new_[9719]_ , \new_[9720]_ ,
    \new_[9721]_ , \new_[9722]_ , \new_[9723]_ , \new_[9725]_ ,
    \new_[9726]_ , \new_[9727]_ , \new_[9728]_ , \new_[9730]_ ,
    \new_[9731]_ , \new_[9732]_ , \new_[9733]_ , \new_[9734]_ ,
    \new_[9735]_ , \new_[9736]_ , \new_[9737]_ , \new_[9738]_ ,
    \new_[9739]_ , \new_[9740]_ , \new_[9741]_ , \new_[9742]_ ,
    \new_[9744]_ , \new_[9745]_ , \new_[9746]_ , \new_[9747]_ ,
    \new_[9748]_ , \new_[9749]_ , \new_[9750]_ , \new_[9751]_ ,
    \new_[9752]_ , \new_[9753]_ , \new_[9755]_ , \new_[9756]_ ,
    \new_[9757]_ , \new_[9758]_ , \new_[9759]_ , \new_[9760]_ ,
    \new_[9766]_ , \new_[9767]_ , \new_[9768]_ , \new_[9769]_ ,
    \new_[9770]_ , \new_[9771]_ , \new_[9772]_ , \new_[9773]_ ,
    \new_[9774]_ , \new_[9775]_ , \new_[9776]_ , \new_[9777]_ ,
    \new_[9778]_ , \new_[9779]_ , \new_[9780]_ , \new_[9781]_ ,
    \new_[9782]_ , \new_[9783]_ , \new_[9784]_ , \new_[9785]_ ,
    \new_[9786]_ , \new_[9787]_ , \new_[9788]_ , \new_[9789]_ ,
    \new_[9790]_ , \new_[9791]_ , \new_[9792]_ , \new_[9793]_ ,
    \new_[9794]_ , \new_[9795]_ , \new_[9796]_ , \new_[9797]_ ,
    \new_[9798]_ , \new_[9799]_ , \new_[9800]_ , \new_[9801]_ ,
    \new_[9802]_ , \new_[9803]_ , \new_[9804]_ , \new_[9805]_ ,
    \new_[9806]_ , \new_[9807]_ , \new_[9808]_ , \new_[9809]_ ,
    \new_[9810]_ , \new_[9811]_ , \new_[9812]_ , \new_[9813]_ ,
    \new_[9814]_ , \new_[9815]_ , \new_[9816]_ , \new_[9817]_ ,
    \new_[9818]_ , \new_[9819]_ , \new_[9820]_ , \new_[9821]_ ,
    \new_[9822]_ , \new_[9823]_ , \new_[9824]_ , \new_[9825]_ ,
    \new_[9826]_ , \new_[9827]_ , \new_[9828]_ , \new_[9830]_ ,
    \new_[9832]_ , \new_[9834]_ , \new_[9835]_ , \new_[9836]_ ,
    \new_[9837]_ , \new_[9838]_ , \new_[9840]_ , \new_[9841]_ ,
    \new_[9842]_ , \new_[9843]_ , \new_[9844]_ , \new_[9845]_ ,
    \new_[9846]_ , \new_[9847]_ , \new_[9848]_ , \new_[9849]_ ,
    \new_[9850]_ , \new_[9851]_ , \new_[9852]_ , \new_[9853]_ ,
    \new_[9854]_ , \new_[9855]_ , \new_[9856]_ , \new_[9857]_ ,
    \new_[9858]_ , \new_[9859]_ , \new_[9860]_ , \new_[9861]_ ,
    \new_[9862]_ , \new_[9863]_ , \new_[9864]_ , \new_[9865]_ ,
    \new_[9866]_ , \new_[9867]_ , \new_[9868]_ , \new_[9869]_ ,
    \new_[9870]_ , \new_[9871]_ , \new_[9872]_ , \new_[9873]_ ,
    \new_[9874]_ , \new_[9876]_ , \new_[9877]_ , \new_[9878]_ ,
    \new_[9879]_ , \new_[9880]_ , \new_[9881]_ , \new_[9882]_ ,
    \new_[9883]_ , \new_[9884]_ , \new_[9885]_ , \new_[9886]_ ,
    \new_[9887]_ , \new_[9888]_ , \new_[9889]_ , \new_[9890]_ ,
    \new_[9891]_ , \new_[9892]_ , \new_[9893]_ , \new_[9894]_ ,
    \new_[9895]_ , \new_[9896]_ , \new_[9897]_ , \new_[9899]_ ,
    \new_[9900]_ , \new_[9901]_ , \new_[9902]_ , \new_[9903]_ ,
    \new_[9904]_ , \new_[9905]_ , \new_[9906]_ , \new_[9907]_ ,
    \new_[9908]_ , \new_[9909]_ , \new_[9910]_ , \new_[9911]_ ,
    \new_[9913]_ , \new_[9914]_ , \new_[9915]_ , \new_[9916]_ ,
    \new_[9919]_ , \new_[9921]_ , \new_[9923]_ , \new_[9925]_ ,
    \new_[9927]_ , \new_[9929]_ , \new_[9930]_ , \new_[9931]_ ,
    \new_[9932]_ , \new_[9933]_ , \new_[9934]_ , \new_[9935]_ ,
    \new_[9936]_ , \new_[9937]_ , \new_[9938]_ , \new_[9939]_ ,
    \new_[9940]_ , \new_[9941]_ , \new_[9942]_ , \new_[9943]_ ,
    \new_[9945]_ , \new_[9946]_ , \new_[9947]_ , \new_[9949]_ ,
    \new_[9951]_ , \new_[9955]_ , \new_[9956]_ , \new_[9957]_ ,
    \new_[9958]_ , \new_[9959]_ , \new_[9960]_ , \new_[9961]_ ,
    \new_[9962]_ , \new_[9963]_ , \new_[9964]_ , \new_[9965]_ ,
    \new_[9966]_ , \new_[9967]_ , \new_[9968]_ , \new_[9969]_ ,
    \new_[9970]_ , \new_[9971]_ , \new_[9972]_ , \new_[9973]_ ,
    \new_[9974]_ , \new_[9975]_ , \new_[9976]_ , \new_[9977]_ ,
    \new_[9978]_ , \new_[9979]_ , \new_[9980]_ , \new_[9981]_ ,
    \new_[9982]_ , \new_[9983]_ , \new_[9984]_ , \new_[9985]_ ,
    \new_[9986]_ , \new_[9987]_ , \new_[9988]_ , \new_[9989]_ ,
    \new_[9990]_ , \new_[9991]_ , \new_[9992]_ , \new_[9993]_ ,
    \new_[9994]_ , \new_[9995]_ , \new_[9996]_ , \new_[9997]_ ,
    \new_[9998]_ , \new_[9999]_ , \new_[10000]_ , \new_[10001]_ ,
    \new_[10002]_ , \new_[10003]_ , \new_[10004]_ , \new_[10005]_ ,
    \new_[10006]_ , \new_[10007]_ , \new_[10008]_ , \new_[10009]_ ,
    \new_[10010]_ , \new_[10012]_ , \new_[10013]_ , \new_[10014]_ ,
    \new_[10015]_ , \new_[10016]_ , \new_[10017]_ , \new_[10018]_ ,
    \new_[10019]_ , \new_[10020]_ , \new_[10021]_ , \new_[10022]_ ,
    \new_[10023]_ , \new_[10024]_ , \new_[10027]_ , \new_[10028]_ ,
    \new_[10029]_ , \new_[10030]_ , \new_[10031]_ , \new_[10032]_ ,
    \new_[10033]_ , \new_[10034]_ , \new_[10035]_ , \new_[10036]_ ,
    \new_[10037]_ , \new_[10038]_ , \new_[10039]_ , \new_[10040]_ ,
    \new_[10041]_ , \new_[10042]_ , \new_[10043]_ , \new_[10044]_ ,
    \new_[10045]_ , \new_[10046]_ , \new_[10047]_ , \new_[10048]_ ,
    \new_[10049]_ , \new_[10050]_ , \new_[10051]_ , \new_[10052]_ ,
    \new_[10053]_ , \new_[10054]_ , \new_[10055]_ , \new_[10056]_ ,
    \new_[10057]_ , \new_[10058]_ , \new_[10063]_ , \new_[10064]_ ,
    \new_[10065]_ , \new_[10066]_ , \new_[10067]_ , \new_[10068]_ ,
    \new_[10069]_ , \new_[10070]_ , \new_[10071]_ , \new_[10072]_ ,
    \new_[10073]_ , \new_[10074]_ , \new_[10075]_ , \new_[10076]_ ,
    \new_[10077]_ , \new_[10078]_ , \new_[10079]_ , \new_[10080]_ ,
    \new_[10081]_ , \new_[10082]_ , \new_[10083]_ , \new_[10084]_ ,
    \new_[10085]_ , \new_[10086]_ , \new_[10087]_ , \new_[10088]_ ,
    \new_[10089]_ , \new_[10090]_ , \new_[10091]_ , \new_[10092]_ ,
    \new_[10093]_ , \new_[10094]_ , \new_[10095]_ , \new_[10096]_ ,
    \new_[10097]_ , \new_[10098]_ , \new_[10099]_ , \new_[10101]_ ,
    \new_[10102]_ , \new_[10103]_ , \new_[10104]_ , \new_[10105]_ ,
    \new_[10106]_ , \new_[10107]_ , \new_[10108]_ , \new_[10110]_ ,
    \new_[10111]_ , \new_[10112]_ , \new_[10113]_ , \new_[10114]_ ,
    \new_[10115]_ , \new_[10116]_ , \new_[10117]_ , \new_[10118]_ ,
    \new_[10120]_ , \new_[10121]_ , \new_[10122]_ , \new_[10123]_ ,
    \new_[10124]_ , \new_[10125]_ , \new_[10126]_ , \new_[10127]_ ,
    \new_[10128]_ , \new_[10129]_ , \new_[10130]_ , \new_[10131]_ ,
    \new_[10132]_ , \new_[10133]_ , \new_[10134]_ , \new_[10135]_ ,
    \new_[10136]_ , \new_[10137]_ , \new_[10138]_ , \new_[10139]_ ,
    \new_[10140]_ , \new_[10141]_ , \new_[10142]_ , \new_[10143]_ ,
    \new_[10144]_ , \new_[10145]_ , \new_[10146]_ , \new_[10147]_ ,
    \new_[10148]_ , \new_[10149]_ , \new_[10150]_ , \new_[10151]_ ,
    \new_[10152]_ , \new_[10153]_ , \new_[10154]_ , \new_[10155]_ ,
    \new_[10156]_ , \new_[10157]_ , \new_[10158]_ , \new_[10159]_ ,
    \new_[10160]_ , \new_[10161]_ , \new_[10162]_ , \new_[10163]_ ,
    \new_[10164]_ , \new_[10165]_ , \new_[10166]_ , \new_[10167]_ ,
    \new_[10168]_ , \new_[10169]_ , \new_[10170]_ , \new_[10171]_ ,
    \new_[10172]_ , \new_[10173]_ , \new_[10174]_ , \new_[10175]_ ,
    \new_[10176]_ , \new_[10177]_ , \new_[10178]_ , \new_[10179]_ ,
    \new_[10180]_ , \new_[10181]_ , \new_[10182]_ , \new_[10183]_ ,
    \new_[10184]_ , \new_[10185]_ , \new_[10186]_ , \new_[10187]_ ,
    \new_[10188]_ , \new_[10189]_ , \new_[10190]_ , \new_[10191]_ ,
    \new_[10192]_ , \new_[10193]_ , \new_[10194]_ , \new_[10195]_ ,
    \new_[10196]_ , \new_[10197]_ , \new_[10198]_ , \new_[10199]_ ,
    \new_[10200]_ , \new_[10201]_ , \new_[10202]_ , \new_[10203]_ ,
    \new_[10204]_ , \new_[10205]_ , \new_[10206]_ , \new_[10207]_ ,
    \new_[10208]_ , \new_[10209]_ , \new_[10210]_ , \new_[10211]_ ,
    \new_[10212]_ , \new_[10213]_ , \new_[10214]_ , \new_[10215]_ ,
    \new_[10216]_ , \new_[10217]_ , \new_[10218]_ , \new_[10219]_ ,
    \new_[10220]_ , \new_[10221]_ , \new_[10222]_ , \new_[10224]_ ,
    \new_[10225]_ , \new_[10226]_ , \new_[10227]_ , \new_[10228]_ ,
    \new_[10229]_ , \new_[10230]_ , \new_[10231]_ , \new_[10233]_ ,
    \new_[10234]_ , \new_[10235]_ , \new_[10236]_ , \new_[10237]_ ,
    \new_[10238]_ , \new_[10239]_ , \new_[10240]_ , \new_[10241]_ ,
    \new_[10242]_ , \new_[10243]_ , \new_[10244]_ , \new_[10245]_ ,
    \new_[10246]_ , \new_[10247]_ , \new_[10248]_ , \new_[10249]_ ,
    \new_[10251]_ , \new_[10252]_ , \new_[10253]_ , \new_[10254]_ ,
    \new_[10255]_ , \new_[10256]_ , \new_[10257]_ , \new_[10258]_ ,
    \new_[10259]_ , \new_[10260]_ , \new_[10261]_ , \new_[10262]_ ,
    \new_[10263]_ , \new_[10264]_ , \new_[10265]_ , \new_[10266]_ ,
    \new_[10267]_ , \new_[10268]_ , \new_[10269]_ , \new_[10270]_ ,
    \new_[10271]_ , \new_[10272]_ , \new_[10273]_ , \new_[10274]_ ,
    \new_[10275]_ , \new_[10276]_ , \new_[10277]_ , \new_[10278]_ ,
    \new_[10279]_ , \new_[10280]_ , \new_[10281]_ , \new_[10282]_ ,
    \new_[10283]_ , \new_[10284]_ , \new_[10285]_ , \new_[10286]_ ,
    \new_[10287]_ , \new_[10288]_ , \new_[10289]_ , \new_[10291]_ ,
    \new_[10292]_ , \new_[10295]_ , \new_[10296]_ , \new_[10297]_ ,
    \new_[10298]_ , \new_[10299]_ , \new_[10300]_ , \new_[10301]_ ,
    \new_[10302]_ , \new_[10303]_ , \new_[10304]_ , \new_[10305]_ ,
    \new_[10306]_ , \new_[10307]_ , \new_[10308]_ , \new_[10309]_ ,
    \new_[10310]_ , \new_[10311]_ , \new_[10313]_ , \new_[10314]_ ,
    \new_[10315]_ , \new_[10316]_ , \new_[10317]_ , \new_[10318]_ ,
    \new_[10319]_ , \new_[10320]_ , \new_[10322]_ , \new_[10323]_ ,
    \new_[10325]_ , \new_[10326]_ , \new_[10327]_ , \new_[10329]_ ,
    \new_[10330]_ , \new_[10331]_ , \new_[10332]_ , \new_[10333]_ ,
    \new_[10334]_ , \new_[10338]_ , \new_[10339]_ , \new_[10340]_ ,
    \new_[10341]_ , \new_[10342]_ , \new_[10344]_ , \new_[10345]_ ,
    \new_[10347]_ , \new_[10348]_ , \new_[10349]_ , \new_[10350]_ ,
    \new_[10351]_ , \new_[10352]_ , \new_[10353]_ , \new_[10354]_ ,
    \new_[10355]_ , \new_[10356]_ , \new_[10357]_ , \new_[10358]_ ,
    \new_[10359]_ , \new_[10360]_ , \new_[10362]_ , \new_[10363]_ ,
    \new_[10364]_ , \new_[10365]_ , \new_[10366]_ , \new_[10368]_ ,
    \new_[10369]_ , \new_[10370]_ , \new_[10371]_ , \new_[10372]_ ,
    \new_[10373]_ , \new_[10375]_ , \new_[10376]_ , \new_[10377]_ ,
    \new_[10378]_ , \new_[10379]_ , \new_[10380]_ , \new_[10381]_ ,
    \new_[10382]_ , \new_[10383]_ , \new_[10384]_ , \new_[10385]_ ,
    \new_[10386]_ , \new_[10387]_ , \new_[10388]_ , \new_[10389]_ ,
    \new_[10390]_ , \new_[10391]_ , \new_[10392]_ , \new_[10393]_ ,
    \new_[10394]_ , \new_[10395]_ , \new_[10396]_ , \new_[10397]_ ,
    \new_[10398]_ , \new_[10399]_ , \new_[10400]_ , \new_[10401]_ ,
    \new_[10402]_ , \new_[10403]_ , \new_[10404]_ , \new_[10405]_ ,
    \new_[10406]_ , \new_[10407]_ , \new_[10408]_ , \new_[10409]_ ,
    \new_[10410]_ , \new_[10411]_ , \new_[10413]_ , \new_[10414]_ ,
    \new_[10415]_ , \new_[10416]_ , \new_[10417]_ , \new_[10418]_ ,
    \new_[10419]_ , \new_[10420]_ , \new_[10421]_ , \new_[10422]_ ,
    \new_[10423]_ , \new_[10424]_ , \new_[10425]_ , \new_[10426]_ ,
    \new_[10427]_ , \new_[10428]_ , \new_[10429]_ , \new_[10430]_ ,
    \new_[10431]_ , \new_[10432]_ , \new_[10433]_ , \new_[10434]_ ,
    \new_[10435]_ , \new_[10436]_ , \new_[10437]_ , \new_[10438]_ ,
    \new_[10439]_ , \new_[10440]_ , \new_[10441]_ , \new_[10442]_ ,
    \new_[10443]_ , \new_[10444]_ , \new_[10445]_ , \new_[10446]_ ,
    \new_[10447]_ , \new_[10448]_ , \new_[10449]_ , \new_[10450]_ ,
    \new_[10451]_ , \new_[10452]_ , \new_[10453]_ , \new_[10454]_ ,
    \new_[10455]_ , \new_[10456]_ , \new_[10457]_ , \new_[10458]_ ,
    \new_[10459]_ , \new_[10460]_ , \new_[10461]_ , \new_[10462]_ ,
    \new_[10463]_ , \new_[10464]_ , \new_[10465]_ , \new_[10466]_ ,
    \new_[10467]_ , \new_[10468]_ , \new_[10469]_ , \new_[10470]_ ,
    \new_[10471]_ , \new_[10472]_ , \new_[10473]_ , \new_[10474]_ ,
    \new_[10475]_ , \new_[10476]_ , \new_[10477]_ , \new_[10478]_ ,
    \new_[10479]_ , \new_[10480]_ , \new_[10481]_ , \new_[10482]_ ,
    \new_[10483]_ , \new_[10484]_ , \new_[10485]_ , \new_[10486]_ ,
    \new_[10487]_ , \new_[10488]_ , \new_[10489]_ , \new_[10490]_ ,
    \new_[10491]_ , \new_[10492]_ , \new_[10493]_ , \new_[10494]_ ,
    \new_[10495]_ , \new_[10496]_ , \new_[10497]_ , \new_[10498]_ ,
    \new_[10499]_ , \new_[10500]_ , \new_[10501]_ , \new_[10502]_ ,
    \new_[10503]_ , \new_[10505]_ , \new_[10506]_ , \new_[10507]_ ,
    \new_[10508]_ , \new_[10509]_ , \new_[10510]_ , \new_[10511]_ ,
    \new_[10512]_ , \new_[10513]_ , \new_[10514]_ , \new_[10515]_ ,
    \new_[10516]_ , \new_[10517]_ , \new_[10518]_ , \new_[10519]_ ,
    \new_[10520]_ , \new_[10521]_ , \new_[10522]_ , \new_[10523]_ ,
    \new_[10524]_ , \new_[10525]_ , \new_[10526]_ , \new_[10527]_ ,
    \new_[10528]_ , \new_[10529]_ , \new_[10530]_ , \new_[10531]_ ,
    \new_[10532]_ , \new_[10533]_ , \new_[10534]_ , \new_[10535]_ ,
    \new_[10536]_ , \new_[10537]_ , \new_[10538]_ , \new_[10539]_ ,
    \new_[10540]_ , \new_[10541]_ , \new_[10542]_ , \new_[10543]_ ,
    \new_[10544]_ , \new_[10545]_ , \new_[10546]_ , \new_[10547]_ ,
    \new_[10548]_ , \new_[10549]_ , \new_[10550]_ , \new_[10551]_ ,
    \new_[10552]_ , \new_[10553]_ , \new_[10554]_ , \new_[10555]_ ,
    \new_[10556]_ , \new_[10557]_ , \new_[10558]_ , \new_[10559]_ ,
    \new_[10560]_ , \new_[10561]_ , \new_[10562]_ , \new_[10563]_ ,
    \new_[10564]_ , \new_[10565]_ , \new_[10566]_ , \new_[10567]_ ,
    \new_[10568]_ , \new_[10569]_ , \new_[10570]_ , \new_[10571]_ ,
    \new_[10572]_ , \new_[10573]_ , \new_[10574]_ , \new_[10575]_ ,
    \new_[10576]_ , \new_[10577]_ , \new_[10578]_ , \new_[10579]_ ,
    \new_[10580]_ , \new_[10581]_ , \new_[10582]_ , \new_[10583]_ ,
    \new_[10584]_ , \new_[10585]_ , \new_[10586]_ , \new_[10587]_ ,
    \new_[10588]_ , \new_[10589]_ , \new_[10590]_ , \new_[10591]_ ,
    \new_[10592]_ , \new_[10593]_ , \new_[10594]_ , \new_[10595]_ ,
    \new_[10596]_ , \new_[10597]_ , \new_[10598]_ , \new_[10599]_ ,
    \new_[10600]_ , \new_[10601]_ , \new_[10602]_ , \new_[10603]_ ,
    \new_[10604]_ , \new_[10605]_ , \new_[10606]_ , \new_[10607]_ ,
    \new_[10608]_ , \new_[10609]_ , \new_[10610]_ , \new_[10611]_ ,
    \new_[10612]_ , \new_[10613]_ , \new_[10614]_ , \new_[10615]_ ,
    \new_[10617]_ , \new_[10618]_ , \new_[10619]_ , \new_[10620]_ ,
    \new_[10621]_ , \new_[10622]_ , \new_[10623]_ , \new_[10624]_ ,
    \new_[10625]_ , \new_[10626]_ , \new_[10627]_ , \new_[10628]_ ,
    \new_[10629]_ , \new_[10630]_ , \new_[10631]_ , \new_[10632]_ ,
    \new_[10633]_ , \new_[10634]_ , \new_[10635]_ , \new_[10636]_ ,
    \new_[10637]_ , \new_[10638]_ , \new_[10639]_ , \new_[10640]_ ,
    \new_[10641]_ , \new_[10642]_ , \new_[10643]_ , \new_[10644]_ ,
    \new_[10645]_ , \new_[10646]_ , \new_[10647]_ , \new_[10648]_ ,
    \new_[10649]_ , \new_[10650]_ , \new_[10651]_ , \new_[10652]_ ,
    \new_[10653]_ , \new_[10654]_ , \new_[10655]_ , \new_[10656]_ ,
    \new_[10657]_ , \new_[10658]_ , \new_[10659]_ , \new_[10660]_ ,
    \new_[10661]_ , \new_[10662]_ , \new_[10663]_ , \new_[10664]_ ,
    \new_[10665]_ , \new_[10666]_ , \new_[10667]_ , \new_[10668]_ ,
    \new_[10669]_ , \new_[10670]_ , \new_[10671]_ , \new_[10672]_ ,
    \new_[10673]_ , \new_[10674]_ , \new_[10675]_ , \new_[10676]_ ,
    \new_[10677]_ , \new_[10678]_ , \new_[10679]_ , \new_[10680]_ ,
    \new_[10681]_ , \new_[10682]_ , \new_[10683]_ , \new_[10684]_ ,
    \new_[10685]_ , \new_[10686]_ , \new_[10687]_ , \new_[10688]_ ,
    \new_[10689]_ , \new_[10690]_ , \new_[10691]_ , \new_[10692]_ ,
    \new_[10693]_ , \new_[10694]_ , \new_[10695]_ , \new_[10696]_ ,
    \new_[10697]_ , \new_[10698]_ , \new_[10699]_ , \new_[10700]_ ,
    \new_[10701]_ , \new_[10702]_ , \new_[10703]_ , \new_[10704]_ ,
    \new_[10705]_ , \new_[10706]_ , \new_[10707]_ , \new_[10708]_ ,
    \new_[10709]_ , \new_[10710]_ , \new_[10711]_ , \new_[10712]_ ,
    \new_[10713]_ , \new_[10714]_ , \new_[10715]_ , \new_[10716]_ ,
    \new_[10717]_ , \new_[10718]_ , \new_[10719]_ , \new_[10720]_ ,
    \new_[10721]_ , \new_[10722]_ , \new_[10723]_ , \new_[10724]_ ,
    \new_[10725]_ , \new_[10726]_ , \new_[10727]_ , \new_[10728]_ ,
    \new_[10729]_ , \new_[10730]_ , \new_[10731]_ , \new_[10732]_ ,
    \new_[10733]_ , \new_[10734]_ , \new_[10735]_ , \new_[10736]_ ,
    \new_[10737]_ , \new_[10738]_ , \new_[10739]_ , \new_[10740]_ ,
    \new_[10741]_ , \new_[10742]_ , \new_[10743]_ , \new_[10744]_ ,
    \new_[10745]_ , \new_[10746]_ , \new_[10747]_ , \new_[10748]_ ,
    \new_[10749]_ , \new_[10750]_ , \new_[10751]_ , \new_[10752]_ ,
    \new_[10753]_ , \new_[10754]_ , \new_[10755]_ , \new_[10756]_ ,
    \new_[10757]_ , \new_[10758]_ , \new_[10759]_ , \new_[10760]_ ,
    \new_[10761]_ , \new_[10762]_ , \new_[10763]_ , \new_[10764]_ ,
    \new_[10766]_ , \new_[10767]_ , \new_[10768]_ , \new_[10769]_ ,
    \new_[10771]_ , \new_[10772]_ , \new_[10773]_ , \new_[10774]_ ,
    \new_[10777]_ , \new_[10778]_ , \new_[10779]_ , \new_[10780]_ ,
    \new_[10785]_ , \new_[10786]_ , \new_[10787]_ , \new_[10788]_ ,
    \new_[10789]_ , \new_[10790]_ , \new_[10791]_ , \new_[10792]_ ,
    \new_[10793]_ , \new_[10794]_ , \new_[10795]_ , \new_[10796]_ ,
    \new_[10797]_ , \new_[10798]_ , \new_[10799]_ , \new_[10800]_ ,
    \new_[10801]_ , \new_[10802]_ , \new_[10803]_ , \new_[10804]_ ,
    \new_[10805]_ , \new_[10806]_ , \new_[10807]_ , \new_[10808]_ ,
    \new_[10809]_ , \new_[10810]_ , \new_[10811]_ , \new_[10812]_ ,
    \new_[10813]_ , \new_[10814]_ , \new_[10815]_ , \new_[10816]_ ,
    \new_[10817]_ , \new_[10818]_ , \new_[10819]_ , \new_[10820]_ ,
    \new_[10821]_ , \new_[10822]_ , \new_[10823]_ , \new_[10824]_ ,
    \new_[10825]_ , \new_[10826]_ , \new_[10827]_ , \new_[10828]_ ,
    \new_[10829]_ , \new_[10830]_ , \new_[10831]_ , \new_[10832]_ ,
    \new_[10833]_ , \new_[10834]_ , \new_[10835]_ , \new_[10836]_ ,
    \new_[10837]_ , \new_[10838]_ , \new_[10839]_ , \new_[10840]_ ,
    \new_[10841]_ , \new_[10842]_ , \new_[10843]_ , \new_[10844]_ ,
    \new_[10845]_ , \new_[10846]_ , \new_[10847]_ , \new_[10848]_ ,
    \new_[10849]_ , \new_[10850]_ , \new_[10851]_ , \new_[10852]_ ,
    \new_[10853]_ , \new_[10854]_ , \new_[10855]_ , \new_[10856]_ ,
    \new_[10857]_ , \new_[10858]_ , \new_[10859]_ , \new_[10860]_ ,
    \new_[10861]_ , \new_[10862]_ , \new_[10863]_ , \new_[10864]_ ,
    \new_[10865]_ , \new_[10866]_ , \new_[10867]_ , \new_[10868]_ ,
    \new_[10869]_ , \new_[10870]_ , \new_[10871]_ , \new_[10872]_ ,
    \new_[10873]_ , \new_[10874]_ , \new_[10875]_ , \new_[10876]_ ,
    \new_[10877]_ , \new_[10878]_ , \new_[10879]_ , \new_[10880]_ ,
    \new_[10881]_ , \new_[10882]_ , \new_[10883]_ , \new_[10884]_ ,
    \new_[10885]_ , \new_[10886]_ , \new_[10887]_ , \new_[10888]_ ,
    \new_[10889]_ , \new_[10890]_ , \new_[10891]_ , \new_[10892]_ ,
    \new_[10893]_ , \new_[10894]_ , \new_[10895]_ , \new_[10896]_ ,
    \new_[10897]_ , \new_[10898]_ , \new_[10899]_ , \new_[10900]_ ,
    \new_[10901]_ , \new_[10902]_ , \new_[10903]_ , \new_[10904]_ ,
    \new_[10905]_ , \new_[10906]_ , \new_[10907]_ , \new_[10908]_ ,
    \new_[10909]_ , \new_[10910]_ , \new_[10911]_ , \new_[10912]_ ,
    \new_[10913]_ , \new_[10914]_ , \new_[10915]_ , \new_[10917]_ ,
    \new_[10918]_ , \new_[10919]_ , \new_[10920]_ , \new_[10921]_ ,
    \new_[10922]_ , \new_[10923]_ , \new_[10924]_ , \new_[10925]_ ,
    \new_[10926]_ , \new_[10927]_ , \new_[10928]_ , \new_[10929]_ ,
    \new_[10930]_ , \new_[10931]_ , \new_[10932]_ , \new_[10933]_ ,
    \new_[10934]_ , \new_[10935]_ , \new_[10936]_ , \new_[10937]_ ,
    \new_[10938]_ , \new_[10939]_ , \new_[10940]_ , \new_[10941]_ ,
    \new_[10942]_ , \new_[10943]_ , \new_[10944]_ , \new_[10945]_ ,
    \new_[10946]_ , \new_[10947]_ , \new_[10948]_ , \new_[10949]_ ,
    \new_[10950]_ , \new_[10951]_ , \new_[10952]_ , \new_[10953]_ ,
    \new_[10954]_ , \new_[10955]_ , \new_[10956]_ , \new_[10957]_ ,
    \new_[10958]_ , \new_[10959]_ , \new_[10960]_ , \new_[10961]_ ,
    \new_[10962]_ , \new_[10963]_ , \new_[10964]_ , \new_[10965]_ ,
    \new_[10966]_ , \new_[10967]_ , \new_[10968]_ , \new_[10969]_ ,
    \new_[10970]_ , \new_[10971]_ , \new_[10972]_ , \new_[10973]_ ,
    \new_[10974]_ , \new_[10975]_ , \new_[10976]_ , \new_[10978]_ ,
    \new_[10979]_ , \new_[10980]_ , \new_[10981]_ , \new_[10982]_ ,
    \new_[10983]_ , \new_[10984]_ , \new_[10985]_ , \new_[10986]_ ,
    \new_[10987]_ , \new_[10988]_ , \new_[10989]_ , \new_[10990]_ ,
    \new_[10991]_ , \new_[10992]_ , \new_[10993]_ , \new_[10994]_ ,
    \new_[10995]_ , \new_[10996]_ , \new_[10997]_ , \new_[10998]_ ,
    \new_[10999]_ , \new_[11000]_ , \new_[11005]_ , \new_[11006]_ ,
    \new_[11007]_ , \new_[11008]_ , \new_[11009]_ , \new_[11010]_ ,
    \new_[11011]_ , \new_[11012]_ , \new_[11013]_ , \new_[11014]_ ,
    \new_[11015]_ , \new_[11016]_ , \new_[11017]_ , \new_[11018]_ ,
    \new_[11019]_ , \new_[11020]_ , \new_[11021]_ , \new_[11022]_ ,
    \new_[11023]_ , \new_[11024]_ , \new_[11025]_ , \new_[11026]_ ,
    \new_[11027]_ , \new_[11028]_ , \new_[11029]_ , \new_[11030]_ ,
    \new_[11035]_ , \new_[11040]_ , \new_[11041]_ , \new_[11042]_ ,
    \new_[11043]_ , \new_[11044]_ , \new_[11045]_ , \new_[11046]_ ,
    \new_[11047]_ , \new_[11048]_ , \new_[11049]_ , \new_[11050]_ ,
    \new_[11051]_ , \new_[11052]_ , \new_[11053]_ , \new_[11054]_ ,
    \new_[11055]_ , \new_[11056]_ , \new_[11057]_ , \new_[11058]_ ,
    \new_[11059]_ , \new_[11060]_ , \new_[11061]_ , \new_[11062]_ ,
    \new_[11063]_ , \new_[11064]_ , \new_[11065]_ , \new_[11066]_ ,
    \new_[11067]_ , \new_[11068]_ , \new_[11069]_ , \new_[11070]_ ,
    \new_[11071]_ , \new_[11072]_ , \new_[11073]_ , \new_[11074]_ ,
    \new_[11075]_ , \new_[11076]_ , \new_[11077]_ , \new_[11078]_ ,
    \new_[11079]_ , \new_[11080]_ , \new_[11081]_ , \new_[11082]_ ,
    \new_[11083]_ , \new_[11084]_ , \new_[11085]_ , \new_[11086]_ ,
    \new_[11087]_ , \new_[11088]_ , \new_[11089]_ , \new_[11091]_ ,
    \new_[11092]_ , \new_[11093]_ , \new_[11094]_ , \new_[11095]_ ,
    \new_[11096]_ , \new_[11097]_ , \new_[11098]_ , \new_[11099]_ ,
    \new_[11100]_ , \new_[11101]_ , \new_[11103]_ , \new_[11104]_ ,
    \new_[11105]_ , \new_[11106]_ , \new_[11107]_ , \new_[11111]_ ,
    \new_[11112]_ , \new_[11113]_ , \new_[11114]_ , \new_[11115]_ ,
    \new_[11116]_ , \new_[11117]_ , \new_[11118]_ , \new_[11119]_ ,
    \new_[11120]_ , \new_[11121]_ , \new_[11122]_ , \new_[11123]_ ,
    \new_[11124]_ , \new_[11125]_ , \new_[11126]_ , \new_[11127]_ ,
    \new_[11128]_ , \new_[11129]_ , \new_[11130]_ , \new_[11131]_ ,
    \new_[11132]_ , \new_[11133]_ , \new_[11134]_ , \new_[11135]_ ,
    \new_[11136]_ , \new_[11137]_ , \new_[11138]_ , \new_[11139]_ ,
    \new_[11140]_ , \new_[11141]_ , \new_[11142]_ , \new_[11143]_ ,
    \new_[11144]_ , \new_[11145]_ , \new_[11146]_ , \new_[11147]_ ,
    \new_[11148]_ , \new_[11149]_ , \new_[11150]_ , \new_[11151]_ ,
    \new_[11152]_ , \new_[11153]_ , \new_[11154]_ , \new_[11155]_ ,
    \new_[11156]_ , \new_[11157]_ , \new_[11158]_ , \new_[11159]_ ,
    \new_[11160]_ , \new_[11161]_ , \new_[11162]_ , \new_[11163]_ ,
    \new_[11164]_ , \new_[11165]_ , \new_[11166]_ , \new_[11167]_ ,
    \new_[11168]_ , \new_[11169]_ , \new_[11170]_ , \new_[11171]_ ,
    \new_[11172]_ , \new_[11173]_ , \new_[11174]_ , \new_[11175]_ ,
    \new_[11176]_ , \new_[11177]_ , \new_[11178]_ , \new_[11179]_ ,
    \new_[11180]_ , \new_[11181]_ , \new_[11182]_ , \new_[11183]_ ,
    \new_[11184]_ , \new_[11185]_ , \new_[11186]_ , \new_[11187]_ ,
    \new_[11188]_ , \new_[11189]_ , \new_[11190]_ , \new_[11191]_ ,
    \new_[11192]_ , \new_[11193]_ , \new_[11194]_ , \new_[11195]_ ,
    \new_[11196]_ , \new_[11197]_ , \new_[11198]_ , \new_[11199]_ ,
    \new_[11200]_ , \new_[11201]_ , \new_[11202]_ , \new_[11203]_ ,
    \new_[11204]_ , \new_[11205]_ , \new_[11206]_ , \new_[11207]_ ,
    \new_[11208]_ , \new_[11209]_ , \new_[11210]_ , \new_[11211]_ ,
    \new_[11212]_ , \new_[11213]_ , \new_[11214]_ , \new_[11215]_ ,
    \new_[11216]_ , \new_[11217]_ , \new_[11218]_ , \new_[11219]_ ,
    \new_[11220]_ , \new_[11221]_ , \new_[11229]_ , \new_[11231]_ ,
    \new_[11232]_ , \new_[11233]_ , \new_[11234]_ , \new_[11235]_ ,
    \new_[11236]_ , \new_[11237]_ , \new_[11238]_ , \new_[11239]_ ,
    \new_[11240]_ , \new_[11241]_ , \new_[11242]_ , \new_[11243]_ ,
    \new_[11244]_ , \new_[11245]_ , \new_[11246]_ , \new_[11248]_ ,
    \new_[11249]_ , \new_[11250]_ , \new_[11251]_ , \new_[11252]_ ,
    \new_[11253]_ , \new_[11255]_ , \new_[11256]_ , \new_[11257]_ ,
    \new_[11259]_ , \new_[11260]_ , \new_[11261]_ , \new_[11263]_ ,
    \new_[11264]_ , \new_[11265]_ , \new_[11266]_ , \new_[11268]_ ,
    \new_[11269]_ , \new_[11270]_ , \new_[11271]_ , \new_[11272]_ ,
    \new_[11273]_ , \new_[11274]_ , \new_[11275]_ , \new_[11276]_ ,
    \new_[11277]_ , \new_[11278]_ , \new_[11280]_ , \new_[11281]_ ,
    \new_[11282]_ , \new_[11283]_ , \new_[11284]_ , \new_[11285]_ ,
    \new_[11286]_ , \new_[11287]_ , \new_[11288]_ , \new_[11289]_ ,
    \new_[11290]_ , \new_[11291]_ , \new_[11292]_ , \new_[11293]_ ,
    \new_[11294]_ , \new_[11295]_ , \new_[11296]_ , \new_[11297]_ ,
    \new_[11298]_ , \new_[11299]_ , \new_[11300]_ , \new_[11301]_ ,
    \new_[11302]_ , \new_[11303]_ , \new_[11304]_ , \new_[11305]_ ,
    \new_[11306]_ , \new_[11307]_ , \new_[11308]_ , \new_[11309]_ ,
    \new_[11310]_ , \new_[11312]_ , \new_[11313]_ , \new_[11314]_ ,
    \new_[11315]_ , \new_[11316]_ , \new_[11318]_ , \new_[11319]_ ,
    \new_[11321]_ , \new_[11322]_ , \new_[11323]_ , \new_[11324]_ ,
    \new_[11325]_ , \new_[11326]_ , \new_[11327]_ , \new_[11328]_ ,
    \new_[11329]_ , \new_[11330]_ , \new_[11331]_ , \new_[11332]_ ,
    \new_[11333]_ , \new_[11334]_ , \new_[11335]_ , \new_[11336]_ ,
    \new_[11337]_ , \new_[11338]_ , \new_[11346]_ , \new_[11349]_ ,
    \new_[11352]_ , \new_[11354]_ , \new_[11355]_ , \new_[11356]_ ,
    \new_[11358]_ , \new_[11362]_ , \new_[11363]_ , \new_[11364]_ ,
    \new_[11365]_ , \new_[11368]_ , \new_[11369]_ , \new_[11371]_ ,
    \new_[11373]_ , \new_[11377]_ , \new_[11378]_ , \new_[11379]_ ,
    \new_[11380]_ , \new_[11381]_ , \new_[11382]_ , \new_[11383]_ ,
    \new_[11384]_ , \new_[11386]_ , \new_[11387]_ , \new_[11388]_ ,
    \new_[11390]_ , \new_[11391]_ , \new_[11392]_ , \new_[11393]_ ,
    \new_[11394]_ , \new_[11395]_ , \new_[11396]_ , \new_[11397]_ ,
    \new_[11398]_ , \new_[11399]_ , \new_[11400]_ , \new_[11403]_ ,
    \new_[11404]_ , \new_[11405]_ , \new_[11406]_ , \new_[11407]_ ,
    \new_[11408]_ , \new_[11410]_ , \new_[11411]_ , \new_[11412]_ ,
    \new_[11413]_ , \new_[11414]_ , \new_[11415]_ , \new_[11417]_ ,
    \new_[11418]_ , \new_[11419]_ , \new_[11420]_ , \new_[11421]_ ,
    \new_[11422]_ , \new_[11423]_ , \new_[11424]_ , \new_[11425]_ ,
    \new_[11426]_ , \new_[11427]_ , \new_[11428]_ , \new_[11429]_ ,
    \new_[11430]_ , \new_[11431]_ , \new_[11432]_ , \new_[11433]_ ,
    \new_[11434]_ , \new_[11435]_ , \new_[11436]_ , \new_[11437]_ ,
    \new_[11438]_ , \new_[11439]_ , \new_[11440]_ , \new_[11441]_ ,
    \new_[11442]_ , \new_[11443]_ , \new_[11444]_ , \new_[11445]_ ,
    \new_[11446]_ , \new_[11447]_ , \new_[11448]_ , \new_[11449]_ ,
    \new_[11450]_ , \new_[11452]_ , \new_[11453]_ , \new_[11454]_ ,
    \new_[11455]_ , \new_[11456]_ , \new_[11457]_ , \new_[11458]_ ,
    \new_[11459]_ , \new_[11460]_ , \new_[11461]_ , \new_[11462]_ ,
    \new_[11463]_ , \new_[11464]_ , \new_[11465]_ , \new_[11466]_ ,
    \new_[11467]_ , \new_[11468]_ , \new_[11469]_ , \new_[11470]_ ,
    \new_[11471]_ , \new_[11472]_ , \new_[11473]_ , \new_[11474]_ ,
    \new_[11475]_ , \new_[11476]_ , \new_[11477]_ , \new_[11478]_ ,
    \new_[11479]_ , \new_[11480]_ , \new_[11481]_ , \new_[11482]_ ,
    \new_[11483]_ , \new_[11484]_ , \new_[11485]_ , \new_[11486]_ ,
    \new_[11487]_ , \new_[11488]_ , \new_[11489]_ , \new_[11490]_ ,
    \new_[11491]_ , \new_[11492]_ , \new_[11493]_ , \new_[11494]_ ,
    \new_[11495]_ , \new_[11496]_ , \new_[11497]_ , \new_[11498]_ ,
    \new_[11499]_ , \new_[11500]_ , \new_[11501]_ , \new_[11502]_ ,
    \new_[11503]_ , \new_[11504]_ , \new_[11505]_ , \new_[11506]_ ,
    \new_[11507]_ , \new_[11508]_ , \new_[11509]_ , \new_[11510]_ ,
    \new_[11511]_ , \new_[11512]_ , \new_[11513]_ , \new_[11514]_ ,
    \new_[11515]_ , \new_[11516]_ , \new_[11517]_ , \new_[11518]_ ,
    \new_[11519]_ , \new_[11520]_ , \new_[11521]_ , \new_[11522]_ ,
    \new_[11523]_ , \new_[11524]_ , \new_[11525]_ , \new_[11526]_ ,
    \new_[11527]_ , \new_[11528]_ , \new_[11529]_ , \new_[11530]_ ,
    \new_[11531]_ , \new_[11532]_ , \new_[11533]_ , \new_[11534]_ ,
    \new_[11535]_ , \new_[11536]_ , \new_[11537]_ , \new_[11538]_ ,
    \new_[11539]_ , \new_[11540]_ , \new_[11541]_ , \new_[11542]_ ,
    \new_[11543]_ , \new_[11544]_ , \new_[11545]_ , \new_[11546]_ ,
    \new_[11547]_ , \new_[11548]_ , \new_[11549]_ , \new_[11550]_ ,
    \new_[11551]_ , \new_[11552]_ , \new_[11553]_ , \new_[11554]_ ,
    \new_[11555]_ , \new_[11556]_ , \new_[11557]_ , \new_[11558]_ ,
    \new_[11559]_ , \new_[11560]_ , \new_[11561]_ , \new_[11562]_ ,
    \new_[11563]_ , \new_[11564]_ , \new_[11565]_ , \new_[11566]_ ,
    \new_[11567]_ , \new_[11568]_ , \new_[11569]_ , \new_[11570]_ ,
    \new_[11571]_ , \new_[11572]_ , \new_[11573]_ , \new_[11574]_ ,
    \new_[11575]_ , \new_[11576]_ , \new_[11577]_ , \new_[11578]_ ,
    \new_[11579]_ , \new_[11580]_ , \new_[11581]_ , \new_[11582]_ ,
    \new_[11583]_ , \new_[11584]_ , \new_[11585]_ , \new_[11586]_ ,
    \new_[11587]_ , \new_[11588]_ , \new_[11589]_ , \new_[11590]_ ,
    \new_[11591]_ , \new_[11592]_ , \new_[11593]_ , \new_[11594]_ ,
    \new_[11595]_ , \new_[11596]_ , \new_[11597]_ , \new_[11598]_ ,
    \new_[11599]_ , \new_[11600]_ , \new_[11601]_ , \new_[11602]_ ,
    \new_[11603]_ , \new_[11604]_ , \new_[11605]_ , \new_[11606]_ ,
    \new_[11607]_ , \new_[11608]_ , \new_[11609]_ , \new_[11610]_ ,
    \new_[11611]_ , \new_[11612]_ , \new_[11613]_ , \new_[11614]_ ,
    \new_[11615]_ , \new_[11616]_ , \new_[11617]_ , \new_[11618]_ ,
    \new_[11619]_ , \new_[11620]_ , \new_[11621]_ , \new_[11622]_ ,
    \new_[11623]_ , \new_[11624]_ , \new_[11625]_ , \new_[11626]_ ,
    \new_[11627]_ , \new_[11628]_ , \new_[11629]_ , \new_[11630]_ ,
    \new_[11631]_ , \new_[11632]_ , \new_[11633]_ , \new_[11634]_ ,
    \new_[11635]_ , \new_[11636]_ , \new_[11637]_ , \new_[11638]_ ,
    \new_[11639]_ , \new_[11640]_ , \new_[11642]_ , \new_[11643]_ ,
    \new_[11644]_ , \new_[11645]_ , \new_[11647]_ , \new_[11648]_ ,
    \new_[11649]_ , \new_[11650]_ , \new_[11651]_ , \new_[11652]_ ,
    \new_[11653]_ , \new_[11654]_ , \new_[11655]_ , \new_[11657]_ ,
    \new_[11658]_ , \new_[11659]_ , \new_[11660]_ , \new_[11661]_ ,
    \new_[11662]_ , \new_[11663]_ , \new_[11664]_ , \new_[11665]_ ,
    \new_[11666]_ , \new_[11668]_ , \new_[11669]_ , \new_[11671]_ ,
    \new_[11672]_ , \new_[11673]_ , \new_[11674]_ , \new_[11675]_ ,
    \new_[11676]_ , \new_[11677]_ , \new_[11678]_ , \new_[11679]_ ,
    \new_[11680]_ , \new_[11681]_ , \new_[11682]_ , \new_[11683]_ ,
    \new_[11684]_ , \new_[11685]_ , \new_[11686]_ , \new_[11687]_ ,
    \new_[11688]_ , \new_[11689]_ , \new_[11690]_ , \new_[11691]_ ,
    \new_[11692]_ , \new_[11693]_ , \new_[11694]_ , \new_[11695]_ ,
    \new_[11696]_ , \new_[11697]_ , \new_[11698]_ , \new_[11699]_ ,
    \new_[11700]_ , \new_[11701]_ , \new_[11702]_ , \new_[11703]_ ,
    \new_[11704]_ , \new_[11705]_ , \new_[11706]_ , \new_[11707]_ ,
    \new_[11708]_ , \new_[11709]_ , \new_[11710]_ , \new_[11711]_ ,
    \new_[11712]_ , \new_[11713]_ , \new_[11714]_ , \new_[11715]_ ,
    \new_[11716]_ , \new_[11718]_ , \new_[11719]_ , \new_[11720]_ ,
    \new_[11721]_ , \new_[11722]_ , \new_[11723]_ , \new_[11724]_ ,
    \new_[11725]_ , \new_[11727]_ , \new_[11728]_ , \new_[11729]_ ,
    \new_[11730]_ , \new_[11731]_ , \new_[11732]_ , \new_[11733]_ ,
    \new_[11734]_ , \new_[11735]_ , \new_[11736]_ , \new_[11737]_ ,
    \new_[11738]_ , \new_[11739]_ , \new_[11740]_ , \new_[11741]_ ,
    \new_[11742]_ , \new_[11743]_ , \new_[11744]_ , \new_[11745]_ ,
    \new_[11746]_ , \new_[11747]_ , \new_[11748]_ , \new_[11749]_ ,
    \new_[11751]_ , \new_[11752]_ , \new_[11753]_ , \new_[11754]_ ,
    \new_[11755]_ , \new_[11756]_ , \new_[11757]_ , \new_[11758]_ ,
    \new_[11759]_ , \new_[11760]_ , \new_[11761]_ , \new_[11762]_ ,
    \new_[11763]_ , \new_[11764]_ , \new_[11765]_ , \new_[11766]_ ,
    \new_[11767]_ , \new_[11768]_ , \new_[11769]_ , \new_[11770]_ ,
    \new_[11771]_ , \new_[11773]_ , \new_[11774]_ , \new_[11775]_ ,
    \new_[11776]_ , \new_[11777]_ , \new_[11778]_ , \new_[11779]_ ,
    \new_[11780]_ , \new_[11781]_ , \new_[11783]_ , \new_[11784]_ ,
    \new_[11785]_ , \new_[11786]_ , \new_[11787]_ , \new_[11788]_ ,
    \new_[11789]_ , \new_[11790]_ , \new_[11791]_ , \new_[11792]_ ,
    \new_[11793]_ , \new_[11794]_ , \new_[11795]_ , \new_[11796]_ ,
    \new_[11797]_ , \new_[11798]_ , \new_[11799]_ , \new_[11800]_ ,
    \new_[11801]_ , \new_[11802]_ , \new_[11803]_ , \new_[11804]_ ,
    \new_[11805]_ , \new_[11806]_ , \new_[11807]_ , \new_[11808]_ ,
    \new_[11809]_ , \new_[11810]_ , \new_[11811]_ , \new_[11812]_ ,
    \new_[11813]_ , \new_[11814]_ , \new_[11815]_ , \new_[11816]_ ,
    \new_[11817]_ , \new_[11818]_ , \new_[11819]_ , \new_[11820]_ ,
    \new_[11821]_ , \new_[11822]_ , \new_[11823]_ , \new_[11824]_ ,
    \new_[11825]_ , \new_[11826]_ , \new_[11827]_ , \new_[11828]_ ,
    \new_[11829]_ , \new_[11830]_ , \new_[11831]_ , \new_[11832]_ ,
    \new_[11833]_ , \new_[11834]_ , \new_[11835]_ , \new_[11836]_ ,
    \new_[11837]_ , \new_[11838]_ , \new_[11839]_ , \new_[11840]_ ,
    \new_[11841]_ , \new_[11842]_ , \new_[11843]_ , \new_[11844]_ ,
    \new_[11845]_ , \new_[11846]_ , \new_[11847]_ , \new_[11848]_ ,
    \new_[11849]_ , \new_[11850]_ , \new_[11851]_ , \new_[11852]_ ,
    \new_[11853]_ , \new_[11854]_ , \new_[11855]_ , \new_[11856]_ ,
    \new_[11857]_ , \new_[11858]_ , \new_[11859]_ , \new_[11860]_ ,
    \new_[11861]_ , \new_[11862]_ , \new_[11863]_ , \new_[11864]_ ,
    \new_[11865]_ , \new_[11866]_ , \new_[11867]_ , \new_[11868]_ ,
    \new_[11869]_ , \new_[11870]_ , \new_[11871]_ , \new_[11872]_ ,
    \new_[11873]_ , \new_[11874]_ , \new_[11875]_ , \new_[11876]_ ,
    \new_[11877]_ , \new_[11878]_ , \new_[11879]_ , \new_[11880]_ ,
    \new_[11881]_ , \new_[11883]_ , \new_[11892]_ , \new_[11900]_ ,
    \new_[11906]_ , \new_[11907]_ , \new_[11908]_ , \new_[11909]_ ,
    \new_[11910]_ , \new_[11911]_ , \new_[11912]_ , \new_[11913]_ ,
    \new_[11914]_ , \new_[11915]_ , \new_[11916]_ , \new_[11917]_ ,
    \new_[11918]_ , \new_[11919]_ , \new_[11920]_ , \new_[11921]_ ,
    \new_[11922]_ , \new_[11923]_ , \new_[11924]_ , \new_[11925]_ ,
    \new_[11926]_ , \new_[11927]_ , \new_[11928]_ , \new_[11929]_ ,
    \new_[11930]_ , \new_[11931]_ , \new_[11932]_ , \new_[11933]_ ,
    \new_[11934]_ , \new_[11936]_ , \new_[11937]_ , \new_[11938]_ ,
    \new_[11939]_ , \new_[11940]_ , \new_[11941]_ , \new_[11942]_ ,
    \new_[11943]_ , \new_[11944]_ , \new_[11945]_ , \new_[11946]_ ,
    \new_[11947]_ , \new_[11948]_ , \new_[11949]_ , \new_[11950]_ ,
    \new_[11951]_ , \new_[11952]_ , \new_[11953]_ , \new_[11954]_ ,
    \new_[11955]_ , \new_[11956]_ , \new_[11957]_ , \new_[11958]_ ,
    \new_[11959]_ , \new_[11960]_ , \new_[11961]_ , \new_[11962]_ ,
    \new_[11963]_ , \new_[11964]_ , \new_[11965]_ , \new_[11966]_ ,
    \new_[11967]_ , \new_[11968]_ , \new_[11969]_ , \new_[11970]_ ,
    \new_[11971]_ , \new_[11972]_ , \new_[11973]_ , \new_[11974]_ ,
    \new_[11975]_ , \new_[11976]_ , \new_[11977]_ , \new_[11978]_ ,
    \new_[11979]_ , \new_[11980]_ , \new_[11981]_ , \new_[11982]_ ,
    \new_[11983]_ , \new_[11984]_ , \new_[11985]_ , \new_[11986]_ ,
    \new_[11987]_ , \new_[11988]_ , \new_[11989]_ , \new_[11990]_ ,
    \new_[11991]_ , \new_[11992]_ , \new_[11993]_ , \new_[11994]_ ,
    \new_[11995]_ , \new_[11996]_ , \new_[11997]_ , \new_[11998]_ ,
    \new_[11999]_ , \new_[12000]_ , \new_[12001]_ , \new_[12002]_ ,
    \new_[12003]_ , \new_[12004]_ , \new_[12005]_ , \new_[12006]_ ,
    \new_[12007]_ , \new_[12008]_ , \new_[12009]_ , \new_[12010]_ ,
    \new_[12011]_ , \new_[12012]_ , \new_[12013]_ , \new_[12014]_ ,
    \new_[12015]_ , \new_[12016]_ , \new_[12017]_ , \new_[12018]_ ,
    \new_[12019]_ , \new_[12020]_ , \new_[12021]_ , \new_[12022]_ ,
    \new_[12023]_ , \new_[12024]_ , \new_[12025]_ , \new_[12026]_ ,
    \new_[12027]_ , \new_[12028]_ , \new_[12029]_ , \new_[12030]_ ,
    \new_[12031]_ , \new_[12032]_ , \new_[12033]_ , \new_[12034]_ ,
    \new_[12035]_ , \new_[12036]_ , \new_[12037]_ , \new_[12038]_ ,
    \new_[12039]_ , \new_[12040]_ , \new_[12041]_ , \new_[12042]_ ,
    \new_[12043]_ , \new_[12044]_ , \new_[12045]_ , \new_[12046]_ ,
    \new_[12047]_ , \new_[12048]_ , \new_[12049]_ , \new_[12050]_ ,
    \new_[12051]_ , \new_[12052]_ , \new_[12053]_ , \new_[12054]_ ,
    \new_[12055]_ , \new_[12056]_ , \new_[12057]_ , \new_[12058]_ ,
    \new_[12059]_ , \new_[12061]_ , \new_[12062]_ , \new_[12063]_ ,
    \new_[12064]_ , \new_[12065]_ , \new_[12066]_ , \new_[12067]_ ,
    \new_[12068]_ , \new_[12069]_ , \new_[12070]_ , \new_[12071]_ ,
    \new_[12072]_ , \new_[12073]_ , \new_[12074]_ , \new_[12075]_ ,
    \new_[12076]_ , \new_[12077]_ , \new_[12078]_ , \new_[12079]_ ,
    \new_[12080]_ , \new_[12081]_ , \new_[12082]_ , \new_[12083]_ ,
    \new_[12084]_ , \new_[12085]_ , \new_[12086]_ , \new_[12087]_ ,
    \new_[12088]_ , \new_[12089]_ , \new_[12090]_ , \new_[12091]_ ,
    \new_[12092]_ , \new_[12093]_ , \new_[12094]_ , \new_[12095]_ ,
    \new_[12096]_ , \new_[12097]_ , \new_[12098]_ , \new_[12099]_ ,
    \new_[12100]_ , \new_[12101]_ , \new_[12102]_ , \new_[12103]_ ,
    \new_[12104]_ , \new_[12105]_ , \new_[12106]_ , \new_[12107]_ ,
    \new_[12108]_ , \new_[12109]_ , \new_[12110]_ , \new_[12111]_ ,
    \new_[12112]_ , \new_[12113]_ , \new_[12114]_ , \new_[12115]_ ,
    \new_[12116]_ , \new_[12117]_ , \new_[12118]_ , \new_[12119]_ ,
    \new_[12120]_ , \new_[12121]_ , \new_[12122]_ , \new_[12123]_ ,
    \new_[12124]_ , \new_[12125]_ , \new_[12126]_ , \new_[12127]_ ,
    \new_[12128]_ , \new_[12129]_ , \new_[12130]_ , \new_[12131]_ ,
    \new_[12132]_ , \new_[12133]_ , \new_[12134]_ , \new_[12135]_ ,
    \new_[12136]_ , \new_[12137]_ , \new_[12138]_ , \new_[12139]_ ,
    \new_[12140]_ , \new_[12141]_ , \new_[12142]_ , \new_[12143]_ ,
    \new_[12144]_ , \new_[12145]_ , \new_[12146]_ , \new_[12147]_ ,
    \new_[12148]_ , \new_[12149]_ , \new_[12150]_ , \new_[12151]_ ,
    \new_[12152]_ , \new_[12153]_ , \new_[12154]_ , \new_[12155]_ ,
    \new_[12156]_ , \new_[12158]_ , \new_[12159]_ , \new_[12160]_ ,
    \new_[12161]_ , \new_[12162]_ , \new_[12163]_ , \new_[12164]_ ,
    \new_[12165]_ , \new_[12166]_ , \new_[12167]_ , \new_[12169]_ ,
    \new_[12170]_ , \new_[12171]_ , \new_[12172]_ , \new_[12175]_ ,
    \new_[12176]_ , \new_[12177]_ , \new_[12178]_ , \new_[12179]_ ,
    \new_[12180]_ , \new_[12181]_ , \new_[12182]_ , \new_[12184]_ ,
    \new_[12185]_ , \new_[12186]_ , \new_[12187]_ , \new_[12188]_ ,
    \new_[12189]_ , \new_[12190]_ , \new_[12191]_ , \new_[12193]_ ,
    \new_[12194]_ , \new_[12195]_ , \new_[12196]_ , \new_[12197]_ ,
    \new_[12198]_ , \new_[12199]_ , \new_[12200]_ , \new_[12201]_ ,
    \new_[12204]_ , \new_[12205]_ , \new_[12206]_ , \new_[12208]_ ,
    \new_[12209]_ , \new_[12210]_ , \new_[12211]_ , \new_[12212]_ ,
    \new_[12213]_ , \new_[12214]_ , \new_[12215]_ , \new_[12216]_ ,
    \new_[12217]_ , \new_[12218]_ , \new_[12219]_ , \new_[12220]_ ,
    \new_[12221]_ , \new_[12222]_ , \new_[12223]_ , \new_[12224]_ ,
    \new_[12225]_ , \new_[12226]_ , \new_[12227]_ , \new_[12228]_ ,
    \new_[12229]_ , \new_[12230]_ , \new_[12231]_ , \new_[12232]_ ,
    \new_[12233]_ , \new_[12234]_ , \new_[12236]_ , \new_[12237]_ ,
    \new_[12238]_ , \new_[12240]_ , \new_[12241]_ , \new_[12242]_ ,
    \new_[12243]_ , \new_[12244]_ , \new_[12245]_ , \new_[12246]_ ,
    \new_[12247]_ , \new_[12248]_ , \new_[12249]_ , \new_[12250]_ ,
    \new_[12251]_ , \new_[12252]_ , \new_[12253]_ , \new_[12254]_ ,
    \new_[12255]_ , \new_[12256]_ , \new_[12257]_ , \new_[12258]_ ,
    \new_[12259]_ , \new_[12260]_ , \new_[12261]_ , \new_[12262]_ ,
    \new_[12263]_ , \new_[12264]_ , \new_[12265]_ , \new_[12266]_ ,
    \new_[12267]_ , \new_[12269]_ , \new_[12270]_ , \new_[12271]_ ,
    \new_[12272]_ , \new_[12274]_ , \new_[12275]_ , \new_[12276]_ ,
    \new_[12277]_ , \new_[12278]_ , \new_[12279]_ , \new_[12280]_ ,
    \new_[12281]_ , \new_[12282]_ , \new_[12283]_ , \new_[12284]_ ,
    \new_[12285]_ , \new_[12286]_ , \new_[12287]_ , \new_[12288]_ ,
    \new_[12289]_ , \new_[12290]_ , \new_[12291]_ , \new_[12292]_ ,
    \new_[12293]_ , \new_[12294]_ , \new_[12295]_ , \new_[12296]_ ,
    \new_[12297]_ , \new_[12298]_ , \new_[12299]_ , \new_[12300]_ ,
    \new_[12301]_ , \new_[12302]_ , \new_[12303]_ , \new_[12304]_ ,
    \new_[12305]_ , \new_[12306]_ , \new_[12307]_ , \new_[12308]_ ,
    \new_[12309]_ , \new_[12310]_ , \new_[12311]_ , \new_[12312]_ ,
    \new_[12313]_ , \new_[12314]_ , \new_[12315]_ , \new_[12316]_ ,
    \new_[12317]_ , \new_[12318]_ , \new_[12319]_ , \new_[12320]_ ,
    \new_[12321]_ , \new_[12322]_ , \new_[12323]_ , \new_[12324]_ ,
    \new_[12325]_ , \new_[12326]_ , \new_[12327]_ , \new_[12328]_ ,
    \new_[12329]_ , \new_[12330]_ , \new_[12331]_ , \new_[12332]_ ,
    \new_[12333]_ , \new_[12334]_ , \new_[12335]_ , \new_[12336]_ ,
    \new_[12337]_ , \new_[12338]_ , \new_[12339]_ , \new_[12340]_ ,
    \new_[12341]_ , \new_[12342]_ , \new_[12343]_ , \new_[12344]_ ,
    \new_[12345]_ , \new_[12346]_ , \new_[12347]_ , \new_[12348]_ ,
    \new_[12349]_ , \new_[12350]_ , \new_[12351]_ , \new_[12352]_ ,
    \new_[12353]_ , \new_[12354]_ , \new_[12355]_ , \new_[12356]_ ,
    \new_[12357]_ , \new_[12358]_ , \new_[12359]_ , \new_[12361]_ ,
    \new_[12362]_ , \new_[12363]_ , \new_[12364]_ , \new_[12365]_ ,
    \new_[12366]_ , \new_[12367]_ , \new_[12368]_ , \new_[12369]_ ,
    \new_[12370]_ , \new_[12371]_ , \new_[12372]_ , \new_[12373]_ ,
    \new_[12374]_ , \new_[12375]_ , \new_[12376]_ , \new_[12377]_ ,
    \new_[12378]_ , \new_[12379]_ , \new_[12380]_ , \new_[12381]_ ,
    \new_[12382]_ , \new_[12383]_ , \new_[12384]_ , \new_[12385]_ ,
    \new_[12386]_ , \new_[12387]_ , \new_[12388]_ , \new_[12389]_ ,
    \new_[12390]_ , \new_[12391]_ , \new_[12392]_ , \new_[12393]_ ,
    \new_[12394]_ , \new_[12395]_ , \new_[12396]_ , \new_[12397]_ ,
    \new_[12398]_ , \new_[12399]_ , \new_[12400]_ , \new_[12401]_ ,
    \new_[12402]_ , \new_[12403]_ , \new_[12404]_ , \new_[12405]_ ,
    \new_[12406]_ , \new_[12407]_ , \new_[12408]_ , \new_[12409]_ ,
    \new_[12410]_ , \new_[12411]_ , \new_[12412]_ , \new_[12413]_ ,
    \new_[12414]_ , \new_[12415]_ , \new_[12416]_ , \new_[12417]_ ,
    \new_[12418]_ , \new_[12419]_ , \new_[12420]_ , \new_[12421]_ ,
    \new_[12422]_ , \new_[12423]_ , \new_[12424]_ , \new_[12425]_ ,
    \new_[12426]_ , \new_[12427]_ , \new_[12428]_ , \new_[12429]_ ,
    \new_[12430]_ , \new_[12431]_ , \new_[12433]_ , \new_[12434]_ ,
    \new_[12435]_ , \new_[12436]_ , \new_[12437]_ , \new_[12438]_ ,
    \new_[12439]_ , \new_[12440]_ , \new_[12441]_ , \new_[12442]_ ,
    \new_[12443]_ , \new_[12444]_ , \new_[12445]_ , \new_[12446]_ ,
    \new_[12447]_ , \new_[12448]_ , \new_[12449]_ , \new_[12450]_ ,
    \new_[12451]_ , \new_[12452]_ , \new_[12454]_ , \new_[12455]_ ,
    \new_[12456]_ , \new_[12457]_ , \new_[12458]_ , \new_[12459]_ ,
    \new_[12460]_ , \new_[12461]_ , \new_[12462]_ , \new_[12463]_ ,
    \new_[12464]_ , \new_[12465]_ , \new_[12466]_ , \new_[12467]_ ,
    \new_[12468]_ , \new_[12469]_ , \new_[12470]_ , \new_[12471]_ ,
    \new_[12472]_ , \new_[12473]_ , \new_[12474]_ , \new_[12475]_ ,
    \new_[12476]_ , \new_[12477]_ , \new_[12478]_ , \new_[12479]_ ,
    \new_[12480]_ , \new_[12481]_ , \new_[12482]_ , \new_[12483]_ ,
    \new_[12484]_ , \new_[12485]_ , \new_[12486]_ , \new_[12487]_ ,
    \new_[12488]_ , \new_[12489]_ , \new_[12491]_ , \new_[12492]_ ,
    \new_[12493]_ , \new_[12494]_ , \new_[12495]_ , \new_[12496]_ ,
    \new_[12497]_ , \new_[12498]_ , \new_[12499]_ , \new_[12500]_ ,
    \new_[12501]_ , \new_[12502]_ , \new_[12503]_ , \new_[12504]_ ,
    \new_[12505]_ , \new_[12506]_ , \new_[12507]_ , \new_[12508]_ ,
    \new_[12509]_ , \new_[12510]_ , \new_[12511]_ , \new_[12512]_ ,
    \new_[12513]_ , \new_[12514]_ , \new_[12515]_ , \new_[12516]_ ,
    \new_[12517]_ , \new_[12518]_ , \new_[12519]_ , \new_[12520]_ ,
    \new_[12521]_ , \new_[12522]_ , \new_[12523]_ , \new_[12524]_ ,
    \new_[12525]_ , \new_[12526]_ , \new_[12527]_ , \new_[12528]_ ,
    \new_[12529]_ , \new_[12530]_ , \new_[12531]_ , \new_[12532]_ ,
    \new_[12533]_ , \new_[12534]_ , \new_[12535]_ , \new_[12537]_ ,
    \new_[12538]_ , \new_[12540]_ , \new_[12541]_ , \new_[12542]_ ,
    \new_[12543]_ , \new_[12544]_ , \new_[12545]_ , \new_[12546]_ ,
    \new_[12547]_ , \new_[12548]_ , \new_[12549]_ , \new_[12550]_ ,
    \new_[12551]_ , \new_[12552]_ , \new_[12553]_ , \new_[12554]_ ,
    \new_[12555]_ , \new_[12556]_ , \new_[12557]_ , \new_[12558]_ ,
    \new_[12559]_ , \new_[12560]_ , \new_[12561]_ , \new_[12562]_ ,
    \new_[12563]_ , \new_[12564]_ , \new_[12565]_ , \new_[12566]_ ,
    \new_[12567]_ , \new_[12568]_ , \new_[12569]_ , \new_[12570]_ ,
    \new_[12571]_ , \new_[12572]_ , \new_[12573]_ , \new_[12574]_ ,
    \new_[12575]_ , \new_[12576]_ , \new_[12577]_ , \new_[12578]_ ,
    \new_[12579]_ , \new_[12580]_ , \new_[12581]_ , \new_[12582]_ ,
    \new_[12583]_ , \new_[12584]_ , \new_[12585]_ , \new_[12586]_ ,
    \new_[12587]_ , \new_[12588]_ , \new_[12589]_ , \new_[12590]_ ,
    \new_[12591]_ , \new_[12592]_ , \new_[12593]_ , \new_[12594]_ ,
    \new_[12595]_ , \new_[12596]_ , \new_[12597]_ , \new_[12598]_ ,
    \new_[12599]_ , \new_[12600]_ , \new_[12601]_ , \new_[12602]_ ,
    \new_[12603]_ , \new_[12604]_ , \new_[12605]_ , \new_[12606]_ ,
    \new_[12607]_ , \new_[12608]_ , \new_[12609]_ , \new_[12610]_ ,
    \new_[12611]_ , \new_[12612]_ , \new_[12613]_ , \new_[12614]_ ,
    \new_[12615]_ , \new_[12616]_ , \new_[12617]_ , \new_[12618]_ ,
    \new_[12619]_ , \new_[12620]_ , \new_[12621]_ , \new_[12622]_ ,
    \new_[12623]_ , \new_[12624]_ , \new_[12625]_ , \new_[12626]_ ,
    \new_[12627]_ , \new_[12628]_ , \new_[12629]_ , \new_[12630]_ ,
    \new_[12631]_ , \new_[12632]_ , \new_[12633]_ , \new_[12634]_ ,
    \new_[12635]_ , \new_[12636]_ , \new_[12637]_ , \new_[12638]_ ,
    \new_[12639]_ , \new_[12640]_ , \new_[12641]_ , \new_[12642]_ ,
    \new_[12643]_ , \new_[12644]_ , \new_[12645]_ , \new_[12646]_ ,
    \new_[12647]_ , \new_[12648]_ , \new_[12649]_ , \new_[12650]_ ,
    \new_[12651]_ , \new_[12652]_ , \new_[12653]_ , \new_[12654]_ ,
    \new_[12655]_ , \new_[12656]_ , \new_[12657]_ , \new_[12658]_ ,
    \new_[12659]_ , \new_[12660]_ , \new_[12661]_ , \new_[12662]_ ,
    \new_[12663]_ , \new_[12664]_ , \new_[12665]_ , \new_[12666]_ ,
    \new_[12667]_ , \new_[12668]_ , \new_[12669]_ , \new_[12670]_ ,
    \new_[12671]_ , \new_[12672]_ , \new_[12673]_ , \new_[12674]_ ,
    \new_[12675]_ , \new_[12676]_ , \new_[12677]_ , \new_[12678]_ ,
    \new_[12679]_ , \new_[12680]_ , \new_[12681]_ , \new_[12682]_ ,
    \new_[12683]_ , \new_[12684]_ , \new_[12685]_ , \new_[12686]_ ,
    \new_[12687]_ , \new_[12688]_ , \new_[12689]_ , \new_[12690]_ ,
    \new_[12691]_ , \new_[12692]_ , \new_[12693]_ , \new_[12694]_ ,
    \new_[12695]_ , \new_[12696]_ , \new_[12697]_ , \new_[12698]_ ,
    \new_[12699]_ , \new_[12700]_ , \new_[12701]_ , \new_[12702]_ ,
    \new_[12703]_ , \new_[12704]_ , \new_[12705]_ , \new_[12706]_ ,
    \new_[12707]_ , \new_[12708]_ , \new_[12709]_ , \new_[12710]_ ,
    \new_[12711]_ , \new_[12712]_ , \new_[12713]_ , \new_[12714]_ ,
    \new_[12715]_ , \new_[12716]_ , \new_[12717]_ , \new_[12718]_ ,
    \new_[12719]_ , \new_[12720]_ , \new_[12721]_ , \new_[12722]_ ,
    \new_[12723]_ , \new_[12724]_ , \new_[12725]_ , \new_[12726]_ ,
    \new_[12727]_ , \new_[12728]_ , \new_[12729]_ , \new_[12730]_ ,
    \new_[12731]_ , \new_[12732]_ , \new_[12733]_ , \new_[12734]_ ,
    \new_[12735]_ , \new_[12736]_ , \new_[12737]_ , \new_[12738]_ ,
    \new_[12739]_ , \new_[12740]_ , \new_[12741]_ , \new_[12742]_ ,
    \new_[12743]_ , \new_[12744]_ , \new_[12745]_ , \new_[12746]_ ,
    \new_[12747]_ , \new_[12748]_ , \new_[12749]_ , \new_[12750]_ ,
    \new_[12751]_ , \new_[12752]_ , \new_[12753]_ , \new_[12754]_ ,
    \new_[12755]_ , \new_[12756]_ , \new_[12757]_ , \new_[12758]_ ,
    \new_[12759]_ , \new_[12760]_ , \new_[12761]_ , \new_[12762]_ ,
    \new_[12763]_ , \new_[12764]_ , \new_[12765]_ , \new_[12766]_ ,
    \new_[12767]_ , \new_[12768]_ , \new_[12769]_ , \new_[12770]_ ,
    \new_[12771]_ , \new_[12772]_ , \new_[12773]_ , \new_[12774]_ ,
    \new_[12775]_ , \new_[12776]_ , \new_[12777]_ , \new_[12778]_ ,
    \new_[12779]_ , \new_[12780]_ , \new_[12781]_ , \new_[12782]_ ,
    \new_[12783]_ , \new_[12784]_ , \new_[12785]_ , \new_[12786]_ ,
    \new_[12787]_ , \new_[12788]_ , \new_[12789]_ , \new_[12790]_ ,
    \new_[12791]_ , \new_[12792]_ , \new_[12793]_ , \new_[12794]_ ,
    \new_[12795]_ , \new_[12796]_ , \new_[12797]_ , \new_[12798]_ ,
    \new_[12800]_ , \new_[12801]_ , \new_[12802]_ , \new_[12803]_ ,
    \new_[12804]_ , \new_[12805]_ , \new_[12806]_ , \new_[12807]_ ,
    \new_[12808]_ , \new_[12809]_ , \new_[12810]_ , \new_[12811]_ ,
    \new_[12812]_ , \new_[12813]_ , \new_[12814]_ , \new_[12815]_ ,
    \new_[12816]_ , \new_[12817]_ , \new_[12818]_ , \new_[12819]_ ,
    \new_[12820]_ , \new_[12821]_ , \new_[12822]_ , \new_[12823]_ ,
    \new_[12824]_ , \new_[12825]_ , \new_[12826]_ , \new_[12827]_ ,
    \new_[12828]_ , \new_[12829]_ , \new_[12830]_ , \new_[12831]_ ,
    \new_[12832]_ , \new_[12833]_ , \new_[12834]_ , \new_[12835]_ ,
    \new_[12836]_ , \new_[12837]_ , \new_[12838]_ , \new_[12839]_ ,
    \new_[12840]_ , \new_[12841]_ , \new_[12842]_ , \new_[12843]_ ,
    \new_[12844]_ , \new_[12845]_ , \new_[12846]_ , \new_[12847]_ ,
    \new_[12848]_ , \new_[12849]_ , \new_[12850]_ , \new_[12851]_ ,
    \new_[12853]_ , \new_[12854]_ , \new_[12855]_ , \new_[12856]_ ,
    \new_[12857]_ , \new_[12858]_ , \new_[12859]_ , \new_[12860]_ ,
    \new_[12861]_ , \new_[12862]_ , \new_[12863]_ , \new_[12864]_ ,
    \new_[12865]_ , \new_[12866]_ , \new_[12867]_ , \new_[12868]_ ,
    \new_[12869]_ , \new_[12870]_ , \new_[12871]_ , \new_[12872]_ ,
    \new_[12873]_ , \new_[12874]_ , \new_[12875]_ , \new_[12876]_ ,
    \new_[12877]_ , \new_[12878]_ , \new_[12879]_ , \new_[12880]_ ,
    \new_[12881]_ , \new_[12882]_ , \new_[12883]_ , \new_[12884]_ ,
    \new_[12885]_ , \new_[12886]_ , \new_[12887]_ , \new_[12888]_ ,
    \new_[12889]_ , \new_[12890]_ , \new_[12891]_ , \new_[12892]_ ,
    \new_[12894]_ , \new_[12895]_ , \new_[12896]_ , \new_[12897]_ ,
    \new_[12898]_ , \new_[12899]_ , \new_[12900]_ , \new_[12901]_ ,
    \new_[12902]_ , \new_[12903]_ , \new_[12904]_ , \new_[12905]_ ,
    \new_[12906]_ , \new_[12908]_ , \new_[12909]_ , \new_[12910]_ ,
    \new_[12911]_ , \new_[12912]_ , \new_[12913]_ , \new_[12914]_ ,
    \new_[12916]_ , \new_[12918]_ , \new_[12919]_ , \new_[12920]_ ,
    \new_[12921]_ , \new_[12922]_ , \new_[12923]_ , \new_[12924]_ ,
    \new_[12925]_ , \new_[12926]_ , \new_[12927]_ , \new_[12928]_ ,
    \new_[12929]_ , \new_[12931]_ , \new_[12932]_ , \new_[12933]_ ,
    \new_[12934]_ , \new_[12935]_ , \new_[12936]_ , \new_[12937]_ ,
    \new_[12938]_ , \new_[12939]_ , \new_[12940]_ , \new_[12941]_ ,
    \new_[12942]_ , \new_[12943]_ , \new_[12944]_ , \new_[12945]_ ,
    \new_[12946]_ , \new_[12947]_ , \new_[12948]_ , \new_[12949]_ ,
    \new_[12950]_ , \new_[12951]_ , \new_[12952]_ , \new_[12953]_ ,
    \new_[12954]_ , \new_[12955]_ , \new_[12956]_ , \new_[12958]_ ,
    \new_[12959]_ , \new_[12960]_ , \new_[12961]_ , \new_[12962]_ ,
    \new_[12963]_ , \new_[12964]_ , \new_[12965]_ , \new_[12966]_ ,
    \new_[12967]_ , \new_[12968]_ , \new_[12969]_ , \new_[12970]_ ,
    \new_[12971]_ , \new_[12972]_ , \new_[12973]_ , \new_[12974]_ ,
    \new_[12975]_ , \new_[12976]_ , \new_[12977]_ , \new_[12978]_ ,
    \new_[12979]_ , \new_[12980]_ , \new_[12981]_ , \new_[12982]_ ,
    \new_[12983]_ , \new_[12984]_ , \new_[12985]_ , \new_[12986]_ ,
    \new_[12987]_ , \new_[12988]_ , \new_[12989]_ , \new_[12990]_ ,
    \new_[12991]_ , \new_[12992]_ , \new_[12993]_ , \new_[12994]_ ,
    \new_[12995]_ , \new_[12996]_ , \new_[12997]_ , \new_[12998]_ ,
    \new_[12999]_ , \new_[13000]_ , \new_[13001]_ , \new_[13002]_ ,
    \new_[13003]_ , \new_[13004]_ , \new_[13005]_ , \new_[13006]_ ,
    \new_[13007]_ , \new_[13008]_ , \new_[13009]_ , \new_[13010]_ ,
    \new_[13011]_ , \new_[13012]_ , \new_[13013]_ , \new_[13014]_ ,
    \new_[13015]_ , \new_[13016]_ , \new_[13017]_ , \new_[13018]_ ,
    \new_[13019]_ , \new_[13020]_ , \new_[13021]_ , \new_[13022]_ ,
    \new_[13023]_ , \new_[13024]_ , \new_[13025]_ , \new_[13026]_ ,
    \new_[13027]_ , \new_[13028]_ , \new_[13029]_ , \new_[13030]_ ,
    \new_[13031]_ , \new_[13032]_ , \new_[13033]_ , \new_[13034]_ ,
    \new_[13035]_ , \new_[13036]_ , \new_[13037]_ , \new_[13038]_ ,
    \new_[13039]_ , \new_[13040]_ , \new_[13041]_ , \new_[13042]_ ,
    \new_[13043]_ , \new_[13044]_ , \new_[13045]_ , \new_[13046]_ ,
    \new_[13047]_ , \new_[13048]_ , \new_[13049]_ , \new_[13050]_ ,
    \new_[13051]_ , \new_[13052]_ , \new_[13053]_ , \new_[13054]_ ,
    \new_[13055]_ , \new_[13056]_ , \new_[13057]_ , \new_[13058]_ ,
    \new_[13059]_ , \new_[13060]_ , \new_[13061]_ , \new_[13062]_ ,
    \new_[13063]_ , \new_[13064]_ , \new_[13065]_ , \new_[13066]_ ,
    \new_[13067]_ , \new_[13068]_ , \new_[13069]_ , \new_[13070]_ ,
    \new_[13071]_ , \new_[13072]_ , \new_[13073]_ , \new_[13074]_ ,
    \new_[13075]_ , \new_[13076]_ , \new_[13077]_ , \new_[13078]_ ,
    \new_[13079]_ , \new_[13080]_ , \new_[13081]_ , \new_[13082]_ ,
    \new_[13083]_ , \new_[13084]_ , \new_[13085]_ , \new_[13086]_ ,
    \new_[13087]_ , \new_[13088]_ , \new_[13089]_ , \new_[13090]_ ,
    \new_[13091]_ , \new_[13092]_ , \new_[13093]_ , \new_[13094]_ ,
    \new_[13095]_ , \new_[13096]_ , \new_[13097]_ , \new_[13098]_ ,
    \new_[13099]_ , \new_[13100]_ , \new_[13101]_ , \new_[13102]_ ,
    \new_[13103]_ , \new_[13104]_ , \new_[13105]_ , \new_[13106]_ ,
    \new_[13107]_ , \new_[13108]_ , \new_[13109]_ , \new_[13110]_ ,
    \new_[13111]_ , \new_[13112]_ , \new_[13113]_ , \new_[13114]_ ,
    \new_[13115]_ , \new_[13116]_ , \new_[13117]_ , \new_[13118]_ ,
    \new_[13119]_ , \new_[13120]_ , \new_[13121]_ , \new_[13122]_ ,
    \new_[13123]_ , \new_[13124]_ , \new_[13125]_ , \new_[13126]_ ,
    \new_[13127]_ , \new_[13128]_ , \new_[13129]_ , \new_[13130]_ ,
    \new_[13131]_ , \new_[13132]_ , \new_[13133]_ , \new_[13134]_ ,
    \new_[13135]_ , \new_[13136]_ , \new_[13137]_ , \new_[13138]_ ,
    \new_[13139]_ , \new_[13140]_ , \new_[13141]_ , \new_[13142]_ ,
    \new_[13143]_ , \new_[13144]_ , \new_[13145]_ , \new_[13147]_ ,
    \new_[13148]_ , \new_[13149]_ , \new_[13150]_ , \new_[13151]_ ,
    \new_[13152]_ , \new_[13153]_ , \new_[13154]_ , \new_[13155]_ ,
    \new_[13156]_ , \new_[13157]_ , \new_[13158]_ , \new_[13159]_ ,
    \new_[13160]_ , \new_[13161]_ , \new_[13162]_ , \new_[13163]_ ,
    \new_[13164]_ , \new_[13165]_ , \new_[13166]_ , \new_[13167]_ ,
    \new_[13168]_ , \new_[13169]_ , \new_[13170]_ , \new_[13171]_ ,
    \new_[13172]_ , \new_[13173]_ , \new_[13174]_ , \new_[13177]_ ,
    \new_[13178]_ , \new_[13179]_ , \new_[13180]_ , \new_[13181]_ ,
    \new_[13182]_ , \new_[13183]_ , \new_[13184]_ , \new_[13185]_ ,
    \new_[13186]_ , \new_[13187]_ , \new_[13188]_ , \new_[13189]_ ,
    \new_[13190]_ , \new_[13191]_ , \new_[13192]_ , \new_[13193]_ ,
    \new_[13194]_ , \new_[13196]_ , \new_[13197]_ , \new_[13198]_ ,
    \new_[13199]_ , \new_[13200]_ , \new_[13201]_ , \new_[13202]_ ,
    \new_[13203]_ , \new_[13204]_ , \new_[13205]_ , \new_[13206]_ ,
    \new_[13207]_ , \new_[13208]_ , \new_[13209]_ , \new_[13211]_ ,
    \new_[13212]_ , \new_[13213]_ , \new_[13214]_ , \new_[13215]_ ,
    \new_[13216]_ , \new_[13217]_ , \new_[13218]_ , \new_[13219]_ ,
    \new_[13220]_ , \new_[13221]_ , \new_[13222]_ , \new_[13223]_ ,
    \new_[13224]_ , \new_[13225]_ , \new_[13226]_ , \new_[13227]_ ,
    \new_[13228]_ , \new_[13229]_ , \new_[13230]_ , \new_[13231]_ ,
    \new_[13232]_ , \new_[13233]_ , \new_[13234]_ , \new_[13235]_ ,
    \new_[13236]_ , \new_[13237]_ , \new_[13238]_ , \new_[13239]_ ,
    \new_[13240]_ , \new_[13241]_ , \new_[13242]_ , \new_[13243]_ ,
    \new_[13244]_ , \new_[13245]_ , \new_[13246]_ , \new_[13247]_ ,
    \new_[13248]_ , \new_[13249]_ , \new_[13250]_ , \new_[13251]_ ,
    \new_[13252]_ , \new_[13253]_ , \new_[13254]_ , \new_[13255]_ ,
    \new_[13256]_ , \new_[13257]_ , \new_[13258]_ , \new_[13259]_ ,
    \new_[13260]_ , \new_[13261]_ , \new_[13262]_ , \new_[13263]_ ,
    \new_[13264]_ , \new_[13265]_ , \new_[13267]_ , \new_[13268]_ ,
    \new_[13270]_ , \new_[13271]_ , \new_[13272]_ , \new_[13274]_ ,
    \new_[13275]_ , \new_[13276]_ , \new_[13277]_ , \new_[13278]_ ,
    \new_[13279]_ , \new_[13280]_ , \new_[13281]_ , \new_[13282]_ ,
    \new_[13283]_ , \new_[13284]_ , \new_[13285]_ , \new_[13286]_ ,
    \new_[13287]_ , \new_[13288]_ , \new_[13289]_ , \new_[13290]_ ,
    \new_[13291]_ , \new_[13292]_ , \new_[13293]_ , \new_[13294]_ ,
    \new_[13296]_ , \new_[13297]_ , \new_[13298]_ , \new_[13299]_ ,
    \new_[13300]_ , \new_[13301]_ , \new_[13302]_ , \new_[13303]_ ,
    \new_[13304]_ , \new_[13305]_ , \new_[13306]_ , \new_[13307]_ ,
    \new_[13308]_ , \new_[13309]_ , \new_[13310]_ , \new_[13311]_ ,
    \new_[13312]_ , \new_[13313]_ , \new_[13314]_ , \new_[13315]_ ,
    \new_[13316]_ , \new_[13317]_ , \new_[13318]_ , \new_[13319]_ ,
    \new_[13320]_ , \new_[13321]_ , \new_[13322]_ , \new_[13323]_ ,
    \new_[13324]_ , \new_[13325]_ , \new_[13326]_ , \new_[13327]_ ,
    \new_[13328]_ , \new_[13330]_ , \new_[13331]_ , \new_[13333]_ ,
    \new_[13334]_ , \new_[13335]_ , \new_[13336]_ , \new_[13337]_ ,
    \new_[13339]_ , \new_[13340]_ , \new_[13341]_ , \new_[13342]_ ,
    \new_[13343]_ , \new_[13344]_ , \new_[13345]_ , \new_[13346]_ ,
    \new_[13347]_ , \new_[13348]_ , \new_[13349]_ , \new_[13350]_ ,
    \new_[13351]_ , \new_[13352]_ , \new_[13353]_ , \new_[13355]_ ,
    \new_[13356]_ , \new_[13357]_ , \new_[13358]_ , \new_[13359]_ ,
    \new_[13360]_ , \new_[13361]_ , \new_[13362]_ , \new_[13363]_ ,
    \new_[13364]_ , \new_[13365]_ , \new_[13366]_ , \new_[13367]_ ,
    \new_[13368]_ , \new_[13369]_ , \new_[13370]_ , \new_[13371]_ ,
    \new_[13372]_ , \new_[13373]_ , \new_[13374]_ , \new_[13375]_ ,
    \new_[13376]_ , \new_[13377]_ , \new_[13378]_ , \new_[13379]_ ,
    \new_[13380]_ , \new_[13381]_ , \new_[13382]_ , \new_[13383]_ ,
    \new_[13384]_ , \new_[13385]_ , \new_[13386]_ , \new_[13387]_ ,
    \new_[13388]_ , \new_[13389]_ , \new_[13390]_ , \new_[13391]_ ,
    \new_[13392]_ , \new_[13393]_ , \new_[13394]_ , \new_[13395]_ ,
    \new_[13396]_ , \new_[13397]_ , \new_[13398]_ , \new_[13399]_ ,
    \new_[13400]_ , \new_[13403]_ , \new_[13405]_ , \new_[13406]_ ,
    \new_[13407]_ , \new_[13408]_ , \new_[13409]_ , \new_[13410]_ ,
    \new_[13411]_ , \new_[13412]_ , \new_[13413]_ , \new_[13415]_ ,
    \new_[13416]_ , \new_[13417]_ , \new_[13418]_ , \new_[13419]_ ,
    \new_[13420]_ , \new_[13421]_ , \new_[13422]_ , \new_[13423]_ ,
    \new_[13424]_ , \new_[13426]_ , \new_[13427]_ , \new_[13428]_ ,
    \new_[13429]_ , \new_[13430]_ , \new_[13431]_ , \new_[13432]_ ,
    \new_[13433]_ , \new_[13434]_ , \new_[13435]_ , \new_[13436]_ ,
    \new_[13437]_ , \new_[13438]_ , \new_[13440]_ , \new_[13441]_ ,
    \new_[13442]_ , \new_[13443]_ , \new_[13444]_ , \new_[13445]_ ,
    \new_[13446]_ , \new_[13447]_ , \new_[13448]_ , \new_[13449]_ ,
    \new_[13450]_ , \new_[13451]_ , \new_[13452]_ , \new_[13453]_ ,
    \new_[13454]_ , \new_[13455]_ , \new_[13456]_ , \new_[13457]_ ,
    \new_[13458]_ , \new_[13459]_ , \new_[13460]_ , \new_[13461]_ ,
    \new_[13462]_ , \new_[13463]_ , \new_[13464]_ , \new_[13465]_ ,
    \new_[13466]_ , \new_[13468]_ , \new_[13469]_ , \new_[13470]_ ,
    \new_[13471]_ , \new_[13472]_ , \new_[13473]_ , \new_[13474]_ ,
    \new_[13476]_ , \new_[13477]_ , \new_[13478]_ , \new_[13479]_ ,
    \new_[13480]_ , \new_[13481]_ , \new_[13482]_ , \new_[13483]_ ,
    \new_[13485]_ , \new_[13486]_ , \new_[13488]_ , \new_[13489]_ ,
    \new_[13490]_ , \new_[13491]_ , \new_[13492]_ , \new_[13493]_ ,
    \new_[13494]_ , \new_[13495]_ , \new_[13496]_ , \new_[13497]_ ,
    \new_[13498]_ , \new_[13499]_ , \new_[13500]_ , \new_[13501]_ ,
    \new_[13502]_ , \new_[13503]_ , \new_[13504]_ , \new_[13505]_ ,
    \new_[13506]_ , \new_[13507]_ , \new_[13508]_ , \new_[13509]_ ,
    \new_[13511]_ , \new_[13512]_ , \new_[13513]_ , \new_[13514]_ ,
    \new_[13515]_ , \new_[13516]_ , \new_[13517]_ , \new_[13518]_ ,
    \new_[13519]_ , \new_[13520]_ , \new_[13521]_ , \new_[13522]_ ,
    \new_[13523]_ , \new_[13524]_ , \new_[13525]_ , \new_[13526]_ ,
    \new_[13527]_ , \new_[13528]_ , \new_[13529]_ , \new_[13530]_ ,
    \new_[13531]_ , \new_[13532]_ , \new_[13533]_ , \new_[13534]_ ,
    \new_[13535]_ , \new_[13536]_ , \new_[13537]_ , \new_[13538]_ ,
    \new_[13539]_ , \new_[13540]_ , \new_[13541]_ , \new_[13542]_ ,
    \new_[13543]_ , \new_[13545]_ , \new_[13546]_ , \new_[13547]_ ,
    \new_[13548]_ , \new_[13549]_ , \new_[13550]_ , \new_[13551]_ ,
    \new_[13552]_ , \new_[13553]_ , \new_[13554]_ , \new_[13555]_ ,
    \new_[13556]_ , \new_[13557]_ , \new_[13558]_ , \new_[13559]_ ,
    \new_[13560]_ , \new_[13561]_ , \new_[13562]_ , \new_[13563]_ ,
    \new_[13564]_ , \new_[13565]_ , \new_[13566]_ , \new_[13567]_ ,
    \new_[13568]_ , \new_[13569]_ , \new_[13570]_ , \new_[13571]_ ,
    \new_[13572]_ , \new_[13573]_ , \new_[13574]_ , \new_[13575]_ ,
    \new_[13576]_ , \new_[13578]_ , \new_[13579]_ , \new_[13580]_ ,
    \new_[13581]_ , \new_[13582]_ , \new_[13583]_ , \new_[13584]_ ,
    \new_[13585]_ , \new_[13586]_ , \new_[13587]_ , \new_[13588]_ ,
    \new_[13589]_ , \new_[13590]_ , \new_[13592]_ , \new_[13593]_ ,
    \new_[13594]_ , \new_[13595]_ , \new_[13596]_ , \new_[13597]_ ,
    \new_[13598]_ , \new_[13599]_ , \new_[13600]_ , \new_[13601]_ ,
    \new_[13602]_ , \new_[13603]_ , \new_[13605]_ , \new_[13606]_ ,
    \new_[13607]_ , \new_[13608]_ , \new_[13609]_ , \new_[13610]_ ,
    \new_[13611]_ , \new_[13612]_ , \new_[13613]_ , \new_[13614]_ ,
    \new_[13615]_ , \new_[13616]_ , \new_[13617]_ , \new_[13618]_ ,
    \new_[13619]_ , \new_[13620]_ , \new_[13621]_ , \new_[13622]_ ,
    \new_[13623]_ , \new_[13624]_ , \new_[13625]_ , \new_[13626]_ ,
    \new_[13627]_ , \new_[13628]_ , \new_[13629]_ , \new_[13630]_ ,
    \new_[13631]_ , \new_[13632]_ , \new_[13633]_ , \new_[13634]_ ,
    \new_[13635]_ , \new_[13637]_ , \new_[13638]_ , \new_[13639]_ ,
    \new_[13640]_ , \new_[13641]_ , \new_[13642]_ , \new_[13643]_ ,
    \new_[13644]_ , \new_[13645]_ , \new_[13646]_ , \new_[13647]_ ,
    \new_[13648]_ , \new_[13649]_ , \new_[13650]_ , \new_[13651]_ ,
    \new_[13652]_ , \new_[13653]_ , \new_[13654]_ , \new_[13655]_ ,
    \new_[13656]_ , \new_[13657]_ , \new_[13658]_ , \new_[13659]_ ,
    \new_[13660]_ , \new_[13661]_ , \new_[13662]_ , \new_[13663]_ ,
    \new_[13664]_ , \new_[13665]_ , \new_[13666]_ , \new_[13667]_ ,
    \new_[13668]_ , \new_[13669]_ , \new_[13670]_ , \new_[13671]_ ,
    \new_[13672]_ , \new_[13673]_ , \new_[13674]_ , \new_[13675]_ ,
    \new_[13676]_ , \new_[13677]_ , \new_[13678]_ , \new_[13679]_ ,
    \new_[13680]_ , \new_[13681]_ , \new_[13682]_ , \new_[13683]_ ,
    \new_[13684]_ , \new_[13685]_ , \new_[13686]_ , \new_[13687]_ ,
    \new_[13688]_ , \new_[13689]_ , \new_[13690]_ , \new_[13691]_ ,
    \new_[13692]_ , \new_[13693]_ , \new_[13694]_ , \new_[13695]_ ,
    \new_[13696]_ , \new_[13697]_ , \new_[13698]_ , \new_[13699]_ ,
    \new_[13700]_ , \new_[13701]_ , \new_[13702]_ , \new_[13703]_ ,
    \new_[13704]_ , \new_[13705]_ , \new_[13706]_ , \new_[13707]_ ,
    \new_[13708]_ , \new_[13709]_ , \new_[13710]_ , \new_[13711]_ ,
    \new_[13712]_ , \new_[13713]_ , \new_[13714]_ , \new_[13715]_ ,
    \new_[13716]_ , \new_[13717]_ , \new_[13718]_ , \new_[13719]_ ,
    \new_[13720]_ , \new_[13721]_ , \new_[13722]_ , \new_[13723]_ ,
    \new_[13724]_ , \new_[13725]_ , \new_[13726]_ , \new_[13727]_ ,
    \new_[13728]_ , \new_[13729]_ , \new_[13730]_ , \new_[13731]_ ,
    \new_[13732]_ , \new_[13733]_ , \new_[13734]_ , \new_[13735]_ ,
    \new_[13736]_ , \new_[13737]_ , \new_[13738]_ , \new_[13739]_ ,
    \new_[13740]_ , \new_[13741]_ , \new_[13742]_ , \new_[13743]_ ,
    \new_[13744]_ , \new_[13745]_ , \new_[13746]_ , \new_[13747]_ ,
    \new_[13748]_ , \new_[13749]_ , \new_[13750]_ , \new_[13751]_ ,
    \new_[13752]_ , \new_[13753]_ , \new_[13754]_ , \new_[13755]_ ,
    \new_[13756]_ , \new_[13757]_ , \new_[13758]_ , \new_[13759]_ ,
    \new_[13760]_ , \new_[13761]_ , \new_[13762]_ , \new_[13763]_ ,
    \new_[13764]_ , \new_[13765]_ , \new_[13766]_ , \new_[13767]_ ,
    \new_[13768]_ , \new_[13769]_ , \new_[13770]_ , \new_[13771]_ ,
    \new_[13772]_ , \new_[13773]_ , \new_[13774]_ , \new_[13775]_ ,
    \new_[13776]_ , \new_[13777]_ , \new_[13778]_ , \new_[13779]_ ,
    \new_[13780]_ , \new_[13782]_ , \new_[13783]_ , \new_[13784]_ ,
    \new_[13785]_ , \new_[13786]_ , \new_[13787]_ , \new_[13788]_ ,
    \new_[13789]_ , \new_[13790]_ , \new_[13791]_ , \new_[13792]_ ,
    \new_[13793]_ , \new_[13794]_ , \new_[13795]_ , \new_[13796]_ ,
    \new_[13797]_ , \new_[13798]_ , \new_[13799]_ , \new_[13800]_ ,
    \new_[13801]_ , \new_[13802]_ , \new_[13803]_ , \new_[13804]_ ,
    \new_[13805]_ , \new_[13806]_ , \new_[13807]_ , \new_[13808]_ ,
    \new_[13809]_ , \new_[13810]_ , \new_[13811]_ , \new_[13812]_ ,
    \new_[13813]_ , \new_[13814]_ , \new_[13815]_ , \new_[13816]_ ,
    \new_[13817]_ , \new_[13818]_ , \new_[13819]_ , \new_[13820]_ ,
    \new_[13821]_ , \new_[13822]_ , \new_[13823]_ , \new_[13824]_ ,
    \new_[13825]_ , \new_[13826]_ , \new_[13827]_ , \new_[13828]_ ,
    \new_[13829]_ , \new_[13830]_ , \new_[13831]_ , \new_[13833]_ ,
    \new_[13834]_ , \new_[13835]_ , \new_[13836]_ , \new_[13837]_ ,
    \new_[13838]_ , \new_[13839]_ , \new_[13840]_ , \new_[13841]_ ,
    \new_[13842]_ , \new_[13843]_ , \new_[13844]_ , \new_[13845]_ ,
    \new_[13846]_ , \new_[13847]_ , \new_[13848]_ , \new_[13849]_ ,
    \new_[13850]_ , \new_[13851]_ , \new_[13852]_ , \new_[13853]_ ,
    \new_[13854]_ , \new_[13855]_ , \new_[13856]_ , \new_[13857]_ ,
    \new_[13858]_ , \new_[13859]_ , \new_[13860]_ , \new_[13861]_ ,
    \new_[13862]_ , \new_[13863]_ , \new_[13864]_ , \new_[13865]_ ,
    \new_[13866]_ , \new_[13867]_ , \new_[13868]_ , \new_[13869]_ ,
    \new_[13870]_ , \new_[13871]_ , \new_[13872]_ , \new_[13873]_ ,
    \new_[13874]_ , \new_[13875]_ , \new_[13876]_ , \new_[13877]_ ,
    \new_[13878]_ , \new_[13879]_ , \new_[13880]_ , \new_[13881]_ ,
    \new_[13882]_ , \new_[13883]_ , \new_[13884]_ , \new_[13885]_ ,
    \new_[13886]_ , \new_[13887]_ , \new_[13888]_ , \new_[13889]_ ,
    \new_[13890]_ , \new_[13891]_ , \new_[13892]_ , \new_[13893]_ ,
    \new_[13894]_ , \new_[13895]_ , \new_[13896]_ , \new_[13897]_ ,
    \new_[13898]_ , \new_[13899]_ , \new_[13900]_ , \new_[13901]_ ,
    \new_[13902]_ , \new_[13903]_ , \new_[13904]_ , \new_[13905]_ ,
    \new_[13906]_ , \new_[13907]_ , \new_[13908]_ , \new_[13909]_ ,
    \new_[13910]_ , \new_[13911]_ , \new_[13912]_ , \new_[13913]_ ,
    \new_[13914]_ , \new_[13915]_ , \new_[13916]_ , \new_[13917]_ ,
    \new_[13918]_ , \new_[13919]_ , \new_[13920]_ , \new_[13921]_ ,
    \new_[13922]_ , \new_[13923]_ , \new_[13924]_ , \new_[13925]_ ,
    \new_[13926]_ , \new_[13927]_ , \new_[13928]_ , \new_[13929]_ ,
    \new_[13930]_ , \new_[13931]_ , \new_[13932]_ , \new_[13933]_ ,
    \new_[13934]_ , \new_[13935]_ , \new_[13936]_ , \new_[13937]_ ,
    \new_[13938]_ , \new_[13939]_ , \new_[13940]_ , \new_[13941]_ ,
    \new_[13942]_ , \new_[13943]_ , \new_[13944]_ , \new_[13945]_ ,
    \new_[13946]_ , \new_[13947]_ , \new_[13948]_ , \new_[13949]_ ,
    \new_[13950]_ , \new_[13951]_ , \new_[13952]_ , \new_[13953]_ ,
    \new_[13954]_ , \new_[13955]_ , \new_[13956]_ , \new_[13957]_ ,
    \new_[13958]_ , \new_[13959]_ , \new_[13961]_ , \new_[13962]_ ,
    \new_[13963]_ , \new_[13964]_ , \new_[13965]_ , \new_[13966]_ ,
    \new_[13967]_ , \new_[13968]_ , \new_[13969]_ , \new_[13970]_ ,
    \new_[13971]_ , \new_[13972]_ , \new_[13973]_ , \new_[13974]_ ,
    \new_[13975]_ , \new_[13976]_ , \new_[13977]_ , \new_[13978]_ ,
    \new_[13979]_ , \new_[13980]_ , \new_[13981]_ , \new_[13982]_ ,
    \new_[13983]_ , \new_[13984]_ , \new_[13985]_ , \new_[13986]_ ,
    \new_[13987]_ , \new_[13988]_ , \new_[13989]_ , \new_[13990]_ ,
    \new_[13991]_ , \new_[13992]_ , \new_[13993]_ , \new_[13994]_ ,
    \new_[13995]_ , \new_[13996]_ , \new_[13997]_ , \new_[13998]_ ,
    \new_[13999]_ , \new_[14000]_ , \new_[14001]_ , \new_[14002]_ ,
    \new_[14003]_ , \new_[14004]_ , \new_[14005]_ , \new_[14006]_ ,
    \new_[14007]_ , \new_[14008]_ , \new_[14009]_ , \new_[14010]_ ,
    \new_[14011]_ , \new_[14012]_ , \new_[14013]_ , \new_[14014]_ ,
    \new_[14015]_ , \new_[14016]_ , \new_[14017]_ , \new_[14018]_ ,
    \new_[14019]_ , \new_[14020]_ , \new_[14021]_ , \new_[14022]_ ,
    \new_[14023]_ , \new_[14024]_ , \new_[14025]_ , \new_[14026]_ ,
    \new_[14027]_ , \new_[14028]_ , \new_[14029]_ , \new_[14030]_ ,
    \new_[14031]_ , \new_[14032]_ , \new_[14033]_ , \new_[14034]_ ,
    \new_[14035]_ , \new_[14036]_ , \new_[14037]_ , \new_[14038]_ ,
    \new_[14039]_ , \new_[14041]_ , \new_[14042]_ , \new_[14043]_ ,
    \new_[14044]_ , \new_[14045]_ , \new_[14046]_ , \new_[14047]_ ,
    \new_[14048]_ , \new_[14049]_ , \new_[14050]_ , \new_[14051]_ ,
    \new_[14052]_ , \new_[14053]_ , \new_[14054]_ , \new_[14055]_ ,
    \new_[14056]_ , \new_[14057]_ , \new_[14058]_ , \new_[14059]_ ,
    \new_[14060]_ , \new_[14061]_ , \new_[14062]_ , \new_[14063]_ ,
    \new_[14064]_ , \new_[14065]_ , \new_[14066]_ , \new_[14067]_ ,
    \new_[14068]_ , \new_[14069]_ , \new_[14070]_ , \new_[14071]_ ,
    \new_[14072]_ , \new_[14073]_ , \new_[14074]_ , \new_[14075]_ ,
    \new_[14076]_ , \new_[14077]_ , \new_[14078]_ , \new_[14079]_ ,
    \new_[14080]_ , \new_[14081]_ , \new_[14082]_ , \new_[14083]_ ,
    \new_[14084]_ , \new_[14085]_ , \new_[14086]_ , \new_[14087]_ ,
    \new_[14088]_ , \new_[14089]_ , \new_[14090]_ , \new_[14091]_ ,
    \new_[14092]_ , \new_[14093]_ , \new_[14094]_ , \new_[14095]_ ,
    \new_[14096]_ , \new_[14097]_ , \new_[14098]_ , \new_[14099]_ ,
    \new_[14100]_ , \new_[14101]_ , \new_[14102]_ , \new_[14103]_ ,
    \new_[14104]_ , \new_[14105]_ , \new_[14106]_ , \new_[14107]_ ,
    \new_[14108]_ , \new_[14109]_ , \new_[14110]_ , \new_[14111]_ ,
    \new_[14112]_ , \new_[14113]_ , \new_[14114]_ , \new_[14115]_ ,
    \new_[14117]_ , \new_[14118]_ , \new_[14119]_ , \new_[14120]_ ,
    \new_[14121]_ , \new_[14122]_ , \new_[14123]_ , \new_[14124]_ ,
    \new_[14125]_ , \new_[14126]_ , \new_[14127]_ , \new_[14128]_ ,
    \new_[14129]_ , \new_[14130]_ , \new_[14131]_ , \new_[14132]_ ,
    \new_[14133]_ , \new_[14134]_ , \new_[14135]_ , \new_[14136]_ ,
    \new_[14137]_ , \new_[14138]_ , \new_[14139]_ , \new_[14140]_ ,
    \new_[14141]_ , \new_[14142]_ , \new_[14143]_ , \new_[14144]_ ,
    \new_[14145]_ , \new_[14146]_ , \new_[14147]_ , \new_[14148]_ ,
    \new_[14149]_ , \new_[14150]_ , \new_[14151]_ , \new_[14152]_ ,
    \new_[14153]_ , \new_[14154]_ , \new_[14155]_ , \new_[14156]_ ,
    \new_[14157]_ , \new_[14158]_ , \new_[14159]_ , \new_[14160]_ ,
    \new_[14161]_ , \new_[14162]_ , \new_[14163]_ , \new_[14164]_ ,
    \new_[14165]_ , \new_[14166]_ , \new_[14167]_ , \new_[14168]_ ,
    \new_[14169]_ , \new_[14170]_ , \new_[14171]_ , \new_[14172]_ ,
    \new_[14173]_ , \new_[14174]_ , \new_[14175]_ , \new_[14176]_ ,
    \new_[14177]_ , \new_[14178]_ , \new_[14179]_ , \new_[14180]_ ,
    \new_[14181]_ , \new_[14182]_ , \new_[14183]_ , \new_[14184]_ ,
    \new_[14185]_ , \new_[14186]_ , \new_[14187]_ , \new_[14188]_ ,
    \new_[14189]_ , \new_[14190]_ , \new_[14191]_ , \new_[14192]_ ,
    \new_[14193]_ , \new_[14194]_ , \new_[14195]_ , \new_[14196]_ ,
    \new_[14197]_ , \new_[14198]_ , \new_[14199]_ , \new_[14200]_ ,
    \new_[14201]_ , \new_[14202]_ , \new_[14203]_ , \new_[14204]_ ,
    \new_[14205]_ , \new_[14206]_ , \new_[14207]_ , \new_[14208]_ ,
    \new_[14209]_ , \new_[14210]_ , \new_[14211]_ , \new_[14212]_ ,
    \new_[14213]_ , \new_[14214]_ , \new_[14215]_ , \new_[14216]_ ,
    \new_[14217]_ , \new_[14218]_ , \new_[14219]_ , \new_[14220]_ ,
    \new_[14221]_ , \new_[14222]_ , \new_[14223]_ , \new_[14224]_ ,
    \new_[14225]_ , \new_[14226]_ , \new_[14227]_ , \new_[14228]_ ,
    \new_[14229]_ , \new_[14230]_ , \new_[14231]_ , \new_[14232]_ ,
    \new_[14233]_ , \new_[14234]_ , \new_[14235]_ , \new_[14236]_ ,
    \new_[14237]_ , \new_[14238]_ , \new_[14239]_ , \new_[14240]_ ,
    \new_[14241]_ , \new_[14242]_ , \new_[14243]_ , \new_[14244]_ ,
    \new_[14245]_ , \new_[14246]_ , \new_[14247]_ , \new_[14248]_ ,
    \new_[14249]_ , \new_[14250]_ , \new_[14251]_ , \new_[14252]_ ,
    \new_[14253]_ , \new_[14254]_ , \new_[14255]_ , \new_[14257]_ ,
    \new_[14258]_ , \new_[14259]_ , \new_[14260]_ , \new_[14261]_ ,
    \new_[14262]_ , \new_[14263]_ , \new_[14264]_ , \new_[14265]_ ,
    \new_[14267]_ , \new_[14268]_ , \new_[14269]_ , \new_[14270]_ ,
    \new_[14271]_ , \new_[14272]_ , \new_[14273]_ , \new_[14274]_ ,
    \new_[14275]_ , \new_[14276]_ , \new_[14277]_ , \new_[14278]_ ,
    \new_[14279]_ , \new_[14280]_ , \new_[14281]_ , \new_[14282]_ ,
    \new_[14283]_ , \new_[14284]_ , \new_[14285]_ , \new_[14286]_ ,
    \new_[14287]_ , \new_[14288]_ , \new_[14289]_ , \new_[14290]_ ,
    \new_[14291]_ , \new_[14292]_ , \new_[14293]_ , \new_[14294]_ ,
    \new_[14295]_ , \new_[14296]_ , \new_[14297]_ , \new_[14298]_ ,
    \new_[14299]_ , \new_[14300]_ , \new_[14301]_ , \new_[14302]_ ,
    \new_[14303]_ , \new_[14304]_ , \new_[14305]_ , \new_[14306]_ ,
    \new_[14307]_ , \new_[14308]_ , \new_[14309]_ , \new_[14310]_ ,
    \new_[14311]_ , \new_[14312]_ , \new_[14313]_ , \new_[14314]_ ,
    \new_[14315]_ , \new_[14316]_ , \new_[14317]_ , \new_[14318]_ ,
    \new_[14319]_ , \new_[14320]_ , \new_[14321]_ , \new_[14322]_ ,
    \new_[14323]_ , \new_[14324]_ , \new_[14325]_ , \new_[14326]_ ,
    \new_[14327]_ , \new_[14328]_ , \new_[14329]_ , \new_[14330]_ ,
    \new_[14331]_ , \new_[14332]_ , \new_[14333]_ , \new_[14334]_ ,
    \new_[14335]_ , \new_[14336]_ , \new_[14337]_ , \new_[14338]_ ,
    \new_[14339]_ , \new_[14340]_ , \new_[14341]_ , \new_[14342]_ ,
    \new_[14343]_ , \new_[14344]_ , \new_[14345]_ , \new_[14346]_ ,
    \new_[14347]_ , \new_[14348]_ , \new_[14349]_ , \new_[14350]_ ,
    \new_[14351]_ , \new_[14352]_ , \new_[14353]_ , \new_[14354]_ ,
    \new_[14355]_ , \new_[14356]_ , \new_[14357]_ , \new_[14358]_ ,
    \new_[14359]_ , \new_[14360]_ , \new_[14361]_ , \new_[14362]_ ,
    \new_[14363]_ , \new_[14364]_ , \new_[14365]_ , \new_[14366]_ ,
    \new_[14367]_ , \new_[14368]_ , \new_[14369]_ , \new_[14370]_ ,
    \new_[14371]_ , \new_[14372]_ , \new_[14373]_ , \new_[14374]_ ,
    \new_[14375]_ , \new_[14376]_ , \new_[14377]_ , \new_[14378]_ ,
    \new_[14379]_ , \new_[14380]_ , \new_[14381]_ , \new_[14382]_ ,
    \new_[14383]_ , \new_[14384]_ , \new_[14385]_ , \new_[14386]_ ,
    \new_[14387]_ , \new_[14388]_ , \new_[14389]_ , \new_[14390]_ ,
    \new_[14391]_ , \new_[14392]_ , \new_[14393]_ , \new_[14394]_ ,
    \new_[14395]_ , \new_[14396]_ , \new_[14397]_ , \new_[14398]_ ,
    \new_[14399]_ , \new_[14400]_ , \new_[14401]_ , \new_[14402]_ ,
    \new_[14403]_ , \new_[14404]_ , \new_[14405]_ , \new_[14406]_ ,
    \new_[14407]_ , \new_[14408]_ , \new_[14409]_ , \new_[14410]_ ,
    \new_[14411]_ , \new_[14412]_ , \new_[14413]_ , \new_[14414]_ ,
    \new_[14415]_ , \new_[14416]_ , \new_[14417]_ , \new_[14418]_ ,
    \new_[14419]_ , \new_[14420]_ , \new_[14421]_ , \new_[14422]_ ,
    \new_[14423]_ , \new_[14424]_ , \new_[14425]_ , \new_[14426]_ ,
    \new_[14427]_ , \new_[14428]_ , \new_[14429]_ , \new_[14430]_ ,
    \new_[14431]_ , \new_[14433]_ , \new_[14434]_ , \new_[14435]_ ,
    \new_[14436]_ , \new_[14437]_ , \new_[14438]_ , \new_[14439]_ ,
    \new_[14440]_ , \new_[14441]_ , \new_[14442]_ , \new_[14443]_ ,
    \new_[14444]_ , \new_[14445]_ , \new_[14446]_ , \new_[14447]_ ,
    \new_[14448]_ , \new_[14449]_ , \new_[14450]_ , \new_[14451]_ ,
    \new_[14452]_ , \new_[14453]_ , \new_[14454]_ , \new_[14455]_ ,
    \new_[14456]_ , \new_[14457]_ , \new_[14458]_ , \new_[14459]_ ,
    \new_[14460]_ , \new_[14461]_ , \new_[14462]_ , \new_[14463]_ ,
    \new_[14464]_ , \new_[14465]_ , \new_[14466]_ , \new_[14467]_ ,
    \new_[14468]_ , \new_[14469]_ , \new_[14470]_ , \new_[14471]_ ,
    \new_[14472]_ , \new_[14473]_ , \new_[14474]_ , \new_[14475]_ ,
    \new_[14476]_ , \new_[14477]_ , \new_[14478]_ , \new_[14479]_ ,
    \new_[14480]_ , \new_[14481]_ , \new_[14482]_ , \new_[14483]_ ,
    \new_[14484]_ , \new_[14485]_ , \new_[14486]_ , \new_[14487]_ ,
    \new_[14488]_ , \new_[14489]_ , \new_[14490]_ , \new_[14491]_ ,
    \new_[14492]_ , \new_[14493]_ , \new_[14494]_ , \new_[14495]_ ,
    \new_[14497]_ , \new_[14498]_ , \new_[14499]_ , \new_[14501]_ ,
    \new_[14502]_ , \new_[14503]_ , \new_[14504]_ , \new_[14505]_ ,
    \new_[14506]_ , \new_[14507]_ , \new_[14508]_ , \new_[14509]_ ,
    \new_[14510]_ , \new_[14511]_ , \new_[14512]_ , \new_[14513]_ ,
    \new_[14514]_ , \new_[14515]_ , \new_[14516]_ , \new_[14517]_ ,
    \new_[14518]_ , \new_[14519]_ , \new_[14520]_ , \new_[14521]_ ,
    \new_[14522]_ , \new_[14523]_ , \new_[14524]_ , \new_[14525]_ ,
    \new_[14526]_ , \new_[14527]_ , \new_[14528]_ , \new_[14529]_ ,
    \new_[14530]_ , \new_[14531]_ , \new_[14532]_ , \new_[14533]_ ,
    \new_[14534]_ , \new_[14535]_ , \new_[14536]_ , \new_[14537]_ ,
    \new_[14538]_ , \new_[14539]_ , \new_[14540]_ , \new_[14541]_ ,
    \new_[14542]_ , \new_[14543]_ , \new_[14544]_ , \new_[14545]_ ,
    \new_[14546]_ , \new_[14547]_ , \new_[14548]_ , \new_[14549]_ ,
    \new_[14550]_ , \new_[14551]_ , \new_[14552]_ , \new_[14553]_ ,
    \new_[14554]_ , \new_[14555]_ , \new_[14556]_ , \new_[14557]_ ,
    \new_[14558]_ , \new_[14559]_ , \new_[14560]_ , \new_[14561]_ ,
    \new_[14562]_ , \new_[14563]_ , \new_[14564]_ , \new_[14565]_ ,
    \new_[14566]_ , \new_[14567]_ , \new_[14568]_ , \new_[14569]_ ,
    \new_[14570]_ , \new_[14571]_ , \new_[14572]_ , \new_[14573]_ ,
    \new_[14574]_ , \new_[14575]_ , \new_[14576]_ , \new_[14577]_ ,
    \new_[14578]_ , \new_[14579]_ , \new_[14580]_ , \new_[14581]_ ,
    \new_[14582]_ , \new_[14583]_ , \new_[14584]_ , \new_[14585]_ ,
    \new_[14586]_ , \new_[14587]_ , \new_[14588]_ , \new_[14589]_ ,
    \new_[14590]_ , \new_[14591]_ , \new_[14592]_ , \new_[14593]_ ,
    \new_[14594]_ , \new_[14595]_ , \new_[14596]_ , \new_[14597]_ ,
    \new_[14598]_ , \new_[14599]_ , \new_[14600]_ , \new_[14601]_ ,
    \new_[14602]_ , \new_[14603]_ , \new_[14604]_ , \new_[14605]_ ,
    \new_[14606]_ , \new_[14607]_ , \new_[14608]_ , \new_[14609]_ ,
    \new_[14610]_ , \new_[14611]_ , \new_[14612]_ , \new_[14613]_ ,
    \new_[14614]_ , \new_[14615]_ , \new_[14616]_ , \new_[14617]_ ,
    \new_[14618]_ , \new_[14619]_ , \new_[14620]_ , \new_[14621]_ ,
    \new_[14622]_ , \new_[14623]_ , \new_[14624]_ , \new_[14625]_ ,
    \new_[14626]_ , \new_[14627]_ , \new_[14628]_ , \new_[14629]_ ,
    \new_[14630]_ , \new_[14631]_ , \new_[14632]_ , \new_[14633]_ ,
    \new_[14634]_ , \new_[14635]_ , \new_[14636]_ , \new_[14637]_ ,
    \new_[14638]_ , \new_[14639]_ , \new_[14640]_ , \new_[14641]_ ,
    \new_[14642]_ , \new_[14643]_ , \new_[14644]_ , \new_[14645]_ ,
    \new_[14646]_ , \new_[14647]_ , \new_[14648]_ , \new_[14649]_ ,
    \new_[14650]_ , \new_[14651]_ , \new_[14652]_ , \new_[14653]_ ,
    \new_[14654]_ , \new_[14655]_ , \new_[14656]_ , \new_[14657]_ ,
    \new_[14658]_ , \new_[14659]_ , \new_[14660]_ , \new_[14661]_ ,
    \new_[14662]_ , \new_[14663]_ , \new_[14664]_ , \new_[14665]_ ,
    \new_[14666]_ , \new_[14667]_ , \new_[14668]_ , \new_[14669]_ ,
    \new_[14670]_ , \new_[14671]_ , \new_[14672]_ , \new_[14673]_ ,
    \new_[14674]_ , \new_[14675]_ , \new_[14676]_ , \new_[14677]_ ,
    \new_[14678]_ , \new_[14679]_ , \new_[14680]_ , \new_[14681]_ ,
    \new_[14682]_ , \new_[14683]_ , \new_[14684]_ , \new_[14685]_ ,
    \new_[14686]_ , \new_[14687]_ , \new_[14688]_ , \new_[14689]_ ,
    \new_[14690]_ , \new_[14691]_ , \new_[14692]_ , \new_[14693]_ ,
    \new_[14694]_ , \new_[14695]_ , \new_[14696]_ , \new_[14697]_ ,
    \new_[14698]_ , \new_[14699]_ , \new_[14700]_ , \new_[14701]_ ,
    \new_[14702]_ , \new_[14703]_ , \new_[14704]_ , \new_[14705]_ ,
    \new_[14706]_ , \new_[14707]_ , \new_[14708]_ , \new_[14709]_ ,
    \new_[14710]_ , \new_[14711]_ , \new_[14712]_ , \new_[14713]_ ,
    \new_[14714]_ , \new_[14715]_ , \new_[14716]_ , \new_[14717]_ ,
    \new_[14718]_ , \new_[14719]_ , \new_[14720]_ , \new_[14721]_ ,
    \new_[14722]_ , \new_[14723]_ , \new_[14724]_ , \new_[14725]_ ,
    \new_[14726]_ , \new_[14727]_ , \new_[14728]_ , \new_[14729]_ ,
    \new_[14730]_ , \new_[14731]_ , \new_[14732]_ , \new_[14733]_ ,
    \new_[14734]_ , \new_[14735]_ , \new_[14736]_ , \new_[14737]_ ,
    \new_[14738]_ , \new_[14739]_ , \new_[14740]_ , \new_[14741]_ ,
    \new_[14742]_ , \new_[14743]_ , \new_[14744]_ , \new_[14745]_ ,
    \new_[14746]_ , \new_[14747]_ , \new_[14748]_ , \new_[14749]_ ,
    \new_[14750]_ , \new_[14751]_ , \new_[14752]_ , \new_[14753]_ ,
    \new_[14754]_ , \new_[14755]_ , \new_[14756]_ , \new_[14757]_ ,
    \new_[14758]_ , \new_[14759]_ , \new_[14760]_ , \new_[14761]_ ,
    \new_[14762]_ , \new_[14763]_ , \new_[14764]_ , \new_[14765]_ ,
    \new_[14766]_ , \new_[14767]_ , \new_[14768]_ , \new_[14769]_ ,
    \new_[14770]_ , \new_[14771]_ , \new_[14772]_ , \new_[14773]_ ,
    \new_[14774]_ , \new_[14775]_ , \new_[14776]_ , \new_[14777]_ ,
    \new_[14778]_ , \new_[14780]_ , \new_[14781]_ , \new_[14782]_ ,
    \new_[14783]_ , \new_[14784]_ , \new_[14785]_ , \new_[14786]_ ,
    \new_[14787]_ , \new_[14788]_ , \new_[14789]_ , \new_[14790]_ ,
    \new_[14791]_ , \new_[14792]_ , \new_[14793]_ , \new_[14794]_ ,
    \new_[14795]_ , \new_[14796]_ , \new_[14797]_ , \new_[14798]_ ,
    \new_[14799]_ , \new_[14800]_ , \new_[14801]_ , \new_[14802]_ ,
    \new_[14803]_ , \new_[14804]_ , \new_[14805]_ , \new_[14806]_ ,
    \new_[14807]_ , \new_[14808]_ , \new_[14809]_ , \new_[14810]_ ,
    \new_[14811]_ , \new_[14812]_ , \new_[14813]_ , \new_[14814]_ ,
    \new_[14815]_ , \new_[14816]_ , \new_[14817]_ , \new_[14818]_ ,
    \new_[14819]_ , \new_[14820]_ , \new_[14821]_ , \new_[14822]_ ,
    \new_[14823]_ , \new_[14824]_ , \new_[14825]_ , \new_[14826]_ ,
    \new_[14827]_ , \new_[14828]_ , \new_[14829]_ , \new_[14830]_ ,
    \new_[14831]_ , \new_[14832]_ , \new_[14833]_ , \new_[14834]_ , n500,
    n505, n510, n515, n520, n525, n530, n535, n540, n545, n550, n555, n560,
    n565, n570, n575, n580, n585, n590, n595, n600, n605, n610, n615, n620,
    n625, n630, n635, n640, n645, n650, n655, n660, n665, n670, n675, n680,
    n685, n690, n695, n700, n705, n710, n715, n720, n725, n730, n735, n740,
    n745, n750, n755, n760, n765, n770, n775, n780, n785, n790, n795, n800,
    n805, n810, n815, n820, n825, n830, n835, n840, n845, n850, n855, n860,
    n865, n870, n875, n880, n885, n890, n895, n900, n905, n910, n915, n920,
    n925, n930, n935, n940, n945, n950, n955, n960, n965, n970, n975, n980,
    n985, n990, n995, n1000, n1005, n1010, n1015, n1020, n1025, n1030,
    n1035, n1040, n1045, n1050, n1055, n1060, n1065, n1070, n1075, n1080,
    n1085, n1090, n1095, n1100, n1105, n1110, n1115, n1120, n1125, n1130,
    n1135, n1140, n1145, n1150, n1155, n1160, n1165, n1170, n1175, n1180,
    n1185, n1190, n1195, n1200, n1205, n1210, n1215, n1220, n1225, n1230,
    n1235, n1240, n1245, n1250, n1255, n1260, n1265, n1270, n1275, n1280,
    n1285, n1290, n1295, n1300, n1305, n1310, n1315, n1320, n1325, n1330,
    n1335, n1340, n1345, n1350, n1355, n1360, n1365, n1370, n1375, n1380,
    n1385, n1390, n1395, n1400, n1405, n1410, n1415, n1420, n1425, n1430,
    n1435, n1440, n1445, n1450, n1455, n1460, n1465, n1470, n1475, n1480,
    n1485, n1490, n1495, n1500, n1505, n1510, n1515, n1520, n1525, n1530,
    n1535, n1540, n1545, n1550, n1555, n1560, n1565, n1570, n1575, n1580,
    n1585, n1590, n1595, n1600, n1605, n1610, n1615, n1620, n1625, n1630,
    n1635, n1640, n1645, n1650, n1655, n1660, n1665, n1670, n1675, n1680,
    n1685, n1690, n1695, n1700, n1705, n1710, n1715, n1720, n1725, n1730,
    n1735, n1740, n1745, n1750, n1755, n1760, n1765, n1770, n1775, n1780,
    n1785, n1790, n1795, n1800, n1805, n1810, n1815, n1820, n1825, n1830,
    n1835, n1840, n1845, n1850, n1855, n1860, n1865, n1870, n1875, n1880,
    n1885, n1890, n1895, n1900, n1905, n1910, n1915, n1920, n1925, n1930,
    n1935, n1940, n1945, n1950, n1955, n1960, n1965, n1970, n1975, n1980,
    n1985, n1990, n1995, n2000, n2005, n2010, n2015, n2020, n2025, n2030,
    n2035, n2040, n2045, n2050, n2055, n2060, n2065, n2070, n2075, n2080,
    n2085, n2090, n2095, n2100, n2105, n2110, n2115, n2120, n2125, n2130,
    n2135, n2140, n2145, n2150, n2155, n2160, n2165, n2170, n2175, n2180,
    n2185, n2190, n2195, n2200, n2205, n2210, n2215, n2220, n2225, n2230,
    n2235, n2240, n2245, n2250, n2255, n2260, n2265, n2270, n2275, n2280,
    n2285, n2290, n2295, n2300, n2305, n2310, n2315, n2320, n2325, n2330,
    n2335, n2340, n2345, n2350, n2355, n2360, n2365, n2370, n2375, n2380,
    n2385, n2390, n2395, n2400, n2405, n2410, n2415, n2420, n2425, n2430,
    n2435, n2440, n2445, n2450, n2455, n2460, n2465, n2470, n2475, n2480,
    n2485, n2490, n2495, n2500, n2505, n2510, n2515, n2520, n2525, n2530,
    n2535, n2540, n2545, n2550, n2555, n2560, n2565, n2570, n2575, n2580,
    n2585, n2590, n2595, n2600, n2605, n2610, n2615, n2620, n2625, n2630,
    n2635, n2640, n2645, n2650, n2655, n2660, n2665, n2670, n2675, n2680,
    n2685, n2690, n2695, n2700, n2705, n2710, n2715, n2720, n2725, n2730,
    n2735, n2740, n2745, n2750, n2755, n2760, n2765, n2770, n2775, n2780,
    n2785, n2790, n2795, n2800, n2805, n2810, n2815, n2820, n2825, n2830,
    n2835, n2840, n2845, n2850, n2855, n2860, n2865, n2870, n2875, n2880,
    n2885, n2890, n2895, n2900, n2905, n2910, n2915, n2920, n2925, n2930,
    n2935, n2940, n2945, n2950, n2955, n2960, n2965, n2970, n2975, n2980,
    n2985, n2990, n2995, n3000, n3005, n3010, n3015, n3020, n3025, n3030,
    n3035, n3040, n3045, n3050, n3055, n3060, n3065, n3070, n3075, n3080,
    n3085, n3090, n3095, n3100, n3105, n3110, n3115, n3120, n3125, n3130,
    n3135, n3140, n3145, n3150, n3155, n3160, n3165, n3170, n3175, n3180,
    n3185, n3190, n3195, n3200, n3205, n3210, n3215, n3220, n3225, n3230,
    n3235, n3240, n3245, n3250, n3255, n3260, n3265, n3270, n3275, n3280,
    n3285, n3290, n3295, n3300, n3305, n3310, n3315, n3320, n3325, n3330,
    n3335, n3340, n3345, n3350, n3355, n3360, n3365, n3370, n3375, n3380,
    n3385, n3390, n3395, n3400, n3405, n3410, n3415, n3420, n3425, n3430,
    n3435, n3440, n3445, n3450, n3455, n3460, n3465, n3470, n3475, n3480,
    n3485, n3490, n3495, n3500, n3505, n3510, n3515, n3520, n3525, n3530,
    n3535, n3540, n3545, n3550, n3555, n3560, n3565, n3570, n3575, n3580,
    n3585, n3590, n3595, n3600, n3605, n3610, n3615, n3620, n3625, n3630,
    n3635, n3640, n3645, n3650, n3655, n3660, n3665, n3670, n3675, n3680,
    n3685, n3690, n3695, n3700, n3705, n3710, n3715, n3720, n3725, n3730,
    n3735, n3740, n3745, n3750, n3755, n3760, n3765, n3770, n3775, n3780,
    n3785, n3790, n3795, n3800, n3805, n3810, n3815, n3820, n3825, n3830,
    n3835, n3840, n3845, n3850, n3855, n3860, n3865, n3870, n3875, n3880,
    n3885, n3890, n3895, n3900, n3905, n3910, n3915, n3920, n3925, n3930,
    n3935, n3940, n3945, n3950, n3955, n3960, n3965, n3970, n3975, n3980,
    n3985, n3990, n3995, n4000, n4005, n4010, n4015, n4020, n4025, n4030,
    n4035, n4040, n4045, n4050, n4055, n4060, n4065, n4070, n4075, n4080,
    n4085, n4090, n4095, n4100, n4105, n4110, n4115, n4120, n4125, n4130,
    n4135, n4140, n4145, n4150, n4155, n4160, n4165, n4170, n4175, n4180,
    n4185, n4190, n4195, n4200, n4205, n4210, n4215, n4220, n4225, n4230,
    n4235, n4240, n4245, n4250, n4255, n4260, n4265, n4270, n4275, n4280,
    n4285, n4290, n4295, n4300, n4305, n4310, n4315, n4320, n4325, n4330,
    n4335, n4340, n4345, n4350, n4355, n4360, n4365, n4370, n4375, n4380,
    n4385, n4390, n4395, n4400, n4405, n4410, n4415, n4420, n4425, n4430,
    n4435, n4440, n4445, n4450, n4455, n4460, n4465, n4470, n4475, n4480,
    n4485, n4490, n4495, n4500, n4505, n4510, n4515, n4520, n4525, n4530,
    n4535, n4540, n4545, n4550, n4555, n4560, n4565, n4570, n4575, n4580,
    n4585, n4590, n4595, n4600, n4605, n4610, n4615, n4620, n4625, n4630,
    n4635, n4640, n4645, n4650, n4655, n4660, n4665, n4670, n4675, n4680,
    n4685, n4690, n4695, n4700, n4705, n4710, n4715, n4720, n4725, n4730,
    n4735, n4740, n4745, n4750, n4755, n4760, n4765, n4770, n4775, n4780,
    n4785, n4790, n4795, n4800, n4805, n4810, n4815, n4820, n4825, n4830,
    n4835, n4840, n4845, n4850, n4855, n4860, n4865, n4870, n4875, n4880,
    n4885, n4890, n4895, n4900, n4905, n4910, n4915, n4920, n4925, n4930,
    n4935, n4940, n4945, n4950, n4955, n4960, n4965, n4970, n4975, n4980,
    n4985, n4990, n4995, n5000, n5005, n5010, n5015, n5020, n5025, n5030,
    n5035, n5040, n5045, n5050, n5055, n5060, n5065, n5070, n5075, n5080,
    n5085, n5090, n5095, n5100, n5105, n5110, n5115, n5120, n5125, n5130,
    n5135, n5140, n5145, n5150, n5155, n5160, n5165, n5170, n5175, n5180,
    n5185, n5190, n5195, n5200, n5205, n5210, n5215, n5220, n5225, n5230,
    n5235, n5240, n5245, n5250, n5255, n5260, n5265, n5270, n5275, n5280,
    n5285, n5290, n5295, n5300, n5305, n5310, n5315, n5320, n5325, n5330,
    n5335, n5340, n5345, n5350, n5355, n5360, n5365, n5370, n5375, n5380,
    n5385, n5390, n5395, n5400, n5405, n5410, n5415, n5420, n5425, n5430,
    n5435, n5440, n5445, n5450, n5455, n5460, n5465, n5470, n5475, n5480,
    n5485, n5490, n5495, n5500, n5505, n5510, n5515, n5520, n5525, n5530,
    n5535, n5540, n5545, n5550, n5555, n5560, n5565, n5570, n5575, n5580,
    n5585, n5590, n5595, n5600, n5605, n5610, n5615, n5620, n5625, n5630,
    n5635, n5640, n5645, n5650, n5655, n5660, n5665, n5670, n5675, n5680,
    n5685, n5690, n5695, n5700, n5705, n5710, n5715, n5720, n5725, n5730,
    n5735, n5740, n5745, n5750, n5755, n5760, n5765, n5770, n5775, n5780,
    n5785, n5790, n5795, n5800, n5805, n5810, n5815, n5820, n5825, n5830,
    n5835, n5840, n5845, n5850, n5855, n5860, n5865, n5870, n5875, n5880,
    n5885, n5890, n5895, n5900, n5905, n5910, n5915, n5920, n5925, n5930,
    n5935, n5940, n5945, n5950, n5955, n5960, n5965, n5970, n5975, n5980,
    n5985, n5990, n5995, n6000, n6005, n6010, n6015, n6020, n6025, n6030,
    n6035, n6040, n6045, n6050, n6055, n6060, n6065, n6070, n6075, n6080,
    n6085, n6090, n6095, n6100, n6105, n6110, n6115, n6120, n6125, n6130,
    n6135, n6140, n6145, n6150, n6155, n6160, n6165, n6170, n6175, n6180,
    n6185, n6190, n6195, n6200, n6205, n6210, n6215, n6220, n6225, n6230,
    n6235, n6240, n6245, n6250, n6255, n6260, n6265, n6270, n6275, n6280,
    n6285, n6290, n6295, n6300, n6305, n6310, n6315, n6320, n6325, n6330,
    n6335, n6340, n6345, n6350, n6355, n6360, n6365, n6370, n6375, n6380,
    n6385, n6390, n6395, n6400, n6405, n6410, n6415, n6420, n6425, n6430,
    n6435, n6440, n6445, n6450, n6455, n6460, n6465, n6470, n6475, n6480,
    n6485, n6490, n6495, n6500, n6505, n6510, n6515, n6520, n6525, n6530,
    n6535, n6540, n6545, n6550, n6555, n6560, n6565, n6570, n6575, n6580,
    n6585, n6590, n6595, n6600, n6605, n6610, n6615, n6620, n6625, n6630,
    n6635, n6640, n6645, n6650, n6655, n6660, n6665, n6670, n6675, n6680,
    n6685, n6690, n6695, n6700, n6705, n6710, n6715, n6720, n6725, n6730,
    n6735, n6740, n6745, n6750, n6755, n6760, n6765, n6770, n6775, n6780,
    n6785, n6790, n6795, n6800, n6805, n6810, n6815, n6820, n6825, n6830,
    n6835, n6840, n6845, n6850, n6855, n6860, n6865, n6870, n6875, n6880,
    n6885, n6890, n6895, n6900, n6905, n6910, n6915, n6920, n6925, n6930,
    n6935, n6940, n6945, n6950, n6955, n6960, n6965, n6970, n6975, n6980,
    n6985, n6990, n6995, n7000, n7005, n7010, n7015, n7020, n7025, n7030,
    n7035, n7040, n7045, n7050, n7055, n7060, n7065, n7070, n7075, n7080,
    n7085, n7090, n7095, n7100, n7105, n7110, n7115, n7120, n7125, n7130,
    n7135, n7140, n7145, n7150, n7155, n7160, n7165, n7170, n7175, n7180,
    n7185, n7190, n7195, n7200, n7205, n7210, n7215, n7220, n7225, n7230,
    n7235, n7240, n7245, n7250, n7255, n7260, n7265, n7270, n7275, n7280,
    n7285, n7290, n7295, n7300, n7305, n7310, n7315, n7320, n7325, n7330,
    n7335, n7340, n7345, n7350, n7355, n7360, n7365, n7370, n7375, n7380,
    n7385, n7390, n7395, n7400, n7405, n7410, n7415, n7420, n7425, n7430,
    n7435, n7440, n7445, n7450, n7455, n7460, n7465, n7470, n7475, n7480,
    n7485, n7490, n7495, n7500, n7505, n7510, n7515, n7520, n7525, n7530,
    n7535, n7540, n7545, n7550, n7555, n7560, n7565, n7570, n7575, n7580,
    n7585, n7590, n7595, n7600, n7605, n7610, n7615, n7620, n7625, n7630,
    n7635, n7640, n7645, n7650, n7655, n7660, n7665, n7670, n7675, n7680,
    n7685, n7690, n7695, n7700, n7705, n7710, n7715, n7720, n7725, n7730,
    n7735, n7740, n7745, n7750, n7755, n7760, n7765, n7770, n7775, n7780,
    n7785, n7790, n7795, n7800, n7805, n7810, n7815, n7820, n7825, n7830,
    n7835, n7840, n7845, n7850, n7855, n7860, n7865, n7870, n7875, n7880,
    n7885, n7890, n7895, n7900, n7905, n7910, n7915, n7920, n7925, n7930,
    n7935, n7940, n7945, n7950, n7955, n7960, n7965, n7970, n7975, n7980,
    n7985, n7990, n7995, n8000, n8005, n8010, n8015, n8020, n8025, n8030,
    n8035, n8040, n8045, n8050, n8055, n8060, n8065, n8070, n8075, n8080,
    n8085, n8090, n8095, n8100, n8105, n8110, n8115, n8120, n8125, n8130,
    n8135, n8140, n8145, n8150, n8155, n8160, n8165, n8170, n8175, n8180,
    n8185, n8190, n8195, n8200, n8205, n8210, n8215, n8220, n8225, n8230,
    n8235, n8240, n8245, n8250, n8255, n8260, n8265, n8270, n8275, n8280,
    n8285, n8290, n8295, n8300, n8305, n8310, n8315, n8320, n8325, n8330,
    n8335, n8340, n8345, n8350, n8355, n8360, n8365, n8370, n8375, n8380,
    n8385, n8390, n8395, n8400, n8405, n8410, n8415, n8420, n8425, n8430,
    n8435, n8440, n8445, n8450, n8455, n8460, n8465, n8470, n8475, n8480,
    n8485, n8490, n8495, n8500, n8505, n8510, n8515, n8520, n8525, n8530,
    n8535, n8540, n8545, n8550, n8555, n8560, n8565, n8570, n8575, n8580,
    n8585, n8590, n8595, n8600, n8605, n8610, n8615, n8620, n8625, n8630,
    n8635, n8640, n8645, n8650, n8655, n8660, n8665, n8670, n8675, n8680,
    n8685, n8690, n8695, n8700, n8705, n8710, n8715, n8720, n8725, n8730,
    n8735, n8740, n8745, n8750, n8755, n8760, n8765, n8770, n8775, n8780,
    n8785, n8790, n8795, n8800, n8805, n8810, n8815, n8820, n8825, n8830,
    n8835, n8840, n8845, n8850, n8855, n8860, n8865, n8870, n8875, n8880,
    n8885, n8890, n8895, n8900, n8905, n8910, n8915, n8920, n8925, n8930,
    n8935, n8940, n8945, n8950, n8955, n8960, n8965, n8970, n8975, n8980,
    n8985, n8990, n8995, n9000, n9005, n9010, n9015, n9020, n9025, n9030,
    n9035, n9040, n9045, n9050, n9055, n9060, n9065, n9070, n9075, n9080,
    n9085, n9090, n9095, n9100, n9105, n9110, n9115, n9120, n9125, n9130,
    n9135, n9140, n9145, n9150, n9155, n9160, n9165, n9170, n9175, n9180,
    n9185, n9190, n9195, n9200, n9205, n9210, n9215, n9220, n9225;
  assign \new_[1995]_  = 1'b0;
  assign \new_[1996]_  = 1'b1;
  assign sram_re_o = \new_[1996]_ ;
  assign \dma_req_o[4]  = \new_[1995]_ ;
  assign \dma_req_o[5]  = \new_[1995]_ ;
  assign \dma_req_o[6]  = \new_[1995]_ ;
  assign \dma_req_o[7]  = \new_[1995]_ ;
  assign \dma_req_o[8]  = \new_[1995]_ ;
  assign \dma_req_o[9]  = \new_[1995]_ ;
  assign \dma_req_o[10]  = \new_[1995]_ ;
  assign \dma_req_o[11]  = \new_[1995]_ ;
  assign \dma_req_o[12]  = \new_[1995]_ ;
  assign \dma_req_o[13]  = \new_[1995]_ ;
  assign \dma_req_o[14]  = \new_[1995]_ ;
  assign \dma_req_o[15]  = \new_[1995]_ ;
  assign \DataOut_pad_o[3]  = \\u0_DataOut_reg[3] ;
  assign \DataOut_pad_o[7]  = \\u0_DataOut_reg[7] ;
  assign n500 = ~\new_[2227]_  | (~\new_[2014]_  & ~\new_[2257]_ );
  assign n505 = ~\new_[2233]_  | (~\new_[2015]_  & ~\new_[2257]_ );
  assign \new_[2014]_  = \new_[2018]_  ? \new_[2328]_  : \new_[2198]_ ;
  assign \new_[2015]_  = \new_[2021]_  ? \new_[2328]_  : \new_[2200]_ ;
  assign \DataOut_pad_o[2]  = \\u0_DataOut_reg[2] ;
  assign \DataOut_pad_o[6]  = \\u0_DataOut_reg[6] ;
  assign \new_[2018]_  = \new_[2022]_  ^ \new_[2027]_ ;
  assign n510 = ~\new_[2226]_  | (~\new_[2023]_  & ~\new_[2257]_ );
  assign n515 = ~\new_[2231]_  | (~\new_[2024]_  & ~\new_[2257]_ );
  assign \new_[2021]_  = \new_[2025]_  ^ \new_[2027]_ ;
  assign \new_[2022]_  = ~\new_[2025]_ ;
  assign \new_[2023]_  = \new_[2027]_  ? \new_[2328]_  : \new_[2197]_ ;
  assign \new_[2024]_  = ~\new_[2159]_  | (~\new_[2328]_  & ~\new_[2027]_ );
  assign \new_[2025]_  = ~\\u1_u3_token_pid_sel_reg[0] ;
  assign n520 = (~\new_[2725]_  & ~\new_[11024]_  & ~\new_[12680]_ ) | (~\new_[2611]_  & ~\new_[2029]_  & ~\new_[11023]_ );
  assign \new_[2027]_  = ~\\u1_u3_token_pid_sel_reg[1] ;
  assign n525 = ~\new_[2572]_  | (~\new_[2030]_  & ~\new_[3243]_ );
  assign \new_[2029]_  = ~\new_[4148]_  & (~\new_[2031]_  | ~\new_[3597]_ );
  assign \new_[2030]_  = \new_[2032]_  | \new_[11023]_ ;
  assign \new_[2031]_  = ~\new_[2032]_ ;
  assign \new_[2032]_  = ~\new_[8959]_  | ~\new_[2036]_  | ~\new_[2033]_ ;
  assign \new_[2033]_  = u1_u3_no_bufs0_reg;
  assign \new_[2034]_  = \\u1_u3_idin_reg[13] ;
  assign n535 = ~\new_[2102]_  | ~\new_[2043]_  | ~\new_[13072]_ ;
  assign \new_[2036]_  = u1_u3_no_bufs1_reg;
  assign n530 = ~\new_[4270]_  | ~\new_[2054]_  | ~\new_[9561]_  | ~\new_[13658]_ ;
  assign \new_[2038]_  = \\u1_u1_crc16_reg[15] ;
  assign \new_[2039]_  = ~\\u1_u1_crc16_reg[1] ;
  assign \new_[2040]_  = \\u1_u3_idin_reg[14] ;
  assign n540 = \new_[2056]_  | \new_[8810]_ ;
  assign \new_[2042]_  = u1_u3_buffer_done_reg;
  assign \new_[2043]_  = ~\new_[14284]_ ;
  assign n550 = ~\new_[6207]_  | ~\new_[2070]_  | ~\new_[10117]_ ;
  assign n555 = \new_[2065]_  ? n9145 : \new_[13594]_ ;
  assign \new_[2046]_  = ~\\u1_u1_crc16_reg[0] ;
  assign \new_[2047]_  = \\u1_u3_idin_reg[12] ;
  assign \new_[2048]_  = \\u1_u3_idin_reg[16] ;
  assign \new_[2049]_  = \\u1_u3_idin_reg[10] ;
  assign n545 = ~\new_[6206]_  | ~\new_[2066]_  | ~\new_[10117]_ ;
  assign \DataOut_pad_o[4]  = \\u0_DataOut_reg[4] ;
  assign \new_[2052]_  = \\u1_u3_idin_reg[15] ;
  assign \new_[2053]_  = \\u1_u3_idin_reg[11] ;
  assign \new_[2054]_  = ~\new_[11573]_  | ~\new_[8261]_  | ~\new_[2072]_ ;
  assign n560 = \new_[2072]_  ? \new_[9036]_  : \new_[2081]_ ;
  assign \new_[2056]_  = \new_[2072]_  ? \new_[8261]_  : \new_[4011]_ ;
  assign n580 = \new_[2099]_  ? n9145 : \new_[14019]_ ;
  assign n570 = \new_[2100]_  ? n9145 : \new_[13921]_ ;
  assign n575 = \new_[2101]_  ? n9145 : \new_[14247]_ ;
  assign \DataOut_pad_o[1]  = \\u0_DataOut_reg[1] ;
  assign \DataOut_pad_o[0]  = \\u0_DataOut_reg[0] ;
  assign \new_[2062]_  = \\u1_u3_idin_reg[9] ;
  assign n565 = ~\new_[6202]_  | ~\new_[10117]_  | ~\new_[2080]_ ;
  assign \new_[2064]_  = \\u1_u3_idin_reg[6] ;
  assign \new_[2065]_  = \new_[4858]_  ^ \new_[2109]_ ;
  assign \new_[2066]_  = ~\new_[6759]_  | ~\new_[14763]_ ;
  assign n585 = ~\new_[2228]_  | ~\new_[2079]_ ;
  assign n590 = ~\new_[13067]_  | (~\new_[2111]_  & ~n9145);
  assign n595 = \new_[14433]_  ? n9145 : \new_[13654]_ ;
  assign \new_[2070]_  = ~\new_[6759]_  | ~\new_[14303]_ ;
  assign n600 = ~\new_[2224]_  | ~\new_[2106]_ ;
  assign \new_[2072]_  = u1_u3_buffer_full_reg;
  assign \new_[2073]_  = ~\\u1_u1_crc16_reg[8] ;
  assign \DataOut_pad_o[5]  = \\u0_DataOut_reg[5] ;
  assign \new_[2075]_  = \\u1_u3_idin_reg[8] ;
  assign \new_[2076]_  = \\u1_u3_idin_reg[5] ;
  assign n605 = ~\new_[2229]_  | ~\new_[2103]_ ;
  assign n610 = \new_[2117]_  ? n9145 : \new_[13628]_ ;
  assign \new_[2079]_  = ~\new_[2112]_  & ~\new_[2225]_ ;
  assign \new_[2080]_  = ~\new_[6759]_  | ~\new_[2113]_ ;
  assign \new_[2081]_  = u1_u3_buffer_empty_reg;
  assign \new_[2082]_  = \\u1_u3_idin_reg[7] ;
  assign \new_[2083]_  = \\u1_u2_adr_cw_reg[11] ;
  assign \new_[2084]_  = \\u1_u2_adr_cw_reg[13] ;
  assign \new_[2085]_  = \\u1_u2_adr_cw_reg[14] ;
  assign \new_[2086]_  = \\u1_u2_adr_cw_reg[5] ;
  assign \new_[2087]_  = \\u1_u2_adr_cw_reg[6] ;
  assign \new_[2088]_  = \\u1_u2_adr_cw_reg[7] ;
  assign \new_[2089]_  = \\u1_u2_adr_cw_reg[8] ;
  assign \new_[2090]_  = \\u1_u2_adr_cw_reg[0] ;
  assign \new_[2091]_  = \\u1_u2_adr_cw_reg[3] ;
  assign \new_[2092]_  = \\u1_u2_adr_cw_reg[2] ;
  assign \new_[2093]_  = \\u1_u2_adr_cw_reg[4] ;
  assign \new_[2094]_  = \\u1_u2_adr_cw_reg[10] ;
  assign \new_[2095]_  = \\u1_u2_adr_cw_reg[12] ;
  assign \new_[2096]_  = \\u1_u2_adr_cw_reg[1] ;
  assign \new_[2097]_  = \\u1_u2_adr_cw_reg[9] ;
  assign n615 = \new_[2140]_  ? n9145 : \new_[13526]_ ;
  assign \new_[2099]_  = \new_[2357]_  ^ \new_[2138]_ ;
  assign \new_[2100]_  = \new_[2466]_  ^ \new_[2139]_ ;
  assign \new_[2101]_  = \new_[4743]_  ^ \new_[2137]_ ;
  assign \new_[2102]_  = ~\new_[2419]_  | ~\new_[2489]_  | ~\new_[14290]_  | ~\new_[2195]_ ;
  assign \new_[2103]_  = ~\new_[2223]_  | (~\new_[2160]_  & ~\new_[2190]_ );
  assign n630 = ~\new_[2230]_  | (~\new_[2162]_  & ~\new_[2204]_ );
  assign n625 = ~\new_[2134]_  | ~\new_[10117]_ ;
  assign \new_[2106]_  = ~\new_[2143]_  & ~\new_[2225]_ ;
  assign n635 = \new_[2164]_  ? n9145 : \new_[13505]_ ;
  assign n620 = \new_[2191]_  | \new_[2142]_ ;
  assign \new_[2109]_  = ~\new_[2141]_  | (~\new_[14359]_  & ~\new_[2324]_ );
  assign n640 = \new_[2166]_  ? n9145 : \new_[14051]_ ;
  assign \new_[2111]_  = \new_[4859]_  ^ \new_[2165]_ ;
  assign \new_[2112]_  = ~\new_[2161]_  & ~\new_[2257]_ ;
  assign \new_[2113]_  = \new_[10362]_  ^ \new_[2170]_ ;
  assign \new_[2114]_  = \\u1_u3_idin_reg[4] ;
  assign TxValid_pad_o = u0_TxValid_reg;
  assign n650 = \new_[2183]_  ? n9145 : \new_[13990]_ ;
  assign \new_[2117]_  = \new_[2298]_  ^ \new_[2181]_ ;
  assign n645 = ~\new_[2168]_  & ~\new_[3393]_ ;
  assign n690 = ~\new_[2144]_  | ~\new_[4490]_ ;
  assign n710 = ~\new_[2145]_  | (~\new_[13330]_  & ~\new_[5774]_ );
  assign n655 = ~\new_[2146]_  | (~\new_[13330]_  & ~\new_[5514]_ );
  assign n715 = ~\new_[2147]_  | (~\new_[13330]_  & ~\new_[5776]_ );
  assign n660 = ~\new_[2148]_  | (~\new_[13330]_  & ~\new_[5777]_ );
  assign n665 = ~\new_[2149]_  | (~\new_[13330]_  & ~\new_[5778]_ );
  assign n720 = ~\new_[2150]_  | (~\new_[13330]_  & ~\new_[5518]_ );
  assign n700 = ~\new_[2151]_  | (~\new_[13330]_  & ~\new_[5519]_ );
  assign n695 = ~\new_[2152]_  | (~\new_[13330]_  & ~\new_[5520]_ );
  assign n705 = ~\new_[2153]_  | (~\new_[13330]_  & ~\new_[5782]_ );
  assign n670 = ~\new_[2154]_  | (~\new_[13330]_  & ~\new_[5783]_ );
  assign n675 = ~\new_[2155]_  | (~\new_[13330]_  & ~\new_[5784]_ );
  assign n680 = ~\new_[2156]_  | (~\new_[13330]_  & ~\new_[5785]_ );
  assign n685 = ~\new_[2157]_  | (~\new_[13330]_  & ~\new_[5525]_ );
  assign n725 = ~\new_[2158]_  | (~\new_[13330]_  & ~\new_[5787]_ );
  assign \new_[2134]_  = (~\new_[7178]_  | ~\new_[13845]_ ) & (~\new_[7436]_  | ~\new_[2189]_ );
  assign \new_[2135]_  = ~\\u1_u1_crc16_reg[6] ;
  assign \new_[2136]_  = \\u1_u3_idin_reg[3] ;
  assign \new_[2137]_  = ~\new_[2185]_  & (~\new_[2245]_  | ~\new_[14632]_ );
  assign \new_[2138]_  = ~\new_[14620]_  | ~\new_[14359]_ ;
  assign \new_[2139]_  = ~\new_[2180]_  | ~\new_[2236]_ ;
  assign \new_[2140]_  = \new_[2295]_  ^ \new_[2194]_ ;
  assign \new_[2141]_  = ~\new_[2388]_  & (~\new_[2203]_  | ~\new_[2420]_ );
  assign \new_[2142]_  = ~\new_[2169]_  & (~\new_[2821]_  | ~\new_[3007]_ );
  assign \new_[2143]_  = ~\new_[2257]_  & (~\new_[2196]_  | ~\new_[2207]_ );
  assign \new_[2144]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[8632]_ ;
  assign \new_[2145]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[8283]_ ;
  assign \new_[2146]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[7871]_ ;
  assign \new_[2147]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[8593]_ ;
  assign \new_[2148]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[8293]_ ;
  assign \new_[2149]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[7282]_ ;
  assign \new_[2150]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[8969]_ ;
  assign \new_[2151]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[8852]_ ;
  assign \new_[2152]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[8668]_ ;
  assign \new_[2153]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[8683]_ ;
  assign \new_[2154]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[8851]_ ;
  assign \new_[2155]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[8680]_ ;
  assign \new_[2156]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[8679]_ ;
  assign \new_[2157]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[8630]_ ;
  assign \new_[2158]_  = ~\new_[13330]_  | ~\new_[14799]_  | ~\new_[9069]_ ;
  assign \new_[2159]_  = ~\new_[2199]_  | ~\new_[2328]_ ;
  assign \new_[2160]_  = ~\new_[2186]_  & (~\new_[2268]_  | ~\new_[7166]_ );
  assign \new_[2161]_  = ~\new_[2187]_  & (~\new_[2252]_  | ~\new_[14681]_ );
  assign \new_[2162]_  = ~\new_[2188]_  & (~\new_[2252]_  | ~\new_[14682]_ );
  assign n730 = \new_[2218]_  ? n9145 : \new_[13523]_ ;
  assign \new_[2164]_  = \new_[2297]_  ^ \new_[14633]_ ;
  assign \new_[2165]_  = ~\new_[2201]_  & (~\new_[2237]_  | ~\new_[14327]_ );
  assign \new_[2166]_  = \new_[2331]_  ^ \new_[2220]_ ;
  assign n735 = \new_[2202]_  & \new_[12158]_ ;
  assign \new_[2168]_  = ~\new_[4491]_  | ~\new_[4013]_  | ~\new_[3632]_  | ~\new_[2208]_ ;
  assign \new_[2169]_  = ~\new_[2744]_  | ~\new_[3002]_  | ~\new_[9945]_  | ~\new_[2239]_ ;
  assign \new_[2170]_  = \new_[14572]_  ? \new_[2270]_  : \new_[2232]_ ;
  assign \new_[2171]_  = ~\\u1_u1_crc16_reg[2] ;
  assign \new_[2172]_  = ~\\u1_u1_crc16_reg[3] ;
  assign \new_[2173]_  = ~\\u1_u1_crc16_reg[4] ;
  assign \new_[2174]_  = \\u1_u1_crc16_reg[7] ;
  assign \new_[2175]_  = \\u1_u1_crc16_reg[9] ;
  assign \new_[2176]_  = \\u1_u1_state_reg[1] ;
  assign \new_[2177]_  = \\u1_u3_idin_reg[2] ;
  assign \new_[2178]_  = \\u1_u3_idin_reg[1] ;
  assign n740 = ~\new_[2206]_  | ~\new_[10117]_ ;
  assign \new_[2180]_  = ~\new_[14632]_  | ~\new_[2264]_ ;
  assign \new_[2181]_  = ~\new_[2242]_  | (~\new_[2240]_  & ~\new_[2274]_ );
  assign n745 = \new_[2221]_  ? \new_[9842]_  : \new_[4694]_ ;
  assign \new_[2183]_  = \new_[2296]_  ^ \new_[14327]_ ;
  assign \new_[2184]_  = \new_[2205]_  | \new_[2293]_ ;
  assign \new_[2185]_  = ~\new_[2335]_  | (~\new_[2236]_  & ~\new_[2368]_ );
  assign \new_[2186]_  = ~\new_[2268]_  & ~\new_[2448]_ ;
  assign \new_[2187]_  = ~\new_[7168]_  & ~\new_[2238]_ ;
  assign \new_[2188]_  = ~\new_[7172]_  & ~\new_[2238]_ ;
  assign \new_[2189]_  = \new_[12676]_  ^ \new_[14607]_ ;
  assign \new_[2190]_  = ~\new_[2207]_ ;
  assign \new_[2191]_  = \new_[2239]_  & \new_[2530]_ ;
  assign \new_[2192]_  = u1_u1_tx_valid_r_reg;
  assign \new_[2193]_  = \\u1_u1_state_reg[0] ;
  assign \new_[2194]_  = ~\new_[14360]_ ;
  assign \new_[2195]_  = ~\new_[2294]_  | ~\new_[2244]_  | ~\new_[2254]_ ;
  assign \new_[2196]_  = (~\new_[2252]_  | ~\new_[14269]_ ) & (~\new_[2268]_  | ~\new_[6753]_ );
  assign \new_[2197]_  = (~\new_[2252]_  | ~\new_[14271]_ ) & (~\new_[2268]_  | ~\new_[5030]_ );
  assign \new_[2198]_  = (~\new_[2252]_  | ~\new_[14272]_ ) & (~\new_[2268]_  | ~\new_[4706]_ );
  assign \new_[2199]_  = (~\new_[2252]_  | ~\new_[14407]_ ) & (~\new_[2268]_  | ~\new_[5031]_ );
  assign \new_[2200]_  = (~\new_[2252]_  | ~\new_[14402]_ ) & (~\new_[2268]_  | ~\new_[4710]_ );
  assign \new_[2201]_  = ~\new_[2299]_  | (~\new_[14438]_  & ~\new_[2387]_ );
  assign \new_[2202]_  = ~\new_[9587]_  | ~\new_[9521]_  | ~\new_[2234]_  | ~\new_[2406]_ ;
  assign \new_[2203]_  = ~\new_[2326]_  | (~\new_[14620]_  & ~\new_[2358]_ );
  assign \new_[2204]_  = ~\new_[2223]_ ;
  assign \new_[2205]_  = ~\new_[2242]_  & ~\new_[2308]_ ;
  assign \new_[2206]_  = (~\new_[7178]_  | ~\new_[13817]_ ) & (~\new_[7436]_  | ~\new_[2262]_ );
  assign \new_[2207]_  = \new_[2252]_  | \new_[7939]_ ;
  assign \new_[2208]_  = ~\new_[2251]_  & ~\new_[6874]_ ;
  assign \new_[2209]_  = ~\\u1_u1_crc16_reg[5] ;
  assign \new_[2210]_  = \\u1_u1_state_reg[4] ;
  assign n775 = ~\new_[12804]_  & (~\new_[9639]_  | ~\new_[2261]_ );
  assign n750 = ~\new_[2243]_  | ~\new_[10117]_ ;
  assign n755 = ~\new_[2247]_  | ~\new_[10117]_ ;
  assign n760 = ~\new_[2248]_  | ~\new_[10117]_ ;
  assign n765 = ~\new_[2249]_  | ~\new_[10117]_ ;
  assign n770 = ~\new_[2250]_  | ~\new_[10117]_ ;
  assign n780 = \new_[2255]_  ? \new_[9842]_  : \new_[4228]_ ;
  assign \new_[2218]_  = \new_[2360]_  ^ \new_[14300]_ ;
  assign n785 = ~\new_[2256]_  | ~\new_[9196]_  | ~\new_[9289]_ ;
  assign \new_[2220]_  = ~\new_[2240]_ ;
  assign \new_[2221]_  = \new_[2329]_  ^ \new_[14319]_ ;
  assign n790 = u1_u1_tx_valid_r1_reg;
  assign \new_[2223]_  = ~\new_[2257]_  & ~\new_[2307]_ ;
  assign \new_[2224]_  = ~\DataOut_pad_o[1]  | ~\new_[2257]_  | ~\new_[11651]_ ;
  assign \new_[2225]_  = ~\new_[2257]_  & ~\new_[2328]_ ;
  assign \new_[2226]_  = ~\DataOut_pad_o[2]  | ~\new_[2257]_  | ~\new_[11651]_ ;
  assign \new_[2227]_  = ~\DataOut_pad_o[3]  | ~\new_[2257]_  | ~\new_[11651]_ ;
  assign \new_[2228]_  = ~\DataOut_pad_o[4]  | ~\new_[2257]_  | ~\new_[11651]_ ;
  assign \new_[2229]_  = ~\DataOut_pad_o[0]  | ~\new_[2257]_  | ~\new_[11651]_ ;
  assign \new_[2230]_  = ~\DataOut_pad_o[5]  | ~\new_[2257]_  | ~\new_[11651]_ ;
  assign \new_[2231]_  = ~\DataOut_pad_o[6]  | ~\new_[2257]_  | ~\new_[11651]_ ;
  assign \new_[2232]_  = ~\new_[14572]_ ;
  assign \new_[2233]_  = ~\DataOut_pad_o[7]  | ~\new_[2257]_  | ~\new_[11651]_ ;
  assign \new_[2234]_  = ~n810 & ~n8245;
  assign n795 = ~\new_[9828]_  | ~\new_[9825]_  | ~\new_[13165]_  | ~\new_[2275]_ ;
  assign \new_[2236]_  = \new_[2260]_  & \new_[2326]_ ;
  assign \new_[2237]_  = ~\new_[2263]_  & ~\new_[2387]_ ;
  assign \new_[2238]_  = ~\new_[2268]_  | ~\new_[7939]_ ;
  assign \new_[2239]_  = \new_[2269]_  & \new_[2375]_ ;
  assign \new_[2240]_  = ~\new_[2254]_ ;
  assign n805 = ~\new_[12849]_  & (~\new_[9832]_  | ~\new_[2288]_ );
  assign \new_[2242]_  = ~\new_[2292]_  & (~\new_[2290]_  | ~\new_[2309]_ );
  assign \new_[2243]_  = (~\new_[7178]_  | ~\new_[13844]_ ) & (~\new_[7436]_  | ~\new_[2280]_ );
  assign \new_[2244]_  = ~\new_[2417]_  & ~\new_[2274]_ ;
  assign \new_[2245]_  = ~\new_[2273]_  & ~\new_[2368]_ ;
  assign \new_[2246]_  = ~\new_[2263]_ ;
  assign \new_[2247]_  = (~\new_[7178]_  | ~\new_[13977]_ ) & (~\new_[7436]_  | ~\new_[2282]_ );
  assign \new_[2248]_  = (~\new_[7178]_  | ~\new_[13823]_ ) & (~\new_[7436]_  | ~\new_[2284]_ );
  assign \new_[2249]_  = (~\new_[7178]_  | ~\new_[2174]_ ) & (~\new_[7436]_  | ~\new_[2289]_ );
  assign \new_[2250]_  = (~\new_[7178]_  | ~\new_[2175]_ ) & (~\new_[7436]_  | ~\new_[2291]_ );
  assign \new_[2251]_  = \new_[2755]_  | \new_[13520]_  | \new_[2749]_  | \new_[2302]_ ;
  assign \new_[2252]_  = ~\new_[2268]_ ;
  assign n800 = ~\new_[2276]_  | ~\new_[10117]_ ;
  assign \new_[2254]_  = ~\new_[2279]_  | ~\new_[2306]_  | ~\new_[2285]_ ;
  assign \new_[2255]_  = \new_[14692]_  ^ \new_[2330]_ ;
  assign \new_[2256]_  = \new_[2283]_  | \new_[9842]_ ;
  assign \new_[2257]_  = ~TxReady_pad_i & (~\new_[2305]_  | ~n840);
  assign \new_[2258]_  = ~\new_[14629]_  & (~\new_[14364]_  | ~\new_[14366]_ );
  assign n810 = ~\new_[10847]_  | ~\new_[11153]_  | ~\new_[2287]_  | ~\new_[11818]_ ;
  assign \new_[2260]_  = ~\new_[14628]_  | ~\new_[14651]_ ;
  assign \new_[2261]_  = ~\new_[10074]_  & (~\new_[11206]_  | ~\new_[2310]_ );
  assign \new_[2262]_  = \new_[14307]_  ^ \new_[2320]_ ;
  assign \new_[2263]_  = ~\new_[2294]_  | ~\new_[2309]_ ;
  assign \new_[2264]_  = ~\new_[2273]_ ;
  assign \new_[2265]_  = \\u1_u3_idin_reg[30] ;
  assign \new_[2266]_  = \\u1_u3_idin_reg[0] ;
  assign \new_[2267]_  = u1_u1_send_token_r_reg;
  assign \new_[2268]_  = ~\new_[9400]_  | ~\new_[11051]_  | ~\new_[2287]_  | ~\new_[11490]_ ;
  assign \new_[2269]_  = ~\new_[2302]_  & ~\new_[13520]_ ;
  assign \new_[2270]_  = ~\new_[2311]_  | ~\new_[2312]_ ;
  assign \new_[2271]_  = ~\new_[2314]_  | ~\new_[2337]_ ;
  assign \new_[2272]_  = ~\new_[14366]_  | ~\new_[14362]_ ;
  assign \new_[2273]_  = ~\new_[14651]_  | ~\new_[14630]_ ;
  assign \new_[2274]_  = ~\new_[14379]_  | ~\new_[2309]_ ;
  assign \new_[2275]_  = ~\new_[13443]_  | ~\new_[2310]_  | ~\new_[2193]_ ;
  assign \new_[2276]_  = (~\new_[7178]_  | ~\new_[14146]_ ) & (~\new_[7436]_  | ~\new_[2323]_ );
  assign \new_[2277]_  = ~\new_[14462]_  | ~\new_[2038]_ ;
  assign \new_[2278]_  = u1_u1_zero_length_r_reg;
  assign \new_[2279]_  = ~\new_[14689]_  | ~\new_[2322]_  | ~\new_[14512]_ ;
  assign \new_[2280]_  = \new_[12645]_  ^ \new_[2379]_ ;
  assign n820 = ~\new_[8950]_  | (~\new_[2361]_  & ~\new_[9842]_ );
  assign \new_[2282]_  = \new_[12903]_  ^ \new_[2381]_ ;
  assign \new_[2283]_  = \new_[14318]_  ^ \new_[2359]_ ;
  assign \new_[2284]_  = \new_[13169]_  ^ \new_[2380]_ ;
  assign \new_[2285]_  = ~\new_[14320]_  | ~\new_[14512]_ ;
  assign n825 = ~\new_[12732]_  & (~\new_[10252]_  | ~\new_[2406]_ );
  assign \new_[2287]_  = ~\new_[10870]_  & ~\new_[2327]_ ;
  assign \new_[2288]_  = ~\new_[10500]_  & ~\new_[2327]_ ;
  assign \new_[2289]_  = \new_[14602]_  ^ \new_[2353]_ ;
  assign \new_[2290]_  = ~\new_[2364]_  | (~\new_[2367]_  & ~\new_[2410]_ );
  assign \new_[2291]_  = \new_[2038]_  ^ \new_[2354]_ ;
  assign \new_[2292]_  = ~\new_[14622]_  | (~\new_[2365]_  & ~\new_[2366]_ );
  assign \new_[2293]_  = ~\new_[2428]_  | (~\new_[14652]_  & ~\new_[14627]_ );
  assign \new_[2294]_  = ~\new_[2308]_ ;
  assign \new_[2295]_  = ~\new_[2364]_  | ~\new_[2334]_ ;
  assign \new_[2296]_  = ~\new_[2332]_  & ~\new_[2363]_ ;
  assign \new_[2297]_  = ~\new_[2333]_  & ~\new_[2366]_ ;
  assign \new_[2298]_  = ~\new_[14623]_  & ~\new_[14626]_ ;
  assign \new_[2299]_  = (~\new_[2469]_  | ~\new_[4858]_ ) & (~\new_[2369]_  | ~\new_[2433]_ );
  assign \new_[2300]_  = ~\new_[14761]_  | ~\new_[14077]_ ;
  assign \new_[2301]_  = \\u1_u3_state_reg[0] ;
  assign \new_[2302]_  = ~\new_[3005]_  | ~\new_[2352]_ ;
  assign n815 = ~\new_[2352]_  & ~n9145;
  assign n830 = ~\new_[9183]_  & (~\new_[9567]_  | ~\new_[2382]_ );
  assign \new_[2305]_  = ~u1_u1_tx_first_r_reg;
  assign \new_[2306]_  = ~\new_[2325]_ ;
  assign \new_[2307]_  = ~\new_[2328]_ ;
  assign \new_[2308]_  = \new_[14652]_  | \new_[14623]_ ;
  assign \new_[2309]_  = ~\new_[2363]_  & ~\new_[2366]_ ;
  assign \new_[2310]_  = ~\new_[11513]_  & ~\new_[2362]_ ;
  assign \new_[2311]_  = ~\new_[2379]_  | ~\new_[14796]_ ;
  assign \new_[2312]_  = ~\new_[14406]_  | ~\new_[2380]_ ;
  assign \new_[2313]_  = \new_[2389]_  ^ \new_[8293]_ ;
  assign \new_[2314]_  = ~\new_[2380]_  | ~\new_[14399]_ ;
  assign \new_[2315]_  = ~\new_[7283]_  | ~\new_[2370]_ ;
  assign \new_[2316]_  = \\u1_u2_sizd_c_reg[10] ;
  assign \new_[2317]_  = \\u1_u2_sizd_c_reg[12] ;
  assign \new_[2318]_  = \\u1_u2_sizd_c_reg[4] ;
  assign \dma_req_o[1]  = u4_u1_dma_req_r_reg;
  assign \new_[2320]_  = ~\new_[14794]_ ;
  assign n835 = ~\new_[2430]_  | ~\new_[9491]_  | ~\new_[3105]_  | ~\new_[4971]_ ;
  assign \new_[2322]_  = ~\new_[2355]_ ;
  assign \new_[2323]_  = \new_[13241]_  ^ \new_[2426]_ ;
  assign \new_[2324]_  = ~\new_[14651]_  | ~\new_[2420]_ ;
  assign \new_[2325]_  = ~\new_[2427]_  | (~\new_[14697]_  & ~\new_[14667]_ );
  assign \new_[2326]_  = ~\new_[2383]_  & ~\new_[2488]_ ;
  assign \new_[2327]_  = ~\new_[11513]_  & ~\new_[2385]_ ;
  assign \new_[2328]_  = ~\new_[2267]_  & ~\new_[2384]_ ;
  assign \new_[2329]_  = ~\new_[14697]_  | ~\new_[14690]_ ;
  assign \new_[2330]_  = \new_[14378]_  & \new_[14689]_ ;
  assign \new_[2331]_  = ~\new_[14444]_  & ~\new_[2386]_ ;
  assign \new_[2332]_  = ~\new_[2365]_ ;
  assign \new_[2333]_  = ~\new_[14622]_ ;
  assign \new_[2334]_  = ~\new_[2367]_ ;
  assign \new_[2335]_  = ~\new_[2388]_  | ~\new_[13376]_ ;
  assign \new_[2336]_  = ~\new_[14406]_  | ~\new_[14405]_ ;
  assign \new_[2337]_  = ~\new_[14796]_  | ~\new_[14407]_ ;
  assign \new_[2338]_  = ~\new_[7282]_  | ~\new_[2390]_ ;
  assign \new_[2339]_  = \\u1_u2_sizd_c_reg[0] ;
  assign \new_[2340]_  = \\u1_u2_sizd_c_reg[11] ;
  assign \new_[2341]_  = \\u1_u2_sizd_c_reg[13] ;
  assign \new_[2342]_  = \\u1_u2_sizd_c_reg[1] ;
  assign \new_[2343]_  = \\u1_u2_sizd_c_reg[2] ;
  assign \new_[2344]_  = \\u1_u2_sizd_c_reg[3] ;
  assign \new_[2345]_  = \\u1_u2_sizd_c_reg[5] ;
  assign \new_[2346]_  = \\u1_u2_sizd_c_reg[6] ;
  assign \new_[2347]_  = \\u1_u2_sizd_c_reg[7] ;
  assign \new_[2348]_  = \\u1_u2_sizd_c_reg[8] ;
  assign \new_[2349]_  = \\u1_u2_sizd_c_reg[9] ;
  assign \dma_req_o[2]  = u4_u2_dma_req_r_reg;
  assign \dma_req_o[0]  = u4_u0_dma_req_r_reg;
  assign \new_[2352]_  = ~\\u1_u3_new_size_reg[13] ;
  assign \new_[2353]_  = \new_[14271]_  ^ \new_[14269]_ ;
  assign \new_[2354]_  = \new_[13561]_  ^ \new_[2448]_ ;
  assign \new_[2355]_  = ~\new_[14318]_  | ~\new_[2407]_ ;
  assign n840 = ~\new_[2406]_  | ~\new_[13443]_ ;
  assign \new_[2357]_  = ~\new_[2411]_  & ~\new_[14652]_ ;
  assign \new_[2358]_  = ~\new_[14651]_ ;
  assign \new_[2359]_  = ~\new_[2407]_  | ~\new_[2408]_ ;
  assign \new_[2360]_  = ~\new_[2427]_  | ~\new_[2409]_ ;
  assign \new_[2361]_  = \new_[5075]_  ^ \new_[2431]_ ;
  assign \new_[2362]_  = ~\new_[2385]_ ;
  assign \new_[2363]_  = ~\new_[2414]_  & ~\new_[4861]_ ;
  assign \new_[2364]_  = ~\new_[2415]_  | ~\new_[4860]_ ;
  assign \new_[2365]_  = ~\new_[2414]_  | ~\new_[4861]_ ;
  assign \new_[2366]_  = ~\new_[2416]_  & ~\new_[4862]_ ;
  assign \new_[2367]_  = ~\new_[2415]_  & ~\new_[4860]_ ;
  assign \new_[2368]_  = ~\new_[2420]_  | ~\new_[13376]_ ;
  assign \new_[2369]_  = \new_[2418]_  | \new_[2514]_ ;
  assign \new_[2370]_  = ~\new_[2390]_ ;
  assign \dma_req_o[3]  = u4_u3_dma_req_r_reg;
  assign \new_[2372]_  = \\u1_u3_state_reg[1] ;
  assign \new_[2373]_  = \\u1_u3_state_reg[4] ;
  assign n860 = ~\new_[2425]_  | (~\new_[11679]_  & ~\new_[10668]_ );
  assign \new_[2375]_  = ~\new_[2753]_  & (~\new_[2434]_  | ~\new_[2754]_ );
  assign n850 = ~\new_[2423]_  | ~\new_[12100]_ ;
  assign n845 = ~\new_[2421]_  | ~\new_[13165]_ ;
  assign n855 = ~\new_[2422]_  | ~\new_[13165]_ ;
  assign \new_[2379]_  = ~\new_[14406]_ ;
  assign \new_[2380]_  = ~\new_[14796]_ ;
  assign \new_[2381]_  = \new_[14682]_  ^ \new_[14407]_ ;
  assign \new_[2382]_  = \new_[2432]_  | \new_[10117]_ ;
  assign \new_[2383]_  = ~\new_[2428]_  & ~\new_[14653]_ ;
  assign \new_[2384]_  = ~\new_[2406]_ ;
  assign \new_[2385]_  = \new_[2432]_  | \new_[13443]_ ;
  assign \new_[2386]_  = ~\new_[2410]_ ;
  assign \new_[2387]_  = ~\new_[2435]_  | ~\new_[2433]_ ;
  assign \new_[2388]_  = ~\new_[2436]_  | ~\new_[2489]_ ;
  assign \new_[2389]_  = \\u1_u2_last_buf_adr_reg[13] ;
  assign \new_[2390]_  = \\u1_u2_last_buf_adr_reg[14] ;
  assign \new_[2391]_  = \new_[2470]_  ^ \new_[8283]_ ;
  assign \new_[2392]_  = \\u1_u3_state_reg[2] ;
  assign n920 = ~\new_[2459]_  | (~\new_[11672]_  & ~\new_[10631]_ );
  assign n925 = ~\new_[2460]_  | (~\new_[11708]_  & ~\new_[10667]_ );
  assign n865 = ~\new_[2437]_  | ~\new_[13165]_ ;
  assign n870 = ~\new_[2446]_  | ~\new_[12067]_ ;
  assign n875 = ~\new_[2447]_  | ~\new_[12100]_ ;
  assign n885 = ~\new_[2438]_  | ~rst_i;
  assign n890 = ~\new_[2439]_  | ~rst_i;
  assign n895 = ~\new_[2440]_  | ~\new_[13165]_ ;
  assign n900 = ~\new_[2444]_  | ~\new_[13165]_ ;
  assign n905 = ~\new_[2441]_  | ~\new_[13165]_ ;
  assign n910 = ~\new_[2442]_  | ~\new_[13165]_ ;
  assign n915 = ~\new_[2443]_  | ~rst_i;
  assign n930 = \new_[2467]_  ^ \new_[3066]_ ;
  assign \new_[2406]_  = ~u1_u3_send_token_reg;
  assign \new_[2407]_  = \new_[14608]_  | \new_[5249]_ ;
  assign \new_[2408]_  = ~\new_[14608]_  | ~\new_[5249]_ ;
  assign \new_[2409]_  = ~\new_[14667]_ ;
  assign \new_[2410]_  = ~\new_[14445]_  | ~\new_[5248]_ ;
  assign \new_[2411]_  = ~\new_[2428]_ ;
  assign n945 = ~\new_[14417]_  & (~\new_[4972]_  | ~\new_[2487]_ );
  assign n940 = ~\new_[14417]_  & (~\new_[5367]_  | ~\new_[2485]_ );
  assign \new_[2414]_  = ~\new_[9282]_  | ~\new_[10034]_  | ~\new_[2496]_ ;
  assign \new_[2415]_  = ~\new_[9274]_  | ~\new_[10036]_  | ~\new_[2497]_ ;
  assign \new_[2416]_  = ~\new_[9529]_  | ~\new_[10044]_  | ~\new_[2498]_ ;
  assign \new_[2417]_  = ~\new_[2435]_ ;
  assign \new_[2418]_  = ~\new_[2468]_  & ~\new_[2515]_ ;
  assign \new_[2419]_  = ~\new_[14292]_  & ~n9145;
  assign \new_[2420]_  = ~\new_[14292]_  & ~\new_[2515]_ ;
  assign \new_[2421]_  = ~\new_[2461]_  & (~\new_[8764]_  | ~\new_[14499]_ );
  assign \new_[2422]_  = ~\new_[2463]_  & (~\new_[8775]_  | ~\new_[14499]_ );
  assign \new_[2423]_  = ~\new_[2462]_  & (~\new_[7747]_  | ~\new_[14499]_ );
  assign n935 = ~\new_[2481]_  | (~\new_[11575]_  & ~\new_[10653]_ );
  assign \new_[2425]_  = ~\new_[11616]_  & (~\new_[2482]_  | ~\new_[13162]_ );
  assign \new_[2426]_  = \new_[14681]_  ^ \new_[14272]_ ;
  assign \new_[2427]_  = ~\new_[14668]_  | ~\new_[4515]_ ;
  assign \new_[2428]_  = ~\new_[2483]_  | ~\new_[4512]_ ;
  assign n960 = ~\new_[14417]_  & (~\new_[5376]_  | ~\new_[2508]_ );
  assign \new_[2430]_  = ~\new_[2484]_  & (~\new_[10376]_  | ~\new_[3243]_ );
  assign \new_[2431]_  = ~\new_[2464]_ ;
  assign \new_[2432]_  = ~u1_u1_send_zero_length_r_reg;
  assign \new_[2433]_  = \new_[14289]_  & \new_[4858]_ ;
  assign \new_[2434]_  = ~\new_[2521]_  | ~\new_[2610]_  | ~\new_[2886]_ ;
  assign \new_[2435]_  = ~\new_[14653]_  & ~\new_[2515]_ ;
  assign \new_[2436]_  = ~\new_[2514]_  | ~\new_[14289]_ ;
  assign \new_[2437]_  = \new_[2798]_  ? \new_[14499]_  : \new_[8720]_ ;
  assign \new_[2438]_  = \new_[2732]_  ? \new_[14499]_  : \new_[8338]_ ;
  assign \new_[2439]_  = \new_[2733]_  ? \new_[14499]_  : \new_[8358]_ ;
  assign \new_[2440]_  = \new_[2736]_  ? \new_[14499]_  : \new_[8371]_ ;
  assign \new_[2441]_  = \new_[2739]_  ? \new_[14499]_  : \new_[8379]_ ;
  assign \new_[2442]_  = \new_[2740]_  ? \new_[14499]_  : \new_[7964]_ ;
  assign \new_[2443]_  = \new_[2742]_  ? \new_[14499]_  : \new_[7731]_ ;
  assign \new_[2444]_  = \new_[2738]_  ? \new_[14499]_  : \new_[8403]_ ;
  assign n950 = \new_[4263]_  ^ \new_[2522]_ ;
  assign \new_[2446]_  = \new_[2818]_  ? \new_[14499]_  : \new_[7173]_ ;
  assign \new_[2447]_  = \new_[2820]_  ? \new_[14499]_  : \new_[7174]_ ;
  assign \new_[2448]_  = ~\new_[14309]_ ;
  assign \new_[2449]_  = \new_[2523]_  ^ \new_[9069]_ ;
  assign n955 = \new_[5776]_  ^ \new_[2528]_ ;
  assign \new_[2451]_  = \new_[2527]_  ^ \new_[7871]_ ;
  assign \new_[2452]_  = \\u1_u3_state_reg[8] ;
  assign \new_[2453]_  = u1_u2_send_zero_length_r_reg;
  assign \new_[2454]_  = u1_u2_rx_dma_en_r_reg;
  assign \new_[2455]_  = ~\\u1_u3_new_sizeb_reg[6] ;
  assign \new_[2456]_  = ~\\u1_u3_new_sizeb_reg[7] ;
  assign \new_[2457]_  = ~\\u1_u3_new_sizeb_reg[8] ;
  assign \new_[2458]_  = ~\\u1_u3_new_sizeb_reg[9] ;
  assign \new_[2459]_  = ~\new_[11728]_  & (~\new_[2506]_  | ~\new_[13162]_ );
  assign \new_[2460]_  = ~\new_[11608]_  & (~\new_[2507]_  | ~\new_[13162]_ );
  assign \new_[2461]_  = ~\new_[14499]_  & ~\new_[2797]_ ;
  assign \new_[2462]_  = ~\new_[14499]_  & ~\new_[2819]_ ;
  assign \new_[2463]_  = ~\new_[14499]_  & ~\new_[2800]_ ;
  assign \new_[2464]_  = ~\new_[10035]_  & (~\new_[2542]_  | ~\new_[14833]_ );
  assign n965 = ~\new_[2572]_  | ~\new_[3358]_  | ~\new_[2540]_ ;
  assign \new_[2466]_  = ~\new_[2514]_  & ~\new_[2515]_ ;
  assign \new_[2467]_  = \new_[2544]_  ^ \new_[14275]_ ;
  assign \new_[2468]_  = ~\new_[2488]_ ;
  assign \new_[2469]_  = ~\new_[2489]_ ;
  assign \new_[2470]_  = ~\\u1_u2_last_buf_adr_reg[10] ;
  assign \new_[2471]_  = ~\\u1_u3_new_sizeb_reg[0] ;
  assign \new_[2472]_  = ~\\u1_u3_new_sizeb_reg[1] ;
  assign \new_[2473]_  = ~\\u1_u3_new_sizeb_reg[2] ;
  assign \new_[2474]_  = ~\\u1_u3_new_sizeb_reg[3] ;
  assign \new_[2475]_  = ~\\u1_u3_new_sizeb_reg[5] ;
  assign \new_[2476]_  = \\u1_u3_state_reg[3] ;
  assign \new_[2477]_  = \\u1_u3_state_reg[5] ;
  assign \new_[2478]_  = \\u1_u3_state_reg[6] ;
  assign \new_[2479]_  = \\u1_u3_state_reg[7] ;
  assign n8990 = \\u1_u3_state_reg[9] ;
  assign \new_[2481]_  = ~\new_[11572]_  & (~\new_[2531]_  | ~\new_[13162]_ );
  assign \new_[2482]_  = ~\new_[9155]_  | ~\new_[2532]_ ;
  assign \new_[2483]_  = ~\new_[9522]_  | (~\new_[2560]_  & ~\new_[14829]_ );
  assign \new_[2484]_  = ~\new_[2539]_  | (~\new_[4667]_  & ~\new_[10801]_ );
  assign \new_[2485]_  = ~\new_[2541]_  & (~\new_[9779]_  | ~\new_[2852]_ );
  assign n975 = ~\new_[14417]_  & (~\new_[2848]_  | ~\new_[2562]_ );
  assign \new_[2487]_  = ~\new_[4959]_  & (~\new_[2563]_  | ~\new_[11106]_ );
  assign \new_[2488]_  = \new_[14654]_  & \new_[4857]_ ;
  assign \new_[2489]_  = ~\new_[2546]_  | ~\new_[4513]_ ;
  assign n980 = ~\new_[8937]_  & ~\new_[2545]_ ;
  assign n985 = ~\new_[2545]_  & ~\new_[8930]_ ;
  assign n990 = ~\new_[9274]_  | ~\new_[10036]_  | ~\new_[2568]_ ;
  assign n995 = ~\new_[9282]_  | ~\new_[10034]_  | ~\new_[2569]_ ;
  assign n1000 = ~\new_[9529]_  | ~\new_[10044]_  | ~\new_[2570]_ ;
  assign n1005 = ~\new_[14408]_  | ~\new_[14337]_  | ~\new_[2571]_ ;
  assign \new_[2496]_  = ~\new_[10116]_  | ~\new_[14833]_  | ~\new_[2564]_ ;
  assign \new_[2497]_  = ~\new_[10116]_  | ~\new_[14833]_  | ~\new_[2565]_ ;
  assign \new_[2498]_  = ~\new_[10116]_  | ~\new_[14833]_  | ~\new_[2566]_ ;
  assign \new_[2499]_  = \\u1_u2_last_buf_adr_reg[12] ;
  assign \new_[2500]_  = \\u4_u2_int_stat_reg[2] ;
  assign \new_[2501]_  = \\u4_u3_int_stat_reg[2] ;
  assign \new_[2502]_  = \\u4_u0_int_stat_reg[2] ;
  assign \new_[2503]_  = ~\\u1_u3_new_sizeb_reg[4] ;
  assign \new_[2504]_  = \\u4_u1_int_stat_reg[2] ;
  assign \new_[2505]_  = ~\\u1_u3_new_sizeb_reg[10] ;
  assign \new_[2506]_  = ~\new_[9148]_  | ~\new_[2556]_ ;
  assign \new_[2507]_  = ~\new_[9153]_  | ~\new_[2557]_ ;
  assign \new_[2508]_  = \new_[2559]_  | \new_[10806]_ ;
  assign n1015 = \new_[2558]_  | \new_[10035]_ ;
  assign n1020 = ~\new_[14612]_  | (~\new_[2591]_  & ~\new_[9834]_ );
  assign n1025 = ~\new_[14831]_  | (~\new_[2592]_  & ~\new_[9834]_ );
  assign n1030 = ~\new_[14516]_  | (~\new_[2593]_  & ~\new_[9834]_ );
  assign n1035 = ~\new_[14447]_  | (~\new_[2594]_  & ~\new_[9834]_ );
  assign \new_[2514]_  = ~\new_[2561]_  & ~\new_[4742]_ ;
  assign \new_[2515]_  = \new_[2561]_  & \new_[4742]_ ;
  assign n1045 = ~\new_[14417]_  & (~\new_[2601]_  | ~\new_[4924]_ );
  assign n1050 = ~\new_[14417]_  & (~\new_[10042]_  | ~\new_[2602]_ );
  assign n1055 = ~\new_[14417]_  & (~\new_[2603]_  | ~\new_[4925]_ );
  assign n1060 = ~\new_[14417]_  & (~\new_[2604]_  | ~\new_[10755]_ );
  assign n1040 = ~\new_[14417]_  & (~\new_[2600]_  | ~\new_[4159]_ );
  assign \new_[2521]_  = (~\new_[3058]_  | ~\new_[2607]_ ) & (~\new_[2889]_  | ~\new_[2607]_ );
  assign \new_[2522]_  = ~\new_[2612]_  | ~\new_[5100]_  | ~\new_[3077]_ ;
  assign \new_[2523]_  = ~\\u1_u2_last_buf_adr_reg[9] ;
  assign \new_[2524]_  = u1_u2_tx_dma_en_r_reg;
  assign \new_[2525]_  = \new_[2613]_  ^ \new_[8630]_ ;
  assign \new_[2526]_  = \new_[2614]_  ^ \new_[8680]_ ;
  assign \new_[2527]_  = ~\\u1_u2_last_buf_adr_reg[11] ;
  assign \new_[2528]_  = ~\new_[3556]_  & (~\new_[3804]_  | ~\new_[14487]_ );
  assign n1010 = \new_[4262]_  ^ \new_[14487]_ ;
  assign \new_[2530]_  = ~\new_[2607]_  | ~\new_[2754]_  | ~\new_[2824]_ ;
  assign \new_[2531]_  = ~\new_[9149]_  | ~\new_[2582]_ ;
  assign \new_[2532]_  = ~\new_[13251]_  | ~\dma_req_o[1]  | ~\new_[2583]_  | ~\new_[9179]_ ;
  assign n1070 = ~\new_[2585]_  & ~\new_[7411]_ ;
  assign n1075 = ~\new_[2586]_  & ~\new_[8124]_ ;
  assign n1080 = ~\new_[2587]_  & ~\new_[7414]_ ;
  assign n1090 = ~\new_[2588]_  & ~\new_[7418]_ ;
  assign n1095 = ~\new_[9522]_  | (~\new_[2628]_  & ~\new_[9834]_ );
  assign n1085 = ~\new_[14672]_  | (~\new_[2629]_  & ~\new_[9834]_ );
  assign \new_[2539]_  = (~\new_[2627]_  | ~\new_[10041]_ ) & (~\new_[10365]_  | ~\new_[2852]_ );
  assign \new_[2540]_  = \new_[2590]_  | \new_[11024]_ ;
  assign \new_[2541]_  = ~\new_[10806]_  & (~\new_[2634]_  | ~\new_[2725]_ );
  assign \new_[2542]_  = ~\new_[2589]_  | ~\new_[9821]_ ;
  assign \new_[2543]_  = ~\new_[9558]_  & (~\new_[2631]_  | ~\new_[14834]_ );
  assign \new_[2544]_  = ~\\u1_u3_new_sizeb_reg[13] ;
  assign \new_[2545]_  = \new_[11775]_  | \new_[2852]_  | \new_[8134]_  | \new_[12680]_ ;
  assign \new_[2546]_  = ~\new_[2596]_  & ~\new_[9834]_ ;
  assign \new_[2547]_  = \\u1_u3_idin_reg[27] ;
  assign \new_[2548]_  = u4_dma_out_buf_avail_reg;
  assign \new_[2549]_  = ~\\u1_u3_new_sizeb_reg[11] ;
  assign \new_[2550]_  = ~\\u1_u3_new_sizeb_reg[12] ;
  assign \new_[2551]_  = \\u4_u2_int_stat_reg[5] ;
  assign \new_[2552]_  = \\u4_u3_int_stat_reg[5] ;
  assign \new_[2553]_  = \\u4_u0_int_stat_reg[5] ;
  assign \new_[2554]_  = \\u4_u1_int_stat_reg[5] ;
  assign n1065 = \new_[4457]_  ^ \new_[2672]_ ;
  assign \new_[2556]_  = ~\new_[13040]_  | ~\dma_req_o[2]  | ~\new_[2620]_  | ~\new_[9178]_ ;
  assign \new_[2557]_  = ~\new_[13124]_  | ~\dma_req_o[0]  | ~\new_[2621]_  | ~\new_[8929]_ ;
  assign \new_[2558]_  = ~\new_[9834]_  & (~\new_[2724]_  | ~\new_[9821]_ );
  assign \new_[2559]_  = (~\new_[2722]_  | ~\new_[7762]_ ) & (~\new_[2852]_  | ~\new_[2392]_ );
  assign \new_[2560]_  = ~\new_[9560]_  & (~\new_[2720]_  | ~\new_[14834]_ );
  assign \new_[2561]_  = ~\new_[9036]_  | ~\new_[9610]_  | ~\new_[2727]_ ;
  assign \new_[2562]_  = (~\new_[4668]_  | ~\new_[7208]_ ) & (~\new_[9500]_  | ~\new_[2852]_ );
  assign \new_[2563]_  = ~\new_[2635]_  & (~\new_[7415]_  | ~\new_[2923]_ );
  assign \new_[2564]_  = \\u1_u3_size_next_r_reg[7] ;
  assign \new_[2565]_  = \\u1_u3_size_next_r_reg[6] ;
  assign \new_[2566]_  = \\u1_u3_size_next_r_reg[8] ;
  assign \new_[2567]_  = \\u1_u3_size_next_r_reg[9] ;
  assign \new_[2568]_  = ~n1165 | ~\new_[8257]_ ;
  assign \new_[2569]_  = ~n1160 | ~\new_[8257]_ ;
  assign \new_[2570]_  = ~n1170 | ~\new_[8257]_ ;
  assign \new_[2571]_  = ~n1175 | ~\new_[8257]_ ;
  assign \new_[2572]_  = ~\new_[12680]_  | ~\new_[2923]_  | ~\new_[10725]_ ;
  assign \new_[2573]_  = \\u4_int_srcb_reg[2] ;
  assign n1100 = \new_[4269]_  ^ \new_[14517]_ ;
  assign n1110 = \new_[4456]_  ^ \new_[2752]_ ;
  assign \new_[2576]_  = ~\new_[2694]_  | ~\new_[2678]_ ;
  assign \new_[2577]_  = ~\new_[2696]_  | ~\new_[2695]_ ;
  assign \new_[2578]_  = ~\new_[2709]_  | ~\new_[2683]_ ;
  assign \new_[2579]_  = ~\new_[2708]_  | ~\new_[2710]_ ;
  assign \new_[2580]_  = ~\new_[2714]_  | ~\new_[2685]_ ;
  assign \new_[2581]_  = ~\new_[2715]_  | ~\new_[2716]_ ;
  assign \new_[2582]_  = ~\new_[13080]_  | ~\dma_req_o[3]  | ~\new_[2674]_  | ~\new_[9462]_ ;
  assign \new_[2583]_  = u4_u1_dma_req_in_hold2_reg;
  assign n1125 = ~\new_[2792]_  | ~\new_[2693]_  | ~\new_[2793]_ ;
  assign \new_[2585]_  = ~\new_[2500]_  & (~\new_[8633]_  | ~\new_[2794]_ );
  assign \new_[2586]_  = ~\new_[2501]_  & (~\new_[2794]_  | ~\new_[8970]_ );
  assign \new_[2587]_  = ~\new_[2502]_  & (~\new_[7866]_  | ~\new_[2794]_ );
  assign \new_[2588]_  = ~\new_[2504]_  & (~\new_[8247]_  | ~\new_[2794]_ );
  assign \new_[2589]_  = ~\new_[2718]_  | ~\new_[14610]_ ;
  assign \new_[2590]_  = \new_[2721]_  & \new_[2725]_ ;
  assign \new_[2591]_  = ~\new_[14611]_  & (~n1240 | ~\new_[9036]_ );
  assign \new_[2592]_  = ~\new_[14828]_  & (~n1250 | ~\new_[9036]_ );
  assign \new_[2593]_  = ~\new_[9558]_  & (~n1245 | ~\new_[9036]_ );
  assign \new_[2594]_  = ~\new_[9559]_  & (~n1255 | ~\new_[9036]_ );
  assign \new_[2595]_  = ~\new_[2726]_  | ~\new_[9036]_ ;
  assign \new_[2596]_  = ~\new_[2728]_  | ~\new_[9036]_ ;
  assign n1130 = ~\new_[2729]_  & ~\new_[9834]_ ;
  assign n1135 = ~\new_[2730]_  & ~\new_[9834]_ ;
  assign n1115 = ~\new_[2731]_  & ~\new_[9834]_ ;
  assign \new_[2600]_  = ~\new_[2476]_  | ~\new_[2852]_  | ~\new_[11106]_ ;
  assign \new_[2601]_  = ~\new_[2477]_  | ~\new_[2852]_  | ~\new_[11106]_ ;
  assign \new_[2602]_  = ~\new_[2478]_  | ~\new_[2852]_  | ~\new_[11106]_ ;
  assign \new_[2603]_  = ~\new_[2479]_  | ~\new_[2852]_  | ~\new_[11106]_ ;
  assign \new_[2604]_  = ~n8990 | ~\new_[2852]_  | ~\new_[11106]_ ;
  assign n1140 = ~\new_[2745]_  & ~\new_[7411]_ ;
  assign n1145 = ~\new_[2746]_  & ~\new_[8124]_ ;
  assign \new_[2607]_  = ~\new_[2887]_  | ~\new_[3047]_  | ~\new_[2888]_  | ~\new_[14452]_ ;
  assign n1150 = ~\new_[2747]_  & ~\new_[7414]_ ;
  assign n1155 = ~\new_[2748]_  & ~\new_[7418]_ ;
  assign \new_[2610]_  = ~\new_[2743]_  & (~\new_[3108]_  | ~\new_[12591]_ );
  assign \new_[2611]_  = u1_u3_abort_reg;
  assign \new_[2612]_  = ~\new_[5101]_  | ~\new_[5099]_  | ~\new_[14517]_  | ~\new_[4454]_ ;
  assign \new_[2613]_  = ~\\u1_u2_last_buf_adr_reg[8] ;
  assign \new_[2614]_  = ~\\u1_u2_last_buf_adr_reg[6] ;
  assign \new_[2615]_  = ~\new_[3011]_  | ~\new_[3447]_  | ~\new_[2894]_  | ~\new_[2827]_ ;
  assign \new_[2616]_  = \new_[2825]_  ^ \new_[8683]_ ;
  assign \new_[2617]_  = \new_[2826]_  ^ \new_[8851]_ ;
  assign n1120 = \new_[2755]_  ? n9145 : \new_[2869]_ ;
  assign \new_[2619]_  = \\u1_u2_dout_r_reg[30] ;
  assign \new_[2620]_  = u4_u2_dma_req_in_hold2_reg;
  assign \new_[2621]_  = u4_u0_dma_req_in_hold2_reg;
  assign \new_[2622]_  = \\u1_u2_dout_r_reg[5] ;
  assign \new_[2623]_  = \\u1_u2_dout_r_reg[27] ;
  assign \new_[2624]_  = \\u1_u2_dout_r_reg[1] ;
  assign \new_[2625]_  = \\u1_u2_dout_r_reg[16] ;
  assign n1180 = ~\new_[6963]_  & (~\new_[2839]_  | ~\new_[13757]_ );
  assign \new_[2627]_  = ~\new_[9457]_  & ~\new_[2795]_ ;
  assign \new_[2628]_  = ~\new_[9560]_  & (~n1445 | ~\new_[9036]_ );
  assign \new_[2629]_  = ~\new_[9312]_  & (~n1440 | ~\new_[9036]_ );
  assign \new_[2630]_  = \\u1_u3_size_next_r_reg[1] ;
  assign \new_[2631]_  = \\u1_u3_size_next_r_reg[3] ;
  assign \new_[2632]_  = \\u1_u3_size_next_r_reg[2] ;
  assign \new_[2633]_  = \\u1_u3_size_next_r_reg[5] ;
  assign \new_[2634]_  = ~\new_[8566]_  | ~\new_[2923]_ ;
  assign \new_[2635]_  = ~\new_[2923]_  & ~\new_[2373]_ ;
  assign \new_[2636]_  = \\u1_u2_adr_cb_reg[0] ;
  assign \new_[2637]_  = \\u1_mfm_cnt_reg[1] ;
  assign \new_[2638]_  = \\u1_u3_idin_reg[25] ;
  assign \new_[2639]_  = \\u1_u3_idin_reg[26] ;
  assign n1165 = ~\new_[2738]_ ;
  assign n1160 = ~\new_[2739]_ ;
  assign n1170 = ~\new_[2740]_ ;
  assign \new_[2643]_  = \\u1_u2_dout_r_reg[0] ;
  assign \new_[2644]_  = \\u1_u2_dout_r_reg[10] ;
  assign \new_[2645]_  = \\u1_u2_dout_r_reg[12] ;
  assign \new_[2646]_  = \\u1_u2_dout_r_reg[11] ;
  assign \new_[2647]_  = \\u1_u2_dout_r_reg[13] ;
  assign \new_[2648]_  = \\u1_u2_dout_r_reg[14] ;
  assign \new_[2649]_  = \\u1_u2_dout_r_reg[15] ;
  assign \new_[2650]_  = \\u1_u2_dout_r_reg[17] ;
  assign \new_[2651]_  = \\u1_u2_dout_r_reg[18] ;
  assign \new_[2652]_  = \\u1_u2_dout_r_reg[19] ;
  assign \new_[2653]_  = \\u1_u2_dout_r_reg[20] ;
  assign \new_[2654]_  = \\u1_u2_dout_r_reg[21] ;
  assign \new_[2655]_  = \\u1_u2_dout_r_reg[22] ;
  assign \new_[2656]_  = \\u1_u2_dout_r_reg[23] ;
  assign \new_[2657]_  = \\u1_u2_dout_r_reg[24] ;
  assign \new_[2658]_  = \\u1_u2_dout_r_reg[25] ;
  assign \new_[2659]_  = \\u1_u2_dout_r_reg[26] ;
  assign \new_[2660]_  = \\u1_u2_dout_r_reg[28] ;
  assign \new_[2661]_  = \\u1_u2_dout_r_reg[29] ;
  assign \new_[2662]_  = \\u1_u2_dout_r_reg[2] ;
  assign \new_[2663]_  = \\u1_u2_dout_r_reg[31] ;
  assign \new_[2664]_  = \\u1_u2_dout_r_reg[3] ;
  assign \new_[2665]_  = \\u1_u2_dout_r_reg[4] ;
  assign \new_[2666]_  = \\u1_u2_dout_r_reg[6] ;
  assign \new_[2667]_  = \\u1_u2_dout_r_reg[7] ;
  assign \new_[2668]_  = \\u1_u2_dout_r_reg[8] ;
  assign \new_[2669]_  = \\u1_u2_dout_r_reg[9] ;
  assign n1175 = ~\new_[2742]_ ;
  assign \new_[2671]_  = \new_[2892]_  ^ \new_[8679]_ ;
  assign \new_[2672]_  = ~\new_[2939]_  | ~\new_[4232]_  | ~\new_[2831]_ ;
  assign \new_[2673]_  = ~u0_u0_me_cnt_100_ms_reg;
  assign \new_[2674]_  = u4_u3_dma_req_in_hold2_reg;
  assign n1185 = ~\new_[2837]_  | ~\new_[2919]_ ;
  assign \new_[2676]_  = ~\new_[2841]_  | ~\new_[10552]_ ;
  assign \new_[2677]_  = ~\new_[14753]_  | ~\new_[11334]_ ;
  assign \new_[2678]_  = ~\new_[2841]_  | ~\new_[10640]_ ;
  assign \new_[2679]_  = ~\new_[2840]_  | ~\new_[11028]_ ;
  assign \new_[2680]_  = ~\new_[2841]_  | ~\new_[10669]_ ;
  assign \new_[2681]_  = ~\new_[2840]_  | ~\new_[11365]_ ;
  assign \new_[2682]_  = ~\new_[2840]_  | ~\new_[11327]_ ;
  assign \new_[2683]_  = ~\new_[2841]_  | ~\new_[10515]_ ;
  assign \new_[2684]_  = ~\new_[2840]_  | ~\new_[11018]_ ;
  assign \new_[2685]_  = ~\new_[2841]_  | ~\new_[10507]_ ;
  assign \new_[2686]_  = ~\new_[14824]_  | ~\new_[10656]_ ;
  assign \new_[2687]_  = ~\new_[2844]_  | ~\new_[11363]_ ;
  assign \new_[2688]_  = ~\new_[2845]_  | ~\new_[11352]_ ;
  assign \new_[2689]_  = ~\new_[2846]_  | ~\new_[10645]_ ;
  assign \new_[2690]_  = ~\new_[14721]_  | ~\new_[11216]_ ;
  assign \new_[2691]_  = ~\new_[14596]_  | ~\new_[10634]_ ;
  assign \new_[2692]_  = ~\new_[2847]_  | ~\new_[10694]_ ;
  assign \new_[2693]_  = ~\new_[2838]_  & (~\new_[7482]_  | ~\new_[2977]_ );
  assign \new_[2694]_  = ~\new_[14824]_  | ~\new_[10646]_ ;
  assign \new_[2695]_  = ~\new_[2845]_  | ~\new_[11391]_ ;
  assign \new_[2696]_  = ~\new_[2844]_  | ~\new_[11218]_ ;
  assign \new_[2697]_  = ~\new_[14596]_  | ~\new_[10664]_ ;
  assign \new_[2698]_  = ~\new_[14566]_  | ~\new_[10636]_ ;
  assign \new_[2699]_  = ~\new_[14721]_  | ~\new_[11381]_ ;
  assign \new_[2700]_  = ~\new_[14596]_  | ~\new_[10644]_ ;
  assign \new_[2701]_  = ~\new_[14566]_  | ~\new_[10695]_ ;
  assign \new_[2702]_  = ~\new_[14824]_  | ~\new_[10568]_ ;
  assign \new_[2703]_  = ~\new_[14721]_  | ~\new_[11380]_ ;
  assign \new_[2704]_  = \\u1_mfm_cnt_reg[3] ;
  assign \new_[2705]_  = ~\new_[14721]_  | ~\new_[11386]_ ;
  assign \new_[2706]_  = ~\new_[2844]_  | ~\new_[11030]_ ;
  assign \new_[2707]_  = ~\new_[2845]_  | ~\new_[11355]_ ;
  assign \new_[2708]_  = ~\new_[14596]_  | ~\new_[10643]_ ;
  assign \new_[2709]_  = ~\new_[14824]_  | ~\new_[10647]_ ;
  assign \new_[2710]_  = ~\new_[14566]_  | ~\new_[10641]_ ;
  assign \new_[2711]_  = ~\new_[14721]_  | ~\new_[11057]_ ;
  assign \new_[2712]_  = ~\new_[2844]_  | ~\new_[11384]_ ;
  assign \new_[2713]_  = ~\new_[2845]_  | ~\new_[11398]_ ;
  assign \new_[2714]_  = ~\new_[14824]_  | ~\new_[10649]_ ;
  assign \new_[2715]_  = ~\new_[14596]_  | ~\new_[10547]_ ;
  assign \new_[2716]_  = ~\new_[14566]_  | ~\new_[10648]_ ;
  assign \new_[2717]_  = \\u1_mfm_cnt_reg[0] ;
  assign \new_[2718]_  = \\u1_u3_size_next_r_reg[0] ;
  assign \new_[2719]_  = \\u1_u3_size_next_r_reg[4] ;
  assign \new_[2720]_  = \\u1_u3_size_next_r_reg[10] ;
  assign \new_[2721]_  = \new_[2852]_  | \new_[10479]_ ;
  assign \new_[2722]_  = ~\new_[2852]_  & ~\new_[9910]_ ;
  assign n1190 = ~\new_[2980]_  | ~\new_[2878]_ ;
  assign \new_[2724]_  = ~n1435 | ~\new_[9036]_ ;
  assign \new_[2725]_  = \new_[9140]_  | \new_[2852]_ ;
  assign \new_[2726]_  = \\u1_u3_size_next_r_reg[11] ;
  assign \new_[2727]_  = \\u1_u3_size_next_r_reg[12] ;
  assign \new_[2728]_  = \\u1_u3_size_next_r_reg[13] ;
  assign \new_[2729]_  = ~n1450 | ~\new_[9036]_ ;
  assign \new_[2730]_  = ~n1455 | ~\new_[9036]_ ;
  assign \new_[2731]_  = ~n1460 | ~\new_[9036]_ ;
  assign \new_[2732]_  = ~n1250;
  assign \new_[2733]_  = ~n1245;
  assign \new_[2734]_  = \\u1_u2_adr_cb_reg[2] ;
  assign \new_[2735]_  = \\u1_u3_idin_reg[29] ;
  assign \new_[2736]_  = ~n1255;
  assign \new_[2737]_  = \\u1_mfm_cnt_reg[2] ;
  assign \new_[2738]_  = ~\new_[2881]_  & (~\new_[3000]_  | ~\new_[4800]_ );
  assign \new_[2739]_  = ~\new_[2882]_  & (~\new_[3000]_  | ~\new_[4801]_ );
  assign \new_[2740]_  = ~\new_[2883]_  & (~\new_[3000]_  | ~\new_[4802]_ );
  assign \new_[2741]_  = u1_u2_word_done_r_reg;
  assign \new_[2742]_  = ~\new_[2884]_  & (~\new_[3000]_  | ~\new_[4651]_ );
  assign \new_[2743]_  = ~\new_[2888]_  & ~\new_[4802]_ ;
  assign \new_[2744]_  = ~\new_[2890]_  | ~\new_[2999]_ ;
  assign \new_[2745]_  = ~\new_[2551]_  & (~\new_[8633]_  | ~\new_[2936]_ );
  assign \new_[2746]_  = ~\new_[2552]_  & (~\new_[2936]_  | ~\new_[8970]_ );
  assign \new_[2747]_  = ~\new_[2553]_  & (~\new_[7866]_  | ~\new_[2936]_ );
  assign \new_[2748]_  = ~\new_[2554]_  & (~\new_[8247]_  | ~\new_[2936]_ );
  assign \new_[2749]_  = ~\new_[3245]_  | ~\new_[3003]_  | ~\new_[3395]_  | ~\new_[3267]_ ;
  assign n1200 = \new_[4034]_  ^ \new_[14495]_ ;
  assign n1195 = \new_[4268]_  ^ \new_[2938]_ ;
  assign \new_[2752]_  = ~\new_[3134]_  | ~\new_[4231]_  | ~\new_[2899]_ ;
  assign \new_[2753]_  = ~\new_[2829]_  & ~\new_[4923]_ ;
  assign \new_[2754]_  = ~\new_[2829]_  | ~\new_[4923]_ ;
  assign \new_[2755]_  = ~\new_[2829]_ ;
  assign n1280 = \new_[2862]_  ? \new_[2960]_  : \new_[2643]_ ;
  assign n1285 = \new_[2804]_  ? \new_[2960]_  : \new_[2644]_ ;
  assign n1295 = \new_[2805]_  ? \new_[2960]_  : \new_[2646]_ ;
  assign n1290 = \new_[2788]_  ? \new_[2960]_  : \new_[2645]_ ;
  assign n1300 = \new_[2806]_  ? \new_[2960]_  : \new_[2647]_ ;
  assign n1305 = \new_[2807]_  ? \new_[2960]_  : \new_[2648]_ ;
  assign n1310 = \new_[2808]_  ? \new_[2960]_  : \new_[2649]_ ;
  assign n1235 = \new_[2833]_  ? \new_[2960]_  : \new_[2625]_ ;
  assign n1315 = \new_[2809]_  ? \new_[2960]_  : \new_[2650]_ ;
  assign n1320 = \new_[2858]_  ? \new_[2960]_  : \new_[2651]_ ;
  assign n1325 = \new_[2830]_  ? \new_[2960]_  : \new_[2652]_ ;
  assign n1230 = \new_[2863]_  ? \new_[2960]_  : \new_[2624]_ ;
  assign n1330 = \new_[2859]_  ? \new_[2960]_  : \new_[2653]_ ;
  assign n1335 = \new_[2860]_  ? \new_[2960]_  : \new_[2654]_ ;
  assign n1340 = \new_[2893]_  ? \new_[2960]_  : \new_[2655]_ ;
  assign n1345 = \new_[2810]_  ? \new_[2960]_  : \new_[2656]_ ;
  assign n1350 = \new_[2812]_  ? \new_[2960]_  : \new_[2657]_ ;
  assign n1355 = \new_[2811]_  ? \new_[2960]_  : \new_[2658]_ ;
  assign n1360 = \new_[2813]_  ? \new_[2960]_  : \new_[2659]_ ;
  assign n1225 = \new_[2814]_  ? \new_[2960]_  : \new_[2623]_ ;
  assign n1365 = \new_[2828]_  ? \new_[2960]_  : \new_[2660]_ ;
  assign n1370 = \new_[2815]_  ? \new_[2960]_  : \new_[2661]_ ;
  assign n1375 = \new_[2895]_  ? \new_[2960]_  : \new_[2662]_ ;
  assign n1205 = \new_[2816]_  ? \new_[2960]_  : \new_[2619]_ ;
  assign n1380 = \new_[2817]_  ? \new_[2960]_  : \new_[2663]_ ;
  assign n1385 = \new_[2868]_  ? \new_[2960]_  : \new_[2664]_ ;
  assign n1390 = \new_[2864]_  ? \new_[2960]_  : \new_[2665]_ ;
  assign n1220 = \new_[2865]_  ? \new_[2960]_  : \new_[2622]_ ;
  assign n1395 = \new_[2866]_  ? \new_[2960]_  : \new_[2666]_ ;
  assign n1400 = \new_[2867]_  ? \new_[2960]_  : \new_[2667]_ ;
  assign n1405 = \new_[2896]_  ? \new_[2960]_  : \new_[2668]_ ;
  assign n1410 = \new_[2861]_  ? \new_[2960]_  : \new_[2669]_ ;
  assign \new_[2788]_  = \\u1_u2_dtmp_r_reg[12] ;
  assign n1210 = ~\new_[2917]_  | ~\new_[2971]_ ;
  assign n1215 = ~\new_[2918]_  | ~\new_[2974]_ ;
  assign n1260 = ~\new_[2931]_  & ~\new_[12804]_ ;
  assign \new_[2792]_  = (~\new_[7483]_  | ~\new_[2548]_ ) & (~n7650 | ~\new_[2975]_ );
  assign \new_[2793]_  = ~\new_[8634]_  | ~\new_[2920]_ ;
  assign \new_[2794]_  = u1_u3_int_upid_set_reg;
  assign \new_[2795]_  = ~\new_[9140]_  | ~\new_[2923]_ ;
  assign n1265 = ~\new_[2994]_  & (~\new_[2998]_  | ~\new_[3046]_ );
  assign \new_[2797]_  = ~n1445;
  assign \new_[2798]_  = ~n1435;
  assign n1245 = \new_[7298]_  ? \new_[14781]_  : \new_[4798]_ ;
  assign \new_[2800]_  = ~n1440;
  assign \new_[2801]_  = \\u1_u2_adr_cb_reg[1] ;
  assign \new_[2802]_  = ~\\u1_u3_new_size_reg[11] ;
  assign n1255 = \new_[7846]_  ? \new_[14781]_  : \new_[4620]_ ;
  assign \new_[2804]_  = \\u1_u2_dtmp_r_reg[10] ;
  assign \new_[2805]_  = \\u1_u2_dtmp_r_reg[11] ;
  assign \new_[2806]_  = \\u1_u2_dtmp_r_reg[13] ;
  assign \new_[2807]_  = \\u1_u2_dtmp_r_reg[14] ;
  assign \new_[2808]_  = \\u1_u2_dtmp_r_reg[15] ;
  assign \new_[2809]_  = \\u1_u2_dtmp_r_reg[17] ;
  assign \new_[2810]_  = \\u1_u2_dtmp_r_reg[23] ;
  assign \new_[2811]_  = \\u1_u2_dtmp_r_reg[25] ;
  assign \new_[2812]_  = \\u1_u2_dtmp_r_reg[24] ;
  assign \new_[2813]_  = \\u1_u2_dtmp_r_reg[26] ;
  assign \new_[2814]_  = \\u1_u2_dtmp_r_reg[27] ;
  assign \new_[2815]_  = \\u1_u2_dtmp_r_reg[29] ;
  assign \new_[2816]_  = \\u1_u2_dtmp_r_reg[30] ;
  assign \new_[2817]_  = \\u1_u2_dtmp_r_reg[31] ;
  assign \new_[2818]_  = ~n1450;
  assign \new_[2819]_  = ~n1455;
  assign \new_[2820]_  = ~n1460;
  assign \new_[2821]_  = ~\new_[2935]_  & (~\new_[3414]_  | ~\new_[13118]_ );
  assign n1270 = \new_[3108]_  ? n9145 : \new_[2857]_ ;
  assign n1275 = ~\new_[13312]_  | (~\new_[3003]_  & ~n9145);
  assign \new_[2824]_  = ~\new_[3059]_  | ~\new_[3124]_  | ~\new_[3061]_  | ~\new_[14582]_ ;
  assign \new_[2825]_  = ~\\u1_u2_last_buf_adr_reg[4] ;
  assign \new_[2826]_  = ~\\u1_u2_last_buf_adr_reg[5] ;
  assign \new_[2827]_  = \new_[2942]_  ^ \new_[8852]_ ;
  assign \new_[2828]_  = \\u1_u2_dtmp_r_reg[28] ;
  assign \new_[2829]_  = ~\\u1_u3_new_size_reg[10] ;
  assign \new_[2830]_  = \\u1_u2_dtmp_r_reg[19] ;
  assign \new_[2831]_  = ~\new_[2973]_  | ~\new_[4453]_ ;
  assign n1480 = ~\new_[2960]_  & ~\new_[2741]_ ;
  assign \new_[2833]_  = \\u1_u2_dtmp_r_reg[16] ;
  assign n1420 = ~\new_[2963]_  | ~\new_[3015]_ ;
  assign n1465 = ~\new_[2978]_  & ~\new_[12804]_ ;
  assign \new_[2836]_  = \\u1_u2_sizu_c_reg[5] ;
  assign \new_[2837]_  = ~\new_[6674]_  | ~\new_[7180]_  | ~\new_[8275]_  | ~\new_[3017]_ ;
  assign \new_[2838]_  = ~\new_[8622]_  & ~\new_[2976]_ ;
  assign \new_[2839]_  = ~u4_nse_err_r_reg;
  assign \new_[2840]_  = ~\new_[14755]_ ;
  assign \new_[2841]_  = ~\new_[2921]_ ;
  assign \new_[2842]_  = ~\new_[2921]_ ;
  assign \new_[2843]_  = ~\new_[2921]_ ;
  assign \new_[2844]_  = ~\new_[14639]_ ;
  assign \new_[2845]_  = ~\new_[14675]_ ;
  assign \new_[2846]_  = ~\new_[14567]_ ;
  assign \new_[2847]_  = ~\new_[14567]_ ;
  assign \new_[2848]_  = ~\new_[2981]_  & (~\new_[10402]_  | ~\new_[5154]_ );
  assign n1430 = ~\new_[3045]_  & ~\new_[2994]_ ;
  assign n1475 = ~\new_[2995]_  & ~\new_[2994]_ ;
  assign n1425 = ~\new_[2996]_  & ~\new_[2994]_ ;
  assign \new_[2852]_  = ~\new_[2923]_ ;
  assign n1435 = \new_[14548]_  ? \new_[3048]_  : \new_[4852]_ ;
  assign n1445 = \new_[14507]_  ? \new_[3048]_  : \new_[4923]_ ;
  assign n1440 = \new_[8602]_  ? \new_[3048]_  : \new_[12760]_ ;
  assign \new_[2856]_  = \\u1_u3_idin_reg[24] ;
  assign \new_[2857]_  = \\u1_u2_sizu_c_reg[8] ;
  assign \new_[2858]_  = \\u1_u2_dtmp_r_reg[18] ;
  assign \new_[2859]_  = \\u1_u2_dtmp_r_reg[20] ;
  assign \new_[2860]_  = \\u1_u2_dtmp_r_reg[21] ;
  assign \new_[2861]_  = \\u1_u2_dtmp_r_reg[9] ;
  assign \new_[2862]_  = \\u1_u2_dtmp_r_reg[0] ;
  assign \new_[2863]_  = \\u1_u2_dtmp_r_reg[1] ;
  assign \new_[2864]_  = \\u1_u2_dtmp_r_reg[4] ;
  assign \new_[2865]_  = \\u1_u2_dtmp_r_reg[5] ;
  assign \new_[2866]_  = \\u1_u2_dtmp_r_reg[6] ;
  assign \new_[2867]_  = \\u1_u2_dtmp_r_reg[7] ;
  assign \new_[2868]_  = \\u1_u2_dtmp_r_reg[3] ;
  assign \new_[2869]_  = \\u1_u2_sizu_c_reg[10] ;
  assign \new_[2870]_  = \\u1_u2_sizu_c_reg[1] ;
  assign \new_[2871]_  = \\u1_u2_sizu_c_reg[2] ;
  assign \new_[2872]_  = \\u1_u2_sizu_c_reg[3] ;
  assign \new_[2873]_  = \\u1_u2_sizu_c_reg[4] ;
  assign \new_[2874]_  = \\u1_u2_sizu_c_reg[6] ;
  assign \new_[2875]_  = \\u1_u2_sizu_c_reg[7] ;
  assign \new_[2876]_  = \\u1_u2_sizu_c_reg[9] ;
  assign n1450 = ~\new_[3000]_  & ~\new_[14270]_ ;
  assign \new_[2878]_  = ~u1_u3_buffer_overflow_reg;
  assign n1455 = ~\new_[14276]_  & ~\new_[3000]_ ;
  assign n1460 = ~\new_[3000]_  & ~\new_[14312]_ ;
  assign \new_[2881]_  = ~\new_[3001]_  & ~\new_[8224]_ ;
  assign \new_[2882]_  = ~\new_[3001]_  & ~\new_[8601]_ ;
  assign \new_[2883]_  = ~\new_[3000]_  & ~\new_[8603]_ ;
  assign \new_[2884]_  = ~\new_[3001]_  & ~\new_[8600]_ ;
  assign n1415 = ~\new_[2934]_ ;
  assign \new_[2886]_  = \new_[3003]_  | \new_[4651]_ ;
  assign \new_[2887]_  = \new_[3003]_  | \new_[4802]_ ;
  assign \new_[2888]_  = \new_[3245]_  | \new_[3003]_ ;
  assign \new_[2889]_  = (~\new_[3061]_  & ~\new_[4800]_ ) | (~\new_[3395]_  & ~\new_[14582]_ );
  assign \new_[2890]_  = ~\new_[3008]_  | (~\new_[3632]_  & ~\new_[4798]_ );
  assign n1470 = ~\new_[3005]_  & ~n9145;
  assign \new_[2892]_  = ~\\u1_u2_last_buf_adr_reg[7] ;
  assign \new_[2893]_  = \\u1_u2_dtmp_r_reg[22] ;
  assign \new_[2894]_  = \new_[3009]_  ^ \new_[8668]_ ;
  assign \new_[2895]_  = \\u1_u2_dtmp_r_reg[2] ;
  assign \new_[2896]_  = \\u1_u2_dtmp_r_reg[8] ;
  assign n1575 = \new_[4033]_  ^ \new_[14471]_ ;
  assign n1580 = \new_[4266]_  ^ \new_[14521]_ ;
  assign \new_[2899]_  = ~\new_[3016]_  | ~\new_[4454]_ ;
  assign n1505 = ~\new_[9335]_  | (~\new_[3085]_  & ~\new_[9914]_ );
  assign n1510 = ~\new_[9315]_  | (~\new_[3086]_  & ~\new_[9914]_ );
  assign n1485 = ~\new_[9319]_  | (~\new_[3087]_  & ~\new_[9914]_ );
  assign n1515 = ~\new_[9320]_  | (~\new_[3088]_  & ~\new_[9914]_ );
  assign n1520 = ~\new_[9339]_  | (~\new_[3089]_  & ~\new_[9914]_ );
  assign n1525 = ~\new_[9340]_  | (~\new_[3090]_  & ~\new_[9914]_ );
  assign n1530 = ~\new_[9323]_  | (~\new_[3091]_  & ~\new_[9914]_ );
  assign n1535 = ~\new_[9330]_  | (~\new_[3092]_  & ~\new_[9914]_ );
  assign n1545 = ~\new_[9341]_  | (~\new_[3093]_  & ~\new_[9914]_ );
  assign n1540 = ~\new_[9342]_  | (~\new_[3094]_  & ~\new_[9914]_ );
  assign n1550 = ~\new_[9344]_  | (~\new_[3095]_  & ~\new_[9914]_ );
  assign n1555 = ~\new_[9331]_  | (~\new_[3096]_  & ~\new_[9914]_ );
  assign n1585 = ~\new_[9322]_  | (~\new_[3097]_  & ~\new_[9914]_ );
  assign n1560 = ~\new_[9345]_  | (~\new_[3098]_  & ~\new_[9914]_ );
  assign n1565 = ~\new_[9317]_  | (~\new_[3099]_  & ~\new_[9914]_ );
  assign n1570 = ~\new_[9329]_  | (~\new_[3100]_  & ~\new_[9914]_ );
  assign n1495 = ~\new_[3020]_  & ~\new_[12804]_ ;
  assign \new_[2917]_  = ~\new_[7390]_  | ~\new_[7734]_  | ~\new_[9026]_  | ~\new_[3070]_ ;
  assign \new_[2918]_  = ~\new_[7071]_  | ~\new_[7437]_  | ~\new_[8656]_  | ~\new_[3071]_ ;
  assign \new_[2919]_  = ~\new_[5543]_  | ~\new_[3017]_ ;
  assign \new_[2920]_  = u4_u1_dma_out_buf_avail_reg;
  assign \new_[2921]_  = ~\new_[3120]_  | ~\new_[14820]_ ;
  assign n1490 = ~\new_[3042]_  & (~\new_[8968]_  | ~\new_[9194]_ );
  assign \new_[2923]_  = ~\new_[3042]_  & (~\new_[4790]_  | ~\new_[13692]_ );
  assign \new_[2924]_  = \\u1_frame_no_r_reg[10] ;
  assign \new_[2925]_  = \\u1_frame_no_r_reg[4] ;
  assign \new_[2926]_  = \\u1_frame_no_r_reg[7] ;
  assign \new_[2927]_  = \\u1_frame_no_r_reg[8] ;
  assign \new_[2928]_  = \\u1_u3_idin_reg[23] ;
  assign \new_[2929]_  = \\u1_frame_no_r_reg[9] ;
  assign wb_ack_o = u5_wb_ack_o_reg;
  assign \new_[2931]_  = ~\new_[4747]_  & (~\new_[14657]_  | ~\new_[13330]_ );
  assign \new_[2932]_  = \\u1_u2_sizu_c_reg[0] ;
  assign \new_[2933]_  = u1_u2_wr_last_reg;
  assign \new_[2934]_  = ~\new_[13608]_  | ~\new_[3050]_  | ~\new_[13694]_ ;
  assign \new_[2935]_  = ~\new_[2999]_ ;
  assign \new_[2936]_  = u1_u3_int_seqerr_set_reg;
  assign n1500 = \new_[6707]_  ^ \new_[3065]_ ;
  assign \new_[2938]_  = ~\new_[3388]_  & (~\new_[14471]_  | ~\new_[3803]_ );
  assign \new_[2939]_  = ~\new_[14489]_  | ~\new_[3803]_  | ~\new_[14471]_  | ~\new_[4453]_ ;
  assign n1725 = \new_[4267]_  ^ \new_[3133]_ ;
  assign n1590 = ~\new_[3067]_  | (~\new_[3615]_  & ~\new_[3413]_ );
  assign \new_[2942]_  = ~\\u1_u2_last_buf_adr_reg[2] ;
  assign n1680 = ~\new_[3068]_  & ~\new_[12681]_ ;
  assign n1600 = ~\new_[9348]_  | (~\new_[3139]_  & ~\new_[9914]_ );
  assign n1625 = ~\new_[9334]_  | (~\new_[3140]_  & ~\new_[9914]_ );
  assign n1595 = ~\new_[9347]_  | (~\new_[3141]_  & ~\new_[9914]_ );
  assign n1630 = ~\new_[9326]_  | (~\new_[3142]_  & ~\new_[9914]_ );
  assign n1635 = ~\new_[9321]_  | (~\new_[3143]_  & ~\new_[9914]_ );
  assign n1730 = ~\new_[9316]_  | (~\new_[3144]_  & ~\new_[9914]_ );
  assign n1740 = ~\new_[9343]_  | (~\new_[3145]_  & ~\new_[9914]_ );
  assign n1640 = ~\new_[9346]_  | (~\new_[3146]_  & ~\new_[9914]_ );
  assign n1645 = \new_[3147]_  ? \new_[9914]_  : \sram_data_i[0] ;
  assign n1650 = \new_[3148]_  ? \new_[9914]_  : \sram_data_i[1] ;
  assign n1735 = \new_[3149]_  ? \new_[9914]_  : \sram_data_i[2] ;
  assign n1675 = \new_[3150]_  ? \new_[9914]_  : \sram_data_i[3] ;
  assign n1655 = \new_[3151]_  ? \new_[9914]_  : \sram_data_i[4] ;
  assign n1660 = \new_[3152]_  ? \new_[9914]_  : \sram_data_i[5] ;
  assign n1665 = \new_[3153]_  ? \new_[9914]_  : \sram_data_i[6] ;
  assign n1670 = \new_[3154]_  ? \new_[9914]_  : \sram_data_i[7] ;
  assign \new_[2960]_  = ~u1_u2_word_done_reg;
  assign \new_[2961]_  = u0_u0_T2_wakeup_reg;
  assign \new_[2962]_  = \\u1_frame_no_r_reg[5] ;
  assign \new_[2963]_  = ~\new_[7391]_  | ~\new_[7737]_  | ~\new_[9027]_  | ~\new_[3136]_ ;
  assign n1690 = ~\new_[3081]_  & ~\new_[12681]_ ;
  assign n1695 = ~\new_[3082]_  & ~\new_[12681]_ ;
  assign n1700 = ~\new_[3083]_  & ~\new_[12681]_ ;
  assign n1605 = ~\new_[3084]_  & ~\new_[12681]_ ;
  assign n1705 = ~\new_[3078]_  & ~\new_[12681]_ ;
  assign n1710 = ~\new_[3079]_  & ~\new_[12681]_ ;
  assign n1715 = ~\new_[3080]_  & ~\new_[12681]_ ;
  assign \new_[2971]_  = ~\new_[4876]_  | ~\new_[3070]_ ;
  assign n1685 = ~\new_[12681]_  & (~\new_[3359]_  | ~\new_[3193]_ );
  assign \new_[2973]_  = ~\new_[3072]_  | ~\new_[14491]_ ;
  assign \new_[2974]_  = ~\new_[4877]_  | ~\new_[3071]_ ;
  assign \new_[2975]_  = u4_u0_dma_out_buf_avail_reg;
  assign \new_[2976]_  = ~u4_u2_dma_out_buf_avail_reg;
  assign \new_[2977]_  = u4_u3_dma_out_buf_avail_reg;
  assign \new_[2978]_  = ~\new_[4748]_  & (~\new_[3248]_  | ~\new_[13330]_ );
  assign n1610 = u1_u3_nse_err_reg;
  assign \new_[2980]_  = (~n2260 | ~\new_[10382]_ ) & (~\new_[3242]_  | ~\new_[4413]_ );
  assign \new_[2981]_  = ~\new_[9803]_  | (~\new_[10726]_  & ~\new_[3243]_ );
  assign \new_[2982]_  = \\u1_hms_cnt_reg[1] ;
  assign \new_[2983]_  = \\u1_frame_no_r_reg[0] ;
  assign \new_[2984]_  = \\u1_frame_no_r_reg[3] ;
  assign \new_[2985]_  = \\u1_frame_no_r_reg[1] ;
  assign \new_[2986]_  = \\u1_frame_no_r_reg[2] ;
  assign \new_[2987]_  = \\u1_frame_no_r_reg[6] ;
  assign \new_[2988]_  = \\u1_hms_cnt_reg[2] ;
  assign \new_[2989]_  = \\u1_hms_cnt_reg[3] ;
  assign \new_[2990]_  = u0_u0_T2_gt_100_uS_reg;
  assign \new_[2991]_  = u0_u0_T2_gt_1_0_mS_reg;
  assign \new_[2992]_  = u0_u0_T2_gt_1_2_mS_reg;
  assign \new_[2993]_  = ~\\u0_u0_me_ps_reg[1] ;
  assign \new_[2994]_  = ~phy_rst_pad_o | (~\new_[4191]_  & ~\new_[3244]_ );
  assign \new_[2995]_  = (~\new_[11449]_  | ~\new_[3244]_ ) & (~\new_[3387]_  | ~\new_[2737]_ );
  assign \new_[2996]_  = (~\new_[10978]_  | ~\new_[3244]_ ) & (~\new_[3387]_  | ~\new_[2704]_ );
  assign n1720 = ~\new_[3113]_  | (~\new_[3571]_  & ~\new_[4554]_ );
  assign \new_[2998]_  = ~\new_[3387]_  | ~\new_[2637]_ ;
  assign \new_[2999]_  = ~\new_[11715]_  | ~\new_[3392]_  | ~\new_[3394]_  | ~\new_[14424]_ ;
  assign \new_[3000]_  = ~\new_[3049]_ ;
  assign \new_[3001]_  = ~\new_[14782]_ ;
  assign \new_[3002]_  = ~\new_[3112]_  & (~\new_[3782]_  | ~\new_[12565]_ );
  assign \new_[3003]_  = ~\\u1_u3_new_size_reg[9] ;
  assign n1615 = ~\new_[13410]_  | (~\new_[3267]_  & ~n9145);
  assign \new_[3005]_  = ~\\u1_u3_new_size_reg[12] ;
  assign n1620 = ~\new_[3064]_  & ~\new_[12681]_ ;
  assign \new_[3007]_  = ~\new_[3278]_  | ~\new_[3598]_  | ~\new_[3279]_  | ~\new_[12932]_ ;
  assign \new_[3008]_  = ~\new_[3599]_  & ~\new_[3129]_ ;
  assign \new_[3009]_  = ~\\u1_u2_last_buf_adr_reg[3] ;
  assign \new_[3010]_  = ~\\u0_u0_me_ps2_reg[5] ;
  assign \new_[3011]_  = \new_[3286]_  ^ \new_[8969]_ ;
  assign \new_[3012]_  = ~\\u0_u0_me_cnt_reg[4] ;
  assign \new_[3013]_  = \\u1_hms_cnt_reg[4] ;
  assign n1785 = ~\new_[3155]_  & ~\new_[12681]_ ;
  assign \new_[3015]_  = ~\new_[5542]_  | ~\new_[3136]_ ;
  assign \new_[3016]_  = ~\new_[3137]_  | ~\new_[14523]_ ;
  assign \new_[3017]_  = ~\new_[3138]_  | (~\new_[5581]_  & ~\new_[4062]_ );
  assign n1790 = ~\new_[3194]_  & ~\new_[5224]_ ;
  assign n1745 = ~\new_[3531]_  | ~\new_[6781]_  | ~\new_[4938]_  | ~\new_[4942]_ ;
  assign \new_[3020]_  = \new_[5511]_  ? \new_[13330]_  : \new_[14774]_ ;
  assign \new_[3021]_  = \\u1_u3_idin_reg[21] ;
  assign \new_[3022]_  = ~\\u0_u0_me_ps2_reg[0] ;
  assign \new_[3023]_  = ~\\u0_u0_me_ps2_reg[1] ;
  assign \new_[3024]_  = ~\\u0_u0_me_ps2_reg[2] ;
  assign \new_[3025]_  = \\u0_u0_me_ps2_reg[3] ;
  assign \new_[3026]_  = ~\\u0_u0_me_ps2_reg[4] ;
  assign \new_[3027]_  = ~\\u0_u0_me_ps2_reg[6] ;
  assign \new_[3028]_  = ~\\u0_u0_me_ps2_reg[7] ;
  assign \new_[3029]_  = ~\\u0_u0_me_ps_reg[0] ;
  assign \new_[3030]_  = ~\\u0_u0_me_ps_reg[2] ;
  assign \new_[3031]_  = ~\\u0_u0_me_ps_reg[4] ;
  assign \new_[3032]_  = ~\\u0_u0_me_ps_reg[5] ;
  assign \new_[3033]_  = ~\\u0_u0_me_ps_reg[6] ;
  assign \new_[3034]_  = \\u1_u3_idin_reg[20] ;
  assign \new_[3035]_  = \\u0_u0_me_cnt_reg[0] ;
  assign \new_[3036]_  = \\u0_u0_me_cnt_reg[1] ;
  assign \new_[3037]_  = \\u0_u0_me_cnt_reg[2] ;
  assign \new_[3038]_  = \\u0_u0_me_cnt_reg[3] ;
  assign \new_[3039]_  = ~\\u0_u0_me_cnt_reg[6] ;
  assign \new_[3040]_  = ~\\u0_u0_me_cnt_reg[7] ;
  assign \new_[3041]_  = ~\\u0_u0_me_cnt_reg[5] ;
  assign \new_[3042]_  = ~\new_[11725]_  | ~\new_[3242]_ ;
  assign sram_we_o = ~\new_[3253]_  | (~\new_[3400]_  & ~\new_[7654]_ );
  assign \new_[3044]_  = ~\new_[3107]_ ;
  assign \new_[3045]_  = \new_[2717]_  ^ \new_[3387]_ ;
  assign \new_[3046]_  = ~\new_[12889]_  | ~\new_[3244]_ ;
  assign \new_[3047]_  = \new_[3245]_  | \new_[4651]_ ;
  assign \new_[3048]_  = \new_[14791]_ ;
  assign \new_[3049]_  = ~\new_[14791]_ ;
  assign \new_[3050]_  = ~\new_[3265]_  & ~\new_[3036]_ ;
  assign n1750 = ~\new_[12245]_  & (~\new_[3402]_  | ~\new_[3576]_ );
  assign n1755 = ~\new_[12732]_  & (~\new_[3403]_  | ~\new_[3583]_ );
  assign n1760 = ~\new_[12849]_  & (~\new_[3404]_  | ~\new_[3588]_ );
  assign n1765 = ~\new_[12505]_  & (~\new_[3405]_  | ~\new_[3589]_ );
  assign n1775 = ~\new_[12505]_  & (~\new_[3406]_  | ~\new_[3590]_ );
  assign n1770 = ~\new_[13362]_  | (~\new_[3395]_  & ~n9145);
  assign n1780 = \new_[3276]_  & \new_[3266]_ ;
  assign \new_[3058]_  = ~\new_[3267]_  & ~\new_[4801]_ ;
  assign \new_[3059]_  = \new_[3267]_  | \new_[4800]_ ;
  assign n1795 = ~\new_[3126]_ ;
  assign \new_[3061]_  = \new_[3395]_  | \new_[3267]_ ;
  assign \new_[3062]_  = ~\\u0_u0_me_ps_reg[3] ;
  assign \new_[3063]_  = ~\\u0_u0_me_ps_reg[7] ;
  assign \new_[3064]_  = ~\new_[3277]_  & (~\new_[4154]_  | ~\new_[2857]_ );
  assign \new_[3065]_  = ~\new_[4201]_  | ~\new_[5623]_  | ~\new_[3420]_ ;
  assign \new_[3066]_  = ~\new_[4373]_  | (~\new_[4969]_  & ~\new_[14613]_ );
  assign \new_[3067]_  = ~\new_[3616]_  & (~\new_[3413]_  | ~\new_[5632]_ );
  assign \new_[3068]_  = ~\new_[3291]_  & (~\new_[4154]_  | ~\new_[2869]_ );
  assign n1800 = \new_[4264]_  ^ \new_[3553]_ ;
  assign \new_[3070]_  = ~\new_[3289]_  | (~\new_[5564]_  & ~\new_[4282]_ );
  assign \new_[3071]_  = ~\new_[3290]_  | (~\new_[5576]_  & ~\new_[4283]_ );
  assign \new_[3072]_  = ~\new_[3388]_  | ~\new_[14489]_ ;
  assign n1805 = \new_[3367]_  | \new_[2933]_ ;
  assign n1830 = ~\new_[3742]_  | ~\new_[7203]_  | ~\new_[4935]_  | ~\new_[4940]_ ;
  assign n1820 = ~\new_[3743]_  | ~\new_[6780]_  | ~\new_[4937]_  | ~\new_[4941]_ ;
  assign n1825 = ~\new_[3744]_  | ~\new_[7204]_  | ~\new_[4939]_  | ~\new_[4943]_ ;
  assign \new_[3077]_  = ~\new_[3389]_  | ~\new_[5101]_ ;
  assign \new_[3078]_  = ~\new_[3364]_  & (~\new_[4154]_  | ~\new_[2874]_ );
  assign \new_[3079]_  = ~\new_[3365]_  & (~\new_[4154]_  | ~\new_[2875]_ );
  assign \new_[3080]_  = ~\new_[3366]_  & (~\new_[4154]_  | ~\new_[2876]_ );
  assign \new_[3081]_  = ~\new_[3360]_  & (~\new_[4154]_  | ~\new_[2871]_ );
  assign \new_[3082]_  = ~\new_[3361]_  & (~\new_[4154]_  | ~\new_[2872]_ );
  assign \new_[3083]_  = ~\new_[3362]_  & (~\new_[4154]_  | ~\new_[2873]_ );
  assign \new_[3084]_  = ~\new_[3363]_  & (~\new_[4154]_  | ~\new_[2836]_ );
  assign \new_[3085]_  = ~\new_[3370]_  & (~\new_[2804]_  | ~\new_[4153]_ );
  assign \new_[3086]_  = ~\new_[3371]_  & (~\new_[2805]_  | ~\new_[4154]_ );
  assign \new_[3087]_  = ~\new_[3372]_  & (~\new_[2788]_  | ~\new_[4154]_ );
  assign \new_[3088]_  = ~\new_[3373]_  & (~\new_[2806]_  | ~\new_[4153]_ );
  assign \new_[3089]_  = ~\new_[3374]_  & (~\new_[2807]_  | ~\new_[4153]_ );
  assign \new_[3090]_  = ~\new_[3375]_  & (~\new_[2808]_  | ~\new_[4153]_ );
  assign \new_[3091]_  = ~\new_[3376]_  & (~\new_[2809]_  | ~\new_[4153]_ );
  assign \new_[3092]_  = ~\new_[3378]_  & (~\new_[2810]_  | ~\new_[4153]_ );
  assign \new_[3093]_  = ~\new_[3379]_  & (~\new_[2812]_  | ~\new_[4154]_ );
  assign \new_[3094]_  = ~\new_[3380]_  & (~\new_[2811]_  | ~\new_[4153]_ );
  assign \new_[3095]_  = ~\new_[3381]_  & (~\new_[2813]_  | ~\new_[4153]_ );
  assign \new_[3096]_  = ~\new_[3382]_  & (~\new_[2814]_  | ~\new_[4154]_ );
  assign \new_[3097]_  = ~\new_[3383]_  & (~\new_[2828]_  | ~\new_[4153]_ );
  assign \new_[3098]_  = ~\new_[3384]_  & (~\new_[2815]_  | ~\new_[4153]_ );
  assign \new_[3099]_  = ~\new_[3385]_  & (~\new_[2816]_  | ~\new_[4153]_ );
  assign \new_[3100]_  = ~\new_[3386]_  & (~\new_[2817]_  | ~\new_[4154]_ );
  assign \new_[3101]_  = \\u1_u2_state_reg[0] ;
  assign \new_[3102]_  = \\u1_u3_idin_reg[18] ;
  assign \new_[3103]_  = ~\\u4_u0_buf0_reg[28] ;
  assign \new_[3104]_  = ~\\u4_u0_buf0_reg[31] ;
  assign \new_[3105]_  = ~\new_[14411]_  & (~\new_[12456]_  | ~\new_[11816]_ );
  assign n1835 = ~\new_[3377]_  & (~\new_[10596]_  | ~\new_[11626]_ );
  assign \new_[3107]_  = ~\new_[14774]_  | ~\new_[14730]_ ;
  assign \new_[3108]_  = ~\new_[3245]_ ;
  assign n1840 = \new_[12891]_  & \new_[3391]_ ;
  assign n1870 = \new_[11720]_  & \new_[3391]_ ;
  assign n1875 = \new_[10975]_  & \new_[3391]_ ;
  assign \new_[3112]_  = ~\new_[3394]_  & ~\new_[12760]_ ;
  assign \new_[3113]_  = ~\new_[7186]_  | ~\new_[4586]_  | ~\new_[3398]_  | ~\new_[4517]_ ;
  assign n1845 = ~\new_[12505]_  & (~\new_[3574]_  | ~\new_[3575]_ );
  assign n1855 = ~\new_[12505]_  & (~\new_[3578]_  | ~\new_[3577]_ );
  assign n1850 = ~\new_[12505]_  & (~\new_[3582]_  | ~\new_[3581]_ );
  assign n1860 = ~\new_[12849]_  & (~\new_[3579]_  | ~\new_[3580]_ );
  assign n1815 = ~\new_[12505]_  & (~\new_[3584]_  | ~\new_[3585]_ );
  assign n1865 = ~\new_[12794]_  & (~\new_[3586]_  | ~\new_[3587]_ );
  assign \new_[3120]_  = ~\new_[14822]_ ;
  assign n1880 = \new_[12271]_  & \new_[3407]_ ;
  assign n1890 = \new_[3396]_  | \new_[3408]_ ;
  assign n1810 = \new_[3397]_  | \new_[3408]_ ;
  assign \new_[3124]_  = \new_[3395]_  | \new_[4801]_ ;
  assign n1895 = \new_[12526]_  & \new_[3401]_ ;
  assign \new_[3126]_  = ~\new_[2373]_  | ~n7590 | ~\new_[5710]_  | ~\new_[3794]_ ;
  assign n1905 = \new_[5984]_  ^ \new_[3591]_ ;
  assign n1900 = \new_[6230]_  ^ \new_[14613]_ ;
  assign \new_[3129]_  = ~\new_[3279]_  & ~\new_[4796]_ ;
  assign n1995 = ~\new_[11675]_  | (~\new_[3632]_  & ~n9145);
  assign \new_[3131]_  = ~\\u4_u0_buf0_reg[9] ;
  assign \new_[3132]_  = ~\\u4_u0_buf0_reg[27] ;
  assign \new_[3133]_  = ~\new_[3555]_  & (~\new_[3618]_  | ~\new_[3764]_ );
  assign \new_[3134]_  = ~\new_[3802]_  | ~\new_[4451]_  | ~\new_[3764]_  | ~\new_[4454]_ ;
  assign n1910 = \new_[4265]_  ^ \new_[3764]_ ;
  assign \new_[3136]_  = ~\new_[3444]_  | (~\new_[6063]_  & ~\new_[4489]_ );
  assign \new_[3137]_  = ~\new_[3555]_  | ~\new_[14526]_ ;
  assign \new_[3138]_  = ~\new_[6081]_  | ~\new_[5858]_  | ~\new_[6114]_  | ~\new_[3672]_ ;
  assign \new_[3139]_  = ~\new_[3545]_  & (~\new_[2833]_  | ~\new_[4154]_ );
  assign \new_[3140]_  = ~\new_[3546]_  & (~\new_[2858]_  | ~\new_[4153]_ );
  assign \new_[3141]_  = ~\new_[3547]_  & (~\new_[2830]_  | ~\new_[4154]_ );
  assign \new_[3142]_  = ~\new_[3548]_  & (~\new_[2859]_  | ~\new_[4154]_ );
  assign \new_[3143]_  = ~\new_[3549]_  & (~\new_[2860]_  | ~\new_[4153]_ );
  assign \new_[3144]_  = ~\new_[3550]_  & (~\new_[2893]_  | ~\new_[4153]_ );
  assign \new_[3145]_  = ~\new_[3551]_  & (~\new_[2896]_  | ~\new_[4153]_ );
  assign \new_[3146]_  = ~\new_[3552]_  & (~\new_[2861]_  | ~\new_[4153]_ );
  assign \new_[3147]_  = \new_[10970]_  ? \new_[4154]_  : \new_[2862]_ ;
  assign \new_[3148]_  = \new_[10979]_  ? \new_[4154]_  : \new_[2863]_ ;
  assign \new_[3149]_  = \new_[10958]_  ? \new_[4154]_  : \new_[2895]_ ;
  assign \new_[3150]_  = \new_[10953]_  ? \new_[4154]_  : \new_[2868]_ ;
  assign \new_[3151]_  = \new_[10964]_  ? \new_[4154]_  : \new_[2864]_ ;
  assign \new_[3152]_  = \new_[10878]_  ? \new_[4154]_  : \new_[2865]_ ;
  assign \new_[3153]_  = \new_[10962]_  ? \new_[4154]_  : \new_[2866]_ ;
  assign \new_[3154]_  = \new_[10980]_  ? \new_[4154]_  : \new_[2867]_ ;
  assign \new_[3155]_  = \new_[4153]_  ^ \new_[2932]_ ;
  assign \new_[3156]_  = ~\\u4_u0_buf0_reg[14] ;
  assign \new_[3157]_  = ~\\u4_u0_buf0_reg[10] ;
  assign \new_[3158]_  = ~\\u4_u0_buf0_reg[13] ;
  assign \new_[3159]_  = ~\\u4_u0_buf1_reg[14] ;
  assign \new_[3160]_  = ~\\u4_u0_buf0_reg[11] ;
  assign \new_[3161]_  = ~\\u4_u0_buf0_reg[15] ;
  assign \new_[3162]_  = ~\\u4_u0_buf0_reg[6] ;
  assign \new_[3163]_  = ~\\u4_u0_buf1_reg[10] ;
  assign \new_[3164]_  = ~\\u4_u0_buf1_reg[13] ;
  assign \new_[3165]_  = ~\\u4_u0_buf0_reg[7] ;
  assign \new_[3166]_  = ~\\u4_u0_buf1_reg[11] ;
  assign \new_[3167]_  = ~\\u4_u0_buf1_reg[15] ;
  assign \new_[3168]_  = ~\\u4_u0_buf1_reg[6] ;
  assign \new_[3169]_  = ~\\u4_u0_buf1_reg[4] ;
  assign \new_[3170]_  = ~\\u4_u0_buf1_reg[5] ;
  assign \new_[3171]_  = ~\\u4_u0_buf1_reg[7] ;
  assign \new_[3172]_  = \\u1_hms_cnt_reg[0] ;
  assign \new_[3173]_  = \\u1_u3_idin_reg[19] ;
  assign \new_[3174]_  = \\u1_u3_new_size_reg[5] ;
  assign \new_[3175]_  = ~\\u4_u0_buf1_reg[28] ;
  assign \new_[3176]_  = ~\\u4_u0_buf1_reg[31] ;
  assign \new_[3177]_  = \\u1_u2_state_reg[3] ;
  assign \new_[3178]_  = ~\\u4_u0_buf0_reg[0] ;
  assign \new_[3179]_  = ~\\u4_u0_buf0_reg[18] ;
  assign \new_[3180]_  = ~\\u4_u0_buf0_reg[19] ;
  assign \new_[3181]_  = ~\\u4_u0_buf0_reg[1] ;
  assign \new_[3182]_  = ~\\u4_u0_buf0_reg[20] ;
  assign \new_[3183]_  = ~\\u4_u0_buf0_reg[21] ;
  assign \new_[3184]_  = ~\\u4_u0_buf0_reg[23] ;
  assign \new_[3185]_  = ~\\u4_u0_buf0_reg[24] ;
  assign \new_[3186]_  = ~\\u4_u0_buf0_reg[25] ;
  assign \new_[3187]_  = ~\\u4_u0_buf0_reg[26] ;
  assign \new_[3188]_  = ~\\u4_u0_buf0_reg[30] ;
  assign \new_[3189]_  = ~\\u4_u0_buf0_reg[3] ;
  assign \new_[3190]_  = ~\\u4_u0_buf0_reg[8] ;
  assign \new_[3191]_  = ~\\u4_u1_buf0_reg[28] ;
  assign \new_[3192]_  = ~\\u4_u1_buf0_reg[31] ;
  assign \new_[3193]_  = ~\new_[11463]_  | ~\new_[4337]_ ;
  assign \new_[3194]_  = \new_[4337]_  | \new_[12130]_ ;
  assign \sram_adr_o[14]  = \new_[2085]_  ? \new_[3611]_  : \wb_addr_i[16] ;
  assign \sram_adr_o[13]  = \new_[2084]_  ? \new_[3608]_  : \wb_addr_i[15] ;
  assign \sram_adr_o[12]  = \new_[2095]_  ? \new_[3603]_  : \wb_addr_i[14] ;
  assign \sram_adr_o[11]  = \new_[2083]_  ? \new_[3603]_  : \wb_addr_i[13] ;
  assign \sram_adr_o[10]  = \new_[2094]_  ? \new_[3609]_  : \wb_addr_i[12] ;
  assign \sram_adr_o[9]  = \new_[2097]_  ? \new_[3610]_  : \wb_addr_i[11] ;
  assign \sram_adr_o[8]  = \new_[2089]_  ? \new_[3605]_  : \wb_addr_i[10] ;
  assign \sram_adr_o[7]  = \new_[2088]_  ? \new_[3605]_  : \wb_addr_i[9] ;
  assign \sram_adr_o[6]  = \new_[2087]_  ? \new_[3613]_  : \wb_addr_i[8] ;
  assign \sram_adr_o[5]  = \new_[2086]_  ? \new_[3607]_  : \wb_addr_i[7] ;
  assign \sram_adr_o[4]  = \new_[2093]_  ? \new_[3612]_  : \wb_addr_i[6] ;
  assign \sram_adr_o[3]  = \new_[2091]_  ? \new_[3603]_  : \wb_addr_i[5] ;
  assign \sram_adr_o[2]  = \new_[2092]_  ? \new_[3603]_  : \wb_addr_i[4] ;
  assign \sram_adr_o[1]  = \new_[2096]_  ? \new_[3609]_  : \wb_addr_i[3] ;
  assign \sram_adr_o[0]  = \new_[2090]_  ? \new_[3607]_  : \wb_addr_i[2] ;
  assign \sram_data_o[31]  = \new_[2663]_  ? \new_[3612]_  : \wb_data_i[31] ;
  assign \sram_data_o[30]  = \new_[2619]_  ? \new_[3609]_  : \wb_data_i[30] ;
  assign \sram_data_o[29]  = \new_[2661]_  ? \new_[3613]_  : \wb_data_i[29] ;
  assign \sram_data_o[28]  = \new_[2660]_  ? \new_[3612]_  : \wb_data_i[28] ;
  assign \sram_data_o[27]  = \new_[2623]_  ? \new_[3613]_  : \wb_data_i[27] ;
  assign \sram_data_o[26]  = \new_[2659]_  ? \new_[3605]_  : \wb_data_i[26] ;
  assign \sram_data_o[25]  = \new_[2658]_  ? \new_[3613]_  : \wb_data_i[25] ;
  assign \sram_data_o[24]  = \new_[2657]_  ? \new_[3610]_  : \wb_data_i[24] ;
  assign \sram_data_o[23]  = \new_[2656]_  ? \new_[3608]_  : \wb_data_i[23] ;
  assign \sram_data_o[22]  = \new_[2655]_  ? \new_[3608]_  : \wb_data_i[22] ;
  assign \sram_data_o[21]  = \new_[2654]_  ? \new_[3603]_  : \wb_data_i[21] ;
  assign \sram_data_o[20]  = \new_[2653]_  ? \new_[3603]_  : \wb_data_i[20] ;
  assign \sram_data_o[19]  = \new_[2652]_  ? \new_[3605]_  : \wb_data_i[19] ;
  assign \sram_data_o[18]  = \new_[2651]_  ? \new_[3608]_  : \wb_data_i[18] ;
  assign \sram_data_o[17]  = \new_[2650]_  ? \new_[3603]_  : \wb_data_i[17] ;
  assign \sram_data_o[16]  = \new_[2625]_  ? \new_[3606]_  : \wb_data_i[16] ;
  assign \sram_data_o[15]  = \new_[2649]_  ? \new_[3611]_  : \wb_data_i[15] ;
  assign \sram_data_o[14]  = \new_[2648]_  ? \new_[3603]_  : \wb_data_i[14] ;
  assign \sram_data_o[13]  = \new_[2647]_  ? \new_[3603]_  : \wb_data_i[13] ;
  assign \sram_data_o[12]  = \new_[2645]_  ? \new_[3609]_  : \wb_data_i[12] ;
  assign \sram_data_o[11]  = \new_[2646]_  ? \new_[3603]_  : \wb_data_i[11] ;
  assign \sram_data_o[10]  = \new_[2644]_  ? \new_[3606]_  : \wb_data_i[10] ;
  assign \sram_data_o[9]  = \new_[2669]_  ? \new_[3612]_  : \wb_data_i[9] ;
  assign \sram_data_o[8]  = \new_[2668]_  ? \new_[3611]_  : \wb_data_i[8] ;
  assign \sram_data_o[7]  = \new_[2667]_  ? \new_[3610]_  : \wb_data_i[7] ;
  assign \sram_data_o[6]  = \new_[2666]_  ? \new_[3611]_  : \wb_data_i[6] ;
  assign \sram_data_o[5]  = \new_[2622]_  ? \new_[3603]_  : \wb_data_i[5] ;
  assign \sram_data_o[4]  = \new_[2665]_  ? \new_[3607]_  : \wb_data_i[4] ;
  assign \sram_data_o[3]  = \new_[2664]_  ? \new_[3607]_  : \wb_data_i[3] ;
  assign \sram_data_o[2]  = \new_[2662]_  ? \new_[3606]_  : \wb_data_i[2] ;
  assign \sram_data_o[1]  = \new_[2624]_  ? \new_[3606]_  : \wb_data_i[1] ;
  assign \sram_data_o[0]  = \new_[2643]_  ? \new_[3610]_  : \wb_data_i[0] ;
  assign \new_[3242]_  = u1_u3_match_r_reg;
  assign \new_[3243]_  = \new_[3573]_  | \new_[4148]_ ;
  assign \new_[3244]_  = ~\new_[3387]_ ;
  assign \new_[3245]_  = ~\\u1_u3_new_size_reg[8] ;
  assign n1925 = ~\new_[10718]_  & ~\new_[3566]_ ;
  assign n1930 = \new_[3782]_  ? n9145 : \new_[2873]_ ;
  assign \new_[3248]_  = ~\new_[14775]_ ;
  assign n1970 = ~\new_[14321]_  & ~\new_[14000]_ ;
  assign n1985 = ~\new_[10845]_  & ~\new_[14321]_ ;
  assign n1990 = ~\new_[10622]_  & ~\new_[14321]_ ;
  assign n2040 = ~\new_[10624]_  & ~\new_[14321]_ ;
  assign \new_[3253]_  = ~\new_[3604]_  | ~\new_[5032]_  | ~\new_[4480]_ ;
  assign n1935 = \new_[12791]_  & \new_[3572]_ ;
  assign n1940 = \new_[11403]_  & \new_[3572]_ ;
  assign n1945 = \new_[10313]_  & \new_[3572]_ ;
  assign n1950 = \new_[9607]_  & \new_[3572]_ ;
  assign n1955 = \new_[9103]_  & \new_[3572]_ ;
  assign n1915 = \new_[9648]_  & \new_[3572]_ ;
  assign n1960 = \new_[8675]_  & \new_[3572]_ ;
  assign n1965 = \new_[8947]_  & \new_[3572]_ ;
  assign n1975 = ~\new_[11056]_  & ~\new_[14321]_ ;
  assign n2035 = ~\new_[10959]_  & ~\new_[14321]_ ;
  assign n1980 = ~\new_[10493]_  & ~\new_[14321]_ ;
  assign \new_[3265]_  = ~\new_[12728]_  | ~\new_[3038]_  | ~\new_[3601]_  | ~\new_[13476]_ ;
  assign \new_[3266]_  = ~u5_wb_ack_s2_reg;
  assign \new_[3267]_  = ~\\u1_u3_new_size_reg[7] ;
  assign n2005 = ~\new_[3602]_  & (~\new_[12583]_  | ~\new_[11774]_ );
  assign n2000 = ~\new_[12397]_  & ~\new_[3602]_ ;
  assign n2010 = ~\new_[9632]_  & ~\new_[3602]_ ;
  assign n2015 = ~\new_[9593]_  & ~\new_[3602]_ ;
  assign n1920 = ~\new_[9081]_  & ~\new_[3602]_ ;
  assign n2030 = ~\new_[9406]_  & ~\new_[3602]_ ;
  assign n2020 = ~\new_[9035]_  & ~\new_[3602]_ ;
  assign n2025 = ~\new_[9165]_  & ~\new_[3602]_ ;
  assign \new_[3276]_  = ~\new_[3630]_  & ~wb_ack_o;
  assign \new_[3277]_  = ~\new_[9882]_  & ~\new_[4154]_ ;
  assign \new_[3278]_  = \new_[3632]_  | \new_[4796]_ ;
  assign \new_[3279]_  = \new_[4013]_  | \new_[3632]_ ;
  assign \new_[3280]_  = ~\\u4_u1_buf0_reg[8] ;
  assign \new_[3281]_  = ~\\u4_u1_buf1_reg[6] ;
  assign \new_[3282]_  = \\u4_u2_dma_in_cnt_reg[9] ;
  assign \new_[3283]_  = \\u4_u3_dma_in_cnt_reg[9] ;
  assign n2050 = \new_[4285]_  ? n9145 : \new_[2870]_ ;
  assign \new_[3285]_  = ~\\u4_u0_buf1_reg[3] ;
  assign \new_[3286]_  = ~\\u1_u2_last_buf_adr_reg[1] ;
  assign n2045 = ~\new_[4717]_  | ~phy_rst_pad_o | ~\new_[3600]_  | ~\new_[7940]_ ;
  assign \new_[3288]_  = ~\\u4_u1_buf0_reg[6] ;
  assign \new_[3289]_  = ~\new_[6566]_  | ~\new_[6071]_  | ~\new_[6617]_  | ~\new_[3859]_ ;
  assign \new_[3290]_  = ~\new_[6589]_  | ~\new_[6072]_  | ~\new_[6618]_  | ~\new_[3860]_ ;
  assign \new_[3291]_  = ~\new_[9397]_  & ~\new_[4154]_ ;
  assign \new_[3292]_  = ~\\u4_u1_buf0_reg[14] ;
  assign \new_[3293]_  = ~\\u4_u1_buf0_reg[10] ;
  assign \new_[3294]_  = ~\\u4_u1_buf0_reg[13] ;
  assign \new_[3295]_  = ~\\u4_u1_buf1_reg[14] ;
  assign \new_[3296]_  = ~\\u4_u1_buf0_reg[11] ;
  assign \new_[3297]_  = ~\\u4_u1_buf0_reg[15] ;
  assign \new_[3298]_  = ~\\u4_u1_buf1_reg[10] ;
  assign \new_[3299]_  = ~\\u4_u1_buf1_reg[13] ;
  assign \new_[3300]_  = ~\\u4_u1_buf0_reg[7] ;
  assign \new_[3301]_  = ~\\u4_u1_buf1_reg[11] ;
  assign \new_[3302]_  = ~\\u4_u1_buf1_reg[15] ;
  assign \new_[3303]_  = ~\\u4_u1_buf1_reg[4] ;
  assign \new_[3304]_  = ~\\u4_u1_buf1_reg[7] ;
  assign \new_[3305]_  = ~\\u4_u1_buf1_reg[5] ;
  assign \new_[3306]_  = ~\\u4_u0_buf1_reg[29] ;
  assign \new_[3307]_  = ~\\u4_u0_buf1_reg[21] ;
  assign \new_[3308]_  = \\u4_u0_dma_in_cnt_reg[9] ;
  assign \new_[3309]_  = \\u4_u1_dma_in_cnt_reg[9] ;
  assign \new_[3310]_  = \\u4_u0_dma_in_cnt_reg[11] ;
  assign \new_[3311]_  = \\u1_u0_state_reg[2] ;
  assign \new_[3312]_  = \\u4_u0_dma_out_cnt_reg[11] ;
  assign \new_[3313]_  = \\u4_u0_dma_out_cnt_reg[9] ;
  assign \new_[3314]_  = u4_dma_in_buf_sz1_reg;
  assign \new_[3315]_  = \\u4_u0_dma_in_cnt_reg[7] ;
  assign \new_[3316]_  = \\u4_u0_dma_in_cnt_reg[6] ;
  assign \new_[3317]_  = \\u4_u0_dma_out_cnt_reg[6] ;
  assign \new_[3318]_  = ~\\u4_u0_buf1_reg[0] ;
  assign \new_[3319]_  = ~\\u4_u0_buf1_reg[12] ;
  assign \new_[3320]_  = ~\\u4_u0_buf1_reg[16] ;
  assign \new_[3321]_  = ~\\u4_u0_buf1_reg[17] ;
  assign \new_[3322]_  = ~\\u4_u0_buf1_reg[19] ;
  assign \new_[3323]_  = ~\\u4_u0_buf1_reg[1] ;
  assign \new_[3324]_  = ~\\u4_u0_buf1_reg[20] ;
  assign \new_[3325]_  = ~\\u4_u0_buf1_reg[22] ;
  assign \new_[3326]_  = ~\\u4_u0_buf1_reg[24] ;
  assign \new_[3327]_  = ~\\u4_u0_buf1_reg[25] ;
  assign \new_[3328]_  = ~\\u4_u0_buf1_reg[23] ;
  assign \new_[3329]_  = ~\\u4_u0_buf1_reg[27] ;
  assign \new_[3330]_  = ~\\u4_u0_buf1_reg[26] ;
  assign \new_[3331]_  = ~\\u4_u0_buf1_reg[2] ;
  assign \new_[3332]_  = ~\\u4_u0_buf1_reg[30] ;
  assign \new_[3333]_  = ~\\u4_u0_buf1_reg[8] ;
  assign \new_[3334]_  = ~\\u4_u0_buf1_reg[9] ;
  assign \new_[3335]_  = ~\\u4_u1_buf1_reg[28] ;
  assign \new_[3336]_  = ~\\u4_u1_buf1_reg[31] ;
  assign \new_[3337]_  = \\u4_u0_dma_in_cnt_reg[0] ;
  assign \new_[3338]_  = \\u1_u2_state_reg[4] ;
  assign \new_[3339]_  = \\u4_u0_dma_out_cnt_reg[0] ;
  assign \new_[3340]_  = \\u4_u0_dma_out_cnt_reg[1] ;
  assign \new_[3341]_  = \\u4_u0_dma_out_cnt_reg[2] ;
  assign \new_[3342]_  = \\u4_u0_dma_out_cnt_reg[3] ;
  assign \new_[3343]_  = ~\\u4_u1_buf0_reg[16] ;
  assign \new_[3344]_  = ~\\u4_u1_buf0_reg[18] ;
  assign \new_[3345]_  = ~\\u4_u1_buf0_reg[19] ;
  assign \new_[3346]_  = ~\\u4_u1_buf0_reg[1] ;
  assign \new_[3347]_  = ~\\u4_u1_buf0_reg[20] ;
  assign \new_[3348]_  = ~\\u4_u1_buf0_reg[21] ;
  assign \new_[3349]_  = ~\\u4_u1_buf0_reg[23] ;
  assign \new_[3350]_  = ~\\u4_u1_buf0_reg[24] ;
  assign \new_[3351]_  = ~\\u4_u1_buf0_reg[25] ;
  assign \new_[3352]_  = ~\\u4_u1_buf0_reg[27] ;
  assign \new_[3353]_  = ~\\u4_u1_buf0_reg[30] ;
  assign \new_[3354]_  = ~\\u4_u1_buf0_reg[3] ;
  assign \new_[3355]_  = ~\\u4_u1_buf0_reg[9] ;
  assign \new_[3356]_  = ~\\u4_u2_buf0_reg[28] ;
  assign \new_[3357]_  = ~\\u4_u2_buf0_reg[31] ;
  assign \new_[3358]_  = \new_[3763]_  | \new_[11023]_ ;
  assign \new_[3359]_  = ~\new_[4154]_  | ~\new_[2870]_ ;
  assign \new_[3360]_  = ~\new_[11035]_  & ~\new_[4154]_ ;
  assign \new_[3361]_  = ~\new_[10665]_  & ~\new_[4154]_ ;
  assign \new_[3362]_  = ~\new_[10118]_  & ~\new_[4154]_ ;
  assign \new_[3363]_  = ~\new_[10065]_  & ~\new_[4154]_ ;
  assign \new_[3364]_  = ~\new_[10071]_  & ~\new_[4154]_ ;
  assign \new_[3365]_  = ~\new_[10286]_  & ~\new_[4154]_ ;
  assign \new_[3366]_  = ~\new_[9492]_  & ~\new_[4154]_ ;
  assign \new_[3367]_  = ~\new_[14314]_  & ~\new_[4154]_ ;
  assign n2055 = ~\new_[8357]_  | ~\new_[13165]_  | ~\new_[3800]_ ;
  assign n2060 = ~\new_[8362]_  | ~\new_[12197]_  | ~\new_[3801]_ ;
  assign \new_[3370]_  = ~\new_[4154]_  & (~\new_[10925]_  | ~\new_[10897]_ );
  assign \new_[3371]_  = ~\new_[4154]_  & (~\new_[10929]_  | ~\new_[10917]_ );
  assign \new_[3372]_  = ~\new_[4154]_  & (~\new_[10926]_  | ~\new_[10900]_ );
  assign \new_[3373]_  = ~\new_[4154]_  & (~\new_[10920]_  | ~\new_[10908]_ );
  assign \new_[3374]_  = ~\new_[4154]_  & (~\new_[10921]_  | ~\new_[10894]_ );
  assign \new_[3375]_  = ~\new_[4154]_  & (~\new_[10932]_  | ~\new_[10918]_ );
  assign \new_[3376]_  = ~\new_[4153]_  & (~\new_[10931]_  | ~\new_[10905]_ );
  assign \new_[3377]_  = ~\new_[14412]_  | ~\new_[6464]_ ;
  assign \new_[3378]_  = ~\new_[4153]_  & (~\new_[10909]_  | ~\new_[10923]_ );
  assign \new_[3379]_  = ~\new_[10671]_  & ~\new_[4153]_ ;
  assign \new_[3380]_  = ~\new_[10567]_  & ~\new_[4153]_ ;
  assign \new_[3381]_  = ~\new_[10565]_  & ~\new_[4153]_ ;
  assign \new_[3382]_  = ~\new_[10670]_  & ~\new_[4153]_ ;
  assign \new_[3383]_  = ~\new_[10563]_  & ~\new_[4153]_ ;
  assign \new_[3384]_  = ~\new_[10564]_  & ~\new_[4153]_ ;
  assign \new_[3385]_  = ~\new_[10562]_  & ~\new_[4153]_ ;
  assign \new_[3386]_  = ~\new_[10655]_  & ~\new_[4153]_ ;
  assign \new_[3387]_  = ~u1_frame_no_same_reg;
  assign \new_[3388]_  = ~\new_[3775]_  | ~\new_[4229]_ ;
  assign \new_[3389]_  = ~\new_[3776]_  | ~\new_[5098]_ ;
  assign \new_[3390]_  = ~\\u4_u0_buf1_reg[18] ;
  assign \new_[3391]_  = ~\new_[3566]_ ;
  assign \new_[3392]_  = ~\new_[3782]_  | ~\new_[13646]_ ;
  assign \new_[3393]_  = \new_[3782]_  | \new_[3174]_ ;
  assign \new_[3394]_  = ~\new_[3782]_  | ~\new_[3174]_ ;
  assign \new_[3395]_  = ~\\u1_u3_new_size_reg[6] ;
  assign \new_[3396]_  = ~\new_[3602]_  & (~\new_[11459]_  | ~\new_[13606]_ );
  assign \new_[3397]_  = ~\new_[10983]_  & ~\new_[3602]_ ;
  assign \new_[3398]_  = ~\new_[3571]_ ;
  assign \new_[3399]_  = ~\\u4_u1_buf0_reg[26] ;
  assign \new_[3400]_  = \new_[3604]_  | \new_[11687]_ ;
  assign \new_[3401]_  = ~\new_[14321]_ ;
  assign \new_[3402]_  = ~\new_[3967]_  | ~\new_[6718]_ ;
  assign \new_[3403]_  = ~\new_[3967]_  | ~\new_[6018]_ ;
  assign \new_[3404]_  = ~\new_[3967]_  | ~\new_[12396]_ ;
  assign \new_[3405]_  = ~\new_[3967]_  | ~\new_[6696]_ ;
  assign \new_[3406]_  = ~\new_[3967]_  | ~\new_[6716]_ ;
  assign \new_[3407]_  = ~\new_[3602]_  & (~\new_[12250]_  | ~\new_[11731]_ );
  assign \new_[3408]_  = ~\new_[3602]_  & (~\new_[12728]_  | ~\new_[12510]_ );
  assign n2075 = ~\new_[8342]_  | ~\new_[12258]_  | ~\new_[4162]_ ;
  assign \new_[3410]_  = \\u1_sof_time_reg[2] ;
  assign n2160 = ~\new_[11662]_  | (~\new_[4013]_  & ~n9145);
  assign n2270 = u5_wb_ack_s1a_reg;
  assign \new_[3413]_  = ~\new_[5721]_  | (~\new_[4057]_  & ~\new_[6220]_ );
  assign \new_[3414]_  = ~\new_[3822]_  & (~\new_[4285]_  | ~\new_[14546]_ );
  assign n2120 = ~\new_[12067]_  | ~\new_[8368]_  | ~\new_[4151]_ ;
  assign \new_[3416]_  = ~\\u4_u0_buf0_reg[2] ;
  assign n2125 = ~\new_[3829]_  | ~phy_rst_pad_o;
  assign n2130 = ~\new_[3830]_  | ~phy_rst_pad_o;
  assign n2135 = ~\new_[3831]_  | ~phy_rst_pad_o;
  assign \new_[3420]_  = ~\new_[3617]_ ;
  assign \new_[3421]_  = ~\\u4_u2_buf0_reg[8] ;
  assign \new_[3422]_  = ~\\u4_u3_buf0_reg[31] ;
  assign \new_[3423]_  = ~\\u4_u0_buf0_reg[22] ;
  assign \new_[3424]_  = ~\\u4_u2_buf0_reg[12] ;
  assign \new_[3425]_  = ~\\u4_u1_buf1_reg[1] ;
  assign n2165 = \new_[5988]_  ^ \new_[14614]_ ;
  assign n2275 = \new_[6228]_  ^ \new_[4029]_ ;
  assign \new_[3428]_  = \\u4_u0_dma_out_cnt_reg[8] ;
  assign \new_[3429]_  = \\u4_u0_dma_out_cnt_reg[4] ;
  assign \new_[3430]_  = ~\\u4_u1_buf1_reg[9] ;
  assign \new_[3431]_  = ~\\u4_u2_buf0_reg[19] ;
  assign \new_[3432]_  = ~\\u4_u1_buf1_reg[27] ;
  assign \new_[3433]_  = ~\\u4_u1_buf1_reg[23] ;
  assign \new_[3434]_  = ~\\u4_u0_buf0_reg[5] ;
  assign \new_[3435]_  = \\u1_sof_time_reg[6] ;
  assign n2210 = ~\new_[8350]_  | ~\new_[12255]_  | ~\new_[3987]_ ;
  assign n2095 = ~\new_[8339]_  | ~\new_[12486]_  | ~\new_[3970]_ ;
  assign n2100 = ~\new_[8343]_  | ~\new_[12339]_  | ~\new_[3971]_ ;
  assign \new_[3439]_  = ~\\u4_u2_buf0_reg[6] ;
  assign \new_[3440]_  = ~\\u4_u2_buf0_reg[11] ;
  assign n2105 = ~\new_[8367]_  | ~\new_[13165]_  | ~\new_[3975]_ ;
  assign \new_[3442]_  = ~\\u4_u2_buf0_reg[10] ;
  assign n2110 = ~\new_[3924]_  | ~phy_rst_pad_o;
  assign \new_[3444]_  = ~\new_[6852]_  | ~\new_[6542]_  | ~\new_[6894]_  | ~\new_[4060]_ ;
  assign n2170 = ~\new_[3920]_  | ~phy_rst_pad_o;
  assign n2175 = ~\new_[3921]_  | ~phy_rst_pad_o;
  assign \new_[3447]_  = \new_[4157]_  ^ \new_[8632]_ ;
  assign \new_[3448]_  = ~\\u4_u2_buf0_reg[14] ;
  assign \new_[3449]_  = ~\\u4_u2_buf0_reg[13] ;
  assign \new_[3450]_  = ~\\u4_u2_buf1_reg[14] ;
  assign \new_[3451]_  = ~\\u4_u2_buf0_reg[15] ;
  assign \new_[3452]_  = ~\\u4_u2_buf1_reg[10] ;
  assign \new_[3453]_  = ~\\u4_u2_buf1_reg[13] ;
  assign \new_[3454]_  = ~\\u4_u0_buf0_reg[4] ;
  assign \new_[3455]_  = ~\\u4_u2_buf0_reg[7] ;
  assign \new_[3456]_  = ~\\u4_u2_buf1_reg[11] ;
  assign \new_[3457]_  = ~\\u4_u2_buf1_reg[6] ;
  assign \new_[3458]_  = ~\\u4_u2_buf1_reg[4] ;
  assign \new_[3459]_  = ~\\u4_u2_buf1_reg[5] ;
  assign \new_[3460]_  = ~\\u4_u2_buf1_reg[7] ;
  assign \new_[3461]_  = ~\\u1_sof_time_reg[11] ;
  assign \new_[3462]_  = \\u4_u0_dma_in_cnt_reg[8] ;
  assign \new_[3463]_  = \\u1_sof_time_reg[7] ;
  assign \new_[3464]_  = \\u4_u1_dma_in_cnt_reg[11] ;
  assign \new_[3465]_  = \\u1_sof_time_reg[0] ;
  assign \new_[3466]_  = \\u4_u0_dma_in_cnt_reg[10] ;
  assign \new_[3467]_  = \\u4_u1_dma_out_cnt_reg[11] ;
  assign \new_[3468]_  = \\u4_u1_dma_out_cnt_reg[9] ;
  assign \new_[3469]_  = \\u1_sof_time_reg[10] ;
  assign \new_[3470]_  = \\u1_sof_time_reg[1] ;
  assign \new_[3471]_  = \\u1_sof_time_reg[3] ;
  assign \new_[3472]_  = \\u1_sof_time_reg[4] ;
  assign \new_[3473]_  = \\u1_sof_time_reg[5] ;
  assign \new_[3474]_  = \\u1_sof_time_reg[9] ;
  assign \new_[3475]_  = \\u1_sof_time_reg[8] ;
  assign \new_[3476]_  = \\u4_u0_dma_in_cnt_reg[5] ;
  assign \new_[3477]_  = \\u4_u0_dma_out_cnt_reg[10] ;
  assign \new_[3478]_  = \\u4_u0_dma_out_cnt_reg[7] ;
  assign \new_[3479]_  = \\u4_u1_dma_in_cnt_reg[7] ;
  assign \new_[3480]_  = \\u4_u0_dma_in_cnt_reg[4] ;
  assign \new_[3481]_  = \\u4_u1_dma_in_cnt_reg[6] ;
  assign \new_[3482]_  = \\u4_u1_dma_out_cnt_reg[6] ;
  assign \new_[3483]_  = ~\\u4_u1_buf1_reg[0] ;
  assign \new_[3484]_  = ~\\u4_u1_buf1_reg[12] ;
  assign \new_[3485]_  = ~\\u4_u1_buf1_reg[16] ;
  assign \new_[3486]_  = ~\\u4_u1_buf1_reg[17] ;
  assign \new_[3487]_  = ~\\u4_u1_buf1_reg[18] ;
  assign \new_[3488]_  = ~\\u4_u1_buf1_reg[19] ;
  assign \new_[3489]_  = ~\\u4_u1_buf1_reg[20] ;
  assign \new_[3490]_  = ~\\u4_u1_buf1_reg[21] ;
  assign \new_[3491]_  = ~\\u4_u1_buf1_reg[22] ;
  assign \new_[3492]_  = ~\\u4_u1_buf1_reg[24] ;
  assign \new_[3493]_  = ~\\u4_u1_buf1_reg[25] ;
  assign \new_[3494]_  = ~\\u4_u1_buf1_reg[26] ;
  assign \new_[3495]_  = ~\\u4_u1_buf1_reg[2] ;
  assign \new_[3496]_  = ~\\u4_u1_buf1_reg[30] ;
  assign \new_[3497]_  = ~\\u4_u1_buf1_reg[29] ;
  assign \new_[3498]_  = ~\\u4_u1_buf1_reg[3] ;
  assign \new_[3499]_  = ~\\u4_u1_buf1_reg[8] ;
  assign \new_[3500]_  = ~\\u4_u2_buf1_reg[28] ;
  assign \new_[3501]_  = ~\\u4_u2_buf1_reg[31] ;
  assign \new_[3502]_  = \\u4_u1_dma_in_cnt_reg[0] ;
  assign \new_[3503]_  = \\u4_u0_dma_in_cnt_reg[1] ;
  assign \new_[3504]_  = \\u4_u0_dma_in_cnt_reg[2] ;
  assign \new_[3505]_  = \\u4_u0_dma_in_cnt_reg[3] ;
  assign \new_[3506]_  = \\u4_u0_dma_out_cnt_reg[5] ;
  assign \new_[3507]_  = \\u4_u1_dma_out_cnt_reg[0] ;
  assign \new_[3508]_  = \\u4_u1_dma_out_cnt_reg[1] ;
  assign \new_[3509]_  = \\u4_u1_dma_out_cnt_reg[2] ;
  assign \new_[3510]_  = \\u4_u1_dma_out_cnt_reg[3] ;
  assign \new_[3511]_  = ~\\u4_u3_buf0_reg[28] ;
  assign \new_[3512]_  = ~\\u4_u0_buf0_reg[12] ;
  assign \new_[3513]_  = ~\\u4_u0_buf0_reg[16] ;
  assign \new_[3514]_  = ~\\u4_u0_buf0_reg[17] ;
  assign \new_[3515]_  = ~\\u4_u0_buf0_reg[29] ;
  assign \new_[3516]_  = ~\\u4_u2_buf0_reg[0] ;
  assign \new_[3517]_  = ~\\u4_u2_buf0_reg[16] ;
  assign \new_[3518]_  = ~\\u4_u2_buf0_reg[17] ;
  assign \new_[3519]_  = ~\\u4_u2_buf0_reg[18] ;
  assign \new_[3520]_  = ~\\u4_u2_buf0_reg[20] ;
  assign \new_[3521]_  = ~\\u4_u2_buf0_reg[22] ;
  assign \new_[3522]_  = ~\\u4_u2_buf0_reg[24] ;
  assign \new_[3523]_  = ~\\u4_u2_buf0_reg[25] ;
  assign \new_[3524]_  = ~\\u4_u2_buf0_reg[29] ;
  assign \new_[3525]_  = ~\\u4_u2_buf0_reg[1] ;
  assign \new_[3526]_  = ~\\u4_u2_buf0_reg[30] ;
  assign \new_[3527]_  = ~\\u4_u2_buf0_reg[3] ;
  assign n2080 = ~\new_[8337]_  | ~\new_[12158]_  | ~\new_[4024]_ ;
  assign n2180 = \new_[3937]_  & \new_[12197]_ ;
  assign n2185 = ~\new_[8336]_  | ~\new_[12255]_  | ~\new_[3981]_ ;
  assign \new_[3531]_  = ~\new_[5924]_  & (~\new_[4129]_  | ~\new_[5922]_ );
  assign n2195 = ~\new_[8347]_  | ~\new_[12255]_  | ~\new_[3984]_ ;
  assign n2200 = ~\new_[8348]_  | ~\new_[12255]_  | ~\new_[3985]_ ;
  assign n2215 = ~\new_[8352]_  | ~\new_[12158]_  | ~\new_[3988]_ ;
  assign n2220 = ~\new_[8353]_  | ~\new_[12197]_  | ~\new_[3989]_ ;
  assign n2225 = ~\new_[8354]_  | ~\new_[12197]_  | ~\new_[3990]_ ;
  assign n2230 = ~\new_[8355]_  | ~\new_[12197]_  | ~\new_[3991]_ ;
  assign n2070 = ~\new_[8356]_  | ~\new_[12197]_  | ~\new_[3992]_ ;
  assign n2235 = ~\new_[8361]_  | ~\new_[12252]_  | ~\new_[3993]_ ;
  assign n2240 = ~\new_[8363]_  | ~\new_[12197]_  | ~\new_[3994]_ ;
  assign n2245 = ~\new_[8369]_  | ~\new_[13165]_  | ~\new_[3995]_ ;
  assign n2065 = ~\new_[8370]_  | ~\new_[13165]_  | ~\new_[3996]_ ;
  assign n2250 = ~\new_[8501]_  | ~\new_[12491]_  | ~\new_[4000]_ ;
  assign n2255 = ~\new_[8133]_  | ~\new_[12491]_  | ~\new_[4001]_ ;
  assign \new_[3545]_  = ~\new_[4153]_  & (~\new_[10785]_  | ~\new_[10919]_ );
  assign \new_[3546]_  = ~\new_[4153]_  & (~\new_[10934]_  | ~\new_[10733]_ );
  assign \new_[3547]_  = ~\new_[4153]_  & (~\new_[10928]_  | ~\new_[10771]_ );
  assign \new_[3548]_  = ~\new_[4153]_  & (~\new_[10924]_  | ~\new_[10910]_ );
  assign \new_[3549]_  = ~\new_[4153]_  & (~\new_[10922]_  | ~\new_[10884]_ );
  assign \new_[3550]_  = ~\new_[4153]_  & (~\new_[10927]_  | ~\new_[10915]_ );
  assign \new_[3551]_  = ~\new_[4153]_  & (~\new_[10822]_  | ~\new_[10930]_ );
  assign \new_[3552]_  = ~\new_[4153]_  & (~\new_[10901]_  | ~\new_[10935]_ );
  assign \new_[3553]_  = ~\new_[3765]_ ;
  assign \new_[3554]_  = ~\new_[5082]_  | ~\new_[3935]_  | ~\new_[4451]_ ;
  assign \new_[3555]_  = \new_[3929]_  | \new_[14525]_ ;
  assign \new_[3556]_  = ~\new_[3936]_  | (~\new_[4232]_  & ~\new_[4260]_ );
  assign n2190 = ~\new_[8346]_  | ~\new_[12258]_  | ~\new_[3983]_ ;
  assign n2115 = ~\new_[3818]_  | ~phy_rst_pad_o;
  assign n2260 = ~\new_[14412]_ ;
  assign n2140 = ~\new_[3958]_  | ~phy_rst_pad_o;
  assign n2145 = ~\new_[3959]_  | ~\new_[12058]_ ;
  assign n2150 = ~\new_[3960]_  | ~phy_rst_pad_o;
  assign \new_[3563]_  = ~\new_[3805]_  | ~\new_[4451]_ ;
  assign \new_[3564]_  = ~\\u4_u2_buf1_reg[15] ;
  assign n2155 = ~\new_[13296]_  & ~\new_[3944]_  & ~\new_[3172]_ ;
  assign \new_[3566]_  = \new_[3944]_  | \new_[12368]_ ;
  assign n2085 = ~\new_[8341]_  | ~\new_[12244]_  | ~\new_[4128]_ ;
  assign n2090 = ~\new_[3862]_  | ~phy_rst_pad_o;
  assign n2205 = ~\new_[8349]_  | ~\new_[12067]_  | ~\new_[3986]_ ;
  assign n2265 = \new_[6229]_  ^ \new_[3977]_ ;
  assign \new_[3571]_  = ~\new_[14274]_  | ~\new_[3797]_  | ~n4870;
  assign \new_[3572]_  = ~\new_[14326]_  & ~\new_[9645]_ ;
  assign \new_[3573]_  = \new_[3794]_  | \new_[2611]_ ;
  assign \new_[3574]_  = ~\new_[3967]_  | ~\new_[6015]_ ;
  assign \new_[3575]_  = ~\new_[4191]_  | ~\new_[2983]_ ;
  assign \new_[3576]_  = ~\new_[4191]_  | ~\new_[2924]_ ;
  assign \new_[3577]_  = ~\new_[4191]_  | ~\new_[2985]_ ;
  assign \new_[3578]_  = ~\new_[3967]_  | ~\new_[6016]_ ;
  assign \new_[3579]_  = ~\new_[3967]_  | ~\new_[6033]_ ;
  assign \new_[3580]_  = ~\new_[4191]_  | ~\new_[2986]_ ;
  assign \new_[3581]_  = ~\new_[4191]_  | ~\new_[2984]_ ;
  assign \new_[3582]_  = ~\new_[3967]_  | ~\new_[6017]_ ;
  assign \new_[3583]_  = ~\new_[4191]_  | ~\new_[2925]_ ;
  assign \new_[3584]_  = ~\new_[3967]_  | ~\new_[6019]_ ;
  assign \new_[3585]_  = ~\new_[4191]_  | ~\new_[2962]_ ;
  assign \new_[3586]_  = ~\new_[3967]_  | ~\new_[5978]_ ;
  assign \new_[3587]_  = ~\new_[4191]_  | ~\new_[2987]_ ;
  assign \new_[3588]_  = ~\new_[4191]_  | ~\new_[2926]_ ;
  assign \new_[3589]_  = ~\new_[4191]_  | ~\new_[2927]_ ;
  assign \new_[3590]_  = ~\new_[4191]_  | ~\new_[2929]_ ;
  assign \new_[3591]_  = ~\new_[7448]_  | ~\new_[4192]_  | ~\new_[3972]_ ;
  assign \new_[3592]_  = \\u4_u1_dma_in_cnt_reg[8] ;
  assign n2315 = ~\new_[8011]_  | ~\new_[13165]_  | ~\new_[4352]_ ;
  assign \new_[3594]_  = ~\\u4_u1_buf0_reg[2] ;
  assign \new_[3595]_  = \\u4_u3_int_stat_reg[0] ;
  assign \new_[3596]_  = ~\\u4_u1_buf0_reg[22] ;
  assign \new_[3597]_  = ~\new_[3794]_ ;
  assign \new_[3598]_  = \new_[4013]_  | \new_[4798]_ ;
  assign \new_[3599]_  = ~\new_[4013]_  & ~\new_[12932]_ ;
  assign \new_[3600]_  = ~\new_[7873]_  & ~\new_[4170]_ ;
  assign \new_[3601]_  = ~\new_[14326]_ ;
  assign \new_[3602]_  = \new_[14322]_ ;
  assign \new_[3603]_  = ~\new_[3798]_ ;
  assign \new_[3604]_  = ~\new_[3798]_ ;
  assign \new_[3605]_  = ~\new_[3798]_ ;
  assign \new_[3606]_  = ~\new_[3798]_ ;
  assign \new_[3607]_  = ~\new_[3798]_ ;
  assign \new_[3608]_  = ~\new_[3798]_ ;
  assign \new_[3609]_  = ~\new_[3798]_ ;
  assign \new_[3610]_  = ~\new_[3798]_ ;
  assign \new_[3611]_  = ~\new_[3798]_ ;
  assign \new_[3612]_  = ~\new_[3798]_ ;
  assign \new_[3613]_  = ~\new_[3798]_ ;
  assign \new_[3614]_  = ~\\u4_u2_buf1_reg[3] ;
  assign \new_[3615]_  = ~\new_[4059]_  | ~\new_[5914]_ ;
  assign \new_[3616]_  = ~\new_[4059]_  & ~\new_[5914]_ ;
  assign \new_[3617]_  = ~\new_[5912]_  & (~\new_[4249]_  | ~\new_[6180]_ );
  assign \new_[3618]_  = \new_[4451]_  & \new_[4031]_ ;
  assign n2355 = ~\new_[8507]_  | ~\new_[12197]_  | ~\new_[4336]_ ;
  assign n2360 = ~\new_[4030]_  | ~\new_[12067]_ ;
  assign \new_[3621]_  = ~\\u4_u2_buf1_reg[20] ;
  assign \new_[3622]_  = ~\\u4_u2_buf1_reg[27] ;
  assign n2365 = ~\new_[4032]_  | ~\new_[12100]_ ;
  assign \new_[3624]_  = ~\\u4_u2_buf1_reg[24] ;
  assign n2285 = ~\new_[4035]_  | ~phy_rst_pad_o;
  assign \new_[3626]_  = \\u4_u1_dma_out_cnt_reg[4] ;
  assign n2655 = \new_[5990]_  ^ \new_[4274]_ ;
  assign \new_[3628]_  = ~\\u4_u3_buf0_reg[29] ;
  assign \new_[3629]_  = ~\\u4_u2_buf1_reg[17] ;
  assign \new_[3630]_  = ~n2670;
  assign \new_[3631]_  = ~\\u4_u3_buf0_reg[25] ;
  assign \new_[3632]_  = ~\\u1_u3_new_size_reg[3] ;
  assign \new_[3633]_  = ~\\u4_u3_buf0_reg[21] ;
  assign \new_[3634]_  = ~\\u4_u3_buf0_reg[5] ;
  assign n2430 = \new_[4058]_  & \new_[6267]_ ;
  assign \new_[3636]_  = ~\\u4_u1_buf0_reg[5] ;
  assign n2565 = \new_[4176]_  & \new_[6267]_ ;
  assign \new_[3638]_  = \\u4_u1_dma_in_cnt_reg[5] ;
  assign \new_[3639]_  = ~\\u4_u3_buf0_reg[6] ;
  assign n2435 = \new_[4124]_  & \new_[6267]_ ;
  assign n2440 = \new_[4125]_  & \new_[6267]_ ;
  assign n2335 = ~\new_[8494]_  | ~\new_[13165]_  | ~\new_[4204]_ ;
  assign n2445 = ~\new_[4130]_  | ~phy_rst_pad_o;
  assign n2450 = ~\new_[4131]_  | ~\new_[12067]_ ;
  assign n2455 = ~\new_[4132]_  | ~\new_[12067]_ ;
  assign n2460 = ~\new_[4133]_  | ~phy_rst_pad_o;
  assign n2650 = ~\new_[4134]_  | ~phy_rst_pad_o;
  assign n2465 = ~\new_[4135]_  | ~\new_[12067]_ ;
  assign n2470 = ~\new_[4136]_  | ~\new_[12067]_ ;
  assign n2475 = ~\new_[4137]_  | ~phy_rst_pad_o;
  assign n2390 = ~\new_[4138]_  | ~phy_rst_pad_o;
  assign n2480 = ~\new_[4139]_  | ~\new_[12067]_ ;
  assign n2495 = ~\new_[4140]_  | ~\new_[12067]_ ;
  assign n2485 = ~\new_[4141]_  | ~phy_rst_pad_o;
  assign n2490 = ~\new_[4142]_  | ~phy_rst_pad_o;
  assign n2505 = ~\new_[4143]_  | ~phy_rst_pad_o;
  assign n2500 = ~\new_[4144]_  | ~phy_rst_pad_o;
  assign n2385 = ~\new_[4145]_  | ~phy_rst_pad_o;
  assign \new_[3659]_  = ~\\u4_u3_buf0_reg[10] ;
  assign n2510 = ~\new_[4146]_  | ~phy_rst_pad_o;
  assign n2515 = ~\new_[4147]_  | ~phy_rst_pad_o;
  assign n2300 = ~\new_[4149]_  | ~phy_rst_pad_o;
  assign n2520 = ~\new_[4150]_  | ~phy_rst_pad_o;
  assign n2555 = \new_[4174]_  & \new_[6267]_ ;
  assign n2525 = ~\new_[4152]_  | ~phy_rst_pad_o;
  assign n2340 = ~\new_[8496]_  | ~\new_[12158]_  | ~\new_[4205]_ ;
  assign n2530 = ~\new_[4126]_  | ~phy_rst_pad_o;
  assign n2535 = ~\new_[4127]_  | ~phy_rst_pad_o;
  assign n2345 = ~\new_[4156]_  | ~phy_rst_pad_o;
  assign n2310 = ~\new_[8505]_  | ~\new_[12387]_  | ~\new_[4222]_ ;
  assign \new_[3671]_  = \\u4_u2_dma_out_cnt_reg[9] ;
  assign \new_[3672]_  = ~\new_[4062]_  & (~\new_[8306]_  | ~\new_[3479]_ );
  assign n2540 = \new_[4171]_  & \new_[6267]_ ;
  assign n2545 = ~\new_[4172]_  & ~\new_[12849]_ ;
  assign n2550 = \new_[4173]_  & \new_[6267]_ ;
  assign \new_[3676]_  = ~\\u4_u3_buf0_reg[14] ;
  assign \new_[3677]_  = ~\\u4_u3_buf0_reg[13] ;
  assign n2560 = \new_[4175]_  & \new_[6267]_ ;
  assign \new_[3679]_  = ~\\u4_u3_buf0_reg[11] ;
  assign \new_[3680]_  = ~\\u4_u3_buf0_reg[15] ;
  assign \new_[3681]_  = ~\\u4_u3_buf0_reg[4] ;
  assign \new_[3682]_  = ~\\u4_u3_buf0_reg[7] ;
  assign \new_[3683]_  = ~\\u4_u1_buf0_reg[4] ;
  assign \new_[3684]_  = \\u4_u1_dma_out_cnt_reg[8] ;
  assign \wb_data_o[1]  = \\u5_wb_data_o_reg[1] ;
  assign \new_[3686]_  = \\u4_u1_dma_in_cnt_reg[10] ;
  assign \new_[3687]_  = \\u4_u2_dma_out_cnt_reg[11] ;
  assign \new_[3688]_  = \\u4_u1_dma_out_cnt_reg[10] ;
  assign \new_[3689]_  = \\u4_u1_dma_out_cnt_reg[7] ;
  assign \new_[3690]_  = \\u4_u2_dma_in_cnt_reg[7] ;
  assign \new_[3691]_  = \\u4_u1_dma_in_cnt_reg[4] ;
  assign \new_[3692]_  = \\u4_u2_dma_out_cnt_reg[6] ;
  assign \new_[3693]_  = \\u4_u2_dma_in_cnt_reg[6] ;
  assign \new_[3694]_  = ~\\u4_u2_buf1_reg[0] ;
  assign \new_[3695]_  = ~\\u4_u2_buf1_reg[12] ;
  assign \new_[3696]_  = ~\\u4_u2_buf1_reg[16] ;
  assign \new_[3697]_  = ~\\u4_u2_buf1_reg[18] ;
  assign \new_[3698]_  = ~\\u4_u2_buf1_reg[19] ;
  assign \new_[3699]_  = ~\\u4_u2_buf1_reg[1] ;
  assign \new_[3700]_  = ~\\u4_u2_buf1_reg[22] ;
  assign \new_[3701]_  = ~\\u4_u2_buf1_reg[23] ;
  assign \new_[3702]_  = ~\\u4_u2_buf1_reg[21] ;
  assign \new_[3703]_  = ~\\u4_u2_buf1_reg[26] ;
  assign \new_[3704]_  = ~\\u4_u2_buf1_reg[25] ;
  assign \new_[3705]_  = ~\\u4_u2_buf1_reg[29] ;
  assign \new_[3706]_  = ~\\u4_u2_buf1_reg[2] ;
  assign \new_[3707]_  = ~\\u4_u2_buf1_reg[30] ;
  assign \new_[3708]_  = ~\\u4_u2_buf1_reg[8] ;
  assign \new_[3709]_  = ~\\u4_u2_buf1_reg[9] ;
  assign \new_[3710]_  = \\u4_u2_dma_in_cnt_reg[0] ;
  assign \new_[3711]_  = \\u4_u1_dma_in_cnt_reg[2] ;
  assign \new_[3712]_  = \\u4_u1_dma_out_cnt_reg[5] ;
  assign \new_[3713]_  = \\u4_u2_dma_out_cnt_reg[1] ;
  assign \new_[3714]_  = \\u4_u2_dma_out_cnt_reg[2] ;
  assign \new_[3715]_  = \\u4_u2_dma_out_cnt_reg[3] ;
  assign \new_[3716]_  = \\u4_u2_int_stat_reg[0] ;
  assign \new_[3717]_  = ~\\u4_u3_buf0_reg[0] ;
  assign \new_[3718]_  = \\u4_u2_dma_out_cnt_reg[0] ;
  assign \new_[3719]_  = ~\\u4_u3_buf0_reg[16] ;
  assign \new_[3720]_  = ~\\u4_u3_buf0_reg[17] ;
  assign \new_[3721]_  = ~\\u4_u3_buf0_reg[18] ;
  assign \new_[3722]_  = ~\\u4_u3_buf0_reg[19] ;
  assign \new_[3723]_  = ~\\u4_u3_buf0_reg[1] ;
  assign \new_[3724]_  = ~\\u4_u3_buf0_reg[20] ;
  assign \new_[3725]_  = ~\\u4_u3_buf0_reg[12] ;
  assign \new_[3726]_  = ~\\u4_u3_buf0_reg[23] ;
  assign \new_[3727]_  = ~\\u4_u3_buf0_reg[24] ;
  assign \new_[3728]_  = ~\\u4_u3_buf0_reg[22] ;
  assign \new_[3729]_  = ~\\u4_u3_buf0_reg[27] ;
  assign \new_[3730]_  = ~\\u4_u3_buf0_reg[26] ;
  assign \new_[3731]_  = ~\\u4_u3_buf0_reg[2] ;
  assign \new_[3732]_  = ~\\u4_u3_buf0_reg[30] ;
  assign \new_[3733]_  = ~\\u4_u3_buf0_reg[3] ;
  assign \new_[3734]_  = ~\\u4_u3_buf0_reg[8] ;
  assign \new_[3735]_  = ~\\u4_u3_buf0_reg[9] ;
  assign \new_[3736]_  = ~\\u4_u1_buf0_reg[0] ;
  assign \new_[3737]_  = ~\\u4_u1_buf0_reg[12] ;
  assign \new_[3738]_  = ~\\u4_u1_buf0_reg[17] ;
  assign \new_[3739]_  = \\u4_u0_int_stat_reg[0] ;
  assign \new_[3740]_  = ~\\u4_u1_buf0_reg[29] ;
  assign \new_[3741]_  = \\u4_u1_int_stat_reg[0] ;
  assign \new_[3742]_  = ~\new_[5918]_  & (~\new_[4309]_  | ~\new_[5916]_ );
  assign \new_[3743]_  = ~\new_[5921]_  & (~\new_[4310]_  | ~\new_[5919]_ );
  assign \new_[3744]_  = ~\new_[5927]_  & (~\new_[4311]_  | ~\new_[5925]_ );
  assign n2320 = ~\new_[8129]_  | ~\new_[12244]_  | ~\new_[4261]_ ;
  assign n2570 = ~\new_[8130]_  | ~\new_[13165]_  | ~\new_[4207]_ ;
  assign n2575 = ~\new_[8497]_  | ~\new_[13165]_  | ~\new_[4208]_ ;
  assign n2580 = ~\new_[8009]_  | ~\new_[13165]_  | ~\new_[4209]_ ;
  assign n2585 = ~\new_[8498]_  | ~\new_[12387]_  | ~\new_[4210]_ ;
  assign n2590 = ~\new_[8016]_  | ~\new_[12387]_  | ~\new_[4211]_ ;
  assign n2595 = ~\new_[8540]_  | ~\new_[13165]_  | ~\new_[4212]_ ;
  assign n2600 = ~\new_[8481]_  | ~\new_[12158]_  | ~\new_[4213]_ ;
  assign n2605 = ~\new_[8466]_  | ~\new_[12387]_  | ~\new_[4214]_ ;
  assign n2610 = ~\new_[8463]_  | ~\new_[12491]_  | ~\new_[4215]_ ;
  assign n2660 = ~\new_[8132]_  | ~\new_[12491]_  | ~\new_[4216]_ ;
  assign n2615 = ~\new_[8500]_  | ~\new_[12491]_  | ~\new_[4217]_ ;
  assign n2620 = ~\new_[8512]_  | ~\new_[12244]_  | ~\new_[4218]_ ;
  assign n2625 = ~\new_[8503]_  | ~\new_[12491]_  | ~\new_[4219]_ ;
  assign n2280 = ~\new_[8508]_  | ~\new_[12158]_  | ~\new_[4220]_ ;
  assign n2630 = ~\new_[8510]_  | ~\new_[12244]_  | ~\new_[4221]_ ;
  assign n2635 = ~\new_[8557]_  | ~\new_[12197]_  | ~\new_[4224]_ ;
  assign n2640 = ~\new_[8546]_  | ~\new_[12197]_  | ~\new_[4225]_ ;
  assign \new_[3763]_  = \new_[4148]_  | \new_[2611]_ ;
  assign \new_[3764]_  = ~\new_[4163]_  | ~\new_[4007]_ ;
  assign \new_[3765]_  = ~\new_[4164]_  | ~\new_[5080]_ ;
  assign n2295 = \new_[4165]_  & \new_[6256]_ ;
  assign n2395 = \new_[4166]_  & \new_[6267]_ ;
  assign n2400 = \new_[4167]_  & \new_[6276]_ ;
  assign n2290 = \new_[4168]_  & \new_[6288]_ ;
  assign n2350 = ~\new_[4017]_  | ~\new_[12067]_ ;
  assign n2305 = \new_[4246]_  ^ \new_[4459]_ ;
  assign n2370 = ~\new_[4184]_  | ~\new_[12100]_ ;
  assign n2380 = ~\new_[3961]_  | ~phy_rst_pad_o;
  assign n2375 = ~\new_[3962]_  | ~phy_rst_pad_o;
  assign \new_[3775]_  = ~\new_[14463]_  | ~\new_[14494]_ ;
  assign \new_[3776]_  = ~\new_[4008]_  | ~\new_[5099]_ ;
  assign \new_[3777]_  = \\u4_u1_dma_in_cnt_reg[1] ;
  assign n2645 = ~\new_[3934]_ ;
  assign n2325 = ~\new_[8432]_  | ~\new_[12244]_  | ~\new_[4312]_ ;
  assign n2330 = ~\new_[4063]_  | ~phy_rst_pad_o;
  assign \new_[3781]_  = \\u5_state_reg[0] ;
  assign \new_[3782]_  = \\u1_u3_new_size_reg[4] ;
  assign n2410 = ~\new_[3978]_  & ~\new_[13296]_ ;
  assign n2405 = \new_[3979]_  & \new_[6267]_ ;
  assign n2415 = \new_[3980]_  & \new_[6267]_ ;
  assign n2420 = \new_[3982]_  & \new_[6267]_ ;
  assign \new_[3787]_  = \\u4_u2_dma_in_cnt_reg[11] ;
  assign \new_[3788]_  = \\u4_u1_dma_in_cnt_reg[3] ;
  assign n2425 = ~\new_[4248]_  | ~\new_[4020]_  | ~\new_[4464]_ ;
  assign \new_[3790]_  = \\u4_u2_dma_in_cnt_reg[8] ;
  assign \new_[3791]_  = ~\\u4_u3_buf1_reg[7] ;
  assign n2690 = ~\new_[8351]_  | ~\new_[12158]_  | ~\new_[4381]_ ;
  assign n2760 = ~\new_[8539]_  | ~\new_[12387]_  | ~\new_[4598]_ ;
  assign \new_[3794]_  = u1_u3_pid_seq_err_reg;
  assign n2790 = ~\new_[8364]_  | ~\new_[12197]_  | ~\new_[4521]_ ;
  assign n2735 = ~\new_[8365]_  | ~\new_[12197]_  | ~\new_[4522]_ ;
  assign \new_[3797]_  = ~\new_[6629]_  & (~\new_[4478]_  | ~\new_[6469]_ );
  assign \new_[3798]_  = ~\new_[4242]_  | ~\new_[7654]_ ;
  assign \new_[3799]_  = ~\\u4_u2_buf0_reg[2] ;
  assign \new_[3800]_  = ~\new_[4275]_  | ~\new_[9380]_ ;
  assign \new_[3801]_  = ~\new_[4276]_  | ~\new_[8877]_ ;
  assign \new_[3802]_  = ~\new_[14528]_  & ~\new_[14527]_ ;
  assign \new_[3803]_  = \new_[14470]_  & \new_[14494]_ ;
  assign \new_[3804]_  = ~\new_[4259]_  & ~\new_[4260]_ ;
  assign \new_[3805]_  = ~\new_[4007]_ ;
  assign \new_[3806]_  = \\u4_u2_dma_out_cnt_reg[4] ;
  assign \new_[3807]_  = ~\\u4_u3_buf1_reg[5] ;
  assign \new_[3808]_  = ~\\u4_u2_buf0_reg[26] ;
  assign n2795 = ~\new_[8555]_  | ~\new_[12216]_  | ~\new_[4551]_ ;
  assign n2800 = ~\new_[4271]_  | ~\new_[12067]_ ;
  assign n2670 = u5_wb_ack_s1_reg;
  assign n3040 = \new_[4360]_  & \new_[6267]_ ;
  assign n3160 = ~\new_[4272]_  | ~phy_rst_pad_o;
  assign n2805 = ~\new_[4273]_  | ~\new_[12058]_ ;
  assign \new_[3815]_  = \\u4_u2_dma_out_cnt_reg[7] ;
  assign \new_[3816]_  = ~\\u4_u2_buf0_reg[4] ;
  assign n2915 = \new_[4278]_  & \new_[6276]_ ;
  assign \new_[3818]_  = ~\new_[4254]_  & (~\new_[9135]_  | ~\wb_data_i[13] );
  assign n2910 = \new_[4279]_  & \new_[6267]_ ;
  assign n2905 = \new_[4280]_  & \new_[6267]_ ;
  assign n2900 = \new_[4281]_  & \new_[6267]_ ;
  assign \new_[3822]_  = ~\new_[6606]_  & (~\new_[4491]_  | ~\new_[4615]_ );
  assign n3055 = \new_[4355]_  & \new_[6276]_ ;
  assign \new_[3824]_  = ~\\u4_u3_buf1_reg[6] ;
  assign n2925 = \new_[4300]_  & \new_[6276]_ ;
  assign n2930 = \new_[4301]_  & \new_[6276]_ ;
  assign n2920 = \new_[4302]_  & \new_[6267]_ ;
  assign n2710 = \new_[4313]_  & \new_[6267]_ ;
  assign \new_[3829]_  = ~\new_[4340]_  & (~\new_[9135]_  | ~\wb_data_i[11] );
  assign \new_[3830]_  = ~\new_[4339]_  & (~\new_[9135]_  | ~\wb_data_i[15] );
  assign \new_[3831]_  = ~\new_[4341]_  & (~\new_[9135]_  | ~\wb_data_i[6] );
  assign \new_[3832]_  = \\u5_state_reg[5] ;
  assign n2935 = ~\new_[4314]_  | ~phy_rst_pad_o;
  assign n2940 = ~\new_[4315]_  | ~phy_rst_pad_o;
  assign n2945 = ~\new_[4316]_  | ~phy_rst_pad_o;
  assign n2950 = ~\new_[4317]_  | ~phy_rst_pad_o;
  assign n2955 = ~\new_[4318]_  | ~phy_rst_pad_o;
  assign n2960 = ~\new_[4319]_  | ~phy_rst_pad_o;
  assign n2700 = ~\new_[4320]_  | ~phy_rst_pad_o;
  assign n2965 = ~\new_[4321]_  | ~phy_rst_pad_o;
  assign n2970 = ~\new_[4322]_  | ~phy_rst_pad_o;
  assign n2975 = ~\new_[4323]_  | ~phy_rst_pad_o;
  assign n2730 = ~\new_[4324]_  | ~phy_rst_pad_o;
  assign n2980 = ~\new_[4325]_  | ~phy_rst_pad_o;
  assign n2985 = ~\new_[4326]_  | ~phy_rst_pad_o;
  assign n2990 = ~\new_[4327]_  | ~\new_[13165]_ ;
  assign n2725 = ~\new_[4328]_  | ~\new_[13165]_ ;
  assign n3005 = ~\new_[4329]_  | ~phy_rst_pad_o;
  assign n2995 = ~\new_[4330]_  | ~\new_[13165]_ ;
  assign n3000 = ~\new_[4331]_  | ~\new_[13165]_ ;
  assign n3010 = ~\new_[4332]_  | ~phy_rst_pad_o;
  assign n3015 = ~\new_[4333]_  | ~phy_rst_pad_o;
  assign n2715 = ~\new_[4334]_  | ~phy_rst_pad_o;
  assign n3020 = ~\new_[4305]_  | ~\new_[12067]_ ;
  assign n3025 = ~\new_[4306]_  | ~phy_rst_pad_o;
  assign n2750 = ~\new_[8439]_  | ~\new_[12158]_  | ~\new_[4412]_ ;
  assign n2775 = ~\new_[8472]_  | ~\new_[12442]_  | ~\new_[4414]_ ;
  assign n2780 = ~\new_[4338]_  | ~phy_rst_pad_o;
  assign \new_[3859]_  = ~\new_[4282]_  & (~\new_[9055]_  | ~\new_[3690]_ );
  assign \new_[3860]_  = ~\new_[4283]_  & (~\new_[8691]_  | ~\new_[3315]_ );
  assign n2745 = ~\new_[8548]_  | ~\new_[12244]_  | ~\new_[4415]_ ;
  assign \new_[3862]_  = ~\new_[4335]_  & (~\new_[9135]_  | ~\wb_data_i[14] );
  assign n3030 = \new_[4354]_  & \new_[6276]_ ;
  assign \new_[3864]_  = ~\\u4_u3_buf1_reg[14] ;
  assign \new_[3865]_  = ~\\u4_u3_buf1_reg[10] ;
  assign \new_[3866]_  = ~\\u4_u3_buf1_reg[13] ;
  assign \new_[3867]_  = ~\\u4_u3_buf1_reg[11] ;
  assign \new_[3868]_  = ~\\u4_u3_buf1_reg[15] ;
  assign \new_[3869]_  = ~\\u4_u2_buf0_reg[5] ;
  assign \new_[3870]_  = ~\\u4_u3_buf1_reg[4] ;
  assign n3060 = \new_[4356]_  & \new_[6276]_ ;
  assign n3065 = \new_[4357]_  & \new_[6276]_ ;
  assign n3070 = \new_[4358]_  & \new_[6276]_ ;
  assign n3045 = \new_[4361]_  & \new_[6267]_ ;
  assign \new_[3875]_  = \\u4_u2_dma_out_cnt_reg[8] ;
  assign \wb_data_o[3]  = \\u5_wb_data_o_reg[3] ;
  assign n3050 = \new_[4362]_  & \new_[6267]_ ;
  assign \new_[3878]_  = \\u4_int_srcb_reg[0] ;
  assign \new_[3879]_  = \\u4_u2_dma_in_cnt_reg[10] ;
  assign \new_[3880]_  = u2_wack_r_reg;
  assign \new_[3881]_  = \\u1_u0_state_reg[3] ;
  assign \new_[3882]_  = \\u4_u2_dma_in_cnt_reg[5] ;
  assign \new_[3883]_  = \\u4_u2_dma_out_cnt_reg[10] ;
  assign \new_[3884]_  = \\u4_u2_dma_in_cnt_reg[4] ;
  assign n3035 = \new_[4366]_  & \new_[6267]_ ;
  assign \new_[3886]_  = ~\\u4_u3_buf1_reg[28] ;
  assign \new_[3887]_  = ~\\u4_u3_buf1_reg[31] ;
  assign \new_[3888]_  = \\u4_u2_dma_in_cnt_reg[2] ;
  assign \new_[3889]_  = \\u4_u2_dma_in_cnt_reg[3] ;
  assign \new_[3890]_  = \\u4_u2_dma_out_cnt_reg[5] ;
  assign \new_[3891]_  = ~\\u4_u2_buf0_reg[21] ;
  assign \new_[3892]_  = ~\\u4_u2_buf0_reg[23] ;
  assign \new_[3893]_  = ~\\u4_u2_buf0_reg[27] ;
  assign \new_[3894]_  = ~\\u4_u2_buf0_reg[9] ;
  assign \new_[3895]_  = \\u1_u2_state_reg[2] ;
  assign n3075 = ~\new_[8554]_  | ~\new_[13165]_  | ~\new_[4375]_ ;
  assign n2685 = ~\new_[8462]_  | ~\new_[12491]_  | ~\new_[4376]_ ;
  assign n3080 = ~\new_[8340]_  | ~\new_[12197]_  | ~\new_[4378]_ ;
  assign n3085 = ~\new_[8344]_  | ~\new_[12197]_  | ~\new_[4379]_ ;
  assign n3090 = ~\new_[8345]_  | ~\new_[12258]_  | ~\new_[4380]_ ;
  assign n3095 = ~\new_[8359]_  | ~\new_[13165]_  | ~\new_[4382]_ ;
  assign n2675 = ~\new_[8360]_  | ~\new_[12252]_  | ~\new_[4383]_ ;
  assign n3100 = ~\new_[8535]_  | ~\new_[12442]_  | ~\new_[4395]_ ;
  assign n2695 = ~\new_[8537]_  | ~\new_[12442]_  | ~\new_[4396]_ ;
  assign n3105 = ~\new_[8471]_  | ~\new_[12197]_  | ~\new_[4397]_ ;
  assign n3110 = ~\new_[8465]_  | ~\new_[12244]_  | ~\new_[4398]_ ;
  assign n2755 = ~\new_[8536]_  | ~\new_[12244]_  | ~\new_[4487]_ ;
  assign n3115 = ~\new_[8532]_  | ~\new_[12244]_  | ~\new_[4399]_ ;
  assign n2720 = ~\new_[8541]_  | ~\new_[12197]_  | ~\new_[4400]_ ;
  assign n3145 = ~\new_[8542]_  | ~\new_[12244]_  | ~\new_[4393]_ ;
  assign n3120 = ~\new_[8511]_  | ~\new_[12244]_  | ~\new_[4401]_ ;
  assign n3125 = ~\new_[8531]_  | ~\new_[13162]_  | ~\new_[4389]_ ;
  assign n3130 = ~\new_[8543]_  | ~\new_[13165]_  | ~\new_[4402]_ ;
  assign n3135 = ~\new_[8457]_  | ~\new_[13165]_  | ~\new_[4403]_ ;
  assign n3140 = ~\new_[8544]_  | ~\new_[12197]_  | ~\new_[4404]_ ;
  assign n3150 = ~\new_[8428]_  | ~\new_[12486]_  | ~\new_[4405]_ ;
  assign n3155 = ~\new_[8556]_  | ~\new_[12197]_  | ~\new_[4394]_ ;
  assign n2680 = ~\new_[8553]_  | ~\new_[12197]_  | ~\new_[4406]_ ;
  assign n2825 = ~\new_[7456]_  & ~\new_[4190]_ ;
  assign \new_[3920]_  = ~\new_[4345]_  & (~\new_[9135]_  | ~\wb_data_i[28] );
  assign \new_[3921]_  = ~\new_[4346]_  & (~\new_[9135]_  | ~\wb_data_i[31] );
  assign n2785 = ~\new_[4243]_  | ~\new_[13165]_ ;
  assign \wb_data_o[0]  = \\u5_wb_data_o_reg[0] ;
  assign \new_[3924]_  = ~\new_[4238]_  & (~\new_[9135]_  | ~\wb_data_i[10] );
  assign n2815 = ~\new_[4186]_  | ~\new_[12100]_ ;
  assign n2820 = ~\new_[4188]_  | ~phy_rst_pad_o;
  assign n2810 = ~\new_[4187]_  | ~phy_rst_pad_o;
  assign n2830 = \new_[4185]_  & \new_[6267]_ ;
  assign \new_[3929]_  = ~\new_[4230]_  & ~\new_[14528]_ ;
  assign \new_[3930]_  = \\u4_u2_dma_in_cnt_reg[1] ;
  assign n2705 = \new_[4189]_  & \new_[6267]_ ;
  assign \new_[3932]_  = \\u4_u3_dma_out_cnt_reg[9] ;
  assign n2835 = ~\new_[8260]_  & ~\new_[4190]_ ;
  assign \new_[3934]_  = ~\new_[10046]_  | ~\new_[10486]_  | ~\new_[10070]_  | ~\new_[4374]_ ;
  assign \new_[3935]_  = ~\new_[4164]_ ;
  assign \new_[3936]_  = ~\new_[4458]_  | ~\new_[4233]_ ;
  assign \new_[3937]_  = ~\new_[8795]_  | ~\new_[4746]_  | ~\new_[6027]_  | ~\new_[10372]_ ;
  assign \new_[3938]_  = \\u4_u3_dma_in_cnt_reg[10] ;
  assign n2840 = \new_[4199]_  & \new_[6276]_ ;
  assign \new_[3940]_  = \\u4_u3_dma_in_cnt_reg[11] ;
  assign n2855 = \new_[4202]_  & \new_[6276]_ ;
  assign n2860 = \new_[4203]_  & \new_[6276]_ ;
  assign n2850 = \new_[4227]_  & \new_[6267]_ ;
  assign \new_[3944]_  = ~\new_[4191]_  | ~\new_[13315]_ ;
  assign n2845 = ~\new_[12046]_  & ~\new_[4190]_ ;
  assign n2765 = ~\new_[8538]_  | ~\new_[12244]_  | ~\new_[4546]_ ;
  assign n2770 = ~\new_[4284]_  | ~phy_rst_pad_o;
  assign n2865 = ~\new_[8945]_  & ~\new_[4190]_ ;
  assign n2870 = ~\new_[11455]_  & ~\new_[4190]_ ;
  assign n2665 = ~\new_[10672]_  & ~\new_[4190]_ ;
  assign n2875 = ~\new_[9878]_  & ~\new_[4190]_ ;
  assign \wb_data_o[2]  = \\u5_wb_data_o_reg[2] ;
  assign n2880 = ~\new_[9379]_  & ~\new_[4190]_ ;
  assign n2885 = ~\new_[9977]_  & ~\new_[4190]_ ;
  assign n2740 = ~\new_[9365]_  & ~\new_[4190]_ ;
  assign n2895 = ~\new_[8689]_  & ~\new_[4190]_ ;
  assign n2890 = ~\new_[9123]_  & ~\new_[4190]_ ;
  assign \new_[3958]_  = ~\new_[4251]_  & (~\new_[9135]_  | ~\wb_data_i[4] );
  assign \new_[3959]_  = ~\new_[4252]_  & (~\new_[9135]_  | ~\wb_data_i[5] );
  assign \new_[3960]_  = ~\new_[4253]_  & (~\new_[9135]_  | ~\wb_data_i[7] );
  assign \new_[3961]_  = ~\new_[4423]_  & (~\new_[9141]_  | ~\wb_data_i[5] );
  assign \new_[3962]_  = ~\new_[4424]_  & (~\new_[9141]_  | ~\wb_data_i[7] );
  assign n3435 = \new_[4592]_  & \new_[6276]_ ;
  assign n3285 = ~\new_[8433]_  | ~\new_[12244]_  | ~\new_[4866]_ ;
  assign n3235 = ~\new_[8478]_  | ~\new_[12244]_  | ~\new_[4867]_ ;
  assign n3290 = ~\new_[8437]_  | ~\new_[12197]_  | ~\new_[4868]_ ;
  assign \new_[3967]_  = ~\new_[4191]_ ;
  assign \new_[3968]_  = ~\\u4_u3_buf1_reg[25] ;
  assign n3490 = ~\new_[8550]_  | ~\new_[12244]_  | ~\new_[4629]_ ;
  assign \new_[3970]_  = ~\new_[4492]_  | ~\new_[8877]_ ;
  assign \new_[3971]_  = ~\new_[4494]_  | ~\new_[9380]_ ;
  assign \new_[3972]_  = (~\new_[4654]_  | ~\new_[7449]_ ) & (~\new_[5191]_  | ~\new_[5355]_ );
  assign n3595 = ~\new_[5156]_  | ~\new_[8916]_  | ~rst_i | ~\new_[11781]_ ;
  assign \new_[3974]_  = ~\\u4_u3_buf1_reg[21] ;
  assign \new_[3975]_  = ~\new_[4499]_  | ~\new_[8877]_ ;
  assign n3505 = ~\new_[8485]_  | ~\new_[12197]_  | ~\new_[4624]_ ;
  assign \new_[3977]_  = ~\new_[5191]_  & (~\new_[4718]_  | ~\new_[5419]_ );
  assign \new_[3978]_  = ~\new_[4418]_  & (~\new_[7542]_  | ~\new_[9021]_ );
  assign \new_[3979]_  = ~\new_[4460]_  | (~\new_[7694]_  & ~\new_[12650]_ );
  assign \new_[3980]_  = ~\new_[4516]_  | (~\new_[8678]_  & ~\new_[12650]_ );
  assign \new_[3981]_  = ~\new_[4463]_  | ~\new_[9380]_ ;
  assign \new_[3982]_  = ~\new_[4420]_  | (~\new_[9962]_  & ~\new_[12650]_ );
  assign \new_[3983]_  = ~\new_[4465]_  | ~\new_[8876]_ ;
  assign \new_[3984]_  = ~\new_[4466]_  | ~\new_[8876]_ ;
  assign \new_[3985]_  = ~\new_[4467]_  | ~\new_[8877]_ ;
  assign \new_[3986]_  = ~\new_[4468]_  | ~\new_[8877]_ ;
  assign \new_[3987]_  = ~\new_[4469]_  | ~\new_[8877]_ ;
  assign \new_[3988]_  = ~\new_[4470]_  | ~\new_[8878]_ ;
  assign \new_[3989]_  = ~\new_[4471]_  | ~\new_[8876]_ ;
  assign \new_[3990]_  = ~\new_[4472]_  | ~\new_[8876]_ ;
  assign \new_[3991]_  = ~\new_[4473]_  | ~\new_[9380]_ ;
  assign \new_[3992]_  = ~\new_[4474]_  | ~\new_[9380]_ ;
  assign \new_[3993]_  = ~\new_[4475]_  | ~\new_[8876]_ ;
  assign \new_[3994]_  = ~\new_[4476]_  | ~\new_[8877]_ ;
  assign \new_[3995]_  = ~\new_[4477]_  | ~\new_[8874]_ ;
  assign \new_[3996]_  = ~\new_[4479]_  | ~\new_[9380]_ ;
  assign \new_[3997]_  = \\u4_u3_dma_out_cnt_reg[3] ;
  assign \new_[3998]_  = ~\\u4_u3_buf1_reg[0] ;
  assign n3295 = ~\new_[8504]_  | ~\new_[12339]_  | ~\new_[4879]_ ;
  assign \new_[4000]_  = ~\new_[4482]_  | ~\new_[9138]_ ;
  assign \new_[4001]_  = ~\new_[4483]_  | ~\new_[9138]_ ;
  assign n3240 = ~\new_[8482]_  | ~\new_[13165]_  | ~\new_[4880]_ ;
  assign \new_[4003]_  = ~\\u4_u3_buf1_reg[18] ;
  assign n3610 = \new_[4594]_  & \new_[6276]_ ;
  assign n3440 = \new_[4595]_  & \new_[6276]_ ;
  assign \new_[4006]_  = ~\new_[4229]_ ;
  assign \new_[4007]_  = ~\new_[5083]_  & (~\new_[5082]_  | ~\new_[4750]_ );
  assign \new_[4008]_  = ~\new_[4231]_ ;
  assign n3600 = \new_[6708]_  ^ \new_[4718]_ ;
  assign n3255 = ~\new_[8455]_  | ~\new_[12491]_  | ~\new_[4693]_ ;
  assign \new_[4011]_  = u1_u3_buf1_st_max_reg;
  assign n3495 = ~\new_[8528]_  | ~\new_[12252]_  | ~\new_[4630]_ ;
  assign \new_[4013]_  = ~\\u1_u3_new_size_reg[2] ;
  assign n3330 = \new_[4481]_  & \new_[6288]_ ;
  assign n3325 = \new_[4484]_  & \new_[6276]_ ;
  assign n3320 = \new_[4485]_  & \new_[6276]_ ;
  assign \new_[4017]_  = ~\new_[4425]_  & (~\new_[9141]_  | ~\wb_data_i[13] );
  assign n3245 = \new_[4486]_  & \new_[6276]_ ;
  assign n3480 = ~\new_[8435]_  | ~\new_[12244]_  | ~\new_[4627]_ ;
  assign \new_[4020]_  = ~\new_[4428]_  & (~\new_[7482]_  | ~\new_[5078]_ );
  assign n3275 = ~\new_[8421]_  | ~\new_[12197]_  | ~\new_[4610]_ ;
  assign n3280 = ~\new_[8424]_  | ~\new_[12486]_  | ~\new_[4611]_ ;
  assign n3250 = ~\new_[8456]_  | ~\new_[12486]_  | ~\new_[4614]_ ;
  assign \new_[4024]_  = ~\new_[4555]_  | ~\new_[8877]_ ;
  assign n3345 = \new_[4518]_  & \new_[6288]_ ;
  assign n3340 = \new_[4519]_  & \new_[6288]_ ;
  assign n3335 = \new_[4520]_  & \new_[6276]_ ;
  assign n3205 = \new_[4523]_  & \new_[6276]_ ;
  assign \new_[4029]_  = ~\new_[4891]_  & (~\new_[5420]_  | ~\new_[4894]_ );
  assign \new_[4030]_  = ~\new_[4547]_  & (~\new_[9141]_  | ~\wb_data_i[11] );
  assign \new_[4031]_  = ~\new_[14528]_ ;
  assign \new_[4032]_  = ~\new_[4548]_  & (~\new_[9141]_  | ~\wb_data_i[15] );
  assign \new_[4033]_  = ~\new_[5086]_  & ~\new_[4764]_ ;
  assign \new_[4034]_  = \new_[5092]_  | \new_[5091]_ ;
  assign \new_[4035]_  = ~\new_[4549]_  & (~\new_[9141]_  | ~\wb_data_i[6] );
  assign n3350 = ~\new_[4525]_  | ~phy_rst_pad_o;
  assign n3355 = ~\new_[4526]_  | ~\new_[12100]_ ;
  assign n3360 = ~\new_[4527]_  | ~phy_rst_pad_o;
  assign n3215 = ~\new_[4528]_  | ~phy_rst_pad_o;
  assign n3365 = ~\new_[4529]_  | ~phy_rst_pad_o;
  assign n3370 = ~\new_[4530]_  | ~\new_[12067]_ ;
  assign n3375 = ~\new_[4531]_  | ~\new_[12067]_ ;
  assign n3190 = ~\new_[4532]_  | ~\new_[12100]_ ;
  assign n3390 = ~\new_[4533]_  | ~\new_[12100]_ ;
  assign n3380 = ~\new_[4534]_  | ~phy_rst_pad_o;
  assign n3385 = ~\new_[4535]_  | ~phy_rst_pad_o;
  assign n3200 = ~\new_[4536]_  | ~phy_rst_pad_o;
  assign n3400 = ~\new_[4537]_  | ~phy_rst_pad_o;
  assign n3395 = ~\new_[4538]_  | ~phy_rst_pad_o;
  assign n3195 = ~\new_[4539]_  | ~phy_rst_pad_o;
  assign n3405 = ~\new_[4540]_  | ~\new_[12067]_ ;
  assign n3410 = ~\new_[4541]_  | ~phy_rst_pad_o;
  assign n3415 = ~\new_[4542]_  | ~\new_[12067]_ ;
  assign n3185 = ~\new_[4543]_  | ~\new_[12067]_ ;
  assign n3420 = ~\new_[4544]_  | ~phy_rst_pad_o;
  assign n3425 = ~\new_[4545]_  | ~phy_rst_pad_o;
  assign \new_[4057]_  = ~\new_[5720]_  & (~\new_[4890]_  | ~\new_[6222]_ );
  assign \new_[4058]_  = ~\new_[4580]_  | (~\new_[9164]_  & ~\new_[12650]_ );
  assign \new_[4059]_  = ~\new_[5029]_  | ~\new_[6222]_  | ~\new_[5575]_  | ~\new_[5981]_ ;
  assign \new_[4060]_  = ~\new_[4489]_  & (~\new_[9054]_  | ~\new_[4070]_ );
  assign n3225 = \new_[5987]_  ^ \new_[4894]_ ;
  assign \new_[4062]_  = ~\new_[5582]_  | ~\new_[5184]_  | ~\new_[5607]_  | ~\new_[6905]_ ;
  assign \new_[4063]_  = ~\new_[4524]_  & (~\new_[9141]_  | ~\wb_data_i[14] );
  assign n3430 = \new_[4587]_  & \new_[6288]_ ;
  assign n3470 = \new_[4588]_  & \new_[6288]_ ;
  assign n3445 = \new_[4589]_  & \new_[6288]_ ;
  assign n3450 = \new_[4590]_  & \new_[6288]_ ;
  assign n3455 = \new_[4591]_  & \new_[6288]_ ;
  assign \new_[4069]_  = \\u4_u3_dma_out_cnt_reg[11] ;
  assign \new_[4070]_  = \\u4_u3_dma_in_cnt_reg[7] ;
  assign \new_[4071]_  = ~u4_u0_r1_reg;
  assign \new_[4072]_  = \\u5_state_reg[4] ;
  assign \new_[4073]_  = \\u4_u3_dma_in_cnt_reg[6] ;
  assign \new_[4074]_  = \\u4_u3_dma_out_cnt_reg[6] ;
  assign \new_[4075]_  = ~\\u4_u3_buf1_reg[12] ;
  assign \new_[4076]_  = ~\\u4_u3_buf1_reg[16] ;
  assign \new_[4077]_  = ~\\u4_u3_buf1_reg[17] ;
  assign \new_[4078]_  = ~\\u4_u3_buf1_reg[19] ;
  assign \new_[4079]_  = ~\\u4_u3_buf1_reg[1] ;
  assign \new_[4080]_  = ~\\u4_u3_buf1_reg[20] ;
  assign \new_[4081]_  = ~\\u4_u3_buf1_reg[22] ;
  assign \new_[4082]_  = ~\\u4_u3_buf1_reg[23] ;
  assign \new_[4083]_  = ~\\u4_u3_buf1_reg[24] ;
  assign n3590 = \new_[4596]_  & \new_[6276]_ ;
  assign \new_[4085]_  = ~\\u4_u3_buf1_reg[27] ;
  assign \new_[4086]_  = ~\\u4_u3_buf1_reg[26] ;
  assign \new_[4087]_  = ~\\u4_u3_buf1_reg[30] ;
  assign \new_[4088]_  = ~\\u4_u3_buf1_reg[2] ;
  assign \new_[4089]_  = ~\\u4_u3_buf1_reg[9] ;
  assign \new_[4090]_  = ~\\u4_u3_buf1_reg[8] ;
  assign \new_[4091]_  = \\u1_u0_state_reg[0] ;
  assign \new_[4092]_  = \\u1_u0_state_reg[1] ;
  assign n3460 = ~\new_[4582]_  & ~\new_[7411]_ ;
  assign n3465 = ~\new_[8427]_  | ~\new_[12197]_  | ~\new_[4652]_ ;
  assign \new_[4095]_  = \\u4_u3_dma_in_cnt_reg[0] ;
  assign \new_[4096]_  = \\u4_u3_dma_out_cnt_reg[1] ;
  assign \new_[4097]_  = \\u4_u3_dma_out_cnt_reg[2] ;
  assign \new_[4098]_  = \\u4_u3_dma_out_cnt_reg[0] ;
  assign n3475 = ~\new_[8425]_  | ~\new_[12244]_  | ~\new_[4625]_ ;
  assign n3485 = ~\new_[8426]_  | ~\new_[12244]_  | ~\new_[4628]_ ;
  assign n3500 = ~\new_[8420]_  | ~\new_[12252]_  | ~\new_[4631]_ ;
  assign n3230 = ~\new_[8477]_  | ~\new_[12339]_  | ~\new_[4632]_ ;
  assign n3520 = ~\new_[8458]_  | ~\new_[12067]_  | ~\new_[4633]_ ;
  assign n3510 = ~\new_[8419]_  | ~\new_[12491]_  | ~\new_[4634]_ ;
  assign n3515 = ~\new_[8474]_  | ~\new_[12491]_  | ~\new_[4635]_ ;
  assign n3220 = ~\new_[8475]_  | ~\new_[12486]_  | ~\new_[4636]_ ;
  assign n3530 = ~\new_[8492]_  | ~\new_[12486]_  | ~\new_[4637]_ ;
  assign n3525 = ~\new_[8429]_  | ~\new_[13165]_  | ~\new_[4639]_ ;
  assign n3210 = ~\new_[8430]_  | ~\new_[12486]_  | ~\new_[4640]_ ;
  assign n3535 = ~\new_[8431]_  | ~\new_[12486]_  | ~\new_[4642]_ ;
  assign n3540 = ~\new_[8488]_  | ~\new_[12491]_  | ~\new_[4644]_ ;
  assign n3545 = ~\new_[8491]_  | ~\new_[12197]_  | ~\new_[4645]_ ;
  assign n3550 = ~\new_[8530]_  | ~\new_[12197]_  | ~\new_[4646]_ ;
  assign n3555 = ~\new_[8434]_  | ~\new_[12258]_  | ~\new_[4647]_ ;
  assign n3175 = ~\new_[4583]_  & ~\new_[8124]_ ;
  assign n3575 = ~\new_[4584]_  & ~\new_[7414]_ ;
  assign n3565 = ~\new_[8495]_  | ~\new_[13165]_  | ~\new_[4656]_ ;
  assign n3560 = ~\new_[8493]_  | ~\new_[13165]_  | ~\new_[4655]_ ;
  assign n3570 = ~\new_[8131]_  | ~\new_[13165]_  | ~\new_[4657]_ ;
  assign n3180 = ~\new_[8489]_  | ~\new_[12158]_  | ~\new_[4658]_ ;
  assign n3580 = ~\new_[8188]_  | ~\new_[12491]_  | ~\new_[4659]_ ;
  assign n3170 = ~\new_[8502]_  | ~\new_[12244]_  | ~\new_[4660]_ ;
  assign n3585 = ~\new_[4585]_  & ~\new_[7418]_ ;
  assign \new_[4124]_  = ~\new_[4579]_  | (~\new_[9676]_  & ~\new_[12650]_ );
  assign \new_[4125]_  = ~\new_[4581]_  | (~\new_[10688]_  & ~\new_[12650]_ );
  assign \new_[4126]_  = ~\new_[4556]_  & (~\new_[9141]_  | ~\wb_data_i[28] );
  assign \new_[4127]_  = ~\new_[4557]_  & (~\new_[9141]_  | ~\wb_data_i[31] );
  assign \new_[4128]_  = ~\new_[4421]_  | ~\new_[8876]_ ;
  assign \new_[4129]_  = ~\new_[4613]_  | ~\new_[5700]_  | ~\new_[6897]_ ;
  assign \new_[4130]_  = ~\new_[4558]_  & (~\new_[9135]_  | ~\wb_data_i[0] );
  assign \new_[4131]_  = ~\new_[4559]_  & (~\new_[9135]_  | ~\wb_data_i[12] );
  assign \new_[4132]_  = ~\new_[4560]_  & (~\new_[9135]_  | ~\wb_data_i[16] );
  assign \new_[4133]_  = ~\new_[4561]_  & (~\new_[9135]_  | ~\wb_data_i[17] );
  assign \new_[4134]_  = ~\new_[4562]_  & (~\new_[9135]_  | ~\wb_data_i[18] );
  assign \new_[4135]_  = ~\new_[4563]_  & (~\new_[9135]_  | ~\wb_data_i[19] );
  assign \new_[4136]_  = ~\new_[4564]_  & (~\new_[9135]_  | ~\wb_data_i[1] );
  assign \new_[4137]_  = ~\new_[4565]_  & (~\new_[9135]_  | ~\wb_data_i[20] );
  assign \new_[4138]_  = ~\new_[4566]_  & (~\new_[9135]_  | ~\wb_data_i[21] );
  assign \new_[4139]_  = ~\new_[4567]_  & (~\new_[9135]_  | ~\wb_data_i[22] );
  assign \new_[4140]_  = ~\new_[4568]_  & (~\new_[9135]_  | ~\wb_data_i[23] );
  assign \new_[4141]_  = ~\new_[4569]_  & (~\new_[9135]_  | ~\wb_data_i[24] );
  assign \new_[4142]_  = ~\new_[4570]_  & (~\new_[9135]_  | ~\wb_data_i[25] );
  assign \new_[4143]_  = ~\new_[4571]_  & (~\new_[9135]_  | ~\wb_data_i[26] );
  assign \new_[4144]_  = ~\new_[4572]_  & (~\new_[9135]_  | ~\wb_data_i[27] );
  assign \new_[4145]_  = ~\new_[4573]_  & (~\new_[9135]_  | ~\wb_data_i[29] );
  assign \new_[4146]_  = ~\new_[4574]_  & (~\new_[9135]_  | ~\wb_data_i[2] );
  assign \new_[4147]_  = ~\new_[4575]_  & (~\new_[9135]_  | ~\wb_data_i[30] );
  assign \new_[4148]_  = \new_[4550]_  | \new_[4413]_ ;
  assign \new_[4149]_  = ~\new_[4576]_  & (~\new_[9135]_  | ~\wb_data_i[3] );
  assign \new_[4150]_  = ~\new_[4577]_  & (~\new_[9135]_  | ~\wb_data_i[8] );
  assign \new_[4151]_  = ~\new_[4410]_  | ~\new_[8877]_ ;
  assign \new_[4152]_  = ~\new_[4578]_  & (~\new_[9135]_  | ~\wb_data_i[9] );
  assign \new_[4153]_  = ~\new_[4337]_ ;
  assign \new_[4154]_  = ~\new_[4337]_ ;
  assign n3270 = ~\new_[8422]_  | ~\new_[12244]_  | ~\new_[4870]_ ;
  assign \new_[4156]_  = ~\new_[4407]_  & (~\new_[9141]_  | ~\wb_data_i[10] );
  assign \new_[4157]_  = ~\\u1_u2_last_buf_adr_reg[0] ;
  assign n3165 = \new_[4369]_  & \new_[6276]_ ;
  assign \new_[4159]_  = (~\new_[4707]_  | ~\new_[6477]_ ) & (~\new_[5509]_  | ~\new_[10402]_ );
  assign n3300 = \new_[4371]_  & \new_[6276]_ ;
  assign \new_[4161]_  = \\u5_state_reg[1] ;
  assign \new_[4162]_  = ~\new_[4411]_  | ~\new_[8877]_ ;
  assign \new_[4163]_  = ~\new_[5082]_  | ~\new_[4604]_  | ~\new_[5105]_ ;
  assign \new_[4164]_  = ~\new_[4604]_  | ~\new_[5105]_ ;
  assign \new_[4165]_  = ~\new_[4599]_  | (~\new_[9201]_  & ~\new_[12840]_ );
  assign \new_[4166]_  = ~\new_[4601]_  | (~\new_[9202]_  & ~\new_[12650]_ );
  assign \new_[4167]_  = ~\new_[4602]_  | (~\new_[9203]_  & ~\new_[12502]_ );
  assign \new_[4168]_  = ~\new_[4603]_  | (~\new_[9204]_  & ~\new_[12835]_ );
  assign n3305 = \new_[4618]_  ? \wb_addr_i[17]  : \sram_data_i[1] ;
  assign \new_[4170]_  = (~\new_[9789]_  & ~\new_[4697]_ ) | (~\new_[11621]_  & ~\new_[10007]_ );
  assign \new_[4171]_  = ~\new_[4384]_  | (~\new_[3337]_  & ~\new_[12650]_ );
  assign \new_[4172]_  = (~\new_[4699]_  | ~\new_[13595]_ ) & (~\new_[9109]_  | ~\new_[13369]_ );
  assign \new_[4173]_  = ~\new_[4388]_  | (~\new_[3339]_  & ~\new_[12650]_ );
  assign \new_[4174]_  = ~\new_[4390]_  | (~\new_[11624]_  & ~\new_[12650]_ );
  assign \new_[4175]_  = ~\new_[4391]_  | (~\new_[11379]_  & ~\new_[12650]_ );
  assign \new_[4176]_  = ~\new_[4392]_  | (~\new_[10660]_  & ~\new_[12650]_ );
  assign n3605 = \new_[4377]_  & \new_[6288]_ ;
  assign n3315 = \new_[4385]_  & \new_[6288]_ ;
  assign n3260 = \new_[4386]_  & \new_[6288]_ ;
  assign n3310 = \new_[4409]_  & \new_[6276]_ ;
  assign \new_[4181]_  = ~\\u4_u3_buf1_reg[3] ;
  assign \new_[4182]_  = ~\\u4_u3_buf1_reg[29] ;
  assign n3265 = ~\new_[8423]_  | ~\new_[12339]_  | ~\new_[4888]_ ;
  assign \new_[4184]_  = ~\new_[4422]_  & (~\new_[9141]_  | ~\wb_data_i[4] );
  assign \new_[4185]_  = \new_[9173]_  ? \new_[12650]_  : \new_[5025]_ ;
  assign \new_[4186]_  = ~\new_[4701]_  & (~\new_[9142]_  | ~\wb_data_i[5] );
  assign \new_[4187]_  = ~\new_[4700]_  & (~\new_[9142]_  | ~\wb_data_i[4] );
  assign \new_[4188]_  = ~\new_[4703]_  & (~\new_[9142]_  | ~\wb_data_i[7] );
  assign \new_[4189]_  = \new_[9726]_  ? \new_[12650]_  : \new_[5026]_ ;
  assign \new_[4190]_  = u1_clr_sof_time_reg;
  assign \new_[4191]_  = ~u1_frame_no_we_r_reg;
  assign \new_[4192]_  = ~\new_[5419]_  | ~\new_[4718]_  | ~\new_[5355]_ ;
  assign n3690 = ~\new_[4711]_  | ~phy_rst_pad_o;
  assign n3695 = ~\new_[4714]_  | ~phy_rst_pad_o;
  assign n3665 = ~\new_[4715]_  | ~phy_rst_pad_o;
  assign n3735 = ~\new_[12732]_  & (~\new_[6831]_  | ~\new_[5042]_ );
  assign \new_[4197]_  = \\u4_u3_dma_out_cnt_reg[5] ;
  assign n3800 = ~\new_[4698]_  & ~\new_[12794]_ ;
  assign \new_[4199]_  = ~\new_[4719]_  | (~\new_[7695]_  & ~\new_[12502]_ );
  assign n3770 = \new_[4928]_  & \new_[6288]_ ;
  assign \new_[4201]_  = ~\new_[6226]_  | ~\new_[14618]_  | ~\new_[4894]_  | ~\new_[5627]_ ;
  assign \new_[4202]_  = ~\new_[4865]_  | (~\new_[8681]_  & ~\new_[12502]_ );
  assign \new_[4203]_  = ~\new_[4689]_  | (~\new_[10325]_  & ~\new_[12502]_ );
  assign \new_[4204]_  = ~\new_[4671]_  | ~\new_[9138]_ ;
  assign \new_[4205]_  = ~\new_[4772]_  | ~\new_[9138]_ ;
  assign \new_[4206]_  = \\u4_u3_dma_in_cnt_reg[3] ;
  assign \new_[4207]_  = ~\new_[4720]_  | ~\new_[9138]_ ;
  assign \new_[4208]_  = ~\new_[4721]_  | ~\new_[9138]_ ;
  assign \new_[4209]_  = ~\new_[4722]_  | ~\new_[9138]_ ;
  assign \new_[4210]_  = ~\new_[4723]_  | ~\new_[9138]_ ;
  assign \new_[4211]_  = ~\new_[4724]_  | ~\new_[9138]_ ;
  assign \new_[4212]_  = ~\new_[4725]_  | ~\new_[9138]_ ;
  assign \new_[4213]_  = ~\new_[4726]_  | ~\new_[8884]_ ;
  assign \new_[4214]_  = ~\new_[4727]_  | ~\new_[9138]_ ;
  assign \new_[4215]_  = ~\new_[4728]_  | ~\new_[9138]_ ;
  assign \new_[4216]_  = ~\new_[4729]_  | ~\new_[9138]_ ;
  assign \new_[4217]_  = ~\new_[4730]_  | ~\new_[9138]_ ;
  assign \new_[4218]_  = ~\new_[4731]_  | ~\new_[9138]_ ;
  assign \new_[4219]_  = ~\new_[4732]_  | ~\new_[9138]_ ;
  assign \new_[4220]_  = ~\new_[4733]_  | ~\new_[9138]_ ;
  assign \new_[4221]_  = ~\new_[4734]_  | ~\new_[9138]_ ;
  assign \new_[4222]_  = ~\new_[4775]_  | ~\new_[9138]_ ;
  assign n3765 = \new_[4927]_  & \new_[6288]_ ;
  assign \new_[4224]_  = ~\new_[4736]_  | ~\new_[8909]_ ;
  assign \new_[4225]_  = ~\new_[4737]_  | ~\new_[8910]_ ;
  assign n3730 = ~\new_[4408]_ ;
  assign \new_[4227]_  = \new_[9050]_  ? \new_[12650]_  : \new_[5073]_ ;
  assign \new_[4228]_  = \new_[5028]_  ? n9145 : \new_[13801]_ ;
  assign \new_[4229]_  = ~\new_[5093]_  & (~\new_[5089]_  | ~\new_[5092]_ );
  assign \new_[4230]_  = ~\new_[5086]_  & (~\new_[5084]_  | ~\new_[5104]_ );
  assign \new_[4231]_  = ~\new_[5097]_  & (~\new_[5096]_  | ~\new_[5095]_ );
  assign \new_[4232]_  = ~\new_[4762]_  & (~\new_[5099]_  | ~\new_[5097]_ );
  assign \new_[4233]_  = (~\new_[14312]_  | ~\new_[5100]_ ) & (~\new_[5102]_  | ~\new_[5103]_ );
  assign n3660 = ~\new_[8552]_  | ~\new_[12244]_  | ~\new_[5189]_ ;
  assign n3700 = ~\new_[8547]_  | ~\new_[12244]_  | ~\new_[5190]_ ;
  assign \new_[4236]_  = \\u4_u3_dma_out_cnt_reg[8] ;
  assign \new_[4237]_  = \\u4_u3_dma_out_cnt_reg[4] ;
  assign \new_[4238]_  = ~\new_[4738]_  & ~\new_[9135]_ ;
  assign n3655 = \new_[4735]_  & \new_[6288]_ ;
  assign n3745 = \new_[4739]_  & \new_[6288]_ ;
  assign n3740 = \new_[4740]_  & \new_[6288]_ ;
  assign \new_[4242]_  = ~\new_[4712]_  | ~\new_[6621]_ ;
  assign \new_[4243]_  = ~\new_[4705]_  & (~\new_[9142]_  | ~\wb_data_i[13] );
  assign n3670 = ~\new_[12842]_  & (~\new_[5158]_  | ~\new_[11464]_ );
  assign \new_[4245]_  = ~u4_u1_r1_reg;
  assign \new_[4246]_  = ~\new_[4604]_ ;
  assign n3625 = (~\new_[5241]_  | ~\new_[5746]_ ) & (~\new_[5240]_  | ~\new_[5475]_ );
  assign \new_[4248]_  = (~\new_[7483]_  | ~\new_[3314]_ ) & (~\new_[9029]_  | ~\new_[5077]_ );
  assign \new_[4249]_  = ~\new_[4891]_  | ~\new_[6225]_ ;
  assign n3680 = ~\new_[4881]_  | ~phy_rst_pad_o;
  assign \new_[4251]_  = ~\new_[4749]_  & ~\new_[9135]_ ;
  assign \new_[4252]_  = ~\new_[4752]_  & ~\new_[9135]_ ;
  assign \new_[4253]_  = ~\new_[4760]_  & ~\new_[9135]_ ;
  assign \new_[4254]_  = ~\new_[4893]_  & ~\new_[9135]_ ;
  assign n3750 = \new_[4869]_  & \new_[6288]_ ;
  assign n3635 = \new_[4874]_  & \new_[6288]_ ;
  assign n3755 = ~\new_[4871]_  | ~phy_rst_pad_o;
  assign n3760 = ~\new_[4872]_  | ~phy_rst_pad_o;
  assign \new_[4259]_  = ~\new_[4453]_ ;
  assign \new_[4260]_  = ~\new_[5101]_  | ~\new_[4763]_ ;
  assign \new_[4261]_  = ~\new_[4916]_  | ~\new_[9138]_ ;
  assign \new_[4262]_  = ~\new_[4761]_  & ~\new_[5097]_ ;
  assign \new_[4263]_  = \new_[5102]_  & \new_[4763]_ ;
  assign \new_[4264]_  = ~\new_[4753]_  | ~\new_[5082]_ ;
  assign \new_[4265]_  = ~\new_[5084]_  & ~\new_[4751]_ ;
  assign \new_[4266]_  = \new_[4754]_  & \new_[5087]_ ;
  assign \new_[4267]_  = ~\new_[4758]_  | ~\new_[5089]_ ;
  assign \new_[4268]_  = ~\new_[4759]_  | ~\new_[5088]_ ;
  assign \new_[4269]_  = ~\new_[4756]_  & ~\new_[5095]_ ;
  assign \new_[4270]_  = \new_[8261]_  | \new_[4745]_ ;
  assign \new_[4271]_  = ~\new_[4884]_  & (~\new_[9142]_  | ~\wb_data_i[11] );
  assign \new_[4272]_  = ~\new_[4885]_  & (~\new_[9142]_  | ~\wb_data_i[15] );
  assign \new_[4273]_  = ~\new_[4887]_  & (~\new_[9142]_  | ~\wb_data_i[6] );
  assign \new_[4274]_  = ~\new_[4890]_  & (~\new_[5575]_  | ~\new_[5029]_ );
  assign \new_[4275]_  = \new_[6198]_  ? \new_[7307]_  : \new_[5186]_ ;
  assign \new_[4276]_  = \new_[13507]_  ? \new_[7307]_  : \new_[5187]_ ;
  assign n3650 = ~\new_[10710]_  | ~\new_[5234]_  | ~\new_[5233]_ ;
  assign \new_[4278]_  = ~\new_[4921]_  | (~\new_[9166]_  & ~\new_[12502]_ );
  assign \new_[4279]_  = \new_[9711]_  ? \new_[12650]_  : \new_[4998]_ ;
  assign \new_[4280]_  = \new_[9937]_  ? \new_[12650]_  : \new_[5244]_ ;
  assign \new_[4281]_  = \new_[9555]_  ? \new_[12650]_  : \new_[5245]_ ;
  assign \new_[4282]_  = ~\new_[5841]_  | ~\new_[5540]_  | ~\new_[5885]_  | ~\new_[7601]_ ;
  assign \new_[4283]_  = ~\new_[5853]_  | ~\new_[5541]_  | ~\new_[5886]_  | ~\new_[7365]_ ;
  assign \new_[4284]_  = ~\new_[4878]_  & (~\new_[9142]_  | ~\wb_data_i[14] );
  assign \new_[4285]_  = ~\new_[4491]_ ;
  assign \new_[4286]_  = \\u4_u3_dma_in_cnt_reg[8] ;
  assign \new_[4287]_  = ~u4_u2_r1_reg;
  assign \new_[4288]_  = \\u4_u3_dma_in_cnt_reg[5] ;
  assign \new_[4289]_  = \\u4_u3_dma_out_cnt_reg[10] ;
  assign \new_[4290]_  = \\u5_state_reg[2] ;
  assign \new_[4291]_  = \\u4_u3_dma_in_cnt_reg[4] ;
  assign \new_[4292]_  = \\u4_u3_dma_in_cnt_reg[1] ;
  assign \new_[4293]_  = \\u4_u3_dma_in_cnt_reg[2] ;
  assign n3780 = ~\new_[8438]_  | ~\new_[12244]_  | ~\new_[4974]_ ;
  assign n3785 = ~\new_[8529]_  | ~\new_[13162]_  | ~\new_[4975]_ ;
  assign n3645 = ~\new_[8486]_  | ~\new_[12197]_  | ~\new_[4976]_ ;
  assign n3790 = ~\new_[8436]_  | ~\new_[12197]_  | ~\new_[4977]_ ;
  assign n3630 = ~\new_[8545]_  | ~\new_[12197]_  | ~\new_[4978]_ ;
  assign n3795 = ~\new_[8549]_  | ~\new_[12197]_  | ~\new_[4979]_ ;
  assign \new_[4300]_  = ~\new_[4920]_  | (~\new_[9638]_  & ~\new_[12502]_ );
  assign \new_[4301]_  = ~\new_[4922]_  | (~\new_[10323]_  & ~\new_[12502]_ );
  assign \new_[4302]_  = \new_[9598]_  ? \new_[12650]_  : \new_[4993]_ ;
  assign n3685 = ~\new_[4679]_  | ~phy_rst_pad_o;
  assign n3705 = ~\new_[4933]_  | ~phy_rst_pad_o;
  assign \new_[4305]_  = ~\new_[4917]_  & (~\new_[9142]_  | ~\wb_data_i[28] );
  assign \new_[4306]_  = ~\new_[4918]_  & (~\new_[9142]_  | ~\wb_data_i[31] );
  assign n3640 = ~\new_[4934]_  | ~\new_[12058]_ ;
  assign n3620 = ~\new_[4936]_  | ~\new_[12058]_ ;
  assign \new_[4309]_  = ~\new_[4947]_  | ~\new_[5929]_  | ~\new_[7346]_ ;
  assign \new_[4310]_  = ~\new_[4948]_  | ~\new_[5930]_  | ~\new_[7345]_ ;
  assign \new_[4311]_  = ~\new_[4949]_  | ~\new_[5931]_  | ~\new_[7348]_ ;
  assign \new_[4312]_  = ~\new_[4696]_  | ~\new_[9138]_ ;
  assign \new_[4313]_  = \new_[10229]_  ? \new_[12650]_  : \new_[4996]_ ;
  assign \new_[4314]_  = ~\new_[4895]_  & (~\new_[9141]_  | ~\wb_data_i[0] );
  assign \new_[4315]_  = ~\new_[4896]_  & (~\new_[9141]_  | ~\wb_data_i[12] );
  assign \new_[4316]_  = ~\new_[4897]_  & (~\new_[9141]_  | ~\wb_data_i[16] );
  assign \new_[4317]_  = ~\new_[4898]_  & (~\new_[9141]_  | ~\wb_data_i[17] );
  assign \new_[4318]_  = ~\new_[4899]_  & (~\new_[9141]_  | ~\wb_data_i[18] );
  assign \new_[4319]_  = ~\new_[4900]_  & (~\new_[9141]_  | ~\wb_data_i[19] );
  assign \new_[4320]_  = ~\new_[4901]_  & (~\new_[9141]_  | ~\wb_data_i[1] );
  assign \new_[4321]_  = ~\new_[4902]_  & (~\new_[9141]_  | ~\wb_data_i[20] );
  assign \new_[4322]_  = ~\new_[4903]_  & (~\new_[9141]_  | ~\wb_data_i[21] );
  assign \new_[4323]_  = ~\new_[4904]_  & (~\new_[9141]_  | ~\wb_data_i[22] );
  assign \new_[4324]_  = ~\new_[4905]_  & (~\new_[9141]_  | ~\wb_data_i[23] );
  assign \new_[4325]_  = ~\new_[4906]_  & (~\new_[9141]_  | ~\wb_data_i[24] );
  assign \new_[4326]_  = ~\new_[4907]_  & (~\new_[9141]_  | ~\wb_data_i[25] );
  assign \new_[4327]_  = ~\new_[4908]_  & (~\new_[9141]_  | ~\wb_data_i[26] );
  assign \new_[4328]_  = ~\new_[4909]_  & (~\new_[9141]_  | ~\wb_data_i[27] );
  assign \new_[4329]_  = ~\new_[4910]_  & (~\new_[9141]_  | ~\wb_data_i[29] );
  assign \new_[4330]_  = ~\new_[4911]_  & (~\new_[9141]_  | ~\wb_data_i[2] );
  assign \new_[4331]_  = ~\new_[4912]_  & (~\new_[9141]_  | ~\wb_data_i[30] );
  assign \new_[4332]_  = ~\new_[4913]_  & (~\new_[9141]_  | ~\wb_data_i[3] );
  assign \new_[4333]_  = ~\new_[4914]_  & (~\new_[9141]_  | ~\wb_data_i[8] );
  assign \new_[4334]_  = ~\new_[4915]_  & (~\new_[9141]_  | ~\wb_data_i[9] );
  assign \new_[4335]_  = ~\new_[4691]_  & ~\new_[9135]_ ;
  assign \new_[4336]_  = ~\new_[4672]_  | ~\new_[9138]_ ;
  assign \new_[4337]_  = ~\new_[14483]_ ;
  assign \new_[4338]_  = ~\new_[4675]_  & (~\new_[9142]_  | ~\wb_data_i[10] );
  assign \new_[4339]_  = ~\new_[4643]_  & ~\new_[9135]_ ;
  assign \new_[4340]_  = ~\new_[4626]_  & ~\new_[9135]_ ;
  assign \new_[4341]_  = ~\new_[4649]_  & ~\new_[9135]_ ;
  assign n3675 = ~\new_[4744]_  | ~phy_rst_pad_o;
  assign n3615 = \new_[4606]_  & \new_[6288]_ ;
  assign n3710 = \new_[4612]_  & \new_[6288]_ ;
  assign \new_[4345]_  = ~\new_[4673]_  & ~\new_[9135]_ ;
  assign \new_[4346]_  = ~\new_[4674]_  & ~\new_[9135]_ ;
  assign \new_[4347]_  = \\u4_u3_dma_out_cnt_reg[7] ;
  assign n3810 = \new_[4932]_  & \new_[6288]_ ;
  assign n3805 = \new_[4952]_  ? \wb_addr_i[17]  : \sram_data_i[0] ;
  assign n3830 = \new_[4954]_  ? \wb_addr_i[17]  : \sram_data_i[2] ;
  assign n3715 = \new_[4955]_  ? \wb_addr_i[17]  : \sram_data_i[3] ;
  assign \new_[4352]_  = ~\new_[4803]_  | ~\new_[9138]_ ;
  assign \new_[4353]_  = ~u4_u3_r1_reg;
  assign \new_[4354]_  = ~\new_[4661]_  | (~\new_[3502]_  & ~\new_[12502]_ );
  assign \new_[4355]_  = ~\new_[4662]_  | (~\new_[3507]_  & ~\new_[12502]_ );
  assign \new_[4356]_  = ~\new_[4663]_  | (~\new_[11633]_  & ~\new_[12502]_ );
  assign \new_[4357]_  = ~\new_[4664]_  | (~\new_[10398]_  & ~\new_[12502]_ );
  assign \new_[4358]_  = ~\new_[4665]_  | (~\new_[10661]_  & ~\new_[12502]_ );
  assign n3825 = \new_[4638]_  & \new_[6256]_ ;
  assign \new_[4360]_  = \new_[10761]_  ? \new_[12650]_  : \new_[5049]_ ;
  assign \new_[4361]_  = \new_[10308]_  ? \new_[12650]_  : \new_[5050]_ ;
  assign \new_[4362]_  = \new_[10066]_  ? \new_[12650]_  : \new_[5055]_ ;
  assign n3815 = \new_[4650]_  & \new_[6256]_ ;
  assign n3820 = \new_[4669]_  & \new_[6256]_ ;
  assign n3725 = \new_[4670]_  & \new_[6288]_ ;
  assign \new_[4366]_  = \new_[12211]_  ? \new_[12650]_  : \new_[5048]_ ;
  assign n3775 = \new_[4929]_  & \new_[6288]_ ;
  assign n3720 = ~\new_[6963]_  & (~\new_[4990]_  | ~\new_[13522]_ );
  assign \new_[4369]_  = \new_[9174]_  ? \new_[12502]_  : \new_[5410]_ ;
  assign \new_[4370]_  = \\u1_u0_crc16_sum_reg[1] ;
  assign \new_[4371]_  = \new_[9727]_  ? \new_[12502]_  : \new_[5411]_ ;
  assign \new_[4372]_  = \\u1_u0_crc16_sum_reg[11] ;
  assign \new_[4373]_  = ~\new_[4962]_  & (~\new_[6702]_  | ~\new_[5726]_ );
  assign \new_[4374]_  = ~\new_[5022]_  & ~\new_[11428]_ ;
  assign \new_[4375]_  = ~\new_[5034]_  | ~\new_[8860]_ ;
  assign \new_[4376]_  = ~\new_[5035]_  | ~\new_[9128]_ ;
  assign \new_[4377]_  = ~\new_[5036]_  | (~\new_[7696]_  & ~\new_[12835]_ );
  assign \new_[4378]_  = ~\new_[5039]_  | ~\new_[8878]_ ;
  assign \new_[4379]_  = ~\new_[5040]_  | ~\new_[8877]_ ;
  assign \new_[4380]_  = ~\new_[5041]_  | ~\new_[8877]_ ;
  assign \new_[4381]_  = ~\new_[5043]_  | ~\new_[8878]_ ;
  assign \new_[4382]_  = ~\new_[5045]_  | ~\new_[9380]_ ;
  assign \new_[4383]_  = ~\new_[5046]_  | ~\new_[8876]_ ;
  assign \new_[4384]_  = ~\new_[5033]_  | ~\new_[12650]_ ;
  assign \new_[4385]_  = ~\new_[5155]_  | (~\new_[8682]_  & ~\new_[12835]_ );
  assign \new_[4386]_  = ~\new_[5023]_  | (~\new_[9965]_  & ~\new_[12835]_ );
  assign \new_[4387]_  = u0_u0_T1_gt_2_5_uS_reg;
  assign \new_[4388]_  = ~\new_[5051]_  | ~\new_[12650]_ ;
  assign \new_[4389]_  = ~\new_[5066]_  | ~\new_[8911]_ ;
  assign \new_[4390]_  = ~\new_[5052]_  | ~\new_[12650]_ ;
  assign \new_[4391]_  = ~\new_[5053]_  | ~\new_[12650]_ ;
  assign \new_[4392]_  = ~\new_[5054]_  | ~\new_[12650]_ ;
  assign \new_[4393]_  = ~\new_[5064]_  | ~\new_[8909]_ ;
  assign \new_[4394]_  = ~\new_[5057]_  | ~\new_[8911]_ ;
  assign \new_[4395]_  = ~\new_[5058]_  | ~\new_[8910]_ ;
  assign \new_[4396]_  = ~\new_[5059]_  | ~\new_[8910]_ ;
  assign \new_[4397]_  = ~\new_[5060]_  | ~\new_[8909]_ ;
  assign \new_[4398]_  = ~\new_[5061]_  | ~\new_[8910]_ ;
  assign \new_[4399]_  = ~\new_[5062]_  | ~\new_[8910]_ ;
  assign \new_[4400]_  = ~\new_[5063]_  | ~\new_[8910]_ ;
  assign \new_[4401]_  = ~\new_[5065]_  | ~\new_[8910]_ ;
  assign \new_[4402]_  = ~\new_[5067]_  | ~\new_[8909]_ ;
  assign \new_[4403]_  = ~\new_[5068]_  | ~\new_[8909]_ ;
  assign \new_[4404]_  = ~\new_[5069]_  | ~\new_[8909]_ ;
  assign \new_[4405]_  = ~\new_[5070]_  | ~\new_[8910]_ ;
  assign \new_[4406]_  = ~\new_[5071]_  | ~\new_[9448]_ ;
  assign \new_[4407]_  = ~\new_[5072]_  & ~\new_[9141]_ ;
  assign \new_[4408]_  = ~\new_[6621]_  | ~phy_rst_pad_o | ~\new_[5032]_  | ~\new_[7654]_ ;
  assign \new_[4409]_  = \new_[9051]_  ? \new_[12502]_  : \new_[5469]_ ;
  assign \new_[4410]_  = \new_[14194]_  ? \new_[7307]_  : \new_[5484]_ ;
  assign \new_[4411]_  = \new_[13967]_  ? \new_[7307]_  : \new_[5403]_ ;
  assign \new_[4412]_  = ~\new_[4945]_  | ~\new_[8910]_ ;
  assign \new_[4413]_  = u1_u3_to_large_reg;
  assign \new_[4414]_  = ~\new_[5146]_  | ~\new_[8909]_ ;
  assign \new_[4415]_  = ~\new_[5152]_  | ~\new_[8909]_ ;
  assign n3875 = \new_[5047]_  & \new_[6256]_ ;
  assign n3885 = ~\new_[12245]_  & (~\new_[11522]_  | ~\new_[5527]_ );
  assign \new_[4418]_  = ~\new_[5056]_  | (~\new_[8267]_  & ~\new_[12099]_ );
  assign n3880 = \new_[5044]_  & \new_[11609]_ ;
  assign \new_[4420]_  = ~\new_[5074]_  | ~\new_[12650]_ ;
  assign \new_[4421]_  = \new_[13855]_  ? \new_[7307]_  : \new_[5567]_ ;
  assign \new_[4422]_  = ~\new_[5106]_  & ~\new_[9141]_ ;
  assign \new_[4423]_  = ~\new_[5107]_  & ~\new_[9141]_ ;
  assign \new_[4424]_  = ~\new_[5000]_  & ~\new_[9141]_ ;
  assign \new_[4425]_  = ~\new_[5192]_  & ~\new_[9141]_ ;
  assign n3890 = \new_[5159]_  & \new_[6256]_ ;
  assign n3895 = \new_[5160]_  & \new_[6256]_ ;
  assign \new_[4428]_  = ~\new_[8622]_  & ~\new_[5079]_ ;
  assign n3850 = ~\new_[5162]_  | ~phy_rst_pad_o;
  assign n3900 = ~\new_[5163]_  | ~phy_rst_pad_o;
  assign n3905 = ~\new_[5164]_  | ~\new_[12058]_ ;
  assign n3910 = ~\new_[5165]_  | ~\new_[12058]_ ;
  assign n3855 = ~\new_[5166]_  | ~phy_rst_pad_o;
  assign n3915 = ~\new_[5167]_  | ~phy_rst_pad_o;
  assign n3920 = ~\new_[5168]_  | ~\new_[12058]_ ;
  assign n3925 = ~\new_[5169]_  | ~\new_[12058]_ ;
  assign n3840 = ~\new_[5170]_  | ~\new_[13165]_ ;
  assign n3930 = ~\new_[5171]_  | ~\new_[13165]_ ;
  assign n3935 = ~\new_[5172]_  | ~phy_rst_pad_o;
  assign n3940 = ~\new_[5173]_  | ~phy_rst_pad_o;
  assign n3835 = ~\new_[5175]_  | ~phy_rst_pad_o;
  assign n3950 = ~\new_[5176]_  | ~phy_rst_pad_o;
  assign n3945 = ~\new_[5177]_  | ~phy_rst_pad_o;
  assign n4020 = ~\new_[5178]_  | ~phy_rst_pad_o;
  assign n3960 = ~\new_[5179]_  | ~phy_rst_pad_o;
  assign n3955 = ~\new_[5180]_  | ~phy_rst_pad_o;
  assign n4015 = ~\new_[5181]_  | ~phy_rst_pad_o;
  assign n3970 = ~\new_[5182]_  | ~phy_rst_pad_o;
  assign n3965 = ~\new_[5183]_  | ~phy_rst_pad_o;
  assign n4010 = ~\new_[5147]_  | (~\new_[8853]_  & ~\new_[12804]_ );
  assign \new_[4451]_  = \new_[5081]_  & \new_[5104]_ ;
  assign n3860 = ~\new_[4716]_ ;
  assign \new_[4453]_  = \new_[5096]_  & \new_[5099]_ ;
  assign \new_[4454]_  = \new_[5096]_  & \new_[5090]_ ;
  assign \new_[4455]_  = ~\new_[5091]_  & ~\new_[5087]_ ;
  assign \new_[4456]_  = \new_[5098]_  & \new_[5099]_ ;
  assign \new_[4457]_  = \new_[5100]_  & \new_[5101]_ ;
  assign \new_[4458]_  = ~\new_[5100]_  | ~\new_[5514]_ ;
  assign \new_[4459]_  = ~\new_[5105]_  | ~\new_[5080]_ ;
  assign \new_[4460]_  = ~\new_[5161]_  | ~\new_[12650]_ ;
  assign n3980 = ~\new_[12794]_  & (~\new_[6832]_  | ~\new_[5586]_ );
  assign n3975 = ~\new_[5618]_  | ~\new_[7199]_  | ~rst_i | ~\new_[7529]_ ;
  assign \new_[4463]_  = \new_[13918]_  ? \new_[7307]_  : \new_[5546]_ ;
  assign \new_[4464]_  = ~\new_[5076]_  | ~\new_[8634]_ ;
  assign \new_[4465]_  = \new_[13808]_  ? \new_[7307]_  : \new_[5547]_ ;
  assign \new_[4466]_  = \new_[6484]_  ? \new_[7307]_  : \new_[5548]_ ;
  assign \new_[4467]_  = \new_[13829]_  ? \new_[7307]_  : \new_[5549]_ ;
  assign \new_[4468]_  = \new_[6168]_  ? \new_[7307]_  : \new_[5550]_ ;
  assign \new_[4469]_  = \new_[6319]_  ? \new_[7307]_  : \new_[5551]_ ;
  assign \new_[4470]_  = \new_[6320]_  ? \new_[7307]_  : \new_[5552]_ ;
  assign \new_[4471]_  = \new_[6238]_  ? \new_[7307]_  : \new_[5553]_ ;
  assign \new_[4472]_  = \new_[6322]_  ? \new_[7307]_  : \new_[5554]_ ;
  assign \new_[4473]_  = \new_[6234]_  ? \new_[7307]_  : \new_[5555]_ ;
  assign \new_[4474]_  = \new_[6323]_  ? \new_[7307]_  : \new_[5556]_ ;
  assign \new_[4475]_  = \new_[6326]_  ? \new_[7307]_  : \new_[5557]_ ;
  assign \new_[4476]_  = \new_[14252]_  ? \new_[7307]_  : \new_[5558]_ ;
  assign \new_[4477]_  = \new_[13559]_  ? \new_[7307]_  : \new_[5559]_ ;
  assign \new_[4478]_  = ~\new_[6687]_  | ~\new_[7183]_  | ~\new_[5603]_ ;
  assign \new_[4479]_  = \new_[14179]_  ? \new_[7307]_  : \new_[5560]_ ;
  assign \new_[4480]_  = ~\new_[5153]_  | (~\new_[10039]_  & ~\new_[11079]_ );
  assign \new_[4481]_  = ~\new_[5231]_  | (~\new_[9167]_  & ~\new_[12835]_ );
  assign \new_[4482]_  = \new_[6512]_  ? \new_[7549]_  : \new_[5544]_ ;
  assign \new_[4483]_  = \new_[14067]_  ? \new_[7549]_  : \new_[5545]_ ;
  assign \new_[4484]_  = \new_[9712]_  ? \new_[12502]_  : \new_[5375]_ ;
  assign \new_[4485]_  = \new_[9647]_  ? \new_[12502]_  : \new_[5599]_ ;
  assign \new_[4486]_  = \new_[9557]_  ? \new_[12502]_  : \new_[5601]_ ;
  assign \new_[4487]_  = ~\new_[5214]_  | ~\new_[8909]_ ;
  assign n3865 = \new_[5481]_  ^ \new_[5575]_ ;
  assign \new_[4489]_  = ~\new_[6064]_  | ~\new_[5796]_  | ~\new_[6085]_  | ~\new_[7602]_ ;
  assign \new_[4490]_  = ~\new_[4748]_ ;
  assign \new_[4491]_  = ~\\u1_u3_new_size_reg[1] ;
  assign \new_[4492]_  = \new_[13857]_  ? \new_[7307]_  : \new_[5342]_ ;
  assign n3985 = \new_[5235]_  & \new_[6256]_ ;
  assign \new_[4494]_  = \new_[13542]_  ? \new_[7307]_  : \new_[5348]_ ;
  assign n4000 = \new_[5236]_  & \new_[6256]_ ;
  assign n3990 = \new_[5237]_  & \new_[6256]_ ;
  assign n3995 = \new_[5238]_  & \new_[6256]_ ;
  assign n3845 = \new_[5239]_  & \new_[6256]_ ;
  assign \new_[4499]_  = \new_[14006]_  ? \new_[7307]_  : \new_[5352]_ ;
  assign \new_[4500]_  = \\u1_u0_crc16_sum_reg[15] ;
  assign \new_[4501]_  = \\u4_int_srcb_reg[6] ;
  assign \new_[4502]_  = \\u1_u0_crc16_sum_reg[0] ;
  assign \new_[4503]_  = \\u1_u0_crc16_sum_reg[10] ;
  assign \new_[4504]_  = \\u1_u0_crc16_sum_reg[12] ;
  assign \new_[4505]_  = \\u1_u0_crc16_sum_reg[14] ;
  assign \new_[4506]_  = \\u1_u0_crc16_sum_reg[3] ;
  assign \new_[4507]_  = \\u1_u0_crc16_sum_reg[4] ;
  assign \new_[4508]_  = \\u1_u0_crc16_sum_reg[5] ;
  assign \new_[4509]_  = \\u1_u0_crc16_sum_reg[7] ;
  assign \new_[4510]_  = \\u1_u0_crc16_sum_reg[8] ;
  assign \new_[4511]_  = \\u1_u0_crc16_sum_reg[9] ;
  assign \new_[4512]_  = \\u1_u3_adr_r_reg[10] ;
  assign \new_[4513]_  = \\u1_u3_adr_r_reg[13] ;
  assign \new_[4514]_  = \\u1_u3_adr_r_reg[3] ;
  assign \new_[4515]_  = \\u1_u3_adr_r_reg[4] ;
  assign \new_[4516]_  = ~\new_[5246]_  | ~\new_[12650]_ ;
  assign \new_[4517]_  = ~\new_[6688]_  & (~\new_[5351]_  | ~\new_[5717]_ );
  assign \new_[4518]_  = ~\new_[5230]_  | (~\new_[9687]_  & ~\new_[12835]_ );
  assign \new_[4519]_  = ~\new_[5232]_  | (~\new_[10689]_  & ~\new_[12835]_ );
  assign \new_[4520]_  = \new_[9599]_  ? \new_[12502]_  : \new_[5370]_ ;
  assign \new_[4521]_  = ~\new_[4984]_  | ~\new_[8876]_ ;
  assign \new_[4522]_  = ~\new_[4985]_  | ~\new_[9380]_ ;
  assign \new_[4523]_  = \new_[10231]_  ? \new_[12502]_  : \new_[5373]_ ;
  assign \new_[4524]_  = ~\new_[5024]_  & ~\new_[9141]_ ;
  assign \new_[4525]_  = ~\new_[5193]_  & (~\new_[9142]_  | ~\wb_data_i[0] );
  assign \new_[4526]_  = ~\new_[5194]_  & (~\new_[9142]_  | ~\wb_data_i[12] );
  assign \new_[4527]_  = ~\new_[5195]_  & (~\new_[9142]_  | ~\wb_data_i[16] );
  assign \new_[4528]_  = ~\new_[5196]_  & (~\new_[9142]_  | ~\wb_data_i[17] );
  assign \new_[4529]_  = ~\new_[5197]_  & (~\new_[9142]_  | ~\wb_data_i[18] );
  assign \new_[4530]_  = ~\new_[5198]_  & (~\new_[9142]_  | ~\wb_data_i[19] );
  assign \new_[4531]_  = ~\new_[5199]_  & (~\new_[9142]_  | ~\wb_data_i[1] );
  assign \new_[4532]_  = ~\new_[5200]_  & (~\new_[9142]_  | ~\wb_data_i[20] );
  assign \new_[4533]_  = ~\new_[5201]_  & (~\new_[9142]_  | ~\wb_data_i[21] );
  assign \new_[4534]_  = ~\new_[5202]_  & (~\new_[9142]_  | ~\wb_data_i[22] );
  assign \new_[4535]_  = ~\new_[5203]_  & (~\new_[9142]_  | ~\wb_data_i[23] );
  assign \new_[4536]_  = ~\new_[5204]_  & (~\new_[9142]_  | ~\wb_data_i[24] );
  assign \new_[4537]_  = ~\new_[5205]_  & (~\new_[9142]_  | ~\wb_data_i[25] );
  assign \new_[4538]_  = ~\new_[5206]_  & (~\new_[9142]_  | ~\wb_data_i[26] );
  assign \new_[4539]_  = ~\new_[5207]_  & (~\new_[9142]_  | ~\wb_data_i[27] );
  assign \new_[4540]_  = ~\new_[5208]_  & (~\new_[9142]_  | ~\wb_data_i[29] );
  assign \new_[4541]_  = ~\new_[5209]_  & (~\new_[9142]_  | ~\wb_data_i[2] );
  assign \new_[4542]_  = ~\new_[5210]_  & (~\new_[9142]_  | ~\wb_data_i[30] );
  assign \new_[4543]_  = ~\new_[5211]_  & (~\new_[9142]_  | ~\wb_data_i[3] );
  assign \new_[4544]_  = ~\new_[5212]_  & (~\new_[9142]_  | ~\wb_data_i[8] );
  assign \new_[4545]_  = ~\new_[5213]_  & (~\new_[9142]_  | ~\wb_data_i[9] );
  assign \new_[4546]_  = ~\new_[5027]_  | ~\new_[8910]_ ;
  assign \new_[4547]_  = ~\new_[4964]_  & ~\new_[9141]_ ;
  assign \new_[4548]_  = ~\new_[4965]_  & ~\new_[9141]_ ;
  assign \new_[4549]_  = ~\new_[4968]_  & ~\new_[9141]_ ;
  assign \new_[4550]_  = u1_u3_to_small_reg;
  assign \new_[4551]_  = ~\new_[4999]_  | ~\new_[8909]_ ;
  assign \new_[4552]_  = \\u1_u0_crc16_sum_reg[13] ;
  assign \new_[4553]_  = \\u1_u0_crc16_sum_reg[6] ;
  assign \new_[4554]_  = \new_[4967]_  & \new_[6469]_ ;
  assign \new_[4555]_  = \new_[13896]_  ? \new_[7307]_  : \new_[5464]_ ;
  assign \new_[4556]_  = ~\new_[4991]_  & ~\new_[9141]_ ;
  assign \new_[4557]_  = ~\new_[4992]_  & ~\new_[9141]_ ;
  assign \new_[4558]_  = ~\new_[5001]_  & ~\new_[9135]_ ;
  assign \new_[4559]_  = ~\new_[5002]_  & ~\new_[9135]_ ;
  assign \new_[4560]_  = ~\new_[5003]_  & ~\new_[9135]_ ;
  assign \new_[4561]_  = ~\new_[5004]_  & ~\new_[9135]_ ;
  assign \new_[4562]_  = ~\new_[5005]_  & ~\new_[9135]_ ;
  assign \new_[4563]_  = ~\new_[5006]_  & ~\new_[9135]_ ;
  assign \new_[4564]_  = ~\new_[5007]_  & ~\new_[9135]_ ;
  assign \new_[4565]_  = ~\new_[5008]_  & ~\new_[9135]_ ;
  assign \new_[4566]_  = ~\new_[5009]_  & ~\new_[9135]_ ;
  assign \new_[4567]_  = ~\new_[5010]_  & ~\new_[9135]_ ;
  assign \new_[4568]_  = ~\new_[5011]_  & ~\new_[9135]_ ;
  assign \new_[4569]_  = ~\new_[5012]_  & ~\new_[9135]_ ;
  assign \new_[4570]_  = ~\new_[5013]_  & ~\new_[9135]_ ;
  assign \new_[4571]_  = ~\new_[5014]_  & ~\new_[9135]_ ;
  assign \new_[4572]_  = ~\new_[5015]_  & ~\new_[9135]_ ;
  assign \new_[4573]_  = ~\new_[5016]_  & ~\new_[9135]_ ;
  assign \new_[4574]_  = ~\new_[5017]_  & ~\new_[9135]_ ;
  assign \new_[4575]_  = ~\new_[5018]_  & ~\new_[9135]_ ;
  assign \new_[4576]_  = ~\new_[5019]_  & ~\new_[9135]_ ;
  assign \new_[4577]_  = ~\new_[5020]_  & ~\new_[9135]_ ;
  assign \new_[4578]_  = ~\new_[5021]_  & ~\new_[9135]_ ;
  assign \new_[4579]_  = ~\new_[4994]_  | ~\new_[12650]_ ;
  assign \new_[4580]_  = ~\new_[4995]_  | ~\new_[12650]_ ;
  assign \new_[4581]_  = ~\new_[4997]_  | ~\new_[12650]_ ;
  assign \new_[4582]_  = ~\new_[3716]_  & (~\new_[5416]_  | ~\new_[8633]_ );
  assign \new_[4583]_  = ~\new_[3595]_  & (~\new_[5416]_  | ~\new_[8970]_ );
  assign \new_[4584]_  = ~\new_[3739]_  & (~\new_[5416]_  | ~\new_[7866]_ );
  assign \new_[4585]_  = ~\new_[3741]_  & (~\new_[5416]_  | ~\new_[8247]_ );
  assign \new_[4586]_  = ~\new_[5717]_  | ~\new_[4958]_  | ~\new_[5423]_ ;
  assign \new_[4587]_  = ~\new_[4973]_  | (~\new_[3710]_  & ~\new_[12835]_ );
  assign \new_[4588]_  = ~\new_[4980]_  | (~\new_[3718]_  & ~\new_[12835]_ );
  assign \new_[4589]_  = ~\new_[4981]_  | (~\new_[11632]_  & ~\new_[12835]_ );
  assign \new_[4590]_  = ~\new_[4982]_  | (~\new_[11044]_  & ~\new_[12835]_ );
  assign \new_[4591]_  = ~\new_[4983]_  | (~\new_[10663]_  & ~\new_[12835]_ );
  assign \new_[4592]_  = \new_[10763]_  ? \new_[12502]_  : \new_[5455]_ ;
  assign n3870 = \new_[4963]_  & \new_[6256]_ ;
  assign \new_[4594]_  = \new_[10310]_  ? \new_[12502]_  : \new_[5456]_ ;
  assign \new_[4595]_  = \new_[10415]_  ? \new_[12502]_  : \new_[5462]_ ;
  assign \new_[4596]_  = \new_[12209]_  ? \new_[12502]_  : \new_[5454]_ ;
  assign \new_[4597]_  = \\u1_u0_crc16_sum_reg[2] ;
  assign \new_[4598]_  = ~\new_[5150]_  | ~\new_[8909]_ ;
  assign \new_[4599]_  = ~\new_[4986]_  | ~\new_[12840]_ ;
  assign \new_[4600]_  = n4965 | \new_[12326]_  | \new_[9790]_  | \new_[11657]_ ;
  assign \new_[4601]_  = ~\new_[4987]_  | ~\new_[12650]_ ;
  assign \new_[4602]_  = ~\new_[4988]_  | ~\new_[12502]_ ;
  assign \new_[4603]_  = ~\new_[4989]_  | ~\new_[12835]_ ;
  assign \new_[4604]_  = \new_[14548]_  & n4975;
  assign n4005 = \new_[14548]_  ^ n4975;
  assign \new_[4606]_  = \new_[9175]_  ? \new_[12835]_  : \new_[5701]_ ;
  assign \new_[4607]_  = \\u1_u1_crc16_reg[14] ;
  assign \new_[4608]_  = \\u4_buf1_reg[25] ;
  assign \new_[4609]_  = \\u4_buf1_reg[29] ;
  assign \new_[4610]_  = ~\new_[5474]_  | ~\new_[8860]_ ;
  assign \new_[4611]_  = ~\new_[5478]_  | ~\new_[8860]_ ;
  assign \new_[4612]_  = \new_[9731]_  ? \new_[12835]_  : \new_[5702]_ ;
  assign \new_[4613]_  = (~\new_[7656]_  | ~\new_[5694]_ ) & (~\new_[6767]_  | ~\new_[5694]_ );
  assign \new_[4614]_  = ~\new_[5483]_  | ~\new_[8860]_ ;
  assign \new_[4615]_  = \\u4_csr_reg[1] ;
  assign \new_[4616]_  = \\u4_buf1_reg[21] ;
  assign \new_[4617]_  = ~\\u4_buf1_reg[14] ;
  assign \new_[4618]_  = \\u4_dout_reg[1] ;
  assign \new_[4619]_  = \\u4_buf1_reg[18] ;
  assign \new_[4620]_  = \\u4_csr_reg[5] ;
  assign \new_[4621]_  = ~\\u4_buf0_reg[3] ;
  assign n4065 = \new_[5404]_  & \new_[11612]_ ;
  assign n4105 = \new_[5405]_  & \new_[11592]_ ;
  assign \new_[4624]_  = ~\new_[5465]_  | ~\new_[8860]_ ;
  assign \new_[4625]_  = ~\new_[5457]_  | ~\new_[8860]_ ;
  assign \new_[4626]_  = ~\new_[5406]_  & (~\new_[6084]_  | ~\new_[13951]_ );
  assign \new_[4627]_  = ~\new_[5438]_  | ~\new_[8860]_ ;
  assign \new_[4628]_  = ~\new_[5433]_  | ~\new_[8860]_ ;
  assign \new_[4629]_  = ~\new_[5435]_  | ~\new_[8860]_ ;
  assign \new_[4630]_  = ~\new_[5434]_  | ~\new_[9128]_ ;
  assign \new_[4631]_  = ~\new_[5429]_  | ~\new_[8860]_ ;
  assign \new_[4632]_  = ~\new_[5452]_  | ~\new_[8860]_ ;
  assign \new_[4633]_  = ~\new_[5430]_  | ~\new_[9128]_ ;
  assign \new_[4634]_  = ~\new_[5437]_  | ~\new_[9128]_ ;
  assign \new_[4635]_  = ~\new_[5451]_  | ~\new_[9128]_ ;
  assign \new_[4636]_  = ~\new_[5442]_  | ~\new_[8860]_ ;
  assign \new_[4637]_  = ~\new_[5463]_  | ~\new_[8860]_ ;
  assign \new_[4638]_  = ~\new_[5422]_  | (~\new_[7693]_  & ~\new_[12840]_ );
  assign \new_[4639]_  = ~\new_[5450]_  | ~\new_[8860]_ ;
  assign \new_[4640]_  = ~\new_[5453]_  | ~\new_[8860]_ ;
  assign \new_[4641]_  = ~\\u4_buf0_reg[7] ;
  assign \new_[4642]_  = ~\new_[5431]_  | ~\new_[8860]_ ;
  assign \new_[4643]_  = ~\new_[5407]_  & (~\new_[6084]_  | ~\new_[14132]_ );
  assign \new_[4644]_  = ~\new_[5440]_  | ~\new_[9128]_ ;
  assign \new_[4645]_  = ~\new_[5441]_  | ~\new_[9128]_ ;
  assign \new_[4646]_  = ~\new_[5432]_  | ~\new_[9425]_ ;
  assign \new_[4647]_  = ~\new_[5428]_  | ~\new_[9425]_ ;
  assign \new_[4648]_  = ~\\u4_buf1_reg[10] ;
  assign \new_[4649]_  = ~\new_[5409]_  & (~\new_[6084]_  | ~\new_[13701]_ );
  assign \new_[4650]_  = ~\new_[5402]_  | (~\new_[9963]_  & ~\new_[12840]_ );
  assign \new_[4651]_  = \\u4_csr_reg[9] ;
  assign \new_[4652]_  = ~\new_[5439]_  | ~\new_[8860]_ ;
  assign \new_[4653]_  = \\u0_u0_state_reg[13] ;
  assign \new_[4654]_  = ~\new_[6631]_  | (~\new_[5721]_  & ~\new_[6904]_ );
  assign \new_[4655]_  = ~\new_[5443]_  | ~\new_[9138]_ ;
  assign \new_[4656]_  = ~\new_[5444]_  | ~\new_[8884]_ ;
  assign \new_[4657]_  = ~\new_[5445]_  | ~\new_[9138]_ ;
  assign \new_[4658]_  = ~\new_[5446]_  | ~\new_[8884]_ ;
  assign \new_[4659]_  = ~\new_[5447]_  | ~\new_[9138]_ ;
  assign \new_[4660]_  = ~\new_[5448]_  | ~\new_[9138]_ ;
  assign \new_[4661]_  = ~\new_[5427]_  | ~\new_[12502]_ ;
  assign \new_[4662]_  = ~\new_[5458]_  | ~\new_[12502]_ ;
  assign \new_[4663]_  = ~\new_[5459]_  | ~\new_[12502]_ ;
  assign \new_[4664]_  = ~\new_[5460]_  | ~\new_[12502]_ ;
  assign \new_[4665]_  = ~\new_[5461]_  | ~\new_[12502]_ ;
  assign \new_[4666]_  = \\u0_u0_idle_cnt1_reg[1] ;
  assign \new_[4667]_  = ~\new_[7471]_  & (~\new_[5748]_  | ~\new_[2301]_ );
  assign \new_[4668]_  = ~\new_[10801]_  & (~\new_[5748]_  | ~\new_[14135]_ );
  assign \new_[4669]_  = \new_[9049]_  ? \new_[12840]_  : \new_[5742]_ ;
  assign \new_[4670]_  = \new_[9052]_  ? \new_[12835]_  : \new_[5743]_ ;
  assign \new_[4671]_  = \new_[13672]_  ? \new_[7549]_  : \new_[5613]_ ;
  assign \new_[4672]_  = \new_[13653]_  ? \new_[7549]_  : \new_[5699]_ ;
  assign \new_[4673]_  = ~\new_[5414]_  & (~\new_[6084]_  | ~\new_[13725]_ );
  assign \new_[4674]_  = ~\new_[5415]_  & (~\new_[6084]_  | ~\new_[13868]_ );
  assign \new_[4675]_  = ~\new_[5471]_  & ~\new_[9142]_ ;
  assign \new_[4676]_  = \\u4_buf0_reg[29] ;
  assign \new_[4677]_  = ~\\u0_u0_ps_cnt_reg[2] ;
  assign \new_[4678]_  = ~\\u0_u0_idle_cnt1_reg[4] ;
  assign \new_[4679]_  = ~\new_[5417]_  & (~\new_[9137]_  | ~\wb_data_i[13] );
  assign n4080 = ~\new_[5467]_  & ~\new_[13296]_ ;
  assign n4100 = \new_[5449]_  & \new_[6256]_ ;
  assign n4075 = \new_[5466]_  & \new_[6256]_ ;
  assign \new_[4683]_  = \\u0_u0_idle_cnt1_reg[6] ;
  assign n4070 = \new_[5468]_  & \new_[6256]_ ;
  assign \new_[4685]_  = ~\\u0_u0_idle_cnt1_reg[7] ;
  assign \new_[4686]_  = \\u4_csr_reg[30] ;
  assign n4055 = \new_[5436]_  & \new_[11439]_ ;
  assign n4030 = ~\new_[5022]_ ;
  assign \new_[4689]_  = ~\new_[5470]_  | ~\new_[12502]_ ;
  assign \new_[4690]_  = \\u4_buf0_reg[30] ;
  assign \new_[4691]_  = ~\new_[5418]_  & (~\new_[6084]_  | ~\new_[13871]_ );
  assign \wb_data_o[23]  = \\u5_wb_data_o_reg[23] ;
  assign \new_[4693]_  = ~\new_[5568]_  | ~\new_[8860]_ ;
  assign \new_[4694]_  = \new_[5753]_  ? n9145 : \new_[13785]_ ;
  assign \new_[4695]_  = \\u4_buf0_reg[21] ;
  assign \new_[4696]_  = \new_[13693]_  ? \new_[7549]_  : \new_[5850]_ ;
  assign \new_[4697]_  = ~\new_[5472]_  & ~\new_[2611]_ ;
  assign \new_[4698]_  = ~\new_[9488]_  & ~\new_[5357]_ ;
  assign \new_[4699]_  = ~\new_[5605]_  & ~\new_[9789]_ ;
  assign \new_[4700]_  = ~\new_[5496]_  & ~\new_[9142]_ ;
  assign \new_[4701]_  = ~\new_[5497]_  & ~\new_[9142]_ ;
  assign \new_[4702]_  = \\u4_csr_reg[27] ;
  assign \new_[4703]_  = ~\new_[5500]_  & ~\new_[9142]_ ;
  assign n4040 = \new_[5589]_  & \new_[6256]_ ;
  assign \new_[4705]_  = ~\new_[5583]_  & ~\new_[9142]_ ;
  assign \new_[4706]_  = \new_[5746]_  ? \new_[7939]_  : \new_[7430]_ ;
  assign \new_[4707]_  = ~\new_[10801]_  & ~\new_[5482]_ ;
  assign n4085 = \new_[5528]_  & \new_[6256]_ ;
  assign \new_[4709]_  = \\u4_buf0_reg[25] ;
  assign \new_[4710]_  = ~\new_[6694]_  | (~\new_[7939]_  & ~\new_[5746]_ );
  assign \new_[4711]_  = ~\new_[5529]_  & (~\new_[9137]_  | ~\wb_data_i[11] );
  assign \new_[4712]_  = ~\new_[5032]_ ;
  assign n4050 = \new_[5534]_  & \new_[6256]_ ;
  assign \new_[4714]_  = ~\new_[5530]_  & (~\new_[9137]_  | ~\wb_data_i[15] );
  assign \new_[4715]_  = ~\new_[5531]_  & (~\new_[9137]_  | ~\wb_data_i[6] );
  assign \new_[4716]_  = ~\new_[5821]_  & (~\new_[9200]_  | ~\new_[5848]_ );
  assign \new_[4717]_  = ~\new_[9992]_  & ~\new_[5473]_ ;
  assign \new_[4718]_  = ~\new_[5719]_  | (~\new_[5849]_  & ~\new_[5747]_ );
  assign \new_[4719]_  = ~\new_[5532]_  | ~\new_[12502]_ ;
  assign \new_[4720]_  = \new_[13637]_  ? \new_[7549]_  : \new_[5806]_ ;
  assign \new_[4721]_  = \new_[13968]_  ? \new_[7549]_  : \new_[5807]_ ;
  assign \new_[4722]_  = \new_[6341]_  ? \new_[7549]_  : \new_[5808]_ ;
  assign \new_[4723]_  = \new_[13892]_  ? \new_[7549]_  : \new_[5809]_ ;
  assign \new_[4724]_  = \new_[6592]_  ? \new_[7549]_  : \new_[5810]_ ;
  assign \new_[4725]_  = \new_[6343]_  ? \new_[7549]_  : \new_[5811]_ ;
  assign \new_[4726]_  = \new_[6345]_  ? \new_[7549]_  : \new_[5812]_ ;
  assign \new_[4727]_  = \new_[6551]_  ? \new_[7549]_  : \new_[5813]_ ;
  assign \new_[4728]_  = \new_[6346]_  ? \new_[7549]_  : \new_[5814]_ ;
  assign \new_[4729]_  = \new_[6347]_  ? \new_[7549]_  : \new_[5815]_ ;
  assign \new_[4730]_  = \new_[6348]_  ? \new_[7549]_  : \new_[5816]_ ;
  assign \new_[4731]_  = \new_[6012]_  ? \new_[7549]_  : \new_[5817]_ ;
  assign \new_[4732]_  = \new_[14066]_  ? \new_[7549]_  : \new_[5818]_ ;
  assign \new_[4733]_  = \new_[13809]_  ? \new_[7549]_  : \new_[5819]_ ;
  assign \new_[4734]_  = \new_[13880]_  ? \new_[7549]_  : \new_[5820]_ ;
  assign \new_[4735]_  = \new_[9716]_  ? \new_[12835]_  : \new_[5634]_ ;
  assign \new_[4736]_  = \new_[6092]_  ? \new_[7857]_  : \new_[5804]_ ;
  assign \new_[4737]_  = \new_[13973]_  ? \new_[7857]_  : \new_[5805]_ ;
  assign \new_[4738]_  = ~\new_[5539]_  & (~\new_[6084]_  | ~\new_[13879]_ );
  assign \new_[4739]_  = \new_[9938]_  ? \new_[12835]_  : \new_[5881]_ ;
  assign \new_[4740]_  = \new_[9556]_  ? \new_[12835]_  : \new_[5884]_ ;
  assign \new_[4741]_  = \\u0_u0_state_reg[11] ;
  assign \new_[4742]_  = ~\\u1_u3_adr_r_reg[12] ;
  assign \new_[4743]_  = ~\\u1_u3_adr_r_reg[16] ;
  assign \new_[4744]_  = ~\new_[5533]_  & (~\new_[9137]_  | ~\wb_data_i[14] );
  assign \new_[4745]_  = ~u1_u3_buf0_st_max_reg;
  assign \new_[4746]_  = ~\new_[9481]_  | ~\new_[5538]_ ;
  assign \new_[4747]_  = ~\new_[13330]_  & ~\new_[5510]_ ;
  assign \new_[4748]_  = ~\new_[13330]_  & ~\new_[5512]_ ;
  assign \new_[4749]_  = ~\new_[5507]_  & (~\new_[6652]_  | ~\new_[13767]_ );
  assign \new_[4750]_  = ~\new_[5080]_ ;
  assign \new_[4751]_  = ~\new_[5081]_ ;
  assign \new_[4752]_  = ~\new_[5506]_  & (~\new_[6084]_  | ~\new_[14138]_ );
  assign \new_[4753]_  = ~\new_[5083]_ ;
  assign \new_[4754]_  = ~\new_[5085]_ ;
  assign \new_[4755]_  = ~\new_[5086]_ ;
  assign \new_[4756]_  = ~\new_[5090]_ ;
  assign \new_[4757]_  = ~\new_[5091]_ ;
  assign \new_[4758]_  = ~\new_[5093]_ ;
  assign \new_[4759]_  = ~\new_[5094]_ ;
  assign \new_[4760]_  = ~\new_[5508]_  & (~\new_[6084]_  | ~\new_[14170]_ );
  assign \new_[4761]_  = ~\new_[5096]_ ;
  assign \new_[4762]_  = ~\new_[5098]_ ;
  assign \new_[4763]_  = ~\new_[5103]_ ;
  assign \new_[4764]_  = ~\new_[5104]_ ;
  assign \new_[4765]_  = \\u1_u1_crc16_reg[10] ;
  assign \new_[4766]_  = \\u1_u1_crc16_reg[13] ;
  assign \new_[4767]_  = \\u1_u1_crc16_reg[12] ;
  assign \new_[4768]_  = \\u4_csr_reg[23] ;
  assign \wb_data_o[22]  = \\u5_wb_data_o_reg[22] ;
  assign n4035 = \new_[5590]_  & \new_[6256]_ ;
  assign n4090 = \new_[5591]_  & \new_[6256]_ ;
  assign \new_[4772]_  = \new_[13677]_  ? \new_[7549]_  : \new_[5614]_ ;
  assign \wb_data_o[7]  = \\u5_wb_data_o_reg[7] ;
  assign \new_[4774]_  = \\u0_u0_idle_cnt1_reg[3] ;
  assign \new_[4775]_  = \new_[13765]_  ? \new_[7549]_  : \new_[5616]_ ;
  assign \wb_data_o[8]  = \\u5_wb_data_o_reg[8] ;
  assign \new_[4777]_  = u0_u0_T1_gt_3_0_mS_reg;
  assign \new_[4778]_  = \\u4_int_srcb_reg[3] ;
  assign \new_[4779]_  = \\u0_u0_idle_cnt1_reg[0] ;
  assign \new_[4780]_  = \\u0_u0_idle_cnt1_reg[2] ;
  assign \new_[4781]_  = ~u1_u0_rxv2_reg;
  assign \new_[4782]_  = ~\\u0_u0_idle_cnt1_reg[5] ;
  assign \new_[4783]_  = ~\\u0_u0_ps_cnt_reg[0] ;
  assign \new_[4784]_  = ~\\u0_u0_ps_cnt_reg[1] ;
  assign \new_[4785]_  = ~\\u0_u0_ps_cnt_reg[3] ;
  assign n9120 = resume_req_r_reg;
  assign \new_[4787]_  = \\u4_csr_reg[12] ;
  assign \new_[4788]_  = \\u4_csr_reg[15] ;
  assign \new_[4789]_  = ~\\u4_csr_reg[17] ;
  assign \new_[4790]_  = \\u4_csr_reg[22] ;
  assign \new_[4791]_  = \\u4_csr_reg[24] ;
  assign \new_[4792]_  = \\u4_csr_reg[25] ;
  assign \new_[4793]_  = \\u4_csr_reg[26] ;
  assign \new_[4794]_  = \\u4_csr_reg[28] ;
  assign \new_[4795]_  = \\u4_csr_reg[29] ;
  assign \new_[4796]_  = \\u4_csr_reg[2] ;
  assign \new_[4797]_  = ~\\u4_csr_reg[31] ;
  assign \new_[4798]_  = \\u4_csr_reg[3] ;
  assign \new_[4799]_  = \\u4_csr_reg[4] ;
  assign \new_[4800]_  = \\u4_csr_reg[6] ;
  assign \new_[4801]_  = \\u4_csr_reg[7] ;
  assign \new_[4802]_  = \\u4_csr_reg[8] ;
  assign \new_[4803]_  = \new_[14128]_  ? \new_[7549]_  : \new_[5698]_ ;
  assign \new_[4804]_  = ~\\u4_buf0_reg[0] ;
  assign \new_[4805]_  = ~\\u4_buf0_reg[10] ;
  assign \new_[4806]_  = ~\\u4_buf0_reg[11] ;
  assign \new_[4807]_  = ~\\u4_buf0_reg[12] ;
  assign \new_[4808]_  = ~\\u4_buf0_reg[13] ;
  assign \new_[4809]_  = ~\\u4_buf0_reg[15] ;
  assign \new_[4810]_  = ~\\u4_buf0_reg[16] ;
  assign \new_[4811]_  = \\u4_buf0_reg[17] ;
  assign \new_[4812]_  = \\u4_buf0_reg[19] ;
  assign \new_[4813]_  = ~\\u4_buf0_reg[1] ;
  assign \new_[4814]_  = \\u4_buf0_reg[20] ;
  assign \new_[4815]_  = \\u4_buf0_reg[22] ;
  assign \new_[4816]_  = \\u4_buf0_reg[23] ;
  assign \new_[4817]_  = \\u4_buf0_reg[24] ;
  assign \new_[4818]_  = \\u4_buf0_reg[26] ;
  assign \new_[4819]_  = \\u4_buf0_reg[27] ;
  assign \new_[4820]_  = \\u4_buf0_reg[28] ;
  assign \new_[4821]_  = ~\\u4_buf0_reg[2] ;
  assign \new_[4822]_  = ~\\u4_buf0_reg[31] ;
  assign \new_[4823]_  = ~\\u4_buf0_reg[4] ;
  assign \new_[4824]_  = ~\\u4_buf0_reg[5] ;
  assign \new_[4825]_  = ~\\u4_buf0_reg[6] ;
  assign \new_[4826]_  = ~\\u4_buf0_reg[8] ;
  assign \new_[4827]_  = ~\\u4_buf0_reg[9] ;
  assign \new_[4828]_  = ~\\u4_buf1_reg[0] ;
  assign \new_[4829]_  = ~\\u4_buf1_reg[11] ;
  assign \new_[4830]_  = ~\\u4_buf1_reg[12] ;
  assign \new_[4831]_  = ~\\u4_buf1_reg[13] ;
  assign \new_[4832]_  = ~\\u4_buf1_reg[15] ;
  assign \new_[4833]_  = ~\\u4_buf1_reg[16] ;
  assign \new_[4834]_  = \\u4_buf1_reg[17] ;
  assign \new_[4835]_  = \\u4_buf1_reg[19] ;
  assign \new_[4836]_  = ~\\u4_buf1_reg[1] ;
  assign \new_[4837]_  = \\u4_buf1_reg[20] ;
  assign \new_[4838]_  = \\u4_buf1_reg[22] ;
  assign \new_[4839]_  = \\u4_buf1_reg[23] ;
  assign \new_[4840]_  = \\u4_buf1_reg[24] ;
  assign \new_[4841]_  = \\u4_buf1_reg[26] ;
  assign \new_[4842]_  = \\u4_buf1_reg[27] ;
  assign \new_[4843]_  = \\u4_buf1_reg[28] ;
  assign \new_[4844]_  = ~\\u4_buf1_reg[2] ;
  assign \new_[4845]_  = \\u4_buf1_reg[30] ;
  assign \new_[4846]_  = ~\\u4_buf1_reg[31] ;
  assign \new_[4847]_  = ~\\u4_buf1_reg[4] ;
  assign \new_[4848]_  = ~\\u4_buf1_reg[5] ;
  assign \new_[4849]_  = ~\\u4_buf1_reg[6] ;
  assign \new_[4850]_  = ~\\u4_buf1_reg[8] ;
  assign \new_[4851]_  = ~\\u4_buf1_reg[9] ;
  assign \new_[4852]_  = \\u4_csr_reg[0] ;
  assign \new_[4853]_  = \\u4_csr_reg[11] ;
  assign \new_[4854]_  = \\u4_u0_uc_bsel_reg[0] ;
  assign \new_[4855]_  = \\u4_u0_uc_bsel_reg[1] ;
  assign \new_[4856]_  = \\u4_u0_uc_dpd_reg[0] ;
  assign \new_[4857]_  = \\u1_u3_adr_r_reg[11] ;
  assign \new_[4858]_  = \\u1_u3_adr_r_reg[14] ;
  assign \new_[4859]_  = \\u1_u3_adr_r_reg[15] ;
  assign \new_[4860]_  = \\u1_u3_adr_r_reg[6] ;
  assign \new_[4861]_  = \\u1_u3_adr_r_reg[7] ;
  assign \new_[4862]_  = \\u1_u3_adr_r_reg[8] ;
  assign \new_[4863]_  = ~\\u4_buf0_reg[14] ;
  assign \new_[4864]_  = \\u4_buf0_reg[18] ;
  assign \new_[4865]_  = ~\new_[5602]_  | ~\new_[12502]_ ;
  assign \new_[4866]_  = ~\new_[5360]_  | ~\new_[8860]_ ;
  assign \new_[4867]_  = ~\new_[5361]_  | ~\new_[8860]_ ;
  assign \new_[4868]_  = ~\new_[5362]_  | ~\new_[9128]_ ;
  assign \new_[4869]_  = \new_[9601]_  ? \new_[12835]_  : \new_[5629]_ ;
  assign \new_[4870]_  = ~\new_[5413]_  | ~\new_[9128]_ ;
  assign \new_[4871]_  = ~\new_[5563]_  & (~\new_[9137]_  | ~\wb_data_i[28] );
  assign \new_[4872]_  = ~\new_[5565]_  & (~\new_[9137]_  | ~\wb_data_i[31] );
  assign \new_[4873]_  = ~u0_u0_T1_gt_5_0_mS_reg;
  assign \new_[4874]_  = \new_[10131]_  ? \new_[12835]_  : \new_[5633]_ ;
  assign \new_[4875]_  = ~\\u4_csr_reg[16] ;
  assign \new_[4876]_  = ~\new_[7669]_  | ~\new_[5890]_  | ~\new_[6565]_  | ~\new_[6883]_ ;
  assign \new_[4877]_  = ~\new_[7672]_  | ~\new_[5892]_  | ~\new_[6586]_  | ~\new_[6884]_ ;
  assign \new_[4878]_  = ~\new_[5412]_  & ~\new_[9142]_ ;
  assign \new_[4879]_  = ~\new_[5365]_  | ~\new_[9138]_ ;
  assign \new_[4880]_  = ~\new_[5366]_  | ~\new_[9138]_ ;
  assign \new_[4881]_  = ~\new_[5260]_  & (~\new_[9137]_  | ~\wb_data_i[10] );
  assign \new_[4882]_  = u1_u2_rx_data_valid_r_reg;
  assign \new_[4883]_  = \\u1_u3_adr_r_reg[9] ;
  assign \new_[4884]_  = ~\new_[5356]_  & ~\new_[9142]_ ;
  assign \new_[4885]_  = ~\new_[5358]_  & ~\new_[9142]_ ;
  assign \new_[4886]_  = \\u4_u0_uc_dpd_reg[1] ;
  assign \new_[4887]_  = ~\new_[5359]_  & ~\new_[9142]_ ;
  assign \new_[4888]_  = ~\new_[5485]_  | ~\new_[8860]_ ;
  assign n4060 = \new_[5250]_  & \new_[6256]_ ;
  assign \new_[4890]_  = ~\new_[5955]_  | (~\new_[5719]_  & ~\new_[6221]_ );
  assign \new_[4891]_  = ~\new_[5957]_  | (~\new_[14617]_  & ~\new_[6224]_ );
  assign n4045 = \new_[5251]_  & \new_[6256]_ ;
  assign \new_[4893]_  = ~\new_[5592]_  & (~\new_[6652]_  | ~\new_[13669]_ );
  assign \new_[4894]_  = ~\new_[5354]_  | ~\new_[5722]_ ;
  assign \new_[4895]_  = ~\new_[5377]_  & ~\new_[9141]_ ;
  assign \new_[4896]_  = ~\new_[5378]_  & ~\new_[9141]_ ;
  assign \new_[4897]_  = ~\new_[5379]_  & ~\new_[9141]_ ;
  assign \new_[4898]_  = ~\new_[5380]_  & ~\new_[9141]_ ;
  assign \new_[4899]_  = ~\new_[5381]_  & ~\new_[9141]_ ;
  assign \new_[4900]_  = ~\new_[5382]_  & ~\new_[9141]_ ;
  assign \new_[4901]_  = ~\new_[5383]_  & ~\new_[9141]_ ;
  assign \new_[4902]_  = ~\new_[5384]_  & ~\new_[9141]_ ;
  assign \new_[4903]_  = ~\new_[5385]_  & ~\new_[9141]_ ;
  assign \new_[4904]_  = ~\new_[5386]_  & ~\new_[9141]_ ;
  assign \new_[4905]_  = ~\new_[5387]_  & ~\new_[9141]_ ;
  assign \new_[4906]_  = ~\new_[5388]_  & ~\new_[9141]_ ;
  assign \new_[4907]_  = ~\new_[5389]_  & ~\new_[9141]_ ;
  assign \new_[4908]_  = ~\new_[5390]_  & ~\new_[9141]_ ;
  assign \new_[4909]_  = ~\new_[5391]_  & ~\new_[9141]_ ;
  assign \new_[4910]_  = ~\new_[5392]_  & ~\new_[9141]_ ;
  assign \new_[4911]_  = ~\new_[5393]_  & ~\new_[9141]_ ;
  assign \new_[4912]_  = ~\new_[5394]_  & ~\new_[9141]_ ;
  assign \new_[4913]_  = ~\new_[5395]_  & ~\new_[9141]_ ;
  assign \new_[4914]_  = ~\new_[5396]_  & ~\new_[9141]_ ;
  assign \new_[4915]_  = ~\new_[5397]_  & ~\new_[9141]_ ;
  assign \new_[4916]_  = \new_[14047]_  ? \new_[7549]_  : \new_[5741]_ ;
  assign \new_[4917]_  = ~\new_[5368]_  & ~\new_[9142]_ ;
  assign \new_[4918]_  = ~\new_[5369]_  & ~\new_[9142]_ ;
  assign n4095 = \new_[5588]_  & \new_[6256]_ ;
  assign \new_[4920]_  = ~\new_[5371]_  | ~\new_[12502]_ ;
  assign \new_[4921]_  = ~\new_[5372]_  | ~\new_[12502]_ ;
  assign \new_[4922]_  = ~\new_[5374]_  | ~\new_[12502]_ ;
  assign \new_[4923]_  = \\u4_csr_reg[10] ;
  assign \new_[4924]_  = (~\new_[8245]_  | ~\new_[5715]_ ) & (~\new_[5798]_  | ~\new_[10402]_ );
  assign \new_[4925]_  = (~\new_[7561]_  | ~\new_[5715]_ ) & (~\new_[5799]_  | ~\new_[10402]_ );
  assign \new_[4926]_  = \\u1_u1_crc16_reg[11] ;
  assign \new_[4927]_  = \new_[10762]_  ? \new_[12835]_  : \new_[5728]_ ;
  assign \new_[4928]_  = \new_[10311]_  ? \new_[12835]_  : \new_[5736]_ ;
  assign \new_[4929]_  = \new_[10054]_  ? \new_[12835]_  : \new_[5740]_ ;
  assign \new_[4930]_  = ~\\u4_buf1_reg[7] ;
  assign \new_[4931]_  = ~\\u4_buf1_reg[3] ;
  assign \new_[4932]_  = \new_[12205]_  ? \new_[12835]_  : \new_[5735]_ ;
  assign \new_[4933]_  = ~\new_[5398]_  & (~\new_[9137]_  | ~\wb_data_i[4] );
  assign \new_[4934]_  = ~\new_[5399]_  & (~\new_[9137]_  | ~\wb_data_i[5] );
  assign \new_[4935]_  = ~\new_[6432]_  | ~\new_[5947]_  | ~\new_[5917]_  | ~\new_[5916]_ ;
  assign \new_[4936]_  = ~\new_[5400]_  & (~\new_[9137]_  | ~\wb_data_i[7] );
  assign \new_[4937]_  = ~\new_[6424]_  | ~\new_[5948]_  | ~\new_[5920]_  | ~\new_[5919]_ ;
  assign \new_[4938]_  = ~\new_[6462]_  | ~\new_[5949]_  | ~\new_[5694]_  | ~\new_[5922]_ ;
  assign \new_[4939]_  = ~\new_[6466]_  | ~\new_[5951]_  | ~\new_[5926]_  | ~\new_[5925]_ ;
  assign \new_[4940]_  = ~\new_[5289]_  & ~\new_[5706]_ ;
  assign \new_[4941]_  = ~\new_[5318]_  & ~\new_[5707]_ ;
  assign \new_[4942]_  = ~\new_[5320]_  & ~\new_[5708]_ ;
  assign \new_[4943]_  = ~\new_[5322]_  & ~\new_[5709]_ ;
  assign n4215 = (~\new_[6673]_  & ~\new_[8204]_  & ~\new_[13878]_ ) | (~\new_[5915]_  & ~\new_[10503]_  & ~\new_[13878]_ );
  assign \new_[4945]_  = \new_[13805]_  ? \new_[7857]_  : \new_[5896]_ ;
  assign n4125 = (~\new_[9653]_  & ~\new_[6171]_  & ~\new_[13963]_ ) | (~\new_[13963]_  & ~\new_[8558]_  & ~\new_[6171]_ );
  assign \new_[4947]_  = (~\new_[7623]_  | ~\new_[5917]_ ) & (~\new_[6764]_  | ~\new_[5917]_ );
  assign \new_[4948]_  = (~\new_[6765]_  | ~\new_[5920]_ ) & (~\new_[7640]_  | ~\new_[5920]_ );
  assign \new_[4949]_  = (~\new_[7637]_  | ~\new_[5926]_ ) & (~\new_[6771]_  | ~\new_[5926]_ );
  assign \new_[4950]_  = ~\\u1_u0_d1_reg[0] ;
  assign \wb_data_o[25]  = \\u5_wb_data_o_reg[25] ;
  assign \new_[4952]_  = \\u4_dout_reg[0] ;
  assign \new_[4953]_  = ~\\u1_u0_d1_reg[4] ;
  assign \new_[4954]_  = \\u4_dout_reg[2] ;
  assign \new_[4955]_  = \\u4_dout_reg[3] ;
  assign \new_[4956]_  = ~\\u1_u0_d0_reg[4] ;
  assign \wb_data_o[26]  = \\u5_wb_data_o_reg[26] ;
  assign \new_[4958]_  = ~\new_[5718]_  | (~\new_[2932]_  & ~\new_[2870]_ );
  assign \new_[4959]_  = ~\new_[5797]_  & ~\new_[10056]_ ;
  assign \new_[4960]_  = ~\\u1_u0_d0_reg[1] ;
  assign \new_[4961]_  = ~\\u1_u0_d0_reg[3] ;
  assign \new_[4962]_  = ~\new_[5623]_  & ~\new_[6227]_ ;
  assign \new_[4963]_  = ~\new_[5789]_  | (~\new_[8677]_  & ~\new_[12840]_ );
  assign \new_[4964]_  = ~\new_[5703]_  & (~\new_[6555]_  | ~\new_[13722]_ );
  assign \new_[4965]_  = ~\new_[5704]_  & (~\new_[6555]_  | ~\new_[13976]_ );
  assign \new_[4966]_  = \\u4_u1_int_stat_reg[4] ;
  assign \new_[4967]_  = \new_[5716]_  & \new_[6175]_ ;
  assign \new_[4968]_  = ~\new_[5705]_  & (~\new_[6555]_  | ~\new_[13955]_ );
  assign \new_[4969]_  = ~\new_[5627]_  | ~\new_[5985]_ ;
  assign \new_[4970]_  = \\u4_u3_int_stat_reg[4] ;
  assign \new_[4971]_  = \new_[5723]_  | \new_[10395]_ ;
  assign \new_[4972]_  = ~\new_[9375]_  | ~\new_[5715]_  | ~\new_[2373]_ ;
  assign \new_[4973]_  = ~\new_[5725]_  | ~\new_[12835]_ ;
  assign \new_[4974]_  = ~\new_[5729]_  | ~\new_[8909]_ ;
  assign \new_[4975]_  = ~\new_[5730]_  | ~\new_[8911]_ ;
  assign \new_[4976]_  = ~\new_[5731]_  | ~\new_[8909]_ ;
  assign \new_[4977]_  = ~\new_[5732]_  | ~\new_[8909]_ ;
  assign \new_[4978]_  = ~\new_[5733]_  | ~\new_[8909]_ ;
  assign \new_[4979]_  = ~\new_[5734]_  | ~\new_[8910]_ ;
  assign \new_[4980]_  = ~\new_[5727]_  | ~\new_[12835]_ ;
  assign \new_[4981]_  = ~\new_[5737]_  | ~\new_[12835]_ ;
  assign \new_[4982]_  = ~\new_[5738]_  | ~\new_[12835]_ ;
  assign \new_[4983]_  = ~\new_[5739]_  | ~\new_[12835]_ ;
  assign \new_[4984]_  = \new_[14258]_  ? \new_[7307]_  : \new_[5991]_ ;
  assign \new_[4985]_  = \new_[14016]_  ? \new_[7307]_  : \new_[5992]_ ;
  assign \new_[4986]_  = \new_[3283]_  ? \new_[7455]_  : \new_[5971]_ ;
  assign \new_[4987]_  = \new_[3308]_  ? \new_[6031]_  : \new_[5972]_ ;
  assign \new_[4988]_  = \new_[3309]_  ? \new_[6476]_  : \new_[5973]_ ;
  assign \new_[4989]_  = \new_[3282]_  ? \new_[6778]_  : \new_[5976]_ ;
  assign \new_[4990]_  = ~u4_crc5_err_r_reg;
  assign \new_[4991]_  = ~\new_[5711]_  & (~\new_[6555]_  | ~\new_[14202]_ );
  assign \new_[4992]_  = ~\new_[5712]_  & (~\new_[6555]_  | ~\new_[13784]_ );
  assign \new_[4993]_  = \new_[3480]_  ? \new_[6031]_  : \new_[9921]_ ;
  assign \new_[4994]_  = \new_[3316]_  ? \new_[6031]_  : \new_[9071]_ ;
  assign \new_[4995]_  = \new_[3315]_  ? \new_[6031]_  : \new_[8710]_ ;
  assign \new_[4996]_  = \new_[3429]_  ? \new_[6031]_  : \new_[9384]_ ;
  assign \new_[4997]_  = \new_[3317]_  ? \new_[6031]_  : \new_[8711]_ ;
  assign \new_[4998]_  = \new_[3478]_  ? \new_[6031]_  : \new_[8712]_ ;
  assign \new_[4999]_  = \new_[14259]_  ? \new_[7857]_  : \new_[5996]_ ;
  assign \new_[5000]_  = ~\new_[5770]_  & (~\new_[6555]_  | ~\new_[13596]_ );
  assign \new_[5001]_  = (~\new_[6652]_  | ~\new_[13562]_ ) & (~\new_[6101]_  | ~\new_[2266]_ );
  assign \new_[5002]_  = (~\new_[6652]_  | ~\new_[13979]_ ) & (~\new_[6101]_  | ~\new_[2047]_ );
  assign \new_[5003]_  = (~\new_[6652]_  | ~\new_[13909]_ ) & (~\new_[6101]_  | ~\new_[2048]_ );
  assign \new_[5004]_  = (~\new_[6084]_  | ~\new_[13671]_ ) & (~\new_[6101]_  | ~\new_[5421]_ );
  assign \new_[5005]_  = (~\new_[6084]_  | ~\new_[13929]_ ) & (~\new_[6101]_  | ~\new_[3102]_ );
  assign \new_[5006]_  = (~\new_[6084]_  | ~\new_[13998]_ ) & (~\new_[6101]_  | ~\new_[3173]_ );
  assign \new_[5007]_  = (~\new_[6084]_  | ~\new_[13773]_ ) & (~\new_[6101]_  | ~\new_[2178]_ );
  assign \new_[5008]_  = (~\new_[6084]_  | ~\new_[14183]_ ) & (~\new_[6101]_  | ~\new_[3034]_ );
  assign \new_[5009]_  = (~\new_[6084]_  | ~\new_[13869]_ ) & (~\new_[6101]_  | ~\new_[3021]_ );
  assign \new_[5010]_  = (~\new_[6084]_  | ~\new_[13890]_ ) & (~\new_[6101]_  | ~\new_[9037]_ );
  assign \new_[5011]_  = (~\new_[6084]_  | ~\new_[14065]_ ) & (~\new_[6101]_  | ~\new_[2928]_ );
  assign \new_[5012]_  = (~\new_[6652]_  | ~\new_[13934]_ ) & (~\new_[6101]_  | ~\new_[2856]_ );
  assign \new_[5013]_  = (~\new_[6652]_  | ~\new_[13762]_ ) & (~\new_[6101]_  | ~\new_[2638]_ );
  assign \new_[5014]_  = (~\new_[6084]_  | ~\new_[13853]_ ) & (~\new_[6101]_  | ~\new_[2639]_ );
  assign \new_[5015]_  = (~\new_[6084]_  | ~\new_[13838]_ ) & (~\new_[6101]_  | ~\new_[2547]_ );
  assign \new_[5016]_  = (~\new_[6652]_  | ~\new_[13935]_ ) & (~\new_[6101]_  | ~\new_[2735]_ );
  assign \new_[5017]_  = (~\new_[6652]_  | ~\new_[14175]_ ) & (~\new_[6101]_  | ~\new_[2177]_ );
  assign \new_[5018]_  = (~\new_[6084]_  | ~\new_[14122]_ ) & (~\new_[6101]_  | ~\new_[2265]_ );
  assign \new_[5019]_  = (~\new_[6084]_  | ~\new_[14014]_ ) & (~\new_[6101]_  | ~\new_[2136]_ );
  assign \new_[5020]_  = (~\new_[6652]_  | ~\new_[13991]_ ) & (~\new_[6101]_  | ~\new_[2075]_ );
  assign \new_[5021]_  = (~\new_[6084]_  | ~\new_[14168]_ ) & (~\new_[6101]_  | ~\new_[2062]_ );
  assign \new_[5022]_  = \new_[5624]_  | n4965;
  assign \new_[5023]_  = ~\new_[5744]_  | ~\new_[12835]_ ;
  assign \new_[5024]_  = ~\new_[5713]_  & (~\new_[6555]_  | ~\new_[14165]_ );
  assign \new_[5025]_  = \new_[3462]_  ? \new_[6031]_  : \new_[8181]_ ;
  assign \new_[5026]_  = \new_[3428]_  ? \new_[6031]_  : \new_[7460]_ ;
  assign \new_[5027]_  = \new_[13783]_  ? \new_[7857]_  : \new_[6068]_ ;
  assign \new_[5028]_  = \\u1_u3_next_dpid_reg[0] ;
  assign \new_[5029]_  = ~\new_[5747]_  & ~\new_[6221]_ ;
  assign \new_[5030]_  = \new_[5928]_  ? \new_[7939]_  : \new_[7429]_ ;
  assign \new_[5031]_  = ~\new_[6692]_  | (~\new_[7939]_  & ~\new_[5928]_ );
  assign \new_[5032]_  = ~\new_[5791]_  | ~\new_[6059]_ ;
  assign \new_[5033]_  = \new_[3337]_  ? \new_[6031]_  : \new_[12032]_ ;
  assign \new_[5034]_  = \new_[6304]_  ? \new_[8608]_  : \new_[6034]_ ;
  assign \new_[5035]_  = \new_[14125]_  ? \new_[8608]_  : \new_[6035]_ ;
  assign \new_[5036]_  = ~\new_[5793]_  | ~\new_[12835]_ ;
  assign n4135 = ~\new_[5801]_  | ~\new_[8661]_ ;
  assign n4110 = ~\new_[5802]_  | ~\new_[8661]_ ;
  assign \new_[5039]_  = \new_[13700]_  ? \new_[7307]_  : \new_[6038]_ ;
  assign \new_[5040]_  = \new_[14080]_  ? \new_[7307]_  : \new_[6039]_ ;
  assign \new_[5041]_  = \new_[14054]_  ? \new_[7307]_  : \new_[6041]_ ;
  assign \new_[5042]_  = ~\new_[7570]_  & (~\new_[7772]_  | ~\new_[6073]_ );
  assign \new_[5043]_  = \new_[6232]_  ? \new_[7307]_  : \new_[6042]_ ;
  assign \new_[5044]_  = ~\new_[10667]_  & (~\new_[9815]_  | ~\new_[6075]_ );
  assign \new_[5045]_  = \new_[6324]_  ? \new_[7307]_  : \new_[6044]_ ;
  assign \new_[5046]_  = \new_[14095]_  ? \new_[7307]_  : \new_[6045]_ ;
  assign \new_[5047]_  = ~\new_[5856]_  | (~\new_[9163]_  & ~\new_[12840]_ );
  assign \new_[5048]_  = \new_[3503]_  ? \new_[6031]_  : \new_[10766]_ ;
  assign \new_[5049]_  = \new_[3504]_  ? \new_[6031]_  : \new_[10570]_ ;
  assign \new_[5050]_  = \new_[3505]_  ? \new_[6031]_  : \new_[9970]_ ;
  assign \new_[5051]_  = \new_[3339]_  ? \new_[6031]_  : \new_[12897]_ ;
  assign \new_[5052]_  = \new_[3340]_  ? \new_[6031]_  : \new_[11453]_ ;
  assign \new_[5053]_  = \new_[3341]_  ? \new_[6031]_  : \new_[9971]_ ;
  assign \new_[5054]_  = \new_[3342]_  ? \new_[6031]_  : \new_[9707]_ ;
  assign \new_[5055]_  = \new_[3506]_  ? \new_[6031]_  : \new_[9116]_ ;
  assign \new_[5056]_  = ~\new_[5767]_  & (~\new_[9852]_  | ~\new_[9313]_ );
  assign \new_[5057]_  = \new_[14243]_  ? \new_[7857]_  : \new_[6056]_ ;
  assign \new_[5058]_  = \new_[13797]_  ? \new_[7857]_  : \new_[6051]_ ;
  assign \new_[5059]_  = \new_[14002]_  ? \new_[7857]_  : \new_[6057]_ ;
  assign \new_[5060]_  = \new_[14101]_  ? \new_[7857]_  : \new_[6052]_ ;
  assign \new_[5061]_  = \new_[13938]_  ? \new_[7857]_  : \new_[6050]_ ;
  assign \new_[5062]_  = \new_[14214]_  ? \new_[7857]_  : \new_[6053]_ ;
  assign \new_[5063]_  = \new_[6365]_  ? \new_[7857]_  : \new_[6054]_ ;
  assign \new_[5064]_  = \new_[14150]_  ? \new_[7857]_  : \new_[6049]_ ;
  assign \new_[5065]_  = \new_[6366]_  ? \new_[7857]_  : \new_[6048]_ ;
  assign \new_[5066]_  = \new_[6368]_  ? \new_[7857]_  : \new_[6046]_ ;
  assign \new_[5067]_  = \new_[6369]_  ? \new_[7857]_  : \new_[6043]_ ;
  assign \new_[5068]_  = \new_[6370]_  ? \new_[7857]_  : \new_[6040]_ ;
  assign \new_[5069]_  = \new_[6461]_  ? \new_[7857]_  : \new_[6055]_ ;
  assign \new_[5070]_  = \new_[6556]_  ? \new_[7857]_  : \new_[6036]_ ;
  assign \new_[5071]_  = \new_[14263]_  ? \new_[7857]_  : \new_[6047]_ ;
  assign \new_[5072]_  = ~\new_[5803]_  & (~\new_[6555]_  | ~\new_[13948]_ );
  assign \new_[5073]_  = \new_[3466]_  ? \new_[6031]_  : \new_[6855]_ ;
  assign \new_[5074]_  = \new_[3313]_  ? \new_[6031]_  : \new_[7304]_ ;
  assign \new_[5075]_  = ~\\u1_u3_adr_r_reg[0] ;
  assign \new_[5076]_  = u4_u1_dma_in_buf_sz1_reg;
  assign \new_[5077]_  = u4_u0_dma_in_buf_sz1_reg;
  assign \new_[5078]_  = u4_u3_dma_in_buf_sz1_reg;
  assign \new_[5079]_  = ~u4_u2_dma_in_buf_sz1_reg;
  assign \new_[5080]_  = ~\new_[14539]_  | ~n5230;
  assign \new_[5081]_  = \new_[8222]_  | n4205;
  assign \new_[5082]_  = \new_[14788]_  | n5200;
  assign \new_[5083]_  = \new_[14787]_  & n5200;
  assign \new_[5084]_  = \new_[7845]_  & n4205;
  assign \new_[5085]_  = ~\new_[14422]_  & ~n5225;
  assign \new_[5086]_  = \new_[8602]_  & n4210;
  assign \new_[5087]_  = ~\new_[7846]_  | ~n5225;
  assign \new_[5088]_  = ~\new_[8603]_  | ~\new_[5784]_ ;
  assign \new_[5089]_  = ~\new_[8601]_  | ~\new_[5783]_ ;
  assign \new_[5090]_  = ~\new_[8600]_  | ~\new_[5785]_ ;
  assign \new_[5091]_  = \new_[8224]_  & \new_[5782]_ ;
  assign \new_[5092]_  = ~\new_[8224]_  & ~\new_[5782]_ ;
  assign \new_[5093]_  = ~\new_[8601]_  & ~\new_[5783]_ ;
  assign \new_[5094]_  = ~\new_[8603]_  & ~\new_[5784]_ ;
  assign \new_[5095]_  = ~\new_[8600]_  & ~\new_[5785]_ ;
  assign \new_[5096]_  = \new_[14507]_  | n4195;
  assign \new_[5097]_  = \new_[14507]_  & n4195;
  assign \new_[5098]_  = \new_[14270]_  | \new_[5787]_ ;
  assign \new_[5099]_  = ~\new_[14270]_  | ~\new_[5787]_ ;
  assign \new_[5100]_  = \new_[14276]_  | \new_[5774]_ ;
  assign \new_[5101]_  = ~\new_[14276]_  | ~\new_[5774]_ ;
  assign \new_[5102]_  = ~\new_[14275]_  | ~n4200;
  assign \new_[5103]_  = ~\new_[14275]_  & ~n4200;
  assign \new_[5104]_  = \new_[14423]_  | n4210;
  assign \new_[5105]_  = \new_[14539]_  | n5230;
  assign \new_[5106]_  = ~\new_[5768]_  & (~\new_[6555]_  | ~\new_[14212]_ );
  assign \new_[5107]_  = ~\new_[5769]_  & (~\new_[7284]_  | ~\new_[13590]_ );
  assign TermSel_pad_o = u0_u0_TermSel_reg;
  assign \new_[5109]_  = \\u4_int_srcb_reg[5] ;
  assign \wb_data_o[4]  = \\u5_wb_data_o_reg[4] ;
  assign \new_[5111]_  = \\u4_u2_int_stat_reg[4] ;
  assign \new_[5112]_  = \\u4_u0_int_stat_reg[4] ;
  assign \wb_data_o[16]  = \\u5_wb_data_o_reg[16] ;
  assign \wb_data_o[24]  = \\u5_wb_data_o_reg[24] ;
  assign \wb_data_o[28]  = \\u5_wb_data_o_reg[28] ;
  assign \wb_data_o[21]  = \\u5_wb_data_o_reg[21] ;
  assign \wb_data_o[20]  = \\u5_wb_data_o_reg[20] ;
  assign \wb_data_o[19]  = \\u5_wb_data_o_reg[19] ;
  assign \wb_data_o[6]  = \\u5_wb_data_o_reg[6] ;
  assign \wb_data_o[5]  = \\u5_wb_data_o_reg[5] ;
  assign \wb_data_o[18]  = \\u5_wb_data_o_reg[18] ;
  assign \wb_data_o[17]  = \\u5_wb_data_o_reg[17] ;
  assign \new_[5123]_  = \\u4_int_srcb_reg[4] ;
  assign \new_[5124]_  = \\u0_u0_state_reg[1] ;
  assign \new_[5125]_  = ~u1_u0_rxv1_reg;
  assign \new_[5126]_  = ~\\u1_u0_d0_reg[0] ;
  assign \new_[5127]_  = ~\\u0_u0_chirp_cnt_reg[1] ;
  assign \new_[5128]_  = ~\\u1_u0_d0_reg[2] ;
  assign \new_[5129]_  = ~\\u0_u0_chirp_cnt_reg[2] ;
  assign \new_[5130]_  = ~\\u1_u0_d0_reg[5] ;
  assign \new_[5131]_  = ~\\u1_u0_d0_reg[6] ;
  assign \new_[5132]_  = ~\\u1_u0_d0_reg[7] ;
  assign \new_[5133]_  = ~\\u1_u0_d1_reg[1] ;
  assign \new_[5134]_  = ~\\u1_u0_d1_reg[2] ;
  assign \new_[5135]_  = ~\\u1_u0_d1_reg[3] ;
  assign \new_[5136]_  = ~\\u1_u0_d1_reg[5] ;
  assign \new_[5137]_  = ~\\u1_u0_d1_reg[6] ;
  assign \new_[5138]_  = ~\\u1_u0_d1_reg[7] ;
  assign \new_[5139]_  = ~\\u1_u0_d2_reg[1] ;
  assign \new_[5140]_  = ~\\u1_u0_d2_reg[2] ;
  assign \new_[5141]_  = ~\\u1_u0_d2_reg[3] ;
  assign \new_[5142]_  = ~\\u1_u0_d2_reg[5] ;
  assign \new_[5143]_  = ~\\u1_u0_d2_reg[6] ;
  assign \new_[5144]_  = ~\\u1_u0_d2_reg[7] ;
  assign \new_[5145]_  = \\u0_u0_state_reg[12] ;
  assign \new_[5146]_  = \new_[14107]_  ? \new_[7857]_  : \new_[5897]_ ;
  assign \new_[5147]_  = ~\new_[13162]_  | ~\new_[5823]_  | ~\new_[4161]_ ;
  assign \new_[5148]_  = \\u4_u1_uc_bsel_reg[0] ;
  assign \new_[5149]_  = \\u4_u1_uc_dpd_reg[0] ;
  assign \new_[5150]_  = \new_[13787]_  ? \new_[7857]_  : \new_[5932]_ ;
  assign \new_[5151]_  = \\u1_u3_adr_r_reg[2] ;
  assign \new_[5152]_  = \new_[14076]_  ? \new_[7857]_  : \new_[5898]_ ;
  assign \new_[5153]_  = ~\new_[4161]_  | ~\new_[11079]_  | ~\new_[6621]_ ;
  assign \new_[5154]_  = ~\new_[5800]_  | (~\new_[6522]_  & ~\new_[12798]_ );
  assign \new_[5155]_  = ~\new_[5883]_  | ~\new_[12835]_ ;
  assign \new_[5156]_  = ~\new_[3781]_  | ~\new_[10852]_  | ~\new_[6621]_ ;
  assign n4140 = ~\new_[6179]_  | ~\new_[5847]_ ;
  assign \new_[5158]_  = ~\new_[13457]_  | ~\new_[10852]_  | ~\new_[6621]_ ;
  assign \new_[5159]_  = ~\new_[5855]_  | (~\new_[9530]_  & ~\new_[12840]_ );
  assign \new_[5160]_  = ~\new_[5857]_  | (~\new_[10687]_  & ~\new_[12840]_ );
  assign \new_[5161]_  = \new_[3310]_  ? \new_[6031]_  : \new_[6902]_ ;
  assign \new_[5162]_  = ~\new_[5824]_  & (~\new_[9137]_  | ~\wb_data_i[0] );
  assign \new_[5163]_  = ~\new_[5825]_  & (~\new_[9137]_  | ~\wb_data_i[12] );
  assign \new_[5164]_  = ~\new_[5826]_  & (~\new_[9137]_  | ~\wb_data_i[16] );
  assign \new_[5165]_  = ~\new_[5827]_  & (~\new_[9137]_  | ~\wb_data_i[17] );
  assign \new_[5166]_  = ~\new_[5828]_  & (~\new_[9137]_  | ~\wb_data_i[18] );
  assign \new_[5167]_  = ~\new_[5829]_  & (~\new_[9137]_  | ~\wb_data_i[19] );
  assign \new_[5168]_  = ~\new_[5830]_  & (~\new_[9137]_  | ~\wb_data_i[1] );
  assign \new_[5169]_  = ~\new_[5831]_  & (~\new_[9137]_  | ~\wb_data_i[20] );
  assign \new_[5170]_  = ~\new_[5832]_  & (~\new_[9137]_  | ~\wb_data_i[21] );
  assign \new_[5171]_  = ~\new_[5833]_  & (~\new_[9137]_  | ~\wb_data_i[22] );
  assign \new_[5172]_  = ~\new_[5834]_  & (~\new_[9137]_  | ~\wb_data_i[23] );
  assign \new_[5173]_  = ~\new_[5835]_  & (~\new_[9137]_  | ~\wb_data_i[24] );
  assign \new_[5174]_  = \\u4_u1_uc_bsel_reg[1] ;
  assign \new_[5175]_  = ~\new_[5836]_  & (~\new_[9137]_  | ~\wb_data_i[25] );
  assign \new_[5176]_  = ~\new_[5837]_  & (~\new_[9137]_  | ~\wb_data_i[26] );
  assign \new_[5177]_  = ~\new_[5838]_  & (~\new_[9137]_  | ~\wb_data_i[27] );
  assign \new_[5178]_  = ~\new_[5839]_  & (~\new_[9137]_  | ~\wb_data_i[29] );
  assign \new_[5179]_  = ~\new_[5840]_  & (~\new_[9137]_  | ~\wb_data_i[2] );
  assign \new_[5180]_  = ~\new_[5842]_  & (~\new_[9137]_  | ~\wb_data_i[30] );
  assign \new_[5181]_  = ~\new_[5843]_  & (~\new_[9137]_  | ~\wb_data_i[3] );
  assign \new_[5182]_  = ~\new_[5844]_  & (~\new_[9137]_  | ~\wb_data_i[8] );
  assign \new_[5183]_  = ~\new_[5845]_  & (~\new_[9137]_  | ~\wb_data_i[9] );
  assign \new_[5184]_  = ~\new_[6080]_  | ~\new_[8314]_  | ~\new_[7389]_ ;
  assign \new_[5185]_  = \\u4_u1_uc_dpd_reg[1] ;
  assign \new_[5186]_  = ~\new_[5851]_  | (~\new_[7548]_  & ~\new_[11733]_ );
  assign \new_[5187]_  = ~\new_[5852]_  | (~\new_[7548]_  & ~\new_[11577]_ );
  assign n4120 = ~\new_[5902]_  | ~\new_[5822]_ ;
  assign \new_[5189]_  = ~\new_[5625]_  | ~\new_[8910]_ ;
  assign \new_[5190]_  = ~\new_[5626]_  | ~\new_[8909]_ ;
  assign \new_[5191]_  = ~\new_[5956]_  | (~\new_[5955]_  & ~\new_[6705]_ );
  assign \new_[5192]_  = ~\new_[5882]_  & (~\new_[6555]_  | ~\new_[13726]_ );
  assign \new_[5193]_  = ~\new_[5674]_  & ~\new_[9142]_ ;
  assign \new_[5194]_  = ~\new_[5675]_  & ~\new_[9142]_ ;
  assign \new_[5195]_  = ~\new_[5676]_  & ~\new_[9142]_ ;
  assign \new_[5196]_  = ~\new_[5693]_  & ~\new_[9142]_ ;
  assign \new_[5197]_  = ~\new_[5677]_  & ~\new_[9142]_ ;
  assign \new_[5198]_  = ~\new_[5678]_  & ~\new_[9142]_ ;
  assign \new_[5199]_  = ~\new_[5679]_  & ~\new_[9142]_ ;
  assign \new_[5200]_  = ~\new_[5680]_  & ~\new_[9142]_ ;
  assign \new_[5201]_  = ~\new_[5681]_  & ~\new_[9142]_ ;
  assign \new_[5202]_  = ~\new_[5682]_  & ~\new_[9142]_ ;
  assign \new_[5203]_  = ~\new_[5683]_  & ~\new_[9142]_ ;
  assign \new_[5204]_  = ~\new_[5684]_  & ~\new_[9142]_ ;
  assign \new_[5205]_  = ~\new_[5685]_  & ~\new_[9142]_ ;
  assign \new_[5206]_  = ~\new_[5686]_  & ~\new_[9142]_ ;
  assign \new_[5207]_  = ~\new_[5687]_  & ~\new_[9142]_ ;
  assign \new_[5208]_  = ~\new_[5688]_  & ~\new_[9142]_ ;
  assign \new_[5209]_  = ~\new_[5673]_  & ~\new_[9142]_ ;
  assign \new_[5210]_  = ~\new_[5689]_  & ~\new_[9142]_ ;
  assign \new_[5211]_  = ~\new_[5690]_  & ~\new_[9142]_ ;
  assign \new_[5212]_  = ~\new_[5691]_  & ~\new_[9142]_ ;
  assign \new_[5213]_  = ~\new_[5692]_  & ~\new_[9142]_ ;
  assign \new_[5214]_  = \new_[14246]_  ? \new_[7857]_  : \new_[5969]_ ;
  assign n4145 = ~\new_[5672]_  | ~\new_[8661]_ ;
  assign n4150 = ~\new_[5635]_  | ~\new_[8661]_ ;
  assign n4115 = ~\new_[5636]_  | ~\new_[8661]_ ;
  assign n4155 = ~\new_[5637]_  | ~\new_[8661]_ ;
  assign n4220 = ~\new_[5638]_  | ~\new_[8661]_ ;
  assign n4160 = ~\new_[5639]_  | ~\new_[8661]_ ;
  assign n4230 = ~\new_[5640]_  | ~\new_[8661]_ ;
  assign n4165 = ~\new_[5641]_  | ~\new_[8661]_ ;
  assign n4170 = ~\new_[5642]_  | ~\new_[8661]_ ;
  assign \new_[5224]_  = ~\new_[5788]_  & (~\new_[11104]_  | ~\new_[9510]_ );
  assign n4175 = ~\new_[5643]_  | ~\new_[8661]_ ;
  assign n4225 = ~\new_[5644]_  | ~\new_[8661]_ ;
  assign n4180 = ~\new_[5645]_  | ~\new_[8661]_ ;
  assign n4185 = ~\new_[5646]_  | ~\new_[8661]_ ;
  assign n4190 = ~\new_[5647]_  | ~\new_[8661]_ ;
  assign \new_[5230]_  = ~\new_[5630]_  | ~\new_[12835]_ ;
  assign \new_[5231]_  = ~\new_[5631]_  | ~\new_[12835]_ ;
  assign \new_[5232]_  = ~\new_[5628]_  | ~\new_[12835]_ ;
  assign \new_[5233]_  = ~\new_[13348]_  | ~\new_[6119]_  | ~\new_[4161]_ ;
  assign \new_[5234]_  = ~\new_[4290]_  | ~\new_[6119]_  | ~\new_[14127]_ ;
  assign \new_[5235]_  = ~\new_[5612]_  | (~\new_[4095]_  & ~\new_[12840]_ );
  assign \new_[5236]_  = ~\new_[5619]_  | (~\new_[4098]_  & ~\new_[12840]_ );
  assign \new_[5237]_  = ~\new_[5620]_  | (~\new_[11636]_  & ~\new_[12840]_ );
  assign \new_[5238]_  = ~\new_[5621]_  | (~\new_[11371]_  & ~\new_[12840]_ );
  assign \new_[5239]_  = ~\new_[5622]_  | (~\new_[10659]_  & ~\new_[12840]_ );
  assign \new_[5240]_  = \new_[11756]_  ? \new_[5928]_  : \new_[11747]_ ;
  assign \new_[5241]_  = \new_[11929]_  ? \new_[5928]_  : \new_[11707]_ ;
  assign \new_[5242]_  = ~\\u1_u0_d2_reg[0] ;
  assign \new_[5243]_  = ~\\u1_u0_d2_reg[4] ;
  assign \new_[5244]_  = \new_[3477]_  ? \new_[6031]_  : \new_[7685]_ ;
  assign \new_[5245]_  = \new_[3476]_  ? \new_[6031]_  : \new_[7912]_ ;
  assign \new_[5246]_  = \new_[3312]_  ? \new_[6031]_  : \new_[7403]_ ;
  assign n4130 = \new_[8417]_  ^ \new_[5986]_ ;
  assign \new_[5248]_  = \\u1_u3_adr_r_reg[5] ;
  assign \new_[5249]_  = \\u1_u3_adr_r_reg[1] ;
  assign \new_[5250]_  = \new_[9172]_  ? \new_[12840]_  : \new_[6161]_ ;
  assign \new_[5251]_  = \new_[9725]_  ? \new_[12840]_  : \new_[6162]_ ;
  assign n4480 = ~\new_[6314]_  | ~\new_[7790]_  | ~\new_[6788]_ ;
  assign n4865 = ~\new_[6321]_  | ~\new_[7505]_  | ~\new_[7209]_ ;
  assign n4775 = ~\new_[6453]_  | ~\new_[7515]_  | ~\new_[7229]_ ;
  assign n4485 = ~\new_[6333]_  | ~\new_[7809]_  | ~\new_[7210]_ ;
  assign n4250 = ~\new_[6349]_  | ~\new_[7802]_  | ~\new_[6791]_ ;
  assign n4490 = ~\new_[6356]_  | ~\new_[7792]_  | ~\new_[7211]_ ;
  assign n4400 = ~\new_[6360]_  | ~\new_[7506]_  | ~\new_[7234]_ ;
  assign n4495 = ~\new_[6395]_  | ~\new_[7487]_  | ~\new_[7221]_ ;
  assign \new_[5260]_  = ~\new_[5967]_  & ~\new_[9137]_ ;
  assign n4500 = ~\new_[6372]_  | ~\new_[7497]_  | ~\new_[6806]_ ;
  assign n4505 = ~\new_[6376]_  | ~\new_[7793]_  | ~\new_[6792]_ ;
  assign n4355 = ~\new_[6529]_  | ~\new_[7794]_  | ~\new_[6793]_ ;
  assign n4510 = ~\new_[6164]_  | ~\new_[7488]_  | ~\new_[7214]_ ;
  assign n4515 = ~\new_[6381]_  | ~\new_[7489]_  | ~\new_[7251]_ ;
  assign n4520 = ~\new_[6596]_  | ~\new_[7808]_  | ~\new_[6794]_ ;
  assign n4335 = ~\new_[6382]_  | ~\new_[7795]_  | ~\new_[6807]_ ;
  assign n4525 = ~\new_[6388]_  | ~\new_[7490]_  | ~\new_[7215]_ ;
  assign n4530 = ~\new_[6389]_  | ~\new_[7491]_  | ~\new_[6795]_ ;
  assign n4535 = ~\new_[6390]_  | ~\new_[7796]_  | ~\new_[6810]_ ;
  assign n4275 = ~\new_[6399]_  | ~\new_[7807]_  | ~\new_[6799]_ ;
  assign n4540 = ~\new_[6455]_  | ~\new_[7511]_  | ~\new_[6812]_ ;
  assign n4545 = ~\new_[6391]_  | ~\new_[7806]_  | ~\new_[6797]_ ;
  assign n4550 = ~\new_[6392]_  | ~\new_[7510]_  | ~\new_[6805]_ ;
  assign n4295 = ~\new_[6393]_  | ~\new_[7797]_  | ~\new_[6796]_ ;
  assign n4735 = ~\new_[6445]_  | ~\new_[7810]_  | ~\new_[6813]_ ;
  assign n4555 = ~\new_[6400]_  | ~\new_[7516]_  | ~\new_[7239]_ ;
  assign n4560 = ~\new_[6401]_  | ~\new_[7517]_  | ~\new_[7240]_ ;
  assign n4565 = ~\new_[6402]_  | ~\new_[7815]_  | ~\new_[7241]_ ;
  assign n4570 = ~\new_[6403]_  | ~\new_[7518]_  | ~\new_[7220]_ ;
  assign n4575 = ~\new_[6404]_  | ~\new_[7519]_  | ~\new_[7242]_ ;
  assign n4850 = ~\new_[6405]_  | ~\new_[7520]_  | ~\new_[7244]_ ;
  assign n4580 = ~\new_[6406]_  | ~\new_[7493]_  | ~\new_[7245]_ ;
  assign n4585 = ~\new_[6208]_  | ~\new_[7507]_  | ~\new_[6798]_ ;
  assign n4590 = ~\new_[6407]_  | ~\new_[7823]_  | ~\new_[6804]_ ;
  assign n4855 = ~\new_[6408]_  | ~\new_[7501]_  | ~\new_[6818]_ ;
  assign n4595 = ~\new_[6397]_  | ~\new_[7821]_  | ~\new_[6789]_ ;
  assign n4780 = ~\new_[6394]_  | ~\new_[7814]_  | ~\new_[7223]_ ;
  assign \new_[5289]_  = \\u4_u3_dma_out_left_reg[10] ;
  assign n4600 = ~\new_[6409]_  | ~\new_[7527]_  | ~\new_[7217]_ ;
  assign n4605 = ~\new_[6410]_  | ~\new_[7822]_  | ~\new_[6801]_ ;
  assign n4350 = ~\new_[6411]_  | ~\new_[7816]_  | ~\new_[6817]_ ;
  assign n4610 = ~\new_[6412]_  | ~\new_[7817]_  | ~\new_[6824]_ ;
  assign n4615 = ~\new_[6413]_  | ~\new_[7818]_  | ~\new_[6814]_ ;
  assign n4620 = ~\new_[6398]_  | ~\new_[7811]_  | ~\new_[6811]_ ;
  assign n4360 = ~\new_[6414]_  | ~\new_[7813]_  | ~\new_[6815]_ ;
  assign n4625 = ~\new_[6415]_  | ~\new_[7803]_  | ~\new_[6816]_ ;
  assign n4630 = ~\new_[6416]_  | ~\new_[7500]_  | ~\new_[7222]_ ;
  assign n4635 = ~\new_[6417]_  | ~\new_[7494]_  | ~\new_[7219]_ ;
  assign n4310 = ~\new_[6418]_  | ~\new_[7825]_  | ~\new_[7246]_ ;
  assign n4640 = ~\new_[6419]_  | ~\new_[7820]_  | ~\new_[7216]_ ;
  assign n4340 = ~\new_[6420]_  | ~\new_[7502]_  | ~\new_[7247]_ ;
  assign n4645 = ~\new_[6421]_  | ~\new_[7504]_  | ~\new_[7225]_ ;
  assign n4280 = ~\new_[6423]_  | ~\new_[7499]_  | ~\new_[7236]_ ;
  assign n4650 = ~\new_[6425]_  | ~\new_[7509]_  | ~\new_[7212]_ ;
  assign n4655 = ~\new_[6426]_  | ~\new_[7495]_  | ~\new_[7256]_ ;
  assign n4660 = ~\new_[6427]_  | ~\new_[7498]_  | ~\new_[6819]_ ;
  assign n4285 = ~\new_[6428]_  | ~\new_[7496]_  | ~\new_[7237]_ ;
  assign n4665 = ~\new_[6429]_  | ~\new_[7805]_  | ~\new_[7231]_ ;
  assign n4670 = ~\new_[6430]_  | ~\new_[7524]_  | ~\new_[7228]_ ;
  assign n4675 = ~\new_[6431]_  | ~\new_[7514]_  | ~\new_[7248]_ ;
  assign n4290 = ~\new_[6575]_  | ~\new_[7521]_  | ~\new_[7235]_ ;
  assign n4680 = ~\new_[6433]_  | ~\new_[7503]_  | ~\new_[7226]_ ;
  assign n4685 = ~\new_[6434]_  | ~\new_[7798]_  | ~\new_[6800]_ ;
  assign n4690 = ~\new_[6435]_  | ~\new_[7799]_  | ~\new_[7218]_ ;
  assign n4260 = ~\new_[6436]_  | ~\new_[7801]_  | ~\new_[7232]_ ;
  assign n4695 = ~\new_[6422]_  | ~\new_[7522]_  | ~\new_[7250]_ ;
  assign \new_[5318]_  = \\u4_u0_dma_out_left_reg[10] ;
  assign n4700 = ~\new_[6437]_  | ~\new_[7828]_  | ~\new_[7233]_ ;
  assign \new_[5320]_  = \\u4_u1_dma_out_left_reg[10] ;
  assign n4705 = ~\new_[6438]_  | ~\new_[7830]_  | ~\new_[6820]_ ;
  assign \new_[5322]_  = \\u4_u2_dma_out_left_reg[10] ;
  assign n4270 = ~\new_[6439]_  | ~\new_[7523]_  | ~\new_[6821]_ ;
  assign n4710 = ~\new_[6440]_  | ~\new_[7833]_  | ~\new_[6803]_ ;
  assign n4715 = ~\new_[6441]_  | ~\new_[7834]_  | ~\new_[7227]_ ;
  assign n4720 = ~\new_[6443]_  | ~\new_[7835]_  | ~\new_[6822]_ ;
  assign n4255 = ~\new_[6444]_  | ~\new_[7836]_  | ~\new_[6823]_ ;
  assign n4725 = ~\new_[6527]_  | ~\new_[7812]_  | ~\new_[6802]_ ;
  assign n4730 = ~\new_[6442]_  | ~\new_[7837]_  | ~\new_[6825]_ ;
  assign n4240 = ~\new_[6446]_  | ~\new_[7800]_  | ~\new_[6808]_ ;
  assign n4900 = ~\new_[6451]_  | ~\new_[7512]_  | ~\new_[7255]_ ;
  assign n4740 = ~\new_[6329]_  | ~\new_[7791]_  | ~\new_[6790]_ ;
  assign n4745 = ~\new_[6396]_  | ~\new_[7819]_  | ~\new_[6826]_ ;
  assign n4750 = ~\new_[6487]_  | ~\new_[7508]_  | ~\new_[7252]_ ;
  assign n4245 = ~\new_[6447]_  | ~\new_[7804]_  | ~\new_[7253]_ ;
  assign n4755 = ~\new_[6448]_  | ~\new_[7525]_  | ~\new_[6827]_ ;
  assign n4760 = ~\new_[6449]_  | ~\new_[7838]_  | ~\new_[7238]_ ;
  assign n4765 = ~\new_[6450]_  | ~\new_[7526]_  | ~\new_[7254]_ ;
  assign n4770 = ~\new_[6452]_  | ~\new_[7829]_  | ~\new_[6828]_ ;
  assign n4895 = ~\new_[6454]_  | ~\new_[7513]_  | ~\new_[7257]_ ;
  assign n4785 = ~\new_[6156]_  | ~\new_[7839]_  | ~\new_[7230]_ ;
  assign \new_[5342]_  = \new_[2053]_  ? \new_[7548]_  : \new_[14166]_ ;
  assign n4790 = ~\new_[6456]_  | ~\new_[7840]_  | ~\new_[7213]_ ;
  assign n4795 = ~\new_[6457]_  | ~\new_[7841]_  | ~\new_[6829]_ ;
  assign n4885 = ~\new_[6458]_  | ~\new_[7528]_  | ~\new_[6830]_ ;
  assign n4800 = ~\new_[6459]_  | ~\new_[7842]_  | ~\new_[7243]_ ;
  assign n4475 = ~\new_[6460]_  | ~\new_[7843]_  | ~\new_[7224]_ ;
  assign \new_[5348]_  = \new_[2052]_  ? \new_[7548]_  : \new_[14198]_ ;
  assign \new_[5349]_  = ~\new_[5939]_  & ~\new_[14640]_ ;
  assign \wb_data_o[30]  = \\u5_wb_data_o_reg[30] ;
  assign \new_[5351]_  = ~\new_[6766]_  | ~\new_[5959]_ ;
  assign \new_[5352]_  = \new_[2064]_  ? \new_[6594]_  : \new_[13589]_ ;
  assign \wb_data_o[31]  = \\u5_wb_data_o_reg[31] ;
  assign \new_[5354]_  = ~\new_[6763]_  | ~\new_[8417]_  | ~\new_[7189]_ ;
  assign \new_[5355]_  = ~\new_[5913]_  & ~\new_[6220]_ ;
  assign \new_[5356]_  = ~\new_[5941]_  & (~\new_[6695]_  | ~\new_[13688]_ );
  assign \new_[5357]_  = ~\new_[8794]_  | (~\new_[6546]_  & ~\new_[11104]_ );
  assign \new_[5358]_  = ~\new_[5942]_  & (~\new_[6695]_  | ~\new_[13883]_ );
  assign \new_[5359]_  = ~\new_[5943]_  & (~\new_[6695]_  | ~\new_[13587]_ );
  assign \new_[5360]_  = \new_[14008]_  ? \new_[8608]_  : \new_[6212]_ ;
  assign \new_[5361]_  = \new_[14223]_  ? \new_[8608]_  : \new_[6216]_ ;
  assign \new_[5362]_  = \new_[14217]_  ? \new_[8608]_  : \new_[6217]_ ;
  assign n4300 = ~\new_[5945]_  & ~n8885;
  assign n4470 = ~\new_[5950]_  & ~\new_[13373]_ ;
  assign \new_[5365]_  = \new_[13728]_  ? \new_[7549]_  : \new_[6173]_ ;
  assign \new_[5366]_  = \new_[14087]_  ? \new_[7549]_  : \new_[6176]_ ;
  assign \new_[5367]_  = ~\new_[2372]_  | ~\new_[10402]_  | ~\new_[6522]_ ;
  assign \new_[5368]_  = ~\new_[5953]_  & (~\new_[6695]_  | ~\new_[13535]_ );
  assign \new_[5369]_  = ~\new_[5954]_  & (~\new_[6695]_  | ~\new_[14027]_ );
  assign \new_[5370]_  = \new_[3691]_  ? \new_[6476]_  : \new_[9923]_ ;
  assign \new_[5371]_  = \new_[3481]_  ? \new_[6476]_  : \new_[9074]_ ;
  assign \new_[5372]_  = \new_[3479]_  ? \new_[6476]_  : \new_[8319]_ ;
  assign \new_[5373]_  = \new_[3626]_  ? \new_[6476]_  : \new_[9385]_ ;
  assign \new_[5374]_  = \new_[3482]_  ? \new_[6476]_  : \new_[8714]_ ;
  assign \new_[5375]_  = \new_[3689]_  ? \new_[6476]_  : \new_[8715]_ ;
  assign \new_[5376]_  = ~\new_[2392]_  | ~\new_[10402]_  | ~\new_[6522]_ ;
  assign \new_[5377]_  = (~\new_[6555]_  | ~\new_[13543]_ ) & (~\new_[6847]_  | ~\new_[2266]_ );
  assign \new_[5378]_  = (~\new_[6555]_  | ~\new_[13786]_ ) & (~\new_[6847]_  | ~\new_[2047]_ );
  assign \new_[5379]_  = (~\new_[6555]_  | ~\new_[13982]_ ) & (~\new_[6847]_  | ~\new_[2048]_ );
  assign \new_[5380]_  = (~\new_[6555]_  | ~\new_[13792]_ ) & (~\new_[6847]_  | ~\new_[5421]_ );
  assign \new_[5381]_  = (~\new_[6555]_  | ~\new_[13652]_ ) & (~\new_[6847]_  | ~\new_[3102]_ );
  assign \new_[5382]_  = (~\new_[6555]_  | ~\new_[14092]_ ) & (~\new_[6847]_  | ~\new_[3173]_ );
  assign \new_[5383]_  = (~\new_[7284]_  | ~\new_[14062]_ ) & (~\new_[6847]_  | ~\new_[2178]_ );
  assign \new_[5384]_  = (~\new_[7284]_  | ~\new_[14154]_ ) & (~\new_[6847]_  | ~\new_[3034]_ );
  assign \new_[5385]_  = (~\new_[6555]_  | ~\new_[14178]_ ) & (~\new_[6847]_  | ~\new_[3021]_ );
  assign \new_[5386]_  = (~\new_[6555]_  | ~\new_[14024]_ ) & (~\new_[6847]_  | ~\new_[9037]_ );
  assign \new_[5387]_  = (~\new_[7284]_  | ~\new_[13854]_ ) & (~\new_[6847]_  | ~\new_[2928]_ );
  assign \new_[5388]_  = (~\new_[6555]_  | ~\new_[13707]_ ) & (~\new_[6847]_  | ~\new_[2856]_ );
  assign \new_[5389]_  = (~\new_[6555]_  | ~\new_[13983]_ ) & (~\new_[6847]_  | ~\new_[2638]_ );
  assign \new_[5390]_  = (~\new_[7284]_  | ~\new_[14113]_ ) & (~\new_[6847]_  | ~\new_[2639]_ );
  assign \new_[5391]_  = (~\new_[7284]_  | ~\new_[14137]_ ) & (~\new_[6847]_  | ~\new_[2547]_ );
  assign \new_[5392]_  = (~\new_[6555]_  | ~\new_[14255]_ ) & (~\new_[6847]_  | ~\new_[2735]_ );
  assign \new_[5393]_  = (~\new_[6555]_  | ~\new_[13739]_ ) & (~\new_[6847]_  | ~\new_[2177]_ );
  assign \new_[5394]_  = (~\new_[6555]_  | ~\new_[14220]_ ) & (~\new_[6847]_  | ~\new_[2265]_ );
  assign \new_[5395]_  = (~\new_[6555]_  | ~\new_[13622]_ ) & (~\new_[6847]_  | ~\new_[2136]_ );
  assign \new_[5396]_  = (~\new_[6555]_  | ~\new_[14145]_ ) & (~\new_[6847]_  | ~\new_[2075]_ );
  assign \new_[5397]_  = (~\new_[6555]_  | ~\new_[13683]_ ) & (~\new_[6847]_  | ~\new_[2062]_ );
  assign \new_[5398]_  = ~\new_[5980]_  & ~\new_[9137]_ ;
  assign \new_[5399]_  = ~\new_[5982]_  & ~\new_[9137]_ ;
  assign \new_[5400]_  = ~\new_[5989]_  & ~\new_[9137]_ ;
  assign n4320 = ~\new_[5895]_  & (~\new_[12287]_  | ~\new_[9080]_ );
  assign \new_[5402]_  = ~\new_[5968]_  | ~\new_[12840]_ ;
  assign \new_[5403]_  = \new_[2040]_  ? \new_[6594]_  : \new_[13524]_ ;
  assign \new_[5404]_  = ~\new_[10631]_  & (~\new_[9813]_  | ~\new_[6480]_ );
  assign \new_[5405]_  = ~\new_[10653]_  & (~\new_[9814]_  | ~\new_[6482]_ );
  assign \new_[5406]_  = ~\new_[6084]_  & ~\new_[14225]_ ;
  assign \new_[5407]_  = ~\new_[6084]_  & ~\new_[14071]_ ;
  assign n4265 = ~\new_[9017]_  | ~\new_[8865]_  | ~\new_[6833]_  | ~\new_[6467]_ ;
  assign \new_[5409]_  = ~\new_[6084]_  & ~\new_[14215]_ ;
  assign \new_[5410]_  = \new_[3592]_  ? \new_[6476]_  : \new_[8189]_ ;
  assign \new_[5411]_  = \new_[3684]_  ? \new_[6476]_  : \new_[7462]_ ;
  assign \new_[5412]_  = ~\new_[5944]_  & (~\new_[6695]_  | ~\new_[13789]_ );
  assign \new_[5413]_  = \new_[13874]_  ? \new_[7544]_  : \new_[6525]_ ;
  assign \new_[5414]_  = ~\new_[6084]_  & ~\new_[11733]_ ;
  assign \new_[5415]_  = ~\new_[6084]_  & ~\new_[11577]_ ;
  assign \new_[5416]_  = ~\new_[5952]_  | ~\new_[6070]_ ;
  assign \new_[5417]_  = ~\new_[6061]_  & ~\new_[9137]_ ;
  assign \new_[5418]_  = ~\new_[6084]_  & ~\new_[14100]_ ;
  assign \new_[5419]_  = ~\new_[6705]_  & ~\new_[6221]_ ;
  assign \new_[5420]_  = ~\new_[5983]_  & ~\new_[6224]_ ;
  assign \new_[5421]_  = \\u1_u3_idin_reg[17] ;
  assign \new_[5422]_  = ~\new_[6029]_  | ~\new_[12840]_ ;
  assign \new_[5423]_  = ~\new_[6768]_  | ~\new_[6769]_  | ~\new_[12085]_  | ~\new_[14329]_ ;
  assign n4330 = ~\new_[5895]_  & (~\new_[12295]_  | ~\new_[8915]_ );
  assign \new_[5425]_  = ~\new_[5722]_ ;
  assign n4365 = ~\new_[5966]_  & ~n8885;
  assign \new_[5427]_  = \new_[3502]_  ? \new_[6476]_  : \new_[12036]_ ;
  assign \new_[5428]_  = \new_[13634]_  ? \new_[8608]_  : \new_[6508]_ ;
  assign \new_[5429]_  = \new_[6602]_  ? \new_[8608]_  : \new_[6496]_ ;
  assign \new_[5430]_  = \new_[6300]_  ? \new_[7544]_  : \new_[6498]_ ;
  assign \new_[5431]_  = \new_[14133]_  ? \new_[8608]_  : \new_[6504]_ ;
  assign \new_[5432]_  = \new_[14210]_  ? \new_[7544]_  : \new_[6507]_ ;
  assign \new_[5433]_  = \new_[13696]_  ? \new_[7544]_  : \new_[6509]_ ;
  assign \new_[5434]_  = \new_[13907]_  ? \new_[7544]_  : \new_[6495]_ ;
  assign \new_[5435]_  = \new_[6733]_  ? \new_[8608]_  : \new_[6494]_ ;
  assign \new_[5436]_  = ~\new_[10668]_  & (~\new_[9816]_  | ~\new_[6558]_ );
  assign \new_[5437]_  = \new_[6301]_  ? \new_[7544]_  : \new_[6499]_ ;
  assign \new_[5438]_  = \new_[13518]_  ? \new_[8608]_  : \new_[6493]_ ;
  assign \new_[5439]_  = \new_[13720]_  ? \new_[7544]_  : \new_[6514]_ ;
  assign \new_[5440]_  = \new_[6305]_  ? \new_[7544]_  : \new_[6505]_ ;
  assign \new_[5441]_  = \new_[14239]_  ? \new_[8608]_  : \new_[6506]_ ;
  assign \new_[5442]_  = \new_[6588]_  ? \new_[8608]_  : \new_[6501]_ ;
  assign \new_[5443]_  = \new_[14160]_  ? \new_[7549]_  : \new_[6515]_ ;
  assign \new_[5444]_  = \new_[14176]_  ? \new_[7549]_  : \new_[6510]_ ;
  assign \new_[5445]_  = \new_[14091]_  ? \new_[7549]_  : \new_[6516]_ ;
  assign \new_[5446]_  = \new_[6344]_  ? \new_[7549]_  : \new_[6517]_ ;
  assign \new_[5447]_  = \new_[6351]_  ? \new_[7549]_  : \new_[6518]_ ;
  assign \new_[5448]_  = \new_[14049]_  ? \new_[7549]_  : \new_[6519]_ ;
  assign \new_[5449]_  = \new_[9708]_  ? \new_[12840]_  : \new_[6133]_ ;
  assign \new_[5450]_  = \new_[6853]_  ? \new_[8608]_  : \new_[6513]_ ;
  assign \new_[5451]_  = \new_[6302]_  ? \new_[7544]_  : \new_[6500]_ ;
  assign \new_[5452]_  = \new_[6299]_  ? \new_[8608]_  : \new_[6497]_ ;
  assign \new_[5453]_  = \new_[6560]_  ? \new_[7544]_  : \new_[6503]_ ;
  assign \new_[5454]_  = \new_[3777]_  ? \new_[6476]_  : \new_[10777]_ ;
  assign \new_[5455]_  = \new_[3711]_  ? \new_[6476]_  : \new_[10698]_ ;
  assign \new_[5456]_  = \new_[3788]_  ? \new_[6476]_  : \new_[9972]_ ;
  assign \new_[5457]_  = \new_[13534]_  ? \new_[7544]_  : \new_[6520]_ ;
  assign \new_[5458]_  = \new_[3507]_  ? \new_[6476]_  : \new_[12885]_ ;
  assign \new_[5459]_  = \new_[3508]_  ? \new_[6476]_  : \new_[11454]_ ;
  assign \new_[5460]_  = \new_[3509]_  ? \new_[6476]_  : \new_[9973]_ ;
  assign \new_[5461]_  = \new_[3510]_  ? \new_[6476]_  : \new_[9709]_ ;
  assign \new_[5462]_  = \new_[3712]_  ? \new_[6476]_  : \new_[9119]_ ;
  assign \new_[5463]_  = \new_[6303]_  ? \new_[7544]_  : \new_[6502]_ ;
  assign \new_[5464]_  = \new_[2049]_  ? \new_[7548]_  : \new_[13538]_ ;
  assign \new_[5465]_  = \new_[14064]_  ? \new_[7544]_  : \new_[6492]_ ;
  assign \new_[5466]_  = \new_[9936]_  ? \new_[12840]_  : \new_[6587]_ ;
  assign \new_[5467]_  = (~\new_[10038]_  | ~\new_[9427]_ ) & (~\new_[6523]_  | ~\new_[4290]_ );
  assign \new_[5468]_  = \new_[9554]_  ? \new_[12840]_  : \new_[6590]_ ;
  assign \new_[5469]_  = \new_[3686]_  ? \new_[6476]_  : \new_[6856]_ ;
  assign \new_[5470]_  = \new_[3468]_  ? \new_[6476]_  : \new_[7305]_ ;
  assign \new_[5471]_  = ~\new_[6037]_  & (~\new_[6695]_  | ~\new_[13856]_ );
  assign \new_[5472]_  = ~\new_[2933]_  & (~\new_[6521]_  | ~\new_[14216]_ );
  assign \new_[5473]_  = ~\new_[11104]_  & (~\new_[6532]_  | ~\new_[13595]_ );
  assign \new_[5474]_  = \new_[13515]_  ? \new_[8608]_  : \new_[6104]_ ;
  assign \new_[5475]_  = ~\new_[5746]_ ;
  assign n4805 = ~\new_[12732]_  & (~\new_[6839]_  | ~\new_[6534]_ );
  assign n4810 = ~\new_[12505]_  & (~\new_[6535]_  | ~\new_[6840]_ );
  assign \new_[5478]_  = \new_[13574]_  ? \new_[8608]_  : \new_[6106]_ ;
  assign n4815 = ~\new_[12794]_  & (~\new_[6841]_  | ~\new_[6531]_ );
  assign n4880 = ~\new_[12849]_  & (~\new_[6536]_  | ~\new_[6835]_ );
  assign \new_[5481]_  = ~\new_[6761]_  & ~\new_[6028]_ ;
  assign \new_[5482]_  = ~\new_[5748]_ ;
  assign \new_[5483]_  = \new_[14260]_  ? \new_[7544]_  : \new_[6108]_ ;
  assign \new_[5484]_  = \new_[2082]_  ? \new_[6594]_  : \new_[14143]_ ;
  assign \new_[5485]_  = \new_[14121]_  ? \new_[7544]_  : \new_[6158]_ ;
  assign \new_[5486]_  = \\u0_u0_state_reg[9] ;
  assign \wb_data_o[27]  = \\u5_wb_data_o_reg[27] ;
  assign \wb_data_o[29]  = \\u5_wb_data_o_reg[29] ;
  assign \new_[5489]_  = \\u4_u3_int_stat_reg[3] ;
  assign \new_[5490]_  = \\u4_u0_int_stat_reg[3] ;
  assign \new_[5491]_  = \\u4_u1_int_stat_reg[3] ;
  assign \new_[5492]_  = u0_u0_T1_st_3_0_mS_reg;
  assign \wb_data_o[11]  = \\u5_wb_data_o_reg[11] ;
  assign \wb_data_o[9]  = \\u5_wb_data_o_reg[9] ;
  assign \new_[5495]_  = ~\\u0_u0_chirp_cnt_reg[0] ;
  assign \new_[5496]_  = ~\new_[6024]_  & (~\new_[6695]_  | ~\new_[13800]_ );
  assign \new_[5497]_  = ~\new_[6025]_  & (~\new_[6695]_  | ~\new_[14159]_ );
  assign \wb_data_o[12]  = \\u5_wb_data_o_reg[12] ;
  assign \new_[5499]_  = \\u4_u0_int_stat_reg[6] ;
  assign \new_[5500]_  = ~\new_[6026]_  & (~\new_[6695]_  | ~\new_[13528]_ );
  assign \new_[5501]_  = \\u0_u0_state_reg[4] ;
  assign \new_[5502]_  = \\u4_u2_uc_bsel_reg[0] ;
  assign \new_[5503]_  = \\u4_u2_uc_bsel_reg[1] ;
  assign \new_[5504]_  = \\u4_u2_uc_dpd_reg[0] ;
  assign n4415 = ~\new_[5895]_  & (~\new_[12399]_  | ~\new_[9591]_ );
  assign \new_[5506]_  = ~\new_[6084]_  & ~\new_[13708]_ ;
  assign \new_[5507]_  = ~\new_[6084]_  & ~\new_[14191]_ ;
  assign \new_[5508]_  = ~\new_[6084]_  & ~\new_[13992]_ ;
  assign \new_[5509]_  = \new_[12798]_  ? \new_[6522]_  : \new_[2476]_ ;
  assign \new_[5510]_  = ~n4975;
  assign \new_[5511]_  = ~n5230;
  assign \new_[5512]_  = ~n5200;
  assign n4370 = ~\new_[5774]_ ;
  assign \new_[5514]_  = ~n4200;
  assign n4825 = ~\new_[5776]_ ;
  assign n4830 = ~\new_[5777]_ ;
  assign n4375 = ~\new_[5778]_ ;
  assign \new_[5518]_  = ~n4205;
  assign \new_[5519]_  = ~n4210;
  assign \new_[5520]_  = ~n5225;
  assign n4835 = ~\new_[5782]_ ;
  assign n4840 = ~\new_[5783]_ ;
  assign n4845 = ~\new_[5784]_ ;
  assign n4875 = ~\new_[5785]_ ;
  assign \new_[5525]_  = ~n4195;
  assign n4820 = ~\new_[5787]_ ;
  assign \new_[5527]_  = ~\new_[10442]_  | (~\new_[6119]_  & ~\new_[13403]_ );
  assign \new_[5528]_  = \new_[9597]_  ? \new_[12840]_  : \new_[6128]_ ;
  assign \new_[5529]_  = ~\new_[5888]_  & ~\new_[9137]_ ;
  assign \new_[5530]_  = ~\new_[5889]_  & ~\new_[9137]_ ;
  assign \new_[5531]_  = ~\new_[5891]_  & ~\new_[9137]_ ;
  assign \new_[5532]_  = \new_[3464]_  ? \new_[6476]_  : \new_[6626]_ ;
  assign \new_[5533]_  = ~\new_[5923]_  & ~\new_[9137]_ ;
  assign \new_[5534]_  = \new_[10228]_  ? \new_[12840]_  : \new_[6131]_ ;
  assign n4405 = \new_[6094]_  ? \wb_addr_i[17]  : \sram_data_i[22] ;
  assign n4345 = \new_[6095]_  ? \wb_addr_i[17]  : \sram_data_i[23] ;
  assign n4410 = \new_[6096]_  ? \wb_addr_i[17]  : \sram_data_i[7] ;
  assign \new_[5538]_  = ~\new_[6058]_  & ~\new_[2933]_ ;
  assign \new_[5539]_  = ~\new_[6084]_  & ~\new_[13927]_ ;
  assign \new_[5540]_  = ~\new_[6565]_  | ~\new_[9065]_  | ~\new_[6649]_ ;
  assign \new_[5541]_  = ~\new_[6586]_  | ~\new_[8693]_  | ~\new_[6660]_ ;
  assign \new_[5542]_  = ~\new_[7904]_  | ~\new_[6612]_  | ~\new_[6851]_  | ~\new_[7321]_ ;
  assign \new_[5543]_  = ~\new_[7680]_  | ~\new_[6613]_  | ~\new_[6080]_  | ~\new_[6614]_ ;
  assign \new_[5544]_  = ~\new_[6067]_  | (~\new_[7858]_  & ~\new_[11733]_ );
  assign \new_[5545]_  = ~\new_[6065]_  | (~\new_[7858]_  & ~\new_[11577]_ );
  assign \new_[5546]_  = \new_[2266]_  ? \new_[6594]_  : \new_[14022]_ ;
  assign \new_[5547]_  = \new_[3102]_  ? \new_[6594]_  : \new_[14112]_ ;
  assign \new_[5548]_  = \new_[3173]_  ? \new_[6594]_  : \new_[13830]_ ;
  assign \new_[5549]_  = \new_[2178]_  ? \new_[6594]_  : \new_[13582]_ ;
  assign \new_[5550]_  = \new_[3034]_  ? \new_[6594]_  : \new_[13775]_ ;
  assign \new_[5551]_  = \new_[3021]_  ? \new_[6594]_  : \new_[14158]_ ;
  assign \new_[5552]_  = \new_[2928]_  ? \new_[6594]_  : \new_[13529]_ ;
  assign \new_[5553]_  = \new_[2856]_  ? \new_[6594]_  : \new_[13685]_ ;
  assign \new_[5554]_  = \new_[2638]_  ? \new_[6594]_  : \new_[14075]_ ;
  assign \new_[5555]_  = \new_[2639]_  ? \new_[6594]_  : \new_[13846]_ ;
  assign \new_[5556]_  = \new_[2547]_  ? \new_[6594]_  : \new_[13678]_ ;
  assign \new_[5557]_  = \new_[2265]_  ? \new_[7548]_  : \new_[13831]_ ;
  assign \new_[5558]_  = \new_[2136]_  ? \new_[6594]_  : \new_[13527]_ ;
  assign \new_[5559]_  = \new_[2075]_  ? \new_[6594]_  : \new_[14249]_ ;
  assign \new_[5560]_  = \new_[2062]_  ? \new_[6594]_  : \new_[13965]_ ;
  assign n4445 = ~\new_[5906]_  & ~\new_[12245]_ ;
  assign \new_[5562]_  = \\u4_u2_int_stat_reg[3] ;
  assign \new_[5563]_  = ~\new_[5907]_  & ~\new_[9137]_ ;
  assign \new_[5564]_  = \new_[5890]_  & \new_[6565]_ ;
  assign \new_[5565]_  = ~\new_[5908]_  & ~\new_[9137]_ ;
  assign n4430 = ~\new_[6177]_  | ~\new_[5905]_ ;
  assign \new_[5567]_  = \new_[2034]_  ? \new_[6594]_  : \new_[14209]_ ;
  assign \new_[5568]_  = \new_[13721]_  ? \new_[7544]_  : \new_[6199]_ ;
  assign n4435 = ~\new_[5895]_  & (~\new_[12293]_  | ~\new_[12024]_ );
  assign n4305 = ~\new_[5895]_  & (~\new_[12461]_  | ~\new_[11041]_ );
  assign n4440 = ~\new_[5895]_  & (~\new_[11946]_  | ~\new_[10307]_ );
  assign n4450 = ~\new_[5895]_  & (~\new_[12296]_  | ~\new_[9446]_ );
  assign n4325 = ~\new_[5895]_  & (~\new_[12266]_  | ~\new_[9039]_ );
  assign n4860 = ~\new_[10854]_  & ~\new_[5903]_ ;
  assign \new_[5575]_  = ~\new_[5849]_ ;
  assign \new_[5576]_  = \new_[5892]_  & \new_[6586]_ ;
  assign n4455 = ~\new_[5899]_  & ~\new_[13679]_ ;
  assign n4460 = ~\new_[5899]_  & (~\new_[12733]_  | ~\new_[12827]_ );
  assign n4315 = ~\new_[11908]_  & ~\new_[5899]_ ;
  assign n4465 = ~\new_[11019]_  & ~\new_[5899]_ ;
  assign \new_[5581]_  = \new_[6613]_  & \new_[6080]_ ;
  assign \new_[5582]_  = ~\new_[3309]_  | ~\new_[6080]_  | ~\new_[8718]_ ;
  assign \new_[5583]_  = ~\new_[6082]_  & (~\new_[6695]_  | ~\new_[13607]_ );
  assign n4380 = ~\new_[5859]_ ;
  assign \new_[5585]_  = \\u0_u0_state_reg[3] ;
  assign \new_[5586]_  = ~\new_[7316]_  & (~\new_[7453]_  | ~\new_[6183]_ );
  assign n4425 = ~\new_[5894]_  & (~\new_[11462]_  | ~\new_[13111]_ );
  assign \new_[5588]_  = \new_[10969]_  ? \new_[12840]_  : \new_[6190]_ ;
  assign \new_[5589]_  = \new_[10309]_  ? \new_[12840]_  : \new_[6191]_ ;
  assign \new_[5590]_  = \new_[10064]_  ? \new_[12840]_  : \new_[6195]_ ;
  assign \new_[5591]_  = \new_[12213]_  ? \new_[12840]_  : \new_[6189]_ ;
  assign \new_[5592]_  = ~\new_[6084]_  & ~\new_[13642]_ ;
  assign n4385 = ~\new_[5960]_  | ~\new_[10117]_ ;
  assign n4890 = ~\new_[5961]_  | ~\new_[10117]_ ;
  assign n4395 = ~\new_[5962]_  | ~\new_[10117]_ ;
  assign n4420 = \new_[6159]_  ? \wb_addr_i[17]  : \sram_data_i[8] ;
  assign n4390 = ~\new_[5964]_  | ~\new_[10117]_ ;
  assign n4235 = ~\new_[5965]_  | ~\new_[10117]_ ;
  assign \new_[5599]_  = \new_[3688]_  ? \new_[6476]_  : \new_[7686]_ ;
  assign \wb_data_o[10]  = \\u5_wb_data_o_reg[10] ;
  assign \new_[5601]_  = \new_[3638]_  ? \new_[6476]_  : \new_[7913]_ ;
  assign \new_[5602]_  = \new_[3467]_  ? \new_[6476]_  : \new_[7404]_ ;
  assign \new_[5603]_  = (~\new_[6185]_  | ~\new_[6175]_ ) & (~\new_[7741]_  | ~\new_[6175]_ );
  assign \new_[5604]_  = \\u4_u2_uc_dpd_reg[1] ;
  assign \new_[5605]_  = ~\new_[2933]_  & (~\new_[6521]_  | ~\new_[13369]_ );
  assign n4870 = u1_u0_data_valid0_reg;
  assign \new_[5607]_  = ~\new_[7417]_  & (~\new_[6648]_  | ~\new_[3686]_ );
  assign XcvSelect_pad_o = u0_u0_XcvSelect_reg;
  assign n5085 = ~\new_[13296]_  & (~\new_[7867]_  | ~\new_[6779]_ );
  assign n5095 = ~\new_[6204]_  & ~\new_[13386]_ ;
  assign n5105 = ~\new_[6205]_  & ~\new_[13386]_ ;
  assign \new_[5612]_  = ~\new_[6186]_  | ~\new_[12840]_ ;
  assign \new_[5613]_  = \new_[2053]_  ? \new_[7858]_  : \new_[14173]_ ;
  assign \new_[5614]_  = \new_[2052]_  ? \new_[7858]_  : \new_[13553]_ ;
  assign \OpMode_pad_o[1]  = \\u0_u0_OpMode_reg[1] ;
  assign \new_[5616]_  = \new_[2064]_  ? \new_[6860]_  : \new_[13958]_ ;
  assign \new_[5617]_  = \\u4_int_srcb_reg[8] ;
  assign \new_[5618]_  = ~\new_[7453]_  | ~\new_[6182]_ ;
  assign \new_[5619]_  = ~\new_[6192]_  | ~\new_[12840]_ ;
  assign \new_[5620]_  = ~\new_[6193]_  | ~\new_[12840]_ ;
  assign \new_[5621]_  = ~\new_[6197]_  | ~\new_[12840]_ ;
  assign \new_[5622]_  = ~\new_[6194]_  | ~\new_[12840]_ ;
  assign \new_[5623]_  = \new_[6134]_  & \new_[6631]_ ;
  assign \new_[5624]_  = ~\new_[12163]_  | ~\new_[6464]_ ;
  assign \new_[5625]_  = \new_[14257]_  ? \new_[7857]_  : \new_[6848]_ ;
  assign \new_[5626]_  = \new_[14017]_  ? \new_[7857]_  : \new_[6628]_ ;
  assign \new_[5627]_  = ~\new_[5912]_ ;
  assign \new_[5628]_  = \new_[3692]_  ? \new_[6778]_  : \new_[8716]_ ;
  assign \new_[5629]_  = \new_[3884]_  ? \new_[6778]_  : \new_[9925]_ ;
  assign \new_[5630]_  = \new_[3693]_  ? \new_[6778]_  : \new_[9072]_ ;
  assign \new_[5631]_  = \new_[3690]_  ? \new_[6778]_  : \new_[8321]_ ;
  assign \new_[5632]_  = ~\new_[5914]_ ;
  assign \new_[5633]_  = \new_[3806]_  ? \new_[6778]_  : \new_[9387]_ ;
  assign \new_[5634]_  = \new_[3815]_  ? \new_[6778]_  : \new_[8709]_ ;
  assign \new_[5635]_  = (~\new_[6779]_  | ~\new_[4503]_ ) & (~\new_[7289]_  | ~\new_[4597]_ );
  assign \new_[5636]_  = (~\new_[6779]_  | ~\new_[4372]_ ) & (~\new_[7289]_  | ~\new_[4506]_ );
  assign \new_[5637]_  = (~\new_[6779]_  | ~\new_[4504]_ ) & (~\new_[7289]_  | ~\new_[4507]_ );
  assign \new_[5638]_  = (~\new_[6779]_  | ~\new_[4552]_ ) & (~\new_[7289]_  | ~\new_[4508]_ );
  assign \new_[5639]_  = (~\new_[6779]_  | ~\new_[4505]_ ) & (~\new_[7289]_  | ~\new_[4553]_ );
  assign \new_[5640]_  = (~\new_[6779]_  | ~\new_[4597]_ ) & (~\new_[7289]_  | ~\new_[11060]_ );
  assign \new_[5641]_  = (~\new_[6779]_  | ~\new_[4506]_ ) & (~\new_[7289]_  | ~\new_[10416]_ );
  assign \new_[5642]_  = (~\new_[6779]_  | ~\new_[4507]_ ) & (~\new_[7289]_  | ~\new_[11061]_ );
  assign \new_[5643]_  = (~\new_[6779]_  | ~\new_[4508]_ ) & (~\new_[7289]_  | ~\new_[10772]_ );
  assign \new_[5644]_  = (~\new_[6779]_  | ~\new_[4553]_ ) & (~\new_[7289]_  | ~\new_[11062]_ );
  assign \new_[5645]_  = (~\new_[6779]_  | ~\new_[4509]_ ) & (~\new_[7289]_  | ~\new_[10773]_ );
  assign \new_[5646]_  = (~\new_[6779]_  | ~\new_[4510]_ ) & (~\new_[7289]_  | ~\new_[10334]_ );
  assign \new_[5647]_  = (~\new_[6779]_  | ~\new_[4511]_ ) & (~\new_[7289]_  | ~\new_[10774]_ );
  assign n5090 = \new_[13166]_  ? \new_[6779]_  : \new_[13630]_ ;
  assign n4945 = \new_[12846]_  ? \new_[6779]_  : \new_[13769]_ ;
  assign n5100 = \new_[12783]_  ? \new_[6779]_  : \new_[13558]_ ;
  assign n4950 = \new_[12870]_  ? \new_[6779]_  : \new_[13572]_ ;
  assign n4935 = \new_[12651]_  ? \new_[6779]_  : \new_[13997]_ ;
  assign n5110 = \new_[12816]_  ? \new_[6779]_  : \new_[13565]_ ;
  assign n5115 = \new_[12916]_  ? \new_[6779]_  : \new_[13567]_ ;
  assign n5120 = \new_[13192]_  ? \new_[6779]_  : \new_[13573]_ ;
  assign n4905 = \new_[13630]_  ? \new_[6779]_  : \new_[13703]_ ;
  assign n5125 = \new_[13769]_  ? \new_[6779]_  : \new_[13715]_ ;
  assign n5130 = \new_[13558]_  ? \new_[6779]_  : \new_[13650]_ ;
  assign n5135 = \new_[13572]_  ? \new_[6779]_  : \new_[13541]_ ;
  assign n4920 = \new_[13997]_  ? \new_[6779]_  : \new_[13906]_ ;
  assign n5140 = \new_[13565]_  ? \new_[6779]_  : \new_[13674]_ ;
  assign n5145 = \new_[13567]_  ? \new_[6779]_  : \new_[13827]_ ;
  assign n5150 = \new_[13573]_  ? \new_[6779]_  : \new_[13851]_ ;
  assign n5215 = \new_[13703]_  ? \new_[6779]_  : n9060;
  assign n5155 = \new_[13715]_  ? \new_[6779]_  : n9080;
  assign n5160 = \new_[13650]_  ? \new_[6779]_  : n9065;
  assign n5165 = \new_[13541]_  ? \new_[6779]_  : n9070;
  assign n5220 = \new_[13906]_  ? \new_[6779]_  : n9045;
  assign n5170 = \new_[13674]_  ? \new_[6779]_  : n9085;
  assign n5175 = \new_[13827]_  ? \new_[6779]_  : n9090;
  assign n5180 = \new_[13851]_  ? \new_[6779]_  : n9055;
  assign \new_[5672]_  = (~\new_[6779]_  | ~\new_[4502]_ ) & (~\new_[7289]_  | ~\new_[9386]_ );
  assign \new_[5673]_  = (~\new_[6695]_  | ~\new_[13511]_ ) & (~\new_[7292]_  | ~\new_[2177]_ );
  assign \new_[5674]_  = (~\new_[6695]_  | ~\new_[13931]_ ) & (~\new_[7292]_  | ~\new_[2266]_ );
  assign \new_[5675]_  = (~\new_[6695]_  | ~\new_[13719]_ ) & (~\new_[7292]_  | ~\new_[2047]_ );
  assign \new_[5676]_  = (~\new_[6695]_  | ~\new_[13836]_ ) & (~\new_[7292]_  | ~\new_[2048]_ );
  assign \new_[5677]_  = (~\new_[7541]_  | ~\new_[13888]_ ) & (~\new_[7292]_  | ~\new_[3102]_ );
  assign \new_[5678]_  = (~\new_[7541]_  | ~\new_[13774]_ ) & (~\new_[7292]_  | ~\new_[3173]_ );
  assign \new_[5679]_  = (~\new_[6695]_  | ~\new_[13730]_ ) & (~\new_[7292]_  | ~\new_[2178]_ );
  assign \new_[5680]_  = (~\new_[6695]_  | ~\new_[13795]_ ) & (~\new_[7292]_  | ~\new_[3034]_ );
  assign \new_[5681]_  = (~\new_[6695]_  | ~\new_[13639]_ ) & (~\new_[7292]_  | ~\new_[3021]_ );
  assign \new_[5682]_  = (~\new_[6695]_  | ~\new_[14021]_ ) & (~\new_[7292]_  | ~\new_[9037]_ );
  assign \new_[5683]_  = (~\new_[6695]_  | ~\new_[13516]_ ) & (~\new_[7292]_  | ~\new_[2928]_ );
  assign \new_[5684]_  = (~\new_[6695]_  | ~\new_[14233]_ ) & (~\new_[7292]_  | ~\new_[2856]_ );
  assign \new_[5685]_  = (~\new_[6695]_  | ~\new_[13612]_ ) & (~\new_[7292]_  | ~\new_[2638]_ );
  assign \new_[5686]_  = (~\new_[6695]_  | ~\new_[13697]_ ) & (~\new_[7292]_  | ~\new_[2639]_ );
  assign \new_[5687]_  = (~\new_[6695]_  | ~\new_[13716]_ ) & (~\new_[7292]_  | ~\new_[2547]_ );
  assign \new_[5688]_  = (~\new_[6695]_  | ~\new_[13959]_ ) & (~\new_[7292]_  | ~\new_[2735]_ );
  assign \new_[5689]_  = (~\new_[6695]_  | ~\new_[14030]_ ) & (~\new_[7292]_  | ~\new_[2265]_ );
  assign \new_[5690]_  = (~\new_[7541]_  | ~\new_[13996]_ ) & (~\new_[7292]_  | ~\new_[2136]_ );
  assign \new_[5691]_  = (~\new_[7541]_  | ~\new_[13952]_ ) & (~\new_[7292]_  | ~\new_[2075]_ );
  assign \new_[5692]_  = (~\new_[6695]_  | ~\new_[13578]_ ) & (~\new_[7292]_  | ~\new_[2062]_ );
  assign \new_[5693]_  = (~\new_[6695]_  | ~\new_[13791]_ ) & (~\new_[7292]_  | ~\new_[5421]_ );
  assign \new_[5694]_  = ~\new_[6896]_  | ~\new_[7425]_  | ~\new_[12713]_  | ~\new_[7176]_ ;
  assign n4915 = ~\new_[8996]_  | ~\new_[8893]_  | ~\new_[7249]_  | ~\new_[6755]_ ;
  assign n4925 = ~\new_[8981]_  | ~\new_[8869]_  | ~\new_[7263]_  | ~\new_[6756]_ ;
  assign n4930 = ~\new_[8994]_  | ~\new_[8870]_  | ~\new_[7266]_  | ~\new_[6757]_ ;
  assign \new_[5698]_  = \new_[2040]_  ? \new_[6860]_  : \new_[14148]_ ;
  assign \new_[5699]_  = \new_[2082]_  ? \new_[6860]_  : \new_[14184]_ ;
  assign \new_[5700]_  = ~\new_[6184]_  & (~\new_[12427]_  | ~\new_[8208]_ );
  assign \new_[5701]_  = \new_[3790]_  ? \new_[6778]_  : \new_[8198]_ ;
  assign \new_[5702]_  = \new_[3875]_  ? \new_[6778]_  : \new_[7464]_ ;
  assign \new_[5703]_  = ~\new_[6555]_  & ~\new_[14225]_ ;
  assign \new_[5704]_  = ~\new_[7284]_  & ~\new_[14071]_ ;
  assign \new_[5705]_  = ~\new_[6555]_  & ~\new_[14215]_ ;
  assign \new_[5706]_  = \\u4_u3_dma_out_left_reg[9] ;
  assign \new_[5707]_  = \\u4_u0_dma_out_left_reg[9] ;
  assign \new_[5708]_  = \\u4_u1_dma_out_left_reg[9] ;
  assign \new_[5709]_  = \\u4_u2_dma_out_left_reg[9] ;
  assign \new_[5710]_  = ~\new_[6219]_  & ~\new_[12798]_ ;
  assign \new_[5711]_  = ~\new_[7284]_  & ~\new_[11733]_ ;
  assign \new_[5712]_  = ~\new_[6555]_  & ~\new_[11577]_ ;
  assign \new_[5713]_  = ~\new_[6555]_  & ~\new_[14100]_ ;
  assign n5185 = ~\new_[6463]_  & ~n8885;
  assign \new_[5715]_  = ~\new_[10395]_  & ~\new_[6219]_ ;
  assign \new_[5716]_  = ~\new_[7184]_  | ~\new_[7441]_  | ~\new_[13319]_  | ~\new_[14586]_ ;
  assign \new_[5717]_  = ~\new_[7440]_  | ~\new_[7185]_  | ~\new_[11671]_  | ~\new_[14421]_ ;
  assign \new_[5718]_  = ~\new_[6127]_  & (~\new_[14539]_  | ~\new_[13258]_ );
  assign \new_[5719]_  = ~\new_[6774]_  & (~\new_[7181]_  | ~\new_[6761]_ );
  assign \new_[5720]_  = ~\new_[5956]_ ;
  assign \new_[5721]_  = \new_[6223]_  & \new_[7182]_ ;
  assign \new_[5722]_  = ~\new_[6761]_  & (~\new_[6763]_  | ~\new_[7190]_ );
  assign \new_[5723]_  = ~\new_[6219]_  & (~\new_[2301]_  | ~\new_[9375]_ );
  assign n4965 = \new_[6758]_  & \new_[6464]_ ;
  assign \new_[5725]_  = \new_[3710]_  ? \new_[6778]_  : \new_[12139]_ ;
  assign \new_[5726]_  = (~\new_[14276]_  | ~\new_[7448]_ ) & (~\new_[7195]_  | ~\new_[6776]_ );
  assign \new_[5727]_  = \new_[3718]_  ? \new_[6778]_  : \new_[12895]_ ;
  assign \new_[5728]_  = \new_[3888]_  ? \new_[6778]_  : \new_[10699]_ ;
  assign \new_[5729]_  = \new_[6367]_  ? \new_[7857]_  : \new_[6785]_ ;
  assign \new_[5730]_  = \new_[6102]_  ? \new_[7857]_  : \new_[6784]_ ;
  assign \new_[5731]_  = \new_[6371]_  ? \new_[7857]_  : \new_[6783]_ ;
  assign \new_[5732]_  = \new_[6091]_  ? \new_[7857]_  : \new_[6786]_ ;
  assign \new_[5733]_  = \new_[14229]_  ? \new_[7857]_  : \new_[6782]_ ;
  assign \new_[5734]_  = \new_[13519]_  ? \new_[7857]_  : \new_[6787]_ ;
  assign \new_[5735]_  = \new_[3930]_  ? \new_[6778]_  : \new_[10769]_ ;
  assign \new_[5736]_  = \new_[3889]_  ? \new_[6778]_  : \new_[9975]_ ;
  assign \new_[5737]_  = \new_[3713]_  ? \new_[6778]_  : \new_[11710]_ ;
  assign \new_[5738]_  = \new_[3714]_  ? \new_[6778]_  : \new_[9974]_ ;
  assign \new_[5739]_  = \new_[3715]_  ? \new_[6778]_  : \new_[9710]_ ;
  assign \new_[5740]_  = \new_[3890]_  ? \new_[6778]_  : \new_[9120]_ ;
  assign \new_[5741]_  = \new_[2049]_  ? \new_[7858]_  : \new_[13840]_ ;
  assign \new_[5742]_  = \new_[3938]_  ? \new_[7455]_  : \new_[6854]_ ;
  assign \new_[5743]_  = \new_[3879]_  ? \new_[6778]_  : \new_[6857]_ ;
  assign \new_[5744]_  = \new_[3671]_  ? \new_[6778]_  : \new_[7306]_ ;
  assign \new_[5745]_  = ~\new_[9590]_  | ~\new_[6465]_ ;
  assign \new_[5746]_  = \\u1_u3_this_dpid_reg[0] ;
  assign \new_[5747]_  = ~\new_[7181]_  | ~\new_[6763]_ ;
  assign \new_[5748]_  = ~\new_[11275]_  | ~\new_[6464]_ ;
  assign n5190 = ~\new_[12794]_  & (~\new_[7279]_  | ~\new_[6843]_ );
  assign n5205 = ~\new_[12245]_  & (~\new_[6844]_  | ~\new_[7267]_ );
  assign n5195 = ~\new_[12732]_  & (~\new_[7268]_  | ~\new_[6845]_ );
  assign n5210 = ~\new_[12245]_  & (~\new_[6836]_  | ~\new_[7280]_ );
  assign \new_[5753]_  = \\u1_u3_next_dpid_reg[1] ;
  assign \new_[5754]_  = \\u0_u0_state_reg[10] ;
  assign \OpMode_pad_o[0]  = \\u0_u0_OpMode_reg[0] ;
  assign \new_[5756]_  = \\u4_int_srcb_reg[7] ;
  assign \new_[5757]_  = \\u4_int_srcb_reg[1] ;
  assign \wb_data_o[13]  = \\u5_wb_data_o_reg[13] ;
  assign \wb_data_o[15]  = \\u5_wb_data_o_reg[15] ;
  assign \new_[5760]_  = \\u4_u1_int_stat_reg[6] ;
  assign \new_[5761]_  = \\u4_u0_int_stat_reg[1] ;
  assign \new_[5762]_  = \\u4_u3_uc_bsel_reg[0] ;
  assign \new_[5763]_  = \\u4_u3_uc_bsel_reg[1] ;
  assign \new_[5764]_  = \\u4_u3_uc_dpd_reg[0] ;
  assign \new_[5765]_  = \\u0_u0_state_reg[6] ;
  assign \new_[5766]_  = u1_u3_buf1_set_reg;
  assign \new_[5767]_  = ~\new_[12605]_  & (~\new_[7771]_  | ~\new_[6619]_ );
  assign \new_[5768]_  = ~\new_[6555]_  & ~\new_[14191]_ ;
  assign \new_[5769]_  = ~\new_[6555]_  & ~\new_[13708]_ ;
  assign \new_[5770]_  = ~\new_[7284]_  & ~\new_[13992]_ ;
  assign n4975 = \\u1_u3_adr_reg[0] ;
  assign n5230 = \\u1_u3_adr_reg[1] ;
  assign n5200 = \\u1_u3_adr_reg[2] ;
  assign \new_[5774]_  = ~\\u1_u3_adr_reg[12] ;
  assign n4200 = \\u1_u3_adr_reg[13] ;
  assign \new_[5776]_  = ~\\u1_u3_adr_reg[14] ;
  assign \new_[5777]_  = ~\\u1_u3_adr_reg[15] ;
  assign \new_[5778]_  = ~\\u1_u3_adr_reg[16] ;
  assign n4205 = \\u1_u3_adr_reg[3] ;
  assign n4210 = \\u1_u3_adr_reg[4] ;
  assign n5225 = \\u1_u3_adr_reg[5] ;
  assign \new_[5782]_  = ~\\u1_u3_adr_reg[6] ;
  assign \new_[5783]_  = ~\\u1_u3_adr_reg[7] ;
  assign \new_[5784]_  = ~\\u1_u3_adr_reg[8] ;
  assign \new_[5785]_  = ~\\u1_u3_adr_reg[9] ;
  assign n4195 = \\u1_u3_adr_reg[10] ;
  assign \new_[5787]_  = ~\\u1_u3_adr_reg[11] ;
  assign \new_[5788]_  = ~\new_[6027]_ ;
  assign \new_[5789]_  = ~\new_[6591]_  | ~\new_[12840]_ ;
  assign n5005 = (~\new_[7406]_  & ~\new_[13760]_  & ~\new_[12849]_ ) | (~\new_[13345]_  & ~\new_[12280]_  & ~\new_[6963]_ );
  assign \new_[5791]_  = ~\new_[6523]_  & (~\new_[10029]_  | ~\new_[10856]_ );
  assign n4970 = ~\new_[7131]_  | ~\new_[7934]_  | ~\new_[7949]_  | ~\new_[8955]_ ;
  assign \new_[5793]_  = \new_[3787]_  ? \new_[6778]_  : \new_[6627]_ ;
  assign n5000 = ~\new_[7706]_  | ~\new_[7724]_  | ~\new_[6623]_ ;
  assign n5010 = \new_[6605]_  ? \new_[13120]_  : \sram_data_i[4] ;
  assign \new_[5796]_  = ~\new_[6851]_  | ~\new_[9059]_  | ~\new_[7386]_ ;
  assign \new_[5797]_  = ~\new_[6522]_  | ~\new_[2373]_ ;
  assign \new_[5798]_  = \new_[6522]_  & \new_[2477]_ ;
  assign \new_[5799]_  = \new_[6522]_  & \new_[2479]_ ;
  assign \new_[5800]_  = ~\new_[6522]_  | ~\new_[2452]_ ;
  assign \new_[5801]_  = (~\new_[6779]_  | ~\new_[4500]_ ) & (~\new_[7289]_  | ~\new_[8285]_ );
  assign \new_[5802]_  = (~\new_[6779]_  | ~\new_[4370]_ ) & (~\new_[7289]_  | ~\new_[8286]_ );
  assign \new_[5803]_  = ~\new_[6555]_  & ~\new_[13927]_ ;
  assign \new_[5804]_  = ~\new_[6540]_  | (~\new_[8233]_  & ~\new_[11733]_ );
  assign \new_[5805]_  = ~\new_[6541]_  | (~\new_[8233]_  & ~\new_[11577]_ );
  assign \new_[5806]_  = \new_[2048]_  ? \new_[6860]_  : \new_[13961]_ ;
  assign \new_[5807]_  = \new_[3102]_  ? \new_[6860]_  : \new_[13641]_ ;
  assign \new_[5808]_  = \new_[3173]_  ? \new_[6860]_  : \new_[13557]_ ;
  assign \new_[5809]_  = \new_[2178]_  ? \new_[6860]_  : \new_[14097]_ ;
  assign \new_[5810]_  = \new_[3034]_  ? \new_[6860]_  : \new_[13887]_ ;
  assign \new_[5811]_  = \new_[3021]_  ? \new_[6860]_  : \new_[14117]_ ;
  assign \new_[5812]_  = \new_[2928]_  ? \new_[6860]_  : \new_[13687]_ ;
  assign \new_[5813]_  = \new_[2856]_  ? \new_[6860]_  : \new_[14140]_ ;
  assign \new_[5814]_  = \new_[2638]_  ? \new_[6860]_  : \new_[13859]_ ;
  assign \new_[5815]_  = \new_[2639]_  ? \new_[6860]_  : \new_[13632]_ ;
  assign \new_[5816]_  = \new_[2547]_  ? \new_[6860]_  : \new_[13545]_ ;
  assign \new_[5817]_  = \new_[2265]_  ? \new_[7858]_  : \new_[13539]_ ;
  assign \new_[5818]_  = \new_[2136]_  ? \new_[6860]_  : \new_[13709]_ ;
  assign \new_[5819]_  = \new_[2075]_  ? \new_[6860]_  : \new_[13806]_ ;
  assign \new_[5820]_  = \new_[2062]_  ? \new_[6860]_  : \new_[14222]_ ;
  assign \new_[5821]_  = ~\new_[6115]_  & (~\new_[9325]_  | ~\new_[10947]_ );
  assign \new_[5822]_  = ~\new_[6683]_  | ~\new_[4774]_  | ~\new_[12143]_ ;
  assign \new_[5823]_  = ~\new_[6059]_ ;
  assign \new_[5824]_  = ~\new_[6135]_  & ~\new_[9137]_ ;
  assign \new_[5825]_  = ~\new_[6136]_  & ~\new_[9137]_ ;
  assign \new_[5826]_  = ~\new_[6137]_  & ~\new_[9137]_ ;
  assign \new_[5827]_  = ~\new_[6138]_  & ~\new_[9137]_ ;
  assign \new_[5828]_  = ~\new_[6139]_  & ~\new_[9137]_ ;
  assign \new_[5829]_  = ~\new_[6140]_  & ~\new_[9137]_ ;
  assign \new_[5830]_  = ~\new_[6141]_  & ~\new_[9137]_ ;
  assign \new_[5831]_  = ~\new_[6142]_  & ~\new_[9137]_ ;
  assign \new_[5832]_  = ~\new_[6143]_  & ~\new_[9137]_ ;
  assign \new_[5833]_  = ~\new_[6144]_  & ~\new_[9137]_ ;
  assign \new_[5834]_  = ~\new_[6145]_  & ~\new_[9137]_ ;
  assign \new_[5835]_  = ~\new_[6146]_  & ~\new_[9137]_ ;
  assign \new_[5836]_  = ~\new_[6147]_  & ~\new_[9137]_ ;
  assign \new_[5837]_  = ~\new_[6148]_  & ~\new_[9137]_ ;
  assign \new_[5838]_  = ~\new_[6149]_  & ~\new_[9137]_ ;
  assign \new_[5839]_  = ~\new_[6150]_  & ~\new_[9137]_ ;
  assign \new_[5840]_  = ~\new_[6151]_  & ~\new_[9137]_ ;
  assign \new_[5841]_  = ~\new_[3282]_  | ~\new_[6565]_  | ~\new_[7942]_ ;
  assign \new_[5842]_  = ~\new_[6152]_  & ~\new_[9137]_ ;
  assign \new_[5843]_  = ~\new_[6153]_  & ~\new_[9137]_ ;
  assign \new_[5844]_  = ~\new_[6154]_  & ~\new_[9137]_ ;
  assign \new_[5845]_  = ~\new_[6155]_  & ~\new_[9137]_ ;
  assign n5075 = ~\new_[6178]_  | ~\new_[6126]_ ;
  assign \new_[5847]_  = ~\new_[6113]_  | ~\new_[13345]_ ;
  assign \new_[5848]_  = ~\new_[8919]_  & ~\new_[6115]_ ;
  assign \new_[5849]_  = ~\new_[6118]_  & ~\new_[7190]_ ;
  assign \new_[5850]_  = \new_[2034]_  ? \new_[6860]_  : \new_[14248]_ ;
  assign \new_[5851]_  = ~\new_[14093]_  | ~\new_[6594]_ ;
  assign \new_[5852]_  = ~\new_[13566]_  | ~\new_[6594]_ ;
  assign \new_[5853]_  = ~\new_[3308]_  | ~\new_[6586]_  | ~\new_[7941]_ ;
  assign n5080 = ~n8885 & (~\new_[6684]_  | ~\new_[9809]_ );
  assign \new_[5855]_  = ~\new_[6129]_  | ~\new_[12840]_ ;
  assign \new_[5856]_  = ~\new_[6130]_  | ~\new_[12840]_ ;
  assign \new_[5857]_  = ~\new_[6132]_  | ~\new_[12840]_ ;
  assign \new_[5858]_  = ~\new_[6614]_  | ~\new_[9112]_  | ~\new_[7879]_ ;
  assign \new_[5859]_  = ~\new_[7269]_  | ~\new_[13581]_  | ~\new_[7538]_  | ~\new_[13336]_ ;
  assign \new_[5860]_  = \\u4_u3_uc_dpd_reg[1] ;
  assign n5015 = ~\new_[6110]_  & ~\new_[7411]_ ;
  assign n4990 = ~\new_[6877]_  | ~\new_[6111]_ ;
  assign n4960 = ~\new_[6112]_  & ~\new_[8124]_ ;
  assign n4985 = ~\new_[7318]_  | ~\new_[6116]_ ;
  assign n5020 = ~\new_[6117]_  & ~\new_[7414]_ ;
  assign n4980 = ~\new_[7319]_  | ~\new_[6120]_ ;
  assign n4955 = ~\new_[6121]_  & ~\new_[7418]_ ;
  assign n4995 = ~\new_[6879]_  | ~\new_[6122]_ ;
  assign n5025 = \new_[6637]_  ? \wb_addr_i[17]  : \sram_data_i[16] ;
  assign n5070 = \new_[6638]_  ? \new_[13120]_  : \sram_data_i[17] ;
  assign n5065 = \new_[6639]_  ? \wb_addr_i[17]  : \sram_data_i[18] ;
  assign n5050 = \new_[6640]_  ? \wb_addr_i[17]  : \sram_data_i[19] ;
  assign n5045 = \new_[6636]_  ? \new_[13120]_  : \sram_data_i[20] ;
  assign n5040 = \new_[6641]_  ? \new_[13120]_  : \sram_data_i[21] ;
  assign n4910 = \new_[6643]_  ? \new_[13120]_  : \sram_data_i[25] ;
  assign n4940 = \new_[6644]_  ? \wb_addr_i[17]  : \sram_data_i[26] ;
  assign n5035 = \new_[6645]_  ? \wb_addr_i[17]  : \sram_data_i[28] ;
  assign n5060 = \new_[6646]_  ? \new_[13120]_  : \sram_data_i[5] ;
  assign n5055 = \new_[6647]_  ? \new_[13120]_  : \sram_data_i[6] ;
  assign n5030 = \new_[6642]_  ? \new_[13120]_  : \sram_data_i[24] ;
  assign \new_[5881]_  = \new_[3883]_  ? \new_[6778]_  : \new_[7687]_ ;
  assign \new_[5882]_  = ~\new_[7284]_  & ~\new_[13642]_ ;
  assign \new_[5883]_  = \new_[3687]_  ? \new_[6778]_  : \new_[7405]_ ;
  assign \new_[5884]_  = \new_[3882]_  ? \new_[6778]_  : \new_[7914]_ ;
  assign \new_[5885]_  = ~\new_[7139]_  & (~\new_[6906]_  | ~\new_[3879]_ );
  assign \new_[5886]_  = ~\new_[7144]_  & (~\new_[6911]_  | ~\new_[3466]_ );
  assign n5315 = ~\new_[6698]_  & ~\new_[13386]_ ;
  assign \new_[5888]_  = ~\new_[6630]_  & (~\new_[7317]_  | ~\new_[13812]_ );
  assign \new_[5889]_  = ~\new_[6632]_  & (~\new_[7317]_  | ~\new_[13706]_ );
  assign \new_[5890]_  = ~\new_[7408]_  | ~\new_[12528]_  | ~\new_[7132]_ ;
  assign \new_[5891]_  = ~\new_[6634]_  & (~\new_[7317]_  | ~\new_[13600]_ );
  assign \new_[5892]_  = ~\new_[7413]_  | ~\new_[13470]_  | ~\new_[7133]_ ;
  assign n5300 = \new_[12190]_  & \new_[6683]_ ;
  assign \new_[5894]_  = ~\new_[12479]_  | ~\new_[6683]_ ;
  assign \new_[5895]_  = ~\new_[6850]_  | ~\new_[6683]_  | ~\new_[13575]_ ;
  assign \new_[5896]_  = \new_[2053]_  ? \new_[8233]_  : \new_[14201]_ ;
  assign \new_[5897]_  = \new_[2052]_  ? \new_[8233]_  : \new_[14207]_ ;
  assign \new_[5898]_  = \new_[2064]_  ? \new_[7309]_  : \new_[13504]_ ;
  assign \new_[5899]_  = ~\new_[6850]_  | ~\new_[6683]_  | ~\new_[14251]_ ;
  assign \new_[5900]_  = \new_[7740]_  & \new_[14418]_ ;
  assign n5355 = ~n8885 & (~\new_[6959]_  | ~\new_[7466]_ );
  assign \new_[5902]_  = ~\new_[11604]_  | ~\new_[6683]_ ;
  assign \new_[5903]_  = ~\new_[6683]_  | (~\new_[12443]_  & ~\new_[11900]_ );
  assign intb_o = u4_intb_reg;
  assign \new_[5905]_  = ~n8875 | ~\new_[12197]_  | ~\new_[11843]_  | ~\new_[7705]_ ;
  assign \new_[5906]_  = (~\new_[7289]_  | ~\new_[14245]_ ) & (~\new_[14186]_  | ~\new_[9375]_ );
  assign \new_[5907]_  = ~\new_[6654]_  & (~\new_[7317]_  | ~\new_[13670]_ );
  assign \new_[5908]_  = ~\new_[6672]_  & (~\new_[7317]_  | ~\new_[13660]_ );
  assign n5360 = \new_[7136]_  ? \new_[13120]_  : \sram_data_i[10] ;
  assign n5305 = \new_[7137]_  ? \wb_addr_i[17]  : \sram_data_i[11] ;
  assign n5310 = \new_[7138]_  ? \new_[13120]_  : \sram_data_i[9] ;
  assign \new_[5912]_  = \new_[6904]_  | \new_[6772]_ ;
  assign \new_[5913]_  = ~\new_[7449]_  | ~\new_[6633]_ ;
  assign \new_[5914]_  = \new_[6631]_  & \new_[6633]_ ;
  assign \new_[5915]_  = \new_[6673]_  | \new_[9519]_ ;
  assign \new_[5916]_  = ~\new_[6661]_  | ~\new_[6247]_ ;
  assign \new_[5917]_  = ~\new_[7323]_  | ~\new_[7361]_  | ~\new_[12865]_  | ~\new_[7434]_ ;
  assign \new_[5918]_  = ~\new_[6661]_  & ~\new_[6247]_ ;
  assign \new_[5919]_  = ~\new_[6662]_  | ~\new_[6264]_ ;
  assign \new_[5920]_  = ~\new_[7344]_  | ~\new_[7424]_  | ~\new_[12530]_  | ~\new_[7433]_ ;
  assign \new_[5921]_  = ~\new_[6662]_  & ~\new_[6264]_ ;
  assign \new_[5922]_  = ~\new_[6666]_  | ~\new_[6272]_ ;
  assign \new_[5923]_  = ~\new_[6663]_  & (~\new_[7317]_  | ~\new_[13939]_ );
  assign \new_[5924]_  = ~\new_[6666]_  & ~\new_[6272]_ ;
  assign \new_[5925]_  = ~\new_[6671]_  | ~\new_[6284]_ ;
  assign \new_[5926]_  = ~\new_[7347]_  | ~\new_[7431]_  | ~\new_[12785]_  | ~\new_[7435]_ ;
  assign \new_[5927]_  = ~\new_[6671]_  & ~\new_[6284]_ ;
  assign \new_[5928]_  = \\u1_u3_this_dpid_reg[1] ;
  assign \new_[5929]_  = ~\new_[6680]_  & (~\new_[12369]_  | ~\new_[8206]_ );
  assign \new_[5930]_  = ~\new_[6681]_  & (~\new_[12373]_  | ~\new_[8207]_ );
  assign \new_[5931]_  = ~\new_[6689]_  & (~\new_[12380]_  | ~\new_[8210]_ );
  assign \new_[5932]_  = \new_[2040]_  ? \new_[7309]_  : \new_[14190]_ ;
  assign n5235 = \new_[12009]_  ^ \new_[7169]_ ;
  assign n5240 = \new_[11967]_  ^ \new_[7170]_ ;
  assign n5245 = \new_[12198]_  ^ \new_[7171]_ ;
  assign n5250 = \new_[12127]_  ^ \new_[7175]_ ;
  assign \new_[5937]_  = ~\new_[6704]_  & ~\new_[6703]_ ;
  assign \new_[5938]_  = \new_[6704]_  & n8645;
  assign \new_[5939]_  = ~\new_[6703]_  | ~\new_[8979]_ ;
  assign n5370 = ~\new_[6779]_  & ~\new_[4781]_ ;
  assign \new_[5941]_  = ~\new_[6695]_  & ~\new_[14225]_ ;
  assign \new_[5942]_  = ~\new_[7541]_  & ~\new_[14071]_ ;
  assign \new_[5943]_  = ~\new_[7541]_  & ~\new_[14215]_ ;
  assign \new_[5944]_  = ~\new_[6695]_  & ~\new_[14100]_ ;
  assign \new_[5945]_  = ~\new_[6625]_  & ~\new_[7201]_ ;
  assign n5330 = ~\new_[6719]_  & ~n8885;
  assign \new_[5947]_  = ~\new_[7281]_  | ~\new_[7352]_  | ~\new_[9053]_ ;
  assign \new_[5948]_  = ~\new_[7287]_  | ~\new_[7353]_  | ~\new_[9056]_ ;
  assign \new_[5949]_  = ~\new_[7288]_  | ~\new_[7354]_  | ~\new_[9061]_ ;
  assign \new_[5950]_  = ~\new_[6700]_  | ~phy_rst_pad_o;
  assign \new_[5951]_  = ~\new_[7290]_  | ~\new_[7355]_  | ~\new_[9063]_ ;
  assign \new_[5952]_  = ~\new_[11805]_  | ~\new_[7471]_  | ~\new_[11448]_  | ~\new_[13655]_ ;
  assign \new_[5953]_  = ~\new_[6695]_  & ~\new_[11733]_ ;
  assign \new_[5954]_  = ~\new_[7541]_  & ~\new_[11577]_ ;
  assign \new_[5955]_  = ~\new_[7193]_  & (~\new_[7446]_  | ~\new_[7192]_ );
  assign \new_[5956]_  = ~\new_[7447]_  & (~\new_[7745]_  | ~\new_[7197]_ );
  assign \new_[5957]_  = ~\new_[7197]_  & (~\new_[7445]_  | ~\new_[7193]_ );
  assign n5325 = ~\new_[7414]_  & (~\new_[7308]_  | ~\new_[13964]_ );
  assign \new_[5959]_  = ~\new_[7143]_  & (~\new_[14787]_  | ~\new_[12488]_ );
  assign \new_[5960]_  = (~\new_[7178]_  | ~\new_[4765]_ ) & (~\new_[7436]_  | ~\new_[13844]_ );
  assign \new_[5961]_  = (~\new_[7178]_  | ~\new_[4926]_ ) & (~\new_[7436]_  | ~\new_[13977]_ );
  assign \new_[5962]_  = (~\new_[7178]_  | ~\new_[4767]_ ) & (~\new_[7436]_  | ~\new_[13823]_ );
  assign n5320 = \new_[7167]_  ? \wb_addr_i[17]  : \sram_data_i[12] ;
  assign \new_[5964]_  = (~\new_[7178]_  | ~\new_[4766]_ ) & (~\new_[7436]_  | ~\new_[14146]_ );
  assign \new_[5965]_  = (~\new_[7178]_  | ~\new_[4607]_ ) & (~\new_[7436]_  | ~\new_[13817]_ );
  assign \new_[5966]_  = ~\new_[6710]_  & (~\new_[8234]_  | ~\new_[9221]_ );
  assign \new_[5967]_  = ~\new_[6760]_  & (~\new_[7317]_  | ~\new_[14241]_ );
  assign \new_[5968]_  = \new_[3932]_  ? \new_[7455]_  : \new_[7303]_ ;
  assign \new_[5969]_  = \new_[2049]_  ? \new_[7309]_  : \new_[14162]_ ;
  assign \new_[5970]_  = ~\new_[6210]_ ;
  assign \new_[5971]_  = \new_[3283]_  ^ \new_[7293]_ ;
  assign \new_[5972]_  = \new_[3308]_  ^ \new_[7294]_ ;
  assign \new_[5973]_  = \new_[3309]_  ^ \new_[7295]_ ;
  assign n5335 = ~\new_[12849]_  & (~\new_[7472]_  | ~\new_[7264]_ );
  assign n5340 = ~\new_[12849]_  & (~\new_[7276]_  | ~\new_[7479]_ );
  assign \new_[5976]_  = \new_[3282]_  ^ \new_[7296]_ ;
  assign n5365 = ~\new_[12849]_  & (~\new_[7265]_  | ~\new_[7476]_ );
  assign \new_[5978]_  = \\u1_u0_token0_reg[6] ;
  assign n5345 = ~\new_[12732]_  & (~\new_[7478]_  | ~\new_[7275]_ );
  assign \new_[5980]_  = ~\new_[6740]_  & (~\new_[7317]_  | ~\new_[13834]_ );
  assign \new_[5981]_  = ~\new_[6220]_ ;
  assign \new_[5982]_  = ~\new_[6741]_  & (~\new_[7317]_  | ~\new_[13899]_ );
  assign \new_[5983]_  = ~\new_[6226]_ ;
  assign \new_[5984]_  = ~\new_[6775]_  & ~\new_[6776]_ ;
  assign \new_[5985]_  = ~\new_[6227]_ ;
  assign \new_[5986]_  = ~\new_[6770]_  & ~\new_[7190]_ ;
  assign \new_[5987]_  = ~\new_[6774]_  & ~\new_[6762]_ ;
  assign \new_[5988]_  = ~\new_[6773]_  & ~\new_[7193]_ ;
  assign \new_[5989]_  = ~\new_[6742]_  & (~\new_[7317]_  | ~\new_[13936]_ );
  assign \new_[5990]_  = ~\new_[6777]_  | ~\new_[7445]_ ;
  assign \new_[5991]_  = \new_[2114]_  ? \new_[7548]_  : \new_[13885]_ ;
  assign \new_[5992]_  = \new_[2076]_  ? \new_[7548]_  : \new_[13713]_ ;
  assign \new_[5993]_  = u1_u2_send_data_r_reg;
  assign \new_[5994]_  = \\u0_u0_state_reg[5] ;
  assign inta_o = u4_inta_reg;
  assign \new_[5996]_  = \new_[2082]_  ? \new_[7309]_  : \new_[14011]_ ;
  assign \new_[5997]_  = \\u0_u0_state_reg[14] ;
  assign \new_[5998]_  = \\u4_u0_csr0_reg[2] ;
  assign \new_[5999]_  = \\u4_u0_csr0_reg[4] ;
  assign \new_[6000]_  = \\u4_u0_csr1_reg[1] ;
  assign \new_[6001]_  = \\u4_u0_csr1_reg[2] ;
  assign \new_[6002]_  = \\u4_u0_csr1_reg[3] ;
  assign \new_[6003]_  = \\u4_u1_csr0_reg[2] ;
  assign \new_[6004]_  = \\u4_u1_csr0_reg[5] ;
  assign \new_[6005]_  = \\u4_u1_csr0_reg[9] ;
  assign \new_[6006]_  = ~\\u4_u1_csr1_reg[10] ;
  assign \new_[6007]_  = ~\\u4_u2_csr0_reg[0] ;
  assign \new_[6008]_  = \\u4_u2_csr0_reg[2] ;
  assign \new_[6009]_  = \\u4_u2_csr0_reg[6] ;
  assign \new_[6010]_  = \\u4_u2_csr0_reg[9] ;
  assign \new_[6011]_  = \\u4_u2_int_stat_reg[1] ;
  assign \new_[6012]_  = \\u4_u1_buf0_orig_reg[30] ;
  assign \new_[6013]_  = \\u4_u1_int_stat_reg[1] ;
  assign n9005 = u0_u0_usb_suspend_reg;
  assign \new_[6015]_  = \\u1_u0_token0_reg[0] ;
  assign \new_[6016]_  = \\u1_u0_token0_reg[1] ;
  assign \new_[6017]_  = \\u1_u0_token0_reg[3] ;
  assign \new_[6018]_  = \\u1_u0_token0_reg[4] ;
  assign \new_[6019]_  = \\u1_u0_token0_reg[5] ;
  assign \new_[6020]_  = \\u1_u0_token0_reg[7] ;
  assign \new_[6021]_  = \\u0_u0_state_reg[7] ;
  assign \new_[6022]_  = \\u0_u0_state_reg[2] ;
  assign \new_[6023]_  = u1_u3_buf0_set_reg;
  assign \new_[6024]_  = ~\new_[6695]_  & ~\new_[14191]_ ;
  assign \new_[6025]_  = ~\new_[6695]_  & ~\new_[13708]_ ;
  assign \new_[6026]_  = ~\new_[7541]_  & ~\new_[13992]_ ;
  assign \new_[6027]_  = ~\new_[13595]_  | ~\new_[10823]_  | ~\new_[7299]_ ;
  assign \new_[6028]_  = ~\new_[6763]_ ;
  assign \new_[6029]_  = \new_[3940]_  ? \new_[7455]_  : \new_[6901]_ ;
  assign n5265 = \new_[6874]_  ? n9145 : \new_[2932]_ ;
  assign \new_[6031]_  = ~\new_[7548]_  | ~\new_[7307]_  | ~\new_[7556]_ ;
  assign \new_[6032]_  = \\u4_u2_int_stat_reg[6] ;
  assign \new_[6033]_  = \\u1_u0_token0_reg[2] ;
  assign \new_[6034]_  = ~\new_[6834]_  | (~\new_[11733]_  & ~\new_[8609]_ );
  assign \new_[6035]_  = ~\new_[6837]_  | (~\new_[11577]_  & ~\new_[8609]_ );
  assign \new_[6036]_  = \new_[2265]_  ? \new_[7309]_  : \new_[13841]_ ;
  assign \new_[6037]_  = ~\new_[7541]_  & ~\new_[13927]_ ;
  assign \new_[6038]_  = \new_[2047]_  ? \new_[7548]_  : \new_[14114]_ ;
  assign \new_[6039]_  = \new_[2048]_  ? \new_[7548]_  : \new_[14235]_ ;
  assign \new_[6040]_  = \new_[2638]_  ? \new_[7309]_  : \new_[13822]_ ;
  assign \new_[6041]_  = \new_[5421]_  ? \new_[7548]_  : \new_[13603]_ ;
  assign \new_[6042]_  = \new_[9037]_  ? \new_[7548]_  : \new_[13651]_ ;
  assign \new_[6043]_  = \new_[2856]_  ? \new_[7309]_  : \new_[14055]_ ;
  assign \new_[6044]_  = \new_[2735]_  ? \new_[7548]_  : \new_[14182]_ ;
  assign \new_[6045]_  = \new_[2177]_  ? \new_[7548]_  : \new_[14068]_ ;
  assign \new_[6046]_  = \new_[9037]_  ? \new_[7309]_  : \new_[13864]_ ;
  assign \new_[6047]_  = \new_[2075]_  ? \new_[7309]_  : \new_[13818]_ ;
  assign \new_[6048]_  = \new_[3034]_  ? \new_[7309]_  : \new_[14056]_ ;
  assign \new_[6049]_  = \new_[2178]_  ? \new_[8233]_  : \new_[13686]_ ;
  assign \new_[6050]_  = \new_[5421]_  ? \new_[7309]_  : \new_[13605]_ ;
  assign \new_[6051]_  = \new_[2266]_  ? \new_[7309]_  : \new_[14250]_ ;
  assign \new_[6052]_  = \new_[2048]_  ? \new_[7309]_  : \new_[13499]_ ;
  assign \new_[6053]_  = \new_[3102]_  ? \new_[7309]_  : \new_[13729]_ ;
  assign \new_[6054]_  = \new_[3173]_  ? \new_[7309]_  : \new_[13867]_ ;
  assign \new_[6055]_  = \new_[2735]_  ? \new_[8233]_  : \new_[13994]_ ;
  assign \new_[6056]_  = \new_[2136]_  ? \new_[7309]_  : \new_[13758]_ ;
  assign \new_[6057]_  = \new_[2047]_  ? \new_[7309]_  : \new_[14240]_ ;
  assign \new_[6058]_  = ~\new_[6521]_ ;
  assign \new_[6059]_  = ~\new_[10852]_  | ~\new_[6621]_ ;
  assign n5350 = ~\new_[6615]_  & ~\new_[7411]_ ;
  assign \new_[6061]_  = ~\new_[6849]_  & (~\new_[7317]_  | ~\new_[14012]_ );
  assign n5285 = ~\new_[6616]_  & ~\new_[8124]_ ;
  assign \new_[6063]_  = \new_[6612]_  & \new_[6851]_ ;
  assign \new_[6064]_  = ~\new_[3283]_  | ~\new_[6851]_  | ~\new_[8717]_ ;
  assign \new_[6065]_  = ~\new_[13580]_  | ~\new_[6860]_ ;
  assign n5290 = ~\new_[6620]_  & ~\new_[7414]_ ;
  assign \new_[6067]_  = ~\new_[14196]_  | ~\new_[6860]_ ;
  assign \new_[6068]_  = \new_[2034]_  ? \new_[7309]_  : \new_[13843]_ ;
  assign n5295 = ~\new_[6622]_  & ~\new_[7418]_ ;
  assign \new_[6070]_  = ~\new_[2373]_  | ~\new_[11805]_  | ~\new_[12089]_  | ~\new_[7207]_ ;
  assign \new_[6071]_  = ~\new_[6883]_  | ~\new_[9646]_  | ~\new_[8036]_ ;
  assign \new_[6072]_  = ~\new_[6884]_  | ~\new_[9411]_  | ~\new_[8221]_ ;
  assign \new_[6073]_  = ~\new_[12605]_  & (~\new_[7134]_  | ~\new_[8610]_ );
  assign n5270 = ~n8885 & (~\new_[7485]_  | ~\new_[7125]_ );
  assign \new_[6075]_  = ~\new_[7320]_  | ~\new_[7605]_  | ~\new_[13044]_  | ~\new_[6267]_ ;
  assign n5275 = \new_[6910]_  ? \wb_addr_i[17]  : \sram_data_i[27] ;
  assign n5280 = \new_[6907]_  ? \wb_addr_i[17]  : \sram_data_i[29] ;
  assign n5255 = \new_[6908]_  ? \wb_addr_i[17]  : \sram_data_i[30] ;
  assign n5260 = \new_[6909]_  ? \new_[13120]_  : \sram_data_i[31] ;
  assign \new_[6080]_  = ~\new_[13417]_  | ~\new_[6624]_  | ~\new_[6912]_ ;
  assign \new_[6081]_  = ~\new_[3638]_  | ~\new_[6614]_  | ~\new_[9418]_ ;
  assign \new_[6082]_  = ~\new_[6695]_  & ~\new_[13642]_ ;
  assign \new_[6083]_  = \\u0_u0_state_reg[8] ;
  assign \new_[6084]_  = ~\new_[6101]_ ;
  assign \new_[6085]_  = ~\new_[7710]_  & (~\new_[7367]_  | ~\new_[3938]_ );
  assign \new_[6086]_  = \\u4_u3_csr1_reg[2] ;
  assign \new_[6087]_  = ~u4_u3_ots_stop_reg;
  assign \new_[6088]_  = ~\\u4_u0_buf0_orig_reg[7] ;
  assign \new_[6089]_  = \\u4_u1_csr1_reg[3] ;
  assign \new_[6090]_  = ~\\u4_u0_buf0_orig_reg[8] ;
  assign \new_[6091]_  = \\u4_u2_buf0_orig_reg[27] ;
  assign \new_[6092]_  = \\u4_u2_buf0_orig_reg[28] ;
  assign \new_[6093]_  = \\u1_u0_pid_reg[6] ;
  assign \new_[6094]_  = \\u4_dout_reg[22] ;
  assign \new_[6095]_  = \\u4_dout_reg[23] ;
  assign \new_[6096]_  = \\u4_dout_reg[7] ;
  assign \new_[6097]_  = ~\\u4_u2_buf0_orig_reg[14] ;
  assign \new_[6098]_  = ~\\u4_u1_buf0_orig_reg[13] ;
  assign \new_[6099]_  = ~\\u4_u2_buf0_orig_reg[1] ;
  assign \new_[6100]_  = ~\\u4_u1_buf0_orig_reg[0] ;
  assign \new_[6101]_  = ~\new_[6652]_ ;
  assign \new_[6102]_  = \\u4_u2_buf0_orig_reg[23] ;
  assign \new_[6103]_  = ~\\u4_u0_buf0_orig_reg[4] ;
  assign \new_[6104]_  = \new_[2053]_  ? \new_[7545]_  : \new_[13738]_ ;
  assign \new_[6105]_  = \\u4_funct_adr_reg[5] ;
  assign \new_[6106]_  = \new_[2052]_  ? \new_[7545]_  : \new_[13957]_ ;
  assign \new_[6107]_  = \\u4_funct_adr_reg[3] ;
  assign \new_[6108]_  = \new_[2064]_  ? \new_[8609]_  : \new_[13824]_ ;
  assign \new_[6109]_  = \\u4_u3_csr1_reg[6] ;
  assign \new_[6110]_  = ~\new_[5111]_  & (~\new_[7370]_  | ~\new_[8633]_ );
  assign \new_[6111]_  = ~\new_[6956]_  | ~\new_[9780]_ ;
  assign \new_[6112]_  = ~\new_[4970]_  & (~\new_[7370]_  | ~\new_[8970]_ );
  assign \new_[6113]_  = ~\new_[11924]_  & ~\new_[6963]_ ;
  assign \new_[6114]_  = ~\new_[8161]_  & (~\new_[7401]_  | ~\new_[3481]_ );
  assign \new_[6115]_  = ~\new_[13956]_  | ~\new_[13265]_  | ~\new_[7400]_ ;
  assign \new_[6116]_  = ~\new_[7016]_  | ~\new_[9784]_ ;
  assign \new_[6117]_  = ~\new_[5112]_  & (~\new_[7370]_  | ~\new_[7866]_ );
  assign \new_[6118]_  = \new_[8417]_  & \new_[7189]_ ;
  assign \new_[6119]_  = ~\new_[6621]_ ;
  assign \new_[6120]_  = ~\new_[7070]_  | ~\new_[9796]_ ;
  assign \new_[6121]_  = ~\new_[4966]_  & (~\new_[7370]_  | ~\new_[8247]_ );
  assign \new_[6122]_  = ~\new_[7123]_  | ~\new_[9792]_ ;
  assign n5435 = ~\new_[6963]_  & (~\new_[9497]_  | ~\new_[14004]_ );
  assign n5430 = ~\new_[6963]_  & (~\new_[10102]_  | ~\new_[13790]_ );
  assign n5385 = ~\new_[6963]_  & (~\new_[9890]_  | ~\new_[13599]_ );
  assign \new_[6126]_  = n8875 | \new_[13296]_  | \new_[11843]_  | \new_[7406]_ ;
  assign \new_[6127]_  = \new_[7187]_  & \new_[14548]_ ;
  assign \new_[6128]_  = \new_[4291]_  ? \new_[7455]_  : \new_[9919]_ ;
  assign \new_[6129]_  = \new_[4073]_  ? \new_[7455]_  : \new_[9070]_ ;
  assign \new_[6130]_  = \new_[4070]_  ? \new_[7455]_  : \new_[8706]_ ;
  assign \new_[6131]_  = \new_[4237]_  ? \new_[7455]_  : \new_[9381]_ ;
  assign \new_[6132]_  = \new_[4074]_  ? \new_[7455]_  : \new_[8705]_ ;
  assign \new_[6133]_  = \new_[4347]_  ? \new_[7455]_  : \new_[8707]_ ;
  assign \new_[6134]_  = \new_[6904]_  | \new_[7182]_ ;
  assign \new_[6135]_  = (~\new_[7317]_  | ~\new_[13717]_ ) & (~\new_[7844]_  | ~\new_[2266]_ );
  assign \new_[6136]_  = (~\new_[7317]_  | ~\new_[13772]_ ) & (~\new_[7844]_  | ~\new_[2047]_ );
  assign \new_[6137]_  = (~\new_[7317]_  | ~\new_[13731]_ ) & (~\new_[7844]_  | ~\new_[2048]_ );
  assign \new_[6138]_  = (~\new_[7317]_  | ~\new_[13736]_ ) & (~\new_[7844]_  | ~\new_[5421]_ );
  assign \new_[6139]_  = (~\new_[7317]_  | ~\new_[13549]_ ) & (~\new_[7844]_  | ~\new_[3102]_ );
  assign \new_[6140]_  = (~\new_[7317]_  | ~\new_[13648]_ ) & (~\new_[7844]_  | ~\new_[3173]_ );
  assign \new_[6141]_  = (~\new_[7317]_  | ~\new_[14048]_ ) & (~\new_[7844]_  | ~\new_[2178]_ );
  assign \new_[6142]_  = (~\new_[7317]_  | ~\new_[14023]_ ) & (~\new_[7844]_  | ~\new_[3034]_ );
  assign \new_[6143]_  = (~\new_[7317]_  | ~\new_[13942]_ ) & (~\new_[7844]_  | ~\new_[3021]_ );
  assign \new_[6144]_  = (~\new_[7317]_  | ~\new_[13826]_ ) & (~\new_[7844]_  | ~\new_[9037]_ );
  assign \new_[6145]_  = (~\new_[7317]_  | ~\new_[14262]_ ) & (~\new_[7844]_  | ~\new_[2928]_ );
  assign \new_[6146]_  = (~\new_[7317]_  | ~\new_[13911]_ ) & (~\new_[7844]_  | ~\new_[2856]_ );
  assign \new_[6147]_  = (~\new_[7317]_  | ~\new_[14025]_ ) & (~\new_[7844]_  | ~\new_[2638]_ );
  assign \new_[6148]_  = (~\new_[7317]_  | ~\new_[14253]_ ) & (~\new_[7844]_  | ~\new_[2639]_ );
  assign \new_[6149]_  = (~\new_[7317]_  | ~\new_[14234]_ ) & (~\new_[7844]_  | ~\new_[2547]_ );
  assign \new_[6150]_  = (~\new_[7317]_  | ~\new_[13860]_ ) & (~\new_[7844]_  | ~\new_[2735]_ );
  assign \new_[6151]_  = (~\new_[7317]_  | ~\new_[13592]_ ) & (~\new_[7844]_  | ~\new_[2177]_ );
  assign \new_[6152]_  = (~\new_[7317]_  | ~\new_[13727]_ ) & (~\new_[7844]_  | ~\new_[2265]_ );
  assign \new_[6153]_  = (~\new_[7317]_  | ~\new_[14193]_ ) & (~\new_[7844]_  | ~\new_[2136]_ );
  assign \new_[6154]_  = (~\new_[7317]_  | ~\new_[13873]_ ) & (~\new_[7844]_  | ~\new_[2075]_ );
  assign \new_[6155]_  = (~\new_[7317]_  | ~\new_[13724]_ ) & (~\new_[7844]_  | ~\new_[2062]_ );
  assign \new_[6156]_  = (~\new_[7782]_  | ~\new_[14053]_ ) & (~\new_[7482]_  | ~\new_[13873]_ );
  assign \new_[6157]_  = ~\\u4_u2_buf0_orig_reg[16] ;
  assign \new_[6158]_  = \new_[2040]_  ? \new_[7545]_  : \new_[14072]_ ;
  assign \new_[6159]_  = \\u4_dout_reg[8] ;
  assign \new_[6160]_  = ~\\u4_u0_buf0_orig_reg[6] ;
  assign \new_[6161]_  = \new_[4286]_  ? \new_[7455]_  : \new_[8165]_ ;
  assign \new_[6162]_  = \new_[4236]_  ? \new_[7455]_  : \new_[7458]_ ;
  assign \new_[6163]_  = \\u4_u3_csr1_reg[10] ;
  assign \new_[6164]_  = (~\new_[7781]_  | ~\new_[4794]_ ) & (~\new_[7482]_  | ~\new_[5764]_ );
  assign \new_[6165]_  = ~\\u4_u0_buf0_orig_reg[31] ;
  assign \new_[6166]_  = \\u4_u1_csr0_reg[8] ;
  assign n5455 = ~\new_[7145]_  & ~\new_[7414]_ ;
  assign \new_[6168]_  = \\u4_u0_buf0_orig_reg[20] ;
  assign \new_[6169]_  = ~\\u4_u1_csr1_reg[1] ;
  assign \new_[6170]_  = \\u1_u0_pid_reg[7] ;
  assign \new_[6171]_  = ~\new_[7486]_  & (~\new_[7480]_  | ~\new_[9097]_ );
  assign \new_[6172]_  = \\u4_u1_csr1_reg[11] ;
  assign \new_[6173]_  = \new_[2114]_  ? \new_[7858]_  : \new_[13737]_ ;
  assign \new_[6174]_  = ~\new_[14477]_ ;
  assign \new_[6175]_  = ~\new_[7743]_  | ~\new_[7742]_  | ~\new_[13397]_  | ~\new_[14450]_ ;
  assign \new_[6176]_  = \new_[2076]_  ? \new_[7858]_  : \new_[14083]_ ;
  assign \new_[6177]_  = ~\new_[13165]_  | ~\new_[7705]_  | ~\new_[4778]_ ;
  assign \new_[6178]_  = ~\new_[13165]_  | ~\new_[7705]_  | ~\new_[5123]_ ;
  assign \new_[6179]_  = ~\new_[13165]_  | ~\new_[7705]_  | ~\new_[4501]_ ;
  assign \new_[6180]_  = ~\new_[7442]_  & (~\new_[7447]_  | ~\new_[7443]_ );
  assign n5450 = ~\new_[7418]_  & (~\new_[7552]_  | ~\new_[13661]_ );
  assign \new_[6182]_  = ~\new_[7141]_  & (~\new_[8568]_  | ~\new_[9889]_ );
  assign \new_[6183]_  = ~\new_[7142]_  & (~\new_[8568]_  | ~\new_[9361]_ );
  assign \new_[6184]_  = ~\new_[7176]_  & ~\new_[6166]_ ;
  assign \new_[6185]_  = (~\new_[8224]_  & ~\new_[13319]_ ) | (~\new_[14586]_  & ~\new_[2874]_ );
  assign \new_[6186]_  = \new_[4095]_  ? \new_[7455]_  : \new_[11734]_ ;
  assign n5440 = \new_[7427]_  ? \new_[13120]_  : \sram_data_i[13] ;
  assign n5445 = \new_[7428]_  ? \wb_addr_i[17]  : \sram_data_i[15] ;
  assign \new_[6189]_  = \new_[4292]_  ? \new_[7455]_  : \new_[10768]_ ;
  assign \new_[6190]_  = \new_[4293]_  ? \new_[7455]_  : \new_[10697]_ ;
  assign \new_[6191]_  = \new_[4206]_  ? \new_[7455]_  : \new_[9881]_ ;
  assign \new_[6192]_  = \new_[4098]_  ? \new_[7455]_  : \new_[12887]_ ;
  assign \new_[6193]_  = \new_[4096]_  ? \new_[7455]_  : \new_[11703]_ ;
  assign \new_[6194]_  = \new_[3997]_  ? \new_[7455]_  : \new_[9705]_ ;
  assign \new_[6195]_  = \new_[4197]_  ? \new_[7455]_  : \new_[9114]_ ;
  assign \new_[6196]_  = \\u4_u3_csr0_reg[7] ;
  assign \new_[6197]_  = \new_[4097]_  ? \new_[7455]_  : \new_[9969]_ ;
  assign \new_[6198]_  = \\u4_u0_buf0_orig_reg[28] ;
  assign \new_[6199]_  = \new_[2049]_  ? \new_[7545]_  : \new_[14090]_ ;
  assign \new_[6200]_  = \\u4_u1_csr0_reg[6] ;
  assign n5420 = ~n8885 & (~\new_[7484]_  | ~\new_[9073]_ );
  assign \new_[6202]_  = ~\new_[7178]_  | ~\new_[14115]_ ;
  assign \new_[6203]_  = ~\\u4_u1_csr0_reg[12] ;
  assign \new_[6204]_  = (~\new_[7765]_  | ~\new_[13815]_ ) & (~\new_[7469]_  | ~\new_[12493]_ );
  assign \new_[6205]_  = (~\new_[7765]_  | ~\new_[13932]_ ) & (~\new_[7469]_  | ~\new_[11054]_ );
  assign \new_[6206]_  = ~\new_[7178]_  | ~\new_[2038]_ ;
  assign \new_[6207]_  = ~\new_[7178]_  | ~\new_[13561]_ ;
  assign \new_[6208]_  = (~\new_[7781]_  | ~\new_[14247]_ ) & (~\new_[7482]_  | ~\new_[13898]_ );
  assign \new_[6209]_  = ~\\u4_u2_buf0_orig_reg[10] ;
  assign \new_[6210]_  = \new_[14283]_  | \new_[14634]_ ;
  assign \new_[6211]_  = ~\\u4_u2_buf0_orig_reg[12] ;
  assign \new_[6212]_  = \new_[2114]_  ? \new_[8609]_  : \new_[13513]_ ;
  assign n5460 = ~\new_[12245]_  & (~\new_[7768]_  | ~\new_[7473]_ );
  assign n5465 = ~\new_[12849]_  & (~\new_[7769]_  | ~\new_[7477]_ );
  assign n5470 = ~\new_[12505]_  & (~\new_[7774]_  | ~\new_[7474]_ );
  assign \new_[6216]_  = \new_[2076]_  ? \new_[7545]_  : \new_[13966]_ ;
  assign \new_[6217]_  = \new_[2082]_  ? \new_[7545]_  : \new_[13984]_ ;
  assign n5570 = ~\new_[12505]_  & (~\new_[7770]_  | ~\new_[7475]_ );
  assign \new_[6219]_  = ~\new_[13595]_  | ~\new_[9162]_  | ~\new_[7470]_ ;
  assign \new_[6220]_  = ~\new_[7443]_  | ~\new_[7191]_ ;
  assign \new_[6221]_  = ~\new_[7744]_  | ~\new_[7192]_ ;
  assign \new_[6222]_  = ~\new_[6705]_ ;
  assign \new_[6223]_  = ~\new_[7442]_  | ~\new_[7191]_ ;
  assign \new_[6224]_  = ~\new_[7192]_  | ~\new_[7445]_ ;
  assign \new_[6225]_  = ~\new_[6706]_ ;
  assign \new_[6226]_  = \new_[7181]_  & \new_[7744]_ ;
  assign \new_[6227]_  = ~\new_[7449]_  | ~\new_[7196]_ ;
  assign \new_[6228]_  = ~\new_[7194]_  | ~\new_[7745]_ ;
  assign \new_[6229]_  = ~\new_[7188]_  | ~\new_[7443]_ ;
  assign \new_[6230]_  = ~\new_[7191]_  | ~\new_[7182]_ ;
  assign \new_[6231]_  = ~\new_[6717]_ ;
  assign \new_[6232]_  = \\u4_u0_buf0_orig_reg[22] ;
  assign \new_[6233]_  = \\u1_u2_state_reg[6] ;
  assign \new_[6234]_  = \\u4_u0_buf0_orig_reg[26] ;
  assign \new_[6235]_  = \\u1_u2_state_reg[1] ;
  assign \new_[6236]_  = \\u1_u2_state_reg[5] ;
  assign \new_[6237]_  = \\u4_u1_csr0_reg[1] ;
  assign \new_[6238]_  = \\u4_u0_buf0_orig_reg[24] ;
  assign \new_[6239]_  = \\u4_funct_adr_reg[0] ;
  assign \new_[6240]_  = \\u4_funct_adr_reg[1] ;
  assign \new_[6241]_  = \\u4_funct_adr_reg[2] ;
  assign \new_[6242]_  = \\u4_funct_adr_reg[4] ;
  assign \new_[6243]_  = \\u4_funct_adr_reg[6] ;
  assign n9145 = u1_u3_out_to_small_r_reg;
  assign \new_[6245]_  = ~u4_u2_ots_stop_reg;
  assign \new_[6246]_  = u1_u2_mack_r_reg;
  assign \new_[6247]_  = \\u4_u3_csr0_reg[10] ;
  assign \new_[6248]_  = ~\\u4_u3_csr0_reg[12] ;
  assign \new_[6249]_  = \\u4_u3_csr0_reg[1] ;
  assign \new_[6250]_  = \\u4_u3_csr0_reg[2] ;
  assign \new_[6251]_  = \\u4_u3_csr0_reg[4] ;
  assign \new_[6252]_  = \\u4_u3_csr0_reg[5] ;
  assign \new_[6253]_  = \\u4_u3_csr0_reg[6] ;
  assign \new_[6254]_  = \\u4_u3_csr0_reg[8] ;
  assign \new_[6255]_  = \\u4_u3_csr0_reg[9] ;
  assign \new_[6256]_  = \\u4_u3_csr1_reg[0] ;
  assign \new_[6257]_  = \\u4_u3_csr1_reg[11] ;
  assign \new_[6258]_  = \\u4_u3_csr1_reg[12] ;
  assign \new_[6259]_  = \\u4_u3_csr1_reg[1] ;
  assign \new_[6260]_  = \\u4_u3_csr1_reg[3] ;
  assign \new_[6261]_  = \\u4_u3_csr1_reg[4] ;
  assign \new_[6262]_  = \\u4_u3_csr1_reg[5] ;
  assign \new_[6263]_  = \\u4_u3_csr1_reg[9] ;
  assign \new_[6264]_  = \\u4_u0_csr0_reg[10] ;
  assign \new_[6265]_  = ~\\u4_u0_csr0_reg[12] ;
  assign \new_[6266]_  = \\u4_u0_csr0_reg[6] ;
  assign \new_[6267]_  = \\u4_u0_csr1_reg[0] ;
  assign \new_[6268]_  = \\u4_u0_csr1_reg[5] ;
  assign \new_[6269]_  = \\u4_u0_csr1_reg[9] ;
  assign \new_[6270]_  = ~u4_u0_ots_stop_reg;
  assign \new_[6271]_  = ~\\u4_u1_csr0_reg[0] ;
  assign \new_[6272]_  = \\u4_u1_csr0_reg[10] ;
  assign \new_[6273]_  = ~\\u4_u1_csr0_reg[11] ;
  assign \new_[6274]_  = \\u4_u1_csr0_reg[4] ;
  assign \new_[6275]_  = \\u4_u1_csr0_reg[7] ;
  assign \new_[6276]_  = \\u4_u1_csr1_reg[0] ;
  assign \new_[6277]_  = \\u4_u1_csr1_reg[12] ;
  assign \new_[6278]_  = ~\\u4_u1_csr1_reg[2] ;
  assign \new_[6279]_  = \\u4_u1_csr1_reg[4] ;
  assign \new_[6280]_  = \\u4_u1_csr1_reg[5] ;
  assign \new_[6281]_  = \\u4_u1_csr1_reg[6] ;
  assign \new_[6282]_  = ~\\u4_u1_csr1_reg[9] ;
  assign \new_[6283]_  = ~u4_u1_ots_stop_reg;
  assign \new_[6284]_  = \\u4_u2_csr0_reg[10] ;
  assign \new_[6285]_  = ~\\u4_u2_csr0_reg[12] ;
  assign \new_[6286]_  = \\u4_u2_csr0_reg[4] ;
  assign \new_[6287]_  = \\u4_u2_csr0_reg[7] ;
  assign \new_[6288]_  = \\u4_u2_csr1_reg[0] ;
  assign \new_[6289]_  = \\u4_u2_csr1_reg[11] ;
  assign \new_[6290]_  = \\u4_u2_csr1_reg[1] ;
  assign \new_[6291]_  = \\u4_u2_csr1_reg[3] ;
  assign \new_[6292]_  = \\u4_u2_csr1_reg[6] ;
  assign \new_[6293]_  = \\u4_u2_csr1_reg[5] ;
  assign \new_[6294]_  = ~\\u4_u3_buf0_orig_reg[0] ;
  assign \new_[6295]_  = ~\\u4_u3_buf0_orig_reg[12] ;
  assign \new_[6296]_  = ~\\u4_u3_buf0_orig_reg[14] ;
  assign \new_[6297]_  = ~\\u4_u3_buf0_orig_reg[15] ;
  assign \new_[6298]_  = ~\\u4_u3_buf0_orig_reg[16] ;
  assign \new_[6299]_  = \\u4_u3_buf0_orig_reg[21] ;
  assign \new_[6300]_  = \\u4_u3_buf0_orig_reg[22] ;
  assign \new_[6301]_  = \\u4_u3_buf0_orig_reg[23] ;
  assign \new_[6302]_  = \\u4_u3_buf0_orig_reg[24] ;
  assign \new_[6303]_  = \\u4_u3_buf0_orig_reg[26] ;
  assign \new_[6304]_  = \\u4_u3_buf0_orig_reg[28] ;
  assign \new_[6305]_  = \\u4_u3_buf0_orig_reg[30] ;
  assign \new_[6306]_  = ~\\u4_u3_buf0_orig_reg[31] ;
  assign \new_[6307]_  = ~\\u4_u3_buf0_orig_reg[5] ;
  assign \new_[6308]_  = ~\\u4_u3_buf0_orig_reg[8] ;
  assign \new_[6309]_  = ~\\u4_u3_csr1_reg[8] ;
  assign \new_[6310]_  = \\u4_u3_int_stat_reg[1] ;
  assign \new_[6311]_  = ~\\u4_u0_buf0_orig_reg[10] ;
  assign \new_[6312]_  = ~\\u4_u0_buf0_orig_reg[11] ;
  assign \new_[6313]_  = ~\\u4_u0_buf0_orig_reg[12] ;
  assign \new_[6314]_  = (~\new_[7781]_  | ~\new_[4788]_ ) & (~\new_[7481]_  | ~\new_[6256]_ );
  assign \new_[6315]_  = ~\\u4_u0_buf0_orig_reg[14] ;
  assign \new_[6316]_  = ~\\u4_u0_buf0_orig_reg[16] ;
  assign \new_[6317]_  = ~\\u4_u0_buf0_orig_reg[18] ;
  assign \new_[6318]_  = ~\\u4_u0_buf0_orig_reg[1] ;
  assign \new_[6319]_  = \\u4_u0_buf0_orig_reg[21] ;
  assign \new_[6320]_  = \\u4_u0_buf0_orig_reg[23] ;
  assign \new_[6321]_  = (~\new_[7783]_  | ~\new_[13878]_ ) & (~\new_[7482]_  | ~\new_[6259]_ );
  assign \new_[6322]_  = \\u4_u0_buf0_orig_reg[25] ;
  assign \new_[6323]_  = \\u4_u0_buf0_orig_reg[27] ;
  assign \new_[6324]_  = \\u4_u0_buf0_orig_reg[29] ;
  assign \new_[6325]_  = ~\\u4_u0_buf0_orig_reg[2] ;
  assign \new_[6326]_  = \\u4_u0_buf0_orig_reg[30] ;
  assign \new_[6327]_  = ~\\u4_u0_buf0_orig_reg[3] ;
  assign \new_[6328]_  = ~\\u4_u0_buf0_orig_reg[5] ;
  assign \new_[6329]_  = (~\new_[7781]_  | ~\new_[4841]_ ) & (~\new_[7481]_  | ~\new_[14253]_ );
  assign \new_[6330]_  = ~\\u4_u0_buf0_orig_reg[9] ;
  assign \new_[6331]_  = ~\\u4_u3_buf0_orig_reg[9] ;
  assign \new_[6332]_  = ~\\u4_u0_csr1_reg[8] ;
  assign \new_[6333]_  = (~\new_[7781]_  | ~\new_[13963]_ ) & (~\new_[7482]_  | ~\new_[6086]_ );
  assign \new_[6334]_  = ~\\u4_u1_buf0_orig_reg[10] ;
  assign \new_[6335]_  = ~\\u4_u1_buf0_orig_reg[11] ;
  assign \new_[6336]_  = ~\\u4_u1_buf0_orig_reg[12] ;
  assign \new_[6337]_  = ~\\u4_u1_buf0_orig_reg[14] ;
  assign \new_[6338]_  = ~\\u4_u1_buf0_orig_reg[15] ;
  assign \new_[6339]_  = ~\\u4_u1_buf0_orig_reg[16] ;
  assign \new_[6340]_  = ~\\u4_u1_buf0_orig_reg[18] ;
  assign \new_[6341]_  = \\u4_u1_buf0_orig_reg[19] ;
  assign \new_[6342]_  = ~\\u4_u1_buf0_orig_reg[1] ;
  assign \new_[6343]_  = \\u4_u1_buf0_orig_reg[21] ;
  assign \new_[6344]_  = \\u4_u1_buf0_orig_reg[22] ;
  assign \new_[6345]_  = \\u4_u1_buf0_orig_reg[23] ;
  assign \new_[6346]_  = \\u4_u1_buf0_orig_reg[25] ;
  assign \new_[6347]_  = \\u4_u1_buf0_orig_reg[26] ;
  assign \new_[6348]_  = \\u4_u1_buf0_orig_reg[27] ;
  assign \new_[6349]_  = (~\new_[7783]_  | ~\new_[4615]_ ) & (~\new_[7482]_  | ~\new_[6249]_ );
  assign \new_[6350]_  = ~\\u4_u1_buf0_orig_reg[2] ;
  assign \new_[6351]_  = \\u4_u1_buf0_orig_reg[29] ;
  assign \new_[6352]_  = ~\\u4_u1_buf0_orig_reg[3] ;
  assign \new_[6353]_  = ~\\u4_u1_buf0_orig_reg[4] ;
  assign \new_[6354]_  = ~\\u4_u1_buf0_orig_reg[5] ;
  assign \new_[6355]_  = ~\\u4_u1_buf0_orig_reg[7] ;
  assign \new_[6356]_  = (~\new_[7782]_  | ~\new_[4790]_ ) & (~\new_[7482]_  | ~\new_[13533]_ );
  assign \new_[6357]_  = ~\\u4_u1_csr1_reg[8] ;
  assign \new_[6358]_  = ~\\u4_u2_buf0_orig_reg[0] ;
  assign \new_[6359]_  = ~\\u4_u2_buf0_orig_reg[11] ;
  assign \new_[6360]_  = (~\new_[7783]_  | ~\new_[4768]_ ) & (~\new_[7482]_  | ~\new_[13902]_ );
  assign \new_[6361]_  = ~\\u4_u2_buf0_orig_reg[13] ;
  assign \new_[6362]_  = ~\\u4_u2_buf0_orig_reg[15] ;
  assign \new_[6363]_  = ~\\u4_u2_buf0_orig_reg[17] ;
  assign \new_[6364]_  = ~\\u4_u2_buf0_orig_reg[18] ;
  assign \new_[6365]_  = \\u4_u2_buf0_orig_reg[19] ;
  assign \new_[6366]_  = \\u4_u2_buf0_orig_reg[20] ;
  assign \new_[6367]_  = \\u4_u2_buf0_orig_reg[21] ;
  assign \new_[6368]_  = \\u4_u2_buf0_orig_reg[22] ;
  assign \new_[6369]_  = \\u4_u2_buf0_orig_reg[24] ;
  assign \new_[6370]_  = \\u4_u2_buf0_orig_reg[25] ;
  assign \new_[6371]_  = \\u4_u2_buf0_orig_reg[26] ;
  assign \new_[6372]_  = (~\new_[7781]_  | ~\new_[4792]_ ) & (~\new_[7482]_  | ~\new_[6163]_ );
  assign \new_[6373]_  = ~\\u4_u2_buf0_orig_reg[2] ;
  assign \new_[6374]_  = ~\\u4_u2_buf0_orig_reg[31] ;
  assign \new_[6375]_  = ~\\u4_u2_buf0_orig_reg[4] ;
  assign \new_[6376]_  = (~\new_[7483]_  | ~\new_[12778]_ ) & (~\new_[8214]_  | ~\new_[6257]_ );
  assign \new_[6377]_  = ~\\u4_u2_buf0_orig_reg[7] ;
  assign \new_[6378]_  = ~\\u4_u2_buf0_orig_reg[9] ;
  assign \new_[6379]_  = ~\\u4_u2_csr1_reg[8] ;
  assign \wb_data_o[14]  = \\u5_wb_data_o_reg[14] ;
  assign \new_[6381]_  = (~\new_[7782]_  | ~\new_[4795]_ ) & (~\new_[7482]_  | ~\new_[5860]_ );
  assign \new_[6382]_  = (~\new_[7483]_  | ~\new_[13284]_ ) & (~\new_[7481]_  | ~\new_[5762]_ );
  assign \new_[6383]_  = \\u1_u0_pid_reg[0] ;
  assign \new_[6384]_  = \\u1_u0_pid_reg[1] ;
  assign \new_[6385]_  = \\u1_u0_pid_reg[2] ;
  assign \new_[6386]_  = \\u1_u0_pid_reg[4] ;
  assign \new_[6387]_  = \\u1_u0_pid_reg[5] ;
  assign \new_[6388]_  = (~\new_[7781]_  | ~\new_[13862]_ ) & (~\new_[7482]_  | ~\new_[5763]_ );
  assign \new_[6389]_  = (~\new_[7783]_  | ~\new_[4798]_ ) & (~\new_[7482]_  | ~\new_[6743]_ );
  assign \new_[6390]_  = (~\new_[7781]_  | ~\new_[12760]_ ) & (~\new_[7481]_  | ~\new_[6251]_ );
  assign \new_[6391]_  = (~\new_[7782]_  | ~\new_[4801]_ ) & (~\new_[7482]_  | ~\new_[6196]_ );
  assign \new_[6392]_  = (~\new_[7782]_  | ~\new_[4802]_ ) & (~\new_[7482]_  | ~\new_[6254]_ );
  assign \new_[6393]_  = (~\new_[7781]_  | ~\new_[4651]_ ) & (~\new_[8214]_  | ~\new_[6255]_ );
  assign \new_[6394]_  = (~\new_[7783]_  | ~\new_[13576]_ ) & (~\new_[7482]_  | ~\new_[13600]_ );
  assign \new_[6395]_  = (~\new_[7781]_  | ~\new_[4791]_ ) & (~\new_[7482]_  | ~\new_[6263]_ );
  assign \new_[6396]_  = (~\new_[7782]_  | ~\new_[4842]_ ) & (~\new_[7482]_  | ~\new_[14234]_ );
  assign \new_[6397]_  = (~\new_[7781]_  | ~\new_[4812]_ ) & (~\new_[8214]_  | ~\new_[14007]_ );
  assign \new_[6398]_  = (~\new_[7483]_  | ~\new_[4817]_ ) & (~\new_[8214]_  | ~\new_[13743]_ );
  assign \new_[6399]_  = (~\new_[7781]_  | ~\new_[4620]_ ) & (~\new_[7481]_  | ~\new_[6252]_ );
  assign \new_[6400]_  = (~\new_[7783]_  | ~\new_[13601]_ ) & (~\new_[7482]_  | ~\new_[14189]_ );
  assign \new_[6401]_  = (~\new_[7783]_  | ~\new_[14019]_ ) & (~\new_[7482]_  | ~\new_[14090]_ );
  assign \new_[6402]_  = (~\new_[7783]_  | ~\new_[13654]_ ) & (~\new_[7482]_  | ~\new_[13738]_ );
  assign \new_[6403]_  = (~\new_[7783]_  | ~\new_[13921]_ ) & (~\new_[7482]_  | ~\new_[13665]_ );
  assign \new_[6404]_  = (~\new_[7783]_  | ~\new_[13502]_ ) & (~\new_[7482]_  | ~\new_[13537]_ );
  assign \new_[6405]_  = (~\new_[7783]_  | ~\new_[13594]_ ) & (~\new_[7482]_  | ~\new_[14072]_ );
  assign \new_[6406]_  = (~\new_[7782]_  | ~\new_[13999]_ ) & (~\new_[7482]_  | ~\new_[13957]_ );
  assign \new_[6407]_  = (~\new_[8215]_  | ~\new_[4811]_ ) & (~\new_[7481]_  | ~\new_[13554]_ );
  assign \new_[6408]_  = (~\new_[7782]_  | ~\new_[4864]_ ) & (~\new_[7482]_  | ~\new_[13954]_ );
  assign \new_[6409]_  = (~\new_[7781]_  | ~\new_[13508]_ ) & (~\new_[7482]_  | ~\new_[13618]_ );
  assign \new_[6410]_  = (~\new_[8215]_  | ~\new_[4814]_ ) & (~\new_[7481]_  | ~\new_[13820]_ );
  assign \new_[6411]_  = (~\new_[7483]_  | ~\new_[4695]_ ) & (~\new_[8214]_  | ~\new_[13910]_ );
  assign \new_[6412]_  = (~\new_[7483]_  | ~\new_[4815]_ ) & (~\new_[7481]_  | ~\new_[13972]_ );
  assign \new_[6413]_  = (~\new_[8215]_  | ~\new_[4816]_ ) & (~\new_[7481]_  | ~\new_[13625]_ );
  assign \new_[6414]_  = (~\new_[7483]_  | ~\new_[4709]_ ) & (~\new_[7481]_  | ~\new_[14177]_ );
  assign \new_[6415]_  = (~\new_[7483]_  | ~\new_[4818]_ ) & (~\new_[7481]_  | ~\new_[14136]_ );
  assign \new_[6416]_  = (~\new_[7782]_  | ~\new_[4819]_ ) & (~\new_[7482]_  | ~\new_[13776]_ );
  assign \new_[6417]_  = (~\new_[7783]_  | ~\new_[4820]_ ) & (~\new_[7482]_  | ~\new_[14227]_ );
  assign \new_[6418]_  = (~\new_[7782]_  | ~\new_[4676]_ ) & (~\new_[7482]_  | ~\new_[13777]_ );
  assign \new_[6419]_  = (~\new_[7782]_  | ~\new_[13801]_ ) & (~\new_[7482]_  | ~\new_[13551]_ );
  assign \new_[6420]_  = (~\new_[8215]_  | ~\new_[4690]_ ) & (~\new_[7482]_  | ~\new_[14044]_ );
  assign \new_[6421]_  = (~\new_[8215]_  | ~\new_[14037]_ ) & (~\new_[7482]_  | ~\new_[14134]_ );
  assign \new_[6422]_  = (~\new_[8215]_  | ~\new_[14124]_ ) & (~\new_[7482]_  | ~\new_[13706]_ );
  assign \new_[6423]_  = (~\new_[7781]_  | ~\new_[13785]_ ) & (~\new_[7482]_  | ~\new_[13745]_ );
  assign \new_[6424]_  = ~\new_[7639]_  | ~\new_[8655]_  | ~\new_[12446]_  | ~\new_[7594]_ ;
  assign \new_[6425]_  = (~\new_[7781]_  | ~\new_[13523]_ ) & (~\new_[7482]_  | ~\new_[13513]_ );
  assign \new_[6426]_  = (~\new_[7782]_  | ~\new_[14051]_ ) & (~\new_[7482]_  | ~\new_[13966]_ );
  assign \new_[6427]_  = (~\new_[7782]_  | ~\new_[13526]_ ) & (~\new_[7482]_  | ~\new_[13824]_ );
  assign \new_[6428]_  = (~\new_[7782]_  | ~\new_[13990]_ ) & (~\new_[7482]_  | ~\new_[13984]_ );
  assign \new_[6429]_  = (~\new_[7782]_  | ~\new_[13505]_ ) & (~\new_[7482]_  | ~\new_[14144]_ );
  assign \new_[6430]_  = (~\new_[7782]_  | ~\new_[13628]_ ) & (~\new_[7482]_  | ~\new_[13684]_ );
  assign \new_[6431]_  = (~\new_[7783]_  | ~\new_[13723]_ ) & (~\new_[7482]_  | ~\new_[13717]_ );
  assign \new_[6432]_  = ~\new_[7622]_  | ~\new_[8653]_  | ~\new_[12483]_  | ~\new_[7593]_ ;
  assign \new_[6433]_  = (~\new_[7782]_  | ~\new_[13530]_ ) & (~\new_[7482]_  | ~\new_[13812]_ );
  assign \new_[6434]_  = (~\new_[7781]_  | ~\new_[13531]_ ) & (~\new_[7482]_  | ~\new_[13772]_ );
  assign \new_[6435]_  = (~\new_[7782]_  | ~\new_[13759]_ ) & (~\new_[7482]_  | ~\new_[14012]_ );
  assign \new_[6436]_  = (~\new_[7783]_  | ~\new_[14105]_ ) & (~\new_[7482]_  | ~\new_[13939]_ );
  assign \new_[6437]_  = (~\new_[7783]_  | ~\new_[13993]_ ) & (~\new_[7482]_  | ~\new_[13731]_ );
  assign \new_[6438]_  = (~\new_[7483]_  | ~\new_[4834]_ ) & (~\new_[7481]_  | ~\new_[13736]_ );
  assign \new_[6439]_  = (~\new_[7783]_  | ~\new_[4619]_ ) & (~\new_[7482]_  | ~\new_[13549]_ );
  assign \new_[6440]_  = (~\new_[7483]_  | ~\new_[4835]_ ) & (~\new_[7481]_  | ~\new_[13648]_ );
  assign \new_[6441]_  = (~\new_[7783]_  | ~\new_[14129]_ ) & (~\new_[7482]_  | ~\new_[14048]_ );
  assign \new_[6442]_  = (~\new_[7781]_  | ~\new_[4839]_ ) & (~\new_[8214]_  | ~\new_[14262]_ );
  assign \new_[6443]_  = (~\new_[7483]_  | ~\new_[4837]_ ) & (~\new_[7481]_  | ~\new_[14023]_ );
  assign \new_[6444]_  = (~\new_[7483]_  | ~\new_[4616]_ ) & (~\new_[7481]_  | ~\new_[13942]_ );
  assign \new_[6445]_  = (~\new_[7781]_  | ~\new_[4840]_ ) & (~\new_[7481]_  | ~\new_[13911]_ );
  assign \new_[6446]_  = (~\new_[7483]_  | ~\new_[4608]_ ) & (~\new_[7481]_  | ~\new_[14025]_ );
  assign \new_[6447]_  = (~\new_[7783]_  | ~\new_[4609]_ ) & (~\new_[7482]_  | ~\new_[13860]_ );
  assign \new_[6448]_  = (~\new_[7783]_  | ~\new_[14029]_ ) & (~\new_[7482]_  | ~\new_[13592]_ );
  assign \new_[6449]_  = (~\new_[7783]_  | ~\new_[4845]_ ) & (~\new_[7482]_  | ~\new_[13727]_ );
  assign \new_[6450]_  = (~\new_[7783]_  | ~\new_[13680]_ ) & (~\new_[7482]_  | ~\new_[13660]_ );
  assign \new_[6451]_  = (~\new_[7783]_  | ~\new_[13676]_ ) & (~\new_[7482]_  | ~\new_[14193]_ );
  assign \new_[6452]_  = (~\new_[7783]_  | ~\new_[14086]_ ) & (~\new_[7482]_  | ~\new_[13834]_ );
  assign \new_[6453]_  = (~\new_[7782]_  | ~\new_[13916]_ ) & (~\new_[7482]_  | ~\new_[13899]_ );
  assign \new_[6454]_  = (~\new_[7782]_  | ~\new_[13847]_ ) & (~\new_[7482]_  | ~\new_[13936]_ );
  assign \new_[6455]_  = (~\new_[8215]_  | ~\new_[4800]_ ) & (~\new_[7481]_  | ~\new_[6253]_ );
  assign \new_[6456]_  = (~\new_[7782]_  | ~\new_[13644]_ ) & (~\new_[7482]_  | ~\new_[13724]_ );
  assign \new_[6457]_  = (~\new_[7782]_  | ~\new_[4852]_ ) & (~\new_[7482]_  | ~\new_[14155]_ );
  assign \new_[6458]_  = (~\new_[7781]_  | ~\new_[4923]_ ) & (~\new_[7482]_  | ~\new_[6247]_ );
  assign \new_[6459]_  = (~\new_[7781]_  | ~\new_[4853]_ ) & (~\new_[7482]_  | ~\new_[13597]_ );
  assign \new_[6460]_  = (~\new_[7782]_  | ~\new_[4787]_ ) & (~\new_[7482]_  | ~\new_[14098]_ );
  assign \new_[6461]_  = \\u4_u2_buf0_orig_reg[29] ;
  assign \new_[6462]_  = ~\new_[7655]_  | ~\new_[8659]_  | ~\new_[12438]_  | ~\new_[7595]_ ;
  assign \new_[6463]_  = ~\new_[6752]_ ;
  assign \new_[6464]_  = u1_u0_token_valid_str1_reg;
  assign \new_[6465]_  = u4_match_r1_reg;
  assign \new_[6466]_  = ~\new_[7671]_  | ~\new_[8660]_  | ~\new_[12445]_  | ~\new_[7596]_ ;
  assign \new_[6467]_  = ~\new_[9248]_  & (~\new_[7322]_  | ~\new_[10475]_ );
  assign \new_[6468]_  = ~\\u4_u0_csr0_reg[0] ;
  assign \new_[6469]_  = ~\new_[14529]_  | ~\new_[2869]_ ;
  assign \new_[6470]_  = \\u1_u0_pid_reg[3] ;
  assign n5405 = ~\new_[7356]_  | ~\new_[7580]_  | ~\new_[7889]_ ;
  assign n5390 = ~\new_[7357]_  | ~\new_[7585]_  | ~\new_[7893]_ ;
  assign n5395 = ~\new_[7358]_  | ~\new_[7588]_  | ~\new_[7897]_ ;
  assign n5400 = ~\new_[7359]_  | ~\new_[7590]_  | ~\new_[7902]_ ;
  assign \new_[6475]_  = ~\\u4_u3_csr0_reg[0] ;
  assign \new_[6476]_  = ~\new_[7858]_  | ~\new_[7549]_  | ~\new_[7558]_ ;
  assign \new_[6477]_  = \new_[2476]_  & \new_[7208]_ ;
  assign \new_[6478]_  = ~\\u4_u1_buf0_orig_reg[31] ;
  assign n5475 = ~n8885 & (~\new_[7553]_  | ~\new_[8960]_ );
  assign \new_[6480]_  = ~\new_[7900]_  | ~\new_[7574]_  | ~\new_[13250]_  | ~\new_[6288]_ ;
  assign \new_[6481]_  = ~\\u4_u0_buf0_orig_reg[13] ;
  assign \new_[6482]_  = ~\new_[7877]_  | ~\new_[7575]_  | ~\new_[13115]_  | ~\new_[6256]_ ;
  assign \new_[6483]_  = ~\\u4_u1_buf0_orig_reg[9] ;
  assign \new_[6484]_  = \\u4_u0_buf0_orig_reg[19] ;
  assign \new_[6485]_  = \\u4_u2_csr1_reg[9] ;
  assign \new_[6486]_  = ~\\u4_u3_csr0_reg[11] ;
  assign \new_[6487]_  = (~\new_[7783]_  | ~\new_[4843]_ ) & (~\new_[7482]_  | ~\new_[13670]_ );
  assign \new_[6488]_  = ~\\u4_u1_buf0_orig_reg[6] ;
  assign \new_[6489]_  = ~\\u4_u1_buf0_orig_reg[8] ;
  assign \new_[6490]_  = ~\\u4_u0_buf0_orig_reg[15] ;
  assign \new_[6491]_  = ~\\u4_u0_buf0_orig_reg[17] ;
  assign \new_[6492]_  = \new_[2047]_  ? \new_[7545]_  : \new_[13665]_ ;
  assign \new_[6493]_  = \new_[5421]_  ? \new_[8609]_  : \new_[13554]_ ;
  assign \new_[6494]_  = \new_[3173]_  ? \new_[8609]_  : \new_[14007]_ ;
  assign \new_[6495]_  = \new_[2178]_  ? \new_[7545]_  : \new_[13618]_ ;
  assign \new_[6496]_  = \new_[3034]_  ? \new_[8609]_  : \new_[13820]_ ;
  assign \new_[6497]_  = \new_[3021]_  ? \new_[8609]_  : \new_[13910]_ ;
  assign \new_[6498]_  = \new_[9037]_  ? \new_[7545]_  : \new_[13972]_ ;
  assign \new_[6499]_  = \new_[2928]_  ? \new_[8609]_  : \new_[13625]_ ;
  assign \new_[6500]_  = \new_[2856]_  ? \new_[7545]_  : \new_[13743]_ ;
  assign \new_[6501]_  = \new_[2638]_  ? \new_[7545]_  : \new_[14177]_ ;
  assign \new_[6502]_  = \new_[2639]_  ? \new_[7545]_  : \new_[14136]_ ;
  assign \new_[6503]_  = \new_[2735]_  ? \new_[7545]_  : \new_[13777]_ ;
  assign \new_[6504]_  = \new_[2177]_  ? \new_[8609]_  : \new_[13551]_ ;
  assign \new_[6505]_  = \new_[2265]_  ? \new_[7545]_  : \new_[14044]_ ;
  assign \new_[6506]_  = \new_[2136]_  ? \new_[7545]_  : \new_[13745]_ ;
  assign \new_[6507]_  = \new_[2075]_  ? \new_[8609]_  : \new_[14144]_ ;
  assign \new_[6508]_  = \new_[2062]_  ? \new_[7545]_  : \new_[13684]_ ;
  assign \new_[6509]_  = \new_[3102]_  ? \new_[7545]_  : \new_[13954]_ ;
  assign \new_[6510]_  = \new_[2047]_  ? \new_[7858]_  : \new_[13498]_ ;
  assign \new_[6511]_  = ~\\u4_u1_buf0_orig_reg[17] ;
  assign \new_[6512]_  = \\u4_u1_buf0_orig_reg[28] ;
  assign \new_[6513]_  = \new_[2547]_  ? \new_[8609]_  : \new_[13776]_ ;
  assign \new_[6514]_  = \new_[2266]_  ? \new_[8609]_  : \new_[14189]_ ;
  assign \new_[6515]_  = \new_[2266]_  ? \new_[7858]_  : \new_[13839]_ ;
  assign \new_[6516]_  = \new_[5421]_  ? \new_[7858]_  : \new_[13619]_ ;
  assign \new_[6517]_  = \new_[9037]_  ? \new_[7858]_  : \new_[14085]_ ;
  assign \new_[6518]_  = \new_[2735]_  ? \new_[7858]_  : \new_[14206]_ ;
  assign \new_[6519]_  = \new_[2177]_  ? \new_[7858]_  : \new_[13536]_ ;
  assign \new_[6520]_  = \new_[2048]_  ? \new_[7545]_  : \new_[13898]_ ;
  assign \new_[6521]_  = ~u1_u2_wr_done_reg;
  assign \new_[6522]_  = ~u1_u2_idma_done_reg;
  assign \new_[6523]_  = ~\new_[11146]_  & ~\new_[6895]_ ;
  assign \new_[6524]_  = \\u4_u0_csr1_reg[10] ;
  assign \new_[6525]_  = \new_[2034]_  ? \new_[8609]_  : \new_[13537]_ ;
  assign \new_[6526]_  = \\u4_u2_csr1_reg[4] ;
  assign \new_[6527]_  = (~\new_[8215]_  | ~\new_[4838]_ ) & (~\new_[7481]_  | ~\new_[13826]_ );
  assign \new_[6528]_  = ~\\u4_u0_buf0_orig_reg[0] ;
  assign \new_[6529]_  = (~\new_[8215]_  | ~\new_[12883]_ ) & (~\new_[7481]_  | ~\new_[6258]_ );
  assign n5375 = ~\new_[6903]_  | (~\new_[9786]_  & ~\new_[10681]_ );
  assign \new_[6531]_  = ~\new_[4856]_  | ~\new_[6861]_ ;
  assign \new_[6532]_  = \new_[7299]_  | \new_[14216]_ ;
  assign n5415 = ~\new_[7934]_  | ~\new_[7146]_  | ~\new_[7398]_ ;
  assign \new_[6534]_  = ~\new_[4854]_  | ~\new_[7313]_ ;
  assign \new_[6535]_  = ~\new_[7313]_  | ~\new_[4855]_ ;
  assign \new_[6536]_  = ~\new_[6861]_  | ~\new_[4886]_ ;
  assign n5425 = ~\new_[6842]_ ;
  assign \new_[6538]_  = \\u4_u2_csr1_reg[2] ;
  assign \new_[6539]_  = \\u4_u0_csr1_reg[11] ;
  assign \new_[6540]_  = ~\new_[14267]_  | ~\new_[7309]_ ;
  assign \new_[6541]_  = ~\new_[13503]_  | ~\new_[7309]_ ;
  assign \new_[6542]_  = ~\new_[7321]_  | ~\new_[9644]_  | ~\new_[8581]_ ;
  assign \new_[6543]_  = \\u4_u0_csr1_reg[12] ;
  assign \new_[6544]_  = \\u4_u2_csr0_reg[5] ;
  assign \new_[6545]_  = \\u4_u2_csr1_reg[12] ;
  assign \new_[6546]_  = \new_[12467]_  | \new_[7299]_ ;
  assign \new_[6547]_  = \\u4_u0_csr1_reg[4] ;
  assign \new_[6548]_  = \\u4_u2_csr1_reg[10] ;
  assign \new_[6549]_  = \\u4_u0_csr1_reg[6] ;
  assign \new_[6550]_  = ~\\u4_u3_buf0_orig_reg[3] ;
  assign \new_[6551]_  = \\u4_u1_buf0_orig_reg[24] ;
  assign \new_[6552]_  = \\u4_u2_csr0_reg[8] ;
  assign n5380 = ~\new_[6898]_  | ~\new_[8205]_ ;
  assign n5410 = ~\new_[7397]_  | ~\new_[6864]_  | ~\new_[9193]_ ;
  assign \new_[6555]_  = ~\new_[6847]_ ;
  assign \new_[6556]_  = \\u4_u2_buf0_orig_reg[30] ;
  assign \new_[6557]_  = \\u4_u0_csr0_reg[9] ;
  assign \new_[6558]_  = ~\new_[7847]_  | ~\new_[7606]_  | ~\new_[13232]_  | ~\new_[6276]_ ;
  assign \new_[6559]_  = ~\\u4_u0_csr0_reg[11] ;
  assign \new_[6560]_  = \\u4_u3_buf0_orig_reg[29] ;
  assign \new_[6561]_  = \\u4_u0_csr0_reg[8] ;
  assign \new_[6562]_  = \\u4_u2_csr0_reg[1] ;
  assign \new_[6563]_  = \\u4_u0_csr0_reg[5] ;
  assign \new_[6564]_  = ~\\u4_u2_csr0_reg[11] ;
  assign \new_[6565]_  = ~\new_[13363]_  | ~\new_[6899]_  | ~\new_[7366]_ ;
  assign \new_[6566]_  = ~\new_[3882]_  | ~\new_[6883]_  | ~\new_[9420]_ ;
  assign \new_[6567]_  = \\u4_u0_csr0_reg[7] ;
  assign n5485 = \new_[13601]_  ? \new_[7869]_  : \new_[13723]_ ;
  assign n5560 = \new_[14019]_  ? \new_[7869]_  : \new_[13547]_ ;
  assign n5565 = \new_[13654]_  ? \new_[7869]_  : \new_[13530]_ ;
  assign n5500 = \new_[13921]_  ? \new_[7869]_  : \new_[13531]_ ;
  assign n5505 = \new_[13502]_  ? \new_[7869]_  : \new_[13759]_ ;
  assign n5510 = \new_[13594]_  ? \new_[7869]_  : \new_[14105]_ ;
  assign n5520 = \new_[14247]_  ? \new_[7869]_  : \new_[13993]_ ;
  assign \new_[6575]_  = (~\new_[7782]_  | ~\new_[13547]_ ) & (~\new_[7482]_  | ~\new_[14241]_ );
  assign n5490 = \new_[13508]_  ? \new_[7869]_  : \new_[14129]_ ;
  assign n5495 = \new_[13801]_  ? \new_[7869]_  : \new_[14029]_ ;
  assign n5525 = \new_[13785]_  ? \new_[7869]_  : \new_[13676]_ ;
  assign n5530 = \new_[13523]_  ? \new_[7869]_  : \new_[14086]_ ;
  assign n5535 = \new_[14051]_  ? \new_[7869]_  : \new_[13916]_ ;
  assign n5540 = \new_[13526]_  ? \new_[7869]_  : \new_[13576]_ ;
  assign n5545 = \new_[13990]_  ? \new_[7869]_  : \new_[13847]_ ;
  assign n5550 = \new_[13505]_  ? \new_[7869]_  : \new_[14053]_ ;
  assign n5555 = \new_[13628]_  ? \new_[7869]_  : \new_[13644]_ ;
  assign n5515 = \new_[13999]_  ? \new_[7869]_  : \new_[14124]_ ;
  assign \new_[6586]_  = ~\new_[13289]_  | ~\new_[6900]_  | ~\new_[7369]_ ;
  assign \new_[6587]_  = \new_[4289]_  ? \new_[7455]_  : \new_[7684]_ ;
  assign \new_[6588]_  = \\u4_u3_buf0_orig_reg[25] ;
  assign \new_[6589]_  = ~\new_[3476]_  | ~\new_[6884]_  | ~\new_[9417]_ ;
  assign \new_[6590]_  = \new_[4288]_  ? \new_[7455]_  : \new_[7911]_ ;
  assign \new_[6591]_  = \new_[4069]_  ? \new_[7455]_  : \new_[7402]_ ;
  assign \new_[6592]_  = \\u4_u1_buf0_orig_reg[20] ;
  assign \new_[6593]_  = \\u4_u0_csr0_reg[3] ;
  assign \new_[6594]_  = ~\new_[6858]_ ;
  assign n5480 = ~\new_[8261]_  & ~\new_[9842]_ ;
  assign \new_[6596]_  = (~\new_[7483]_  | ~\new_[4796]_ ) & (~\new_[8214]_  | ~\new_[6250]_ );
  assign \new_[6597]_  = ~\\u4_u2_buf0_orig_reg[6] ;
  assign \new_[6598]_  = ~\\u4_u2_buf0_orig_reg[8] ;
  assign \new_[6599]_  = \\u4_u0_csr0_reg[1] ;
  assign \new_[6600]_  = ~\\u4_u2_buf0_orig_reg[5] ;
  assign \new_[6601]_  = ~\\u4_u2_buf0_orig_reg[3] ;
  assign \new_[6602]_  = \\u4_u3_buf0_orig_reg[20] ;
  assign \new_[6603]_  = ~\\u4_u3_buf0_orig_reg[18] ;
  assign \new_[6604]_  = \\u1_u0_token1_reg[6] ;
  assign \new_[6605]_  = \\u4_dout_reg[4] ;
  assign \new_[6606]_  = ~\new_[6874]_ ;
  assign \new_[6607]_  = ~\\u4_inta_msk_reg[8] ;
  assign \new_[6608]_  = ~\\u4_intb_msk_reg[3] ;
  assign \new_[6609]_  = \\u4_inta_msk_reg[2] ;
  assign \new_[6610]_  = \\u4_inta_msk_reg[4] ;
  assign \new_[6611]_  = \\u4_inta_msk_reg[0] ;
  assign \new_[6612]_  = ~\new_[7936]_  | ~\new_[12628]_  | ~\new_[7689]_ ;
  assign \new_[6613]_  = ~\new_[7935]_  | ~\new_[13286]_  | ~\new_[7691]_ ;
  assign \new_[6614]_  = ~\new_[13355]_  | ~\new_[7379]_  | ~\new_[7692]_ ;
  assign \new_[6615]_  = ~\new_[5562]_  & (~\new_[7712]_  | ~\new_[8633]_ );
  assign \new_[6616]_  = ~\new_[5489]_  & (~\new_[7712]_  | ~\new_[8970]_ );
  assign \new_[6617]_  = ~\new_[7757]_  & (~\new_[7688]_  | ~\new_[3693]_ );
  assign \new_[6618]_  = ~\new_[7758]_  & (~\new_[7690]_  | ~\new_[3316]_ );
  assign \new_[6619]_  = ~\new_[9850]_  | ~\new_[7396]_  | ~\new_[8610]_ ;
  assign \new_[6620]_  = ~\new_[5490]_  & (~\new_[7712]_  | ~\new_[7866]_ );
  assign \new_[6621]_  = ~\new_[6895]_ ;
  assign \new_[6622]_  = ~\new_[5491]_  & (~\new_[7712]_  | ~\new_[8247]_ );
  assign \new_[6623]_  = ~\new_[7368]_  & (~\new_[7750]_  | ~\new_[10945]_ );
  assign \new_[6624]_  = (~\new_[7653]_  | ~\new_[3686]_ ) & (~\new_[8323]_  | ~\new_[3464]_ );
  assign \new_[6625]_  = (~\new_[7777]_  & ~\new_[9276]_ ) | (~\new_[9808]_  & ~\new_[8977]_ );
  assign \new_[6626]_  = ~\new_[7388]_  | (~\new_[7878]_  & ~\new_[3464]_ );
  assign \new_[6627]_  = ~\new_[7394]_  | (~\new_[7870]_  & ~\new_[3787]_ );
  assign \new_[6628]_  = \new_[2076]_  ? \new_[8233]_  : \new_[13560]_ ;
  assign \new_[6629]_  = ~\new_[7465]_  & (~\new_[14270]_  | ~\new_[2869]_ );
  assign \new_[6630]_  = ~\new_[7317]_  & ~\new_[14225]_ ;
  assign \new_[6631]_  = ~\new_[14507]_  | ~\new_[2505]_ ;
  assign \new_[6632]_  = ~\new_[7317]_  & ~\new_[14071]_ ;
  assign \new_[6633]_  = ~\new_[6904]_ ;
  assign \new_[6634]_  = ~\new_[7317]_  & ~\new_[14215]_ ;
  assign \new_[6635]_  = ~\\u4_u3_buf0_orig_reg[1] ;
  assign \new_[6636]_  = \\u4_dout_reg[20] ;
  assign \new_[6637]_  = \\u4_dout_reg[16] ;
  assign \new_[6638]_  = \\u4_dout_reg[17] ;
  assign \new_[6639]_  = \\u4_dout_reg[18] ;
  assign \new_[6640]_  = \\u4_dout_reg[19] ;
  assign \new_[6641]_  = \\u4_dout_reg[21] ;
  assign \new_[6642]_  = \\u4_dout_reg[24] ;
  assign \new_[6643]_  = \\u4_dout_reg[25] ;
  assign \new_[6644]_  = \\u4_dout_reg[26] ;
  assign \new_[6645]_  = \\u4_dout_reg[28] ;
  assign \new_[6646]_  = \\u4_dout_reg[5] ;
  assign \new_[6647]_  = \\u4_dout_reg[6] ;
  assign \new_[6648]_  = ~\new_[6912]_ ;
  assign \new_[6649]_  = ~\new_[7408]_  | ~\new_[12528]_ ;
  assign n5675 = ~\new_[7714]_  & ~\new_[7411]_ ;
  assign \new_[6651]_  = ~\new_[7465]_  & (~\new_[14270]_  | ~\new_[13092]_ );
  assign \new_[6652]_  = ~\new_[7550]_  & (~\new_[7866]_  | ~\new_[5766]_ );
  assign \new_[6653]_  = ~\\u4_u3_buf0_orig_reg[17] ;
  assign \new_[6654]_  = ~\new_[7317]_  & ~\new_[11733]_ ;
  assign n5610 = ~\new_[12849]_  & (~\new_[7726]_  | ~\new_[8087]_ );
  assign n5615 = ~\new_[12849]_  & (~\new_[7727]_  | ~\new_[8089]_ );
  assign n5620 = ~\new_[12505]_  & (~\new_[7728]_  | ~\new_[8099]_ );
  assign n5625 = ~\new_[12505]_  & (~\new_[7729]_  | ~\new_[8100]_ );
  assign n5630 = ~\new_[12505]_  & (~\new_[7730]_  | ~\new_[8101]_ );
  assign \new_[6660]_  = ~\new_[7413]_  | ~\new_[13470]_ ;
  assign \new_[6661]_  = ~\\u4_u3_dma_out_left_reg[8] ;
  assign \new_[6662]_  = ~\\u4_u0_dma_out_left_reg[8] ;
  assign \new_[6663]_  = ~\new_[7317]_  & ~\new_[14100]_ ;
  assign n5680 = ~\new_[8512]_  | ~phy_rst_pad_o | ~\new_[7733]_ ;
  assign n5590 = ~\new_[12804]_  & (~\new_[7719]_  | ~\new_[12092]_ );
  assign \new_[6666]_  = ~\\u4_u1_dma_out_left_reg[8] ;
  assign n5635 = ~\new_[12849]_  & (~\new_[7756]_  | ~\new_[8076]_ );
  assign n5640 = ~\new_[12505]_  & (~\new_[7759]_  | ~\new_[8074]_ );
  assign n5645 = ~\new_[12245]_  & (~\new_[7760]_  | ~\new_[8039]_ );
  assign n5650 = ~\new_[12505]_  & (~\new_[7761]_  | ~\new_[8148]_ );
  assign \new_[6671]_  = ~\\u4_u2_dma_out_left_reg[8] ;
  assign \new_[6672]_  = ~\new_[7317]_  & ~\new_[11577]_ ;
  assign \new_[6673]_  = ~\new_[7492]_  & (~\new_[7775]_  | ~\new_[9395]_ );
  assign \new_[6674]_  = ~\new_[9640]_  | ~\new_[7426]_ ;
  assign n5685 = ~\new_[7420]_  & ~\new_[7418]_ ;
  assign n5655 = ~\new_[12849]_  & (~\new_[7732]_  | ~\new_[8121]_ );
  assign n5660 = ~\new_[12849]_  & (~\new_[7738]_  | ~\new_[8079]_ );
  assign n5665 = ~\new_[12505]_  & (~\new_[7725]_  | ~\new_[8190]_ );
  assign n5670 = ~\new_[12849]_  & (~\new_[7739]_  | ~\new_[8014]_ );
  assign \new_[6680]_  = ~\new_[7434]_  & ~\new_[6254]_ ;
  assign \new_[6681]_  = ~\new_[7433]_  & ~\new_[6561]_ ;
  assign n5605 = ~\new_[7416]_  & ~n8885;
  assign \new_[6683]_  = ~\new_[7423]_  & (~\new_[8578]_  | ~\new_[9232]_ );
  assign \new_[6684]_  = ~\new_[7419]_  & (~\new_[11676]_  | ~\new_[8625]_ );
  assign n5740 = ~\new_[7411]_  & (~\new_[7852]_  | ~\new_[13753]_ );
  assign n5690 = ~n7075 & (~\new_[7766]_  | ~\new_[13803]_ );
  assign \new_[6687]_  = ~\new_[7412]_  & (~\new_[14451]_  | ~\new_[12975]_ );
  assign \new_[6688]_  = ~\new_[7454]_  | (~\new_[14421]_  & ~\new_[2873]_ );
  assign \new_[6689]_  = ~\new_[7435]_  & ~\new_[6552]_ ;
  assign \new_[6690]_  = \\u4_u1_csr0_reg[3] ;
  assign \new_[6691]_  = ~\\u4_u3_buf0_orig_reg[11] ;
  assign \new_[6692]_  = ~\new_[7939]_  | (~\new_[8125]_  & ~\new_[7752]_ );
  assign \new_[6693]_  = ~\\u4_u3_buf0_orig_reg[13] ;
  assign \new_[6694]_  = ~\new_[7939]_  | (~\new_[8128]_  & ~\new_[7753]_ );
  assign \new_[6695]_  = ~\new_[7292]_ ;
  assign \new_[6696]_  = \\u1_u0_token1_reg[0] ;
  assign \new_[6697]_  = \\u4_u3_int_stat_reg[6] ;
  assign \new_[6698]_  = \new_[13732]_  ^ \new_[7765]_ ;
  assign \new_[6699]_  = \new_[14640]_  ^ \new_[14635]_ ;
  assign \new_[6700]_  = ~suspend_clr_wr_reg;
  assign \new_[6701]_  = ~\\u4_u3_buf0_orig_reg[10] ;
  assign \new_[6702]_  = ~\new_[7448]_  | ~\new_[13953]_ ;
  assign \new_[6703]_  = \new_[14341]_  & \new_[14634]_ ;
  assign \new_[6704]_  = ~\new_[14341]_  & ~\new_[14634]_ ;
  assign \new_[6705]_  = ~\new_[7745]_  | ~\new_[7445]_ ;
  assign \new_[6706]_  = ~\new_[7745]_  | ~\new_[7443]_ ;
  assign \new_[6707]_  = \new_[7448]_  & \new_[7449]_ ;
  assign \new_[6708]_  = ~\new_[7446]_  & ~\new_[7444]_ ;
  assign n5580 = ~\new_[7787]_  | ~\new_[8217]_  | ~\new_[9503]_ ;
  assign \new_[6710]_  = (~\new_[7776]_  & ~\new_[11698]_ ) | (~\new_[11377]_  & ~\new_[9817]_ );
  assign n5750 = ~n8885 & (~\new_[7788]_  | ~\new_[9781]_ );
  assign n5600 = ~\new_[7883]_  | ~\new_[13022]_  | ~\new_[12627]_  | ~\new_[12631]_ ;
  assign n5595 = ~n8885 & (~\new_[8239]_  | ~\new_[7779]_ );
  assign n5725 = ~n8885 & (~\new_[8624]_  | ~\new_[7785]_ );
  assign n5575 = ~\new_[7884]_  | ~\new_[12507]_  | ~\new_[12829]_  | ~\new_[12634]_ ;
  assign \new_[6716]_  = \\u1_u0_token1_reg[1] ;
  assign \new_[6717]_  = ~\new_[14344]_  | ~\new_[9781]_  | ~\new_[7432]_  | ~\new_[14345]_ ;
  assign \new_[6718]_  = \\u1_u0_token1_reg[2] ;
  assign \new_[6719]_  = ~\new_[7468]_  & (~\new_[9187]_  | ~\new_[9229]_ );
  assign n5730 = ~n8885 & (~\new_[7559]_  | ~\new_[8596]_ );
  assign \new_[6721]_  = \\u4_inta_msk_reg[1] ;
  assign \new_[6722]_  = \\u4_inta_msk_reg[3] ;
  assign \new_[6723]_  = \\u4_inta_msk_reg[5] ;
  assign \new_[6724]_  = \\u4_inta_msk_reg[6] ;
  assign \new_[6725]_  = ~\\u4_inta_msk_reg[7] ;
  assign \new_[6726]_  = ~\\u4_intb_msk_reg[0] ;
  assign \new_[6727]_  = ~\\u4_intb_msk_reg[1] ;
  assign \new_[6728]_  = ~\\u4_intb_msk_reg[2] ;
  assign \new_[6729]_  = ~\\u4_intb_msk_reg[4] ;
  assign \new_[6730]_  = ~\\u4_intb_msk_reg[5] ;
  assign \new_[6731]_  = ~\\u4_intb_msk_reg[6] ;
  assign \new_[6732]_  = ~\\u4_intb_msk_reg[8] ;
  assign \new_[6733]_  = \\u4_u3_buf0_orig_reg[19] ;
  assign \new_[6734]_  = ~\\u4_u3_buf0_orig_reg[4] ;
  assign \new_[6735]_  = ~\\u4_u3_buf0_orig_reg[7] ;
  assign \new_[6736]_  = \\u1_u0_token1_reg[3] ;
  assign \new_[6737]_  = \\u1_u0_token1_reg[4] ;
  assign \new_[6738]_  = \\u1_u0_token1_reg[5] ;
  assign \new_[6739]_  = \\u1_u0_token1_reg[7] ;
  assign \new_[6740]_  = ~\new_[7317]_  & ~\new_[14191]_ ;
  assign \new_[6741]_  = ~\new_[7317]_  & ~\new_[13708]_ ;
  assign \new_[6742]_  = ~\new_[7317]_  & ~\new_[13992]_ ;
  assign \new_[6743]_  = \\u4_u3_csr0_reg[3] ;
  assign n5695 = \new_[13166]_  ? \new_[7773]_  : \new_[6015]_ ;
  assign n5700 = \new_[12846]_  ? \new_[7773]_  : \new_[6016]_ ;
  assign n5745 = \new_[12783]_  ? \new_[7773]_  : \new_[6033]_ ;
  assign n5705 = \new_[12870]_  ? \new_[7773]_  : \new_[6017]_ ;
  assign n5710 = \new_[12651]_  ? \new_[7773]_  : \new_[6018]_ ;
  assign n5715 = \new_[12816]_  ? \new_[7773]_  : \new_[6019]_ ;
  assign n5585 = \new_[12916]_  ? \new_[7773]_  : \new_[5978]_ ;
  assign n5720 = \new_[13192]_  ? \new_[7773]_  : \new_[12396]_ ;
  assign \new_[6752]_  = (~\new_[8620]_  & ~\new_[11698]_  & ~\new_[10811]_ ) | (~\new_[11698]_  & ~\new_[7865]_  & ~\new_[9276]_ );
  assign \new_[6753]_  = ~\new_[7452]_  | (~\new_[8202]_  & ~\new_[4607]_ );
  assign \new_[6754]_  = ~\\u4_intb_msk_reg[7] ;
  assign \new_[6755]_  = ~\new_[9265]_  & (~\new_[7581]_  | ~\new_[10475]_ );
  assign \new_[6756]_  = ~\new_[9296]_  & (~\new_[7583]_  | ~\new_[10475]_ );
  assign \new_[6757]_  = ~\new_[9254]_  & (~\new_[7584]_  | ~\new_[10475]_ );
  assign \new_[6758]_  = ~\new_[7906]_  | ~\new_[7933]_  | ~\new_[9122]_  | ~\new_[8312]_ ;
  assign \new_[6759]_  = ~\new_[7178]_ ;
  assign \new_[6760]_  = ~\new_[7317]_  & ~\new_[13927]_ ;
  assign \new_[6761]_  = ~\new_[14792]_  & ~\new_[13837]_ ;
  assign \new_[6762]_  = ~\new_[7181]_ ;
  assign \new_[6763]_  = ~\new_[14792]_  | ~\new_[13837]_ ;
  assign \new_[6764]_  = (~\new_[12483]_  & ~\new_[9367]_ ) | (~\new_[7593]_  & ~\new_[6253]_ );
  assign \new_[6765]_  = (~\new_[7594]_  & ~\new_[6266]_ ) | (~\new_[12446]_  & ~\new_[9368]_ );
  assign \new_[6766]_  = \new_[7540]_  | \new_[2872]_ ;
  assign \new_[6767]_  = (~\new_[12438]_  & ~\new_[9369]_ ) | (~\new_[7595]_  & ~\new_[6200]_ );
  assign \new_[6768]_  = \new_[14792]_  | \new_[2872]_ ;
  assign \new_[6769]_  = \new_[7540]_  | \new_[2871]_ ;
  assign \new_[6770]_  = ~\new_[7189]_ ;
  assign \new_[6771]_  = (~\new_[12445]_  & ~\new_[9370]_ ) | (~\new_[7596]_  & ~\new_[6009]_ );
  assign \new_[6772]_  = ~\new_[7191]_ ;
  assign \new_[6773]_  = ~\new_[7192]_ ;
  assign \new_[6774]_  = ~\new_[7540]_  & ~\new_[13917]_ ;
  assign \new_[6775]_  = ~\new_[7195]_ ;
  assign \new_[6776]_  = ~\new_[7196]_ ;
  assign \new_[6777]_  = ~\new_[7197]_ ;
  assign \new_[6778]_  = ~\new_[8233]_  | ~\new_[7857]_  | ~\new_[7864]_ ;
  assign \new_[6779]_  = ~\new_[7289]_ ;
  assign \new_[6780]_  = ~\\u4_u0_dma_out_left_reg[11] ;
  assign \new_[6781]_  = ~\\u4_u1_dma_out_left_reg[11] ;
  assign \new_[6782]_  = \new_[2177]_  ? \new_[8233]_  : \new_[14010]_ ;
  assign \new_[6783]_  = \new_[2639]_  ? \new_[8233]_  : \new_[13714]_ ;
  assign \new_[6784]_  = \new_[2928]_  ? \new_[8233]_  : \new_[13640]_ ;
  assign \new_[6785]_  = \new_[3021]_  ? \new_[8233]_  : \new_[13662]_ ;
  assign \new_[6786]_  = \new_[2547]_  ? \new_[8233]_  : \new_[13833]_ ;
  assign \new_[6787]_  = \new_[2062]_  ? \new_[8233]_  : \new_[13782]_ ;
  assign \new_[6788]_  = ~\new_[8236]_  | ~\new_[6288]_ ;
  assign \new_[6789]_  = ~\new_[8236]_  | ~\new_[13867]_ ;
  assign \new_[6790]_  = ~\new_[8236]_  | ~\new_[13697]_ ;
  assign \new_[6791]_  = ~\new_[8236]_  | ~\new_[6562]_ ;
  assign \new_[6792]_  = ~\new_[8236]_  | ~\new_[6289]_ ;
  assign \new_[6793]_  = ~\new_[8236]_  | ~\new_[6545]_ ;
  assign \new_[6794]_  = ~\new_[8236]_  | ~\new_[6008]_ ;
  assign \new_[6795]_  = ~\new_[8236]_  | ~\new_[6809]_ ;
  assign \new_[6796]_  = ~\new_[8236]_  | ~\new_[6010]_ ;
  assign \new_[6797]_  = ~\new_[8236]_  | ~\new_[6287]_ ;
  assign \new_[6798]_  = ~\new_[8236]_  | ~\new_[13499]_ ;
  assign \new_[6799]_  = ~\new_[8236]_  | ~\new_[6544]_ ;
  assign \new_[6800]_  = ~\new_[8236]_  | ~\new_[13719]_ ;
  assign \new_[6801]_  = ~\new_[8236]_  | ~\new_[14056]_ ;
  assign \new_[6802]_  = ~\new_[8236]_  | ~\new_[14021]_ ;
  assign \new_[6803]_  = ~\new_[8236]_  | ~\new_[13774]_ ;
  assign \new_[6804]_  = ~\new_[8236]_  | ~\new_[13605]_ ;
  assign \new_[6805]_  = ~\new_[8236]_  | ~\new_[6552]_ ;
  assign \new_[6806]_  = ~\new_[8236]_  | ~\new_[6548]_ ;
  assign \new_[6807]_  = ~\new_[8236]_  | ~\new_[5502]_ ;
  assign \new_[6808]_  = ~\new_[8236]_  | ~\new_[13612]_ ;
  assign \new_[6809]_  = \\u4_u2_csr0_reg[3] ;
  assign \new_[6810]_  = ~\new_[8236]_  | ~\new_[6286]_ ;
  assign \new_[6811]_  = ~\new_[8236]_  | ~\new_[14055]_ ;
  assign \new_[6812]_  = ~\new_[8236]_  | ~\new_[6009]_ ;
  assign \new_[6813]_  = ~\new_[8236]_  | ~\new_[14233]_ ;
  assign \new_[6814]_  = ~\new_[8236]_  | ~\new_[13640]_ ;
  assign \new_[6815]_  = ~\new_[8236]_  | ~\new_[13822]_ ;
  assign \new_[6816]_  = ~\new_[8236]_  | ~\new_[13714]_ ;
  assign \new_[6817]_  = ~\new_[8236]_  | ~\new_[13662]_ ;
  assign \new_[6818]_  = ~\new_[8236]_  | ~\new_[13729]_ ;
  assign \new_[6819]_  = ~\new_[8236]_  | ~\new_[13504]_ ;
  assign \new_[6820]_  = ~\new_[8236]_  | ~\new_[13791]_ ;
  assign \new_[6821]_  = ~\new_[8236]_  | ~\new_[13888]_ ;
  assign \new_[6822]_  = ~\new_[8236]_  | ~\new_[13795]_ ;
  assign \new_[6823]_  = ~\new_[8236]_  | ~\new_[13639]_ ;
  assign \new_[6824]_  = ~\new_[8236]_  | ~\new_[13864]_ ;
  assign \new_[6825]_  = ~\new_[8236]_  | ~\new_[13516]_ ;
  assign \new_[6826]_  = ~\new_[8236]_  | ~\new_[13716]_ ;
  assign \new_[6827]_  = ~\new_[8236]_  | ~\new_[13511]_ ;
  assign \new_[6828]_  = ~\new_[8236]_  | ~\new_[13800]_ ;
  assign \new_[6829]_  = ~\new_[8236]_  | ~\new_[13848]_ ;
  assign \new_[6830]_  = ~\new_[8236]_  | ~\new_[6284]_ ;
  assign \new_[6831]_  = ~\new_[7542]_  | ~\new_[8648]_ ;
  assign \new_[6832]_  = ~\new_[7542]_  | ~\new_[8650]_ ;
  assign \new_[6833]_  = ~\new_[7322]_  | ~\new_[10849]_ ;
  assign \new_[6834]_  = ~\new_[14227]_  | ~\new_[7545]_ ;
  assign \new_[6835]_  = ~\new_[7314]_  | ~\new_[2136]_ ;
  assign \new_[6836]_  = ~\new_[7555]_  | ~\new_[5185]_ ;
  assign \new_[6837]_  = ~\new_[14134]_  | ~\new_[7545]_ ;
  assign \new_[6838]_  = ~\\u4_u3_buf0_orig_reg[6] ;
  assign \new_[6839]_  = ~\new_[7554]_  | ~\new_[2266]_ ;
  assign \new_[6840]_  = ~\new_[7554]_  | ~\new_[2178]_ ;
  assign \new_[6841]_  = ~\new_[7314]_  | ~\new_[2177]_ ;
  assign \new_[6842]_  = ~\OpMode_pad_o[0]  | ~\new_[8205]_  | ~\new_[7678]_ ;
  assign \new_[6843]_  = ~\new_[5148]_  | ~\new_[7315]_ ;
  assign \new_[6844]_  = ~\new_[7315]_  | ~\new_[5174]_ ;
  assign \new_[6845]_  = ~\new_[5149]_  | ~\new_[7555]_ ;
  assign \new_[6846]_  = ~\\u4_u3_buf0_orig_reg[2] ;
  assign \new_[6847]_  = ~\new_[7284]_ ;
  assign \new_[6848]_  = \new_[2114]_  ? \new_[8233]_  : \new_[13986]_ ;
  assign \new_[6849]_  = ~\new_[7317]_  & ~\new_[13642]_ ;
  assign \new_[6850]_  = u0_u0_idle_long_reg;
  assign \new_[6851]_  = ~\new_[13326]_  | ~\new_[7350]_  | ~\new_[7603]_ ;
  assign \new_[6852]_  = ~\new_[4288]_  | ~\new_[7321]_  | ~\new_[9651]_ ;
  assign \new_[6853]_  = \\u4_u3_buf0_orig_reg[27] ;
  assign \new_[6854]_  = \new_[3938]_  ^ \new_[7674]_ ;
  assign \new_[6855]_  = \new_[3466]_  ^ \new_[7675]_ ;
  assign \new_[6856]_  = \new_[3686]_  ^ \new_[7676]_ ;
  assign \new_[6857]_  = \new_[3879]_  ^ \new_[7677]_ ;
  assign \new_[6858]_  = ~\new_[7548]_ ;
  assign n5735 = ~\new_[7869]_  & ~\new_[9842]_ ;
  assign \new_[6860]_  = ~\new_[7311]_ ;
  assign \new_[6861]_  = ~\new_[7314]_ ;
  assign \new_[6862]_  = ~\\u4_u3_ienb_reg[5] ;
  assign \new_[6863]_  = ~\\u4_u3_iena_reg[3] ;
  assign \new_[6864]_  = ~\new_[9517]_  | ~\new_[7573]_ ;
  assign \new_[6865]_  = ~\\u4_u1_iena_reg[4] ;
  assign \new_[6866]_  = ~\\u4_u3_ienb_reg[2] ;
  assign \new_[6867]_  = ~\\u4_u3_ienb_reg[4] ;
  assign \new_[6868]_  = ~\\u4_u1_iena_reg[5] ;
  assign \new_[6869]_  = ~\\u4_u3_iena_reg[4] ;
  assign \new_[6870]_  = ~\\u4_u3_ienb_reg[3] ;
  assign \new_[6871]_  = ~\\u4_u3_ienb_reg[1] ;
  assign \new_[6872]_  = ~\\u4_u3_iena_reg[5] ;
  assign \new_[6873]_  = ~\\u4_u3_ienb_reg[0] ;
  assign \new_[6874]_  = \\u1_u3_new_size_reg[0] ;
  assign \new_[6875]_  = ~\\u4_u1_iena_reg[0] ;
  assign \new_[6876]_  = ~\\u4_u0_csr1_reg[7] ;
  assign \new_[6877]_  = ~\new_[10105]_  | ~\new_[8333]_  | ~\new_[10842]_  | ~\new_[13194]_ ;
  assign \new_[6878]_  = ~\\u4_u3_csr1_reg[7] ;
  assign \new_[6879]_  = ~\new_[9600]_  | ~\new_[8413]_  | ~\new_[10834]_  | ~\new_[13001]_ ;
  assign \new_[6880]_  = ~\\u4_u1_iena_reg[1] ;
  assign \new_[6881]_  = ~\\u4_u3_iena_reg[1] ;
  assign \new_[6882]_  = ~\\u4_u1_iena_reg[3] ;
  assign \new_[6883]_  = ~\new_[13461]_  | ~\new_[7619]_  | ~\new_[7908]_ ;
  assign \new_[6884]_  = ~\new_[13324]_  | ~\new_[7620]_  | ~\new_[7910]_ ;
  assign n5950 = ~\new_[7586]_  & ~\new_[12842]_ ;
  assign n5955 = ~\new_[12849]_  & (~\new_[8041]_  | ~\new_[9359]_ );
  assign n5970 = ~\new_[7698]_  & ~\new_[12245]_ ;
  assign n5975 = ~\new_[7699]_  & ~\new_[12245]_ ;
  assign n5980 = ~\new_[7700]_  & ~\new_[12245]_ ;
  assign n5845 = ~\new_[7701]_  & ~\new_[12245]_ ;
  assign n5985 = ~\new_[7702]_  & ~\new_[12245]_ ;
  assign n5840 = ~\new_[7703]_  & ~\new_[12245]_ ;
  assign n5990 = ~\new_[7704]_  & ~\new_[12245]_ ;
  assign \new_[6894]_  = ~\new_[8440]_  & (~\new_[7909]_  | ~\new_[4073]_ );
  assign \new_[6895]_  = \new_[7654]_  & \new_[3880]_ ;
  assign \new_[6896]_  = ~\new_[7604]_  | ~\new_[14139]_ ;
  assign \new_[6897]_  = ~\new_[7604]_  | ~\new_[13364]_ ;
  assign \new_[6898]_  = ~\new_[7678]_  | ~\OpMode_pad_o[1] ;
  assign \new_[6899]_  = (~\new_[8292]_  | ~\new_[3879]_ ) & (~\new_[7948]_  | ~\new_[3787]_ );
  assign \new_[6900]_  = (~\new_[7899]_  | ~\new_[3466]_ ) & (~\new_[7944]_  | ~\new_[3310]_ );
  assign \new_[6901]_  = ~\new_[7621]_  | (~\new_[8262]_  & ~\new_[3940]_ );
  assign \new_[6902]_  = ~\new_[7638]_  | (~\new_[8284]_  & ~\new_[3310]_ );
  assign \new_[6903]_  = ~\new_[7636]_  & (~\new_[10484]_  | ~\new_[13298]_ );
  assign \new_[6904]_  = ~\new_[14507]_  & ~\new_[2505]_ ;
  assign \new_[6905]_  = ~\new_[7653]_  | ~\new_[3464]_ ;
  assign \new_[6906]_  = ~\new_[7366]_ ;
  assign \new_[6907]_  = \\u4_dout_reg[29] ;
  assign \new_[6908]_  = \\u4_dout_reg[30] ;
  assign \new_[6909]_  = \\u4_dout_reg[31] ;
  assign \new_[6910]_  = \\u4_dout_reg[27] ;
  assign \new_[6911]_  = ~\new_[7369]_ ;
  assign \new_[6912]_  = ~\new_[7653]_  | ~\new_[8323]_ ;
  assign n6000 = ~\new_[12849]_  & (~\new_[8120]_  | ~\new_[8396]_ );
  assign n6415 = ~\new_[8434]_  | ~\new_[12197]_  | ~\new_[7970]_ ;
  assign n6245 = ~\new_[8427]_  | ~\new_[12197]_  | ~\new_[7952]_ ;
  assign n6250 = ~\new_[8485]_  | ~\new_[12339]_  | ~\new_[7968]_ ;
  assign n6255 = ~\new_[8423]_  | ~\new_[12339]_  | ~\new_[7969]_ ;
  assign n6260 = ~\new_[8424]_  | ~\new_[13165]_  | ~\new_[7966]_ ;
  assign n6265 = ~\new_[8425]_  | ~\new_[13165]_  | ~\new_[7961]_ ;
  assign n6275 = ~\new_[8458]_  | ~\new_[13165]_  | ~\new_[7953]_ ;
  assign n6280 = ~\new_[8419]_  | ~\new_[12067]_  | ~\new_[7959]_ ;
  assign n6285 = ~\new_[8474]_  | ~\new_[12067]_  | ~\new_[7954]_ ;
  assign n6875 = ~\new_[8475]_  | ~\new_[12387]_  | ~\new_[7955]_ ;
  assign n6290 = ~\new_[8492]_  | ~\new_[12158]_  | ~\new_[7956]_ ;
  assign n6295 = ~\new_[8554]_  | ~\new_[12244]_  | ~\new_[7957]_ ;
  assign n6845 = ~\new_[8430]_  | ~phy_rst_pad_o | ~\new_[8001]_ ;
  assign n6300 = ~\new_[8488]_  | ~\new_[12158]_  | ~\new_[7958]_ ;
  assign n6305 = ~\new_[8462]_  | ~\new_[12442]_  | ~\new_[7960]_ ;
  assign n6815 = ~\new_[8491]_  | ~\new_[12442]_  | ~\new_[7962]_ ;
  assign n6310 = ~\new_[8478]_  | ~\new_[12244]_  | ~\new_[7965]_ ;
  assign n6215 = ~\new_[12505]_  & (~\new_[8192]_  | ~\new_[8332]_ );
  assign n6685 = ~\new_[12505]_  & (~\new_[8441]_  | ~\new_[8122]_ );
  assign n6010 = ~\new_[12505]_  & (~\new_[8442]_  | ~\new_[8015]_ );
  assign \new_[6934]_  = ~\\u4_u1_csr1_reg[7] ;
  assign n6715 = ~\new_[12804]_  & (~\new_[8483]_  | ~\new_[8115]_ );
  assign n6015 = ~\new_[12849]_  & (~\new_[8480]_  | ~\new_[8017]_ );
  assign n6020 = ~\new_[12505]_  & (~\new_[8443]_  | ~\new_[8018]_ );
  assign n6025 = ~\new_[12849]_  & (~\new_[8444]_  | ~\new_[8113]_ );
  assign n6030 = ~\new_[12804]_  & (~\new_[8445]_  | ~\new_[8157]_ );
  assign n6035 = ~\new_[12804]_  & (~\new_[8446]_  | ~\new_[8117]_ );
  assign n6040 = ~\new_[12804]_  & (~\new_[8447]_  | ~\new_[8114]_ );
  assign n5905 = ~\new_[12505]_  & (~\new_[8490]_  | ~\new_[8019]_ );
  assign n6045 = ~\new_[12804]_  & (~\new_[8509]_  | ~\new_[8020]_ );
  assign n6050 = ~\new_[12849]_  & (~\new_[8448]_  | ~\new_[8135]_ );
  assign n6055 = ~\new_[12505]_  & (~\new_[8021]_  | ~\new_[8479]_ );
  assign n5870 = ~\new_[12849]_  & (~\new_[8449]_  | ~\new_[8022]_ );
  assign n6060 = ~\new_[12849]_  & (~\new_[8023]_  | ~\new_[8418]_ );
  assign n6065 = ~\new_[12505]_  & (~\new_[8024]_  | ~\new_[8468]_ );
  assign n6070 = ~\new_[12849]_  & (~\new_[8450]_  | ~\new_[8127]_ );
  assign n5755 = ~\new_[12505]_  & (~\new_[8499]_  | ~\new_[8118]_ );
  assign n6075 = ~\new_[12505]_  & (~\new_[8459]_  | ~\new_[8025]_ );
  assign n6080 = ~\new_[12245]_  & (~\new_[8451]_  | ~\new_[8123]_ );
  assign n6085 = ~\new_[12505]_  & (~\new_[8452]_  | ~\new_[8119]_ );
  assign n5850 = ~\new_[12505]_  & (~\new_[8484]_  | ~\new_[8026]_ );
  assign n6090 = ~\new_[12849]_  & (~\new_[8454]_  | ~\new_[8027]_ );
  assign \new_[6956]_  = \new_[8560]_  | \new_[12412]_  | \new_[3938]_  | \new_[3940]_ ;
  assign n5795 = ~\new_[9988]_  | ~\new_[8587]_  | ~\new_[8946]_  | ~\new_[9010]_ ;
  assign n6315 = ~\new_[8530]_  | ~\new_[12442]_  | ~\new_[7999]_ ;
  assign \new_[6959]_  = ~\new_[8160]_  & (~\new_[8235]_  | ~\new_[11649]_ );
  assign n6325 = ~\new_[7715]_  & ~\new_[8124]_ ;
  assign n5760 = ~\new_[12505]_  & (~\new_[8075]_  | ~\new_[8460]_ );
  assign n5805 = ~\new_[9736]_  | ~\new_[8585]_  | ~\new_[8616]_  | ~\new_[8644]_ ;
  assign \new_[6963]_  = ~\new_[7705]_  | ~rst_i;
  assign n6770 = ~\new_[8336]_  | ~\new_[12442]_  | ~\new_[8042]_ ;
  assign n6330 = ~\new_[8337]_  | ~\new_[12244]_  | ~\new_[8043]_ ;
  assign n6335 = ~\new_[8339]_  | ~\new_[12244]_  | ~\new_[8044]_ ;
  assign n6340 = ~\new_[8340]_  | ~\new_[12244]_  | ~\new_[8045]_ ;
  assign n6695 = ~\new_[8341]_  | ~\new_[12244]_  | ~\new_[8046]_ ;
  assign n6345 = ~\new_[8342]_  | ~\new_[12244]_  | ~\new_[8047]_ ;
  assign n6730 = ~\new_[8343]_  | ~\new_[12244]_  | ~\new_[8048]_ ;
  assign n6350 = ~\new_[8344]_  | ~\new_[12197]_  | ~\new_[8049]_ ;
  assign n6735 = ~\new_[8345]_  | ~\new_[12258]_  | ~\new_[8050]_ ;
  assign n6355 = ~\new_[8346]_  | ~\new_[12258]_  | ~\new_[8051]_ ;
  assign n6705 = ~\new_[8347]_  | ~\new_[12252]_  | ~\new_[8052]_ ;
  assign n6360 = ~\new_[8348]_  | ~\new_[12258]_  | ~\new_[8053]_ ;
  assign n5885 = ~\new_[8349]_  | ~\new_[12258]_  | ~\new_[8054]_ ;
  assign n6365 = ~\new_[12067]_  | ~\new_[8350]_  | ~\new_[8055]_ ;
  assign n5935 = ~\new_[8351]_  | ~\new_[13162]_  | ~\new_[8056]_ ;
  assign n6370 = ~\new_[8352]_  | ~\new_[13162]_  | ~\new_[8057]_ ;
  assign n5965 = ~\new_[8353]_  | ~\new_[12252]_  | ~\new_[8058]_ ;
  assign n6375 = ~\new_[8354]_  | ~\new_[12197]_  | ~\new_[8059]_ ;
  assign n5945 = ~\new_[12067]_  | ~\new_[8355]_  | ~\new_[8060]_ ;
  assign n6380 = ~\new_[12067]_  | ~\new_[8356]_  | ~\new_[8061]_ ;
  assign n5910 = ~\new_[8357]_  | ~\new_[12067]_  | ~\new_[8062]_ ;
  assign n6385 = ~\new_[8359]_  | ~phy_rst_pad_o | ~\new_[8063]_ ;
  assign n6390 = ~\new_[12067]_  | ~\new_[8360]_  | ~\new_[8064]_ ;
  assign n6395 = ~\new_[8361]_  | ~\new_[12158]_  | ~\new_[8065]_ ;
  assign n5875 = ~\new_[8362]_  | ~\new_[13165]_  | ~\new_[8066]_ ;
  assign n6400 = ~\new_[8363]_  | ~\new_[13165]_  | ~\new_[8067]_ ;
  assign n5835 = ~\new_[8364]_  | ~\new_[13165]_  | ~\new_[8068]_ ;
  assign n6405 = ~\new_[8365]_  | ~\new_[12244]_  | ~\new_[8069]_ ;
  assign n5865 = ~\new_[8367]_  | ~\new_[12244]_  | ~\new_[8070]_ ;
  assign n5765 = ~\new_[8368]_  | ~\new_[12197]_  | ~\new_[8071]_ ;
  assign n5775 = ~\new_[8369]_  | ~\new_[12158]_  | ~\new_[8072]_ ;
  assign n6410 = ~\new_[8370]_  | ~\new_[12158]_  | ~\new_[8073]_ ;
  assign n5800 = ~\new_[9990]_  | ~\new_[8584]_  | ~\new_[8940]_  | ~\new_[8643]_ ;
  assign n6675 = ~\new_[12505]_  & (~\new_[8374]_  | ~\new_[8082]_ );
  assign n6095 = ~\new_[12849]_  & (~\new_[8375]_  | ~\new_[8083]_ );
  assign n6840 = ~\new_[12849]_  & (~\new_[8376]_  | ~\new_[8084]_ );
  assign n6100 = ~\new_[12849]_  & (~\new_[8377]_  | ~\new_[8085]_ );
  assign n6900 = ~\new_[12849]_  & (~\new_[8378]_  | ~\new_[8086]_ );
  assign n6885 = ~\new_[12842]_  & (~\new_[8380]_  | ~\new_[8088]_ );
  assign n6860 = ~\new_[12505]_  & (~\new_[8381]_  | ~\new_[8090]_ );
  assign n6105 = ~\new_[12245]_  & (~\new_[8382]_  | ~\new_[8091]_ );
  assign n6870 = ~\new_[12849]_  & (~\new_[8383]_  | ~\new_[8092]_ );
  assign n6850 = ~\new_[12505]_  & (~\new_[8384]_  | ~\new_[8093]_ );
  assign n6835 = ~\new_[12804]_  & (~\new_[8385]_  | ~\new_[8116]_ );
  assign n6110 = ~\new_[12849]_  & (~\new_[8095]_  | ~\new_[8386]_ );
  assign n6760 = ~\new_[12505]_  & (~\new_[8387]_  | ~\new_[8096]_ );
  assign n6780 = ~\new_[12849]_  & (~\new_[8097]_  | ~\new_[8388]_ );
  assign n6785 = ~\new_[12849]_  & (~\new_[8098]_  | ~\new_[8389]_ );
  assign n6800 = ~\new_[12505]_  & (~\new_[8390]_  | ~\new_[8102]_ );
  assign n6115 = ~\new_[12505]_  & (~\new_[8391]_  | ~\new_[8103]_ );
  assign n6810 = ~\new_[12505]_  & (~\new_[8392]_  | ~\new_[8104]_ );
  assign n6120 = ~\new_[12849]_  & (~\new_[8393]_  | ~\new_[8105]_ );
  assign \new_[7016]_  = \new_[8563]_  | \new_[12290]_  | \new_[3466]_  | \new_[3310]_ ;
  assign n6270 = ~\new_[8477]_  | ~\new_[12244]_  | ~\new_[7967]_ ;
  assign n6125 = ~\new_[12849]_  & (~\new_[8126]_  | ~\new_[8399]_ );
  assign n5825 = ~\new_[8493]_  | ~\new_[12244]_  | ~\new_[7971]_ ;
  assign n6425 = ~\new_[8129]_  | ~\new_[12244]_  | ~\new_[7972]_ ;
  assign n6430 = ~\new_[8494]_  | ~\new_[12197]_  | ~\new_[7973]_ ;
  assign n6435 = ~\new_[8495]_  | ~\new_[12197]_  | ~\new_[7974]_ ;
  assign n5815 = ~\new_[8432]_  | ~\new_[12255]_  | ~\new_[7975]_ ;
  assign n6440 = ~\new_[8011]_  | ~\new_[12255]_  | ~\new_[7976]_ ;
  assign n6445 = ~\new_[8496]_  | ~\new_[12067]_  | ~\new_[7977]_ ;
  assign n6450 = ~\new_[8130]_  | ~\new_[12067]_  | ~\new_[7978]_ ;
  assign n6740 = ~\new_[8131]_  | ~\new_[12244]_  | ~\new_[7979]_ ;
  assign n6455 = ~\new_[8497]_  | ~\new_[12067]_  | ~\new_[7980]_ ;
  assign n6460 = ~\new_[8009]_  | ~\new_[12158]_  | ~\new_[7981]_ ;
  assign n6465 = ~\new_[8498]_  | ~\new_[12158]_  | ~\new_[7982]_ ;
  assign n6880 = ~\new_[8016]_  | ~\new_[12216]_  | ~\new_[7951]_ ;
  assign n6470 = ~\new_[8540]_  | ~\new_[12067]_  | ~\new_[7983]_ ;
  assign n6475 = ~\new_[8489]_  | ~\new_[13162]_  | ~\new_[8000]_ ;
  assign n6480 = ~\new_[8481]_  | ~\new_[13162]_  | ~\new_[7984]_ ;
  assign n6820 = ~\new_[8466]_  | ~\new_[13165]_  | ~\new_[7985]_ ;
  assign n6485 = ~\new_[8463]_  | ~\new_[13165]_  | ~\new_[7986]_ ;
  assign n6490 = ~\new_[8132]_  | ~\new_[12216]_  | ~\new_[7987]_ ;
  assign n6495 = ~\new_[8500]_  | ~\new_[12216]_  | ~\new_[7988]_ ;
  assign n6745 = ~\new_[8501]_  | ~\new_[12216]_  | ~\new_[7989]_ ;
  assign n6505 = ~\new_[8188]_  | ~phy_rst_pad_o | ~\new_[7990]_ ;
  assign n6500 = ~\new_[8502]_  | ~\new_[12216]_  | ~\new_[8002]_ ;
  assign n6690 = ~\new_[8133]_  | ~\new_[12216]_  | ~\new_[7991]_ ;
  assign n6510 = ~\new_[8503]_  | ~\new_[12216]_  | ~\new_[7992]_ ;
  assign n6515 = ~\new_[8504]_  | ~\new_[12197]_  | ~\new_[7993]_ ;
  assign n6520 = ~\new_[8482]_  | ~\new_[12197]_  | ~\new_[7994]_ ;
  assign n6720 = ~\new_[8505]_  | ~\new_[12255]_  | ~\new_[7995]_ ;
  assign n6525 = ~\new_[8507]_  | ~\new_[12255]_  | ~\new_[7996]_ ;
  assign n6725 = ~\new_[8508]_  | ~\new_[12244]_  | ~\new_[7997]_ ;
  assign n6700 = ~\new_[8510]_  | ~\new_[12244]_  | ~\new_[7998]_ ;
  assign n6005 = ~\new_[7654]_ ;
  assign n6130 = ~\new_[12849]_  & (~\new_[8513]_  | ~\new_[8137]_ );
  assign n6135 = ~\new_[12849]_  & (~\new_[8514]_  | ~\new_[8138]_ );
  assign n6140 = ~\new_[12849]_  & (~\new_[8515]_  | ~\new_[8110]_ );
  assign n5920 = ~\new_[12505]_  & (~\new_[8139]_  | ~\new_[8140]_ );
  assign n5960 = ~\new_[12804]_  & (~\new_[8141]_  | ~\new_[8107]_ );
  assign n6145 = ~\new_[12505]_  & (~\new_[8517]_  | ~\new_[8142]_ );
  assign n5915 = ~\new_[12505]_  & (~\new_[8470]_  | ~\new_[8143]_ );
  assign n6150 = ~\new_[12849]_  & (~\new_[8145]_  | ~\new_[8144]_ );
  assign n5880 = ~\new_[12849]_  & (~\new_[8518]_  | ~\new_[8146]_ );
  assign n6155 = ~\new_[12505]_  & (~\new_[8147]_  | ~\new_[8519]_ );
  assign n5900 = ~\new_[12505]_  & (~\new_[8038]_  | ~\new_[8520]_ );
  assign n6160 = ~\new_[12505]_  & (~\new_[8149]_  | ~\new_[8467]_ );
  assign n5890 = ~\new_[12505]_  & (~\new_[8521]_  | ~\new_[8150]_ );
  assign n6165 = ~\new_[12804]_  & (~\new_[8152]_  | ~\new_[8151]_ );
  assign n5770 = ~\new_[12849]_  & (~\new_[8464]_  | ~\new_[8153]_ );
  assign n6170 = ~\new_[12505]_  & (~\new_[8154]_  | ~\new_[8035]_ );
  assign n6175 = ~\new_[12505]_  & (~\new_[8522]_  | ~\new_[8155]_ );
  assign n6180 = ~\new_[12849]_  & (~\new_[8524]_  | ~\new_[8029]_ );
  assign n6185 = ~\new_[12505]_  & (~\new_[8526]_  | ~\new_[8156]_ );
  assign \new_[7070]_  = \new_[8565]_  | \new_[12473]_  | \new_[3686]_  | \new_[3464]_ ;
  assign \new_[7071]_  = ~\new_[9152]_  | ~\new_[7720]_ ;
  assign n6190 = ~\new_[12849]_  & (~\new_[8163]_  | ~\new_[8534]_ );
  assign n6535 = ~\new_[8535]_  | ~\new_[12158]_  | ~\new_[8164]_ ;
  assign n5925 = ~\new_[8536]_  | ~\new_[12158]_  | ~\new_[8166]_ ;
  assign n6540 = ~\new_[8439]_  | ~\new_[12197]_  | ~\new_[8167]_ ;
  assign n5930 = ~\new_[8537]_  | ~\new_[12339]_  | ~\new_[8168]_ ;
  assign n6545 = ~\new_[8538]_  | ~\new_[12197]_  | ~\new_[8169]_ ;
  assign n5810 = ~\new_[8539]_  | ~\new_[12244]_  | ~\new_[8170]_ ;
  assign n6550 = ~\new_[8472]_  | ~\new_[12244]_  | ~\new_[8171]_ ;
  assign n5855 = ~\new_[8471]_  | ~\new_[12197]_  | ~\new_[8172]_ ;
  assign n6555 = ~\new_[8465]_  | ~\new_[12244]_  | ~\new_[8173]_ ;
  assign n6560 = ~\new_[8532]_  | ~\new_[12244]_  | ~\new_[8174]_ ;
  assign n6565 = ~\new_[8541]_  | ~\new_[12244]_  | ~\new_[8175]_ ;
  assign n5820 = ~\new_[8542]_  | ~\new_[12244]_  | ~\new_[8176]_ ;
  assign n6570 = ~\new_[8511]_  | ~\new_[12387]_  | ~\new_[8078]_ ;
  assign n6575 = ~\new_[8438]_  | ~\new_[12387]_  | ~\new_[8177]_ ;
  assign n6580 = ~\new_[8531]_  | ~\new_[13162]_  | ~\new_[8028]_ ;
  assign n5830 = ~\new_[8529]_  | ~\new_[13162]_  | ~\new_[8178]_ ;
  assign n6585 = ~\new_[8543]_  | ~\new_[12491]_  | ~\new_[8111]_ ;
  assign n6590 = ~\new_[8457]_  | ~\new_[12491]_  | ~\new_[8179]_ ;
  assign n6595 = ~\new_[8486]_  | ~\new_[12491]_  | ~\new_[8196]_ ;
  assign n5780 = ~\new_[8436]_  | ~\new_[12158]_  | ~\new_[8180]_ ;
  assign n5785 = ~\new_[8557]_  | ~\new_[12491]_  | ~\new_[8195]_ ;
  assign n6660 = ~\new_[8544]_  | ~phy_rst_pad_o | ~\new_[8182]_ ;
  assign n6600 = ~\new_[8545]_  | ~\new_[12158]_  | ~\new_[8108]_ ;
  assign n6830 = ~\new_[8428]_  | ~\new_[12158]_  | ~\new_[8077]_ ;
  assign n6605 = ~\new_[8546]_  | ~\new_[12158]_  | ~\new_[8183]_ ;
  assign n6910 = ~\new_[8556]_  | ~\new_[12197]_  | ~\new_[8184]_ ;
  assign n6610 = ~\new_[8552]_  | ~\new_[12197]_  | ~\new_[8185]_ ;
  assign n6905 = ~\new_[8547]_  | ~\new_[13165]_  | ~\new_[8186]_ ;
  assign n6890 = ~\new_[8548]_  | ~\new_[13165]_  | ~\new_[8031]_ ;
  assign n6615 = ~\new_[8555]_  | ~\new_[12252]_  | ~\new_[8159]_ ;
  assign n6895 = ~\new_[8553]_  | ~\new_[12252]_  | ~\new_[8197]_ ;
  assign n6620 = ~\new_[8549]_  | ~\new_[13165]_  | ~\new_[8187]_ ;
  assign n6195 = ~\new_[12849]_  & (~\new_[8394]_  | ~\new_[8112]_ );
  assign n6865 = ~\new_[12849]_  & (~\new_[8003]_  | ~\new_[8106]_ );
  assign n6200 = ~\new_[12849]_  & (~\new_[8373]_  | ~\new_[8081]_ );
  assign n6855 = ~\new_[12849]_  & (~\new_[8372]_  | ~\new_[8080]_ );
  assign n6205 = ~\new_[12245]_  & (~\new_[7963]_  | ~\new_[8032]_ );
  assign n6790 = ~\new_[12849]_  & (~\new_[8407]_  | ~\new_[8033]_ );
  assign n6210 = ~\new_[12849]_  & (~\new_[8004]_  | ~\new_[8030]_ );
  assign n6825 = ~\new_[12505]_  & (~\new_[8334]_  | ~\new_[8191]_ );
  assign n6805 = ~\new_[12505]_  & (~\new_[8005]_  | ~\new_[8013]_ );
  assign n6220 = ~\new_[12505]_  & (~\new_[8012]_  | ~\new_[8331]_ );
  assign n6795 = ~\new_[12849]_  & (~\new_[8193]_  | ~\new_[8408]_ );
  assign n6225 = ~\new_[12849]_  & (~\new_[8409]_  | ~\new_[8158]_ );
  assign n6775 = ~\new_[12849]_  & (~\new_[8410]_  | ~\new_[8010]_ );
  assign n6230 = ~\new_[12245]_  & (~\new_[8405]_  | ~\new_[8109]_ );
  assign n6765 = ~\new_[12505]_  & (~\new_[8411]_  | ~\new_[8034]_ );
  assign n6240 = ~\new_[12849]_  & (~\new_[8006]_  | ~\new_[8136]_ );
  assign n6235 = ~\new_[12505]_  & (~\new_[8412]_  | ~\new_[8094]_ );
  assign n6710 = ~\new_[12849]_  & (~\new_[8404]_  | ~\new_[8194]_ );
  assign \new_[7123]_  = \new_[8567]_  | \new_[12470]_  | \new_[3879]_  | \new_[3787]_ ;
  assign n5995 = ~\new_[8259]_  & (~\new_[8199]_  | ~\new_[9337]_ );
  assign \new_[7125]_  = ~\new_[7937]_  & (~\new_[10944]_  | ~\new_[8238]_ );
  assign n6420 = ~\new_[7600]_  | (~\new_[9429]_  & ~\new_[12259]_ );
  assign n6625 = ~\new_[7592]_  | (~\new_[9445]_  & ~\new_[12259]_ );
  assign n6320 = ~\new_[7717]_  | (~\new_[12259]_  & ~\new_[9426]_ );
  assign n6530 = ~\new_[7599]_  | (~\new_[9430]_  & ~\new_[12259]_ );
  assign \new_[7130]_  = \\u1_u2_state_reg[7] ;
  assign \new_[7131]_  = (~\new_[8218]_  | ~\new_[8631]_ ) & (~\new_[8827]_  | ~\new_[8652]_ );
  assign \new_[7132]_  = ~\new_[9065]_  | (~\new_[7942]_  & ~\new_[3282]_ );
  assign \new_[7133]_  = ~\new_[8693]_  | (~\new_[7941]_  & ~\new_[3308]_ );
  assign \new_[7134]_  = (~\new_[8203]_  | ~\new_[3881]_ ) & (~\new_[8568]_  | ~\new_[9602]_ );
  assign n5940 = ~\new_[7716]_  & ~\new_[12849]_ ;
  assign \new_[7136]_  = \\u4_dout_reg[10] ;
  assign \new_[7137]_  = \\u4_dout_reg[11] ;
  assign \new_[7138]_  = \\u4_dout_reg[9] ;
  assign \new_[7139]_  = ~\new_[7723]_  & ~\new_[13363]_ ;
  assign n5860 = \new_[8586]_  | \new_[9005]_  | \new_[9271]_  | \new_[9004]_ ;
  assign \new_[7141]_  = ~\new_[8568]_  & ~\new_[4091]_ ;
  assign \new_[7142]_  = ~\new_[8568]_  & ~\new_[4092]_ ;
  assign \new_[7143]_  = ~\new_[14329]_  & ~\new_[2871]_ ;
  assign \new_[7144]_  = ~\new_[7722]_  & ~\new_[13289]_ ;
  assign \new_[7145]_  = ~\new_[5761]_  & (~\new_[8914]_  | ~\new_[7866]_ );
  assign \new_[7146]_  = ~\new_[10491]_  | ~\new_[4791]_  | ~\new_[7736]_  | ~\new_[10126]_ ;
  assign \new_[7147]_  = ~\\u4_u2_iena_reg[1] ;
  assign \new_[7148]_  = ~\\u4_u2_iena_reg[3] ;
  assign \new_[7149]_  = ~\\u4_u2_iena_reg[5] ;
  assign \new_[7150]_  = ~\\u4_u2_ienb_reg[0] ;
  assign \new_[7151]_  = ~\\u4_u2_ienb_reg[1] ;
  assign \new_[7152]_  = ~\\u4_u2_ienb_reg[4] ;
  assign \new_[7153]_  = ~\\u4_u2_ienb_reg[3] ;
  assign \new_[7154]_  = ~\\u4_u3_iena_reg[0] ;
  assign \new_[7155]_  = ~\\u4_u3_iena_reg[2] ;
  assign \new_[7156]_  = ~\\u4_u0_iena_reg[1] ;
  assign \new_[7157]_  = ~\\u4_u0_iena_reg[2] ;
  assign \new_[7158]_  = ~\\u4_u0_iena_reg[3] ;
  assign \new_[7159]_  = ~\\u4_u0_iena_reg[5] ;
  assign \new_[7160]_  = ~\\u4_u0_ienb_reg[1] ;
  assign \new_[7161]_  = ~\\u4_u0_ienb_reg[4] ;
  assign \new_[7162]_  = ~\\u4_u0_ienb_reg[3] ;
  assign \new_[7163]_  = ~\\u4_u1_iena_reg[2] ;
  assign \new_[7164]_  = ~\\u4_u1_ienb_reg[4] ;
  assign n6630 = \new_[8209]_  ? \wb_addr_i[17]  : \sram_data_i[14] ;
  assign \new_[7166]_  = \new_[2038]_  ? \new_[8202]_  : \new_[2174]_ ;
  assign \new_[7167]_  = \\u4_dout_reg[12] ;
  assign \new_[7168]_  = \new_[4926]_  ? \new_[8202]_  : \new_[13977]_ ;
  assign \new_[7169]_  = ~\new_[7826]_  | ~\new_[12501]_ ;
  assign \new_[7170]_  = ~\new_[7827]_  | ~\new_[12440]_ ;
  assign \new_[7171]_  = ~\new_[7831]_  | ~\new_[12618]_ ;
  assign \new_[7172]_  = \new_[4765]_  ? \new_[8202]_  : \new_[13844]_ ;
  assign \new_[7173]_  = ~\new_[7754]_  & (~\new_[14636]_  | ~\new_[2340]_ );
  assign \new_[7174]_  = ~\new_[7755]_  & (~\new_[14636]_  | ~\new_[2341]_ );
  assign \new_[7175]_  = ~\new_[7832]_  | ~\new_[12673]_ ;
  assign \new_[7176]_  = ~\new_[8208]_  | ~\new_[7604]_ ;
  assign \new_[7177]_  = ~\\u4_u0_ienb_reg[5] ;
  assign \new_[7178]_  = ~\new_[7436]_ ;
  assign \new_[7179]_  = ~\\u4_u1_ienb_reg[0] ;
  assign \new_[7180]_  = ~\new_[8162]_  & (~\new_[7875]_  | ~\new_[3711]_ );
  assign \new_[7181]_  = \new_[7845]_  | \new_[2474]_ ;
  assign \new_[7182]_  = \new_[8600]_  | \new_[13796]_ ;
  assign \new_[7183]_  = \new_[8600]_  | \new_[2876]_ ;
  assign \new_[7184]_  = \new_[8224]_  | \new_[2875]_ ;
  assign \new_[7185]_  = ~\new_[7846]_  | ~\new_[14205]_ ;
  assign \new_[7186]_  = ~\new_[7846]_  | ~\new_[13568]_ ;
  assign \new_[7187]_  = ~\new_[7848]_  | ~\new_[2870]_ ;
  assign \new_[7188]_  = ~\new_[7442]_ ;
  assign \new_[7189]_  = ~\new_[7848]_  | ~\new_[14174]_ ;
  assign \new_[7190]_  = ~\new_[7848]_  & ~\new_[14174]_ ;
  assign \new_[7191]_  = ~\new_[8600]_  | ~\new_[13796]_ ;
  assign \new_[7192]_  = \new_[14422]_  | \new_[2475]_ ;
  assign \new_[7193]_  = \new_[7846]_  & \new_[2475]_ ;
  assign \new_[7194]_  = ~\new_[7447]_ ;
  assign \new_[7195]_  = \new_[14276]_  | \new_[13953]_ ;
  assign \new_[7196]_  = ~\new_[14276]_  | ~\new_[13953]_ ;
  assign \new_[7197]_  = ~\new_[8224]_  & ~\new_[13811]_ ;
  assign \new_[7198]_  = ~\\u4_u0_ienb_reg[2] ;
  assign \new_[7199]_  = ~\new_[7786]_  & ~n7635;
  assign \new_[7200]_  = ~\\u4_u0_iena_reg[4] ;
  assign \new_[7201]_  = ~\new_[7778]_  & ~\new_[9275]_ ;
  assign \new_[7202]_  = ~\\u4_u0_ienb_reg[0] ;
  assign \new_[7203]_  = ~\\u4_u3_dma_out_left_reg[11] ;
  assign \new_[7204]_  = ~\\u4_u2_dma_out_left_reg[11] ;
  assign \new_[7205]_  = ~\\u4_u2_iena_reg[0] ;
  assign \new_[7206]_  = \\u5_state_reg[3] ;
  assign \new_[7207]_  = ~\new_[7470]_ ;
  assign \new_[7208]_  = ~\new_[7471]_ ;
  assign \new_[7209]_  = ~\new_[8236]_  | ~\new_[6290]_ ;
  assign \new_[7210]_  = ~\new_[8236]_  | ~\new_[6538]_ ;
  assign \new_[7211]_  = ~\new_[8236]_  | ~\new_[14244]_ ;
  assign \new_[7212]_  = ~\new_[8236]_  | ~\new_[13986]_ ;
  assign \new_[7213]_  = ~\new_[8236]_  | ~\new_[13578]_ ;
  assign \new_[7214]_  = ~\new_[8236]_  | ~\new_[5504]_ ;
  assign \new_[7215]_  = ~\new_[8236]_  | ~\new_[5503]_ ;
  assign \new_[7216]_  = ~\new_[8236]_  | ~\new_[14010]_ ;
  assign \new_[7217]_  = ~\new_[8236]_  | ~\new_[13686]_ ;
  assign \new_[7218]_  = ~\new_[8236]_  | ~\new_[13607]_ ;
  assign \new_[7219]_  = ~\new_[8236]_  | ~\new_[14267]_ ;
  assign \new_[7220]_  = ~\new_[8236]_  | ~\new_[14240]_ ;
  assign \new_[7221]_  = ~\new_[8236]_  | ~\new_[6485]_ ;
  assign \new_[7222]_  = ~\new_[8236]_  | ~\new_[13833]_ ;
  assign \new_[7223]_  = ~\new_[8236]_  | ~\new_[13587]_ ;
  assign \new_[7224]_  = ~\new_[8236]_  | ~\new_[13922]_ ;
  assign \new_[7225]_  = ~\new_[8236]_  | ~\new_[13503]_ ;
  assign \new_[7226]_  = ~\new_[8236]_  | ~\new_[13688]_ ;
  assign \new_[7227]_  = ~\new_[8236]_  | ~\new_[13730]_ ;
  assign \new_[7228]_  = ~\new_[8236]_  | ~\new_[13782]_ ;
  assign \new_[7229]_  = ~\new_[8236]_  | ~\new_[14159]_ ;
  assign \new_[7230]_  = ~\new_[8236]_  | ~\new_[13952]_ ;
  assign \new_[7231]_  = ~\new_[8236]_  | ~\new_[13818]_ ;
  assign \new_[7232]_  = ~\new_[8236]_  | ~\new_[13789]_ ;
  assign \new_[7233]_  = ~\new_[8236]_  | ~\new_[13836]_ ;
  assign \new_[7234]_  = ~\new_[8236]_  | ~\new_[13609]_ ;
  assign \new_[7235]_  = ~\new_[8236]_  | ~\new_[13856]_ ;
  assign \new_[7236]_  = ~\new_[8236]_  | ~\new_[13758]_ ;
  assign \new_[7237]_  = ~\new_[8236]_  | ~\new_[14011]_ ;
  assign \new_[7238]_  = ~\new_[8236]_  | ~\new_[14030]_ ;
  assign \new_[7239]_  = ~\new_[8236]_  | ~\new_[14250]_ ;
  assign \new_[7240]_  = ~\new_[8236]_  | ~\new_[14162]_ ;
  assign \new_[7241]_  = ~\new_[8236]_  | ~\new_[14201]_ ;
  assign \new_[7242]_  = ~\new_[8236]_  | ~\new_[13843]_ ;
  assign \new_[7243]_  = ~\new_[8236]_  | ~\new_[13750]_ ;
  assign \new_[7244]_  = ~\new_[8236]_  | ~\new_[14190]_ ;
  assign \new_[7245]_  = ~\new_[8236]_  | ~\new_[14207]_ ;
  assign \new_[7246]_  = ~\new_[8236]_  | ~\new_[13994]_ ;
  assign \new_[7247]_  = ~\new_[8236]_  | ~\new_[13841]_ ;
  assign \new_[7248]_  = ~\new_[8236]_  | ~\new_[13931]_ ;
  assign \new_[7249]_  = ~\new_[7581]_  | ~\new_[10849]_ ;
  assign \new_[7250]_  = ~\new_[8236]_  | ~\new_[13883]_ ;
  assign \new_[7251]_  = ~\new_[8236]_  | ~\new_[5604]_ ;
  assign \new_[7252]_  = ~\new_[8236]_  | ~\new_[13535]_ ;
  assign \new_[7253]_  = ~\new_[8236]_  | ~\new_[13959]_ ;
  assign \new_[7254]_  = ~\new_[8236]_  | ~\new_[14027]_ ;
  assign \new_[7255]_  = ~\new_[8236]_  | ~\new_[13996]_ ;
  assign \new_[7256]_  = ~\new_[8236]_  | ~\new_[13560]_ ;
  assign \new_[7257]_  = ~\new_[8236]_  | ~\new_[13528]_ ;
  assign \new_[7258]_  = ~\\u4_u1_ienb_reg[1] ;
  assign n6635 = ~\new_[7563]_  & ~\new_[12794]_ ;
  assign n6640 = ~\new_[7562]_  & ~\new_[12794]_ ;
  assign n6645 = ~\new_[7564]_  & ~\new_[12794]_ ;
  assign n6680 = ~\new_[7565]_  & ~\new_[12794]_ ;
  assign \new_[7263]_  = ~\new_[7583]_  | ~\new_[10849]_ ;
  assign \new_[7264]_  = ~\new_[5502]_  | ~\new_[7860]_ ;
  assign \new_[7265]_  = ~\new_[7557]_  | ~\new_[5604]_ ;
  assign \new_[7266]_  = ~\new_[7584]_  | ~\new_[10849]_ ;
  assign \new_[7267]_  = ~\new_[7560]_  | ~\new_[2178]_ ;
  assign \new_[7268]_  = ~\new_[7859]_  | ~\new_[2177]_ ;
  assign \new_[7269]_  = ~\new_[7764]_  & (~\new_[4819]_  | ~\new_[14508]_ );
  assign n6650 = ~\new_[7566]_  | ~phy_rst_pad_o;
  assign n6655 = ~\new_[7567]_  | ~phy_rst_pad_o;
  assign n5790 = ~\new_[7568]_  | ~phy_rst_pad_o;
  assign n5895 = ~\new_[7569]_  | ~phy_rst_pad_o;
  assign n6665 = \new_[9313]_  | \new_[7849]_ ;
  assign \new_[7275]_  = ~\new_[5504]_  | ~\new_[7557]_ ;
  assign \new_[7276]_  = ~\new_[7860]_  | ~\new_[5503]_ ;
  assign \new_[7277]_  = ~\\u4_u2_ienb_reg[5] ;
  assign \new_[7278]_  = ~\\u4_u0_iena_reg[0] ;
  assign \new_[7279]_  = ~\new_[7560]_  | ~\new_[2266]_ ;
  assign \new_[7280]_  = ~\new_[7859]_  | ~\new_[2136]_ ;
  assign \new_[7281]_  = ~\new_[7582]_  | (~\new_[9665]_  & ~\new_[9407]_ );
  assign \new_[7282]_  = ~\new_[8639]_  | (~\new_[7872]_  & ~\new_[9857]_ );
  assign \new_[7283]_  = \new_[8639]_  & \new_[7850]_ ;
  assign \new_[7284]_  = ~\new_[7855]_  & (~\new_[8247]_  | ~\new_[5766]_ );
  assign \new_[7285]_  = ~\\u4_u2_ienb_reg[2] ;
  assign \new_[7286]_  = ~\\u4_u2_iena_reg[2] ;
  assign \new_[7287]_  = ~\new_[7587]_  | (~\new_[9673]_  & ~\new_[9408]_ );
  assign \new_[7288]_  = ~\new_[7589]_  | (~\new_[9674]_  & ~\new_[9409]_ );
  assign \new_[7289]_  = (~\new_[8216]_  & ~\new_[8610]_ ) | (~\new_[12383]_  & ~\new_[9032]_ );
  assign \new_[7290]_  = ~\new_[7591]_  | (~\new_[9678]_  & ~\new_[9410]_ );
  assign \new_[7291]_  = ~\\u4_u2_iena_reg[4] ;
  assign \new_[7292]_  = ~\new_[7541]_ ;
  assign \new_[7293]_  = ~\new_[7576]_  & (~\new_[11159]_  | ~\new_[10455]_ );
  assign \new_[7294]_  = ~\new_[7577]_  & (~\new_[10857]_  | ~\new_[10701]_ );
  assign \new_[7295]_  = ~\new_[7578]_  & (~\new_[10861]_  | ~\new_[10456]_ );
  assign \new_[7296]_  = ~\new_[7579]_  & (~\new_[10853]_  | ~\new_[10459]_ );
  assign \new_[7297]_  = ~\\u4_u1_ienb_reg[2] ;
  assign \new_[7298]_  = ~\new_[7540]_ ;
  assign \new_[7299]_  = u1_u2_rx_data_done_r2_reg;
  assign n6750 = u1_u2_wr_done_r_reg;
  assign \new_[7301]_  = ~\\u4_u1_ienb_reg[3] ;
  assign \new_[7302]_  = ~\\u4_u1_ienb_reg[5] ;
  assign \new_[7303]_  = \new_[3932]_  ^ \new_[7885]_ ;
  assign \new_[7304]_  = \new_[3313]_  ^ \new_[7887]_ ;
  assign \new_[7305]_  = \new_[3468]_  ^ \new_[7888]_ ;
  assign \new_[7306]_  = \new_[3671]_  ^ \new_[7886]_ ;
  assign \new_[7307]_  = ~\new_[7546]_ ;
  assign \new_[7308]_  = ~\new_[7550]_ ;
  assign \new_[7309]_  = ~\new_[7551]_ ;
  assign \new_[7310]_  = ~\\u4_u2_csr1_reg[7] ;
  assign \new_[7311]_  = ~\new_[7858]_ ;
  assign n6755 = n8235 | n7550;
  assign \new_[7313]_  = ~\new_[7554]_ ;
  assign \new_[7314]_  = \new_[7866]_  & \new_[12812]_ ;
  assign \new_[7315]_  = ~\new_[7560]_ ;
  assign \new_[7316]_  = ~\new_[8636]_  | (~\new_[8266]_  & ~\new_[12099]_ );
  assign \new_[7317]_  = ~\new_[7844]_ ;
  assign \new_[7318]_  = ~\new_[9885]_  | ~\new_[8734]_  | ~\new_[10889]_  | ~\new_[12969]_ ;
  assign \new_[7319]_  = ~\new_[9592]_  | ~\new_[8749]_  | ~\new_[10836]_  | ~\new_[13243]_ ;
  assign \new_[7320]_  = ~\new_[8913]_  | ~\new_[11502]_  | ~\new_[11078]_  | ~\new_[11809]_ ;
  assign \new_[7321]_  = ~\new_[13413]_  | ~\new_[7891]_  | ~\new_[8297]_ ;
  assign \new_[7322]_  = ~\new_[10462]_  | ~\new_[11492]_  | ~\new_[7907]_  | ~\new_[11794]_ ;
  assign \new_[7323]_  = ~\new_[7880]_  | ~\new_[13649]_ ;
  assign n6955 = ~\new_[7915]_  & ~\new_[12842]_ ;
  assign n7095 = ~\new_[7916]_  & ~\new_[12842]_ ;
  assign n6945 = ~\new_[7917]_  & ~\new_[13296]_ ;
  assign n7100 = ~\new_[7918]_  & ~\new_[12245]_ ;
  assign n6950 = ~\new_[7919]_  & ~\new_[12842]_ ;
  assign n7105 = ~\new_[7920]_  & ~\new_[12842]_ ;
  assign n7110 = ~\new_[7921]_  & ~\new_[12842]_ ;
  assign n7115 = ~\new_[7922]_  & ~\new_[12245]_ ;
  assign n6935 = ~\new_[7923]_  & ~\new_[12842]_ ;
  assign n7120 = ~\new_[7924]_  & ~\new_[12842]_ ;
  assign n7125 = ~\new_[7925]_  & ~\new_[12245]_ ;
  assign n7130 = ~\new_[7926]_  & ~\new_[13296]_ ;
  assign n6940 = ~\new_[7927]_  & ~\new_[12245]_ ;
  assign n7135 = ~\new_[7928]_  & ~\new_[13296]_ ;
  assign n7140 = ~\new_[7929]_  & ~\new_[13296]_ ;
  assign n7145 = ~\new_[7930]_  & ~\new_[13296]_ ;
  assign n7195 = ~\new_[7931]_  & ~\new_[12842]_ ;
  assign n7150 = ~\new_[7932]_  & ~\new_[13296]_ ;
  assign n6990 = ~\new_[8997]_  | ~\new_[8896]_  | ~\new_[9993]_  | ~\new_[8582]_ ;
  assign n7020 = ~\new_[9001]_  | ~\new_[8872]_  | ~\new_[9735]_  | ~\new_[8589]_ ;
  assign \new_[7344]_  = ~\new_[7881]_  | ~\new_[14001]_ ;
  assign \new_[7345]_  = ~\new_[7881]_  | ~\new_[13264]_ ;
  assign \new_[7346]_  = ~\new_[7880]_  | ~\new_[13372]_ ;
  assign \new_[7347]_  = ~\new_[7882]_  | ~\new_[13926]_ ;
  assign \new_[7348]_  = ~\new_[7882]_  | ~\new_[13440]_ ;
  assign n6965 = ~\new_[8988]_  | ~\new_[8866]_  | ~\new_[9999]_  | ~\new_[8579]_ ;
  assign \new_[7350]_  = (~\new_[8291]_  | ~\new_[3938]_ ) & (~\new_[8719]_  | ~\new_[3940]_ );
  assign n7200 = ~\new_[7896]_  | (~\new_[8692]_  & ~\new_[12423]_ );
  assign \new_[7352]_  = ~\new_[7892]_  & (~\new_[12088]_  | ~\new_[10297]_ );
  assign \new_[7353]_  = ~\new_[7895]_  & (~\new_[12079]_  | ~\new_[10296]_ );
  assign \new_[7354]_  = ~\new_[7901]_  & (~\new_[12165]_  | ~\new_[10295]_ );
  assign \new_[7355]_  = ~\new_[7905]_  & (~\new_[11876]_  | ~\new_[10298]_ );
  assign \new_[7356]_  = \new_[7890]_  & \new_[9679]_ ;
  assign \new_[7357]_  = \new_[7894]_  & \new_[9666]_ ;
  assign \new_[7358]_  = \new_[7898]_  & \new_[9670]_ ;
  assign \new_[7359]_  = \new_[7903]_  & \new_[9440]_ ;
  assign n7205 = \new_[12337]_  ^ \new_[8310]_ ;
  assign \new_[7361]_  = ~\new_[8206]_  | ~\new_[13372]_ ;
  assign n7070 = ~\new_[8124]_  & (~\new_[8618]_  | ~\new_[14119]_ );
  assign n7000 = ~\new_[9012]_  | ~\new_[8867]_  | ~\new_[9772]_  | ~\new_[8942]_ ;
  assign n6970 = ~\new_[9008]_  | ~\new_[8863]_  | ~\new_[9775]_  | ~\new_[8611]_ ;
  assign \new_[7365]_  = ~\new_[7899]_  | ~\new_[3310]_ ;
  assign \new_[7366]_  = ~\new_[8292]_  | ~\new_[7948]_ ;
  assign \new_[7367]_  = ~\new_[7603]_ ;
  assign \new_[7368]_  = ~\new_[8861]_  & (~\new_[8469]_  | ~\new_[9086]_ );
  assign \new_[7369]_  = ~\new_[7899]_  | ~\new_[7944]_ ;
  assign \new_[7370]_  = ~\new_[7824]_ ;
  assign n7165 = ~\new_[8437]_  | ~\new_[12197]_  | ~\new_[8330]_ ;
  assign n7080 = ~\new_[8455]_  | ~\new_[12197]_  | ~\new_[8335]_ ;
  assign n7055 = ~\new_[8421]_  | ~\new_[12339]_  | ~\new_[8402]_ ;
  assign n7025 = ~\new_[8435]_  | ~\new_[13165]_  | ~\new_[8397]_ ;
  assign n6920 = ~\new_[8426]_  | ~\new_[12158]_  | ~\new_[8414]_ ;
  assign n7155 = ~\new_[8550]_  | ~\new_[12067]_  | ~\new_[8415]_ ;
  assign n6960 = ~\new_[8528]_  | ~\new_[12067]_  | ~\new_[8327]_ ;
  assign n6915 = ~\new_[8420]_  | ~\new_[13165]_  | ~\new_[8328]_ ;
  assign \new_[7379]_  = (~\new_[8306]_  | ~\new_[3481]_ ) & (~\new_[9126]_  | ~\new_[3479]_ );
  assign n7230 = ~\new_[8429]_  | ~\new_[12244]_  | ~\new_[8400]_ ;
  assign n7220 = ~\new_[8431]_  | ~\new_[12442]_  | ~\new_[8329]_ ;
  assign n7160 = ~\new_[8433]_  | ~\new_[12244]_  | ~\new_[8401]_ ;
  assign n7215 = ~\new_[8456]_  | ~\new_[12244]_  | ~\new_[8325]_ ;
  assign n7190 = ~\new_[12842]_  & (~\new_[8461]_  | ~\new_[8779]_ );
  assign n7060 = ~\new_[8422]_  | ~\new_[12158]_  | ~\new_[8326]_ ;
  assign \new_[7386]_  = ~\new_[7936]_  | ~\new_[12628]_ ;
  assign n7050 = ~\new_[12842]_  & (~\new_[8516]_  | ~\new_[8797]_ );
  assign \new_[7388]_  = ~\new_[7878]_  | ~\new_[3464]_ ;
  assign \new_[7389]_  = ~\new_[7935]_  | ~\new_[13286]_ ;
  assign \new_[7390]_  = ~\new_[9147]_  | ~\new_[7938]_ ;
  assign \new_[7391]_  = ~\new_[9151]_  | ~\new_[8211]_ ;
  assign n7210 = ~\new_[12842]_  & (~\new_[8406]_  | ~\new_[8801]_ );
  assign n7010 = ~\new_[9019]_  | ~\new_[8897]_  | ~\new_[9773]_  | ~\new_[8943]_ ;
  assign \new_[7394]_  = ~\new_[7870]_  | ~\new_[3787]_ ;
  assign n6930 = ~\new_[8998]_  | ~\new_[8900]_  | ~\new_[9669]_  | ~\new_[8846]_ ;
  assign \new_[7396]_  = \new_[3311]_  ? \new_[8568]_  : \new_[9852]_ ;
  assign \new_[7397]_  = (~\new_[8533]_  | ~\new_[12416]_ ) & (~\new_[9197]_  | ~\new_[8978]_ );
  assign \new_[7398]_  = (~\new_[8827]_  | ~\new_[8269]_ ) & (~\new_[9516]_  | ~\new_[9218]_ );
  assign n6980 = ~\new_[8986]_  | ~\new_[8894]_  | ~\new_[9770]_  | ~\new_[8613]_ ;
  assign \new_[7400]_  = ~\new_[8201]_  & (~\new_[4842]_  | ~\new_[14508]_ );
  assign \new_[7401]_  = ~\new_[7692]_ ;
  assign \new_[7402]_  = \new_[4069]_  ^ \new_[8571]_ ;
  assign \new_[7403]_  = \new_[3312]_  ^ \new_[8570]_ ;
  assign \new_[7404]_  = \new_[3467]_  ^ \new_[8572]_ ;
  assign \new_[7405]_  = \new_[3687]_  ^ \new_[8573]_ ;
  assign \new_[7406]_  = ~\new_[7705]_ ;
  assign n7225 = ~\new_[12849]_  & (~\new_[8951]_  | ~\new_[8576]_ );
  assign \new_[7408]_  = ~\new_[7942]_  | ~\new_[3790]_ ;
  assign \new_[7409]_  = ~\new_[14421]_  & ~\new_[4799]_ ;
  assign \new_[7410]_  = ~\new_[14450]_  & ~\new_[4802]_ ;
  assign \new_[7411]_  = ~\new_[7945]_  | ~phy_rst_pad_o;
  assign \new_[7412]_  = ~\new_[14450]_  & ~\new_[2857]_ ;
  assign \new_[7413]_  = ~\new_[7941]_  | ~\new_[3462]_ ;
  assign \new_[7414]_  = ~\new_[7946]_  | ~phy_rst_pad_o;
  assign \new_[7415]_  = ~\new_[9463]_  | ~\new_[9140]_  | ~\new_[10097]_  | ~\new_[9565]_ ;
  assign \new_[7416]_  = ~\new_[7950]_  & (~\new_[9526]_  | ~\new_[8591]_ );
  assign \new_[7417]_  = ~\new_[7947]_  & ~\new_[13417]_ ;
  assign \new_[7418]_  = ~\new_[7943]_  | ~phy_rst_pad_o;
  assign \new_[7419]_  = ~\new_[8592]_  | ~\new_[9184]_  | ~\new_[8621]_ ;
  assign \new_[7420]_  = ~\new_[6013]_  & (~\new_[8914]_  | ~\new_[8247]_ );
  assign n7015 = ~\new_[8999]_  | ~\new_[8871]_  | ~\new_[9734]_  | ~\new_[8901]_ ;
  assign n6985 = ~\new_[8987]_  | ~\new_[8895]_  | ~\new_[9777]_  | ~\new_[8939]_ ;
  assign \new_[7423]_  = ~\new_[8588]_  | (~\new_[8605]_  & ~\new_[8965]_ );
  assign \new_[7424]_  = ~\new_[8207]_  | ~\new_[13264]_ ;
  assign \new_[7425]_  = ~\new_[8208]_  | ~\new_[13364]_ ;
  assign \new_[7426]_  = ~\new_[12911]_  | ~\new_[8220]_  | ~\new_[8282]_ ;
  assign \new_[7427]_  = \\u4_dout_reg[13] ;
  assign \new_[7428]_  = \\u4_dout_reg[15] ;
  assign \new_[7429]_  = ~\new_[8037]_  | (~\new_[9106]_  & ~\new_[4766]_ );
  assign \new_[7430]_  = ~\new_[8040]_  | (~\new_[9106]_  & ~\new_[4767]_ );
  assign \new_[7431]_  = ~\new_[8210]_  | ~\new_[13440]_ ;
  assign \new_[7432]_  = ~\new_[14634]_  & ~\new_[8638]_ ;
  assign \new_[7433]_  = ~\new_[8207]_  | ~\new_[7881]_ ;
  assign \new_[7434]_  = ~\new_[8206]_  | ~\new_[7880]_ ;
  assign \new_[7435]_  = ~\new_[8210]_  | ~\new_[7882]_ ;
  assign \new_[7436]_  = ~\new_[7735]_ ;
  assign \new_[7437]_  = ~\new_[8487]_  & (~\new_[8281]_  | ~\new_[3504]_ );
  assign \new_[7438]_  = \new_[8225]_  | \new_[4798]_ ;
  assign \new_[7439]_  = ~\new_[8222]_  | ~\new_[14790]_ ;
  assign \new_[7440]_  = ~\new_[8602]_  | ~\new_[13568]_ ;
  assign \new_[7441]_  = \new_[8601]_  | \new_[2874]_ ;
  assign \new_[7442]_  = ~\new_[8603]_  & ~\new_[14264]_ ;
  assign \new_[7443]_  = ~\new_[8603]_  | ~\new_[14264]_ ;
  assign \new_[7444]_  = ~\new_[7744]_ ;
  assign \new_[7445]_  = ~\new_[8224]_  | ~\new_[13811]_ ;
  assign \new_[7446]_  = \new_[8602]_  & \new_[2503]_ ;
  assign \new_[7447]_  = ~\new_[8601]_  & ~\new_[13919]_ ;
  assign \new_[7448]_  = \new_[14270]_  | \new_[13667]_ ;
  assign \new_[7449]_  = ~\new_[14270]_  | ~\new_[13667]_ ;
  assign \new_[7450]_  = ~\new_[14792]_  & ~\new_[4796]_ ;
  assign n7075 = ~\new_[8219]_  | ~\new_[9146]_ ;
  assign \new_[7452]_  = ~\new_[8202]_  | ~\new_[2135]_ ;
  assign \new_[7453]_  = ~\new_[8216]_  & ~\new_[8230]_ ;
  assign \new_[7454]_  = ~\new_[8602]_  | ~\new_[12172]_ ;
  assign \new_[7455]_  = ~\new_[8609]_  | ~\new_[8608]_  | ~\new_[8619]_ ;
  assign \new_[7456]_  = \new_[3461]_  ? \new_[11727]_  : \new_[8244]_ ;
  assign n7045 = \new_[10971]_  ^ \new_[8263]_ ;
  assign \new_[7458]_  = \new_[12302]_  ^ \new_[8277]_ ;
  assign n7030 = \new_[12406]_  ^ \new_[8264]_ ;
  assign \new_[7460]_  = \new_[12304]_  ^ \new_[8278]_ ;
  assign n7035 = \new_[11290]_  ^ \new_[8271]_ ;
  assign \new_[7462]_  = \new_[12285]_  ^ \new_[8279]_ ;
  assign n7040 = \new_[11999]_  ^ \new_[8274]_ ;
  assign \new_[7464]_  = \new_[12284]_  ^ \new_[8280]_ ;
  assign \new_[7465]_  = \new_[8226]_  & \new_[14529]_ ;
  assign \new_[7466]_  = ~\new_[9229]_  | ~\new_[13257]_  | ~\new_[9186]_  | ~\new_[11801]_ ;
  assign \new_[7467]_  = ~\new_[10828]_  | ~\new_[14635]_ ;
  assign \new_[7468]_  = (~\new_[10833]_  & ~\new_[14642]_ ) | (~\new_[10990]_  & ~\new_[8964]_ );
  assign \new_[7469]_  = ~\new_[7765]_ ;
  assign \new_[7470]_  = ~u1_u3_tx_data_to_reg;
  assign \new_[7471]_  = u1_u3_rx_ack_to_reg;
  assign \new_[7472]_  = ~\new_[8241]_  | ~\new_[2266]_ ;
  assign \new_[7473]_  = ~\new_[2266]_  | ~\new_[7861]_ ;
  assign \new_[7474]_  = ~\new_[2177]_  | ~\new_[8240]_ ;
  assign \new_[7475]_  = ~\new_[2136]_  | ~\new_[8240]_ ;
  assign \new_[7476]_  = ~\new_[7862]_  | ~\new_[2136]_ ;
  assign \new_[7477]_  = ~\new_[2178]_  | ~\new_[7861]_ ;
  assign \new_[7478]_  = ~\new_[7862]_  | ~\new_[2177]_ ;
  assign \new_[7479]_  = ~\new_[8241]_  | ~\new_[2178]_ ;
  assign \new_[7480]_  = ~\new_[7876]_  & ~\new_[12402]_ ;
  assign \new_[7481]_  = ~\new_[7780]_ ;
  assign \new_[7482]_  = ~\new_[7780]_ ;
  assign \new_[7483]_  = ~n6670;
  assign \new_[7484]_  = ~\new_[8238]_  | (~\new_[2991]_  & ~\new_[13386]_ );
  assign \new_[7485]_  = ~\new_[7789]_ ;
  assign \new_[7486]_  = ~\new_[7876]_  & (~\new_[11011]_  | ~\new_[9835]_ );
  assign \new_[7487]_  = (~\new_[9029]_  | ~\new_[6269]_ ) & (~\new_[8634]_  | ~\new_[14009]_ );
  assign \new_[7488]_  = (~\new_[9029]_  | ~\new_[4856]_ ) & (~\new_[8634]_  | ~\new_[5149]_ );
  assign \new_[7489]_  = (~\new_[9029]_  | ~\new_[4886]_ ) & (~\new_[8634]_  | ~\new_[5185]_ );
  assign \new_[7490]_  = (~\new_[9029]_  | ~\new_[4855]_ ) & (~\new_[8634]_  | ~\new_[5174]_ );
  assign \new_[7491]_  = (~\new_[9030]_  | ~\new_[6593]_ ) & (~\new_[8634]_  | ~\new_[6690]_ );
  assign \new_[7492]_  = ~\new_[7874]_  & (~\new_[11014]_  | ~\new_[9578]_ );
  assign \new_[7493]_  = (~\new_[9029]_  | ~\new_[14198]_ ) & (~\new_[8634]_  | ~\new_[13553]_ );
  assign \new_[7494]_  = (~\new_[9029]_  | ~\new_[14093]_ ) & (~\new_[8634]_  | ~\new_[14196]_ );
  assign \new_[7495]_  = (~\new_[9029]_  | ~\new_[13713]_ ) & (~\new_[8634]_  | ~\new_[14083]_ );
  assign \new_[7496]_  = (~\new_[9029]_  | ~\new_[14143]_ ) & (~\new_[8634]_  | ~\new_[14184]_ );
  assign \new_[7497]_  = (~\new_[9029]_  | ~\new_[6524]_ ) & (~\new_[8634]_  | ~\new_[13946]_ );
  assign \new_[7498]_  = (~\new_[9029]_  | ~\new_[13589]_ ) & (~\new_[8634]_  | ~\new_[13958]_ );
  assign \new_[7499]_  = (~\new_[9030]_  | ~\new_[13527]_ ) & (~\new_[8634]_  | ~\new_[13709]_ );
  assign \new_[7500]_  = (~\new_[9029]_  | ~\new_[13678]_ ) & (~\new_[8634]_  | ~\new_[13545]_ );
  assign \new_[7501]_  = (~\new_[9029]_  | ~\new_[14112]_ ) & (~\new_[8634]_  | ~\new_[13641]_ );
  assign \new_[7502]_  = (~\new_[9030]_  | ~\new_[13831]_ ) & (~\new_[8634]_  | ~\new_[13539]_ );
  assign \new_[7503]_  = (~\new_[9029]_  | ~\new_[13951]_ ) & (~\new_[8634]_  | ~\new_[13722]_ );
  assign \new_[7504]_  = (~\new_[9029]_  | ~\new_[13566]_ ) & (~\new_[8634]_  | ~\new_[13580]_ );
  assign \new_[7505]_  = (~\new_[9029]_  | ~\new_[6000]_ ) & (~\new_[8634]_  | ~\new_[13610]_ );
  assign \new_[7506]_  = (~\new_[9029]_  | ~\new_[14181]_ ) & (~\new_[8634]_  | ~\new_[13668]_ );
  assign \new_[7507]_  = (~\new_[9029]_  | ~\new_[14235]_ ) & (~\new_[8634]_  | ~\new_[13961]_ );
  assign \new_[7508]_  = (~\new_[9029]_  | ~\new_[13725]_ ) & (~\new_[8634]_  | ~\new_[14202]_ );
  assign \new_[7509]_  = (~\new_[9029]_  | ~\new_[13885]_ ) & (~\new_[8634]_  | ~\new_[13737]_ );
  assign \new_[7510]_  = (~\new_[9030]_  | ~\new_[6561]_ ) & (~\new_[8634]_  | ~\new_[6166]_ );
  assign \new_[7511]_  = (~\new_[9030]_  | ~\new_[6266]_ ) & (~\new_[8634]_  | ~\new_[6200]_ );
  assign \new_[7512]_  = (~\new_[9029]_  | ~\new_[14014]_ ) & (~\new_[8634]_  | ~\new_[13622]_ );
  assign \new_[7513]_  = (~\new_[9029]_  | ~\new_[14170]_ ) & (~\new_[8634]_  | ~\new_[13596]_ );
  assign \new_[7514]_  = (~\new_[9029]_  | ~\new_[13562]_ ) & (~\new_[8634]_  | ~\new_[13543]_ );
  assign \new_[7515]_  = (~\new_[9030]_  | ~\new_[14138]_ ) & (~\new_[8634]_  | ~\new_[13590]_ );
  assign \new_[7516]_  = (~\new_[9029]_  | ~\new_[14022]_ ) & (~\new_[8634]_  | ~\new_[13839]_ );
  assign \new_[7517]_  = (~\new_[9029]_  | ~\new_[13538]_ ) & (~\new_[8634]_  | ~\new_[13840]_ );
  assign \new_[7518]_  = (~\new_[9030]_  | ~\new_[14114]_ ) & (~\new_[8634]_  | ~\new_[13498]_ );
  assign \new_[7519]_  = (~\new_[9030]_  | ~\new_[14209]_ ) & (~\new_[8634]_  | ~\new_[14248]_ );
  assign \new_[7520]_  = (~\new_[9029]_  | ~\new_[13524]_ ) & (~\new_[8634]_  | ~\new_[14148]_ );
  assign \new_[7521]_  = (~\new_[9029]_  | ~\new_[13879]_ ) & (~\new_[8634]_  | ~\new_[13948]_ );
  assign \new_[7522]_  = (~\new_[9029]_  | ~\new_[14132]_ ) & (~\new_[8634]_  | ~\new_[13976]_ );
  assign \new_[7523]_  = (~\new_[9029]_  | ~\new_[13929]_ ) & (~\new_[8634]_  | ~\new_[13652]_ );
  assign \new_[7524]_  = (~\new_[9029]_  | ~\new_[13965]_ ) & (~\new_[8634]_  | ~\new_[14222]_ );
  assign \new_[7525]_  = (~\new_[9029]_  | ~\new_[14175]_ ) & (~\new_[8634]_  | ~\new_[13739]_ );
  assign \new_[7526]_  = (~\new_[9029]_  | ~\new_[13868]_ ) & (~\new_[8634]_  | ~\new_[13784]_ );
  assign \new_[7527]_  = (~\new_[9029]_  | ~\new_[13582]_ ) & (~\new_[8634]_  | ~\new_[14097]_ );
  assign \new_[7528]_  = (~\new_[9030]_  | ~\new_[6264]_ ) & (~\new_[8634]_  | ~\new_[6272]_ );
  assign \new_[7529]_  = ~\new_[8232]_  & (~\new_[9595]_  | ~\new_[9313]_ );
  assign n7065 = \new_[6696]_  ? n7635 : \new_[13166]_ ;
  assign n7085 = \new_[6716]_  ? n7635 : \new_[12846]_ ;
  assign n7090 = \new_[6718]_  ? n7635 : \new_[12783]_ ;
  assign n7170 = \new_[6736]_  ? n7635 : \new_[12870]_ ;
  assign n7175 = \new_[6737]_  ? n7635 : \new_[12651]_ ;
  assign n7180 = \new_[6738]_  ? n7635 : \new_[12816]_ ;
  assign n6925 = \new_[6604]_  ? n7635 : \new_[12916]_ ;
  assign n7185 = \new_[6739]_  ? n7635 : \new_[13192]_ ;
  assign \new_[7538]_  = ~\new_[9594]_  | ~\new_[10279]_  | ~\new_[8200]_  | ~\new_[10620]_ ;
  assign n7005 = ~\new_[8982]_  | ~\new_[8879]_  | ~\new_[9774]_  | ~\new_[8963]_ ;
  assign \new_[7540]_  = ~\new_[7845]_ ;
  assign \new_[7541]_  = ~\new_[8231]_  & (~\new_[8633]_  | ~\new_[5766]_ );
  assign \new_[7542]_  = ~\new_[12383]_  | ~\new_[7868]_ ;
  assign n6995 = ~\new_[8991]_  | ~\new_[8882]_  | ~\new_[9733]_  | ~\new_[8580]_ ;
  assign \new_[7544]_  = ~\new_[8229]_ ;
  assign \new_[7545]_  = ~\new_[7851]_ ;
  assign \new_[7546]_  = \new_[7866]_  & \new_[9611]_ ;
  assign n6975 = ~\new_[8985]_  | ~\new_[8864]_  | ~\new_[9778]_  | ~\new_[8612]_ ;
  assign \new_[7548]_  = ~\new_[7866]_  | ~\new_[6023]_ ;
  assign \new_[7549]_  = ~\new_[7854]_ ;
  assign \new_[7550]_  = \new_[7866]_  & \new_[13370]_ ;
  assign \new_[7551]_  = ~\new_[8233]_ ;
  assign \new_[7552]_  = ~\new_[7855]_ ;
  assign \new_[7553]_  = ~\new_[8638]_  | (~\new_[13267]_  & ~n8645);
  assign \new_[7554]_  = \new_[7866]_  & \new_[12838]_ ;
  assign \new_[7555]_  = ~\new_[7859]_ ;
  assign \new_[7556]_  = ~\new_[10468]_  | ~\new_[7866]_ ;
  assign \new_[7557]_  = ~\new_[7862]_ ;
  assign \new_[7558]_  = ~\new_[10469]_  | ~\new_[8247]_ ;
  assign \new_[7559]_  = ~\new_[7863]_ ;
  assign \new_[7560]_  = \new_[8247]_  & \new_[12838]_ ;
  assign \new_[7561]_  = ~\new_[8258]_  & (~\new_[12798]_  | ~n7590);
  assign \new_[7562]_  = ~\new_[8249]_  & (~\new_[9031]_  | ~\new_[13496]_ );
  assign \new_[7563]_  = ~\new_[8248]_  & (~\new_[9031]_  | ~\new_[13302]_ );
  assign \new_[7564]_  = ~\new_[8250]_  & (~\new_[9031]_  | ~\new_[6385]_ );
  assign \new_[7565]_  = ~\new_[8251]_  & (~\new_[9031]_  | ~\new_[6470]_ );
  assign \new_[7566]_  = ~\new_[8252]_  & (~\new_[9031]_  | ~\new_[6386]_ );
  assign \new_[7567]_  = ~\new_[8253]_  & (~\new_[9031]_  | ~\new_[6387]_ );
  assign \new_[7568]_  = ~\new_[8254]_  & (~\new_[9031]_  | ~\new_[6093]_ );
  assign \new_[7569]_  = ~\new_[8255]_  & (~\new_[9031]_  | ~\new_[6170]_ );
  assign \new_[7570]_  = ~\new_[8637]_  | (~\new_[8657]_  & ~\new_[12099]_ );
  assign n7550 = u1_u2_rx_data_done_r_reg;
  assign \new_[7572]_  = ~\\u4_utmi_vend_ctrl_r_reg[2] ;
  assign \new_[7573]_  = ~\new_[8652]_  | ~\new_[8269]_ ;
  assign \new_[7574]_  = ~\new_[8289]_  | (~\new_[10447]_  & ~\new_[9633]_ );
  assign \new_[7575]_  = ~\new_[8290]_  | (~\new_[10446]_  & ~\new_[9634]_ );
  assign \new_[7576]_  = ~\new_[11852]_  | (~\new_[8922]_  & ~\new_[12014]_ );
  assign \new_[7577]_  = ~\new_[11846]_  | (~\new_[8662]_  & ~\new_[12472]_ );
  assign \new_[7578]_  = ~\new_[11867]_  | (~\new_[8918]_  & ~\new_[12307]_ );
  assign \new_[7579]_  = ~\new_[11869]_  | (~\new_[8663]_  & ~\new_[12328]_ );
  assign \new_[7580]_  = ~\new_[10342]_  | ~\new_[11485]_  | ~\new_[8684]_ ;
  assign \new_[7581]_  = ~\new_[11092]_  | ~\new_[11508]_  | ~\new_[8294]_  | ~\new_[11795]_ ;
  assign \new_[7582]_  = ~\new_[9060]_  | ~\new_[9616]_  | ~\new_[12441]_  | ~\new_[8672]_ ;
  assign \new_[7583]_  = ~\new_[11091]_  | ~\new_[11500]_  | ~\new_[8295]_  | ~\new_[12094]_ ;
  assign \new_[7584]_  = ~\new_[11094]_  | ~\new_[11494]_  | ~\new_[8296]_  | ~\new_[11493]_ ;
  assign \new_[7585]_  = ~\new_[10345]_  | ~\new_[11629]_  | ~\new_[8685]_ ;
  assign \new_[7586]_  = ~\new_[8562]_  & (~\new_[11599]_  | ~\new_[9363]_ );
  assign \new_[7587]_  = ~\new_[9057]_  | ~\new_[9618]_  | ~\new_[12375]_  | ~\new_[8651]_ ;
  assign \new_[7588]_  = ~\new_[10348]_  | ~\new_[11619]_  | ~\new_[8686]_ ;
  assign \new_[7589]_  = ~\new_[9062]_  | ~\new_[9621]_  | ~\new_[12371]_  | ~\new_[8699]_ ;
  assign \new_[7590]_  = ~\new_[10005]_  | ~\new_[11638]_  | ~\new_[8687]_ ;
  assign \new_[7591]_  = ~\new_[9064]_  | ~\new_[9623]_  | ~\new_[12430]_  | ~\new_[8671]_ ;
  assign \new_[7592]_  = ~\new_[13609]_  | ~\new_[8527]_  | ~\new_[13091]_ ;
  assign \new_[7593]_  = \new_[9367]_  | \new_[8299]_ ;
  assign \new_[7594]_  = \new_[9368]_  | \new_[8298]_ ;
  assign \new_[7595]_  = \new_[9369]_  | \new_[8300]_ ;
  assign \new_[7596]_  = \new_[9370]_  | \new_[8301]_ ;
  assign n7490 = \new_[12347]_  ^ \new_[8690]_ ;
  assign n7495 = \new_[12478]_  ^ \new_[8694]_ ;
  assign \new_[7599]_  = ~\new_[13668]_  | ~\new_[8525]_  | ~\new_[13098]_ ;
  assign \new_[7600]_  = ~\new_[14181]_  | ~\new_[8473]_  | ~\new_[13149]_ ;
  assign \new_[7601]_  = ~\new_[8292]_  | ~\new_[3787]_ ;
  assign \new_[7602]_  = ~\new_[8291]_  | ~\new_[3940]_ ;
  assign \new_[7603]_  = ~\new_[8291]_  | ~\new_[8719]_ ;
  assign \new_[7604]_  = \\u4_u1_dma_out_left_reg[7] ;
  assign \new_[7605]_  = ~\new_[8307]_  | (~\new_[10864]_  & ~\new_[9671]_ );
  assign \new_[7606]_  = ~\new_[8311]_  | (~\new_[10797]_  & ~\new_[9677]_ );
  assign n7500 = ~\new_[12505]_  & (~\new_[8761]_  | ~\new_[8762]_ );
  assign n7370 = ~\new_[12505]_  & (~\new_[8798]_  | ~\new_[8763]_ );
  assign n7530 = ~\new_[12732]_  & (~\new_[8766]_  | ~\new_[8765]_ );
  assign n7375 = ~\new_[12245]_  & (~\new_[8767]_  | ~\new_[8802]_ );
  assign n7535 = ~\new_[12732]_  & (~\new_[8768]_  | ~\new_[8796]_ );
  assign n7380 = ~\new_[12505]_  & (~\new_[8793]_  | ~\new_[8769]_ );
  assign n7385 = ~\new_[12849]_  & (~\new_[8770]_  | ~\new_[8789]_ );
  assign n7390 = ~\new_[12732]_  & (~\new_[8782]_  | ~\new_[8781]_ );
  assign n7525 = ~\new_[12732]_  & (~\new_[8771]_  | ~\new_[8843]_ );
  assign n7400 = ~\new_[12245]_  & (~\new_[8804]_  | ~\new_[8772]_ );
  assign n7395 = ~\new_[12505]_  & (~\new_[8773]_  | ~\new_[8760]_ );
  assign n7515 = ~\new_[12732]_  & (~\new_[8774]_  | ~\new_[8784]_ );
  assign \new_[7619]_  = (~\new_[9055]_  | ~\new_[3693]_ ) & (~\new_[8858]_  | ~\new_[3690]_ );
  assign \new_[7620]_  = (~\new_[8691]_  | ~\new_[3316]_ ) & (~\new_[8856]_  | ~\new_[3315]_ );
  assign \new_[7621]_  = ~\new_[8262]_  | ~\new_[3940]_ ;
  assign \new_[7622]_  = \new_[8299]_  | \new_[6253]_ ;
  assign \new_[7623]_  = ~\new_[8299]_  & ~\new_[6196]_ ;
  assign n7405 = ~\new_[12505]_  & (~\new_[8725]_  | ~\new_[8776]_ );
  assign n7315 = ~\new_[12732]_  & (~\new_[8759]_  | ~\new_[8785]_ );
  assign n7410 = ~\new_[12732]_  & (~\new_[8726]_  | ~\new_[8823]_ );
  assign n7240 = ~\new_[12732]_  & (~\new_[8727]_  | ~\new_[8828]_ );
  assign n7265 = ~\new_[12849]_  & (~\new_[8748]_  | ~\new_[8831]_ );
  assign n7280 = ~\new_[12732]_  & (~\new_[8732]_  | ~\new_[8786]_ );
  assign n7285 = ~\new_[12732]_  & (~\new_[8733]_  | ~\new_[8800]_ );
  assign n7250 = ~\new_[12849]_  & (~\new_[8724]_  | ~\new_[8787]_ );
  assign n7270 = ~\new_[12732]_  & (~\new_[8747]_  | ~\new_[8788]_ );
  assign n7275 = ~\new_[12849]_  & (~\new_[8728]_  | ~\new_[8799]_ );
  assign n7255 = ~\new_[12732]_  & (~\new_[8729]_  | ~\new_[8777]_ );
  assign n7235 = ~\new_[12732]_  & (~\new_[8730]_  | ~\new_[8825]_ );
  assign \new_[7636]_  = ~\new_[8790]_  | ~\new_[9208]_  | ~\new_[10032]_ ;
  assign \new_[7637]_  = ~\new_[8301]_  & ~\new_[6287]_ ;
  assign \new_[7638]_  = ~\new_[8284]_  | ~\new_[3310]_ ;
  assign \new_[7639]_  = \new_[8298]_  | \new_[6266]_ ;
  assign \new_[7640]_  = ~\new_[8298]_  & ~\new_[6567]_ ;
  assign n7520 = ~\new_[12849]_  & (~\new_[8811]_  | ~\new_[8735]_ );
  assign n7415 = ~\new_[12849]_  & (~\new_[8812]_  | ~\new_[8736]_ );
  assign n7420 = ~\new_[12849]_  & (~\new_[8813]_  | ~\new_[8737]_ );
  assign n7425 = ~\new_[12849]_  & (~\new_[8814]_  | ~\new_[8738]_ );
  assign n7480 = ~\new_[12849]_  & (~\new_[8815]_  | ~\new_[8739]_ );
  assign n7430 = ~\new_[12245]_  & (~\new_[8816]_  | ~\new_[8740]_ );
  assign n7485 = ~\new_[12732]_  & (~\new_[8817]_  | ~\new_[8741]_ );
  assign n7435 = ~\new_[12732]_  & (~\new_[8818]_  | ~\new_[8742]_ );
  assign n7475 = ~\new_[12732]_  & (~\new_[8819]_  | ~\new_[8743]_ );
  assign n7445 = ~\new_[12732]_  & (~\new_[8808]_  | ~\new_[8744]_ );
  assign n7440 = ~\new_[12732]_  & (~\new_[8820]_  | ~\new_[8745]_ );
  assign n7465 = ~\new_[12849]_  & (~\new_[8806]_  | ~\new_[8746]_ );
  assign \new_[7653]_  = ~\\u4_u1_buf0_orig_m3_reg[11] ;
  assign \new_[7654]_  = ~\new_[8308]_  & ~\new_[2741]_ ;
  assign \new_[7655]_  = \new_[8300]_  | \new_[6200]_ ;
  assign \new_[7656]_  = ~\new_[8300]_  & ~\new_[6275]_ ;
  assign n7295 = ~\new_[12732]_  & (~\new_[8750]_  | ~\new_[8832]_ );
  assign n7310 = ~\new_[12732]_  & (~\new_[8751]_  | ~\new_[8833]_ );
  assign n7450 = ~\new_[12849]_  & (~\new_[8752]_  | ~\new_[8783]_ );
  assign n7320 = ~\new_[12732]_  & (~\new_[8753]_  | ~\new_[8834]_ );
  assign n7245 = ~\new_[12505]_  & (~\new_[8754]_  | ~\new_[8835]_ );
  assign n7260 = ~\new_[12505]_  & (~\new_[8722]_  | ~\new_[8836]_ );
  assign n7470 = ~\new_[12732]_  & (~\new_[8755]_  | ~\new_[8778]_ );
  assign n7510 = ~\new_[12732]_  & (~\new_[8723]_  | ~\new_[8837]_ );
  assign n7540 = ~\new_[12732]_  & (~\new_[8721]_  | ~\new_[8838]_ );
  assign n7555 = ~\new_[12732]_  & (~\new_[8756]_  | ~\new_[8839]_ );
  assign n7455 = ~\new_[12849]_  & (~\new_[8757]_  | ~\new_[8824]_ );
  assign n7560 = ~\new_[12732]_  & (~\new_[8758]_  | ~\new_[8840]_ );
  assign \new_[7669]_  = ~\new_[8606]_  | ~\new_[8366]_ ;
  assign \new_[7670]_  = \\u1_u1_state_reg[2] ;
  assign \new_[7671]_  = \new_[8301]_  | \new_[6009]_ ;
  assign \new_[7672]_  = ~\new_[8597]_  | ~\new_[8395]_ ;
  assign \new_[7673]_  = ~\\u4_utmi_vend_ctrl_r_reg[1] ;
  assign \new_[7674]_  = ~\new_[8304]_  & (~\new_[11156]_  | ~\new_[10716]_ );
  assign \new_[7675]_  = ~\new_[8305]_  & (~\new_[11165]_  | ~\new_[11013]_ );
  assign \new_[7676]_  = ~\new_[8309]_  & (~\new_[11180]_  | ~\new_[10717]_ );
  assign \new_[7677]_  = ~\new_[8313]_  & (~\new_[11177]_  | ~\new_[10355]_ );
  assign \new_[7678]_  = ~\new_[8303]_  & (~\new_[13469]_  | ~n8645);
  assign n7305 = (~\new_[11917]_  & ~\new_[8780]_ ) | (~\new_[12231]_  & ~\new_[9426]_ );
  assign \new_[7680]_  = ~\new_[8287]_  | ~\new_[8398]_ ;
  assign n7300 = (~\new_[11880]_  & ~\new_[8803]_ ) | (~\new_[8880]_  & ~\new_[12231]_ );
  assign n7345 = (~\new_[11907]_  & ~\new_[8829]_ ) | (~\new_[9430]_  & ~\new_[12231]_ );
  assign n7565 = (~\new_[12274]_  & ~\new_[8830]_ ) | (~\new_[9445]_  & ~\new_[12231]_ );
  assign \new_[7684]_  = \new_[4289]_  ^ \new_[8847]_ ;
  assign \new_[7685]_  = \new_[3477]_  ^ \new_[8848]_ ;
  assign \new_[7686]_  = \new_[3688]_  ^ \new_[8849]_ ;
  assign \new_[7687]_  = \new_[3883]_  ^ \new_[8850]_ ;
  assign \new_[7688]_  = ~\new_[7908]_ ;
  assign \new_[7689]_  = ~\new_[9059]_  | (~\new_[8717]_  & ~\new_[3283]_ );
  assign \new_[7690]_  = ~\new_[7910]_ ;
  assign \new_[7691]_  = ~\new_[8314]_  | (~\new_[8718]_  & ~\new_[3309]_ );
  assign \new_[7692]_  = ~\new_[8306]_  | ~\new_[9126]_ ;
  assign \new_[7693]_  = \new_[3940]_  ^ \new_[8890]_ ;
  assign \new_[7694]_  = \new_[3310]_  ^ \new_[8904]_ ;
  assign \new_[7695]_  = \new_[3464]_  ^ \new_[8906]_ ;
  assign \new_[7696]_  = \new_[3787]_  ^ \new_[8912]_ ;
  assign n7350 = ~\new_[12842]_  & (~\new_[8807]_  | ~\new_[10347]_ );
  assign \new_[7698]_  = (~\new_[8791]_  | ~\wb_data_i[0] ) & (~\new_[9087]_  | ~\new_[6239]_ );
  assign \new_[7699]_  = (~\new_[8791]_  | ~\wb_data_i[1] ) & (~\new_[9087]_  | ~\new_[6240]_ );
  assign \new_[7700]_  = (~\new_[8791]_  | ~\wb_data_i[2] ) & (~\new_[9087]_  | ~\new_[6241]_ );
  assign \new_[7701]_  = (~\new_[8791]_  | ~\wb_data_i[3] ) & (~\new_[9087]_  | ~\new_[6107]_ );
  assign \new_[7702]_  = (~\new_[8791]_  | ~\wb_data_i[4] ) & (~\new_[9087]_  | ~\new_[6242]_ );
  assign \new_[7703]_  = (~\new_[8791]_  | ~\wb_data_i[5] ) & (~\new_[9087]_  | ~\new_[6105]_ );
  assign \new_[7704]_  = (~\new_[8791]_  | ~\wb_data_i[6] ) & (~\new_[9087]_  | ~\new_[6243]_ );
  assign \new_[7705]_  = ~u4_int_src_re_reg;
  assign \new_[7706]_  = ~\new_[13327]_  | ~\new_[13858]_  | ~\new_[8577]_  | ~\new_[2961]_ ;
  assign n7335 = ~\new_[8992]_  | ~\new_[8615]_  | ~\new_[8899]_ ;
  assign n7330 = ~\new_[9013]_  | ~\new_[8944]_  | ~\new_[8905]_ ;
  assign n7325 = ~\new_[8903]_  | ~\new_[8590]_  | ~\new_[9015]_ ;
  assign \new_[7710]_  = ~\new_[8322]_  & ~\new_[13326]_ ;
  assign n7340 = ~\new_[8868]_  | ~\new_[8607]_  | ~\new_[9007]_ ;
  assign \new_[7712]_  = ~\new_[8821]_  & ~\new_[8261]_ ;
  assign n7290 = ~\new_[8416]_  | ~\new_[8417]_ ;
  assign \new_[7714]_  = ~\new_[6011]_  & (~\new_[8914]_  | ~\new_[8633]_ );
  assign \new_[7715]_  = ~\new_[6310]_  & (~\new_[8914]_  | ~\new_[8970]_ );
  assign \new_[7716]_  = ~\new_[9957]_  & (~\new_[8844]_  | ~\new_[10028]_ );
  assign \new_[7717]_  = ~\new_[13902]_  | ~\new_[8453]_  | ~\new_[13151]_ ;
  assign \new_[7718]_  = ~\\u4_utmi_vend_ctrl_r_reg[0] ;
  assign \new_[7719]_  = ~\new_[5993]_  | ~\new_[8523]_  | ~\new_[10720]_ ;
  assign \new_[7720]_  = ~\new_[13350]_  | ~\new_[8598]_  | ~\new_[8666]_ ;
  assign n7505 = ~\new_[10067]_  & (~\new_[8898]_  | ~\new_[10425]_ );
  assign \new_[7722]_  = ~\new_[7944]_ ;
  assign \new_[7723]_  = ~\new_[7948]_ ;
  assign \new_[7724]_  = ~\new_[8577]_  | ~TermSel_pad_o;
  assign \new_[7725]_  = ~\new_[9145]_  | ~\wb_data_i[6] ;
  assign \new_[7726]_  = ~\new_[9047]_  | ~\wb_data_i[2] ;
  assign \new_[7727]_  = ~\new_[9047]_  | ~\wb_data_i[4] ;
  assign \new_[7728]_  = ~\new_[9047]_  | ~\wb_data_i[16] ;
  assign \new_[7729]_  = ~\new_[9047]_  | ~\wb_data_i[17] ;
  assign \new_[7730]_  = ~\new_[9047]_  | ~\wb_data_i[18] ;
  assign \new_[7731]_  = ~\new_[8476]_  & (~\new_[14636]_  | ~\new_[2349]_ );
  assign \new_[7732]_  = ~\new_[9145]_  | ~\wb_data_i[0] ;
  assign \new_[7733]_  = ~\new_[9138]_  | ~\new_[6012]_ ;
  assign \new_[7734]_  = ~\new_[8792]_  & (~\new_[8664]_  | ~\new_[3888]_ );
  assign \new_[7735]_  = (~\new_[10106]_  | ~\new_[9846]_ ) & (~\new_[9106]_  | ~\new_[10572]_ );
  assign \new_[7736]_  = ~\new_[8604]_  & ~\new_[9218]_ ;
  assign \new_[7737]_  = ~\new_[9095]_  & (~\new_[8665]_  | ~\new_[4293]_ );
  assign \new_[7738]_  = ~\new_[9145]_  | ~\wb_data_i[2] ;
  assign \new_[7739]_  = ~\new_[9145]_  | ~\wb_data_i[9] ;
  assign \new_[7740]_  = ~\new_[8599]_  | ~\new_[4798]_ ;
  assign \new_[7741]_  = ~\new_[8601]_  & ~\new_[2875]_ ;
  assign \new_[7742]_  = \new_[8600]_  | \new_[2857]_ ;
  assign \new_[7743]_  = \new_[8603]_  | \new_[2876]_ ;
  assign \new_[7744]_  = \new_[8602]_  | \new_[2503]_ ;
  assign \new_[7745]_  = ~\new_[8601]_  | ~\new_[13919]_ ;
  assign \new_[7746]_  = ~\new_[8599]_  & ~\new_[4798]_ ;
  assign \new_[7747]_  = \new_[8688]_  ? \new_[14636]_  : \new_[2317]_ ;
  assign n7355 = ~\new_[8645]_  | ~\new_[8949]_  | ~\new_[8934]_ ;
  assign n7360 = ~\new_[8983]_  | ~\new_[8958]_  | ~\new_[8935]_ ;
  assign \new_[7750]_  = \new_[10484]_  & \new_[8577]_ ;
  assign n7365 = ~\new_[9006]_  | ~\new_[8948]_  | ~\new_[8933]_ ;
  assign \new_[7752]_  = ~\new_[8564]_  & ~\new_[13561]_ ;
  assign \new_[7753]_  = ~\new_[8564]_  & ~\new_[14115]_ ;
  assign \new_[7754]_  = ~\new_[14636]_  & ~\new_[8595]_ ;
  assign \new_[7755]_  = ~\new_[8288]_  & ~\new_[14636]_ ;
  assign \new_[7756]_  = ~\new_[9048]_  | ~\wb_data_i[2] ;
  assign \new_[7757]_  = ~\new_[8575]_  & ~\new_[13461]_ ;
  assign \new_[7758]_  = ~\new_[8574]_  & ~\new_[13324]_ ;
  assign \new_[7759]_  = ~\new_[9048]_  | ~\wb_data_i[5] ;
  assign \new_[7760]_  = ~\new_[9048]_  | ~\wb_data_i[9] ;
  assign \new_[7761]_  = ~\new_[9048]_  | ~\wb_data_i[25] ;
  assign \new_[7762]_  = ~\new_[8583]_  & (~\new_[9476]_  | ~\new_[10097]_ );
  assign \new_[7763]_  = ~\\u4_utmi_vend_ctrl_r_reg[3] ;
  assign \new_[7764]_  = ~\new_[11000]_  & (~\new_[8629]_  | ~\new_[9605]_ );
  assign \new_[7765]_  = (~\new_[8932]_  | ~\new_[10371]_ ) & (~\new_[8931]_  | ~\new_[9800]_ );
  assign \new_[7766]_  = ~\new_[8594]_  & (~\new_[10496]_  | ~\new_[12606]_ );
  assign n7460 = \new_[9303]_  | \new_[8984]_  | \new_[9009]_  | \new_[9011]_ ;
  assign \new_[7768]_  = ~\new_[5762]_  | ~\new_[8242]_ ;
  assign \new_[7769]_  = ~\new_[8242]_  | ~\new_[5763]_ ;
  assign \new_[7770]_  = ~\new_[8627]_  | ~\new_[5860]_ ;
  assign \new_[7771]_  = ~\new_[8614]_  | ~\new_[9850]_ ;
  assign \new_[7772]_  = ~\new_[8614]_  & ~\new_[10277]_ ;
  assign \new_[7773]_  = ~\new_[9574]_  | ~\new_[8614]_ ;
  assign \new_[7774]_  = ~\new_[5764]_  | ~\new_[8627]_ ;
  assign \new_[7775]_  = \new_[8272]_  & \new_[12350]_ ;
  assign \new_[7776]_  = \new_[8246]_  | \new_[9275]_ ;
  assign \new_[7777]_  = ~\new_[11698]_  & (~\new_[8641]_  | ~\new_[11430]_ );
  assign \new_[7778]_  = ~\new_[11698]_  & (~\new_[8641]_  | ~\new_[10452]_ );
  assign \new_[7779]_  = ~\new_[9229]_  | ~\new_[9190]_  | ~\new_[11430]_ ;
  assign \new_[7780]_  = ~\new_[8214]_ ;
  assign \new_[7781]_  = \new_[8215]_ ;
  assign \new_[7782]_  = \new_[8215]_ ;
  assign \new_[7783]_  = \new_[8215]_ ;
  assign n6670 = ~\new_[8215]_ ;
  assign \new_[7785]_  = ~\new_[13456]_  | ~\new_[8623]_  | ~\new_[13450]_ ;
  assign \new_[7786]_  = (~\new_[8654]_  & ~\new_[12099]_ ) | (~\new_[8649]_  & ~\new_[12125]_ );
  assign \new_[7787]_  = ~\new_[4791]_  | ~\new_[12416]_  | ~\new_[8243]_  | ~\new_[13293]_ ;
  assign \new_[7788]_  = ~\new_[13135]_  | ~\new_[8625]_  | ~\new_[2673]_ ;
  assign \new_[7789]_  = ~\new_[14346]_  & (~\new_[9528]_  | ~\new_[9229]_ );
  assign \new_[7790]_  = (~\new_[9029]_  | ~\new_[6267]_ ) & (~\new_[8634]_  | ~\new_[6276]_ );
  assign \new_[7791]_  = (~\new_[9029]_  | ~\new_[13853]_ ) & (~\new_[8634]_  | ~\new_[14113]_ );
  assign \new_[7792]_  = (~n7650 | ~\new_[13615]_ ) & (~\new_[8634]_  | ~\new_[13741]_ );
  assign \new_[7793]_  = (~\new_[9029]_  | ~\new_[6539]_ ) & (~\new_[8634]_  | ~\new_[6172]_ );
  assign \new_[7794]_  = (~\new_[9029]_  | ~\new_[6543]_ ) & (~\new_[8634]_  | ~\new_[6277]_ );
  assign \new_[7795]_  = (~\new_[9029]_  | ~\new_[4854]_ ) & (~\new_[8634]_  | ~\new_[5148]_ );
  assign \new_[7796]_  = (~\new_[9029]_  | ~\new_[5999]_ ) & (~\new_[8634]_  | ~\new_[6274]_ );
  assign \new_[7797]_  = (~\new_[9029]_  | ~\new_[6557]_ ) & (~\new_[8634]_  | ~\new_[6005]_ );
  assign \new_[7798]_  = (~n7650 | ~\new_[13979]_ ) & (~\new_[8634]_  | ~\new_[13786]_ );
  assign \new_[7799]_  = (~n7650 | ~\new_[13669]_ ) & (~\new_[8634]_  | ~\new_[13726]_ );
  assign \new_[7800]_  = (~\new_[9029]_  | ~\new_[13762]_ ) & (~\new_[8634]_  | ~\new_[13983]_ );
  assign \new_[7801]_  = (~\new_[9030]_  | ~\new_[13871]_ ) & (~\new_[8634]_  | ~\new_[14165]_ );
  assign \new_[7802]_  = (~\new_[9030]_  | ~\new_[6599]_ ) & (~\new_[8634]_  | ~\new_[6237]_ );
  assign \new_[7803]_  = (~\new_[9029]_  | ~\new_[13846]_ ) & (~\new_[8634]_  | ~\new_[13632]_ );
  assign \new_[7804]_  = (~n7650 | ~\new_[13935]_ ) & (~\new_[8634]_  | ~\new_[14255]_ );
  assign \new_[7805]_  = (~\new_[9030]_  | ~\new_[14249]_ ) & (~\new_[8634]_  | ~\new_[13806]_ );
  assign \new_[7806]_  = (~\new_[9030]_  | ~\new_[6567]_ ) & (~\new_[8634]_  | ~\new_[6275]_ );
  assign \new_[7807]_  = (~\new_[9029]_  | ~\new_[6563]_ ) & (~\new_[8634]_  | ~\new_[6004]_ );
  assign \new_[7808]_  = (~\new_[9029]_  | ~\new_[5998]_ ) & (~\new_[8634]_  | ~\new_[6003]_ );
  assign \new_[7809]_  = (~n7650 | ~\new_[6001]_ ) & (~\new_[8634]_  | ~\new_[14172]_ );
  assign \new_[7810]_  = (~\new_[9620]_  | ~\new_[13934]_ ) & (~\new_[8634]_  | ~\new_[13707]_ );
  assign \new_[7811]_  = (~\new_[9029]_  | ~\new_[13685]_ ) & (~\new_[8634]_  | ~\new_[14140]_ );
  assign \new_[7812]_  = (~\new_[9029]_  | ~\new_[13890]_ ) & (~\new_[8634]_  | ~\new_[14024]_ );
  assign \new_[7813]_  = (~\new_[9029]_  | ~\new_[14075]_ ) & (~\new_[8634]_  | ~\new_[13859]_ );
  assign \new_[7814]_  = (~n7650 | ~\new_[13701]_ ) & (~\new_[8634]_  | ~\new_[13955]_ );
  assign \new_[7815]_  = (~n7650 | ~\new_[14166]_ ) & (~\new_[8634]_  | ~\new_[14173]_ );
  assign \new_[7816]_  = (~\new_[9029]_  | ~\new_[14158]_ ) & (~\new_[8634]_  | ~\new_[14117]_ );
  assign \new_[7817]_  = (~\new_[9029]_  | ~\new_[13651]_ ) & (~\new_[8634]_  | ~\new_[14085]_ );
  assign \new_[7818]_  = (~\new_[9029]_  | ~\new_[13529]_ ) & (~\new_[8634]_  | ~\new_[13687]_ );
  assign \new_[7819]_  = (~n7650 | ~\new_[13838]_ ) & (~\new_[8634]_  | ~\new_[14137]_ );
  assign \new_[7820]_  = (~n7650 | ~\new_[14068]_ ) & (~\new_[8634]_  | ~\new_[13536]_ );
  assign \new_[7821]_  = (~\new_[9029]_  | ~\new_[13830]_ ) & (~\new_[8634]_  | ~\new_[13557]_ );
  assign \new_[7822]_  = (~\new_[9029]_  | ~\new_[13775]_ ) & (~\new_[8634]_  | ~\new_[13887]_ );
  assign \new_[7823]_  = (~\new_[9620]_  | ~\new_[13603]_ ) & (~\new_[8634]_  | ~\new_[13619]_ );
  assign \new_[7824]_  = ~\new_[9415]_  | ~\new_[2042]_  | ~\new_[8261]_  | ~\new_[2452]_ ;
  assign \new_[7825]_  = (~\new_[9030]_  | ~\new_[14182]_ ) & (~\new_[8634]_  | ~\new_[14206]_ );
  assign \new_[7826]_  = ~\new_[8265]_  & (~\new_[10744]_  | ~\new_[12359]_ );
  assign \new_[7827]_  = ~\new_[8270]_  & (~\new_[10743]_  | ~\new_[12612]_ );
  assign \new_[7828]_  = (~n7650 | ~\new_[13909]_ ) & (~\new_[8634]_  | ~\new_[13982]_ );
  assign \new_[7829]_  = (~n7650 | ~\new_[13767]_ ) & (~\new_[8634]_  | ~\new_[14212]_ );
  assign \new_[7830]_  = (~\new_[9029]_  | ~\new_[13671]_ ) & (~\new_[8634]_  | ~\new_[13792]_ );
  assign \new_[7831]_  = ~\new_[8273]_  & (~\new_[10411]_  | ~\new_[12294]_ );
  assign \new_[7832]_  = ~\new_[8276]_  & (~\new_[10413]_  | ~\new_[12272]_ );
  assign \new_[7833]_  = (~\new_[9029]_  | ~\new_[13998]_ ) & (~\new_[8634]_  | ~\new_[14092]_ );
  assign \new_[7834]_  = (~n7650 | ~\new_[13773]_ ) & (~\new_[8634]_  | ~\new_[14062]_ );
  assign \new_[7835]_  = (~\new_[9029]_  | ~\new_[14183]_ ) & (~\new_[8634]_  | ~\new_[14154]_ );
  assign \new_[7836]_  = (~\new_[9029]_  | ~\new_[13869]_ ) & (~\new_[8634]_  | ~\new_[14178]_ );
  assign \new_[7837]_  = (~\new_[9029]_  | ~\new_[14065]_ ) & (~\new_[8634]_  | ~\new_[13854]_ );
  assign \new_[7838]_  = (~n7650 | ~\new_[14122]_ ) & (~\new_[8634]_  | ~\new_[14220]_ );
  assign \new_[7839]_  = (~n7650 | ~\new_[13991]_ ) & (~\new_[8634]_  | ~\new_[14145]_ );
  assign \new_[7840]_  = (~\new_[9030]_  | ~\new_[14168]_ ) & (~\new_[8634]_  | ~\new_[13683]_ );
  assign \new_[7841]_  = (~\new_[9030]_  | ~\new_[13500]_ ) & (~\new_[8634]_  | ~\new_[13764]_ );
  assign \new_[7842]_  = (~\new_[9030]_  | ~\new_[14123]_ ) & (~\new_[8634]_  | ~\new_[13807]_ );
  assign \new_[7843]_  = (~n7650 | ~\new_[13894]_ ) & (~\new_[8634]_  | ~\new_[14192]_ );
  assign \new_[7844]_  = ~\new_[8559]_  | ~\new_[8618]_ ;
  assign \new_[7845]_  = \new_[8222]_ ;
  assign \new_[7846]_  = ~\new_[8223]_ ;
  assign \new_[7847]_  = ~\new_[9161]_  | ~\new_[11434]_  | ~\new_[11086]_  | ~\new_[11752]_ ;
  assign \new_[7848]_  = ~\new_[14539]_ ;
  assign \new_[7849]_  = u1_u0_token_valid_r1_reg;
  assign \new_[7850]_  = ~\new_[8268]_  | ~\new_[9576]_ ;
  assign \new_[7851]_  = ~\new_[8609]_ ;
  assign \new_[7852]_  = ~\new_[8231]_ ;
  assign \new_[7853]_  = ~u4_utmi_vend_wr_r_reg;
  assign \new_[7854]_  = \new_[8247]_  & \new_[9611]_ ;
  assign \new_[7855]_  = \new_[8247]_  & \new_[13370]_ ;
  assign \new_[7856]_  = \\u1_u1_state_reg[3] ;
  assign \new_[7857]_  = ~\new_[8237]_ ;
  assign \new_[7858]_  = ~\new_[8247]_  | ~\new_[6023]_ ;
  assign \new_[7859]_  = \new_[8247]_  & \new_[12812]_ ;
  assign \new_[7860]_  = ~\new_[8241]_ ;
  assign \new_[7861]_  = ~\new_[8242]_ ;
  assign \new_[7862]_  = \new_[8633]_  & \new_[12812]_ ;
  assign \new_[7863]_  = ~\new_[9232]_  & (~\new_[10495]_  | ~\new_[10282]_ );
  assign \new_[7864]_  = ~\new_[10466]_  | ~\new_[8633]_ ;
  assign \new_[7865]_  = ~\new_[8640]_  & (~\new_[11006]_  | ~\new_[10096]_ );
  assign \new_[7866]_  = u4_u0_ep_match_r_reg;
  assign \new_[7867]_  = ~\new_[14245]_  | ~\new_[9375]_ ;
  assign \new_[7868]_  = \new_[12125]_  | \new_[9352]_ ;
  assign \new_[7869]_  = ~\new_[8261]_ ;
  assign \new_[7870]_  = ~\new_[9472]_  | ~\new_[11869]_  | ~\new_[10352]_  | ~\new_[13299]_ ;
  assign \new_[7871]_  = ~\new_[9220]_  | (~\new_[9046]_  & ~\new_[9857]_ );
  assign \new_[7872]_  = ~\new_[8268]_ ;
  assign \new_[7873]_  = ~\new_[8667]_  | (~\new_[9782]_  & ~\new_[11621]_ );
  assign \new_[7874]_  = ~\new_[8272]_ ;
  assign \new_[7875]_  = ~\new_[8282]_ ;
  assign \new_[7876]_  = ~\new_[13117]_  | ~\new_[10483]_  | ~\new_[9066]_ ;
  assign \new_[7877]_  = ~\new_[9206]_  | ~\new_[11133]_  | ~\new_[10369]_  | ~\new_[11142]_ ;
  assign \new_[7878]_  = ~\new_[9483]_  | ~\new_[11867]_  | ~\new_[10012]_  | ~\new_[13379]_ ;
  assign \new_[7879]_  = ~\new_[8287]_ ;
  assign \new_[7880]_  = \\u4_u3_dma_out_left_reg[7] ;
  assign \new_[7881]_  = \\u4_u0_dma_out_left_reg[7] ;
  assign \new_[7882]_  = \\u4_u2_dma_out_left_reg[7] ;
  assign \new_[7883]_  = ~\new_[8859]_  & ~\new_[12836]_ ;
  assign \new_[7884]_  = ~\new_[8928]_  & ~\new_[12336]_ ;
  assign \new_[7885]_  = ~\new_[8695]_  | (~\new_[11135]_  & ~\new_[10408]_ );
  assign \new_[7886]_  = ~\new_[8698]_  | (~\new_[11137]_  & ~\new_[10410]_ );
  assign \new_[7887]_  = ~\new_[8696]_  | (~\new_[11154]_  & ~\new_[10409]_ );
  assign \new_[7888]_  = ~\new_[8697]_  | (~\new_[11136]_  & ~\new_[10406]_ );
  assign \new_[7889]_  = \new_[8684]_  | \new_[12673]_ ;
  assign \new_[7890]_  = \new_[8684]_  | \new_[12272]_ ;
  assign \new_[7891]_  = (~\new_[9054]_  | ~\new_[4073]_ ) & (~\new_[9419]_  | ~\new_[4070]_ );
  assign \new_[7892]_  = ~\new_[8672]_  & ~\new_[6251]_ ;
  assign \new_[7893]_  = \new_[8685]_  | \new_[12359]_ ;
  assign \new_[7894]_  = \new_[8685]_  | \new_[12501]_ ;
  assign \new_[7895]_  = ~\new_[8651]_  & ~\new_[5999]_ ;
  assign \new_[7896]_  = ~\new_[8692]_  | ~\new_[12423]_ ;
  assign \new_[7897]_  = \new_[8686]_  | \new_[12440]_ ;
  assign \new_[7898]_  = \new_[8686]_  | \new_[12612]_ ;
  assign \new_[7899]_  = ~\\u4_u0_buf0_orig_m3_reg[11] ;
  assign \new_[7900]_  = ~\new_[9205]_  | ~\new_[11128]_  | ~\new_[10366]_  | ~\new_[11150]_ ;
  assign \new_[7901]_  = ~\new_[8699]_  & ~\new_[6274]_ ;
  assign \new_[7902]_  = \new_[8687]_  | \new_[12294]_ ;
  assign \new_[7903]_  = \new_[8687]_  | \new_[12618]_ ;
  assign \new_[7904]_  = ~\new_[8676]_  | ~\new_[8731]_ ;
  assign \new_[7905]_  = ~\new_[8671]_  & ~\new_[6286]_ ;
  assign \new_[7906]_  = \new_[6738]_  ^ \new_[9110]_ ;
  assign \new_[7907]_  = (~\new_[12587]_  | ~\new_[11942]_ ) & (~\new_[9075]_  | ~\new_[12519]_ );
  assign \new_[7908]_  = ~\new_[9055]_  | ~\new_[8858]_ ;
  assign \new_[7909]_  = ~\new_[8297]_ ;
  assign \new_[7910]_  = ~\new_[8691]_  | ~\new_[8856]_ ;
  assign \new_[7911]_  = \new_[11994]_  ^ \new_[9076]_ ;
  assign \new_[7912]_  = \new_[11825]_  ^ \new_[9078]_ ;
  assign \new_[7913]_  = \new_[11983]_  ^ \new_[9077]_ ;
  assign \new_[7914]_  = \new_[11767]_  ^ \new_[9079]_ ;
  assign \new_[7915]_  = (~\new_[9104]_  | ~\wb_data_i[0] ) & (~\new_[9402]_  | ~\new_[6611]_ );
  assign \new_[7916]_  = (~\new_[9104]_  | ~\wb_data_i[1] ) & (~\new_[9402]_  | ~\new_[6721]_ );
  assign \new_[7917]_  = (~\new_[9104]_  | ~\wb_data_i[2] ) & (~\new_[9402]_  | ~\new_[6609]_ );
  assign \new_[7918]_  = (~\new_[9104]_  | ~\wb_data_i[3] ) & (~\new_[9402]_  | ~\new_[6722]_ );
  assign \new_[7919]_  = (~\new_[9104]_  | ~\wb_data_i[4] ) & (~\new_[9402]_  | ~\new_[6610]_ );
  assign \new_[7920]_  = (~\new_[9104]_  | ~\wb_data_i[5] ) & (~\new_[9402]_  | ~\new_[6723]_ );
  assign \new_[7921]_  = (~\new_[9104]_  | ~\wb_data_i[6] ) & (~\new_[9402]_  | ~\new_[6724]_ );
  assign \new_[7922]_  = (~\new_[9104]_  | ~\wb_data_i[7] ) & (~\new_[9402]_  | ~\new_[13995]_ );
  assign \new_[7923]_  = (~\new_[9104]_  | ~\wb_data_i[8] ) & (~\new_[9402]_  | ~\new_[14074]_ );
  assign \new_[7924]_  = (~\new_[9104]_  | ~\wb_data_i[16] ) & (~\new_[9402]_  | ~\new_[13702]_ );
  assign \new_[7925]_  = (~\new_[9104]_  | ~\wb_data_i[17] ) & (~\new_[9402]_  | ~\new_[14164]_ );
  assign \new_[7926]_  = (~\new_[9104]_  | ~\wb_data_i[18] ) & (~\new_[9402]_  | ~\new_[13512]_ );
  assign \new_[7927]_  = (~\new_[9104]_  | ~\wb_data_i[19] ) & (~\new_[9402]_  | ~\new_[13734]_ );
  assign \new_[7928]_  = (~\new_[9104]_  | ~\wb_data_i[20] ) & (~\new_[9402]_  | ~\new_[13712]_ );
  assign \new_[7929]_  = (~\new_[9104]_  | ~\wb_data_i[21] ) & (~\new_[9402]_  | ~\new_[14110]_ );
  assign \new_[7930]_  = (~\new_[9104]_  | ~\wb_data_i[22] ) & (~\new_[9402]_  | ~\new_[14081]_ );
  assign \new_[7931]_  = (~\new_[9104]_  | ~\wb_data_i[23] ) & (~\new_[9402]_  | ~\new_[14208]_ );
  assign \new_[7932]_  = (~\new_[9104]_  | ~\wb_data_i[24] ) & (~\new_[9402]_  | ~\new_[13763]_ );
  assign \new_[7933]_  = \new_[6737]_  ^ \new_[9121]_ ;
  assign \new_[7934]_  = ~\new_[8827]_  | ~\new_[9191]_ ;
  assign \new_[7935]_  = ~\new_[8718]_  | ~\new_[3592]_ ;
  assign \new_[7936]_  = ~\new_[8717]_  | ~\new_[4286]_ ;
  assign \new_[7937]_  = \new_[8628]_  | \new_[8841]_ ;
  assign \new_[7938]_  = ~\new_[12690]_  | ~\new_[8923]_  | ~\new_[9033]_ ;
  assign \new_[7939]_  = ~\new_[9106]_  | ~\new_[11490]_  | ~\new_[11255]_ ;
  assign \new_[7940]_  = \new_[8822]_  | \new_[10796]_ ;
  assign \new_[7941]_  = ~\\u4_u0_buf0_orig_m3_reg[9] ;
  assign \new_[7942]_  = ~\\u4_u2_buf0_orig_m3_reg[9] ;
  assign \new_[7943]_  = ~u4_u1_int_re_reg;
  assign \new_[7944]_  = ~\\u4_u0_buf0_orig_m3_reg[10] ;
  assign \new_[7945]_  = ~u4_u2_int_re_reg;
  assign \new_[7946]_  = ~u4_u0_int_re_reg;
  assign \new_[7947]_  = ~\new_[8323]_ ;
  assign \new_[7948]_  = ~\\u4_u2_buf0_orig_m3_reg[10] ;
  assign \new_[7949]_  = ~\new_[8921]_  | ~\new_[10087]_ ;
  assign \new_[7950]_  = ~\new_[9276]_  & (~\new_[9478]_  | ~\new_[8974]_ );
  assign \new_[7951]_  = ~\new_[8886]_  | ~\new_[6592]_ ;
  assign \new_[7952]_  = ~\new_[13720]_  | ~\new_[8860]_ ;
  assign \new_[7953]_  = ~\new_[8860]_  | ~\new_[6300]_ ;
  assign \new_[7954]_  = ~\new_[8860]_  | ~\new_[6302]_ ;
  assign \new_[7955]_  = ~\new_[8860]_  | ~\new_[6588]_ ;
  assign \new_[7956]_  = ~\new_[8860]_  | ~\new_[6303]_ ;
  assign \new_[7957]_  = ~\new_[8860]_  | ~\new_[6304]_ ;
  assign \new_[7958]_  = ~\new_[8860]_  | ~\new_[6305]_ ;
  assign \new_[7959]_  = ~\new_[8860]_  | ~\new_[6301]_ ;
  assign \new_[7960]_  = ~\new_[14125]_  | ~\new_[8860]_ ;
  assign \new_[7961]_  = ~\new_[13534]_  | ~\new_[8860]_ ;
  assign \new_[7962]_  = ~\new_[14239]_  | ~\new_[8860]_ ;
  assign \new_[7963]_  = ~\new_[9145]_  | ~\wb_data_i[4] ;
  assign \new_[7964]_  = ~\new_[8805]_  & (~\new_[14636]_  | ~\new_[2348]_ );
  assign \new_[7965]_  = ~\new_[14223]_  | ~\new_[8860]_ ;
  assign \new_[7966]_  = ~\new_[13574]_  | ~\new_[8860]_ ;
  assign \new_[7967]_  = ~\new_[8860]_  | ~\new_[6299]_ ;
  assign \new_[7968]_  = ~\new_[14064]_  | ~\new_[8860]_ ;
  assign \new_[7969]_  = ~\new_[14121]_  | ~\new_[8860]_ ;
  assign \new_[7970]_  = ~\new_[8860]_  | ~\new_[13634]_ ;
  assign \new_[7971]_  = ~\new_[14160]_  | ~\new_[8884]_ ;
  assign \new_[7972]_  = ~\new_[14047]_  | ~\new_[9138]_ ;
  assign \new_[7973]_  = ~\new_[13672]_  | ~\new_[9138]_ ;
  assign \new_[7974]_  = ~\new_[14176]_  | ~\new_[9138]_ ;
  assign \new_[7975]_  = ~\new_[13693]_  | ~\new_[9138]_ ;
  assign \new_[7976]_  = ~\new_[14128]_  | ~\new_[8885]_ ;
  assign \new_[7977]_  = ~\new_[13677]_  | ~\new_[9138]_ ;
  assign \new_[7978]_  = ~\new_[13637]_  | ~\new_[9138]_ ;
  assign \new_[7979]_  = ~\new_[14091]_  | ~\new_[8884]_ ;
  assign \new_[7980]_  = ~\new_[13968]_  | ~\new_[8885]_ ;
  assign \new_[7981]_  = ~\new_[8886]_  | ~\new_[6341]_ ;
  assign \new_[7982]_  = ~\new_[13892]_  | ~\new_[8885]_ ;
  assign \new_[7983]_  = ~\new_[8886]_  | ~\new_[6343]_ ;
  assign \new_[7984]_  = ~\new_[8884]_  | ~\new_[6345]_ ;
  assign \new_[7985]_  = ~\new_[8886]_  | ~\new_[6551]_ ;
  assign \new_[7986]_  = ~\new_[8884]_  | ~\new_[6346]_ ;
  assign \new_[7987]_  = ~\new_[8886]_  | ~\new_[6347]_ ;
  assign \new_[7988]_  = ~\new_[8884]_  | ~\new_[6348]_ ;
  assign \new_[7989]_  = ~\new_[8884]_  | ~\new_[6512]_ ;
  assign \new_[7990]_  = ~\new_[9138]_  | ~\new_[6351]_ ;
  assign \new_[7991]_  = ~\new_[14067]_  | ~\new_[8885]_ ;
  assign \new_[7992]_  = ~\new_[14066]_  | ~\new_[8885]_ ;
  assign \new_[7993]_  = ~\new_[13728]_  | ~\new_[9138]_ ;
  assign \new_[7994]_  = ~\new_[14087]_  | ~\new_[9138]_ ;
  assign \new_[7995]_  = ~\new_[13765]_  | ~\new_[8885]_ ;
  assign \new_[7996]_  = ~\new_[13653]_  | ~\new_[9138]_ ;
  assign \new_[7997]_  = ~\new_[13809]_  | ~\new_[9138]_ ;
  assign \new_[7998]_  = ~\new_[8884]_  | ~\new_[13880]_ ;
  assign \new_[7999]_  = ~\new_[14210]_  | ~\new_[8860]_ ;
  assign \new_[8000]_  = ~\new_[8884]_  | ~\new_[6344]_ ;
  assign \new_[8001]_  = ~\new_[8860]_  | ~\new_[6560]_ ;
  assign \new_[8002]_  = ~\new_[14049]_  | ~\new_[9138]_ ;
  assign \new_[8003]_  = ~\new_[9145]_  | ~\wb_data_i[11] ;
  assign \new_[8004]_  = ~\new_[9145]_  | ~\wb_data_i[7] ;
  assign \new_[8005]_  = ~\new_[9145]_  | ~\wb_data_i[25] ;
  assign \new_[8006]_  = ~\new_[9145]_  | ~\wb_data_i[20] ;
  assign \new_[8007]_  = \new_[14427]_  | \new_[4800]_ ;
  assign \new_[8008]_  = \new_[14587]_  & \new_[4801]_ ;
  assign \new_[8009]_  = ~\new_[9434]_  | ~\wb_data_i[19] ;
  assign \new_[8010]_  = ~\new_[6538]_  | ~\new_[9445]_ ;
  assign \new_[8011]_  = ~\new_[9434]_  | ~\wb_data_i[14] ;
  assign \new_[8012]_  = ~\new_[9445]_  | ~\new_[6289]_ ;
  assign \new_[8013]_  = ~\new_[6548]_  | ~\new_[8889]_ ;
  assign \new_[8014]_  = ~\new_[6010]_  | ~\new_[8889]_ ;
  assign \new_[8015]_  = ~\new_[6247]_  | ~\new_[8862]_ ;
  assign \new_[8016]_  = ~\new_[9434]_  | ~\wb_data_i[20] ;
  assign \new_[8017]_  = ~\new_[14098]_  | ~\new_[9426]_ ;
  assign \new_[8018]_  = ~\new_[6249]_  | ~\new_[8862]_ ;
  assign \new_[8019]_  = ~\new_[6196]_  | ~\new_[8862]_ ;
  assign \new_[8020]_  = ~\new_[6254]_  | ~\new_[8862]_ ;
  assign \new_[8021]_  = ~\new_[9426]_  | ~\new_[6256]_ ;
  assign \new_[8022]_  = ~\new_[6163]_  | ~\new_[8862]_ ;
  assign \new_[8023]_  = ~\new_[9426]_  | ~\new_[6257]_ ;
  assign \new_[8024]_  = ~\new_[9426]_  | ~\new_[6258]_ ;
  assign \new_[8025]_  = ~\new_[6260]_  | ~\new_[8862]_ ;
  assign \new_[8026]_  = ~\new_[6109]_  | ~\new_[9426]_ ;
  assign \new_[8027]_  = ~\new_[6263]_  | ~\new_[9426]_ ;
  assign \new_[8028]_  = ~\new_[8908]_  | ~\new_[6368]_ ;
  assign \new_[8029]_  = ~\new_[6281]_  | ~\new_[8881]_ ;
  assign \new_[8030]_  = ~\new_[6287]_  | ~\new_[8889]_ ;
  assign \new_[8031]_  = ~\new_[14076]_  | ~\new_[9448]_ ;
  assign \new_[8032]_  = ~\new_[6286]_  | ~\new_[8889]_ ;
  assign \new_[8033]_  = ~\new_[6544]_  | ~\new_[8889]_ ;
  assign \new_[8034]_  = ~\new_[6526]_  | ~\new_[9445]_ ;
  assign \new_[8035]_  = ~\new_[6279]_  | ~\new_[8881]_ ;
  assign \new_[8036]_  = ~\new_[8606]_ ;
  assign \new_[8037]_  = ~\new_[9106]_  | ~\new_[2209]_ ;
  assign \new_[8038]_  = ~\new_[9430]_  | ~\new_[6172]_ ;
  assign \new_[8039]_  = ~\new_[6005]_  | ~\new_[8881]_ ;
  assign \new_[8040]_  = ~\new_[9106]_  | ~\new_[2173]_ ;
  assign \new_[8041]_  = ~\new_[13438]_  | ~\new_[12420]_  | ~\new_[10285]_ ;
  assign \new_[8042]_  = ~\new_[13918]_  | ~\new_[8873]_ ;
  assign \new_[8043]_  = ~\new_[13896]_  | ~\new_[8873]_ ;
  assign \new_[8044]_  = ~\new_[13857]_  | ~\new_[8878]_ ;
  assign \new_[8045]_  = ~\new_[13700]_  | ~\new_[8874]_ ;
  assign \new_[8046]_  = ~\new_[13855]_  | ~\new_[8873]_ ;
  assign \new_[8047]_  = ~\new_[13967]_  | ~\new_[8874]_ ;
  assign \new_[8048]_  = ~\new_[13542]_  | ~\new_[8874]_ ;
  assign \new_[8049]_  = ~\new_[14080]_  | ~\new_[8874]_ ;
  assign \new_[8050]_  = ~\new_[14054]_  | ~\new_[8873]_ ;
  assign \new_[8051]_  = ~\new_[13808]_  | ~\new_[8878]_ ;
  assign \new_[8052]_  = ~\new_[8878]_  | ~\new_[6484]_ ;
  assign \new_[8053]_  = ~\new_[13829]_  | ~\new_[9380]_ ;
  assign \new_[8054]_  = ~\new_[8878]_  | ~\new_[6168]_ ;
  assign \new_[8055]_  = ~\new_[8875]_  | ~\new_[6319]_ ;
  assign \new_[8056]_  = ~\new_[8875]_  | ~\new_[6232]_ ;
  assign \new_[8057]_  = ~\new_[8875]_  | ~\new_[6320]_ ;
  assign \new_[8058]_  = ~\new_[8878]_  | ~\new_[6238]_ ;
  assign \new_[8059]_  = ~\new_[8878]_  | ~\new_[6322]_ ;
  assign \new_[8060]_  = ~\new_[8875]_  | ~\new_[6234]_ ;
  assign \new_[8061]_  = ~\new_[8875]_  | ~\new_[6323]_ ;
  assign \new_[8062]_  = ~\new_[8878]_  | ~\new_[6198]_ ;
  assign \new_[8063]_  = ~\new_[8877]_  | ~\new_[6324]_ ;
  assign \new_[8064]_  = ~\new_[14095]_  | ~\new_[9380]_ ;
  assign \new_[8065]_  = ~\new_[8877]_  | ~\new_[6326]_ ;
  assign \new_[8066]_  = ~\new_[13507]_  | ~\new_[9380]_ ;
  assign \new_[8067]_  = ~\new_[14252]_  | ~\new_[8873]_ ;
  assign \new_[8068]_  = ~\new_[14258]_  | ~\new_[8874]_ ;
  assign \new_[8069]_  = ~\new_[14016]_  | ~\new_[9380]_ ;
  assign \new_[8070]_  = ~\new_[14006]_  | ~\new_[9380]_ ;
  assign \new_[8071]_  = ~\new_[14194]_  | ~\new_[8873]_ ;
  assign \new_[8072]_  = ~\new_[13559]_  | ~\new_[9380]_ ;
  assign \new_[8073]_  = ~\new_[8875]_  | ~\new_[14179]_ ;
  assign \new_[8074]_  = ~\new_[6004]_  | ~\new_[8881]_ ;
  assign \new_[8075]_  = ~\new_[9426]_  | ~\new_[13884]_ ;
  assign \new_[8076]_  = ~\new_[6003]_  | ~\new_[8881]_ ;
  assign \new_[8077]_  = ~\new_[8910]_  | ~\new_[6556]_ ;
  assign \new_[8078]_  = ~\new_[8911]_  | ~\new_[6366]_ ;
  assign \new_[8079]_  = ~\new_[6008]_  | ~\new_[8889]_ ;
  assign \new_[8080]_  = ~\new_[6562]_  | ~\new_[8889]_ ;
  assign \new_[8081]_  = ~\new_[13922]_  | ~\new_[9445]_ ;
  assign \new_[8082]_  = ~\new_[13500]_  | ~\new_[9429]_ ;
  assign \new_[8083]_  = ~\new_[6264]_  | ~\new_[8880]_ ;
  assign \new_[8084]_  = ~\new_[14123]_  | ~\new_[8880]_ ;
  assign \new_[8085]_  = ~\new_[13894]_  | ~\new_[8880]_ ;
  assign \new_[8086]_  = ~\new_[6599]_  | ~\new_[9429]_ ;
  assign \new_[8087]_  = ~\new_[5998]_  | ~\new_[9429]_ ;
  assign \new_[8088]_  = ~\new_[6593]_  | ~\new_[8880]_ ;
  assign \new_[8089]_  = ~\new_[5999]_  | ~\new_[8880]_ ;
  assign \new_[8090]_  = ~\new_[6563]_  | ~\new_[9429]_ ;
  assign \new_[8091]_  = ~\new_[6266]_  | ~\new_[8880]_ ;
  assign \new_[8092]_  = ~\new_[6567]_  | ~\new_[9429]_ ;
  assign \new_[8093]_  = ~\new_[6561]_  | ~\new_[8880]_ ;
  assign \new_[8094]_  = ~\new_[6292]_  | ~\new_[9445]_ ;
  assign \new_[8095]_  = ~\new_[8880]_  | ~\new_[6267]_ ;
  assign \new_[8096]_  = ~\new_[6524]_  | ~\new_[8880]_ ;
  assign \new_[8097]_  = ~\new_[8880]_  | ~\new_[6539]_ ;
  assign \new_[8098]_  = ~\new_[8880]_  | ~\new_[6543]_ ;
  assign \new_[8099]_  = ~\new_[6000]_  | ~\new_[9429]_ ;
  assign \new_[8100]_  = ~\new_[6001]_  | ~\new_[8880]_ ;
  assign \new_[8101]_  = ~\new_[6002]_  | ~\new_[8880]_ ;
  assign \new_[8102]_  = ~\new_[6547]_  | ~\new_[8880]_ ;
  assign \new_[8103]_  = ~\new_[6268]_  | ~\new_[8880]_ ;
  assign \new_[8104]_  = ~\new_[6549]_  | ~\new_[9429]_ ;
  assign \new_[8105]_  = ~\new_[6269]_  | ~\new_[8880]_ ;
  assign \new_[8106]_  = ~\new_[13750]_  | ~\new_[8889]_ ;
  assign \new_[8107]_  = ~\new_[6237]_  | ~\new_[9430]_ ;
  assign \new_[8108]_  = ~\new_[14229]_  | ~\new_[8907]_ ;
  assign \new_[8109]_  = ~\new_[6291]_  | ~\new_[8889]_ ;
  assign \new_[8110]_  = ~\new_[13807]_  | ~\new_[9430]_ ;
  assign \new_[8111]_  = ~\new_[8911]_  | ~\new_[6369]_ ;
  assign \new_[8112]_  = ~\new_[6284]_  | ~\new_[8889]_ ;
  assign \new_[8113]_  = ~\new_[6250]_  | ~\new_[8862]_ ;
  assign \new_[8114]_  = ~\new_[6253]_  | ~\new_[8862]_ ;
  assign \new_[8115]_  = ~\new_[13597]_  | ~\new_[8862]_ ;
  assign \new_[8116]_  = ~\new_[6557]_  | ~\new_[9429]_ ;
  assign \new_[8117]_  = ~\new_[6252]_  | ~\new_[8862]_ ;
  assign \new_[8118]_  = ~\new_[6086]_  | ~\new_[8862]_ ;
  assign \new_[8119]_  = ~\new_[6262]_  | ~\new_[9426]_ ;
  assign \new_[8120]_  = ~\new_[9445]_  | ~\new_[13711]_ ;
  assign \new_[8121]_  = ~\new_[13848]_  | ~\new_[9445]_ ;
  assign \new_[8122]_  = ~\new_[14155]_  | ~\new_[8862]_ ;
  assign \new_[8123]_  = ~\new_[6261]_  | ~\new_[9426]_ ;
  assign \new_[8124]_  = ~\new_[8855]_  | ~phy_rst_pad_o;
  assign \new_[8125]_  = ~\new_[9106]_  & ~\new_[2175]_ ;
  assign \new_[8126]_  = ~\new_[8880]_  | ~\new_[13768]_ ;
  assign \new_[8127]_  = ~\new_[6259]_  | ~\new_[8862]_ ;
  assign \new_[8128]_  = ~\new_[9106]_  & ~\new_[13845]_ ;
  assign \new_[8129]_  = ~\new_[9434]_  | ~\wb_data_i[10] ;
  assign \new_[8130]_  = ~\new_[9434]_  | ~\wb_data_i[16] ;
  assign \new_[8131]_  = ~\new_[9434]_  | ~\wb_data_i[17] ;
  assign \new_[8132]_  = ~\new_[9434]_  | ~\wb_data_i[26] ;
  assign \new_[8133]_  = ~\new_[9434]_  | ~\wb_data_i[31] ;
  assign \new_[8134]_  = ~\new_[9140]_  | ~\new_[10479]_ ;
  assign \new_[8135]_  = ~\new_[6255]_  | ~\new_[9426]_ ;
  assign \new_[8136]_  = ~\new_[6293]_  | ~\new_[9445]_ ;
  assign \new_[8137]_  = ~\new_[13764]_  | ~\new_[9430]_ ;
  assign \new_[8138]_  = ~\new_[6272]_  | ~\new_[8881]_ ;
  assign \new_[8139]_  = ~\new_[9048]_  | ~\wb_data_i[12] ;
  assign \new_[8140]_  = ~\new_[14192]_  | ~\new_[9430]_ ;
  assign \new_[8141]_  = ~\new_[9048]_  | ~\wb_data_i[1] ;
  assign \new_[8142]_  = ~\new_[6274]_  | ~\new_[8881]_ ;
  assign \new_[8143]_  = ~\new_[6200]_  | ~\new_[8881]_ ;
  assign \new_[8144]_  = ~\new_[6275]_  | ~\new_[8881]_ ;
  assign \new_[8145]_  = ~\new_[9048]_  | ~\wb_data_i[7] ;
  assign \new_[8146]_  = ~\new_[6166]_  | ~\new_[8881]_ ;
  assign \new_[8147]_  = ~\new_[9430]_  | ~\new_[6276]_ ;
  assign \new_[8148]_  = ~\new_[13946]_  | ~\new_[9430]_ ;
  assign \new_[8149]_  = ~\new_[9430]_  | ~\new_[6277]_ ;
  assign \new_[8150]_  = ~\new_[13610]_  | ~\new_[9430]_ ;
  assign \new_[8151]_  = ~\new_[14172]_  | ~\new_[8881]_ ;
  assign \new_[8152]_  = ~\new_[9048]_  | ~\wb_data_i[17] ;
  assign \new_[8153]_  = ~\new_[6089]_  | ~\new_[9430]_ ;
  assign \new_[8154]_  = ~\new_[9048]_  | ~\wb_data_i[19] ;
  assign \new_[8155]_  = ~\new_[6280]_  | ~\new_[9430]_ ;
  assign \new_[8156]_  = ~\new_[14009]_  | ~\new_[8881]_ ;
  assign \new_[8157]_  = ~\new_[6251]_  | ~\new_[8862]_ ;
  assign \new_[8158]_  = ~\new_[6290]_  | ~\new_[9445]_ ;
  assign \new_[8159]_  = ~\new_[14259]_  | ~\new_[9448]_ ;
  assign \new_[8160]_  = ~\new_[9213]_  & (~\new_[9185]_  | ~\new_[9189]_ );
  assign \new_[8161]_  = ~\new_[8857]_  & ~\new_[13355]_ ;
  assign \new_[8162]_  = ~\new_[8854]_  & ~\new_[12911]_ ;
  assign \new_[8163]_  = ~\new_[9430]_  | ~\new_[14078]_ ;
  assign \new_[8164]_  = ~\new_[13797]_  | ~\new_[8907]_ ;
  assign \new_[8165]_  = \new_[11291]_  ^ \new_[9022]_ ;
  assign \new_[8166]_  = ~\new_[14246]_  | ~\new_[9448]_ ;
  assign \new_[8167]_  = ~\new_[13805]_  | ~\new_[9448]_ ;
  assign \new_[8168]_  = ~\new_[14002]_  | ~\new_[8911]_ ;
  assign \new_[8169]_  = ~\new_[13783]_  | ~\new_[8907]_ ;
  assign \new_[8170]_  = ~\new_[13787]_  | ~\new_[9448]_ ;
  assign \new_[8171]_  = ~\new_[14107]_  | ~\new_[8907]_ ;
  assign \new_[8172]_  = ~\new_[14101]_  | ~\new_[9448]_ ;
  assign \new_[8173]_  = ~\new_[13938]_  | ~\new_[9448]_ ;
  assign \new_[8174]_  = ~\new_[14214]_  | ~\new_[8907]_ ;
  assign \new_[8175]_  = ~\new_[8911]_  | ~\new_[6365]_ ;
  assign \new_[8176]_  = ~\new_[14150]_  | ~\new_[8907]_ ;
  assign \new_[8177]_  = ~\new_[8911]_  | ~\new_[6367]_ ;
  assign \new_[8178]_  = ~\new_[8908]_  | ~\new_[6102]_ ;
  assign \new_[8179]_  = ~\new_[8911]_  | ~\new_[6370]_ ;
  assign \new_[8180]_  = ~\new_[8908]_  | ~\new_[6091]_ ;
  assign \new_[8181]_  = \new_[11288]_  ^ \new_[9023]_ ;
  assign \new_[8182]_  = ~\new_[9448]_  | ~\new_[6461]_ ;
  assign \new_[8183]_  = ~\new_[13973]_  | ~\new_[9448]_ ;
  assign \new_[8184]_  = ~\new_[14243]_  | ~\new_[9448]_ ;
  assign \new_[8185]_  = ~\new_[14257]_  | ~\new_[8911]_ ;
  assign \new_[8186]_  = ~\new_[14017]_  | ~\new_[9448]_ ;
  assign \new_[8187]_  = ~\new_[8908]_  | ~\new_[13519]_ ;
  assign \new_[8188]_  = ~\new_[9434]_  | ~\wb_data_i[29] ;
  assign \new_[8189]_  = \new_[11293]_  ^ \new_[9024]_ ;
  assign \new_[8190]_  = ~\new_[6009]_  | ~\new_[8889]_ ;
  assign \new_[8191]_  = ~\new_[6552]_  | ~\new_[8889]_ ;
  assign \new_[8192]_  = ~\new_[9445]_  | ~\new_[6288]_ ;
  assign \new_[8193]_  = ~\new_[9445]_  | ~\new_[6545]_ ;
  assign \new_[8194]_  = ~\new_[6485]_  | ~\new_[9445]_ ;
  assign \new_[8195]_  = ~\new_[8908]_  | ~\new_[6092]_ ;
  assign \new_[8196]_  = ~\new_[8908]_  | ~\new_[6371]_ ;
  assign \new_[8197]_  = ~\new_[14263]_  | ~\new_[9448]_ ;
  assign \new_[8198]_  = \new_[11292]_  ^ \new_[9025]_ ;
  assign \new_[8199]_  = ~\new_[8891]_  & ~\new_[8975]_ ;
  assign \new_[8200]_  = ~\new_[9915]_  | ~\new_[9546]_  | ~\new_[8966]_ ;
  assign \new_[8201]_  = ~\new_[11330]_  & (~\new_[8967]_  | ~\new_[10130]_ );
  assign \new_[8202]_  = ~\new_[8564]_ ;
  assign \new_[8203]_  = ~\new_[8568]_ ;
  assign \new_[8204]_  = ~\new_[8569]_ ;
  assign \new_[8205]_  = ~\new_[8892]_  & (~\new_[2961]_  | ~\new_[13327]_ );
  assign \new_[8206]_  = \\u4_u3_dma_out_left_reg[6] ;
  assign \new_[8207]_  = \\u4_u0_dma_out_left_reg[6] ;
  assign \new_[8208]_  = \\u4_u1_dma_out_left_reg[6] ;
  assign \new_[8209]_  = \\u4_dout_reg[14] ;
  assign \new_[8210]_  = \\u4_u2_dma_out_left_reg[6] ;
  assign \new_[8211]_  = ~\new_[12524]_  | ~\new_[8924]_  | ~\new_[9034]_ ;
  assign n7570 = ~\new_[8952]_  | ~\new_[8953]_ ;
  assign n7575 = ~\new_[8956]_  | ~\new_[8938]_ ;
  assign \new_[8214]_  = \new_[8961]_  & \new_[9562]_ ;
  assign \new_[8215]_  = \new_[8936]_  & \new_[9562]_ ;
  assign \new_[8216]_  = ~\new_[9574]_  | ~\new_[8941]_ ;
  assign \new_[8217]_  = ~\new_[10095]_  | ~\new_[4791]_  | ~\new_[12114]_  | ~\new_[8978]_ ;
  assign \new_[8218]_  = ~\new_[8957]_  & ~\new_[9218]_ ;
  assign \new_[8219]_  = (~\new_[9769]_  | ~\new_[10840]_ ) & (~\new_[8979]_  | ~\new_[13257]_ );
  assign \new_[8220]_  = (~\new_[9125]_  | ~\new_[3788]_ ) & (~\new_[9038]_  | ~\new_[3711]_ );
  assign \new_[8221]_  = ~\new_[8597]_ ;
  assign \new_[8222]_  = ~\new_[8599]_ ;
  assign \new_[8223]_  = ~\new_[14422]_ ;
  assign \new_[8224]_  = ~\new_[14585]_ ;
  assign \new_[8225]_  = ~\new_[14788]_ ;
  assign \new_[8226]_  = (~\new_[9020]_  | ~\new_[4820]_ ) & (~\new_[14537]_  | ~\new_[4843]_ );
  assign n7585 = \new_[8646]_  & \new_[9900]_ ;
  assign n7580 = \new_[8647]_  & \new_[9901]_ ;
  assign \new_[8229]_  = ~\new_[8608]_ ;
  assign \new_[8230]_  = ~\new_[8610]_ ;
  assign \new_[8231]_  = \new_[8633]_  & \new_[13370]_ ;
  assign \new_[8232]_  = ~\new_[8649]_  & ~\new_[12383]_ ;
  assign \new_[8233]_  = ~\new_[8633]_  | ~\new_[6023]_ ;
  assign \new_[8234]_  = ~\new_[9276]_  & ~\new_[8642]_ ;
  assign \new_[8235]_  = ~\new_[9232]_  & (~\new_[11598]_  | ~\new_[13084]_ );
  assign \new_[8236]_  = ~\new_[8622]_ ;
  assign \new_[8237]_  = \new_[8633]_  & \new_[9611]_ ;
  assign \new_[8238]_  = ~\new_[14345]_ ;
  assign \new_[8239]_  = ~\new_[13327]_  | ~\new_[8635]_  | ~\new_[13436]_ ;
  assign \new_[8240]_  = ~\new_[8627]_ ;
  assign \new_[8241]_  = \new_[8633]_  & \new_[12838]_ ;
  assign \new_[8242]_  = ~\new_[12838]_  | ~\new_[8970]_ ;
  assign \new_[8243]_  = \new_[10491]_  & \new_[8978]_ ;
  assign \new_[8244]_  = \new_[14268]_  ^ \new_[9364]_ ;
  assign \new_[8245]_  = \new_[12798]_  ? \new_[9375]_  : \new_[2477]_ ;
  assign \new_[8246]_  = ~\new_[8980]_  & (~\new_[10811]_  | ~\new_[10096]_ );
  assign \new_[8247]_  = u4_u1_ep_match_r_reg;
  assign \new_[8248]_  = ~\new_[9031]_  & ~\new_[13418]_ ;
  assign \new_[8249]_  = ~\new_[9031]_  & ~\new_[13453]_ ;
  assign \new_[8250]_  = ~\new_[9031]_  & ~\new_[13328]_ ;
  assign \new_[8251]_  = ~\new_[9031]_  & ~\new_[13349]_ ;
  assign \new_[8252]_  = ~\new_[9031]_  & ~\new_[13449]_ ;
  assign \new_[8253]_  = ~\new_[9031]_  & ~\new_[13433]_ ;
  assign \new_[8254]_  = ~\new_[9031]_  & ~\new_[13446]_ ;
  assign \new_[8255]_  = ~\new_[9031]_  & ~\new_[13343]_ ;
  assign n7635 = ~\new_[12125]_  & ~\new_[9032]_ ;
  assign \new_[8257]_  = \new_[9610]_  & \new_[9036]_ ;
  assign \new_[8258]_  = ~\new_[2479]_  & ~n7590;
  assign \new_[8259]_  = ~\new_[9834]_  | ~n8990;
  assign \new_[8260]_  = (~\new_[9371]_  | ~\new_[11727]_ ) & (~\new_[13315]_  | ~\new_[3463]_ );
  assign \new_[8261]_  = ~\new_[14313]_ ;
  assign \new_[8262]_  = ~\new_[9728]_  | ~\new_[11852]_  | ~\new_[10350]_  | ~\new_[13454]_ ;
  assign \new_[8263]_  = ~\new_[9045]_  | ~\new_[11569]_ ;
  assign \new_[8264]_  = ~\new_[9041]_  | ~\new_[11856]_ ;
  assign \new_[8265]_  = ~\new_[9041]_  & ~\new_[11623]_ ;
  assign \new_[8266]_  = ~\new_[9603]_  & ~\new_[4092]_ ;
  assign \new_[8267]_  = \new_[9603]_  | \new_[13778]_ ;
  assign \new_[8268]_  = \new_[14094]_  ? \new_[9377]_  : \new_[2085]_ ;
  assign \new_[8269]_  = ~\new_[9036]_  | ~\new_[4795]_ ;
  assign \new_[8270]_  = ~\new_[9042]_  & ~\new_[11628]_ ;
  assign \new_[8271]_  = ~\new_[9042]_  | ~\new_[12050]_ ;
  assign \new_[8272]_  = ~\new_[10859]_  & ~\new_[9043]_ ;
  assign \new_[8273]_  = ~\new_[9044]_  & ~\new_[11630]_ ;
  assign \new_[8274]_  = ~\new_[9044]_  | ~\new_[11561]_ ;
  assign \new_[8275]_  = ~\new_[9038]_  | ~\new_[3788]_ ;
  assign \new_[8276]_  = ~\new_[9045]_  & ~\new_[11289]_ ;
  assign \new_[8277]_  = ~\new_[11912]_  & (~\new_[9460]_  | ~\new_[12291]_ );
  assign \new_[8278]_  = ~\new_[11827]_  & (~\new_[9353]_  | ~\new_[11952]_ );
  assign \new_[8279]_  = ~\new_[11829]_  & (~\new_[9350]_  | ~\new_[12738]_ );
  assign \new_[8280]_  = ~\new_[11831]_  & (~\new_[9306]_  | ~\new_[12305]_ );
  assign \new_[8281]_  = ~\new_[8666]_ ;
  assign \new_[8282]_  = ~\new_[9125]_  | ~\new_[9038]_ ;
  assign \new_[8283]_  = ~\new_[9215]_  | (~\new_[9378]_  & ~\new_[9857]_ );
  assign \new_[8284]_  = ~\new_[9739]_  | ~\new_[11846]_  | ~\new_[10351]_  | ~\new_[13388]_ ;
  assign \new_[8285]_  = \new_[10331]_  ^ \new_[9382]_ ;
  assign \new_[8286]_  = \new_[10333]_  ^ \new_[9383]_ ;
  assign \new_[8287]_  = ~\new_[12987]_  & (~\new_[9418]_  | ~\new_[3691]_ );
  assign \new_[8288]_  = \new_[2341]_  ^ \new_[9458]_ ;
  assign \new_[8289]_  = ~\new_[10377]_  | ~\new_[10024]_  | ~\new_[8971]_  | ~\new_[11523]_ ;
  assign \new_[8290]_  = ~\new_[10625]_  | ~\new_[10023]_  | ~\new_[9040]_  | ~\new_[11709]_ ;
  assign \new_[8291]_  = ~\\u4_u3_buf0_orig_m3_reg[11] ;
  assign \new_[8292]_  = ~\\u4_u2_buf0_orig_m3_reg[11] ;
  assign \new_[8293]_  = ~\new_[9222]_  | (~\new_[9643]_  & ~\new_[9857]_ );
  assign \new_[8294]_  = (~\new_[12614]_  | ~\new_[11942]_ ) & (~\new_[9388]_  | ~\new_[12519]_ );
  assign \new_[8295]_  = (~\new_[12559]_  | ~\new_[11942]_ ) & (~\new_[9392]_  | ~\new_[12519]_ );
  assign \new_[8296]_  = (~\new_[12848]_  | ~\new_[11942]_ ) & (~\new_[12519]_  | ~\new_[9389]_ );
  assign \new_[8297]_  = ~\new_[9054]_  | ~\new_[9419]_ ;
  assign \new_[8298]_  = ~\\u4_u0_dma_out_left_reg[5] ;
  assign \new_[8299]_  = ~\\u4_u3_dma_out_left_reg[5] ;
  assign \new_[8300]_  = ~\\u4_u1_dma_out_left_reg[5] ;
  assign \new_[8301]_  = ~\\u4_u2_dma_out_left_reg[5] ;
  assign n7640 = ~\new_[13296]_  & (~\new_[13346]_  | ~\new_[9431]_ );
  assign \new_[8303]_  = ~\new_[9085]_  & ~\new_[13469]_ ;
  assign \new_[8304]_  = \new_[9083]_  | \new_[12412]_ ;
  assign \new_[8305]_  = \new_[9094]_  | \new_[12290]_ ;
  assign \new_[8306]_  = ~\\u4_u1_buf0_orig_m3_reg[7] ;
  assign \new_[8307]_  = ~\new_[10373]_  | ~\new_[10022]_  | ~\new_[9107]_  | ~\new_[11525]_ ;
  assign \new_[8308]_  = ~\new_[6246]_  & (~\new_[9437]_  | ~\new_[9469]_ );
  assign \new_[8309]_  = \new_[9096]_  | \new_[12473]_ ;
  assign \new_[8310]_  = \new_[9105]_  & \new_[9810]_ ;
  assign \new_[8311]_  = ~\new_[10379]_  | ~\new_[10021]_  | ~\new_[9108]_  | ~\new_[11518]_ ;
  assign \new_[8312]_  = ~\new_[9642]_  & ~\new_[9111]_ ;
  assign \new_[8313]_  = \new_[9099]_  | \new_[12470]_ ;
  assign \new_[8314]_  = ~\\u4_u1_buf0_orig_m3_reg[8] ;
  assign n7625 = \wb_data_i[0]  ? \new_[9431]_  : n9040;
  assign n7615 = \wb_data_i[1]  ? \new_[9431]_  : n9075;
  assign n7630 = \wb_data_i[3]  ? \new_[9431]_  : n9030;
  assign n7595 = \wb_data_i[2]  ? \new_[9431]_  : n9050;
  assign \new_[8319]_  = \new_[11969]_  ^ \new_[9452]_ ;
  assign n7600 = \new_[11631]_  ^ \new_[9451]_ ;
  assign \new_[8321]_  = \new_[11972]_  ^ \new_[9453]_ ;
  assign \new_[8322]_  = ~\new_[8719]_ ;
  assign \new_[8323]_  = ~\\u4_u1_buf0_orig_m3_reg[10] ;
  assign n7645 = ~\new_[9154]_  & ~\new_[12842]_ ;
  assign \new_[8325]_  = ~\new_[14260]_  | ~\new_[9425]_ ;
  assign \new_[8326]_  = ~\new_[13874]_  | ~\new_[9425]_ ;
  assign \new_[8327]_  = ~\new_[13907]_  | ~\new_[9425]_ ;
  assign \new_[8328]_  = ~\new_[9128]_  | ~\new_[6602]_ ;
  assign \new_[8329]_  = ~\new_[14133]_  | ~\new_[9425]_ ;
  assign \new_[8330]_  = ~\new_[14217]_  | ~\new_[9425]_ ;
  assign \new_[8331]_  = ~\new_[9144]_  | ~\wb_data_i[26] ;
  assign \new_[8332]_  = ~\new_[9144]_  | ~\wb_data_i[15] ;
  assign \new_[8333]_  = \new_[9159]_  & \new_[9780]_ ;
  assign \new_[8334]_  = ~\new_[9143]_  | ~\wb_data_i[8] ;
  assign \new_[8335]_  = ~\new_[13721]_  | ~\new_[9425]_ ;
  assign \new_[8336]_  = ~\new_[9068]_  | ~\wb_data_i[0] ;
  assign \new_[8337]_  = ~\new_[9134]_  | ~\wb_data_i[10] ;
  assign \new_[8338]_  = ~\new_[9089]_  & (~\new_[14636]_  | ~\new_[2343]_ );
  assign \new_[8339]_  = ~\new_[9134]_  | ~\wb_data_i[11] ;
  assign \new_[8340]_  = ~\new_[9068]_  | ~\wb_data_i[12] ;
  assign \new_[8341]_  = ~\new_[9134]_  | ~\wb_data_i[13] ;
  assign \new_[8342]_  = ~\new_[9134]_  | ~\wb_data_i[14] ;
  assign \new_[8343]_  = ~\new_[9133]_  | ~\wb_data_i[15] ;
  assign \new_[8344]_  = ~\new_[9067]_  | ~\wb_data_i[16] ;
  assign \new_[8345]_  = ~\new_[9067]_  | ~\wb_data_i[17] ;
  assign \new_[8346]_  = ~\new_[9067]_  | ~\wb_data_i[18] ;
  assign \new_[8347]_  = ~\new_[9132]_  | ~\wb_data_i[19] ;
  assign \new_[8348]_  = ~\new_[9067]_  | ~\wb_data_i[1] ;
  assign \new_[8349]_  = ~\new_[9132]_  | ~\wb_data_i[20] ;
  assign \new_[8350]_  = ~\new_[9134]_  | ~\wb_data_i[21] ;
  assign \new_[8351]_  = ~\new_[9133]_  | ~\wb_data_i[22] ;
  assign \new_[8352]_  = ~\new_[9133]_  | ~\wb_data_i[23] ;
  assign \new_[8353]_  = ~\new_[9133]_  | ~\wb_data_i[24] ;
  assign \new_[8354]_  = ~\new_[9067]_  | ~\wb_data_i[25] ;
  assign \new_[8355]_  = ~\new_[9133]_  | ~\wb_data_i[26] ;
  assign \new_[8356]_  = ~\new_[9133]_  | ~\wb_data_i[27] ;
  assign \new_[8357]_  = ~\new_[9068]_  | ~\wb_data_i[28] ;
  assign \new_[8358]_  = ~\new_[9090]_  & (~\new_[14636]_  | ~\new_[2344]_ );
  assign \new_[8359]_  = ~\new_[9132]_  | ~\wb_data_i[29] ;
  assign \new_[8360]_  = ~\new_[9134]_  | ~\wb_data_i[2] ;
  assign \new_[8361]_  = ~\new_[9132]_  | ~\wb_data_i[30] ;
  assign \new_[8362]_  = ~\new_[9134]_  | ~\wb_data_i[31] ;
  assign \new_[8363]_  = ~\new_[9067]_  | ~\wb_data_i[3] ;
  assign \new_[8364]_  = ~\new_[9133]_  | ~\wb_data_i[4] ;
  assign \new_[8365]_  = ~\new_[9133]_  | ~\wb_data_i[5] ;
  assign \new_[8366]_  = ~\new_[9646]_  | (~\new_[9420]_  & ~\new_[3882]_ );
  assign \new_[8367]_  = ~\new_[9067]_  | ~\wb_data_i[6] ;
  assign \new_[8368]_  = ~\new_[9067]_  | ~\wb_data_i[7] ;
  assign \new_[8369]_  = ~\new_[9068]_  | ~\wb_data_i[8] ;
  assign \new_[8370]_  = ~\new_[9134]_  | ~\wb_data_i[9] ;
  assign \new_[8371]_  = ~\new_[9091]_  & (~\new_[14636]_  | ~\new_[2345]_ );
  assign \new_[8372]_  = ~\new_[9143]_  | ~\wb_data_i[1] ;
  assign \new_[8373]_  = ~\new_[9143]_  | ~\wb_data_i[12] ;
  assign \new_[8374]_  = ~\new_[9047]_  | ~\wb_data_i[0] ;
  assign \new_[8375]_  = ~\new_[9047]_  | ~\wb_data_i[10] ;
  assign \new_[8376]_  = ~\new_[9047]_  | ~\wb_data_i[11] ;
  assign \new_[8377]_  = ~\new_[9047]_  | ~\wb_data_i[12] ;
  assign \new_[8378]_  = ~\new_[9047]_  | ~\wb_data_i[1] ;
  assign \new_[8379]_  = ~\new_[9093]_  & (~\new_[14636]_  | ~\new_[2347]_ );
  assign \new_[8380]_  = ~\new_[9047]_  | ~\wb_data_i[3] ;
  assign \new_[8381]_  = ~\new_[9047]_  | ~\wb_data_i[5] ;
  assign \new_[8382]_  = ~\new_[9047]_  | ~\wb_data_i[6] ;
  assign \new_[8383]_  = ~\new_[9047]_  | ~\wb_data_i[7] ;
  assign \new_[8384]_  = ~\new_[9047]_  | ~\wb_data_i[8] ;
  assign \new_[8385]_  = ~\new_[9047]_  | ~\wb_data_i[9] ;
  assign \new_[8386]_  = ~\new_[9047]_  | ~\wb_data_i[15] ;
  assign \new_[8387]_  = ~\new_[9047]_  | ~\wb_data_i[25] ;
  assign \new_[8388]_  = ~\new_[9047]_  | ~\wb_data_i[26] ;
  assign \new_[8389]_  = ~\new_[9047]_  | ~\wb_data_i[27] ;
  assign \new_[8390]_  = ~\new_[9047]_  | ~\wb_data_i[19] ;
  assign \new_[8391]_  = ~\new_[9047]_  | ~\wb_data_i[20] ;
  assign \new_[8392]_  = ~\new_[9047]_  | ~\wb_data_i[21] ;
  assign \new_[8393]_  = ~\new_[9047]_  | ~\wb_data_i[24] ;
  assign \new_[8394]_  = ~\new_[9143]_  | ~\wb_data_i[10] ;
  assign \new_[8395]_  = ~\new_[9411]_  | (~\new_[9417]_  & ~\new_[3476]_ );
  assign \new_[8396]_  = ~\new_[9144]_  | ~\wb_data_i[13] ;
  assign \new_[8397]_  = ~\new_[13518]_  | ~\new_[9425]_ ;
  assign \new_[8398]_  = ~\new_[9112]_  | (~\new_[9418]_  & ~\new_[3638]_ );
  assign \new_[8399]_  = ~\new_[9047]_  | ~\wb_data_i[13] ;
  assign \new_[8400]_  = ~\new_[9128]_  | ~\new_[6853]_ ;
  assign \new_[8401]_  = ~\new_[14008]_  | ~\new_[9425]_ ;
  assign \new_[8402]_  = ~\new_[13515]_  | ~\new_[9425]_ ;
  assign \new_[8403]_  = ~\new_[9092]_  & (~\new_[14636]_  | ~\new_[2346]_ );
  assign \new_[8404]_  = ~\new_[9143]_  | ~\wb_data_i[24] ;
  assign \new_[8405]_  = ~\new_[9144]_  | ~\wb_data_i[18] ;
  assign \new_[8406]_  = ~\new_[9144]_  | ~\wb_data_i[3] ;
  assign \new_[8407]_  = ~\new_[9143]_  | ~\wb_data_i[5] ;
  assign \new_[8408]_  = ~\new_[9144]_  | ~\wb_data_i[27] ;
  assign \new_[8409]_  = ~\new_[9143]_  | ~\wb_data_i[16] ;
  assign \new_[8410]_  = ~\new_[9143]_  | ~\wb_data_i[17] ;
  assign \new_[8411]_  = ~\new_[9144]_  | ~\wb_data_i[19] ;
  assign \new_[8412]_  = ~\new_[9144]_  | ~\wb_data_i[21] ;
  assign \new_[8413]_  = \new_[9160]_  & \new_[9792]_ ;
  assign \new_[8414]_  = ~\new_[13696]_  | ~\new_[9425]_ ;
  assign \new_[8415]_  = ~\new_[9128]_  | ~\new_[6733]_ ;
  assign \new_[8416]_  = ~\new_[14548]_  | ~\new_[2471]_ ;
  assign \new_[8417]_  = \new_[14548]_  | \new_[2471]_ ;
  assign \new_[8418]_  = ~\new_[9131]_  | ~\wb_data_i[26] ;
  assign \new_[8419]_  = ~\new_[9129]_  | ~\wb_data_i[23] ;
  assign \new_[8420]_  = ~\new_[9129]_  | ~\wb_data_i[20] ;
  assign \new_[8421]_  = ~\new_[9130]_  | ~\wb_data_i[11] ;
  assign \new_[8422]_  = ~\new_[9129]_  | ~\wb_data_i[13] ;
  assign \new_[8423]_  = ~\new_[9129]_  | ~\wb_data_i[14] ;
  assign \new_[8424]_  = ~\new_[9130]_  | ~\wb_data_i[15] ;
  assign \new_[8425]_  = ~\new_[9129]_  | ~\wb_data_i[16] ;
  assign \new_[8426]_  = ~\new_[9129]_  | ~\wb_data_i[18] ;
  assign \new_[8427]_  = ~\new_[9130]_  | ~\wb_data_i[0] ;
  assign \new_[8428]_  = ~\new_[9156]_  | ~\wb_data_i[30] ;
  assign \new_[8429]_  = ~\new_[9082]_  | ~\wb_data_i[27] ;
  assign \new_[8430]_  = ~\new_[9129]_  | ~\wb_data_i[29] ;
  assign \new_[8431]_  = ~\new_[9082]_  | ~\wb_data_i[2] ;
  assign \new_[8432]_  = ~\new_[9139]_  | ~\wb_data_i[13] ;
  assign \new_[8433]_  = ~\new_[9082]_  | ~\wb_data_i[4] ;
  assign \new_[8434]_  = ~\new_[9129]_  | ~\wb_data_i[9] ;
  assign \new_[8435]_  = ~\new_[9129]_  | ~\wb_data_i[17] ;
  assign \new_[8436]_  = ~\new_[9158]_  | ~\wb_data_i[27] ;
  assign \new_[8437]_  = ~\new_[9082]_  | ~\wb_data_i[7] ;
  assign \new_[8438]_  = ~\new_[9156]_  | ~\wb_data_i[21] ;
  assign \new_[8439]_  = ~\new_[9157]_  | ~\wb_data_i[11] ;
  assign \new_[8440]_  = ~\new_[9127]_  & ~\new_[13413]_ ;
  assign \new_[8441]_  = ~\new_[9131]_  | ~\wb_data_i[0] ;
  assign \new_[8442]_  = ~\new_[9131]_  | ~\wb_data_i[10] ;
  assign \new_[8443]_  = ~\new_[9131]_  | ~\wb_data_i[1] ;
  assign \new_[8444]_  = ~\new_[9131]_  | ~\wb_data_i[2] ;
  assign \new_[8445]_  = ~\new_[9131]_  | ~\wb_data_i[4] ;
  assign \new_[8446]_  = ~\new_[9131]_  | ~\wb_data_i[5] ;
  assign \new_[8447]_  = ~\new_[9131]_  | ~\wb_data_i[6] ;
  assign \new_[8448]_  = ~\new_[9131]_  | ~\wb_data_i[9] ;
  assign \new_[8449]_  = ~\new_[9131]_  | ~\wb_data_i[25] ;
  assign \new_[8450]_  = ~\new_[9131]_  | ~\wb_data_i[16] ;
  assign \new_[8451]_  = ~\new_[9131]_  | ~\wb_data_i[19] ;
  assign \new_[8452]_  = ~\new_[9131]_  | ~\wb_data_i[20] ;
  assign \new_[8453]_  = ~\new_[8780]_ ;
  assign \new_[8454]_  = ~\new_[9131]_  | ~\wb_data_i[24] ;
  assign \new_[8455]_  = ~\new_[9130]_  | ~\wb_data_i[10] ;
  assign \new_[8456]_  = ~\new_[9129]_  | ~\wb_data_i[6] ;
  assign \new_[8457]_  = ~\new_[9101]_  | ~\wb_data_i[25] ;
  assign \new_[8458]_  = ~\new_[9130]_  | ~\wb_data_i[22] ;
  assign \new_[8459]_  = ~\new_[9131]_  | ~\wb_data_i[18] ;
  assign \new_[8460]_  = ~\new_[9131]_  | ~\wb_data_i[13] ;
  assign \new_[8461]_  = ~\new_[9131]_  | ~\wb_data_i[3] ;
  assign \new_[8462]_  = ~\new_[9082]_  | ~\wb_data_i[31] ;
  assign \new_[8463]_  = ~\new_[9139]_  | ~\wb_data_i[25] ;
  assign \new_[8464]_  = ~\new_[9136]_  | ~\wb_data_i[18] ;
  assign \new_[8465]_  = ~\new_[9156]_  | ~\wb_data_i[17] ;
  assign \new_[8466]_  = ~\new_[9139]_  | ~\wb_data_i[24] ;
  assign \new_[8467]_  = ~\new_[9136]_  | ~\wb_data_i[27] ;
  assign \new_[8468]_  = ~\new_[9131]_  | ~\wb_data_i[27] ;
  assign \new_[8469]_  = ~\new_[9509]_  | ~\new_[10574]_  | ~\new_[11643]_  | ~\new_[10489]_ ;
  assign \new_[8470]_  = ~\new_[9048]_  | ~\wb_data_i[6] ;
  assign \new_[8471]_  = ~\new_[9101]_  | ~\wb_data_i[16] ;
  assign \new_[8472]_  = ~\new_[9157]_  | ~\wb_data_i[15] ;
  assign \new_[8473]_  = ~\new_[8803]_ ;
  assign \new_[8474]_  = ~\new_[9129]_  | ~\wb_data_i[24] ;
  assign \new_[8475]_  = ~\new_[9130]_  | ~\wb_data_i[25] ;
  assign \new_[8476]_  = ~\new_[14637]_  & ~\new_[9084]_ ;
  assign \new_[8477]_  = ~\new_[9129]_  | ~\wb_data_i[21] ;
  assign \new_[8478]_  = ~\new_[9129]_  | ~\wb_data_i[5] ;
  assign \new_[8479]_  = ~\new_[9131]_  | ~\wb_data_i[15] ;
  assign \new_[8480]_  = ~\new_[9131]_  | ~\wb_data_i[12] ;
  assign \new_[8481]_  = ~\new_[9139]_  | ~\wb_data_i[23] ;
  assign \new_[8482]_  = ~\new_[9139]_  | ~\wb_data_i[5] ;
  assign \new_[8483]_  = ~\new_[9131]_  | ~\wb_data_i[11] ;
  assign \new_[8484]_  = ~\new_[9131]_  | ~\wb_data_i[21] ;
  assign \new_[8485]_  = ~\new_[9082]_  | ~\wb_data_i[12] ;
  assign \new_[8486]_  = ~\new_[9158]_  | ~\wb_data_i[26] ;
  assign \new_[8487]_  = ~\new_[9124]_  & ~\new_[13350]_ ;
  assign \new_[8488]_  = ~\new_[9129]_  | ~\wb_data_i[30] ;
  assign \new_[8489]_  = ~\new_[9139]_  | ~\wb_data_i[22] ;
  assign \new_[8490]_  = ~\new_[9131]_  | ~\wb_data_i[7] ;
  assign \new_[8491]_  = ~\new_[9130]_  | ~\wb_data_i[3] ;
  assign \new_[8492]_  = ~\new_[9129]_  | ~\wb_data_i[26] ;
  assign \new_[8493]_  = ~\new_[9139]_  | ~\wb_data_i[0] ;
  assign \new_[8494]_  = ~\new_[9139]_  | ~\wb_data_i[11] ;
  assign \new_[8495]_  = ~\new_[9139]_  | ~\wb_data_i[12] ;
  assign \new_[8496]_  = ~\new_[9139]_  | ~\wb_data_i[15] ;
  assign \new_[8497]_  = ~\new_[9139]_  | ~\wb_data_i[18] ;
  assign \new_[8498]_  = ~\new_[9139]_  | ~\wb_data_i[1] ;
  assign \new_[8499]_  = ~\new_[9131]_  | ~\wb_data_i[17] ;
  assign \new_[8500]_  = ~\new_[9139]_  | ~\wb_data_i[27] ;
  assign \new_[8501]_  = ~\new_[9139]_  | ~\wb_data_i[28] ;
  assign \new_[8502]_  = ~\new_[9139]_  | ~\wb_data_i[2] ;
  assign \new_[8503]_  = ~\new_[9139]_  | ~\wb_data_i[3] ;
  assign \new_[8504]_  = ~\new_[9139]_  | ~\wb_data_i[4] ;
  assign \new_[8505]_  = ~\new_[9139]_  | ~\wb_data_i[6] ;
  assign n7610 = ~\new_[12804]_  & (~\new_[9199]_  | ~\new_[9939]_ );
  assign \new_[8507]_  = ~\new_[9139]_  | ~\wb_data_i[7] ;
  assign \new_[8508]_  = ~\new_[9139]_  | ~\wb_data_i[8] ;
  assign \new_[8509]_  = ~\new_[9131]_  | ~\wb_data_i[8] ;
  assign \new_[8510]_  = ~\new_[9139]_  | ~\wb_data_i[9] ;
  assign \new_[8511]_  = ~\new_[9156]_  | ~\wb_data_i[20] ;
  assign \new_[8512]_  = ~\new_[9434]_  | ~\wb_data_i[30] ;
  assign \new_[8513]_  = ~\new_[9048]_  | ~\wb_data_i[0] ;
  assign \new_[8514]_  = ~\new_[9048]_  | ~\wb_data_i[10] ;
  assign \new_[8515]_  = ~\new_[9048]_  | ~\wb_data_i[11] ;
  assign \new_[8516]_  = ~\new_[9136]_  | ~\wb_data_i[3] ;
  assign \new_[8517]_  = ~\new_[9048]_  | ~\wb_data_i[4] ;
  assign \new_[8518]_  = ~\new_[9048]_  | ~\wb_data_i[8] ;
  assign \new_[8519]_  = ~\new_[9136]_  | ~\wb_data_i[15] ;
  assign \new_[8520]_  = ~\new_[9136]_  | ~\wb_data_i[26] ;
  assign \new_[8521]_  = ~\new_[9048]_  | ~\wb_data_i[16] ;
  assign \new_[8522]_  = ~\new_[9136]_  | ~\wb_data_i[20] ;
  assign \new_[8523]_  = ~\new_[9654]_  | ~\new_[2339]_  | ~\new_[11595]_  | ~\new_[12277]_ ;
  assign \new_[8524]_  = ~\new_[9136]_  | ~\wb_data_i[21] ;
  assign \new_[8525]_  = ~\new_[8829]_ ;
  assign \new_[8526]_  = ~\new_[9048]_  | ~\wb_data_i[24] ;
  assign \new_[8527]_  = ~\new_[8830]_ ;
  assign \new_[8528]_  = ~\new_[9130]_  | ~\wb_data_i[1] ;
  assign \new_[8529]_  = ~\new_[9101]_  | ~\wb_data_i[23] ;
  assign \new_[8530]_  = ~\new_[9082]_  | ~\wb_data_i[8] ;
  assign \new_[8531]_  = ~\new_[9156]_  | ~\wb_data_i[22] ;
  assign \new_[8532]_  = ~\new_[9156]_  | ~\wb_data_i[18] ;
  assign \new_[8533]_  = ~\new_[9226]_  & (~\new_[10123]_  | ~\new_[9480]_ );
  assign \new_[8534]_  = ~\new_[9136]_  | ~\wb_data_i[13] ;
  assign \new_[8535]_  = ~\new_[9101]_  | ~\wb_data_i[0] ;
  assign \new_[8536]_  = ~\new_[9156]_  | ~\wb_data_i[10] ;
  assign \new_[8537]_  = ~\new_[9156]_  | ~\wb_data_i[12] ;
  assign \new_[8538]_  = ~\new_[9156]_  | ~\wb_data_i[13] ;
  assign \new_[8539]_  = ~\new_[9157]_  | ~\wb_data_i[14] ;
  assign \new_[8540]_  = ~\new_[9139]_  | ~\wb_data_i[21] ;
  assign \new_[8541]_  = ~\new_[9101]_  | ~\wb_data_i[19] ;
  assign \new_[8542]_  = ~\new_[9156]_  | ~\wb_data_i[1] ;
  assign \new_[8543]_  = ~\new_[9101]_  | ~\wb_data_i[24] ;
  assign \new_[8544]_  = ~\new_[9156]_  | ~\wb_data_i[29] ;
  assign \new_[8545]_  = ~\new_[9157]_  | ~\wb_data_i[2] ;
  assign \new_[8546]_  = ~\new_[9158]_  | ~\wb_data_i[31] ;
  assign \new_[8547]_  = ~\new_[9101]_  | ~\wb_data_i[5] ;
  assign \new_[8548]_  = ~\new_[9156]_  | ~\wb_data_i[6] ;
  assign \new_[8549]_  = ~\new_[9101]_  | ~\wb_data_i[9] ;
  assign \new_[8550]_  = ~\new_[9129]_  | ~\wb_data_i[19] ;
  assign n7605 = \new_[6012]_  ^ \new_[9338]_ ;
  assign \new_[8552]_  = ~\new_[9158]_  | ~\wb_data_i[4] ;
  assign \new_[8553]_  = ~\new_[9157]_  | ~\wb_data_i[8] ;
  assign \new_[8554]_  = ~\new_[9082]_  | ~\wb_data_i[28] ;
  assign \new_[8555]_  = ~\new_[9157]_  | ~\wb_data_i[7] ;
  assign \new_[8556]_  = ~\new_[9157]_  | ~\wb_data_i[3] ;
  assign \new_[8557]_  = ~\new_[9157]_  | ~\wb_data_i[28] ;
  assign \new_[8558]_  = ~\new_[8845]_ ;
  assign \new_[8559]_  = ~\new_[5766]_  | ~\new_[8970]_ ;
  assign \new_[8560]_  = ~\new_[12830]_  & (~\new_[9485]_  | ~\new_[11199]_ );
  assign n7620 = ~\new_[11958]_  & ~\new_[9150]_ ;
  assign \new_[8562]_  = ~\new_[11603]_  & (~\new_[9782]_  | ~\new_[10007]_ );
  assign \new_[8563]_  = ~\new_[12656]_  & (~\new_[9489]_  | ~\new_[11197]_ );
  assign \new_[8564]_  = ~\new_[9106]_ ;
  assign \new_[8565]_  = ~\new_[12754]_  & (~\new_[9198]_  | ~\new_[11209]_ );
  assign \new_[8566]_  = ~\new_[10479]_  | ~\new_[12960]_  | ~\new_[9479]_ ;
  assign \new_[8567]_  = ~\new_[12668]_  & (~\new_[9486]_  | ~\new_[11195]_ );
  assign \new_[8568]_  = ~\new_[10125]_  | (~\new_[9477]_  & ~\new_[9804]_ );
  assign \new_[8569]_  = ~\new_[9578]_  | ~\new_[10013]_  | ~\new_[11014]_  | ~\new_[10353]_ ;
  assign \new_[8570]_  = ~\new_[9169]_  | (~\new_[10612]_  & ~\new_[10394]_ );
  assign \new_[8571]_  = ~\new_[9168]_  | (~\new_[10436]_  & ~\new_[10387]_ );
  assign \new_[8572]_  = ~\new_[9170]_  | (~\new_[10437]_  & ~\new_[10397]_ );
  assign \new_[8573]_  = ~\new_[9171]_  | (~\new_[10450]_  & ~\new_[10404]_ );
  assign \new_[8574]_  = ~\new_[8856]_ ;
  assign \new_[8575]_  = ~\new_[8858]_ ;
  assign \new_[8576]_  = ~n7975 | (~\new_[9211]_  & ~\new_[6850]_ );
  assign \new_[8577]_  = ~\new_[8861]_ ;
  assign \new_[8578]_  = ~\new_[9213]_  & ~\new_[9189]_ ;
  assign \new_[8579]_  = ~\new_[9014]_  & (~\new_[10731]_  | ~\new_[10475]_ );
  assign \new_[8580]_  = ~\new_[8990]_  & (~\new_[10732]_  | ~\new_[10475]_ );
  assign \new_[8581]_  = ~\new_[8676]_ ;
  assign \new_[8582]_  = ~\new_[8989]_  & (~\new_[10729]_  | ~\new_[10475]_ );
  assign \new_[8583]_  = ~\new_[9140]_ ;
  assign \new_[8584]_  = ~\new_[9016]_  & (~\new_[10730]_  | ~\new_[10475]_ );
  assign \new_[8585]_  = ~\new_[9002]_  & (~\new_[10050]_  | ~\new_[10475]_ );
  assign \new_[8586]_  = ~\new_[9192]_  | (~\new_[11098]_  & ~\new_[11149]_ );
  assign \new_[8587]_  = ~\new_[8995]_  & (~\new_[10734]_  | ~\new_[10475]_ );
  assign \new_[8588]_  = ~\new_[10496]_  | ~\new_[9523]_  | ~\new_[9213]_ ;
  assign \new_[8589]_  = ~\new_[9000]_  & (~\new_[10031]_  | ~\new_[10475]_ );
  assign \new_[8590]_  = ~\new_[9235]_  & (~\new_[9309]_  | ~\new_[10839]_ );
  assign \new_[8591]_  = ~\new_[8974]_  | (~\new_[9225]_  & ~\new_[11698]_ );
  assign \new_[8592]_  = ~\new_[11944]_  | ~\new_[12797]_  | ~\new_[9523]_  | ~\new_[11649]_ ;
  assign \new_[8593]_  = \new_[9360]_  ? \new_[9857]_  : \new_[2095]_ ;
  assign \new_[8594]_  = ~\new_[9189]_  & ~\new_[12588]_ ;
  assign \new_[8595]_  = \new_[2340]_  ^ \new_[9373]_ ;
  assign \new_[8596]_  = ~\new_[10270]_  | ~\new_[13481]_  | ~\new_[9501]_  | ~\new_[9506]_ ;
  assign \new_[8597]_  = ~\new_[13466]_  & (~\new_[9417]_  | ~\new_[3480]_ );
  assign \new_[8598]_  = (~\new_[9413]_  | ~\new_[3505]_ ) & (~\new_[9366]_  | ~\new_[3504]_ );
  assign \new_[8599]_  = ~\new_[14330]_ ;
  assign \new_[8600]_  = ~\new_[8927]_ ;
  assign \new_[8601]_  = \new_[14587]_ ;
  assign \new_[8602]_  = \new_[14423]_ ;
  assign \new_[8603]_  = ~\new_[14451]_ ;
  assign \new_[8604]_  = ~\new_[8631]_ ;
  assign \new_[8605]_  = \new_[14389]_  ^ \new_[9213]_ ;
  assign \new_[8606]_  = ~\new_[13351]_  & (~\new_[9420]_  | ~\new_[3884]_ );
  assign \new_[8607]_  = ~\new_[9018]_  & (~\new_[11954]_  | ~\new_[10086]_ );
  assign \new_[8608]_  = ~\new_[9611]_  | ~\new_[8970]_ ;
  assign \new_[8609]_  = ~\new_[6023]_  | ~\new_[8970]_ ;
  assign \new_[8610]_  = \new_[9806]_  | \new_[9032]_ ;
  assign \new_[8611]_  = ~\new_[9502]_  & (~\new_[9314]_  | ~\new_[10835]_ );
  assign \new_[8612]_  = ~\new_[9514]_  & (~\new_[9332]_  | ~\new_[10835]_ );
  assign \new_[8613]_  = ~\new_[9504]_  & (~\new_[9324]_  | ~\new_[10835]_ );
  assign \new_[8614]_  = ~\new_[8941]_ ;
  assign \new_[8615]_  = ~\new_[8993]_  & (~\new_[9732]_  | ~\new_[10839]_ );
  assign \new_[8616]_  = ~\new_[9270]_  & (~\new_[9473]_  | ~\new_[10839]_ );
  assign n9130 = u0_u0_usb_attached_reg;
  assign \new_[8618]_  = ~\new_[13370]_  | ~\new_[8970]_ ;
  assign \new_[8619]_  = ~\new_[10642]_  | ~\new_[8970]_ ;
  assign \new_[8620]_  = \new_[9275]_  | \new_[8976]_ ;
  assign \new_[8621]_  = \new_[8973]_  | \new_[9808]_ ;
  assign \new_[8622]_  = ~n7795 | ~\new_[9824]_  | ~\new_[9836]_ ;
  assign \new_[8623]_  = ~\new_[8964]_ ;
  assign \new_[8624]_  = \new_[12096]_  | \new_[14643]_ ;
  assign \new_[8625]_  = ~\new_[8965]_ ;
  assign \new_[8626]_  = u1_u3_in_token_reg;
  assign \new_[8627]_  = ~\new_[12812]_  | ~\new_[8970]_ ;
  assign \new_[8628]_  = ~\new_[9232]_  & (~\new_[11148]_  | ~\new_[11649]_ );
  assign \new_[8629]_  = ~\new_[9310]_  & (~\new_[4818]_  | ~\new_[14453]_ );
  assign \new_[8630]_  = ~\new_[9231]_  | (~\new_[9884]_  & ~\new_[9857]_ );
  assign \new_[8631]_  = \new_[9230]_  & \new_[9219]_ ;
  assign \new_[8632]_  = \new_[2090]_  ^ \new_[9576]_ ;
  assign \new_[8633]_  = u4_u2_ep_match_r_reg;
  assign \new_[8634]_  = ~\new_[8972]_ ;
  assign \new_[8635]_  = ~\new_[14643]_ ;
  assign \new_[8636]_  = ~\new_[9596]_  | ~\new_[9313]_ ;
  assign \new_[8637]_  = ~\new_[9602]_  | ~\new_[9313]_ ;
  assign \new_[8638]_  = ~\new_[14642]_ ;
  assign \new_[8639]_  = ~\new_[9857]_  | ~\new_[2085]_ ;
  assign \new_[8640]_  = ~\new_[8976]_ ;
  assign \new_[8641]_  = ~\new_[8977]_ ;
  assign \new_[8642]_  = ~\new_[8980]_ ;
  assign \new_[8643]_  = ~\new_[9357]_  | ~\new_[10839]_ ;
  assign \new_[8644]_  = ~\new_[9003]_ ;
  assign \new_[8645]_  = ~\new_[9351]_  | ~\new_[10839]_ ;
  assign \new_[8646]_  = ~\new_[9376]_  & ~\new_[9894]_ ;
  assign \new_[8647]_  = ~\new_[9333]_  & ~\new_[9897]_ ;
  assign \new_[8648]_  = \new_[9602]_  ? \new_[10125]_  : \new_[3881]_ ;
  assign \new_[8649]_  = ~\new_[9327]_  & (~\new_[4091]_  | ~\new_[10125]_ );
  assign \new_[8650]_  = \new_[9596]_  ? \new_[10125]_  : \new_[4092]_ ;
  assign \new_[8651]_  = ~\new_[10296]_  | ~\new_[9391]_ ;
  assign \new_[8652]_  = ~\new_[14409]_  | ~\new_[4794]_ ;
  assign \new_[8653]_  = \new_[9367]_  | \new_[6196]_ ;
  assign \new_[8654]_  = ~\new_[9955]_  | ~\new_[4091]_ ;
  assign \new_[8655]_  = \new_[9368]_  | \new_[6567]_ ;
  assign \new_[8656]_  = ~\new_[9366]_  | ~\new_[3505]_ ;
  assign \new_[8657]_  = ~\new_[9955]_  | ~\new_[3881]_ ;
  assign \new_[8658]_  = \\u1_u3_tx_data_to_cnt_reg[4] ;
  assign \new_[8659]_  = \new_[9369]_  | \new_[6275]_ ;
  assign \new_[8660]_  = \new_[9370]_  | \new_[6287]_ ;
  assign \new_[8661]_  = ~\new_[9358]_  | ~n7980;
  assign \new_[8662]_  = ~\new_[11207]_  & (~\new_[9690]_  | ~\new_[12128]_ );
  assign \new_[8663]_  = ~\new_[11211]_  & (~\new_[9693]_  | ~\new_[11966]_ );
  assign \new_[8664]_  = ~\new_[9033]_ ;
  assign \new_[8665]_  = ~\new_[9034]_ ;
  assign \new_[8666]_  = ~\new_[9413]_  | ~\new_[9366]_ ;
  assign \new_[8667]_  = ~\new_[13494]_  | ~\new_[9363]_  | ~\new_[12353]_ ;
  assign \new_[8668]_  = ~\new_[9217]_  | (~\new_[11396]_  & ~\new_[9857]_ );
  assign n7730 = \new_[12120]_  ^ \new_[9624]_ ;
  assign n7710 = \new_[11987]_  ^ \new_[9617]_ ;
  assign \new_[8671]_  = ~\new_[10298]_  | ~\new_[9394]_ ;
  assign \new_[8672]_  = ~\new_[10297]_  | ~\new_[9390]_ ;
  assign n7715 = \new_[11981]_  ^ \new_[9619]_ ;
  assign n7720 = \new_[12025]_  ^ \new_[9622]_ ;
  assign \new_[8675]_  = \new_[13666]_  ? \new_[10715]_  : \new_[9635]_ ;
  assign \new_[8676]_  = ~\new_[13268]_  & (~\new_[9651]_  | ~\new_[4291]_ );
  assign \new_[8677]_  = \new_[4069]_  ^ \new_[9661]_ ;
  assign \new_[8678]_  = \new_[3312]_  ^ \new_[9668]_ ;
  assign \new_[8679]_  = ~\new_[9216]_  | (~\new_[9967]_  & ~\new_[9857]_ );
  assign \new_[8680]_  = ~\new_[9223]_  | (~\new_[9968]_  & ~\new_[9857]_ );
  assign \new_[8681]_  = \new_[3467]_  ^ \new_[9672]_ ;
  assign \new_[8682]_  = \new_[3687]_  ^ \new_[9512]_ ;
  assign \new_[8683]_  = ~\new_[9214]_  | (~\new_[10121]_  & ~\new_[9857]_ );
  assign \new_[8684]_  = ~\new_[11204]_  & (~\new_[9684]_  | ~\new_[11974]_ );
  assign \new_[8685]_  = ~\new_[11568]_  & (~\new_[9688]_  | ~\new_[12323]_ );
  assign \new_[8686]_  = ~\new_[11565]_  & (~\new_[9691]_  | ~\new_[12321]_ );
  assign \new_[8687]_  = ~\new_[11564]_  & (~\new_[9692]_  | ~\new_[12199]_ );
  assign \new_[8688]_  = \new_[2317]_  ^ \new_[9663]_ ;
  assign \new_[8689]_  = (~\new_[9704]_  | ~\new_[11727]_ ) & (~\new_[13315]_  | ~\new_[3475]_ );
  assign \new_[8690]_  = \new_[9401]_  & \new_[9805]_ ;
  assign \new_[8691]_  = ~\\u4_u0_buf0_orig_m3_reg[7] ;
  assign \new_[8692]_  = ~\new_[10997]_  | ~\new_[9403]_  | ~\new_[10430]_ ;
  assign \new_[8693]_  = ~\\u4_u0_buf0_orig_m3_reg[8] ;
  assign \new_[8694]_  = \new_[9404]_  & \new_[9899]_ ;
  assign \new_[8695]_  = ~\new_[11826]_  & (~\new_[9698]_  | ~\new_[12857]_ );
  assign \new_[8696]_  = ~\new_[11828]_  & (~\new_[9699]_  | ~\new_[12620]_ );
  assign \new_[8697]_  = ~\new_[11830]_  & (~\new_[9700]_  | ~\new_[12563]_ );
  assign \new_[8698]_  = ~\new_[11832]_  & (~\new_[9701]_  | ~\new_[12615]_ );
  assign \new_[8699]_  = ~\new_[10295]_  | ~\new_[9393]_ ;
  assign \new_[8700]_  = \\u1_u3_tx_data_to_cnt_reg[6] ;
  assign \new_[8701]_  = \\u1_u3_tx_data_to_cnt_reg[2] ;
  assign \new_[8702]_  = \\u1_u3_tx_data_to_cnt_reg[1] ;
  assign \new_[8703]_  = \\u1_u3_tx_data_to_cnt_reg[0] ;
  assign n7665 = \new_[12119]_  ^ \new_[9697]_ ;
  assign \new_[8705]_  = \new_[12435]_  ^ \new_[9680]_ ;
  assign \new_[8706]_  = \new_[12008]_  ^ \new_[9702]_ ;
  assign \new_[8707]_  = \new_[11951]_  ^ \new_[9657]_ ;
  assign n7655 = \new_[12007]_  ^ \new_[9694]_ ;
  assign \new_[8709]_  = \new_[12159]_  ^ \new_[9658]_ ;
  assign \new_[8710]_  = \new_[12006]_  ^ \new_[9703]_ ;
  assign \new_[8711]_  = \new_[12226]_  ^ \new_[9681]_ ;
  assign \new_[8712]_  = \new_[11920]_  ^ \new_[9659]_ ;
  assign n7660 = \new_[12388]_  ^ \new_[9695]_ ;
  assign \new_[8714]_  = \new_[11960]_  ^ \new_[9682]_ ;
  assign \new_[8715]_  = \new_[12187]_  ^ \new_[9660]_ ;
  assign \new_[8716]_  = \new_[12389]_  ^ \new_[9683]_ ;
  assign \new_[8717]_  = ~\\u4_u3_buf0_orig_m3_reg[9] ;
  assign \new_[8718]_  = ~\\u4_u1_buf0_orig_m3_reg[9] ;
  assign \new_[8719]_  = ~\\u4_u3_buf0_orig_m3_reg[10] ;
  assign \new_[8720]_  = \new_[2339]_  ^ \new_[14637]_ ;
  assign \new_[8721]_  = \new_[9441]_  | \new_[7297]_ ;
  assign \new_[8722]_  = \new_[9441]_  | \new_[6868]_ ;
  assign \new_[8723]_  = \new_[9441]_  | \new_[7258]_ ;
  assign \new_[8724]_  = \new_[9444]_  | \new_[6866]_ ;
  assign \new_[8725]_  = \new_[9444]_  | \new_[7154]_ ;
  assign \new_[8726]_  = \new_[9444]_  | \new_[7155]_ ;
  assign \new_[8727]_  = \new_[9444]_  | \new_[6863]_ ;
  assign \new_[8728]_  = \new_[9444]_  | \new_[6871]_ ;
  assign \new_[8729]_  = \new_[9444]_  | \new_[6867]_ ;
  assign \new_[8730]_  = \new_[9444]_  | \new_[6862]_ ;
  assign \new_[8731]_  = ~\new_[9644]_  | (~\new_[9651]_  & ~\new_[4288]_ );
  assign \new_[8732]_  = \new_[9444]_  | \new_[6872]_ ;
  assign \new_[8733]_  = \new_[9444]_  | \new_[6873]_ ;
  assign \new_[8734]_  = \new_[9449]_  & \new_[9784]_ ;
  assign \new_[8735]_  = ~\new_[9432]_  | ~\wb_data_i[24] ;
  assign \new_[8736]_  = ~\new_[9432]_  | ~\wb_data_i[25] ;
  assign \new_[8737]_  = ~\new_[9432]_  | ~\wb_data_i[26] ;
  assign \new_[8738]_  = ~\new_[9432]_  | ~\wb_data_i[27] ;
  assign \new_[8739]_  = ~\new_[9432]_  | ~\wb_data_i[28] ;
  assign \new_[8740]_  = ~\new_[9432]_  | ~\wb_data_i[29] ;
  assign \new_[8741]_  = ~\new_[9432]_  | ~\wb_data_i[16] ;
  assign \new_[8742]_  = ~\new_[9432]_  | ~\wb_data_i[17] ;
  assign \new_[8743]_  = ~\new_[9432]_  | ~\wb_data_i[18] ;
  assign \new_[8744]_  = ~\new_[9432]_  | ~\wb_data_i[19] ;
  assign \new_[8745]_  = ~\new_[9432]_  | ~\wb_data_i[20] ;
  assign \new_[8746]_  = ~\new_[9432]_  | ~\wb_data_i[21] ;
  assign \new_[8747]_  = \new_[9444]_  | \new_[6870]_ ;
  assign \new_[8748]_  = \new_[9444]_  | \new_[6869]_ ;
  assign \new_[8749]_  = \new_[9450]_  & \new_[9796]_ ;
  assign \new_[8750]_  = \new_[9441]_  | \new_[6875]_ ;
  assign \new_[8751]_  = \new_[9441]_  | \new_[6880]_ ;
  assign \new_[8752]_  = \new_[9441]_  | \new_[7163]_ ;
  assign \new_[8753]_  = \new_[9441]_  | \new_[6882]_ ;
  assign \new_[8754]_  = \new_[9441]_  | \new_[6865]_ ;
  assign \new_[8755]_  = \new_[9441]_  | \new_[7179]_ ;
  assign \new_[8756]_  = \new_[9441]_  | \new_[7301]_ ;
  assign \new_[8757]_  = \new_[9441]_  | \new_[7164]_ ;
  assign \new_[8758]_  = \new_[9441]_  | \new_[7302]_ ;
  assign \new_[8759]_  = \new_[9444]_  | \new_[6881]_ ;
  assign \new_[8760]_  = ~\new_[9447]_  | ~\wb_data_i[20] ;
  assign \new_[8761]_  = \new_[9447]_  | \new_[7205]_ ;
  assign \new_[8762]_  = ~\new_[9447]_  | ~\wb_data_i[24] ;
  assign \new_[8763]_  = ~\new_[9447]_  | ~\wb_data_i[25] ;
  assign \new_[8764]_  = \new_[9913]_  ? \new_[14637]_  : \new_[2316]_ ;
  assign \new_[8765]_  = ~\new_[9447]_  | ~\wb_data_i[26] ;
  assign \new_[8766]_  = \new_[9447]_  | \new_[7286]_ ;
  assign \new_[8767]_  = \new_[9447]_  | \new_[7148]_ ;
  assign \new_[8768]_  = \new_[9447]_  | \new_[7291]_ ;
  assign \new_[8769]_  = ~\new_[9447]_  | ~\wb_data_i[29] ;
  assign \new_[8770]_  = \new_[9447]_  | \new_[7150]_ ;
  assign \new_[8771]_  = \new_[9447]_  | \new_[7285]_ ;
  assign \new_[8772]_  = ~\new_[9447]_  | ~\wb_data_i[19] ;
  assign \new_[8773]_  = \new_[9447]_  | \new_[7152]_ ;
  assign \new_[8774]_  = \new_[9447]_  | \new_[7277]_ ;
  assign \new_[8775]_  = \new_[10225]_  ? \new_[14637]_  : \new_[2318]_ ;
  assign \new_[8776]_  = ~\new_[9444]_  | ~\wb_data_i[24] ;
  assign \new_[8777]_  = ~\new_[9444]_  | ~\wb_data_i[20] ;
  assign \new_[8778]_  = ~\new_[9441]_  | ~\wb_data_i[16] ;
  assign \new_[8779]_  = ~\new_[6743]_  | ~\new_[9426]_ ;
  assign \new_[8780]_  = ~\new_[9426]_  | ~\new_[12197]_ ;
  assign \new_[8781]_  = ~\new_[9447]_  | ~\wb_data_i[17] ;
  assign \new_[8782]_  = \new_[9447]_  | \new_[7151]_ ;
  assign \new_[8783]_  = ~\new_[9441]_  | ~\wb_data_i[26] ;
  assign \new_[8784]_  = ~\new_[9447]_  | ~\wb_data_i[21] ;
  assign \new_[8785]_  = ~\new_[9444]_  | ~\wb_data_i[25] ;
  assign \new_[8786]_  = ~\new_[9444]_  | ~\wb_data_i[29] ;
  assign \new_[8787]_  = ~\new_[9444]_  | ~\wb_data_i[18] ;
  assign \new_[8788]_  = ~\new_[9444]_  | ~\wb_data_i[19] ;
  assign \new_[8789]_  = ~\new_[9447]_  | ~\wb_data_i[16] ;
  assign \new_[8790]_  = ~\new_[10786]_  | ~XcvSelect_pad_o | ~\new_[9750]_ ;
  assign \new_[8791]_  = ~\new_[9087]_ ;
  assign \new_[8792]_  = ~\new_[9414]_  & ~\new_[12690]_ ;
  assign \new_[8793]_  = \new_[9447]_  | \new_[7149]_ ;
  assign \new_[8794]_  = ~\new_[3895]_  | ~\new_[12420]_  | ~\new_[10285]_ ;
  assign \new_[8795]_  = ~\new_[3177]_  | ~\new_[12420]_  | ~\new_[10285]_ ;
  assign \new_[8796]_  = ~\new_[9447]_  | ~\wb_data_i[28] ;
  assign \new_[8797]_  = ~\new_[6690]_  | ~\new_[9430]_ ;
  assign \new_[8798]_  = \new_[9447]_  | \new_[7147]_ ;
  assign \new_[8799]_  = ~\new_[9444]_  | ~\wb_data_i[17] ;
  assign \new_[8800]_  = ~\new_[9444]_  | ~\wb_data_i[16] ;
  assign \new_[8801]_  = ~\new_[6809]_  | ~\new_[9445]_ ;
  assign \new_[8802]_  = ~\new_[9447]_  | ~\wb_data_i[27] ;
  assign \new_[8803]_  = ~\new_[9429]_  | ~\new_[12197]_ ;
  assign \new_[8804]_  = \new_[9447]_  | \new_[7153]_ ;
  assign \new_[8805]_  = ~\new_[14637]_  & ~\new_[9396]_ ;
  assign \new_[8806]_  = \new_[9432]_  | \new_[7177]_ ;
  assign \new_[8807]_  = ~\new_[13138]_  | ~\new_[10028]_  | ~\new_[9656]_ ;
  assign \new_[8808]_  = \new_[9432]_  | \new_[7162]_ ;
  assign \new_[8809]_  = u1_u3_buf0_na_reg;
  assign \new_[8810]_  = u1_u3_buf1_na_reg;
  assign \new_[8811]_  = \new_[9432]_  | \new_[7278]_ ;
  assign \new_[8812]_  = \new_[9432]_  | \new_[7156]_ ;
  assign \new_[8813]_  = \new_[9432]_  | \new_[7157]_ ;
  assign \new_[8814]_  = \new_[9432]_  | \new_[7158]_ ;
  assign \new_[8815]_  = \new_[9432]_  | \new_[7200]_ ;
  assign \new_[8816]_  = \new_[9432]_  | \new_[7159]_ ;
  assign \new_[8817]_  = \new_[9432]_  | \new_[7202]_ ;
  assign \new_[8818]_  = \new_[9432]_  | \new_[7160]_ ;
  assign \new_[8819]_  = \new_[9432]_  | \new_[7198]_ ;
  assign \new_[8820]_  = \new_[9432]_  | \new_[7161]_ ;
  assign \new_[8821]_  = \new_[9416]_  | \new_[12756]_ ;
  assign \new_[8822]_  = ~\new_[12688]_  & (~\new_[9656]_  | ~\new_[13494]_ );
  assign \new_[8823]_  = ~\new_[9444]_  | ~\wb_data_i[26] ;
  assign \new_[8824]_  = ~\new_[9441]_  | ~\wb_data_i[20] ;
  assign \new_[8825]_  = ~\new_[9444]_  | ~\wb_data_i[21] ;
  assign \new_[8826]_  = \\u1_u3_tx_data_to_cnt_reg[3] ;
  assign \new_[8827]_  = ~\new_[10087]_  & ~\new_[9219]_ ;
  assign \new_[8828]_  = ~\new_[9444]_  | ~\wb_data_i[27] ;
  assign \new_[8829]_  = ~\new_[9430]_  | ~\new_[12197]_ ;
  assign \new_[8830]_  = ~\new_[9445]_  | ~rst_i;
  assign \new_[8831]_  = ~\new_[9444]_  | ~\wb_data_i[28] ;
  assign \new_[8832]_  = ~\new_[9441]_  | ~\wb_data_i[24] ;
  assign \new_[8833]_  = ~\new_[9441]_  | ~\wb_data_i[25] ;
  assign \new_[8834]_  = ~\new_[9441]_  | ~\wb_data_i[27] ;
  assign \new_[8835]_  = ~\new_[9441]_  | ~\wb_data_i[28] ;
  assign \new_[8836]_  = ~\new_[9441]_  | ~\wb_data_i[29] ;
  assign \new_[8837]_  = ~\new_[9441]_  | ~\wb_data_i[17] ;
  assign \new_[8838]_  = ~\new_[9441]_  | ~\wb_data_i[18] ;
  assign \new_[8839]_  = ~\new_[9441]_  | ~\wb_data_i[19] ;
  assign \new_[8840]_  = ~\new_[9441]_  | ~\wb_data_i[21] ;
  assign \new_[8841]_  = ~\new_[9213]_  & (~\new_[9738]_  | ~\new_[9506]_ );
  assign n7670 = \new_[6326]_  ^ \new_[9566]_ ;
  assign \new_[8843]_  = ~\new_[9447]_  | ~\wb_data_i[18] ;
  assign \new_[8844]_  = \new_[9422]_  | \new_[13464]_ ;
  assign \new_[8845]_  = ~\new_[9835]_  | ~\new_[10002]_  | ~\new_[11011]_  | ~\new_[10712]_ ;
  assign \new_[8846]_  = ~\new_[9258]_  & (~\new_[10344]_  | ~\new_[10475]_ );
  assign \new_[8847]_  = ~\new_[9730]_  | ~\new_[9987]_  | ~\new_[10877]_ ;
  assign \new_[8848]_  = ~\new_[9741]_  | ~\new_[9996]_  | ~\new_[10752]_ ;
  assign \new_[8849]_  = ~\new_[9744]_  | ~\new_[9986]_  | ~\new_[10753]_ ;
  assign \new_[8850]_  = ~\new_[9746]_  | ~\new_[10009]_  | ~\new_[10751]_ ;
  assign \new_[8851]_  = ~\new_[9224]_  | (~\new_[11015]_  & ~\new_[9857]_ );
  assign \new_[8852]_  = ~\new_[9227]_  | (~\new_[11751]_  & ~\new_[9857]_ );
  assign \new_[8853]_  = ~\new_[10010]_  | ~\new_[11077]_  | ~\new_[10425]_  | ~\new_[10802]_ ;
  assign \new_[8854]_  = ~\new_[9125]_ ;
  assign \new_[8855]_  = ~u4_u3_int_re_reg;
  assign \new_[8856]_  = ~\\u4_u0_buf0_orig_m3_reg[6] ;
  assign \new_[8857]_  = ~\new_[9126]_ ;
  assign \new_[8858]_  = ~\\u4_u2_buf0_orig_m3_reg[6] ;
  assign \new_[8859]_  = ~\new_[9966]_  | ~\new_[10702]_  | ~\new_[10704]_  | ~\new_[10705]_ ;
  assign \new_[8860]_  = ~\new_[9129]_ ;
  assign \new_[8861]_  = ~\new_[10786]_  | (~\new_[9513]_  & ~\new_[11335]_ );
  assign \new_[8862]_  = ~\new_[9131]_ ;
  assign \new_[8863]_  = ~\new_[9283]_  & (~\new_[9545]_  | ~\new_[11143]_ );
  assign \new_[8864]_  = ~\new_[9286]_  & (~\new_[9550]_  | ~\new_[11143]_ );
  assign \new_[8865]_  = ~\new_[9277]_  & (~\new_[9539]_  | ~\new_[11143]_ );
  assign \new_[8866]_  = ~\new_[9302]_  & (~\new_[9535]_  | ~\new_[11143]_ );
  assign \new_[8867]_  = ~\new_[9263]_  & (~\new_[9538]_  | ~\new_[11143]_ );
  assign \new_[8868]_  = ~\new_[9301]_  & (~\new_[9548]_  | ~\new_[10829]_ );
  assign \new_[8869]_  = ~\new_[9300]_  & (~\new_[9547]_  | ~\new_[11143]_ );
  assign \new_[8870]_  = ~\new_[9256]_  & (~\new_[9540]_  | ~\new_[11143]_ );
  assign \new_[8871]_  = ~\new_[9266]_  & (~\new_[9542]_  | ~\new_[11143]_ );
  assign \new_[8872]_  = ~\new_[9269]_  & (~\new_[9543]_  | ~\new_[11143]_ );
  assign \new_[8873]_  = ~\new_[9132]_ ;
  assign \new_[8874]_  = ~\new_[9132]_ ;
  assign \new_[8875]_  = ~\new_[9132]_ ;
  assign \new_[8876]_  = ~\new_[9132]_ ;
  assign \new_[8877]_  = ~\new_[9132]_ ;
  assign \new_[8878]_  = ~\new_[9068]_ ;
  assign \new_[8879]_  = ~\new_[9278]_  & (~\new_[9537]_  | ~\new_[11143]_ );
  assign \new_[8880]_  = ~\new_[9047]_ ;
  assign \new_[8881]_  = ~\new_[9136]_ ;
  assign \new_[8882]_  = ~\new_[9268]_  & (~\new_[9536]_  | ~\new_[11143]_ );
  assign n7700 = ~\new_[11504]_  & ~\new_[9490]_ ;
  assign \new_[8884]_  = ~\new_[9434]_ ;
  assign \new_[8885]_  = ~\new_[9434]_ ;
  assign \new_[8886]_  = ~\new_[9139]_ ;
  assign n7685 = ~\new_[11877]_  & ~\new_[9490]_ ;
  assign \new_[8888]_  = \\u1_u3_tx_data_to_cnt_reg[7] ;
  assign \new_[8889]_  = ~\new_[9144]_ ;
  assign \new_[8890]_  = ~\new_[4070]_  | ~\new_[9354]_  | ~\new_[3938]_ ;
  assign \new_[8891]_  = ~\new_[9886]_  | ~\new_[10804]_  | ~\new_[9903]_  | ~\new_[10273]_ ;
  assign \new_[8892]_  = ~\new_[9484]_  & ~\new_[11323]_ ;
  assign \new_[8893]_  = ~\new_[9294]_  & (~\new_[9544]_  | ~\new_[10839]_ );
  assign \new_[8894]_  = ~\new_[9240]_  & (~\new_[9551]_  | ~\new_[10839]_ );
  assign \new_[8895]_  = ~\new_[9242]_  & (~\new_[9534]_  | ~\new_[10839]_ );
  assign \new_[8896]_  = ~\new_[9244]_  & (~\new_[9549]_  | ~\new_[10839]_ );
  assign \new_[8897]_  = ~\new_[9249]_  & (~\new_[9818]_  | ~\new_[10839]_ );
  assign \new_[8898]_  = \new_[9468]_  & \new_[11077]_ ;
  assign \new_[8899]_  = ~\new_[9252]_  & (~\new_[9819]_  | ~\new_[2704]_ );
  assign \new_[8900]_  = ~\new_[9261]_  & (~\new_[9541]_  | ~\new_[10839]_ );
  assign \new_[8901]_  = ~\new_[9262]_  & (~\new_[10030]_  | ~\new_[10475]_ );
  assign n7695 = ~\new_[9490]_  & ~\new_[11488]_ ;
  assign \new_[8903]_  = ~\new_[9290]_  & (~\new_[9819]_  | ~\new_[2637]_ );
  assign \new_[8904]_  = ~\new_[3315]_  | ~\new_[9336]_  | ~\new_[3466]_ ;
  assign \new_[8905]_  = ~\new_[9250]_  & (~\new_[9819]_  | ~\new_[2737]_ );
  assign \new_[8906]_  = ~\new_[3479]_  | ~\new_[9349]_  | ~\new_[3686]_ ;
  assign \new_[8907]_  = ~\new_[9102]_ ;
  assign \new_[8908]_  = ~\new_[9102]_ ;
  assign \new_[8909]_  = ~\new_[9102]_ ;
  assign \new_[8910]_  = ~\new_[9156]_ ;
  assign \new_[8911]_  = ~\new_[9158]_ ;
  assign \new_[8912]_  = ~\new_[3690]_  | ~\new_[9356]_  | ~\new_[3879]_ ;
  assign \new_[8913]_  = ~\new_[9207]_  & (~\new_[11933]_  | ~\new_[11736]_ );
  assign \new_[8914]_  = ~\new_[9162]_ ;
  assign \new_[8915]_  = ~\new_[9475]_  | ~\new_[13238]_ ;
  assign \new_[8916]_  = ~\new_[11077]_  | ~\new_[10425]_  | ~\new_[9721]_  | ~\new_[10856]_ ;
  assign n7675 = ~\new_[9474]_  | (~\new_[9802]_  & ~\new_[6198]_ );
  assign \new_[8918]_  = ~\new_[11210]_  & (~\new_[9689]_  | ~\new_[11971]_ );
  assign \new_[8919]_  = ~\new_[9195]_  | (~\new_[13478]_  & ~\new_[4620]_ );
  assign n7680 = ~\new_[9482]_  | (~\new_[9801]_  & ~\new_[6092]_ );
  assign \new_[8921]_  = \new_[9516]_  ? \new_[9823]_  : \new_[9794]_ ;
  assign \new_[8922]_  = ~\new_[11214]_  & (~\new_[9685]_  | ~\new_[12000]_ );
  assign \new_[8923]_  = (~\new_[9649]_  | ~\new_[3889]_ ) & (~\new_[9609]_  | ~\new_[3888]_ );
  assign \new_[8924]_  = (~\new_[9946]_  | ~\new_[4206]_ ) & (~\new_[9608]_  | ~\new_[4293]_ );
  assign n7705 = \new_[6461]_  ^ \new_[9520]_ ;
  assign n7690 = \new_[6324]_  ^ \new_[9511]_ ;
  assign \new_[8927]_  = ~\new_[9466]_  | ~\new_[9723]_ ;
  assign \new_[8928]_  = ~\new_[9956]_  | ~\new_[10692]_  | ~\new_[10691]_  | ~\new_[10706]_ ;
  assign \new_[8929]_  = u4_u0_dma_req_in_hold_reg;
  assign \new_[8930]_  = ~\new_[9531]_  | ~\new_[10097]_ ;
  assign \new_[8931]_  = \new_[9526]_  & \new_[9276]_ ;
  assign \new_[8932]_  = ~\new_[9526]_  & ~\new_[9276]_ ;
  assign \new_[8933]_  = ~\new_[9272]_  & (~\new_[11125]_  | ~\new_[10086]_ );
  assign \new_[8934]_  = ~\new_[9291]_  & (~\new_[11113]_  | ~\new_[10086]_ );
  assign \new_[8935]_  = ~\new_[9279]_  & (~\new_[10826]_  | ~\new_[10086]_ );
  assign \new_[8936]_  = ~n7900 & ~\new_[9228]_ ;
  assign \new_[8937]_  = ~\new_[14508]_  | ~\new_[12610]_  | ~\new_[9589]_  | ~\new_[9563]_ ;
  assign \new_[8938]_  = ~\new_[9292]_  & (~\new_[9581]_  | ~\new_[10835]_ );
  assign \new_[8939]_  = ~\new_[9505]_  & (~\new_[9573]_  | ~\new_[10835]_ );
  assign \new_[8940]_  = ~\new_[9246]_  & (~\new_[9580]_  | ~\new_[11143]_ );
  assign \new_[8941]_  = ~\new_[9804]_  | ~\new_[9352]_ ;
  assign \new_[8942]_  = ~\new_[9507]_  & (~\new_[9564]_  | ~\new_[10835]_ );
  assign \new_[8943]_  = ~\new_[9508]_  & (~\new_[9571]_  | ~\new_[10835]_ );
  assign \new_[8944]_  = ~\new_[9251]_  & (~\new_[9737]_  | ~\new_[10839]_ );
  assign \new_[8945]_  = (~\new_[9615]_  | ~\new_[11727]_ ) & (~\new_[13315]_  | ~\new_[3469]_ );
  assign \new_[8946]_  = ~\new_[9245]_  & (~\new_[9585]_  | ~\new_[10839]_ );
  assign \new_[8947]_  = \new_[13819]_  ? \new_[10715]_  : \new_[9614]_ ;
  assign \new_[8948]_  = ~\new_[9273]_  & (~\new_[9655]_  | ~\new_[10835]_ );
  assign \new_[8949]_  = ~\new_[9295]_  & (~\new_[9583]_  | ~\new_[10835]_ );
  assign \new_[8950]_  = ~\new_[9308]_  | ~\new_[9842]_ ;
  assign \new_[8951]_  = ~\new_[9211]_  | ~\new_[6850]_ ;
  assign \new_[8952]_  = ~\new_[9285]_  & (~\new_[9675]_  | ~\new_[10839]_ );
  assign \new_[8953]_  = ~\new_[9237]_  & (~\new_[9584]_  | ~\new_[10835]_ );
  assign \new_[8954]_  = \\u1_u3_tx_data_to_cnt_reg[5] ;
  assign \new_[8955]_  = ~\new_[9794]_  | ~\new_[9218]_ ;
  assign \new_[8956]_  = ~\new_[9284]_  & (~\new_[9586]_  | ~\new_[10839]_ );
  assign \new_[8957]_  = ~\new_[9311]_  & (~\new_[11955]_  | ~\new_[13740]_ );
  assign \new_[8958]_  = ~\new_[9298]_  & (~\new_[9582]_  | ~\new_[10835]_ );
  assign \new_[8959]_  = u0_u0_mode_hs_reg;
  assign \new_[8960]_  = ~\new_[13267]_  | ~\new_[9233]_  | ~\new_[14060]_ ;
  assign \new_[8961]_  = ~\new_[9837]_  & ~\new_[9228]_ ;
  assign n7725 = \new_[9304]_  | \new_[9305]_ ;
  assign \new_[8963]_  = ~\new_[9515]_  & (~\new_[9572]_  | ~\new_[10835]_ );
  assign \new_[8964]_  = ~\new_[14383]_  | ~\new_[13456]_  | ~\new_[11586]_  | ~\new_[14739]_ ;
  assign \new_[8965]_  = ~\new_[13135]_  | ~\new_[14347]_  | ~\new_[13155]_ ;
  assign \new_[8966]_  = ~\new_[9552]_  & (~\new_[4815]_  | ~\new_[13646]_ );
  assign \new_[8967]_  = ~\new_[9553]_  & (~\new_[4841]_  | ~\new_[14453]_ );
  assign \new_[8968]_  = (~\new_[9951]_  | ~\new_[10465]_ ) & (~\new_[10467]_  | ~\new_[12056]_ );
  assign \new_[8969]_  = \new_[12643]_  ? \new_[9857]_  : \new_[2096]_ ;
  assign \new_[8970]_  = u4_u3_ep_match_r_reg;
  assign \new_[8971]_  = ~\new_[9633]_  & (~\new_[3690]_  | ~\new_[13913]_ );
  assign \new_[8972]_  = ~\new_[9824]_  | ~n7735;
  assign \new_[8973]_  = \new_[13858]_  & \new_[10096]_ ;
  assign \new_[8974]_  = \new_[11698]_  | \new_[10096]_ ;
  assign \new_[8975]_  = \new_[12124]_  | \new_[11328]_  | \new_[11300]_  | \new_[9892]_ ;
  assign \new_[8976]_  = ~\new_[13311]_  | ~\new_[10096]_ ;
  assign \new_[8977]_  = ~\new_[13288]_  | ~\new_[10096]_ ;
  assign \new_[8978]_  = ~\new_[9226]_ ;
  assign \new_[8979]_  = ~\new_[9229]_ ;
  assign \new_[8980]_  = \new_[13398]_  & \new_[10096]_ ;
  assign \new_[8981]_  = ~\new_[9234]_ ;
  assign \new_[8982]_  = ~\new_[9236]_ ;
  assign \new_[8983]_  = ~\new_[9588]_  | ~\new_[10839]_ ;
  assign \new_[8984]_  = ~\new_[11587]_  & (~\new_[10597]_  | ~\new_[9859]_ );
  assign \new_[8985]_  = ~\new_[9238]_ ;
  assign \new_[8986]_  = ~\new_[9239]_ ;
  assign \new_[8987]_  = ~\new_[9241]_ ;
  assign \new_[8988]_  = ~\new_[9243]_ ;
  assign \new_[8989]_  = ~\new_[10272]_  & (~\new_[9873]_  | ~\new_[10155]_ );
  assign \new_[8990]_  = ~\new_[10272]_  & (~\new_[9868]_  | ~\new_[10240]_ );
  assign \new_[8991]_  = ~\new_[9247]_ ;
  assign \new_[8992]_  = ~\new_[9253]_ ;
  assign \new_[8993]_  = ~\new_[10272]_  & (~\new_[10256]_  | ~\new_[9863]_ );
  assign \new_[8994]_  = ~\new_[9255]_ ;
  assign \new_[8995]_  = ~\new_[10272]_  & (~\new_[10592]_  | ~\new_[9861]_ );
  assign \new_[8996]_  = ~\new_[9257]_ ;
  assign \new_[8997]_  = ~\new_[9259]_ ;
  assign \new_[8998]_  = ~\new_[9260]_ ;
  assign \new_[8999]_  = ~\new_[9264]_ ;
  assign \new_[9000]_  = ~\new_[10272]_  & (~\new_[9864]_  | ~\new_[10183]_ );
  assign \new_[9001]_  = ~\new_[9267]_ ;
  assign \new_[9002]_  = ~\new_[10272]_  & (~\new_[10603]_  | ~\new_[9865]_ );
  assign \new_[9003]_  = ~\new_[11587]_  & (~\new_[10579]_  | ~\new_[9866]_ );
  assign \new_[9004]_  = ~\new_[11123]_  & (~\new_[10591]_  | ~\new_[9880]_ );
  assign \new_[9005]_  = ~\new_[11130]_  & (~\new_[10589]_  | ~\new_[9867]_ );
  assign \new_[9006]_  = ~\new_[9579]_  | ~\new_[10839]_ ;
  assign \new_[9007]_  = ~\new_[9568]_  | ~\new_[10835]_ ;
  assign \new_[9008]_  = ~\new_[9280]_ ;
  assign \new_[9009]_  = ~\new_[10272]_  & (~\new_[10595]_  | ~\new_[9872]_ );
  assign \new_[9010]_  = ~\new_[9281]_ ;
  assign \new_[9011]_  = ~\new_[11130]_  & (~\new_[10586]_  | ~\new_[9862]_ );
  assign \new_[9012]_  = ~\new_[9287]_ ;
  assign \new_[9013]_  = ~\new_[9288]_ ;
  assign \new_[9014]_  = ~\new_[10272]_  & (~\new_[9877]_  | ~\new_[10170]_ );
  assign \new_[9015]_  = ~\new_[9570]_  | ~\new_[10835]_ ;
  assign \new_[9016]_  = ~\new_[10272]_  & (~\new_[10584]_  | ~\new_[9879]_ );
  assign \new_[9017]_  = ~\new_[9297]_ ;
  assign \new_[9018]_  = ~\new_[11587]_  & (~\new_[9858]_  | ~\new_[10538]_ );
  assign \new_[9019]_  = ~\new_[9299]_ ;
  assign \new_[9020]_  = ~\new_[14537]_ ;
  assign \new_[9021]_  = \new_[9852]_  ? \new_[10125]_  : \new_[3311]_ ;
  assign \new_[9022]_  = ~\new_[12131]_  | (~\new_[9883]_  & ~\new_[12390]_ );
  assign \new_[9023]_  = ~\new_[12116]_  | (~\new_[9851]_  & ~\new_[12241]_ );
  assign \new_[9024]_  = ~\new_[11836]_  | (~\new_[9930]_  & ~\new_[12319]_ );
  assign \new_[9025]_  = ~\new_[11838]_  | (~\new_[9757]_  & ~\new_[12225]_ );
  assign \new_[9026]_  = ~\new_[9609]_  | ~\new_[3889]_ ;
  assign \new_[9027]_  = ~\new_[9608]_  | ~\new_[4206]_ ;
  assign \new_[9028]_  = ~\new_[9620]_ ;
  assign \new_[9029]_  = ~\new_[9028]_ ;
  assign \new_[9030]_  = ~\new_[9028]_ ;
  assign \new_[9031]_  = ~\new_[13778]_  | ~\new_[9603]_  | ~\new_[12562]_ ;
  assign \new_[9032]_  = ~\new_[9352]_ ;
  assign \new_[9033]_  = ~\new_[9649]_  | ~\new_[9609]_ ;
  assign \new_[9034]_  = ~\new_[9946]_  | ~\new_[9608]_ ;
  assign \new_[9035]_  = ~\new_[9612]_  & (~\new_[13694]_  | ~\new_[13297]_ );
  assign \new_[9036]_  = ~\new_[14409]_ ;
  assign \new_[9037]_  = \\u1_u3_idin_reg[22] ;
  assign \new_[9038]_  = ~\\u4_u1_buf0_orig_m3_reg[3] ;
  assign \new_[9039]_  = ~\new_[9627]_  | ~\new_[13238]_ ;
  assign \new_[9040]_  = ~\new_[9634]_  & (~\new_[4070]_  | ~\new_[13904]_ );
  assign \new_[9041]_  = ~\new_[13249]_  | ~\new_[9617]_  | ~\new_[13034]_ ;
  assign \new_[9042]_  = ~\new_[13094]_  | ~\new_[9619]_  | ~\new_[13063]_ ;
  assign \new_[9043]_  = ~\new_[9625]_  | ~\new_[12913]_ ;
  assign \new_[9044]_  = ~\new_[12544]_  | ~\new_[9622]_  | ~\new_[13103]_ ;
  assign \new_[9045]_  = ~\new_[12613]_  | ~\new_[9624]_  | ~\new_[13017]_ ;
  assign \new_[9046]_  = \new_[2083]_  ^ \new_[9958]_ ;
  assign \new_[9047]_  = ~\new_[9429]_ ;
  assign \new_[9048]_  = ~\new_[9430]_ ;
  assign \new_[9049]_  = \new_[3938]_  ^ \new_[9927]_ ;
  assign \new_[9050]_  = \new_[3466]_  ^ \new_[9929]_ ;
  assign \new_[9051]_  = \new_[3686]_  ^ \new_[9933]_ ;
  assign \new_[9052]_  = \new_[3879]_  ^ \new_[9931]_ ;
  assign \new_[9053]_  = \new_[9628]_  | \new_[6252]_ ;
  assign \new_[9054]_  = ~\\u4_u3_buf0_orig_m3_reg[7] ;
  assign \new_[9055]_  = ~\\u4_u2_buf0_orig_m3_reg[7] ;
  assign \new_[9056]_  = \new_[9629]_  | \new_[6563]_ ;
  assign \new_[9057]_  = \new_[9629]_  | \new_[5999]_ ;
  assign n7650 = ~\new_[9028]_ ;
  assign \new_[9059]_  = ~\\u4_u3_buf0_orig_m3_reg[8] ;
  assign \new_[9060]_  = \new_[9628]_  | \new_[6251]_ ;
  assign \new_[9061]_  = \new_[9630]_  | \new_[6004]_ ;
  assign \new_[9062]_  = \new_[9630]_  | \new_[6274]_ ;
  assign \new_[9063]_  = \new_[9631]_  | \new_[6544]_ ;
  assign \new_[9064]_  = \new_[9631]_  | \new_[6286]_ ;
  assign \new_[9065]_  = ~\\u4_u2_buf0_orig_m3_reg[8] ;
  assign \new_[9066]_  = (~\new_[9964]_  | ~\new_[4801]_ ) & (~\new_[11011]_  | ~\new_[11328]_ );
  assign \new_[9067]_  = ~\new_[9380]_ ;
  assign \new_[9068]_  = ~\new_[9380]_ ;
  assign \new_[9069]_  = \new_[10693]_  ? \new_[9857]_  : \new_[2097]_ ;
  assign \new_[9070]_  = \new_[11807]_  ^ \new_[9941]_ ;
  assign \new_[9071]_  = \new_[12178]_  ^ \new_[9942]_ ;
  assign \new_[9072]_  = \new_[12026]_  ^ \new_[9940]_ ;
  assign \new_[9073]_  = ~\new_[13386]_  | ~\new_[9532]_  | ~\new_[13659]_ ;
  assign \new_[9074]_  = \new_[11980]_  ^ \new_[9943]_ ;
  assign \new_[9075]_  = \\u4_int_srca_reg[1] ;
  assign \new_[9076]_  = \new_[9685]_  | \new_[10455]_ ;
  assign \new_[9077]_  = \new_[9689]_  | \new_[10456]_ ;
  assign \new_[9078]_  = \new_[9690]_  | \new_[10701]_ ;
  assign \new_[9079]_  = \new_[9693]_  | \new_[10459]_ ;
  assign \new_[9080]_  = ~\new_[9641]_  | ~\new_[13238]_ ;
  assign \new_[9081]_  = ~\new_[9667]_  & (~\new_[13970]_  | ~\new_[13297]_ );
  assign \new_[9082]_  = ~\new_[9425]_ ;
  assign \new_[9083]_  = ~\new_[12830]_  & (~\new_[9998]_  | ~\new_[12131]_ );
  assign \new_[9084]_  = \new_[2349]_  ^ \new_[9822]_ ;
  assign \new_[9085]_  = ~\new_[10063]_  | ~\new_[12082]_  | ~\new_[10814]_  | ~\new_[14167]_ ;
  assign \new_[9086]_  = ~\new_[10609]_  | ~\new_[12113]_  | ~\new_[9749]_  | ~\new_[11643]_ ;
  assign \new_[9087]_  = ~\wb_addr_i[2]  | ~\new_[12718]_  | ~\new_[9991]_ ;
  assign \new_[9088]_  = ~\new_[11988]_  & ~\new_[14637]_ ;
  assign \new_[9089]_  = ~\new_[11441]_  & ~\new_[14637]_ ;
  assign \new_[9090]_  = ~\new_[10305]_  & ~\new_[14637]_ ;
  assign \new_[9091]_  = ~\new_[14637]_  & ~\new_[10115]_ ;
  assign \new_[9092]_  = ~\new_[14637]_  & ~\new_[10360]_ ;
  assign \new_[9093]_  = ~\new_[14637]_  & ~\new_[9613]_ ;
  assign \new_[9094]_  = ~\new_[12656]_  & (~\new_[10001]_  | ~\new_[12116]_ );
  assign \new_[9095]_  = ~\new_[9650]_  & ~\new_[12524]_ ;
  assign \new_[9096]_  = ~\new_[12754]_  & (~\new_[10000]_  | ~\new_[11836]_ );
  assign \new_[9097]_  = ~\new_[9662]_  & (~\new_[11266]_  | ~\new_[4620]_ );
  assign n7740 = \new_[6305]_  ^ \new_[9820]_ ;
  assign \new_[9099]_  = ~\new_[12668]_  & (~\new_[10008]_  | ~\new_[11838]_ );
  assign n7745 = \new_[6556]_  ^ \new_[9976]_ ;
  assign \new_[9101]_  = ~\new_[9448]_ ;
  assign \new_[9102]_  = ~\new_[9448]_ ;
  assign \new_[9103]_  = \new_[14211]_  ? \new_[10715]_  : \new_[9856]_ ;
  assign \new_[9104]_  = ~\new_[9402]_ ;
  assign \new_[9105]_  = ~\new_[12294]_  | ~\new_[12199]_  | ~\new_[9696]_  | ~\new_[13046]_ ;
  assign \new_[9106]_  = ~\new_[9499]_  & ~\new_[9652]_ ;
  assign \new_[9107]_  = ~\new_[9671]_  & (~\new_[3315]_  | ~\new_[13718]_ );
  assign \new_[9108]_  = ~\new_[9677]_  & (~\new_[3479]_  | ~\new_[13548]_ );
  assign \new_[9109]_  = ~\new_[9664]_  | (~\new_[10370]_  & ~\new_[6246]_ );
  assign \new_[9110]_  = \new_[12153]_  ? \new_[9853]_  : \new_[12458]_ ;
  assign \new_[9111]_  = \new_[6604]_  ^ \new_[9760]_ ;
  assign \new_[9112]_  = ~\\u4_u1_buf0_orig_m3_reg[4] ;
  assign n7760 = \new_[11975]_  ^ \new_[9981]_ ;
  assign \new_[9114]_  = \new_[12112]_  ^ \new_[9989]_ ;
  assign n7755 = \new_[11986]_  ^ \new_[9980]_ ;
  assign \new_[9116]_  = \new_[11947]_  ^ \new_[9997]_ ;
  assign n7750 = \new_[12012]_  ^ \new_[9982]_ ;
  assign n7765 = \new_[11802]_  ^ \new_[9979]_ ;
  assign \new_[9119]_  = \new_[11813]_  ^ \new_[9932]_ ;
  assign \new_[9120]_  = \new_[11945]_  ^ \new_[10006]_ ;
  assign \new_[9121]_  = \new_[11760]_  ? \new_[9759]_  : \new_[11640]_ ;
  assign \new_[9122]_  = \new_[6739]_  ^ \new_[9758]_ ;
  assign \new_[9123]_  = (~\new_[9756]_  | ~\new_[11727]_ ) & (~\new_[13315]_  | ~\new_[3474]_ );
  assign \new_[9124]_  = ~\new_[9413]_ ;
  assign \new_[9125]_  = ~\\u4_u1_buf0_orig_m3_reg[2] ;
  assign \new_[9126]_  = ~\\u4_u1_buf0_orig_m3_reg[6] ;
  assign \new_[9127]_  = ~\new_[9419]_ ;
  assign \new_[9128]_  = \new_[9425]_ ;
  assign \new_[9129]_  = ~\new_[9425]_ ;
  assign \new_[9130]_  = ~\new_[9425]_ ;
  assign \new_[9131]_  = ~\new_[9426]_ ;
  assign \new_[9132]_  = ~\new_[9380]_ ;
  assign \new_[9133]_  = ~\new_[9380]_ ;
  assign \new_[9134]_  = ~\new_[9380]_ ;
  assign \new_[9135]_  = ~\new_[9428]_ ;
  assign \new_[9136]_  = ~\new_[9430]_ ;
  assign \new_[9137]_  = ~\new_[9433]_ ;
  assign \new_[9138]_  = ~\new_[9434]_ ;
  assign \new_[9139]_  = \new_[9434]_ ;
  assign \new_[9140]_  = \new_[9493]_  & \new_[9561]_ ;
  assign \new_[9141]_  = ~\new_[9436]_ ;
  assign \new_[9142]_  = ~\new_[9443]_ ;
  assign \new_[9143]_  = ~\new_[9445]_ ;
  assign \new_[9144]_  = ~\new_[9445]_ ;
  assign \new_[9145]_  = ~\new_[9445]_ ;
  assign \new_[9146]_  = ~\new_[13205]_  | ~\new_[11688]_  | ~\new_[9811]_ ;
  assign \new_[9147]_  = ~\new_[9791]_  | ~\new_[9751]_ ;
  assign \new_[9148]_  = ~\dma_req_o[2]  | ~\new_[9714]_  | ~\new_[12640]_ ;
  assign \new_[9149]_  = ~\dma_req_o[3]  | ~\new_[9715]_  | ~\new_[12506]_ ;
  assign \new_[9150]_  = ~\wb_addr_i[2]  | ~\new_[12771]_  | ~\new_[9787]_ ;
  assign \new_[9151]_  = ~\new_[9783]_  | ~\new_[9752]_ ;
  assign \new_[9152]_  = ~\new_[9795]_  | ~\new_[9753]_ ;
  assign \new_[9153]_  = ~\dma_req_o[0]  | ~\new_[9717]_  | ~\new_[12763]_ ;
  assign \new_[9154]_  = ~\new_[10261]_  & (~\new_[9771]_  | ~\new_[7856]_ );
  assign \new_[9155]_  = ~\dma_req_o[1]  | ~\new_[9718]_  | ~\new_[12543]_ ;
  assign \new_[9156]_  = ~\new_[9448]_ ;
  assign \new_[9157]_  = ~\new_[9448]_ ;
  assign \new_[9158]_  = ~\new_[9448]_ ;
  assign \new_[9159]_  = ~\new_[12871]_  | ~\new_[9719]_  | ~\new_[10508]_ ;
  assign \new_[9160]_  = ~\new_[12657]_  | ~\new_[9720]_  | ~\new_[10509]_ ;
  assign \new_[9161]_  = ~\new_[9494]_  & (~\new_[11941]_  | ~\new_[11642]_ );
  assign \new_[9162]_  = ~n7590 | (~\new_[11442]_  & ~\new_[11810]_ );
  assign \new_[9163]_  = \new_[4070]_  ^ \new_[9905]_ ;
  assign \new_[9164]_  = \new_[3315]_  ^ \new_[9906]_ ;
  assign \new_[9165]_  = ~\new_[9575]_  & (~\new_[13297]_  | ~\new_[13608]_ );
  assign \new_[9166]_  = \new_[3479]_  ^ \new_[9908]_ ;
  assign \new_[9167]_  = \new_[3690]_  ^ \new_[9909]_ ;
  assign \new_[9168]_  = ~\new_[9637]_  & (~\new_[11826]_  | ~\new_[13382]_ );
  assign \new_[9169]_  = ~\new_[9742]_  & (~\new_[11828]_  | ~\new_[13473]_ );
  assign \new_[9170]_  = ~\new_[9745]_  & (~\new_[11830]_  | ~\new_[13300]_ );
  assign \new_[9171]_  = ~\new_[9747]_  & (~\new_[11832]_  | ~\new_[13459]_ );
  assign \new_[9172]_  = \new_[4286]_  ^ \new_[9888]_ ;
  assign \new_[9173]_  = \new_[3462]_  ^ \new_[9891]_ ;
  assign \new_[9174]_  = \new_[3592]_  ^ \new_[9902]_ ;
  assign \new_[9175]_  = \new_[3790]_  ^ \new_[9887]_ ;
  assign n7780 = \new_[6351]_  ^ \new_[9793]_ ;
  assign n7770 = \new_[6347]_  ^ \new_[9893]_ ;
  assign \new_[9178]_  = u4_u2_dma_req_in_hold_reg;
  assign \new_[9179]_  = u4_u1_dma_req_in_hold_reg;
  assign n7790 = ~\new_[12804]_  & (~\new_[9827]_  | ~\new_[11626]_ );
  assign n7785 = ~\new_[11973]_  & (~\new_[9854]_  | ~\new_[9838]_ );
  assign n7775 = \new_[6348]_  ^ \new_[9895]_ ;
  assign \new_[9183]_  = ~\new_[9521]_  | ~\new_[13165]_ ;
  assign \new_[9184]_  = \new_[12075]_  | \new_[9524]_ ;
  assign \new_[9185]_  = ~\new_[9506]_  | ~\new_[13257]_ ;
  assign \new_[9186]_  = ~\new_[14346]_  & ~\new_[11006]_ ;
  assign \new_[9187]_  = ~\new_[14346]_  & (~\new_[10805]_  | ~\new_[11430]_ );
  assign \new_[9188]_  = u1_u3_out_token_reg;
  assign \new_[9189]_  = ~\new_[9506]_  | ~\new_[9799]_ ;
  assign \new_[9190]_  = ~\new_[14346]_  & (~\new_[11801]_  | ~\new_[14167]_ );
  assign \new_[9191]_  = u1_u3_setup_token_reg;
  assign \new_[9192]_  = ~\new_[10033]_  & (~\new_[9841]_  | ~\new_[10835]_ );
  assign \new_[9193]_  = \new_[9518]_  | \new_[11747]_ ;
  assign \new_[9194]_  = ~\new_[10630]_  | ~\new_[12573]_  | ~\new_[9843]_  | ~\new_[10465]_ ;
  assign \new_[9195]_  = ~\new_[10506]_  & (~\new_[10461]_  | ~\new_[10112]_ );
  assign \new_[9196]_  = ~\new_[10480]_  | ~\new_[9842]_  | ~\new_[11105]_ ;
  assign \new_[9197]_  = (~\new_[10099]_  & ~\new_[12778]_ ) | (~\new_[12363]_  & ~\new_[4791]_ );
  assign \new_[9198]_  = ~\new_[13028]_  & (~\new_[10088]_  | ~\new_[10836]_ );
  assign \new_[9199]_  = ~\new_[9776]_  & (~\new_[11517]_  | ~\new_[7670]_ );
  assign \new_[9200]_  = ~\new_[10112]_  | ~\new_[9855]_  | ~\new_[10427]_ ;
  assign \new_[9201]_  = \new_[3283]_  ^ \new_[10283]_ ;
  assign \new_[9202]_  = \new_[3308]_  ^ \new_[10092]_ ;
  assign \new_[9203]_  = \new_[3309]_  ^ \new_[10249]_ ;
  assign \new_[9204]_  = \new_[3282]_  ^ \new_[10079]_ ;
  assign \new_[9205]_  = ~\new_[9766]_  | (~\new_[6368]_  & ~\new_[13912]_ );
  assign \new_[9206]_  = ~\new_[9767]_  | (~\new_[6300]_  & ~\new_[13623]_ );
  assign \new_[9207]_  = ~\new_[9768]_  & (~\new_[14043]_  | ~\new_[3505]_ );
  assign \new_[9208]_  = ~\new_[11674]_  | ~\new_[11588]_  | ~\new_[9838]_  | ~\new_[10574]_ ;
  assign n7870 = \new_[6322]_  ^ \new_[10081]_ ;
  assign n7875 = \new_[6370]_  ^ \new_[10091]_ ;
  assign \new_[9211]_  = u0_u0_ls_idle_r_reg;
  assign n7895 = \new_[9911]_  & \new_[9845]_ ;
  assign \new_[9213]_  = ~\new_[9501]_ ;
  assign \new_[9214]_  = ~\new_[9857]_  | ~\new_[2093]_ ;
  assign \new_[9215]_  = ~\new_[9857]_  | ~\new_[2094]_ ;
  assign \new_[9216]_  = ~\new_[9857]_  | ~\new_[2088]_ ;
  assign \new_[9217]_  = ~\new_[9857]_  | ~\new_[2091]_ ;
  assign \new_[9218]_  = ~\new_[9823]_  & ~\new_[10087]_ ;
  assign \new_[9219]_  = ~\new_[9823]_  | ~\new_[10440]_ ;
  assign \new_[9220]_  = ~\new_[9857]_  | ~\new_[2083]_ ;
  assign \new_[9221]_  = ~\new_[11698]_  & ~\new_[11006]_ ;
  assign \new_[9222]_  = ~\new_[9857]_  | ~\new_[2084]_ ;
  assign \new_[9223]_  = ~\new_[9857]_  | ~\new_[2087]_ ;
  assign \new_[9224]_  = ~\new_[9857]_  | ~\new_[2086]_ ;
  assign \new_[9225]_  = ~\new_[10452]_  | ~\new_[13407]_ ;
  assign \new_[9226]_  = ~\new_[10089]_  | ~\new_[9830]_ ;
  assign \new_[9227]_  = ~\new_[9857]_  | ~\new_[2092]_ ;
  assign \new_[9228]_  = ~\new_[9824]_  | ~\new_[9836]_ ;
  assign \new_[9229]_  = ~\new_[9844]_  | ~\new_[4387]_ ;
  assign \new_[9230]_  = \new_[9823]_  | \new_[10440]_ ;
  assign \new_[9231]_  = ~\new_[9857]_  | ~\new_[2089]_ ;
  assign \new_[9232]_  = ~\new_[9523]_ ;
  assign \new_[9233]_  = ~\new_[9524]_ ;
  assign \new_[9234]_  = ~\new_[11123]_  & (~\new_[10234]_  | ~\new_[10533]_ );
  assign \new_[9235]_  = ~\new_[11123]_  & (~\new_[10241]_  | ~\new_[10551]_ );
  assign \new_[9236]_  = ~\new_[11123]_  & (~\new_[10152]_  | ~\new_[10198]_ );
  assign \new_[9237]_  = ~\new_[11123]_  & (~\new_[10314]_  | ~\new_[10136]_ );
  assign \new_[9238]_  = ~\new_[11123]_  & (~\new_[10194]_  | ~\new_[10147]_ );
  assign \new_[9239]_  = ~\new_[11123]_  & (~\new_[10150]_  | ~\new_[10151]_ );
  assign \new_[9240]_  = ~\new_[11587]_  & (~\new_[10137]_  | ~\new_[10516]_ );
  assign \new_[9241]_  = ~\new_[11123]_  & (~\new_[10149]_  | ~\new_[10546]_ );
  assign \new_[9242]_  = ~\new_[11587]_  & (~\new_[10182]_  | ~\new_[10517]_ );
  assign \new_[9243]_  = ~\new_[11123]_  & (~\new_[10238]_  | ~\new_[10196]_ );
  assign \new_[9244]_  = ~\new_[11587]_  & (~\new_[10247]_  | ~\new_[10545]_ );
  assign \new_[9245]_  = ~\new_[11123]_  & (~\new_[10604]_  | ~\new_[10237]_ );
  assign \new_[9246]_  = ~\new_[11123]_  & (~\new_[10407]_  | ~\new_[10157]_ );
  assign \new_[9247]_  = ~\new_[11123]_  & (~\new_[10220]_  | ~\new_[10158]_ );
  assign \new_[9248]_  = ~\new_[10272]_  & (~\new_[10148]_  | ~\new_[10199]_ );
  assign \new_[9249]_  = ~\new_[11587]_  & (~\new_[10202]_  | ~\new_[10540]_ );
  assign \new_[9250]_  = ~\new_[11587]_  & (~\new_[10594]_  | ~\new_[10208]_ );
  assign \new_[9251]_  = ~\new_[10272]_  & (~\new_[10287]_  | ~\new_[10166]_ );
  assign \new_[9252]_  = ~\new_[11587]_  & (~\new_[10585]_  | ~\new_[10167]_ );
  assign \new_[9253]_  = ~\new_[11123]_  & (~\new_[10257]_  | ~\new_[10168]_ );
  assign \new_[9254]_  = ~\new_[10272]_  & (~\new_[10143]_  | ~\new_[10156]_ );
  assign \new_[9255]_  = ~\new_[11123]_  & (~\new_[10153]_  | ~\new_[10522]_ );
  assign \new_[9256]_  = ~\new_[11130]_  & (~\new_[10171]_  | ~\new_[10523]_ );
  assign \new_[9257]_  = ~\new_[11123]_  & (~\new_[10224]_  | ~\new_[10561]_ );
  assign \new_[9258]_  = ~\new_[10272]_  & (~\new_[10173]_  | ~\new_[10174]_ );
  assign \new_[9259]_  = ~\new_[11123]_  & (~\new_[10146]_  | ~\new_[10219]_ );
  assign \new_[9260]_  = ~\new_[11123]_  & (~\new_[10175]_  | ~\new_[10176]_ );
  assign \new_[9261]_  = ~\new_[11587]_  & (~\new_[10177]_  | ~\new_[10178]_ );
  assign \new_[9262]_  = ~\new_[10272]_  & (~\new_[10179]_  | ~\new_[10180]_ );
  assign \new_[9263]_  = ~\new_[11130]_  & (~\new_[10161]_  | ~\new_[10511]_ );
  assign \new_[9264]_  = ~\new_[11123]_  & (~\new_[10133]_  | ~\new_[10525]_ );
  assign \new_[9265]_  = ~\new_[10272]_  & (~\new_[10172]_  | ~\new_[10134]_ );
  assign \new_[9266]_  = ~\new_[11130]_  & (~\new_[10132]_  | ~\new_[10526]_ );
  assign \new_[9267]_  = ~\new_[11123]_  & (~\new_[10185]_  | ~\new_[10528]_ );
  assign \new_[9268]_  = ~\new_[11130]_  & (~\new_[10159]_  | ~\new_[10531]_ );
  assign \new_[9269]_  = ~\new_[11130]_  & (~\new_[10186]_  | ~\new_[10529]_ );
  assign \new_[9270]_  = ~\new_[11123]_  & (~\new_[10578]_  | ~\new_[10187]_ );
  assign \new_[9271]_  = ~\new_[11587]_  & (~\new_[10601]_  | ~\new_[10188]_ );
  assign \new_[9272]_  = ~\new_[11587]_  & (~\new_[10700]_  | ~\new_[10189]_ );
  assign \new_[9273]_  = ~\new_[11123]_  & (~\new_[10265]_  | ~\new_[10230]_ );
  assign \new_[9274]_  = ~\new_[2874]_  | ~\new_[14830]_  | ~\new_[10490]_ ;
  assign \new_[9275]_  = ~\new_[9526]_ ;
  assign \new_[9276]_  = ~\new_[14156]_  | ~\new_[13398]_  | ~\new_[9826]_  | ~\new_[14385]_ ;
  assign \new_[9277]_  = ~\new_[11130]_  & (~\new_[10184]_  | ~\new_[10536]_ );
  assign \new_[9278]_  = ~\new_[11130]_  & (~\new_[10068]_  | ~\new_[10518]_ );
  assign \new_[9279]_  = ~\new_[11587]_  & (~\new_[10588]_  | ~\new_[10138]_ );
  assign \new_[9280]_  = ~\new_[11123]_  & (~\new_[10245]_  | ~\new_[10215]_ );
  assign \new_[9281]_  = ~\new_[11587]_  & (~\new_[10587]_  | ~\new_[10203]_ );
  assign \new_[9282]_  = ~\new_[2875]_  | ~\new_[14830]_  | ~\new_[10490]_ ;
  assign \new_[9283]_  = ~\new_[11130]_  & (~\new_[10209]_  | ~\new_[10513]_ );
  assign \new_[9284]_  = ~\new_[11587]_  & (~\new_[10253]_  | ~\new_[10181]_ );
  assign \new_[9285]_  = ~\new_[11587]_  & (~\new_[10269]_  | ~\new_[10140]_ );
  assign \new_[9286]_  = ~\new_[11130]_  & (~\new_[10233]_  | ~\new_[10514]_ );
  assign \new_[9287]_  = ~\new_[11123]_  & (~\new_[10135]_  | ~\new_[10144]_ );
  assign \new_[9288]_  = ~\new_[11123]_  & (~\new_[10260]_  | ~\new_[10207]_ );
  assign \new_[9289]_  = ~\new_[13508]_  | ~\new_[9842]_  | ~n9145;
  assign \new_[9290]_  = ~\new_[11587]_  & (~\new_[10213]_  | ~\new_[10957]_ );
  assign \new_[9291]_  = ~\new_[11587]_  & (~\new_[10598]_  | ~\new_[10227]_ );
  assign \new_[9292]_  = ~\new_[11123]_  & (~\new_[10259]_  | ~\new_[10195]_ );
  assign n7885 = \new_[9840]_  & \new_[13044]_ ;
  assign \new_[9294]_  = ~\new_[11587]_  & (~\new_[10210]_  | ~\new_[10519]_ );
  assign \new_[9295]_  = ~\new_[11123]_  & (~\new_[10255]_  | ~\new_[10162]_ );
  assign \new_[9296]_  = ~\new_[10272]_  & (~\new_[10214]_  | ~\new_[10164]_ );
  assign \new_[9297]_  = ~\new_[11123]_  & (~\new_[10212]_  | ~\new_[10541]_ );
  assign \new_[9298]_  = ~\new_[11123]_  & (~\new_[10254]_  | ~\new_[10211]_ );
  assign \new_[9299]_  = ~\new_[11123]_  & (~\new_[10218]_  | ~\new_[10204]_ );
  assign \new_[9300]_  = ~\new_[11130]_  & (~\new_[10142]_  | ~\new_[10520]_ );
  assign \new_[9301]_  = ~\new_[11130]_  & (~\new_[10193]_  | ~\new_[10139]_ );
  assign \new_[9302]_  = ~\new_[11130]_  & (~\new_[10244]_  | ~\new_[10534]_ );
  assign \new_[9303]_  = ~\new_[11123]_  & (~\new_[10268]_  | ~\new_[10226]_ );
  assign \new_[9304]_  = (~\new_[10200]_  & ~\new_[11587]_ ) | (~\new_[10163]_  & ~\new_[11130]_ );
  assign \new_[9305]_  = (~\new_[10205]_  & ~\new_[11123]_ ) | (~\new_[10192]_  & ~\new_[10272]_ );
  assign \new_[9306]_  = ~\new_[11192]_  | (~\new_[10322]_  & ~\new_[11618]_ );
  assign \new_[9307]_  = ~\new_[14332]_ ;
  assign \new_[9308]_  = ~\new_[9533]_ ;
  assign \new_[9309]_  = ~\new_[10222]_  | ~\new_[10581]_  | ~\new_[10722]_ ;
  assign \new_[9310]_  = ~\new_[9849]_  & (~\new_[11356]_  | ~\new_[11203]_ );
  assign \new_[9311]_  = (~\new_[4791]_  & ~\new_[4794]_  & ~\new_[12883]_ ) | (~\new_[10124]_  & ~\new_[13426]_  & ~\new_[12883]_ );
  assign \new_[9312]_  = ~\new_[14834]_  & ~\new_[14205]_ ;
  assign \new_[9313]_  = ~\new_[12605]_  & ~\new_[9850]_ ;
  assign \new_[9314]_  = ~\new_[9860]_  | ~\new_[10555]_ ;
  assign \new_[9315]_  = ~\new_[9914]_  | ~\sram_data_i[11] ;
  assign \new_[9316]_  = ~\new_[9914]_  | ~\sram_data_i[22] ;
  assign \new_[9317]_  = ~\new_[9914]_  | ~\sram_data_i[30] ;
  assign n7795 = ~\new_[9562]_ ;
  assign \new_[9319]_  = ~\new_[9914]_  | ~\sram_data_i[12] ;
  assign \new_[9320]_  = ~\new_[9914]_  | ~\sram_data_i[13] ;
  assign \new_[9321]_  = ~\new_[9914]_  | ~\sram_data_i[21] ;
  assign \new_[9322]_  = ~\new_[9914]_  | ~\sram_data_i[28] ;
  assign \new_[9323]_  = ~\new_[9914]_  | ~\sram_data_i[17] ;
  assign \new_[9324]_  = ~\new_[9869]_  | ~\new_[10557]_ ;
  assign \new_[9325]_  = ~\new_[10111]_  & (~\new_[11602]_  | ~\new_[10275]_ );
  assign \new_[9326]_  = ~\new_[9914]_  | ~\sram_data_i[20] ;
  assign \new_[9327]_  = ~\new_[9889]_  & ~\new_[10125]_ ;
  assign n7825 = ~\new_[12646]_  & ~n7980;
  assign \new_[9329]_  = ~\new_[9914]_  | ~\sram_data_i[31] ;
  assign \new_[9330]_  = ~\new_[9914]_  | ~\sram_data_i[23] ;
  assign \new_[9331]_  = ~\new_[9914]_  | ~\sram_data_i[27] ;
  assign \new_[9332]_  = ~\new_[9871]_  | ~\new_[10550]_ ;
  assign \new_[9333]_  = ~\new_[13802]_  | ~\new_[8701]_  | ~\new_[9848]_  | ~\new_[14061]_ ;
  assign \new_[9334]_  = ~\new_[9914]_  | ~\sram_data_i[18] ;
  assign \new_[9335]_  = ~\new_[9914]_  | ~\sram_data_i[10] ;
  assign \new_[9336]_  = ~\new_[9906]_  & ~\new_[13470]_ ;
  assign \new_[9337]_  = ~\new_[9896]_  & ~\new_[10608]_ ;
  assign \new_[9338]_  = \new_[11333]_  & \new_[9893]_ ;
  assign \new_[9339]_  = ~\new_[9914]_  | ~\sram_data_i[14] ;
  assign \new_[9340]_  = ~\new_[9914]_  | ~\sram_data_i[15] ;
  assign \new_[9341]_  = ~\new_[9914]_  | ~\sram_data_i[24] ;
  assign \new_[9342]_  = ~\new_[9914]_  | ~\sram_data_i[25] ;
  assign \new_[9343]_  = ~\new_[9914]_  | ~\sram_data_i[8] ;
  assign \new_[9344]_  = ~\new_[9914]_  | ~\sram_data_i[26] ;
  assign \new_[9345]_  = ~\new_[9914]_  | ~\sram_data_i[29] ;
  assign \new_[9346]_  = ~\new_[9914]_  | ~\sram_data_i[9] ;
  assign \new_[9347]_  = ~\new_[9914]_  | ~\sram_data_i[19] ;
  assign \new_[9348]_  = ~\new_[9914]_  | ~\sram_data_i[16] ;
  assign \new_[9349]_  = ~\new_[9908]_  & ~\new_[13286]_ ;
  assign \new_[9350]_  = ~\new_[11190]_  | (~\new_[10317]_  & ~\new_[11590]_ );
  assign \new_[9351]_  = ~\new_[10251]_  | ~\new_[9874]_ ;
  assign \new_[9352]_  = ~\new_[9955]_  & ~n8240;
  assign \new_[9353]_  = ~\new_[11191]_  | (~\new_[10320]_  & ~\new_[11601]_ );
  assign \new_[9354]_  = ~\new_[9905]_  & ~\new_[12628]_ ;
  assign n7880 = ~\new_[10952]_  & ~n7980;
  assign \new_[9356]_  = ~\new_[9909]_  & ~\new_[12528]_ ;
  assign \new_[9357]_  = ~\new_[9876]_  | (~\new_[6379]_  & ~\new_[13047]_ );
  assign \new_[9358]_  = ~u1_u0_rx_active_r_reg;
  assign \new_[9359]_  = \new_[11338]_  | \new_[9788]_ ;
  assign \new_[9360]_  = \new_[2095]_  ^ \new_[10280]_ ;
  assign \new_[9361]_  = ~\new_[9596]_ ;
  assign n7830 = ~\new_[8703]_  & ~n7980;
  assign \new_[9363]_  = ~\new_[9788]_  & ~\new_[12251]_ ;
  assign \new_[9364]_  = ~\new_[3463]_  | ~\new_[9904]_  | ~\new_[3469]_ ;
  assign \new_[9365]_  = (~\new_[10281]_  | ~\new_[11727]_ ) & (~\new_[13315]_  | ~\new_[3435]_ );
  assign \new_[9366]_  = ~\\u4_u0_buf0_orig_m3_reg[3] ;
  assign \new_[9367]_  = ~\\u4_u3_dma_out_left_reg[4] ;
  assign \new_[9368]_  = ~\\u4_u0_dma_out_left_reg[4] ;
  assign \new_[9369]_  = ~\\u4_u1_dma_out_left_reg[4] ;
  assign \new_[9370]_  = ~\\u4_u2_dma_out_left_reg[4] ;
  assign \new_[9371]_  = ~\new_[9907]_  | (~\new_[10650]_  & ~\new_[3463]_ );
  assign \new_[9372]_  = \\u1_u3_rx_ack_to_cnt_reg[4] ;
  assign \new_[9373]_  = ~\new_[13279]_  | ~\new_[13406]_  | ~\new_[10300]_ ;
  assign n7860 = ~\new_[11397]_  & ~n7980;
  assign \new_[9375]_  = ~n7590;
  assign \new_[9376]_  = ~\new_[14171]_  | ~\new_[9412]_  | ~\new_[9847]_  | ~\new_[14219]_ ;
  assign \new_[9377]_  = ~\new_[2095]_  | ~\new_[2084]_  | ~\new_[9949]_  | ~\new_[13432]_ ;
  assign \new_[9378]_  = \new_[2094]_  ^ \new_[10316]_ ;
  assign \new_[9379]_  = (~\new_[10113]_  | ~\new_[11727]_ ) & (~\new_[13315]_  | ~\new_[3472]_ );
  assign \new_[9380]_  = \new_[13167]_  | \new_[9994]_ ;
  assign \new_[9381]_  = \new_[11607]_  ^ \new_[10318]_ ;
  assign \new_[9382]_  = \new_[11788]_  ^ \new_[10330]_ ;
  assign \new_[9383]_  = \new_[13186]_  ^ \new_[10332]_ ;
  assign \new_[9384]_  = \new_[11611]_  ^ \new_[10320]_ ;
  assign \new_[9385]_  = \new_[11605]_  ^ \new_[10317]_ ;
  assign \new_[9386]_  = \new_[10719]_  ^ \new_[10329]_ ;
  assign \new_[9387]_  = \new_[11706]_  ^ \new_[10322]_ ;
  assign \new_[9388]_  = \\u4_int_srca_reg[0] ;
  assign \new_[9389]_  = \\u4_int_srca_reg[3] ;
  assign \new_[9390]_  = ~\new_[9628]_ ;
  assign \new_[9391]_  = ~\new_[9629]_ ;
  assign \new_[9392]_  = \\u4_int_srca_reg[2] ;
  assign \new_[9393]_  = ~\new_[9630]_ ;
  assign \new_[9394]_  = ~\new_[9631]_ ;
  assign \new_[9395]_  = ~\new_[10501]_  & (~\new_[10090]_  | ~\new_[10353]_ );
  assign \new_[9396]_  = \new_[2348]_  ^ \new_[10248]_ ;
  assign \new_[9397]_  = \new_[2869]_  ^ \new_[10108]_ ;
  assign n7855 = n8050 | \new_[13680]_ ;
  assign n7815 = ~\new_[10968]_  & ~n7980;
  assign \new_[9400]_  = \new_[11153]_  & \new_[9939]_ ;
  assign \new_[9401]_  = ~\new_[12359]_  | ~\new_[12323]_  | ~\new_[9959]_  | ~\new_[12906]_ ;
  assign \new_[9402]_  = \new_[10375]_  | \wb_addr_i[2]  | \new_[11958]_  | \new_[13129]_ ;
  assign \new_[9403]_  = ~\new_[12612]_  | ~\new_[12321]_  | ~\new_[9960]_  | ~\new_[13029]_ ;
  assign \new_[9404]_  = ~\new_[12272]_  | ~\new_[11974]_  | ~\new_[9961]_  | ~\new_[13206]_ ;
  assign \new_[9405]_  = \\u1_u3_rx_ack_to_cnt_reg[3] ;
  assign \new_[9406]_  = ~\new_[9947]_  & (~\new_[14185]_  | ~\new_[13297]_ );
  assign \new_[9407]_  = (~\new_[10778]_  | ~\new_[6250]_ ) & (~\new_[10341]_  | ~\new_[6743]_ );
  assign \new_[9408]_  = (~\new_[10780]_  | ~\new_[5998]_ ) & (~\new_[10340]_  | ~\new_[6593]_ );
  assign \new_[9409]_  = (~\new_[10981]_  | ~\new_[6003]_ ) & (~\new_[10338]_  | ~\new_[6690]_ );
  assign \new_[9410]_  = (~\new_[10779]_  | ~\new_[6008]_ ) & (~\new_[10326]_  | ~\new_[6809]_ );
  assign \new_[9411]_  = ~\\u4_u0_buf0_orig_m3_reg[4] ;
  assign \new_[9412]_  = \\u1_u3_rx_ack_to_cnt_reg[2] ;
  assign \new_[9413]_  = ~\\u4_u0_buf0_orig_m3_reg[2] ;
  assign \new_[9414]_  = ~\new_[9649]_ ;
  assign \new_[9415]_  = ~u1_u3_buf1_not_aloc_reg;
  assign \new_[9416]_  = u1_u3_buf0_not_aloc_reg;
  assign \new_[9417]_  = ~\\u4_u0_buf0_orig_m3_reg[5] ;
  assign \new_[9418]_  = ~\\u4_u1_buf0_orig_m3_reg[5] ;
  assign \new_[9419]_  = ~\\u4_u3_buf0_orig_m3_reg[6] ;
  assign \new_[9420]_  = ~\\u4_u2_buf0_orig_m3_reg[5] ;
  assign \new_[9421]_  = \\u1_u3_rx_ack_to_cnt_reg[6] ;
  assign \new_[9422]_  = ~\new_[9656]_ ;
  assign n7850 = n8055 | \new_[14037]_ ;
  assign \new_[9424]_  = \\u1_u3_rx_ack_to_cnt_reg[0] ;
  assign \new_[9425]_  = \new_[13167]_  | \new_[9995]_ ;
  assign \new_[9426]_  = \new_[13047]_  | \new_[9995]_ ;
  assign \new_[9427]_  = ~\new_[10291]_  & (~\new_[10040]_  | ~\new_[10802]_ );
  assign \new_[9428]_  = \new_[9994]_  | \new_[13427]_ ;
  assign \new_[9429]_  = \new_[9994]_  | \new_[13047]_ ;
  assign \new_[9430]_  = \new_[13047]_  | \new_[9934]_ ;
  assign \new_[9431]_  = ~\new_[11942]_  | ~\new_[9991]_ ;
  assign \new_[9432]_  = ~\new_[9994]_  & ~\new_[13116]_ ;
  assign \new_[9433]_  = \new_[13427]_  | \new_[9995]_ ;
  assign \new_[9434]_  = ~\new_[9934]_  & ~\new_[13167]_ ;
  assign n7800 = ~\new_[10851]_  & ~n7980;
  assign \new_[9436]_  = \new_[9934]_  | \new_[13427]_ ;
  assign \new_[9437]_  = ~\new_[9782]_  | ~\new_[10285]_ ;
  assign n7820 = ~\new_[11452]_  & ~n7980;
  assign n7890 = ~\new_[11017]_  & ~n7980;
  assign \new_[9440]_  = \new_[11638]_  | \new_[10005]_ ;
  assign \new_[9441]_  = ~\new_[9934]_  & ~\new_[13116]_ ;
  assign \new_[9442]_  = \\u1_u3_rx_ack_to_cnt_reg[1] ;
  assign \new_[9443]_  = \new_[9755]_  | \new_[13427]_ ;
  assign \new_[9444]_  = ~\new_[9995]_  & ~\new_[13116]_ ;
  assign \new_[9445]_  = \new_[9755]_  | \new_[13047]_ ;
  assign \new_[9446]_  = ~\new_[9978]_  | ~\new_[13238]_ ;
  assign \new_[9447]_  = ~\new_[9755]_  & ~\new_[13116]_ ;
  assign \new_[9448]_  = \new_[13167]_  | \new_[9755]_ ;
  assign \new_[9449]_  = ~\new_[12814]_  | ~\new_[9983]_  | ~\new_[10505]_ ;
  assign \new_[9450]_  = ~\new_[13027]_  | ~\new_[9984]_  | ~\new_[10502]_ ;
  assign \new_[9451]_  = ~\new_[9696]_ ;
  assign \new_[9452]_  = ~\new_[9797]_  & (~\new_[10745]_  | ~\new_[11531]_ );
  assign \new_[9453]_  = ~\new_[9798]_  & (~\new_[10747]_  | ~\new_[11519]_ );
  assign n7835 = ~\new_[10004]_  | (~\new_[10381]_  & ~\new_[6304]_ );
  assign n7840 = ~\new_[9985]_  | (~\new_[10383]_  & ~\new_[6512]_ );
  assign \new_[9456]_  = \\u1_u3_rx_ack_to_cnt_reg[7] ;
  assign \new_[9457]_  = ~\new_[10479]_  | ~\new_[2301]_  | ~\new_[9812]_  | ~\new_[10097]_ ;
  assign \new_[9458]_  = ~\new_[13279]_  | ~\new_[13344]_  | ~\new_[10072]_ ;
  assign n7845 = \new_[6560]_  ^ \new_[10043]_ ;
  assign \new_[9460]_  = ~\new_[11193]_  | (~\new_[10318]_  & ~\new_[11514]_ );
  assign n7805 = \new_[6234]_  ^ \new_[10262]_ ;
  assign \new_[9462]_  = u4_u3_dma_req_in_hold_reg;
  assign \new_[9463]_  = ~\new_[9812]_  | ~\new_[13655]_ ;
  assign \new_[9464]_  = ~\new_[14331]_  | ~\new_[4838]_ ;
  assign \new_[9465]_  = ~\new_[14331]_  | ~\new_[4608]_ ;
  assign \new_[9466]_  = ~\new_[14331]_  | ~\new_[4841]_ ;
  assign \new_[9467]_  = ~\new_[14331]_  | ~\new_[4616]_ ;
  assign \new_[9468]_  = ~\new_[9785]_  | ~\new_[7206]_ ;
  assign \new_[9469]_  = \new_[9782]_  | \new_[2611]_ ;
  assign n7810 = \new_[6323]_  ^ \new_[10264]_ ;
  assign \new_[9471]_  = \\u1_u3_rx_ack_to_cnt_reg[5] ;
  assign \new_[9472]_  = ~\new_[9798]_  | ~\new_[12028]_ ;
  assign \new_[9473]_  = ~\new_[10590]_  | ~\new_[9870]_ ;
  assign \new_[9474]_  = ~\new_[9802]_  | ~\new_[6198]_ ;
  assign \new_[9475]_  = \\u0_u0_idle_cnt1_next_reg[7] ;
  assign \new_[9476]_  = ~\new_[9812]_  | ~\new_[2392]_ ;
  assign \new_[9477]_  = ~\new_[9806]_  | ~\new_[10939]_ ;
  assign \new_[9478]_  = ~\new_[13407]_  | ~\new_[14230]_  | ~\new_[11430]_ ;
  assign \new_[9479]_  = ~\new_[2372]_  | ~\new_[9812]_  | ~\new_[10097]_ ;
  assign \new_[9480]_  = ~\new_[4794]_  | (~\new_[10075]_  & ~\new_[13740]_ );
  assign \new_[9481]_  = ~\new_[9789]_  & ~\new_[12457]_ ;
  assign \new_[9482]_  = ~\new_[9801]_  | ~\new_[6092]_ ;
  assign \new_[9483]_  = ~\new_[9797]_  | ~\new_[12188]_ ;
  assign \new_[9484]_  = ~\new_[11229]_  | ~\new_[10478]_  | ~\new_[12082]_  | ~\new_[10073]_ ;
  assign \new_[9485]_  = ~\new_[12954]_  & (~\new_[10077]_  | ~\new_[10842]_ );
  assign \new_[9486]_  = ~\new_[13107]_  & (~\new_[10078]_  | ~\new_[10834]_ );
  assign n7865 = \new_[10444]_  & \new_[9787]_ ;
  assign \new_[9488]_  = ~\new_[9782]_  & (~\new_[12467]_  | ~\new_[11658]_ );
  assign \new_[9489]_  = ~\new_[13253]_  & (~\new_[10082]_  | ~\new_[10889]_ );
  assign \new_[9490]_  = ~\new_[9787]_  | ~\new_[12415]_ ;
  assign \new_[9491]_  = (~\new_[10448]_  | ~\new_[13187]_ ) & (~\new_[10813]_  | ~\new_[2611]_ );
  assign \new_[9492]_  = \new_[2876]_  ^ \new_[10707]_ ;
  assign \new_[9493]_  = (~\new_[10463]_  | ~\new_[12573]_ ) & (~\new_[8810]_  | ~\new_[13415]_ );
  assign \new_[9494]_  = ~\new_[10027]_  & (~\new_[13897]_  | ~\new_[3788]_ );
  assign n7950 = \new_[6346]_  ^ \new_[10443]_ ;
  assign n7945 = ~\new_[9807]_ ;
  assign \new_[9497]_  = ~u4_pid_cs_err_r_reg;
  assign n7965 = ~\new_[12849]_  & (~\new_[10843]_  | ~\new_[10596]_ );
  assign \new_[9499]_  = ~\new_[10084]_  | ~\new_[11153]_ ;
  assign \new_[9500]_  = ~\new_[10806]_  & ~\new_[14135]_ ;
  assign \new_[9501]_  = ~\new_[14344]_ ;
  assign \new_[9502]_  = ~\new_[11099]_  & ~\new_[10827]_ ;
  assign \new_[9503]_  = ~\new_[10083]_  | ~\new_[11325]_ ;
  assign \new_[9504]_  = ~\new_[11093]_  & ~\new_[10827]_ ;
  assign \new_[9505]_  = ~\new_[11100]_  & ~\new_[10827]_ ;
  assign \new_[9506]_  = \new_[14060]_  | \new_[10096]_ ;
  assign \new_[9507]_  = ~\new_[11693]_  & ~\new_[10827]_ ;
  assign \new_[9508]_  = ~\new_[11471]_  & ~\new_[10827]_ ;
  assign \new_[9509]_  = \new_[10069]_  & \new_[11688]_ ;
  assign \new_[9510]_  = ~\new_[9789]_ ;
  assign \new_[9511]_  = \new_[11126]_  & \new_[10081]_ ;
  assign \new_[9512]_  = ~\new_[12695]_  | ~\new_[13281]_  | ~\new_[10621]_ ;
  assign \new_[9513]_  = ~\new_[11119]_  | ~\new_[11118]_  | ~\new_[10478]_ ;
  assign \new_[9514]_  = ~\new_[11101]_  & ~\new_[10827]_ ;
  assign \new_[9515]_  = ~\new_[11474]_  & ~\new_[10827]_ ;
  assign \new_[9516]_  = \new_[10085]_  & \new_[11707]_ ;
  assign \new_[9517]_  = ~\new_[9191]_  & ~\new_[10089]_ ;
  assign \new_[9518]_  = ~\new_[10083]_  | ~\new_[11589]_ ;
  assign \new_[9519]_  = \new_[10098]_  | \new_[11232]_ ;
  assign \new_[9520]_  = \new_[11117]_  & \new_[10091]_ ;
  assign \new_[9521]_  = ~\new_[10948]_  & ~\new_[10261]_ ;
  assign \new_[9522]_  = ~\new_[14832]_  | ~\new_[4923]_ ;
  assign \new_[9523]_  = ~\new_[14389]_ ;
  assign \new_[9524]_  = ~\new_[13267]_  | ~\new_[13744]_  | ~\new_[10076]_  | ~\new_[12570]_ ;
  assign n7955 = \new_[10094]_  & \new_[13250]_ ;
  assign \new_[9526]_  = ~\new_[10080]_  & ~\new_[10855]_ ;
  assign n7960 = \new_[10093]_  & \new_[13232]_ ;
  assign \new_[9528]_  = ~n8390 | ~\new_[11430]_  | ~\new_[11801]_ ;
  assign \new_[9529]_  = ~\new_[2857]_  | ~\new_[14830]_  | ~\new_[10490]_ ;
  assign \new_[9530]_  = \new_[4073]_  ^ \new_[10682]_ ;
  assign \new_[9531]_  = ~\new_[9812]_ ;
  assign \new_[9532]_  = ~\new_[9817]_ ;
  assign \new_[9533]_  = (~\new_[12345]_  | ~\new_[10480]_ ) & (~n9145 | ~\new_[13601]_ );
  assign \new_[9534]_  = ~\new_[10556]_  | ~\new_[10956]_  | ~\new_[10906]_ ;
  assign \new_[9535]_  = ~\new_[10558]_  | ~\new_[10886]_  | ~\new_[11274]_ ;
  assign \new_[9536]_  = ~\new_[10560]_  | ~\new_[10895]_  | ~\new_[11251]_ ;
  assign \new_[9537]_  = ~\new_[10535]_  | ~\new_[10913]_  | ~\new_[11280]_ ;
  assign \new_[9538]_  = ~\new_[10543]_  | ~\new_[10760]_  | ~\new_[11281]_ ;
  assign \new_[9539]_  = ~\new_[10537]_  | ~\new_[10885]_  | ~\new_[10891]_ ;
  assign \new_[9540]_  = ~\new_[10524]_  | ~\new_[11249]_  | ~\new_[10904]_ ;
  assign \new_[9541]_  = ~\new_[10512]_  | ~\new_[10887]_  | ~\new_[10892]_ ;
  assign \new_[9542]_  = ~\new_[10527]_  | ~\new_[10789]_  | ~\new_[10883]_ ;
  assign \new_[9543]_  = ~\new_[10530]_  | ~\new_[10899]_  | ~\new_[10876]_ ;
  assign \new_[9544]_  = ~\new_[10548]_  | ~\new_[10907]_  | ~\new_[10911]_ ;
  assign \new_[9545]_  = ~\new_[10542]_  | ~\new_[10999]_  | ~\new_[11369]_ ;
  assign \new_[9546]_  = ~\new_[10488]_  | ~\new_[10426]_  | ~\new_[10487]_ ;
  assign \new_[9547]_  = ~\new_[10510]_  | ~\new_[11265]_  | ~\new_[10903]_ ;
  assign \new_[9548]_  = ~\new_[10544]_  | ~\new_[10593]_  | ~\new_[11270]_ ;
  assign \new_[9549]_  = ~\new_[10521]_  | ~\new_[10890]_  | ~\new_[11259]_ ;
  assign \new_[9550]_  = ~\new_[10873]_  | ~\new_[10266]_  | ~\new_[10880]_ ;
  assign \new_[9551]_  = ~\new_[10559]_  | ~\new_[10912]_  | ~\new_[11252]_ ;
  assign \new_[9552]_  = ~\new_[10110]_  & (~\new_[11202]_  | ~\new_[12805]_ );
  assign \new_[9553]_  = ~\new_[10111]_  & (~\new_[12061]_  | ~\new_[11205]_ );
  assign \new_[9554]_  = \new_[4288]_  ^ \new_[10470]_ ;
  assign \new_[9555]_  = \new_[3476]_  ^ \new_[10471]_ ;
  assign \new_[9556]_  = \new_[3882]_  ^ \new_[10472]_ ;
  assign \new_[9557]_  = \new_[3638]_  ^ \new_[10473]_ ;
  assign \new_[9558]_  = ~\new_[10116]_  & ~\new_[13978]_ ;
  assign \new_[9559]_  = ~\new_[14834]_  & ~\new_[13568]_ ;
  assign \new_[9560]_  = \new_[14409]_  & \new_[2869]_ ;
  assign \new_[9561]_  = ~\new_[10129]_  | ~\new_[14664]_ ;
  assign \new_[9562]_  = \new_[11298]_  | \new_[10936]_  | \new_[10938]_  | \new_[10937]_ ;
  assign \new_[9563]_  = ~\new_[10221]_  & ~\new_[4852]_ ;
  assign \new_[9564]_  = ~\new_[10160]_  | ~\new_[10554]_ ;
  assign \new_[9565]_  = ~\new_[9910]_ ;
  assign \new_[9566]_  = \new_[11116]_  & \new_[10262]_ ;
  assign \new_[9567]_  = ~\new_[10117]_  | ~\new_[2278]_ ;
  assign \new_[9568]_  = ~\new_[10242]_  | ~\new_[10553]_ ;
  assign n7590 = ~\new_[12383]_  & ~\new_[10125]_ ;
  assign \new_[9570]_  = ~\new_[10216]_  | ~\new_[10539]_ ;
  assign \new_[9571]_  = ~\new_[10217]_  | ~\new_[10872]_ ;
  assign \new_[9572]_  = ~\new_[10243]_  | ~\new_[10871]_ ;
  assign \new_[9573]_  = ~\new_[10154]_  | ~\new_[10549]_ ;
  assign \new_[9574]_  = ~\new_[12605]_  & ~\new_[10277]_ ;
  assign \new_[9575]_  = ~\new_[10284]_  & ~\new_[13297]_ ;
  assign \new_[9576]_  = ~\new_[9857]_ ;
  assign n7900 = ~\new_[9837]_ ;
  assign \new_[9578]_  = \new_[10128]_  | \new_[13012]_ ;
  assign \new_[9579]_  = ~\new_[10190]_  | (~\new_[13440]_  & ~\new_[13047]_ );
  assign \new_[9580]_  = ~\new_[10145]_  | (~\new_[6309]_  & ~\new_[13047]_ );
  assign \new_[9581]_  = ~\new_[10263]_  | ~\new_[10201]_ ;
  assign \new_[9582]_  = ~\new_[10197]_  | (~\new_[6559]_  & ~\new_[13047]_ );
  assign \new_[9583]_  = ~\new_[10600]_  | ~\new_[10127]_ ;
  assign \new_[9584]_  = ~\new_[10141]_  | (~\new_[6270]_  & ~\new_[13047]_ );
  assign \new_[9585]_  = ~\new_[10239]_  | (~\new_[7310]_  & ~\new_[13047]_ );
  assign \new_[9586]_  = ~\new_[10267]_  | ~\new_[10235]_ ;
  assign \new_[9587]_  = ~TxValid_pad_o | ~\new_[10103]_  | ~\new_[13842]_ ;
  assign \new_[9588]_  = ~\new_[10206]_  | (~\new_[6564]_  & ~\new_[13047]_ );
  assign \new_[9589]_  = ~\new_[10097]_ ;
  assign \new_[9590]_  = ~\new_[10107]_  & (~\new_[12711]_  | ~\new_[12566]_ );
  assign \new_[9591]_  = ~\new_[10246]_  | ~\new_[13238]_ ;
  assign \new_[9592]_  = ~\new_[13365]_  | ~\new_[10274]_  | ~\new_[12438]_ ;
  assign \new_[9593]_  = ~\new_[10271]_  & (~\new_[3038]_  | ~\new_[13297]_ );
  assign \new_[9594]_  = ~\new_[14582]_  | ~\new_[10289]_  | ~\new_[13424]_ ;
  assign \new_[9595]_  = ~\new_[9889]_ ;
  assign \new_[9596]_  = \new_[4092]_  & n7980;
  assign \new_[9597]_  = \new_[4291]_  ^ \new_[10675]_ ;
  assign \new_[9598]_  = \new_[3480]_  ^ \new_[10676]_ ;
  assign \new_[9599]_  = \new_[3691]_  ^ \new_[10678]_ ;
  assign \new_[9600]_  = ~\new_[13011]_  | ~\new_[10276]_  | ~\new_[12445]_ ;
  assign \new_[9601]_  = \new_[3884]_  ^ \new_[10679]_ ;
  assign \new_[9602]_  = \new_[3881]_  & n7980;
  assign \new_[9603]_  = ~\new_[9955]_ ;
  assign n7735 = ~\new_[9836]_ ;
  assign \new_[9605]_  = ~\new_[10258]_  & (~\new_[12591]_  | ~\new_[4709]_ );
  assign n7940 = \new_[6345]_  ^ \new_[10677]_ ;
  assign \new_[9607]_  = \new_[3025]_  ? \new_[10715]_  : \new_[10666]_ ;
  assign \new_[9608]_  = ~\\u4_u3_buf0_orig_m3_reg[3] ;
  assign \new_[9609]_  = ~\\u4_u2_buf0_orig_m3_reg[3] ;
  assign \new_[9610]_  = ~\new_[9834]_ ;
  assign \new_[9611]_  = u1_u3_buf0_rl_reg;
  assign \new_[9612]_  = ~\new_[10319]_  & ~\new_[13297]_ ;
  assign \new_[9613]_  = \new_[2347]_  ^ \new_[10654]_ ;
  assign \new_[9614]_  = ~\new_[10288]_  | (~\new_[10973]_  & ~\new_[13819]_ );
  assign \new_[9615]_  = \new_[3469]_  ^ \new_[10657]_ ;
  assign \new_[9616]_  = ~\new_[10297]_  | ~\new_[14195]_ ;
  assign \new_[9617]_  = ~\new_[10299]_  | ~\new_[11841]_ ;
  assign \new_[9618]_  = ~\new_[10296]_  | ~\new_[13914]_ ;
  assign \new_[9619]_  = ~\new_[10301]_  | ~\new_[11849]_ ;
  assign \new_[9620]_  = ~\new_[9824]_ ;
  assign \new_[9621]_  = ~\new_[10295]_  | ~\new_[13980]_ ;
  assign \new_[9622]_  = ~\new_[10304]_  | ~\new_[11862]_ ;
  assign \new_[9623]_  = ~\new_[10298]_  | ~\new_[13617]_ ;
  assign \new_[9624]_  = ~\new_[10303]_  | ~\new_[11871]_ ;
  assign \new_[9625]_  = (~\new_[10686]_  | ~\new_[12610]_ ) & (~\new_[11014]_  | ~\new_[12124]_ );
  assign n7910 = ~\new_[9935]_ ;
  assign \new_[9627]_  = \\u0_u0_idle_cnt1_next_reg[6] ;
  assign \new_[9628]_  = ~\\u4_u3_dma_out_left_reg[3] ;
  assign \new_[9629]_  = ~\\u4_u0_dma_out_left_reg[3] ;
  assign \new_[9630]_  = ~\\u4_u1_dma_out_left_reg[3] ;
  assign \new_[9631]_  = ~\\u4_u2_dma_out_left_reg[3] ;
  assign \new_[9632]_  = ~\new_[10315]_  & (~\new_[3037]_  | ~\new_[13297]_ );
  assign \new_[9633]_  = ~\new_[11081]_  | ~\new_[10750]_  | ~\new_[11835]_  | ~\new_[13123]_ ;
  assign \new_[9634]_  = ~\new_[11319]_  | ~\new_[10749]_  | ~\new_[12118]_  | ~\new_[12908]_ ;
  assign \new_[9635]_  = ~\new_[10302]_  | (~\new_[10992]_  & ~\new_[13666]_ );
  assign n7905 = \new_[3174]_  ? n9145 : \new_[2836]_ ;
  assign \new_[9637]_  = ~\new_[10048]_  & ~\new_[11799]_ ;
  assign \new_[9638]_  = \new_[3481]_  ^ \new_[10684]_ ;
  assign \new_[9639]_  = ~\new_[12678]_  | ~\new_[11517]_  | ~\new_[10680]_ ;
  assign \new_[9640]_  = ~\new_[10378]_  | ~\new_[10014]_ ;
  assign \new_[9641]_  = \\u0_u0_idle_cnt1_next_reg[4] ;
  assign \new_[9642]_  = \new_[6736]_  ^ \new_[10357]_ ;
  assign \new_[9643]_  = \new_[2084]_  ^ \new_[10354]_ ;
  assign \new_[9644]_  = ~\\u4_u3_buf0_orig_m3_reg[4] ;
  assign \new_[9645]_  = u0_u0_me_ps2_0_5_ms_reg;
  assign \new_[9646]_  = ~\\u4_u2_buf0_orig_m3_reg[4] ;
  assign \new_[9647]_  = \new_[3688]_  ^ \new_[10709]_ ;
  assign \new_[9648]_  = \new_[14036]_  ? \new_[10715]_  : \new_[10356]_ ;
  assign \new_[9649]_  = ~\\u4_u2_buf0_orig_m3_reg[2] ;
  assign \new_[9650]_  = ~\new_[9946]_ ;
  assign \new_[9651]_  = ~\\u4_u3_buf0_orig_m3_reg[5] ;
  assign \new_[9652]_  = ~\new_[9939]_ ;
  assign \new_[9653]_  = ~\new_[10101]_  | (~\new_[12361]_  & ~\new_[10399]_ );
  assign \new_[9654]_  = ~\new_[2342]_  & ~\new_[14273]_ ;
  assign \new_[9655]_  = ~\new_[10191]_  | (~\new_[13264]_  & ~\new_[13047]_ );
  assign \new_[9656]_  = \new_[14273]_  | \new_[14314]_ ;
  assign \new_[9657]_  = ~\new_[10048]_  | (~\new_[10387]_  & ~\new_[11321]_ );
  assign \new_[9658]_  = ~\new_[10049]_  | (~\new_[10404]_  & ~\new_[11151]_ );
  assign \new_[9659]_  = ~\new_[10053]_  | (~\new_[10394]_  & ~\new_[11231]_ );
  assign \new_[9660]_  = ~\new_[10057]_  | (~\new_[10397]_  & ~\new_[11134]_ );
  assign \new_[9661]_  = ~\new_[12509]_  | ~\new_[13462]_  | ~\new_[10583]_ ;
  assign \new_[9662]_  = ~\new_[10292]_  & (~\new_[10497]_  | ~\new_[11911]_ );
  assign \new_[9663]_  = ~\new_[12520]_  & ~\new_[10248]_ ;
  assign \new_[9664]_  = ~\new_[12420]_  | ~\new_[10285]_ ;
  assign \new_[9665]_  = ~\new_[10341]_  & ~\new_[6743]_ ;
  assign \new_[9666]_  = \new_[11629]_  | \new_[10345]_ ;
  assign \new_[9667]_  = ~\new_[10120]_  & ~\new_[13297]_ ;
  assign \new_[9668]_  = ~\new_[12701]_  | ~\new_[13485]_  | ~\new_[10605]_ ;
  assign \new_[9669]_  = ~\new_[10344]_  | ~\new_[10849]_ ;
  assign \new_[9670]_  = \new_[11619]_  | \new_[10348]_ ;
  assign \new_[9671]_  = ~\new_[10018]_  | ~\new_[11854]_ ;
  assign \new_[9672]_  = ~\new_[12787]_  | ~\new_[13435]_  | ~\new_[10614]_ ;
  assign \new_[9673]_  = ~\new_[10340]_  & ~\new_[6593]_ ;
  assign \new_[9674]_  = ~\new_[10338]_  & ~\new_[6690]_ ;
  assign \new_[9675]_  = ~\new_[10236]_  | (~\new_[6245]_  & ~\new_[13047]_ );
  assign \new_[9676]_  = \new_[3316]_  ^ \new_[10683]_ ;
  assign \new_[9677]_  = ~\new_[10016]_  | ~\new_[11865]_ ;
  assign \new_[9678]_  = ~\new_[10326]_  & ~\new_[6809]_ ;
  assign \new_[9679]_  = \new_[11485]_  | \new_[10342]_ ;
  assign \new_[9680]_  = ~\new_[10047]_  | (~\new_[10737]_  & ~\new_[11131]_ );
  assign \new_[9681]_  = ~\new_[10052]_  | (~\new_[10735]_  & ~\new_[11144]_ );
  assign \new_[9682]_  = ~\new_[10055]_  | (~\new_[10736]_  & ~\new_[11127]_ );
  assign \new_[9683]_  = ~\new_[10058]_  | (~\new_[10738]_  & ~\new_[11129]_ );
  assign \new_[9684]_  = ~\new_[12117]_  | (~\new_[10384]_  & ~\new_[12318]_ );
  assign \new_[9685]_  = ~\new_[10015]_  & (~\new_[11839]_  | ~\new_[12322]_ );
  assign n7935 = ~\new_[10339]_  | ~\new_[10327]_ ;
  assign \new_[9687]_  = \new_[3693]_  ^ \new_[10685]_ ;
  assign \new_[9688]_  = ~\new_[11857]_  | (~\new_[10391]_  & ~\new_[12407]_ );
  assign \new_[9689]_  = ~\new_[10019]_  & (~\new_[11860]_  | ~\new_[12054]_ );
  assign \new_[9690]_  = ~\new_[10017]_  & (~\new_[11845]_  | ~\new_[12394]_ );
  assign \new_[9691]_  = ~\new_[11851]_  | (~\new_[10401]_  & ~\new_[12234]_ );
  assign \new_[9692]_  = ~\new_[11834]_  | (~\new_[10385]_  & ~\new_[12230]_ );
  assign \new_[9693]_  = ~\new_[10020]_  & (~\new_[11868]_  | ~\new_[12005]_ );
  assign \new_[9694]_  = ~\new_[9959]_ ;
  assign \new_[9695]_  = ~\new_[9960]_ ;
  assign \new_[9696]_  = ~\new_[11834]_  | ~\new_[10349]_  | ~\new_[11085]_ ;
  assign \new_[9697]_  = ~\new_[9961]_ ;
  assign \new_[9698]_  = ~\new_[11545]_  | (~\new_[10390]_  & ~\new_[12289]_ );
  assign \new_[9699]_  = ~\new_[11538]_  | (~\new_[10389]_  & ~\new_[12301]_ );
  assign \new_[9700]_  = ~\new_[11544]_  | (~\new_[10400]_  & ~\new_[12292]_ );
  assign \new_[9701]_  = ~\new_[11539]_  | (~\new_[10405]_  & ~\new_[12282]_ );
  assign \new_[9702]_  = ~\new_[10045]_  & (~\new_[10739]_  | ~\new_[11532]_ );
  assign \new_[9703]_  = ~\new_[10037]_  & (~\new_[10741]_  | ~\new_[11529]_ );
  assign \new_[9704]_  = \new_[3475]_  ^ \new_[10582]_ ;
  assign \new_[9705]_  = \new_[12254]_  ^ \new_[10387]_ ;
  assign n7915 = \new_[6303]_  ^ \new_[10571]_ ;
  assign \new_[9707]_  = \new_[11614]_  ^ \new_[10394]_ ;
  assign \new_[9708]_  = \new_[4347]_  ^ \new_[10583]_ ;
  assign \new_[9709]_  = \new_[11610]_  ^ \new_[10397]_ ;
  assign \new_[9710]_  = \new_[12286]_  ^ \new_[10404]_ ;
  assign \new_[9711]_  = \new_[3478]_  ^ \new_[10605]_ ;
  assign \new_[9712]_  = \new_[3689]_  ^ \new_[10614]_ ;
  assign n7920 = \new_[6371]_  ^ \new_[10618]_ ;
  assign \new_[9714]_  = u4_u2_dma_req_out_hold_reg;
  assign \new_[9715]_  = u4_u3_dma_req_out_hold_reg;
  assign \new_[9716]_  = \new_[3815]_  ^ \new_[10621]_ ;
  assign \new_[9717]_  = u4_u0_dma_req_out_hold_reg;
  assign \new_[9718]_  = u4_u1_dma_req_out_hold_reg;
  assign \new_[9719]_  = ~\new_[10122]_  | ~\new_[11048]_ ;
  assign \new_[9720]_  = ~\new_[10114]_  | ~\new_[11049]_ ;
  assign \new_[9721]_  = ~\new_[10029]_  & ~\new_[13771]_ ;
  assign \new_[9722]_  = ~\new_[14533]_  | ~\new_[4709]_ ;
  assign \new_[9723]_  = ~\new_[14533]_  | ~\new_[4818]_ ;
  assign n7925 = \new_[6853]_  ^ \new_[10617]_ ;
  assign \new_[9725]_  = \new_[4236]_  ^ \new_[10575]_ ;
  assign \new_[9726]_  = \new_[3428]_  ^ \new_[10606]_ ;
  assign \new_[9727]_  = \new_[3684]_  ^ \new_[10615]_ ;
  assign \new_[9728]_  = ~\new_[10045]_  | ~\new_[12327]_ ;
  assign n7930 = \new_[6091]_  ^ \new_[10619]_ ;
  assign \new_[9730]_  = \new_[10047]_  | \new_[11503]_ ;
  assign \new_[9731]_  = \new_[3875]_  ^ \new_[10569]_ ;
  assign \new_[9732]_  = ~\new_[10577]_  | ~\new_[10169]_ ;
  assign \new_[9733]_  = ~\new_[10732]_  | ~\new_[10849]_ ;
  assign \new_[9734]_  = ~\new_[10030]_  | ~\new_[10849]_ ;
  assign \new_[9735]_  = ~\new_[10031]_  | ~\new_[10849]_ ;
  assign \new_[9736]_  = ~\new_[10050]_  | ~\new_[10849]_ ;
  assign \new_[9737]_  = ~\new_[10580]_  | ~\new_[10165]_ ;
  assign \new_[9738]_  = ~\new_[10270]_  | ~n8390;
  assign \new_[9739]_  = ~\new_[10037]_  | ~\new_[11976]_ ;
  assign \new_[9740]_  = ~\new_[14533]_  | ~\new_[4695]_ ;
  assign \new_[9741]_  = \new_[10052]_  | \new_[11141]_ ;
  assign \new_[9742]_  = ~\new_[10053]_  & ~\new_[11808]_ ;
  assign n7970 = ~\new_[12849]_  & (~\new_[10576]_  | ~\new_[11702]_ );
  assign \new_[9744]_  = \new_[10055]_  | \new_[12029]_ ;
  assign \new_[9745]_  = ~\new_[10057]_  & ~\new_[11803]_ ;
  assign \new_[9746]_  = \new_[10058]_  | \new_[11515]_ ;
  assign \new_[9747]_  = ~\new_[10049]_  & ~\new_[11814]_ ;
  assign \new_[9748]_  = ~\new_[14533]_  | ~\new_[4815]_ ;
  assign \new_[9749]_  = (~\new_[10424]_  & ~\new_[13155]_  & ~\new_[12437]_ ) | (~\new_[11115]_  & ~n8390 & ~\new_[12437]_ );
  assign \new_[9750]_  = ~\new_[12113]_  | ~\new_[13205]_  | ~\new_[10464]_  | ~\new_[10609]_ ;
  assign \new_[9751]_  = (~\new_[12869]_  & ~\new_[3710]_ ) | (~\new_[10419]_  & ~\new_[3930]_ );
  assign \new_[9752]_  = (~\new_[12874]_  & ~\new_[4095]_ ) | (~\new_[10418]_  & ~\new_[4292]_ );
  assign \new_[9753]_  = (~\new_[12862]_  & ~\new_[3337]_ ) | (~\new_[10417]_  & ~\new_[3503]_ );
  assign n8055 = ~\new_[10364]_  & ~\new_[13159]_ ;
  assign \new_[9755]_  = \new_[11488]_  | \new_[10375]_ ;
  assign \new_[9756]_  = ~\new_[10368]_  | (~\new_[11089]_  & ~\new_[3474]_ );
  assign \new_[9757]_  = ~\new_[11570]_  & (~\new_[10996]_  | ~\new_[11637]_ );
  assign \new_[9758]_  = ~\new_[10380]_  | (~\new_[11107]_  & ~\new_[12346]_ );
  assign \new_[9759]_  = \new_[12346]_  ? \new_[10960]_  : \new_[12048]_ ;
  assign \new_[9760]_  = \new_[6716]_  ^ \new_[10824]_ ;
  assign n8060 = \new_[6238]_  ^ \new_[10790]_ ;
  assign n8070 = \new_[6588]_  ^ \new_[10792]_ ;
  assign n8065 = \new_[6551]_  ^ \new_[10800]_ ;
  assign n8075 = \new_[6369]_  ^ \new_[10808]_ ;
  assign n8045 = ~\new_[10051]_ ;
  assign \new_[9766]_  = ~\new_[10420]_  & ~\new_[11201]_ ;
  assign \new_[9767]_  = ~\new_[10421]_  & ~\new_[11198]_ ;
  assign \new_[9768]_  = ~\new_[11200]_  | (~\new_[11171]_  & ~\new_[10841]_ );
  assign \new_[9769]_  = ~\new_[10451]_  & ~\new_[11235]_ ;
  assign \new_[9770]_  = \new_[11093]_  | \new_[11149]_ ;
  assign \new_[9771]_  = ~\new_[10438]_  | ~\new_[10847]_ ;
  assign \new_[9772]_  = \new_[11693]_  | \new_[11149]_ ;
  assign \new_[9773]_  = \new_[11471]_  | \new_[11149]_ ;
  assign \new_[9774]_  = \new_[11474]_  | \new_[11149]_ ;
  assign \new_[9775]_  = \new_[11099]_  | \new_[11149]_ ;
  assign \new_[9776]_  = ~\new_[11153]_  | (~\new_[10759]_  & ~\new_[10847]_ );
  assign \new_[9777]_  = \new_[11100]_  | \new_[11149]_ ;
  assign \new_[9778]_  = \new_[11101]_  | \new_[11149]_ ;
  assign \new_[9779]_  = \new_[11106]_  & \new_[2372]_ ;
  assign \new_[9780]_  = ~\new_[11238]_  | ~\new_[12033]_  | ~\new_[11236]_  | ~\new_[11482]_ ;
  assign \new_[9781]_  = ~\new_[10449]_  | ~\new_[11588]_ ;
  assign \new_[9782]_  = ~\new_[6235]_  | ~\new_[10432]_  | ~\new_[14216]_ ;
  assign \new_[9783]_  = ~\new_[10418]_  | ~\new_[4292]_ ;
  assign \new_[9784]_  = ~\new_[11219]_  | ~\new_[12074]_  | ~\new_[11239]_  | ~\new_[11678]_ ;
  assign \new_[9785]_  = ~\new_[10029]_ ;
  assign \new_[9786]_  = ~\new_[11119]_  | ~\new_[10478]_  | ~\new_[11926]_ ;
  assign \new_[9787]_  = ~\new_[10425]_  & ~\new_[11079]_ ;
  assign \new_[9788]_  = ~\new_[13645]_  | ~\new_[10432]_  | ~\new_[13494]_ ;
  assign \new_[9789]_  = ~\new_[3177]_  | ~\new_[13218]_  | ~\new_[10850]_ ;
  assign \new_[9790]_  = ~\new_[10875]_  | ~\new_[11716]_  | ~\new_[10863]_ ;
  assign \new_[9791]_  = ~\new_[10419]_  | ~\new_[3930]_ ;
  assign \new_[9792]_  = ~\new_[11243]_  | ~\new_[12151]_  | ~\new_[10882]_  | ~\new_[11580]_ ;
  assign \new_[9793]_  = \new_[11121]_  & \new_[10443]_ ;
  assign \new_[9794]_  = \new_[10440]_  & \new_[11707]_ ;
  assign \new_[9795]_  = ~\new_[10417]_  | ~\new_[3503]_ ;
  assign \new_[9796]_  = ~\new_[11173]_  | ~\new_[12098]_  | ~\new_[10820]_  | ~\new_[11584]_ ;
  assign \new_[9797]_  = ~\new_[10673]_  | ~\new_[11559]_ ;
  assign \new_[9798]_  = ~\new_[10453]_  | ~\new_[11560]_ ;
  assign \new_[9799]_  = ~\new_[10270]_ ;
  assign \new_[9800]_  = ~\new_[11698]_  & ~\new_[10452]_ ;
  assign \new_[9801]_  = ~\new_[12084]_  | ~\new_[14197]_  | ~\new_[10481]_  | ~\new_[12722]_ ;
  assign \new_[9802]_  = ~\new_[12097]_  | ~\new_[14149]_  | ~\new_[10482]_  | ~\new_[12557]_ ;
  assign \new_[9803]_  = ~\new_[14106]_  | ~\new_[10448]_  | ~\new_[2479]_ ;
  assign \new_[9804]_  = ~\new_[11168]_  | ~\new_[11697]_  | ~\new_[11702]_  | ~\new_[11597]_ ;
  assign \new_[9805]_  = ~\new_[10458]_  & (~\new_[11634]_  | ~\new_[11568]_ );
  assign \new_[9806]_  = ~\new_[10441]_  & ~\new_[11707]_ ;
  assign \new_[9807]_  = \new_[10422]_  & \new_[11067]_ ;
  assign \new_[9808]_  = ~\new_[10837]_  | ~\new_[10844]_  | ~\new_[12364]_ ;
  assign \new_[9809]_  = ~\new_[11705]_  | ~\new_[10844]_  | ~\new_[10837]_ ;
  assign \new_[9810]_  = ~\new_[10457]_  & (~\new_[11639]_  | ~\new_[11564]_ );
  assign \new_[9811]_  = ~\new_[11627]_  & ~\new_[10451]_ ;
  assign \new_[9812]_  = ~\new_[14665]_  & (~\new_[10838]_  | ~\new_[12573]_ );
  assign \new_[9813]_  = ~\new_[6288]_  | ~\new_[10428]_  | ~\new_[12640]_ ;
  assign \new_[9814]_  = ~\new_[6256]_  | ~\new_[10423]_  | ~\new_[12506]_ ;
  assign \new_[9815]_  = ~\new_[6267]_  | ~\new_[10431]_  | ~\new_[12763]_ ;
  assign \new_[9816]_  = ~\new_[6276]_  | ~\new_[10433]_  | ~\new_[12543]_ ;
  assign \new_[9817]_  = ~\new_[13386]_  | ~\new_[12617]_  | ~\new_[10474]_  | ~\new_[11237]_ ;
  assign \new_[9818]_  = ~\new_[10963]_  | ~\new_[10898]_  | ~\new_[10881]_ ;
  assign \new_[9819]_  = ~\new_[12278]_  & (~\new_[10827]_  | ~\new_[11149]_ );
  assign \new_[9820]_  = \new_[11120]_  & \new_[10571]_ ;
  assign \new_[9821]_  = ~\new_[10490]_  | ~\new_[2932]_ ;
  assign \new_[9822]_  = ~\new_[10072]_ ;
  assign \new_[9823]_  = ~\new_[10498]_  | ~\new_[14666]_ ;
  assign \new_[9824]_  = \new_[11294]_  | \new_[11304]_  | \new_[11420]_  | \new_[12035]_ ;
  assign \new_[9825]_  = ~\new_[12404]_  | ~\new_[10494]_  | ~\new_[2193]_ ;
  assign \new_[9826]_  = ~\new_[10080]_ ;
  assign \new_[9827]_  = ~\new_[10596]_  | ~\new_[8626]_ ;
  assign \new_[9828]_  = \new_[10599]_  | \new_[11490]_ ;
  assign n7975 = ~\new_[11145]_  | (~\new_[12782]_  & ~\new_[8959]_ );
  assign \new_[9830]_  = ~\new_[10083]_ ;
  assign n8090 = ~\new_[12876]_  & ~\new_[10629]_ ;
  assign \new_[9832]_  = ~\new_[12404]_  | ~\new_[11324]_  | ~\new_[2210]_ ;
  assign n8085 = ~\new_[10629]_  & ~\new_[9424]_ ;
  assign \new_[9834]_  = \new_[14829]_ ;
  assign \new_[9835]_  = ~\new_[10499]_  | ~\new_[11404]_ ;
  assign \new_[9836]_  = \new_[11742]_  | \new_[11295]_  | \new_[11303]_  | \new_[11302]_ ;
  assign \new_[9837]_  = \new_[11296]_  | \new_[11648]_  | \new_[11299]_  | \new_[11424]_ ;
  assign \new_[9838]_  = \new_[10476]_  & \new_[10825]_ ;
  assign n8095 = ~\new_[10951]_  & ~\new_[10629]_ ;
  assign \new_[9840]_  = ~\new_[11241]_  | ~\new_[14043]_  | ~\new_[11256]_  | ~\new_[13272]_ ;
  assign \new_[9841]_  = ~\new_[10532]_  | (~\new_[14001]_  & ~\new_[13047]_ );
  assign \new_[9842]_  = ~\new_[10477]_  | ~\new_[2452]_ ;
  assign \new_[9843]_  = \new_[10467]_  & \new_[10628]_ ;
  assign \new_[9844]_  = ~\new_[10096]_ ;
  assign \new_[9845]_  = ~\new_[11688]_  | ~\new_[11213]_  | ~\new_[10574]_  | ~\new_[11229]_ ;
  assign \new_[9846]_  = ~u1_u1_send_data_r2_reg;
  assign \new_[9847]_  = ~\new_[13493]_  & ~\new_[10610]_ ;
  assign \new_[9848]_  = ~\new_[13452]_  & ~\new_[10607]_ ;
  assign \new_[9849]_  = ~\new_[10279]_ ;
  assign \new_[9850]_  = ~\new_[10277]_ ;
  assign \new_[9851]_  = ~\new_[11554]_  & (~\new_[10994]_  | ~\new_[11991]_ );
  assign \new_[9852]_  = ~\new_[13778]_  & ~\new_[10893]_ ;
  assign \new_[9853]_  = \new_[12343]_  ? \new_[10817]_  : \new_[12497]_ ;
  assign \new_[9854]_  = \new_[10574]_  & \new_[11688]_ ;
  assign \new_[9855]_  = ~\new_[12932]_  | ~\new_[10611]_  | ~\new_[13460]_ ;
  assign \new_[9856]_  = \new_[14211]_  ^ \new_[10985]_ ;
  assign \new_[9857]_  = ~\new_[10626]_  | ~\new_[6246]_ ;
  assign \new_[9858]_  = (~\new_[13776]_  | ~\new_[11489]_ ) & (~\new_[14234]_  | ~\new_[12970]_ );
  assign \new_[9859]_  = (~\new_[13665]_  | ~\new_[11489]_ ) & (~\new_[13772]_  | ~\new_[12970]_ );
  assign \new_[9860]_  = (~\new_[14235]_  | ~\new_[11476]_ ) & (~\new_[13909]_  | ~\new_[12970]_ );
  assign \new_[9861]_  = (~\new_[13651]_  | ~\new_[11476]_ ) & (~\new_[13890]_  | ~\new_[12970]_ );
  assign \new_[9862]_  = (~\new_[14240]_  | ~\new_[11484]_ ) & (~\new_[13719]_  | ~\new_[12970]_ );
  assign \new_[9863]_  = (~\new_[13566]_  | ~\new_[11489]_ ) & (~\new_[13868]_  | ~\new_[12970]_ );
  assign \new_[9864]_  = (~\new_[13589]_  | ~\new_[11484]_ ) & (~\new_[13701]_  | ~\new_[12970]_ );
  assign \new_[9865]_  = (~\new_[14143]_  | ~\new_[11476]_ ) & (~\new_[14170]_  | ~\new_[12970]_ );
  assign \new_[9866]_  = (~\new_[13984]_  | ~\new_[11489]_ ) & (~\new_[13936]_  | ~\new_[12970]_ );
  assign \new_[9867]_  = (~\new_[13818]_  | ~\new_[11489]_ ) & (~\new_[13952]_  | ~\new_[12970]_ );
  assign \new_[9868]_  = (~\new_[13685]_  | ~\new_[11484]_ ) & (~\new_[13934]_  | ~\new_[12970]_ );
  assign \new_[9869]_  = (~\new_[14112]_  | ~\new_[11476]_ ) & (~\new_[13929]_  | ~\new_[12970]_ );
  assign \new_[9870]_  = (~\new_[14011]_  | ~\new_[11484]_ ) & (~\new_[13528]_  | ~\new_[12970]_ );
  assign \new_[9871]_  = (~\new_[13603]_  | ~\new_[11476]_ ) & (~\new_[13671]_  | ~\new_[12970]_ );
  assign \new_[9872]_  = (~\new_[14114]_  | ~\new_[11476]_ ) & (~\new_[13979]_  | ~\new_[12970]_ );
  assign \new_[9873]_  = (~\new_[14158]_  | ~\new_[11484]_ ) & (~\new_[13869]_  | ~\new_[12970]_ );
  assign \new_[9874]_  = (~\new_[14162]_  | ~\new_[11489]_ ) & (~\new_[13856]_  | ~\new_[12970]_ );
  assign n8035 = \new_[6320]_  ^ \new_[10984]_ ;
  assign \new_[9876]_  = (~\new_[13640]_  | ~\new_[11489]_ ) & (~\new_[13516]_  | ~\new_[12970]_ );
  assign \new_[9877]_  = (~\new_[13775]_  | ~\new_[11484]_ ) & (~\new_[14183]_  | ~\new_[12970]_ );
  assign \new_[9878]_  = (~\new_[10974]_  | ~\new_[11727]_ ) & (~\new_[13315]_  | ~\new_[3471]_ );
  assign \new_[9879]_  = (~\new_[13529]_  | ~\new_[11476]_ ) & (~\new_[14065]_  | ~\new_[12970]_ );
  assign \new_[9880]_  = (~\new_[13806]_  | ~\new_[11484]_ ) & (~\new_[14145]_  | ~\new_[12970]_ );
  assign \new_[9881]_  = \new_[11990]_  ^ \new_[10739]_ ;
  assign \new_[9882]_  = \new_[2857]_  ^ \new_[10965]_ ;
  assign \new_[9883]_  = ~\new_[11553]_  & (~\new_[10991]_  | ~\new_[11620]_ );
  assign \new_[9884]_  = \new_[2089]_  ^ \new_[10966]_ ;
  assign \new_[9885]_  = ~\new_[13221]_  | ~\new_[10613]_  | ~\new_[12446]_ ;
  assign \new_[9886]_  = ~\new_[11301]_  & ~\new_[10696]_ ;
  assign \new_[9887]_  = \new_[12459]_  & \new_[10679]_ ;
  assign \new_[9888]_  = \new_[12481]_  & \new_[10675]_ ;
  assign \new_[9889]_  = ~\new_[4091]_  & ~\new_[10893]_ ;
  assign \new_[9890]_  = ~u4_usb_reset_r_reg;
  assign \new_[9891]_  = \new_[12410]_  & \new_[10676]_ ;
  assign \new_[9892]_  = \new_[2876]_  ^ \new_[4651]_ ;
  assign \new_[9893]_  = \new_[12107]_  & \new_[10677]_ ;
  assign \new_[9894]_  = \new_[9372]_  ^ \new_[8959]_ ;
  assign \new_[9895]_  = \new_[11272]_  & \new_[10677]_ ;
  assign \new_[9896]_  = \new_[2875]_  ^ \new_[4801]_ ;
  assign \new_[9897]_  = \new_[8658]_  ^ \new_[8959]_ ;
  assign n8030 = ~\new_[11395]_  & ~\new_[10629]_ ;
  assign \new_[9899]_  = ~\new_[10454]_  & (~\new_[11635]_  | ~\new_[11204]_ );
  assign \new_[9900]_  = \new_[9471]_  ^ \new_[8959]_ ;
  assign \new_[9901]_  = \new_[8954]_  ^ \new_[8959]_ ;
  assign \new_[9902]_  = \new_[12166]_  & \new_[10678]_ ;
  assign \new_[9903]_  = ~\new_[10278]_ ;
  assign \new_[9904]_  = ~\new_[10650]_  & ~\new_[13378]_ ;
  assign \new_[9905]_  = ~\new_[4073]_  | ~\new_[10675]_  | ~\new_[13268]_ ;
  assign \new_[9906]_  = ~\new_[3316]_  | ~\new_[10676]_  | ~\new_[13466]_ ;
  assign \new_[9907]_  = ~\new_[10650]_  | ~\new_[3463]_ ;
  assign \new_[9908]_  = ~\new_[3481]_  | ~\new_[10678]_  | ~\new_[12987]_ ;
  assign \new_[9909]_  = ~\new_[3693]_  | ~\new_[10679]_  | ~\new_[13351]_ ;
  assign \new_[9910]_  = ~\new_[10479]_  | ~\new_[12960]_ ;
  assign \new_[9911]_  = ~\new_[13598]_  | ~\new_[13901]_ ;
  assign n8110 = ~\new_[10627]_  | (~\new_[11392]_  & ~\new_[14261]_ );
  assign \new_[9913]_  = \new_[2316]_  ^ \new_[10723]_ ;
  assign \new_[9914]_  = ~\new_[10626]_ ;
  assign \new_[9915]_  = ~\new_[10602]_  & (~\new_[12565]_  | ~\new_[4695]_ );
  assign \new_[9916]_  = u0_u0_idle_cnt1_clr_reg;
  assign n8100 = \new_[10396]_  & \new_[13115]_ ;
  assign n8005 = \new_[12020]_  ^ \new_[10989]_ ;
  assign \new_[9919]_  = \new_[11984]_  ^ \new_[10991]_ ;
  assign n7990 = \new_[11992]_  ^ \new_[10986]_ ;
  assign \new_[9921]_  = \new_[12021]_  ^ \new_[10994]_ ;
  assign n7995 = \new_[12001]_  ^ \new_[10987]_ ;
  assign \new_[9923]_  = \new_[12161]_  ^ \new_[10995]_ ;
  assign n8000 = \new_[11287]_  ^ \new_[10988]_ ;
  assign \new_[9925]_  = \new_[12018]_  ^ \new_[10996]_ ;
  assign n7985 = ~\new_[10306]_ ;
  assign \new_[9927]_  = ~\new_[12176]_  & ~\new_[10682]_ ;
  assign n8080 = ~\new_[10998]_  & ~\new_[10629]_ ;
  assign \new_[9929]_  = ~\new_[12611]_  & ~\new_[10683]_ ;
  assign \new_[9930]_  = ~\new_[11546]_  & (~\new_[10995]_  | ~\new_[12051]_ );
  assign \new_[9931]_  = ~\new_[11964]_  & ~\new_[10685]_ ;
  assign \new_[9932]_  = ~\new_[10400]_  | ~\new_[10406]_ ;
  assign \new_[9933]_  = ~\new_[12773]_  & ~\new_[10684]_ ;
  assign \new_[9934]_  = \new_[11877]_  | \new_[10375]_ ;
  assign \new_[9935]_  = ~\new_[10677]_  & (~\new_[11067]_  | ~\new_[6344]_ );
  assign \new_[9936]_  = \new_[4289]_  ^ \new_[11008]_ ;
  assign \new_[9937]_  = \new_[3477]_  ^ \new_[11010]_ ;
  assign \new_[9938]_  = \new_[3883]_  ^ \new_[10972]_ ;
  assign \new_[9939]_  = \new_[11818]_  | \new_[10680]_ ;
  assign \new_[9940]_  = ~\new_[10386]_  & ~\new_[10355]_ ;
  assign \new_[9941]_  = ~\new_[10429]_  & ~\new_[10716]_ ;
  assign \new_[9942]_  = ~\new_[10392]_  & ~\new_[11013]_ ;
  assign \new_[9943]_  = ~\new_[10388]_  & ~\new_[10717]_ ;
  assign n8105 = ~\new_[11233]_  & ~\new_[10629]_ ;
  assign \new_[9945]_  = ~\new_[3174]_  | ~\new_[13646]_ ;
  assign \new_[9946]_  = ~\\u4_u3_buf0_orig_m3_reg[2] ;
  assign \new_[9947]_  = ~\new_[10566]_  & ~\new_[13297]_ ;
  assign n8010 = ~\new_[10846]_  & ~\new_[10629]_ ;
  assign \new_[9949]_  = ~\new_[10316]_ ;
  assign n8040 = ~\new_[11450]_  & ~\new_[10629]_ ;
  assign \new_[9951]_  = \new_[10630]_  & \new_[14665]_ ;
  assign n8015 = ~\new_[10702]_  | ~\new_[10692]_ ;
  assign n8025 = ~\new_[10704]_  | ~\new_[10691]_ ;
  assign n8020 = ~\new_[10705]_  | ~\new_[10706]_ ;
  assign \new_[9955]_  = \new_[10573]_  | \new_[10893]_ ;
  assign \new_[9956]_  = ~\new_[10690]_  & (~\new_[5757]_  | ~\new_[14164]_ );
  assign \new_[9957]_  = (~\new_[11053]_  & ~\new_[11103]_ ) | (~\new_[11591]_  & ~\new_[10728]_ );
  assign \new_[9958]_  = ~\new_[2097]_  | ~\new_[2094]_  | ~\new_[10623]_  | ~\new_[13209]_ ;
  assign \new_[9959]_  = ~\new_[11857]_  | ~\new_[10708]_  | ~\new_[11329]_ ;
  assign \new_[9960]_  = ~\new_[11851]_  | ~\new_[10713]_  | ~\new_[11084]_ ;
  assign \new_[9961]_  = ~\new_[12117]_  | ~\new_[10711]_  | ~\new_[11076]_ ;
  assign \new_[9962]_  = \new_[3313]_  ^ \new_[10724]_ ;
  assign \new_[9963]_  = \new_[3932]_  ^ \new_[10721]_ ;
  assign \new_[9964]_  = ~\new_[10714]_  & (~\new_[13423]_  | ~\new_[11404]_ );
  assign \new_[9965]_  = \new_[3671]_  ^ \new_[10914]_ ;
  assign \new_[9966]_  = ~\new_[10703]_  & (~\new_[6721]_  | ~\new_[5757]_ );
  assign \new_[9967]_  = \new_[2088]_  ^ \new_[10949]_ ;
  assign \new_[9968]_  = \new_[2087]_  ^ \new_[10950]_ ;
  assign \new_[9969]_  = \new_[11684]_  ^ \new_[10737]_ ;
  assign \new_[9970]_  = \new_[11982]_  ^ \new_[10741]_ ;
  assign \new_[9971]_  = \new_[11456]_  ^ \new_[10735]_ ;
  assign \new_[9972]_  = \new_[12306]_  ^ \new_[10745]_ ;
  assign \new_[9973]_  = \new_[11440]_  ^ \new_[10736]_ ;
  assign \new_[9974]_  = \new_[11719]_  ^ \new_[10738]_ ;
  assign \new_[9975]_  = \new_[11837]_  ^ \new_[10747]_ ;
  assign \new_[9976]_  = \new_[11114]_  & \new_[10618]_ ;
  assign \new_[9977]_  = (~\new_[10767]_  | ~\new_[11727]_ ) & (~\new_[13315]_  | ~\new_[3473]_ );
  assign \new_[9978]_  = \\u0_u0_idle_cnt1_next_reg[5] ;
  assign \new_[9979]_  = ~\new_[10384]_  | ~\new_[10754]_ ;
  assign \new_[9980]_  = ~\new_[10391]_  | ~\new_[10756]_ ;
  assign \new_[9981]_  = ~\new_[10385]_  | ~\new_[10414]_ ;
  assign \new_[9982]_  = ~\new_[10401]_  | ~\new_[10757]_ ;
  assign \new_[9983]_  = ~\new_[10485]_  | ~\new_[11050]_ ;
  assign \new_[9984]_  = ~\new_[10492]_  | ~\new_[11052]_ ;
  assign \new_[9985]_  = ~\new_[10383]_  | ~\new_[6512]_ ;
  assign \new_[9986]_  = ~\new_[10434]_  | ~\new_[11046]_ ;
  assign \new_[9987]_  = ~\new_[10435]_  | ~\new_[11047]_ ;
  assign \new_[9988]_  = ~\new_[10734]_  | ~\new_[10849]_ ;
  assign \new_[9989]_  = ~\new_[10390]_  | ~\new_[10408]_ ;
  assign \new_[9990]_  = ~\new_[10730]_  | ~\new_[10849]_ ;
  assign \new_[9991]_  = ~\new_[11957]_  & ~\new_[10375]_ ;
  assign \new_[9992]_  = ~\new_[10370]_  & (~\new_[13930]_  | ~\new_[14216]_ );
  assign \new_[9993]_  = ~\new_[10729]_  | ~\new_[10849]_ ;
  assign \new_[9994]_  = \new_[11504]_  | \new_[10375]_ ;
  assign \new_[9995]_  = \new_[11800]_  | \new_[10375]_ ;
  assign \new_[9996]_  = ~\new_[10439]_  | ~\new_[11045]_ ;
  assign \new_[9997]_  = ~\new_[10389]_  | ~\new_[10409]_ ;
  assign \new_[9998]_  = ~\new_[10429]_  | ~\new_[11753]_ ;
  assign \new_[9999]_  = ~\new_[10731]_  | ~\new_[10849]_ ;
  assign \new_[10000]_  = ~\new_[10388]_  | ~\new_[12016]_ ;
  assign \new_[10001]_  = ~\new_[10392]_  | ~\new_[12027]_ ;
  assign \new_[10002]_  = ~\new_[10393]_  | ~\new_[12057]_ ;
  assign \new_[10003]_  = u1_u2_sizd_is_zero_reg;
  assign \new_[10004]_  = ~\new_[10381]_  | ~\new_[6304]_ ;
  assign \new_[10005]_  = \new_[11400]_  | \new_[10414]_ ;
  assign \new_[10006]_  = ~\new_[10405]_  | ~\new_[10410]_ ;
  assign \new_[10007]_  = ~\new_[10285]_ ;
  assign \new_[10008]_  = ~\new_[10386]_  | ~\new_[12022]_ ;
  assign \new_[10009]_  = ~\new_[10445]_  | ~\new_[11318]_ ;
  assign \new_[10010]_  = ~\new_[11163]_  & (~\new_[14127]_  | ~\new_[10787]_ );
  assign n8050 = ~\new_[10363]_  & ~\new_[13013]_ ;
  assign \new_[10012]_  = ~\new_[12188]_  | ~\new_[10745]_  | ~\new_[11531]_ ;
  assign \new_[10013]_  = \new_[10727]_  | \new_[12070]_ ;
  assign \new_[10014]_  = (~\new_[12452]_  & ~\new_[3502]_ ) | (~\new_[11066]_  & ~\new_[3777]_ );
  assign \new_[10015]_  = ~\new_[11524]_  | ~\new_[10740]_ ;
  assign \new_[10016]_  = ~\new_[11005]_  & (~\new_[3464]_  | ~\new_[14073]_ );
  assign \new_[10017]_  = ~\new_[11526]_  | ~\new_[10742]_ ;
  assign \new_[10018]_  = ~\new_[10764]_  & (~\new_[3310]_  | ~\new_[14120]_ );
  assign \new_[10019]_  = ~\new_[11183]_  | ~\new_[10746]_ ;
  assign \new_[10020]_  = ~\new_[11181]_  | ~\new_[10748]_ ;
  assign \new_[10021]_  = ~\new_[3691]_  | ~\new_[11754]_  | ~\new_[11086]_ ;
  assign \new_[10022]_  = ~\new_[3480]_  | ~\new_[12299]_  | ~\new_[11078]_ ;
  assign \new_[10023]_  = ~\new_[4291]_  | ~\new_[12281]_  | ~\new_[11073]_ ;
  assign \new_[10024]_  = ~\new_[3884]_  | ~\new_[12303]_  | ~\new_[11072]_ ;
  assign n8185 = \new_[6302]_  ^ \new_[11132]_ ;
  assign n8180 = ~\new_[10403]_ ;
  assign \new_[10027]_  = ~\new_[11212]_  | (~\new_[11182]_  & ~\new_[11152]_ );
  assign \new_[10028]_  = ~\new_[10796]_  & ~\new_[12688]_ ;
  assign \new_[10029]_  = ~\new_[10787]_  | ~\new_[10802]_ ;
  assign \new_[10030]_  = ~\new_[10815]_  | ~\new_[11096]_ ;
  assign \new_[10031]_  = ~\new_[10816]_  | ~\new_[11097]_ ;
  assign \new_[10032]_  = ~XcvSelect_pad_o | ~\new_[10786]_  | ~\new_[13469]_ ;
  assign \new_[10033]_  = ~\new_[11098]_  & ~\new_[10827]_ ;
  assign \new_[10034]_  = ~\new_[14829]_  | ~\new_[4801]_ ;
  assign \new_[10035]_  = \new_[14829]_  & \new_[4852]_ ;
  assign \new_[10036]_  = ~\new_[14829]_  | ~\new_[4800]_ ;
  assign \new_[10037]_  = ~\new_[10812]_  | ~\new_[11555]_ ;
  assign \new_[10038]_  = \new_[10856]_  & \new_[11077]_ ;
  assign \new_[10039]_  = \new_[4161]_  | \new_[10787]_ ;
  assign \new_[10040]_  = ~\new_[4290]_  | ~\new_[10787]_ ;
  assign \new_[10041]_  = ~\new_[10806]_  & ~\new_[12680]_ ;
  assign \new_[10042]_  = ~\new_[10813]_  | ~\new_[13595]_ ;
  assign \new_[10043]_  = \new_[11111]_  & \new_[10792]_ ;
  assign \new_[10044]_  = ~\new_[14829]_  | ~\new_[4802]_ ;
  assign \new_[10045]_  = ~\new_[11012]_  | ~\new_[11571]_ ;
  assign \new_[10046]_  = ~\new_[10810]_  & ~\new_[11419]_ ;
  assign \new_[10047]_  = \new_[10794]_  & \new_[11193]_ ;
  assign \new_[10048]_  = \new_[10807]_  & \new_[11545]_ ;
  assign \new_[10049]_  = \new_[10793]_  & \new_[11539]_ ;
  assign \new_[10050]_  = ~\new_[10818]_  | (~\new_[12152]_  & ~\new_[6725]_ );
  assign \new_[10051]_  = \new_[10788]_  & \new_[11457]_ ;
  assign \new_[10052]_  = \new_[10798]_  & \new_[11191]_ ;
  assign \new_[10053]_  = \new_[10799]_  & \new_[11538]_ ;
  assign \new_[10054]_  = ~\new_[10896]_  | (~\new_[11509]_  & ~\new_[3890]_ );
  assign \new_[10055]_  = \new_[10795]_  & \new_[11190]_ ;
  assign \new_[10056]_  = ~\new_[10402]_ ;
  assign \new_[10057]_  = \new_[10862]_  & \new_[11544]_ ;
  assign \new_[10058]_  = \new_[10809]_  & \new_[11192]_ ;
  assign n8190 = ~\new_[13040]_  & (~\new_[11155]_  | ~\new_[12693]_ );
  assign n8200 = ~\new_[13124]_  & (~\new_[11174]_  | ~\new_[12710]_ );
  assign n8195 = ~\new_[13080]_  & (~\new_[11172]_  | ~\new_[12556]_ );
  assign n8205 = ~\new_[13251]_  & (~\new_[11178]_  | ~\new_[13055]_ );
  assign \new_[10063]_  = ~\new_[10933]_  & ~\new_[11075]_ ;
  assign \new_[10064]_  = ~\new_[10803]_  | (~\new_[11506]_  & ~\new_[4197]_ );
  assign \new_[10065]_  = \new_[2836]_  ^ \new_[11138]_ ;
  assign \new_[10066]_  = ~\new_[10791]_  | (~\new_[11498]_  & ~\new_[3506]_ );
  assign \new_[10067]_  = ~\new_[10856]_  | ~\new_[13165]_ ;
  assign \new_[10068]_  = (~\new_[13714]_  | ~\new_[11797]_ ) & (~\new_[13697]_  | ~\new_[12970]_ );
  assign \new_[10069]_  = ~\new_[10424]_ ;
  assign \new_[10070]_  = ~\new_[10832]_  & ~\new_[12477]_ ;
  assign \new_[10071]_  = \new_[2874]_  ^ \new_[11427]_ ;
  assign \new_[10072]_  = \new_[10967]_  & \new_[12264]_ ;
  assign \new_[10073]_  = \new_[10825]_  & \new_[13882]_ ;
  assign \new_[10074]_  = ~\new_[10888]_  & ~\new_[11490]_ ;
  assign \new_[10075]_  = ~\new_[11147]_  & ~\new_[4792]_ ;
  assign \new_[10076]_  = ~\new_[14737]_  & ~\new_[14386]_ ;
  assign \new_[10077]_  = ~\new_[10868]_  | ~\new_[12926]_ ;
  assign \new_[10078]_  = ~\new_[10866]_  | ~\new_[12977]_ ;
  assign \new_[10079]_  = ~\new_[3790]_  | ~\new_[3710]_  | ~\new_[12552]_  | ~\new_[11306]_ ;
  assign \new_[10080]_  = ~\new_[10837]_  | ~\new_[12694]_ ;
  assign \new_[10081]_  = \new_[10831]_  & \new_[12557]_ ;
  assign \new_[10082]_  = ~\new_[10865]_  | ~\new_[13235]_ ;
  assign \new_[10083]_  = ~\new_[10858]_  & ~\new_[12573]_ ;
  assign \new_[10084]_  = ~\new_[10848]_  | ~\new_[12404]_ ;
  assign \new_[10085]_  = ~\new_[10440]_ ;
  assign \new_[10086]_  = ~\new_[10827]_  | ~\new_[11149]_ ;
  assign \new_[10087]_  = ~\new_[12573]_  & (~\new_[11246]_  | ~\new_[11244]_ );
  assign \new_[10088]_  = ~\new_[10867]_  | ~\new_[13227]_ ;
  assign \new_[10089]_  = ~\new_[10858]_  | ~\new_[12573]_ ;
  assign \new_[10090]_  = ~\new_[11659]_  | (~\new_[11282]_  & ~\new_[4798]_ );
  assign \new_[10091]_  = \new_[10830]_  & \new_[12722]_ ;
  assign \new_[10092]_  = ~\new_[3462]_  | ~\new_[3337]_  | ~\new_[12594]_  | ~\new_[11307]_ ;
  assign \new_[10093]_  = ~\new_[11581]_  | ~\new_[13897]_  | ~\new_[11272]_  | ~\new_[13256]_ ;
  assign \new_[10094]_  = ~\new_[11574]_  | ~\new_[13788]_  | ~\new_[11310]_  | ~\new_[12834]_ ;
  assign \new_[10095]_  = ~\new_[11147]_  | (~\new_[13426]_  & ~\new_[4794]_ );
  assign \new_[10096]_  = ~n8645 | ~\new_[10961]_ ;
  assign \new_[10097]_  = \new_[10460]_ ;
  assign \new_[10098]_  = (~\new_[11278]_  | ~\new_[11314]_ ) & (~\new_[13569]_  | ~\new_[4852]_ );
  assign \new_[10099]_  = (~\new_[13333]_  | ~\new_[12249]_ ) & (~\new_[12941]_  | ~\new_[12135]_ );
  assign n8115 = ~\new_[11685]_  | ~\new_[12341]_  | ~\new_[12045]_  | ~\new_[12344]_ ;
  assign \new_[10101]_  = (~\new_[11316]_  | ~\new_[4615]_ ) & (~\new_[13367]_  | ~\new_[4796]_ );
  assign \new_[10102]_  = ~u4_rx_err_r_reg;
  assign \new_[10103]_  = ~u0_drive_k_r_reg;
  assign \new_[10104]_  = ~\new_[14736]_ ;
  assign \new_[10105]_  = ~\new_[12921]_  | ~\new_[10955]_  | ~\new_[12483]_ ;
  assign \new_[10106]_  = ~\new_[10869]_  & ~\new_[2278]_ ;
  assign \new_[10107]_  = ~\new_[11597]_  & ~\new_[8959]_ ;
  assign \new_[10108]_  = ~\new_[2876]_  | ~\new_[13012]_  | ~\new_[10993]_  | ~\new_[2874]_ ;
  assign n8130 = ~\new_[12756]_  & ~\new_[11573]_ ;
  assign \new_[10110]_  = ~\new_[10488]_ ;
  assign \new_[10111]_  = \new_[11263]_  & \new_[10941]_ ;
  assign \new_[10112]_  = ~\new_[14424]_  | ~\new_[10943]_  | ~\new_[13229]_ ;
  assign \new_[10113]_  = \new_[3472]_  ^ \new_[11412]_ ;
  assign \new_[10114]_  = ~\new_[12690]_  | ~\new_[10940]_  | ~\new_[12430]_ ;
  assign \new_[10115]_  = ~\new_[10967]_  & (~\new_[11696]_  | ~\new_[2345]_ );
  assign \new_[10116]_  = ~\new_[10490]_ ;
  assign \new_[10117]_  = ~n8625 | ~\new_[10869]_ ;
  assign \new_[10118]_  = \new_[2873]_  ^ \new_[11373]_ ;
  assign n8160 = \new_[13664]_  ^ \new_[11408]_ ;
  assign \new_[10120]_  = \new_[13970]_  ^ \new_[11410]_ ;
  assign \new_[10121]_  = \new_[2093]_  ^ \new_[12185]_ ;
  assign \new_[10122]_  = ~\new_[12524]_  | ~\new_[10874]_  | ~\new_[12441]_ ;
  assign \new_[10123]_  = ~\new_[12135]_  | ~\new_[12249]_  | ~\new_[13293]_ ;
  assign \new_[10124]_  = ~\new_[10879]_  | ~\new_[13293]_ ;
  assign \new_[10125]_  = ~n8240 & ~\new_[10893]_ ;
  assign \new_[10126]_  = ~\new_[10946]_  & ~\new_[4792]_ ;
  assign \new_[10127]_  = (~\new_[13538]_  | ~\new_[11489]_ ) & (~\new_[13879]_  | ~\new_[12970]_ );
  assign \new_[10128]_  = ~\new_[12062]_  | (~\new_[11328]_  & ~\new_[4801]_ );
  assign \new_[10129]_  = \new_[10902]_  | \new_[11250]_ ;
  assign \new_[10130]_  = (~\new_[12821]_  | ~\new_[14200]_ ) & (~\new_[12591]_  | ~\new_[4608]_ );
  assign \new_[10131]_  = \new_[3806]_  ^ \new_[11406]_ ;
  assign \new_[10132]_  = (~\new_[13560]_  | ~\new_[11797]_ ) & (~\new_[14159]_  | ~\new_[12970]_ );
  assign \new_[10133]_  = (~\new_[14083]_  | ~\new_[11484]_ ) & (~\new_[13590]_  | ~\new_[12970]_ );
  assign \new_[10134]_  = (~\new_[13500]_  | ~\new_[12811]_ ) & (~\new_[3739]_  | ~\new_[12415]_ );
  assign \new_[10135]_  = (~\new_[13859]_  | ~\new_[11797]_ ) & (~\new_[13983]_  | ~\new_[12970]_ );
  assign \new_[10136]_  = (~\new_[14248]_  | ~\new_[11476]_ ) & (~\new_[13726]_  | ~\new_[12970]_ );
  assign \new_[10137]_  = (~\new_[13954]_  | ~\new_[11797]_ ) & (~\new_[13549]_  | ~\new_[12970]_ );
  assign \new_[10138]_  = (~\new_[13738]_  | ~\new_[11489]_ ) & (~\new_[13812]_  | ~\new_[12970]_ );
  assign \new_[10139]_  = (~\new_[14153]_  | ~\new_[12415]_ ) & (~\new_[6545]_  | ~\new_[12811]_ );
  assign \new_[10140]_  = (~\new_[13537]_  | ~\new_[11476]_ ) & (~\new_[14012]_  | ~\new_[12970]_ );
  assign \new_[10141]_  = (~\new_[14209]_  | ~\new_[11489]_ ) & (~\new_[13669]_  | ~\new_[12970]_ );
  assign \new_[10142]_  = (~\new_[14010]_  | ~\new_[11797]_ ) & (~\new_[13511]_  | ~\new_[12970]_ );
  assign \new_[10143]_  = (~\new_[13527]_  | ~\new_[11476]_ ) & (~\new_[14014]_  | ~\new_[12970]_ );
  assign \new_[10144]_  = (~\new_[13946]_  | ~\new_[12811]_ ) & (~\new_[13638]_  | ~\new_[12415]_ );
  assign \new_[10145]_  = (~\new_[13625]_  | ~\new_[11797]_ ) & (~\new_[14262]_  | ~\new_[12970]_ );
  assign \new_[10146]_  = (~\new_[14117]_  | ~\new_[11484]_ ) & (~\new_[14178]_  | ~\new_[12970]_ );
  assign \new_[10147]_  = (~\new_[14172]_  | ~\new_[12811]_ ) & (~\new_[13525]_  | ~\new_[12415]_ );
  assign \new_[10148]_  = (~\new_[13582]_  | ~\new_[11476]_ ) & (~\new_[13773]_  | ~\new_[12970]_ );
  assign \new_[10149]_  = (~\new_[13557]_  | ~\new_[11484]_ ) & (~\new_[14092]_  | ~\new_[12970]_ );
  assign \new_[10150]_  = (~\new_[13641]_  | ~\new_[11484]_ ) & (~\new_[13652]_  | ~\new_[12970]_ );
  assign \new_[10151]_  = (~\new_[6089]_  | ~\new_[12811]_ ) & (~\new_[14130]_  | ~\new_[12415]_ );
  assign \new_[10152]_  = (~\new_[13632]_  | ~\new_[11797]_ ) & (~\new_[14113]_  | ~\new_[12970]_ );
  assign \new_[10153]_  = (~\new_[13709]_  | ~\new_[11484]_ ) & (~\new_[13622]_  | ~\new_[12970]_ );
  assign \new_[10154]_  = (~\new_[13830]_  | ~\new_[11797]_ ) & (~\new_[13998]_  | ~\new_[12970]_ );
  assign \new_[10155]_  = (~\new_[6549]_  | ~\new_[12811]_ ) & (~\new_[14103]_  | ~\new_[12415]_ );
  assign \new_[10156]_  = (~\new_[6593]_  | ~\new_[12811]_ ) & (~\new_[5490]_  | ~\new_[12415]_ );
  assign \new_[10157]_  = (~\new_[13687]_  | ~\new_[11476]_ ) & (~\new_[13854]_  | ~\new_[12970]_ );
  assign \new_[10158]_  = (~\new_[14009]_  | ~\new_[12811]_ ) & (~\new_[14059]_  | ~\new_[12415]_ );
  assign \new_[10159]_  = (~\new_[14055]_  | ~\new_[11797]_ ) & (~\new_[14233]_  | ~\new_[12970]_ );
  assign \new_[10160]_  = (~\new_[14075]_  | ~\new_[11797]_ ) & (~\new_[13762]_  | ~\new_[12970]_ );
  assign \new_[10161]_  = (~\new_[13822]_  | ~\new_[11797]_ ) & (~\new_[13612]_  | ~\new_[12970]_ );
  assign \new_[10162]_  = (~\new_[13840]_  | ~\new_[11484]_ ) & (~\new_[13948]_  | ~\new_[12970]_ );
  assign \new_[10163]_  = (~\new_[14190]_  | ~\new_[11797]_ ) & (~\new_[13789]_  | ~\new_[12970]_ );
  assign \new_[10164]_  = (~\new_[5998]_  | ~\new_[12811]_ ) & (~\new_[2502]_  | ~\new_[12415]_ );
  assign \new_[10165]_  = (~\new_[13841]_  | ~\new_[11489]_ ) & (~\new_[14030]_  | ~\new_[12970]_ );
  assign \new_[10166]_  = (~\new_[13831]_  | ~\new_[11484]_ ) & (~\new_[14122]_  | ~\new_[12970]_ );
  assign \new_[10167]_  = (~\new_[14134]_  | ~\new_[11489]_ ) & (~\new_[13660]_  | ~\new_[12970]_ );
  assign \new_[10168]_  = (~\new_[13580]_  | ~\new_[11484]_ ) & (~\new_[13784]_  | ~\new_[12970]_ );
  assign \new_[10169]_  = (~\new_[13503]_  | ~\new_[11489]_ ) & (~\new_[14027]_  | ~\new_[12970]_ );
  assign \new_[10170]_  = (~\new_[6268]_  | ~\new_[12811]_ ) & (~\new_[14099]_  | ~\new_[12415]_ );
  assign \new_[10171]_  = (~\new_[13758]_  | ~\new_[11797]_ ) & (~\new_[13996]_  | ~\new_[12970]_ );
  assign \new_[10172]_  = (~\new_[14022]_  | ~\new_[11476]_ ) & (~\new_[13562]_  | ~\new_[12970]_ );
  assign \new_[10173]_  = (~\new_[13885]_  | ~\new_[11797]_ ) & (~\new_[13767]_  | ~\new_[12970]_ );
  assign \new_[10174]_  = (~\new_[5999]_  | ~\new_[12811]_ ) & (~\new_[5112]_  | ~\new_[12415]_ );
  assign \new_[10175]_  = (~\new_[13737]_  | ~\new_[11484]_ ) & (~\new_[14212]_  | ~\new_[12970]_ );
  assign \new_[10176]_  = (~\new_[6274]_  | ~\new_[12811]_ ) & (~\new_[4966]_  | ~\new_[12415]_ );
  assign \new_[10177]_  = (~\new_[13513]_  | ~\new_[11797]_ ) & (~\new_[13834]_  | ~\new_[12970]_ );
  assign \new_[10178]_  = (~\new_[6251]_  | ~\new_[12811]_ ) & (~\new_[4970]_  | ~\new_[12415]_ );
  assign \new_[10179]_  = (~\new_[13713]_  | ~\new_[11476]_ ) & (~\new_[14138]_  | ~\new_[12970]_ );
  assign \new_[10180]_  = (~\new_[6563]_  | ~\new_[12811]_ ) & (~\new_[2553]_  | ~\new_[12415]_ );
  assign \new_[10181]_  = (~\new_[13957]_  | ~\new_[11476]_ ) & (~\new_[13706]_  | ~\new_[12970]_ );
  assign \new_[10182]_  = (~\new_[14007]_  | ~\new_[11797]_ ) & (~\new_[13648]_  | ~\new_[12970]_ );
  assign \new_[10183]_  = (~\new_[6266]_  | ~\new_[12811]_ ) & (~\new_[5499]_  | ~\new_[12415]_ );
  assign \new_[10184]_  = (~\new_[13686]_  | ~\new_[11797]_ ) & (~\new_[13730]_  | ~\new_[12970]_ );
  assign \new_[10185]_  = (~\new_[13958]_  | ~\new_[11484]_ ) & (~\new_[13955]_  | ~\new_[12970]_ );
  assign \new_[10186]_  = (~\new_[13504]_  | ~\new_[11797]_ ) & (~\new_[13587]_  | ~\new_[12970]_ );
  assign \new_[10187]_  = (~\new_[14184]_  | ~\new_[11476]_ ) & (~\new_[13596]_  | ~\new_[12970]_ );
  assign \new_[10188]_  = (~\new_[14144]_  | ~\new_[11797]_ ) & (~\new_[13873]_  | ~\new_[12970]_ );
  assign \new_[10189]_  = (~\new_[11489]_  | ~\new_[13684]_ ) & (~\new_[12970]_  | ~\new_[13724]_ );
  assign \new_[10190]_  = (~\new_[13782]_  | ~\new_[11489]_ ) & (~\new_[13578]_  | ~\new_[12970]_ );
  assign \new_[10191]_  = (~\new_[13965]_  | ~\new_[11476]_ ) & (~\new_[14168]_  | ~\new_[12970]_ );
  assign \new_[10192]_  = (~\new_[13524]_  | ~\new_[11797]_ ) & (~\new_[13871]_  | ~\new_[12970]_ );
  assign \new_[10193]_  = (~\new_[13833]_  | ~\new_[11489]_ ) & (~\new_[13716]_  | ~\new_[12970]_ );
  assign \new_[10194]_  = (~\new_[13619]_  | ~\new_[11484]_ ) & (~\new_[13792]_  | ~\new_[12970]_ );
  assign \new_[10195]_  = (~\new_[13553]_  | ~\new_[11476]_ ) & (~\new_[13976]_  | ~\new_[12970]_ );
  assign \new_[10196]_  = (~\new_[6280]_  | ~\new_[12811]_ ) & (~\new_[13586]_  | ~\new_[12415]_ );
  assign \new_[10197]_  = (~\new_[14166]_  | ~\new_[11476]_ ) & (~\new_[13951]_  | ~\new_[12970]_ );
  assign \new_[10198]_  = (~\new_[14232]_  | ~\new_[12415]_ ) & (~\new_[6172]_  | ~\new_[12811]_ );
  assign \new_[10199]_  = (~\new_[6599]_  | ~\new_[12811]_ ) & (~\new_[5761]_  | ~\new_[12415]_ );
  assign \new_[10200]_  = (~\new_[14072]_  | ~\new_[11489]_ ) & (~\new_[13939]_  | ~\new_[12970]_ );
  assign \new_[10201]_  = (~\new_[14198]_  | ~\new_[11484]_ ) & (~\new_[14132]_  | ~\new_[12970]_ );
  assign \new_[10202]_  = (~\new_[14227]_  | ~\new_[11797]_ ) & (~\new_[13670]_  | ~\new_[12970]_ );
  assign \new_[10203]_  = (~\new_[13972]_  | ~\new_[11476]_ ) & (~\new_[13826]_  | ~\new_[12970]_ );
  assign \new_[10204]_  = (~\new_[13611]_  | ~\new_[12415]_ ) & (~\new_[5149]_  | ~\new_[12811]_ );
  assign \new_[10205]_  = (~\new_[14148]_  | ~\new_[11476]_ ) & (~\new_[14165]_  | ~\new_[12970]_ );
  assign \new_[10206]_  = (~\new_[14201]_  | ~\new_[11489]_ ) & (~\new_[13688]_  | ~\new_[12970]_ );
  assign \new_[10207]_  = (~\new_[13539]_  | ~\new_[11484]_ ) & (~\new_[14220]_  | ~\new_[12970]_ );
  assign \new_[10208]_  = (~\new_[14044]_  | ~\new_[11489]_ ) & (~\new_[13727]_  | ~\new_[12970]_ );
  assign \new_[10209]_  = (~\new_[13499]_  | ~\new_[11797]_ ) & (~\new_[13836]_  | ~\new_[12970]_ );
  assign \new_[10210]_  = (~\new_[14189]_  | ~\new_[11797]_ ) & (~\new_[13717]_  | ~\new_[12970]_ );
  assign \new_[10211]_  = (~\new_[14173]_  | ~\new_[11484]_ ) & (~\new_[13722]_  | ~\new_[12970]_ );
  assign \new_[10212]_  = (~\new_[14097]_  | ~\new_[11484]_ ) & (~\new_[14062]_  | ~\new_[12970]_ );
  assign \new_[10213]_  = (~\new_[13777]_  | ~\new_[11489]_ ) & (~\new_[13860]_  | ~\new_[12970]_ );
  assign \new_[10214]_  = (~\new_[14068]_  | ~\new_[11476]_ ) & (~\new_[14175]_  | ~\new_[12970]_ );
  assign \new_[10215]_  = (~\new_[13610]_  | ~\new_[12811]_ ) & (~\new_[14104]_  | ~\new_[12415]_ );
  assign \new_[10216]_  = (~\new_[14182]_  | ~\new_[11476]_ ) & (~\new_[13935]_  | ~\new_[12970]_ );
  assign \new_[10217]_  = (~\new_[14093]_  | ~\new_[11797]_ ) & (~\new_[13725]_  | ~\new_[12970]_ );
  assign \new_[10218]_  = (~\new_[14196]_  | ~\new_[11797]_ ) & (~\new_[14202]_  | ~\new_[12970]_ );
  assign \new_[10219]_  = (~\new_[6281]_  | ~\new_[12811]_ ) & (~\new_[14265]_  | ~\new_[12415]_ );
  assign \new_[10220]_  = (~\new_[14140]_  | ~\new_[11484]_ ) & (~\new_[13707]_  | ~\new_[12970]_ );
  assign \new_[10221]_  = ~\new_[11677]_  | ~\new_[12080]_  | ~\new_[12565]_  | ~\new_[12591]_ ;
  assign \new_[10222]_  = (~\new_[13994]_  | ~\new_[11489]_ ) & (~\new_[13959]_  | ~\new_[12970]_ );
  assign n8165 = \new_[6301]_  ^ \new_[11388]_ ;
  assign \new_[10224]_  = (~\new_[13839]_  | ~\new_[11484]_ ) & (~\new_[13543]_  | ~\new_[12970]_ );
  assign \new_[10225]_  = \new_[2318]_  ^ \new_[11407]_ ;
  assign \new_[10226]_  = (~\new_[13498]_  | ~\new_[11489]_ ) & (~\new_[13786]_  | ~\new_[12970]_ );
  assign \new_[10227]_  = (~\new_[14090]_  | ~\new_[11489]_ ) & (~\new_[14241]_  | ~\new_[12970]_ );
  assign \new_[10228]_  = \new_[4237]_  ^ \new_[11413]_ ;
  assign \new_[10229]_  = \new_[3429]_  ^ \new_[11411]_ ;
  assign \new_[10230]_  = (~\new_[14222]_  | ~\new_[11484]_ ) & (~\new_[13683]_  | ~\new_[12970]_ );
  assign \new_[10231]_  = \new_[3626]_  ^ \new_[11414]_ ;
  assign n8175 = \new_[6102]_  ^ \new_[11415]_ ;
  assign \new_[10233]_  = (~\new_[13605]_  | ~\new_[11797]_ ) & (~\new_[13791]_  | ~\new_[12970]_ );
  assign \new_[10234]_  = (~\new_[13536]_  | ~\new_[11489]_ ) & (~\new_[13739]_  | ~\new_[12970]_ );
  assign \new_[10235]_  = (~\new_[14207]_  | ~\new_[11489]_ ) & (~\new_[13883]_  | ~\new_[12970]_ );
  assign \new_[10236]_  = (~\new_[13843]_  | ~\new_[11489]_ ) & (~\new_[13607]_  | ~\new_[12970]_ );
  assign \new_[10237]_  = (~\new_[14085]_  | ~\new_[11476]_ ) & (~\new_[14024]_  | ~\new_[12970]_ );
  assign \new_[10238]_  = (~\new_[13887]_  | ~\new_[11484]_ ) & (~\new_[14154]_  | ~\new_[12970]_ );
  assign \new_[10239]_  = (~\new_[13864]_  | ~\new_[11797]_ ) & (~\new_[14021]_  | ~\new_[12970]_ );
  assign \new_[10240]_  = (~\new_[6269]_  | ~\new_[12811]_ ) & (~\new_[13579]_  | ~\new_[12415]_ );
  assign \new_[10241]_  = (~\new_[14206]_  | ~\new_[11484]_ ) & (~\new_[14255]_  | ~\new_[12970]_ );
  assign \new_[10242]_  = (~\new_[13678]_  | ~\new_[11476]_ ) & (~\new_[13838]_  | ~\new_[12970]_ );
  assign \new_[10243]_  = (~\new_[13846]_  | ~\new_[11797]_ ) & (~\new_[13853]_  | ~\new_[12970]_ );
  assign \new_[10244]_  = (~\new_[14056]_  | ~\new_[11797]_ ) & (~\new_[13795]_  | ~\new_[12970]_ );
  assign \new_[10245]_  = (~\new_[13961]_  | ~\new_[11797]_ ) & (~\new_[13982]_  | ~\new_[12970]_ );
  assign \new_[10246]_  = \\u0_u0_idle_cnt1_next_reg[3] ;
  assign \new_[10247]_  = (~\new_[13910]_  | ~\new_[11797]_ ) & (~\new_[13942]_  | ~\new_[12970]_ );
  assign \new_[10248]_  = ~\new_[13002]_  | ~\new_[13341]_  | ~\new_[11407]_ ;
  assign \new_[10249]_  = ~\new_[3592]_  | ~\new_[3502]_  | ~\new_[12595]_  | ~\new_[11308]_ ;
  assign n7980 = ~\new_[10893]_ ;
  assign \new_[10251]_  = ~\new_[6284]_  | ~\new_[12811]_ ;
  assign \new_[10252]_  = ~\new_[2267]_  | ~\new_[12404]_ ;
  assign \new_[10253]_  = ~\new_[12811]_  | ~\new_[6256]_ ;
  assign \new_[10254]_  = ~\new_[13807]_  | ~\new_[12811]_ ;
  assign \new_[10255]_  = ~\new_[6272]_  | ~\new_[12811]_ ;
  assign \new_[10256]_  = ~\new_[4855]_  | ~\new_[12811]_ ;
  assign \new_[10257]_  = ~\new_[5174]_  | ~\new_[12811]_ ;
  assign \new_[10258]_  = ~\new_[13122]_  & ~\new_[4802]_ ;
  assign \new_[10259]_  = ~\new_[6276]_  | ~\new_[12811]_ ;
  assign \new_[10260]_  = ~\new_[5148]_  | ~\new_[12811]_ ;
  assign \new_[10261]_  = ~\new_[10847]_  & ~\new_[12404]_ ;
  assign \new_[10262]_  = \new_[11579]_  & \new_[10984]_ ;
  assign \new_[10263]_  = ~\new_[6267]_  | ~\new_[12811]_ ;
  assign \new_[10264]_  = \new_[11256]_  & \new_[10984]_ ;
  assign \new_[10265]_  = ~\new_[6005]_  | ~\new_[12811]_ ;
  assign \new_[10266]_  = ~\new_[13554]_  | ~\new_[11476]_ ;
  assign \new_[10267]_  = ~\new_[6288]_  | ~\new_[12811]_ ;
  assign \new_[10268]_  = ~\new_[14192]_  | ~\new_[12811]_ ;
  assign \new_[10269]_  = ~\new_[12811]_  | ~\new_[13884]_ ;
  assign \new_[10270]_  = ~\new_[10811]_  | ~\new_[2990]_ ;
  assign \new_[10271]_  = ~\new_[10976]_  & ~\new_[13297]_ ;
  assign \new_[10272]_  = ~\new_[10835]_ ;
  assign \new_[10273]_  = \new_[14205]_  ^ \new_[12760]_ ;
  assign \new_[10274]_  = (~\new_[14221]_  | ~\new_[3638]_ ) & (~\new_[14082]_  | ~\new_[3691]_ );
  assign \new_[10275]_  = (~\new_[4839]_  | ~\new_[12610]_ ) & (~\new_[4840]_  | ~\new_[13756]_ );
  assign \new_[10276]_  = (~\new_[14069]_  | ~\new_[3882]_ ) & (~\new_[13924]_  | ~\new_[3884]_ );
  assign \new_[10277]_  = ~\new_[11716]_  & ~n8240;
  assign \new_[10278]_  = \new_[13568]_  ^ \new_[13646]_ ;
  assign \new_[10279]_  = ~\new_[14452]_  | ~\new_[10942]_  | ~\new_[13122]_ ;
  assign \new_[10280]_  = ~\new_[12298]_  & ~\new_[10966]_ ;
  assign \new_[10281]_  = \new_[3435]_  ^ \new_[11422]_ ;
  assign \new_[10282]_  = ~\new_[10484]_ ;
  assign \new_[10283]_  = ~\new_[4286]_  | ~\new_[4095]_  | ~\new_[12589]_  | ~\new_[11305]_ ;
  assign \new_[10284]_  = \new_[13608]_  ^ \new_[11393]_ ;
  assign \new_[10285]_  = ~\new_[11103]_  | ~\new_[10728]_ ;
  assign \new_[10286]_  = \new_[2875]_  ^ \new_[11417]_ ;
  assign \new_[10287]_  = ~\new_[4854]_  | ~\new_[12811]_ ;
  assign \new_[10288]_  = ~\new_[10973]_  | ~\new_[13819]_ ;
  assign \new_[10289]_  = (~\new_[4816]_  | ~\new_[12610]_ ) & (~\new_[4817]_  | ~\new_[13756]_ );
  assign n9215 = u4_u2_dma_ack_wr1_reg;
  assign \new_[10291]_  = ~\new_[10425]_ ;
  assign \new_[10292]_  = ~\new_[10712]_ ;
  assign n8125 = ~\new_[10662]_ ;
  assign n8120 = ~\new_[10658]_ ;
  assign \new_[10295]_  = \\u4_u1_dma_out_left_reg[2] ;
  assign \new_[10296]_  = \\u4_u0_dma_out_left_reg[2] ;
  assign \new_[10297]_  = \\u4_u3_dma_out_left_reg[2] ;
  assign \new_[10298]_  = \\u4_u2_dma_out_left_reg[2] ;
  assign \new_[10299]_  = ~\new_[12946]_  | ~\new_[10986]_  | ~\new_[13000]_ ;
  assign \new_[10300]_  = ~\new_[10654]_ ;
  assign \new_[10301]_  = ~\new_[12904]_  | ~\new_[10987]_  | ~\new_[12924]_ ;
  assign \new_[10302]_  = ~\new_[10992]_  | ~\new_[13666]_ ;
  assign \new_[10303]_  = ~\new_[13101]_  | ~\new_[10989]_  | ~\new_[13039]_ ;
  assign \new_[10304]_  = ~\new_[12912]_  | ~\new_[10988]_  | ~\new_[13212]_ ;
  assign \new_[10305]_  = ~\new_[11407]_  & (~\new_[12195]_  | ~\new_[2344]_ );
  assign \new_[10306]_  = ~\new_[10984]_  & (~\new_[11457]_  | ~\new_[6232]_ );
  assign \new_[10307]_  = ~\new_[10982]_  | ~\new_[13238]_ ;
  assign \new_[10308]_  = \new_[3505]_  ^ \new_[11368]_ ;
  assign \new_[10309]_  = \new_[11071]_  ^ \new_[4206]_ ;
  assign \new_[10310]_  = \new_[3788]_  ^ \new_[11068]_ ;
  assign \new_[10311]_  = \new_[11070]_  ^ \new_[3889]_ ;
  assign n9150 = u4_u1_dma_ack_wr1_reg;
  assign \new_[10313]_  = \new_[14089]_  ? \new_[10715]_  : \new_[11055]_ ;
  assign \new_[10314]_  = ~\new_[14078]_  | ~\new_[12811]_ ;
  assign \new_[10315]_  = ~\new_[10758]_  & ~\new_[13297]_ ;
  assign \new_[10316]_  = ~\new_[12934]_  | ~\new_[13069]_  | ~\new_[11332]_ ;
  assign \new_[10317]_  = ~\new_[11535]_  & (~\new_[11046]_  | ~\new_[11921]_ );
  assign \new_[10318]_  = ~\new_[11547]_  & (~\new_[11047]_  | ~\new_[12186]_ );
  assign \new_[10319]_  = \new_[13694]_  ^ \new_[11423]_ ;
  assign \new_[10320]_  = ~\new_[11541]_  & (~\new_[11045]_  | ~\new_[11939]_ );
  assign n8170 = ~\new_[11007]_  & ~\new_[12463]_ ;
  assign \new_[10322]_  = ~\new_[11550]_  & (~\new_[11318]_  | ~\new_[11956]_ );
  assign \new_[10323]_  = \new_[3482]_  ^ \new_[11025]_ ;
  assign n8135 = ~\new_[11009]_  | (~\new_[11445]_  & ~\new_[4683]_ );
  assign \new_[10325]_  = \new_[3468]_  ^ \new_[11026]_ ;
  assign \new_[10326]_  = ~\\u4_u2_dma_out_left_reg[1] ;
  assign \new_[10327]_  = ~\new_[10690]_ ;
  assign n8140 = \new_[12115]_  ^ \new_[11021]_ ;
  assign \new_[10329]_  = \new_[11064]_  ^ \new_[11063]_ ;
  assign \new_[10330]_  = \new_[12971]_  ^ \new_[11421]_ ;
  assign \new_[10331]_  = \new_[11059]_  ^ \new_[11058]_ ;
  assign \new_[10332]_  = \new_[13026]_  ^ \new_[11064]_ ;
  assign \new_[10333]_  = \new_[11789]_  ^ \new_[11065]_ ;
  assign \new_[10334]_  = \new_[12931]_  ^ \new_[11421]_ ;
  assign n8145 = \new_[12013]_  ^ \new_[11022]_ ;
  assign n8150 = \new_[11978]_  ^ \new_[11027]_ ;
  assign n8155 = \new_[12181]_  ^ \new_[11029]_ ;
  assign \new_[10338]_  = ~\\u4_u1_dma_out_left_reg[1] ;
  assign \new_[10339]_  = ~\new_[10703]_ ;
  assign \new_[10340]_  = ~\\u4_u0_dma_out_left_reg[1] ;
  assign \new_[10341]_  = ~\\u4_u3_dma_out_left_reg[1] ;
  assign \new_[10342]_  = \new_[11170]_  | \new_[10754]_ ;
  assign n9170 = u4_u0_dma_ack_wr1_reg;
  assign \new_[10344]_  = ~\new_[11095]_  | ~\new_[10819]_  | ~\new_[11796]_ ;
  assign \new_[10345]_  = \new_[11161]_  | \new_[10756]_ ;
  assign n9140 = u4_u3_dma_ack_wr1_reg;
  assign \new_[10347]_  = \new_[11297]_  | \new_[10728]_ ;
  assign \new_[10348]_  = \new_[11176]_  | \new_[10757]_ ;
  assign \new_[10349]_  = ~\new_[11027]_  | ~\new_[10860]_ ;
  assign \new_[10350]_  = ~\new_[12327]_  | ~\new_[10739]_  | ~\new_[11532]_ ;
  assign \new_[10351]_  = ~\new_[11976]_  | ~\new_[10741]_  | ~\new_[11529]_ ;
  assign \new_[10352]_  = ~\new_[12028]_  | ~\new_[10747]_  | ~\new_[11519]_ ;
  assign \new_[10353]_  = \new_[11020]_  | \new_[12147]_ ;
  assign \new_[10354]_  = ~\new_[2083]_  | ~\new_[2095]_  | ~\new_[11042]_  | ~\new_[2094]_ ;
  assign \new_[10355]_  = ~\new_[11184]_  & ~\new_[11738]_ ;
  assign \new_[10356]_  = \new_[14036]_  ^ \new_[11469]_ ;
  assign \new_[10357]_  = \new_[12346]_  ^ \new_[11690]_ ;
  assign \new_[10358]_  = \\u1_u2_rd_buf1_reg[19] ;
  assign \new_[10359]_  = \\u1_u2_rd_buf1_reg[1] ;
  assign \new_[10360]_  = \new_[2346]_  ^ \new_[11466]_ ;
  assign n8225 = ~\new_[10954]_ ;
  assign \new_[10362]_  = \new_[11790]_  ^ \new_[11481]_ ;
  assign \new_[10363]_  = ~\new_[11516]_  | ~\new_[14029]_  | ~\new_[11497]_ ;
  assign \new_[10364]_  = ~\new_[11511]_  | ~\new_[13801]_  | ~\new_[11512]_ ;
  assign \new_[10365]_  = \new_[11106]_  & \new_[2301]_ ;
  assign \new_[10366]_  = \new_[11072]_  & \new_[11815]_ ;
  assign n8235 = ~\new_[10720]_ ;
  assign \new_[10368]_  = ~\new_[11089]_  | ~\new_[3474]_ ;
  assign \new_[10369]_  = \new_[11073]_  & \new_[11806]_ ;
  assign \new_[10370]_  = ~\new_[13369]_  | ~\new_[12267]_  | ~\new_[11507]_ ;
  assign \new_[10371]_  = ~\new_[11698]_  & ~\new_[11430]_ ;
  assign \new_[10372]_  = \new_[11104]_  | \new_[12457]_ ;
  assign \new_[10373]_  = ~\new_[14149]_  | ~\new_[11078]_  | ~\new_[3476]_ ;
  assign n8220 = ~\new_[11088]_  & ~\new_[12444]_ ;
  assign \new_[10375]_  = \new_[11077]_  | \new_[11079]_ ;
  assign \new_[10376]_  = ~\new_[10726]_ ;
  assign \new_[10377]_  = ~\new_[14197]_  | ~\new_[11072]_  | ~\new_[3882]_ ;
  assign \new_[10378]_  = ~\new_[11066]_  | ~\new_[3777]_ ;
  assign \new_[10379]_  = ~\new_[13584]_  | ~\new_[11086]_  | ~\new_[3638]_ ;
  assign \new_[10380]_  = ~\new_[11107]_  | ~\new_[12346]_ ;
  assign \new_[10381]_  = ~\new_[12077]_  | ~\new_[13675]_  | ~\new_[11483]_  | ~\new_[12720]_ ;
  assign \new_[10382]_  = ~\new_[13937]_  | ~\new_[11805]_  | ~\new_[13099]_  | ~\new_[13339]_ ;
  assign \new_[10383]_  = ~\new_[12066]_  | ~\new_[13584]_  | ~\new_[11112]_  | ~\new_[11681]_ ;
  assign \new_[10384]_  = ~\new_[11552]_  & (~\new_[11551]_  | ~\new_[12454]_ );
  assign \new_[10385]_  = ~\new_[11563]_  & (~\new_[11562]_  | ~\new_[12189]_ );
  assign \new_[10386]_  = \new_[11087]_  | \new_[11570]_ ;
  assign \new_[10387]_  = ~\new_[11548]_  & (~\new_[11615]_  | ~\new_[12886]_ );
  assign \new_[10388]_  = \new_[11082]_  | \new_[11546]_ ;
  assign \new_[10389]_  = ~\new_[11540]_  & (~\new_[11549]_  | ~\new_[12111]_ );
  assign \new_[10390]_  = ~\new_[11537]_  & (~\new_[11548]_  | ~\new_[11757]_ );
  assign \new_[10391]_  = ~\new_[11567]_  & (~\new_[11558]_  | ~\new_[12311]_ );
  assign \new_[10392]_  = \new_[11194]_  | \new_[11554]_ ;
  assign \new_[10393]_  = ~\new_[12068]_  & (~\new_[11659]_  | ~\new_[4798]_ );
  assign \new_[10394]_  = ~\new_[11549]_  & (~\new_[11689]_  | ~\new_[12896]_ );
  assign \new_[10395]_  = ~\new_[13532]_  | ~\new_[11242]_  | ~\new_[2373]_ ;
  assign \new_[10396]_  = ~\new_[11874]_  | ~\new_[13962]_  | ~\new_[11245]_  | ~\new_[12712]_ ;
  assign \new_[10397]_  = ~\new_[11543]_  & (~\new_[11600]_  | ~\new_[12884]_ );
  assign \new_[10398]_  = \new_[11362]_  & \new_[11769]_ ;
  assign \new_[10399]_  = ~\new_[11316]_  & (~\new_[11692]_  | ~\new_[4615]_ );
  assign \new_[10400]_  = ~\new_[11701]_  & (~\new_[11543]_  | ~\new_[12162]_ );
  assign \new_[10401]_  = ~\new_[11566]_  & (~\new_[11556]_  | ~\new_[12237]_ );
  assign \new_[10402]_  = \new_[12993]_  & \new_[11242]_ ;
  assign \new_[10403]_  = \new_[11069]_  & \new_[11768]_ ;
  assign \new_[10404]_  = ~\new_[11536]_  & (~\new_[11594]_  | ~\new_[12894]_ );
  assign \new_[10405]_  = ~\new_[11542]_  & (~\new_[11536]_  | ~\new_[12105]_ );
  assign \new_[10406]_  = ~\new_[13463]_  | ~\new_[12162]_  | ~\new_[12884]_  | ~\new_[12455]_ ;
  assign \new_[10407]_  = ~\new_[13668]_  | ~\new_[12811]_ ;
  assign \new_[10408]_  = ~\new_[13325]_  | ~\new_[11757]_  | ~\new_[12886]_  | ~\new_[12370]_ ;
  assign \new_[10409]_  = ~\new_[13381]_  | ~\new_[12111]_  | ~\new_[12896]_  | ~\new_[12482]_ ;
  assign \new_[10410]_  = ~\new_[13285]_  | ~\new_[12105]_  | ~\new_[12894]_  | ~\new_[12352]_ ;
  assign \new_[10411]_  = ~\new_[13024]_  | (~\new_[11561]_  & ~\new_[12533]_ );
  assign n8230 = ~\new_[11080]_  | (~\new_[11875]_  & ~\new_[13710]_ );
  assign \new_[10413]_  = ~\new_[12335]_  | (~\new_[11569]_  & ~\new_[12719]_ );
  assign \new_[10414]_  = ~\new_[13025]_  | ~\new_[12189]_  | ~\new_[13119]_  | ~\new_[13141]_ ;
  assign \new_[10415]_  = ~\new_[11309]_  | (~\new_[11817]_  & ~\new_[3712]_ );
  assign \new_[10416]_  = \new_[13226]_  ^ \new_[11576]_ ;
  assign \new_[10417]_  = ~\\u4_u0_buf0_orig_m3_reg[1] ;
  assign \new_[10418]_  = ~\\u4_u3_buf0_orig_m3_reg[1] ;
  assign \new_[10419]_  = ~\\u4_u2_buf0_orig_m3_reg[1] ;
  assign \new_[10420]_  = ~\new_[11157]_  & (~\new_[11593]_  | ~\new_[11650]_ );
  assign \new_[10421]_  = ~\new_[11166]_  & (~\new_[11936]_  | ~\new_[11654]_ );
  assign \new_[10422]_  = ~\new_[12206]_  | ~\new_[6343]_ ;
  assign \new_[10423]_  = ~\new_[14169]_  | ~\new_[11172]_  | ~\new_[12401]_ ;
  assign \new_[10424]_  = ~\new_[11118]_  | ~\new_[13598]_ ;
  assign \new_[10425]_  = \new_[11140]_  | \wb_addr_i[17] ;
  assign \new_[10426]_  = ~\new_[11188]_  | ~\new_[13118]_ ;
  assign \new_[10427]_  = ~\new_[11189]_  | ~\new_[13118]_ ;
  assign \new_[10428]_  = ~\new_[13804]_  | ~\new_[11155]_  | ~\new_[12466]_ ;
  assign \new_[10429]_  = \new_[11074]_  | \new_[11553]_ ;
  assign \new_[10430]_  = ~\new_[11446]_  | ~\new_[11326]_ ;
  assign \new_[10431]_  = ~\new_[13943]_  | ~\new_[11174]_  | ~\new_[12256]_ ;
  assign \new_[10432]_  = ~\new_[11432]_  & ~\new_[3177]_ ;
  assign \new_[10433]_  = ~\new_[13794]_  | ~\new_[11178]_  | ~\new_[12776]_ ;
  assign \new_[10434]_  = ~\new_[12029]_  & ~\new_[11127]_ ;
  assign \new_[10435]_  = ~\new_[11503]_  & ~\new_[11131]_ ;
  assign \new_[10436]_  = \new_[11799]_  | \new_[11321]_ ;
  assign \new_[10437]_  = \new_[11803]_  | \new_[11134]_ ;
  assign \new_[10438]_  = ~\new_[10948]_ ;
  assign \new_[10439]_  = ~\new_[11141]_  & ~\new_[11144]_ ;
  assign \new_[10440]_  = \new_[11147]_  | \new_[11811]_ ;
  assign \new_[10441]_  = ~\new_[11617]_  | ~\new_[11325]_ ;
  assign \new_[10442]_  = ~\new_[11158]_  | ~\new_[11146]_ ;
  assign \new_[10443]_  = \new_[11122]_  & \new_[11681]_ ;
  assign \new_[10444]_  = ~\new_[11800]_  & ~\new_[13116]_ ;
  assign \new_[10445]_  = ~\new_[11515]_  & ~\new_[11129]_ ;
  assign \new_[10446]_  = \new_[11133]_  & \new_[11806]_ ;
  assign \new_[10447]_  = \new_[11128]_  & \new_[11815]_ ;
  assign \new_[10448]_  = ~\new_[12548]_  & ~\new_[11124]_ ;
  assign \new_[10449]_  = \new_[11237]_  & \new_[11721]_ ;
  assign \new_[10450]_  = \new_[11814]_  | \new_[11151]_ ;
  assign \new_[10451]_  = ~\new_[12500]_  | ~\new_[12617]_  | ~\new_[11487]_  | ~\new_[12700]_ ;
  assign \new_[10452]_  = ~\new_[10811]_ ;
  assign \new_[10453]_  = \new_[11185]_  | \new_[11993]_ ;
  assign \new_[10454]_  = ~\new_[11221]_  & (~\new_[12673]_  | ~\new_[3883]_ );
  assign \new_[10455]_  = \new_[11164]_  & \new_[13182]_ ;
  assign \new_[10456]_  = \new_[11162]_  & \new_[13057]_ ;
  assign \new_[10457]_  = ~\new_[11405]_  & (~\new_[12618]_  | ~\new_[3688]_ );
  assign \new_[10458]_  = ~\new_[11220]_  & (~\new_[12501]_  | ~\new_[4289]_ );
  assign \new_[10459]_  = \new_[11175]_  & \new_[13074]_ ;
  assign \new_[10460]_  = ~\new_[12056]_  & (~\new_[12126]_  | ~\new_[12573]_ );
  assign \new_[10461]_  = ~\new_[11208]_  | (~\new_[14088]_  & ~\new_[4798]_ );
  assign \new_[10462]_  = (~\new_[8959]_  | ~\new_[12349]_ ) & (~\new_[12275]_  | ~\new_[6240]_ );
  assign \new_[10463]_  = ~\new_[10821]_ ;
  assign \new_[10464]_  = (~\new_[11723]_  & ~\new_[13407]_  & ~\new_[13155]_ ) | (~\new_[11444]_  & ~\new_[12146]_  & ~\new_[13398]_ );
  assign \new_[10465]_  = ~u1_u3_pid_OUT_r_reg;
  assign \new_[10466]_  = u4_u2_set_r_reg;
  assign \new_[10467]_  = ~u1_u3_pid_IN_r_reg;
  assign \new_[10468]_  = u4_u0_set_r_reg;
  assign \new_[10469]_  = u4_u1_set_r_reg;
  assign \new_[10470]_  = \new_[11305]_  & \new_[4095]_ ;
  assign \new_[10471]_  = \new_[11307]_  & \new_[3337]_ ;
  assign \new_[10472]_  = \new_[11306]_  & \new_[3710]_ ;
  assign \new_[10473]_  = \new_[11308]_  & \new_[3502]_ ;
  assign \new_[10474]_  = ~\new_[11426]_  & ~\new_[13456]_ ;
  assign \new_[10475]_  = ~\new_[10827]_ ;
  assign \new_[10476]_  = \new_[11229]_  & \new_[13155]_ ;
  assign \new_[10477]_  = ~\new_[14664]_  | ~\new_[2042]_ ;
  assign \new_[10478]_  = ~\new_[11235]_  & ~\new_[13481]_ ;
  assign \new_[10479]_  = ~n8410 | ~\new_[8959]_ ;
  assign \new_[10480]_  = ~n9145 & ~\new_[14806]_ ;
  assign \new_[10481]_  = ~\new_[11240]_  & ~\new_[6091]_ ;
  assign \new_[10482]_  = ~\new_[11418]_  & ~\new_[6323]_ ;
  assign \new_[10483]_  = \new_[11683]_  | \new_[14453]_ ;
  assign \new_[10484]_  = \new_[11268]_  & \new_[11649]_ ;
  assign \new_[10485]_  = ~\new_[13350]_  | ~\new_[11337]_  | ~\new_[12375]_ ;
  assign \new_[10486]_  = ~\new_[11447]_  & ~\new_[11322]_ ;
  assign \new_[10487]_  = ~\new_[12932]_  | ~\new_[11315]_  | ~\new_[13347]_ ;
  assign \new_[10488]_  = ~\new_[14424]_  | ~\new_[11313]_  | ~\new_[13220]_ ;
  assign \new_[10489]_  = ~\new_[11425]_  & ~\new_[13456]_ ;
  assign \new_[10490]_  = ~\new_[14827]_ ;
  assign \new_[10491]_  = ~\new_[11147]_ ;
  assign \new_[10492]_  = ~\new_[12911]_  | ~\new_[11312]_  | ~\new_[12371]_ ;
  assign \new_[10493]_  = \new_[13908]_  ^ \new_[11713]_ ;
  assign \new_[10494]_  = ~\new_[10847]_ ;
  assign \new_[10495]_  = ~\new_[13481]_  | ~\new_[11649]_  | ~\new_[13084]_ ;
  assign \new_[10496]_  = ~\new_[11358]_  & ~\new_[13084]_ ;
  assign \new_[10497]_  = ~\new_[11248]_  | ~\new_[4798]_ ;
  assign \new_[10498]_  = ~\new_[4795]_  | ~\new_[12883]_  | ~\new_[11257]_  | ~\new_[4791]_ ;
  assign \new_[10499]_  = \new_[11394]_  & \new_[13423]_ ;
  assign \new_[10500]_  = ~\new_[11196]_  & ~\new_[11513]_ ;
  assign \new_[10501]_  = ~\new_[4620]_  & (~\new_[12882]_  | ~\new_[11660]_ );
  assign \new_[10502]_  = ~\new_[11276]_  & (~\new_[12165]_  | ~\new_[3711]_ );
  assign \new_[10503]_  = ~\new_[11284]_  | (~\new_[13150]_  & ~\new_[4615]_ );
  assign n8210 = ~\new_[10869]_ ;
  assign \new_[10505]_  = ~\new_[11253]_  & (~\new_[12079]_  | ~\new_[3504]_ );
  assign \new_[10506]_  = ~\new_[11264]_  | (~\new_[13229]_  & ~\new_[12760]_ );
  assign \new_[10507]_  = \\u1_u2_rd_buf1_reg[31] ;
  assign \new_[10508]_  = ~\new_[11271]_  & (~\new_[12088]_  | ~\new_[4293]_ );
  assign \new_[10509]_  = ~\new_[11261]_  & (~\new_[11876]_  | ~\new_[3888]_ );
  assign \new_[10510]_  = (~\new_[13551]_  | ~\new_[11489]_ ) & (~\new_[13592]_  | ~\new_[12970]_ );
  assign \new_[10511]_  = (~\new_[6548]_  | ~\new_[12811]_ ) & (~\new_[13949]_  | ~\new_[12415]_ );
  assign \new_[10512]_  = (~\new_[13986]_  | ~\new_[11489]_ ) & (~\new_[13800]_  | ~\new_[12970]_ );
  assign \new_[10513]_  = (~\new_[6290]_  | ~\new_[12811]_ ) & (~\new_[14042]_  | ~\new_[12415]_ );
  assign \new_[10514]_  = (~\new_[6538]_  | ~\new_[12811]_ ) & (~\new_[14038]_  | ~\new_[12415]_ );
  assign \new_[10515]_  = \\u1_u2_rd_buf1_reg[30] ;
  assign \new_[10516]_  = (~\new_[6260]_  | ~\new_[12811]_ ) & (~\new_[14224]_  | ~\new_[12415]_ );
  assign \new_[10517]_  = (~\new_[6261]_  | ~\new_[12811]_ ) & (~\new_[14057]_  | ~\new_[12415]_ );
  assign \new_[10518]_  = (~\new_[14236]_  | ~\new_[12415]_ ) & (~\new_[6289]_  | ~\new_[12811]_ );
  assign \new_[10519]_  = (~\new_[14155]_  | ~\new_[12811]_ ) & (~\new_[3595]_  | ~\new_[12415]_ );
  assign \new_[10520]_  = (~\new_[6008]_  | ~\new_[12811]_ ) & (~\new_[2500]_  | ~\new_[12415]_ );
  assign \new_[10521]_  = (~\new_[13662]_  | ~\new_[11489]_ ) & (~\new_[13639]_  | ~\new_[12970]_ );
  assign \new_[10522]_  = (~\new_[6690]_  | ~\new_[12811]_ ) & (~\new_[5491]_  | ~\new_[12415]_ );
  assign \new_[10523]_  = (~\new_[6809]_  | ~\new_[12811]_ ) & (~\new_[5562]_  | ~\new_[12415]_ );
  assign \new_[10524]_  = (~\new_[13745]_  | ~\new_[11484]_ ) & (~\new_[14193]_  | ~\new_[12970]_ );
  assign \new_[10525]_  = (~\new_[6004]_  | ~\new_[12811]_ ) & (~\new_[2554]_  | ~\new_[12415]_ );
  assign \new_[10526]_  = (~\new_[6544]_  | ~\new_[12811]_ ) & (~\new_[2551]_  | ~\new_[12415]_ );
  assign \new_[10527]_  = (~\new_[13966]_  | ~\new_[11489]_ ) & (~\new_[13899]_  | ~\new_[12970]_ );
  assign \new_[10528]_  = (~\new_[6200]_  | ~\new_[12811]_ ) & (~\new_[5760]_  | ~\new_[12415]_ );
  assign \new_[10529]_  = (~\new_[6009]_  | ~\new_[12811]_ ) & (~\new_[6032]_  | ~\new_[12415]_ );
  assign \new_[10530]_  = (~\new_[13824]_  | ~\new_[11489]_ ) & (~\new_[13600]_  | ~\new_[12970]_ );
  assign \new_[10531]_  = (~\new_[6485]_  | ~\new_[12811]_ ) & (~\new_[14109]_  | ~\new_[12415]_ );
  assign \new_[10532]_  = (~\new_[14249]_  | ~\new_[11484]_ ) & (~\new_[13991]_  | ~\new_[12970]_ );
  assign \new_[10533]_  = (~\new_[6003]_  | ~\new_[12811]_ ) & (~\new_[2504]_  | ~\new_[12415]_ );
  assign \new_[10534]_  = (~\new_[6293]_  | ~\new_[12811]_ ) & (~\new_[14157]_  | ~\new_[12415]_ );
  assign \new_[10535]_  = (~\new_[14136]_  | ~\new_[11489]_ ) & (~\new_[14253]_  | ~\new_[12970]_ );
  assign \new_[10536]_  = (~\new_[6562]_  | ~\new_[12811]_ ) & (~\new_[6011]_  | ~\new_[12415]_ );
  assign \new_[10537]_  = (~\new_[13618]_  | ~\new_[11489]_ ) & (~\new_[14048]_  | ~\new_[12970]_ );
  assign \new_[10538]_  = (~\new_[14063]_  | ~\new_[12415]_ ) & (~\new_[12811]_  | ~\new_[6258]_ );
  assign \new_[10539]_  = (~\new_[13925]_  | ~\new_[12415]_ ) & (~\new_[4886]_  | ~\new_[12811]_ );
  assign \new_[10540]_  = (~\new_[13681]_  | ~\new_[12415]_ ) & (~\new_[12811]_  | ~\new_[5764]_ );
  assign \new_[10541]_  = (~\new_[6237]_  | ~\new_[12811]_ ) & (~\new_[6013]_  | ~\new_[12415]_ );
  assign \new_[10542]_  = (~\new_[13898]_  | ~\new_[11489]_ ) & (~\new_[13731]_  | ~\new_[12970]_ );
  assign \new_[10543]_  = (~\new_[14177]_  | ~\new_[11484]_ ) & (~\new_[14025]_  | ~\new_[12970]_ );
  assign \new_[10544]_  = (~\new_[13545]_  | ~\new_[11489]_ ) & (~\new_[14137]_  | ~\new_[12970]_ );
  assign \new_[10545]_  = (~\new_[6109]_  | ~\new_[12811]_ ) & (~\new_[13602]_  | ~\new_[12415]_ );
  assign \new_[10546]_  = (~\new_[6279]_  | ~\new_[12811]_ ) & (~\new_[14218]_  | ~\new_[12415]_ );
  assign \new_[10547]_  = \\u1_u2_rd_buf1_reg[7] ;
  assign \new_[10548]_  = (~\new_[14250]_  | ~\new_[11484]_ ) & (~\new_[13931]_  | ~\new_[12970]_ );
  assign \new_[10549]_  = (~\new_[6547]_  | ~\new_[12811]_ ) & (~\new_[13780]_  | ~\new_[12415]_ );
  assign \new_[10550]_  = (~\new_[6001]_  | ~\new_[12811]_ ) & (~\new_[14033]_  | ~\new_[12415]_ );
  assign \new_[10551]_  = (~\new_[14131]_  | ~\new_[12415]_ ) & (~\new_[5185]_  | ~\new_[12811]_ );
  assign \new_[10552]_  = \\u1_u2_rd_buf1_reg[24] ;
  assign \new_[10553]_  = (~\new_[13881]_  | ~\new_[12415]_ ) & (~\new_[6543]_  | ~\new_[12811]_ );
  assign \new_[10554]_  = (~\new_[6524]_  | ~\new_[12811]_ ) & (~\new_[13509]_  | ~\new_[12415]_ );
  assign \new_[10555]_  = (~\new_[6000]_  | ~\new_[12811]_ ) & (~\new_[14180]_  | ~\new_[12415]_ );
  assign \new_[10556]_  = (~\new_[13867]_  | ~\new_[11489]_ ) & (~\new_[13774]_  | ~\new_[12970]_ );
  assign \new_[10557]_  = (~\new_[6002]_  | ~\new_[12811]_ ) & (~\new_[14039]_  | ~\new_[12415]_ );
  assign \new_[10558]_  = (~\new_[13820]_  | ~\new_[11489]_ ) & (~\new_[14023]_  | ~\new_[12970]_ );
  assign \new_[10559]_  = (~\new_[13729]_  | ~\new_[11484]_ ) & (~\new_[13888]_  | ~\new_[12970]_ );
  assign \new_[10560]_  = (~\new_[13743]_  | ~\new_[11489]_ ) & (~\new_[13911]_  | ~\new_[12970]_ );
  assign \new_[10561]_  = (~\new_[13764]_  | ~\new_[12811]_ ) & (~\new_[3741]_  | ~\new_[12415]_ );
  assign \new_[10562]_  = ~\new_[11277]_  & (~\new_[2816]_  | ~\new_[14314]_ );
  assign \new_[10563]_  = ~\new_[11285]_  & (~\new_[2828]_  | ~\new_[14314]_ );
  assign \new_[10564]_  = ~\new_[11040]_  & (~\new_[2815]_  | ~\new_[14314]_ );
  assign \new_[10565]_  = ~\new_[11283]_  & (~\new_[2813]_  | ~\new_[14314]_ );
  assign \new_[10566]_  = \new_[14185]_  ^ \new_[11722]_ ;
  assign \new_[10567]_  = ~\new_[11336]_  & (~\new_[2811]_  | ~\new_[14314]_ );
  assign \new_[10568]_  = \\u1_u2_rd_buf1_reg[21] ;
  assign \new_[10569]_  = \new_[11406]_  & \new_[12569]_ ;
  assign \new_[10570]_  = \new_[12004]_  ^ \new_[11740]_ ;
  assign \new_[10571]_  = \new_[11918]_  & \new_[11388]_ ;
  assign \new_[10572]_  = ~\new_[14273]_ ;
  assign \new_[10573]_  = ~\new_[10939]_ ;
  assign \new_[10574]_  = \new_[11331]_  & \new_[14167]_ ;
  assign \new_[10575]_  = \new_[11413]_  & \new_[12757]_ ;
  assign \new_[10576]_  = ~\new_[11626]_  | ~\new_[9191]_  | ~\new_[11697]_ ;
  assign \new_[10577]_  = ~\new_[5503]_  | ~\new_[12811]_ ;
  assign \new_[10578]_  = ~\new_[6275]_  | ~\new_[12811]_ ;
  assign \new_[10579]_  = ~\new_[6196]_  | ~\new_[12811]_ ;
  assign \new_[10580]_  = ~\new_[5502]_  | ~\new_[12811]_ ;
  assign \new_[10581]_  = ~\new_[5604]_  | ~\new_[12811]_ ;
  assign \new_[10582]_  = \new_[12485]_  & \new_[11412]_ ;
  assign \new_[10583]_  = \new_[11413]_  & \new_[12421]_ ;
  assign \new_[10584]_  = ~\new_[14181]_  | ~\new_[12811]_ ;
  assign \new_[10585]_  = ~\new_[12811]_  | ~\new_[5763]_ ;
  assign \new_[10586]_  = ~\new_[13922]_  | ~\new_[12811]_ ;
  assign \new_[10587]_  = ~\new_[13533]_  | ~\new_[12811]_ ;
  assign \new_[10588]_  = ~\new_[13597]_  | ~\new_[12811]_ ;
  assign \new_[10589]_  = ~\new_[6552]_  | ~\new_[12811]_ ;
  assign \new_[10590]_  = ~\new_[6287]_  | ~\new_[12811]_ ;
  assign \new_[10591]_  = ~\new_[6166]_  | ~\new_[12811]_ ;
  assign \new_[10592]_  = ~\new_[13615]_  | ~\new_[12811]_ ;
  assign \new_[10593]_  = ~\new_[6277]_  | ~\new_[12811]_ ;
  assign \new_[10594]_  = ~\new_[12811]_  | ~\new_[5762]_ ;
  assign \new_[10595]_  = ~\new_[13894]_  | ~\new_[12811]_ ;
  assign \new_[10596]_  = ~\new_[10838]_ ;
  assign \new_[10597]_  = ~\new_[14098]_  | ~\new_[12811]_ ;
  assign \new_[10598]_  = ~\new_[6247]_  | ~\new_[12811]_ ;
  assign \new_[10599]_  = ~\new_[2193]_  & ~\new_[12160]_ ;
  assign \new_[10600]_  = ~\new_[6264]_  | ~\new_[12811]_ ;
  assign \new_[10601]_  = ~\new_[6254]_  | ~\new_[12811]_ ;
  assign \new_[10602]_  = ~\new_[13220]_  & ~\new_[12760]_ ;
  assign \new_[10603]_  = ~\new_[6567]_  | ~\new_[12811]_ ;
  assign \new_[10604]_  = ~\new_[13741]_  | ~\new_[12811]_ ;
  assign \new_[10605]_  = \new_[11411]_  & \new_[12419]_ ;
  assign \new_[10606]_  = \new_[11411]_  & \new_[12511]_ ;
  assign \new_[10607]_  = \new_[8702]_  ^ \new_[8959]_ ;
  assign \new_[10608]_  = \new_[2874]_  ^ \new_[4800]_ ;
  assign \new_[10609]_  = ~\new_[11235]_  & ~\new_[12414]_ ;
  assign \new_[10610]_  = \new_[9442]_  ^ \new_[8959]_ ;
  assign \new_[10611]_  = (~\new_[4835]_  | ~\new_[13861]_ ) & (~\new_[4837]_  | ~\new_[14790]_ );
  assign \new_[10612]_  = \new_[11808]_  | \new_[11231]_ ;
  assign \new_[10613]_  = (~\new_[13552]_  | ~\new_[3476]_ ) & (~\new_[14199]_  | ~\new_[3480]_ );
  assign \new_[10614]_  = \new_[11414]_  & \new_[12247]_ ;
  assign \new_[10615]_  = \new_[11414]_  & \new_[12518]_ ;
  assign n8215 = u0_u0_usb_reset_reg;
  assign \new_[10617]_  = \new_[11245]_  & \new_[11388]_ ;
  assign \new_[10618]_  = \new_[11914]_  & \new_[11415]_ ;
  assign \new_[10619]_  = \new_[11310]_  & \new_[11415]_ ;
  assign \new_[10620]_  = ~\new_[11000]_ ;
  assign \new_[10621]_  = \new_[11406]_  & \new_[12297]_ ;
  assign \new_[10622]_  = \new_[13870]_  ^ \new_[11718]_ ;
  assign \new_[10623]_  = ~\new_[10949]_ ;
  assign \new_[10624]_  = \new_[14041]_  ^ \new_[11704]_ ;
  assign \new_[10625]_  = ~\new_[13675]_  | ~\new_[11073]_  | ~\new_[4288]_ ;
  assign \new_[10626]_  = ~u1_u2_dtmp_sel_r_reg;
  assign \new_[10627]_  = ~\new_[11392]_  | ~\new_[14261]_ ;
  assign \new_[10628]_  = ~u1_u3_pid_SETUP_r_reg;
  assign \new_[10629]_  = u1_u3_rx_ack_to_clr_reg;
  assign \new_[10630]_  = ~u1_u3_pid_PING_r_reg;
  assign \new_[10631]_  = u4_u2_r2_reg;
  assign \new_[10632]_  = \\u1_u2_rd_buf1_reg[26] ;
  assign \new_[10633]_  = \\u1_u2_rd_buf1_reg[27] ;
  assign \new_[10634]_  = \\u1_u2_rd_buf1_reg[3] ;
  assign \new_[10635]_  = \\u1_u2_rd_buf1_reg[0] ;
  assign \new_[10636]_  = \\u1_u2_rd_buf1_reg[12] ;
  assign \new_[10637]_  = \\u1_u2_rd_buf1_reg[2] ;
  assign \new_[10638]_  = \\u1_u2_rd_buf1_reg[8] ;
  assign \new_[10639]_  = \\u1_u2_rd_buf1_reg[18] ;
  assign \new_[10640]_  = \\u1_u2_rd_buf1_reg[28] ;
  assign \new_[10641]_  = \\u1_u2_rd_buf1_reg[14] ;
  assign \new_[10642]_  = u4_u3_set_r_reg;
  assign \new_[10643]_  = \\u1_u2_rd_buf1_reg[6] ;
  assign \new_[10644]_  = \\u1_u2_rd_buf1_reg[5] ;
  assign \new_[10645]_  = \\u1_u2_rd_buf1_reg[9] ;
  assign \new_[10646]_  = \\u1_u2_rd_buf1_reg[20] ;
  assign \new_[10647]_  = \\u1_u2_rd_buf1_reg[22] ;
  assign \new_[10648]_  = \\u1_u2_rd_buf1_reg[15] ;
  assign \new_[10649]_  = \\u1_u2_rd_buf1_reg[23] ;
  assign \new_[10650]_  = ~\new_[3473]_  | ~\new_[3435]_  | ~\new_[11412]_  | ~\new_[3472]_ ;
  assign \new_[10651]_  = \\u1_u2_rd_buf1_reg[25] ;
  assign \new_[10652]_  = \\u1_u2_rd_buf1_reg[17] ;
  assign \new_[10653]_  = u4_u3_r2_reg;
  assign \new_[10654]_  = ~\new_[13002]_  | ~\new_[12978]_  | ~\new_[12429]_ ;
  assign \new_[10655]_  = ~\new_[11286]_  & (~\new_[2817]_  | ~\new_[14314]_ );
  assign \new_[10656]_  = \\u1_u2_rd_buf1_reg[16] ;
  assign \new_[10657]_  = \new_[12825]_  & \new_[11422]_ ;
  assign \new_[10658]_  = ~\new_[11388]_  & (~\new_[11762]_  | ~\new_[6300]_ );
  assign \new_[10659]_  = ~\new_[11413]_  & (~\new_[12141]_  | ~\new_[3997]_ );
  assign \new_[10660]_  = ~\new_[11411]_  & (~\new_[12136]_  | ~\new_[3342]_ );
  assign \new_[10661]_  = ~\new_[11414]_  & (~\new_[11769]_  | ~\new_[3510]_ );
  assign \new_[10662]_  = ~\new_[11415]_  & (~\new_[11768]_  | ~\new_[6368]_ );
  assign \new_[10663]_  = ~\new_[11406]_  & (~\new_[11765]_  | ~\new_[3715]_ );
  assign \new_[10664]_  = \\u1_u2_rd_buf1_reg[4] ;
  assign \new_[10665]_  = \new_[2872]_  ^ \new_[12227]_ ;
  assign \new_[10666]_  = \new_[3025]_  ^ \new_[11458]_ ;
  assign \new_[10667]_  = u4_u0_r2_reg;
  assign \new_[10668]_  = u4_u1_r2_reg;
  assign \new_[10669]_  = \\u1_u2_rd_buf1_reg[29] ;
  assign \new_[10670]_  = ~\new_[11273]_  & (~\new_[2814]_  | ~\new_[14314]_ );
  assign \new_[10671]_  = ~\new_[11269]_  & (~\new_[2812]_  | ~\new_[14314]_ );
  assign \new_[10672]_  = (~\new_[11700]_  | ~\new_[11727]_ ) & (~\new_[13315]_  | ~\new_[3410]_ );
  assign \new_[10673]_  = \new_[11179]_  | \new_[12215]_ ;
  assign \new_[10674]_  = \\u1_u2_rd_buf1_reg[10] ;
  assign \new_[10675]_  = \new_[11071]_  & \new_[4206]_ ;
  assign \new_[10676]_  = \new_[11368]_  & \new_[3505]_ ;
  assign \new_[10677]_  = ~\new_[11067]_  & ~\new_[6344]_ ;
  assign \new_[10678]_  = \new_[11068]_  & \new_[3788]_ ;
  assign \new_[10679]_  = \new_[11070]_  & \new_[3889]_ ;
  assign \new_[10680]_  = ~\new_[13443]_  | ~\new_[11429]_ ;
  assign \new_[10681]_  = ~\new_[13858]_  | ~\new_[12082]_  | ~\new_[13407]_ ;
  assign \new_[10682]_  = ~\new_[13268]_  | ~\new_[11071]_  | ~\new_[4206]_ ;
  assign \new_[10683]_  = ~\new_[13466]_  | ~\new_[11368]_  | ~\new_[3505]_ ;
  assign \new_[10684]_  = ~\new_[12987]_  | ~\new_[11068]_  | ~\new_[3788]_ ;
  assign \new_[10685]_  = ~\new_[13351]_  | ~\new_[11070]_  | ~\new_[3889]_ ;
  assign \new_[10686]_  = \new_[11260]_  & \new_[11014]_ ;
  assign \new_[10687]_  = \new_[4074]_  ^ \new_[11435]_ ;
  assign \new_[10688]_  = \new_[3317]_  ^ \new_[11436]_ ;
  assign \new_[10689]_  = \new_[3692]_  ^ \new_[11438]_ ;
  assign \new_[10690]_  = u4_u1_intb_reg;
  assign \new_[10691]_  = ~u4_u2_intb_reg;
  assign \new_[10692]_  = ~u4_u0_intb_reg;
  assign \new_[10693]_  = \new_[2097]_  ^ \new_[11433]_ ;
  assign \new_[10694]_  = \\u1_u2_rd_buf1_reg[11] ;
  assign \new_[10695]_  = \\u1_u2_rd_buf1_reg[13] ;
  assign \new_[10696]_  = (~\new_[13367]_  | ~\new_[14790]_ ) & (~\new_[2871]_  | ~\new_[4796]_ );
  assign \new_[10697]_  = \new_[11979]_  ^ \new_[11735]_ ;
  assign \new_[10698]_  = \new_[11985]_  ^ \new_[11741]_ ;
  assign \new_[10699]_  = \new_[12023]_  ^ \new_[11738]_ ;
  assign \new_[10700]_  = ~\new_[6255]_  | ~\new_[12811]_ ;
  assign \new_[10701]_  = \new_[11167]_  & \new_[13006]_ ;
  assign \new_[10702]_  = ~u4_u0_inta_reg;
  assign \new_[10703]_  = u4_u1_inta_reg;
  assign \new_[10704]_  = ~u4_u2_inta_reg;
  assign \new_[10705]_  = ~u4_u3_inta_reg;
  assign \new_[10706]_  = ~u4_u3_intb_reg;
  assign \new_[10707]_  = ~\new_[13012]_  | ~\new_[2932]_  | ~\new_[11139]_  | ~\new_[2836]_ ;
  assign \new_[10708]_  = ~\new_[11021]_  | ~\new_[11160]_ ;
  assign \new_[10709]_  = ~\new_[12104]_  & ~\new_[11025]_ ;
  assign \new_[10710]_  = ~\new_[7206]_  | ~\new_[13771]_  | ~\new_[11234]_  | ~\new_[11779]_ ;
  assign \new_[10711]_  = ~\new_[11029]_  | ~\new_[11187]_ ;
  assign \new_[10712]_  = ~\new_[11043]_  | ~\new_[12053]_ ;
  assign \new_[10713]_  = ~\new_[11022]_  | ~\new_[11169]_ ;
  assign \new_[10714]_  = ~\new_[11011]_ ;
  assign \new_[10715]_  = u0_u0_me_ps_2_5_us_reg;
  assign \new_[10716]_  = ~\new_[11186]_  & ~\new_[11735]_ ;
  assign \new_[10717]_  = ~\new_[11533]_  & ~\new_[11741]_ ;
  assign \new_[10718]_  = \new_[3013]_  ^ \new_[11786]_ ;
  assign \new_[10719]_  = \new_[12129]_  ^ \new_[11787]_ ;
  assign \new_[10720]_  = \new_[11491]_  | \new_[11466]_ ;
  assign \new_[10721]_  = \new_[13472]_  | \new_[4074]_  | \new_[11506]_  | \new_[4236]_ ;
  assign \new_[10722]_  = ~\new_[13647]_  | ~\new_[12415]_ ;
  assign \new_[10723]_  = ~\new_[11466]_  & ~\new_[12806]_ ;
  assign \new_[10724]_  = \new_[13468]_  | \new_[3317]_  | \new_[11498]_  | \new_[3428]_ ;
  assign \new_[10725]_  = ~\new_[11024]_ ;
  assign \new_[10726]_  = ~\new_[2478]_  | ~\new_[11916]_  | ~\new_[12059]_ ;
  assign \new_[10727]_  = \new_[11465]_  | \new_[12956]_ ;
  assign \new_[10728]_  = ~\new_[6233]_  | ~\new_[14118]_  | ~\new_[11507]_  | ~\new_[13933]_ ;
  assign \new_[10729]_  = ~\new_[11478]_  | (~\new_[12152]_  & ~\new_[6730]_ );
  assign \new_[10730]_  = ~\new_[11473]_  | (~\new_[12152]_  & ~\new_[6754]_ );
  assign \new_[10731]_  = ~\new_[11475]_  | (~\new_[12152]_  & ~\new_[6729]_ );
  assign \new_[10732]_  = ~\new_[11472]_  | (~\new_[12152]_  & ~\new_[6732]_ );
  assign \new_[10733]_  = ~\new_[2858]_  | ~\new_[11437]_ ;
  assign \new_[10734]_  = ~\new_[11477]_  | (~\new_[12152]_  & ~\new_[6731]_ );
  assign \new_[10735]_  = ~\new_[11045]_ ;
  assign \new_[10736]_  = ~\new_[11046]_ ;
  assign \new_[10737]_  = ~\new_[11047]_ ;
  assign \new_[10738]_  = ~\new_[11318]_ ;
  assign \new_[10739]_  = ~\new_[11470]_  | ~\new_[11839]_ ;
  assign \new_[10740]_  = ~\new_[12315]_  | (~\new_[11839]_  & ~\new_[12468]_ );
  assign \new_[10741]_  = ~\new_[11467]_  | ~\new_[11845]_ ;
  assign \new_[10742]_  = ~\new_[11995]_  | (~\new_[11845]_  & ~\new_[12248]_ );
  assign \new_[10743]_  = ~\new_[12945]_  | (~\new_[12050]_  & ~\new_[12749]_ );
  assign \new_[10744]_  = ~\new_[13168]_  | (~\new_[11856]_  & ~\new_[12682]_ );
  assign \new_[10745]_  = ~\new_[11714]_  | ~\new_[11860]_ ;
  assign \new_[10746]_  = ~\new_[12215]_  | (~\new_[11860]_  & ~\new_[12400]_ );
  assign \new_[10747]_  = ~\new_[11468]_  | ~\new_[11868]_ ;
  assign \new_[10748]_  = ~\new_[11993]_  | (~\new_[11868]_  & ~\new_[12224]_ );
  assign \new_[10749]_  = ~\new_[4286]_  | ~\new_[12434]_  | ~\new_[11806]_ ;
  assign \new_[10750]_  = ~\new_[3790]_  | ~\new_[12300]_  | ~\new_[11815]_ ;
  assign \new_[10751]_  = (~\new_[12963]_  | ~\new_[3671]_ ) & (~\new_[11831]_  | ~\new_[12747]_ );
  assign \new_[10752]_  = (~\new_[13112]_  | ~\new_[3313]_ ) & (~\new_[11827]_  | ~\new_[12593]_ );
  assign \new_[10753]_  = (~\new_[13158]_  | ~\new_[3468]_ ) & (~\new_[11829]_  | ~\new_[12868]_ );
  assign \new_[10754]_  = ~\new_[13087]_  | ~\new_[12454]_  | ~\new_[12995]_  | ~\new_[12984]_ ;
  assign \new_[10755]_  = ~\new_[13987]_  | ~\new_[2452]_  | ~\new_[12059]_  | ~\new_[13228]_ ;
  assign \new_[10756]_  = ~\new_[13004]_  | ~\new_[12311]_  | ~\new_[13142]_  | ~\new_[12968]_ ;
  assign \new_[10757]_  = ~\new_[12992]_  | ~\new_[12237]_  | ~\new_[12959]_  | ~\new_[13105]_ ;
  assign \new_[10758]_  = \new_[3037]_  ^ \new_[12103]_ ;
  assign \new_[10759]_  = ~\new_[7670]_  | ~\new_[12404]_ ;
  assign \new_[10760]_  = ~\new_[6163]_  | ~\new_[12811]_ ;
  assign \new_[10761]_  = \new_[12210]_  ^ \new_[3504]_ ;
  assign \new_[10762]_  = \new_[12204]_  ^ \new_[3888]_ ;
  assign \new_[10763]_  = \new_[12208]_  ^ \new_[3711]_ ;
  assign \new_[10764]_  = ~\new_[11501]_  & (~\new_[11853]_  | ~\new_[13174]_ );
  assign n8285 = \new_[12995]_  ^ \new_[11989]_ ;
  assign \new_[10766]_  = \new_[13006]_  ^ \new_[11776]_ ;
  assign \new_[10767]_  = \new_[3473]_  ^ \new_[11793]_ ;
  assign \new_[10768]_  = \new_[13182]_  ^ \new_[12003]_ ;
  assign \new_[10769]_  = \new_[13074]_  ^ \new_[11977]_ ;
  assign n8300 = \new_[13142]_  ^ \new_[11755]_ ;
  assign \new_[10771]_  = ~\new_[2830]_  | ~\new_[11437]_ ;
  assign \new_[10772]_  = \new_[13061]_  ^ \new_[12110]_ ;
  assign \new_[10773]_  = \new_[12971]_  ^ \new_[11910]_ ;
  assign \new_[10774]_  = \new_[4500]_  ^ \new_[11909]_ ;
  assign n8295 = \new_[12959]_  ^ \new_[11777]_ ;
  assign n8290 = \new_[13119]_  ^ \new_[11968]_ ;
  assign \new_[10777]_  = \new_[13057]_  ^ \new_[11961]_ ;
  assign \new_[10778]_  = ~\\u4_u3_dma_out_left_reg[0] ;
  assign \new_[10779]_  = ~\\u4_u2_dma_out_left_reg[0] ;
  assign \new_[10780]_  = ~\\u4_u0_dma_out_left_reg[0] ;
  assign n8310 = ~\new_[11520]_  & ~\new_[13296]_ ;
  assign n8305 = ~\new_[11527]_  & ~\new_[13296]_ ;
  assign n8280 = ~\new_[11521]_  & ~\new_[13296]_ ;
  assign n8255 = ~\new_[11534]_  & ~\new_[13296]_ ;
  assign \new_[10785]_  = \new_[11437]_  | \new_[13156]_ ;
  assign \new_[10786]_  = ~\new_[11499]_  | ~\new_[13469]_ ;
  assign \new_[10787]_  = ~\new_[11495]_  | ~\wb_addr_i[17] ;
  assign \new_[10788]_  = \new_[12557]_  | \new_[13761]_ ;
  assign \new_[10789]_  = ~\new_[6252]_  | ~\new_[12811]_ ;
  assign \new_[10790]_  = \new_[12557]_  & \new_[11578]_ ;
  assign \new_[10791]_  = ~\new_[11498]_  | ~\new_[3506]_ ;
  assign \new_[10792]_  = \new_[11486]_  & \new_[12720]_ ;
  assign \new_[10793]_  = ~\new_[11542]_  | ~\new_[12872]_ ;
  assign \new_[10794]_  = ~\new_[11547]_  | ~\new_[11780]_ ;
  assign \new_[10795]_  = ~\new_[11535]_  | ~\new_[12177]_ ;
  assign \new_[10796]_  = ~\new_[13138]_  | ~\new_[11507]_  | ~\new_[12696]_ ;
  assign \new_[10797]_  = \new_[11752]_  & \new_[11434]_ ;
  assign \new_[10798]_  = ~\new_[11541]_  | ~\new_[11937]_ ;
  assign \new_[10799]_  = ~\new_[11540]_  | ~\new_[12521]_ ;
  assign \new_[10800]_  = \new_[11681]_  & \new_[11583]_ ;
  assign \new_[10801]_  = ~\new_[11448]_  | ~\new_[11505]_ ;
  assign \new_[10802]_  = ~\new_[11496]_  | ~\wb_addr_i[17] ;
  assign \new_[10803]_  = ~\new_[11506]_  | ~\new_[4197]_ ;
  assign \new_[10804]_  = ~\new_[11647]_  & ~\new_[12448]_ ;
  assign \new_[10805]_  = ~\new_[11801]_  | ~\new_[13469]_ ;
  assign \new_[10806]_  = ~\new_[11106]_ ;
  assign \new_[10807]_  = ~\new_[11537]_  | ~\new_[12600]_ ;
  assign \new_[10808]_  = \new_[12722]_  & \new_[11557]_ ;
  assign \new_[10809]_  = ~\new_[11550]_  | ~\new_[11965]_ ;
  assign \new_[10810]_  = \new_[12325]_  | \new_[12476]_  | \new_[11644]_  | \new_[12480]_ ;
  assign \new_[10811]_  = ~\new_[12782]_  & ~\new_[11686]_ ;
  assign \new_[10812]_  = \new_[11530]_  | \new_[11995]_ ;
  assign \new_[10813]_  = \new_[11798]_  & \new_[11505]_ ;
  assign \new_[10814]_  = ~\new_[11669]_  & ~\new_[13481]_ ;
  assign \new_[10815]_  = (~\new_[12549]_  | ~\new_[11942]_ ) & (~\new_[12275]_  | ~\new_[6105]_ );
  assign \new_[10816]_  = (~\new_[12275]_  | ~\new_[6243]_ ) & (~\new_[12691]_  | ~\new_[11942]_ );
  assign \new_[10817]_  = \new_[12048]_  ? \new_[12047]_  : \new_[12346]_ ;
  assign \new_[10818]_  = (~\new_[3463]_  | ~\new_[12671]_ ) & (~\new_[12599]_  | ~\new_[11942]_ );
  assign \new_[10819]_  = (~\new_[12602]_  | ~\new_[11942]_ ) & (~\new_[12349]_  | ~\new_[13465]_ );
  assign \new_[10820]_  = ~\new_[11668]_  & ~\new_[6003]_ ;
  assign \new_[10821]_  = (~n8340 | ~\new_[13415]_ ) & (~\new_[12126]_  | ~\new_[8810]_ );
  assign \new_[10822]_  = ~\new_[2896]_  | ~\new_[11663]_ ;
  assign \new_[10823]_  = ~\new_[11104]_ ;
  assign \new_[10824]_  = \new_[12180]_  ^ \new_[12648]_ ;
  assign \new_[10825]_  = ~\new_[11582]_  & ~\new_[13407]_ ;
  assign \new_[10826]_  = ~\new_[3461]_  & ~\new_[12278]_ ;
  assign \new_[10827]_  = ~\new_[11613]_  | ~\wb_addr_i[4] ;
  assign \new_[10828]_  = ~\new_[11606]_  | ~\new_[11649]_ ;
  assign \new_[10829]_  = ~\new_[11123]_ ;
  assign \new_[10830]_  = \new_[11557]_  & \new_[14197]_ ;
  assign \new_[10831]_  = \new_[11578]_  & \new_[14149]_ ;
  assign \new_[10832]_  = \new_[11645]_  | \new_[12253]_ ;
  assign \new_[10833]_  = ~\new_[13469]_  | ~\new_[12101]_ ;
  assign \new_[10834]_  = ~\new_[13461]_  | ~\new_[11653]_  | ~\new_[12785]_ ;
  assign \new_[10835]_  = ~\new_[11596]_  & ~\wb_addr_i[4] ;
  assign \new_[10836]_  = ~\new_[13355]_  | ~\new_[11682]_  | ~\new_[12713]_ ;
  assign \new_[10837]_  = \new_[14739]_  & \new_[11585]_ ;
  assign \new_[10838]_  = ~\new_[11702]_  | ~\new_[11697]_ ;
  assign \new_[10839]_  = ~\new_[11130]_ ;
  assign \new_[10840]_  = \new_[11588]_  & \new_[13744]_ ;
  assign \new_[10841]_  = \new_[11680]_  & \new_[12071]_ ;
  assign \new_[10842]_  = ~\new_[13413]_  | ~\new_[11655]_  | ~\new_[12865]_ ;
  assign \new_[10843]_  = ~\new_[9188]_  | ~\new_[11626]_ ;
  assign \new_[10844]_  = \new_[12715]_  & \new_[14385]_ ;
  assign \new_[10845]_  = \new_[14003]_  ^ \new_[11791]_ ;
  assign \new_[10846]_  = \new_[9372]_  ^ \new_[12155]_ ;
  assign \new_[10847]_  = \new_[11051]_ ;
  assign \new_[10848]_  = ~\new_[11051]_ ;
  assign \new_[10849]_  = ~\new_[11149]_ ;
  assign \new_[10850]_  = ~\new_[11432]_ ;
  assign \new_[10851]_  = \new_[8658]_  ^ \new_[12184]_ ;
  assign \new_[10852]_  = ~\new_[11158]_ ;
  assign \new_[10853]_  = ~\new_[12365]_  & ~\new_[12328]_ ;
  assign \new_[10854]_  = ~\new_[14261]_  & (~\new_[12144]_  | ~\new_[4683]_ );
  assign \new_[10855]_  = ~\new_[13920]_  | ~\new_[14385]_  | ~\new_[13311]_ ;
  assign \new_[10856]_  = ~\new_[11163]_ ;
  assign \new_[10857]_  = ~\new_[12313]_  & ~\new_[12472]_ ;
  assign \new_[10858]_  = ~\new_[13426]_  | ~\new_[11666]_  | ~\new_[12135]_ ;
  assign \new_[10859]_  = ~\new_[4651]_  & (~\new_[13489]_  | ~\new_[13083]_ );
  assign \new_[10860]_  = ~\new_[11622]_  & ~\new_[12230]_ ;
  assign \new_[10861]_  = ~\new_[12484]_  & ~\new_[12307]_ ;
  assign \new_[10862]_  = ~\new_[11701]_  | ~\new_[12542]_ ;
  assign \new_[10863]_  = ~\new_[12366]_  | (~\new_[12717]_  & ~\new_[12566]_ );
  assign \new_[10864]_  = \new_[11809]_  & \new_[11502]_ ;
  assign \new_[10865]_  = ~\new_[11881]_  & (~\new_[12086]_  | ~\new_[3480]_ );
  assign \new_[10866]_  = ~\new_[11461]_  & (~\new_[12069]_  | ~\new_[3884]_ );
  assign \new_[10867]_  = ~\new_[11729]_  & (~\new_[12148]_  | ~\new_[3691]_ );
  assign \new_[10868]_  = ~\new_[12170]_  & (~\new_[11823]_  | ~\new_[4291]_ );
  assign \new_[10869]_  = ~u1_u1_send_data_r_reg;
  assign \new_[10870]_  = ~\new_[11513]_  & ~\new_[13443]_ ;
  assign \new_[10871]_  = (~\new_[13821]_  | ~\new_[12415]_ ) & (~\new_[6539]_  | ~\new_[12811]_ );
  assign \new_[10872]_  = (~\new_[13849]_  | ~\new_[12415]_ ) & (~\new_[4856]_  | ~\new_[12811]_ );
  assign \new_[10873]_  = (~\new_[6086]_  | ~\new_[12811]_ ) & (~\new_[14102]_  | ~\new_[12415]_ );
  assign \new_[10874]_  = (~\new_[13629]_  | ~\new_[4206]_ ) & (~\new_[14195]_  | ~\new_[4293]_ );
  assign \new_[10875]_  = (~\new_[12366]_  | ~\new_[12374]_ ) & (~\new_[12717]_  | ~\new_[12711]_ );
  assign \new_[10876]_  = ~\new_[6697]_  | ~\new_[12415]_ ;
  assign \new_[10877]_  = (~\new_[13190]_  | ~\new_[3932]_ ) & (~\new_[11912]_  | ~\new_[12706]_ );
  assign \new_[10878]_  = \new_[2865]_  ? \new_[12130]_  : \new_[12837]_ ;
  assign \new_[10879]_  = ~\new_[11665]_  | ~\new_[4795]_ ;
  assign \new_[10880]_  = ~\new_[13736]_  | ~\new_[12970]_ ;
  assign \new_[10881]_  = ~\new_[13535]_  | ~\new_[12970]_ ;
  assign \new_[10882]_  = ~\new_[11691]_  & ~\new_[6008]_ ;
  assign \new_[10883]_  = ~\new_[2552]_  | ~\new_[12415]_ ;
  assign \new_[10884]_  = ~\new_[2860]_  | ~\new_[11437]_ ;
  assign \new_[10885]_  = ~\new_[6249]_  | ~\new_[12811]_ ;
  assign \new_[10886]_  = ~\new_[6262]_  | ~\new_[12811]_ ;
  assign \new_[10887]_  = ~\new_[6286]_  | ~\new_[12811]_ ;
  assign \new_[10888]_  = ~\new_[12404]_  | ~\new_[12678]_ ;
  assign \new_[10889]_  = ~\new_[13324]_  | ~\new_[11652]_  | ~\new_[12530]_ ;
  assign \new_[10890]_  = ~\new_[6292]_  | ~\new_[12811]_ ;
  assign \new_[10891]_  = ~\new_[6310]_  | ~\new_[12415]_ ;
  assign \new_[10892]_  = ~\new_[5111]_  | ~\new_[12415]_ ;
  assign \new_[10893]_  = ~u0_rx_active_reg;
  assign \new_[10894]_  = ~\new_[2807]_  | ~\new_[11663]_ ;
  assign \new_[10895]_  = ~\new_[6263]_  | ~\new_[12811]_ ;
  assign \new_[10896]_  = ~\new_[11509]_  | ~\new_[3890]_ ;
  assign \new_[10897]_  = ~\new_[2804]_  | ~\new_[11663]_ ;
  assign \new_[10898]_  = ~\new_[14267]_  | ~\new_[11489]_ ;
  assign \new_[10899]_  = ~\new_[6253]_  | ~\new_[12811]_ ;
  assign \new_[10900]_  = ~\new_[2788]_  | ~\new_[11663]_ ;
  assign \new_[10901]_  = ~\new_[11663]_  | ~\new_[2861]_ ;
  assign \new_[10902]_  = ~\new_[11711]_  & ~\new_[3314]_ ;
  assign \new_[10903]_  = ~\new_[2501]_  | ~\new_[12415]_ ;
  assign \new_[10904]_  = ~\new_[5489]_  | ~\new_[12415]_ ;
  assign \new_[10905]_  = ~\new_[2809]_  | ~\new_[11437]_ ;
  assign \new_[10906]_  = ~\new_[14079]_  | ~\new_[12415]_ ;
  assign \new_[10907]_  = ~\new_[13848]_  | ~\new_[12811]_ ;
  assign \new_[10908]_  = ~\new_[2806]_  | ~\new_[11663]_ ;
  assign \new_[10909]_  = ~\new_[11437]_  | ~\new_[2810]_ ;
  assign \new_[10910]_  = ~\new_[2859]_  | ~\new_[11437]_ ;
  assign \new_[10911]_  = ~\new_[3716]_  | ~\new_[12415]_ ;
  assign \new_[10912]_  = ~\new_[6291]_  | ~\new_[12811]_ ;
  assign \new_[10913]_  = ~\new_[12811]_  | ~\new_[6257]_ ;
  assign \new_[10914]_  = \new_[13471]_  | \new_[3692]_  | \new_[11509]_  | \new_[3875]_ ;
  assign \new_[10915]_  = ~\new_[2893]_  | ~\new_[11437]_ ;
  assign n8240 = u0_rx_err_reg;
  assign \new_[10917]_  = ~\new_[2805]_  | ~\new_[11663]_ ;
  assign \new_[10918]_  = ~\new_[2808]_  | ~\new_[11663]_ ;
  assign \new_[10919]_  = ~\new_[2833]_  | ~\new_[11437]_ ;
  assign \new_[10920]_  = \new_[13203]_  | \new_[11663]_ ;
  assign \new_[10921]_  = \new_[13204]_  | \new_[11663]_ ;
  assign \new_[10922]_  = \new_[11437]_  | \new_[13203]_ ;
  assign \new_[10923]_  = \new_[11437]_  | \new_[13132]_ ;
  assign \new_[10924]_  = \new_[11437]_  | \new_[12952]_ ;
  assign \new_[10925]_  = \new_[13164]_  | \new_[11663]_ ;
  assign \new_[10926]_  = \new_[12952]_  | \new_[11663]_ ;
  assign \new_[10927]_  = \new_[11437]_  | \new_[13204]_ ;
  assign \new_[10928]_  = \new_[11437]_  | \new_[13170]_ ;
  assign \new_[10929]_  = \new_[13170]_  | \new_[11663]_ ;
  assign \new_[10930]_  = \new_[13156]_  | \new_[11663]_ ;
  assign \new_[10931]_  = \new_[11437]_  | \new_[13185]_ ;
  assign \new_[10932]_  = \new_[13132]_  | \new_[11663]_ ;
  assign \new_[10933]_  = ~\new_[12364]_  & ~\new_[11705]_ ;
  assign \new_[10934]_  = \new_[11437]_  | \new_[13164]_ ;
  assign \new_[10935]_  = \new_[13185]_  | \new_[11663]_ ;
  assign \new_[10936]_  = ~\new_[11664]_  & (~\new_[6526]_  | ~\new_[6696]_ );
  assign \new_[10937]_  = ~\new_[11661]_  & (~\new_[6292]_  | ~\new_[6718]_ );
  assign \new_[10938]_  = ~\new_[11673]_  & (~\new_[6291]_  | ~\new_[12396]_ );
  assign \new_[10939]_  = u0_rx_valid_reg;
  assign \new_[10940]_  = (~\new_[13621]_  | ~\new_[3889]_ ) & (~\new_[13617]_  | ~\new_[3888]_ );
  assign \new_[10941]_  = (~\new_[4608]_  | ~\new_[14453]_ ) & (~\new_[4841]_  | ~\new_[14200]_ );
  assign \new_[10942]_  = (~\new_[4709]_  | ~\new_[14453]_ ) & (~\new_[4818]_  | ~\new_[14200]_ );
  assign \new_[10943]_  = (~\new_[4616]_  | ~\new_[13646]_ ) & (~\new_[4838]_  | ~\new_[13895]_ );
  assign \new_[10944]_  = ~\new_[2991]_  & ~\new_[13155]_ ;
  assign \new_[10945]_  = ~\new_[13327]_  & ~\new_[13858]_ ;
  assign \new_[10946]_  = ~\new_[4794]_  | ~\new_[12416]_ ;
  assign \new_[10947]_  = ~\new_[11330]_ ;
  assign \new_[10948]_  = ~\new_[11490]_  & ~\new_[12160]_ ;
  assign \new_[10949]_  = ~\new_[12592]_  | ~\new_[11695]_ ;
  assign \new_[10950]_  = ~\new_[11332]_ ;
  assign \new_[10951]_  = \new_[9456]_  ^ \new_[12169]_ ;
  assign \new_[10952]_  = \new_[8888]_  ^ \new_[12145]_ ;
  assign \new_[10953]_  = \new_[2868]_  ? \new_[12130]_  : \new_[12807]_ ;
  assign \new_[10954]_  = \new_[11460]_  & \new_[11762]_ ;
  assign \new_[10955]_  = (~\new_[13751]_  | ~\new_[4288]_ ) & (~\new_[13656]_  | ~\new_[4291]_ );
  assign \new_[10956]_  = ~\new_[6526]_  | ~\new_[12811]_ ;
  assign \new_[10957]_  = (~\new_[13742]_  | ~\new_[12415]_ ) & (~\new_[12811]_  | ~\new_[5860]_ );
  assign \new_[10958]_  = \new_[2895]_  ? \new_[12130]_  : \new_[12817]_ ;
  assign \new_[10959]_  = \new_[13409]_  ^ \new_[12194]_ ;
  assign \new_[10960]_  = \new_[5978]_  ? \new_[12047]_  : \new_[13889]_ ;
  assign \new_[10961]_  = u0_u0_ls_se0_r_reg;
  assign \new_[10962]_  = \new_[2866]_  ? \new_[12130]_  : \new_[12652]_ ;
  assign \new_[10963]_  = (~\new_[14070]_  | ~\new_[12415]_ ) & (~\new_[5504]_  | ~\new_[12811]_ );
  assign \new_[10964]_  = \new_[2864]_  ? \new_[12130]_  : \new_[12831]_ ;
  assign \new_[10965]_  = ~\new_[12236]_  | ~\new_[2875]_  | ~\new_[11712]_  | ~\new_[2873]_ ;
  assign \new_[10966]_  = ~\new_[13069]_  | ~\new_[2086]_  | ~\new_[11695]_  | ~\new_[2093]_ ;
  assign \new_[10967]_  = ~\new_[11696]_  & ~\new_[2345]_ ;
  assign \new_[10968]_  = \new_[8700]_  ^ \new_[11749]_ ;
  assign \new_[10969]_  = \new_[12212]_  ^ \new_[4293]_ ;
  assign \new_[10970]_  = \new_[2862]_  ? \new_[12130]_  : \new_[12802]_ ;
  assign \new_[10971]_  = ~\new_[12038]_  & ~\new_[12719]_ ;
  assign \new_[10972]_  = ~\new_[12150]_  & ~\new_[11438]_ ;
  assign \new_[10973]_  = ~\new_[14036]_  | ~\new_[13666]_  | ~\new_[11458]_  | ~\new_[13219]_ ;
  assign \new_[10974]_  = \new_[3471]_  ^ \new_[12140]_ ;
  assign \new_[10975]_  = \new_[2989]_  ^ \new_[11761]_ ;
  assign \new_[10976]_  = \new_[13606]_  ^ \new_[12133]_ ;
  assign n8250 = \new_[4774]_  ^ \new_[12138]_ ;
  assign \new_[10978]_  = \new_[2704]_  ^ \new_[12134]_ ;
  assign \new_[10979]_  = \new_[2863]_  ? \new_[12130]_  : \new_[12822]_ ;
  assign \new_[10980]_  = \new_[2867]_  ? \new_[12130]_  : \new_[12775]_ ;
  assign \new_[10981]_  = ~\\u4_u1_dma_out_left_reg[0] ;
  assign \new_[10982]_  = \\u0_u0_idle_cnt1_next_reg[2] ;
  assign \new_[10983]_  = \new_[11459]_  | \new_[13606]_ ;
  assign \new_[10984]_  = ~\new_[11457]_  & ~\new_[6232]_ ;
  assign \new_[10985]_  = \new_[11458]_  & \new_[3025]_ ;
  assign \new_[10986]_  = ~\new_[11840]_  | (~\new_[11739]_  & ~\new_[12395]_ );
  assign \new_[10987]_  = ~\new_[11848]_  | (~\new_[11744]_  & ~\new_[12232]_ );
  assign \new_[10988]_  = ~\new_[11861]_  | (~\new_[11743]_  & ~\new_[12424]_ );
  assign \new_[10989]_  = ~\new_[11870]_  | (~\new_[11928]_  & ~\new_[12405]_ );
  assign \new_[10990]_  = ~\new_[2991]_  & ~\new_[13469]_ ;
  assign \new_[10991]_  = ~\new_[11859]_  | (~\new_[11735]_  & ~\new_[12223]_ );
  assign \new_[10992]_  = ~\new_[14211]_  | ~\new_[14036]_  | ~\new_[11458]_  | ~\new_[3025]_ ;
  assign \new_[10993]_  = ~\new_[11427]_ ;
  assign \new_[10994]_  = ~\new_[11844]_  | (~\new_[11740]_  & ~\new_[12320]_ );
  assign \new_[10995]_  = ~\new_[11906]_  | (~\new_[11741]_  & ~\new_[12233]_ );
  assign \new_[10996]_  = ~\new_[11833]_  | (~\new_[11738]_  & ~\new_[12309]_ );
  assign \new_[10997]_  = ~\new_[12612]_  | ~\new_[11565]_  | ~\new_[13029]_ ;
  assign \new_[10998]_  = \new_[9421]_  ^ \new_[11748]_ ;
  assign \new_[10999]_  = ~\new_[6259]_  | ~\new_[12811]_ ;
  assign \new_[11000]_  = ~\new_[4819]_  & ~\new_[14508]_ ;
  assign n8270 = \new_[11764]_  ^ \new_[11739]_ ;
  assign n8265 = \new_[12010]_  ^ \new_[11744]_ ;
  assign n8260 = \new_[11785]_  ^ \new_[11743]_ ;
  assign n8275 = \new_[12002]_  ^ \new_[11928]_ ;
  assign \new_[11005]_  = ~\new_[11510]_  & (~\new_[11847]_  | ~\new_[13036]_ );
  assign \new_[11006]_  = ~\new_[11430]_ ;
  assign \new_[11007]_  = ~\new_[12745]_  | ~\new_[14050]_  | ~\new_[3025]_  | ~\new_[11915]_ ;
  assign \new_[11008]_  = ~\new_[11919]_  & ~\new_[11435]_ ;
  assign \new_[11009]_  = ~\new_[11445]_  | ~\new_[4683]_ ;
  assign \new_[11010]_  = ~\new_[11953]_  & ~\new_[11436]_ ;
  assign \new_[11011]_  = ~\new_[11443]_  | ~\new_[12809]_ ;
  assign \new_[11012]_  = \new_[11694]_  | \new_[12315]_ ;
  assign \new_[11013]_  = ~\new_[11528]_  & ~\new_[11740]_ ;
  assign \new_[11014]_  = ~\new_[13489]_  | ~\new_[13083]_  | ~\new_[12238]_ ;
  assign \new_[11015]_  = \new_[2086]_  ^ \new_[12242]_ ;
  assign \new_[11016]_  = \\u1_u2_rd_buf0_reg[2] ;
  assign \new_[11017]_  = \new_[8954]_  ^ \new_[12243]_ ;
  assign \new_[11018]_  = \\u1_u2_rd_buf0_reg[31] ;
  assign \new_[11019]_  = \new_[14204]_  ^ \new_[12260]_ ;
  assign \new_[11020]_  = ~\new_[12882]_  | (~\new_[12402]_  & ~\new_[4620]_ );
  assign \new_[11021]_  = ~\new_[11783]_  | ~\new_[11858]_ ;
  assign \new_[11022]_  = ~\new_[12167]_  | ~\new_[11850]_ ;
  assign \new_[11023]_  = ~\new_[11775]_  | ~\new_[2478]_ ;
  assign \new_[11024]_  = \new_[11775]_  | \new_[2478]_ ;
  assign \new_[11025]_  = ~\new_[13055]_  | ~\new_[13309]_  | ~\new_[12376]_ ;
  assign \new_[11026]_  = \new_[13287]_  | \new_[3482]_  | \new_[11817]_  | \new_[3684]_ ;
  assign \new_[11027]_  = ~\new_[11784]_  | ~\new_[11863]_ ;
  assign \new_[11028]_  = \\u1_u2_rd_buf0_reg[28] ;
  assign \new_[11029]_  = ~\new_[12179]_  | ~\new_[12132]_ ;
  assign \new_[11030]_  = \\u1_u2_rd_buf0_reg[6] ;
  assign n8595 = ~\new_[12751]_  | ~\new_[12942]_  | ~\new_[12761]_  | ~\new_[12839]_ ;
  assign n8600 = ~\new_[12638]_  | ~\new_[12999]_  | ~\new_[12639]_  | ~\new_[12629]_ ;
  assign n8565 = ~\new_[12766]_  | ~\new_[13071]_  | ~\new_[12503]_  | ~\new_[12808]_ ;
  assign n8580 = ~\new_[12843]_  | ~\new_[12958]_  | ~\new_[12633]_  | ~\new_[12768]_ ;
  assign \new_[11035]_  = \new_[13258]_  ^ \new_[2871]_ ;
  assign n8585 = ~\new_[12762]_  | ~\new_[13234]_  | ~\new_[12632]_  | ~\new_[12867]_ ;
  assign n8555 = ~\new_[12743]_  | ~\new_[12961]_  | ~\new_[12636]_  | ~\new_[12764]_ ;
  assign n8560 = ~\new_[12750]_  | ~\new_[12988]_  | ~\new_[12767]_  | ~\new_[12635]_ ;
  assign n8590 = ~\new_[12630]_  | ~\new_[12927]_  | ~\new_[12795]_  | ~\new_[12744]_ ;
  assign \new_[11040]_  = ~\new_[13203]_  & ~\new_[14314]_ ;
  assign \new_[11041]_  = ~\new_[11758]_  | ~\new_[13238]_ ;
  assign \new_[11042]_  = ~\new_[11970]_  & ~\new_[12242]_ ;
  assign \new_[11043]_  = ~\new_[12531]_  & (~\new_[12350]_  | ~\new_[4620]_ );
  assign \new_[11044]_  = \new_[11770]_  & \new_[11765]_ ;
  assign \new_[11045]_  = ~\new_[12106]_  | ~\new_[13479]_ ;
  assign \new_[11046]_  = ~\new_[11878]_  | ~\new_[13335]_ ;
  assign \new_[11047]_  = ~\new_[11773]_  | ~\new_[13334]_ ;
  assign \new_[11048]_  = ~\new_[11735]_ ;
  assign \new_[11049]_  = ~\new_[11738]_ ;
  assign \new_[11050]_  = ~\new_[11740]_ ;
  assign \new_[11051]_  = ~\new_[13940]_  | ~\new_[11771]_  | ~\new_[7670]_ ;
  assign \new_[11052]_  = ~\new_[11741]_ ;
  assign \new_[11053]_  = ~\new_[11892]_  & (~\new_[13595]_  | ~\new_[13464]_ );
  assign \new_[11054]_  = \new_[13932]_  ^ \new_[12492]_ ;
  assign \new_[11055]_  = \new_[14089]_  ^ \new_[12494]_ ;
  assign \new_[11056]_  = \new_[14163]_  ^ \new_[13068]_ ;
  assign \new_[11057]_  = \\u1_u2_rd_buf0_reg[23] ;
  assign \new_[11058]_  = \new_[13236]_  ^ \new_[12393]_ ;
  assign \new_[11059]_  = \new_[12391]_  ^ \new_[12392]_ ;
  assign \new_[11060]_  = \new_[12928]_  ^ \new_[12393]_ ;
  assign \new_[11061]_  = \new_[13230]_  ^ \new_[12392]_ ;
  assign \new_[11062]_  = \new_[13186]_  ^ \new_[12391]_ ;
  assign \new_[11063]_  = \new_[12393]_  ^ \new_[12392]_ ;
  assign \new_[11064]_  = \new_[12269]_  ^ \new_[12391]_ ;
  assign \new_[11065]_  = \new_[12916]_  ^ \new_[12392]_ ;
  assign \new_[11066]_  = ~\\u4_u1_buf0_orig_m3_reg[1] ;
  assign \new_[11067]_  = \new_[12206]_  | \new_[6343]_ ;
  assign \new_[11068]_  = \new_[12208]_  & \new_[3711]_ ;
  assign \new_[11069]_  = \new_[12722]_  | \new_[13989]_ ;
  assign \new_[11070]_  = \new_[12204]_  & \new_[3888]_ ;
  assign \new_[11071]_  = \new_[12212]_  & \new_[4293]_ ;
  assign \new_[11072]_  = ~\new_[13461]_  | ~\new_[13038]_  | ~\new_[12312]_ ;
  assign \new_[11073]_  = ~\new_[13413]_  | ~\new_[13242]_  | ~\new_[12310]_ ;
  assign \new_[11074]_  = ~\new_[11859]_  & ~\new_[11812]_ ;
  assign \new_[11075]_  = ~\new_[12500]_  | ~\new_[13155]_  | ~\new_[12113]_  | ~\new_[14156]_ ;
  assign \new_[11076]_  = \new_[11842]_  | \new_[12318]_ ;
  assign \new_[11077]_  = \new_[11804]_  | \wb_addr_i[17] ;
  assign \new_[11078]_  = ~\new_[13324]_  | ~\new_[13143]_  | ~\new_[12489]_ ;
  assign \new_[11079]_  = ~\new_[13246]_  | ~\new_[12193]_ ;
  assign \new_[11080]_  = ~\new_[11875]_  | ~\new_[13710]_ ;
  assign \new_[11081]_  = ~\new_[13947]_  | ~\new_[11815]_  | ~\new_[3282]_ ;
  assign \new_[11082]_  = ~\new_[11906]_  & ~\new_[12351]_ ;
  assign \new_[11083]_  = \\u1_u2_rd_buf0_reg[19] ;
  assign \new_[11084]_  = \new_[11866]_  | \new_[12234]_ ;
  assign \new_[11085]_  = \new_[11864]_  | \new_[12230]_ ;
  assign \new_[11086]_  = ~\new_[13355]_  | ~\new_[13010]_  | ~\new_[12447]_ ;
  assign \new_[11087]_  = ~\new_[11833]_  & ~\new_[12017]_ ;
  assign \new_[11088]_  = ~\new_[4683]_  | ~\new_[14261]_  | ~\new_[4666]_  | ~\new_[12362]_ ;
  assign \new_[11089]_  = ~\new_[3463]_  | ~\new_[3475]_  | ~\new_[11737]_  | ~\new_[3435]_ ;
  assign n8325 = n9010 ^ \new_[13891]_ ;
  assign \new_[11091]_  = (~n9130 | ~\new_[12349]_ ) & (~\new_[12275]_  | ~\new_[6241]_ );
  assign \new_[11092]_  = (~\new_[12349]_  | ~n9005) & (~\new_[12275]_  | ~\new_[6239]_ );
  assign \new_[11093]_  = (~\new_[2986]_  | ~\new_[12671]_ ) & (~\new_[12418]_  | ~\new_[13512]_ );
  assign \new_[11094]_  = (~\new_[3471]_  | ~\new_[12671]_ ) & (~\new_[12275]_  | ~\new_[6107]_ );
  assign \new_[11095]_  = (~\new_[12275]_  | ~\new_[6242]_ ) & (~\new_[12418]_  | ~\new_[6610]_ );
  assign \new_[11096]_  = (~\new_[3473]_  | ~\new_[12671]_ ) & (~\new_[12418]_  | ~\new_[6723]_ );
  assign \new_[11097]_  = (~\new_[3435]_  | ~\new_[12671]_ ) & (~\new_[12418]_  | ~\new_[6724]_ );
  assign \new_[11098]_  = (~\new_[12418]_  | ~\new_[14074]_ ) & (~\new_[3475]_  | ~\new_[12671]_ );
  assign \new_[11099]_  = (~\new_[2983]_  | ~\new_[12671]_ ) & (~\new_[12418]_  | ~\new_[13702]_ );
  assign \new_[11100]_  = (~\new_[2984]_  | ~\new_[12671]_ ) & (~\new_[12418]_  | ~\new_[13734]_ );
  assign \new_[11101]_  = (~\new_[2985]_  | ~\new_[12671]_ ) & (~\new_[12418]_  | ~\new_[14164]_ );
  assign SuspendM_pad_o = ~\new_[11479]_ ;
  assign \new_[11103]_  = ~\new_[14118]_  | ~\new_[13438]_  | ~\new_[11963]_  | ~\new_[12696]_ ;
  assign \new_[11104]_  = ~\new_[3895]_  | ~\new_[13501]_  | ~\new_[12109]_  | ~\new_[13218]_ ;
  assign \new_[11105]_  = \new_[13862]_  ? \new_[2042]_  : \new_[12340]_ ;
  assign \new_[11106]_  = \new_[11816]_  & \new_[13099]_ ;
  assign \new_[11107]_  = \new_[12514]_  ^ \new_[12218]_ ;
  assign n8415 = ~\new_[12622]_  & ~\new_[13296]_ ;
  assign n8520 = ~\new_[12803]_  & ~\new_[13296]_ ;
  assign n8540 = ~\new_[12777]_  & ~\new_[13296]_ ;
  assign \new_[11111]_  = ~\new_[11925]_  & ~\new_[6588]_ ;
  assign \new_[11112]_  = ~\new_[11855]_  & ~\new_[6348]_ ;
  assign \new_[11113]_  = \new_[3469]_  & \new_[12671]_ ;
  assign \new_[11114]_  = ~\new_[11820]_  & ~\new_[6461]_ ;
  assign \new_[11115]_  = ~\new_[11926]_  | ~\new_[13407]_ ;
  assign \new_[11116]_  = ~\new_[11913]_  & ~\new_[6324]_ ;
  assign \new_[11117]_  = ~\new_[11820]_  & ~\new_[6370]_ ;
  assign \new_[11118]_  = ~\new_[12052]_  & ~\new_[13407]_ ;
  assign \new_[11119]_  = \new_[12113]_  & \new_[13155]_ ;
  assign \new_[11120]_  = ~\new_[11925]_  & ~\new_[6560]_ ;
  assign \new_[11121]_  = ~\new_[11931]_  & ~\new_[6346]_ ;
  assign \new_[11122]_  = ~\new_[11855]_  & ~\new_[6551]_ ;
  assign \new_[11123]_  = ~\new_[12191]_  | ~\wb_addr_i[4] ;
  assign \new_[11124]_  = ~\new_[11916]_  | ~\new_[13987]_ ;
  assign \new_[11125]_  = \new_[12671]_  & \new_[3474]_ ;
  assign \new_[11126]_  = ~\new_[11913]_  & ~\new_[6322]_ ;
  assign \new_[11127]_  = ~\new_[11921]_  | ~\new_[12177]_ ;
  assign \new_[11128]_  = ~\new_[13172]_  | ~\new_[12031]_  | ~\new_[12528]_ ;
  assign \new_[11129]_  = ~\new_[11956]_  | ~\new_[11965]_ ;
  assign \new_[11130]_  = \new_[12164]_  | \wb_addr_i[4] ;
  assign \new_[11131]_  = ~\new_[12186]_  | ~\new_[11780]_ ;
  assign \new_[11132]_  = \new_[12720]_  & \new_[11922]_ ;
  assign \new_[11133]_  = ~\new_[12964]_  | ~\new_[11759]_  | ~\new_[12628]_ ;
  assign \new_[11134]_  = ~\new_[12162]_  | ~\new_[12542]_ ;
  assign \new_[11135]_  = ~\new_[12600]_  | ~\new_[12857]_ ;
  assign \new_[11136]_  = ~\new_[12542]_  | ~\new_[12563]_ ;
  assign \new_[11137]_  = ~\new_[12872]_  | ~\new_[12615]_ ;
  assign \new_[11138]_  = ~\new_[11883]_  | ~\new_[2932]_ ;
  assign \new_[11139]_  = \new_[11883]_  & \new_[2874]_ ;
  assign \new_[11140]_  = ~\new_[11496]_ ;
  assign \new_[11141]_  = ~\new_[12593]_  | ~\new_[11952]_ ;
  assign \new_[11142]_  = ~\new_[13222]_  | ~\new_[12030]_  | ~\new_[12921]_ ;
  assign \new_[11143]_  = ~\new_[11587]_ ;
  assign \new_[11144]_  = ~\new_[11939]_  | ~\new_[11937]_ ;
  assign \new_[11145]_  = ~\new_[11499]_ ;
  assign \new_[11146]_  = ~\new_[4290]_  | ~\new_[12193]_  | ~\new_[13458]_ ;
  assign \new_[11147]_  = \new_[12603]_  | \new_[12135]_ ;
  assign \new_[11148]_  = ~n8390 | ~\new_[12797]_  | ~\new_[13084]_ ;
  assign \new_[11149]_  = \new_[11957]_  | \wb_addr_i[4] ;
  assign \new_[11150]_  = ~\new_[13198]_  | ~\new_[12034]_  | ~\new_[13011]_ ;
  assign \new_[11151]_  = ~\new_[12105]_  | ~\new_[12872]_ ;
  assign \new_[11152]_  = \new_[11959]_  & \new_[12043]_ ;
  assign \new_[11153]_  = ~\new_[2210]_  | ~\new_[11771]_  | ~\new_[14034]_ ;
  assign \new_[11154]_  = ~\new_[12521]_  | ~\new_[12620]_ ;
  assign \new_[11155]_  = \new_[12569]_  & \new_[11927]_ ;
  assign \new_[11156]_  = ~\new_[12390]_  & ~\new_[12830]_ ;
  assign \new_[11157]_  = ~\new_[12039]_  & (~\new_[13540]_  | ~\new_[3930]_ );
  assign \new_[11158]_  = ~\new_[13771]_  | ~\new_[12200]_  | ~\new_[4161]_ ;
  assign \new_[11159]_  = \new_[12000]_  & \new_[12327]_ ;
  assign \new_[11160]_  = ~\new_[12175]_  & ~\new_[12407]_ ;
  assign \new_[11161]_  = ~\new_[11997]_  | ~\new_[12323]_ ;
  assign \new_[11162]_  = ~\new_[12400]_  & ~\new_[12049]_ ;
  assign \new_[11163]_  = ~\new_[3781]_  | ~\new_[12200]_  | ~\new_[14127]_ ;
  assign \new_[11164]_  = ~\new_[12468]_  & ~\new_[11998]_ ;
  assign \new_[11165]_  = ~\new_[12241]_  & ~\new_[12656]_ ;
  assign \new_[11166]_  = ~\new_[12108]_  & (~\new_[13571]_  | ~\new_[4292]_ );
  assign \new_[11167]_  = ~\new_[12248]_  & ~\new_[11996]_ ;
  assign \new_[11168]_  = ~\new_[12126]_  & ~\new_[12163]_ ;
  assign \new_[11169]_  = ~\new_[11778]_  & ~\new_[12234]_ ;
  assign \new_[11170]_  = ~\new_[12011]_  | ~\new_[11974]_ ;
  assign \new_[11171]_  = ~\new_[12042]_  & (~\new_[13891]_  | ~\new_[3503]_ );
  assign \new_[11172]_  = \new_[12757]_  & \new_[11950]_ ;
  assign \new_[11173]_  = ~\new_[13764]_  & ~\new_[12713]_ ;
  assign \new_[11174]_  = \new_[12511]_  & \new_[11745]_ ;
  assign \new_[11175]_  = ~\new_[12224]_  & ~\new_[11732]_ ;
  assign \new_[11176]_  = ~\new_[12015]_  | ~\new_[12321]_ ;
  assign \new_[11177]_  = ~\new_[12225]_  & ~\new_[12668]_ ;
  assign \new_[11178]_  = \new_[12518]_  & \new_[11962]_ ;
  assign \new_[11179]_  = \new_[12054]_  | \new_[12484]_ ;
  assign \new_[11180]_  = ~\new_[12319]_  & ~\new_[12754]_ ;
  assign \new_[11181]_  = ~\new_[12005]_  | ~\new_[12224]_ ;
  assign \new_[11182]_  = ~\new_[12044]_  & (~\new_[13872]_  | ~\new_[3777]_ );
  assign \new_[11183]_  = ~\new_[12054]_  | ~\new_[12400]_ ;
  assign \new_[11184]_  = \new_[12309]_  | \new_[12017]_ ;
  assign \new_[11185]_  = \new_[12005]_  | \new_[12365]_ ;
  assign \new_[11186]_  = \new_[12223]_  | \new_[11812]_ ;
  assign \new_[11187]_  = \new_[12454]_  & \new_[12011]_ ;
  assign \new_[11188]_  = (~\new_[12354]_  | ~\new_[4811]_ ) & (~\new_[14546]_  | ~\new_[4864]_ );
  assign \new_[11189]_  = (~\new_[12356]_  | ~\new_[4834]_ ) & (~\new_[14546]_  | ~\new_[4619]_ );
  assign \new_[11190]_  = ~\new_[12538]_  & (~\new_[12263]_  | ~\new_[13153]_ );
  assign \new_[11191]_  = ~\new_[12702]_  & (~\new_[12436]_  | ~\new_[13114]_ );
  assign \new_[11192]_  = ~\new_[12707]_  & (~\new_[12257]_  | ~\new_[13331]_ );
  assign \new_[11193]_  = ~\new_[11943]_  & ~\new_[12789]_ ;
  assign \new_[11194]_  = ~\new_[11844]_  & ~\new_[12425]_ ;
  assign \new_[11195]_  = ~\new_[12279]_  & (~\new_[12380]_  | ~\new_[3693]_ );
  assign \new_[11196]_  = ~\new_[2210]_  | ~\new_[13443]_ ;
  assign \new_[11197]_  = ~\new_[12219]_  & (~\new_[12373]_  | ~\new_[3316]_ );
  assign \new_[11198]_  = ~\new_[11949]_  | (~\new_[6299]_  & ~\new_[12524]_ );
  assign \new_[11199]_  = ~\new_[12367]_  & (~\new_[12369]_  | ~\new_[4073]_ );
  assign \new_[11200]_  = ~\new_[11934]_  & (~\new_[12779]_  | ~\new_[3504]_ );
  assign \new_[11201]_  = ~\new_[11746]_  | (~\new_[6367]_  & ~\new_[12690]_ );
  assign \new_[11202]_  = ~\new_[11938]_  & (~\new_[12832]_  | ~\new_[4812]_ );
  assign \new_[11203]_  = ~\new_[12102]_  & (~\new_[12796]_  | ~\new_[4816]_ );
  assign \new_[11204]_  = ~\new_[12335]_  | (~\new_[12985]_  & ~\new_[12719]_ );
  assign \new_[11205]_  = ~\new_[11940]_  & (~\new_[12796]_  | ~\new_[4839]_ );
  assign \new_[11206]_  = ~\new_[13443]_  | ~\new_[13189]_ ;
  assign \new_[11207]_  = ~\new_[11555]_ ;
  assign \new_[11208]_  = ~\new_[11879]_  & (~\new_[12832]_  | ~\new_[4835]_ );
  assign \new_[11209]_  = ~\new_[12451]_  & (~\new_[12427]_  | ~\new_[3481]_ );
  assign \new_[11210]_  = ~\new_[11559]_ ;
  assign \new_[11211]_  = ~\new_[11560]_ ;
  assign \new_[11212]_  = ~\new_[11948]_  & (~\new_[12496]_  | ~\new_[3711]_ );
  assign \new_[11213]_  = ~\new_[11582]_ ;
  assign \new_[11214]_  = ~\new_[11571]_ ;
  assign \new_[11215]_  = \\u1_u2_rd_buf0_reg[24] ;
  assign \new_[11216]_  = \\u1_u2_rd_buf0_reg[18] ;
  assign \new_[11217]_  = \\u1_u2_rd_buf0_reg[10] ;
  assign \new_[11218]_  = \\u1_u2_rd_buf0_reg[4] ;
  assign \new_[11219]_  = ~\new_[13500]_  & ~\new_[12530]_ ;
  assign \new_[11220]_  = ~\new_[11872]_  | (~\new_[13078]_  & ~\new_[12906]_ );
  assign \new_[11221]_  = ~\new_[11873]_  | (~\new_[12955]_  & ~\new_[13206]_ );
  assign n8450 = \sram_data_i[8]  ? \new_[12381]_  : \new_[10638]_ ;
  assign n8455 = \sram_data_i[18]  ? \new_[12381]_  : \new_[10639]_ ;
  assign n8495 = \sram_data_i[22]  ? \new_[12381]_  : \new_[10647]_ ;
  assign n8525 = \sram_data_i[16]  ? \new_[12381]_  : \new_[10656]_ ;
  assign n8500 = \sram_data_i[15]  ? \new_[12381]_  : \new_[10648]_ ;
  assign n8505 = \sram_data_i[23]  ? \new_[12381]_  : \new_[10649]_ ;
  assign n8480 = \sram_data_i[5]  ? \new_[12381]_  : \new_[10644]_ ;
  assign \new_[11229]_  = ~\new_[12149]_  & ~\new_[13456]_ ;
  assign n8465 = \sram_data_i[14]  ? \new_[12381]_  : \new_[10641]_ ;
  assign \new_[11231]_  = ~\new_[12111]_  | ~\new_[12521]_ ;
  assign \new_[11232]_  = ~\new_[11692]_ ;
  assign \new_[11233]_  = \new_[9471]_  ^ \new_[12403]_ ;
  assign \new_[11234]_  = ~\new_[11625]_ ;
  assign \new_[11235]_  = ~\new_[14167]_  | ~\new_[12182]_ ;
  assign \new_[11236]_  = ~\new_[12142]_  & ~\new_[6250]_ ;
  assign \new_[11237]_  = ~\new_[14740]_  & ~\new_[11930]_ ;
  assign \new_[11238]_  = ~\new_[14155]_  & ~\new_[12865]_ ;
  assign \new_[11239]_  = ~\new_[12076]_  & ~\new_[5998]_ ;
  assign \new_[11240]_  = ~\new_[11557]_ ;
  assign \new_[11241]_  = ~\new_[6319]_  & ~\new_[13134]_ ;
  assign \new_[11242]_  = \new_[12462]_  & \new_[12089]_ ;
  assign \new_[11243]_  = ~\new_[13848]_  & ~\new_[12785]_ ;
  assign \new_[11244]_  = \new_[12135]_  | \new_[4794]_ ;
  assign \new_[11245]_  = \new_[12077]_  & \new_[12727]_ ;
  assign \new_[11246]_  = ~\new_[11811]_  & ~\new_[13426]_ ;
  assign n8470 = ~\new_[12840]_  & ~\new_[13263]_ ;
  assign \new_[11248]_  = ~\new_[12372]_  | ~\new_[12057]_ ;
  assign \new_[11249]_  = ~\new_[6743]_  | ~\new_[12811]_ ;
  assign \new_[11250]_  = ~\new_[12121]_  & ~\new_[2548]_ ;
  assign \new_[11251]_  = ~\new_[14142]_  | ~\new_[12415]_ ;
  assign \new_[11252]_  = ~\new_[13863]_  | ~\new_[12415]_ ;
  assign \new_[11253]_  = ~\new_[5999]_  & ~\new_[13350]_ ;
  assign n8355 = ~\new_[12650]_  & ~\new_[13263]_ ;
  assign \new_[11255]_  = ~\new_[7670]_  | ~\new_[12160]_ ;
  assign \new_[11256]_  = \new_[12097]_  & \new_[12752]_ ;
  assign \new_[11257]_  = ~\new_[12135]_  & ~\new_[13426]_ ;
  assign n8400 = ~\new_[11702]_ ;
  assign \new_[11259]_  = ~\new_[13614]_  | ~\new_[12415]_ ;
  assign \new_[11260]_  = ~\new_[12062]_  | ~\new_[13359]_ ;
  assign \new_[11261]_  = ~\new_[6286]_  & ~\new_[12690]_ ;
  assign n8345 = ~\new_[12835]_  & ~\new_[13263]_ ;
  assign \new_[11263]_  = ~\new_[12821]_  & ~\new_[12591]_ ;
  assign \new_[11264]_  = ~\new_[12565]_  | ~\new_[4616]_ ;
  assign \new_[11265]_  = ~\new_[6250]_  | ~\new_[12811]_ ;
  assign \new_[11266]_  = ~\new_[12377]_  | ~\new_[12053]_ ;
  assign n8405 = \new_[12040]_  | TxValid_pad_o;
  assign \new_[11268]_  = ~\new_[11606]_ ;
  assign \new_[11269]_  = ~\new_[13156]_  & ~\new_[14314]_ ;
  assign \new_[11270]_  = ~\new_[14231]_  | ~\new_[12415]_ ;
  assign \new_[11271]_  = ~\new_[6251]_  & ~\new_[12524]_ ;
  assign \new_[11272]_  = \new_[12066]_  & \new_[12358]_ ;
  assign \new_[11273]_  = ~\new_[13170]_  & ~\new_[14314]_ ;
  assign \new_[11274]_  = ~\new_[14151]_  | ~\new_[12415]_ ;
  assign \new_[11275]_  = ~\new_[11716]_ ;
  assign \new_[11276]_  = ~\new_[6274]_  & ~\new_[12911]_ ;
  assign \new_[11277]_  = ~\new_[13204]_  & ~\new_[14314]_ ;
  assign \new_[11278]_  = ~\new_[12080]_  & ~\new_[12574]_ ;
  assign n8360 = ~\new_[12502]_  & ~\new_[13263]_ ;
  assign \new_[11280]_  = ~\new_[13564]_  | ~\new_[12415]_ ;
  assign \new_[11281]_  = ~\new_[13704]_  | ~\new_[12415]_ ;
  assign \new_[11282]_  = ~\new_[12956]_  & ~\new_[12070]_ ;
  assign \new_[11283]_  = ~\new_[13164]_  & ~\new_[14314]_ ;
  assign \new_[11284]_  = ~\new_[12080]_  | ~\new_[2870]_ ;
  assign \new_[11285]_  = ~\new_[12952]_  & ~\new_[14314]_ ;
  assign \new_[11286]_  = ~\new_[13132]_  & ~\new_[14314]_ ;
  assign \new_[11287]_  = ~\new_[13048]_  & ~\new_[12864]_ ;
  assign \new_[11288]_  = ~\new_[13161]_  & ~\new_[12656]_ ;
  assign \new_[11289]_  = ~\new_[12272]_  | ~\new_[12087]_ ;
  assign \new_[11290]_  = ~\new_[12855]_  & ~\new_[12749]_ ;
  assign \new_[11291]_  = ~\new_[13056]_  & ~\new_[12830]_ ;
  assign \new_[11292]_  = ~\new_[13244]_  & ~\new_[12668]_ ;
  assign \new_[11293]_  = ~\new_[12923]_  & ~\new_[12754]_ ;
  assign \new_[11294]_  = ~\new_[12091]_  & (~\new_[6549]_  | ~\new_[6718]_ );
  assign \new_[11295]_  = ~\new_[12083]_  & (~\new_[6279]_  | ~\new_[6696]_ );
  assign \new_[11296]_  = ~\new_[12063]_  & (~\new_[6696]_  | ~\new_[6261]_ );
  assign \new_[11297]_  = ~\new_[11892]_  & (~\new_[13595]_  | ~\new_[13138]_ );
  assign \new_[11298]_  = ~\new_[12065]_  & (~\new_[6293]_  | ~\new_[6716]_ );
  assign \new_[11299]_  = ~\new_[12123]_  & (~\new_[6020]_  | ~\new_[6260]_ );
  assign \new_[11300]_  = \new_[2869]_  ^ \new_[4923]_ ;
  assign \new_[11301]_  = \new_[2872]_  ^ \new_[4798]_ ;
  assign \new_[11302]_  = ~\new_[12081]_  & (~\new_[6281]_  | ~\new_[6718]_ );
  assign \new_[11303]_  = ~\new_[12072]_  & (~\new_[6089]_  | ~\new_[6020]_ );
  assign \new_[11304]_  = ~\new_[12093]_  & (~\new_[6547]_  | ~\new_[6696]_ );
  assign \new_[11305]_  = ~\new_[12154]_  & ~\new_[12078]_ ;
  assign \new_[11306]_  = ~\new_[12095]_  & ~\new_[12064]_ ;
  assign \new_[11307]_  = ~\new_[12041]_  & ~\new_[13361]_ ;
  assign \new_[11308]_  = ~\new_[12171]_  & ~\new_[13430]_ ;
  assign \new_[11309]_  = ~\new_[11817]_  | ~\new_[3712]_ ;
  assign \new_[11310]_  = \new_[12084]_  & \new_[12545]_ ;
  assign n8245 = ~\new_[11651]_ ;
  assign \new_[11312]_  = (~\new_[13631]_  | ~\new_[3788]_ ) & (~\new_[13980]_  | ~\new_[3711]_ );
  assign \new_[11313]_  = (~\new_[4695]_  | ~\new_[13646]_ ) & (~\new_[4815]_  | ~\new_[13895]_ );
  assign \new_[11314]_  = (~\new_[2870]_  | ~\new_[14790]_ ) & (~\new_[2871]_  | ~\new_[13096]_ );
  assign \new_[11315]_  = (~\new_[4812]_  | ~\new_[13861]_ ) & (~\new_[4814]_  | ~\new_[14790]_ );
  assign \new_[11316]_  = ~\new_[2870]_  & (~\new_[14790]_  | ~\new_[2871]_ );
  assign n8330 = n9020 ^ \new_[13571]_ ;
  assign \new_[11318]_  = ~\new_[12055]_  | ~\new_[13294]_ ;
  assign \new_[11319]_  = ~\new_[13754]_  | ~\new_[11806]_  | ~\new_[3283]_ ;
  assign n8335 = n9015 ^ \new_[13540]_ ;
  assign \new_[11321]_  = ~\new_[11757]_  | ~\new_[12600]_ ;
  assign \new_[11322]_  = \new_[2927]_  ^ \new_[6696]_ ;
  assign \new_[11323]_  = ~\new_[14167]_  | ~n8390;
  assign \new_[11324]_  = ~\new_[11490]_ ;
  assign \new_[11325]_  = ~\new_[11756]_  & ~\new_[11929]_ ;
  assign \new_[11326]_  = ~\new_[12246]_  & (~\new_[12440]_  | ~\new_[3477]_ );
  assign \new_[11327]_  = \\u1_u2_rd_buf0_reg[30] ;
  assign \new_[11328]_  = ~\new_[2857]_  & ~\new_[14200]_ ;
  assign \new_[11329]_  = \new_[11822]_  | \new_[12407]_ ;
  assign \new_[11330]_  = ~\new_[4842]_  & ~\new_[14508]_ ;
  assign \new_[11331]_  = ~\new_[13469]_  & ~\new_[13267]_ ;
  assign \new_[11332]_  = ~\new_[13247]_  & ~\new_[12185]_ ;
  assign \new_[11333]_  = ~\new_[11931]_  & ~\new_[6351]_ ;
  assign \new_[11334]_  = \\u1_u2_rd_buf0_reg[27] ;
  assign \new_[11335]_  = ~\new_[13288]_  | ~\new_[12082]_  | ~\new_[13616]_ ;
  assign \new_[11336]_  = ~\new_[13185]_  & ~\new_[14314]_ ;
  assign \new_[11337]_  = (~\new_[14015]_  | ~\new_[3505]_ ) & (~\new_[13914]_  | ~\new_[3504]_ );
  assign \new_[11338]_  = ~\new_[12251]_  & (~\new_[12353]_  | ~\new_[13438]_ );
  assign n8460 = \sram_data_i[28]  ? \new_[12381]_  : \new_[10640]_ ;
  assign n8570 = \sram_data_i[11]  ? \new_[12381]_  : \new_[10694]_ ;
  assign n8385 = \sram_data_i[21]  ? \new_[12381]_  : \new_[10568]_ ;
  assign n8380 = \sram_data_i[24]  ? \new_[12381]_  : \new_[10552]_ ;
  assign n8425 = \sram_data_i[27]  ? \new_[12381]_  : \new_[10633]_ ;
  assign n8550 = \sram_data_i[10]  ? \new_[12381]_  : \new_[10674]_ ;
  assign n8535 = ~\new_[12621]_  & ~\new_[13296]_ ;
  assign \new_[11346]_  = \\u1_u2_rd_buf0_reg[3] ;
  assign n8485 = \sram_data_i[9]  ? \new_[12381]_  : \new_[10645]_ ;
  assign n8430 = \sram_data_i[3]  ? \new_[12381]_  : \new_[10634]_ ;
  assign \new_[11349]_  = \\u1_u2_rd_buf0_reg[5] ;
  assign n8395 = ~\new_[11603]_ ;
  assign n8475 = \sram_data_i[6]  ? \new_[12381]_  : \new_[10643]_ ;
  assign \new_[11352]_  = \\u1_u2_rd_buf0_reg[8] ;
  assign n8370 = \sram_data_i[30]  ? \new_[12381]_  : \new_[10515]_ ;
  assign \new_[11354]_  = \\u1_u2_rd_buf0_reg[26] ;
  assign \new_[11355]_  = \\u1_u2_rd_buf0_reg[14] ;
  assign \new_[11356]_  = ~\new_[4817]_  | ~\new_[12610]_ ;
  assign n8350 = ~\new_[11626]_ ;
  assign \new_[11358]_  = ~\new_[11649]_ ;
  assign n8365 = \sram_data_i[31]  ? \new_[12381]_  : \new_[10507]_ ;
  assign n8320 = \sram_data_i[1]  ? \new_[12381]_  : \new_[10359]_ ;
  assign n8445 = \sram_data_i[2]  ? \new_[12381]_  : \new_[10637]_ ;
  assign \new_[11362]_  = ~\new_[12740]_  | ~\new_[3509]_ ;
  assign \new_[11363]_  = \\u1_u2_rd_buf0_reg[0] ;
  assign \new_[11364]_  = \\u1_u2_rd_buf0_reg[1] ;
  assign \new_[11365]_  = \\u1_u2_rd_buf0_reg[29] ;
  assign n8375 = \sram_data_i[7]  ? \new_[12381]_  : \new_[10547]_ ;
  assign n8490 = \sram_data_i[20]  ? \new_[12381]_  : \new_[10646]_ ;
  assign \new_[11368]_  = \new_[12210]_  & \new_[3504]_ ;
  assign \new_[11369]_  = ~\new_[13563]_  | ~\new_[12415]_ ;
  assign n8530 = \sram_data_i[4]  ? \new_[12381]_  : \new_[10664]_ ;
  assign \new_[11371]_  = \new_[11763]_  & \new_[12141]_ ;
  assign n8515 = \sram_data_i[17]  ? \new_[12381]_  : \new_[10652]_ ;
  assign \new_[11373]_  = ~\new_[11712]_ ;
  assign n8545 = \sram_data_i[29]  ? \new_[12381]_  : \new_[10669]_ ;
  assign n8435 = \sram_data_i[0]  ? \new_[12381]_  : \new_[10635]_ ;
  assign n8315 = \sram_data_i[19]  ? \new_[12381]_  : \new_[10358]_ ;
  assign \new_[11377]_  = ~\new_[2992]_  & ~\new_[13398]_ ;
  assign \new_[11378]_  = \\u1_u2_rd_buf0_reg[9] ;
  assign \new_[11379]_  = \new_[11766]_  & \new_[12136]_ ;
  assign \new_[11380]_  = \\u1_u2_rd_buf0_reg[21] ;
  assign \new_[11381]_  = \\u1_u2_rd_buf0_reg[20] ;
  assign \new_[11382]_  = \\u1_u2_rd_buf0_reg[16] ;
  assign \new_[11383]_  = \\u1_u2_rd_buf0_reg[17] ;
  assign \new_[11384]_  = \\u1_u2_rd_buf0_reg[7] ;
  assign n8575 = \sram_data_i[13]  ? \new_[12381]_  : \new_[10695]_ ;
  assign \new_[11386]_  = \\u1_u2_rd_buf0_reg[22] ;
  assign \new_[11387]_  = \\u1_u2_rd_buf0_reg[13] ;
  assign \new_[11388]_  = ~\new_[11762]_  & ~\new_[6300]_ ;
  assign n8510 = \sram_data_i[25]  ? \new_[12381]_  : \new_[10651]_ ;
  assign \new_[11390]_  = \\u1_u2_rd_buf0_reg[25] ;
  assign \new_[11391]_  = \\u1_u2_rd_buf0_reg[12] ;
  assign \new_[11392]_  = ~\new_[13710]_  | ~\new_[4683]_  | ~\new_[12138]_  | ~\new_[13140]_ ;
  assign \new_[11393]_  = ~\new_[14185]_  | ~\new_[13694]_  | ~\new_[12133]_  | ~\new_[13121]_ ;
  assign \new_[11394]_  = \new_[12124]_  | \new_[12610]_ ;
  assign \new_[11395]_  = \new_[9405]_  ^ \new_[12217]_ ;
  assign \new_[11396]_  = \new_[2091]_  ^ \new_[13139]_ ;
  assign \new_[11397]_  = \new_[8826]_  ^ \new_[12475]_ ;
  assign \new_[11398]_  = \\u1_u2_rd_buf0_reg[15] ;
  assign \new_[11399]_  = \\u1_u2_rd_buf0_reg[11] ;
  assign \new_[11400]_  = ~\new_[12019]_  | ~\new_[12199]_ ;
  assign n8440 = \sram_data_i[12]  ? \new_[12381]_  : \new_[10636]_ ;
  assign n8420 = \sram_data_i[26]  ? \new_[12381]_  : \new_[10632]_ ;
  assign \new_[11403]_  = \new_[13799]_  ? \new_[10715]_  : \new_[12495]_ ;
  assign \new_[11404]_  = \new_[2875]_  | \new_[14200]_ ;
  assign \new_[11405]_  = ~\new_[11932]_  | (~\new_[13035]_  & ~\new_[13046]_ );
  assign \new_[11406]_  = ~\new_[11765]_  & ~\new_[3715]_ ;
  assign \new_[11407]_  = ~\new_[12195]_  & ~\new_[2344]_ ;
  assign \new_[11408]_  = \new_[12138]_  & \new_[4774]_ ;
  assign n8410 = ~\new_[11597]_ ;
  assign \new_[11410]_  = ~\new_[12133]_  | ~\new_[3038]_ ;
  assign \new_[11411]_  = ~\new_[12136]_  & ~\new_[3342]_ ;
  assign \new_[11412]_  = \new_[12140]_  & \new_[3471]_ ;
  assign \new_[11413]_  = ~\new_[12141]_  & ~\new_[3997]_ ;
  assign \new_[11414]_  = ~\new_[11769]_  & ~\new_[3510]_ ;
  assign \new_[11415]_  = ~\new_[11768]_  & ~\new_[6368]_ ;
  assign n8605 = ~\new_[11724]_ ;
  assign \new_[11417]_  = ~\new_[12236]_  | ~\new_[12196]_  | ~\new_[12956]_ ;
  assign \new_[11418]_  = ~\new_[11578]_ ;
  assign \new_[11419]_  = \new_[2924]_  ^ \new_[6718]_ ;
  assign \new_[11420]_  = ~\new_[12090]_  & (~\new_[6002]_  | ~\new_[6020]_ );
  assign \new_[11421]_  = \new_[4500]_  ^ \new_[12269]_ ;
  assign \new_[11422]_  = \new_[12578]_  & \new_[12140]_ ;
  assign \new_[11423]_  = ~\new_[13970]_  | ~\new_[14185]_  | ~\new_[12133]_  | ~\new_[3038]_ ;
  assign \new_[11424]_  = ~\new_[12037]_  & (~\new_[6718]_  | ~\new_[6109]_ );
  assign \new_[11425]_  = ~\new_[12617]_  | ~\new_[12437]_ ;
  assign \new_[11426]_  = ~\new_[11585]_ ;
  assign \new_[11427]_  = ~\new_[2836]_  | ~\new_[12196]_  | ~\new_[12956]_ ;
  assign \new_[11428]_  = \new_[2926]_  ^ \new_[12396]_ ;
  assign \new_[11429]_  = ~\new_[14315]_ ;
  assign \new_[11430]_  = ~n8870 | ~\new_[11792]_ ;
  assign \new_[11431]_  = u0_u0_ps_cnt_clr_reg;
  assign \new_[11432]_  = ~\new_[12109]_  | ~\new_[13514]_ ;
  assign \new_[11433]_  = ~\new_[12242]_  & ~\new_[12316]_ ;
  assign \new_[11434]_  = ~\new_[13108]_  | ~\new_[12385]_  | ~\new_[13286]_ ;
  assign \new_[11435]_  = ~\new_[12556]_  | ~\new_[13391]_  | ~\new_[12582]_ ;
  assign \new_[11436]_  = ~\new_[12710]_  | ~\new_[13276]_  | ~\new_[12788]_ ;
  assign \new_[11437]_  = ~\new_[11730]_ ;
  assign \new_[11438]_  = ~\new_[12693]_  | ~\new_[13318]_  | ~\new_[12723]_ ;
  assign \new_[11439]_  = ~n8945 & ~\new_[12471]_ ;
  assign \new_[11440]_  = ~\new_[12725]_  | ~\new_[12455]_ ;
  assign \new_[11441]_  = ~\new_[12429]_  & (~\new_[2343]_  | ~\new_[13020]_ );
  assign \new_[11442]_  = ~\new_[12920]_  | ~\new_[13303]_  | ~\new_[13323]_  | ~\new_[13474]_ ;
  assign \new_[11443]_  = ~\new_[13392]_  & (~\new_[12913]_  | ~\new_[4651]_ );
  assign \new_[11444]_  = ~\new_[12364]_  | ~\new_[14156]_ ;
  assign \new_[11445]_  = ~\new_[4780]_  | ~\new_[4774]_  | ~\new_[12861]_  | ~\new_[12892]_ ;
  assign \new_[11446]_  = ~\new_[12440]_  | ~\new_[13643]_ ;
  assign \new_[11447]_  = \new_[2929]_  ^ \new_[6716]_ ;
  assign \new_[11448]_  = ~\new_[12487]_  & ~\new_[2477]_ ;
  assign \new_[11449]_  = \new_[2737]_  ^ \new_[12888]_ ;
  assign \new_[11450]_  = \new_[9412]_  ^ \new_[12585]_ ;
  assign n8655 = \new_[4780]_  ^ \new_[12892]_ ;
  assign \new_[11452]_  = \new_[8701]_  ^ \new_[12554]_ ;
  assign \new_[11453]_  = \new_[12896]_  ^ \new_[12584]_ ;
  assign \new_[11454]_  = \new_[12884]_  ^ \new_[12555]_ ;
  assign \new_[11455]_  = (~\new_[12901]_  | ~\new_[11727]_ ) & (~\new_[13315]_  | ~\new_[3470]_ );
  assign \new_[11456]_  = ~\new_[12687]_  | ~\new_[12482]_ ;
  assign \new_[11457]_  = ~\new_[12557]_  | ~\new_[13761]_ ;
  assign \new_[11458]_  = \new_[12494]_  & \new_[14089]_ ;
  assign \new_[11459]_  = ~\new_[12898]_  & ~\new_[3037]_ ;
  assign \new_[11460]_  = \new_[12720]_  | \new_[13747]_ ;
  assign \new_[11461]_  = ~\new_[6009]_  & ~\new_[13011]_ ;
  assign \new_[11462]_  = ~\new_[11900]_ ;
  assign \new_[11463]_  = \new_[2870]_  ^ \new_[2932]_ ;
  assign \new_[11464]_  = ~\new_[13403]_  | ~\new_[12860]_  | ~\new_[12540]_ ;
  assign \new_[11465]_  = ~\new_[12262]_  & ~\new_[4798]_ ;
  assign \new_[11466]_  = \new_[12474]_  | \new_[13020]_ ;
  assign \new_[11467]_  = ~\new_[13006]_  | ~\new_[12214]_ ;
  assign \new_[11468]_  = ~\new_[13074]_  | ~\new_[12317]_ ;
  assign \new_[11469]_  = \new_[12270]_  & \new_[12494]_ ;
  assign \new_[11470]_  = ~\new_[13182]_  | ~\new_[12409]_ ;
  assign \new_[11471]_  = (~\new_[2717]_  | ~\new_[12671]_ ) & (~\new_[12519]_  | ~\new_[5617]_ );
  assign \new_[11472]_  = (~\new_[2927]_  | ~\new_[12671]_ ) & (~\new_[12519]_  | ~\new_[5123]_ );
  assign \new_[11473]_  = (~\new_[2926]_  | ~\new_[12671]_ ) & (~\new_[12519]_  | ~\new_[4778]_ );
  assign \new_[11474]_  = (~\new_[2924]_  | ~\new_[12671]_ ) & (~\new_[12519]_  | ~\new_[4501]_ );
  assign \new_[11475]_  = (~\new_[2925]_  | ~\new_[12671]_ ) & (~\new_[12519]_  | ~\new_[3878]_ );
  assign \new_[11476]_  = ~\new_[13167]_ ;
  assign \new_[11477]_  = (~\new_[2987]_  | ~\new_[12671]_ ) & (~\new_[12519]_  | ~\new_[2573]_ );
  assign \new_[11478]_  = (~\new_[2962]_  | ~\new_[12671]_ ) & (~\new_[12519]_  | ~\new_[5757]_ );
  assign \new_[11479]_  = (~\new_[13699]_  | ~\LineState_pad_i[1] ) & (~\new_[12586]_  | ~n9005);
  assign \new_[11480]_  = ~\new_[12122]_ ;
  assign \new_[11481]_  = \new_[12645]_  ^ \new_[13169]_ ;
  assign \new_[11482]_  = ~\new_[6249]_  & ~\new_[12441]_ ;
  assign \new_[11483]_  = ~\new_[12276]_  & ~\new_[6853]_ ;
  assign \new_[11484]_  = ~\new_[13167]_ ;
  assign \new_[11485]_  = \new_[12673]_  & \new_[12272]_ ;
  assign \new_[11486]_  = ~\new_[12276]_  & ~\new_[6302]_ ;
  assign \new_[11487]_  = ~\new_[12417]_  & ~\new_[13407]_ ;
  assign \new_[11488]_  = ~\new_[12261]_  | ~\new_[13366]_ ;
  assign \new_[11489]_  = ~\new_[13167]_ ;
  assign \new_[11490]_  = ~\new_[7856]_  | ~\new_[13419]_  | ~\new_[12800]_ ;
  assign \new_[11491]_  = ~\new_[12277]_  | ~\new_[12625]_ ;
  assign \new_[11492]_  = ~\new_[12418]_  | ~\new_[6721]_ ;
  assign \new_[11493]_  = ~\new_[13408]_  | ~\new_[12349]_ ;
  assign \new_[11494]_  = ~\new_[12418]_  | ~\new_[6722]_ ;
  assign \new_[11495]_  = ~\new_[11804]_ ;
  assign \new_[11496]_  = ~wb_we_i & ~\new_[12324]_ ;
  assign \new_[11497]_  = ~\new_[12331]_  & ~\new_[12332]_ ;
  assign \new_[11498]_  = ~\new_[12561]_  | ~\new_[12256]_ ;
  assign \new_[11499]_  = n8645 & \new_[8959]_ ;
  assign \new_[11500]_  = ~\new_[12418]_  | ~\new_[6609]_ ;
  assign \new_[11501]_  = ~\new_[11809]_ ;
  assign \new_[11502]_  = ~\new_[12919]_  | ~\new_[12355]_  | ~\new_[13470]_ ;
  assign \new_[11503]_  = ~\new_[12706]_  | ~\new_[12291]_ ;
  assign \new_[11504]_  = ~\new_[13128]_  | ~\new_[12261]_ ;
  assign \new_[11505]_  = \new_[12462]_  & \new_[13395]_ ;
  assign \new_[11506]_  = ~\new_[12881]_  | ~\new_[12401]_ ;
  assign \new_[11507]_  = ~\new_[12288]_  & ~\new_[13438]_ ;
  assign \new_[11508]_  = ~\new_[12418]_  | ~\new_[6611]_ ;
  assign \new_[11509]_  = ~\new_[12714]_  | ~\new_[12466]_ ;
  assign \new_[11510]_  = ~\new_[11752]_ ;
  assign \new_[11511]_  = ~\new_[12972]_  & ~\new_[12330]_ ;
  assign \new_[11512]_  = ~\new_[12329]_  & ~\new_[12220]_ ;
  assign \new_[11513]_  = ~\new_[13850]_  | ~\new_[13189]_  | ~\new_[13419]_  | ~\new_[2193]_ ;
  assign \new_[11514]_  = ~\new_[11780]_ ;
  assign \new_[11515]_  = ~\new_[12747]_  | ~\new_[12305]_ ;
  assign \new_[11516]_  = ~\new_[13211]_  & ~\new_[12333]_ ;
  assign \new_[11517]_  = ~\new_[11818]_ ;
  assign \new_[11518]_  = ~\new_[11819]_ ;
  assign \new_[11519]_  = ~\new_[12224]_  & ~\new_[12365]_ ;
  assign \new_[11520]_  = ~\dma_ack_i[3]  & (~\new_[12833]_  | ~n9140);
  assign \new_[11521]_  = ~\dma_ack_i[1]  & (~\new_[12649]_  | ~n9150);
  assign \new_[11522]_  = ~\new_[7206]_  | ~\new_[12540]_  | ~\new_[12684]_ ;
  assign \new_[11523]_  = ~\new_[12201]_ ;
  assign \new_[11524]_  = ~\new_[12322]_  | ~\new_[12468]_ ;
  assign \new_[11525]_  = ~\new_[12156]_ ;
  assign \new_[11526]_  = ~\new_[12394]_  | ~\new_[12248]_ ;
  assign \new_[11527]_  = ~\dma_ack_i[0]  & (~\new_[12653]_  | ~n9170);
  assign \new_[11528]_  = \new_[12320]_  | \new_[12425]_ ;
  assign \new_[11529]_  = ~\new_[12248]_  & ~\new_[12313]_ ;
  assign \new_[11530]_  = \new_[12394]_  | \new_[12313]_ ;
  assign \new_[11531]_  = ~\new_[12400]_  & ~\new_[12484]_ ;
  assign \new_[11532]_  = ~\new_[12468]_  & ~\new_[12411]_ ;
  assign \new_[11533]_  = \new_[12233]_  | \new_[12351]_ ;
  assign \new_[11534]_  = ~\dma_ack_i[2]  & (~\new_[12790]_  | ~n9215);
  assign \new_[11535]_  = ~\new_[12697]_  | (~\new_[12725]_  & ~\new_[12873]_ );
  assign \new_[11536]_  = ~\new_[12850]_  | (~\new_[13294]_  & ~\new_[12703]_ );
  assign \new_[11537]_  = ~\new_[12550]_  | (~\new_[13304]_  & ~\new_[12547]_ );
  assign \new_[11538]_  = ~\new_[13400]_  & (~\new_[12702]_  | ~\new_[13254]_ );
  assign \new_[11539]_  = ~\new_[13321]_  & (~\new_[12707]_  | ~\new_[13399]_ );
  assign \new_[11540]_  = ~\new_[12793]_  | (~\new_[12535]_  & ~\new_[12786]_ );
  assign \new_[11541]_  = ~\new_[12535]_  | (~\new_[12687]_  & ~\new_[12667]_ );
  assign \new_[11542]_  = ~\new_[12699]_  | (~\new_[13280]_  & ~\new_[12847]_ );
  assign \new_[11543]_  = ~\new_[12725]_  | (~\new_[13335]_  & ~\new_[12851]_ );
  assign \new_[11544]_  = ~\new_[13308]_  & (~\new_[12538]_  | ~\new_[12989]_ );
  assign \new_[11545]_  = ~\new_[13380]_  & (~\new_[12789]_  | ~\new_[13488]_ );
  assign \new_[11546]_  = ~\new_[13227]_  | (~\new_[12516]_  & ~\new_[12576]_ );
  assign \new_[11547]_  = ~\new_[13304]_  | (~\new_[12758]_  & ~\new_[13360]_ );
  assign \new_[11548]_  = ~\new_[12758]_  | (~\new_[13334]_  & ~\new_[12686]_ );
  assign \new_[11549]_  = ~\new_[12687]_  | (~\new_[13479]_  & ~\new_[12608]_ );
  assign \new_[11550]_  = ~\new_[13280]_  | (~\new_[12850]_  & ~\new_[13342]_ );
  assign \new_[11551]_  = ~\new_[12132]_ ;
  assign \new_[11552]_  = ~\new_[11842]_ ;
  assign \new_[11553]_  = ~\new_[12926]_  | (~\new_[12672]_  & ~\new_[12604]_ );
  assign \new_[11554]_  = ~\new_[13235]_  | (~\new_[12598]_  & ~\new_[12564]_ );
  assign \new_[11555]_  = ~\new_[12905]_  & (~\new_[12823]_  | ~\new_[13245]_ );
  assign \new_[11556]_  = ~\new_[11850]_ ;
  assign \new_[11557]_  = ~\new_[12357]_  & ~\new_[6102]_ ;
  assign \new_[11558]_  = ~\new_[11858]_ ;
  assign \new_[11559]_  = ~\new_[13041]_  & (~\new_[12853]_  | ~\new_[13064]_ );
  assign \new_[11560]_  = ~\new_[13127]_  & (~\new_[12623]_  | ~\new_[12997]_ );
  assign \new_[11561]_  = ~\new_[13008]_  & (~\new_[12936]_  | ~\new_[12544]_ );
  assign \new_[11562]_  = ~\new_[11863]_ ;
  assign \new_[11563]_  = ~\new_[11864]_ ;
  assign \new_[11564]_  = ~\new_[12314]_  | ~\new_[13024]_ ;
  assign \new_[11565]_  = ~\new_[12945]_  | (~\new_[12939]_  & ~\new_[12749]_ );
  assign \new_[11566]_  = ~\new_[11866]_ ;
  assign \new_[11567]_  = ~\new_[11822]_ ;
  assign \new_[11568]_  = ~\new_[12308]_  | ~\new_[13168]_ ;
  assign \new_[11569]_  = ~\new_[12819]_  & (~\new_[13077]_  | ~\new_[12613]_ );
  assign \new_[11570]_  = ~\new_[12977]_  | (~\new_[13052]_  & ~\new_[12739]_ );
  assign \new_[11571]_  = ~\new_[12943]_  & (~\new_[12726]_  | ~\new_[13097]_ );
  assign \new_[11572]_  = ~\new_[12386]_  & ~\dma_ack_i[3] ;
  assign \new_[11573]_  = ~\new_[14664]_ ;
  assign \new_[11574]_  = ~\new_[6367]_  & ~\new_[12981]_ ;
  assign \new_[11575]_  = ~\new_[13556]_  | ~\new_[13162]_ ;
  assign \new_[11576]_  = \new_[13433]_  ^ \new_[13446]_ ;
  assign \new_[11577]_  = ~\\u1_u3_idin_reg[31] ;
  assign \new_[11578]_  = ~\new_[12426]_  & ~\new_[6320]_ ;
  assign \new_[11579]_  = ~\new_[13223]_  & ~\new_[6322]_ ;
  assign \new_[11580]_  = ~\new_[6562]_  & ~\new_[12430]_ ;
  assign \new_[11581]_  = ~\new_[6343]_  & ~\new_[13160]_ ;
  assign \new_[11582]_  = ~\new_[12700]_  | ~\new_[13920]_ ;
  assign \new_[11583]_  = ~\new_[11855]_ ;
  assign \new_[11584]_  = ~\new_[6237]_  & ~\new_[12371]_ ;
  assign \new_[11585]_  = ~\new_[11821]_ ;
  assign \new_[11586]_  = ~\new_[13386]_  & ~\new_[12967]_ ;
  assign \new_[11587]_  = ~\new_[12450]_  | ~\wb_addr_i[4] ;
  assign \new_[11588]_  = ~\new_[12414]_  & ~\new_[13205]_ ;
  assign \new_[11589]_  = ~\new_[11756]_ ;
  assign \new_[11590]_  = ~\new_[12177]_ ;
  assign \new_[11591]_  = ~\new_[12420]_  | ~\new_[13464]_ ;
  assign \new_[11592]_  = ~n8995 & ~\new_[12348]_ ;
  assign \new_[11593]_  = \new_[12357]_  & \new_[12690]_ ;
  assign \new_[11594]_  = \new_[12352]_  & \new_[13285]_ ;
  assign \new_[11595]_  = ~\new_[12398]_  & ~\new_[12474]_ ;
  assign \new_[11596]_  = ~\new_[12191]_ ;
  assign \new_[11597]_  = ~\new_[12711]_  | ~\new_[12374]_ ;
  assign \new_[11598]_  = ~\new_[12797]_  | ~\new_[13257]_ ;
  assign \new_[11599]_  = ~\new_[12353]_  | ~\new_[13645]_ ;
  assign \new_[11600]_  = \new_[12455]_  & \new_[13463]_ ;
  assign \new_[11601]_  = ~\new_[11937]_ ;
  assign \new_[11602]_  = \new_[13434]_  & \new_[14582]_ ;
  assign \new_[11603]_  = ~\new_[12420]_  | ~\new_[6235]_ ;
  assign \new_[11604]_  = ~\new_[12428]_  | ~\new_[13111]_ ;
  assign \new_[11605]_  = \new_[12263]_  | \new_[12856]_ ;
  assign \new_[11606]_  = ~\new_[12431]_  | ~\new_[13084]_ ;
  assign \new_[11607]_  = ~\new_[12550]_  | ~\new_[12379]_ ;
  assign \new_[11608]_  = ~\new_[12334]_  & ~\dma_ack_i[0] ;
  assign \new_[11609]_  = ~n8955 & ~\new_[12460]_ ;
  assign \new_[11610]_  = ~\new_[12697]_  | ~\new_[12378]_ ;
  assign \new_[11611]_  = \new_[12436]_  | \new_[12786]_ ;
  assign \new_[11612]_  = ~n8985 & ~\new_[12449]_ ;
  assign \new_[11613]_  = ~\new_[11957]_ ;
  assign \new_[11614]_  = ~\new_[12535]_  | ~\new_[12382]_ ;
  assign \new_[11615]_  = \new_[12370]_  & \new_[13325]_ ;
  assign \new_[11616]_  = ~\new_[12469]_  & ~\dma_ack_i[1] ;
  assign \new_[11617]_  = ~\new_[11747]_ ;
  assign \new_[11618]_  = ~\new_[11965]_ ;
  assign \new_[11619]_  = \new_[12440]_  & \new_[12612]_ ;
  assign \new_[11620]_  = ~\new_[11812]_ ;
  assign \new_[11621]_  = ~\new_[2611]_  & (~\new_[13930]_  | ~\new_[13494]_ );
  assign \new_[11622]_  = ~\new_[12189]_ ;
  assign \new_[11623]_  = ~\new_[12359]_  | ~\new_[13051]_ ;
  assign \new_[11624]_  = ~\new_[12788]_  & (~\new_[3340]_  | ~\new_[3339]_ );
  assign \new_[11625]_  = ~\new_[13246]_  & (~\new_[4161]_  | ~\new_[4290]_ );
  assign \new_[11626]_  = ~\new_[12126]_ ;
  assign \new_[11627]_  = ~\new_[12433]_  & ~\new_[14387]_ ;
  assign \new_[11628]_  = ~\new_[12612]_  | ~\new_[13109]_ ;
  assign \new_[11629]_  = \new_[12501]_  & \new_[12359]_ ;
  assign \new_[11630]_  = ~\new_[12294]_  | ~\new_[13196]_ ;
  assign \new_[11631]_  = \new_[13008]_  | \new_[13147]_ ;
  assign \new_[11632]_  = ~\new_[12723]_  & (~\new_[3713]_  | ~\new_[3718]_ );
  assign \new_[11633]_  = ~\new_[12376]_  & (~\new_[3508]_  | ~\new_[3507]_ );
  assign \new_[11634]_  = \new_[12906]_  & \new_[12359]_ ;
  assign \new_[11635]_  = \new_[13206]_  & \new_[12272]_ ;
  assign \new_[11636]_  = ~\new_[12582]_  & (~\new_[4096]_  | ~\new_[4098]_ );
  assign \new_[11637]_  = ~\new_[12017]_ ;
  assign \new_[11638]_  = \new_[12618]_  & \new_[12294]_ ;
  assign \new_[11639]_  = \new_[13046]_  & \new_[12294]_ ;
  assign \new_[11640]_  = ~\new_[11760]_ ;
  assign n8620 = ~\new_[12959]_  | (~n9010 & ~\new_[3339]_ );
  assign \new_[11642]_  = ~\new_[12228]_  & (~\new_[3691]_  | ~\new_[13584]_ );
  assign \new_[11643]_  = \new_[13298]_  ^ \new_[14167]_ ;
  assign \new_[11644]_  = \new_[2984]_  ^ \new_[6017]_ ;
  assign \new_[11645]_  = \new_[2925]_  ^ \new_[6018]_ ;
  assign n8615 = ~\new_[12995]_  | (~n9015 & ~\new_[3718]_ );
  assign \new_[11647]_  = \new_[2870]_  ^ \new_[4615]_ ;
  assign \new_[11648]_  = ~\new_[12265]_  & (~\new_[6716]_  | ~\new_[6262]_ );
  assign \new_[11649]_  = ~\new_[4387]_  | ~\new_[13901]_  | ~\new_[14031]_  | ~\new_[5492]_ ;
  assign \new_[11650]_  = (~\new_[13788]_  | ~\new_[3888]_ ) & (~\new_[13989]_  | ~\new_[3889]_ );
  assign \new_[11651]_  = ~u0_u0_drive_k_reg;
  assign \new_[11652]_  = (~\new_[14001]_  | ~\new_[3315]_ ) & (~\new_[13264]_  | ~\new_[3316]_ );
  assign \new_[11653]_  = (~\new_[13926]_  | ~\new_[3690]_ ) & (~\new_[13440]_  | ~\new_[3693]_ );
  assign \new_[11654]_  = (~\new_[13962]_  | ~\new_[4293]_ ) & (~\new_[13747]_  | ~\new_[4206]_ );
  assign \new_[11655]_  = (~\new_[13649]_  | ~\new_[4070]_ ) & (~\new_[13372]_  | ~\new_[4073]_ );
  assign n8630 = RxActive_pad_i & rst_i;
  assign \new_[11657]_  = \new_[6242]_  ^ \new_[6018]_ ;
  assign \new_[11658]_  = ~\new_[11892]_ ;
  assign \new_[11659]_  = ~\new_[2873]_  | ~\new_[13895]_ ;
  assign \new_[11660]_  = ~\new_[12147]_ ;
  assign \new_[11661]_  = ~\new_[6292]_  & ~\new_[6718]_ ;
  assign \new_[11662]_  = ~n9145 | ~\new_[2871]_ ;
  assign \new_[11663]_  = ~\new_[12073]_ ;
  assign \new_[11664]_  = ~\new_[6526]_  & ~\new_[6696]_ ;
  assign \new_[11665]_  = ~\new_[12135]_ ;
  assign \new_[11666]_  = ~\new_[11811]_ ;
  assign n8635 = RxError_pad_i & rst_i;
  assign \new_[11668]_  = \new_[6690]_  | \new_[6200]_ ;
  assign \new_[11669]_  = ~\new_[12182]_ ;
  assign n8640 = RxValid_pad_i & rst_i;
  assign \new_[11671]_  = ~\new_[12172]_ ;
  assign \new_[11672]_  = ~\new_[14237]_  | ~\new_[13162]_ ;
  assign \new_[11673]_  = ~\new_[6291]_  & ~\new_[12396]_ ;
  assign \new_[11674]_  = ~\new_[13298]_  & ~\new_[13257]_ ;
  assign \new_[11675]_  = ~n9145 | ~\new_[2872]_ ;
  assign \new_[11676]_  = ~\new_[2673]_  | ~\new_[13858]_ ;
  assign \new_[11677]_  = ~\new_[4798]_  & ~\new_[4800]_ ;
  assign \new_[11678]_  = ~\new_[6599]_  & ~\new_[12375]_ ;
  assign \new_[11679]_  = ~\new_[14152]_  | ~\new_[13162]_ ;
  assign \new_[11680]_  = \new_[12426]_  & \new_[13350]_ ;
  assign \new_[11681]_  = ~\new_[12206]_ ;
  assign \new_[11682]_  = (~\new_[14139]_  | ~\new_[3479]_ ) & (~\new_[13364]_  | ~\new_[3481]_ );
  assign \new_[11683]_  = ~\new_[13392]_  & ~\new_[12439]_ ;
  assign \new_[11684]_  = ~\new_[12758]_  | ~\new_[12370]_ ;
  assign \new_[11685]_  = \new_[6387]_  ^ \new_[13496]_ ;
  assign \new_[11686]_  = ~u0_u0_ls_j_r_reg;
  assign \new_[11687]_  = ~u1_u2_mwe_reg;
  assign \new_[11688]_  = ~\new_[12414]_  & ~\new_[13257]_ ;
  assign \new_[11689]_  = \new_[12482]_  & \new_[13381]_ ;
  assign \new_[11690]_  = \new_[12644]_  ^ \new_[12596]_ ;
  assign \new_[11691]_  = \new_[6809]_  | \new_[6009]_ ;
  assign \new_[11692]_  = ~\new_[2871]_  | ~\new_[14790]_ ;
  assign \new_[11693]_  = (~\new_[2929]_  | ~\new_[12671]_ ) & (~\new_[12519]_  | ~\new_[5109]_ );
  assign \new_[11694]_  = \new_[12322]_  | \new_[12411]_ ;
  assign \new_[11695]_  = ~\new_[12185]_ ;
  assign \new_[11696]_  = ~\new_[12774]_  | ~\new_[12429]_ ;
  assign \new_[11697]_  = ~n8340;
  assign \new_[11698]_  = u0_u0_chirp_cnt_is_6_reg;
  assign \new_[11699]_  = \new_[6107]_  ^ \new_[6017]_ ;
  assign \new_[11700]_  = \new_[3410]_  ^ \new_[12900]_ ;
  assign \new_[11701]_  = ~\new_[12746]_  | (~\new_[12697]_  & ~\new_[12856]_ );
  assign \new_[11702]_  = ~\new_[12717]_  | ~\new_[12342]_ ;
  assign \new_[11703]_  = \new_[12886]_  ^ \new_[12527]_ ;
  assign \new_[11704]_  = ~\new_[14003]_  | ~\new_[13870]_  | ~\new_[12229]_  | ~\new_[13416]_ ;
  assign \new_[11705]_  = \new_[13407]_  & \new_[13598]_ ;
  assign \new_[11706]_  = \new_[12257]_  | \new_[12847]_ ;
  assign \new_[11707]_  = ~\new_[12384]_  & ~\new_[12704]_ ;
  assign \new_[11708]_  = ~\new_[13521]_  | ~\new_[13162]_ ;
  assign \new_[11709]_  = ~\new_[11824]_ ;
  assign \new_[11710]_  = \new_[12894]_  ^ \new_[12689]_ ;
  assign \new_[11711]_  = ~\new_[12056]_ ;
  assign \new_[11712]_  = ~\new_[12227]_  & ~\new_[13978]_ ;
  assign \new_[11713]_  = ~\new_[12229]_  | ~\new_[13409]_ ;
  assign \new_[11714]_  = ~\new_[13057]_  | ~\new_[12338]_ ;
  assign \new_[11715]_  = ~\new_[3174]_  | ~\new_[13895]_ ;
  assign \new_[11716]_  = ~\new_[12366]_  | ~\new_[12408]_ ;
  assign n8650 = ~\new_[13119]_  | (~n8890 & ~\new_[3507]_ );
  assign \new_[11718]_  = ~\new_[13908]_  | ~\new_[14003]_  | ~\new_[12229]_  | ~\new_[13409]_ ;
  assign \new_[11719]_  = ~\new_[12850]_  | ~\new_[12352]_ ;
  assign \new_[11720]_  = \new_[2988]_  ^ \new_[12890]_ ;
  assign \new_[11721]_  = ~\new_[14386]_ ;
  assign \new_[11722]_  = ~\new_[13121]_  | ~\new_[12898]_  | ~\new_[3037]_ ;
  assign \new_[11723]_  = ~\new_[11926]_ ;
  assign \new_[11724]_  = \new_[13870]_  | \new_[3063]_  | \new_[12240]_  | \new_[14003]_ ;
  assign \new_[11725]_  = ~\new_[12163]_ ;
  assign n8610 = ~\new_[13142]_  | (~n9020 & ~\new_[4098]_ );
  assign \new_[11727]_  = u1_hms_clk_reg;
  assign \new_[11728]_  = ~\new_[12413]_  & ~\dma_ack_i[2] ;
  assign \new_[11729]_  = ~\new_[6200]_  & ~\new_[13365]_ ;
  assign \new_[11730]_  = ~\new_[14678]_ ;
  assign \new_[11731]_  = ~\new_[3025]_  | (~\new_[12965]_  & ~\new_[14089]_ );
  assign \new_[11732]_  = ~\new_[12317]_ ;
  assign \new_[11733]_  = ~\\u1_u3_idin_reg[28] ;
  assign \new_[11734]_  = ~\new_[13182]_  | (~\new_[6250]_  & ~\new_[13393]_ );
  assign \new_[11735]_  = ~\new_[13225]_  & (~\new_[13182]_  | ~\new_[13059]_ );
  assign \new_[11736]_  = ~\new_[12818]_  & (~\new_[3480]_  | ~\new_[14149]_ );
  assign \new_[11737]_  = ~\new_[13411]_  & ~\new_[12637]_ ;
  assign \new_[11738]_  = ~\new_[13014]_  & (~\new_[13074]_  | ~\new_[13086]_ );
  assign \new_[11739]_  = ~\new_[12979]_  & (~\new_[13142]_  | ~\new_[13004]_ );
  assign \new_[11740]_  = ~\new_[12910]_  & (~\new_[13006]_  | ~\new_[13233]_ );
  assign \new_[11741]_  = ~\new_[12944]_  & (~\new_[13057]_  | ~\new_[12918]_ );
  assign \new_[11742]_  = ~\new_[12845]_  & (~\new_[6280]_  | ~\new_[6716]_ );
  assign \new_[11743]_  = ~\new_[13015]_  & (~\new_[13119]_  | ~\new_[13025]_ );
  assign \new_[11744]_  = ~\new_[13053]_  & (~\new_[12959]_  | ~\new_[12992]_ );
  assign \new_[11745]_  = \new_[13486]_  & \new_[12701]_ ;
  assign \new_[11746]_  = ~\new_[12663]_  | ~\new_[3888]_ ;
  assign \new_[11747]_  = ~\new_[12704]_  & ~\new_[12674]_ ;
  assign \new_[11748]_  = ~\new_[13316]_  | ~\new_[9412]_  | ~\new_[13495]_  | ~\new_[9405]_ ;
  assign \new_[11749]_  = ~\new_[13383]_  | ~\new_[8701]_  | ~\new_[13356]_  | ~\new_[8826]_ ;
  assign n8665 = \sram_data_i[31]  ? \new_[13178]_  : \new_[11018]_ ;
  assign \new_[11751]_  = \new_[2092]_  ^ \new_[12973]_ ;
  assign \new_[11752]_  = ~\new_[13160]_  | ~\new_[12641]_  | ~\new_[13417]_ ;
  assign \new_[11753]_  = ~\new_[12390]_ ;
  assign \new_[11754]_  = ~\new_[12665]_  | ~\new_[12525]_ ;
  assign \new_[11755]_  = ~\new_[12979]_  & ~\new_[12597]_ ;
  assign \new_[11756]_  = ~\new_[12704]_  & ~\new_[12553]_ ;
  assign \new_[11757]_  = ~\new_[13360]_  & ~\new_[12547]_ ;
  assign \new_[11758]_  = \\u0_u0_idle_cnt1_next_reg[1] ;
  assign \new_[11759]_  = ~\new_[12765]_  & (~\new_[4286]_  | ~\new_[13754]_ );
  assign \new_[11760]_  = ~\new_[12724]_  & (~\new_[6716]_  | ~\new_[6020]_ );
  assign \new_[11761]_  = \new_[12890]_  & \new_[2988]_ ;
  assign \new_[11762]_  = ~\new_[12720]_  | ~\new_[13747]_ ;
  assign \new_[11763]_  = \new_[12582]_  | \new_[13421]_ ;
  assign \new_[11764]_  = ~\new_[12670]_  | ~\new_[12968]_ ;
  assign \new_[11765]_  = ~\new_[12723]_  | ~\new_[13271]_ ;
  assign \new_[11766]_  = \new_[12788]_  | \new_[13497]_ ;
  assign \new_[11767]_  = ~\new_[12623]_  & ~\new_[12739]_ ;
  assign \new_[11768]_  = ~\new_[12722]_  | ~\new_[13989]_ ;
  assign \new_[11769]_  = \new_[12740]_  | \new_[3509]_ ;
  assign \new_[11770]_  = \new_[12723]_  | \new_[13271]_ ;
  assign \new_[11771]_  = \new_[12800]_  & \new_[13850]_ ;
  assign n8730 = \sram_data_i[5]  ? \new_[13178]_  : \new_[11349]_ ;
  assign \new_[11773]_  = ~\new_[12886]_  | ~\new_[13325]_ ;
  assign \new_[11774]_  = ~\new_[12899]_  | ~\new_[13144]_ ;
  assign \new_[11775]_  = ~\new_[13385]_  | ~\new_[13937]_  | ~\new_[12609]_  | ~\new_[13339]_ ;
  assign \new_[11776]_  = ~\new_[12910]_  & ~\new_[12863]_ ;
  assign \new_[11777]_  = ~\new_[13053]_  & ~\new_[12577]_ ;
  assign \new_[11778]_  = ~\new_[12237]_ ;
  assign \new_[11779]_  = \new_[13246]_  & \new_[12684]_ ;
  assign \new_[11780]_  = ~\new_[12547]_  & ~\new_[12983]_ ;
  assign \new_[11781]_  = ~\new_[13457]_  | ~\new_[13389]_  | ~\new_[12540]_  | ~\new_[13137]_ ;
  assign n8825 = ~\new_[13181]_  & ~\new_[12733]_ ;
  assign \new_[11783]_  = ~\new_[13004]_  | ~\new_[13142]_  | ~\new_[12968]_ ;
  assign \new_[11784]_  = ~\new_[13025]_  | ~\new_[13119]_  | ~\new_[13141]_ ;
  assign \new_[11785]_  = ~\new_[12815]_  | ~\new_[13141]_ ;
  assign \new_[11786]_  = ~\new_[2989]_  | ~\new_[12890]_  | ~\new_[2988]_ ;
  assign \new_[11787]_  = \new_[13026]_  ^ \new_[13186]_ ;
  assign \new_[11788]_  = \new_[13061]_  ^ \new_[13226]_ ;
  assign \new_[11789]_  = \new_[4511]_  ^ \new_[13230]_ ;
  assign \new_[11790]_  = \new_[14308]_  ^ \new_[14571]_ ;
  assign \new_[11791]_  = ~\new_[13416]_  | ~\new_[12735]_  | ~\new_[14163]_ ;
  assign \new_[11792]_  = u0_u0_ls_k_r_reg;
  assign \new_[11793]_  = ~\new_[12637]_  & ~\new_[14096]_ ;
  assign \new_[11794]_  = ~\new_[3470]_  | ~\new_[12671]_ ;
  assign \new_[11795]_  = ~\new_[3465]_  | ~\new_[12671]_ ;
  assign \new_[11796]_  = ~\new_[3472]_  | ~\new_[12671]_ ;
  assign \new_[11797]_  = ~\new_[13167]_ ;
  assign \new_[11798]_  = \new_[12580]_  & \new_[2477]_ ;
  assign \new_[11799]_  = ~\new_[13382]_  | ~\new_[12857]_ ;
  assign \new_[11800]_  = ~\new_[13366]_  | ~\new_[12551]_ ;
  assign \new_[11801]_  = \new_[4873]_  | \new_[12586]_ ;
  assign \new_[11802]_  = ~\new_[13215]_  & ~\new_[12748]_ ;
  assign \new_[11803]_  = ~\new_[13300]_  | ~\new_[12563]_ ;
  assign \new_[11804]_  = ~wb_we_i | ~\new_[12626]_ ;
  assign \new_[11805]_  = \new_[12609]_  & \new_[13532]_ ;
  assign \new_[11806]_  = ~\new_[13237]_  | ~\new_[12647]_  | ~\new_[13326]_ ;
  assign \new_[11807]_  = ~\new_[12721]_  | ~\new_[13097]_ ;
  assign \new_[11808]_  = ~\new_[13473]_  | ~\new_[12620]_ ;
  assign \new_[11809]_  = ~\new_[13134]_  | ~\new_[12567]_  | ~\new_[13289]_ ;
  assign \new_[11810]_  = \new_[4508]_  | \new_[4507]_  | \new_[12770]_  | \new_[13314]_ ;
  assign \new_[11811]_  = ~\new_[4791]_  | ~\new_[12883]_ ;
  assign \new_[11812]_  = \new_[12731]_  | \new_[12604]_ ;
  assign \new_[11813]_  = ~\new_[12538]_  & ~\new_[13307]_ ;
  assign \new_[11814]_  = ~\new_[13459]_  | ~\new_[12615]_ ;
  assign \new_[11815]_  = ~\new_[12981]_  | ~\new_[12642]_  | ~\new_[13363]_ ;
  assign \new_[11816]_  = ~\new_[12619]_  & ~\new_[12548]_ ;
  assign \new_[11817]_  = ~\new_[12558]_  | ~\new_[12776]_ ;
  assign \new_[11818]_  = ~\new_[13850]_  | ~\new_[13320]_  | ~\new_[13419]_  | ~\new_[13657]_ ;
  assign \new_[11819]_  = ~\new_[6346]_  & (~\new_[13355]_  | ~\new_[13010]_ );
  assign \new_[11820]_  = ~\new_[12834]_  | ~\new_[13913]_ ;
  assign \new_[11821]_  = ~\new_[12560]_  | ~\new_[13588]_ ;
  assign \new_[11822]_  = ~\new_[13019]_  & (~\new_[12998]_  | ~\new_[13000]_ );
  assign \new_[11823]_  = ~\new_[12483]_ ;
  assign \new_[11824]_  = ~\new_[6588]_  & (~\new_[13413]_  | ~\new_[13242]_ );
  assign \new_[11825]_  = ~\new_[12823]_  & ~\new_[12564]_ ;
  assign \new_[11826]_  = ~\new_[13491]_  | (~\new_[13073]_  & ~\new_[13270]_ );
  assign \new_[11827]_  = ~\new_[13003]_  | (~\new_[13184]_  & ~\new_[13277]_ );
  assign \new_[11828]_  = ~\new_[13384]_  | (~\new_[13003]_  & ~\new_[13260]_ );
  assign \new_[11829]_  = ~\new_[13130]_  | (~\new_[13152]_  & ~\new_[13444]_ );
  assign \new_[11830]_  = ~\new_[13259]_  | (~\new_[13130]_  & ~\new_[13275]_ );
  assign \new_[11831]_  = ~\new_[13216]_  | (~\new_[13179]_  & ~\new_[13480]_ );
  assign \new_[11832]_  = ~\new_[13306]_  | (~\new_[13216]_  & ~\new_[13274]_ );
  assign \new_[11833]_  = ~\new_[13202]_  & (~\new_[12940]_  | ~\new_[13088]_ );
  assign \new_[11834]_  = ~\new_[12936]_  & (~\new_[13005]_  | ~\new_[13103]_ );
  assign \new_[11835]_  = ~\new_[12590]_  & (~\new_[3879]_  | ~\new_[13337]_ );
  assign \new_[11836]_  = ~\new_[13028]_  & (~\new_[13041]_  | ~\new_[13106]_ );
  assign \new_[11837]_  = \new_[12657]_  & \new_[13088]_ ;
  assign \new_[11838]_  = ~\new_[13107]_  & (~\new_[13127]_  | ~\new_[13009]_ );
  assign \new_[11839]_  = ~\new_[13208]_  & (~\new_[13225]_  | ~\new_[13090]_ );
  assign \new_[11840]_  = ~\new_[12998]_  & (~\new_[13173]_  | ~\new_[13131]_ );
  assign \new_[11841]_  = ~\new_[12937]_  & (~\new_[13019]_  | ~\new_[12946]_ );
  assign \new_[11842]_  = ~\new_[12980]_  & (~\new_[12902]_  | ~\new_[13039]_ );
  assign \new_[11843]_  = ~u4_suspend_r1_reg;
  assign \new_[11844]_  = ~\new_[12996]_  & (~\new_[13049]_  | ~\new_[12935]_ );
  assign \new_[11845]_  = ~\new_[13049]_  & (~\new_[12910]_  | ~\new_[13076]_ );
  assign \new_[11846]_  = ~\new_[13161]_  & (~\new_[13253]_  | ~\new_[12969]_ );
  assign \new_[11847]_  = ~\new_[12513]_  & (~\new_[3592]_  | ~\new_[13256]_ );
  assign \new_[11848]_  = ~\new_[13045]_  & (~\new_[13104]_  | ~\new_[13066]_ );
  assign \new_[11849]_  = ~\new_[13145]_  & (~\new_[12986]_  | ~\new_[12904]_ );
  assign \new_[11850]_  = ~\new_[13104]_  & (~\new_[13053]_  | ~\new_[13105]_ );
  assign \new_[11851]_  = ~\new_[13180]_  & (~\new_[13145]_  | ~\new_[13063]_ );
  assign \new_[11852]_  = ~\new_[13056]_  & (~\new_[12954]_  | ~\new_[13194]_ );
  assign \new_[11853]_  = ~\new_[12607]_  & (~\new_[3462]_  | ~\new_[13272]_ );
  assign \new_[11854]_  = ~\new_[12616]_  & (~\new_[3466]_  | ~\new_[13301]_ );
  assign \new_[11855]_  = ~\new_[12496]_  | ~\new_[14108]_ ;
  assign \new_[11856]_  = ~\new_[13033]_  & (~\new_[12925]_  | ~\new_[13249]_ );
  assign \new_[11857]_  = ~\new_[12925]_  & (~\new_[12937]_  | ~\new_[13034]_ );
  assign \new_[11858]_  = ~\new_[13173]_  & (~\new_[12979]_  | ~\new_[12968]_ );
  assign \new_[11859]_  = ~\new_[13239]_  & (~\new_[13208]_  | ~\new_[12990]_ );
  assign \new_[11860]_  = ~\new_[13093]_  & (~\new_[12944]_  | ~\new_[13213]_ );
  assign \new_[11861]_  = ~\new_[13199]_  & (~\new_[13177]_  | ~\new_[12909]_ );
  assign \new_[11862]_  = ~\new_[13005]_  & (~\new_[13048]_  | ~\new_[12912]_ );
  assign \new_[11863]_  = ~\new_[13177]_  & (~\new_[13015]_  | ~\new_[13141]_ );
  assign \new_[11864]_  = ~\new_[13048]_  & (~\new_[13199]_  | ~\new_[13212]_ );
  assign \new_[11865]_  = ~\new_[12512]_  & (~\new_[3686]_  | ~\new_[13255]_ );
  assign \new_[11866]_  = ~\new_[12986]_  & (~\new_[13045]_  | ~\new_[12924]_ );
  assign \new_[11867]_  = ~\new_[12923]_  & (~\new_[13028]_  | ~\new_[13243]_ );
  assign \new_[11868]_  = ~\new_[12940]_  & (~\new_[13014]_  | ~\new_[13133]_ );
  assign \new_[11869]_  = ~\new_[13244]_  & (~\new_[13107]_  | ~\new_[13001]_ );
  assign \new_[11870]_  = ~\new_[12902]_  & (~\new_[13154]_  | ~\new_[13082]_ );
  assign \new_[11871]_  = ~\new_[13215]_  & (~\new_[12980]_  | ~\new_[13101]_ );
  assign \new_[11872]_  = ~\new_[12501]_  | ~\new_[13752]_ ;
  assign \new_[11873]_  = ~\new_[12673]_  | ~\new_[13506]_ ;
  assign \new_[11874]_  = ~\new_[6299]_  & ~\new_[13237]_ ;
  assign \new_[11875]_  = ~\new_[4666]_  | ~\new_[4780]_  | ~\new_[13140]_  | ~\new_[4779]_ ;
  assign \new_[11876]_  = ~\new_[12430]_ ;
  assign \new_[11877]_  = ~\new_[13128]_  | ~\new_[12551]_ ;
  assign \new_[11878]_  = ~\new_[12884]_  | ~\new_[13463]_ ;
  assign \new_[11879]_  = ~\new_[13460]_  & ~\new_[4796]_ ;
  assign \new_[11880]_  = ~\new_[13615]_  & ~\new_[12575]_ ;
  assign \new_[11881]_  = ~\new_[6266]_  & ~\new_[13221]_ ;
  assign n8805 = \sram_data_i[25]  ? \new_[13178]_  : \new_[11390]_ ;
  assign \new_[11883]_  = ~\new_[12529]_  & ~\new_[13150]_ ;
  assign n8820 = \sram_data_i[11]  ? \new_[13178]_  : \new_[11399]_ ;
  assign n8790 = \sram_data_i[7]  ? \new_[13178]_  : \new_[11384]_ ;
  assign n8765 = \sram_data_i[9]  ? \new_[13178]_  : \new_[11378]_ ;
  assign n8725 = \sram_data_i[3]  ? \new_[13178]_  : \new_[11346]_ ;
  assign n8750 = \sram_data_i[0]  ? \new_[13178]_  : \new_[11363]_ ;
  assign n8810 = \sram_data_i[12]  ? \new_[13178]_  : \new_[11391]_ ;
  assign n8710 = \sram_data_i[4]  ? \new_[13178]_  : \new_[11218]_ ;
  assign n8780 = \sram_data_i[16]  ? \new_[13178]_  : \new_[11382]_ ;
  assign \new_[11892]_  = ~\new_[13930]_  & ~\new_[2611]_ ;
  assign n8705 = \sram_data_i[10]  ? \new_[13178]_  : \new_[11217]_ ;
  assign n8770 = \sram_data_i[21]  ? \new_[13178]_  : \new_[11380]_ ;
  assign n8700 = \sram_data_i[18]  ? \new_[13178]_  : \new_[11216]_ ;
  assign n8720 = \sram_data_i[27]  ? \new_[13178]_  : \new_[11334]_ ;
  assign n8755 = \sram_data_i[1]  ? \new_[13178]_  : \new_[11364]_ ;
  assign n8715 = \sram_data_i[30]  ? \new_[13178]_  : \new_[11327]_ ;
  assign n8660 = \sram_data_i[2]  ? \new_[13178]_  : \new_[11016]_ ;
  assign \new_[11900]_  = \new_[4780]_  | \new_[4774]_  | \new_[4779]_  | \new_[4666]_ ;
  assign n8760 = \sram_data_i[29]  ? \new_[13178]_  : \new_[11365]_ ;
  assign n8680 = \sram_data_i[23]  ? \new_[13178]_  : \new_[11057]_ ;
  assign n8775 = \sram_data_i[20]  ? \new_[13178]_  : \new_[11381]_ ;
  assign n8675 = \sram_data_i[6]  ? \new_[13178]_  : \new_[11030]_ ;
  assign n8695 = \sram_data_i[24]  ? \new_[13178]_  : \new_[11215]_ ;
  assign \new_[11906]_  = ~\new_[12742]_  & (~\new_[13093]_  | ~\new_[13023]_ );
  assign \new_[11907]_  = ~\new_[13741]_  & ~\new_[12877]_ ;
  assign \new_[11908]_  = \new_[13749]_  ^ \new_[13085]_ ;
  assign \new_[11909]_  = \new_[4370]_  ^ \new_[13166]_ ;
  assign \new_[11910]_  = \new_[13453]_  ^ \new_[13328]_ ;
  assign \new_[11911]_  = ~\new_[12262]_ ;
  assign \new_[11912]_  = ~\new_[13073]_  | (~\new_[13113]_  & ~\new_[13291]_ );
  assign \new_[11913]_  = ~\new_[13272]_  | ~\new_[13718]_ ;
  assign \new_[11914]_  = ~\new_[13198]_  & ~\new_[6370]_ ;
  assign \new_[11915]_  = ~\new_[12498]_  & ~\new_[14089]_ ;
  assign \new_[11916]_  = ~\new_[13261]_  & ~\new_[2452]_ ;
  assign \new_[11917]_  = ~\new_[13533]_  & ~\new_[12859]_ ;
  assign \new_[11918]_  = ~\new_[13222]_  & ~\new_[6588]_ ;
  assign \new_[11919]_  = ~\new_[12509]_  | ~\new_[13368]_ ;
  assign \new_[11920]_  = ~\new_[12572]_  & ~\new_[13277]_ ;
  assign \new_[11921]_  = ~\new_[12851]_  & ~\new_[12873]_ ;
  assign \new_[11922]_  = ~\new_[12276]_ ;
  assign \new_[11923]_  = ~\new_[12588]_  & ~\new_[12437]_ ;
  assign \new_[11924]_  = ~\new_[12280]_ ;
  assign \new_[11925]_  = ~\new_[12712]_  | ~\new_[13904]_ ;
  assign \new_[11926]_  = \new_[12700]_  & \new_[12500]_ ;
  assign \new_[11927]_  = \new_[13283]_  & \new_[12695]_ ;
  assign \new_[11928]_  = ~\new_[13016]_  & (~\new_[12995]_  | ~\new_[13087]_ );
  assign \new_[11929]_  = ~\new_[12704]_  & ~\new_[12982]_ ;
  assign \new_[11930]_  = ~\new_[12283]_ ;
  assign \new_[11931]_  = ~\new_[13256]_  | ~\new_[13548]_ ;
  assign \new_[11932]_  = ~\new_[12618]_  | ~\new_[13981]_ ;
  assign \new_[11933]_  = ~\new_[13466]_  & ~\new_[12752]_ ;
  assign \new_[11934]_  = ~\new_[6319]_  & ~\new_[13350]_ ;
  assign n8340 = ~\new_[12553]_  & ~\new_[12824]_ ;
  assign \new_[11936]_  = \new_[12948]_  & \new_[12524]_ ;
  assign \new_[11937]_  = ~\new_[12786]_  & ~\new_[13387]_ ;
  assign \new_[11938]_  = ~\new_[13347]_  & ~\new_[4796]_ ;
  assign \new_[11939]_  = ~\new_[12608]_  & ~\new_[12667]_ ;
  assign \new_[11940]_  = ~\new_[13434]_  & ~\new_[4800]_ ;
  assign \new_[11941]_  = \new_[13365]_  & \new_[12525]_ ;
  assign \new_[11942]_  = \new_[12415]_  & \wb_addr_i[4] ;
  assign \new_[11943]_  = ~\new_[12550]_  & ~\new_[12983]_ ;
  assign \new_[11944]_  = \new_[13084]_  & \new_[13298]_ ;
  assign \new_[11945]_  = ~\new_[12707]_  & ~\new_[13126]_ ;
  assign \new_[11946]_  = ~\new_[4780]_  | ~\new_[13428]_ ;
  assign \new_[11947]_  = ~\new_[12702]_  & ~\new_[13387]_ ;
  assign \new_[11948]_  = ~\new_[6343]_  & ~\new_[12911]_ ;
  assign \new_[11949]_  = ~\new_[12523]_  | ~\new_[4293]_ ;
  assign \new_[11950]_  = \new_[13290]_  & \new_[12509]_ ;
  assign \new_[11951]_  = ~\new_[12878]_  & ~\new_[13291]_ ;
  assign \new_[11952]_  = ~\new_[13396]_  & ~\new_[13277]_ ;
  assign \new_[11953]_  = ~\new_[12701]_  | ~\new_[13358]_ ;
  assign \new_[11954]_  = \new_[12519]_  & \new_[5756]_ ;
  assign \new_[11955]_  = ~\new_[4794]_  & ~\new_[12778]_ ;
  assign \new_[11956]_  = ~\new_[12703]_  & ~\new_[13342]_ ;
  assign \new_[11957]_  = ~\new_[12541]_  | ~\new_[13431]_ ;
  assign \new_[11958]_  = \wb_addr_i[6]  | \wb_addr_i[7]  | \wb_addr_i[4]  | \wb_addr_i[8] ;
  assign \new_[11959]_  = ~\new_[12496]_  & ~\new_[13492]_ ;
  assign \new_[11960]_  = ~\new_[13308]_  & ~\new_[13482]_ ;
  assign \new_[11961]_  = ~\new_[12944]_  & ~\new_[12675]_ ;
  assign \new_[11962]_  = \new_[13310]_  & \new_[12787]_ ;
  assign \new_[11963]_  = ~\new_[12288]_ ;
  assign \new_[11964]_  = \new_[12528]_  | \new_[13461]_ ;
  assign \new_[11965]_  = ~\new_[12847]_  & ~\new_[13126]_ ;
  assign \new_[11966]_  = ~\new_[12365]_ ;
  assign \new_[11967]_  = \new_[12579]_  & \new_[13029]_ ;
  assign \new_[11968]_  = ~\new_[13015]_  & ~\new_[12669]_ ;
  assign \new_[11969]_  = ~\new_[12499]_  | ~\new_[13106]_ ;
  assign \new_[11970]_  = ~\new_[12534]_  | ~\new_[2097]_ ;
  assign \new_[11971]_  = ~\new_[12484]_ ;
  assign \new_[11972]_  = ~\new_[12772]_  | ~\new_[13009]_ ;
  assign \new_[11973]_  = ~n9130 & (~\new_[13570]_  | ~\new_[13135]_ );
  assign \new_[11974]_  = ~\new_[12719]_  & ~\new_[13157]_ ;
  assign \new_[11975]_  = ~\new_[13005]_  & ~\new_[12508]_ ;
  assign \new_[11976]_  = ~\new_[12472]_ ;
  assign \new_[11977]_  = ~\new_[13014]_  & ~\new_[12866]_ ;
  assign \new_[11978]_  = ~\new_[13199]_  & ~\new_[12546]_ ;
  assign \new_[11979]_  = ~\new_[12664]_  | ~\new_[13090]_ ;
  assign \new_[11980]_  = ~\new_[12660]_  | ~\new_[13064]_ ;
  assign \new_[11981]_  = ~\new_[13180]_  & ~\new_[12683]_ ;
  assign \new_[11982]_  = \new_[12814]_  & \new_[12935]_ ;
  assign \new_[11983]_  = ~\new_[12853]_  & ~\new_[12576]_ ;
  assign \new_[11984]_  = ~\new_[13102]_  & ~\new_[12731]_ ;
  assign \new_[11985]_  = ~\new_[12741]_  | ~\new_[13213]_ ;
  assign \new_[11986]_  = ~\new_[12937]_  & ~\new_[12854]_ ;
  assign \new_[11987]_  = ~\new_[12925]_  & ~\new_[12666]_ ;
  assign \new_[11988]_  = ~\new_[12708]_  & (~\new_[2339]_  | ~\new_[2342]_ );
  assign \new_[11989]_  = ~\new_[13016]_  & ~\new_[12826]_ ;
  assign \new_[11990]_  = \new_[12871]_  & \new_[12990]_ ;
  assign \new_[11991]_  = ~\new_[12425]_ ;
  assign \new_[11992]_  = ~\new_[13019]_  & ~\new_[12730]_ ;
  assign \new_[11993]_  = \new_[12657]_  & \new_[13052]_ ;
  assign \new_[11994]_  = ~\new_[12726]_  & ~\new_[12604]_ ;
  assign \new_[11995]_  = \new_[12814]_  & \new_[12598]_ ;
  assign \new_[11996]_  = ~\new_[12214]_ ;
  assign \new_[11997]_  = ~\new_[12407]_ ;
  assign \new_[11998]_  = ~\new_[12409]_ ;
  assign \new_[11999]_  = ~\new_[12841]_  & ~\new_[12533]_ ;
  assign \new_[12000]_  = ~\new_[12411]_ ;
  assign \new_[12001]_  = ~\new_[12986]_  & ~\new_[12844]_ ;
  assign \new_[12002]_  = ~\new_[12792]_  | ~\new_[12984]_ ;
  assign \new_[12003]_  = ~\new_[13225]_  & ~\new_[12677]_ ;
  assign \new_[12004]_  = ~\new_[12858]_  | ~\new_[13076]_ ;
  assign \new_[12005]_  = \new_[13052]_  & \new_[12685]_ ;
  assign \new_[12006]_  = ~\new_[12658]_  | ~\new_[13217]_ ;
  assign \new_[12007]_  = ~\new_[12659]_  | ~\new_[13249]_ ;
  assign \new_[12008]_  = ~\new_[12880]_  | ~\new_[13050]_ ;
  assign \new_[12009]_  = ~\new_[13078]_  & ~\new_[12504]_ ;
  assign \new_[12010]_  = ~\new_[12801]_  | ~\new_[13105]_ ;
  assign \new_[12011]_  = ~\new_[12318]_ ;
  assign \new_[12012]_  = ~\new_[13145]_  & ~\new_[12581]_ ;
  assign \new_[12013]_  = ~\new_[13045]_  & ~\new_[12662]_ ;
  assign \new_[12014]_  = ~\new_[12327]_ ;
  assign \new_[12015]_  = ~\new_[12234]_ ;
  assign \new_[12016]_  = ~\new_[12319]_ ;
  assign \new_[12017]_  = \new_[12685]_  | \new_[12739]_ ;
  assign \new_[12018]_  = ~\new_[12705]_  & ~\new_[12685]_ ;
  assign \new_[12019]_  = ~\new_[12230]_ ;
  assign \new_[12020]_  = ~\new_[12980]_  & ~\new_[12813]_ ;
  assign \new_[12021]_  = \new_[12598]_  & \new_[12938]_ ;
  assign \new_[12022]_  = ~\new_[12225]_ ;
  assign \new_[12023]_  = ~\new_[12517]_  | ~\new_[13133]_ ;
  assign \new_[12024]_  = ~\new_[12875]_  | ~\new_[13238]_ ;
  assign \new_[12025]_  = ~\new_[12936]_  & ~\new_[12737]_ ;
  assign \new_[12026]_  = ~\new_[12769]_  | ~\new_[12997]_ ;
  assign \new_[12027]_  = ~\new_[12241]_ ;
  assign \new_[12028]_  = ~\new_[12328]_ ;
  assign \new_[12029]_  = ~\new_[12868]_  | ~\new_[12738]_ ;
  assign \new_[12030]_  = ~\new_[12820]_  & (~\new_[4291]_  | ~\new_[13675]_ );
  assign \new_[12031]_  = ~\new_[12729]_  & (~\new_[3790]_  | ~\new_[13947]_ );
  assign \new_[12032]_  = ~\new_[13006]_  | (~\new_[5998]_  & ~\new_[13262]_ );
  assign \new_[12033]_  = ~\new_[6196]_  & ~\new_[6247]_ ;
  assign \new_[12034]_  = ~\new_[12601]_  & (~\new_[3884]_  | ~\new_[14197]_ );
  assign \new_[12035]_  = ~\new_[12522]_  & (~\new_[6268]_  | ~\new_[6716]_ );
  assign \new_[12036]_  = ~\new_[13057]_  | (~\new_[6003]_  & ~\new_[13422]_ );
  assign \new_[12037]_  = ~\new_[6718]_  & ~\new_[6109]_ ;
  assign \new_[12038]_  = ~\new_[12335]_ ;
  assign \new_[12039]_  = (~\new_[13371]_  | ~\new_[6365]_ ) & (~\new_[6366]_  | ~\new_[13865]_ );
  assign \new_[12040]_  = ~\new_[2476]_  & ~\new_[2392]_ ;
  assign \new_[12041]_  = ~\new_[3503]_  | ~\new_[3504]_ ;
  assign \new_[12042]_  = (~\new_[13262]_  | ~\new_[6484]_ ) & (~\new_[6168]_  | ~\new_[14045]_ );
  assign \new_[12043]_  = (~\new_[13897]_  | ~\new_[3711]_ ) & (~\new_[13905]_  | ~\new_[3788]_ );
  assign \new_[12044]_  = (~\new_[13422]_  | ~\new_[6341]_ ) & (~\new_[6592]_  | ~\new_[13798]_ );
  assign \new_[12045]_  = \new_[6170]_  ^ \new_[6470]_ ;
  assign \new_[12046]_  = (~\new_[13315]_  | ~\new_[3465]_ ) & (~\new_[11727]_  | ~\new_[14096]_ );
  assign \new_[12047]_  = ~\new_[12709]_  | ~\new_[13248]_ ;
  assign \new_[12048]_  = ~\new_[12346]_ ;
  assign \new_[12049]_  = ~\new_[12338]_ ;
  assign \new_[12050]_  = ~\new_[12698]_  & (~\new_[13180]_  | ~\new_[13094]_ );
  assign \new_[12051]_  = ~\new_[12351]_ ;
  assign \new_[12052]_  = ~\new_[14156]_  | ~\new_[12500]_ ;
  assign \new_[12053]_  = ~\new_[13568]_  | ~\new_[4800]_ ;
  assign \new_[12054]_  = \new_[13027]_  & \new_[12516]_ ;
  assign \new_[12055]_  = ~\new_[12894]_  | ~\new_[13285]_ ;
  assign \new_[12056]_  = ~\new_[12464]_ ;
  assign \new_[12057]_  = ~\new_[13978]_  | ~\new_[4799]_ ;
  assign \new_[12058]_  = ~\new_[12368]_ ;
  assign \new_[12059]_  = ~\new_[12548]_  & ~\new_[12966]_ ;
  assign n8745 = \sram_data_i[14]  ? \new_[13178]_  : \new_[11355]_ ;
  assign \new_[12061]_  = ~\new_[4840]_  | ~\new_[12610]_ ;
  assign \new_[12062]_  = ~\new_[2875]_  | ~\new_[14200]_ ;
  assign \new_[12063]_  = ~\new_[6696]_  & ~\new_[6261]_ ;
  assign \new_[12064]_  = ~\new_[3889]_  | ~\new_[3884]_ ;
  assign \new_[12065]_  = ~\new_[6293]_  & ~\new_[6716]_ ;
  assign \new_[12066]_  = ~\new_[6346]_  & ~\new_[6347]_ ;
  assign \new_[12067]_  = ~\new_[12368]_ ;
  assign \new_[12068]_  = ~\new_[12372]_ ;
  assign \new_[12069]_  = ~\new_[12445]_ ;
  assign \new_[12070]_  = ~\new_[13978]_  & ~\new_[12760]_ ;
  assign \new_[12071]_  = (~\new_[14043]_  | ~\new_[3504]_ ) & (~\new_[13761]_  | ~\new_[3505]_ );
  assign \new_[12072]_  = ~\new_[6089]_  & ~\new_[6020]_ ;
  assign \new_[12073]_  = ~\new_[14679]_ ;
  assign \new_[12074]_  = ~\new_[6567]_  & ~\new_[6264]_ ;
  assign \new_[12075]_  = ~\new_[2990]_  & ~\new_[13298]_ ;
  assign \new_[12076]_  = \new_[6593]_  | \new_[6266]_ ;
  assign \new_[12077]_  = ~\new_[6588]_  & ~\new_[6303]_ ;
  assign \new_[12078]_  = ~\new_[4206]_  | ~\new_[4291]_ ;
  assign \new_[12079]_  = ~\new_[12375]_ ;
  assign \new_[12080]_  = ~\new_[4615]_  & ~\new_[4796]_ ;
  assign \new_[12081]_  = ~\new_[6281]_  & ~\new_[6718]_ ;
  assign \new_[12082]_  = ~\new_[13298]_  & ~\new_[12437]_ ;
  assign \new_[12083]_  = ~\new_[6279]_  & ~\new_[6696]_ ;
  assign \new_[12084]_  = ~\new_[6370]_  & ~\new_[6371]_ ;
  assign \new_[12085]_  = ~\new_[12488]_ ;
  assign \new_[12086]_  = ~\new_[12446]_ ;
  assign \new_[12087]_  = ~\new_[12719]_ ;
  assign \new_[12088]_  = ~\new_[12441]_ ;
  assign \new_[12089]_  = \new_[12580]_  & \new_[13937]_ ;
  assign \new_[12090]_  = ~\new_[6002]_  & ~\new_[6020]_ ;
  assign \new_[12091]_  = ~\new_[6549]_  & ~\new_[6718]_ ;
  assign \new_[12092]_  = ~\new_[12422]_ ;
  assign \new_[12093]_  = ~\new_[6547]_  & ~\new_[6696]_ ;
  assign \new_[12094]_  = ~\new_[3410]_  | ~\new_[12671]_ ;
  assign \new_[12095]_  = ~\new_[3930]_  | ~\new_[3888]_ ;
  assign \new_[12096]_  = ~\new_[2961]_  & ~\new_[13456]_ ;
  assign \new_[12097]_  = ~\new_[6322]_  & ~\new_[6234]_ ;
  assign \new_[12098]_  = ~\new_[6275]_  & ~\new_[6272]_ ;
  assign \new_[12099]_  = ~\new_[4091]_  | ~\new_[12562]_  | ~\new_[13778]_ ;
  assign \new_[12100]_  = ~\new_[12368]_ ;
  assign \new_[12101]_  = ~n8645;
  assign \new_[12102]_  = ~\new_[13424]_  & ~\new_[4800]_ ;
  assign \new_[12103]_  = ~\new_[12898]_ ;
  assign \new_[12104]_  = ~\new_[12787]_  | ~\new_[13357]_ ;
  assign \new_[12105]_  = ~\new_[13342]_  & ~\new_[12847]_ ;
  assign \new_[12106]_  = ~\new_[12896]_  | ~\new_[13381]_ ;
  assign \new_[12107]_  = ~\new_[12525]_  & ~\new_[6346]_ ;
  assign \new_[12108]_  = (~\new_[13393]_  | ~\new_[6733]_ ) & (~\new_[6602]_  | ~\new_[13733]_ );
  assign \new_[12109]_  = \new_[12929]_  & \new_[12696]_ ;
  assign \new_[12110]_  = \new_[13349]_  ^ \new_[13449]_ ;
  assign \new_[12111]_  = ~\new_[12667]_  & ~\new_[12786]_ ;
  assign \new_[12112]_  = ~\new_[12789]_  & ~\new_[12983]_ ;
  assign \new_[12113]_  = \new_[12780]_  & \new_[14348]_ ;
  assign \new_[12114]_  = ~\new_[4792]_  & ~\new_[12778]_ ;
  assign \new_[12115]_  = ~\new_[12998]_  & ~\new_[12759]_ ;
  assign \new_[12116]_  = ~\new_[13253]_  & (~\new_[12905]_  | ~\new_[13217]_ );
  assign \new_[12117]_  = ~\new_[13077]_  & (~\new_[13215]_  | ~\new_[13017]_ );
  assign \new_[12118]_  = ~\new_[12571]_  & (~\new_[3938]_  | ~\new_[13317]_ );
  assign \new_[12119]_  = ~\new_[12985]_  | ~\new_[12613]_ ;
  assign \new_[12120]_  = ~\new_[13077]_  & ~\new_[12655]_ ;
  assign \new_[12121]_  = ~\new_[14665]_ ;
  assign \new_[12122]_  = \new_[2175]_  ^ \new_[13169]_ ;
  assign \new_[12123]_  = ~\new_[6020]_  & ~\new_[6260]_ ;
  assign \new_[12124]_  = \new_[2857]_  & \new_[14200]_ ;
  assign \new_[12125]_  = ~\new_[14203]_  | ~\new_[12562]_  | ~\new_[3311]_ ;
  assign \new_[12126]_  = ~\new_[12982]_  & ~\new_[12824]_ ;
  assign \new_[12127]_  = ~\new_[12955]_  & ~\new_[12661]_ ;
  assign \new_[12128]_  = ~\new_[12313]_ ;
  assign \new_[12129]_  = \new_[12928]_  ^ \new_[13230]_ ;
  assign \new_[12130]_  = ~\new_[14700]_  & ~\new_[12734]_ ;
  assign \new_[12131]_  = ~\new_[12954]_  & (~\new_[12943]_  | ~\new_[13050]_ );
  assign \new_[12132]_  = ~\new_[13154]_  & (~\new_[13016]_  | ~\new_[12984]_ );
  assign \new_[12133]_  = \new_[12898]_  & \new_[3037]_ ;
  assign \new_[12134]_  = \new_[12888]_  & \new_[2737]_ ;
  assign \new_[12135]_  = ~\new_[4853]_  | ~\new_[8959]_ ;
  assign \new_[12136]_  = ~\new_[12788]_  | ~\new_[13497]_ ;
  assign \new_[12137]_  = ~\new_[12755]_  | (~\new_[6019]_  & ~\new_[6105]_ );
  assign \new_[12138]_  = \new_[12892]_  & \new_[4780]_ ;
  assign \new_[12139]_  = ~\new_[13074]_  | (~\new_[6008]_  & ~\new_[13371]_ );
  assign \new_[12140]_  = \new_[12900]_  & \new_[3410]_ ;
  assign \new_[12141]_  = ~\new_[12582]_  | ~\new_[13421]_ ;
  assign \new_[12142]_  = \new_[6743]_  | \new_[6253]_ ;
  assign \new_[12143]_  = \new_[12892]_  | \new_[4780]_ ;
  assign \new_[12144]_  = ~\new_[12428]_ ;
  assign \new_[12145]_  = ~\new_[13383]_  | ~\new_[8826]_  | ~\new_[12784]_  | ~\new_[8700]_ ;
  assign \new_[12146]_  = \new_[13386]_  | n8390;
  assign \new_[12147]_  = ~\new_[13568]_  & ~\new_[4800]_ ;
  assign \new_[12148]_  = ~\new_[12438]_ ;
  assign \new_[12149]_  = \new_[13386]_  | \new_[13135]_ ;
  assign \new_[12150]_  = ~\new_[12695]_  | ~\new_[13447]_ ;
  assign \new_[12151]_  = ~\new_[6287]_  & ~\new_[6284]_ ;
  assign \new_[12152]_  = ~\new_[12418]_ ;
  assign \new_[12153]_  = ~\new_[12458]_ ;
  assign \new_[12154]_  = ~\new_[4292]_  | ~\new_[4293]_ ;
  assign \new_[12155]_  = ~\new_[12781]_  | ~\new_[9405]_ ;
  assign \new_[12156]_  = ~\new_[6322]_  & (~\new_[13324]_  | ~\new_[13143]_ );
  assign n8815 = \sram_data_i[15]  ? \new_[13178]_  : \new_[11398]_ ;
  assign \new_[12158]_  = ~\new_[12842]_ ;
  assign \new_[12159]_  = ~\new_[12568]_  & ~\new_[13480]_ ;
  assign \new_[12160]_  = ~\new_[12404]_ ;
  assign \new_[12161]_  = \new_[12516]_  & \new_[13043]_ ;
  assign \new_[12162]_  = ~\new_[12873]_  & ~\new_[12856]_ ;
  assign \new_[12163]_  = ~\new_[12824]_  & ~\new_[12674]_ ;
  assign \new_[12164]_  = ~\new_[12450]_ ;
  assign \new_[12165]_  = ~\new_[12371]_ ;
  assign \new_[12166]_  = ~\new_[13365]_  & ~\new_[13355]_ ;
  assign \new_[12167]_  = ~\new_[12992]_  | ~\new_[12959]_  | ~\new_[13105]_ ;
  assign n8795 = \sram_data_i[22]  ? \new_[13178]_  : \new_[11386]_ ;
  assign \new_[12169]_  = ~\new_[13316]_  | ~\new_[9405]_  | ~\new_[12781]_  | ~\new_[9421]_ ;
  assign \new_[12170]_  = ~\new_[6253]_  & ~\new_[12921]_ ;
  assign \new_[12171]_  = ~\new_[3777]_  | ~\new_[3711]_ ;
  assign \new_[12172]_  = ~\new_[2873]_  & ~\new_[2836]_ ;
  assign n8785 = \sram_data_i[17]  ? \new_[13178]_  : \new_[11383]_ ;
  assign n8735 = \sram_data_i[8]  ? \new_[13178]_  : \new_[11352]_ ;
  assign \new_[12175]_  = ~\new_[12311]_ ;
  assign \new_[12176]_  = \new_[12628]_  | \new_[13413]_ ;
  assign \new_[12177]_  = ~\new_[12856]_  & ~\new_[13307]_ ;
  assign \new_[12178]_  = ~\new_[12679]_  | ~\new_[13245]_ ;
  assign \new_[12179]_  = ~\new_[13087]_  | ~\new_[12995]_  | ~\new_[12984]_ ;
  assign \new_[12180]_  = \new_[14026]_  ^ \new_[14058]_ ;
  assign \new_[12181]_  = ~\new_[12902]_  & ~\new_[12736]_ ;
  assign \new_[12182]_  = ~\new_[13469]_  & ~\new_[13257]_ ;
  assign n8690 = \sram_data_i[19]  ? \new_[13178]_  : \new_[11083]_ ;
  assign \new_[12184]_  = ~\new_[12784]_  | ~\new_[8826]_ ;
  assign \new_[12185]_  = ~\new_[12879]_  | ~\new_[2091]_ ;
  assign \new_[12186]_  = ~\new_[12686]_  & ~\new_[13360]_ ;
  assign \new_[12187]_  = ~\new_[12537]_  & ~\new_[13444]_ ;
  assign \new_[12188]_  = ~\new_[12307]_ ;
  assign \new_[12189]_  = ~\new_[12864]_  & ~\new_[12546]_ ;
  assign \new_[12190]_  = ~\new_[12479]_ ;
  assign \new_[12191]_  = \new_[13128]_  & \new_[13431]_ ;
  assign n8740 = \sram_data_i[26]  ? \new_[13178]_  : \new_[11354]_ ;
  assign \new_[12193]_  = \new_[12684]_  & \new_[13389]_ ;
  assign \new_[12194]_  = ~\new_[12229]_ ;
  assign \new_[12195]_  = ~\new_[12429]_ ;
  assign \new_[12196]_  = ~\new_[12227]_ ;
  assign \new_[12197]_  = ~\new_[13296]_ ;
  assign \new_[12198]_  = ~\new_[13035]_  & ~\new_[12515]_ ;
  assign \new_[12199]_  = ~\new_[12533]_  & ~\new_[13147]_ ;
  assign \new_[12200]_  = \new_[12949]_  & \new_[12684]_ ;
  assign \new_[12201]_  = ~\new_[6370]_  & (~\new_[13461]_  | ~\new_[13038]_ );
  assign n8800 = \sram_data_i[13]  ? \new_[13178]_  : \new_[11387]_ ;
  assign n8670 = \sram_data_i[28]  ? \new_[13178]_  : \new_[11028]_ ;
  assign \new_[12204]_  = \new_[3710]_  & \new_[3930]_ ;
  assign \new_[12205]_  = \new_[3710]_  ^ \new_[3930]_ ;
  assign \new_[12206]_  = \new_[6341]_  & \new_[6592]_ ;
  assign n8685 = \new_[6341]_  ^ \new_[6592]_ ;
  assign \new_[12208]_  = \new_[3502]_  & \new_[3777]_ ;
  assign \new_[12209]_  = \new_[3502]_  ^ \new_[3777]_ ;
  assign \new_[12210]_  = \new_[3337]_  & \new_[3503]_ ;
  assign \new_[12211]_  = \new_[3337]_  ^ \new_[3503]_ ;
  assign \new_[12212]_  = \new_[4095]_  & \new_[4292]_ ;
  assign \new_[12213]_  = \new_[4095]_  ^ \new_[4292]_ ;
  assign \new_[12214]_  = \new_[13076]_  & \new_[13233]_ ;
  assign \new_[12215]_  = ~\new_[13207]_  & ~\new_[13043]_ ;
  assign \new_[12216]_  = ~\new_[14503]_ ;
  assign \new_[12217]_  = ~\new_[12781]_ ;
  assign \new_[12218]_  = \new_[6019]_  ? \new_[6018]_  : \new_[13770]_ ;
  assign \new_[12219]_  = ~\new_[6561]_  & ~\new_[13324]_ ;
  assign \new_[12220]_  = ~\new_[13990]_  | ~\new_[13505]_  | ~\new_[14051]_  | ~\new_[13526]_ ;
  assign \new_[12221]_  = \new_[6239]_  ^ \new_[6015]_ ;
  assign \new_[12222]_  = \new_[6241]_  ^ \new_[6033]_ ;
  assign \new_[12223]_  = ~\new_[12990]_  | ~\new_[13090]_ ;
  assign \new_[12224]_  = ~\new_[13054]_  | ~\new_[13088]_ ;
  assign \new_[12225]_  = ~\new_[12997]_  | ~\new_[13009]_ ;
  assign \new_[12226]_  = \new_[13184]_  & \new_[13254]_ ;
  assign \new_[12227]_  = ~\new_[13081]_  | ~\new_[2871]_ ;
  assign \new_[12228]_  = ~\new_[12665]_ ;
  assign \new_[12229]_  = ~\new_[13068]_  & ~\new_[3030]_ ;
  assign \new_[12230]_  = ~\new_[12912]_  | ~\new_[13103]_ ;
  assign \new_[12231]_  = ~\wb_data_i[22]  | ~\new_[13162]_ ;
  assign \new_[12232]_  = ~\new_[13105]_  | ~\new_[13066]_ ;
  assign \new_[12233]_  = ~\new_[13023]_  | ~\new_[13213]_ ;
  assign \new_[12234]_  = ~\new_[12904]_  | ~\new_[13063]_ ;
  assign n8645 = ~\new_[13448]_  & ~\new_[13197]_ ;
  assign \new_[12236]_  = ~\new_[12882]_ ;
  assign \new_[12237]_  = \new_[12924]_  & \new_[13066]_ ;
  assign \new_[12238]_  = ~\new_[13117]_  | ~\new_[14453]_ ;
  assign n8855 = ~\new_[12532]_ ;
  assign \new_[12240]_  = ~\new_[3062]_  | ~\new_[13908]_  | ~\new_[13224]_  | ~\new_[14163]_ ;
  assign \new_[12241]_  = ~\new_[13245]_  | ~\new_[13217]_ ;
  assign \new_[12242]_  = ~\new_[2091]_  | ~\new_[2093]_  | ~\new_[13278]_  | ~\new_[2092]_ ;
  assign \new_[12243]_  = ~\new_[8701]_  | ~\new_[8658]_  | ~\new_[13356]_  | ~\new_[8826]_ ;
  assign \new_[12244]_  = ~\new_[14503]_ ;
  assign \new_[12245]_  = ~phy_rst_pad_o;
  assign \new_[12246]_  = ~\new_[13007]_  & ~\new_[13029]_ ;
  assign \new_[12247]_  = ~\new_[13037]_  & ~\new_[3482]_ ;
  assign \new_[12248]_  = ~\new_[12938]_  | ~\new_[12935]_ ;
  assign \new_[12249]_  = ~\new_[13426]_  & ~\new_[13740]_ ;
  assign \new_[12250]_  = ~\new_[12991]_  & ~\new_[14211]_ ;
  assign \new_[12251]_  = ~\new_[13030]_  & ~\new_[2453]_ ;
  assign \new_[12252]_  = ~\new_[14503]_ ;
  assign \new_[12253]_  = \new_[2962]_  ^ \new_[6019]_ ;
  assign \new_[12254]_  = ~\new_[13304]_  | ~\new_[13021]_ ;
  assign \new_[12255]_  = ~\new_[14503]_ ;
  assign \new_[12256]_  = ~\new_[3340]_  & ~\new_[13065]_ ;
  assign \new_[12257]_  = ~\new_[12699]_ ;
  assign \new_[12258]_  = ~\new_[14503]_ ;
  assign \new_[12259]_  = ~\wb_data_i[23]  | ~\new_[12197]_ ;
  assign \new_[12260]_  = \new_[13085]_  | \new_[4677]_ ;
  assign \new_[12261]_  = ~\new_[12914]_  & ~\wb_addr_i[4] ;
  assign \new_[12262]_  = ~\new_[2873]_  & ~\new_[13895]_ ;
  assign \new_[12263]_  = ~\new_[12746]_ ;
  assign \new_[12264]_  = ~\new_[13193]_  & ~\new_[2348]_ ;
  assign \new_[12265]_  = ~\new_[6716]_  & ~\new_[6262]_ ;
  assign \new_[12266]_  = ~\new_[4683]_  | ~\new_[13428]_ ;
  assign \new_[12267]_  = ~\new_[13464]_  & ~\new_[13138]_ ;
  assign n8850 = ~\new_[12976]_  & ~\new_[13732]_ ;
  assign \new_[12269]_  = \new_[13418]_  ^ \new_[13453]_ ;
  assign \new_[12270]_  = \new_[14089]_  & \new_[13219]_ ;
  assign \new_[12271]_  = \new_[12991]_  | \new_[14036]_ ;
  assign \new_[12272]_  = ~\new_[13947]_  | ~\new_[3671]_ ;
  assign n8845 = ~\new_[13089]_  | ~\new_[13933]_ ;
  assign \new_[12274]_  = \new_[7310]_  & \new_[13091]_ ;
  assign \new_[12275]_  = ~\new_[13116]_  & ~\wb_addr_i[4] ;
  assign \new_[12276]_  = \new_[12948]_  | \new_[6301]_ ;
  assign \new_[12277]_  = ~\new_[12806]_ ;
  assign \new_[12278]_  = ~\new_[12671]_ ;
  assign \new_[12279]_  = ~\new_[6552]_  & ~\new_[13461]_ ;
  assign \new_[12280]_  = u4_attach_r1_reg;
  assign \new_[12281]_  = ~\new_[13191]_  | ~\new_[13222]_ ;
  assign \new_[12282]_  = ~\new_[12872]_ ;
  assign \new_[12283]_  = ~\new_[13171]_  & ~\new_[13240]_ ;
  assign \new_[12284]_  = \new_[12963]_  | \new_[13274]_ ;
  assign \new_[12285]_  = \new_[13158]_  | \new_[13275]_ ;
  assign \new_[12286]_  = ~\new_[13280]_  | ~\new_[12950]_ ;
  assign \new_[12287]_  = ~\new_[13664]_  | ~\new_[13428]_ ;
  assign \new_[12288]_  = ~\new_[13218]_  | ~\new_[13089]_ ;
  assign \new_[12289]_  = ~\new_[12600]_ ;
  assign \new_[12290]_  = \new_[13161]_  | \new_[3308]_ ;
  assign \new_[12291]_  = ~\new_[13062]_  & ~\new_[13291]_ ;
  assign \new_[12292]_  = ~\new_[12542]_ ;
  assign \new_[12293]_  = ~\new_[4779]_  | ~\new_[13428]_ ;
  assign \new_[12294]_  = ~\new_[13941]_  | ~\new_[3468]_ ;
  assign \new_[12295]_  = ~\new_[13428]_  | ~\new_[14261]_ ;
  assign \new_[12296]_  = ~\new_[13710]_  | ~\new_[13428]_ ;
  assign \new_[12297]_  = ~\new_[13060]_  & ~\new_[3692]_ ;
  assign \new_[12298]_  = ~\new_[13432]_  | ~\new_[12934]_ ;
  assign \new_[12299]_  = ~\new_[13183]_  | ~\new_[13223]_ ;
  assign \new_[12300]_  = ~\new_[13100]_  | ~\new_[13172]_ ;
  assign \new_[12301]_  = ~\new_[12521]_ ;
  assign \new_[12302]_  = \new_[13190]_  | \new_[13270]_ ;
  assign \new_[12303]_  = ~\new_[13148]_  | ~\new_[13198]_ ;
  assign \new_[12304]_  = \new_[13112]_  | \new_[13260]_ ;
  assign \new_[12305]_  = ~\new_[12962]_  & ~\new_[13480]_ ;
  assign \new_[12306]_  = \new_[13027]_  & \new_[13023]_ ;
  assign \new_[12307]_  = ~\new_[13243]_  | ~\new_[13106]_ ;
  assign \new_[12308]_  = ~\new_[13033]_  | ~\new_[13051]_ ;
  assign \new_[12309]_  = ~\new_[13088]_  | ~\new_[13133]_ ;
  assign \new_[12310]_  = ~\new_[12692]_ ;
  assign \new_[12311]_  = \new_[13000]_  & \new_[13131]_ ;
  assign \new_[12312]_  = ~\new_[12810]_ ;
  assign \new_[12313]_  = ~\new_[13032]_  | ~\new_[13245]_ ;
  assign \new_[12314]_  = ~\new_[13008]_  | ~\new_[13196]_ ;
  assign \new_[12315]_  = ~\new_[13239]_  & ~\new_[13102]_ ;
  assign \new_[12316]_  = ~\new_[12534]_ ;
  assign \new_[12317]_  = \new_[13133]_  & \new_[13086]_ ;
  assign \new_[12318]_  = ~\new_[13101]_  | ~\new_[13017]_ ;
  assign \new_[12319]_  = ~\new_[13064]_  | ~\new_[13106]_ ;
  assign \new_[12320]_  = ~\new_[12935]_  | ~\new_[13076]_ ;
  assign \new_[12321]_  = \new_[13109]_  & \new_[13094]_ ;
  assign \new_[12322]_  = ~\new_[13102]_  & ~\new_[12994]_ ;
  assign \new_[12323]_  = \new_[13051]_  & \new_[13249]_ ;
  assign \new_[12324]_  = ~\new_[12626]_ ;
  assign \new_[12325]_  = \new_[2983]_  ^ \new_[6015]_ ;
  assign \new_[12326]_  = \new_[6243]_  ^ \new_[5978]_ ;
  assign \new_[12327]_  = \new_[13194]_  & \new_[13050]_ ;
  assign \new_[12328]_  = ~\new_[13001]_  | ~\new_[13009]_ ;
  assign \new_[12329]_  = ~\new_[13999]_  | ~\new_[14247]_  | ~\new_[13502]_  | ~\new_[13594]_ ;
  assign \new_[12330]_  = ~\new_[13921]_  | ~\new_[13628]_  | ~\new_[14019]_  | ~\new_[13654]_ ;
  assign \new_[12331]_  = ~\new_[13847]_  | ~\new_[14053]_  | ~\new_[13916]_  | ~\new_[13576]_ ;
  assign \new_[12332]_  = ~\new_[14124]_  | ~\new_[13993]_  | ~\new_[13759]_  | ~\new_[14105]_ ;
  assign \new_[12333]_  = ~\new_[13531]_  | ~\new_[13644]_  | ~\new_[13547]_  | ~\new_[13530]_ ;
  assign \new_[12334]_  = ~\new_[12197]_  | ~\dma_req_o[0] ;
  assign \new_[12335]_  = ~\new_[6091]_  | ~\new_[13746]_ ;
  assign \new_[12336]_  = ~\new_[12753]_ ;
  assign \new_[12337]_  = \new_[3467]_  ^ \new_[6012]_ ;
  assign \new_[12338]_  = \new_[13213]_  & \new_[12918]_ ;
  assign \new_[12339]_  = ~\new_[14503]_ ;
  assign \new_[12340]_  = \new_[13284]_  ^ \new_[13862]_ ;
  assign \new_[12341]_  = \new_[6386]_  ^ \new_[13302]_ ;
  assign \new_[12342]_  = ~\new_[12824]_ ;
  assign \new_[12343]_  = ~\new_[12497]_ ;
  assign \new_[12344]_  = \new_[6093]_  ^ \new_[6385]_ ;
  assign \new_[12345]_  = \new_[13284]_  ^ \new_[2042]_ ;
  assign \new_[12346]_  = ~\new_[13031]_  | ~\new_[13079]_ ;
  assign \new_[12347]_  = \new_[4069]_  ^ \new_[6305]_ ;
  assign \new_[12348]_  = ~\new_[12840]_ ;
  assign \new_[12349]_  = ~\new_[13047]_  & ~\wb_addr_i[4] ;
  assign \new_[12350]_  = ~\new_[2874]_  | ~\new_[13756]_ ;
  assign \new_[12351]_  = ~\new_[13043]_  | ~\new_[13042]_ ;
  assign \new_[12352]_  = ~\new_[12703]_ ;
  assign \new_[12353]_  = ~\new_[2454]_  | ~\new_[13595]_ ;
  assign \new_[12354]_  = \new_[4864]_  | \new_[13096]_ ;
  assign \new_[12355]_  = (~\new_[3462]_  | ~\new_[13866]_ ) & (~\new_[3308]_  | ~\new_[13779]_ );
  assign \new_[12356]_  = \new_[4619]_  | \new_[13096]_ ;
  assign \new_[12357]_  = ~\new_[12663]_ ;
  assign \new_[12358]_  = ~\new_[12525]_ ;
  assign \new_[12359]_  = ~\new_[13754]_  | ~\new_[3932]_ ;
  assign n8830 = ~n9145 & ~\new_[14242]_ ;
  assign \new_[12361]_  = ~\new_[13569]_  & ~\new_[4852]_ ;
  assign \new_[12362]_  = ~\new_[13214]_  & ~\new_[4779]_ ;
  assign \new_[12363]_  = ~\new_[4794]_  | ~\new_[13136]_ ;
  assign \new_[12364]_  = ~\new_[5997]_  & ~\new_[13598]_ ;
  assign \new_[12365]_  = ~\new_[13075]_  | ~\new_[12997]_ ;
  assign \new_[12366]_  = ~\new_[13302]_  & ~\new_[14254]_ ;
  assign \new_[12367]_  = ~\new_[6254]_  & ~\new_[13413]_ ;
  assign \new_[12368]_  = ~rst_i;
  assign \new_[12369]_  = ~\new_[12865]_ ;
  assign \new_[12370]_  = ~\new_[12686]_ ;
  assign \new_[12371]_  = ~\new_[13631]_  | ~\new_[13980]_ ;
  assign \new_[12372]_  = ~\new_[13978]_  | ~\new_[14205]_ ;
  assign \new_[12373]_  = ~\new_[12530]_ ;
  assign \new_[12374]_  = ~\new_[12674]_ ;
  assign \new_[12375]_  = ~\new_[14015]_  | ~\new_[13914]_ ;
  assign \new_[12376]_  = ~\new_[12740]_ ;
  assign \new_[12377]_  = ~\new_[12531]_ ;
  assign \new_[12378]_  = ~\new_[12873]_ ;
  assign \new_[12379]_  = ~\new_[12547]_ ;
  assign \new_[12380]_  = ~\new_[12785]_ ;
  assign \new_[12381]_  = ~\new_[2090]_  | ~\new_[6246]_ ;
  assign \new_[12382]_  = ~\new_[12667]_ ;
  assign \new_[12383]_  = ~\new_[3881]_  | ~\new_[13429]_  | ~\new_[13682]_ ;
  assign \new_[12384]_  = ~\new_[12717]_ ;
  assign \new_[12385]_  = (~\new_[3592]_  | ~\new_[13941]_ ) & (~\new_[3309]_  | ~\new_[13624]_ );
  assign \new_[12386]_  = ~\new_[12197]_  | ~\dma_req_o[3] ;
  assign \new_[12387]_  = ~\new_[14503]_ ;
  assign \new_[12388]_  = ~\new_[12939]_  | ~\new_[13094]_ ;
  assign \new_[12389]_  = \new_[13179]_  & \new_[13399]_ ;
  assign \new_[12390]_  = ~\new_[13097]_  | ~\new_[13050]_ ;
  assign \new_[12391]_  = \new_[13328]_  ^ \new_[13349]_ ;
  assign \new_[12392]_  = \new_[13449]_  ^ \new_[13433]_ ;
  assign \new_[12393]_  = \new_[13446]_  ^ \new_[13343]_ ;
  assign \new_[12394]_  = ~\new_[12922]_  & ~\new_[12938]_ ;
  assign \new_[12395]_  = ~\new_[12968]_  | ~\new_[13131]_ ;
  assign \new_[12396]_  = \new_[6020]_ ;
  assign \new_[12397]_  = \new_[3035]_  ^ \new_[13297]_ ;
  assign \new_[12398]_  = ~\new_[12625]_ ;
  assign \new_[12399]_  = ~\new_[4774]_  | ~\new_[13428]_ ;
  assign \new_[12400]_  = ~\new_[13043]_  | ~\new_[13023]_ ;
  assign \new_[12401]_  = ~\new_[4096]_  & ~\new_[13070]_ ;
  assign \new_[12402]_  = ~\new_[2874]_  & ~\new_[13756]_ ;
  assign \new_[12403]_  = ~\new_[9412]_  | ~\new_[9372]_  | ~\new_[13495]_  | ~\new_[9405]_ ;
  assign \new_[12404]_  = ~\new_[12654]_ ;
  assign \new_[12405]_  = ~\new_[12984]_  | ~\new_[13082]_ ;
  assign \new_[12406]_  = \new_[13168]_  & \new_[13051]_ ;
  assign \new_[12407]_  = ~\new_[12946]_  | ~\new_[13034]_ ;
  assign \new_[12408]_  = ~\new_[12553]_ ;
  assign \new_[12409]_  = \new_[13090]_  & \new_[13059]_ ;
  assign \new_[12410]_  = ~\new_[13221]_  & ~\new_[13324]_ ;
  assign \new_[12411]_  = ~\new_[13095]_  | ~\new_[13097]_ ;
  assign \new_[12412]_  = \new_[13056]_  | \new_[3283]_ ;
  assign \new_[12413]_  = ~\new_[12197]_  | ~\dma_req_o[2] ;
  assign \new_[12414]_  = ~\new_[12560]_ ;
  assign \new_[12415]_  = ~\new_[13116]_ ;
  assign \new_[12416]_  = ~\new_[12883]_ ;
  assign \new_[12417]_  = ~\new_[12780]_ ;
  assign \new_[12418]_  = ~\new_[13167]_  & ~\wb_addr_i[4] ;
  assign \new_[12419]_  = ~\new_[12974]_  & ~\new_[3317]_ ;
  assign \new_[12420]_  = ~\new_[6246]_  & ~\new_[2611]_ ;
  assign \new_[12421]_  = ~\new_[12951]_  & ~\new_[4074]_ ;
  assign \new_[12422]_  = ~\new_[13930]_  & ~\new_[14084]_ ;
  assign \new_[12423]_  = \new_[3312]_  ^ \new_[6326]_ ;
  assign \new_[12424]_  = ~\new_[13141]_  | ~\new_[12909]_ ;
  assign \new_[12425]_  = ~\new_[12938]_  | ~\new_[13032]_ ;
  assign \new_[12426]_  = ~\new_[12779]_ ;
  assign \new_[12427]_  = ~\new_[12713]_ ;
  assign \new_[12428]_  = ~\new_[13664]_  & ~\new_[13710]_ ;
  assign \new_[12429]_  = ~\new_[2343]_  & ~\new_[13020]_ ;
  assign \new_[12430]_  = ~\new_[13621]_  | ~\new_[13617]_ ;
  assign \new_[12431]_  = ~\new_[12797]_ ;
  assign n8390 = ~\new_[13155]_ ;
  assign \new_[12433]_  = ~\new_[13327]_  & ~\new_[13616]_ ;
  assign \new_[12434]_  = ~\new_[13125]_  | ~\new_[12964]_ ;
  assign \new_[12435]_  = \new_[13113]_  & \new_[13488]_ ;
  assign \new_[12436]_  = ~\new_[12793]_ ;
  assign \new_[12437]_  = \\u0_u0_state_reg[0] ;
  assign \new_[12438]_  = ~\new_[14221]_  | ~\new_[14082]_ ;
  assign \new_[12439]_  = ~\new_[12809]_ ;
  assign \new_[12440]_  = ~\new_[6198]_  | ~\new_[14147]_ ;
  assign \new_[12441]_  = ~\new_[13629]_  | ~\new_[14195]_ ;
  assign \new_[12442]_  = ~\new_[14503]_ ;
  assign \new_[12443]_  = \new_[13710]_  | \new_[14261]_ ;
  assign \new_[12444]_  = ~\new_[14046]_  | ~\new_[4774]_ ;
  assign \new_[12445]_  = ~\new_[14069]_  | ~\new_[13924]_ ;
  assign \new_[12446]_  = ~\new_[13552]_  | ~\new_[14199]_ ;
  assign \new_[12447]_  = ~\new_[12828]_ ;
  assign \new_[12448]_  = \new_[2932]_  ^ \new_[4852]_ ;
  assign \new_[12449]_  = ~\new_[12835]_ ;
  assign \new_[12450]_  = ~\new_[12947]_  & ~\new_[12914]_ ;
  assign \new_[12451]_  = ~\new_[6166]_  & ~\new_[13355]_ ;
  assign \new_[12452]_  = ~\\u4_u1_buf0_orig_m3_reg[0] ;
  assign n8835 = ~\new_[14738]_ ;
  assign \new_[12454]_  = \new_[13039]_  & \new_[13082]_ ;
  assign \new_[12455]_  = ~\new_[12851]_ ;
  assign \new_[12456]_  = \new_[2372]_  & \new_[13813]_ ;
  assign \new_[12457]_  = ~\new_[13595]_  | ~\new_[3177]_ ;
  assign \new_[12458]_  = \new_[6718]_  ^ \new_[6696]_ ;
  assign \new_[12459]_  = ~\new_[13011]_  & ~\new_[13461]_ ;
  assign \new_[12460]_  = ~\new_[12650]_ ;
  assign \new_[12461]_  = ~\new_[4666]_  | ~\new_[13428]_ ;
  assign \new_[12462]_  = ~\new_[12619]_ ;
  assign \new_[12463]_  = ~\new_[13666]_  | ~\new_[13819]_ ;
  assign \new_[12464]_  = ~\new_[13018]_  | ~\new_[13442]_ ;
  assign \new_[12465]_  = \new_[6240]_  ^ \new_[6016]_ ;
  assign \new_[12466]_  = ~\new_[3713]_  & ~\new_[13188]_ ;
  assign \new_[12467]_  = ~\new_[13595]_  | ~\new_[3895]_ ;
  assign \new_[12468]_  = ~\new_[12994]_  | ~\new_[12990]_ ;
  assign \new_[12469]_  = ~\new_[12197]_  | ~\dma_req_o[1] ;
  assign \new_[12470]_  = \new_[13244]_  | \new_[3282]_ ;
  assign \new_[12471]_  = ~\new_[12502]_ ;
  assign \new_[12472]_  = ~\new_[12969]_  | ~\new_[13217]_ ;
  assign \new_[12473]_  = \new_[12923]_  | \new_[3309]_ ;
  assign \new_[12474]_  = ~\new_[13292]_  | ~\new_[13002]_ ;
  assign \new_[12475]_  = ~\new_[12784]_ ;
  assign \new_[12476]_  = \new_[2985]_  ^ \new_[6016]_ ;
  assign \new_[12477]_  = \new_[2987]_  ^ \new_[5978]_ ;
  assign \new_[12478]_  = \new_[3687]_  ^ \new_[6556]_ ;
  assign \new_[12479]_  = ~\new_[13111]_  | ~\new_[13214]_ ;
  assign \new_[12480]_  = \new_[2986]_  ^ \new_[6033]_ ;
  assign \new_[12481]_  = ~\new_[12921]_  & ~\new_[13413]_ ;
  assign \new_[12482]_  = ~\new_[12608]_ ;
  assign \new_[12483]_  = ~\new_[13751]_  | ~\new_[13656]_ ;
  assign \new_[12484]_  = ~\new_[13042]_  | ~\new_[13064]_ ;
  assign \new_[12485]_  = ~\new_[12933]_  & ~\new_[13445]_ ;
  assign \new_[12486]_  = ~\new_[14503]_ ;
  assign \new_[12487]_  = ~\new_[13228]_  | ~\new_[2476]_ ;
  assign \new_[12488]_  = ~\new_[2872]_  & ~\new_[2871]_ ;
  assign \new_[12489]_  = ~\new_[12624]_ ;
  assign n8840 = ~\new_[12782]_ ;
  assign \new_[12491]_  = ~\new_[14503]_ ;
  assign \new_[12492]_  = \new_[13732]_  & \new_[13815]_ ;
  assign \new_[12493]_  = \new_[13732]_  ^ \new_[13815]_ ;
  assign \new_[12494]_  = \new_[13735]_  & \new_[13799]_ ;
  assign \new_[12495]_  = \new_[13735]_  ^ \new_[13799]_ ;
  assign \new_[12496]_  = ~\new_[6344]_  & ~\new_[6343]_ ;
  assign \new_[12497]_  = \new_[14018]_  ^ \new_[14032]_ ;
  assign \new_[12498]_  = \new_[14211]_  | \new_[14036]_ ;
  assign \new_[12499]_  = ~\new_[13028]_ ;
  assign \new_[12500]_  = ~\new_[13398]_  & ~\new_[13386]_ ;
  assign \new_[12501]_  = ~\new_[6304]_  | ~\new_[13550]_ ;
  assign \new_[12502]_  = ~u4_u1_r5_reg;
  assign \new_[12503]_  = (~\new_[14033]_  | ~\new_[5761]_ ) & (~\new_[14180]_  | ~\new_[3739]_ );
  assign \new_[12504]_  = ~\new_[12906]_ ;
  assign \new_[12505]_  = ~\new_[13162]_ ;
  assign \new_[12506]_  = ~\new_[13080]_ ;
  assign \new_[12507]_  = (~\new_[2573]_  | ~\new_[13512]_ ) & (~\new_[4778]_  | ~\new_[13734]_ );
  assign \new_[12508]_  = ~\new_[12912]_ ;
  assign \new_[12509]_  = ~\new_[4236]_  & ~\new_[3932]_ ;
  assign \new_[12510]_  = ~\new_[13694]_  & ~\new_[13608]_ ;
  assign \new_[12511]_  = \new_[13276]_  & \new_[13358]_ ;
  assign \new_[12512]_  = ~\new_[13417]_  & ~\new_[6351]_ ;
  assign \new_[12513]_  = ~\new_[13286]_  & ~\new_[6348]_ ;
  assign \new_[12514]_  = \new_[13886]_  ^ \new_[14018]_ ;
  assign \new_[12515]_  = ~\new_[13046]_ ;
  assign \new_[12516]_  = ~\new_[13207]_ ;
  assign \new_[12517]_  = ~\new_[12940]_ ;
  assign \new_[12518]_  = \new_[13309]_  & \new_[13357]_ ;
  assign \new_[12519]_  = ~\new_[13427]_  & ~\wb_addr_i[4] ;
  assign \new_[12520]_  = ~\new_[13313]_  | ~\new_[13420]_ ;
  assign \new_[12521]_  = ~\new_[13387]_  & ~\new_[13396]_ ;
  assign \new_[12522]_  = ~\new_[6268]_  & ~\new_[6716]_ ;
  assign \new_[12523]_  = ~\new_[12948]_ ;
  assign \new_[12524]_  = ~\new_[4293]_  | ~\new_[4206]_ ;
  assign \new_[12525]_  = ~\new_[13584]_  | ~\new_[14108]_ ;
  assign \new_[12526]_  = \new_[13620]_  ^ \new_[14000]_ ;
  assign \new_[12527]_  = \new_[13334]_  & \new_[13325]_ ;
  assign \new_[12528]_  = ~\new_[3790]_  | ~\new_[3282]_ ;
  assign \new_[12529]_  = ~\new_[12956]_ ;
  assign \new_[12530]_  = ~\new_[14001]_  | ~\new_[13264]_ ;
  assign \new_[12531]_  = ~\new_[2874]_  & ~\new_[2836]_ ;
  assign \new_[12532]_  = ~\new_[2989]_  | ~\new_[3013]_  | ~\new_[13483]_  | ~\new_[2988]_ ;
  assign \new_[12533]_  = ~\new_[13196]_ ;
  assign \new_[12534]_  = ~\new_[13353]_  & ~\new_[13375]_ ;
  assign \new_[12535]_  = ~\new_[6563]_  | ~\new_[3342]_ ;
  assign n8870 = ~\new_[13448]_  & ~\new_[13441]_ ;
  assign \new_[12537]_  = ~\new_[13130]_ ;
  assign \new_[12538]_  = \new_[6275]_  & \new_[3712]_ ;
  assign n8875 = u4_suspend_r_reg;
  assign \new_[12540]_  = \new_[13458]_  & \new_[13348]_ ;
  assign \new_[12541]_  = ~\wb_addr_i[5]  & ~\wb_addr_i[6] ;
  assign \new_[12542]_  = ~\new_[13307]_  & ~\new_[13482]_ ;
  assign \new_[12543]_  = ~\new_[13251]_ ;
  assign \new_[12544]_  = ~\new_[13147]_ ;
  assign \new_[12545]_  = ~\new_[13198]_ ;
  assign \new_[12546]_  = ~\new_[12909]_ ;
  assign \new_[12547]_  = ~\new_[6253]_  & ~\new_[4237]_ ;
  assign \new_[12548]_  = ~\new_[13305]_  | ~\new_[13395]_ ;
  assign \new_[12549]_  = \\u4_utmi_vend_stat_r_reg[5] ;
  assign \new_[12550]_  = ~\new_[6253]_  | ~\new_[4237]_ ;
  assign \new_[12551]_  = \new_[13431]_  & \wb_addr_i[4] ;
  assign \new_[12552]_  = ~\new_[13322]_  & ~\new_[13461]_ ;
  assign \new_[12553]_  = ~\new_[13282]_  | ~\new_[13923]_ ;
  assign \new_[12554]_  = ~\new_[13356]_ ;
  assign \new_[12555]_  = \new_[13335]_  & \new_[13463]_ ;
  assign \new_[12556]_  = ~\new_[13070]_ ;
  assign \new_[12557]_  = ~\new_[6484]_  | ~\new_[6168]_ ;
  assign \new_[12558]_  = ~\new_[3507]_  & ~\new_[3626]_ ;
  assign \new_[12559]_  = \\u4_utmi_vend_stat_r_reg[2] ;
  assign \new_[12560]_  = ~\new_[13110]_ ;
  assign \new_[12561]_  = ~\new_[3339]_  & ~\new_[3429]_ ;
  assign \new_[12562]_  = ~\new_[4092]_  & ~\new_[3881]_ ;
  assign \new_[12563]_  = ~\new_[13444]_  & ~\new_[13275]_ ;
  assign \new_[12564]_  = ~\new_[13032]_ ;
  assign \new_[12565]_  = ~\new_[14424]_ ;
  assign \new_[12566]_  = ~\new_[12982]_ ;
  assign \new_[12567]_  = (~\new_[3466]_  | ~\new_[14120]_ ) & (~\new_[3310]_  | ~\new_[13643]_ );
  assign \new_[12568]_  = ~\new_[13216]_ ;
  assign \new_[12569]_  = \new_[13318]_  & \new_[13447]_ ;
  assign \new_[12570]_  = ~\new_[13200]_ ;
  assign \new_[12571]_  = ~\new_[13326]_  & ~\new_[6560]_ ;
  assign \new_[12572]_  = ~\new_[13003]_ ;
  assign \new_[12573]_  = ~\new_[14666]_ ;
  assign \new_[12574]_  = ~\new_[13150]_ ;
  assign \new_[12575]_  = ~\new_[13149]_ ;
  assign \new_[12576]_  = ~\new_[13042]_ ;
  assign \new_[12577]_  = ~\new_[12992]_ ;
  assign \new_[12578]_  = \new_[13412]_  & \new_[3471]_ ;
  assign \new_[12579]_  = ~\new_[13007]_ ;
  assign \new_[12580]_  = ~\new_[13261]_  & ~\new_[2476]_ ;
  assign \new_[12581]_  = ~\new_[12904]_ ;
  assign \new_[12582]_  = ~\new_[4096]_  & ~\new_[4098]_ ;
  assign \new_[12583]_  = ~\new_[3036]_  | ~\new_[13297]_ ;
  assign \new_[12584]_  = \new_[13479]_  & \new_[13381]_ ;
  assign \new_[12585]_  = ~\new_[13495]_ ;
  assign \new_[12586]_  = ~u0_u0_resume_req_s_reg;
  assign \new_[12587]_  = \\u4_utmi_vend_stat_r_reg[1] ;
  assign \new_[12588]_  = ~\new_[13858]_  | ~\new_[13481]_ ;
  assign \new_[12589]_  = ~\new_[13374]_  & ~\new_[13413]_ ;
  assign \new_[12590]_  = ~\new_[13363]_  & ~\new_[6461]_ ;
  assign \new_[12591]_  = ~\new_[14452]_ ;
  assign \new_[12592]_  = ~\new_[13353]_  & ~\new_[14035]_ ;
  assign \new_[12593]_  = ~\new_[13260]_  & ~\new_[14147]_ ;
  assign \new_[12594]_  = ~\new_[13490]_  & ~\new_[13324]_ ;
  assign \new_[12595]_  = ~\new_[13405]_  & ~\new_[13355]_ ;
  assign \new_[12596]_  = \new_[14028]_  ^ \new_[13889]_ ;
  assign \new_[12597]_  = ~\new_[13004]_ ;
  assign \new_[12598]_  = ~\new_[12922]_ ;
  assign \new_[12599]_  = \\u4_utmi_vend_stat_r_reg[7] ;
  assign \new_[12600]_  = \new_[13455]_  & \new_[13488]_ ;
  assign \new_[12601]_  = ~\new_[13148]_ ;
  assign \new_[12602]_  = \\u4_utmi_vend_stat_r_reg[4] ;
  assign \new_[12603]_  = \new_[13426]_  | \new_[4795]_ ;
  assign \new_[12604]_  = ~\new_[13095]_ ;
  assign \new_[12605]_  = ~\new_[13593]_  | ~\new_[13429]_  | ~\new_[4092]_ ;
  assign \new_[12606]_  = ~\new_[13858]_  & ~\new_[13481]_ ;
  assign \new_[12607]_  = ~\new_[13470]_  & ~\new_[6323]_ ;
  assign \new_[12608]_  = ~\new_[5999]_  & ~\new_[3341]_ ;
  assign \new_[12609]_  = \new_[13451]_  & \new_[13390]_ ;
  assign \new_[12610]_  = ~\new_[4801]_ ;
  assign \new_[12611]_  = \new_[13470]_  | \new_[13324]_ ;
  assign \new_[12612]_  = ~\new_[13866]_  | ~\new_[3313]_ ;
  assign \new_[12613]_  = ~\new_[13157]_ ;
  assign \new_[12614]_  = \\u4_utmi_vend_stat_r_reg[0] ;
  assign \new_[12615]_  = ~\new_[13480]_  & ~\new_[13274]_ ;
  assign \new_[12616]_  = ~\new_[13289]_  & ~\new_[6324]_ ;
  assign \new_[12617]_  = ~\new_[12967]_ ;
  assign \new_[12618]_  = ~\new_[6512]_  | ~\new_[13928]_ ;
  assign \new_[12619]_  = ~\new_[14135]_  | ~\new_[13437]_  | ~\new_[13987]_ ;
  assign \new_[12620]_  = ~\new_[13277]_  & ~\new_[13260]_ ;
  assign \new_[12621]_  = ~\new_[13521]_  & (~\new_[10667]_  | ~\new_[14020]_ );
  assign \new_[12622]_  = ~\new_[14237]_  & (~\new_[10631]_  | ~\new_[14126]_ );
  assign \new_[12623]_  = ~\new_[12977]_ ;
  assign \new_[12624]_  = ~\new_[6322]_  & (~\new_[13893]_  | ~\new_[6234]_ );
  assign \new_[12625]_  = \new_[13377]_  & \new_[13420]_ ;
  assign \new_[12626]_  = u5_wb_req_s1_reg;
  assign \new_[12627]_  = (~\new_[14074]_  | ~\new_[5617]_ ) & (~\new_[6611]_  | ~\new_[3878]_ );
  assign \new_[12628]_  = ~\new_[4286]_  | ~\new_[3283]_ ;
  assign \new_[12629]_  = (~\new_[14057]_  | ~\new_[5489]_ ) & (~\new_[14224]_  | ~\new_[2501]_ );
  assign \new_[12630]_  = (~\new_[14070]_  | ~\new_[2551]_ ) & (~\new_[13647]_  | ~\new_[6032]_ );
  assign \new_[12631]_  = (~\new_[13995]_  | ~\new_[5756]_ ) & (~\new_[6724]_  | ~\new_[4501]_ );
  assign \new_[12632]_  = (~\new_[13638]_  | ~\new_[6013]_ ) & (~\new_[14059]_  | ~\new_[3741]_ );
  assign \new_[12633]_  = (~\new_[13821]_  | ~\new_[2502]_ ) & (~\new_[13881]_  | ~\new_[5490]_ );
  assign \new_[12634]_  = (~\new_[5756]_  | ~\new_[14208]_ ) & (~\new_[4501]_  | ~\new_[14081]_ );
  assign \new_[12635]_  = (~\new_[14079]_  | ~\new_[5562]_ ) & (~\new_[13863]_  | ~\new_[2500]_ );
  assign \new_[12636]_  = (~\new_[14218]_  | ~\new_[5491]_ ) & (~\new_[14130]_  | ~\new_[2504]_ );
  assign \new_[12637]_  = ~\new_[3471]_  | ~\new_[3472]_  | ~\new_[3470]_  | ~\new_[3410]_ ;
  assign \new_[12638]_  = (~\new_[14151]_  | ~\new_[2552]_ ) & (~\new_[4970]_  | ~\new_[14057]_ );
  assign \new_[12639]_  = (~\new_[14102]_  | ~\new_[6310]_ ) & (~\new_[13563]_  | ~\new_[3595]_ );
  assign \new_[12640]_  = ~\new_[13040]_ ;
  assign \new_[12641]_  = (~\new_[3686]_  | ~\new_[14073]_ ) & (~\new_[3464]_  | ~\new_[13981]_ );
  assign \new_[12642]_  = (~\new_[3879]_  | ~\new_[13705]_ ) & (~\new_[3787]_  | ~\new_[13506]_ );
  assign \new_[12643]_  = \new_[2096]_  ^ \new_[2090]_ ;
  assign \new_[12644]_  = \new_[13944]_  ^ \new_[13770]_ ;
  assign \new_[12645]_  = \new_[2175]_  ^ \new_[13845]_ ;
  assign \new_[12646]_  = \new_[8702]_  ^ \new_[14061]_ ;
  assign \new_[12647]_  = (~\new_[3938]_  | ~\new_[13555]_ ) & (~\new_[3940]_  | ~\new_[13752]_ );
  assign \new_[12648]_  = \new_[14032]_  ^ \new_[13889]_ ;
  assign \new_[12649]_  = ~u4_u1_dma_ack_clr1_reg;
  assign \new_[12650]_  = ~u4_u0_r5_reg;
  assign \new_[12651]_  = ~\new_[13449]_ ;
  assign \new_[12652]_  = ~\new_[13204]_ ;
  assign \new_[12653]_  = ~u4_u0_dma_ack_clr1_reg;
  assign \new_[12654]_  = u0_tx_ready_reg;
  assign \new_[12655]_  = ~\new_[13017]_ ;
  assign \new_[12656]_  = ~\new_[12969]_ ;
  assign \new_[12657]_  = ~\new_[13202]_ ;
  assign \new_[12658]_  = ~\new_[13253]_ ;
  assign \new_[12659]_  = ~\new_[13033]_ ;
  assign \new_[12660]_  = ~\new_[13041]_ ;
  assign \new_[12661]_  = ~\new_[13206]_ ;
  assign \new_[12662]_  = ~\new_[13066]_ ;
  assign \new_[12663]_  = ~\new_[6368]_  & ~\new_[6367]_ ;
  assign \new_[12664]_  = ~\new_[13208]_ ;
  assign \new_[12665]_  = ~\new_[3638]_  | ~\new_[14108]_ ;
  assign \new_[12666]_  = ~\new_[13034]_ ;
  assign \new_[12667]_  = ~\new_[6563]_  & ~\new_[3342]_ ;
  assign \new_[12668]_  = ~\new_[13001]_ ;
  assign \new_[12669]_  = ~\new_[13025]_ ;
  assign \new_[12670]_  = ~\new_[13173]_ ;
  assign \new_[12671]_  = \new_[13352]_  & \wb_addr_i[4] ;
  assign \new_[12672]_  = ~\new_[13102]_ ;
  assign \new_[12673]_  = ~\new_[6092]_  | ~\new_[14213]_ ;
  assign \new_[12674]_  = ~\new_[13282]_  | ~\new_[6385]_ ;
  assign \new_[12675]_  = ~\new_[12918]_ ;
  assign \new_[12676]_  = \new_[14115]_  ^ \new_[4607]_ ;
  assign \new_[12677]_  = ~\new_[13059]_ ;
  assign \new_[12678]_  = ~\new_[13189]_ ;
  assign \new_[12679]_  = ~\new_[12905]_ ;
  assign \new_[12680]_  = ~\new_[12960]_ ;
  assign \new_[12681]_  = \new_[2454]_  | \new_[12368]_ ;
  assign \new_[12682]_  = ~\new_[13051]_ ;
  assign \new_[12683]_  = ~\new_[13063]_ ;
  assign \new_[12684]_  = ~\new_[13231]_ ;
  assign \new_[12685]_  = ~\new_[13054]_ ;
  assign \new_[12686]_  = ~\new_[6251]_  & ~\new_[4097]_ ;
  assign \new_[12687]_  = ~\new_[5999]_  | ~\new_[3341]_ ;
  assign \new_[12688]_  = \new_[10003]_  | \new_[2611]_ ;
  assign \new_[12689]_  = \new_[13294]_  & \new_[13285]_ ;
  assign \new_[12690]_  = ~\new_[3888]_  | ~\new_[3889]_ ;
  assign \new_[12691]_  = \\u4_utmi_vend_stat_r_reg[6] ;
  assign \new_[12692]_  = ~\new_[6588]_  & (~\new_[13689]_  | ~\new_[6303]_ );
  assign \new_[12693]_  = ~\new_[13188]_ ;
  assign \new_[12694]_  = ~\new_[13171]_ ;
  assign \new_[12695]_  = ~\new_[3875]_  & ~\new_[3671]_ ;
  assign \new_[12696]_  = ~\new_[13058]_ ;
  assign \new_[12697]_  = ~\new_[6004]_  | ~\new_[3510]_ ;
  assign \new_[12698]_  = ~\new_[12939]_ ;
  assign \new_[12699]_  = ~\new_[6009]_  | ~\new_[3806]_ ;
  assign \new_[12700]_  = ~\new_[13311]_  & ~\new_[13288]_ ;
  assign \new_[12701]_  = ~\new_[3428]_  & ~\new_[3313]_ ;
  assign \new_[12702]_  = \new_[6567]_  & \new_[3506]_ ;
  assign \new_[12703]_  = ~\new_[6286]_  & ~\new_[3714]_ ;
  assign \new_[12704]_  = ~\new_[13163]_ ;
  assign \new_[12705]_  = ~\new_[13052]_ ;
  assign \new_[12706]_  = ~\new_[13270]_  & ~\new_[13550]_ ;
  assign \new_[12707]_  = \new_[6287]_  & \new_[3890]_ ;
  assign \new_[12708]_  = ~\new_[13020]_ ;
  assign \new_[12709]_  = ~\new_[6017]_  | ~\new_[13944]_ ;
  assign \new_[12710]_  = ~\new_[13065]_ ;
  assign \new_[12711]_  = ~\new_[13302]_  & ~\new_[13496]_ ;
  assign \new_[12712]_  = ~\new_[12964]_ ;
  assign \new_[12713]_  = ~\new_[14139]_  | ~\new_[13364]_ ;
  assign \new_[12714]_  = ~\new_[3718]_  & ~\new_[3806]_ ;
  assign \new_[12715]_  = ~\new_[13240]_ ;
  assign \new_[12716]_  = ~\new_[12953]_ ;
  assign \new_[12717]_  = ~\new_[13282]_  & ~\new_[13923]_ ;
  assign \new_[12718]_  = ~\wb_addr_i[3]  & ~\wb_addr_i[4] ;
  assign \new_[12719]_  = ~\new_[6091]_  & ~\new_[13746]_ ;
  assign \new_[12720]_  = ~\new_[6733]_  | ~\new_[6602]_ ;
  assign \new_[12721]_  = ~\new_[12943]_ ;
  assign \new_[12722]_  = ~\new_[6365]_  | ~\new_[6366]_ ;
  assign \new_[12723]_  = ~\new_[3713]_  & ~\new_[3718]_ ;
  assign \new_[12724]_  = ~\new_[6716]_  & ~\new_[6020]_ ;
  assign \new_[12725]_  = ~\new_[6274]_  | ~\new_[3509]_ ;
  assign \new_[12726]_  = ~\new_[12926]_ ;
  assign \new_[12727]_  = ~\new_[13222]_ ;
  assign \new_[12728]_  = ~\new_[13970]_  & ~\new_[14185]_ ;
  assign \new_[12729]_  = ~\new_[13100]_ ;
  assign \new_[12730]_  = ~\new_[13000]_ ;
  assign \new_[12731]_  = ~\new_[12994]_ ;
  assign \new_[12732]_  = ~\new_[12197]_ ;
  assign \new_[12733]_  = \new_[4783]_  | \new_[13755]_ ;
  assign \new_[12734]_  = ~\new_[14373]_ ;
  assign \new_[12735]_  = ~\new_[13068]_ ;
  assign \new_[12736]_  = ~\new_[13082]_ ;
  assign \new_[12737]_  = ~\new_[13103]_ ;
  assign \new_[12738]_  = ~\new_[13482]_  & ~\new_[13444]_ ;
  assign \new_[12739]_  = ~\new_[13075]_ ;
  assign \new_[12740]_  = \new_[3508]_  | \new_[3507]_ ;
  assign \new_[12741]_  = ~\new_[13093]_ ;
  assign \new_[12742]_  = ~\new_[13027]_ ;
  assign \new_[12743]_  = (~\new_[13586]_  | ~\new_[2554]_ ) & (~\new_[4966]_  | ~\new_[14218]_ );
  assign \new_[12744]_  = (~\new_[14236]_  | ~\new_[2500]_ ) & (~\new_[14153]_  | ~\new_[5562]_ );
  assign \new_[12745]_  = ~\new_[12965]_ ;
  assign \new_[12746]_  = ~\new_[6200]_  | ~\new_[3626]_ ;
  assign \new_[12747]_  = ~\new_[13274]_  & ~\new_[14213]_ ;
  assign \new_[12748]_  = ~\new_[13101]_ ;
  assign \new_[12749]_  = ~\new_[13109]_ ;
  assign \new_[12750]_  = (~\new_[14157]_  | ~\new_[2551]_ ) & (~\new_[5111]_  | ~\new_[14079]_ );
  assign \new_[12751]_  = (~\new_[13681]_  | ~\new_[2552]_ ) & (~\new_[13742]_  | ~\new_[6697]_ );
  assign \new_[12752]_  = ~\new_[13223]_ ;
  assign \new_[12753]_  = (~\new_[5109]_  | ~\new_[14110]_ ) & (~\new_[5123]_  | ~\new_[13712]_ );
  assign \new_[12754]_  = ~\new_[13243]_ ;
  assign \new_[12755]_  = ~\new_[6019]_  | ~\new_[6105]_ ;
  assign \new_[12756]_  = ~\new_[2452]_  | ~\new_[2042]_ ;
  assign \new_[12757]_  = \new_[13391]_  & \new_[13368]_ ;
  assign \new_[12758]_  = ~\new_[6251]_  | ~\new_[4097]_ ;
  assign \new_[12759]_  = ~\new_[13131]_ ;
  assign \new_[12760]_  = ~\new_[13895]_ ;
  assign \new_[12761]_  = (~\new_[13704]_  | ~\new_[6310]_ ) & (~\new_[14142]_  | ~\new_[3595]_ );
  assign \new_[12762]_  = (~\new_[13611]_  | ~\new_[2554]_ ) & (~\new_[14131]_  | ~\new_[5760]_ );
  assign \new_[12763]_  = ~\new_[13124]_ ;
  assign \new_[12764]_  = (~\new_[13525]_  | ~\new_[6013]_ ) & (~\new_[14104]_  | ~\new_[3741]_ );
  assign \new_[12765]_  = ~\new_[13125]_ ;
  assign \new_[12766]_  = (~\new_[5490]_  | ~\new_[13780]_ ) & (~\new_[14039]_  | ~\new_[2502]_ );
  assign \new_[12767]_  = (~\new_[14038]_  | ~\new_[6011]_ ) & (~\new_[14042]_  | ~\new_[3716]_ );
  assign \new_[12768]_  = (~\new_[13509]_  | ~\new_[5761]_ ) & (~\new_[13579]_  | ~\new_[3739]_ );
  assign \new_[12769]_  = ~\new_[13127]_ ;
  assign \new_[12770]_  = ~\new_[4597]_  | ~\new_[4506]_  | ~\new_[14013]_  | ~\new_[4502]_ ;
  assign \new_[12771]_  = ~\new_[13129]_ ;
  assign \new_[12772]_  = ~\new_[13107]_ ;
  assign \new_[12773]_  = \new_[13286]_  | \new_[13355]_ ;
  assign \new_[12774]_  = ~\new_[2318]_  & ~\new_[2344]_ ;
  assign \new_[12775]_  = ~\new_[13132]_ ;
  assign \new_[12776]_  = ~\new_[3508]_  & ~\new_[13340]_ ;
  assign \new_[12777]_  = ~\new_[14152]_  & (~\new_[10668]_  | ~\new_[13626]_ );
  assign \new_[12778]_  = ~\new_[13136]_ ;
  assign \new_[12779]_  = ~\new_[6232]_  & ~\new_[6319]_ ;
  assign \new_[12780]_  = ~\new_[13456]_  & ~\new_[13267]_ ;
  assign \new_[12781]_  = \new_[13495]_  & \new_[9412]_ ;
  assign \new_[12782]_  = ~\new_[13448]_  | ~\new_[13441]_ ;
  assign \new_[12783]_  = ~\new_[13328]_ ;
  assign \new_[12784]_  = \new_[13356]_  & \new_[8701]_ ;
  assign \new_[12785]_  = ~\new_[13926]_  | ~\new_[13440]_ ;
  assign \new_[12786]_  = ~\new_[6266]_  & ~\new_[3429]_ ;
  assign \new_[12787]_  = ~\new_[3684]_  & ~\new_[3468]_ ;
  assign \new_[12788]_  = ~\new_[3340]_  & ~\new_[3339]_ ;
  assign \new_[12789]_  = \new_[6196]_  & \new_[4197]_ ;
  assign \new_[12790]_  = ~u4_u2_dma_ack_clr1_reg;
  assign \new_[12791]_  = \new_[13735]_  ^ \new_[10715]_ ;
  assign \new_[12792]_  = ~\new_[13154]_ ;
  assign \new_[12793]_  = ~\new_[6266]_  | ~\new_[3429]_ ;
  assign \new_[12794]_  = ~\new_[13165]_ ;
  assign \new_[12795]_  = (~\new_[13949]_  | ~\new_[6011]_ ) & (~\new_[14109]_  | ~\new_[3716]_ );
  assign \new_[12796]_  = ~\new_[14582]_ ;
  assign \new_[12797]_  = ~\new_[4777]_  | ~\new_[8959]_ ;
  assign \new_[12798]_  = ~\new_[12941]_ ;
  assign n8860 = ~\new_[2802]_  & ~n9145;
  assign \new_[12800]_  = ~\new_[2193]_  & ~\new_[13320]_ ;
  assign \new_[12801]_  = ~\new_[13104]_ ;
  assign \new_[12802]_  = ~\new_[13156]_ ;
  assign \new_[12803]_  = ~\new_[13556]_  & (~\new_[10653]_  | ~\new_[13971]_ );
  assign \new_[12804]_  = ~\new_[13162]_ ;
  assign \new_[12805]_  = ~\new_[4814]_  | ~\new_[13861]_ ;
  assign \new_[12806]_  = ~\new_[13341]_  | ~\new_[13313]_ ;
  assign \new_[12807]_  = ~\new_[13170]_ ;
  assign \new_[12808]_  = (~\new_[14099]_  | ~\new_[2553]_ ) & (~\new_[13780]_  | ~\new_[5112]_ );
  assign \new_[12809]_  = \new_[2876]_  | \new_[14508]_ ;
  assign \new_[12810]_  = ~\new_[6370]_  & (~\new_[13876]_  | ~\new_[6371]_ );
  assign \new_[12811]_  = ~\new_[13047]_ ;
  assign \new_[12812]_  = u1_u3_uc_dpd_set_reg;
  assign \new_[12813]_  = ~\new_[13039]_ ;
  assign \new_[12814]_  = ~\new_[12996]_ ;
  assign \new_[12815]_  = ~\new_[13177]_ ;
  assign \new_[12816]_  = ~\new_[13433]_ ;
  assign \new_[12817]_  = ~\new_[13164]_ ;
  assign \new_[12818]_  = ~\new_[13183]_ ;
  assign \new_[12819]_  = ~\new_[12985]_ ;
  assign \new_[12820]_  = ~\new_[13191]_ ;
  assign \new_[12821]_  = \new_[4608]_  & \new_[4841]_ ;
  assign \new_[12822]_  = ~\new_[13185]_ ;
  assign \new_[12823]_  = ~\new_[13235]_ ;
  assign \new_[12824]_  = ~\new_[6383]_  | ~\new_[14254]_ ;
  assign \new_[12825]_  = ~\new_[13378]_  & ~\new_[13445]_ ;
  assign \new_[12826]_  = ~\new_[13087]_ ;
  assign \new_[12827]_  = ~\new_[4783]_  | ~\new_[13755]_ ;
  assign \new_[12828]_  = ~\new_[6346]_  & (~\new_[13814]_  | ~\new_[6347]_ );
  assign \new_[12829]_  = (~\new_[5617]_  | ~\new_[13763]_ ) & (~\new_[3878]_  | ~\new_[13702]_ );
  assign \new_[12830]_  = ~\new_[13194]_ ;
  assign \new_[12831]_  = ~\new_[12952]_ ;
  assign \new_[12832]_  = ~\new_[12932]_ ;
  assign \new_[12833]_  = ~u4_u3_dma_ack_clr1_reg;
  assign \new_[12834]_  = ~\new_[13172]_ ;
  assign \new_[12835]_  = ~u4_u2_r5_reg;
  assign \new_[12836]_  = ~\new_[13201]_ ;
  assign \new_[12837]_  = ~\new_[13203]_ ;
  assign \new_[12838]_  = u1_u3_uc_bsel_set_reg;
  assign \new_[12839]_  = (~\new_[13564]_  | ~\new_[2501]_ ) & (~\new_[14063]_  | ~\new_[5489]_ );
  assign \new_[12840]_  = ~u4_u3_r5_reg;
  assign \new_[12841]_  = ~\new_[13024]_ ;
  assign \new_[12842]_  = ~\new_[12197]_ ;
  assign \new_[12843]_  = (~\new_[13849]_  | ~\new_[2553]_ ) & (~\new_[13925]_  | ~\new_[5499]_ );
  assign \new_[12844]_  = ~\new_[12924]_ ;
  assign \new_[12845]_  = ~\new_[6280]_  & ~\new_[6716]_ ;
  assign \new_[12846]_  = ~\new_[13453]_ ;
  assign \new_[12847]_  = ~\new_[6009]_  & ~\new_[3806]_ ;
  assign \new_[12848]_  = \\u4_utmi_vend_stat_r_reg[3] ;
  assign \new_[12849]_  = ~\new_[13162]_ ;
  assign \new_[12850]_  = ~\new_[6286]_  | ~\new_[3714]_ ;
  assign \new_[12851]_  = ~\new_[6274]_  & ~\new_[3509]_ ;
  assign susp_o = susp_o_reg;
  assign \new_[12853]_  = ~\new_[13227]_ ;
  assign \new_[12854]_  = ~\new_[12946]_ ;
  assign \new_[12855]_  = ~\new_[12945]_ ;
  assign \new_[12856]_  = ~\new_[6200]_  & ~\new_[3626]_ ;
  assign \new_[12857]_  = ~\new_[13291]_  & ~\new_[13270]_ ;
  assign \new_[12858]_  = ~\new_[13049]_ ;
  assign \new_[12859]_  = ~\new_[13151]_ ;
  assign \new_[12860]_  = ~\new_[13457]_  & ~\new_[7206]_ ;
  assign \new_[12861]_  = ~\new_[13214]_ ;
  assign \new_[12862]_  = ~\\u4_u0_buf0_orig_m3_reg[0] ;
  assign \new_[12863]_  = ~\new_[13233]_ ;
  assign \new_[12864]_  = ~\new_[13212]_ ;
  assign \new_[12865]_  = ~\new_[13649]_  | ~\new_[13372]_ ;
  assign \new_[12866]_  = ~\new_[13086]_ ;
  assign \new_[12867]_  = (~\new_[14232]_  | ~\new_[2504]_ ) & (~\new_[14231]_  | ~\new_[5491]_ );
  assign \new_[12868]_  = ~\new_[13275]_  & ~\new_[13928]_ ;
  assign \new_[12869]_  = ~\\u4_u2_buf0_orig_m3_reg[0] ;
  assign \new_[12870]_  = ~\new_[13349]_ ;
  assign \new_[12871]_  = ~\new_[13239]_ ;
  assign \new_[12872]_  = \new_[13331]_  & \new_[13399]_ ;
  assign \new_[12873]_  = ~\new_[6004]_  & ~\new_[3510]_ ;
  assign \new_[12874]_  = ~\\u4_u3_buf0_orig_m3_reg[0] ;
  assign \new_[12875]_  = \\u0_u0_idle_cnt1_next_reg[0] ;
  assign \new_[12876]_  = \new_[9442]_  ^ \new_[14219]_ ;
  assign \new_[12877]_  = ~\new_[13098]_ ;
  assign \new_[12878]_  = ~\new_[13073]_ ;
  assign \new_[12879]_  = ~\new_[13139]_ ;
  assign \new_[12880]_  = ~\new_[12954]_ ;
  assign \new_[12881]_  = ~\new_[4098]_  & ~\new_[4237]_ ;
  assign \new_[12882]_  = ~\new_[2874]_  | ~\new_[2836]_ ;
  assign \new_[12883]_  = ~\new_[13018]_ ;
  assign \new_[12884]_  = \new_[6003]_  & \new_[3507]_ ;
  assign \new_[12885]_  = \new_[6003]_  ^ \new_[3507]_ ;
  assign \new_[12886]_  = \new_[6250]_  & \new_[4098]_ ;
  assign \new_[12887]_  = \new_[6250]_  ^ \new_[4098]_ ;
  assign \new_[12888]_  = \new_[2717]_  & \new_[2637]_ ;
  assign \new_[12889]_  = \new_[2717]_  ^ \new_[2637]_ ;
  assign \new_[12890]_  = \new_[3172]_  & \new_[2982]_ ;
  assign \new_[12891]_  = \new_[3172]_  ^ \new_[2982]_ ;
  assign \new_[12892]_  = \new_[4779]_  & \new_[4666]_ ;
  assign n8865 = \new_[4779]_  ^ \new_[4666]_ ;
  assign \new_[12894]_  = \new_[6008]_  & \new_[3718]_ ;
  assign \new_[12895]_  = \new_[6008]_  ^ \new_[3718]_ ;
  assign \new_[12896]_  = \new_[5998]_  & \new_[3339]_ ;
  assign \new_[12897]_  = \new_[5998]_  ^ \new_[3339]_ ;
  assign \new_[12898]_  = \new_[3035]_  & \new_[3036]_ ;
  assign \new_[12899]_  = \new_[3035]_  ^ \new_[3036]_ ;
  assign \new_[12900]_  = \new_[3465]_  & \new_[3470]_ ;
  assign \new_[12901]_  = \new_[3465]_  ^ \new_[3470]_ ;
  assign \new_[12902]_  = ~\new_[13788]_  & ~\new_[3715]_ ;
  assign \new_[12903]_  = \new_[4765]_  ^ \new_[2175]_ ;
  assign \new_[12904]_  = ~\new_[14149]_  | ~\new_[3506]_ ;
  assign \new_[12905]_  = \new_[14001]_  & \new_[3316]_ ;
  assign \new_[12906]_  = ~\new_[13752]_  | ~\new_[4289]_ ;
  assign \VControl_pad_o[3]  = \\u4_utmi_vend_ctrl_reg[3] ;
  assign \new_[12908]_  = ~\new_[3940]_  | ~\new_[13555]_ ;
  assign \new_[12909]_  = ~\new_[13897]_  | ~\new_[3510]_ ;
  assign \new_[12910]_  = ~\new_[6593]_  & ~\new_[14045]_ ;
  assign \new_[12911]_  = ~\new_[13492]_ ;
  assign \new_[12912]_  = ~\new_[13584]_  | ~\new_[3712]_ ;
  assign \new_[12913]_  = ~\new_[2869]_  | ~\new_[14508]_ ;
  assign \new_[12914]_  = ~\new_[13431]_ ;
  assign VControl_Load_pad_o = u4_utmi_vend_wr_reg;
  assign \new_[12916]_  = ~\new_[13446]_ ;
  assign \VControl_pad_o[0]  = \\u4_utmi_vend_ctrl_reg[0] ;
  assign \new_[12918]_  = ~\new_[6690]_  | ~\new_[13798]_ ;
  assign \new_[12919]_  = ~\new_[13272]_ ;
  assign \new_[12920]_  = ~\new_[4504]_  & ~\new_[13663]_ ;
  assign \new_[12921]_  = ~\new_[13268]_ ;
  assign \new_[12922]_  = \new_[13552]_  & \new_[3480]_ ;
  assign \new_[12923]_  = ~\new_[6272]_  & ~\new_[13816]_ ;
  assign \new_[12924]_  = ~\new_[13517]_  | ~\new_[3429]_ ;
  assign \new_[12925]_  = ~\new_[13793]_  & ~\new_[4074]_ ;
  assign \new_[12926]_  = ~\new_[13656]_  | ~\new_[4288]_ ;
  assign \new_[12927]_  = ~\new_[14153]_  | ~\new_[5111]_ ;
  assign \new_[12928]_  = \new_[4510]_  ^ \new_[4511]_ ;
  assign \new_[12929]_  = \new_[14118]_  & \new_[14084]_ ;
  assign n8885 = usb_vbus_pad_i | \new_[12368]_ ;
  assign \new_[12931]_  = \new_[4502]_  ^ \new_[4505]_ ;
  assign \new_[12932]_  = ~\new_[14790]_  | ~\new_[13861]_ ;
  assign \new_[12933]_  = ~\new_[13412]_ ;
  assign \new_[12934]_  = ~\new_[14111]_  & ~\new_[13766]_ ;
  assign \new_[12935]_  = \new_[13914]_  | \new_[3505]_ ;
  assign \new_[12936]_  = ~\new_[13875]_  & ~\new_[3482]_ ;
  assign \new_[12937]_  = ~\new_[13675]_  & ~\new_[4197]_ ;
  assign \new_[12938]_  = \new_[13552]_  | \new_[3480]_ ;
  assign \new_[12939]_  = \new_[13718]_  | \new_[3478]_ ;
  assign \new_[12940]_  = \new_[13621]_  & \new_[3888]_ ;
  assign \new_[12941]_  = ~\new_[13740]_  & ~\new_[4792]_ ;
  assign \new_[12942]_  = ~\new_[14063]_  | ~\new_[4970]_ ;
  assign \new_[12943]_  = \new_[13649]_  & \new_[4073]_ ;
  assign \new_[12944]_  = ~\new_[6690]_  & ~\new_[13798]_ ;
  assign \new_[12945]_  = \new_[13779]_  | \new_[3428]_ ;
  assign \new_[12946]_  = ~\new_[13675]_  | ~\new_[4197]_ ;
  assign \new_[12947]_  = ~\new_[13366]_ ;
  assign \new_[12948]_  = ~\new_[13962]_  | ~\new_[13747]_ ;
  assign \new_[12949]_  = ~\new_[7206]_  & ~\new_[4290]_ ;
  assign \new_[12950]_  = ~\new_[13342]_ ;
  assign \new_[12951]_  = ~\new_[13391]_ ;
  assign \new_[12952]_  = ~\\u1_u2_rx_data_st_r_reg[4] ;
  assign \new_[12953]_  = \new_[13882]_  & \new_[13744]_ ;
  assign \new_[12954]_  = ~\new_[6255]_  & ~\new_[13689]_ ;
  assign \new_[12955]_  = ~\new_[13506]_  & ~\new_[3883]_ ;
  assign \new_[12956]_  = ~\new_[13978]_  & ~\new_[14205]_ ;
  assign \VControl_pad_o[2]  = \\u4_utmi_vend_ctrl_reg[2] ;
  assign \new_[12958]_  = ~\new_[13881]_  | ~\new_[5112]_ ;
  assign \new_[12959]_  = ~n9010 | ~\new_[3339]_ ;
  assign \new_[12960]_  = \new_[4790]_  | \new_[13692]_ ;
  assign \new_[12961]_  = ~\new_[14265]_  | ~\new_[5760]_ ;
  assign \new_[12962]_  = ~\new_[13399]_ ;
  assign \new_[12963]_  = ~\new_[13306]_ ;
  assign \new_[12964]_  = ~\new_[13754]_  | ~\new_[14052]_ ;
  assign \new_[12965]_  = \new_[13735]_  | \new_[13799]_ ;
  assign \new_[12966]_  = ~\new_[13437]_ ;
  assign \new_[12967]_  = ~\new_[14342]_  | ~\new_[14348]_ ;
  assign \new_[12968]_  = ~\new_[13747]_  | ~\new_[4097]_ ;
  assign \new_[12969]_  = ~\new_[6264]_  | ~\new_[14188]_ ;
  assign \new_[12970]_  = ~\new_[13427]_ ;
  assign \new_[12971]_  = \new_[4552]_  ^ \new_[4505]_ ;
  assign \new_[12972]_  = ~\new_[13601]_  | ~\new_[13508]_ ;
  assign \new_[12973]_  = ~\new_[13278]_ ;
  assign \new_[12974]_  = ~\new_[13276]_ ;
  assign \new_[12975]_  = ~\new_[13397]_ ;
  assign \new_[12976]_  = ~\new_[13815]_  | ~\new_[13932]_ ;
  assign \new_[12977]_  = ~\new_[13924]_  | ~\new_[3882]_ ;
  assign \new_[12978]_  = ~\new_[2344]_  & ~\new_[2346]_ ;
  assign \new_[12979]_  = ~\new_[13571]_  & ~\new_[4096]_ ;
  assign \new_[12980]_  = ~\new_[13915]_  & ~\new_[3806]_ ;
  assign \new_[12981]_  = ~\new_[13337]_ ;
  assign \new_[12982]_  = ~\new_[6470]_  | ~\new_[13969]_ ;
  assign \new_[12983]_  = ~\new_[13455]_ ;
  assign \new_[12984]_  = ~\new_[13989]_  | ~\new_[3714]_ ;
  assign \new_[12985]_  = \new_[13913]_  | \new_[3815]_ ;
  assign \new_[12986]_  = ~\new_[13517]_  & ~\new_[3429]_ ;
  assign \new_[12987]_  = ~\new_[13365]_ ;
  assign \new_[12988]_  = ~\new_[13614]_  | ~\new_[6032]_ ;
  assign \new_[12989]_  = ~\new_[13482]_ ;
  assign \new_[12990]_  = ~\new_[6252]_  | ~\new_[13623]_ ;
  assign \new_[12991]_  = \new_[13666]_  | \new_[13819]_ ;
  assign \new_[12992]_  = ~\new_[13891]_  | ~\new_[3340]_ ;
  assign \new_[12993]_  = ~\new_[2373]_  & ~\new_[13532]_ ;
  assign \new_[12994]_  = \new_[13751]_  | \new_[4291]_ ;
  assign \new_[12995]_  = ~n9015 | ~\new_[3718]_ ;
  assign \new_[12996]_  = \new_[13914]_  & \new_[3505]_ ;
  assign \new_[12997]_  = \new_[13926]_  | \new_[3693]_ ;
  assign \new_[12998]_  = ~\new_[13962]_  & ~\new_[3997]_ ;
  assign \new_[12999]_  = ~\new_[13602]_  | ~\new_[6697]_ ;
  assign \new_[13000]_  = ~\new_[13613]_  | ~\new_[4237]_ ;
  assign \new_[13001]_  = ~\new_[6284]_  | ~\new_[13635]_ ;
  assign \new_[13002]_  = \new_[13585]_  & \new_[14187]_ ;
  assign \new_[13003]_  = ~\new_[6557]_  | ~\new_[3478]_ ;
  assign \new_[13004]_  = ~\new_[13571]_  | ~\new_[4096]_ ;
  assign \new_[13005]_  = ~\new_[13584]_  & ~\new_[3712]_ ;
  assign \new_[13006]_  = ~\new_[5998]_  | ~\new_[13262]_ ;
  assign \new_[13007]_  = ~\new_[13643]_  & ~\new_[3477]_ ;
  assign \new_[13008]_  = ~\new_[13548]_  & ~\new_[3689]_ ;
  assign \new_[13009]_  = ~\new_[6010]_  | ~\new_[13876]_ ;
  assign \new_[13010]_  = ~\new_[3481]_  | ~\new_[13548]_ ;
  assign \new_[13011]_  = ~\new_[13351]_ ;
  assign \new_[13012]_  = ~\new_[13359]_ ;
  assign \new_[13013]_  = ~\new_[13676]_  | ~\new_[14086]_ ;
  assign \new_[13014]_  = ~\new_[6809]_  & ~\new_[13865]_ ;
  assign \new_[13015]_  = ~\new_[13872]_  & ~\new_[3508]_ ;
  assign \new_[13016]_  = ~\new_[13540]_  & ~\new_[3713]_ ;
  assign \new_[13017]_  = ~\new_[13903]_  | ~\new_[3692]_ ;
  assign \new_[13018]_  = ~\new_[13394]_ ;
  assign \new_[13019]_  = ~\new_[13613]_  & ~\new_[4237]_ ;
  assign \new_[13020]_  = ~\new_[13900]_  | ~\new_[13698]_ ;
  assign \new_[13021]_  = ~\new_[13360]_ ;
  assign \new_[13022]_  = (~\new_[6609]_  | ~\new_[2573]_ ) & (~\new_[6722]_  | ~\new_[4778]_ );
  assign \new_[13023]_  = \new_[13980]_  | \new_[3788]_ ;
  assign \new_[13024]_  = \new_[13624]_  | \new_[3684]_ ;
  assign \new_[13025]_  = ~\new_[13872]_  | ~\new_[3508]_ ;
  assign \new_[13026]_  = \new_[4500]_  ^ \new_[4505]_ ;
  assign \new_[13027]_  = ~\new_[13980]_  | ~\new_[3788]_ ;
  assign \new_[13028]_  = ~\new_[6005]_  & ~\new_[13814]_ ;
  assign \new_[13029]_  = ~\new_[13643]_  | ~\new_[3477]_ ;
  assign \new_[13030]_  = ~\new_[2524]_  | ~\new_[13595]_ ;
  assign \new_[13031]_  = ~\new_[6016]_  | ~\new_[13633]_ ;
  assign \new_[13032]_  = ~\new_[6567]_  | ~\new_[13490]_ ;
  assign \new_[13033]_  = ~\new_[13904]_  & ~\new_[4347]_ ;
  assign \new_[13034]_  = ~\new_[13793]_  | ~\new_[4074]_ ;
  assign \new_[13035]_  = ~\new_[13981]_  & ~\new_[3688]_ ;
  assign \new_[13036]_  = ~\new_[3309]_  | ~\new_[13941]_ ;
  assign \new_[13037]_  = ~\new_[13309]_ ;
  assign \new_[13038]_  = ~\new_[3693]_  | ~\new_[13913]_ ;
  assign \new_[13039]_  = ~\new_[13915]_  | ~\new_[3806]_ ;
  assign \new_[13040]_  = ~\new_[13985]_  | ~\new_[6545]_ ;
  assign \new_[13041]_  = \new_[14139]_  & \new_[3481]_ ;
  assign \new_[13042]_  = ~\new_[6275]_  | ~\new_[13405]_ ;
  assign \new_[13043]_  = \new_[14221]_  | \new_[3691]_ ;
  assign \new_[13044]_  = ~\new_[14238]_  & ~\new_[6543]_ ;
  assign \new_[13045]_  = ~\new_[14043]_  & ~\new_[3342]_ ;
  assign \new_[13046]_  = ~\new_[13981]_  | ~\new_[3688]_ ;
  assign \new_[13047]_  = ~\new_[13352]_ ;
  assign \new_[13048]_  = ~\new_[14108]_  & ~\new_[3626]_ ;
  assign \new_[13049]_  = \new_[14015]_  & \new_[3504]_ ;
  assign \new_[13050]_  = ~\new_[6255]_  | ~\new_[13689]_ ;
  assign \new_[13051]_  = ~\new_[14052]_  | ~\new_[4236]_ ;
  assign \new_[13052]_  = ~\new_[14069]_  | ~\new_[3884]_ ;
  assign \new_[13053]_  = ~\new_[13891]_  & ~\new_[3340]_ ;
  assign \new_[13054]_  = \new_[14069]_  | \new_[3884]_ ;
  assign \new_[13055]_  = ~\new_[13340]_ ;
  assign \new_[13056]_  = ~\new_[6247]_  & ~\new_[14005]_ ;
  assign \new_[13057]_  = ~\new_[6003]_  | ~\new_[13422]_ ;
  assign \new_[13058]_  = ~\new_[13933]_  | ~\new_[14226]_ ;
  assign \new_[13059]_  = ~\new_[6743]_  | ~\new_[13733]_ ;
  assign \new_[13060]_  = ~\new_[13318]_ ;
  assign \new_[13061]_  = \new_[4372]_  ^ \new_[4504]_ ;
  assign \new_[13062]_  = ~\new_[13488]_ ;
  assign \new_[13063]_  = ~\new_[13945]_  | ~\new_[3317]_ ;
  assign \new_[13064]_  = \new_[14139]_  | \new_[3481]_ ;
  assign \new_[13065]_  = \new_[3342]_  | \new_[3341]_ ;
  assign \new_[13066]_  = ~\new_[14043]_  | ~\new_[3342]_ ;
  assign \new_[13067]_  = ~n9145 | ~\new_[13999]_ ;
  assign \new_[13068]_  = ~\new_[14000]_  | ~\new_[13620]_ ;
  assign \new_[13069]_  = ~\new_[13583]_  & ~\new_[13828]_ ;
  assign \new_[13070]_  = \new_[3997]_  | \new_[4097]_ ;
  assign \new_[13071]_  = ~\new_[14103]_  | ~\new_[5499]_ ;
  assign \new_[13072]_  = ~n9145 | ~\new_[13502]_ ;
  assign \new_[13073]_  = ~\new_[6255]_  | ~\new_[4347]_ ;
  assign \new_[13074]_  = ~\new_[6008]_  | ~\new_[13371]_ ;
  assign \new_[13075]_  = ~\new_[6287]_  | ~\new_[13322]_ ;
  assign \new_[13076]_  = \new_[14015]_  | \new_[3504]_ ;
  assign \new_[13077]_  = ~\new_[13903]_  & ~\new_[3692]_ ;
  assign \new_[13078]_  = ~\new_[13752]_  & ~\new_[4289]_ ;
  assign \new_[13079]_  = ~\new_[13988]_  | ~\new_[6015]_ ;
  assign \new_[13080]_  = ~\new_[13627]_  | ~\new_[6258]_ ;
  assign \new_[13081]_  = ~\new_[13258]_ ;
  assign \new_[13082]_  = ~\new_[13788]_  | ~\new_[3715]_ ;
  assign \new_[13083]_  = ~\new_[2876]_  | ~\new_[14508]_ ;
  assign \new_[13084]_  = ~\new_[4777]_  | ~\new_[13901]_ ;
  assign \new_[13085]_  = ~\new_[13679]_  | ~\new_[13755]_ ;
  assign \new_[13086]_  = ~\new_[6809]_  | ~\new_[13865]_ ;
  assign \new_[13087]_  = ~\new_[13540]_  | ~\new_[3713]_ ;
  assign \new_[13088]_  = ~\new_[6544]_  | ~\new_[13912]_ ;
  assign \new_[13089]_  = \new_[13514]_  & \new_[13501]_ ;
  assign \new_[13090]_  = \new_[13629]_  | \new_[4293]_ ;
  assign \new_[13091]_  = ~\new_[13711]_  | ~\new_[13370]_ ;
  assign \new_[13092]_  = ~\new_[14508]_ ;
  assign \new_[13093]_  = \new_[13631]_  & \new_[3711]_ ;
  assign \new_[13094]_  = ~\new_[13718]_  | ~\new_[3478]_ ;
  assign \new_[13095]_  = ~\new_[6196]_  | ~\new_[13374]_ ;
  assign \new_[13096]_  = ~\new_[4615]_ ;
  assign \new_[13097]_  = \new_[13649]_  | \new_[4073]_ ;
  assign \new_[13098]_  = ~\new_[14078]_  | ~\new_[13370]_ ;
  assign \new_[13099]_  = ~\new_[2372]_  & ~\new_[13813]_ ;
  assign \new_[13100]_  = ~\new_[3282]_  | ~\new_[13825]_ ;
  assign \new_[13101]_  = ~\new_[14197]_  | ~\new_[3890]_ ;
  assign \new_[13102]_  = \new_[13751]_  & \new_[4291]_ ;
  assign \new_[13103]_  = ~\new_[13875]_  | ~\new_[3482]_ ;
  assign \new_[13104]_  = ~\new_[13761]_  & ~\new_[3341]_ ;
  assign \new_[13105]_  = ~\new_[13761]_  | ~\new_[3341]_ ;
  assign \new_[13106]_  = ~\new_[6005]_  | ~\new_[13814]_ ;
  assign \new_[13107]_  = ~\new_[6010]_  & ~\new_[13876]_ ;
  assign \new_[13108]_  = ~\new_[13256]_ ;
  assign \new_[13109]_  = ~\new_[13779]_  | ~\new_[3428]_ ;
  assign \new_[13110]_  = ~\new_[13852]_  | ~\new_[13748]_ ;
  assign \new_[13111]_  = ~\new_[4683]_  & ~\new_[14261]_ ;
  assign \new_[13112]_  = ~\new_[13384]_ ;
  assign \new_[13113]_  = ~\new_[13380]_ ;
  assign \new_[13114]_  = ~\new_[13387]_ ;
  assign \new_[13115]_  = ~\new_[13627]_  & ~\new_[6258]_ ;
  assign \new_[13116]_  = ~\wb_addr_i[2]  | ~\new_[13695]_ ;
  assign \new_[13117]_  = \new_[2869]_  | \new_[14508]_ ;
  assign \new_[13118]_  = \new_[4852]_  | \new_[4615]_ ;
  assign \new_[13119]_  = ~n8890 | ~\new_[3507]_ ;
  assign \new_[13120]_  = ~\new_[13477]_ ;
  assign \new_[13121]_  = ~\new_[13606]_  & ~\new_[3012]_ ;
  assign \new_[13122]_  = ~\new_[4709]_  | ~\new_[4818]_ ;
  assign \new_[13123]_  = ~\new_[3787]_  | ~\new_[13705]_ ;
  assign \new_[13124]_  = ~\new_[14238]_  | ~\new_[6543]_ ;
  assign \new_[13125]_  = ~\new_[3283]_  | ~\new_[14052]_ ;
  assign \new_[13126]_  = ~\new_[13331]_ ;
  assign \new_[13127]_  = \new_[13926]_  & \new_[3693]_ ;
  assign \new_[13128]_  = ~\wb_addr_i[5]  & ~\new_[13974]_ ;
  assign \new_[13129]_  = \new_[13695]_  | \wb_addr_i[5] ;
  assign \new_[13130]_  = ~\new_[6005]_  | ~\new_[3689]_ ;
  assign \new_[13131]_  = ~\new_[13962]_  | ~\new_[3997]_ ;
  assign \new_[13132]_  = ~\\u1_u2_rx_data_st_r_reg[7] ;
  assign \new_[13133]_  = \new_[13621]_  | \new_[3888]_ ;
  assign \new_[13134]_  = ~\new_[13301]_ ;
  assign \new_[13135]_  = ~\new_[14348]_ ;
  assign \new_[13136]_  = ~\new_[13442]_ ;
  assign \new_[13137]_  = ~\new_[13403]_ ;
  assign \new_[13138]_  = ~\new_[14118]_ ;
  assign \new_[13139]_  = ~\new_[2096]_  | ~\new_[2092]_  | ~\new_[2090]_ ;
  assign \new_[13140]_  = \new_[4774]_  & \new_[13664]_ ;
  assign \new_[13141]_  = ~\new_[13905]_  | ~\new_[3509]_ ;
  assign \new_[13142]_  = ~n9020 | ~\new_[4098]_ ;
  assign \new_[13143]_  = ~\new_[3316]_  | ~\new_[13718]_ ;
  assign \new_[13144]_  = ~\new_[13297]_ ;
  assign \new_[13145]_  = ~\new_[14149]_  & ~\new_[3506]_ ;
  assign phy_rst_pad_o = ~\new_[14503]_ ;
  assign \new_[13147]_  = \new_[13548]_  & \new_[3689]_ ;
  assign \new_[13148]_  = ~\new_[3882]_  | ~\new_[13915]_ ;
  assign \new_[13149]_  = ~\new_[13768]_  | ~\new_[13370]_ ;
  assign \new_[13150]_  = ~\new_[2870]_  | ~\new_[2871]_ ;
  assign \new_[13151]_  = ~\new_[13370]_  | ~\new_[13884]_ ;
  assign \new_[13152]_  = ~\new_[13308]_ ;
  assign \new_[13153]_  = ~\new_[13307]_ ;
  assign \new_[13154]_  = ~\new_[13989]_  & ~\new_[3714]_ ;
  assign \new_[13155]_  = ~\new_[5486]_ ;
  assign \new_[13156]_  = ~\\u1_u2_rx_data_st_r_reg[0] ;
  assign \new_[13157]_  = \new_[13913]_  & \new_[3815]_ ;
  assign \new_[13158]_  = ~\new_[13259]_ ;
  assign \new_[13159]_  = ~\new_[13785]_  | ~\new_[13523]_ ;
  assign \new_[13160]_  = ~\new_[13255]_ ;
  assign \new_[13161]_  = ~\new_[6264]_  & ~\new_[14188]_ ;
  assign \new_[13162]_  = ~\new_[12368]_ ;
  assign \new_[13163]_  = ~\new_[14161]_  & ~\new_[14254]_ ;
  assign \new_[13164]_  = ~\\u1_u2_rx_data_st_r_reg[2] ;
  assign \new_[13165]_  = ~\new_[12368]_ ;
  assign \new_[13166]_  = ~\new_[13418]_ ;
  assign \new_[13167]_  = \wb_addr_i[2]  | \new_[13695]_ ;
  assign \new_[13168]_  = \new_[14052]_  | \new_[4236]_ ;
  assign \new_[13169]_  = \new_[4926]_  ^ \new_[4765]_ ;
  assign \new_[13170]_  = ~\\u1_u2_rx_data_st_r_reg[3] ;
  assign \new_[13171]_  = ~\new_[13691]_  | ~\new_[13598]_ ;
  assign \new_[13172]_  = ~\new_[13947]_  | ~\new_[13825]_ ;
  assign \new_[13173]_  = ~\new_[13747]_  & ~\new_[4097]_ ;
  assign \new_[13174]_  = ~\new_[3308]_  | ~\new_[13866]_ ;
  assign \VControl_pad_o[1]  = \\u4_utmi_vend_ctrl_reg[1] ;
  assign n8880 = ~\new_[13345]_ ;
  assign \new_[13177]_  = ~\new_[13905]_  & ~\new_[3509]_ ;
  assign \new_[13178]_  = \new_[2090]_  | \new_[13930]_ ;
  assign \new_[13179]_  = ~\new_[13321]_ ;
  assign \new_[13180]_  = ~\new_[13945]_  & ~\new_[3317]_ ;
  assign \new_[13181]_  = ~\new_[13749]_  | ~\new_[14204]_ ;
  assign \new_[13182]_  = ~\new_[6250]_  | ~\new_[13393]_ ;
  assign \new_[13183]_  = ~\new_[3476]_  | ~\new_[13517]_ ;
  assign \new_[13184]_  = ~\new_[13400]_ ;
  assign \new_[13185]_  = ~\\u1_u2_rx_data_st_r_reg[1] ;
  assign \new_[13186]_  = \new_[4552]_  ^ \new_[4504]_ ;
  assign \new_[13187]_  = ~\new_[2479]_  & ~\new_[14106]_ ;
  assign \new_[13188]_  = \new_[3715]_  | \new_[3714]_ ;
  assign \new_[13189]_  = ~\new_[13320]_ ;
  assign \new_[13190]_  = ~\new_[13491]_ ;
  assign \new_[13191]_  = ~\new_[4288]_  | ~\new_[13613]_ ;
  assign \new_[13192]_  = ~\new_[13343]_ ;
  assign \new_[13193]_  = ~\new_[13341]_ ;
  assign \new_[13194]_  = ~\new_[6247]_  | ~\new_[14005]_ ;
  assign n8625 = ~\new_[13443]_ ;
  assign \new_[13196]_  = ~\new_[13624]_  | ~\new_[3684]_ ;
  assign \new_[13197]_  = ~\new_[13441]_ ;
  assign \new_[13198]_  = ~\new_[14197]_  | ~\new_[13915]_ ;
  assign \new_[13199]_  = ~\new_[13897]_  & ~\new_[3510]_ ;
  assign \new_[13200]_  = ~\new_[13673]_  | ~\new_[13616]_ ;
  assign \new_[13201]_  = (~\new_[6723]_  | ~\new_[5109]_ ) & (~\new_[6610]_  | ~\new_[5123]_ );
  assign \new_[13202]_  = ~\new_[6544]_  & ~\new_[13912]_ ;
  assign \new_[13203]_  = ~\\u1_u2_rx_data_st_r_reg[5] ;
  assign \new_[13204]_  = ~\\u1_u2_rx_data_st_r_reg[6] ;
  assign \new_[13205]_  = ~\new_[12437]_ ;
  assign \new_[13206]_  = ~\new_[13506]_  | ~\new_[3883]_ ;
  assign \new_[13207]_  = \new_[14221]_  & \new_[3691]_ ;
  assign \new_[13208]_  = \new_[13629]_  & \new_[4293]_ ;
  assign \new_[13209]_  = ~\new_[13375]_ ;
  assign n8890 = ~\new_[6341]_ ;
  assign \new_[13211]_  = ~\new_[13723]_  | ~\new_[14129]_ ;
  assign \new_[13212]_  = ~\new_[14108]_  | ~\new_[3626]_ ;
  assign \new_[13213]_  = \new_[13631]_  | \new_[3711]_ ;
  assign \new_[13214]_  = ~\new_[13664]_  | ~\new_[13710]_ ;
  assign \new_[13215]_  = ~\new_[14197]_  & ~\new_[3890]_ ;
  assign \new_[13216]_  = ~\new_[6010]_  | ~\new_[3815]_ ;
  assign \new_[13217]_  = ~\new_[6557]_  | ~\new_[13893]_ ;
  assign \new_[13218]_  = \new_[14216]_  & \new_[13645]_ ;
  assign \new_[13219]_  = \new_[3025]_  & \new_[14211]_ ;
  assign \new_[13220]_  = ~\new_[4695]_  | ~\new_[4815]_ ;
  assign \new_[13221]_  = ~\new_[13466]_ ;
  assign \new_[13222]_  = ~\new_[13675]_  | ~\new_[13613]_ ;
  assign \new_[13223]_  = ~\new_[14149]_  | ~\new_[13517]_ ;
  assign \new_[13224]_  = ~\new_[14000]_  & ~\new_[13620]_ ;
  assign \new_[13225]_  = ~\new_[6743]_  & ~\new_[13733]_ ;
  assign \new_[13226]_  = \new_[4503]_  ^ \new_[4511]_ ;
  assign \new_[13227]_  = ~\new_[14082]_  | ~\new_[3638]_ ;
  assign \new_[13228]_  = ~\new_[13261]_ ;
  assign \new_[13229]_  = ~\new_[4616]_  | ~\new_[4838]_ ;
  assign \new_[13230]_  = \new_[4372]_  ^ \new_[4503]_ ;
  assign \new_[13231]_  = ~\new_[14141]_  | ~\new_[13835]_ ;
  assign \new_[13232]_  = ~\new_[14228]_  & ~\new_[6277]_ ;
  assign \new_[13233]_  = ~\new_[6593]_  | ~\new_[14045]_ ;
  assign \new_[13234]_  = ~\new_[14231]_  | ~\new_[4966]_ ;
  assign \new_[13235]_  = ~\new_[14199]_  | ~\new_[3476]_ ;
  assign \new_[13236]_  = \new_[4509]_  ^ \new_[4510]_ ;
  assign \new_[13237]_  = ~\new_[13317]_ ;
  assign \new_[13238]_  = ~\new_[13428]_ ;
  assign \new_[13239]_  = ~\new_[6252]_  & ~\new_[13623]_ ;
  assign \new_[13240]_  = ~\new_[14156]_  | ~\new_[13920]_ ;
  assign \new_[13241]_  = \new_[4767]_  ^ \new_[4926]_ ;
  assign \new_[13242]_  = ~\new_[4073]_  | ~\new_[13904]_ ;
  assign \new_[13243]_  = ~\new_[6272]_  | ~\new_[13816]_ ;
  assign \new_[13244]_  = ~\new_[6284]_  & ~\new_[13635]_ ;
  assign \new_[13245]_  = \new_[14001]_  | \new_[3316]_ ;
  assign \new_[13246]_  = \new_[13810]_  & \new_[13348]_ ;
  assign \new_[13247]_  = \new_[14035]_  | \new_[13975]_ ;
  assign \new_[13248]_  = ~\new_[14058]_  | ~\new_[6033]_ ;
  assign \new_[13249]_  = ~\new_[13904]_  | ~\new_[4347]_ ;
  assign \new_[13250]_  = ~\new_[13985]_  & ~\new_[6545]_ ;
  assign \new_[13251]_  = ~\new_[14228]_  | ~\new_[6277]_ ;
  assign \new_[13252]_  = ~\new_[13394]_ ;
  assign \new_[13253]_  = ~\new_[6557]_  & ~\new_[13893]_ ;
  assign \new_[13254]_  = ~\new_[13396]_ ;
  assign \new_[13255]_  = ~\new_[6351]_  & ~\new_[6012]_ ;
  assign \new_[13256]_  = ~\new_[6348]_  & ~\new_[6512]_ ;
  assign \new_[13257]_  = ~\new_[13744]_ ;
  assign \new_[13258]_  = ~\new_[2932]_  | ~\new_[2870]_ ;
  assign \new_[13259]_  = ~\new_[6272]_  | ~\new_[3684]_ ;
  assign \new_[13260]_  = ~\new_[6264]_  & ~\new_[3428]_ ;
  assign \new_[13261]_  = \new_[2372]_  | \new_[2301]_ ;
  assign \new_[13262]_  = ~\new_[3337]_ ;
  assign \new_[13263]_  = ~\new_[9611]_  & ~\new_[6023]_ ;
  assign \new_[13264]_  = ~\new_[6557]_ ;
  assign \new_[13265]_  = ~\new_[4609]_  & ~\new_[4845]_ ;
  assign n8905 = \\VStatus_r_reg[5] ;
  assign \new_[13267]_  = ~\new_[13882]_ ;
  assign \new_[13268]_  = \new_[4291]_  & \new_[4288]_ ;
  assign n8920 = \\VStatus_r_reg[1] ;
  assign \new_[13270]_  = ~\new_[6247]_  & ~\new_[4236]_ ;
  assign \new_[13271]_  = ~\new_[3714]_ ;
  assign \new_[13272]_  = ~\new_[6323]_  & ~\new_[6198]_ ;
  assign n9025 = ~\new_[4779]_ ;
  assign \new_[13274]_  = ~\new_[6284]_  & ~\new_[3875]_ ;
  assign \new_[13275]_  = ~\new_[6272]_  & ~\new_[3684]_ ;
  assign \new_[13276]_  = ~\new_[3429]_  & ~\new_[3506]_ ;
  assign \new_[13277]_  = ~\new_[6557]_  & ~\new_[3478]_ ;
  assign \new_[13278]_  = \new_[2090]_  & \new_[2096]_ ;
  assign \new_[13279]_  = ~\new_[2349]_  & ~\new_[2316]_ ;
  assign \new_[13280]_  = ~\new_[6544]_  | ~\new_[3715]_ ;
  assign \new_[13281]_  = ~\new_[3883]_  & ~\new_[3815]_ ;
  assign \new_[13282]_  = ~\new_[6470]_ ;
  assign \new_[13283]_  = ~\new_[3883]_  & ~\new_[3687]_ ;
  assign \new_[13284]_  = ~\new_[13690]_ ;
  assign \new_[13285]_  = \new_[6809]_  | \new_[3713]_ ;
  assign \new_[13286]_  = ~\new_[3592]_  | ~\new_[3309]_ ;
  assign \new_[13287]_  = \new_[3689]_  | \new_[3712]_ ;
  assign \new_[13288]_  = ~\new_[13598]_ ;
  assign \new_[13289]_  = ~\new_[3466]_  | ~\new_[3310]_ ;
  assign \new_[13290]_  = ~\new_[4289]_  & ~\new_[4069]_ ;
  assign \new_[13291]_  = ~\new_[6255]_  & ~\new_[4347]_ ;
  assign \new_[13292]_  = ~\new_[2344]_  & ~\new_[2343]_ ;
  assign \new_[13293]_  = ~\new_[4792]_  & ~\new_[4794]_ ;
  assign \new_[13294]_  = ~\new_[6809]_  | ~\new_[3713]_ ;
  assign n9000 = \\VStatus_r_reg[3] ;
  assign \new_[13296]_  = ~rst_i;
  assign \new_[13297]_  = ~\new_[9645]_  | ~\new_[2673]_ ;
  assign \new_[13298]_  = ~\new_[13858]_ ;
  assign \new_[13299]_  = ~\new_[3282]_  & ~\new_[3879]_ ;
  assign \new_[13300]_  = \new_[3468]_  & \new_[3688]_ ;
  assign \new_[13301]_  = ~\new_[6324]_  & ~\new_[6326]_ ;
  assign \new_[13302]_  = ~\new_[14161]_ ;
  assign \new_[13303]_  = ~\new_[4505]_  & ~\new_[4552]_ ;
  assign \new_[13304]_  = ~\new_[6252]_  | ~\new_[3997]_ ;
  assign \new_[13305]_  = ~\new_[2477]_  & ~\new_[2476]_ ;
  assign \new_[13306]_  = ~\new_[6284]_  | ~\new_[3875]_ ;
  assign \new_[13307]_  = ~\new_[6275]_  & ~\new_[3712]_ ;
  assign \new_[13308]_  = \new_[6166]_  & \new_[3482]_ ;
  assign \new_[13309]_  = ~\new_[3626]_  & ~\new_[3712]_ ;
  assign \new_[13310]_  = ~\new_[3688]_  & ~\new_[3467]_ ;
  assign \new_[13311]_  = ~\new_[14156]_ ;
  assign \new_[13312]_  = ~n9145 | ~\new_[2876]_ ;
  assign \new_[13313]_  = ~\new_[2348]_  & ~\new_[2349]_ ;
  assign \new_[13314]_  = \new_[4509]_  | \new_[4553]_ ;
  assign \new_[13315]_  = ~\new_[11727]_ ;
  assign \new_[13316]_  = \new_[9372]_  & \new_[9471]_ ;
  assign \new_[13317]_  = ~\new_[6560]_  & ~\new_[6305]_ ;
  assign \new_[13318]_  = ~\new_[3806]_  & ~\new_[3890]_ ;
  assign \new_[13319]_  = \new_[2874]_  | \new_[2875]_ ;
  assign \new_[13320]_  = ~\new_[14317]_ ;
  assign \new_[13321]_  = \new_[6552]_  & \new_[3692]_ ;
  assign \new_[13322]_  = ~\new_[3882]_ ;
  assign \new_[13323]_  = ~\new_[4510]_  & ~\new_[4503]_ ;
  assign \new_[13324]_  = ~\new_[3316]_  | ~\new_[3315]_ ;
  assign \new_[13325]_  = \new_[6743]_  | \new_[4096]_ ;
  assign \new_[13326]_  = ~\new_[3938]_  | ~\new_[3940]_ ;
  assign \new_[13327]_  = ~\new_[14167]_ ;
  assign \new_[13328]_  = ~\\u0_rx_data_reg[2] ;
  assign n8910 = \\VStatus_r_reg[2] ;
  assign \new_[13330]_  = ~\new_[2524]_  & ~\new_[2454]_ ;
  assign \new_[13331]_  = \new_[6287]_  | \new_[3890]_ ;
  assign n8915 = u0_u0_resume_req_s1_reg;
  assign \new_[13333]_  = ~\new_[4792]_  & ~\new_[4795]_ ;
  assign \new_[13334]_  = ~\new_[6743]_  | ~\new_[4096]_ ;
  assign \new_[13335]_  = ~\new_[6690]_  | ~\new_[3508]_ ;
  assign \new_[13336]_  = ~\new_[4676]_  & ~\new_[4690]_ ;
  assign \new_[13337]_  = ~\new_[6461]_  & ~\new_[6556]_ ;
  assign n8940 = wb_cyc_i & wb_stb_i;
  assign \new_[13339]_  = ~\new_[2476]_  & ~\new_[2373]_ ;
  assign \new_[13340]_  = \new_[3510]_  | \new_[3509]_ ;
  assign \new_[13341]_  = ~\new_[2347]_  & ~\new_[2346]_ ;
  assign \new_[13342]_  = ~\new_[6544]_  & ~\new_[3715]_ ;
  assign \new_[13343]_  = ~\\u0_rx_data_reg[7] ;
  assign \new_[13344]_  = ~\new_[2340]_  & ~\new_[2317]_ ;
  assign \new_[13345]_  = ~u4_attach_r_reg;
  assign \new_[13346]_  = \new_[7853]_  | VControl_Load_pad_o;
  assign \new_[13347]_  = ~\new_[4812]_  | ~\new_[4814]_ ;
  assign \new_[13348]_  = ~\new_[4290]_ ;
  assign \new_[13349]_  = ~\\u0_rx_data_reg[3] ;
  assign \new_[13350]_  = ~\new_[3504]_  | ~\new_[3505]_ ;
  assign \new_[13351]_  = \new_[3884]_  & \new_[3882]_ ;
  assign \new_[13352]_  = ~\wb_addr_i[2]  & ~\wb_addr_i[3] ;
  assign \new_[13353]_  = ~\new_[2086]_  | ~\new_[2087]_ ;
  assign n8995 = u4_u3_r4_reg;
  assign \new_[13355]_  = ~\new_[3481]_  | ~\new_[3479]_ ;
  assign \new_[13356]_  = \new_[8703]_  & \new_[8702]_ ;
  assign \new_[13357]_  = ~\new_[3482]_  & ~\new_[3689]_ ;
  assign \new_[13358]_  = ~\new_[3317]_  & ~\new_[3478]_ ;
  assign \new_[13359]_  = ~\new_[2875]_  | ~\new_[2857]_ ;
  assign \new_[13360]_  = ~\new_[6252]_  & ~\new_[3997]_ ;
  assign \new_[13361]_  = ~\new_[3505]_  | ~\new_[3480]_ ;
  assign \new_[13362]_  = ~n9145 | ~\new_[2874]_ ;
  assign \new_[13363]_  = ~\new_[3879]_  | ~\new_[3787]_ ;
  assign \new_[13364]_  = ~\new_[6005]_ ;
  assign \new_[13365]_  = ~\new_[3691]_  | ~\new_[3638]_ ;
  assign \new_[13366]_  = \wb_addr_i[5]  & \wb_addr_i[6] ;
  assign \new_[13367]_  = ~\new_[2871]_ ;
  assign \new_[13368]_  = ~\new_[4074]_  & ~\new_[4347]_ ;
  assign \new_[13369]_  = ~\new_[13933]_ ;
  assign \new_[13370]_  = u1_u3_out_to_small_reg;
  assign \new_[13371]_  = ~\new_[3710]_ ;
  assign \new_[13372]_  = ~\new_[6255]_ ;
  assign \new_[13373]_  = ~resume_req_i & ~n9120;
  assign \new_[13374]_  = ~\new_[4288]_ ;
  assign \new_[13375]_  = ~\new_[2088]_  | ~\new_[2089]_ ;
  assign \new_[13376]_  = \new_[4858]_  & \new_[4859]_ ;
  assign \new_[13377]_  = ~\new_[2317]_  & ~\new_[2341]_ ;
  assign \new_[13378]_  = ~\new_[3475]_  | ~\new_[3474]_ ;
  assign \new_[13379]_  = ~\new_[3309]_  & ~\new_[3686]_ ;
  assign \new_[13380]_  = \new_[6254]_  & \new_[4074]_ ;
  assign \new_[13381]_  = \new_[6593]_  | \new_[3340]_ ;
  assign \new_[13382]_  = \new_[3932]_  & \new_[4289]_ ;
  assign \new_[13383]_  = \new_[8658]_  & \new_[8954]_ ;
  assign \new_[13384]_  = ~\new_[6264]_  | ~\new_[3428]_ ;
  assign \new_[13385]_  = ~\new_[2372]_  & ~\new_[2392]_ ;
  assign \new_[13386]_  = ~\new_[13950]_ ;
  assign \new_[13387]_  = ~\new_[6567]_  & ~\new_[3506]_ ;
  assign \new_[13388]_  = ~\new_[3308]_  & ~\new_[3466]_ ;
  assign \new_[13389]_  = ~\new_[7206]_ ;
  assign \new_[13390]_  = ~n8990 & ~\new_[2452]_ ;
  assign \new_[13391]_  = ~\new_[4237]_  & ~\new_[4197]_ ;
  assign \new_[13392]_  = ~\new_[2876]_  & ~\new_[2869]_ ;
  assign \new_[13393]_  = ~\new_[4095]_ ;
  assign \new_[13394]_  = ~\new_[14485]_ ;
  assign \new_[13395]_  = ~\new_[2373]_  & ~\new_[2392]_ ;
  assign \new_[13396]_  = ~\new_[6561]_  & ~\new_[3317]_ ;
  assign \new_[13397]_  = \new_[2876]_  | \new_[2857]_ ;
  assign \new_[13398]_  = ~\new_[13920]_ ;
  assign \new_[13399]_  = \new_[6552]_  | \new_[3692]_ ;
  assign \new_[13400]_  = \new_[6561]_  & \new_[3317]_ ;
  assign n9010 = ~\new_[6484]_ ;
  assign n9020 = ~\new_[6733]_ ;
  assign \new_[13403]_  = ~\new_[14141]_ ;
  assign n8945 = u4_u1_r4_reg;
  assign \new_[13405]_  = ~\new_[3638]_ ;
  assign \new_[13406]_  = ~\new_[2348]_  & ~\new_[2347]_ ;
  assign \new_[13407]_  = ~\new_[13691]_ ;
  assign \new_[13408]_  = \\LineState_r_reg[0] ;
  assign \new_[13409]_  = ~\new_[3062]_ ;
  assign \new_[13410]_  = ~n9145 | ~\new_[2875]_ ;
  assign \new_[13411]_  = ~\new_[3465]_  | ~\new_[3473]_ ;
  assign \new_[13412]_  = \new_[3472]_  & \new_[3473]_ ;
  assign \new_[13413]_  = ~\new_[4073]_  | ~\new_[4070]_ ;
  assign n8930 = \\VStatus_r_reg[4] ;
  assign \new_[13415]_  = ~\new_[13658]_ ;
  assign \new_[13416]_  = ~\new_[3062]_  & ~\new_[3031]_ ;
  assign \new_[13417]_  = ~\new_[3686]_  | ~\new_[3464]_ ;
  assign \new_[13418]_  = ~\\u0_rx_data_reg[0] ;
  assign \new_[13419]_  = ~\new_[7670]_  & ~\new_[2210]_ ;
  assign \new_[13420]_  = ~\new_[2340]_  & ~\new_[2316]_ ;
  assign \new_[13421]_  = ~\new_[4097]_ ;
  assign \new_[13422]_  = ~\new_[3502]_ ;
  assign \new_[13423]_  = \new_[2875]_  | \new_[2857]_ ;
  assign \new_[13424]_  = ~\new_[4816]_  | ~\new_[4817]_ ;
  assign n8955 = u4_u0_r4_reg;
  assign \new_[13426]_  = ~\new_[4787]_  | ~\new_[8959]_ ;
  assign \new_[13427]_  = ~\wb_addr_i[2]  | ~\wb_addr_i[3] ;
  assign \new_[13428]_  = ~\new_[11431]_  | ~\new_[4873]_ ;
  assign \new_[13429]_  = ~\new_[3311]_  & ~\new_[4091]_ ;
  assign \new_[13430]_  = ~\new_[3788]_  | ~\new_[3691]_ ;
  assign \new_[13431]_  = ~\wb_addr_i[7]  & ~\wb_addr_i[8] ;
  assign \new_[13432]_  = \new_[2094]_  & \new_[2083]_ ;
  assign \new_[13433]_  = ~\\u0_rx_data_reg[5] ;
  assign \new_[13434]_  = ~\new_[4839]_  | ~\new_[4840]_ ;
  assign \new_[13435]_  = ~\new_[3688]_  & ~\new_[3689]_ ;
  assign \new_[13436]_  = ~\new_[2961]_ ;
  assign \new_[13437]_  = ~\new_[2479]_  & ~n8990;
  assign \new_[13438]_  = ~\new_[14084]_ ;
  assign n8925 = \\VStatus_r_reg[7] ;
  assign \new_[13440]_  = ~\new_[6010]_ ;
  assign \new_[13441]_  = ~\\u0_u0_line_state_r_reg[1] ;
  assign \new_[13442]_  = ~\new_[14486]_ ;
  assign \new_[13443]_  = ~\new_[5993]_  & ~\new_[2453]_ ;
  assign \new_[13444]_  = ~\new_[6005]_  & ~\new_[3689]_ ;
  assign \new_[13445]_  = ~\new_[3435]_  | ~\new_[3463]_ ;
  assign \new_[13446]_  = ~\\u0_rx_data_reg[6] ;
  assign \new_[13447]_  = ~\new_[3692]_  & ~\new_[3815]_ ;
  assign \new_[13448]_  = \\u0_u0_line_state_r_reg[0] ;
  assign \new_[13449]_  = ~\\u0_rx_data_reg[4] ;
  assign \new_[13450]_  = ~\new_[2991]_ ;
  assign \new_[13451]_  = ~\new_[2478]_  & ~\new_[2479]_ ;
  assign \new_[13452]_  = \new_[8700]_  | \new_[8888]_ ;
  assign \new_[13453]_  = ~\\u0_rx_data_reg[1] ;
  assign \new_[13454]_  = ~\new_[3283]_  & ~\new_[3938]_ ;
  assign \new_[13455]_  = \new_[6196]_  | \new_[4197]_ ;
  assign \new_[13456]_  = ~\new_[13877]_ ;
  assign \new_[13457]_  = ~\new_[13835]_ ;
  assign \new_[13458]_  = ~\new_[4161]_  & ~\new_[3781]_ ;
  assign \new_[13459]_  = \new_[3671]_  & \new_[3883]_ ;
  assign \new_[13460]_  = ~\new_[4835]_  | ~\new_[4837]_ ;
  assign \new_[13461]_  = ~\new_[3693]_  | ~\new_[3690]_ ;
  assign \new_[13462]_  = ~\new_[4289]_  & ~\new_[4347]_ ;
  assign \new_[13463]_  = \new_[6690]_  | \new_[3508]_ ;
  assign \new_[13464]_  = ~\new_[14226]_ ;
  assign \new_[13465]_  = \\LineState_r_reg[1] ;
  assign \new_[13466]_  = \new_[3480]_  & \new_[3476]_ ;
  assign n8985 = u4_u2_r4_reg;
  assign \new_[13468]_  = \new_[3478]_  | \new_[3506]_ ;
  assign \new_[13469]_  = ~\new_[13616]_ ;
  assign \new_[13470]_  = ~\new_[3462]_  | ~\new_[3308]_ ;
  assign \new_[13471]_  = \new_[3815]_  | \new_[3890]_ ;
  assign \new_[13472]_  = \new_[4347]_  | \new_[4197]_ ;
  assign \new_[13473]_  = \new_[3313]_  & \new_[3477]_ ;
  assign \new_[13474]_  = ~\new_[4511]_  & ~\new_[4372]_ ;
  assign n9015 = ~\new_[6365]_ ;
  assign \new_[13476]_  = ~\new_[3035]_  & ~\new_[3037]_ ;
  assign \new_[13477]_  = ~\wb_addr_i[17] ;
  assign \new_[13478]_  = ~\new_[4838]_ ;
  assign \new_[13479]_  = ~\new_[6593]_  | ~\new_[3340]_ ;
  assign \new_[13480]_  = ~\new_[6010]_  & ~\new_[3815]_ ;
  assign \new_[13481]_  = ~\new_[13748]_ ;
  assign \new_[13482]_  = ~\new_[6166]_  & ~\new_[3482]_ ;
  assign \new_[13483]_  = ~\new_[3172]_  & ~\new_[2982]_ ;
  assign n8965 = \\VStatus_r_reg[6] ;
  assign \new_[13485]_  = ~\new_[3477]_  & ~\new_[3478]_ ;
  assign \new_[13486]_  = ~\new_[3477]_  & ~\new_[3312]_ ;
  assign n8935 = \\VStatus_r_reg[0] ;
  assign \new_[13488]_  = \new_[6254]_  | \new_[4074]_ ;
  assign \new_[13489]_  = ~\new_[2876]_  | ~\new_[2869]_ ;
  assign \new_[13490]_  = ~\new_[3476]_ ;
  assign \new_[13491]_  = ~\new_[6247]_  | ~\new_[4236]_ ;
  assign \new_[13492]_  = \new_[3711]_  & \new_[3788]_ ;
  assign \new_[13493]_  = \new_[9421]_  | \new_[9456]_ ;
  assign \new_[13494]_  = ~\new_[14216]_ ;
  assign \new_[13495]_  = \new_[9424]_  & \new_[9442]_ ;
  assign \new_[13496]_  = ~\new_[14254]_ ;
  assign \new_[13497]_  = ~\new_[3341]_ ;
  assign \new_[13498]_  = ~\new_[3737]_ ;
  assign \new_[13499]_  = ~\new_[3517]_ ;
  assign \new_[13500]_  = ~\new_[6468]_ ;
  assign \new_[13501]_  = ~\new_[3177]_ ;
  assign \new_[13502]_  = ~\new_[4808]_ ;
  assign \new_[13503]_  = ~\new_[3357]_ ;
  assign \new_[13504]_  = ~\new_[3439]_ ;
  assign \new_[13505]_  = ~\new_[4826]_ ;
  assign \new_[13506]_  = ~\new_[6461]_ ;
  assign \new_[13507]_  = ~\new_[6165]_ ;
  assign \new_[13508]_  = ~\new_[4813]_ ;
  assign \new_[13509]_  = ~\new_[7156]_ ;
  assign n9065 = ~\new_[5140]_ ;
  assign \new_[13511]_  = ~\new_[3706]_ ;
  assign \new_[13512]_  = ~\new_[6728]_ ;
  assign \new_[13513]_  = ~\new_[3681]_ ;
  assign \new_[13514]_  = ~\new_[3895]_ ;
  assign \new_[13515]_  = ~\new_[6691]_ ;
  assign \new_[13516]_  = ~\new_[3701]_ ;
  assign \new_[13517]_  = ~\new_[6320]_ ;
  assign \new_[13518]_  = ~\new_[6653]_ ;
  assign \new_[13519]_  = ~\new_[6378]_ ;
  assign \new_[13520]_  = ~\new_[2802]_ ;
  assign \new_[13521]_  = ~\new_[4071]_ ;
  assign \new_[13522]_  = ~\new_[3878]_ ;
  assign \new_[13523]_  = ~\new_[4823]_ ;
  assign \new_[13524]_  = ~\new_[3156]_ ;
  assign \new_[13525]_  = ~\new_[7258]_ ;
  assign \new_[13526]_  = ~\new_[4825]_ ;
  assign \new_[13527]_  = ~\new_[3189]_ ;
  assign \new_[13528]_  = ~\new_[3460]_ ;
  assign \new_[13529]_  = ~\new_[3184]_ ;
  assign \new_[13530]_  = ~\new_[4829]_ ;
  assign \new_[13531]_  = ~\new_[4830]_ ;
  assign \new_[13532]_  = ~\new_[2392]_ ;
  assign \new_[13533]_  = ~\new_[6878]_ ;
  assign \new_[13534]_  = ~\new_[6298]_ ;
  assign \new_[13535]_  = ~\new_[3500]_ ;
  assign \new_[13536]_  = ~\new_[3594]_ ;
  assign \new_[13537]_  = ~\new_[3677]_ ;
  assign \new_[13538]_  = ~\new_[3157]_ ;
  assign \new_[13539]_  = ~\new_[3353]_ ;
  assign \new_[13540]_  = ~\new_[6366]_ ;
  assign \new_[13541]_  = ~\new_[5135]_ ;
  assign \new_[13542]_  = ~\new_[6490]_ ;
  assign \new_[13543]_  = ~\new_[3483]_ ;
  assign n9035 = ~\new_[7853]_ ;
  assign \new_[13545]_  = ~\new_[3352]_ ;
  assign \new_[13546]_  = ~\new_[4766]_ ;
  assign \new_[13547]_  = ~\new_[4648]_ ;
  assign \new_[13548]_  = ~\new_[6347]_ ;
  assign \new_[13549]_  = ~\new_[4003]_ ;
  assign \new_[13550]_  = ~\new_[3932]_ ;
  assign \new_[13551]_  = ~\new_[3731]_ ;
  assign \new_[13552]_  = ~\new_[6266]_ ;
  assign \new_[13553]_  = ~\new_[3297]_ ;
  assign \new_[13554]_  = ~\new_[3720]_ ;
  assign \new_[13555]_  = ~\new_[6305]_ ;
  assign \new_[13556]_  = ~\new_[4353]_ ;
  assign \new_[13557]_  = ~\new_[3345]_ ;
  assign \new_[13558]_  = ~\new_[5128]_ ;
  assign \new_[13559]_  = ~\new_[6090]_ ;
  assign \new_[13560]_  = ~\new_[3869]_ ;
  assign \new_[13561]_  = ~\new_[2039]_ ;
  assign \new_[13562]_  = ~\new_[3318]_ ;
  assign \new_[13563]_  = ~\new_[6873]_ ;
  assign \new_[13564]_  = ~\new_[7155]_ ;
  assign \new_[13565]_  = ~\new_[5130]_ ;
  assign \new_[13566]_  = ~\new_[3104]_ ;
  assign \new_[13567]_  = ~\new_[5131]_ ;
  assign \new_[13568]_  = ~\new_[2836]_ ;
  assign \new_[13569]_  = ~\new_[2932]_ ;
  assign \new_[13570]_  = ~\new_[2673]_ ;
  assign \new_[13571]_  = ~\new_[6602]_ ;
  assign \new_[13572]_  = ~\new_[4961]_ ;
  assign \new_[13573]_  = ~\new_[5132]_ ;
  assign \new_[13574]_  = ~\new_[6297]_ ;
  assign \new_[13575]_  = ~\new_[9916]_ ;
  assign \new_[13576]_  = ~\new_[4849]_ ;
  assign n9030 = ~\new_[7763]_ ;
  assign \new_[13578]_  = ~\new_[3709]_ ;
  assign \new_[13579]_  = ~\new_[7278]_ ;
  assign \new_[13580]_  = ~\new_[3192]_ ;
  assign \new_[13581]_  = ~\new_[4820]_ ;
  assign \new_[13582]_  = ~\new_[3181]_ ;
  assign \new_[13583]_  = ~\new_[2087]_ ;
  assign \new_[13584]_  = ~\new_[6551]_ ;
  assign \new_[13585]_  = ~\new_[2345]_ ;
  assign \new_[13586]_  = ~\new_[7164]_ ;
  assign \new_[13587]_  = ~\new_[3457]_ ;
  assign \new_[13588]_  = ~\new_[12437]_ ;
  assign \new_[13589]_  = ~\new_[3162]_ ;
  assign \new_[13590]_  = ~\new_[3305]_ ;
  assign n9090 = ~\new_[5143]_ ;
  assign \new_[13592]_  = ~\new_[4088]_ ;
  assign \new_[13593]_  = ~\new_[3881]_ ;
  assign \new_[13594]_  = ~\new_[4863]_ ;
  assign \new_[13595]_  = ~\new_[2611]_ ;
  assign \new_[13596]_  = ~\new_[3304]_ ;
  assign \new_[13597]_  = ~\new_[6486]_ ;
  assign \new_[13598]_  = ~\new_[4653]_ ;
  assign \new_[13599]_  = ~\new_[5617]_ ;
  assign \new_[13600]_  = ~\new_[3824]_ ;
  assign \new_[13601]_  = ~\new_[4804]_ ;
  assign \new_[13602]_  = ~\new_[6862]_ ;
  assign \new_[13603]_  = ~\new_[3514]_ ;
  assign n9085 = ~\new_[5142]_ ;
  assign \new_[13605]_  = ~\new_[3518]_ ;
  assign \new_[13606]_  = ~\new_[3038]_ ;
  assign \new_[13607]_  = ~\new_[3453]_ ;
  assign \new_[13608]_  = ~\new_[3040]_ ;
  assign \new_[13609]_  = ~\new_[6379]_ ;
  assign \new_[13610]_  = ~\new_[6169]_ ;
  assign \new_[13611]_  = ~\new_[6865]_ ;
  assign \new_[13612]_  = ~\new_[3704]_ ;
  assign \new_[13613]_  = ~\new_[6301]_ ;
  assign \new_[13614]_  = ~\new_[7277]_ ;
  assign \new_[13615]_  = ~\new_[6876]_ ;
  assign \new_[13616]_  = ~\new_[5501]_ ;
  assign \new_[13617]_  = ~\new_[6544]_ ;
  assign \new_[13618]_  = ~\new_[3723]_ ;
  assign \new_[13619]_  = ~\new_[3738]_ ;
  assign \new_[13620]_  = ~\new_[2993]_ ;
  assign \new_[13621]_  = ~\new_[6286]_ ;
  assign \new_[13622]_  = ~\new_[3498]_ ;
  assign \new_[13623]_  = ~\new_[4206]_ ;
  assign \new_[13624]_  = ~\new_[6348]_ ;
  assign \new_[13625]_  = ~\new_[3726]_ ;
  assign \new_[13626]_  = ~n8945;
  assign \new_[13627]_  = ~\new_[6257]_ ;
  assign \new_[13628]_  = ~\new_[4827]_ ;
  assign \new_[13629]_  = ~\new_[6251]_ ;
  assign \new_[13630]_  = ~\new_[5126]_ ;
  assign \new_[13631]_  = ~\new_[6274]_ ;
  assign \new_[13632]_  = ~\new_[3399]_ ;
  assign \new_[13633]_  = ~\new_[6015]_ ;
  assign \new_[13634]_  = ~\new_[6331]_ ;
  assign \new_[13635]_  = ~\new_[3790]_ ;
  assign n9080 = ~\new_[5139]_ ;
  assign \new_[13637]_  = ~\new_[6339]_ ;
  assign \new_[13638]_  = ~\new_[6880]_ ;
  assign \new_[13639]_  = ~\new_[3702]_ ;
  assign \new_[13640]_  = ~\new_[3892]_ ;
  assign \new_[13641]_  = ~\new_[3344]_ ;
  assign \new_[13642]_  = ~\new_[2034]_ ;
  assign \new_[13643]_  = ~\new_[6324]_ ;
  assign \new_[13644]_  = ~\new_[4851]_ ;
  assign \new_[13645]_  = ~\new_[6235]_ ;
  assign \new_[13646]_  = ~\new_[4620]_ ;
  assign \new_[13647]_  = ~\new_[7149]_ ;
  assign \new_[13648]_  = ~\new_[4078]_ ;
  assign \new_[13649]_  = ~\new_[6254]_ ;
  assign \new_[13650]_  = ~\new_[5134]_ ;
  assign \new_[13651]_  = ~\new_[3423]_ ;
  assign \new_[13652]_  = ~\new_[3487]_ ;
  assign \new_[13653]_  = ~\new_[6355]_ ;
  assign \new_[13654]_  = ~\new_[4806]_ ;
  assign \new_[13655]_  = ~\new_[2373]_ ;
  assign \new_[13656]_  = ~\new_[6196]_ ;
  assign \new_[13657]_  = ~\new_[2193]_ ;
  assign \new_[13658]_  = ~\new_[8809]_ ;
  assign \new_[13659]_  = ~\new_[2992]_ ;
  assign \new_[13660]_  = ~\new_[3887]_ ;
  assign \new_[13661]_  = ~\new_[5760]_ ;
  assign \new_[13662]_  = ~\new_[3891]_ ;
  assign \new_[13663]_  = ~\new_[4500]_ ;
  assign \new_[13664]_  = ~\new_[4678]_ ;
  assign \new_[13665]_  = ~\new_[3725]_ ;
  assign \new_[13666]_  = ~\new_[3027]_ ;
  assign \new_[13667]_  = ~\new_[2549]_ ;
  assign \new_[13668]_  = ~\new_[6357]_ ;
  assign \new_[13669]_  = ~\new_[3164]_ ;
  assign \new_[13670]_  = ~\new_[3886]_ ;
  assign \new_[13671]_  = ~\new_[3321]_ ;
  assign \new_[13672]_  = ~\new_[6335]_ ;
  assign \new_[13673]_  = ~\new_[5994]_ ;
  assign \new_[13674]_  = ~\new_[5136]_ ;
  assign \new_[13675]_  = ~\new_[6302]_ ;
  assign \new_[13676]_  = ~\new_[4931]_ ;
  assign \new_[13677]_  = ~\new_[6338]_ ;
  assign \new_[13678]_  = ~\new_[3132]_ ;
  assign \new_[13679]_  = ~\new_[4783]_ ;
  assign \new_[13680]_  = ~\new_[4846]_ ;
  assign \new_[13681]_  = ~\new_[6869]_ ;
  assign \new_[13682]_  = ~\new_[4092]_ ;
  assign \new_[13683]_  = ~\new_[3430]_ ;
  assign \new_[13684]_  = ~\new_[3735]_ ;
  assign \new_[13685]_  = ~\new_[3185]_ ;
  assign \new_[13686]_  = ~\new_[3525]_ ;
  assign \new_[13687]_  = ~\new_[3349]_ ;
  assign \new_[13688]_  = ~\new_[3456]_ ;
  assign \new_[13689]_  = ~\new_[4070]_ ;
  assign \new_[13690]_  = ~\new_[4686]_ ;
  assign \new_[13691]_  = ~\new_[5997]_ ;
  assign \new_[13692]_  = ~\new_[4768]_ ;
  assign \new_[13693]_  = ~\new_[6098]_ ;
  assign \new_[13694]_  = ~\new_[3039]_ ;
  assign \new_[13695]_  = ~\wb_addr_i[3] ;
  assign \new_[13696]_  = ~\new_[6603]_ ;
  assign \new_[13697]_  = ~\new_[3703]_ ;
  assign \new_[13698]_  = ~\new_[2342]_ ;
  assign \new_[13699]_  = ~\LineState_pad_i[0] ;
  assign \new_[13700]_  = ~\new_[6313]_ ;
  assign \new_[13701]_  = ~\new_[3168]_ ;
  assign \new_[13702]_  = ~\new_[6726]_ ;
  assign \new_[13703]_  = ~\new_[4950]_ ;
  assign \new_[13704]_  = ~\new_[6881]_ ;
  assign \new_[13705]_  = ~\new_[6556]_ ;
  assign \new_[13706]_  = ~\new_[3868]_ ;
  assign \new_[13707]_  = ~\new_[3492]_ ;
  assign \new_[13708]_  = ~\new_[2076]_ ;
  assign \new_[13709]_  = ~\new_[3354]_ ;
  assign \new_[13710]_  = ~\new_[4782]_ ;
  assign \new_[13711]_  = ~\new_[6245]_ ;
  assign \new_[13712]_  = ~\new_[6729]_ ;
  assign \new_[13713]_  = ~\new_[3434]_ ;
  assign \new_[13714]_  = ~\new_[3808]_ ;
  assign \new_[13715]_  = ~\new_[5133]_ ;
  assign \new_[13716]_  = ~\new_[3622]_ ;
  assign \new_[13717]_  = ~\new_[3998]_ ;
  assign \new_[13718]_  = ~\new_[6234]_ ;
  assign \new_[13719]_  = ~\new_[3695]_ ;
  assign \new_[13720]_  = ~\new_[6294]_ ;
  assign \new_[13721]_  = ~\new_[6701]_ ;
  assign \new_[13722]_  = ~\new_[3301]_ ;
  assign \new_[13723]_  = ~\new_[4828]_ ;
  assign \new_[13724]_  = ~\new_[4089]_ ;
  assign \new_[13725]_  = ~\new_[3175]_ ;
  assign \new_[13726]_  = ~\new_[3299]_ ;
  assign \new_[13727]_  = ~\new_[4087]_ ;
  assign \new_[13728]_  = ~\new_[6353]_ ;
  assign \new_[13729]_  = ~\new_[3519]_ ;
  assign \new_[13730]_  = ~\new_[3699]_ ;
  assign \new_[13731]_  = ~\new_[4076]_ ;
  assign \new_[13732]_  = ~\new_[5495]_ ;
  assign \new_[13733]_  = ~\new_[4292]_ ;
  assign \new_[13734]_  = ~\new_[6608]_ ;
  assign \new_[13735]_  = ~\new_[3022]_ ;
  assign \new_[13736]_  = ~\new_[4077]_ ;
  assign \new_[13737]_  = ~\new_[3683]_ ;
  assign \new_[13738]_  = ~\new_[3679]_ ;
  assign \new_[13739]_  = ~\new_[3495]_ ;
  assign \new_[13740]_  = ~\new_[4791]_ ;
  assign \new_[13741]_  = ~\new_[6934]_ ;
  assign \new_[13742]_  = ~\new_[6872]_ ;
  assign \new_[13743]_  = ~\new_[3727]_ ;
  assign \new_[13744]_  = ~\new_[5585]_ ;
  assign \new_[13745]_  = ~\new_[3733]_ ;
  assign \new_[13746]_  = ~\new_[3875]_ ;
  assign \new_[13747]_  = ~\new_[6299]_ ;
  assign \new_[13748]_  = ~\new_[6022]_ ;
  assign \new_[13749]_  = ~\new_[4677]_ ;
  assign \new_[13750]_  = ~\new_[6564]_ ;
  assign \new_[13751]_  = ~\new_[6253]_ ;
  assign \new_[13752]_  = ~\new_[6560]_ ;
  assign \new_[13753]_  = ~\new_[6032]_ ;
  assign \new_[13754]_  = ~\new_[6304]_ ;
  assign \new_[13755]_  = ~\new_[4784]_ ;
  assign \new_[13756]_  = ~\new_[4800]_ ;
  assign \new_[13757]_  = ~\new_[2573]_ ;
  assign \new_[13758]_  = ~\new_[3527]_ ;
  assign \new_[13759]_  = ~\new_[4831]_ ;
  assign \new_[13760]_  = ~\new_[5109]_ ;
  assign \new_[13761]_  = ~\new_[6319]_ ;
  assign \new_[13762]_  = ~\new_[3327]_ ;
  assign \new_[13763]_  = ~\new_[6732]_ ;
  assign \new_[13764]_  = ~\new_[6271]_ ;
  assign \new_[13765]_  = ~\new_[6488]_ ;
  assign \new_[13766]_  = ~\new_[2097]_ ;
  assign \new_[13767]_  = ~\new_[3169]_ ;
  assign \new_[13768]_  = ~\new_[6270]_ ;
  assign \new_[13769]_  = ~\new_[4960]_ ;
  assign \new_[13770]_  = ~\new_[6019]_ ;
  assign \new_[13771]_  = ~\new_[3781]_ ;
  assign \new_[13772]_  = ~\new_[4075]_ ;
  assign \new_[13773]_  = ~\new_[3323]_ ;
  assign \new_[13774]_  = ~\new_[3698]_ ;
  assign \new_[13775]_  = ~\new_[3182]_ ;
  assign \new_[13776]_  = ~\new_[3729]_ ;
  assign \new_[13777]_  = ~\new_[3628]_ ;
  assign \new_[13778]_  = ~\new_[3311]_ ;
  assign \new_[13779]_  = ~\new_[6323]_ ;
  assign \new_[13780]_  = ~\new_[7162]_ ;
  assign n9070 = ~\new_[5141]_ ;
  assign \new_[13782]_  = ~\new_[3894]_ ;
  assign \new_[13783]_  = ~\new_[6361]_ ;
  assign \new_[13784]_  = ~\new_[3336]_ ;
  assign \new_[13785]_  = ~\new_[4621]_ ;
  assign \new_[13786]_  = ~\new_[3484]_ ;
  assign \new_[13787]_  = ~\new_[6097]_ ;
  assign \new_[13788]_  = ~\new_[6368]_ ;
  assign \new_[13789]_  = ~\new_[3450]_ ;
  assign \new_[13790]_  = ~\new_[5756]_ ;
  assign \new_[13791]_  = ~\new_[3629]_ ;
  assign \new_[13792]_  = ~\new_[3486]_ ;
  assign \new_[13793]_  = ~\new_[6588]_ ;
  assign \new_[13794]_  = ~\new_[3507]_ ;
  assign \new_[13795]_  = ~\new_[3621]_ ;
  assign \new_[13796]_  = ~\new_[2458]_ ;
  assign \new_[13797]_  = ~\new_[6358]_ ;
  assign \new_[13798]_  = ~\new_[3777]_ ;
  assign \new_[13799]_  = ~\new_[3023]_ ;
  assign \new_[13800]_  = ~\new_[3458]_ ;
  assign \new_[13801]_  = ~\new_[4821]_ ;
  assign \new_[13802]_  = ~\new_[8826]_ ;
  assign \new_[13803]_  = ~n9005;
  assign \new_[13804]_  = ~\new_[3718]_ ;
  assign \new_[13805]_  = ~\new_[6359]_ ;
  assign \new_[13806]_  = ~\new_[3280]_ ;
  assign \new_[13807]_  = ~\new_[6273]_ ;
  assign \new_[13808]_  = ~\new_[6317]_ ;
  assign \new_[13809]_  = ~\new_[6489]_ ;
  assign \new_[13810]_  = ~\new_[4161]_ ;
  assign \new_[13811]_  = ~\new_[2455]_ ;
  assign \new_[13812]_  = ~\new_[3867]_ ;
  assign \new_[13813]_  = ~\new_[2301]_ ;
  assign \new_[13814]_  = ~\new_[3479]_ ;
  assign \new_[13815]_  = ~\new_[5127]_ ;
  assign \new_[13816]_  = ~\new_[3592]_ ;
  assign \new_[13817]_  = ~\new_[2135]_ ;
  assign \new_[13818]_  = ~\new_[3421]_ ;
  assign \new_[13819]_  = ~\new_[3028]_ ;
  assign \new_[13820]_  = ~\new_[3724]_ ;
  assign \new_[13821]_  = ~\new_[7157]_ ;
  assign \new_[13822]_  = ~\new_[3523]_ ;
  assign \new_[13823]_  = ~\new_[2173]_ ;
  assign \new_[13824]_  = ~\new_[3639]_ ;
  assign \new_[13825]_  = ~\new_[6091]_ ;
  assign \new_[13826]_  = ~\new_[4081]_ ;
  assign \new_[13827]_  = ~\new_[5137]_ ;
  assign \new_[13828]_  = ~\new_[2088]_ ;
  assign \new_[13829]_  = ~\new_[6318]_ ;
  assign \new_[13830]_  = ~\new_[3180]_ ;
  assign \new_[13831]_  = ~\new_[3188]_ ;
  assign n9060 = ~\new_[5242]_ ;
  assign \new_[13833]_  = ~\new_[3893]_ ;
  assign \new_[13834]_  = ~\new_[3870]_ ;
  assign \new_[13835]_  = ~\new_[3832]_ ;
  assign \new_[13836]_  = ~\new_[3696]_ ;
  assign \new_[13837]_  = ~\new_[2473]_ ;
  assign \new_[13838]_  = ~\new_[3329]_ ;
  assign \new_[13839]_  = ~\new_[3736]_ ;
  assign \new_[13840]_  = ~\new_[3293]_ ;
  assign \new_[13841]_  = ~\new_[3526]_ ;
  assign \new_[13842]_  = ~TxReady_pad_i;
  assign \new_[13843]_  = ~\new_[3449]_ ;
  assign \new_[13844]_  = ~\new_[2171]_ ;
  assign \new_[13845]_  = ~\new_[2073]_ ;
  assign \new_[13846]_  = ~\new_[3187]_ ;
  assign \new_[13847]_  = ~\new_[4930]_ ;
  assign \new_[13848]_  = ~\new_[6007]_ ;
  assign \new_[13849]_  = ~\new_[7200]_ ;
  assign \new_[13850]_  = ~\new_[7856]_ ;
  assign \new_[13851]_  = ~\new_[5138]_ ;
  assign \new_[13852]_  = ~\new_[5124]_ ;
  assign \new_[13853]_  = ~\new_[3330]_ ;
  assign \new_[13854]_  = ~\new_[3433]_ ;
  assign \new_[13855]_  = ~\new_[6481]_ ;
  assign \new_[13856]_  = ~\new_[3452]_ ;
  assign \new_[13857]_  = ~\new_[6312]_ ;
  assign \new_[13858]_  = ~\new_[5124]_ ;
  assign \new_[13859]_  = ~\new_[3351]_ ;
  assign \new_[13860]_  = ~\new_[4182]_ ;
  assign \new_[13861]_  = ~\new_[4798]_ ;
  assign \new_[13862]_  = ~\new_[4797]_ ;
  assign \new_[13863]_  = ~\new_[7285]_ ;
  assign \new_[13864]_  = ~\new_[3521]_ ;
  assign \new_[13865]_  = ~\new_[3930]_ ;
  assign \new_[13866]_  = ~\new_[6198]_ ;
  assign \new_[13867]_  = ~\new_[3431]_ ;
  assign \new_[13868]_  = ~\new_[3176]_ ;
  assign \new_[13869]_  = ~\new_[3307]_ ;
  assign \new_[13870]_  = ~\new_[3033]_ ;
  assign \new_[13871]_  = ~\new_[3159]_ ;
  assign \new_[13872]_  = ~\new_[6592]_ ;
  assign \new_[13873]_  = ~\new_[4090]_ ;
  assign \new_[13874]_  = ~\new_[6693]_ ;
  assign \new_[13875]_  = ~\new_[6346]_ ;
  assign \new_[13876]_  = ~\new_[3690]_ ;
  assign \new_[13877]_  = ~\new_[6021]_ ;
  assign \new_[13878]_  = ~\new_[4875]_ ;
  assign \new_[13879]_  = ~\new_[3163]_ ;
  assign \new_[13880]_  = ~\new_[6483]_ ;
  assign \new_[13881]_  = ~\new_[7158]_ ;
  assign \new_[13882]_  = ~\new_[5765]_ ;
  assign \new_[13883]_  = ~\new_[3564]_ ;
  assign \new_[13884]_  = ~\new_[6087]_ ;
  assign \new_[13885]_  = ~\new_[3454]_ ;
  assign \new_[13886]_  = ~\new_[6718]_ ;
  assign \new_[13887]_  = ~\new_[3347]_ ;
  assign \new_[13888]_  = ~\new_[3697]_ ;
  assign \new_[13889]_  = ~\new_[5978]_ ;
  assign \new_[13890]_  = ~\new_[3325]_ ;
  assign \new_[13891]_  = ~\new_[6168]_ ;
  assign \new_[13892]_  = ~\new_[6342]_ ;
  assign \new_[13893]_  = ~\new_[3315]_ ;
  assign \new_[13894]_  = ~\new_[6265]_ ;
  assign \new_[13895]_  = ~\new_[4799]_ ;
  assign \new_[13896]_  = ~\new_[6311]_ ;
  assign \new_[13897]_  = ~\new_[6344]_ ;
  assign \new_[13898]_  = ~\new_[3719]_ ;
  assign \new_[13899]_  = ~\new_[3807]_ ;
  assign \new_[13900]_  = ~\new_[2339]_ ;
  assign \new_[13901]_  = ~\new_[8959]_ ;
  assign \new_[13902]_  = ~\new_[6309]_ ;
  assign \new_[13903]_  = ~\new_[6370]_ ;
  assign \new_[13904]_  = ~\new_[6303]_ ;
  assign \new_[13905]_  = ~\new_[6343]_ ;
  assign \new_[13906]_  = ~\new_[4953]_ ;
  assign \new_[13907]_  = ~\new_[6635]_ ;
  assign \new_[13908]_  = ~\new_[3031]_ ;
  assign \new_[13909]_  = ~\new_[3320]_ ;
  assign \new_[13910]_  = ~\new_[3633]_ ;
  assign \new_[13911]_  = ~\new_[4083]_ ;
  assign \new_[13912]_  = ~\new_[3889]_ ;
  assign \new_[13913]_  = ~\new_[6371]_ ;
  assign \new_[13914]_  = ~\new_[6563]_ ;
  assign \new_[13915]_  = ~\new_[6102]_ ;
  assign \new_[13916]_  = ~\new_[4848]_ ;
  assign \new_[13917]_  = ~\new_[2474]_ ;
  assign \new_[13918]_  = ~\new_[6528]_ ;
  assign \new_[13919]_  = ~\new_[2456]_ ;
  assign \new_[13920]_  = ~\new_[4741]_ ;
  assign \new_[13921]_  = ~\new_[4807]_ ;
  assign \new_[13922]_  = ~\new_[6285]_ ;
  assign \new_[13923]_  = ~\new_[6385]_ ;
  assign \new_[13924]_  = ~\new_[6287]_ ;
  assign \new_[13925]_  = ~\new_[7159]_ ;
  assign \new_[13926]_  = ~\new_[6552]_ ;
  assign \new_[13927]_  = ~\new_[2049]_ ;
  assign \new_[13928]_  = ~\new_[3468]_ ;
  assign \new_[13929]_  = ~\new_[3390]_ ;
  assign \new_[13930]_  = ~\new_[6246]_ ;
  assign \new_[13931]_  = ~\new_[3694]_ ;
  assign \new_[13932]_  = ~\new_[5129]_ ;
  assign \new_[13933]_  = ~\new_[3338]_ ;
  assign \new_[13934]_  = ~\new_[3326]_ ;
  assign \new_[13935]_  = ~\new_[3306]_ ;
  assign \new_[13936]_  = ~\new_[3791]_ ;
  assign \new_[13937]_  = ~\new_[2477]_ ;
  assign \new_[13938]_  = ~\new_[6363]_ ;
  assign \new_[13939]_  = ~\new_[3864]_ ;
  assign \new_[13940]_  = ~\new_[2210]_ ;
  assign \new_[13941]_  = ~\new_[6512]_ ;
  assign \new_[13942]_  = ~\new_[3974]_ ;
  assign \new_[13943]_  = ~\new_[3339]_ ;
  assign \new_[13944]_  = ~\new_[6033]_ ;
  assign \new_[13945]_  = ~\new_[6322]_ ;
  assign \new_[13946]_  = ~\new_[6006]_ ;
  assign \new_[13947]_  = ~\new_[6092]_ ;
  assign \new_[13948]_  = ~\new_[3298]_ ;
  assign \new_[13949]_  = ~\new_[7147]_ ;
  assign \new_[13950]_  = ~\new_[5754]_ ;
  assign \new_[13951]_  = ~\new_[3166]_ ;
  assign \new_[13952]_  = ~\new_[3708]_ ;
  assign \new_[13953]_  = ~\new_[2550]_ ;
  assign \new_[13954]_  = ~\new_[3721]_ ;
  assign \new_[13955]_  = ~\new_[3281]_ ;
  assign \new_[13956]_  = ~\new_[4843]_ ;
  assign \new_[13957]_  = ~\new_[3680]_ ;
  assign \new_[13958]_  = ~\new_[3288]_ ;
  assign \new_[13959]_  = ~\new_[3705]_ ;
  assign n9055 = ~\new_[5144]_ ;
  assign \new_[13961]_  = ~\new_[3343]_ ;
  assign \new_[13962]_  = ~\new_[6300]_ ;
  assign \new_[13963]_  = ~\new_[4789]_ ;
  assign \new_[13964]_  = ~\new_[5499]_ ;
  assign \new_[13965]_  = ~\new_[3131]_ ;
  assign \new_[13966]_  = ~\new_[3634]_ ;
  assign \new_[13967]_  = ~\new_[6315]_ ;
  assign \new_[13968]_  = ~\new_[6340]_ ;
  assign \new_[13969]_  = ~\new_[6385]_ ;
  assign \new_[13970]_  = ~\new_[3012]_ ;
  assign \new_[13971]_  = ~n8995;
  assign \new_[13972]_  = ~\new_[3728]_ ;
  assign \new_[13973]_  = ~\new_[6374]_ ;
  assign \new_[13974]_  = ~\wb_addr_i[6] ;
  assign \new_[13975]_  = ~\new_[2086]_ ;
  assign \new_[13976]_  = ~\new_[3302]_ ;
  assign \new_[13977]_  = ~\new_[2172]_ ;
  assign \new_[13978]_  = ~\new_[2872]_ ;
  assign \new_[13979]_  = ~\new_[3319]_ ;
  assign \new_[13980]_  = ~\new_[6004]_ ;
  assign \new_[13981]_  = ~\new_[6351]_ ;
  assign \new_[13982]_  = ~\new_[3485]_ ;
  assign \new_[13983]_  = ~\new_[3493]_ ;
  assign \new_[13984]_  = ~\new_[3682]_ ;
  assign \new_[13985]_  = ~\new_[6289]_ ;
  assign \new_[13986]_  = ~\new_[3816]_ ;
  assign \new_[13987]_  = ~\new_[2478]_ ;
  assign \new_[13988]_  = ~\new_[6016]_ ;
  assign \new_[13989]_  = ~\new_[6367]_ ;
  assign \new_[13990]_  = ~\new_[4641]_ ;
  assign \new_[13991]_  = ~\new_[3333]_ ;
  assign \new_[13992]_  = ~\new_[2082]_ ;
  assign \new_[13993]_  = ~\new_[4833]_ ;
  assign \new_[13994]_  = ~\new_[3524]_ ;
  assign \new_[13995]_  = ~\new_[6725]_ ;
  assign \new_[13996]_  = ~\new_[3614]_ ;
  assign \new_[13997]_  = ~\new_[4956]_ ;
  assign \new_[13998]_  = ~\new_[3322]_ ;
  assign \new_[13999]_  = ~\new_[4809]_ ;
  assign \new_[14000]_  = ~\new_[3029]_ ;
  assign \new_[14001]_  = ~\new_[6561]_ ;
  assign \new_[14002]_  = ~\new_[6211]_ ;
  assign \new_[14003]_  = ~\new_[3032]_ ;
  assign \new_[14004]_  = ~\new_[5757]_ ;
  assign \new_[14005]_  = ~\new_[4286]_ ;
  assign \new_[14006]_  = ~\new_[6160]_ ;
  assign \new_[14007]_  = ~\new_[3722]_ ;
  assign \new_[14008]_  = ~\new_[6734]_ ;
  assign \new_[14009]_  = ~\new_[6282]_ ;
  assign \new_[14010]_  = ~\new_[3799]_ ;
  assign \new_[14011]_  = ~\new_[3455]_ ;
  assign \new_[14012]_  = ~\new_[3866]_ ;
  assign \new_[14013]_  = ~\new_[4370]_ ;
  assign \new_[14014]_  = ~\new_[3285]_ ;
  assign \new_[14015]_  = ~\new_[5999]_ ;
  assign \new_[14016]_  = ~\new_[6328]_ ;
  assign \new_[14017]_  = ~\new_[6600]_ ;
  assign \new_[14018]_  = ~\new_[6020]_ ;
  assign \new_[14019]_  = ~\new_[4805]_ ;
  assign \new_[14020]_  = ~n8955;
  assign \new_[14021]_  = ~\new_[3700]_ ;
  assign \new_[14022]_  = ~\new_[3178]_ ;
  assign \new_[14023]_  = ~\new_[4080]_ ;
  assign \new_[14024]_  = ~\new_[3491]_ ;
  assign \new_[14025]_  = ~\new_[3968]_ ;
  assign \new_[14026]_  = ~\new_[6015]_ ;
  assign \new_[14027]_  = ~\new_[3501]_ ;
  assign \new_[14028]_  = ~\new_[6696]_ ;
  assign \new_[14029]_  = ~\new_[4844]_ ;
  assign \new_[14030]_  = ~\new_[3707]_ ;
  assign \new_[14031]_  = ~\new_[6850]_ ;
  assign \new_[14032]_  = ~\new_[6018]_ ;
  assign \new_[14033]_  = ~\new_[7160]_ ;
  assign \new_[14034]_  = ~\new_[7670]_ ;
  assign \new_[14035]_  = ~\new_[2093]_ ;
  assign \new_[14036]_  = ~\new_[3010]_ ;
  assign \new_[14037]_  = ~\new_[4822]_ ;
  assign \new_[14038]_  = ~\new_[7151]_ ;
  assign \new_[14039]_  = ~\new_[7198]_ ;
  assign n9050 = ~\new_[7572]_ ;
  assign \new_[14041]_  = ~\new_[3063]_ ;
  assign \new_[14042]_  = ~\new_[7150]_ ;
  assign \new_[14043]_  = ~\new_[6232]_ ;
  assign \new_[14044]_  = ~\new_[3732]_ ;
  assign \new_[14045]_  = ~\new_[3503]_ ;
  assign \new_[14046]_  = ~\new_[4780]_ ;
  assign \new_[14047]_  = ~\new_[6334]_ ;
  assign \new_[14048]_  = ~\new_[4079]_ ;
  assign \new_[14049]_  = ~\new_[6350]_ ;
  assign \new_[14050]_  = ~\new_[9645]_ ;
  assign \new_[14051]_  = ~\new_[4824]_ ;
  assign \new_[14052]_  = ~\new_[6853]_ ;
  assign \new_[14053]_  = ~\new_[4850]_ ;
  assign \new_[14054]_  = ~\new_[6491]_ ;
  assign \new_[14055]_  = ~\new_[3522]_ ;
  assign \new_[14056]_  = ~\new_[3520]_ ;
  assign \new_[14057]_  = ~\new_[6870]_ ;
  assign \new_[14058]_  = ~\new_[6017]_ ;
  assign \new_[14059]_  = ~\new_[6875]_ ;
  assign \new_[14060]_  = ~\new_[2990]_ ;
  assign \new_[14061]_  = ~\new_[8703]_ ;
  assign \new_[14062]_  = ~\new_[3425]_ ;
  assign \new_[14063]_  = ~\new_[6863]_ ;
  assign \new_[14064]_  = ~\new_[6295]_ ;
  assign \new_[14065]_  = ~\new_[3328]_ ;
  assign \new_[14066]_  = ~\new_[6352]_ ;
  assign \new_[14067]_  = ~\new_[6478]_ ;
  assign \new_[14068]_  = ~\new_[3416]_ ;
  assign \new_[14069]_  = ~\new_[6009]_ ;
  assign \new_[14070]_  = ~\new_[7291]_ ;
  assign \new_[14071]_  = ~\new_[2052]_ ;
  assign \new_[14072]_  = ~\new_[3676]_ ;
  assign \new_[14073]_  = ~\new_[6012]_ ;
  assign \new_[14074]_  = ~\new_[6607]_ ;
  assign \new_[14075]_  = ~\new_[3186]_ ;
  assign \new_[14076]_  = ~\new_[6597]_ ;
  assign \new_[14077]_  = ~\new_[2038]_ ;
  assign \new_[14078]_  = ~\new_[6283]_ ;
  assign \new_[14079]_  = ~\new_[7153]_ ;
  assign \new_[14080]_  = ~\new_[6316]_ ;
  assign \new_[14081]_  = ~\new_[6731]_ ;
  assign \new_[14082]_  = ~\new_[6275]_ ;
  assign \new_[14083]_  = ~\new_[3636]_ ;
  assign \new_[14084]_  = ~\new_[6236]_ ;
  assign \new_[14085]_  = ~\new_[3596]_ ;
  assign \new_[14086]_  = ~\new_[4847]_ ;
  assign \new_[14087]_  = ~\new_[6354]_ ;
  assign \new_[14088]_  = ~\new_[4837]_ ;
  assign \new_[14089]_  = ~\new_[3024]_ ;
  assign \new_[14090]_  = ~\new_[3659]_ ;
  assign \new_[14091]_  = ~\new_[6511]_ ;
  assign \new_[14092]_  = ~\new_[3488]_ ;
  assign \new_[14093]_  = ~\new_[3103]_ ;
  assign \new_[14094]_  = ~\new_[2085]_ ;
  assign \new_[14095]_  = ~\new_[6325]_ ;
  assign \new_[14096]_  = ~\new_[3465]_ ;
  assign \new_[14097]_  = ~\new_[3346]_ ;
  assign \new_[14098]_  = ~\new_[6248]_ ;
  assign \new_[14099]_  = ~\new_[7161]_ ;
  assign \new_[14100]_  = ~\new_[2040]_ ;
  assign \new_[14101]_  = ~\new_[6157]_ ;
  assign \new_[14102]_  = ~\new_[6871]_ ;
  assign \new_[14103]_  = ~\new_[7177]_ ;
  assign \new_[14104]_  = ~\new_[7179]_ ;
  assign \new_[14105]_  = ~\new_[4617]_ ;
  assign \new_[14106]_  = ~n8990;
  assign \new_[14107]_  = ~\new_[6362]_ ;
  assign \new_[14108]_  = ~\new_[6345]_ ;
  assign \new_[14109]_  = ~\new_[7205]_ ;
  assign \new_[14110]_  = ~\new_[6730]_ ;
  assign \new_[14111]_  = ~\new_[2089]_ ;
  assign \new_[14112]_  = ~\new_[3179]_ ;
  assign \new_[14113]_  = ~\new_[3494]_ ;
  assign \new_[14114]_  = ~\new_[3512]_ ;
  assign \new_[14115]_  = ~\new_[2046]_ ;
  assign n9040 = ~\new_[7718]_ ;
  assign \new_[14117]_  = ~\new_[3348]_ ;
  assign \new_[14118]_  = ~\new_[7130]_ ;
  assign \new_[14119]_  = ~\new_[6697]_ ;
  assign \new_[14120]_  = ~\new_[6326]_ ;
  assign \new_[14121]_  = ~\new_[6296]_ ;
  assign \new_[14122]_  = ~\new_[3332]_ ;
  assign \new_[14123]_  = ~\new_[6559]_ ;
  assign \new_[14124]_  = ~\new_[4832]_ ;
  assign \new_[14125]_  = ~\new_[6306]_ ;
  assign \new_[14126]_  = ~n8985;
  assign \new_[14127]_  = ~\new_[4161]_ ;
  assign \new_[14128]_  = ~\new_[6337]_ ;
  assign \new_[14129]_  = ~\new_[4836]_ ;
  assign \new_[14130]_  = ~\new_[7297]_ ;
  assign \new_[14131]_  = ~\new_[6868]_ ;
  assign \new_[14132]_  = ~\new_[3167]_ ;
  assign \new_[14133]_  = ~\new_[6846]_ ;
  assign \new_[14134]_  = ~\new_[3422]_ ;
  assign \new_[14135]_  = ~\new_[2452]_ ;
  assign \new_[14136]_  = ~\new_[3730]_ ;
  assign \new_[14137]_  = ~\new_[3432]_ ;
  assign \new_[14138]_  = ~\new_[3170]_ ;
  assign \new_[14139]_  = ~\new_[6166]_ ;
  assign \new_[14140]_  = ~\new_[3350]_ ;
  assign \new_[14141]_  = ~\new_[4072]_ ;
  assign \new_[14142]_  = ~\new_[7154]_ ;
  assign \new_[14143]_  = ~\new_[3165]_ ;
  assign \new_[14144]_  = ~\new_[3734]_ ;
  assign \new_[14145]_  = ~\new_[3499]_ ;
  assign \new_[14146]_  = ~\new_[2209]_ ;
  assign \new_[14147]_  = ~\new_[3313]_ ;
  assign \new_[14148]_  = ~\new_[3292]_ ;
  assign \new_[14149]_  = ~\new_[6238]_ ;
  assign \new_[14150]_  = ~\new_[6099]_ ;
  assign \new_[14151]_  = ~\new_[6867]_ ;
  assign \new_[14152]_  = ~\new_[4245]_ ;
  assign \new_[14153]_  = ~\new_[7148]_ ;
  assign \new_[14154]_  = ~\new_[3489]_ ;
  assign \new_[14155]_  = ~\new_[6475]_ ;
  assign \new_[14156]_  = ~\new_[5145]_ ;
  assign \new_[14157]_  = ~\new_[7152]_ ;
  assign \new_[14158]_  = ~\new_[3183]_ ;
  assign \new_[14159]_  = ~\new_[3459]_ ;
  assign \new_[14160]_  = ~\new_[6100]_ ;
  assign \new_[14161]_  = ~\new_[6383]_ ;
  assign \new_[14162]_  = ~\new_[3442]_ ;
  assign \new_[14163]_  = ~\new_[3030]_ ;
  assign \new_[14164]_  = ~\new_[6727]_ ;
  assign \new_[14165]_  = ~\new_[3295]_ ;
  assign \new_[14166]_  = ~\new_[3160]_ ;
  assign \new_[14167]_  = ~\new_[5994]_ ;
  assign \new_[14168]_  = ~\new_[3334]_ ;
  assign \new_[14169]_  = ~\new_[4098]_ ;
  assign \new_[14170]_  = ~\new_[3171]_ ;
  assign \new_[14171]_  = ~\new_[9405]_ ;
  assign \new_[14172]_  = ~\new_[6278]_ ;
  assign \new_[14173]_  = ~\new_[3296]_ ;
  assign \new_[14174]_  = ~\new_[2472]_ ;
  assign \new_[14175]_  = ~\new_[3331]_ ;
  assign \new_[14176]_  = ~\new_[6336]_ ;
  assign \new_[14177]_  = ~\new_[3631]_ ;
  assign \new_[14178]_  = ~\new_[3490]_ ;
  assign \new_[14179]_  = ~\new_[6330]_ ;
  assign \new_[14180]_  = ~\new_[7202]_ ;
  assign \new_[14181]_  = ~\new_[6332]_ ;
  assign \new_[14182]_  = ~\new_[3515]_ ;
  assign \new_[14183]_  = ~\new_[3324]_ ;
  assign \new_[14184]_  = ~\new_[3300]_ ;
  assign \new_[14185]_  = ~\new_[3041]_ ;
  assign \new_[14186]_  = ~\new_[4781]_ ;
  assign \new_[14187]_  = ~\new_[2318]_ ;
  assign \new_[14188]_  = ~\new_[3462]_ ;
  assign \new_[14189]_  = ~\new_[3717]_ ;
  assign \new_[14190]_  = ~\new_[3448]_ ;
  assign \new_[14191]_  = ~\new_[2114]_ ;
  assign \new_[14192]_  = ~\new_[6203]_ ;
  assign \new_[14193]_  = ~\new_[4181]_ ;
  assign \new_[14194]_  = ~\new_[6088]_ ;
  assign \new_[14195]_  = ~\new_[6252]_ ;
  assign \new_[14196]_  = ~\new_[3191]_ ;
  assign \new_[14197]_  = ~\new_[6369]_ ;
  assign \new_[14198]_  = ~\new_[3161]_ ;
  assign \new_[14199]_  = ~\new_[6567]_ ;
  assign \new_[14200]_  = ~\new_[4802]_ ;
  assign \new_[14201]_  = ~\new_[3440]_ ;
  assign \new_[14202]_  = ~\new_[3335]_ ;
  assign \new_[14203]_  = ~\new_[4091]_ ;
  assign \new_[14204]_  = ~\new_[4785]_ ;
  assign \new_[14205]_  = ~\new_[2873]_ ;
  assign \new_[14206]_  = ~\new_[3740]_ ;
  assign \new_[14207]_  = ~\new_[3451]_ ;
  assign \new_[14208]_  = ~\new_[6754]_ ;
  assign \new_[14209]_  = ~\new_[3158]_ ;
  assign \new_[14210]_  = ~\new_[6308]_ ;
  assign \new_[14211]_  = ~\new_[3026]_ ;
  assign \new_[14212]_  = ~\new_[3303]_ ;
  assign \new_[14213]_  = ~\new_[3671]_ ;
  assign \new_[14214]_  = ~\new_[6364]_ ;
  assign \new_[14215]_  = ~\new_[2064]_ ;
  assign \new_[14216]_  = ~\new_[3101]_ ;
  assign \new_[14217]_  = ~\new_[6735]_ ;
  assign \new_[14218]_  = ~\new_[7301]_ ;
  assign \new_[14219]_  = ~\new_[9424]_ ;
  assign \new_[14220]_  = ~\new_[3496]_ ;
  assign \new_[14221]_  = ~\new_[6200]_ ;
  assign \new_[14222]_  = ~\new_[3355]_ ;
  assign \new_[14223]_  = ~\new_[6307]_ ;
  assign \new_[14224]_  = ~\new_[6866]_ ;
  assign \new_[14225]_  = ~\new_[2053]_ ;
  assign \new_[14226]_  = ~\new_[6233]_ ;
  assign \new_[14227]_  = ~\new_[3511]_ ;
  assign \new_[14228]_  = ~\new_[6172]_ ;
  assign \new_[14229]_  = ~\new_[6373]_ ;
  assign \new_[14230]_  = ~\new_[11698]_ ;
  assign \new_[14231]_  = ~\new_[6882]_ ;
  assign \new_[14232]_  = ~\new_[7163]_ ;
  assign \new_[14233]_  = ~\new_[3624]_ ;
  assign \new_[14234]_  = ~\new_[4085]_ ;
  assign \new_[14235]_  = ~\new_[3513]_ ;
  assign \new_[14236]_  = ~\new_[7286]_ ;
  assign \new_[14237]_  = ~\new_[4287]_ ;
  assign \new_[14238]_  = ~\new_[6539]_ ;
  assign \new_[14239]_  = ~\new_[6550]_ ;
  assign \new_[14240]_  = ~\new_[3424]_ ;
  assign \new_[14241]_  = ~\new_[3865]_ ;
  assign \new_[14242]_  = ~\new_[2042]_ ;
  assign \new_[14243]_  = ~\new_[6601]_ ;
  assign \new_[14244]_  = ~\new_[7310]_ ;
  assign \new_[14245]_  = ~\new_[5125]_ ;
  assign \new_[14246]_  = ~\new_[6209]_ ;
  assign \new_[14247]_  = ~\new_[4810]_ ;
  assign \new_[14248]_  = ~\new_[3294]_ ;
  assign \new_[14249]_  = ~\new_[3190]_ ;
  assign \new_[14250]_  = ~\new_[3516]_ ;
  assign \new_[14251]_  = ~\new_[11431]_ ;
  assign \new_[14252]_  = ~\new_[6327]_ ;
  assign \new_[14253]_  = ~\new_[4086]_ ;
  assign \new_[14254]_  = ~\new_[6384]_ ;
  assign \new_[14255]_  = ~\new_[3497]_ ;
  assign n9075 = ~\new_[7673]_ ;
  assign \new_[14257]_  = ~\new_[6375]_ ;
  assign \new_[14258]_  = ~\new_[6103]_ ;
  assign \new_[14259]_  = ~\new_[6377]_ ;
  assign \new_[14260]_  = ~\new_[6838]_ ;
  assign \new_[14261]_  = ~\new_[4685]_ ;
  assign \new_[14262]_  = ~\new_[4082]_ ;
  assign \new_[14263]_  = ~\new_[6598]_ ;
  assign \new_[14264]_  = ~\new_[2457]_ ;
  assign \new_[14265]_  = ~\new_[7302]_ ;
  assign n9045 = ~\new_[5243]_ ;
  assign \new_[14267]_  = ~\new_[3356]_ ;
  assign \new_[14268]_  = ~\new_[3461]_ ;
  assign \new_[14269]_  = ~\new_[14340]_ ;
  assign \new_[14270]_  = \new_[8226]_ ;
  assign \new_[14271]_  = ~\new_[14368]_ ;
  assign \new_[14272]_  = ~\new_[14349]_ ;
  assign \new_[14273]_  = \new_[14315]_  | \new_[14317]_ ;
  assign \new_[14274]_  = ~\new_[14310]_ ;
  assign \new_[14275]_  = ~\new_[14312]_ ;
  assign \new_[14276]_  = \new_[14311]_ ;
  assign \new_[14277]_  = \new_[5970]_  & \new_[2991]_ ;
  assign \new_[14278]_  = \new_[14279]_  | \new_[5349]_ ;
  assign \new_[14279]_  = ~\new_[14341]_  & (~\new_[14280]_  | ~\new_[14281]_ );
  assign \new_[14280]_  = \new_[14640]_  | \new_[7467]_ ;
  assign \new_[14281]_  = ~\new_[2961]_  | ~\new_[14640]_  | ~\new_[14635]_ ;
  assign \new_[14282]_  = (~\new_[6210]_  & ~\new_[14640]_  & ~\new_[9506]_ ) | (~\new_[5937]_  & ~\new_[6231]_  & ~\new_[6699]_ );
  assign \new_[14283]_  = ~\new_[14341]_ ;
  assign \new_[14284]_  = \new_[14285]_  & \new_[14288]_ ;
  assign \new_[14285]_  = ~\new_[14287]_  | ~\new_[14286]_  | ~\new_[2195]_ ;
  assign \new_[14286]_  = ~\new_[2184]_  | ~\new_[2435]_ ;
  assign \new_[14287]_  = ~\new_[2369]_ ;
  assign \new_[14288]_  = ~n9145 & (~\new_[2489]_  | ~\new_[14289]_ );
  assign \new_[14289]_  = \new_[4513]_  | \new_[2546]_ ;
  assign \new_[14290]_  = ~\new_[2369]_  & ~\new_[14291]_ ;
  assign \new_[14291]_  = ~\new_[14286]_ ;
  assign \new_[14292]_  = ~\new_[14289]_ ;
  assign \new_[14293]_  = ~\new_[13118]_  | ~\new_[14538]_ ;
  assign \new_[14294]_  = ~\new_[7438]_  | ~\new_[7439]_  | ~\new_[14295]_ ;
  assign \new_[14295]_  = \new_[14329]_  & \new_[12932]_ ;
  assign \new_[14296]_  = ~\new_[7409]_ ;
  assign \new_[14297]_  = (~\new_[13646]_  | ~\new_[14422]_ ) & (~\new_[8602]_  | ~\new_[12565]_ );
  assign \new_[14298]_  = ~\new_[14825]_ ;
  assign \new_[14299]_  = ~\new_[5151]_ ;
  assign \new_[14300]_  = \new_[14367]_ ;
  assign \new_[14301]_  = ~\new_[14689]_ ;
  assign \new_[14302]_  = \new_[14640]_ ;
  assign \new_[14303]_  = \new_[14304]_  ^ \new_[14305]_ ;
  assign \new_[14304]_  = \new_[12122]_  ? \new_[2271]_  : \new_[11480]_ ;
  assign \new_[14305]_  = \new_[14306]_  ? \new_[14569]_  : \new_[14307]_ ;
  assign \new_[14306]_  = ~\new_[14307]_ ;
  assign \new_[14307]_  = \new_[14308]_ ;
  assign \new_[14308]_  = \new_[4767]_  ^ \new_[4766]_ ;
  assign \new_[14309]_  = ~\new_[14713]_ ;
  assign \new_[14310]_  = ~\new_[14311]_  | ~\new_[14312]_ ;
  assign \new_[14311]_  = (~\new_[4676]_  | ~\new_[14530]_ ) & (~\new_[14313]_  | ~\new_[4609]_ );
  assign \new_[14312]_  = (~\new_[14530]_  & ~\new_[4845]_ ) | (~\new_[14313]_  & ~\new_[4690]_ );
  assign \new_[14313]_  = ~\new_[14530]_ ;
  assign \new_[14314]_  = ~\new_[14461]_ ;
  assign \new_[14315]_  = \new_[14316]_ ;
  assign \new_[14316]_  = ~\new_[12654]_  | ~\new_[2192]_ ;
  assign \new_[14317]_  = ~\new_[2176]_ ;
  assign \new_[14318]_  = ~\new_[5075]_  & ~\new_[2464]_ ;
  assign \new_[14319]_  = ~\new_[14375]_ ;
  assign \new_[14320]_  = ~\new_[14377]_  | ~\new_[14378]_ ;
  assign \new_[14321]_  = \new_[14322]_  | \new_[10715]_ ;
  assign \new_[14322]_  = ~\new_[14325]_  | ~\new_[14323]_  | ~\new_[14324]_ ;
  assign \new_[14323]_  = ~\new_[14282]_ ;
  assign \new_[14324]_  = ~\new_[14302]_  | (~\new_[14277]_  & ~\new_[5938]_ );
  assign \new_[14325]_  = ~\new_[14278]_ ;
  assign \new_[14326]_  = \new_[14322]_ ;
  assign \new_[14327]_  = ~\new_[14374]_  | ~\new_[14328]_ ;
  assign \new_[14328]_  = ~\new_[2290]_  & (~\new_[2325]_  | ~\new_[14379]_ );
  assign \new_[14329]_  = ~\new_[14330]_  | ~\new_[14788]_ ;
  assign \new_[14330]_  = \new_[4837]_  ? \new_[14531]_  : \new_[4814]_ ;
  assign \new_[14331]_  = ~\new_[14533]_ ;
  assign \new_[14332]_  = ~\new_[14331]_ ;
  assign \new_[14333]_  = ~\new_[14335]_  | ~\new_[14334]_  | ~\new_[14408]_ ;
  assign \new_[14334]_  = ~\new_[14671]_  | ~\new_[2567]_  | ~\new_[9036]_ ;
  assign \new_[14335]_  = ~\new_[4883]_ ;
  assign \new_[14336]_  = ~\new_[14337]_ ;
  assign \new_[14337]_  = ~\new_[4651]_  | ~\new_[14829]_ ;
  assign \new_[14338]_  = ~\new_[14408]_  | ~\new_[14337]_  | ~\new_[14334]_ ;
  assign \new_[14339]_  = ~\new_[14484]_  | ~\new_[8626]_ ;
  assign \new_[14340]_  = ~\new_[14590]_ ;
  assign \new_[14341]_  = ~\new_[14344]_  | ~\new_[14733]_  | ~\new_[14390]_ ;
  assign \new_[14342]_  = ~\new_[5486]_ ;
  assign \new_[14343]_  = \new_[13257]_  & \new_[13882]_ ;
  assign \new_[14344]_  = ~\new_[11923]_  | ~\new_[10449]_ ;
  assign \new_[14345]_  = \new_[14733]_ ;
  assign \new_[14346]_  = \new_[14390]_ ;
  assign \new_[14347]_  = \new_[14734]_  & \new_[14739]_ ;
  assign \new_[14348]_  = ~\new_[6083]_ ;
  assign \new_[14349]_  = ~\new_[14712]_ ;
  assign \new_[14350]_  = ~\new_[2579]_  & ~\new_[14351]_ ;
  assign \new_[14351]_  = ~\new_[2707]_ ;
  assign \new_[14352]_  = \new_[2682]_  & \new_[2706]_ ;
  assign \new_[14353]_  = ~\new_[2578]_ ;
  assign \new_[14354]_  = ~\new_[2711]_ ;
  assign \new_[14355]_  = ~\new_[2713]_ ;
  assign \new_[14356]_  = ~\new_[14355]_  & ~\new_[14354]_ ;
  assign \new_[14357]_  = ~\new_[2581]_  & ~\new_[2580]_ ;
  assign \new_[14358]_  = \new_[2712]_  & \new_[2684]_ ;
  assign \new_[14359]_  = ~\new_[14360]_  | ~\new_[14365]_ ;
  assign \new_[14360]_  = ~\new_[14361]_  | ~\new_[14363]_ ;
  assign \new_[14361]_  = ~\new_[14685]_  | ~\new_[14362]_ ;
  assign \new_[14362]_  = ~\new_[14444]_  & ~\new_[14667]_ ;
  assign \new_[14363]_  = ~\new_[14364]_ ;
  assign \new_[14364]_  = ~\new_[2410]_  | (~\new_[2427]_  & ~\new_[14444]_ );
  assign \new_[14365]_  = \new_[14630]_  & \new_[14366]_ ;
  assign \new_[14366]_  = ~\new_[2367]_  & ~\new_[2363]_ ;
  assign \new_[14367]_  = ~\new_[14685]_ ;
  assign \new_[14368]_  = ~\new_[14549]_ ;
  assign \new_[14369]_  = \new_[14532]_  & \new_[4840]_ ;
  assign \new_[14370]_  = \new_[4839]_  & \new_[14532]_ ;
  assign \new_[14371]_  = ~\new_[14673]_  | ~\new_[11378]_ ;
  assign \new_[14372]_  = ~\new_[14673]_  | ~\new_[11399]_ ;
  assign \new_[14373]_  = ~\new_[14559]_ ;
  assign \new_[14374]_  = ~\new_[14379]_  | ~\new_[14375]_  | ~\new_[14512]_ ;
  assign \new_[14375]_  = ~\new_[14378]_  | ~\new_[14376]_  | ~\new_[14377]_ ;
  assign \new_[14376]_  = ~\new_[14318]_  | ~\new_[14689]_  | ~\new_[2407]_ ;
  assign \new_[14377]_  = \new_[2408]_  | \new_[14301]_ ;
  assign \new_[14378]_  = ~\new_[5151]_  | ~\new_[14825]_ ;
  assign \new_[14379]_  = ~\new_[2367]_  & ~\new_[14444]_ ;
  assign \new_[14380]_  = ~\new_[8810]_  & ~\new_[4788]_ ;
  assign \new_[14381]_  = ~\new_[13658]_  | ~\new_[13690]_ ;
  assign \new_[14382]_  = ~\new_[14388]_  | ~\new_[14383]_  | ~\new_[14384]_ ;
  assign \new_[14383]_  = ~\new_[10104]_ ;
  assign \new_[14384]_  = \new_[14385]_  & \new_[14387]_ ;
  assign \new_[14385]_  = ~\new_[14386]_ ;
  assign \new_[14386]_  = ~\new_[12617]_  | ~\new_[14738]_ ;
  assign \new_[14387]_  = ~\new_[13469]_  & ~\new_[14167]_ ;
  assign \new_[14388]_  = ~\new_[12716]_ ;
  assign \new_[14389]_  = ~\new_[13588]_  | ~\new_[10449]_  | ~\new_[12606]_ ;
  assign \new_[14390]_  = ~\new_[12570]_  | ~\new_[10076]_  | ~\new_[14343]_ ;
  assign \new_[14391]_  = ~\new_[10104]_  & ~\new_[12716]_ ;
  assign \new_[14392]_  = ~\new_[2543]_  & ~\new_[14832]_ ;
  assign \new_[14393]_  = ~\new_[14394]_  | ~\new_[14516]_ ;
  assign \new_[14394]_  = ~\new_[14392]_ ;
  assign \new_[14395]_  = ~\new_[14396]_  | ~\new_[14404]_ ;
  assign \new_[14396]_  = ~\new_[14397]_ ;
  assign \new_[14397]_  = ~\new_[14398]_  | ~\new_[14403]_ ;
  assign \new_[14398]_  = ~\new_[14399]_  | ~\new_[14401]_ ;
  assign \new_[14399]_  = ~\new_[14400]_ ;
  assign \new_[14400]_  = ~\new_[2705]_  | ~\new_[14352]_  | ~\new_[14350]_  | ~\new_[14353]_ ;
  assign \new_[14401]_  = ~\new_[14402]_ ;
  assign \new_[14402]_  = ~\new_[14358]_  | ~\new_[14356]_  | ~\new_[14357]_ ;
  assign \new_[14403]_  = ~\new_[14402]_  | ~\new_[14400]_ ;
  assign \new_[14404]_  = ~\new_[14405]_ ;
  assign \new_[14405]_  = \new_[2174]_  ^ \new_[13845]_ ;
  assign \new_[14406]_  = ~\new_[14403]_  | ~\new_[14398]_ ;
  assign \new_[14407]_  = ~\new_[14399]_ ;
  assign \new_[14408]_  = ~\new_[2876]_  | ~\new_[14671]_  | ~\new_[14409]_ ;
  assign \new_[14409]_  = ~\new_[14610]_ ;
  assign \new_[14410]_  = ~\new_[14411]_ ;
  assign \new_[14411]_  = ~rst_i | ~\new_[14412]_ ;
  assign \new_[14412]_  = \new_[14413]_  | \new_[4600]_ ;
  assign \new_[14413]_  = \new_[14414]_  | \new_[5745]_ ;
  assign \new_[14414]_  = ~\new_[6464]_  | ~\new_[12137]_  | ~\new_[14415]_  | ~\new_[14416]_ ;
  assign \new_[14415]_  = ~\new_[12222]_  & ~\new_[11699]_ ;
  assign \new_[14416]_  = ~\new_[12221]_  & ~\new_[12465]_ ;
  assign \new_[14417]_  = ~\new_[14410]_ ;
  assign \new_[14418]_  = \new_[14419]_  & \new_[14420]_ ;
  assign \new_[14419]_  = ~\new_[4620]_  | ~\new_[9464]_  | ~\new_[9748]_ ;
  assign \new_[14420]_  = ~\new_[9467]_  | ~\new_[4799]_  | ~\new_[9740]_ ;
  assign \new_[14421]_  = ~\new_[14422]_  | ~\new_[14423]_ ;
  assign \new_[14422]_  = ~\new_[9464]_  | ~\new_[9748]_ ;
  assign \new_[14423]_  = ~\new_[9467]_  | ~\new_[9740]_ ;
  assign \new_[14424]_  = ~\new_[13646]_  | ~\new_[13895]_ ;
  assign \new_[14425]_  = ~\new_[14370]_ ;
  assign \new_[14426]_  = ~\new_[14531]_  | ~\new_[4816]_ ;
  assign \new_[14427]_  = \new_[14425]_  & \new_[14426]_ ;
  assign \new_[14428]_  = ~\new_[2524]_ ;
  assign \new_[14429]_  = \new_[2795]_  | \new_[14430]_ ;
  assign \new_[14430]_  = \new_[14431]_  | \new_[9910]_ ;
  assign \new_[14431]_  = \new_[11775]_  | \new_[10460]_ ;
  assign n1105 = ~\new_[14429]_ ;
  assign \new_[14433]_  = \new_[14434]_  ? \new_[14436]_  : \new_[14435]_ ;
  assign \new_[14434]_  = ~\new_[14653]_  & ~\new_[2488]_ ;
  assign \new_[14435]_  = ~\new_[14434]_ ;
  assign \new_[14436]_  = ~\new_[14437]_  | ~\new_[14438]_ ;
  assign \new_[14437]_  = ~\new_[2246]_  | ~\new_[14327]_ ;
  assign \new_[14438]_  = ~\new_[2293]_  & (~\new_[2292]_  | ~\new_[2294]_ );
  assign \new_[14439]_  = ~\new_[14440]_  & ~\new_[14442]_ ;
  assign \new_[14440]_  = ~\new_[14441]_  | ~\new_[2692]_ ;
  assign \new_[14441]_  = ~\new_[2842]_  | ~\new_[10633]_ ;
  assign \new_[14442]_  = ~\new_[14443]_  | ~\new_[2691]_ ;
  assign \new_[14443]_  = ~\new_[14824]_  | ~\new_[10358]_ ;
  assign \new_[14444]_  = ~\new_[5248]_  & ~\new_[14445]_ ;
  assign \new_[14445]_  = ~\new_[14447]_  | (~\new_[14446]_  & ~\new_[14829]_ );
  assign \new_[14446]_  = ~\new_[9559]_  & (~\new_[2633]_  | ~\new_[14610]_ );
  assign \new_[14447]_  = ~\new_[14829]_  | ~\new_[4620]_ ;
  assign \new_[14448]_  = ~\new_[14200]_  & ~\new_[14449]_ ;
  assign \new_[14449]_  = ~\new_[9722]_ ;
  assign \new_[14450]_  = ~\new_[14451]_  | ~\new_[8927]_ ;
  assign \new_[14451]_  = ~\new_[9465]_  | ~\new_[9722]_ ;
  assign \new_[14452]_  = ~\new_[14200]_  | ~\new_[14453]_ ;
  assign \new_[14453]_  = ~\new_[4651]_ ;
  assign \new_[14454]_  = ~\new_[14455]_  & ~\new_[14456]_ ;
  assign \new_[14455]_  = ~\new_[2677]_  | ~\new_[14372]_ ;
  assign \new_[14456]_  = ~\new_[14457]_  | ~\new_[14458]_ ;
  assign \new_[14457]_  = ~\new_[14721]_  | ~\new_[11083]_ ;
  assign \new_[14458]_  = ~\new_[14557]_  | ~\new_[11346]_ ;
  assign \new_[14459]_  = ~\new_[2734]_ ;
  assign \new_[14460]_  = ~\new_[2801]_  | ~\new_[2636]_ ;
  assign \new_[14461]_  = ~\new_[14460]_ ;
  assign \new_[14462]_  = \new_[14588]_  & \new_[14589]_ ;
  assign \new_[14463]_  = ~\new_[5087]_  | (~\new_[4755]_  & ~\new_[5085]_ );
  assign \new_[14464]_  = ~\new_[14468]_  & (~\new_[14465]_  | ~\new_[14466]_ );
  assign \new_[14465]_  = ~\new_[3765]_  | ~\new_[5082]_ ;
  assign \new_[14466]_  = ~\new_[5083]_  & ~\new_[14467]_ ;
  assign \new_[14467]_  = \new_[5084]_ ;
  assign \new_[14468]_  = ~\new_[14470]_  | (~\new_[14467]_  & ~\new_[14469]_ );
  assign \new_[14469]_  = \new_[5081]_ ;
  assign \new_[14470]_  = ~\new_[5085]_  & ~\new_[4764]_ ;
  assign \new_[14471]_  = ~\new_[14472]_  | ~\new_[14473]_ ;
  assign \new_[14472]_  = ~\new_[14467]_  & (~\new_[14469]_  | ~\new_[5083]_ );
  assign \new_[14473]_  = ~\new_[5082]_  | ~\new_[3765]_  | ~\new_[14469]_ ;
  assign \new_[14474]_  = ~\new_[14476]_  | (~\new_[14475]_  & ~\new_[8007]_ );
  assign \new_[14475]_  = \new_[8008]_  | \new_[6174]_ ;
  assign \new_[14476]_  = ~\new_[14480]_  & (~\new_[14477]_  | ~\new_[14479]_ );
  assign \new_[14477]_  = ~\new_[14478]_  & (~\new_[8600]_  | ~\new_[4651]_ );
  assign \new_[14478]_  = \new_[14448]_  & \new_[9465]_ ;
  assign \new_[14479]_  = ~\new_[14587]_  & ~\new_[4801]_ ;
  assign \new_[14480]_  = ~\new_[14481]_  | ~\new_[14482]_ ;
  assign \new_[14481]_  = ~\new_[7410]_ ;
  assign \new_[14482]_  = (~\new_[14453]_  | ~\new_[8927]_ ) & (~\new_[14451]_  | ~\new_[12591]_ );
  assign \new_[14483]_  = ~\new_[4882]_ ;
  assign \new_[14484]_  = ~\new_[14663]_ ;
  assign \new_[14485]_  = ~\new_[4702]_ ;
  assign \new_[14486]_  = ~\new_[4793]_ ;
  assign \new_[14487]_  = ~\new_[14488]_  | ~\new_[14492]_ ;
  assign \new_[14488]_  = ~\new_[14490]_  & (~\new_[4006]_  | ~\new_[14489]_ );
  assign \new_[14489]_  = \new_[5090]_  & \new_[5088]_ ;
  assign \new_[14490]_  = ~\new_[14491]_ ;
  assign \new_[14491]_  = ~\new_[5095]_  & (~\new_[5094]_  | ~\new_[5090]_ );
  assign \new_[14492]_  = ~\new_[14493]_  | (~\new_[14464]_  & ~\new_[14463]_ );
  assign \new_[14493]_  = \new_[14494]_  & \new_[14489]_ ;
  assign \new_[14494]_  = \new_[4757]_  & \new_[5089]_ ;
  assign \new_[14495]_  = ~\new_[14464]_  & ~\new_[14463]_ ;
  assign n880 = ~\new_[14497]_  | ~rst_i;
  assign \new_[14497]_  = ~\new_[14501]_  & (~\new_[14498]_  | ~n1240);
  assign \new_[14498]_  = ~\new_[14499]_ ;
  assign \new_[14499]_  = \new_[14429]_  & \new_[14428]_ ;
  assign n1240 = \new_[14539]_  ? \new_[3001]_  : \new_[4615]_ ;
  assign \new_[14501]_  = ~\new_[14498]_  & ~\new_[14502]_ ;
  assign \new_[14502]_  = ~\new_[9088]_  & (~\new_[14637]_  | ~\new_[2342]_ );
  assign \new_[14503]_  = ~rst_i;
  assign \new_[14504]_  = \new_[14648]_  & \new_[14704]_ ;
  assign \new_[14505]_  = ~\new_[14631]_  & ~\new_[14506]_ ;
  assign \new_[14506]_  = ~\new_[14729]_ ;
  assign \new_[14507]_  = ~\new_[14529]_ ;
  assign \new_[14508]_  = ~\new_[4923]_ ;
  assign \new_[14509]_  = ~\new_[14677]_  | ~\new_[14679]_  | ~\new_[14678]_ ;
  assign \new_[14510]_  = ~\new_[14511]_  | ~\new_[14373]_ ;
  assign \new_[14511]_  = ~\new_[14703]_ ;
  assign \new_[14512]_  = ~\new_[14698]_  & ~\new_[14667]_ ;
  assign \new_[14513]_  = ~\new_[14514]_ ;
  assign \new_[14514]_  = ~\new_[4514]_  & ~\new_[14515]_ ;
  assign \new_[14515]_  = \new_[14829]_  & \new_[4798]_ ;
  assign \new_[14516]_  = ~\new_[14515]_ ;
  assign \new_[14517]_  = ~\new_[14518]_  | ~\new_[14522]_ ;
  assign \new_[14518]_  = ~\new_[14519]_  | ~\new_[14521]_ ;
  assign \new_[14519]_  = ~\new_[14520]_ ;
  assign \new_[14520]_  = ~\new_[5088]_  | ~\new_[5089]_  | ~\new_[4757]_  | ~\new_[4754]_ ;
  assign \new_[14521]_  = ~\new_[4230]_  | ~\new_[3563]_  | ~\new_[3554]_ ;
  assign \new_[14522]_  = \new_[14523]_  & \new_[14524]_ ;
  assign \new_[14523]_  = ~\new_[5094]_  & (~\new_[5093]_  | ~\new_[5088]_ );
  assign \new_[14524]_  = ~\new_[14525]_  | ~\new_[14526]_ ;
  assign \new_[14525]_  = \new_[5092]_  | \new_[4455]_ ;
  assign \new_[14526]_  = \new_[5089]_  & \new_[5088]_ ;
  assign \new_[14527]_  = ~\new_[14526]_ ;
  assign \new_[14528]_  = ~\new_[4757]_  | ~\new_[4754]_ ;
  assign \new_[14529]_  = (~\new_[4819]_  | ~\new_[14530]_ ) & (~\new_[14537]_  | ~\new_[4842]_ );
  assign \new_[14530]_  = \new_[14531]_ ;
  assign \new_[14531]_  = ~\new_[14532]_ ;
  assign \new_[14532]_  = ~\new_[14533]_ ;
  assign \new_[14533]_  = ~\new_[14534]_ ;
  assign \new_[14534]_  = ~\new_[14535]_  | ~\new_[14536]_ ;
  assign \new_[14535]_  = ~\new_[14484]_  | ~\new_[8626]_ ;
  assign \new_[14536]_  = ~\new_[14663]_  | ~\new_[14380]_  | ~\new_[14381]_ ;
  assign \new_[14537]_  = ~\new_[14531]_ ;
  assign \new_[14538]_  = ~\new_[14545]_  | (~\new_[14539]_  & ~\new_[14540]_ );
  assign \new_[14539]_  = \new_[4864]_  ? \new_[9307]_  : \new_[4619]_ ;
  assign \new_[14540]_  = ~\new_[14541]_  & ~\new_[14543]_ ;
  assign \new_[14541]_  = \new_[14542]_  & \new_[14532]_ ;
  assign \new_[14542]_  = ~\new_[4834]_ ;
  assign \new_[14543]_  = \new_[4615]_  | \new_[14544]_ ;
  assign \new_[14544]_  = ~\new_[14532]_  & ~\new_[4811]_ ;
  assign \new_[14545]_  = \new_[14546]_  | \new_[14547]_ ;
  assign \new_[14546]_  = ~\new_[4615]_  | ~\new_[4852]_ ;
  assign \new_[14547]_  = ~\new_[14544]_  & ~\new_[14541]_ ;
  assign \new_[14548]_  = ~\new_[14544]_  & ~\new_[14541]_ ;
  assign \new_[14549]_  = ~\new_[14553]_  | ~\new_[14550]_  | ~\new_[14552]_ ;
  assign \new_[14550]_  = ~\new_[14750]_  & ~\new_[14551]_ ;
  assign \new_[14551]_  = ~\new_[14749]_  | ~\new_[14728]_ ;
  assign \new_[14552]_  = \new_[14726]_  & \new_[2690]_ ;
  assign \new_[14553]_  = \new_[14748]_  & \new_[14556]_ ;
  assign \new_[14554]_  = ~\new_[2681]_  | ~\new_[2703]_ ;
  assign \new_[14555]_  = ~\new_[2702]_  | ~\new_[2680]_ ;
  assign \new_[14556]_  = ~\new_[14557]_  | ~\new_[11016]_ ;
  assign \new_[14557]_  = ~\new_[14638]_ ;
  assign \new_[14558]_  = \new_[14775]_  & \new_[14774]_ ;
  assign \new_[14559]_  = \new_[2801]_ ;
  assign \new_[14560]_  = ~\new_[14561]_  & (~\new_[5900]_  | ~\new_[7450]_ );
  assign \new_[14561]_  = ~\new_[14296]_  | ~\new_[14297]_  | ~\new_[14562]_ ;
  assign \new_[14562]_  = ~\new_[7746]_  | ~\new_[14418]_ ;
  assign \new_[14563]_  = ~\new_[14418]_  | ~\new_[14294]_  | ~\new_[14293]_ ;
  assign \new_[14564]_  = ~\new_[14568]_  | ~\new_[14565]_ ;
  assign \new_[14565]_  = ~\new_[14566]_  | ~\new_[10638]_ ;
  assign \new_[14566]_  = ~\new_[14567]_ ;
  assign \new_[14567]_  = ~\new_[3120]_  | ~\new_[3044]_ ;
  assign \new_[14568]_  = ~\new_[11382]_  | ~\new_[14721]_ ;
  assign \new_[14569]_  = \new_[14570]_  ? \new_[14592]_  : \new_[14571]_ ;
  assign \new_[14570]_  = ~\new_[14571]_ ;
  assign \new_[14571]_  = \new_[2038]_  ^ \new_[4607]_ ;
  assign \new_[14572]_  = ~\new_[14593]_  | ~\new_[14756]_ ;
  assign \new_[14573]_  = ~\new_[2577]_  & ~\new_[2576]_ ;
  assign \new_[14574]_  = ~\new_[14575]_  & ~\new_[14576]_ ;
  assign \new_[14575]_  = ~\new_[2699]_  | ~\new_[2679]_ ;
  assign \new_[14576]_  = ~\new_[2697]_  | ~\new_[2698]_ ;
  assign \new_[14577]_  = \new_[14578]_  & \new_[14582]_ ;
  assign \new_[14578]_  = ~\new_[13756]_  | ~\new_[14579]_ ;
  assign \new_[14579]_  = ~\new_[14580]_  | ~\new_[14581]_ ;
  assign \new_[14580]_  = ~\new_[14369]_ ;
  assign \new_[14581]_  = ~\new_[14332]_  | ~\new_[4817]_ ;
  assign \new_[14582]_  = ~\new_[12610]_  | ~\new_[13756]_ ;
  assign \new_[14583]_  = ~\new_[14585]_  | (~\new_[14584]_  & ~\new_[14369]_ );
  assign \new_[14584]_  = ~\new_[14581]_  | ~\new_[4801]_ ;
  assign \new_[14585]_  = ~\new_[14426]_  | ~\new_[14425]_ ;
  assign \new_[14586]_  = ~\new_[14585]_  | ~\new_[14579]_ ;
  assign \new_[14587]_  = ~\new_[14579]_ ;
  assign \new_[14588]_  = ~\new_[14713]_  | ~\new_[14504]_ ;
  assign \new_[14589]_  = ~\new_[14591]_  | ~\new_[14590]_  | ~\new_[14718]_ ;
  assign \new_[14590]_  = ~\new_[14704]_  | ~\new_[14648]_ ;
  assign \new_[14591]_  = ~\new_[14564]_  & ~\new_[14594]_ ;
  assign \new_[14592]_  = ~\new_[14593]_  | ~\new_[14756]_ ;
  assign \new_[14593]_  = ~\new_[14462]_  | ~\new_[14795]_ ;
  assign \new_[14594]_  = ~\new_[14595]_  | ~\new_[14598]_ ;
  assign \new_[14595]_  = ~\new_[14596]_  | ~\new_[10635]_ ;
  assign \new_[14596]_  = ~\new_[14597]_ ;
  assign \new_[14597]_  = ~\new_[3044]_  | ~\new_[14822]_ ;
  assign \new_[14598]_  = ~\new_[2840]_  | ~\new_[11215]_ ;
  assign \new_[14599]_  = ~\new_[14600]_ ;
  assign \new_[14600]_  = \new_[13241]_  ^ \new_[12903]_ ;
  assign \new_[14601]_  = \new_[14602]_  ? \new_[14606]_  : \new_[14605]_ ;
  assign \new_[14602]_  = ~\new_[14604]_  & (~\new_[14603]_  | ~\new_[13546]_ );
  assign \new_[14603]_  = ~\new_[4607]_ ;
  assign \new_[14604]_  = ~\new_[14603]_  & ~\new_[13546]_ ;
  assign \new_[14605]_  = ~\new_[14602]_ ;
  assign \new_[14606]_  = ~\new_[2277]_  | ~\new_[2300]_ ;
  assign \new_[14607]_  = \new_[14606]_ ;
  assign \new_[14608]_  = ~\new_[14612]_  | (~\new_[14609]_  & ~\new_[14829]_ );
  assign \new_[14609]_  = ~\new_[14611]_  & (~\new_[14610]_  | ~\new_[2630]_ );
  assign \new_[14610]_  = \new_[14827]_ ;
  assign \new_[14611]_  = \new_[10490]_  & \new_[2870]_ ;
  assign \new_[14612]_  = ~\new_[14829]_  | ~\new_[4615]_ ;
  assign \new_[14613]_  = ~\new_[14619]_  & (~\new_[14614]_  | ~\new_[14618]_ );
  assign \new_[14614]_  = ~\new_[14615]_  | ~\new_[14617]_ ;
  assign \new_[14615]_  = ~\new_[6226]_  | (~\new_[14616]_  & ~\new_[5425]_ );
  assign \new_[14616]_  = \new_[6118]_  & \new_[6763]_ ;
  assign \new_[14617]_  = ~\new_[7446]_  & (~\new_[7744]_  | ~\new_[6774]_ );
  assign \new_[14618]_  = ~\new_[6224]_  & ~\new_[6706]_ ;
  assign \new_[14619]_  = ~\new_[6180]_  | (~\new_[5957]_  & ~\new_[6706]_ );
  assign \new_[14620]_  = ~\new_[14626]_  & (~\new_[14621]_  | ~\new_[14624]_ );
  assign \new_[14621]_  = ~\new_[14623]_  & (~\new_[2366]_  | ~\new_[14622]_ );
  assign \new_[14622]_  = ~\new_[2416]_  | ~\new_[4862]_ ;
  assign \new_[14623]_  = ~\new_[14336]_  & ~\new_[14333]_ ;
  assign \new_[14624]_  = ~\new_[14622]_  | ~\new_[14625]_  | ~\new_[2365]_ ;
  assign \new_[14625]_  = \new_[2364]_  | \new_[2363]_ ;
  assign \new_[14626]_  = ~\new_[14627]_ ;
  assign \new_[14627]_  = ~\new_[14338]_  | ~\new_[4883]_ ;
  assign \new_[14628]_  = ~\new_[14627]_  | (~\new_[14623]_  & ~\new_[14622]_ );
  assign \new_[14629]_  = ~\new_[14625]_  | ~\new_[2365]_ ;
  assign \new_[14630]_  = ~\new_[2366]_  & ~\new_[14623]_ ;
  assign \new_[14631]_  = ~\new_[14742]_  & ~\new_[14732]_ ;
  assign \new_[14632]_  = ~\new_[2258]_  | (~\new_[14367]_  & ~\new_[2272]_ );
  assign \new_[14633]_  = ~\new_[2258]_  | (~\new_[14367]_  & ~\new_[2272]_ );
  assign \new_[14634]_  = ~\new_[14390]_  | ~\new_[14382]_  | ~\new_[14389]_ ;
  assign \new_[14635]_  = ~\new_[14390]_  | ~\new_[14382]_  | ~\new_[14389]_ ;
  assign \new_[14636]_  = ~\new_[12422]_  & (~\new_[10720]_  | ~\new_[10572]_ );
  assign \new_[14637]_  = ~\new_[12422]_  & (~\new_[10720]_  | ~\new_[10572]_ );
  assign \new_[14638]_  = ~\new_[14773]_  | ~\new_[14658]_ ;
  assign \new_[14639]_  = ~\new_[14773]_  | ~\new_[14658]_ ;
  assign \new_[14640]_  = ~\new_[14641]_  | ~\new_[14643]_ ;
  assign \new_[14641]_  = \new_[14642]_  & \new_[14733]_ ;
  assign \new_[14642]_  = ~\new_[12433]_  | ~\new_[14391]_  | ~\new_[14385]_ ;
  assign \new_[14643]_  = ~\new_[14388]_  | ~\new_[14383]_  | ~\new_[14384]_ ;
  assign \new_[14644]_  = ~\new_[14645]_  | ~\new_[14646]_ ;
  assign \new_[14645]_  = ~\new_[2845]_  | ~\new_[11387]_ ;
  assign \new_[14646]_  = ~\new_[11349]_  | ~\new_[2844]_ ;
  assign \new_[14647]_  = ~\new_[2700]_  | ~\new_[2701]_ ;
  assign \new_[14648]_  = ~\new_[14649]_  & ~\new_[14719]_ ;
  assign \new_[14649]_  = ~\new_[14371]_  | ~\new_[14655]_ ;
  assign \new_[14650]_  = ~\new_[2192]_  | ~\new_[12654]_  | ~\new_[2176]_ ;
  assign \new_[14651]_  = ~\new_[14652]_  & ~\new_[14653]_ ;
  assign \new_[14652]_  = ~\new_[4512]_  & ~\new_[2483]_ ;
  assign \new_[14653]_  = ~\new_[4857]_  & ~\new_[14654]_ ;
  assign \new_[14654]_  = ~\new_[9834]_  & ~\new_[2595]_ ;
  assign \new_[14655]_  = ~\new_[14753]_  | ~\new_[11390]_ ;
  assign \new_[14656]_  = ~\new_[14631]_  & ~\new_[14506]_ ;
  assign \new_[14657]_  = ~\new_[14658]_ ;
  assign \new_[14658]_  = \new_[14823]_ ;
  assign \new_[14659]_  = ~\new_[14660]_  | ~\new_[14661]_ ;
  assign \new_[14660]_  = \new_[13442]_  | \new_[13252]_ ;
  assign \new_[14661]_  = ~\new_[14662]_  | ~\new_[9188]_ ;
  assign \new_[14662]_  = ~\new_[14663]_ ;
  assign \new_[14663]_  = ~\new_[14485]_  | ~\new_[14486]_ ;
  assign \new_[14664]_  = \new_[4788]_  & \new_[14663]_ ;
  assign \new_[14665]_  = ~\new_[14660]_ ;
  assign \new_[14666]_  = ~\new_[14662]_ ;
  assign \new_[14667]_  = ~\new_[4515]_  & ~\new_[14668]_ ;
  assign \new_[14668]_  = ~\new_[14669]_  | ~\new_[14672]_ ;
  assign \new_[14669]_  = ~\new_[14671]_  | (~\new_[9312]_  & ~\new_[14670]_ );
  assign \new_[14670]_  = \new_[2719]_  & \new_[9036]_ ;
  assign \new_[14671]_  = ~\new_[14829]_ ;
  assign \new_[14672]_  = ~\new_[14832]_  | ~\new_[4799]_ ;
  assign \new_[14673]_  = ~\new_[14674]_ ;
  assign \new_[14674]_  = ~\new_[14558]_  | ~\new_[14657]_ ;
  assign \new_[14675]_  = ~\new_[14558]_  | ~\new_[14657]_ ;
  assign \new_[14676]_  = \new_[14677]_  & \new_[14678]_ ;
  assign \new_[14677]_  = ~\new_[14483]_  | ~\new_[14650]_ ;
  assign \new_[14678]_  = ~\new_[14559]_  | ~\new_[14701]_ ;
  assign \new_[14679]_  = ~\new_[14373]_  | ~\new_[14700]_ ;
  assign \new_[14680]_  = ~\new_[14677]_  & ~\new_[12734]_ ;
  assign \new_[14681]_  = ~\new_[14573]_  | ~\new_[14574]_ ;
  assign \new_[14682]_  = ~\new_[14683]_  | ~\new_[14684]_ ;
  assign \new_[14683]_  = ~\new_[14647]_  & ~\new_[14555]_ ;
  assign \new_[14684]_  = ~\new_[14554]_  & ~\new_[14644]_ ;
  assign \new_[14685]_  = ~\new_[14686]_  | ~\new_[14693]_ ;
  assign \new_[14686]_  = ~\new_[14687]_  | ~\new_[14692]_ ;
  assign \new_[14687]_  = ~\new_[14688]_ ;
  assign \new_[14688]_  = ~\new_[14689]_  | ~\new_[14690]_ ;
  assign \new_[14689]_  = ~\new_[14298]_  | ~\new_[14299]_ ;
  assign \new_[14690]_  = ~\new_[14691]_ ;
  assign \new_[14691]_  = ~\new_[14513]_  & ~\new_[14392]_ ;
  assign \new_[14692]_  = ~\new_[2355]_  | ~\new_[2408]_ ;
  assign \new_[14693]_  = ~\new_[14694]_ ;
  assign \new_[14694]_  = ~\new_[14695]_  | ~\new_[14697]_ ;
  assign \new_[14695]_  = ~\new_[14696]_  | ~\new_[14690]_ ;
  assign \new_[14696]_  = ~\new_[14378]_ ;
  assign \new_[14697]_  = ~\new_[14393]_  | ~\new_[4514]_ ;
  assign \new_[14698]_  = ~\new_[14690]_ ;
  assign \new_[14699]_  = ~\new_[14511]_  | ~\new_[14701]_ ;
  assign \new_[14700]_  = ~\new_[14701]_ ;
  assign \new_[14701]_  = ~\new_[2636]_ ;
  assign \new_[14702]_  = ~\new_[14703]_  | ~\new_[14700]_ ;
  assign \new_[14703]_  = ~\new_[14483]_  | ~\new_[14650]_ ;
  assign \new_[14704]_  = ~\new_[14705]_  & ~\new_[14707]_ ;
  assign \new_[14705]_  = ~\new_[14706]_  | ~\new_[2689]_ ;
  assign \new_[14706]_  = ~\new_[2843]_  | ~\new_[10651]_ ;
  assign \new_[14707]_  = ~\new_[14817]_  | ~\new_[14708]_ ;
  assign \new_[14708]_  = ~\new_[14596]_  | ~\new_[10359]_ ;
  assign \new_[14709]_  = ~\new_[14744]_  & ~\new_[14710]_ ;
  assign \new_[14710]_  = ~\new_[14317]_  & ~\new_[14316]_ ;
  assign \new_[14711]_  = \new_[14724]_  & \new_[14746]_ ;
  assign \new_[14712]_  = ~\new_[14454]_  | ~\new_[14439]_ ;
  assign \new_[14713]_  = ~\new_[14714]_  | ~\new_[14717]_ ;
  assign \new_[14714]_  = ~\new_[14716]_  & ~\new_[14715]_ ;
  assign \new_[14715]_  = ~\new_[2688]_  | ~\new_[2676]_ ;
  assign \new_[14716]_  = ~\new_[2687]_  | ~\new_[2686]_ ;
  assign \new_[14717]_  = ~\new_[14564]_  & ~\new_[14594]_ ;
  assign \new_[14718]_  = ~\new_[14715]_  & ~\new_[14716]_ ;
  assign \new_[14719]_  = ~\new_[14720]_  | ~\new_[14723]_ ;
  assign \new_[14720]_  = ~\new_[14721]_  | ~\new_[11383]_ ;
  assign \new_[14721]_  = ~\new_[14722]_ ;
  assign \new_[14722]_  = ~\new_[14505]_  | ~\new_[14658]_ ;
  assign \new_[14723]_  = ~\new_[14557]_  | ~\new_[11364]_ ;
  assign \new_[14724]_  = ~\new_[14725]_  & ~\new_[14727]_ ;
  assign \new_[14725]_  = ~\new_[14556]_  | ~\new_[14726]_ ;
  assign \new_[14726]_  = ~\new_[14824]_  | ~\new_[10639]_ ;
  assign \new_[14727]_  = ~\new_[2690]_  | ~\new_[14728]_ ;
  assign \new_[14728]_  = ~\new_[14596]_  | ~\new_[10637]_ ;
  assign \new_[14729]_  = ~\new_[14680]_  & (~\new_[14676]_  | ~\new_[14679]_ );
  assign \new_[14730]_  = ~\new_[14742]_  & ~\new_[14731]_ ;
  assign \new_[14731]_  = ~\new_[14777]_  & ~\new_[14709]_ ;
  assign \new_[14732]_  = ~\new_[14709]_  & ~\new_[14777]_ ;
  assign \new_[14733]_  = ~\new_[14741]_  | ~\new_[14734]_  | ~\new_[14739]_ ;
  assign \new_[14734]_  = ~\new_[14735]_ ;
  assign \new_[14735]_  = ~\new_[14736]_  | ~\new_[14738]_ ;
  assign \new_[14736]_  = ~\new_[14737]_ ;
  assign \new_[14737]_  = ~\new_[11585]_  | ~\new_[12283]_ ;
  assign \new_[14738]_  = \new_[13950]_  & \new_[13877]_ ;
  assign \new_[14739]_  = ~\new_[14740]_ ;
  assign \new_[14740]_  = ~\new_[12953]_  | ~\new_[12570]_ ;
  assign \new_[14741]_  = ~\new_[6083]_  & ~\new_[14342]_ ;
  assign \new_[14742]_  = ~\new_[14743]_  & ~\new_[14745]_ ;
  assign \new_[14743]_  = \new_[2734]_  | \new_[14744]_ ;
  assign \new_[14744]_  = \new_[4882]_ ;
  assign \new_[14745]_  = ~\new_[14316]_  & ~\new_[14317]_ ;
  assign \new_[14746]_  = ~\new_[14750]_  & ~\new_[14747]_ ;
  assign \new_[14747]_  = ~\new_[14748]_  | ~\new_[14749]_ ;
  assign \new_[14748]_  = ~\new_[2842]_  | ~\new_[10632]_ ;
  assign \new_[14749]_  = ~\new_[2847]_  | ~\new_[10674]_ ;
  assign \new_[14750]_  = ~\new_[14751]_  | ~\new_[14752]_ ;
  assign \new_[14751]_  = ~\new_[14673]_  | ~\new_[11217]_ ;
  assign \new_[14752]_  = ~\new_[14753]_  | ~\new_[11354]_ ;
  assign \new_[14753]_  = ~\new_[14754]_ ;
  assign \new_[14754]_  = ~\new_[14657]_  | ~\new_[14656]_ ;
  assign \new_[14755]_  = ~\new_[14657]_  | ~\new_[14656]_ ;
  assign \new_[14756]_  = ~\new_[14757]_  | ~\new_[14761]_ ;
  assign \new_[14757]_  = ~\new_[14758]_ ;
  assign \new_[14758]_  = ~\new_[14759]_  | ~\new_[14760]_ ;
  assign \new_[14759]_  = ~\new_[14439]_  | ~\new_[14549]_  | ~\new_[14454]_ ;
  assign \new_[14760]_  = ~\new_[14711]_  | ~\new_[14712]_ ;
  assign \new_[14761]_  = ~\new_[14588]_  | ~\new_[14589]_ ;
  assign \new_[14762]_  = ~\new_[14529]_  | ~\new_[4923]_ ;
  assign \new_[14763]_  = \new_[14764]_  ^ \new_[14767]_ ;
  assign \new_[14764]_  = \new_[14765]_  ? \new_[14793]_  : \new_[14766]_ ;
  assign \new_[14765]_  = ~\new_[14766]_ ;
  assign \new_[14766]_  = ~\new_[14395]_  | ~\new_[2336]_ ;
  assign \new_[14767]_  = \new_[14599]_  ? \new_[14601]_  : \new_[14600]_ ;
  assign \new_[14768]_  = ~\new_[14560]_  | ~\new_[14563]_ ;
  assign \new_[14769]_  = \new_[14762]_  & \new_[14477]_ ;
  assign \new_[14770]_  = \new_[14771]_  | \new_[14772]_ ;
  assign \new_[14771]_  = ~\new_[14583]_ ;
  assign \new_[14772]_  = ~\new_[14577]_ ;
  assign \new_[14773]_  = \new_[14775]_  & \new_[14774]_ ;
  assign \new_[14774]_  = ~\new_[14510]_  | ~\new_[14509]_ ;
  assign \new_[14775]_  = \new_[14776]_  ? \new_[14778]_  : \new_[14459]_ ;
  assign \new_[14776]_  = ~\new_[14777]_ ;
  assign \new_[14777]_  = \new_[14459]_  ? \new_[14460]_  : \new_[2734]_ ;
  assign \new_[14778]_  = ~\new_[4882]_  & ~\new_[14745]_ ;
  assign n1250 = (~\new_[14780]_  | ~\new_[14792]_ ) & (~\new_[14789]_  | ~\new_[14790]_ );
  assign \new_[14780]_  = ~\new_[14781]_ ;
  assign \new_[14781]_  = ~\new_[14782]_ ;
  assign \new_[14782]_  = ~\new_[14783]_ ;
  assign \new_[14783]_  = ~\new_[14786]_  | ~\new_[14784]_  | ~\new_[14785]_ ;
  assign \new_[14784]_  = ~\new_[14769]_  | ~\new_[14768]_  | ~\new_[14770]_ ;
  assign \new_[14785]_  = ~\new_[14474]_  | ~\new_[14762]_ ;
  assign \new_[14786]_  = ~\new_[6651]_  & ~\new_[14310]_ ;
  assign \new_[14787]_  = \new_[14788]_ ;
  assign \new_[14788]_  = \new_[4812]_  ? \new_[14331]_  : \new_[4835]_ ;
  assign \new_[14789]_  = ~\new_[14782]_ ;
  assign \new_[14790]_  = ~\new_[4796]_ ;
  assign \new_[14791]_  = ~\new_[14786]_  | ~\new_[14784]_  | ~\new_[14785]_ ;
  assign \new_[14792]_  = ~\new_[14787]_ ;
  assign \new_[14793]_  = \new_[14794]_  ? \new_[14796]_  : \new_[2320]_ ;
  assign \new_[14794]_  = ~\new_[14795]_ ;
  assign \new_[14795]_  = ~\new_[14759]_  | ~\new_[14760]_ ;
  assign \new_[14796]_  = ~\new_[14797]_  | ~\new_[14798]_ ;
  assign \new_[14797]_  = \new_[14681]_  | \new_[14682]_ ;
  assign \new_[14798]_  = ~\new_[14682]_  | ~\new_[14681]_ ;
  assign \new_[14799]_  = ~\new_[14800]_ ;
  assign \new_[14800]_  = ~\new_[14801]_ ;
  assign \new_[14801]_  = ~\new_[14807]_  | ~\new_[14802]_  | ~\new_[14803]_ ;
  assign \new_[14802]_  = ~\new_[2615]_  & (~\new_[2338]_  | ~\new_[2315]_ );
  assign \new_[14803]_  = ~\new_[14804]_ ;
  assign \new_[14804]_  = ~\new_[14806]_  | ~\new_[14805]_  | ~\new_[2451]_ ;
  assign \new_[14805]_  = ~\new_[2313]_ ;
  assign \new_[14806]_  = ~\new_[11573]_ ;
  assign \new_[14807]_  = ~\new_[14808]_  & ~\new_[14812]_ ;
  assign \new_[14808]_  = ~\new_[14809]_  | ~\new_[14810]_ ;
  assign \new_[14809]_  = \new_[2391]_  & \new_[2449]_ ;
  assign \new_[14810]_  = \new_[14811]_  ? \new_[8593]_  : \new_[2499]_ ;
  assign \new_[14811]_  = ~\new_[2499]_ ;
  assign \new_[14812]_  = ~\new_[14813]_  | ~\new_[14816]_ ;
  assign \new_[14813]_  = ~\new_[14814]_  & ~\new_[14815]_ ;
  assign \new_[14814]_  = ~\new_[2671]_ ;
  assign \new_[14815]_  = ~\new_[2526]_  | ~\new_[2616]_ ;
  assign \new_[14816]_  = \new_[2525]_  & \new_[2617]_ ;
  assign \new_[14817]_  = ~\new_[14818]_  | ~\new_[10652]_ ;
  assign \new_[14818]_  = ~\new_[14819]_ ;
  assign \new_[14819]_  = ~\new_[14820]_  | ~\new_[14822]_ ;
  assign \new_[14820]_  = ~\new_[14821]_ ;
  assign \new_[14821]_  = ~\new_[14730]_  | ~\new_[14729]_ ;
  assign \new_[14822]_  = \new_[14823]_ ;
  assign \new_[14823]_  = ~\new_[14699]_  | ~\new_[14702]_ ;
  assign \new_[14824]_  = ~\new_[14819]_ ;
  assign \new_[14825]_  = ~\new_[14831]_  | (~\new_[14826]_  & ~\new_[14829]_ );
  assign \new_[14826]_  = ~\new_[14828]_  & (~\new_[14834]_  | ~\new_[2632]_ );
  assign \new_[14827]_  = ~\new_[14339]_  | ~\new_[12464]_ ;
  assign \new_[14828]_  = \new_[10490]_  & \new_[2871]_ ;
  assign \new_[14829]_  = ~\new_[14830]_ ;
  assign \new_[14830]_  = ~\new_[14659]_  | ~\new_[14664]_ ;
  assign \new_[14831]_  = ~\new_[14829]_  | ~\new_[4796]_ ;
  assign \new_[14832]_  = ~\new_[14833]_ ;
  assign \new_[14833]_  = ~\new_[14829]_ ;
  assign \new_[14834]_  = ~\new_[10490]_ ;
  assign n970 = n980;
  assign n1885 = n1890;
  assign n4025 = n4030;
  assign n7545 = n7550;
  assign n8895 = n8945;
  assign n8900 = n9005;
  assign n8950 = n8955;
  assign n8960 = TxReady_pad_i;
  assign n8970 = n8985;
  assign n8975 = n8990;
  assign n8980 = n8995;
  assign n9095 = \VStatus_pad_i[5] ;
  assign n9100 = \VStatus_pad_i[1] ;
  assign n9105 = \VStatus_pad_i[3] ;
  assign n9110 = \DataIn_pad_i[2] ;
  assign n9115 = \VStatus_pad_i[2] ;
  assign n9125 = \DataIn_pad_i[7] ;
  assign n9135 = \DataIn_pad_i[3] ;
  assign n9155 = \LineState_pad_i[0] ;
  assign n9160 = \VStatus_pad_i[4] ;
  assign n9165 = \DataIn_pad_i[0] ;
  assign n9175 = \DataIn_pad_i[5] ;
  assign n9180 = \VStatus_pad_i[7] ;
  assign n9185 = \LineState_pad_i[1] ;
  assign n9190 = \DataIn_pad_i[6] ;
  assign n9195 = \LineState_pad_i[0] ;
  assign n9200 = \DataIn_pad_i[4] ;
  assign n9205 = \DataIn_pad_i[1] ;
  assign n9210 = \LineState_pad_i[1] ;
  assign n9220 = \VStatus_pad_i[6] ;
  assign n9225 = \VStatus_pad_i[0] ;
  always @ (posedge clock) begin
    \\u0_DataOut_reg[3]  <= n500;
    \\u0_DataOut_reg[7]  <= n505;
    \\u0_DataOut_reg[2]  <= n510;
    \\u0_DataOut_reg[6]  <= n515;
    \\u1_u3_token_pid_sel_reg[0]  <= n520;
    \\u1_u3_token_pid_sel_reg[1]  <= n525;
    u1_u3_no_bufs0_reg <= n530;
    \\u1_u3_idin_reg[13]  <= n535;
    u1_u3_no_bufs1_reg <= n540;
    \\u1_u1_crc16_reg[15]  <= n545;
    \\u1_u1_crc16_reg[1]  <= n550;
    \\u1_u3_idin_reg[14]  <= n555;
    u1_u3_buffer_done_reg <= n560;
    \\u1_u1_crc16_reg[0]  <= n565;
    \\u1_u3_idin_reg[12]  <= n570;
    \\u1_u3_idin_reg[16]  <= n575;
    \\u1_u3_idin_reg[10]  <= n580;
    \\u0_DataOut_reg[4]  <= n585;
    \\u1_u3_idin_reg[15]  <= n590;
    \\u1_u3_idin_reg[11]  <= n595;
    \\u0_DataOut_reg[1]  <= n600;
    \\u0_DataOut_reg[0]  <= n605;
    \\u1_u3_idin_reg[9]  <= n610;
    \\u1_u3_idin_reg[6]  <= n615;
    u1_u3_buffer_full_reg <= n620;
    \\u1_u1_crc16_reg[8]  <= n625;
    \\u0_DataOut_reg[5]  <= n630;
    \\u1_u3_idin_reg[8]  <= n635;
    \\u1_u3_idin_reg[5]  <= n640;
    u1_u3_buffer_empty_reg <= n645;
    \\u1_u3_idin_reg[7]  <= n650;
    \\u1_u2_adr_cw_reg[11]  <= n655;
    \\u1_u2_adr_cw_reg[13]  <= n660;
    \\u1_u2_adr_cw_reg[14]  <= n665;
    \\u1_u2_adr_cw_reg[5]  <= n670;
    \\u1_u2_adr_cw_reg[6]  <= n675;
    \\u1_u2_adr_cw_reg[7]  <= n680;
    \\u1_u2_adr_cw_reg[8]  <= n685;
    \\u1_u2_adr_cw_reg[0]  <= n690;
    \\u1_u2_adr_cw_reg[3]  <= n695;
    \\u1_u2_adr_cw_reg[2]  <= n700;
    \\u1_u2_adr_cw_reg[4]  <= n705;
    \\u1_u2_adr_cw_reg[10]  <= n710;
    \\u1_u2_adr_cw_reg[12]  <= n715;
    \\u1_u2_adr_cw_reg[1]  <= n720;
    \\u1_u2_adr_cw_reg[9]  <= n725;
    \\u1_u3_idin_reg[4]  <= n730;
    u0_TxValid_reg <= n735;
    \\u1_u1_crc16_reg[6]  <= n740;
    \\u1_u3_idin_reg[3]  <= n745;
    \\u1_u1_crc16_reg[2]  <= n750;
    \\u1_u1_crc16_reg[3]  <= n755;
    \\u1_u1_crc16_reg[4]  <= n760;
    \\u1_u1_crc16_reg[7]  <= n765;
    \\u1_u1_crc16_reg[9]  <= n770;
    \\u1_u1_state_reg[1]  <= n775;
    \\u1_u3_idin_reg[2]  <= n780;
    \\u1_u3_idin_reg[1]  <= n785;
    u1_u1_tx_valid_r_reg <= n790;
    \\u1_u1_state_reg[0]  <= n795;
    \\u1_u1_crc16_reg[5]  <= n800;
    \\u1_u1_state_reg[4]  <= n805;
    u1_u1_tx_valid_r1_reg <= n810;
    \\u1_u3_idin_reg[30]  <= n815;
    \\u1_u3_idin_reg[0]  <= n820;
    u1_u1_send_token_r_reg <= n825;
    u1_u1_zero_length_r_reg <= n830;
    \\u1_u3_state_reg[0]  <= n835;
    u1_u1_tx_first_r_reg <= n840;
    \\u1_u2_sizd_c_reg[10]  <= n845;
    \\u1_u2_sizd_c_reg[12]  <= n850;
    \\u1_u2_sizd_c_reg[4]  <= n855;
    u4_u1_dma_req_r_reg <= n860;
    \\u1_u2_sizd_c_reg[0]  <= n865;
    \\u1_u2_sizd_c_reg[11]  <= n870;
    \\u1_u2_sizd_c_reg[13]  <= n875;
    \\u1_u2_sizd_c_reg[1]  <= n880;
    \\u1_u2_sizd_c_reg[2]  <= n885;
    \\u1_u2_sizd_c_reg[3]  <= n890;
    \\u1_u2_sizd_c_reg[5]  <= n895;
    \\u1_u2_sizd_c_reg[6]  <= n900;
    \\u1_u2_sizd_c_reg[7]  <= n905;
    \\u1_u2_sizd_c_reg[8]  <= n910;
    \\u1_u2_sizd_c_reg[9]  <= n915;
    u4_u2_dma_req_r_reg <= n920;
    u4_u0_dma_req_r_reg <= n925;
    \\u1_u3_new_size_reg[13]  <= n930;
    u4_u3_dma_req_r_reg <= n935;
    \\u1_u3_state_reg[1]  <= n940;
    \\u1_u3_state_reg[4]  <= n945;
    \\u1_u2_last_buf_adr_reg[13]  <= n950;
    \\u1_u2_last_buf_adr_reg[14]  <= n955;
    \\u1_u3_state_reg[2]  <= n960;
    u1_u3_send_token_reg <= n965;
    u1_u1_send_zero_length_r_reg <= n970;
    \\u1_u3_state_reg[8]  <= n975;
    u1_u2_send_zero_length_r_reg <= n980;
    u1_u2_rx_dma_en_r_reg <= n985;
    \\u1_u3_new_sizeb_reg[6]  <= n990;
    \\u1_u3_new_sizeb_reg[7]  <= n995;
    \\u1_u3_new_sizeb_reg[8]  <= n1000;
    \\u1_u3_new_sizeb_reg[9]  <= n1005;
    \\u1_u2_last_buf_adr_reg[10]  <= n1010;
    \\u1_u3_new_sizeb_reg[0]  <= n1015;
    \\u1_u3_new_sizeb_reg[1]  <= n1020;
    \\u1_u3_new_sizeb_reg[2]  <= n1025;
    \\u1_u3_new_sizeb_reg[3]  <= n1030;
    \\u1_u3_new_sizeb_reg[5]  <= n1035;
    \\u1_u3_state_reg[3]  <= n1040;
    \\u1_u3_state_reg[5]  <= n1045;
    \\u1_u3_state_reg[6]  <= n1050;
    \\u1_u3_state_reg[7]  <= n1055;
    \\u1_u3_state_reg[9]  <= n1060;
    \\u1_u2_last_buf_adr_reg[12]  <= n1065;
    \\u4_u2_int_stat_reg[2]  <= n1070;
    \\u4_u3_int_stat_reg[2]  <= n1075;
    \\u4_u0_int_stat_reg[2]  <= n1080;
    \\u1_u3_new_sizeb_reg[4]  <= n1085;
    \\u4_u1_int_stat_reg[2]  <= n1090;
    \\u1_u3_new_sizeb_reg[10]  <= n1095;
    \\u1_u2_last_buf_adr_reg[9]  <= n1100;
    u1_u2_tx_dma_en_r_reg <= n1105;
    \\u1_u2_last_buf_adr_reg[11]  <= n1110;
    \\u1_u3_new_sizeb_reg[13]  <= n1115;
    \\u1_u3_idin_reg[27]  <= n1120;
    u4_dma_out_buf_avail_reg <= n1125;
    \\u1_u3_new_sizeb_reg[11]  <= n1130;
    \\u1_u3_new_sizeb_reg[12]  <= n1135;
    \\u4_u2_int_stat_reg[5]  <= n1140;
    \\u4_u3_int_stat_reg[5]  <= n1145;
    \\u4_u0_int_stat_reg[5]  <= n1150;
    \\u4_u1_int_stat_reg[5]  <= n1155;
    \\u1_u3_size_next_r_reg[7]  <= n1160;
    \\u1_u3_size_next_r_reg[6]  <= n1165;
    \\u1_u3_size_next_r_reg[8]  <= n1170;
    \\u1_u3_size_next_r_reg[9]  <= n1175;
    \\u4_int_srcb_reg[2]  <= n1180;
    u4_u1_dma_req_in_hold2_reg <= n1185;
    u1_u3_abort_reg <= n1190;
    \\u1_u2_last_buf_adr_reg[8]  <= n1195;
    \\u1_u2_last_buf_adr_reg[6]  <= n1200;
    \\u1_u2_dout_r_reg[30]  <= n1205;
    u4_u2_dma_req_in_hold2_reg <= n1210;
    u4_u0_dma_req_in_hold2_reg <= n1215;
    \\u1_u2_dout_r_reg[5]  <= n1220;
    \\u1_u2_dout_r_reg[27]  <= n1225;
    \\u1_u2_dout_r_reg[1]  <= n1230;
    \\u1_u2_dout_r_reg[16]  <= n1235;
    \\u1_u3_size_next_r_reg[1]  <= n1240;
    \\u1_u3_size_next_r_reg[3]  <= n1245;
    \\u1_u3_size_next_r_reg[2]  <= n1250;
    \\u1_u3_size_next_r_reg[5]  <= n1255;
    \\u1_u2_adr_cb_reg[0]  <= n1260;
    \\u1_mfm_cnt_reg[1]  <= n1265;
    \\u1_u3_idin_reg[25]  <= n1270;
    \\u1_u3_idin_reg[26]  <= n1275;
    \\u1_u2_dout_r_reg[0]  <= n1280;
    \\u1_u2_dout_r_reg[10]  <= n1285;
    \\u1_u2_dout_r_reg[12]  <= n1290;
    \\u1_u2_dout_r_reg[11]  <= n1295;
    \\u1_u2_dout_r_reg[13]  <= n1300;
    \\u1_u2_dout_r_reg[14]  <= n1305;
    \\u1_u2_dout_r_reg[15]  <= n1310;
    \\u1_u2_dout_r_reg[17]  <= n1315;
    \\u1_u2_dout_r_reg[18]  <= n1320;
    \\u1_u2_dout_r_reg[19]  <= n1325;
    \\u1_u2_dout_r_reg[20]  <= n1330;
    \\u1_u2_dout_r_reg[21]  <= n1335;
    \\u1_u2_dout_r_reg[22]  <= n1340;
    \\u1_u2_dout_r_reg[23]  <= n1345;
    \\u1_u2_dout_r_reg[24]  <= n1350;
    \\u1_u2_dout_r_reg[25]  <= n1355;
    \\u1_u2_dout_r_reg[26]  <= n1360;
    \\u1_u2_dout_r_reg[28]  <= n1365;
    \\u1_u2_dout_r_reg[29]  <= n1370;
    \\u1_u2_dout_r_reg[2]  <= n1375;
    \\u1_u2_dout_r_reg[31]  <= n1380;
    \\u1_u2_dout_r_reg[3]  <= n1385;
    \\u1_u2_dout_r_reg[4]  <= n1390;
    \\u1_u2_dout_r_reg[6]  <= n1395;
    \\u1_u2_dout_r_reg[7]  <= n1400;
    \\u1_u2_dout_r_reg[8]  <= n1405;
    \\u1_u2_dout_r_reg[9]  <= n1410;
    u0_u0_me_cnt_100_ms_reg <= n1415;
    u4_u3_dma_req_in_hold2_reg <= n1420;
    \\u1_mfm_cnt_reg[3]  <= n1425;
    \\u1_mfm_cnt_reg[0]  <= n1430;
    \\u1_u3_size_next_r_reg[0]  <= n1435;
    \\u1_u3_size_next_r_reg[4]  <= n1440;
    \\u1_u3_size_next_r_reg[10]  <= n1445;
    \\u1_u3_size_next_r_reg[11]  <= n1450;
    \\u1_u3_size_next_r_reg[12]  <= n1455;
    \\u1_u3_size_next_r_reg[13]  <= n1460;
    \\u1_u2_adr_cb_reg[2]  <= n1465;
    \\u1_u3_idin_reg[29]  <= n1470;
    \\u1_mfm_cnt_reg[2]  <= n1475;
    u1_u2_word_done_r_reg <= n1480;
    \\u1_u2_dtmp_r_reg[12]  <= n1485;
    u1_u3_int_upid_set_reg <= n1490;
    \\u1_u2_adr_cb_reg[1]  <= n1495;
    \\u1_u3_new_size_reg[11]  <= n1500;
    \\u1_u2_dtmp_r_reg[10]  <= n1505;
    \\u1_u2_dtmp_r_reg[11]  <= n1510;
    \\u1_u2_dtmp_r_reg[13]  <= n1515;
    \\u1_u2_dtmp_r_reg[14]  <= n1520;
    \\u1_u2_dtmp_r_reg[15]  <= n1525;
    \\u1_u2_dtmp_r_reg[17]  <= n1530;
    \\u1_u2_dtmp_r_reg[23]  <= n1535;
    \\u1_u2_dtmp_r_reg[25]  <= n1540;
    \\u1_u2_dtmp_r_reg[24]  <= n1545;
    \\u1_u2_dtmp_r_reg[26]  <= n1550;
    \\u1_u2_dtmp_r_reg[27]  <= n1555;
    \\u1_u2_dtmp_r_reg[29]  <= n1560;
    \\u1_u2_dtmp_r_reg[30]  <= n1565;
    \\u1_u2_dtmp_r_reg[31]  <= n1570;
    \\u1_u2_last_buf_adr_reg[4]  <= n1575;
    \\u1_u2_last_buf_adr_reg[5]  <= n1580;
    \\u1_u2_dtmp_r_reg[28]  <= n1585;
    \\u1_u3_new_size_reg[10]  <= n1590;
    \\u1_u2_dtmp_r_reg[19]  <= n1595;
    \\u1_u2_dtmp_r_reg[16]  <= n1600;
    \\u1_u2_sizu_c_reg[5]  <= n1605;
    u4_nse_err_r_reg <= n1610;
    \\u1_u3_idin_reg[24]  <= n1615;
    \\u1_u2_sizu_c_reg[8]  <= n1620;
    \\u1_u2_dtmp_r_reg[18]  <= n1625;
    \\u1_u2_dtmp_r_reg[20]  <= n1630;
    \\u1_u2_dtmp_r_reg[21]  <= n1635;
    \\u1_u2_dtmp_r_reg[9]  <= n1640;
    \\u1_u2_dtmp_r_reg[0]  <= n1645;
    \\u1_u2_dtmp_r_reg[1]  <= n1650;
    \\u1_u2_dtmp_r_reg[4]  <= n1655;
    \\u1_u2_dtmp_r_reg[5]  <= n1660;
    \\u1_u2_dtmp_r_reg[6]  <= n1665;
    \\u1_u2_dtmp_r_reg[7]  <= n1670;
    \\u1_u2_dtmp_r_reg[3]  <= n1675;
    \\u1_u2_sizu_c_reg[10]  <= n1680;
    \\u1_u2_sizu_c_reg[1]  <= n1685;
    \\u1_u2_sizu_c_reg[2]  <= n1690;
    \\u1_u2_sizu_c_reg[3]  <= n1695;
    \\u1_u2_sizu_c_reg[4]  <= n1700;
    \\u1_u2_sizu_c_reg[6]  <= n1705;
    \\u1_u2_sizu_c_reg[7]  <= n1710;
    \\u1_u2_sizu_c_reg[9]  <= n1715;
    u1_u3_buffer_overflow_reg <= n1720;
    \\u1_u2_last_buf_adr_reg[7]  <= n1725;
    \\u1_u2_dtmp_r_reg[22]  <= n1730;
    \\u1_u2_dtmp_r_reg[2]  <= n1735;
    \\u1_u2_dtmp_r_reg[8]  <= n1740;
    u4_u1_dma_out_buf_avail_reg <= n1745;
    \\u1_frame_no_r_reg[10]  <= n1750;
    \\u1_frame_no_r_reg[4]  <= n1755;
    \\u1_frame_no_r_reg[7]  <= n1760;
    \\u1_frame_no_r_reg[8]  <= n1765;
    \\u1_u3_idin_reg[23]  <= n1770;
    \\u1_frame_no_r_reg[9]  <= n1775;
    u5_wb_ack_o_reg <= n1780;
    \\u1_u2_sizu_c_reg[0]  <= n1785;
    u1_u2_wr_last_reg <= n1790;
    u1_u3_int_seqerr_set_reg <= n1795;
    \\u1_u2_last_buf_adr_reg[2]  <= n1800;
    u1_u2_word_done_reg <= n1805;
    u0_u0_T2_wakeup_reg <= n1810;
    \\u1_frame_no_r_reg[5]  <= n1815;
    u4_u0_dma_out_buf_avail_reg <= n1820;
    u4_u2_dma_out_buf_avail_reg <= n1825;
    u4_u3_dma_out_buf_avail_reg <= n1830;
    u1_u3_nse_err_reg <= n1835;
    \\u1_hms_cnt_reg[1]  <= n1840;
    \\u1_frame_no_r_reg[0]  <= n1845;
    \\u1_frame_no_r_reg[3]  <= n1850;
    \\u1_frame_no_r_reg[1]  <= n1855;
    \\u1_frame_no_r_reg[2]  <= n1860;
    \\u1_frame_no_r_reg[6]  <= n1865;
    \\u1_hms_cnt_reg[2]  <= n1870;
    \\u1_hms_cnt_reg[3]  <= n1875;
    u0_u0_T2_gt_100_uS_reg <= n1880;
    u0_u0_T2_gt_1_0_mS_reg <= n1885;
    u0_u0_T2_gt_1_2_mS_reg <= n1890;
    \\u0_u0_me_ps_reg[1]  <= n1895;
    \\u1_u3_new_size_reg[9]  <= n1900;
    \\u1_u3_new_size_reg[12]  <= n1905;
    \\u1_u2_last_buf_adr_reg[3]  <= n1910;
    \\u0_u0_me_ps2_reg[5]  <= n1915;
    \\u0_u0_me_cnt_reg[4]  <= n1920;
    \\u1_hms_cnt_reg[4]  <= n1925;
    \\u1_u3_idin_reg[21]  <= n1930;
    \\u0_u0_me_ps2_reg[0]  <= n1935;
    \\u0_u0_me_ps2_reg[1]  <= n1940;
    \\u0_u0_me_ps2_reg[2]  <= n1945;
    \\u0_u0_me_ps2_reg[3]  <= n1950;
    \\u0_u0_me_ps2_reg[4]  <= n1955;
    \\u0_u0_me_ps2_reg[6]  <= n1960;
    \\u0_u0_me_ps2_reg[7]  <= n1965;
    \\u0_u0_me_ps_reg[0]  <= n1970;
    \\u0_u0_me_ps_reg[2]  <= n1975;
    \\u0_u0_me_ps_reg[4]  <= n1980;
    \\u0_u0_me_ps_reg[5]  <= n1985;
    \\u0_u0_me_ps_reg[6]  <= n1990;
    \\u1_u3_idin_reg[20]  <= n1995;
    \\u0_u0_me_cnt_reg[0]  <= n2000;
    \\u0_u0_me_cnt_reg[1]  <= n2005;
    \\u0_u0_me_cnt_reg[2]  <= n2010;
    \\u0_u0_me_cnt_reg[3]  <= n2015;
    \\u0_u0_me_cnt_reg[6]  <= n2020;
    \\u0_u0_me_cnt_reg[7]  <= n2025;
    \\u0_u0_me_cnt_reg[5]  <= n2030;
    \\u0_u0_me_ps_reg[3]  <= n2035;
    \\u0_u0_me_ps_reg[7]  <= n2040;
    \\u1_u2_state_reg[0]  <= n2045;
    \\u1_u3_idin_reg[18]  <= n2050;
    \\u4_u0_buf0_reg[28]  <= n2055;
    \\u4_u0_buf0_reg[31]  <= n2060;
    \\u4_u0_buf0_reg[9]  <= n2065;
    \\u4_u0_buf0_reg[27]  <= n2070;
    \\u4_u0_buf0_reg[14]  <= n2075;
    \\u4_u0_buf0_reg[10]  <= n2080;
    \\u4_u0_buf0_reg[13]  <= n2085;
    \\u4_u0_buf1_reg[14]  <= n2090;
    \\u4_u0_buf0_reg[11]  <= n2095;
    \\u4_u0_buf0_reg[15]  <= n2100;
    \\u4_u0_buf0_reg[6]  <= n2105;
    \\u4_u0_buf1_reg[10]  <= n2110;
    \\u4_u0_buf1_reg[13]  <= n2115;
    \\u4_u0_buf0_reg[7]  <= n2120;
    \\u4_u0_buf1_reg[11]  <= n2125;
    \\u4_u0_buf1_reg[15]  <= n2130;
    \\u4_u0_buf1_reg[6]  <= n2135;
    \\u4_u0_buf1_reg[4]  <= n2140;
    \\u4_u0_buf1_reg[5]  <= n2145;
    \\u4_u0_buf1_reg[7]  <= n2150;
    \\u1_hms_cnt_reg[0]  <= n2155;
    \\u1_u3_idin_reg[19]  <= n2160;
    \\u1_u3_new_size_reg[5]  <= n2165;
    \\u4_u0_buf1_reg[28]  <= n2170;
    \\u4_u0_buf1_reg[31]  <= n2175;
    \\u1_u2_state_reg[3]  <= n2180;
    \\u4_u0_buf0_reg[0]  <= n2185;
    \\u4_u0_buf0_reg[18]  <= n2190;
    \\u4_u0_buf0_reg[19]  <= n2195;
    \\u4_u0_buf0_reg[1]  <= n2200;
    \\u4_u0_buf0_reg[20]  <= n2205;
    \\u4_u0_buf0_reg[21]  <= n2210;
    \\u4_u0_buf0_reg[23]  <= n2215;
    \\u4_u0_buf0_reg[24]  <= n2220;
    \\u4_u0_buf0_reg[25]  <= n2225;
    \\u4_u0_buf0_reg[26]  <= n2230;
    \\u4_u0_buf0_reg[30]  <= n2235;
    \\u4_u0_buf0_reg[3]  <= n2240;
    \\u4_u0_buf0_reg[8]  <= n2245;
    \\u4_u1_buf0_reg[28]  <= n2250;
    \\u4_u1_buf0_reg[31]  <= n2255;
    u1_u3_match_r_reg <= n2260;
    \\u1_u3_new_size_reg[8]  <= n2265;
    u5_wb_ack_s2_reg <= n2270;
    \\u1_u3_new_size_reg[7]  <= n2275;
    \\u4_u1_buf0_reg[8]  <= n2280;
    \\u4_u1_buf1_reg[6]  <= n2285;
    \\u4_u2_dma_in_cnt_reg[9]  <= n2290;
    \\u4_u3_dma_in_cnt_reg[9]  <= n2295;
    \\u4_u0_buf1_reg[3]  <= n2300;
    \\u1_u2_last_buf_adr_reg[1]  <= n2305;
    \\u4_u1_buf0_reg[6]  <= n2310;
    \\u4_u1_buf0_reg[14]  <= n2315;
    \\u4_u1_buf0_reg[10]  <= n2320;
    \\u4_u1_buf0_reg[13]  <= n2325;
    \\u4_u1_buf1_reg[14]  <= n2330;
    \\u4_u1_buf0_reg[11]  <= n2335;
    \\u4_u1_buf0_reg[15]  <= n2340;
    \\u4_u1_buf1_reg[10]  <= n2345;
    \\u4_u1_buf1_reg[13]  <= n2350;
    \\u4_u1_buf0_reg[7]  <= n2355;
    \\u4_u1_buf1_reg[11]  <= n2360;
    \\u4_u1_buf1_reg[15]  <= n2365;
    \\u4_u1_buf1_reg[4]  <= n2370;
    \\u4_u1_buf1_reg[7]  <= n2375;
    \\u4_u1_buf1_reg[5]  <= n2380;
    \\u4_u0_buf1_reg[29]  <= n2385;
    \\u4_u0_buf1_reg[21]  <= n2390;
    \\u4_u0_dma_in_cnt_reg[9]  <= n2395;
    \\u4_u1_dma_in_cnt_reg[9]  <= n2400;
    \\u4_u0_dma_in_cnt_reg[11]  <= n2405;
    \\u1_u0_state_reg[2]  <= n2410;
    \\u4_u0_dma_out_cnt_reg[11]  <= n2415;
    \\u4_u0_dma_out_cnt_reg[9]  <= n2420;
    u4_dma_in_buf_sz1_reg <= n2425;
    \\u4_u0_dma_in_cnt_reg[7]  <= n2430;
    \\u4_u0_dma_in_cnt_reg[6]  <= n2435;
    \\u4_u0_dma_out_cnt_reg[6]  <= n2440;
    \\u4_u0_buf1_reg[0]  <= n2445;
    \\u4_u0_buf1_reg[12]  <= n2450;
    \\u4_u0_buf1_reg[16]  <= n2455;
    \\u4_u0_buf1_reg[17]  <= n2460;
    \\u4_u0_buf1_reg[19]  <= n2465;
    \\u4_u0_buf1_reg[1]  <= n2470;
    \\u4_u0_buf1_reg[20]  <= n2475;
    \\u4_u0_buf1_reg[22]  <= n2480;
    \\u4_u0_buf1_reg[24]  <= n2485;
    \\u4_u0_buf1_reg[25]  <= n2490;
    \\u4_u0_buf1_reg[23]  <= n2495;
    \\u4_u0_buf1_reg[27]  <= n2500;
    \\u4_u0_buf1_reg[26]  <= n2505;
    \\u4_u0_buf1_reg[2]  <= n2510;
    \\u4_u0_buf1_reg[30]  <= n2515;
    \\u4_u0_buf1_reg[8]  <= n2520;
    \\u4_u0_buf1_reg[9]  <= n2525;
    \\u4_u1_buf1_reg[28]  <= n2530;
    \\u4_u1_buf1_reg[31]  <= n2535;
    \\u4_u0_dma_in_cnt_reg[0]  <= n2540;
    \\u1_u2_state_reg[4]  <= n2545;
    \\u4_u0_dma_out_cnt_reg[0]  <= n2550;
    \\u4_u0_dma_out_cnt_reg[1]  <= n2555;
    \\u4_u0_dma_out_cnt_reg[2]  <= n2560;
    \\u4_u0_dma_out_cnt_reg[3]  <= n2565;
    \\u4_u1_buf0_reg[16]  <= n2570;
    \\u4_u1_buf0_reg[18]  <= n2575;
    \\u4_u1_buf0_reg[19]  <= n2580;
    \\u4_u1_buf0_reg[1]  <= n2585;
    \\u4_u1_buf0_reg[20]  <= n2590;
    \\u4_u1_buf0_reg[21]  <= n2595;
    \\u4_u1_buf0_reg[23]  <= n2600;
    \\u4_u1_buf0_reg[24]  <= n2605;
    \\u4_u1_buf0_reg[25]  <= n2610;
    \\u4_u1_buf0_reg[27]  <= n2615;
    \\u4_u1_buf0_reg[30]  <= n2620;
    \\u4_u1_buf0_reg[3]  <= n2625;
    \\u4_u1_buf0_reg[9]  <= n2630;
    \\u4_u2_buf0_reg[28]  <= n2635;
    \\u4_u2_buf0_reg[31]  <= n2640;
    u1_frame_no_same_reg <= n2645;
    \\u4_u0_buf1_reg[18]  <= n2650;
    \\u1_u3_new_size_reg[6]  <= n2655;
    \\u4_u1_buf0_reg[26]  <= n2660;
    \\u1_sof_time_reg[2]  <= n2665;
    u5_wb_ack_s1a_reg <= n2670;
    \\u4_u0_buf0_reg[2]  <= n2675;
    \\u4_u2_buf0_reg[8]  <= n2680;
    \\u4_u3_buf0_reg[31]  <= n2685;
    \\u4_u0_buf0_reg[22]  <= n2690;
    \\u4_u2_buf0_reg[12]  <= n2695;
    \\u4_u1_buf1_reg[1]  <= n2700;
    \\u4_u0_dma_out_cnt_reg[8]  <= n2705;
    \\u4_u0_dma_out_cnt_reg[4]  <= n2710;
    \\u4_u1_buf1_reg[9]  <= n2715;
    \\u4_u2_buf0_reg[19]  <= n2720;
    \\u4_u1_buf1_reg[27]  <= n2725;
    \\u4_u1_buf1_reg[23]  <= n2730;
    \\u4_u0_buf0_reg[5]  <= n2735;
    \\u1_sof_time_reg[6]  <= n2740;
    \\u4_u2_buf0_reg[6]  <= n2745;
    \\u4_u2_buf0_reg[11]  <= n2750;
    \\u4_u2_buf0_reg[10]  <= n2755;
    \\u4_u2_buf0_reg[14]  <= n2760;
    \\u4_u2_buf0_reg[13]  <= n2765;
    \\u4_u2_buf1_reg[14]  <= n2770;
    \\u4_u2_buf0_reg[15]  <= n2775;
    \\u4_u2_buf1_reg[10]  <= n2780;
    \\u4_u2_buf1_reg[13]  <= n2785;
    \\u4_u0_buf0_reg[4]  <= n2790;
    \\u4_u2_buf0_reg[7]  <= n2795;
    \\u4_u2_buf1_reg[11]  <= n2800;
    \\u4_u2_buf1_reg[6]  <= n2805;
    \\u4_u2_buf1_reg[4]  <= n2810;
    \\u4_u2_buf1_reg[5]  <= n2815;
    \\u4_u2_buf1_reg[7]  <= n2820;
    \\u1_sof_time_reg[11]  <= n2825;
    \\u4_u0_dma_in_cnt_reg[8]  <= n2830;
    \\u1_sof_time_reg[7]  <= n2835;
    \\u4_u1_dma_in_cnt_reg[11]  <= n2840;
    \\u1_sof_time_reg[0]  <= n2845;
    \\u4_u0_dma_in_cnt_reg[10]  <= n2850;
    \\u4_u1_dma_out_cnt_reg[11]  <= n2855;
    \\u4_u1_dma_out_cnt_reg[9]  <= n2860;
    \\u1_sof_time_reg[10]  <= n2865;
    \\u1_sof_time_reg[1]  <= n2870;
    \\u1_sof_time_reg[3]  <= n2875;
    \\u1_sof_time_reg[4]  <= n2880;
    \\u1_sof_time_reg[5]  <= n2885;
    \\u1_sof_time_reg[9]  <= n2890;
    \\u1_sof_time_reg[8]  <= n2895;
    \\u4_u0_dma_in_cnt_reg[5]  <= n2900;
    \\u4_u0_dma_out_cnt_reg[10]  <= n2905;
    \\u4_u0_dma_out_cnt_reg[7]  <= n2910;
    \\u4_u1_dma_in_cnt_reg[7]  <= n2915;
    \\u4_u0_dma_in_cnt_reg[4]  <= n2920;
    \\u4_u1_dma_in_cnt_reg[6]  <= n2925;
    \\u4_u1_dma_out_cnt_reg[6]  <= n2930;
    \\u4_u1_buf1_reg[0]  <= n2935;
    \\u4_u1_buf1_reg[12]  <= n2940;
    \\u4_u1_buf1_reg[16]  <= n2945;
    \\u4_u1_buf1_reg[17]  <= n2950;
    \\u4_u1_buf1_reg[18]  <= n2955;
    \\u4_u1_buf1_reg[19]  <= n2960;
    \\u4_u1_buf1_reg[20]  <= n2965;
    \\u4_u1_buf1_reg[21]  <= n2970;
    \\u4_u1_buf1_reg[22]  <= n2975;
    \\u4_u1_buf1_reg[24]  <= n2980;
    \\u4_u1_buf1_reg[25]  <= n2985;
    \\u4_u1_buf1_reg[26]  <= n2990;
    \\u4_u1_buf1_reg[2]  <= n2995;
    \\u4_u1_buf1_reg[30]  <= n3000;
    \\u4_u1_buf1_reg[29]  <= n3005;
    \\u4_u1_buf1_reg[3]  <= n3010;
    \\u4_u1_buf1_reg[8]  <= n3015;
    \\u4_u2_buf1_reg[28]  <= n3020;
    \\u4_u2_buf1_reg[31]  <= n3025;
    \\u4_u1_dma_in_cnt_reg[0]  <= n3030;
    \\u4_u0_dma_in_cnt_reg[1]  <= n3035;
    \\u4_u0_dma_in_cnt_reg[2]  <= n3040;
    \\u4_u0_dma_in_cnt_reg[3]  <= n3045;
    \\u4_u0_dma_out_cnt_reg[5]  <= n3050;
    \\u4_u1_dma_out_cnt_reg[0]  <= n3055;
    \\u4_u1_dma_out_cnt_reg[1]  <= n3060;
    \\u4_u1_dma_out_cnt_reg[2]  <= n3065;
    \\u4_u1_dma_out_cnt_reg[3]  <= n3070;
    \\u4_u3_buf0_reg[28]  <= n3075;
    \\u4_u0_buf0_reg[12]  <= n3080;
    \\u4_u0_buf0_reg[16]  <= n3085;
    \\u4_u0_buf0_reg[17]  <= n3090;
    \\u4_u0_buf0_reg[29]  <= n3095;
    \\u4_u2_buf0_reg[0]  <= n3100;
    \\u4_u2_buf0_reg[16]  <= n3105;
    \\u4_u2_buf0_reg[17]  <= n3110;
    \\u4_u2_buf0_reg[18]  <= n3115;
    \\u4_u2_buf0_reg[20]  <= n3120;
    \\u4_u2_buf0_reg[22]  <= n3125;
    \\u4_u2_buf0_reg[24]  <= n3130;
    \\u4_u2_buf0_reg[25]  <= n3135;
    \\u4_u2_buf0_reg[29]  <= n3140;
    \\u4_u2_buf0_reg[1]  <= n3145;
    \\u4_u2_buf0_reg[30]  <= n3150;
    \\u4_u2_buf0_reg[3]  <= n3155;
    \\u4_u2_buf1_reg[15]  <= n3160;
    \\u4_u1_dma_in_cnt_reg[8]  <= n3165;
    \\u4_u1_buf0_reg[2]  <= n3170;
    \\u4_u3_int_stat_reg[0]  <= n3175;
    \\u4_u1_buf0_reg[22]  <= n3180;
    \\u4_u2_buf1_reg[3]  <= n3185;
    \\u4_u2_buf1_reg[20]  <= n3190;
    \\u4_u2_buf1_reg[27]  <= n3195;
    \\u4_u2_buf1_reg[24]  <= n3200;
    \\u4_u1_dma_out_cnt_reg[4]  <= n3205;
    \\u4_u3_buf0_reg[29]  <= n3210;
    \\u4_u2_buf1_reg[17]  <= n3215;
    \\u4_u3_buf0_reg[25]  <= n3220;
    \\u1_u3_new_size_reg[3]  <= n3225;
    \\u4_u3_buf0_reg[21]  <= n3230;
    \\u4_u3_buf0_reg[5]  <= n3235;
    \\u4_u1_buf0_reg[5]  <= n3240;
    \\u4_u1_dma_in_cnt_reg[5]  <= n3245;
    \\u4_u3_buf0_reg[6]  <= n3250;
    \\u4_u3_buf0_reg[10]  <= n3255;
    \\u4_u2_dma_out_cnt_reg[9]  <= n3260;
    \\u4_u3_buf0_reg[14]  <= n3265;
    \\u4_u3_buf0_reg[13]  <= n3270;
    \\u4_u3_buf0_reg[11]  <= n3275;
    \\u4_u3_buf0_reg[15]  <= n3280;
    \\u4_u3_buf0_reg[4]  <= n3285;
    \\u4_u3_buf0_reg[7]  <= n3290;
    \\u4_u1_buf0_reg[4]  <= n3295;
    \\u4_u1_dma_out_cnt_reg[8]  <= n3300;
    \\u5_wb_data_o_reg[1]  <= n3305;
    \\u4_u1_dma_in_cnt_reg[10]  <= n3310;
    \\u4_u2_dma_out_cnt_reg[11]  <= n3315;
    \\u4_u1_dma_out_cnt_reg[10]  <= n3320;
    \\u4_u1_dma_out_cnt_reg[7]  <= n3325;
    \\u4_u2_dma_in_cnt_reg[7]  <= n3330;
    \\u4_u1_dma_in_cnt_reg[4]  <= n3335;
    \\u4_u2_dma_out_cnt_reg[6]  <= n3340;
    \\u4_u2_dma_in_cnt_reg[6]  <= n3345;
    \\u4_u2_buf1_reg[0]  <= n3350;
    \\u4_u2_buf1_reg[12]  <= n3355;
    \\u4_u2_buf1_reg[16]  <= n3360;
    \\u4_u2_buf1_reg[18]  <= n3365;
    \\u4_u2_buf1_reg[19]  <= n3370;
    \\u4_u2_buf1_reg[1]  <= n3375;
    \\u4_u2_buf1_reg[22]  <= n3380;
    \\u4_u2_buf1_reg[23]  <= n3385;
    \\u4_u2_buf1_reg[21]  <= n3390;
    \\u4_u2_buf1_reg[26]  <= n3395;
    \\u4_u2_buf1_reg[25]  <= n3400;
    \\u4_u2_buf1_reg[29]  <= n3405;
    \\u4_u2_buf1_reg[2]  <= n3410;
    \\u4_u2_buf1_reg[30]  <= n3415;
    \\u4_u2_buf1_reg[8]  <= n3420;
    \\u4_u2_buf1_reg[9]  <= n3425;
    \\u4_u2_dma_in_cnt_reg[0]  <= n3430;
    \\u4_u1_dma_in_cnt_reg[2]  <= n3435;
    \\u4_u1_dma_out_cnt_reg[5]  <= n3440;
    \\u4_u2_dma_out_cnt_reg[1]  <= n3445;
    \\u4_u2_dma_out_cnt_reg[2]  <= n3450;
    \\u4_u2_dma_out_cnt_reg[3]  <= n3455;
    \\u4_u2_int_stat_reg[0]  <= n3460;
    \\u4_u3_buf0_reg[0]  <= n3465;
    \\u4_u2_dma_out_cnt_reg[0]  <= n3470;
    \\u4_u3_buf0_reg[16]  <= n3475;
    \\u4_u3_buf0_reg[17]  <= n3480;
    \\u4_u3_buf0_reg[18]  <= n3485;
    \\u4_u3_buf0_reg[19]  <= n3490;
    \\u4_u3_buf0_reg[1]  <= n3495;
    \\u4_u3_buf0_reg[20]  <= n3500;
    \\u4_u3_buf0_reg[12]  <= n3505;
    \\u4_u3_buf0_reg[23]  <= n3510;
    \\u4_u3_buf0_reg[24]  <= n3515;
    \\u4_u3_buf0_reg[22]  <= n3520;
    \\u4_u3_buf0_reg[27]  <= n3525;
    \\u4_u3_buf0_reg[26]  <= n3530;
    \\u4_u3_buf0_reg[2]  <= n3535;
    \\u4_u3_buf0_reg[30]  <= n3540;
    \\u4_u3_buf0_reg[3]  <= n3545;
    \\u4_u3_buf0_reg[8]  <= n3550;
    \\u4_u3_buf0_reg[9]  <= n3555;
    \\u4_u1_buf0_reg[0]  <= n3560;
    \\u4_u1_buf0_reg[12]  <= n3565;
    \\u4_u1_buf0_reg[17]  <= n3570;
    \\u4_u0_int_stat_reg[0]  <= n3575;
    \\u4_u1_buf0_reg[29]  <= n3580;
    \\u4_u1_int_stat_reg[0]  <= n3585;
    \\u4_u1_dma_in_cnt_reg[1]  <= n3590;
    \\u5_state_reg[0]  <= n3595;
    \\u1_u3_new_size_reg[4]  <= n3600;
    \\u4_u2_dma_in_cnt_reg[11]  <= n3605;
    \\u4_u1_dma_in_cnt_reg[3]  <= n3610;
    \\u4_u2_dma_in_cnt_reg[8]  <= n3615;
    \\u4_u3_buf1_reg[7]  <= n3620;
    u1_u3_pid_seq_err_reg <= n3625;
    \\u4_u2_buf0_reg[2]  <= n3630;
    \\u4_u2_dma_out_cnt_reg[4]  <= n3635;
    \\u4_u3_buf1_reg[5]  <= n3640;
    \\u4_u2_buf0_reg[26]  <= n3645;
    u5_wb_ack_s1_reg <= n3650;
    \\u4_u2_dma_out_cnt_reg[7]  <= n3655;
    \\u4_u2_buf0_reg[4]  <= n3660;
    \\u4_u3_buf1_reg[6]  <= n3665;
    \\u5_state_reg[5]  <= n3670;
    \\u4_u3_buf1_reg[14]  <= n3675;
    \\u4_u3_buf1_reg[10]  <= n3680;
    \\u4_u3_buf1_reg[13]  <= n3685;
    \\u4_u3_buf1_reg[11]  <= n3690;
    \\u4_u3_buf1_reg[15]  <= n3695;
    \\u4_u2_buf0_reg[5]  <= n3700;
    \\u4_u3_buf1_reg[4]  <= n3705;
    \\u4_u2_dma_out_cnt_reg[8]  <= n3710;
    \\u5_wb_data_o_reg[3]  <= n3715;
    \\u4_int_srcb_reg[0]  <= n3720;
    \\u4_u2_dma_in_cnt_reg[10]  <= n3725;
    u2_wack_r_reg <= n3730;
    \\u1_u0_state_reg[3]  <= n3735;
    \\u4_u2_dma_in_cnt_reg[5]  <= n3740;
    \\u4_u2_dma_out_cnt_reg[10]  <= n3745;
    \\u4_u2_dma_in_cnt_reg[4]  <= n3750;
    \\u4_u3_buf1_reg[28]  <= n3755;
    \\u4_u3_buf1_reg[31]  <= n3760;
    \\u4_u2_dma_in_cnt_reg[2]  <= n3765;
    \\u4_u2_dma_in_cnt_reg[3]  <= n3770;
    \\u4_u2_dma_out_cnt_reg[5]  <= n3775;
    \\u4_u2_buf0_reg[21]  <= n3780;
    \\u4_u2_buf0_reg[23]  <= n3785;
    \\u4_u2_buf0_reg[27]  <= n3790;
    \\u4_u2_buf0_reg[9]  <= n3795;
    \\u1_u2_state_reg[2]  <= n3800;
    \\u5_wb_data_o_reg[0]  <= n3805;
    \\u4_u2_dma_in_cnt_reg[1]  <= n3810;
    \\u4_u3_dma_out_cnt_reg[9]  <= n3815;
    \\u4_u3_dma_in_cnt_reg[10]  <= n3820;
    \\u4_u3_dma_in_cnt_reg[11]  <= n3825;
    \\u5_wb_data_o_reg[2]  <= n3830;
    \\u4_u3_buf1_reg[25]  <= n3835;
    \\u4_u3_buf1_reg[21]  <= n3840;
    \\u4_u3_dma_out_cnt_reg[3]  <= n3845;
    \\u4_u3_buf1_reg[0]  <= n3850;
    \\u4_u3_buf1_reg[18]  <= n3855;
    u1_u3_buf1_st_max_reg <= n3860;
    \\u1_u3_new_size_reg[2]  <= n3865;
    \\u4_u3_dma_out_cnt_reg[11]  <= n3870;
    \\u4_u3_dma_in_cnt_reg[7]  <= n3875;
    u4_u0_r1_reg <= n3880;
    \\u5_state_reg[4]  <= n3885;
    \\u4_u3_dma_in_cnt_reg[6]  <= n3890;
    \\u4_u3_dma_out_cnt_reg[6]  <= n3895;
    \\u4_u3_buf1_reg[12]  <= n3900;
    \\u4_u3_buf1_reg[16]  <= n3905;
    \\u4_u3_buf1_reg[17]  <= n3910;
    \\u4_u3_buf1_reg[19]  <= n3915;
    \\u4_u3_buf1_reg[1]  <= n3920;
    \\u4_u3_buf1_reg[20]  <= n3925;
    \\u4_u3_buf1_reg[22]  <= n3930;
    \\u4_u3_buf1_reg[23]  <= n3935;
    \\u4_u3_buf1_reg[24]  <= n3940;
    \\u4_u3_buf1_reg[27]  <= n3945;
    \\u4_u3_buf1_reg[26]  <= n3950;
    \\u4_u3_buf1_reg[30]  <= n3955;
    \\u4_u3_buf1_reg[2]  <= n3960;
    \\u4_u3_buf1_reg[9]  <= n3965;
    \\u4_u3_buf1_reg[8]  <= n3970;
    \\u1_u0_state_reg[0]  <= n3975;
    \\u1_u0_state_reg[1]  <= n3980;
    \\u4_u3_dma_in_cnt_reg[0]  <= n3985;
    \\u4_u3_dma_out_cnt_reg[1]  <= n3990;
    \\u4_u3_dma_out_cnt_reg[2]  <= n3995;
    \\u4_u3_dma_out_cnt_reg[0]  <= n4000;
    \\u1_u2_last_buf_adr_reg[0]  <= n4005;
    \\u5_state_reg[1]  <= n4010;
    \\u4_u3_buf1_reg[3]  <= n4015;
    \\u4_u3_buf1_reg[29]  <= n4020;
    u1_clr_sof_time_reg <= n4025;
    u1_frame_no_we_r_reg <= n4030;
    \\u4_u3_dma_out_cnt_reg[5]  <= n4035;
    \\u4_u3_dma_in_cnt_reg[3]  <= n4040;
    \\u4_u3_dma_out_cnt_reg[8]  <= n4045;
    \\u4_u3_dma_out_cnt_reg[4]  <= n4050;
    u4_u1_r1_reg <= n4055;
    \\u4_u3_dma_in_cnt_reg[8]  <= n4060;
    u4_u2_r1_reg <= n4065;
    \\u4_u3_dma_in_cnt_reg[5]  <= n4070;
    \\u4_u3_dma_out_cnt_reg[10]  <= n4075;
    \\u5_state_reg[2]  <= n4080;
    \\u4_u3_dma_in_cnt_reg[4]  <= n4085;
    \\u4_u3_dma_in_cnt_reg[1]  <= n4090;
    \\u4_u3_dma_in_cnt_reg[2]  <= n4095;
    \\u4_u3_dma_out_cnt_reg[7]  <= n4100;
    u4_u3_r1_reg <= n4105;
    \\u1_u0_crc16_sum_reg[1]  <= n4110;
    \\u1_u0_crc16_sum_reg[11]  <= n4115;
    u0_u0_T1_gt_2_5_uS_reg <= n4120;
    u1_u3_to_large_reg <= n4125;
    \\u1_u3_new_size_reg[1]  <= n4130;
    \\u1_u0_crc16_sum_reg[15]  <= n4135;
    \\u4_int_srcb_reg[6]  <= n4140;
    \\u1_u0_crc16_sum_reg[0]  <= n4145;
    \\u1_u0_crc16_sum_reg[10]  <= n4150;
    \\u1_u0_crc16_sum_reg[12]  <= n4155;
    \\u1_u0_crc16_sum_reg[14]  <= n4160;
    \\u1_u0_crc16_sum_reg[3]  <= n4165;
    \\u1_u0_crc16_sum_reg[4]  <= n4170;
    \\u1_u0_crc16_sum_reg[5]  <= n4175;
    \\u1_u0_crc16_sum_reg[7]  <= n4180;
    \\u1_u0_crc16_sum_reg[8]  <= n4185;
    \\u1_u0_crc16_sum_reg[9]  <= n4190;
    \\u1_u3_adr_r_reg[10]  <= n4195;
    \\u1_u3_adr_r_reg[13]  <= n4200;
    \\u1_u3_adr_r_reg[3]  <= n4205;
    \\u1_u3_adr_r_reg[4]  <= n4210;
    u1_u3_to_small_reg <= n4215;
    \\u1_u0_crc16_sum_reg[13]  <= n4220;
    \\u1_u0_crc16_sum_reg[6]  <= n4225;
    \\u1_u0_crc16_sum_reg[2]  <= n4230;
    \\u1_u1_crc16_reg[14]  <= n4235;
    \\u4_buf1_reg[25]  <= n4240;
    \\u4_buf1_reg[29]  <= n4245;
    \\u4_csr_reg[1]  <= n4250;
    \\u4_buf1_reg[21]  <= n4255;
    \\u4_buf1_reg[14]  <= n4260;
    \\u4_dout_reg[1]  <= n4265;
    \\u4_buf1_reg[18]  <= n4270;
    \\u4_csr_reg[5]  <= n4275;
    \\u4_buf0_reg[3]  <= n4280;
    \\u4_buf0_reg[7]  <= n4285;
    \\u4_buf1_reg[10]  <= n4290;
    \\u4_csr_reg[9]  <= n4295;
    \\u0_u0_state_reg[13]  <= n4300;
    \\u0_u0_idle_cnt1_reg[1]  <= n4305;
    \\u4_buf0_reg[29]  <= n4310;
    \\u0_u0_ps_cnt_reg[2]  <= n4315;
    \\u0_u0_idle_cnt1_reg[4]  <= n4320;
    \\u0_u0_idle_cnt1_reg[6]  <= n4325;
    \\u0_u0_idle_cnt1_reg[7]  <= n4330;
    \\u4_csr_reg[30]  <= n4335;
    \\u4_buf0_reg[30]  <= n4340;
    \\u5_wb_data_o_reg[23]  <= n4345;
    \\u4_buf0_reg[21]  <= n4350;
    \\u4_csr_reg[27]  <= n4355;
    \\u4_buf0_reg[25]  <= n4360;
    \\u0_u0_state_reg[11]  <= n4365;
    \\u1_u3_adr_r_reg[12]  <= n4370;
    \\u1_u3_adr_r_reg[16]  <= n4375;
    u1_u3_buf0_st_max_reg <= n4380;
    \\u1_u1_crc16_reg[10]  <= n4385;
    \\u1_u1_crc16_reg[13]  <= n4390;
    \\u1_u1_crc16_reg[12]  <= n4395;
    \\u4_csr_reg[23]  <= n4400;
    \\u5_wb_data_o_reg[22]  <= n4405;
    \\u5_wb_data_o_reg[7]  <= n4410;
    \\u0_u0_idle_cnt1_reg[3]  <= n4415;
    \\u5_wb_data_o_reg[8]  <= n4420;
    u0_u0_T1_gt_3_0_mS_reg <= n4425;
    \\u4_int_srcb_reg[3]  <= n4430;
    \\u0_u0_idle_cnt1_reg[0]  <= n4435;
    \\u0_u0_idle_cnt1_reg[2]  <= n4440;
    u1_u0_rxv2_reg <= n4445;
    \\u0_u0_idle_cnt1_reg[5]  <= n4450;
    \\u0_u0_ps_cnt_reg[0]  <= n4455;
    \\u0_u0_ps_cnt_reg[1]  <= n4460;
    \\u0_u0_ps_cnt_reg[3]  <= n4465;
    resume_req_r_reg <= n4470;
    \\u4_csr_reg[12]  <= n4475;
    \\u4_csr_reg[15]  <= n4480;
    \\u4_csr_reg[17]  <= n4485;
    \\u4_csr_reg[22]  <= n4490;
    \\u4_csr_reg[24]  <= n4495;
    \\u4_csr_reg[25]  <= n4500;
    \\u4_csr_reg[26]  <= n4505;
    \\u4_csr_reg[28]  <= n4510;
    \\u4_csr_reg[29]  <= n4515;
    \\u4_csr_reg[2]  <= n4520;
    \\u4_csr_reg[31]  <= n4525;
    \\u4_csr_reg[3]  <= n4530;
    \\u4_csr_reg[4]  <= n4535;
    \\u4_csr_reg[6]  <= n4540;
    \\u4_csr_reg[7]  <= n4545;
    \\u4_csr_reg[8]  <= n4550;
    \\u4_buf0_reg[0]  <= n4555;
    \\u4_buf0_reg[10]  <= n4560;
    \\u4_buf0_reg[11]  <= n4565;
    \\u4_buf0_reg[12]  <= n4570;
    \\u4_buf0_reg[13]  <= n4575;
    \\u4_buf0_reg[15]  <= n4580;
    \\u4_buf0_reg[16]  <= n4585;
    \\u4_buf0_reg[17]  <= n4590;
    \\u4_buf0_reg[19]  <= n4595;
    \\u4_buf0_reg[1]  <= n4600;
    \\u4_buf0_reg[20]  <= n4605;
    \\u4_buf0_reg[22]  <= n4610;
    \\u4_buf0_reg[23]  <= n4615;
    \\u4_buf0_reg[24]  <= n4620;
    \\u4_buf0_reg[26]  <= n4625;
    \\u4_buf0_reg[27]  <= n4630;
    \\u4_buf0_reg[28]  <= n4635;
    \\u4_buf0_reg[2]  <= n4640;
    \\u4_buf0_reg[31]  <= n4645;
    \\u4_buf0_reg[4]  <= n4650;
    \\u4_buf0_reg[5]  <= n4655;
    \\u4_buf0_reg[6]  <= n4660;
    \\u4_buf0_reg[8]  <= n4665;
    \\u4_buf0_reg[9]  <= n4670;
    \\u4_buf1_reg[0]  <= n4675;
    \\u4_buf1_reg[11]  <= n4680;
    \\u4_buf1_reg[12]  <= n4685;
    \\u4_buf1_reg[13]  <= n4690;
    \\u4_buf1_reg[15]  <= n4695;
    \\u4_buf1_reg[16]  <= n4700;
    \\u4_buf1_reg[17]  <= n4705;
    \\u4_buf1_reg[19]  <= n4710;
    \\u4_buf1_reg[1]  <= n4715;
    \\u4_buf1_reg[20]  <= n4720;
    \\u4_buf1_reg[22]  <= n4725;
    \\u4_buf1_reg[23]  <= n4730;
    \\u4_buf1_reg[24]  <= n4735;
    \\u4_buf1_reg[26]  <= n4740;
    \\u4_buf1_reg[27]  <= n4745;
    \\u4_buf1_reg[28]  <= n4750;
    \\u4_buf1_reg[2]  <= n4755;
    \\u4_buf1_reg[30]  <= n4760;
    \\u4_buf1_reg[31]  <= n4765;
    \\u4_buf1_reg[4]  <= n4770;
    \\u4_buf1_reg[5]  <= n4775;
    \\u4_buf1_reg[6]  <= n4780;
    \\u4_buf1_reg[8]  <= n4785;
    \\u4_buf1_reg[9]  <= n4790;
    \\u4_csr_reg[0]  <= n4795;
    \\u4_csr_reg[11]  <= n4800;
    \\u4_u0_uc_bsel_reg[0]  <= n4805;
    \\u4_u0_uc_bsel_reg[1]  <= n4810;
    \\u4_u0_uc_dpd_reg[0]  <= n4815;
    \\u1_u3_adr_r_reg[11]  <= n4820;
    \\u1_u3_adr_r_reg[14]  <= n4825;
    \\u1_u3_adr_r_reg[15]  <= n4830;
    \\u1_u3_adr_r_reg[6]  <= n4835;
    \\u1_u3_adr_r_reg[7]  <= n4840;
    \\u1_u3_adr_r_reg[8]  <= n4845;
    \\u4_buf0_reg[14]  <= n4850;
    \\u4_buf0_reg[18]  <= n4855;
    u0_u0_T1_gt_5_0_mS_reg <= n4860;
    \\u4_csr_reg[16]  <= n4865;
    u1_u2_rx_data_valid_r_reg <= n4870;
    \\u1_u3_adr_r_reg[9]  <= n4875;
    \\u4_u0_uc_dpd_reg[1]  <= n4880;
    \\u4_csr_reg[10]  <= n4885;
    \\u1_u1_crc16_reg[11]  <= n4890;
    \\u4_buf1_reg[7]  <= n4895;
    \\u4_buf1_reg[3]  <= n4900;
    \\u1_u0_d1_reg[0]  <= n4905;
    \\u5_wb_data_o_reg[25]  <= n4910;
    \\u4_dout_reg[0]  <= n4915;
    \\u1_u0_d1_reg[4]  <= n4920;
    \\u4_dout_reg[2]  <= n4925;
    \\u4_dout_reg[3]  <= n4930;
    \\u1_u0_d0_reg[4]  <= n4935;
    \\u5_wb_data_o_reg[26]  <= n4940;
    \\u1_u0_d0_reg[1]  <= n4945;
    \\u1_u0_d0_reg[3]  <= n4950;
    \\u4_u1_int_stat_reg[4]  <= n4955;
    \\u4_u3_int_stat_reg[4]  <= n4960;
    u4_crc5_err_r_reg <= n4965;
    \\u1_u3_next_dpid_reg[0]  <= n4970;
    \\u1_u3_adr_r_reg[0]  <= n4975;
    u4_u1_dma_in_buf_sz1_reg <= n4980;
    u4_u0_dma_in_buf_sz1_reg <= n4985;
    u4_u3_dma_in_buf_sz1_reg <= n4990;
    u4_u2_dma_in_buf_sz1_reg <= n4995;
    u0_u0_TermSel_reg <= n5000;
    \\u4_int_srcb_reg[5]  <= n5005;
    \\u5_wb_data_o_reg[4]  <= n5010;
    \\u4_u2_int_stat_reg[4]  <= n5015;
    \\u4_u0_int_stat_reg[4]  <= n5020;
    \\u5_wb_data_o_reg[16]  <= n5025;
    \\u5_wb_data_o_reg[24]  <= n5030;
    \\u5_wb_data_o_reg[28]  <= n5035;
    \\u5_wb_data_o_reg[21]  <= n5040;
    \\u5_wb_data_o_reg[20]  <= n5045;
    \\u5_wb_data_o_reg[19]  <= n5050;
    \\u5_wb_data_o_reg[6]  <= n5055;
    \\u5_wb_data_o_reg[5]  <= n5060;
    \\u5_wb_data_o_reg[18]  <= n5065;
    \\u5_wb_data_o_reg[17]  <= n5070;
    \\u4_int_srcb_reg[4]  <= n5075;
    \\u0_u0_state_reg[1]  <= n5080;
    u1_u0_rxv1_reg <= n5085;
    \\u1_u0_d0_reg[0]  <= n5090;
    \\u0_u0_chirp_cnt_reg[1]  <= n5095;
    \\u1_u0_d0_reg[2]  <= n5100;
    \\u0_u0_chirp_cnt_reg[2]  <= n5105;
    \\u1_u0_d0_reg[5]  <= n5110;
    \\u1_u0_d0_reg[6]  <= n5115;
    \\u1_u0_d0_reg[7]  <= n5120;
    \\u1_u0_d1_reg[1]  <= n5125;
    \\u1_u0_d1_reg[2]  <= n5130;
    \\u1_u0_d1_reg[3]  <= n5135;
    \\u1_u0_d1_reg[5]  <= n5140;
    \\u1_u0_d1_reg[6]  <= n5145;
    \\u1_u0_d1_reg[7]  <= n5150;
    \\u1_u0_d2_reg[1]  <= n5155;
    \\u1_u0_d2_reg[2]  <= n5160;
    \\u1_u0_d2_reg[3]  <= n5165;
    \\u1_u0_d2_reg[5]  <= n5170;
    \\u1_u0_d2_reg[6]  <= n5175;
    \\u1_u0_d2_reg[7]  <= n5180;
    \\u0_u0_state_reg[12]  <= n5185;
    \\u4_u1_uc_bsel_reg[0]  <= n5190;
    \\u4_u1_uc_dpd_reg[0]  <= n5195;
    \\u1_u3_adr_r_reg[2]  <= n5200;
    \\u4_u1_uc_bsel_reg[1]  <= n5205;
    \\u4_u1_uc_dpd_reg[1]  <= n5210;
    \\u1_u0_d2_reg[0]  <= n5215;
    \\u1_u0_d2_reg[4]  <= n5220;
    \\u1_u3_adr_r_reg[5]  <= n5225;
    \\u1_u3_adr_r_reg[1]  <= n5230;
    \\u4_u3_dma_out_left_reg[10]  <= n5235;
    \\u4_u0_dma_out_left_reg[10]  <= n5240;
    \\u4_u1_dma_out_left_reg[10]  <= n5245;
    \\u4_u2_dma_out_left_reg[10]  <= n5250;
    \\u5_wb_data_o_reg[30]  <= n5255;
    \\u5_wb_data_o_reg[31]  <= n5260;
    \\u1_u3_idin_reg[17]  <= n5265;
    \\u0_u0_state_reg[9]  <= n5270;
    \\u5_wb_data_o_reg[27]  <= n5275;
    \\u5_wb_data_o_reg[29]  <= n5280;
    \\u4_u3_int_stat_reg[3]  <= n5285;
    \\u4_u0_int_stat_reg[3]  <= n5290;
    \\u4_u1_int_stat_reg[3]  <= n5295;
    u0_u0_T1_st_3_0_mS_reg <= n5300;
    \\u5_wb_data_o_reg[11]  <= n5305;
    \\u5_wb_data_o_reg[9]  <= n5310;
    \\u0_u0_chirp_cnt_reg[0]  <= n5315;
    \\u5_wb_data_o_reg[12]  <= n5320;
    \\u4_u0_int_stat_reg[6]  <= n5325;
    \\u0_u0_state_reg[4]  <= n5330;
    \\u4_u2_uc_bsel_reg[0]  <= n5335;
    \\u4_u2_uc_bsel_reg[1]  <= n5340;
    \\u4_u2_uc_dpd_reg[0]  <= n5345;
    \\u4_u2_int_stat_reg[3]  <= n5350;
    \\u0_u0_state_reg[3]  <= n5355;
    \\u5_wb_data_o_reg[10]  <= n5360;
    \\u4_u2_uc_dpd_reg[1]  <= n5365;
    u1_u0_data_valid0_reg <= n5370;
    u0_u0_XcvSelect_reg <= n5375;
    \\u0_u0_OpMode_reg[1]  <= n5380;
    \\u4_int_srcb_reg[8]  <= n5385;
    \\u4_u3_dma_out_left_reg[9]  <= n5390;
    \\u4_u0_dma_out_left_reg[9]  <= n5395;
    \\u4_u1_dma_out_left_reg[9]  <= n5400;
    \\u4_u2_dma_out_left_reg[9]  <= n5405;
    \\u1_u3_this_dpid_reg[0]  <= n5410;
    \\u1_u3_next_dpid_reg[1]  <= n5415;
    \\u0_u0_state_reg[10]  <= n5420;
    \\u0_u0_OpMode_reg[0]  <= n5425;
    \\u4_int_srcb_reg[7]  <= n5430;
    \\u4_int_srcb_reg[1]  <= n5435;
    \\u5_wb_data_o_reg[13]  <= n5440;
    \\u5_wb_data_o_reg[15]  <= n5445;
    \\u4_u1_int_stat_reg[6]  <= n5450;
    \\u4_u0_int_stat_reg[1]  <= n5455;
    \\u4_u3_uc_bsel_reg[0]  <= n5460;
    \\u4_u3_uc_bsel_reg[1]  <= n5465;
    \\u4_u3_uc_dpd_reg[0]  <= n5470;
    \\u0_u0_state_reg[6]  <= n5475;
    u1_u3_buf1_set_reg <= n5480;
    \\u1_u3_adr_reg[0]  <= n5485;
    \\u1_u3_adr_reg[1]  <= n5490;
    \\u1_u3_adr_reg[2]  <= n5495;
    \\u1_u3_adr_reg[12]  <= n5500;
    \\u1_u3_adr_reg[13]  <= n5505;
    \\u1_u3_adr_reg[14]  <= n5510;
    \\u1_u3_adr_reg[15]  <= n5515;
    \\u1_u3_adr_reg[16]  <= n5520;
    \\u1_u3_adr_reg[3]  <= n5525;
    \\u1_u3_adr_reg[4]  <= n5530;
    \\u1_u3_adr_reg[5]  <= n5535;
    \\u1_u3_adr_reg[6]  <= n5540;
    \\u1_u3_adr_reg[7]  <= n5545;
    \\u1_u3_adr_reg[8]  <= n5550;
    \\u1_u3_adr_reg[9]  <= n5555;
    \\u1_u3_adr_reg[10]  <= n5560;
    \\u1_u3_adr_reg[11]  <= n5565;
    \\u4_u3_uc_dpd_reg[1]  <= n5570;
    u4_intb_reg <= n5575;
    \\u1_u3_this_dpid_reg[1]  <= n5580;
    \\u1_u0_token0_reg[6]  <= n5585;
    u1_u2_send_data_r_reg <= n5590;
    \\u0_u0_state_reg[5]  <= n5595;
    u4_inta_reg <= n5600;
    \\u0_u0_state_reg[14]  <= n5605;
    \\u4_u0_csr0_reg[2]  <= n5610;
    \\u4_u0_csr0_reg[4]  <= n5615;
    \\u4_u0_csr1_reg[1]  <= n5620;
    \\u4_u0_csr1_reg[2]  <= n5625;
    \\u4_u0_csr1_reg[3]  <= n5630;
    \\u4_u1_csr0_reg[2]  <= n5635;
    \\u4_u1_csr0_reg[5]  <= n5640;
    \\u4_u1_csr0_reg[9]  <= n5645;
    \\u4_u1_csr1_reg[10]  <= n5650;
    \\u4_u2_csr0_reg[0]  <= n5655;
    \\u4_u2_csr0_reg[2]  <= n5660;
    \\u4_u2_csr0_reg[6]  <= n5665;
    \\u4_u2_csr0_reg[9]  <= n5670;
    \\u4_u2_int_stat_reg[1]  <= n5675;
    \\u4_u1_buf0_orig_reg[30]  <= n5680;
    \\u4_u1_int_stat_reg[1]  <= n5685;
    u0_u0_usb_suspend_reg <= n5690;
    \\u1_u0_token0_reg[0]  <= n5695;
    \\u1_u0_token0_reg[1]  <= n5700;
    \\u1_u0_token0_reg[3]  <= n5705;
    \\u1_u0_token0_reg[4]  <= n5710;
    \\u1_u0_token0_reg[5]  <= n5715;
    \\u1_u0_token0_reg[7]  <= n5720;
    \\u0_u0_state_reg[7]  <= n5725;
    \\u0_u0_state_reg[2]  <= n5730;
    u1_u3_buf0_set_reg <= n5735;
    \\u4_u2_int_stat_reg[6]  <= n5740;
    \\u1_u0_token0_reg[2]  <= n5745;
    \\u0_u0_state_reg[8]  <= n5750;
    \\u4_u3_csr1_reg[2]  <= n5755;
    u4_u3_ots_stop_reg <= n5760;
    \\u4_u0_buf0_orig_reg[7]  <= n5765;
    \\u4_u1_csr1_reg[3]  <= n5770;
    \\u4_u0_buf0_orig_reg[8]  <= n5775;
    \\u4_u2_buf0_orig_reg[27]  <= n5780;
    \\u4_u2_buf0_orig_reg[28]  <= n5785;
    \\u1_u0_pid_reg[6]  <= n5790;
    \\u4_dout_reg[22]  <= n5795;
    \\u4_dout_reg[23]  <= n5800;
    \\u4_dout_reg[7]  <= n5805;
    \\u4_u2_buf0_orig_reg[14]  <= n5810;
    \\u4_u1_buf0_orig_reg[13]  <= n5815;
    \\u4_u2_buf0_orig_reg[1]  <= n5820;
    \\u4_u1_buf0_orig_reg[0]  <= n5825;
    \\u4_u2_buf0_orig_reg[23]  <= n5830;
    \\u4_u0_buf0_orig_reg[4]  <= n5835;
    \\u4_funct_adr_reg[5]  <= n5840;
    \\u4_funct_adr_reg[3]  <= n5845;
    \\u4_u3_csr1_reg[6]  <= n5850;
    \\u4_u2_buf0_orig_reg[16]  <= n5855;
    \\u4_dout_reg[8]  <= n5860;
    \\u4_u0_buf0_orig_reg[6]  <= n5865;
    \\u4_u3_csr1_reg[10]  <= n5870;
    \\u4_u0_buf0_orig_reg[31]  <= n5875;
    \\u4_u1_csr0_reg[8]  <= n5880;
    \\u4_u0_buf0_orig_reg[20]  <= n5885;
    \\u4_u1_csr1_reg[1]  <= n5890;
    \\u1_u0_pid_reg[7]  <= n5895;
    \\u4_u1_csr1_reg[11]  <= n5900;
    \\u4_u3_csr0_reg[7]  <= n5905;
    \\u4_u0_buf0_orig_reg[28]  <= n5910;
    \\u4_u1_csr0_reg[6]  <= n5915;
    \\u4_u1_csr0_reg[12]  <= n5920;
    \\u4_u2_buf0_orig_reg[10]  <= n5925;
    \\u4_u2_buf0_orig_reg[12]  <= n5930;
    \\u4_u0_buf0_orig_reg[22]  <= n5935;
    \\u1_u2_state_reg[6]  <= n5940;
    \\u4_u0_buf0_orig_reg[26]  <= n5945;
    \\u1_u2_state_reg[1]  <= n5950;
    \\u1_u2_state_reg[5]  <= n5955;
    \\u4_u1_csr0_reg[1]  <= n5960;
    \\u4_u0_buf0_orig_reg[24]  <= n5965;
    \\u4_funct_adr_reg[0]  <= n5970;
    \\u4_funct_adr_reg[1]  <= n5975;
    \\u4_funct_adr_reg[2]  <= n5980;
    \\u4_funct_adr_reg[4]  <= n5985;
    \\u4_funct_adr_reg[6]  <= n5990;
    u1_u3_out_to_small_r_reg <= n5995;
    u4_u2_ots_stop_reg <= n6000;
    u1_u2_mack_r_reg <= n6005;
    \\u4_u3_csr0_reg[10]  <= n6010;
    \\u4_u3_csr0_reg[12]  <= n6015;
    \\u4_u3_csr0_reg[1]  <= n6020;
    \\u4_u3_csr0_reg[2]  <= n6025;
    \\u4_u3_csr0_reg[4]  <= n6030;
    \\u4_u3_csr0_reg[5]  <= n6035;
    \\u4_u3_csr0_reg[6]  <= n6040;
    \\u4_u3_csr0_reg[8]  <= n6045;
    \\u4_u3_csr0_reg[9]  <= n6050;
    \\u4_u3_csr1_reg[0]  <= n6055;
    \\u4_u3_csr1_reg[11]  <= n6060;
    \\u4_u3_csr1_reg[12]  <= n6065;
    \\u4_u3_csr1_reg[1]  <= n6070;
    \\u4_u3_csr1_reg[3]  <= n6075;
    \\u4_u3_csr1_reg[4]  <= n6080;
    \\u4_u3_csr1_reg[5]  <= n6085;
    \\u4_u3_csr1_reg[9]  <= n6090;
    \\u4_u0_csr0_reg[10]  <= n6095;
    \\u4_u0_csr0_reg[12]  <= n6100;
    \\u4_u0_csr0_reg[6]  <= n6105;
    \\u4_u0_csr1_reg[0]  <= n6110;
    \\u4_u0_csr1_reg[5]  <= n6115;
    \\u4_u0_csr1_reg[9]  <= n6120;
    u4_u0_ots_stop_reg <= n6125;
    \\u4_u1_csr0_reg[0]  <= n6130;
    \\u4_u1_csr0_reg[10]  <= n6135;
    \\u4_u1_csr0_reg[11]  <= n6140;
    \\u4_u1_csr0_reg[4]  <= n6145;
    \\u4_u1_csr0_reg[7]  <= n6150;
    \\u4_u1_csr1_reg[0]  <= n6155;
    \\u4_u1_csr1_reg[12]  <= n6160;
    \\u4_u1_csr1_reg[2]  <= n6165;
    \\u4_u1_csr1_reg[4]  <= n6170;
    \\u4_u1_csr1_reg[5]  <= n6175;
    \\u4_u1_csr1_reg[6]  <= n6180;
    \\u4_u1_csr1_reg[9]  <= n6185;
    u4_u1_ots_stop_reg <= n6190;
    \\u4_u2_csr0_reg[10]  <= n6195;
    \\u4_u2_csr0_reg[12]  <= n6200;
    \\u4_u2_csr0_reg[4]  <= n6205;
    \\u4_u2_csr0_reg[7]  <= n6210;
    \\u4_u2_csr1_reg[0]  <= n6215;
    \\u4_u2_csr1_reg[11]  <= n6220;
    \\u4_u2_csr1_reg[1]  <= n6225;
    \\u4_u2_csr1_reg[3]  <= n6230;
    \\u4_u2_csr1_reg[6]  <= n6235;
    \\u4_u2_csr1_reg[5]  <= n6240;
    \\u4_u3_buf0_orig_reg[0]  <= n6245;
    \\u4_u3_buf0_orig_reg[12]  <= n6250;
    \\u4_u3_buf0_orig_reg[14]  <= n6255;
    \\u4_u3_buf0_orig_reg[15]  <= n6260;
    \\u4_u3_buf0_orig_reg[16]  <= n6265;
    \\u4_u3_buf0_orig_reg[21]  <= n6270;
    \\u4_u3_buf0_orig_reg[22]  <= n6275;
    \\u4_u3_buf0_orig_reg[23]  <= n6280;
    \\u4_u3_buf0_orig_reg[24]  <= n6285;
    \\u4_u3_buf0_orig_reg[26]  <= n6290;
    \\u4_u3_buf0_orig_reg[28]  <= n6295;
    \\u4_u3_buf0_orig_reg[30]  <= n6300;
    \\u4_u3_buf0_orig_reg[31]  <= n6305;
    \\u4_u3_buf0_orig_reg[5]  <= n6310;
    \\u4_u3_buf0_orig_reg[8]  <= n6315;
    \\u4_u3_csr1_reg[8]  <= n6320;
    \\u4_u3_int_stat_reg[1]  <= n6325;
    \\u4_u0_buf0_orig_reg[10]  <= n6330;
    \\u4_u0_buf0_orig_reg[11]  <= n6335;
    \\u4_u0_buf0_orig_reg[12]  <= n6340;
    \\u4_u0_buf0_orig_reg[14]  <= n6345;
    \\u4_u0_buf0_orig_reg[16]  <= n6350;
    \\u4_u0_buf0_orig_reg[18]  <= n6355;
    \\u4_u0_buf0_orig_reg[1]  <= n6360;
    \\u4_u0_buf0_orig_reg[21]  <= n6365;
    \\u4_u0_buf0_orig_reg[23]  <= n6370;
    \\u4_u0_buf0_orig_reg[25]  <= n6375;
    \\u4_u0_buf0_orig_reg[27]  <= n6380;
    \\u4_u0_buf0_orig_reg[29]  <= n6385;
    \\u4_u0_buf0_orig_reg[2]  <= n6390;
    \\u4_u0_buf0_orig_reg[30]  <= n6395;
    \\u4_u0_buf0_orig_reg[3]  <= n6400;
    \\u4_u0_buf0_orig_reg[5]  <= n6405;
    \\u4_u0_buf0_orig_reg[9]  <= n6410;
    \\u4_u3_buf0_orig_reg[9]  <= n6415;
    \\u4_u0_csr1_reg[8]  <= n6420;
    \\u4_u1_buf0_orig_reg[10]  <= n6425;
    \\u4_u1_buf0_orig_reg[11]  <= n6430;
    \\u4_u1_buf0_orig_reg[12]  <= n6435;
    \\u4_u1_buf0_orig_reg[14]  <= n6440;
    \\u4_u1_buf0_orig_reg[15]  <= n6445;
    \\u4_u1_buf0_orig_reg[16]  <= n6450;
    \\u4_u1_buf0_orig_reg[18]  <= n6455;
    \\u4_u1_buf0_orig_reg[19]  <= n6460;
    \\u4_u1_buf0_orig_reg[1]  <= n6465;
    \\u4_u1_buf0_orig_reg[21]  <= n6470;
    \\u4_u1_buf0_orig_reg[22]  <= n6475;
    \\u4_u1_buf0_orig_reg[23]  <= n6480;
    \\u4_u1_buf0_orig_reg[25]  <= n6485;
    \\u4_u1_buf0_orig_reg[26]  <= n6490;
    \\u4_u1_buf0_orig_reg[27]  <= n6495;
    \\u4_u1_buf0_orig_reg[2]  <= n6500;
    \\u4_u1_buf0_orig_reg[29]  <= n6505;
    \\u4_u1_buf0_orig_reg[3]  <= n6510;
    \\u4_u1_buf0_orig_reg[4]  <= n6515;
    \\u4_u1_buf0_orig_reg[5]  <= n6520;
    \\u4_u1_buf0_orig_reg[7]  <= n6525;
    \\u4_u1_csr1_reg[8]  <= n6530;
    \\u4_u2_buf0_orig_reg[0]  <= n6535;
    \\u4_u2_buf0_orig_reg[11]  <= n6540;
    \\u4_u2_buf0_orig_reg[13]  <= n6545;
    \\u4_u2_buf0_orig_reg[15]  <= n6550;
    \\u4_u2_buf0_orig_reg[17]  <= n6555;
    \\u4_u2_buf0_orig_reg[18]  <= n6560;
    \\u4_u2_buf0_orig_reg[19]  <= n6565;
    \\u4_u2_buf0_orig_reg[20]  <= n6570;
    \\u4_u2_buf0_orig_reg[21]  <= n6575;
    \\u4_u2_buf0_orig_reg[22]  <= n6580;
    \\u4_u2_buf0_orig_reg[24]  <= n6585;
    \\u4_u2_buf0_orig_reg[25]  <= n6590;
    \\u4_u2_buf0_orig_reg[26]  <= n6595;
    \\u4_u2_buf0_orig_reg[2]  <= n6600;
    \\u4_u2_buf0_orig_reg[31]  <= n6605;
    \\u4_u2_buf0_orig_reg[4]  <= n6610;
    \\u4_u2_buf0_orig_reg[7]  <= n6615;
    \\u4_u2_buf0_orig_reg[9]  <= n6620;
    \\u4_u2_csr1_reg[8]  <= n6625;
    \\u5_wb_data_o_reg[14]  <= n6630;
    \\u1_u0_pid_reg[0]  <= n6635;
    \\u1_u0_pid_reg[1]  <= n6640;
    \\u1_u0_pid_reg[2]  <= n6645;
    \\u1_u0_pid_reg[4]  <= n6650;
    \\u1_u0_pid_reg[5]  <= n6655;
    \\u4_u2_buf0_orig_reg[29]  <= n6660;
    u1_u0_token_valid_str1_reg <= n6665;
    u4_match_r1_reg <= n6670;
    \\u4_u0_csr0_reg[0]  <= n6675;
    \\u1_u0_pid_reg[3]  <= n6680;
    \\u4_u3_csr0_reg[0]  <= n6685;
    \\u4_u1_buf0_orig_reg[31]  <= n6690;
    \\u4_u0_buf0_orig_reg[13]  <= n6695;
    \\u4_u1_buf0_orig_reg[9]  <= n6700;
    \\u4_u0_buf0_orig_reg[19]  <= n6705;
    \\u4_u2_csr1_reg[9]  <= n6710;
    \\u4_u3_csr0_reg[11]  <= n6715;
    \\u4_u1_buf0_orig_reg[6]  <= n6720;
    \\u4_u1_buf0_orig_reg[8]  <= n6725;
    \\u4_u0_buf0_orig_reg[15]  <= n6730;
    \\u4_u0_buf0_orig_reg[17]  <= n6735;
    \\u4_u1_buf0_orig_reg[17]  <= n6740;
    \\u4_u1_buf0_orig_reg[28]  <= n6745;
    u1_u2_wr_done_reg <= n6750;
    u1_u2_idma_done_reg <= n6755;
    \\u4_u0_csr1_reg[10]  <= n6760;
    \\u4_u2_csr1_reg[4]  <= n6765;
    \\u4_u0_buf0_orig_reg[0]  <= n6770;
    \\u4_u2_csr1_reg[2]  <= n6775;
    \\u4_u0_csr1_reg[11]  <= n6780;
    \\u4_u0_csr1_reg[12]  <= n6785;
    \\u4_u2_csr0_reg[5]  <= n6790;
    \\u4_u2_csr1_reg[12]  <= n6795;
    \\u4_u0_csr1_reg[4]  <= n6800;
    \\u4_u2_csr1_reg[10]  <= n6805;
    \\u4_u0_csr1_reg[6]  <= n6810;
    \\u4_u3_buf0_orig_reg[3]  <= n6815;
    \\u4_u1_buf0_orig_reg[24]  <= n6820;
    \\u4_u2_csr0_reg[8]  <= n6825;
    \\u4_u2_buf0_orig_reg[30]  <= n6830;
    \\u4_u0_csr0_reg[9]  <= n6835;
    \\u4_u0_csr0_reg[11]  <= n6840;
    \\u4_u3_buf0_orig_reg[29]  <= n6845;
    \\u4_u0_csr0_reg[8]  <= n6850;
    \\u4_u2_csr0_reg[1]  <= n6855;
    \\u4_u0_csr0_reg[5]  <= n6860;
    \\u4_u2_csr0_reg[11]  <= n6865;
    \\u4_u0_csr0_reg[7]  <= n6870;
    \\u4_u3_buf0_orig_reg[25]  <= n6875;
    \\u4_u1_buf0_orig_reg[20]  <= n6880;
    \\u4_u0_csr0_reg[3]  <= n6885;
    \\u4_u2_buf0_orig_reg[6]  <= n6890;
    \\u4_u2_buf0_orig_reg[8]  <= n6895;
    \\u4_u0_csr0_reg[1]  <= n6900;
    \\u4_u2_buf0_orig_reg[5]  <= n6905;
    \\u4_u2_buf0_orig_reg[3]  <= n6910;
    \\u4_u3_buf0_orig_reg[20]  <= n6915;
    \\u4_u3_buf0_orig_reg[18]  <= n6920;
    \\u1_u0_token1_reg[6]  <= n6925;
    \\u4_dout_reg[4]  <= n6930;
    \\u4_inta_msk_reg[8]  <= n6935;
    \\u4_intb_msk_reg[3]  <= n6940;
    \\u4_inta_msk_reg[2]  <= n6945;
    \\u4_inta_msk_reg[4]  <= n6950;
    \\u4_inta_msk_reg[0]  <= n6955;
    \\u4_u3_buf0_orig_reg[1]  <= n6960;
    \\u4_dout_reg[20]  <= n6965;
    \\u4_dout_reg[16]  <= n6970;
    \\u4_dout_reg[17]  <= n6975;
    \\u4_dout_reg[18]  <= n6980;
    \\u4_dout_reg[19]  <= n6985;
    \\u4_dout_reg[21]  <= n6990;
    \\u4_dout_reg[24]  <= n6995;
    \\u4_dout_reg[25]  <= n7000;
    \\u4_dout_reg[26]  <= n7005;
    \\u4_dout_reg[28]  <= n7010;
    \\u4_dout_reg[5]  <= n7015;
    \\u4_dout_reg[6]  <= n7020;
    \\u4_u3_buf0_orig_reg[17]  <= n7025;
    \\u4_u3_dma_out_left_reg[8]  <= n7030;
    \\u4_u0_dma_out_left_reg[8]  <= n7035;
    \\u4_u1_dma_out_left_reg[8]  <= n7040;
    \\u4_u2_dma_out_left_reg[8]  <= n7045;
    \\u4_u1_csr0_reg[3]  <= n7050;
    \\u4_u3_buf0_orig_reg[11]  <= n7055;
    \\u4_u3_buf0_orig_reg[13]  <= n7060;
    \\u1_u0_token1_reg[0]  <= n7065;
    \\u4_u3_int_stat_reg[6]  <= n7070;
    suspend_clr_wr_reg <= n7075;
    \\u4_u3_buf0_orig_reg[10]  <= n7080;
    \\u1_u0_token1_reg[1]  <= n7085;
    \\u1_u0_token1_reg[2]  <= n7090;
    \\u4_inta_msk_reg[1]  <= n7095;
    \\u4_inta_msk_reg[3]  <= n7100;
    \\u4_inta_msk_reg[5]  <= n7105;
    \\u4_inta_msk_reg[6]  <= n7110;
    \\u4_inta_msk_reg[7]  <= n7115;
    \\u4_intb_msk_reg[0]  <= n7120;
    \\u4_intb_msk_reg[1]  <= n7125;
    \\u4_intb_msk_reg[2]  <= n7130;
    \\u4_intb_msk_reg[4]  <= n7135;
    \\u4_intb_msk_reg[5]  <= n7140;
    \\u4_intb_msk_reg[6]  <= n7145;
    \\u4_intb_msk_reg[8]  <= n7150;
    \\u4_u3_buf0_orig_reg[19]  <= n7155;
    \\u4_u3_buf0_orig_reg[4]  <= n7160;
    \\u4_u3_buf0_orig_reg[7]  <= n7165;
    \\u1_u0_token1_reg[3]  <= n7170;
    \\u1_u0_token1_reg[4]  <= n7175;
    \\u1_u0_token1_reg[5]  <= n7180;
    \\u1_u0_token1_reg[7]  <= n7185;
    \\u4_u3_csr0_reg[3]  <= n7190;
    \\u4_intb_msk_reg[7]  <= n7195;
    \\u4_u0_dma_out_left_reg[11]  <= n7200;
    \\u4_u1_dma_out_left_reg[11]  <= n7205;
    \\u4_u2_csr0_reg[3]  <= n7210;
    \\u4_u3_buf0_orig_reg[6]  <= n7215;
    \\u4_u3_buf0_orig_reg[2]  <= n7220;
    u0_u0_idle_long_reg <= n7225;
    \\u4_u3_buf0_orig_reg[27]  <= n7230;
    \\u4_u3_ienb_reg[5]  <= n7235;
    \\u4_u3_iena_reg[3]  <= n7240;
    \\u4_u1_iena_reg[4]  <= n7245;
    \\u4_u3_ienb_reg[2]  <= n7250;
    \\u4_u3_ienb_reg[4]  <= n7255;
    \\u4_u1_iena_reg[5]  <= n7260;
    \\u4_u3_iena_reg[4]  <= n7265;
    \\u4_u3_ienb_reg[3]  <= n7270;
    \\u4_u3_ienb_reg[1]  <= n7275;
    \\u4_u3_iena_reg[5]  <= n7280;
    \\u4_u3_ienb_reg[0]  <= n7285;
    \\u1_u3_new_size_reg[0]  <= n7290;
    \\u4_u1_iena_reg[0]  <= n7295;
    \\u4_u0_csr1_reg[7]  <= n7300;
    \\u4_u3_csr1_reg[7]  <= n7305;
    \\u4_u1_iena_reg[1]  <= n7310;
    \\u4_u3_iena_reg[1]  <= n7315;
    \\u4_u1_iena_reg[3]  <= n7320;
    \\u4_dout_reg[29]  <= n7325;
    \\u4_dout_reg[30]  <= n7330;
    \\u4_dout_reg[31]  <= n7335;
    \\u4_dout_reg[27]  <= n7340;
    \\u4_u1_csr1_reg[7]  <= n7345;
    \\u1_u2_state_reg[7]  <= n7350;
    \\u4_dout_reg[10]  <= n7355;
    \\u4_dout_reg[11]  <= n7360;
    \\u4_dout_reg[9]  <= n7365;
    \\u4_u2_iena_reg[1]  <= n7370;
    \\u4_u2_iena_reg[3]  <= n7375;
    \\u4_u2_iena_reg[5]  <= n7380;
    \\u4_u2_ienb_reg[0]  <= n7385;
    \\u4_u2_ienb_reg[1]  <= n7390;
    \\u4_u2_ienb_reg[4]  <= n7395;
    \\u4_u2_ienb_reg[3]  <= n7400;
    \\u4_u3_iena_reg[0]  <= n7405;
    \\u4_u3_iena_reg[2]  <= n7410;
    \\u4_u0_iena_reg[1]  <= n7415;
    \\u4_u0_iena_reg[2]  <= n7420;
    \\u4_u0_iena_reg[3]  <= n7425;
    \\u4_u0_iena_reg[5]  <= n7430;
    \\u4_u0_ienb_reg[1]  <= n7435;
    \\u4_u0_ienb_reg[4]  <= n7440;
    \\u4_u0_ienb_reg[3]  <= n7445;
    \\u4_u1_iena_reg[2]  <= n7450;
    \\u4_u1_ienb_reg[4]  <= n7455;
    \\u4_dout_reg[12]  <= n7460;
    \\u4_u0_ienb_reg[5]  <= n7465;
    \\u4_u1_ienb_reg[0]  <= n7470;
    \\u4_u0_ienb_reg[2]  <= n7475;
    \\u4_u0_iena_reg[4]  <= n7480;
    \\u4_u0_ienb_reg[0]  <= n7485;
    \\u4_u3_dma_out_left_reg[11]  <= n7490;
    \\u4_u2_dma_out_left_reg[11]  <= n7495;
    \\u4_u2_iena_reg[0]  <= n7500;
    \\u5_state_reg[3]  <= n7505;
    \\u4_u1_ienb_reg[1]  <= n7510;
    \\u4_u2_ienb_reg[5]  <= n7515;
    \\u4_u0_iena_reg[0]  <= n7520;
    \\u4_u2_ienb_reg[2]  <= n7525;
    \\u4_u2_iena_reg[2]  <= n7530;
    \\u4_u2_iena_reg[4]  <= n7535;
    \\u4_u1_ienb_reg[2]  <= n7540;
    u1_u2_rx_data_done_r2_reg <= n7545;
    u1_u2_wr_done_r_reg <= n7550;
    \\u4_u1_ienb_reg[3]  <= n7555;
    \\u4_u1_ienb_reg[5]  <= n7560;
    \\u4_u2_csr1_reg[7]  <= n7565;
    \\u4_dout_reg[13]  <= n7570;
    \\u4_dout_reg[15]  <= n7575;
    u1_u3_tx_data_to_reg <= n7580;
    u1_u3_rx_ack_to_reg <= n7585;
    u1_u2_rx_data_done_r_reg <= n7590;
    \\u4_utmi_vend_ctrl_r_reg[2]  <= n7595;
    \\u4_u1_dma_out_left_reg[7]  <= n7600;
    \\u4_u1_buf0_orig_m3_reg[11]  <= n7605;
    \\u1_u1_state_reg[2]  <= n7610;
    \\u4_utmi_vend_ctrl_r_reg[1]  <= n7615;
    u4_int_src_re_reg <= n7620;
    \\u4_utmi_vend_ctrl_r_reg[0]  <= n7625;
    \\u4_utmi_vend_ctrl_r_reg[3]  <= n7630;
    u1_u0_token_valid_r1_reg <= n7635;
    u4_utmi_vend_wr_r_reg <= n7640;
    \\u1_u1_state_reg[3]  <= n7645;
    u4_u0_ep_match_r_reg <= n7650;
    \\u4_u3_dma_out_left_reg[7]  <= n7655;
    \\u4_u0_dma_out_left_reg[7]  <= n7660;
    \\u4_u2_dma_out_left_reg[7]  <= n7665;
    \\u4_u0_buf0_orig_m3_reg[11]  <= n7670;
    \\u4_u0_buf0_orig_m3_reg[9]  <= n7675;
    \\u4_u2_buf0_orig_m3_reg[9]  <= n7680;
    u4_u1_int_re_reg <= n7685;
    \\u4_u0_buf0_orig_m3_reg[10]  <= n7690;
    u4_u2_int_re_reg <= n7695;
    u4_u0_int_re_reg <= n7700;
    \\u4_u2_buf0_orig_m3_reg[10]  <= n7705;
    \\u4_u3_dma_out_left_reg[6]  <= n7710;
    \\u4_u0_dma_out_left_reg[6]  <= n7715;
    \\u4_u1_dma_out_left_reg[6]  <= n7720;
    \\u4_dout_reg[14]  <= n7725;
    \\u4_u2_dma_out_left_reg[6]  <= n7730;
    u4_u1_ep_match_r_reg <= n7735;
    \\u4_u3_buf0_orig_m3_reg[11]  <= n7740;
    \\u4_u2_buf0_orig_m3_reg[11]  <= n7745;
    \\u4_u0_dma_out_left_reg[5]  <= n7750;
    \\u4_u3_dma_out_left_reg[5]  <= n7755;
    \\u4_u1_dma_out_left_reg[5]  <= n7760;
    \\u4_u2_dma_out_left_reg[5]  <= n7765;
    \\u4_u1_buf0_orig_m3_reg[7]  <= n7770;
    \\u4_u1_buf0_orig_m3_reg[8]  <= n7775;
    \\u4_u1_buf0_orig_m3_reg[10]  <= n7780;
    u0_u0_usb_attached_reg <= n7785;
    u1_u3_in_token_reg <= n7790;
    u4_u2_ep_match_r_reg <= n7795;
    \\u1_u3_tx_data_to_cnt_reg[4]  <= n7800;
    \\u4_u0_buf0_orig_m3_reg[7]  <= n7805;
    \\u4_u0_buf0_orig_m3_reg[8]  <= n7810;
    \\u1_u3_tx_data_to_cnt_reg[6]  <= n7815;
    \\u1_u3_tx_data_to_cnt_reg[2]  <= n7820;
    \\u1_u3_tx_data_to_cnt_reg[1]  <= n7825;
    \\u1_u3_tx_data_to_cnt_reg[0]  <= n7830;
    \\u4_u3_buf0_orig_m3_reg[9]  <= n7835;
    \\u4_u1_buf0_orig_m3_reg[9]  <= n7840;
    \\u4_u3_buf0_orig_m3_reg[10]  <= n7845;
    u1_u3_buf0_na_reg <= n7850;
    u1_u3_buf1_na_reg <= n7855;
    \\u1_u3_tx_data_to_cnt_reg[3]  <= n7860;
    u4_u3_int_re_reg <= n7865;
    \\u4_u0_buf0_orig_m3_reg[6]  <= n7870;
    \\u4_u2_buf0_orig_m3_reg[6]  <= n7875;
    \\u1_u3_tx_data_to_cnt_reg[7]  <= n7880;
    u4_u0_dma_req_in_hold_reg <= n7885;
    \\u1_u3_tx_data_to_cnt_reg[5]  <= n7890;
    u0_u0_mode_hs_reg <= n7895;
    u4_u3_ep_match_r_reg <= n7900;
    \\u1_u3_idin_reg[22]  <= n7905;
    \\u4_u1_buf0_orig_m3_reg[3]  <= n7910;
    \\u4_u3_buf0_orig_m3_reg[7]  <= n7915;
    \\u4_u2_buf0_orig_m3_reg[7]  <= n7920;
    \\u4_u3_buf0_orig_m3_reg[8]  <= n7925;
    \\u4_u2_buf0_orig_m3_reg[8]  <= n7930;
    \\u4_int_srca_reg[1]  <= n7935;
    \\u4_u1_buf0_orig_m3_reg[4]  <= n7940;
    \\u4_u1_buf0_orig_m3_reg[2]  <= n7945;
    \\u4_u1_buf0_orig_m3_reg[6]  <= n7950;
    u4_u2_dma_req_in_hold_reg <= n7955;
    u4_u1_dma_req_in_hold_reg <= n7960;
    u1_u3_out_token_reg <= n7965;
    u1_u3_setup_token_reg <= n7970;
    u0_u0_ls_idle_r_reg <= n7975;
    u1_u0_rx_active_r_reg <= n7980;
    \\u4_u0_buf0_orig_m3_reg[3]  <= n7985;
    \\u4_u3_dma_out_left_reg[4]  <= n7990;
    \\u4_u0_dma_out_left_reg[4]  <= n7995;
    \\u4_u1_dma_out_left_reg[4]  <= n8000;
    \\u4_u2_dma_out_left_reg[4]  <= n8005;
    \\u1_u3_rx_ack_to_cnt_reg[4]  <= n8010;
    \\u4_int_srca_reg[0]  <= n8015;
    \\u4_int_srca_reg[3]  <= n8020;
    \\u4_int_srca_reg[2]  <= n8025;
    \\u1_u3_rx_ack_to_cnt_reg[3]  <= n8030;
    \\u4_u0_buf0_orig_m3_reg[4]  <= n8035;
    \\u1_u3_rx_ack_to_cnt_reg[2]  <= n8040;
    \\u4_u0_buf0_orig_m3_reg[2]  <= n8045;
    u1_u3_buf1_not_aloc_reg <= n8050;
    u1_u3_buf0_not_aloc_reg <= n8055;
    \\u4_u0_buf0_orig_m3_reg[5]  <= n8060;
    \\u4_u1_buf0_orig_m3_reg[5]  <= n8065;
    \\u4_u3_buf0_orig_m3_reg[6]  <= n8070;
    \\u4_u2_buf0_orig_m3_reg[5]  <= n8075;
    \\u1_u3_rx_ack_to_cnt_reg[6]  <= n8080;
    \\u1_u3_rx_ack_to_cnt_reg[0]  <= n8085;
    \\u1_u3_rx_ack_to_cnt_reg[1]  <= n8090;
    \\u1_u3_rx_ack_to_cnt_reg[7]  <= n8095;
    u4_u3_dma_req_in_hold_reg <= n8100;
    \\u1_u3_rx_ack_to_cnt_reg[5]  <= n8105;
    \\u0_u0_idle_cnt1_next_reg[7]  <= n8110;
    u4_pid_cs_err_r_reg <= n8115;
    \\u4_u3_buf0_orig_m3_reg[3]  <= n8120;
    \\u4_u2_buf0_orig_m3_reg[3]  <= n8125;
    u1_u3_buf0_rl_reg <= n8130;
    \\u0_u0_idle_cnt1_next_reg[6]  <= n8135;
    \\u4_u3_dma_out_left_reg[3]  <= n8140;
    \\u4_u0_dma_out_left_reg[3]  <= n8145;
    \\u4_u1_dma_out_left_reg[3]  <= n8150;
    \\u4_u2_dma_out_left_reg[3]  <= n8155;
    \\u0_u0_idle_cnt1_next_reg[4]  <= n8160;
    \\u4_u3_buf0_orig_m3_reg[4]  <= n8165;
    u0_u0_me_ps2_0_5_ms_reg <= n8170;
    \\u4_u2_buf0_orig_m3_reg[4]  <= n8175;
    \\u4_u2_buf0_orig_m3_reg[2]  <= n8180;
    \\u4_u3_buf0_orig_m3_reg[5]  <= n8185;
    u4_u2_dma_req_out_hold_reg <= n8190;
    u4_u3_dma_req_out_hold_reg <= n8195;
    u4_u0_dma_req_out_hold_reg <= n8200;
    u4_u1_dma_req_out_hold_reg <= n8205;
    u1_u1_send_data_r2_reg <= n8210;
    u4_usb_reset_r_reg <= n8215;
    u0_u0_idle_cnt1_clr_reg <= n8220;
    \\u4_u3_buf0_orig_m3_reg[2]  <= n8225;
    \\u0_u0_idle_cnt1_next_reg[5]  <= n8230;
    u1_u2_sizd_is_zero_reg <= n8235;
    u4_rx_err_r_reg <= n8240;
    u0_drive_k_r_reg <= n8245;
    \\u0_u0_idle_cnt1_next_reg[3]  <= n8250;
    u4_u2_dma_ack_wr1_reg <= n8255;
    \\u4_u1_dma_out_left_reg[2]  <= n8260;
    \\u4_u0_dma_out_left_reg[2]  <= n8265;
    \\u4_u3_dma_out_left_reg[2]  <= n8270;
    \\u4_u2_dma_out_left_reg[2]  <= n8275;
    u4_u1_dma_ack_wr1_reg <= n8280;
    \\u4_u2_dma_out_left_reg[1]  <= n8285;
    \\u4_u1_dma_out_left_reg[1]  <= n8290;
    \\u4_u0_dma_out_left_reg[1]  <= n8295;
    \\u4_u3_dma_out_left_reg[1]  <= n8300;
    u4_u0_dma_ack_wr1_reg <= n8305;
    u4_u3_dma_ack_wr1_reg <= n8310;
    \\u1_u2_rd_buf1_reg[19]  <= n8315;
    \\u1_u2_rd_buf1_reg[1]  <= n8320;
    \\u4_u0_buf0_orig_m3_reg[1]  <= n8325;
    \\u4_u3_buf0_orig_m3_reg[1]  <= n8330;
    \\u4_u2_buf0_orig_m3_reg[1]  <= n8335;
    u1_u3_pid_OUT_r_reg <= n8340;
    u4_u2_set_r_reg <= n8345;
    u1_u3_pid_IN_r_reg <= n8350;
    u4_u0_set_r_reg <= n8355;
    u4_u1_set_r_reg <= n8360;
    \\u1_u2_rd_buf1_reg[31]  <= n8365;
    \\u1_u2_rd_buf1_reg[30]  <= n8370;
    \\u1_u2_rd_buf1_reg[7]  <= n8375;
    \\u1_u2_rd_buf1_reg[24]  <= n8380;
    \\u1_u2_rd_buf1_reg[21]  <= n8385;
    u0_u0_usb_reset_reg <= n8390;
    u1_u2_dtmp_sel_r_reg <= n8395;
    u1_u3_pid_SETUP_r_reg <= n8400;
    u1_u3_rx_ack_to_clr_reg <= n8405;
    u1_u3_pid_PING_r_reg <= n8410;
    u4_u2_r2_reg <= n8415;
    \\u1_u2_rd_buf1_reg[26]  <= n8420;
    \\u1_u2_rd_buf1_reg[27]  <= n8425;
    \\u1_u2_rd_buf1_reg[3]  <= n8430;
    \\u1_u2_rd_buf1_reg[0]  <= n8435;
    \\u1_u2_rd_buf1_reg[12]  <= n8440;
    \\u1_u2_rd_buf1_reg[2]  <= n8445;
    \\u1_u2_rd_buf1_reg[8]  <= n8450;
    \\u1_u2_rd_buf1_reg[18]  <= n8455;
    \\u1_u2_rd_buf1_reg[28]  <= n8460;
    \\u1_u2_rd_buf1_reg[14]  <= n8465;
    u4_u3_set_r_reg <= n8470;
    \\u1_u2_rd_buf1_reg[6]  <= n8475;
    \\u1_u2_rd_buf1_reg[5]  <= n8480;
    \\u1_u2_rd_buf1_reg[9]  <= n8485;
    \\u1_u2_rd_buf1_reg[20]  <= n8490;
    \\u1_u2_rd_buf1_reg[22]  <= n8495;
    \\u1_u2_rd_buf1_reg[15]  <= n8500;
    \\u1_u2_rd_buf1_reg[23]  <= n8505;
    \\u1_u2_rd_buf1_reg[25]  <= n8510;
    \\u1_u2_rd_buf1_reg[17]  <= n8515;
    u4_u3_r2_reg <= n8520;
    \\u1_u2_rd_buf1_reg[16]  <= n8525;
    \\u1_u2_rd_buf1_reg[4]  <= n8530;
    u4_u0_r2_reg <= n8535;
    u4_u1_r2_reg <= n8540;
    \\u1_u2_rd_buf1_reg[29]  <= n8545;
    \\u1_u2_rd_buf1_reg[10]  <= n8550;
    u4_u1_intb_reg <= n8555;
    u4_u2_intb_reg <= n8560;
    u4_u0_intb_reg <= n8565;
    \\u1_u2_rd_buf1_reg[11]  <= n8570;
    \\u1_u2_rd_buf1_reg[13]  <= n8575;
    u4_u0_inta_reg <= n8580;
    u4_u1_inta_reg <= n8585;
    u4_u2_inta_reg <= n8590;
    u4_u3_inta_reg <= n8595;
    u4_u3_intb_reg <= n8600;
    u0_u0_me_ps_2_5_us_reg <= n8605;
    \\u4_u3_dma_out_left_reg[0]  <= n8610;
    \\u4_u2_dma_out_left_reg[0]  <= n8615;
    \\u4_u0_dma_out_left_reg[0]  <= n8620;
    u1_u1_send_data_r_reg <= n8625;
    u0_rx_active_reg <= n8630;
    u0_rx_err_reg <= n8635;
    u0_rx_valid_reg <= n8640;
    u0_u0_ls_se0_r_reg <= n8645;
    \\u4_u1_dma_out_left_reg[0]  <= n8650;
    \\u0_u0_idle_cnt1_next_reg[2]  <= n8655;
    \\u1_u2_rd_buf0_reg[2]  <= n8660;
    \\u1_u2_rd_buf0_reg[31]  <= n8665;
    \\u1_u2_rd_buf0_reg[28]  <= n8670;
    \\u1_u2_rd_buf0_reg[6]  <= n8675;
    \\u1_u2_rd_buf0_reg[23]  <= n8680;
    \\u4_u1_buf0_orig_m3_reg[1]  <= n8685;
    \\u1_u2_rd_buf0_reg[19]  <= n8690;
    \\u1_u2_rd_buf0_reg[24]  <= n8695;
    \\u1_u2_rd_buf0_reg[18]  <= n8700;
    \\u1_u2_rd_buf0_reg[10]  <= n8705;
    \\u1_u2_rd_buf0_reg[4]  <= n8710;
    \\u1_u2_rd_buf0_reg[30]  <= n8715;
    \\u1_u2_rd_buf0_reg[27]  <= n8720;
    \\u1_u2_rd_buf0_reg[3]  <= n8725;
    \\u1_u2_rd_buf0_reg[5]  <= n8730;
    \\u1_u2_rd_buf0_reg[8]  <= n8735;
    \\u1_u2_rd_buf0_reg[26]  <= n8740;
    \\u1_u2_rd_buf0_reg[14]  <= n8745;
    \\u1_u2_rd_buf0_reg[0]  <= n8750;
    \\u1_u2_rd_buf0_reg[1]  <= n8755;
    \\u1_u2_rd_buf0_reg[29]  <= n8760;
    \\u1_u2_rd_buf0_reg[9]  <= n8765;
    \\u1_u2_rd_buf0_reg[21]  <= n8770;
    \\u1_u2_rd_buf0_reg[20]  <= n8775;
    \\u1_u2_rd_buf0_reg[16]  <= n8780;
    \\u1_u2_rd_buf0_reg[17]  <= n8785;
    \\u1_u2_rd_buf0_reg[7]  <= n8790;
    \\u1_u2_rd_buf0_reg[22]  <= n8795;
    \\u1_u2_rd_buf0_reg[13]  <= n8800;
    \\u1_u2_rd_buf0_reg[25]  <= n8805;
    \\u1_u2_rd_buf0_reg[12]  <= n8810;
    \\u1_u2_rd_buf0_reg[15]  <= n8815;
    \\u1_u2_rd_buf0_reg[11]  <= n8820;
    u0_u0_ps_cnt_clr_reg <= n8825;
    \\u1_u3_idin_reg[31]  <= n8830;
    u0_u0_drive_k_reg <= n8835;
    u0_u0_ls_j_r_reg <= n8840;
    u1_u2_mwe_reg <= n8845;
    u0_u0_chirp_cnt_is_6_reg <= n8850;
    u1_hms_clk_reg <= n8855;
    \\u1_u3_idin_reg[28]  <= n8860;
    \\u0_u0_idle_cnt1_next_reg[1]  <= n8865;
    u0_u0_ls_k_r_reg <= n8870;
    u4_suspend_r1_reg <= n8875;
    u4_attach_r1_reg <= n8880;
    \\u0_u0_state_reg[0]  <= n8885;
    \\u4_u1_buf0_orig_m3_reg[0]  <= n8890;
    u4_u1_r5_reg <= n8895;
    u4_suspend_r_reg <= n8900;
    \\u4_utmi_vend_stat_r_reg[5]  <= n8905;
    \\u4_utmi_vend_stat_r_reg[2]  <= n8910;
    u0_u0_resume_req_s_reg <= n8915;
    \\u4_utmi_vend_stat_r_reg[1]  <= n8920;
    \\u4_utmi_vend_stat_r_reg[7]  <= n8925;
    \\u4_utmi_vend_stat_r_reg[4]  <= n8930;
    \\u4_utmi_vend_stat_r_reg[0]  <= n8935;
    u5_wb_req_s1_reg <= n8940;
    u4_u1_dma_ack_clr1_reg <= n8945;
    u4_u0_r5_reg <= n8950;
    u4_u0_dma_ack_clr1_reg <= n8955;
    u0_tx_ready_reg <= n8960;
    \\u4_utmi_vend_stat_r_reg[6]  <= n8965;
    u4_u2_dma_ack_clr1_reg <= n8970;
    u1_u3_uc_dpd_set_reg <= n8975;
    u4_u3_dma_ack_clr1_reg <= n8980;
    u4_u2_r5_reg <= n8985;
    u1_u3_uc_bsel_set_reg <= n8990;
    u4_u3_r5_reg <= n8995;
    \\u4_utmi_vend_stat_r_reg[3]  <= n9000;
    susp_o_reg <= n9005;
    \\u4_u0_buf0_orig_m3_reg[0]  <= n9010;
    \\u4_u2_buf0_orig_m3_reg[0]  <= n9015;
    \\u4_u3_buf0_orig_m3_reg[0]  <= n9020;
    \\u0_u0_idle_cnt1_next_reg[0]  <= n9025;
    \\u4_utmi_vend_ctrl_reg[3]  <= n9030;
    u4_utmi_vend_wr_reg <= n9035;
    \\u4_utmi_vend_ctrl_reg[0]  <= n9040;
    \\u1_u2_rx_data_st_r_reg[4]  <= n9045;
    \\u4_utmi_vend_ctrl_reg[2]  <= n9050;
    \\u1_u2_rx_data_st_r_reg[7]  <= n9055;
    \\u1_u2_rx_data_st_r_reg[0]  <= n9060;
    \\u1_u2_rx_data_st_r_reg[2]  <= n9065;
    \\u1_u2_rx_data_st_r_reg[3]  <= n9070;
    \\u4_utmi_vend_ctrl_reg[1]  <= n9075;
    \\u1_u2_rx_data_st_r_reg[1]  <= n9080;
    \\u1_u2_rx_data_st_r_reg[5]  <= n9085;
    \\u1_u2_rx_data_st_r_reg[6]  <= n9090;
    \\VStatus_r_reg[5]  <= n9095;
    \\VStatus_r_reg[1]  <= n9100;
    \\VStatus_r_reg[3]  <= n9105;
    \\u0_rx_data_reg[2]  <= n9110;
    \\VStatus_r_reg[2]  <= n9115;
    u0_u0_resume_req_s1_reg <= n9120;
    \\u0_rx_data_reg[7]  <= n9125;
    u4_attach_r_reg <= n9130;
    \\u0_rx_data_reg[3]  <= n9135;
    u4_u3_r4_reg <= n9140;
    u1_u3_out_to_small_reg <= n9145;
    u4_u1_r4_reg <= n9150;
    \\LineState_r_reg[0]  <= n9155;
    \\VStatus_r_reg[4]  <= n9160;
    \\u0_rx_data_reg[0]  <= n9165;
    u4_u0_r4_reg <= n9170;
    \\u0_rx_data_reg[5]  <= n9175;
    \\VStatus_r_reg[7]  <= n9180;
    \\u0_u0_line_state_r_reg[1]  <= n9185;
    \\u0_rx_data_reg[6]  <= n9190;
    \\u0_u0_line_state_r_reg[0]  <= n9195;
    \\u0_rx_data_reg[4]  <= n9200;
    \\u0_rx_data_reg[1]  <= n9205;
    \\LineState_r_reg[1]  <= n9210;
    u4_u2_r4_reg <= n9215;
    \\VStatus_r_reg[6]  <= n9220;
    \\VStatus_r_reg[0]  <= n9225;
  end
endmodule


