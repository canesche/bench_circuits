module top ( clock, 
    p_30, p_20, p_10, p_12, p_23, p_11, p_24, p_33, pclk, p_14, p_21, p_32,
    p_13, p_22, p_31, p_16, p_27, p_15, p_28, p_9, p_18, p_25, p_8, p_17,
    p_26, p_7, p_6, p_19, p_5, p_29, p_4, p_3, p_2, p_1,
    p_140, p_151, p_130, p_152, p_153, p_133, p_144, p_134, p_143, p_124,
    p_131, p_142, p_132, p_141, p_150, p_126, p_137, p_148, p_125, p_138,
    p_147, p_128, p_135, p_146, p_127, p_136, p_145, p_129, p_139, p_149  );
  input  clock;
  input  p_30, p_20, p_10, p_12, p_23, p_11, p_24, p_33, pclk, p_14,
    p_21, p_32, p_13, p_22, p_31, p_16, p_27, p_15, p_28, p_9, p_18, p_25,
    p_8, p_17, p_26, p_7, p_6, p_19, p_5, p_29, p_4, p_3, p_2, p_1;
  output p_140, p_151, p_130, p_152, p_153, p_133, p_144, p_134, p_143, p_124,
    p_131, p_142, p_132, p_141, p_150, p_126, p_137, p_148, p_125, p_138,
    p_147, p_128, p_135, p_146, p_127, p_136, p_145, p_129, p_139, p_149;
  reg n_43, n_39, n_40, n_41, n_42, n_35, n_36, n_37, n_38, n_84, n_95,
    n_106, n_117, n_85, n_94, n_107, n_116, n_86, n_97, n_104, n_115, n_34,
    n_87, n_96, n_105, n_114, n_44, n_55, n_66, n_77, n_45, n_54, n_67,
    n_76, n_46, n_57, n_64, n_75, n_47, n_56, n_65, n_74, n_48, n_59, n_70,
    n_81, n_92, n_103, n_49, n_58, n_71, n_80, n_93, n_102, n_50, n_61,
    n_68, n_79, n_112, n_123, n_51, n_60, n_69, n_78, n_113, n_122, n_52,
    n_63, n_88, n_99, n_110, n_121, n_53, n_62, n_89, n_98, n_111, n_120,
    n_72, n_83, n_90, n_101, n_108, n_119, n_73, n_82, n_91, n_100, n_109,
    n_118;
  wire new_n335_1_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_1_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_1_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_1_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_1_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_1_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_1_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_1_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_1_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_1_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_1_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_1_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_1_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_1_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_1_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_1_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_1_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_1_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_1_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_1_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_1_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_1_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_1_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_1_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_1_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_1_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_1_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_1_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_1_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_1_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_1_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_1_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_1_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_1_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_1_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_1_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_1_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_1_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_1_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_1_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_1_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_1_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_1_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_1_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_1_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_1_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_1_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_1_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_1_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_,
    new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1224_, new_n1225_,
    new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_,
    new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1320_,
    new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_,
    new_n1334_, new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_,
    new_n1340_, new_n1341_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1479_, new_n1480_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_,
    new_n1493_, new_n1494_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_, new_n1518_,
    new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_, new_n1524_,
    new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1530_, new_n1531_,
    new_n1532_, new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_,
    new_n1538_, new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_,
    new_n1544_, new_n1545_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1581_, new_n1583_,
    new_n1585_, new_n1587_, new_n1589_, new_n1591_, new_n1593_, new_n1595_,
    new_n1597_, new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_,
    new_n1605_, new_n1606_, new_n1608_, new_n1609_, new_n1611_, new_n1612_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1620_,
    new_n1621_, new_n1623_, new_n1624_, new_n1626_, new_n1627_, new_n1629_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1635_, new_n1636_,
    new_n1638_, new_n1639_, new_n1641_, new_n1642_, new_n1644_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1652_, new_n1653_,
    new_n1655_, new_n1656_, new_n1658_, new_n1659_, new_n1661_, new_n1663_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1677_, new_n1679_,
    new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1693_, new_n1695_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1709_, new_n1711_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1719_,
    new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1725_, new_n1727_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1735_,
    new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1747_, new_n1748_, new_n1750_,
    new_n1752_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1772_, new_n1773_,
    new_n1775_, new_n1777_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_,
    new_n1791_, new_n1792_, new_n1794_, new_n1795_, new_n1797_, new_n1799_,
    new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1813_, new_n1814_,
    new_n1816_, new_n1817_, new_n1819_, new_n1821_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1829_, new_n1830_, new_n1832_,
    new_n1833_, new_n1835_, new_n1836_, new_n1838_, new_n1840_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1848_, new_n1849_,
    new_n1851_, new_n1852_, new_n1854_, new_n1855_, new_n1857_, new_n1858_,
    new_n1859_, new_n1860_, new_n1861_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1869_, new_n1870_, new_n1871_, new_n1872_,
    new_n1873_, new_n1875_, new_n1876_, new_n1878_, new_n1879_, new_n1881_,
    new_n1882_, new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1896_,
    new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1902_, new_n1903_,
    new_n1905_, new_n1906_, new_n1908_, new_n1909_, n130, n135, n140, n145,
    n150, n155, n160, n165, n170, n175, n180, n185, n190, n195, n200, n205,
    n210, n215, n220, n225, n230, n235, n240, n245, n250, n255, n260, n265,
    n270, n275, n280, n285, n290, n295, n300, n305, n310, n315, n320, n325,
    n330, n335, n340, n345, n350, n355, n360, n365, n370, n375, n380, n385,
    n390, n395, n400, n405, n410, n415, n420, n425, n430, n435, n440, n445,
    n450, n455, n460, n465, n470, n475, n480, n485, n490, n495, n500, n505,
    n510, n515, n520, n525, n530, n535, n540, n545, n550, n555, n560, n565,
    n570, n575;
  assign new_n335_1_ = ~p_3 & p_2;
  assign new_n336_ = ~p_1 & new_n335_1_;
  assign new_n337_ = ~p_4 & n_94;
  assign new_n338_ = p_4 & ~n_94;
  assign new_n339_ = ~new_n337_ & ~new_n338_;
  assign new_n340_1_ = p_4 & ~new_n339_;
  assign new_n341_ = ~p_5 & n_95;
  assign new_n342_ = p_5 & ~n_95;
  assign new_n343_ = ~new_n341_ & ~new_n342_;
  assign new_n344_ = new_n340_1_ & new_n343_;
  assign new_n345_1_ = p_5 & ~new_n343_;
  assign new_n346_ = ~new_n344_ & ~new_n345_1_;
  assign new_n347_ = ~p_6 & n_96;
  assign new_n348_ = p_6 & ~n_96;
  assign new_n349_ = ~new_n347_ & ~new_n348_;
  assign new_n350_1_ = ~new_n346_ & new_n349_;
  assign new_n351_ = p_6 & ~new_n349_;
  assign new_n352_ = ~new_n350_1_ & ~new_n351_;
  assign new_n353_ = ~p_7 & n_97;
  assign new_n354_ = p_7 & ~n_97;
  assign new_n355_1_ = ~new_n353_ & ~new_n354_;
  assign new_n356_ = ~new_n352_ & new_n355_1_;
  assign new_n357_ = p_7 & ~new_n355_1_;
  assign new_n358_ = ~new_n356_ & ~new_n357_;
  assign new_n359_ = ~p_8 & n_98;
  assign new_n360_1_ = p_8 & ~n_98;
  assign new_n361_ = ~new_n359_ & ~new_n360_1_;
  assign new_n362_ = ~new_n358_ & new_n361_;
  assign new_n363_ = p_8 & ~new_n361_;
  assign new_n364_ = ~new_n362_ & ~new_n363_;
  assign new_n365_1_ = ~p_9 & n_99;
  assign new_n366_ = p_9 & ~n_99;
  assign new_n367_ = ~new_n365_1_ & ~new_n366_;
  assign new_n368_ = ~new_n364_ & new_n367_;
  assign new_n369_ = p_9 & ~new_n367_;
  assign new_n370_1_ = ~new_n368_ & ~new_n369_;
  assign new_n371_ = ~p_10 & n_100;
  assign new_n372_ = p_10 & ~n_100;
  assign new_n373_ = ~new_n371_ & ~new_n372_;
  assign new_n374_ = ~new_n370_1_ & new_n373_;
  assign new_n375_1_ = p_10 & ~new_n373_;
  assign new_n376_ = ~new_n374_ & ~new_n375_1_;
  assign new_n377_ = ~p_11 & n_101;
  assign new_n378_ = p_11 & ~n_101;
  assign new_n379_ = ~new_n377_ & ~new_n378_;
  assign new_n380_1_ = ~new_n376_ & new_n379_;
  assign new_n381_ = p_11 & ~new_n379_;
  assign new_n382_ = ~new_n380_1_ & ~new_n381_;
  assign new_n383_ = ~p_12 & n_102;
  assign new_n384_ = p_12 & ~n_102;
  assign new_n385_1_ = ~new_n383_ & ~new_n384_;
  assign new_n386_ = ~new_n382_ & new_n385_1_;
  assign new_n387_ = p_12 & ~new_n385_1_;
  assign new_n388_ = ~new_n386_ & ~new_n387_;
  assign new_n389_ = ~p_13 & n_103;
  assign new_n390_1_ = p_13 & ~n_103;
  assign new_n391_ = ~new_n389_ & ~new_n390_1_;
  assign new_n392_ = ~new_n388_ & new_n391_;
  assign new_n393_ = p_13 & ~new_n391_;
  assign new_n394_ = ~new_n392_ & ~new_n393_;
  assign new_n395_1_ = ~p_14 & n_104;
  assign new_n396_ = p_14 & ~n_104;
  assign new_n397_ = ~new_n395_1_ & ~new_n396_;
  assign new_n398_ = ~new_n394_ & new_n397_;
  assign new_n399_ = p_14 & ~new_n397_;
  assign new_n400_1_ = ~new_n398_ & ~new_n399_;
  assign new_n401_ = ~p_15 & n_105;
  assign new_n402_ = p_15 & ~n_105;
  assign new_n403_ = ~new_n401_ & ~new_n402_;
  assign new_n404_ = ~new_n400_1_ & new_n403_;
  assign new_n405_1_ = p_15 & ~new_n403_;
  assign new_n406_ = ~new_n404_ & ~new_n405_1_;
  assign new_n407_ = ~p_16 & n_106;
  assign new_n408_ = p_16 & ~n_106;
  assign new_n409_ = ~new_n407_ & ~new_n408_;
  assign new_n410_1_ = ~new_n406_ & new_n409_;
  assign new_n411_ = p_16 & ~new_n409_;
  assign new_n412_ = ~new_n410_1_ & ~new_n411_;
  assign new_n413_ = ~p_17 & n_107;
  assign new_n414_ = p_17 & ~n_107;
  assign new_n415_1_ = ~new_n413_ & ~new_n414_;
  assign new_n416_ = ~new_n412_ & new_n415_1_;
  assign new_n417_ = p_17 & ~new_n415_1_;
  assign new_n418_ = ~new_n416_ & ~new_n417_;
  assign new_n419_ = ~p_18 & n_108;
  assign new_n420_1_ = p_18 & ~n_108;
  assign new_n421_ = ~new_n419_ & ~new_n420_1_;
  assign new_n422_ = ~new_n418_ & new_n421_;
  assign new_n423_ = p_18 & ~new_n421_;
  assign new_n424_ = ~new_n422_ & ~new_n423_;
  assign new_n425_1_ = ~p_19 & n_109;
  assign new_n426_ = p_19 & ~n_109;
  assign new_n427_ = ~new_n425_1_ & ~new_n426_;
  assign new_n428_ = ~new_n424_ & new_n427_;
  assign new_n429_ = p_19 & ~new_n427_;
  assign new_n430_1_ = ~new_n428_ & ~new_n429_;
  assign new_n431_ = ~p_20 & n_110;
  assign new_n432_ = p_20 & ~n_110;
  assign new_n433_ = ~new_n431_ & ~new_n432_;
  assign new_n434_ = ~new_n430_1_ & new_n433_;
  assign new_n435_1_ = p_20 & ~new_n433_;
  assign new_n436_ = ~new_n434_ & ~new_n435_1_;
  assign new_n437_ = ~p_21 & n_111;
  assign new_n438_ = p_21 & ~n_111;
  assign new_n439_ = ~new_n437_ & ~new_n438_;
  assign new_n440_1_ = ~new_n436_ & new_n439_;
  assign new_n441_ = p_21 & ~new_n439_;
  assign new_n442_ = ~new_n440_1_ & ~new_n441_;
  assign new_n443_ = ~p_22 & n_112;
  assign new_n444_ = p_22 & ~n_112;
  assign new_n445_1_ = ~new_n443_ & ~new_n444_;
  assign new_n446_ = ~new_n442_ & new_n445_1_;
  assign new_n447_ = p_22 & ~new_n445_1_;
  assign new_n448_ = ~new_n446_ & ~new_n447_;
  assign new_n449_ = ~p_23 & n_113;
  assign new_n450_1_ = p_23 & ~n_113;
  assign new_n451_ = ~new_n449_ & ~new_n450_1_;
  assign new_n452_ = ~new_n448_ & new_n451_;
  assign new_n453_ = p_23 & ~new_n451_;
  assign new_n454_ = ~new_n452_ & ~new_n453_;
  assign new_n455_1_ = ~p_24 & n_114;
  assign new_n456_ = p_24 & ~n_114;
  assign new_n457_ = ~new_n455_1_ & ~new_n456_;
  assign new_n458_ = ~new_n454_ & new_n457_;
  assign new_n459_ = p_24 & ~new_n457_;
  assign new_n460_1_ = ~new_n458_ & ~new_n459_;
  assign new_n461_ = ~p_25 & n_115;
  assign new_n462_ = p_25 & ~n_115;
  assign new_n463_ = ~new_n461_ & ~new_n462_;
  assign new_n464_ = ~new_n460_1_ & new_n463_;
  assign new_n465_1_ = p_25 & ~new_n463_;
  assign new_n466_ = ~new_n464_ & ~new_n465_1_;
  assign new_n467_ = ~p_26 & n_116;
  assign new_n468_ = p_26 & ~n_116;
  assign new_n469_ = ~new_n467_ & ~new_n468_;
  assign new_n470_1_ = ~new_n466_ & new_n469_;
  assign new_n471_ = p_26 & ~new_n469_;
  assign new_n472_ = ~new_n470_1_ & ~new_n471_;
  assign new_n473_ = ~p_27 & n_117;
  assign new_n474_ = p_27 & ~n_117;
  assign new_n475_1_ = ~new_n473_ & ~new_n474_;
  assign new_n476_ = ~new_n472_ & new_n475_1_;
  assign new_n477_ = p_27 & ~new_n475_1_;
  assign new_n478_ = ~new_n476_ & ~new_n477_;
  assign new_n479_ = ~p_28 & n_118;
  assign new_n480_1_ = p_28 & ~n_118;
  assign new_n481_ = ~new_n479_ & ~new_n480_1_;
  assign new_n482_ = ~new_n478_ & new_n481_;
  assign new_n483_ = p_28 & ~new_n481_;
  assign new_n484_ = ~new_n482_ & ~new_n483_;
  assign new_n485_1_ = ~p_29 & n_119;
  assign new_n486_ = p_29 & ~n_119;
  assign new_n487_ = ~new_n485_1_ & ~new_n486_;
  assign new_n488_ = ~new_n484_ & new_n487_;
  assign new_n489_ = p_29 & ~new_n487_;
  assign new_n490_1_ = ~new_n488_ & ~new_n489_;
  assign new_n491_ = ~p_30 & n_120;
  assign new_n492_ = p_30 & ~n_120;
  assign new_n493_ = ~new_n491_ & ~new_n492_;
  assign new_n494_ = ~new_n490_1_ & new_n493_;
  assign new_n495_1_ = p_30 & ~new_n493_;
  assign new_n496_ = ~new_n494_ & ~new_n495_1_;
  assign new_n497_ = ~p_31 & n_121;
  assign new_n498_ = p_31 & ~n_121;
  assign new_n499_ = ~new_n497_ & ~new_n498_;
  assign new_n500_1_ = ~new_n496_ & new_n499_;
  assign new_n501_ = p_31 & ~new_n499_;
  assign new_n502_ = ~new_n500_1_ & ~new_n501_;
  assign new_n503_ = ~p_32 & n_122;
  assign new_n504_ = p_32 & ~n_122;
  assign new_n505_1_ = ~new_n503_ & ~new_n504_;
  assign new_n506_ = ~new_n502_ & new_n505_1_;
  assign new_n507_ = p_32 & ~new_n505_1_;
  assign new_n508_ = ~new_n506_ & ~new_n507_;
  assign new_n509_ = ~p_33 & n_123;
  assign new_n510_1_ = p_33 & ~n_123;
  assign new_n511_ = ~new_n509_ & ~new_n510_1_;
  assign new_n512_ = ~new_n508_ & new_n511_;
  assign new_n513_ = p_33 & ~new_n511_;
  assign new_n514_ = ~new_n512_ & ~new_n513_;
  assign new_n515_1_ = new_n336_ & ~new_n514_;
  assign new_n516_ = n_111 & ~new_n515_1_;
  assign new_n517_ = p_21 & new_n515_1_;
  assign new_n518_ = ~new_n516_ & ~new_n517_;
  assign new_n519_ = new_n336_ & ~new_n518_;
  assign new_n520_1_ = ~p_4 & n_64;
  assign new_n521_ = p_4 & ~n_64;
  assign new_n522_ = ~new_n520_1_ & ~new_n521_;
  assign new_n523_ = p_4 & ~new_n522_;
  assign new_n524_ = ~p_5 & n_65;
  assign new_n525_1_ = p_5 & ~n_65;
  assign new_n526_ = ~new_n524_ & ~new_n525_1_;
  assign new_n527_ = new_n523_ & new_n526_;
  assign new_n528_ = p_5 & ~new_n526_;
  assign new_n529_ = ~new_n527_ & ~new_n528_;
  assign new_n530_1_ = ~p_6 & n_66;
  assign new_n531_ = p_6 & ~n_66;
  assign new_n532_ = ~new_n530_1_ & ~new_n531_;
  assign new_n533_ = ~new_n529_ & new_n532_;
  assign new_n534_ = p_6 & ~new_n532_;
  assign new_n535_1_ = ~new_n533_ & ~new_n534_;
  assign new_n536_ = ~p_7 & n_67;
  assign new_n537_ = p_7 & ~n_67;
  assign new_n538_ = ~new_n536_ & ~new_n537_;
  assign new_n539_ = ~new_n535_1_ & new_n538_;
  assign new_n540_1_ = p_7 & ~new_n538_;
  assign new_n541_ = ~new_n539_ & ~new_n540_1_;
  assign new_n542_ = ~p_8 & n_68;
  assign new_n543_ = p_8 & ~n_68;
  assign new_n544_ = ~new_n542_ & ~new_n543_;
  assign new_n545_1_ = ~new_n541_ & new_n544_;
  assign new_n546_ = p_8 & ~new_n544_;
  assign new_n547_ = ~new_n545_1_ & ~new_n546_;
  assign new_n548_ = ~p_9 & n_69;
  assign new_n549_ = p_9 & ~n_69;
  assign new_n550_1_ = ~new_n548_ & ~new_n549_;
  assign new_n551_ = ~new_n547_ & new_n550_1_;
  assign new_n552_ = p_9 & ~new_n550_1_;
  assign new_n553_ = ~new_n551_ & ~new_n552_;
  assign new_n554_ = ~p_10 & n_70;
  assign new_n555_1_ = p_10 & ~n_70;
  assign new_n556_ = ~new_n554_ & ~new_n555_1_;
  assign new_n557_ = ~new_n553_ & new_n556_;
  assign new_n558_ = p_10 & ~new_n556_;
  assign new_n559_ = ~new_n557_ & ~new_n558_;
  assign new_n560_1_ = ~p_11 & n_71;
  assign new_n561_ = p_11 & ~n_71;
  assign new_n562_ = ~new_n560_1_ & ~new_n561_;
  assign new_n563_ = ~new_n559_ & new_n562_;
  assign new_n564_ = p_11 & ~new_n562_;
  assign new_n565_1_ = ~new_n563_ & ~new_n564_;
  assign new_n566_ = ~p_12 & n_72;
  assign new_n567_ = p_12 & ~n_72;
  assign new_n568_ = ~new_n566_ & ~new_n567_;
  assign new_n569_ = ~new_n565_1_ & new_n568_;
  assign new_n570_1_ = p_12 & ~new_n568_;
  assign new_n571_ = ~new_n569_ & ~new_n570_1_;
  assign new_n572_ = ~p_13 & n_73;
  assign new_n573_ = p_13 & ~n_73;
  assign new_n574_ = ~new_n572_ & ~new_n573_;
  assign new_n575_1_ = ~new_n571_ & new_n574_;
  assign new_n576_ = p_13 & ~new_n574_;
  assign new_n577_ = ~new_n575_1_ & ~new_n576_;
  assign new_n578_ = ~p_14 & n_74;
  assign new_n579_ = p_14 & ~n_74;
  assign new_n580_ = ~new_n578_ & ~new_n579_;
  assign new_n581_ = ~new_n577_ & new_n580_;
  assign new_n582_ = p_14 & ~new_n580_;
  assign new_n583_ = ~new_n581_ & ~new_n582_;
  assign new_n584_ = ~p_15 & n_75;
  assign new_n585_ = p_15 & ~n_75;
  assign new_n586_ = ~new_n584_ & ~new_n585_;
  assign new_n587_ = ~new_n583_ & new_n586_;
  assign new_n588_ = p_15 & ~new_n586_;
  assign new_n589_ = ~new_n587_ & ~new_n588_;
  assign new_n590_ = ~p_16 & n_76;
  assign new_n591_ = p_16 & ~n_76;
  assign new_n592_ = ~new_n590_ & ~new_n591_;
  assign new_n593_ = ~new_n589_ & new_n592_;
  assign new_n594_ = p_16 & ~new_n592_;
  assign new_n595_ = ~new_n593_ & ~new_n594_;
  assign new_n596_ = ~p_17 & n_77;
  assign new_n597_ = p_17 & ~n_77;
  assign new_n598_ = ~new_n596_ & ~new_n597_;
  assign new_n599_ = ~new_n595_ & new_n598_;
  assign new_n600_ = p_17 & ~new_n598_;
  assign new_n601_ = ~new_n599_ & ~new_n600_;
  assign new_n602_ = ~p_18 & n_78;
  assign new_n603_ = p_18 & ~n_78;
  assign new_n604_ = ~new_n602_ & ~new_n603_;
  assign new_n605_ = ~new_n601_ & new_n604_;
  assign new_n606_ = p_18 & ~new_n604_;
  assign new_n607_ = ~new_n605_ & ~new_n606_;
  assign new_n608_ = ~p_19 & n_79;
  assign new_n609_ = p_19 & ~n_79;
  assign new_n610_ = ~new_n608_ & ~new_n609_;
  assign new_n611_ = ~new_n607_ & new_n610_;
  assign new_n612_ = p_19 & ~new_n610_;
  assign new_n613_ = ~new_n611_ & ~new_n612_;
  assign new_n614_ = ~p_20 & n_80;
  assign new_n615_ = p_20 & ~n_80;
  assign new_n616_ = ~new_n614_ & ~new_n615_;
  assign new_n617_ = ~new_n613_ & new_n616_;
  assign new_n618_ = p_20 & ~new_n616_;
  assign new_n619_ = ~new_n617_ & ~new_n618_;
  assign new_n620_ = ~p_21 & n_81;
  assign new_n621_ = p_21 & ~n_81;
  assign new_n622_ = ~new_n620_ & ~new_n621_;
  assign new_n623_ = ~new_n619_ & new_n622_;
  assign new_n624_ = p_21 & ~new_n622_;
  assign new_n625_ = ~new_n623_ & ~new_n624_;
  assign new_n626_ = ~p_22 & n_82;
  assign new_n627_ = p_22 & ~n_82;
  assign new_n628_ = ~new_n626_ & ~new_n627_;
  assign new_n629_ = ~new_n625_ & new_n628_;
  assign new_n630_ = p_22 & ~new_n628_;
  assign new_n631_ = ~new_n629_ & ~new_n630_;
  assign new_n632_ = ~p_23 & n_83;
  assign new_n633_ = p_23 & ~n_83;
  assign new_n634_ = ~new_n632_ & ~new_n633_;
  assign new_n635_ = ~new_n631_ & new_n634_;
  assign new_n636_ = p_23 & ~new_n634_;
  assign new_n637_ = ~new_n635_ & ~new_n636_;
  assign new_n638_ = ~p_24 & n_84;
  assign new_n639_ = p_24 & ~n_84;
  assign new_n640_ = ~new_n638_ & ~new_n639_;
  assign new_n641_ = ~new_n637_ & new_n640_;
  assign new_n642_ = p_24 & ~new_n640_;
  assign new_n643_ = ~new_n641_ & ~new_n642_;
  assign new_n644_ = ~p_25 & n_85;
  assign new_n645_ = p_25 & ~n_85;
  assign new_n646_ = ~new_n644_ & ~new_n645_;
  assign new_n647_ = ~new_n643_ & new_n646_;
  assign new_n648_ = p_25 & ~new_n646_;
  assign new_n649_ = ~new_n647_ & ~new_n648_;
  assign new_n650_ = ~p_26 & n_86;
  assign new_n651_ = p_26 & ~n_86;
  assign new_n652_ = ~new_n650_ & ~new_n651_;
  assign new_n653_ = ~new_n649_ & new_n652_;
  assign new_n654_ = p_26 & ~new_n652_;
  assign new_n655_ = ~new_n653_ & ~new_n654_;
  assign new_n656_ = ~p_27 & n_87;
  assign new_n657_ = p_27 & ~n_87;
  assign new_n658_ = ~new_n656_ & ~new_n657_;
  assign new_n659_ = ~new_n655_ & new_n658_;
  assign new_n660_ = p_27 & ~new_n658_;
  assign new_n661_ = ~new_n659_ & ~new_n660_;
  assign new_n662_ = ~p_28 & n_88;
  assign new_n663_ = p_28 & ~n_88;
  assign new_n664_ = ~new_n662_ & ~new_n663_;
  assign new_n665_ = ~new_n661_ & new_n664_;
  assign new_n666_ = p_28 & ~new_n664_;
  assign new_n667_ = ~new_n665_ & ~new_n666_;
  assign new_n668_ = ~p_29 & n_89;
  assign new_n669_ = p_29 & ~n_89;
  assign new_n670_ = ~new_n668_ & ~new_n669_;
  assign new_n671_ = ~new_n667_ & new_n670_;
  assign new_n672_ = p_29 & ~new_n670_;
  assign new_n673_ = ~new_n671_ & ~new_n672_;
  assign new_n674_ = ~p_30 & n_90;
  assign new_n675_ = p_30 & ~n_90;
  assign new_n676_ = ~new_n674_ & ~new_n675_;
  assign new_n677_ = ~new_n673_ & new_n676_;
  assign new_n678_ = p_30 & ~new_n676_;
  assign new_n679_ = ~new_n677_ & ~new_n678_;
  assign new_n680_ = ~p_31 & n_91;
  assign new_n681_ = p_31 & ~n_91;
  assign new_n682_ = ~new_n680_ & ~new_n681_;
  assign new_n683_ = ~new_n679_ & new_n682_;
  assign new_n684_ = p_31 & ~new_n682_;
  assign new_n685_ = ~new_n683_ & ~new_n684_;
  assign new_n686_ = ~p_32 & n_92;
  assign new_n687_ = p_32 & ~n_92;
  assign new_n688_ = ~new_n686_ & ~new_n687_;
  assign new_n689_ = ~new_n685_ & new_n688_;
  assign new_n690_ = p_32 & ~new_n688_;
  assign new_n691_ = ~new_n689_ & ~new_n690_;
  assign new_n692_ = ~p_33 & n_93;
  assign new_n693_ = p_33 & ~n_93;
  assign new_n694_ = ~new_n692_ & ~new_n693_;
  assign new_n695_ = ~new_n691_ & new_n694_;
  assign new_n696_ = p_33 & ~new_n694_;
  assign new_n697_ = ~new_n695_ & ~new_n696_;
  assign new_n698_ = new_n336_ & ~new_n697_;
  assign new_n699_ = n_81 & new_n698_;
  assign new_n700_ = p_21 & ~new_n698_;
  assign new_n701_ = ~new_n699_ & ~new_n700_;
  assign new_n702_ = new_n336_ & ~new_n701_;
  assign new_n703_ = n_80 & new_n698_;
  assign new_n704_ = p_20 & ~new_n698_;
  assign new_n705_ = ~new_n703_ & ~new_n704_;
  assign new_n706_ = new_n336_ & ~new_n705_;
  assign new_n707_ = n_110 & ~new_n515_1_;
  assign new_n708_ = p_20 & new_n515_1_;
  assign new_n709_ = ~new_n707_ & ~new_n708_;
  assign new_n710_ = new_n336_ & ~new_n709_;
  assign new_n711_ = new_n706_ & new_n710_;
  assign new_n712_ = n_79 & new_n698_;
  assign new_n713_ = p_19 & ~new_n698_;
  assign new_n714_ = ~new_n712_ & ~new_n713_;
  assign new_n715_ = new_n336_ & ~new_n714_;
  assign new_n716_ = n_109 & ~new_n515_1_;
  assign new_n717_ = p_19 & new_n515_1_;
  assign new_n718_ = ~new_n716_ & ~new_n717_;
  assign new_n719_ = new_n336_ & ~new_n718_;
  assign new_n720_ = new_n715_ & new_n719_;
  assign new_n721_ = n_78 & new_n698_;
  assign new_n722_ = p_18 & ~new_n698_;
  assign new_n723_ = ~new_n721_ & ~new_n722_;
  assign new_n724_ = new_n336_ & ~new_n723_;
  assign new_n725_ = n_108 & ~new_n515_1_;
  assign new_n726_ = p_18 & new_n515_1_;
  assign new_n727_ = ~new_n725_ & ~new_n726_;
  assign new_n728_ = new_n336_ & ~new_n727_;
  assign new_n729_ = new_n724_ & new_n728_;
  assign new_n730_ = n_77 & new_n698_;
  assign new_n731_ = p_17 & ~new_n698_;
  assign new_n732_ = ~new_n730_ & ~new_n731_;
  assign new_n733_ = new_n336_ & ~new_n732_;
  assign new_n734_ = n_107 & ~new_n515_1_;
  assign new_n735_ = p_17 & new_n515_1_;
  assign new_n736_ = ~new_n734_ & ~new_n735_;
  assign new_n737_ = new_n336_ & ~new_n736_;
  assign new_n738_ = new_n733_ & new_n737_;
  assign new_n739_ = n_76 & new_n698_;
  assign new_n740_ = p_16 & ~new_n698_;
  assign new_n741_ = ~new_n739_ & ~new_n740_;
  assign new_n742_ = new_n336_ & ~new_n741_;
  assign new_n743_ = n_106 & ~new_n515_1_;
  assign new_n744_ = p_16 & new_n515_1_;
  assign new_n745_ = ~new_n743_ & ~new_n744_;
  assign new_n746_ = new_n336_ & ~new_n745_;
  assign new_n747_ = new_n742_ & new_n746_;
  assign new_n748_ = n_75 & new_n698_;
  assign new_n749_ = p_15 & ~new_n698_;
  assign new_n750_ = ~new_n748_ & ~new_n749_;
  assign new_n751_ = new_n336_ & ~new_n750_;
  assign new_n752_ = n_105 & ~new_n515_1_;
  assign new_n753_ = p_15 & new_n515_1_;
  assign new_n754_ = ~new_n752_ & ~new_n753_;
  assign new_n755_ = new_n336_ & ~new_n754_;
  assign new_n756_ = new_n751_ & new_n755_;
  assign new_n757_ = n_74 & new_n698_;
  assign new_n758_ = p_14 & ~new_n698_;
  assign new_n759_ = ~new_n757_ & ~new_n758_;
  assign new_n760_ = new_n336_ & ~new_n759_;
  assign new_n761_ = n_104 & ~new_n515_1_;
  assign new_n762_ = p_14 & new_n515_1_;
  assign new_n763_ = ~new_n761_ & ~new_n762_;
  assign new_n764_ = new_n336_ & ~new_n763_;
  assign new_n765_ = new_n760_ & new_n764_;
  assign new_n766_ = n_73 & new_n698_;
  assign new_n767_ = p_13 & ~new_n698_;
  assign new_n768_ = ~new_n766_ & ~new_n767_;
  assign new_n769_ = new_n336_ & ~new_n768_;
  assign new_n770_ = n_103 & ~new_n515_1_;
  assign new_n771_ = p_13 & new_n515_1_;
  assign new_n772_ = ~new_n770_ & ~new_n771_;
  assign new_n773_ = new_n336_ & ~new_n772_;
  assign new_n774_ = new_n769_ & new_n773_;
  assign new_n775_ = n_72 & new_n698_;
  assign new_n776_ = p_12 & ~new_n698_;
  assign new_n777_ = ~new_n775_ & ~new_n776_;
  assign new_n778_ = new_n336_ & ~new_n777_;
  assign new_n779_ = n_102 & ~new_n515_1_;
  assign new_n780_ = p_12 & new_n515_1_;
  assign new_n781_ = ~new_n779_ & ~new_n780_;
  assign new_n782_ = new_n336_ & ~new_n781_;
  assign new_n783_ = new_n778_ & new_n782_;
  assign new_n784_ = n_71 & new_n698_;
  assign new_n785_ = p_11 & ~new_n698_;
  assign new_n786_ = ~new_n784_ & ~new_n785_;
  assign new_n787_ = new_n336_ & ~new_n786_;
  assign new_n788_ = n_101 & ~new_n515_1_;
  assign new_n789_ = p_11 & new_n515_1_;
  assign new_n790_ = ~new_n788_ & ~new_n789_;
  assign new_n791_ = new_n336_ & ~new_n790_;
  assign new_n792_ = new_n787_ & new_n791_;
  assign new_n793_ = n_70 & new_n698_;
  assign new_n794_ = p_10 & ~new_n698_;
  assign new_n795_ = ~new_n793_ & ~new_n794_;
  assign new_n796_ = new_n336_ & ~new_n795_;
  assign new_n797_ = n_100 & ~new_n515_1_;
  assign new_n798_ = p_10 & new_n515_1_;
  assign new_n799_ = ~new_n797_ & ~new_n798_;
  assign new_n800_ = new_n336_ & ~new_n799_;
  assign new_n801_ = new_n796_ & new_n800_;
  assign new_n802_ = n_69 & new_n698_;
  assign new_n803_ = p_9 & ~new_n698_;
  assign new_n804_ = ~new_n802_ & ~new_n803_;
  assign new_n805_ = new_n336_ & ~new_n804_;
  assign new_n806_ = n_99 & ~new_n515_1_;
  assign new_n807_ = p_9 & new_n515_1_;
  assign new_n808_ = ~new_n806_ & ~new_n807_;
  assign new_n809_ = new_n336_ & ~new_n808_;
  assign new_n810_ = new_n805_ & new_n809_;
  assign new_n811_ = n_68 & new_n698_;
  assign new_n812_ = p_8 & ~new_n698_;
  assign new_n813_ = ~new_n811_ & ~new_n812_;
  assign new_n814_ = new_n336_ & ~new_n813_;
  assign new_n815_ = n_98 & ~new_n515_1_;
  assign new_n816_ = p_8 & new_n515_1_;
  assign new_n817_ = ~new_n815_ & ~new_n816_;
  assign new_n818_ = new_n336_ & ~new_n817_;
  assign new_n819_ = new_n814_ & new_n818_;
  assign new_n820_ = n_67 & new_n698_;
  assign new_n821_ = p_7 & ~new_n698_;
  assign new_n822_ = ~new_n820_ & ~new_n821_;
  assign new_n823_ = new_n336_ & ~new_n822_;
  assign new_n824_ = n_97 & ~new_n515_1_;
  assign new_n825_ = p_7 & new_n515_1_;
  assign new_n826_ = ~new_n824_ & ~new_n825_;
  assign new_n827_ = new_n336_ & ~new_n826_;
  assign new_n828_ = new_n823_ & new_n827_;
  assign new_n829_ = n_66 & new_n698_;
  assign new_n830_ = p_6 & ~new_n698_;
  assign new_n831_ = ~new_n829_ & ~new_n830_;
  assign new_n832_ = new_n336_ & ~new_n831_;
  assign new_n833_ = n_96 & ~new_n515_1_;
  assign new_n834_ = p_6 & new_n515_1_;
  assign new_n835_ = ~new_n833_ & ~new_n834_;
  assign new_n836_ = new_n336_ & ~new_n835_;
  assign new_n837_ = new_n832_ & new_n836_;
  assign new_n838_ = n_65 & new_n698_;
  assign new_n839_ = p_5 & ~new_n698_;
  assign new_n840_ = ~new_n838_ & ~new_n839_;
  assign new_n841_ = new_n336_ & ~new_n840_;
  assign new_n842_ = n_95 & ~new_n515_1_;
  assign new_n843_ = p_5 & new_n515_1_;
  assign new_n844_ = ~new_n842_ & ~new_n843_;
  assign new_n845_ = new_n336_ & ~new_n844_;
  assign new_n846_ = new_n841_ & new_n845_;
  assign new_n847_ = n_64 & new_n698_;
  assign new_n848_ = p_4 & ~new_n698_;
  assign new_n849_ = ~new_n847_ & ~new_n848_;
  assign new_n850_ = new_n336_ & ~new_n849_;
  assign new_n851_ = n_94 & ~new_n515_1_;
  assign new_n852_ = p_4 & new_n515_1_;
  assign new_n853_ = ~new_n851_ & ~new_n852_;
  assign new_n854_ = new_n336_ & ~new_n853_;
  assign new_n855_ = new_n850_ & new_n854_;
  assign new_n856_ = new_n845_ & new_n855_;
  assign new_n857_ = new_n841_ & new_n855_;
  assign new_n858_ = ~new_n846_ & ~new_n856_;
  assign new_n859_ = ~new_n857_ & new_n858_;
  assign new_n860_ = new_n836_ & ~new_n859_;
  assign new_n861_ = new_n832_ & ~new_n859_;
  assign new_n862_ = ~new_n837_ & ~new_n860_;
  assign new_n863_ = ~new_n861_ & new_n862_;
  assign new_n864_ = new_n827_ & ~new_n863_;
  assign new_n865_ = new_n823_ & ~new_n863_;
  assign new_n866_ = ~new_n828_ & ~new_n864_;
  assign new_n867_ = ~new_n865_ & new_n866_;
  assign new_n868_ = new_n818_ & ~new_n867_;
  assign new_n869_ = new_n814_ & ~new_n867_;
  assign new_n870_ = ~new_n819_ & ~new_n868_;
  assign new_n871_ = ~new_n869_ & new_n870_;
  assign new_n872_ = new_n809_ & ~new_n871_;
  assign new_n873_ = new_n805_ & ~new_n871_;
  assign new_n874_ = ~new_n810_ & ~new_n872_;
  assign new_n875_ = ~new_n873_ & new_n874_;
  assign new_n876_ = new_n800_ & ~new_n875_;
  assign new_n877_ = new_n796_ & ~new_n875_;
  assign new_n878_ = ~new_n801_ & ~new_n876_;
  assign new_n879_ = ~new_n877_ & new_n878_;
  assign new_n880_ = new_n791_ & ~new_n879_;
  assign new_n881_ = new_n787_ & ~new_n879_;
  assign new_n882_ = ~new_n792_ & ~new_n880_;
  assign new_n883_ = ~new_n881_ & new_n882_;
  assign new_n884_ = new_n782_ & ~new_n883_;
  assign new_n885_ = new_n778_ & ~new_n883_;
  assign new_n886_ = ~new_n783_ & ~new_n884_;
  assign new_n887_ = ~new_n885_ & new_n886_;
  assign new_n888_ = new_n773_ & ~new_n887_;
  assign new_n889_ = new_n769_ & ~new_n887_;
  assign new_n890_ = ~new_n774_ & ~new_n888_;
  assign new_n891_ = ~new_n889_ & new_n890_;
  assign new_n892_ = new_n764_ & ~new_n891_;
  assign new_n893_ = new_n760_ & ~new_n891_;
  assign new_n894_ = ~new_n765_ & ~new_n892_;
  assign new_n895_ = ~new_n893_ & new_n894_;
  assign new_n896_ = new_n755_ & ~new_n895_;
  assign new_n897_ = new_n751_ & ~new_n895_;
  assign new_n898_ = ~new_n756_ & ~new_n896_;
  assign new_n899_ = ~new_n897_ & new_n898_;
  assign new_n900_ = new_n746_ & ~new_n899_;
  assign new_n901_ = new_n742_ & ~new_n899_;
  assign new_n902_ = ~new_n747_ & ~new_n900_;
  assign new_n903_ = ~new_n901_ & new_n902_;
  assign new_n904_ = new_n737_ & ~new_n903_;
  assign new_n905_ = new_n733_ & ~new_n903_;
  assign new_n906_ = ~new_n738_ & ~new_n904_;
  assign new_n907_ = ~new_n905_ & new_n906_;
  assign new_n908_ = new_n728_ & ~new_n907_;
  assign new_n909_ = new_n724_ & ~new_n907_;
  assign new_n910_ = ~new_n729_ & ~new_n908_;
  assign new_n911_ = ~new_n909_ & new_n910_;
  assign new_n912_ = new_n719_ & ~new_n911_;
  assign new_n913_ = new_n715_ & ~new_n911_;
  assign new_n914_ = ~new_n720_ & ~new_n912_;
  assign new_n915_ = ~new_n913_ & new_n914_;
  assign new_n916_ = new_n710_ & ~new_n915_;
  assign new_n917_ = new_n706_ & ~new_n915_;
  assign new_n918_ = ~new_n711_ & ~new_n916_;
  assign new_n919_ = ~new_n917_ & new_n918_;
  assign new_n920_ = new_n519_ & new_n702_;
  assign new_n921_ = ~new_n919_ & new_n920_;
  assign new_n922_ = ~new_n519_ & new_n702_;
  assign new_n923_ = new_n919_ & new_n922_;
  assign new_n924_ = new_n519_ & ~new_n702_;
  assign new_n925_ = new_n919_ & new_n924_;
  assign new_n926_ = ~new_n519_ & ~new_n702_;
  assign new_n927_ = ~new_n919_ & new_n926_;
  assign new_n928_ = ~new_n921_ & ~new_n923_;
  assign new_n929_ = ~new_n925_ & ~new_n927_;
  assign new_n930_ = new_n928_ & new_n929_;
  assign new_n931_ = ~p_3 & ~new_n930_;
  assign new_n932_ = p_20 & p_3;
  assign new_n933_ = ~new_n931_ & ~new_n932_;
  assign new_n934_ = p_2 & ~new_n933_;
  assign new_n935_ = ~p_2 & n_50;
  assign new_n936_ = ~new_n934_ & ~new_n935_;
  assign p_140 = ~p_1 & ~new_n936_;
  assign new_n938_ = n_122 & ~new_n515_1_;
  assign new_n939_ = p_32 & new_n515_1_;
  assign new_n940_ = ~new_n938_ & ~new_n939_;
  assign new_n941_ = new_n336_ & ~new_n940_;
  assign new_n942_ = n_92 & new_n698_;
  assign new_n943_ = p_32 & ~new_n698_;
  assign new_n944_ = ~new_n942_ & ~new_n943_;
  assign new_n945_ = new_n336_ & ~new_n944_;
  assign new_n946_ = n_91 & new_n698_;
  assign new_n947_ = p_31 & ~new_n698_;
  assign new_n948_ = ~new_n946_ & ~new_n947_;
  assign new_n949_ = new_n336_ & ~new_n948_;
  assign new_n950_ = n_121 & ~new_n515_1_;
  assign new_n951_ = p_31 & new_n515_1_;
  assign new_n952_ = ~new_n950_ & ~new_n951_;
  assign new_n953_ = new_n336_ & ~new_n952_;
  assign new_n954_ = new_n949_ & new_n953_;
  assign new_n955_ = n_90 & new_n698_;
  assign new_n956_ = p_30 & ~new_n698_;
  assign new_n957_ = ~new_n955_ & ~new_n956_;
  assign new_n958_ = new_n336_ & ~new_n957_;
  assign new_n959_ = n_120 & ~new_n515_1_;
  assign new_n960_ = p_30 & new_n515_1_;
  assign new_n961_ = ~new_n959_ & ~new_n960_;
  assign new_n962_ = new_n336_ & ~new_n961_;
  assign new_n963_ = new_n958_ & new_n962_;
  assign new_n964_ = n_89 & new_n698_;
  assign new_n965_ = p_29 & ~new_n698_;
  assign new_n966_ = ~new_n964_ & ~new_n965_;
  assign new_n967_ = new_n336_ & ~new_n966_;
  assign new_n968_ = n_119 & ~new_n515_1_;
  assign new_n969_ = p_29 & new_n515_1_;
  assign new_n970_ = ~new_n968_ & ~new_n969_;
  assign new_n971_ = new_n336_ & ~new_n970_;
  assign new_n972_ = new_n967_ & new_n971_;
  assign new_n973_ = n_88 & new_n698_;
  assign new_n974_ = p_28 & ~new_n698_;
  assign new_n975_ = ~new_n973_ & ~new_n974_;
  assign new_n976_ = new_n336_ & ~new_n975_;
  assign new_n977_ = n_118 & ~new_n515_1_;
  assign new_n978_ = p_28 & new_n515_1_;
  assign new_n979_ = ~new_n977_ & ~new_n978_;
  assign new_n980_ = new_n336_ & ~new_n979_;
  assign new_n981_ = new_n976_ & new_n980_;
  assign new_n982_ = n_87 & new_n698_;
  assign new_n983_ = p_27 & ~new_n698_;
  assign new_n984_ = ~new_n982_ & ~new_n983_;
  assign new_n985_ = new_n336_ & ~new_n984_;
  assign new_n986_ = n_117 & ~new_n515_1_;
  assign new_n987_ = p_27 & new_n515_1_;
  assign new_n988_ = ~new_n986_ & ~new_n987_;
  assign new_n989_ = new_n336_ & ~new_n988_;
  assign new_n990_ = new_n985_ & new_n989_;
  assign new_n991_ = n_86 & new_n698_;
  assign new_n992_ = p_26 & ~new_n698_;
  assign new_n993_ = ~new_n991_ & ~new_n992_;
  assign new_n994_ = new_n336_ & ~new_n993_;
  assign new_n995_ = n_116 & ~new_n515_1_;
  assign new_n996_ = p_26 & new_n515_1_;
  assign new_n997_ = ~new_n995_ & ~new_n996_;
  assign new_n998_ = new_n336_ & ~new_n997_;
  assign new_n999_ = new_n994_ & new_n998_;
  assign new_n1000_ = n_85 & new_n698_;
  assign new_n1001_ = p_25 & ~new_n698_;
  assign new_n1002_ = ~new_n1000_ & ~new_n1001_;
  assign new_n1003_ = new_n336_ & ~new_n1002_;
  assign new_n1004_ = n_115 & ~new_n515_1_;
  assign new_n1005_ = p_25 & new_n515_1_;
  assign new_n1006_ = ~new_n1004_ & ~new_n1005_;
  assign new_n1007_ = new_n336_ & ~new_n1006_;
  assign new_n1008_ = new_n1003_ & new_n1007_;
  assign new_n1009_ = n_84 & new_n698_;
  assign new_n1010_ = p_24 & ~new_n698_;
  assign new_n1011_ = ~new_n1009_ & ~new_n1010_;
  assign new_n1012_ = new_n336_ & ~new_n1011_;
  assign new_n1013_ = n_114 & ~new_n515_1_;
  assign new_n1014_ = p_24 & new_n515_1_;
  assign new_n1015_ = ~new_n1013_ & ~new_n1014_;
  assign new_n1016_ = new_n336_ & ~new_n1015_;
  assign new_n1017_ = new_n1012_ & new_n1016_;
  assign new_n1018_ = n_83 & new_n698_;
  assign new_n1019_ = p_23 & ~new_n698_;
  assign new_n1020_ = ~new_n1018_ & ~new_n1019_;
  assign new_n1021_ = new_n336_ & ~new_n1020_;
  assign new_n1022_ = n_113 & ~new_n515_1_;
  assign new_n1023_ = p_23 & new_n515_1_;
  assign new_n1024_ = ~new_n1022_ & ~new_n1023_;
  assign new_n1025_ = new_n336_ & ~new_n1024_;
  assign new_n1026_ = new_n1021_ & new_n1025_;
  assign new_n1027_ = n_82 & new_n698_;
  assign new_n1028_ = p_22 & ~new_n698_;
  assign new_n1029_ = ~new_n1027_ & ~new_n1028_;
  assign new_n1030_ = new_n336_ & ~new_n1029_;
  assign new_n1031_ = n_112 & ~new_n515_1_;
  assign new_n1032_ = p_22 & new_n515_1_;
  assign new_n1033_ = ~new_n1031_ & ~new_n1032_;
  assign new_n1034_ = new_n336_ & ~new_n1033_;
  assign new_n1035_ = new_n1030_ & new_n1034_;
  assign new_n1036_ = new_n519_ & ~new_n919_;
  assign new_n1037_ = new_n702_ & ~new_n919_;
  assign new_n1038_ = ~new_n920_ & ~new_n1036_;
  assign new_n1039_ = ~new_n1037_ & new_n1038_;
  assign new_n1040_ = new_n1034_ & ~new_n1039_;
  assign new_n1041_ = new_n1030_ & ~new_n1039_;
  assign new_n1042_ = ~new_n1035_ & ~new_n1040_;
  assign new_n1043_ = ~new_n1041_ & new_n1042_;
  assign new_n1044_ = new_n1025_ & ~new_n1043_;
  assign new_n1045_ = new_n1021_ & ~new_n1043_;
  assign new_n1046_ = ~new_n1026_ & ~new_n1044_;
  assign new_n1047_ = ~new_n1045_ & new_n1046_;
  assign new_n1048_ = new_n1016_ & ~new_n1047_;
  assign new_n1049_ = new_n1012_ & ~new_n1047_;
  assign new_n1050_ = ~new_n1017_ & ~new_n1048_;
  assign new_n1051_ = ~new_n1049_ & new_n1050_;
  assign new_n1052_ = new_n1007_ & ~new_n1051_;
  assign new_n1053_ = new_n1003_ & ~new_n1051_;
  assign new_n1054_ = ~new_n1008_ & ~new_n1052_;
  assign new_n1055_ = ~new_n1053_ & new_n1054_;
  assign new_n1056_ = new_n998_ & ~new_n1055_;
  assign new_n1057_ = new_n994_ & ~new_n1055_;
  assign new_n1058_ = ~new_n999_ & ~new_n1056_;
  assign new_n1059_ = ~new_n1057_ & new_n1058_;
  assign new_n1060_ = new_n989_ & ~new_n1059_;
  assign new_n1061_ = new_n985_ & ~new_n1059_;
  assign new_n1062_ = ~new_n990_ & ~new_n1060_;
  assign new_n1063_ = ~new_n1061_ & new_n1062_;
  assign new_n1064_ = new_n980_ & ~new_n1063_;
  assign new_n1065_ = new_n976_ & ~new_n1063_;
  assign new_n1066_ = ~new_n981_ & ~new_n1064_;
  assign new_n1067_ = ~new_n1065_ & new_n1066_;
  assign new_n1068_ = new_n971_ & ~new_n1067_;
  assign new_n1069_ = new_n967_ & ~new_n1067_;
  assign new_n1070_ = ~new_n972_ & ~new_n1068_;
  assign new_n1071_ = ~new_n1069_ & new_n1070_;
  assign new_n1072_ = new_n962_ & ~new_n1071_;
  assign new_n1073_ = new_n958_ & ~new_n1071_;
  assign new_n1074_ = ~new_n963_ & ~new_n1072_;
  assign new_n1075_ = ~new_n1073_ & new_n1074_;
  assign new_n1076_ = new_n953_ & ~new_n1075_;
  assign new_n1077_ = new_n949_ & ~new_n1075_;
  assign new_n1078_ = ~new_n954_ & ~new_n1076_;
  assign new_n1079_ = ~new_n1077_ & new_n1078_;
  assign new_n1080_ = new_n941_ & new_n945_;
  assign new_n1081_ = ~new_n1079_ & new_n1080_;
  assign new_n1082_ = ~new_n941_ & new_n945_;
  assign new_n1083_ = new_n1079_ & new_n1082_;
  assign new_n1084_ = new_n941_ & ~new_n945_;
  assign new_n1085_ = new_n1079_ & new_n1084_;
  assign new_n1086_ = ~new_n941_ & ~new_n945_;
  assign new_n1087_ = ~new_n1079_ & new_n1086_;
  assign new_n1088_ = ~new_n1081_ & ~new_n1083_;
  assign new_n1089_ = ~new_n1085_ & ~new_n1087_;
  assign new_n1090_ = new_n1088_ & new_n1089_;
  assign new_n1091_ = ~p_3 & ~new_n1090_;
  assign new_n1092_ = p_31 & p_3;
  assign new_n1093_ = ~new_n1091_ & ~new_n1092_;
  assign new_n1094_ = p_2 & ~new_n1093_;
  assign new_n1095_ = ~p_2 & n_61;
  assign new_n1096_ = ~new_n1094_ & ~new_n1095_;
  assign p_151 = ~p_1 & ~new_n1096_;
  assign new_n1098_ = new_n792_ & ~new_n879_;
  assign new_n1099_ = new_n787_ & ~new_n791_;
  assign new_n1100_ = new_n879_ & new_n1099_;
  assign new_n1101_ = ~new_n787_ & new_n791_;
  assign new_n1102_ = new_n879_ & new_n1101_;
  assign new_n1103_ = ~new_n787_ & ~new_n791_;
  assign new_n1104_ = ~new_n879_ & new_n1103_;
  assign new_n1105_ = ~new_n1098_ & ~new_n1100_;
  assign new_n1106_ = ~new_n1102_ & ~new_n1104_;
  assign new_n1107_ = new_n1105_ & new_n1106_;
  assign new_n1108_ = ~p_3 & ~new_n1107_;
  assign new_n1109_ = p_10 & p_3;
  assign new_n1110_ = ~new_n1108_ & ~new_n1109_;
  assign new_n1111_ = p_2 & ~new_n1110_;
  assign new_n1112_ = ~p_2 & n_40;
  assign new_n1113_ = ~new_n1111_ & ~new_n1112_;
  assign p_130 = ~p_1 & ~new_n1113_;
  assign new_n1115_ = n_123 & ~new_n515_1_;
  assign new_n1116_ = p_33 & new_n515_1_;
  assign new_n1117_ = ~new_n1115_ & ~new_n1116_;
  assign new_n1118_ = new_n336_ & ~new_n1117_;
  assign new_n1119_ = n_93 & new_n698_;
  assign new_n1120_ = p_33 & ~new_n698_;
  assign new_n1121_ = ~new_n1119_ & ~new_n1120_;
  assign new_n1122_ = new_n336_ & ~new_n1121_;
  assign new_n1123_ = new_n941_ & ~new_n1079_;
  assign new_n1124_ = new_n945_ & ~new_n1079_;
  assign new_n1125_ = ~new_n1080_ & ~new_n1123_;
  assign new_n1126_ = ~new_n1124_ & new_n1125_;
  assign new_n1127_ = new_n1118_ & new_n1122_;
  assign new_n1128_ = ~new_n1126_ & new_n1127_;
  assign new_n1129_ = ~new_n1118_ & new_n1122_;
  assign new_n1130_ = new_n1126_ & new_n1129_;
  assign new_n1131_ = new_n1118_ & ~new_n1122_;
  assign new_n1132_ = new_n1126_ & new_n1131_;
  assign new_n1133_ = ~new_n1118_ & ~new_n1122_;
  assign new_n1134_ = ~new_n1126_ & new_n1133_;
  assign new_n1135_ = ~new_n1128_ & ~new_n1130_;
  assign new_n1136_ = ~new_n1132_ & ~new_n1134_;
  assign new_n1137_ = new_n1135_ & new_n1136_;
  assign new_n1138_ = ~p_3 & ~new_n1137_;
  assign new_n1139_ = p_32 & p_3;
  assign new_n1140_ = ~new_n1138_ & ~new_n1139_;
  assign new_n1141_ = p_2 & ~new_n1140_;
  assign new_n1142_ = ~p_2 & n_62;
  assign new_n1143_ = ~new_n1141_ & ~new_n1142_;
  assign p_152 = ~p_1 & ~new_n1143_;
  assign new_n1145_ = new_n1118_ & ~new_n1126_;
  assign new_n1146_ = new_n1122_ & ~new_n1126_;
  assign new_n1147_ = ~new_n1127_ & ~new_n1145_;
  assign new_n1148_ = ~new_n1146_ & new_n1147_;
  assign new_n1149_ = ~p_3 & ~new_n1148_;
  assign new_n1150_ = p_33 & p_3;
  assign new_n1151_ = ~new_n1149_ & ~new_n1150_;
  assign new_n1152_ = p_2 & ~new_n1151_;
  assign new_n1153_ = ~p_2 & n_63;
  assign new_n1154_ = ~new_n1152_ & ~new_n1153_;
  assign p_153 = ~p_1 & ~new_n1154_;
  assign new_n1156_ = new_n765_ & ~new_n891_;
  assign new_n1157_ = new_n760_ & ~new_n764_;
  assign new_n1158_ = new_n891_ & new_n1157_;
  assign new_n1159_ = ~new_n760_ & new_n764_;
  assign new_n1160_ = new_n891_ & new_n1159_;
  assign new_n1161_ = ~new_n760_ & ~new_n764_;
  assign new_n1162_ = ~new_n891_ & new_n1161_;
  assign new_n1163_ = ~new_n1156_ & ~new_n1158_;
  assign new_n1164_ = ~new_n1160_ & ~new_n1162_;
  assign new_n1165_ = new_n1163_ & new_n1164_;
  assign new_n1166_ = ~p_3 & ~new_n1165_;
  assign new_n1167_ = p_13 & p_3;
  assign new_n1168_ = ~new_n1166_ & ~new_n1167_;
  assign new_n1169_ = p_2 & ~new_n1168_;
  assign new_n1170_ = ~p_2 & n_43;
  assign new_n1171_ = ~new_n1169_ & ~new_n1170_;
  assign p_133 = ~p_1 & ~new_n1171_;
  assign new_n1173_ = new_n1008_ & ~new_n1051_;
  assign new_n1174_ = new_n1003_ & ~new_n1007_;
  assign new_n1175_ = new_n1051_ & new_n1174_;
  assign new_n1176_ = ~new_n1003_ & new_n1007_;
  assign new_n1177_ = new_n1051_ & new_n1176_;
  assign new_n1178_ = ~new_n1003_ & ~new_n1007_;
  assign new_n1179_ = ~new_n1051_ & new_n1178_;
  assign new_n1180_ = ~new_n1173_ & ~new_n1175_;
  assign new_n1181_ = ~new_n1177_ & ~new_n1179_;
  assign new_n1182_ = new_n1180_ & new_n1181_;
  assign new_n1183_ = ~p_3 & ~new_n1182_;
  assign new_n1184_ = p_24 & p_3;
  assign new_n1185_ = ~new_n1183_ & ~new_n1184_;
  assign new_n1186_ = p_2 & ~new_n1185_;
  assign new_n1187_ = ~p_2 & n_54;
  assign new_n1188_ = ~new_n1186_ & ~new_n1187_;
  assign p_144 = ~p_1 & ~new_n1188_;
  assign new_n1190_ = new_n756_ & ~new_n895_;
  assign new_n1191_ = new_n751_ & ~new_n755_;
  assign new_n1192_ = new_n895_ & new_n1191_;
  assign new_n1193_ = ~new_n751_ & new_n755_;
  assign new_n1194_ = new_n895_ & new_n1193_;
  assign new_n1195_ = ~new_n751_ & ~new_n755_;
  assign new_n1196_ = ~new_n895_ & new_n1195_;
  assign new_n1197_ = ~new_n1190_ & ~new_n1192_;
  assign new_n1198_ = ~new_n1194_ & ~new_n1196_;
  assign new_n1199_ = new_n1197_ & new_n1198_;
  assign new_n1200_ = ~p_3 & ~new_n1199_;
  assign new_n1201_ = p_14 & p_3;
  assign new_n1202_ = ~new_n1200_ & ~new_n1201_;
  assign new_n1203_ = p_2 & ~new_n1202_;
  assign new_n1204_ = ~p_2 & n_44;
  assign new_n1205_ = ~new_n1203_ & ~new_n1204_;
  assign p_134 = ~p_1 & ~new_n1205_;
  assign new_n1207_ = new_n1017_ & ~new_n1047_;
  assign new_n1208_ = new_n1012_ & ~new_n1016_;
  assign new_n1209_ = new_n1047_ & new_n1208_;
  assign new_n1210_ = ~new_n1012_ & new_n1016_;
  assign new_n1211_ = new_n1047_ & new_n1210_;
  assign new_n1212_ = ~new_n1012_ & ~new_n1016_;
  assign new_n1213_ = ~new_n1047_ & new_n1212_;
  assign new_n1214_ = ~new_n1207_ & ~new_n1209_;
  assign new_n1215_ = ~new_n1211_ & ~new_n1213_;
  assign new_n1216_ = new_n1214_ & new_n1215_;
  assign new_n1217_ = ~p_3 & ~new_n1216_;
  assign new_n1218_ = p_23 & p_3;
  assign new_n1219_ = ~new_n1217_ & ~new_n1218_;
  assign new_n1220_ = p_2 & ~new_n1219_;
  assign new_n1221_ = ~p_2 & n_53;
  assign new_n1222_ = ~new_n1220_ & ~new_n1221_;
  assign p_143 = ~p_1 & ~new_n1222_;
  assign new_n1224_ = new_n846_ & new_n855_;
  assign new_n1225_ = new_n841_ & ~new_n845_;
  assign new_n1226_ = ~new_n855_ & new_n1225_;
  assign new_n1227_ = ~new_n841_ & new_n845_;
  assign new_n1228_ = ~new_n855_ & new_n1227_;
  assign new_n1229_ = ~new_n841_ & ~new_n845_;
  assign new_n1230_ = new_n855_ & new_n1229_;
  assign new_n1231_ = ~new_n1224_ & ~new_n1226_;
  assign new_n1232_ = ~new_n1228_ & ~new_n1230_;
  assign new_n1233_ = new_n1231_ & new_n1232_;
  assign new_n1234_ = ~p_3 & ~new_n1233_;
  assign new_n1235_ = p_4 & p_3;
  assign new_n1236_ = ~new_n1234_ & ~new_n1235_;
  assign new_n1237_ = p_2 & ~new_n1236_;
  assign new_n1238_ = ~p_2 & n_34;
  assign new_n1239_ = ~new_n1237_ & ~new_n1238_;
  assign p_124 = ~p_1 & ~new_n1239_;
  assign new_n1241_ = new_n783_ & ~new_n883_;
  assign new_n1242_ = new_n778_ & ~new_n782_;
  assign new_n1243_ = new_n883_ & new_n1242_;
  assign new_n1244_ = ~new_n778_ & new_n782_;
  assign new_n1245_ = new_n883_ & new_n1244_;
  assign new_n1246_ = ~new_n778_ & ~new_n782_;
  assign new_n1247_ = ~new_n883_ & new_n1246_;
  assign new_n1248_ = ~new_n1241_ & ~new_n1243_;
  assign new_n1249_ = ~new_n1245_ & ~new_n1247_;
  assign new_n1250_ = new_n1248_ & new_n1249_;
  assign new_n1251_ = ~p_3 & ~new_n1250_;
  assign new_n1252_ = p_11 & p_3;
  assign new_n1253_ = ~new_n1251_ & ~new_n1252_;
  assign new_n1254_ = p_2 & ~new_n1253_;
  assign new_n1255_ = ~p_2 & n_41;
  assign new_n1256_ = ~new_n1254_ & ~new_n1255_;
  assign p_131 = ~p_1 & ~new_n1256_;
  assign new_n1258_ = new_n1026_ & ~new_n1043_;
  assign new_n1259_ = new_n1021_ & ~new_n1025_;
  assign new_n1260_ = new_n1043_ & new_n1259_;
  assign new_n1261_ = ~new_n1021_ & new_n1025_;
  assign new_n1262_ = new_n1043_ & new_n1261_;
  assign new_n1263_ = ~new_n1021_ & ~new_n1025_;
  assign new_n1264_ = ~new_n1043_ & new_n1263_;
  assign new_n1265_ = ~new_n1258_ & ~new_n1260_;
  assign new_n1266_ = ~new_n1262_ & ~new_n1264_;
  assign new_n1267_ = new_n1265_ & new_n1266_;
  assign new_n1268_ = ~p_3 & ~new_n1267_;
  assign new_n1269_ = p_22 & p_3;
  assign new_n1270_ = ~new_n1268_ & ~new_n1269_;
  assign new_n1271_ = p_2 & ~new_n1270_;
  assign new_n1272_ = ~p_2 & n_52;
  assign new_n1273_ = ~new_n1271_ & ~new_n1272_;
  assign p_142 = ~p_1 & ~new_n1273_;
  assign new_n1275_ = new_n774_ & ~new_n887_;
  assign new_n1276_ = new_n769_ & ~new_n773_;
  assign new_n1277_ = new_n887_ & new_n1276_;
  assign new_n1278_ = ~new_n769_ & new_n773_;
  assign new_n1279_ = new_n887_ & new_n1278_;
  assign new_n1280_ = ~new_n769_ & ~new_n773_;
  assign new_n1281_ = ~new_n887_ & new_n1280_;
  assign new_n1282_ = ~new_n1275_ & ~new_n1277_;
  assign new_n1283_ = ~new_n1279_ & ~new_n1281_;
  assign new_n1284_ = new_n1282_ & new_n1283_;
  assign new_n1285_ = ~p_3 & ~new_n1284_;
  assign new_n1286_ = p_12 & p_3;
  assign new_n1287_ = ~new_n1285_ & ~new_n1286_;
  assign new_n1288_ = p_2 & ~new_n1287_;
  assign new_n1289_ = ~p_2 & n_42;
  assign new_n1290_ = ~new_n1288_ & ~new_n1289_;
  assign p_132 = ~p_1 & ~new_n1290_;
  assign new_n1292_ = new_n1035_ & ~new_n1039_;
  assign new_n1293_ = new_n1030_ & ~new_n1034_;
  assign new_n1294_ = new_n1039_ & new_n1293_;
  assign new_n1295_ = ~new_n1030_ & new_n1034_;
  assign new_n1296_ = new_n1039_ & new_n1295_;
  assign new_n1297_ = ~new_n1030_ & ~new_n1034_;
  assign new_n1298_ = ~new_n1039_ & new_n1297_;
  assign new_n1299_ = ~new_n1292_ & ~new_n1294_;
  assign new_n1300_ = ~new_n1296_ & ~new_n1298_;
  assign new_n1301_ = new_n1299_ & new_n1300_;
  assign new_n1302_ = ~p_3 & ~new_n1301_;
  assign new_n1303_ = p_21 & p_3;
  assign new_n1304_ = ~new_n1302_ & ~new_n1303_;
  assign new_n1305_ = p_2 & ~new_n1304_;
  assign new_n1306_ = ~p_2 & n_51;
  assign new_n1307_ = ~new_n1305_ & ~new_n1306_;
  assign p_141 = ~p_1 & ~new_n1307_;
  assign new_n1309_ = new_n954_ & ~new_n1075_;
  assign new_n1310_ = new_n949_ & ~new_n953_;
  assign new_n1311_ = new_n1075_ & new_n1310_;
  assign new_n1312_ = ~new_n949_ & new_n953_;
  assign new_n1313_ = new_n1075_ & new_n1312_;
  assign new_n1314_ = ~new_n949_ & ~new_n953_;
  assign new_n1315_ = ~new_n1075_ & new_n1314_;
  assign new_n1316_ = ~new_n1309_ & ~new_n1311_;
  assign new_n1317_ = ~new_n1313_ & ~new_n1315_;
  assign new_n1318_ = new_n1316_ & new_n1317_;
  assign new_n1319_ = ~p_3 & ~new_n1318_;
  assign new_n1320_ = p_30 & p_3;
  assign new_n1321_ = ~new_n1319_ & ~new_n1320_;
  assign new_n1322_ = p_2 & ~new_n1321_;
  assign new_n1323_ = ~p_2 & n_60;
  assign new_n1324_ = ~new_n1322_ & ~new_n1323_;
  assign p_150 = ~p_1 & ~new_n1324_;
  assign new_n1326_ = new_n828_ & ~new_n863_;
  assign new_n1327_ = new_n823_ & ~new_n827_;
  assign new_n1328_ = new_n863_ & new_n1327_;
  assign new_n1329_ = ~new_n823_ & new_n827_;
  assign new_n1330_ = new_n863_ & new_n1329_;
  assign new_n1331_ = ~new_n823_ & ~new_n827_;
  assign new_n1332_ = ~new_n863_ & new_n1331_;
  assign new_n1333_ = ~new_n1326_ & ~new_n1328_;
  assign new_n1334_ = ~new_n1330_ & ~new_n1332_;
  assign new_n1335_ = new_n1333_ & new_n1334_;
  assign new_n1336_ = ~p_3 & ~new_n1335_;
  assign new_n1337_ = p_6 & p_3;
  assign new_n1338_ = ~new_n1336_ & ~new_n1337_;
  assign new_n1339_ = p_2 & ~new_n1338_;
  assign new_n1340_ = ~p_2 & n_36;
  assign new_n1341_ = ~new_n1339_ & ~new_n1340_;
  assign p_126 = ~p_1 & ~new_n1341_;
  assign new_n1343_ = new_n729_ & ~new_n907_;
  assign new_n1344_ = new_n724_ & ~new_n728_;
  assign new_n1345_ = new_n907_ & new_n1344_;
  assign new_n1346_ = ~new_n724_ & new_n728_;
  assign new_n1347_ = new_n907_ & new_n1346_;
  assign new_n1348_ = ~new_n724_ & ~new_n728_;
  assign new_n1349_ = ~new_n907_ & new_n1348_;
  assign new_n1350_ = ~new_n1343_ & ~new_n1345_;
  assign new_n1351_ = ~new_n1347_ & ~new_n1349_;
  assign new_n1352_ = new_n1350_ & new_n1351_;
  assign new_n1353_ = ~p_3 & ~new_n1352_;
  assign new_n1354_ = p_17 & p_3;
  assign new_n1355_ = ~new_n1353_ & ~new_n1354_;
  assign new_n1356_ = p_2 & ~new_n1355_;
  assign new_n1357_ = ~p_2 & n_47;
  assign new_n1358_ = ~new_n1356_ & ~new_n1357_;
  assign p_137 = ~p_1 & ~new_n1358_;
  assign new_n1360_ = new_n972_ & ~new_n1067_;
  assign new_n1361_ = new_n967_ & ~new_n971_;
  assign new_n1362_ = new_n1067_ & new_n1361_;
  assign new_n1363_ = ~new_n967_ & new_n971_;
  assign new_n1364_ = new_n1067_ & new_n1363_;
  assign new_n1365_ = ~new_n967_ & ~new_n971_;
  assign new_n1366_ = ~new_n1067_ & new_n1365_;
  assign new_n1367_ = ~new_n1360_ & ~new_n1362_;
  assign new_n1368_ = ~new_n1364_ & ~new_n1366_;
  assign new_n1369_ = new_n1367_ & new_n1368_;
  assign new_n1370_ = ~p_3 & ~new_n1369_;
  assign new_n1371_ = p_28 & p_3;
  assign new_n1372_ = ~new_n1370_ & ~new_n1371_;
  assign new_n1373_ = p_2 & ~new_n1372_;
  assign new_n1374_ = ~p_2 & n_58;
  assign new_n1375_ = ~new_n1373_ & ~new_n1374_;
  assign p_148 = ~p_1 & ~new_n1375_;
  assign new_n1377_ = new_n837_ & ~new_n859_;
  assign new_n1378_ = new_n832_ & ~new_n836_;
  assign new_n1379_ = new_n859_ & new_n1378_;
  assign new_n1380_ = ~new_n832_ & new_n836_;
  assign new_n1381_ = new_n859_ & new_n1380_;
  assign new_n1382_ = ~new_n832_ & ~new_n836_;
  assign new_n1383_ = ~new_n859_ & new_n1382_;
  assign new_n1384_ = ~new_n1377_ & ~new_n1379_;
  assign new_n1385_ = ~new_n1381_ & ~new_n1383_;
  assign new_n1386_ = new_n1384_ & new_n1385_;
  assign new_n1387_ = ~p_3 & ~new_n1386_;
  assign new_n1388_ = p_5 & p_3;
  assign new_n1389_ = ~new_n1387_ & ~new_n1388_;
  assign new_n1390_ = p_2 & ~new_n1389_;
  assign new_n1391_ = ~p_2 & n_35;
  assign new_n1392_ = ~new_n1390_ & ~new_n1391_;
  assign p_125 = ~p_1 & ~new_n1392_;
  assign new_n1394_ = new_n720_ & ~new_n911_;
  assign new_n1395_ = new_n715_ & ~new_n719_;
  assign new_n1396_ = new_n911_ & new_n1395_;
  assign new_n1397_ = ~new_n715_ & new_n719_;
  assign new_n1398_ = new_n911_ & new_n1397_;
  assign new_n1399_ = ~new_n715_ & ~new_n719_;
  assign new_n1400_ = ~new_n911_ & new_n1399_;
  assign new_n1401_ = ~new_n1394_ & ~new_n1396_;
  assign new_n1402_ = ~new_n1398_ & ~new_n1400_;
  assign new_n1403_ = new_n1401_ & new_n1402_;
  assign new_n1404_ = ~p_3 & ~new_n1403_;
  assign new_n1405_ = p_18 & p_3;
  assign new_n1406_ = ~new_n1404_ & ~new_n1405_;
  assign new_n1407_ = p_2 & ~new_n1406_;
  assign new_n1408_ = ~p_2 & n_48;
  assign new_n1409_ = ~new_n1407_ & ~new_n1408_;
  assign p_138 = ~p_1 & ~new_n1409_;
  assign new_n1411_ = new_n981_ & ~new_n1063_;
  assign new_n1412_ = new_n976_ & ~new_n980_;
  assign new_n1413_ = new_n1063_ & new_n1412_;
  assign new_n1414_ = ~new_n976_ & new_n980_;
  assign new_n1415_ = new_n1063_ & new_n1414_;
  assign new_n1416_ = ~new_n976_ & ~new_n980_;
  assign new_n1417_ = ~new_n1063_ & new_n1416_;
  assign new_n1418_ = ~new_n1411_ & ~new_n1413_;
  assign new_n1419_ = ~new_n1415_ & ~new_n1417_;
  assign new_n1420_ = new_n1418_ & new_n1419_;
  assign new_n1421_ = ~p_3 & ~new_n1420_;
  assign new_n1422_ = p_27 & p_3;
  assign new_n1423_ = ~new_n1421_ & ~new_n1422_;
  assign new_n1424_ = p_2 & ~new_n1423_;
  assign new_n1425_ = ~p_2 & n_57;
  assign new_n1426_ = ~new_n1424_ & ~new_n1425_;
  assign p_147 = ~p_1 & ~new_n1426_;
  assign new_n1428_ = new_n810_ & ~new_n871_;
  assign new_n1429_ = new_n805_ & ~new_n809_;
  assign new_n1430_ = new_n871_ & new_n1429_;
  assign new_n1431_ = ~new_n805_ & new_n809_;
  assign new_n1432_ = new_n871_ & new_n1431_;
  assign new_n1433_ = ~new_n805_ & ~new_n809_;
  assign new_n1434_ = ~new_n871_ & new_n1433_;
  assign new_n1435_ = ~new_n1428_ & ~new_n1430_;
  assign new_n1436_ = ~new_n1432_ & ~new_n1434_;
  assign new_n1437_ = new_n1435_ & new_n1436_;
  assign new_n1438_ = ~p_3 & ~new_n1437_;
  assign new_n1439_ = p_8 & p_3;
  assign new_n1440_ = ~new_n1438_ & ~new_n1439_;
  assign new_n1441_ = p_2 & ~new_n1440_;
  assign new_n1442_ = ~p_2 & n_38;
  assign new_n1443_ = ~new_n1441_ & ~new_n1442_;
  assign p_128 = ~p_1 & ~new_n1443_;
  assign new_n1445_ = new_n747_ & ~new_n899_;
  assign new_n1446_ = new_n742_ & ~new_n746_;
  assign new_n1447_ = new_n899_ & new_n1446_;
  assign new_n1448_ = ~new_n742_ & new_n746_;
  assign new_n1449_ = new_n899_ & new_n1448_;
  assign new_n1450_ = ~new_n742_ & ~new_n746_;
  assign new_n1451_ = ~new_n899_ & new_n1450_;
  assign new_n1452_ = ~new_n1445_ & ~new_n1447_;
  assign new_n1453_ = ~new_n1449_ & ~new_n1451_;
  assign new_n1454_ = new_n1452_ & new_n1453_;
  assign new_n1455_ = ~p_3 & ~new_n1454_;
  assign new_n1456_ = p_15 & p_3;
  assign new_n1457_ = ~new_n1455_ & ~new_n1456_;
  assign new_n1458_ = p_2 & ~new_n1457_;
  assign new_n1459_ = ~p_2 & n_45;
  assign new_n1460_ = ~new_n1458_ & ~new_n1459_;
  assign p_135 = ~p_1 & ~new_n1460_;
  assign new_n1462_ = new_n990_ & ~new_n1059_;
  assign new_n1463_ = new_n985_ & ~new_n989_;
  assign new_n1464_ = new_n1059_ & new_n1463_;
  assign new_n1465_ = ~new_n985_ & new_n989_;
  assign new_n1466_ = new_n1059_ & new_n1465_;
  assign new_n1467_ = ~new_n985_ & ~new_n989_;
  assign new_n1468_ = ~new_n1059_ & new_n1467_;
  assign new_n1469_ = ~new_n1462_ & ~new_n1464_;
  assign new_n1470_ = ~new_n1466_ & ~new_n1468_;
  assign new_n1471_ = new_n1469_ & new_n1470_;
  assign new_n1472_ = ~p_3 & ~new_n1471_;
  assign new_n1473_ = p_26 & p_3;
  assign new_n1474_ = ~new_n1472_ & ~new_n1473_;
  assign new_n1475_ = p_2 & ~new_n1474_;
  assign new_n1476_ = ~p_2 & n_56;
  assign new_n1477_ = ~new_n1475_ & ~new_n1476_;
  assign p_146 = ~p_1 & ~new_n1477_;
  assign new_n1479_ = new_n819_ & ~new_n867_;
  assign new_n1480_ = new_n814_ & ~new_n818_;
  assign new_n1481_ = new_n867_ & new_n1480_;
  assign new_n1482_ = ~new_n814_ & new_n818_;
  assign new_n1483_ = new_n867_ & new_n1482_;
  assign new_n1484_ = ~new_n814_ & ~new_n818_;
  assign new_n1485_ = ~new_n867_ & new_n1484_;
  assign new_n1486_ = ~new_n1479_ & ~new_n1481_;
  assign new_n1487_ = ~new_n1483_ & ~new_n1485_;
  assign new_n1488_ = new_n1486_ & new_n1487_;
  assign new_n1489_ = ~p_3 & ~new_n1488_;
  assign new_n1490_ = p_7 & p_3;
  assign new_n1491_ = ~new_n1489_ & ~new_n1490_;
  assign new_n1492_ = p_2 & ~new_n1491_;
  assign new_n1493_ = ~p_2 & n_37;
  assign new_n1494_ = ~new_n1492_ & ~new_n1493_;
  assign p_127 = ~p_1 & ~new_n1494_;
  assign new_n1496_ = new_n738_ & ~new_n903_;
  assign new_n1497_ = new_n733_ & ~new_n737_;
  assign new_n1498_ = new_n903_ & new_n1497_;
  assign new_n1499_ = ~new_n733_ & new_n737_;
  assign new_n1500_ = new_n903_ & new_n1499_;
  assign new_n1501_ = ~new_n733_ & ~new_n737_;
  assign new_n1502_ = ~new_n903_ & new_n1501_;
  assign new_n1503_ = ~new_n1496_ & ~new_n1498_;
  assign new_n1504_ = ~new_n1500_ & ~new_n1502_;
  assign new_n1505_ = new_n1503_ & new_n1504_;
  assign new_n1506_ = ~p_3 & ~new_n1505_;
  assign new_n1507_ = p_16 & p_3;
  assign new_n1508_ = ~new_n1506_ & ~new_n1507_;
  assign new_n1509_ = p_2 & ~new_n1508_;
  assign new_n1510_ = ~p_2 & n_46;
  assign new_n1511_ = ~new_n1509_ & ~new_n1510_;
  assign p_136 = ~p_1 & ~new_n1511_;
  assign new_n1513_ = new_n999_ & ~new_n1055_;
  assign new_n1514_ = new_n994_ & ~new_n998_;
  assign new_n1515_ = new_n1055_ & new_n1514_;
  assign new_n1516_ = ~new_n994_ & new_n998_;
  assign new_n1517_ = new_n1055_ & new_n1516_;
  assign new_n1518_ = ~new_n994_ & ~new_n998_;
  assign new_n1519_ = ~new_n1055_ & new_n1518_;
  assign new_n1520_ = ~new_n1513_ & ~new_n1515_;
  assign new_n1521_ = ~new_n1517_ & ~new_n1519_;
  assign new_n1522_ = new_n1520_ & new_n1521_;
  assign new_n1523_ = ~p_3 & ~new_n1522_;
  assign new_n1524_ = p_25 & p_3;
  assign new_n1525_ = ~new_n1523_ & ~new_n1524_;
  assign new_n1526_ = p_2 & ~new_n1525_;
  assign new_n1527_ = ~p_2 & n_55;
  assign new_n1528_ = ~new_n1526_ & ~new_n1527_;
  assign p_145 = ~p_1 & ~new_n1528_;
  assign new_n1530_ = new_n801_ & ~new_n875_;
  assign new_n1531_ = new_n796_ & ~new_n800_;
  assign new_n1532_ = new_n875_ & new_n1531_;
  assign new_n1533_ = ~new_n796_ & new_n800_;
  assign new_n1534_ = new_n875_ & new_n1533_;
  assign new_n1535_ = ~new_n796_ & ~new_n800_;
  assign new_n1536_ = ~new_n875_ & new_n1535_;
  assign new_n1537_ = ~new_n1530_ & ~new_n1532_;
  assign new_n1538_ = ~new_n1534_ & ~new_n1536_;
  assign new_n1539_ = new_n1537_ & new_n1538_;
  assign new_n1540_ = ~p_3 & ~new_n1539_;
  assign new_n1541_ = p_9 & p_3;
  assign new_n1542_ = ~new_n1540_ & ~new_n1541_;
  assign new_n1543_ = p_2 & ~new_n1542_;
  assign new_n1544_ = ~p_2 & n_39;
  assign new_n1545_ = ~new_n1543_ & ~new_n1544_;
  assign p_129 = ~p_1 & ~new_n1545_;
  assign new_n1547_ = new_n711_ & ~new_n915_;
  assign new_n1548_ = new_n706_ & ~new_n710_;
  assign new_n1549_ = new_n915_ & new_n1548_;
  assign new_n1550_ = ~new_n706_ & new_n710_;
  assign new_n1551_ = new_n915_ & new_n1550_;
  assign new_n1552_ = ~new_n706_ & ~new_n710_;
  assign new_n1553_ = ~new_n915_ & new_n1552_;
  assign new_n1554_ = ~new_n1547_ & ~new_n1549_;
  assign new_n1555_ = ~new_n1551_ & ~new_n1553_;
  assign new_n1556_ = new_n1554_ & new_n1555_;
  assign new_n1557_ = ~p_3 & ~new_n1556_;
  assign new_n1558_ = p_19 & p_3;
  assign new_n1559_ = ~new_n1557_ & ~new_n1558_;
  assign new_n1560_ = p_2 & ~new_n1559_;
  assign new_n1561_ = ~p_2 & n_49;
  assign new_n1562_ = ~new_n1560_ & ~new_n1561_;
  assign p_139 = ~p_1 & ~new_n1562_;
  assign new_n1564_ = new_n963_ & ~new_n1071_;
  assign new_n1565_ = new_n958_ & ~new_n962_;
  assign new_n1566_ = new_n1071_ & new_n1565_;
  assign new_n1567_ = ~new_n958_ & new_n962_;
  assign new_n1568_ = new_n1071_ & new_n1567_;
  assign new_n1569_ = ~new_n958_ & ~new_n962_;
  assign new_n1570_ = ~new_n1071_ & new_n1569_;
  assign new_n1571_ = ~new_n1564_ & ~new_n1566_;
  assign new_n1572_ = ~new_n1568_ & ~new_n1570_;
  assign new_n1573_ = new_n1571_ & new_n1572_;
  assign new_n1574_ = ~p_3 & ~new_n1573_;
  assign new_n1575_ = p_29 & p_3;
  assign new_n1576_ = ~new_n1574_ & ~new_n1575_;
  assign new_n1577_ = p_2 & ~new_n1576_;
  assign new_n1578_ = ~p_2 & n_59;
  assign new_n1579_ = ~new_n1577_ & ~new_n1578_;
  assign p_149 = ~p_1 & ~new_n1579_;
  assign new_n1581_ = p_13 & p_2;
  assign n130 = ~p_1 & new_n1581_;
  assign new_n1583_ = p_9 & p_2;
  assign n135 = ~p_1 & new_n1583_;
  assign new_n1585_ = p_10 & p_2;
  assign n140 = ~p_1 & new_n1585_;
  assign new_n1587_ = p_11 & p_2;
  assign n145 = ~p_1 & new_n1587_;
  assign new_n1589_ = p_12 & p_2;
  assign n150 = ~p_1 & new_n1589_;
  assign new_n1591_ = p_5 & p_2;
  assign n155 = ~p_1 & new_n1591_;
  assign new_n1593_ = p_6 & p_2;
  assign n160 = ~p_1 & new_n1593_;
  assign new_n1595_ = p_7 & p_2;
  assign n165 = ~p_1 & new_n1595_;
  assign new_n1597_ = p_8 & p_2;
  assign n170 = ~p_1 & new_n1597_;
  assign new_n1599_ = ~p_3 & new_n1012_;
  assign new_n1600_ = ~p_3 & ~new_n1599_;
  assign new_n1601_ = p_2 & ~new_n1600_;
  assign new_n1602_ = p_2 & ~new_n1601_;
  assign new_n1603_ = ~p_1 & ~new_n1602_;
  assign n175 = p_1 | new_n1603_;
  assign new_n1605_ = ~p_3 & new_n845_;
  assign new_n1606_ = p_2 & new_n1605_;
  assign n180 = ~p_1 & new_n1606_;
  assign new_n1608_ = ~p_3 & new_n746_;
  assign new_n1609_ = p_2 & new_n1608_;
  assign n185 = ~p_1 & new_n1609_;
  assign new_n1611_ = ~p_3 & new_n989_;
  assign new_n1612_ = p_2 & new_n1611_;
  assign n190 = ~p_1 & new_n1612_;
  assign new_n1614_ = ~p_3 & new_n1003_;
  assign new_n1615_ = ~p_3 & ~new_n1614_;
  assign new_n1616_ = p_2 & ~new_n1615_;
  assign new_n1617_ = p_2 & ~new_n1616_;
  assign new_n1618_ = ~p_1 & ~new_n1617_;
  assign n195 = p_1 | new_n1618_;
  assign new_n1620_ = ~p_3 & new_n854_;
  assign new_n1621_ = p_2 & new_n1620_;
  assign n200 = ~p_1 & new_n1621_;
  assign new_n1623_ = ~p_3 & new_n737_;
  assign new_n1624_ = p_2 & new_n1623_;
  assign n205 = ~p_1 & new_n1624_;
  assign new_n1626_ = ~p_3 & new_n998_;
  assign new_n1627_ = p_2 & new_n1626_;
  assign n210 = ~p_1 & new_n1627_;
  assign new_n1629_ = ~p_3 & new_n994_;
  assign new_n1630_ = ~p_3 & ~new_n1629_;
  assign new_n1631_ = p_2 & ~new_n1630_;
  assign new_n1632_ = p_2 & ~new_n1631_;
  assign new_n1633_ = ~p_1 & ~new_n1632_;
  assign n215 = p_1 | new_n1633_;
  assign new_n1635_ = ~p_3 & new_n827_;
  assign new_n1636_ = p_2 & new_n1635_;
  assign n220 = ~p_1 & new_n1636_;
  assign new_n1638_ = ~p_3 & new_n764_;
  assign new_n1639_ = p_2 & new_n1638_;
  assign n225 = ~p_1 & new_n1639_;
  assign new_n1641_ = ~p_3 & new_n1007_;
  assign new_n1642_ = p_2 & new_n1641_;
  assign n230 = ~p_1 & new_n1642_;
  assign new_n1644_ = p_4 & p_2;
  assign n235 = ~p_1 & new_n1644_;
  assign new_n1646_ = ~p_3 & new_n985_;
  assign new_n1647_ = ~p_3 & ~new_n1646_;
  assign new_n1648_ = p_2 & ~new_n1647_;
  assign new_n1649_ = p_2 & ~new_n1648_;
  assign new_n1650_ = ~p_1 & ~new_n1649_;
  assign n240 = p_1 | new_n1650_;
  assign new_n1652_ = ~p_3 & new_n836_;
  assign new_n1653_ = p_2 & new_n1652_;
  assign n245 = ~p_1 & new_n1653_;
  assign new_n1655_ = ~p_3 & new_n755_;
  assign new_n1656_ = p_2 & new_n1655_;
  assign n250 = ~p_1 & new_n1656_;
  assign new_n1658_ = ~p_3 & new_n1016_;
  assign new_n1659_ = p_2 & new_n1658_;
  assign n255 = ~p_1 & new_n1659_;
  assign new_n1661_ = p_14 & p_2;
  assign n260 = ~p_1 & new_n1661_;
  assign new_n1663_ = p_25 & p_2;
  assign n265 = ~p_1 & new_n1663_;
  assign new_n1665_ = ~p_3 & new_n832_;
  assign new_n1666_ = ~p_3 & ~new_n1665_;
  assign new_n1667_ = p_2 & ~new_n1666_;
  assign new_n1668_ = p_2 & ~new_n1667_;
  assign new_n1669_ = ~p_1 & ~new_n1668_;
  assign n270 = p_1 | new_n1669_;
  assign new_n1671_ = ~p_3 & new_n733_;
  assign new_n1672_ = ~p_3 & ~new_n1671_;
  assign new_n1673_ = p_2 & ~new_n1672_;
  assign new_n1674_ = p_2 & ~new_n1673_;
  assign new_n1675_ = ~p_1 & ~new_n1674_;
  assign n275 = p_1 | new_n1675_;
  assign new_n1677_ = p_15 & p_2;
  assign n280 = ~p_1 & new_n1677_;
  assign new_n1679_ = p_24 & p_2;
  assign n285 = ~p_1 & new_n1679_;
  assign new_n1681_ = ~p_3 & new_n823_;
  assign new_n1682_ = ~p_3 & ~new_n1681_;
  assign new_n1683_ = p_2 & ~new_n1682_;
  assign new_n1684_ = p_2 & ~new_n1683_;
  assign new_n1685_ = ~p_1 & ~new_n1684_;
  assign n290 = p_1 | new_n1685_;
  assign new_n1687_ = ~p_3 & new_n742_;
  assign new_n1688_ = ~p_3 & ~new_n1687_;
  assign new_n1689_ = p_2 & ~new_n1688_;
  assign new_n1690_ = p_2 & ~new_n1689_;
  assign new_n1691_ = ~p_1 & ~new_n1690_;
  assign n295 = p_1 | new_n1691_;
  assign new_n1693_ = p_16 & p_2;
  assign n300 = ~p_1 & new_n1693_;
  assign new_n1695_ = p_27 & p_2;
  assign n305 = ~p_1 & new_n1695_;
  assign new_n1697_ = ~p_3 & new_n850_;
  assign new_n1698_ = ~p_3 & ~new_n1697_;
  assign new_n1699_ = p_2 & ~new_n1698_;
  assign new_n1700_ = p_2 & ~new_n1699_;
  assign new_n1701_ = ~p_1 & ~new_n1700_;
  assign n310 = p_1 | new_n1701_;
  assign new_n1703_ = ~p_3 & new_n751_;
  assign new_n1704_ = ~p_3 & ~new_n1703_;
  assign new_n1705_ = p_2 & ~new_n1704_;
  assign new_n1706_ = p_2 & ~new_n1705_;
  assign new_n1707_ = ~p_1 & ~new_n1706_;
  assign n315 = p_1 | new_n1707_;
  assign new_n1709_ = p_17 & p_2;
  assign n320 = ~p_1 & new_n1709_;
  assign new_n1711_ = p_26 & p_2;
  assign n325 = ~p_1 & new_n1711_;
  assign new_n1713_ = ~p_3 & new_n841_;
  assign new_n1714_ = ~p_3 & ~new_n1713_;
  assign new_n1715_ = p_2 & ~new_n1714_;
  assign new_n1716_ = p_2 & ~new_n1715_;
  assign new_n1717_ = ~p_1 & ~new_n1716_;
  assign n330 = p_1 | new_n1717_;
  assign new_n1719_ = ~p_3 & new_n760_;
  assign new_n1720_ = ~p_3 & ~new_n1719_;
  assign new_n1721_ = p_2 & ~new_n1720_;
  assign new_n1722_ = p_2 & ~new_n1721_;
  assign new_n1723_ = ~p_1 & ~new_n1722_;
  assign n335 = p_1 | new_n1723_;
  assign new_n1725_ = p_18 & p_2;
  assign n340 = ~p_1 & new_n1725_;
  assign new_n1727_ = p_29 & p_2;
  assign n345 = ~p_1 & new_n1727_;
  assign new_n1729_ = ~p_3 & new_n796_;
  assign new_n1730_ = ~p_3 & ~new_n1729_;
  assign new_n1731_ = p_2 & ~new_n1730_;
  assign new_n1732_ = p_2 & ~new_n1731_;
  assign new_n1733_ = ~p_1 & ~new_n1732_;
  assign n350 = p_1 | new_n1733_;
  assign new_n1735_ = ~p_3 & new_n702_;
  assign new_n1736_ = ~p_3 & ~new_n1735_;
  assign new_n1737_ = p_2 & ~new_n1736_;
  assign new_n1738_ = p_2 & ~new_n1737_;
  assign new_n1739_ = ~p_1 & ~new_n1738_;
  assign n355 = p_1 | new_n1739_;
  assign new_n1741_ = ~p_3 & new_n945_;
  assign new_n1742_ = ~p_3 & ~new_n1741_;
  assign new_n1743_ = p_2 & ~new_n1742_;
  assign new_n1744_ = p_2 & ~new_n1743_;
  assign new_n1745_ = ~p_1 & ~new_n1744_;
  assign n360 = p_1 | new_n1745_;
  assign new_n1747_ = ~p_3 & new_n773_;
  assign new_n1748_ = p_2 & new_n1747_;
  assign n365 = ~p_1 & new_n1748_;
  assign new_n1750_ = p_19 & p_2;
  assign n370 = ~p_1 & new_n1750_;
  assign new_n1752_ = p_28 & p_2;
  assign n375 = ~p_1 & new_n1752_;
  assign new_n1754_ = ~p_3 & new_n787_;
  assign new_n1755_ = ~p_3 & ~new_n1754_;
  assign new_n1756_ = p_2 & ~new_n1755_;
  assign new_n1757_ = p_2 & ~new_n1756_;
  assign new_n1758_ = ~p_1 & ~new_n1757_;
  assign n380 = p_1 | new_n1758_;
  assign new_n1760_ = ~p_3 & new_n706_;
  assign new_n1761_ = ~p_3 & ~new_n1760_;
  assign new_n1762_ = p_2 & ~new_n1761_;
  assign new_n1763_ = p_2 & ~new_n1762_;
  assign new_n1764_ = ~p_1 & ~new_n1763_;
  assign n385 = p_1 | new_n1764_;
  assign new_n1766_ = ~p_3 & new_n1122_;
  assign new_n1767_ = ~p_3 & ~new_n1766_;
  assign new_n1768_ = p_2 & ~new_n1767_;
  assign new_n1769_ = p_2 & ~new_n1768_;
  assign new_n1770_ = ~p_1 & ~new_n1769_;
  assign n390 = p_1 | new_n1770_;
  assign new_n1772_ = ~p_3 & new_n782_;
  assign new_n1773_ = p_2 & new_n1772_;
  assign n395 = ~p_1 & new_n1773_;
  assign new_n1775_ = p_20 & p_2;
  assign n400 = ~p_1 & new_n1775_;
  assign new_n1777_ = p_31 & p_2;
  assign n405 = ~p_1 & new_n1777_;
  assign new_n1779_ = ~p_3 & new_n814_;
  assign new_n1780_ = ~p_3 & ~new_n1779_;
  assign new_n1781_ = p_2 & ~new_n1780_;
  assign new_n1782_ = p_2 & ~new_n1781_;
  assign new_n1783_ = ~p_1 & ~new_n1782_;
  assign n410 = p_1 | new_n1783_;
  assign new_n1785_ = ~p_3 & new_n715_;
  assign new_n1786_ = ~p_3 & ~new_n1785_;
  assign new_n1787_ = p_2 & ~new_n1786_;
  assign new_n1788_ = p_2 & ~new_n1787_;
  assign new_n1789_ = ~p_1 & ~new_n1788_;
  assign n415 = p_1 | new_n1789_;
  assign new_n1791_ = ~p_3 & new_n1034_;
  assign new_n1792_ = p_2 & new_n1791_;
  assign n420 = ~p_1 & new_n1792_;
  assign new_n1794_ = ~p_3 & new_n1118_;
  assign new_n1795_ = p_2 & new_n1794_;
  assign n425 = ~p_1 & new_n1795_;
  assign new_n1797_ = p_21 & p_2;
  assign n430 = ~p_1 & new_n1797_;
  assign new_n1799_ = p_30 & p_2;
  assign n435 = ~p_1 & new_n1799_;
  assign new_n1801_ = ~p_3 & new_n805_;
  assign new_n1802_ = ~p_3 & ~new_n1801_;
  assign new_n1803_ = p_2 & ~new_n1802_;
  assign new_n1804_ = p_2 & ~new_n1803_;
  assign new_n1805_ = ~p_1 & ~new_n1804_;
  assign n440 = p_1 | new_n1805_;
  assign new_n1807_ = ~p_3 & new_n724_;
  assign new_n1808_ = ~p_3 & ~new_n1807_;
  assign new_n1809_ = p_2 & ~new_n1808_;
  assign new_n1810_ = p_2 & ~new_n1809_;
  assign new_n1811_ = ~p_1 & ~new_n1810_;
  assign n445 = p_1 | new_n1811_;
  assign new_n1813_ = ~p_3 & new_n1025_;
  assign new_n1814_ = p_2 & new_n1813_;
  assign n450 = ~p_1 & new_n1814_;
  assign new_n1816_ = ~p_3 & new_n941_;
  assign new_n1817_ = p_2 & new_n1816_;
  assign n455 = ~p_1 & new_n1817_;
  assign new_n1819_ = p_22 & p_2;
  assign n460 = ~p_1 & new_n1819_;
  assign new_n1821_ = p_33 & p_2;
  assign n465 = ~p_1 & new_n1821_;
  assign new_n1823_ = ~p_3 & new_n976_;
  assign new_n1824_ = ~p_3 & ~new_n1823_;
  assign new_n1825_ = p_2 & ~new_n1824_;
  assign new_n1826_ = p_2 & ~new_n1825_;
  assign new_n1827_ = ~p_1 & ~new_n1826_;
  assign n470 = p_1 | new_n1827_;
  assign new_n1829_ = ~p_3 & new_n809_;
  assign new_n1830_ = p_2 & new_n1829_;
  assign n475 = ~p_1 & new_n1830_;
  assign new_n1832_ = ~p_3 & new_n710_;
  assign new_n1833_ = p_2 & new_n1832_;
  assign n480 = ~p_1 & new_n1833_;
  assign new_n1835_ = ~p_3 & new_n953_;
  assign new_n1836_ = p_2 & new_n1835_;
  assign n485 = ~p_1 & new_n1836_;
  assign new_n1838_ = p_23 & p_2;
  assign n490 = ~p_1 & new_n1838_;
  assign new_n1840_ = p_32 & p_2;
  assign n495 = ~p_1 & new_n1840_;
  assign new_n1842_ = ~p_3 & new_n967_;
  assign new_n1843_ = ~p_3 & ~new_n1842_;
  assign new_n1844_ = p_2 & ~new_n1843_;
  assign new_n1845_ = p_2 & ~new_n1844_;
  assign new_n1846_ = ~p_1 & ~new_n1845_;
  assign n500 = p_1 | new_n1846_;
  assign new_n1848_ = ~p_3 & new_n818_;
  assign new_n1849_ = p_2 & new_n1848_;
  assign n505 = ~p_1 & new_n1849_;
  assign new_n1851_ = ~p_3 & new_n519_;
  assign new_n1852_ = p_2 & new_n1851_;
  assign n510 = ~p_1 & new_n1852_;
  assign new_n1854_ = ~p_3 & new_n962_;
  assign new_n1855_ = p_2 & new_n1854_;
  assign n515 = ~p_1 & new_n1855_;
  assign new_n1857_ = ~p_3 & new_n778_;
  assign new_n1858_ = ~p_3 & ~new_n1857_;
  assign new_n1859_ = p_2 & ~new_n1858_;
  assign new_n1860_ = p_2 & ~new_n1859_;
  assign new_n1861_ = ~p_1 & ~new_n1860_;
  assign n520 = p_1 | new_n1861_;
  assign new_n1863_ = ~p_3 & new_n1021_;
  assign new_n1864_ = ~p_3 & ~new_n1863_;
  assign new_n1865_ = p_2 & ~new_n1864_;
  assign new_n1866_ = p_2 & ~new_n1865_;
  assign new_n1867_ = ~p_1 & ~new_n1866_;
  assign n525 = p_1 | new_n1867_;
  assign new_n1869_ = ~p_3 & new_n958_;
  assign new_n1870_ = ~p_3 & ~new_n1869_;
  assign new_n1871_ = p_2 & ~new_n1870_;
  assign new_n1872_ = p_2 & ~new_n1871_;
  assign new_n1873_ = ~p_1 & ~new_n1872_;
  assign n530 = p_1 | new_n1873_;
  assign new_n1875_ = ~p_3 & new_n791_;
  assign new_n1876_ = p_2 & new_n1875_;
  assign n535 = ~p_1 & new_n1876_;
  assign new_n1878_ = ~p_3 & new_n728_;
  assign new_n1879_ = p_2 & new_n1878_;
  assign n540 = ~p_1 & new_n1879_;
  assign new_n1881_ = ~p_3 & new_n971_;
  assign new_n1882_ = p_2 & new_n1881_;
  assign n545 = ~p_1 & new_n1882_;
  assign new_n1884_ = ~p_3 & new_n769_;
  assign new_n1885_ = ~p_3 & ~new_n1884_;
  assign new_n1886_ = p_2 & ~new_n1885_;
  assign new_n1887_ = p_2 & ~new_n1886_;
  assign new_n1888_ = ~p_1 & ~new_n1887_;
  assign n550 = p_1 | new_n1888_;
  assign new_n1890_ = ~p_3 & new_n1030_;
  assign new_n1891_ = ~p_3 & ~new_n1890_;
  assign new_n1892_ = p_2 & ~new_n1891_;
  assign new_n1893_ = p_2 & ~new_n1892_;
  assign new_n1894_ = ~p_1 & ~new_n1893_;
  assign n555 = p_1 | new_n1894_;
  assign new_n1896_ = ~p_3 & new_n949_;
  assign new_n1897_ = ~p_3 & ~new_n1896_;
  assign new_n1898_ = p_2 & ~new_n1897_;
  assign new_n1899_ = p_2 & ~new_n1898_;
  assign new_n1900_ = ~p_1 & ~new_n1899_;
  assign n560 = p_1 | new_n1900_;
  assign new_n1902_ = ~p_3 & new_n800_;
  assign new_n1903_ = p_2 & new_n1902_;
  assign n565 = ~p_1 & new_n1903_;
  assign new_n1905_ = ~p_3 & new_n719_;
  assign new_n1906_ = p_2 & new_n1905_;
  assign n570 = ~p_1 & new_n1906_;
  assign new_n1908_ = ~p_3 & new_n980_;
  assign new_n1909_ = p_2 & new_n1908_;
  assign n575 = ~p_1 & new_n1909_;
  always @ (posedge clock) begin
    n_43 <= n130;
    n_39 <= n135;
    n_40 <= n140;
    n_41 <= n145;
    n_42 <= n150;
    n_35 <= n155;
    n_36 <= n160;
    n_37 <= n165;
    n_38 <= n170;
    n_84 <= n175;
    n_95 <= n180;
    n_106 <= n185;
    n_117 <= n190;
    n_85 <= n195;
    n_94 <= n200;
    n_107 <= n205;
    n_116 <= n210;
    n_86 <= n215;
    n_97 <= n220;
    n_104 <= n225;
    n_115 <= n230;
    n_34 <= n235;
    n_87 <= n240;
    n_96 <= n245;
    n_105 <= n250;
    n_114 <= n255;
    n_44 <= n260;
    n_55 <= n265;
    n_66 <= n270;
    n_77 <= n275;
    n_45 <= n280;
    n_54 <= n285;
    n_67 <= n290;
    n_76 <= n295;
    n_46 <= n300;
    n_57 <= n305;
    n_64 <= n310;
    n_75 <= n315;
    n_47 <= n320;
    n_56 <= n325;
    n_65 <= n330;
    n_74 <= n335;
    n_48 <= n340;
    n_59 <= n345;
    n_70 <= n350;
    n_81 <= n355;
    n_92 <= n360;
    n_103 <= n365;
    n_49 <= n370;
    n_58 <= n375;
    n_71 <= n380;
    n_80 <= n385;
    n_93 <= n390;
    n_102 <= n395;
    n_50 <= n400;
    n_61 <= n405;
    n_68 <= n410;
    n_79 <= n415;
    n_112 <= n420;
    n_123 <= n425;
    n_51 <= n430;
    n_60 <= n435;
    n_69 <= n440;
    n_78 <= n445;
    n_113 <= n450;
    n_122 <= n455;
    n_52 <= n460;
    n_63 <= n465;
    n_88 <= n470;
    n_99 <= n475;
    n_110 <= n480;
    n_121 <= n485;
    n_53 <= n490;
    n_62 <= n495;
    n_89 <= n500;
    n_98 <= n505;
    n_111 <= n510;
    n_120 <= n515;
    n_72 <= n520;
    n_83 <= n525;
    n_90 <= n530;
    n_101 <= n535;
    n_108 <= n540;
    n_119 <= n545;
    n_73 <= n550;
    n_82 <= n555;
    n_91 <= n560;
    n_100 <= n565;
    n_109 <= n570;
    n_118 <= n575;
  end
endmodule

