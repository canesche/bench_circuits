module top ( 
    pp, pa0, pq, pr, ps, pt, pu, pv, pw, px, py, pz, pa, pb, pc, pd, pe,
    pf, pg, ph, pj, pk, pl, pm, pn, po,
    pb0, pc0, pd0, pe0, pf0, pg0, ph0, pi0, pj0, pk0, pl0, pm0, pn0, po0,
    pp0, pq0, pr0, ps0, pt0  );
  input  pp, pa0, pq, pr, ps, pt, pu, pv, pw, px, py, pz, pa, pb, pc, pd,
    pe, pf, pg, ph, pj, pk, pl, pm, pn, po;
  output pb0, pc0, pd0, pe0, pf0, pg0, ph0, pi0, pj0, pk0, pl0, pm0, pn0, po0,
    pp0, pq0, pr0, ps0, pt0;
  wire new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_,
    new_n54_, new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_,
    new_n61_, new_n62_, new_n63_, new_n64_, new_n66_, new_n67_, new_n68_,
    new_n69_, new_n70_, new_n71_, new_n73_, new_n74_, new_n75_, new_n76_,
    new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n83_,
    new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_,
    new_n91_, new_n92_, new_n93_, new_n98_, new_n99_, new_n101_, new_n102_,
    new_n104_, new_n105_, new_n106_, new_n107_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n120_, new_n121_, new_n122_, new_n123_,
    new_n124_, new_n125_, new_n126_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_,
    new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_;
  assign pb0 = ~pr & pj;
  assign new_n47_ = pt & ~pv;
  assign new_n48_ = pu & ~pv;
  assign new_n49_ = ps & ~pv;
  assign new_n50_ = ~new_n47_ & ~new_n48_;
  assign new_n51_ = ~new_n49_ & new_n50_;
  assign new_n52_ = pw & new_n51_;
  assign new_n53_ = px & new_n52_;
  assign new_n54_ = ~py & ~new_n53_;
  assign new_n55_ = ~pa0 & new_n54_;
  assign new_n56_ = ~pf & ~ph;
  assign new_n57_ = pa0 & new_n56_;
  assign new_n58_ = ~pe & ~ph;
  assign new_n59_ = pa0 & new_n58_;
  assign new_n60_ = pz & new_n56_;
  assign new_n61_ = pz & new_n58_;
  assign new_n62_ = ~new_n57_ & ~new_n59_;
  assign new_n63_ = ~new_n60_ & ~new_n61_;
  assign new_n64_ = new_n62_ & new_n63_;
  assign pc0 = new_n55_ | new_n64_;
  assign new_n66_ = px & pz;
  assign new_n67_ = new_n51_ & new_n66_;
  assign new_n68_ = pw & new_n67_;
  assign new_n69_ = ~pa0 & ~pz;
  assign new_n70_ = ~pa0 & ~py;
  assign new_n71_ = ~new_n69_ & ~new_n70_;
  assign pe0 = ~new_n68_ & ~new_n71_;
  assign new_n73_ = pc & ~pm;
  assign new_n74_ = pd & ~pn;
  assign new_n75_ = ~pc & pm;
  assign new_n76_ = ~pd & pn;
  assign new_n77_ = ~pb & pl;
  assign new_n78_ = ~new_n75_ & ~new_n76_;
  assign new_n79_ = ~new_n77_ & new_n78_;
  assign new_n80_ = pa & new_n79_;
  assign new_n81_ = ~pk & new_n79_;
  assign new_n82_ = ~new_n80_ & ~new_n81_;
  assign new_n83_ = ~new_n73_ & ~new_n74_;
  assign new_n84_ = ~new_n82_ & new_n83_;
  assign new_n85_ = ~pb & new_n84_;
  assign new_n86_ = ~pa & new_n85_;
  assign new_n87_ = pl & new_n84_;
  assign new_n88_ = ~pa & new_n87_;
  assign new_n89_ = pk & new_n85_;
  assign new_n90_ = pk & new_n87_;
  assign new_n91_ = ~new_n86_ & ~new_n88_;
  assign new_n92_ = ~new_n89_ & ~new_n90_;
  assign new_n93_ = new_n91_ & new_n92_;
  assign pf0 = ~pj & new_n93_;
  assign pg0 = ~pj & ~po;
  assign ph0 = pp & ~pj;
  assign pi0 = ~pg | pj;
  assign new_n98_ = pe & pf;
  assign new_n99_ = ~ph & new_n98_;
  assign pk0 = ~pq & new_n99_;
  assign new_n101_ = ~pq & ~new_n98_;
  assign new_n102_ = ~ph & new_n101_;
  assign pl0 = ~ps & new_n102_;
  assign new_n104_ = ~pt & new_n102_;
  assign new_n105_ = ps & new_n104_;
  assign new_n106_ = pt & new_n102_;
  assign new_n107_ = ~ps & new_n106_;
  assign pm0 = new_n105_ | new_n107_;
  assign new_n109_ = ps & pt;
  assign new_n110_ = pu & new_n109_;
  assign new_n111_ = ~pq & ~ph;
  assign new_n112_ = ~pf & new_n111_;
  assign new_n113_ = ~pe & new_n111_;
  assign new_n114_ = ~new_n112_ & ~new_n113_;
  assign new_n115_ = ~new_n110_ & ~new_n114_;
  assign new_n116_ = pt & new_n115_;
  assign new_n117_ = ps & new_n116_;
  assign new_n118_ = pu & new_n115_;
  assign pn0 = new_n117_ | new_n118_;
  assign new_n120_ = ~pv & new_n110_;
  assign new_n121_ = ~pq & ~new_n120_;
  assign new_n122_ = ~pe & new_n121_;
  assign new_n123_ = ~pf & new_n121_;
  assign new_n124_ = ~new_n122_ & ~new_n123_;
  assign new_n125_ = pv & ~new_n110_;
  assign new_n126_ = ~new_n124_ & ~new_n125_;
  assign po0 = ph | ~new_n126_;
  assign new_n128_ = ~pw & new_n120_;
  assign new_n129_ = ~pq & ~new_n128_;
  assign new_n130_ = ~pe & new_n129_;
  assign new_n131_ = ~pf & new_n129_;
  assign new_n132_ = ~new_n130_ & ~new_n131_;
  assign new_n133_ = ps & new_n48_;
  assign new_n134_ = pt & new_n133_;
  assign new_n135_ = pw & ~new_n134_;
  assign new_n136_ = ~new_n132_ & ~new_n135_;
  assign pp0 = ph | ~new_n136_;
  assign new_n138_ = ~pw & new_n134_;
  assign new_n139_ = ~px & new_n138_;
  assign new_n140_ = ~pq & ~new_n139_;
  assign new_n141_ = ~pe & new_n140_;
  assign new_n142_ = ~pf & new_n140_;
  assign new_n143_ = ~new_n141_ & ~new_n142_;
  assign new_n144_ = ~pw & new_n48_;
  assign new_n145_ = ps & new_n144_;
  assign new_n146_ = pt & new_n145_;
  assign new_n147_ = px & ~new_n146_;
  assign new_n148_ = ~new_n143_ & ~new_n147_;
  assign pq0 = ph | ~new_n148_;
  assign new_n150_ = ~px & new_n146_;
  assign new_n151_ = ~py & new_n150_;
  assign new_n152_ = ~pq & ~new_n151_;
  assign new_n153_ = ~pe & new_n152_;
  assign new_n154_ = ~pf & new_n152_;
  assign new_n155_ = ~new_n153_ & ~new_n154_;
  assign new_n156_ = pt & pu;
  assign new_n157_ = ~pv & ~pw;
  assign new_n158_ = ~px & new_n157_;
  assign new_n159_ = new_n156_ & new_n158_;
  assign new_n160_ = ps & new_n159_;
  assign new_n161_ = py & ~new_n160_;
  assign new_n162_ = ~new_n155_ & ~new_n161_;
  assign pr0 = ph | ~new_n162_;
  assign new_n164_ = ~py & new_n160_;
  assign new_n165_ = ~pz & new_n164_;
  assign new_n166_ = ~pq & ~new_n165_;
  assign new_n167_ = ~pe & new_n166_;
  assign new_n168_ = ~pf & new_n166_;
  assign new_n169_ = ~new_n167_ & ~new_n168_;
  assign new_n170_ = ~pv & new_n156_;
  assign new_n171_ = ~pw & ~px;
  assign new_n172_ = ~py & new_n171_;
  assign new_n173_ = new_n170_ & new_n172_;
  assign new_n174_ = ps & new_n173_;
  assign new_n175_ = pz & ~new_n174_;
  assign new_n176_ = ~new_n169_ & ~new_n175_;
  assign ps0 = ph | ~new_n176_;
  assign new_n178_ = ~pz & new_n174_;
  assign new_n179_ = ~pa0 & new_n178_;
  assign new_n180_ = ~pq & ~new_n179_;
  assign new_n181_ = ~pe & new_n180_;
  assign new_n182_ = ~pf & new_n180_;
  assign new_n183_ = ~new_n181_ & ~new_n182_;
  assign new_n184_ = ~px & ~py;
  assign new_n185_ = ~pz & new_n184_;
  assign new_n186_ = new_n144_ & new_n185_;
  assign new_n187_ = new_n109_ & new_n186_;
  assign new_n188_ = pa0 & ~new_n187_;
  assign new_n189_ = ~new_n183_ & ~new_n188_;
  assign pt0 = ph | ~new_n189_;
  assign pj0 = ~pe0;
  assign pd0 = pr;
endmodule

