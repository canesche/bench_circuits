module top ( 
    pv16_9_, pv40_15_, pv88_6_, pv28_10_, pv88_7_, pv109_1_, pv118_3_,
    pv2_0_, pv40_13_, pv52_10_, pv109_2_, pv128_3_, pv2_1_, pv40_14_,
    pv52_11_, pv88_9_, pv109_3_, pv16_5_, pv40_11_, pv76_3_, pv88_2_,
    pv88_15_, pv100_14_, pv128_1_, pv16_13_, pv52_13_, pv76_2_, pv88_3_,
    pv100_13_, pv128_2_, pv16_7_, pv16_14_, pv52_14_, pv76_1_, pv88_13_,
    pv118_2_, pv16_6_, pv16_15_, pv40_10_, pv52_15_, pv88_5_, pv88_14_,
    pv100_15_, pv118_1_, pv128_0_, pv4_0_, pv52_9_, pv88_11_, pv100_3_,
    pv100_10_, pv121_2_, pv132_0_, pv4_1_, pv28_9_, pv64_1_, pv121_3_,
    pv16_10_, pv28_6_, pv100_5_, pv16_11_, pv28_7_, pv88_10_, pv100_6_,
    pv100_11_, pv121_1_, pv76_14_, pv28_5_, pv64_5_, pv76_15_, pv28_2_,
    pv64_2_, pv100_1_, pv28_3_, pv64_3_, pv100_2_, pv52_1_, pv76_10_,
    pv103_2_, pv124_1_, pv28_1_, pv64_9_, pv76_11_, pv103_3_, pv124_2_,
    pv52_3_, pv64_6_, pv64_15_, pv52_2_, pv64_7_, pv76_13_, pv52_5_,
    pv100_7_, pv112_2_, pv112_1_, pv132_3_, pv133_0_, pv52_7_, pv100_9_,
    pv132_2_, pv40_1_, pv52_6_, pv103_1_, pv112_3_, pv132_1_, pv16_1_,
    pv40_2_, pv76_7_, pv106_1_, pv40_3_, pv64_10_, pv76_6_, pv106_2_,
    pv16_3_, pv28_15_, pv76_5_, pv106_3_, pv16_2_, pv40_5_, pv88_1_,
    pv28_13_, pv40_6_, pv64_13_, pv115_1_, pv28_14_, pv40_7_, pv64_14_,
    pv28_11_, pv64_11_, pv76_9_, pv115_3_, pv124_3_, pv40_9_, pv115_2_,
    pv167_11_, pv199_9_, pv167_12_, pv199_8_, pv167_13_, pv167_14_,
    pv151_1_, pv199_5_, pv151_0_, pv183_10_, pv199_4_, pv151_3_, pv183_11_,
    pv199_7_, pv151_2_, pv167_10_, pv183_12_, pv199_6_, pv167_4_, pv199_1_,
    pv167_5_, pv199_0_, pv167_2_, pv199_3_, pv167_3_, pv199_2_, pv167_8_,
    pv199_14_, pv167_9_, pv199_15_, pv167_6_, pv199_12_, pv167_7_,
    pv199_13_, pv199_10_, pv199_11_, pv167_0_, pv183_6_, pv167_1_,
    pv183_7_, pv183_8_, pv183_9_, pv151_5_, pv151_14_, pv183_2_, pv183_13_,
    pv151_4_, pv151_15_, pv183_3_, pv183_14_, pv151_7_, pv151_12_,
    pv183_4_, pv183_15_, pv151_6_, pv151_13_, pv183_5_, pv151_9_,
    pv151_10_, pv167_15_, pv151_8_, pv151_11_, pv135_1_, pv183_0_,
    pv135_0_, pv183_1_  );
  input  pv16_9_, pv40_15_, pv88_6_, pv28_10_, pv88_7_, pv109_1_,
    pv118_3_, pv2_0_, pv40_13_, pv52_10_, pv109_2_, pv128_3_, pv2_1_,
    pv40_14_, pv52_11_, pv88_9_, pv109_3_, pv16_5_, pv40_11_, pv76_3_,
    pv88_2_, pv88_15_, pv100_14_, pv128_1_, pv16_13_, pv52_13_, pv76_2_,
    pv88_3_, pv100_13_, pv128_2_, pv16_7_, pv16_14_, pv52_14_, pv76_1_,
    pv88_13_, pv118_2_, pv16_6_, pv16_15_, pv40_10_, pv52_15_, pv88_5_,
    pv88_14_, pv100_15_, pv118_1_, pv128_0_, pv4_0_, pv52_9_, pv88_11_,
    pv100_3_, pv100_10_, pv121_2_, pv132_0_, pv4_1_, pv28_9_, pv64_1_,
    pv121_3_, pv16_10_, pv28_6_, pv100_5_, pv16_11_, pv28_7_, pv88_10_,
    pv100_6_, pv100_11_, pv121_1_, pv76_14_, pv28_5_, pv64_5_, pv76_15_,
    pv28_2_, pv64_2_, pv100_1_, pv28_3_, pv64_3_, pv100_2_, pv52_1_,
    pv76_10_, pv103_2_, pv124_1_, pv28_1_, pv64_9_, pv76_11_, pv103_3_,
    pv124_2_, pv52_3_, pv64_6_, pv64_15_, pv52_2_, pv64_7_, pv76_13_,
    pv52_5_, pv100_7_, pv112_2_, pv112_1_, pv132_3_, pv133_0_, pv52_7_,
    pv100_9_, pv132_2_, pv40_1_, pv52_6_, pv103_1_, pv112_3_, pv132_1_,
    pv16_1_, pv40_2_, pv76_7_, pv106_1_, pv40_3_, pv64_10_, pv76_6_,
    pv106_2_, pv16_3_, pv28_15_, pv76_5_, pv106_3_, pv16_2_, pv40_5_,
    pv88_1_, pv28_13_, pv40_6_, pv64_13_, pv115_1_, pv28_14_, pv40_7_,
    pv64_14_, pv28_11_, pv64_11_, pv76_9_, pv115_3_, pv124_3_, pv40_9_,
    pv115_2_;
  output pv167_11_, pv199_9_, pv167_12_, pv199_8_, pv167_13_, pv167_14_,
    pv151_1_, pv199_5_, pv151_0_, pv183_10_, pv199_4_, pv151_3_, pv183_11_,
    pv199_7_, pv151_2_, pv167_10_, pv183_12_, pv199_6_, pv167_4_, pv199_1_,
    pv167_5_, pv199_0_, pv167_2_, pv199_3_, pv167_3_, pv199_2_, pv167_8_,
    pv199_14_, pv167_9_, pv199_15_, pv167_6_, pv199_12_, pv167_7_,
    pv199_13_, pv199_10_, pv199_11_, pv167_0_, pv183_6_, pv167_1_,
    pv183_7_, pv183_8_, pv183_9_, pv151_5_, pv151_14_, pv183_2_, pv183_13_,
    pv151_4_, pv151_15_, pv183_3_, pv183_14_, pv151_7_, pv151_12_,
    pv183_4_, pv183_15_, pv151_6_, pv151_13_, pv183_5_, pv151_9_,
    pv151_10_, pv167_15_, pv151_8_, pv151_11_, pv135_1_, pv183_0_,
    pv135_0_, pv183_1_;
  wire new_n200_, new_n201_, new_n202_, new_n203_, new_n205_, new_n207_,
    new_n209_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_,
    new_n230_, new_n231_, new_n232_, new_n234_, new_n235_, new_n236_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_,
    new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_,
    new_n284_, new_n285_, new_n287_, new_n289_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n304_, new_n306_, new_n308_,
    new_n310_, new_n311_, new_n312_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n319_, new_n320_, new_n321_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_,
    new_n338_, new_n339_, new_n341_, new_n342_, new_n343_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n354_, new_n355_, new_n356_, new_n357_, new_n359_,
    new_n361_, new_n363_, new_n364_, new_n365_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n380_, new_n382_, new_n383_,
    new_n384_, new_n386_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n396_, new_n397_, new_n398_,
    new_n400_, new_n402_, new_n403_, new_n404_, new_n405_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n420_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n430_, new_n431_, new_n432_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n470_, new_n472_,
    new_n474_, new_n475_, new_n476_, new_n478_, new_n480_, new_n482_,
    new_n484_, new_n485_, new_n486_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n513_, new_n514_, new_n515_, new_n517_, new_n519_,
    new_n521_, new_n523_, new_n524_, new_n525_, new_n526_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_;
  assign new_n200_ = pv132_3_ & pv132_2_;
  assign new_n201_ = pv133_0_ & new_n200_;
  assign new_n202_ = pv128_3_ & pv132_2_;
  assign new_n203_ = ~pv128_2_ & ~new_n201_;
  assign pv183_0_ = new_n202_ | ~new_n203_;
  assign new_n205_ = pv112_3_ & pv183_0_;
  assign pv167_12_ = pv109_3_ | new_n205_;
  assign new_n207_ = pv52_11_ & pv167_12_;
  assign pv167_11_ = pv40_11_ | new_n207_;
  assign new_n209_ = pv133_0_ & pv124_3_;
  assign pv199_12_ = pv121_3_ | new_n209_;
  assign new_n211_ = pv100_10_ & pv100_11_;
  assign new_n212_ = pv100_9_ & new_n211_;
  assign new_n213_ = pv199_12_ & new_n212_;
  assign new_n214_ = pv88_10_ & pv100_9_;
  assign new_n215_ = pv88_11_ & pv100_9_;
  assign new_n216_ = pv100_10_ & new_n215_;
  assign new_n217_ = ~pv88_9_ & ~new_n213_;
  assign new_n218_ = ~new_n214_ & ~new_n216_;
  assign pv199_9_ = ~new_n217_ | ~new_n218_;
  assign new_n220_ = pv124_2_ & pv124_3_;
  assign new_n221_ = pv133_0_ & new_n220_;
  assign new_n222_ = pv121_3_ & pv124_2_;
  assign new_n223_ = ~pv121_2_ & ~new_n221_;
  assign pv199_8_ = new_n222_ | ~new_n223_;
  assign new_n225_ = pv52_14_ & pv52_15_;
  assign new_n226_ = pv52_13_ & new_n225_;
  assign new_n227_ = pv183_0_ & new_n226_;
  assign new_n228_ = pv40_14_ & pv52_13_;
  assign new_n229_ = pv40_15_ & pv52_13_;
  assign new_n230_ = pv52_14_ & new_n229_;
  assign new_n231_ = ~pv40_13_ & ~new_n227_;
  assign new_n232_ = ~new_n228_ & ~new_n230_;
  assign pv167_13_ = ~new_n231_ | ~new_n232_;
  assign new_n234_ = pv183_0_ & new_n225_;
  assign new_n235_ = pv40_15_ & pv52_14_;
  assign new_n236_ = ~pv40_14_ & ~new_n234_;
  assign pv167_14_ = new_n235_ | ~new_n236_;
  assign new_n238_ = pv132_1_ & new_n200_;
  assign new_n239_ = pv133_0_ & new_n238_;
  assign new_n240_ = pv128_2_ & pv132_1_;
  assign new_n241_ = pv128_3_ & pv132_1_;
  assign new_n242_ = pv132_2_ & new_n241_;
  assign new_n243_ = ~pv128_1_ & ~new_n239_;
  assign new_n244_ = ~new_n240_ & ~new_n242_;
  assign pv167_0_ = ~new_n243_ | ~new_n244_;
  assign new_n246_ = pv106_2_ & pv106_3_;
  assign new_n247_ = pv106_1_ & new_n246_;
  assign new_n248_ = pv167_0_ & new_n247_;
  assign new_n249_ = pv103_2_ & pv106_1_;
  assign new_n250_ = pv103_3_ & pv106_1_;
  assign new_n251_ = pv106_2_ & new_n250_;
  assign new_n252_ = ~pv103_1_ & ~new_n248_;
  assign new_n253_ = ~new_n249_ & ~new_n251_;
  assign pv151_4_ = ~new_n252_ | ~new_n253_;
  assign new_n255_ = pv28_2_ & pv28_3_;
  assign new_n256_ = pv28_1_ & new_n255_;
  assign new_n257_ = pv151_4_ & new_n256_;
  assign new_n258_ = pv28_1_ & pv16_2_;
  assign new_n259_ = pv28_1_ & pv16_3_;
  assign new_n260_ = pv28_2_ & new_n259_;
  assign new_n261_ = ~pv16_1_ & ~new_n257_;
  assign new_n262_ = ~new_n258_ & ~new_n260_;
  assign pv151_1_ = ~new_n261_ | ~new_n262_;
  assign new_n264_ = pv100_6_ & pv100_7_;
  assign new_n265_ = pv100_5_ & new_n264_;
  assign new_n266_ = pv199_8_ & new_n265_;
  assign new_n267_ = pv88_6_ & pv100_5_;
  assign new_n268_ = pv88_7_ & pv100_5_;
  assign new_n269_ = pv100_6_ & new_n268_;
  assign new_n270_ = ~pv88_5_ & ~new_n266_;
  assign new_n271_ = ~new_n267_ & ~new_n269_;
  assign pv199_5_ = ~new_n270_ | ~new_n271_;
  assign new_n273_ = pv128_2_ & pv132_0_;
  assign new_n274_ = pv132_1_ & new_n273_;
  assign new_n275_ = pv132_3_ & pv132_1_;
  assign new_n276_ = pv132_2_ & new_n275_;
  assign new_n277_ = pv132_0_ & new_n276_;
  assign new_n278_ = pv133_0_ & new_n277_;
  assign new_n279_ = pv128_1_ & pv132_0_;
  assign new_n280_ = pv132_0_ & pv132_1_;
  assign new_n281_ = pv128_3_ & new_n280_;
  assign new_n282_ = pv132_2_ & new_n281_;
  assign new_n283_ = ~new_n274_ & ~new_n278_;
  assign new_n284_ = ~new_n279_ & new_n283_;
  assign new_n285_ = ~pv128_0_ & ~new_n282_;
  assign pv151_0_ = ~new_n284_ | ~new_n285_;
  assign new_n287_ = pv132_3_ & pv133_0_;
  assign pv199_0_ = pv128_3_ | new_n287_;
  assign new_n289_ = pv118_3_ & pv199_0_;
  assign pv183_12_ = pv115_3_ | new_n289_;
  assign new_n291_ = pv76_10_ & pv76_11_;
  assign new_n292_ = pv183_12_ & new_n291_;
  assign new_n293_ = pv76_10_ & pv64_11_;
  assign new_n294_ = ~pv64_10_ & ~new_n292_;
  assign pv183_10_ = new_n293_ | ~new_n294_;
  assign new_n296_ = pv124_1_ & new_n220_;
  assign new_n297_ = pv133_0_ & new_n296_;
  assign new_n298_ = pv121_2_ & pv124_1_;
  assign new_n299_ = pv121_3_ & pv124_1_;
  assign new_n300_ = pv124_2_ & new_n299_;
  assign new_n301_ = ~pv121_1_ & ~new_n297_;
  assign new_n302_ = ~new_n298_ & ~new_n300_;
  assign pv199_4_ = ~new_n301_ | ~new_n302_;
  assign new_n304_ = pv28_3_ & pv151_4_;
  assign pv151_3_ = pv16_3_ | new_n304_;
  assign new_n306_ = pv76_11_ & pv183_12_;
  assign pv183_11_ = pv64_11_ | new_n306_;
  assign new_n308_ = pv100_7_ & pv199_8_;
  assign pv199_7_ = pv88_7_ | new_n308_;
  assign new_n310_ = pv151_4_ & new_n255_;
  assign new_n311_ = pv28_2_ & pv16_3_;
  assign new_n312_ = ~pv16_2_ & ~new_n310_;
  assign pv151_2_ = new_n311_ | ~new_n312_;
  assign new_n314_ = pv52_10_ & pv52_11_;
  assign new_n315_ = pv167_12_ & new_n314_;
  assign new_n316_ = pv52_10_ & pv40_11_;
  assign new_n317_ = ~pv40_10_ & ~new_n315_;
  assign pv167_10_ = new_n316_ | ~new_n317_;
  assign new_n319_ = pv199_8_ & new_n264_;
  assign new_n320_ = pv88_7_ & pv100_6_;
  assign new_n321_ = ~pv88_6_ & ~new_n319_;
  assign pv199_6_ = new_n320_ | ~new_n321_;
  assign new_n323_ = pv112_2_ & pv112_3_;
  assign new_n324_ = pv112_1_ & new_n323_;
  assign new_n325_ = pv183_0_ & new_n324_;
  assign new_n326_ = pv109_2_ & pv112_1_;
  assign new_n327_ = pv109_3_ & pv112_1_;
  assign new_n328_ = pv112_2_ & new_n327_;
  assign new_n329_ = ~pv109_1_ & ~new_n325_;
  assign new_n330_ = ~new_n326_ & ~new_n328_;
  assign pv167_4_ = ~new_n329_ | ~new_n330_;
  assign new_n332_ = pv100_3_ & pv100_2_;
  assign new_n333_ = pv100_1_ & new_n332_;
  assign new_n334_ = pv199_4_ & new_n333_;
  assign new_n335_ = pv88_2_ & pv100_1_;
  assign new_n336_ = pv88_3_ & pv100_1_;
  assign new_n337_ = pv100_2_ & new_n336_;
  assign new_n338_ = ~pv88_1_ & ~new_n334_;
  assign new_n339_ = ~new_n335_ & ~new_n337_;
  assign pv199_1_ = ~new_n338_ | ~new_n339_;
  assign new_n341_ = pv183_0_ & new_n323_;
  assign new_n342_ = pv109_3_ & pv112_2_;
  assign new_n343_ = ~pv109_2_ & ~new_n341_;
  assign pv167_8_ = new_n342_ | ~new_n343_;
  assign new_n345_ = pv52_7_ & pv52_6_;
  assign new_n346_ = pv52_5_ & new_n345_;
  assign new_n347_ = pv167_8_ & new_n346_;
  assign new_n348_ = pv52_5_ & pv40_6_;
  assign new_n349_ = pv52_5_ & pv40_7_;
  assign new_n350_ = pv52_6_ & new_n349_;
  assign new_n351_ = ~pv40_5_ & ~new_n347_;
  assign new_n352_ = ~new_n348_ & ~new_n350_;
  assign pv167_5_ = ~new_n351_ | ~new_n352_;
  assign new_n354_ = pv52_3_ & pv52_2_;
  assign new_n355_ = pv167_4_ & new_n354_;
  assign new_n356_ = pv52_2_ & pv40_3_;
  assign new_n357_ = ~pv40_2_ & ~new_n355_;
  assign pv167_2_ = new_n356_ | ~new_n357_;
  assign new_n359_ = pv100_3_ & pv199_4_;
  assign pv199_3_ = pv88_3_ | new_n359_;
  assign new_n361_ = pv52_3_ & pv167_4_;
  assign pv167_3_ = pv40_3_ | new_n361_;
  assign new_n363_ = pv199_4_ & new_n332_;
  assign new_n364_ = pv88_3_ & pv100_2_;
  assign new_n365_ = ~pv88_2_ & ~new_n363_;
  assign pv199_2_ = new_n364_ | ~new_n365_;
  assign new_n367_ = pv100_14_ & pv100_15_;
  assign new_n368_ = pv133_0_ & new_n367_;
  assign new_n369_ = pv88_15_ & pv100_14_;
  assign new_n370_ = ~pv88_14_ & ~new_n368_;
  assign pv199_14_ = new_n369_ | ~new_n370_;
  assign new_n372_ = pv52_9_ & new_n314_;
  assign new_n373_ = pv167_12_ & new_n372_;
  assign new_n374_ = pv40_10_ & pv52_9_;
  assign new_n375_ = pv40_11_ & pv52_9_;
  assign new_n376_ = pv52_10_ & new_n375_;
  assign new_n377_ = ~pv40_9_ & ~new_n373_;
  assign new_n378_ = ~new_n374_ & ~new_n376_;
  assign pv167_9_ = ~new_n377_ | ~new_n378_;
  assign new_n380_ = pv100_15_ & pv133_0_;
  assign pv199_15_ = pv88_15_ | new_n380_;
  assign new_n382_ = pv167_8_ & new_n345_;
  assign new_n383_ = pv52_6_ & pv40_7_;
  assign new_n384_ = ~pv40_6_ & ~new_n382_;
  assign pv167_6_ = new_n383_ | ~new_n384_;
  assign new_n386_ = pv52_7_ & pv167_8_;
  assign pv167_7_ = pv40_7_ | new_n386_;
  assign new_n388_ = pv100_13_ & new_n367_;
  assign new_n389_ = pv133_0_ & new_n388_;
  assign new_n390_ = pv100_13_ & pv88_14_;
  assign new_n391_ = pv88_15_ & pv100_13_;
  assign new_n392_ = pv100_14_ & new_n391_;
  assign new_n393_ = ~pv88_13_ & ~new_n389_;
  assign new_n394_ = ~new_n390_ & ~new_n392_;
  assign pv199_13_ = ~new_n393_ | ~new_n394_;
  assign new_n396_ = pv199_12_ & new_n211_;
  assign new_n397_ = pv88_11_ & pv100_10_;
  assign new_n398_ = ~pv88_10_ & ~new_n396_;
  assign pv199_10_ = new_n397_ | ~new_n398_;
  assign new_n400_ = pv100_11_ & pv199_12_;
  assign pv199_11_ = pv88_11_ | new_n400_;
  assign new_n402_ = pv118_3_ & pv118_2_;
  assign new_n403_ = pv199_0_ & new_n402_;
  assign new_n404_ = pv118_2_ & pv115_3_;
  assign new_n405_ = ~pv115_2_ & ~new_n403_;
  assign pv183_8_ = new_n404_ | ~new_n405_;
  assign new_n407_ = pv76_7_ & pv76_6_;
  assign new_n408_ = pv183_8_ & new_n407_;
  assign new_n409_ = pv64_7_ & pv76_6_;
  assign new_n410_ = ~pv64_6_ & ~new_n408_;
  assign pv183_6_ = new_n409_ | ~new_n410_;
  assign new_n412_ = pv52_1_ & new_n354_;
  assign new_n413_ = pv167_4_ & new_n412_;
  assign new_n414_ = pv52_1_ & pv40_2_;
  assign new_n415_ = pv52_1_ & pv40_3_;
  assign new_n416_ = pv52_2_ & new_n415_;
  assign new_n417_ = ~pv40_1_ & ~new_n413_;
  assign new_n418_ = ~new_n414_ & ~new_n416_;
  assign pv167_1_ = ~new_n417_ | ~new_n418_;
  assign new_n420_ = pv76_7_ & pv183_8_;
  assign pv183_7_ = pv64_7_ | new_n420_;
  assign new_n422_ = pv76_9_ & new_n291_;
  assign new_n423_ = pv183_12_ & new_n422_;
  assign new_n424_ = pv64_10_ & pv76_9_;
  assign new_n425_ = pv64_11_ & pv76_9_;
  assign new_n426_ = pv76_10_ & new_n425_;
  assign new_n427_ = ~pv64_9_ & ~new_n423_;
  assign new_n428_ = ~new_n424_ & ~new_n426_;
  assign pv183_9_ = ~new_n427_ | ~new_n428_;
  assign new_n430_ = pv167_0_ & new_n246_;
  assign new_n431_ = pv103_3_ & pv106_2_;
  assign new_n432_ = ~pv103_2_ & ~new_n430_;
  assign pv151_8_ = new_n431_ | ~new_n432_;
  assign new_n434_ = pv28_6_ & pv28_7_;
  assign new_n435_ = pv28_5_ & new_n434_;
  assign new_n436_ = pv151_8_ & new_n435_;
  assign new_n437_ = pv16_6_ & pv28_5_;
  assign new_n438_ = pv16_7_ & pv28_5_;
  assign new_n439_ = pv28_6_ & new_n438_;
  assign new_n440_ = ~pv16_5_ & ~new_n436_;
  assign new_n441_ = ~new_n437_ & ~new_n439_;
  assign pv151_5_ = ~new_n440_ | ~new_n441_;
  assign new_n443_ = pv28_15_ & pv28_14_;
  assign new_n444_ = pv167_0_ & new_n443_;
  assign new_n445_ = pv16_15_ & pv28_14_;
  assign new_n446_ = ~pv16_14_ & ~new_n444_;
  assign pv151_14_ = new_n445_ | ~new_n446_;
  assign new_n448_ = pv118_1_ & new_n402_;
  assign new_n449_ = pv199_0_ & new_n448_;
  assign new_n450_ = pv118_1_ & pv115_2_;
  assign new_n451_ = pv118_1_ & pv115_3_;
  assign new_n452_ = pv118_2_ & new_n451_;
  assign new_n453_ = ~pv115_1_ & ~new_n449_;
  assign new_n454_ = ~new_n450_ & ~new_n452_;
  assign pv183_4_ = ~new_n453_ | ~new_n454_;
  assign new_n456_ = pv76_3_ & pv76_2_;
  assign new_n457_ = pv183_4_ & new_n456_;
  assign new_n458_ = pv76_2_ & pv64_3_;
  assign new_n459_ = ~pv64_2_ & ~new_n457_;
  assign pv183_2_ = new_n458_ | ~new_n459_;
  assign new_n461_ = pv76_14_ & pv76_15_;
  assign new_n462_ = pv76_13_ & new_n461_;
  assign new_n463_ = pv199_0_ & new_n462_;
  assign new_n464_ = pv76_13_ & pv64_14_;
  assign new_n465_ = pv64_15_ & pv76_13_;
  assign new_n466_ = pv76_14_ & new_n465_;
  assign new_n467_ = ~pv64_13_ & ~new_n463_;
  assign new_n468_ = ~new_n464_ & ~new_n466_;
  assign pv183_13_ = ~new_n467_ | ~new_n468_;
  assign new_n470_ = pv28_15_ & pv167_0_;
  assign pv151_15_ = pv16_15_ | new_n470_;
  assign new_n472_ = pv76_3_ & pv183_4_;
  assign pv183_3_ = pv64_3_ | new_n472_;
  assign new_n474_ = pv199_0_ & new_n461_;
  assign new_n475_ = pv76_14_ & pv64_15_;
  assign new_n476_ = ~pv64_14_ & ~new_n474_;
  assign pv183_14_ = new_n475_ | ~new_n476_;
  assign new_n478_ = pv28_7_ & pv151_8_;
  assign pv151_7_ = pv16_7_ | new_n478_;
  assign new_n480_ = pv106_3_ & pv167_0_;
  assign pv151_12_ = pv103_3_ | new_n480_;
  assign new_n482_ = pv76_15_ & pv199_0_;
  assign pv183_15_ = pv64_15_ | new_n482_;
  assign new_n484_ = pv151_8_ & new_n434_;
  assign new_n485_ = pv16_7_ & pv28_6_;
  assign new_n486_ = ~pv16_6_ & ~new_n484_;
  assign pv151_6_ = new_n485_ | ~new_n486_;
  assign new_n488_ = pv28_13_ & new_n443_;
  assign new_n489_ = pv167_0_ & new_n488_;
  assign new_n490_ = pv16_14_ & pv28_13_;
  assign new_n491_ = pv16_15_ & pv28_13_;
  assign new_n492_ = pv28_14_ & new_n491_;
  assign new_n493_ = ~pv16_13_ & ~new_n489_;
  assign new_n494_ = ~new_n490_ & ~new_n492_;
  assign pv151_13_ = ~new_n493_ | ~new_n494_;
  assign new_n496_ = pv76_5_ & new_n407_;
  assign new_n497_ = pv183_8_ & new_n496_;
  assign new_n498_ = pv64_6_ & pv76_5_;
  assign new_n499_ = pv64_7_ & pv76_5_;
  assign new_n500_ = pv76_6_ & new_n499_;
  assign new_n501_ = ~pv64_5_ & ~new_n497_;
  assign new_n502_ = ~new_n498_ & ~new_n500_;
  assign pv183_5_ = ~new_n501_ | ~new_n502_;
  assign new_n504_ = pv28_10_ & pv28_11_;
  assign new_n505_ = pv28_9_ & new_n504_;
  assign new_n506_ = pv151_12_ & new_n505_;
  assign new_n507_ = pv28_9_ & pv16_10_;
  assign new_n508_ = pv28_9_ & pv16_11_;
  assign new_n509_ = pv28_10_ & new_n508_;
  assign new_n510_ = ~pv16_9_ & ~new_n506_;
  assign new_n511_ = ~new_n507_ & ~new_n509_;
  assign pv151_9_ = ~new_n510_ | ~new_n511_;
  assign new_n513_ = pv151_12_ & new_n504_;
  assign new_n514_ = pv28_10_ & pv16_11_;
  assign new_n515_ = ~pv16_10_ & ~new_n513_;
  assign pv151_10_ = new_n514_ | ~new_n515_;
  assign new_n517_ = pv52_15_ & pv183_0_;
  assign pv167_15_ = pv40_15_ | new_n517_;
  assign new_n519_ = pv28_11_ & pv151_12_;
  assign pv151_11_ = pv16_11_ | new_n519_;
  assign new_n521_ = pv4_1_ & pv151_0_;
  assign pv135_1_ = pv2_1_ | new_n521_;
  assign new_n523_ = pv4_0_ & pv4_1_;
  assign new_n524_ = pv151_0_ & new_n523_;
  assign new_n525_ = pv2_1_ & pv4_0_;
  assign new_n526_ = ~pv2_0_ & ~new_n524_;
  assign pv135_0_ = new_n525_ | ~new_n526_;
  assign new_n528_ = pv76_1_ & new_n456_;
  assign new_n529_ = pv183_4_ & new_n528_;
  assign new_n530_ = pv76_1_ & pv64_2_;
  assign new_n531_ = pv76_1_ & pv64_3_;
  assign new_n532_ = pv76_2_ & new_n531_;
  assign new_n533_ = ~pv64_1_ & ~new_n529_;
  assign new_n534_ = ~new_n530_ & ~new_n532_;
  assign pv183_1_ = ~new_n533_ | ~new_n534_;
endmodule

