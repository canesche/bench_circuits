// Benchmark "aes_core" written by ABC on Thu Oct  8 22:03:22 2020

module aes_core ( clock, 
    clk, rst, ld, \key[0] , \key[1] , \key[2] , \key[3] , \key[4] ,
    \key[5] , \key[6] , \key[7] , \key[8] , \key[9] , \key[10] , \key[11] ,
    \key[12] , \key[13] , \key[14] , \key[15] , \key[16] , \key[17] ,
    \key[18] , \key[19] , \key[20] , \key[21] , \key[22] , \key[23] ,
    \key[24] , \key[25] , \key[26] , \key[27] , \key[28] , \key[29] ,
    \key[30] , \key[31] , \key[32] , \key[33] , \key[34] , \key[35] ,
    \key[36] , \key[37] , \key[38] , \key[39] , \key[40] , \key[41] ,
    \key[42] , \key[43] , \key[44] , \key[45] , \key[46] , \key[47] ,
    \key[48] , \key[49] , \key[50] , \key[51] , \key[52] , \key[53] ,
    \key[54] , \key[55] , \key[56] , \key[57] , \key[58] , \key[59] ,
    \key[60] , \key[61] , \key[62] , \key[63] , \key[64] , \key[65] ,
    \key[66] , \key[67] , \key[68] , \key[69] , \key[70] , \key[71] ,
    \key[72] , \key[73] , \key[74] , \key[75] , \key[76] , \key[77] ,
    \key[78] , \key[79] , \key[80] , \key[81] , \key[82] , \key[83] ,
    \key[84] , \key[85] , \key[86] , \key[87] , \key[88] , \key[89] ,
    \key[90] , \key[91] , \key[92] , \key[93] , \key[94] , \key[95] ,
    \key[96] , \key[97] , \key[98] , \key[99] , \key[100] , \key[101] ,
    \key[102] , \key[103] , \key[104] , \key[105] , \key[106] , \key[107] ,
    \key[108] , \key[109] , \key[110] , \key[111] , \key[112] , \key[113] ,
    \key[114] , \key[115] , \key[116] , \key[117] , \key[118] , \key[119] ,
    \key[120] , \key[121] , \key[122] , \key[123] , \key[124] , \key[125] ,
    \key[126] , \key[127] , \text_in[0] , \text_in[1] , \text_in[2] ,
    \text_in[3] , \text_in[4] , \text_in[5] , \text_in[6] , \text_in[7] ,
    \text_in[8] , \text_in[9] , \text_in[10] , \text_in[11] ,
    \text_in[12] , \text_in[13] , \text_in[14] , \text_in[15] ,
    \text_in[16] , \text_in[17] , \text_in[18] , \text_in[19] ,
    \text_in[20] , \text_in[21] , \text_in[22] , \text_in[23] ,
    \text_in[24] , \text_in[25] , \text_in[26] , \text_in[27] ,
    \text_in[28] , \text_in[29] , \text_in[30] , \text_in[31] ,
    \text_in[32] , \text_in[33] , \text_in[34] , \text_in[35] ,
    \text_in[36] , \text_in[37] , \text_in[38] , \text_in[39] ,
    \text_in[40] , \text_in[41] , \text_in[42] , \text_in[43] ,
    \text_in[44] , \text_in[45] , \text_in[46] , \text_in[47] ,
    \text_in[48] , \text_in[49] , \text_in[50] , \text_in[51] ,
    \text_in[52] , \text_in[53] , \text_in[54] , \text_in[55] ,
    \text_in[56] , \text_in[57] , \text_in[58] , \text_in[59] ,
    \text_in[60] , \text_in[61] , \text_in[62] , \text_in[63] ,
    \text_in[64] , \text_in[65] , \text_in[66] , \text_in[67] ,
    \text_in[68] , \text_in[69] , \text_in[70] , \text_in[71] ,
    \text_in[72] , \text_in[73] , \text_in[74] , \text_in[75] ,
    \text_in[76] , \text_in[77] , \text_in[78] , \text_in[79] ,
    \text_in[80] , \text_in[81] , \text_in[82] , \text_in[83] ,
    \text_in[84] , \text_in[85] , \text_in[86] , \text_in[87] ,
    \text_in[88] , \text_in[89] , \text_in[90] , \text_in[91] ,
    \text_in[92] , \text_in[93] , \text_in[94] , \text_in[95] ,
    \text_in[96] , \text_in[97] , \text_in[98] , \text_in[99] ,
    \text_in[100] , \text_in[101] , \text_in[102] , \text_in[103] ,
    \text_in[104] , \text_in[105] , \text_in[106] , \text_in[107] ,
    \text_in[108] , \text_in[109] , \text_in[110] , \text_in[111] ,
    \text_in[112] , \text_in[113] , \text_in[114] , \text_in[115] ,
    \text_in[116] , \text_in[117] , \text_in[118] , \text_in[119] ,
    \text_in[120] , \text_in[121] , \text_in[122] , \text_in[123] ,
    \text_in[124] , \text_in[125] , \text_in[126] , \text_in[127] ,
    done, \text_out[0] , \text_out[1] , \text_out[2] , \text_out[3] ,
    \text_out[4] , \text_out[5] , \text_out[6] , \text_out[7] ,
    \text_out[8] , \text_out[9] , \text_out[10] , \text_out[11] ,
    \text_out[12] , \text_out[13] , \text_out[14] , \text_out[15] ,
    \text_out[16] , \text_out[17] , \text_out[18] , \text_out[19] ,
    \text_out[20] , \text_out[21] , \text_out[22] , \text_out[23] ,
    \text_out[24] , \text_out[25] , \text_out[26] , \text_out[27] ,
    \text_out[28] , \text_out[29] , \text_out[30] , \text_out[31] ,
    \text_out[32] , \text_out[33] , \text_out[34] , \text_out[35] ,
    \text_out[36] , \text_out[37] , \text_out[38] , \text_out[39] ,
    \text_out[40] , \text_out[41] , \text_out[42] , \text_out[43] ,
    \text_out[44] , \text_out[45] , \text_out[46] , \text_out[47] ,
    \text_out[48] , \text_out[49] , \text_out[50] , \text_out[51] ,
    \text_out[52] , \text_out[53] , \text_out[54] , \text_out[55] ,
    \text_out[56] , \text_out[57] , \text_out[58] , \text_out[59] ,
    \text_out[60] , \text_out[61] , \text_out[62] , \text_out[63] ,
    \text_out[64] , \text_out[65] , \text_out[66] , \text_out[67] ,
    \text_out[68] , \text_out[69] , \text_out[70] , \text_out[71] ,
    \text_out[72] , \text_out[73] , \text_out[74] , \text_out[75] ,
    \text_out[76] , \text_out[77] , \text_out[78] , \text_out[79] ,
    \text_out[80] , \text_out[81] , \text_out[82] , \text_out[83] ,
    \text_out[84] , \text_out[85] , \text_out[86] , \text_out[87] ,
    \text_out[88] , \text_out[89] , \text_out[90] , \text_out[91] ,
    \text_out[92] , \text_out[93] , \text_out[94] , \text_out[95] ,
    \text_out[96] , \text_out[97] , \text_out[98] , \text_out[99] ,
    \text_out[100] , \text_out[101] , \text_out[102] , \text_out[103] ,
    \text_out[104] , \text_out[105] , \text_out[106] , \text_out[107] ,
    \text_out[108] , \text_out[109] , \text_out[110] , \text_out[111] ,
    \text_out[112] , \text_out[113] , \text_out[114] , \text_out[115] ,
    \text_out[116] , \text_out[117] , \text_out[118] , \text_out[119] ,
    \text_out[120] , \text_out[121] , \text_out[122] , \text_out[123] ,
    \text_out[124] , \text_out[125] , \text_out[126] , \text_out[127]   );
  input  clock;
  input  clk, rst, ld, \key[0] , \key[1] , \key[2] , \key[3] , \key[4] ,
    \key[5] , \key[6] , \key[7] , \key[8] , \key[9] , \key[10] , \key[11] ,
    \key[12] , \key[13] , \key[14] , \key[15] , \key[16] , \key[17] ,
    \key[18] , \key[19] , \key[20] , \key[21] , \key[22] , \key[23] ,
    \key[24] , \key[25] , \key[26] , \key[27] , \key[28] , \key[29] ,
    \key[30] , \key[31] , \key[32] , \key[33] , \key[34] , \key[35] ,
    \key[36] , \key[37] , \key[38] , \key[39] , \key[40] , \key[41] ,
    \key[42] , \key[43] , \key[44] , \key[45] , \key[46] , \key[47] ,
    \key[48] , \key[49] , \key[50] , \key[51] , \key[52] , \key[53] ,
    \key[54] , \key[55] , \key[56] , \key[57] , \key[58] , \key[59] ,
    \key[60] , \key[61] , \key[62] , \key[63] , \key[64] , \key[65] ,
    \key[66] , \key[67] , \key[68] , \key[69] , \key[70] , \key[71] ,
    \key[72] , \key[73] , \key[74] , \key[75] , \key[76] , \key[77] ,
    \key[78] , \key[79] , \key[80] , \key[81] , \key[82] , \key[83] ,
    \key[84] , \key[85] , \key[86] , \key[87] , \key[88] , \key[89] ,
    \key[90] , \key[91] , \key[92] , \key[93] , \key[94] , \key[95] ,
    \key[96] , \key[97] , \key[98] , \key[99] , \key[100] , \key[101] ,
    \key[102] , \key[103] , \key[104] , \key[105] , \key[106] , \key[107] ,
    \key[108] , \key[109] , \key[110] , \key[111] , \key[112] , \key[113] ,
    \key[114] , \key[115] , \key[116] , \key[117] , \key[118] , \key[119] ,
    \key[120] , \key[121] , \key[122] , \key[123] , \key[124] , \key[125] ,
    \key[126] , \key[127] , \text_in[0] , \text_in[1] , \text_in[2] ,
    \text_in[3] , \text_in[4] , \text_in[5] , \text_in[6] , \text_in[7] ,
    \text_in[8] , \text_in[9] , \text_in[10] , \text_in[11] ,
    \text_in[12] , \text_in[13] , \text_in[14] , \text_in[15] ,
    \text_in[16] , \text_in[17] , \text_in[18] , \text_in[19] ,
    \text_in[20] , \text_in[21] , \text_in[22] , \text_in[23] ,
    \text_in[24] , \text_in[25] , \text_in[26] , \text_in[27] ,
    \text_in[28] , \text_in[29] , \text_in[30] , \text_in[31] ,
    \text_in[32] , \text_in[33] , \text_in[34] , \text_in[35] ,
    \text_in[36] , \text_in[37] , \text_in[38] , \text_in[39] ,
    \text_in[40] , \text_in[41] , \text_in[42] , \text_in[43] ,
    \text_in[44] , \text_in[45] , \text_in[46] , \text_in[47] ,
    \text_in[48] , \text_in[49] , \text_in[50] , \text_in[51] ,
    \text_in[52] , \text_in[53] , \text_in[54] , \text_in[55] ,
    \text_in[56] , \text_in[57] , \text_in[58] , \text_in[59] ,
    \text_in[60] , \text_in[61] , \text_in[62] , \text_in[63] ,
    \text_in[64] , \text_in[65] , \text_in[66] , \text_in[67] ,
    \text_in[68] , \text_in[69] , \text_in[70] , \text_in[71] ,
    \text_in[72] , \text_in[73] , \text_in[74] , \text_in[75] ,
    \text_in[76] , \text_in[77] , \text_in[78] , \text_in[79] ,
    \text_in[80] , \text_in[81] , \text_in[82] , \text_in[83] ,
    \text_in[84] , \text_in[85] , \text_in[86] , \text_in[87] ,
    \text_in[88] , \text_in[89] , \text_in[90] , \text_in[91] ,
    \text_in[92] , \text_in[93] , \text_in[94] , \text_in[95] ,
    \text_in[96] , \text_in[97] , \text_in[98] , \text_in[99] ,
    \text_in[100] , \text_in[101] , \text_in[102] , \text_in[103] ,
    \text_in[104] , \text_in[105] , \text_in[106] , \text_in[107] ,
    \text_in[108] , \text_in[109] , \text_in[110] , \text_in[111] ,
    \text_in[112] , \text_in[113] , \text_in[114] , \text_in[115] ,
    \text_in[116] , \text_in[117] , \text_in[118] , \text_in[119] ,
    \text_in[120] , \text_in[121] , \text_in[122] , \text_in[123] ,
    \text_in[124] , \text_in[125] , \text_in[126] , \text_in[127] ;
  output done, \text_out[0] , \text_out[1] , \text_out[2] , \text_out[3] ,
    \text_out[4] , \text_out[5] , \text_out[6] , \text_out[7] ,
    \text_out[8] , \text_out[9] , \text_out[10] , \text_out[11] ,
    \text_out[12] , \text_out[13] , \text_out[14] , \text_out[15] ,
    \text_out[16] , \text_out[17] , \text_out[18] , \text_out[19] ,
    \text_out[20] , \text_out[21] , \text_out[22] , \text_out[23] ,
    \text_out[24] , \text_out[25] , \text_out[26] , \text_out[27] ,
    \text_out[28] , \text_out[29] , \text_out[30] , \text_out[31] ,
    \text_out[32] , \text_out[33] , \text_out[34] , \text_out[35] ,
    \text_out[36] , \text_out[37] , \text_out[38] , \text_out[39] ,
    \text_out[40] , \text_out[41] , \text_out[42] , \text_out[43] ,
    \text_out[44] , \text_out[45] , \text_out[46] , \text_out[47] ,
    \text_out[48] , \text_out[49] , \text_out[50] , \text_out[51] ,
    \text_out[52] , \text_out[53] , \text_out[54] , \text_out[55] ,
    \text_out[56] , \text_out[57] , \text_out[58] , \text_out[59] ,
    \text_out[60] , \text_out[61] , \text_out[62] , \text_out[63] ,
    \text_out[64] , \text_out[65] , \text_out[66] , \text_out[67] ,
    \text_out[68] , \text_out[69] , \text_out[70] , \text_out[71] ,
    \text_out[72] , \text_out[73] , \text_out[74] , \text_out[75] ,
    \text_out[76] , \text_out[77] , \text_out[78] , \text_out[79] ,
    \text_out[80] , \text_out[81] , \text_out[82] , \text_out[83] ,
    \text_out[84] , \text_out[85] , \text_out[86] , \text_out[87] ,
    \text_out[88] , \text_out[89] , \text_out[90] , \text_out[91] ,
    \text_out[92] , \text_out[93] , \text_out[94] , \text_out[95] ,
    \text_out[96] , \text_out[97] , \text_out[98] , \text_out[99] ,
    \text_out[100] , \text_out[101] , \text_out[102] , \text_out[103] ,
    \text_out[104] , \text_out[105] , \text_out[106] , \text_out[107] ,
    \text_out[108] , \text_out[109] , \text_out[110] , \text_out[111] ,
    \text_out[112] , \text_out[113] , \text_out[114] , \text_out[115] ,
    \text_out[116] , \text_out[117] , \text_out[118] , \text_out[119] ,
    \text_out[120] , \text_out[121] , \text_out[122] , \text_out[123] ,
    \text_out[124] , \text_out[125] , \text_out[126] , \text_out[127] ;
  reg \\sa22_reg[4] , \\sa02_reg[1] , \\sa01_reg[1] , \\sa00_reg[1] ,
    \\sa03_reg[4] , \\sa03_reg[3] , \\sa33_reg[0] , \\sa02_reg[4] ,
    \\sa12_reg[3] , \\sa32_reg[3] , \\sa32_reg[0] , \\sa22_reg[3] ,
    \\sa31_reg[0] , \\sa02_reg[3] , \\sa20_reg[3] , \\sa30_reg[0] ,
    \\sa00_reg[4] , \\sa10_reg[0] , \\sa03_reg[0] , \\sa33_reg[3] ,
    \\sa13_reg[0] , \\sa02_reg[6] , \\sa22_reg[5] , \\sa13_reg[4] ,
    \\sa03_reg[1] , \\sa32_reg[5] , \\sa12_reg[1] , \\sa13_reg[3] ,
    \\sa23_reg[3] , \\sa02_reg[0] , \\sa12_reg[0] , \\sa21_reg[4] ,
    \\sa01_reg[4] , \\sa31_reg[5] , \\sa11_reg[1] , \\sa21_reg[3] ,
    \\sa01_reg[0] , \\sa21_reg[5] , \\sa11_reg[0] , \\sa10_reg[1] ,
    \\sa20_reg[1] , \\sa00_reg[5] , \\sa30_reg[6] , \\sa10_reg[3] ,
    \\sa00_reg[0] , \\sa00_reg[7] , \\sa23_reg[6] , \\sa13_reg[6] ,
    \\sa13_reg[1] , \\sa33_reg[4] , \\sa23_reg[7] , \\sa33_reg[7] ,
    \\sa03_reg[6] , \\sa23_reg[0] , \\sa02_reg[5] , \\sa32_reg[6] ,
    \\sa12_reg[6] , \\sa22_reg[6] , \\sa22_reg[1] , \\sa12_reg[4] ,
    \\sa22_reg[0] , \\sa01_reg[6] , \\sa11_reg[6] , \\sa31_reg[6] ,
    \\sa01_reg[5] , \\sa21_reg[1] , \\sa11_reg[3] , \\sa01_reg[3] ,
    \\sa21_reg[0] , \\sa31_reg[3] , \\sa10_reg[5] , \\sa30_reg[5] ,
    \\sa20_reg[5] , \\sa30_reg[1] , \\sa00_reg[3] , \\sa30_reg[4] ,
    \\sa10_reg[4] , \\sa10_reg[6] , \\sa20_reg[0] , \\sa30_reg[3] ,
    \\sa30_reg[2] , \\sa00_reg[6] , \\sa20_reg[6] , \\sa20_reg[2] ,
    \\sa03_reg[5] , \\sa23_reg[4] , \\sa33_reg[5] , \\sa23_reg[5] ,
    \\sa33_reg[1] , \\sa23_reg[1] , \\sa33_reg[2] , \\sa03_reg[2] ,
    \\sa23_reg[2] , \\sa13_reg[7] , \\sa03_reg[7] , \\sa12_reg[5] ,
    \\sa32_reg[1] , \\sa22_reg[7] , \\sa02_reg[7] , \\sa12_reg[7] ,
    \\sa21_reg[6] , \\sa11_reg[5] , \\sa31_reg[1] , \\sa11_reg[4] ,
    \\sa31_reg[2] , \\sa01_reg[7] , \\sa21_reg[2] , \\sa20_reg[4] ,
    \\sa20_reg[7] , \\sa10_reg[7] , \\sa30_reg[7] , \\sa13_reg[5] ,
    \\sa33_reg[6] , \\sa32_reg[2] , \\sa02_reg[2] , \\sa12_reg[2] ,
    \\sa22_reg[2] , \\sa01_reg[2] , \\sa11_reg[2] , \\sa11_reg[7] ,
    \\sa00_reg[2] , \\u0_w_reg[2][19] , \\sa10_reg[2] , \\sa13_reg[2] ,
    \\sa32_reg[7] , \\sa32_reg[4] , \\sa31_reg[7] , \\sa31_reg[4] ,
    \\sa21_reg[7] , \\u0_w_reg[3][29] , \\u0_w_reg[0][19] ,
    \\u0_w_reg[1][19] , \\u0_w_reg[3][19] , \\u0_w_reg[2][21] ,
    \\u0_w_reg[0][27] , \\u0_w_reg[1][27] , \\u0_w_reg[2][27] ,
    \\u0_w_reg[2][11] , \\u0_w_reg[3][27] , \\u0_w_reg[3][24] ,
    \\u0_w_reg[2][29] , \\u0_w_reg[0][29] , \\u0_w_reg[2][5] ,
    \\u0_w_reg[2][3] , \\u0_w_reg[1][29] , \\u0_w_reg[0][30] ,
    \\u0_w_reg[1][30] , \\u0_w_reg[3][30] , \\u0_w_reg[0][21] ,
    \\u0_w_reg[1][21] , \\u0_w_reg[2][0] , \\u0_w_reg[2][10] ,
    \\u0_w_reg[2][14] , \\u0_w_reg[2][30] , \\u0_w_reg[2][16] ,
    \\u0_w_reg[2][8] , \\u0_w_reg[2][15] , \\u0_w_reg[3][21] ,
    \\text_out_reg[12] , \\u0_w_reg[2][12] , \\u0_w_reg[0][24] ,
    \\u0_w_reg[0][31] , \\u0_w_reg[1][24] , \\u0_w_reg[1][31] ,
    \\u0_w_reg[2][24] , \\u0_w_reg[2][31] , \\u0_w_reg[3][31] ,
    \\u0_w_reg[0][5] , \\u0_w_reg[2][22] , \\u0_w_reg[2][6] ,
    \\u0_w_reg[3][5] , \\u0_w_reg[0][11] , \\u0_w_reg[1][11] ,
    \\u0_w_reg[2][17] , \\u0_w_reg[2][9] , \\u0_w_reg[3][11] ,
    \\text_out_reg[125] , \\text_out_reg[44] , \\u0_w_reg[1][5] ,
    \\u0_w_reg[2][13] , \\u0_w_reg[1][3] , \\u0_w_reg[0][3] ,
    \\u0_w_reg[3][3] , \\u0_w_reg[2][4] , \\u0_w_reg[1][28] ,
    \\u0_w_reg[3][28] , \\text_out_reg[93] , \\u0_w_reg[0][0] ,
    \\text_out_reg[61] , \\u0_w_reg[0][16] , \\u0_w_reg[1][0] ,
    \\u0_w_reg[3][0] , \\u0_w_reg[1][16] , \\u0_w_reg[3][16] ,
    \\text_out_reg[101] , \\text_out_reg[108] , \\text_out_reg[43] ,
    \\text_out_reg[109] , \\text_out_reg[117] , \\text_out_reg[76] ,
    \\text_out_reg[111] , \\text_out_reg[48] , \\text_out_reg[80] ,
    \\text_out_reg[112] , \\text_out_reg[46] , \\text_out_reg[126] ,
    \\text_out_reg[10] , \\u0_w_reg[3][26] , \\u0_w_reg[1][26] ,
    \\u0_w_reg[2][26] , \\u0_w_reg[0][26] , \\text_out_reg[0] ,
    \\text_out_reg[4] , \\text_out_reg[6] , \\text_out_reg[32] ,
    \\u0_w_reg[3][14] , \\text_out_reg[64] , \\u0_w_reg[2][18] ,
    \\u0_w_reg[2][2] , \\u0_w_reg[2][23] , \\u0_w_reg[2][20] ,
    \\u0_w_reg[2][28] , \\u0_w_reg[0][10] , \\u0_w_reg[0][13] ,
    \\u0_w_reg[0][15] , \\u0_w_reg[0][8] , \\u0_w_reg[1][13] ,
    \\u0_w_reg[1][14] , \\u0_w_reg[1][15] , \\u0_w_reg[1][10] ,
    \\u0_w_reg[1][8] , \\u0_w_reg[3][10] , \\u0_w_reg[3][13] ,
    \\u0_w_reg[3][15] , \\u0_w_reg[3][8] , \\text_out_reg[29] ,
    \\text_out_reg[51] , \\text_out_reg[45] , \\text_out_reg[105] ,
    \\text_out_reg[104] , \\text_out_reg[77] , \\text_out_reg[13] ,
    \\text_out_reg[115] , \\text_out_reg[19] , \\text_out_reg[47] ,
    \\text_out_reg[42] , \\text_out_reg[79] , \\text_out_reg[74] ,
    \\text_out_reg[100] , \\text_out_reg[62] , \\text_out_reg[94] ,
    \\text_out_reg[110] , \\text_out_reg[78] , \\text_out_reg[121] ,
    \\text_out_reg[124] , \\u0_w_reg[0][28] , \\u0_w_reg[0][14] ,
    \\u0_w_reg[2][1] , \\u0_w_reg[2][7] , \\text_out_reg[21] ,
    \\text_out_reg[120] , \\text_out_reg[16] , \\text_out_reg[5] ,
    \\text_out_reg[37] , \\text_out_reg[35] , \\text_out_reg[69] ,
    \\text_out_reg[67] , \\u0_w_reg[2][25] , \\u0_w_reg[1][25] ,
    \\u0_w_reg[0][12] , \\u0_w_reg[3][12] , \\u0_w_reg[0][22] ,
    \\u0_w_reg[0][6] , \\u0_w_reg[1][22] , \\u0_w_reg[1][6] ,
    \\u0_w_reg[3][22] , \\u0_w_reg[3][6] , \\text_out_reg[56] ,
    \\u0_w_reg[0][17] , \\text_out_reg[88] , \\u0_w_reg[0][9] ,
    \\u0_w_reg[1][17] , \\text_out_reg[53] , \\u0_w_reg[1][9] ,
    \\u0_w_reg[3][17] , \\u0_w_reg[3][9] , \\text_out_reg[85] ,
    \\text_out_reg[83] , \\text_out_reg[24] , \\text_out_reg[75] ,
    \\text_out_reg[123] , \\text_out_reg[73] , \\text_out_reg[106] ,
    \\text_out_reg[82] , \\text_out_reg[30] , \\text_out_reg[23] ,
    \\text_out_reg[18] , \\text_out_reg[114] , \\text_out_reg[57] ,
    \\text_out_reg[89] , \\text_out_reg[60] , \\u0_w_reg[1][12] ,
    \\u0_w_reg[3][25] , \\u0_w_reg[0][25] , \\text_out_reg[41] ,
    \\text_out_reg[1] , \\text_out_reg[7] , \\text_out_reg[38] ,
    \\text_out_reg[36] , \\text_out_reg[33] , \\text_out_reg[39] ,
    \\text_out_reg[68] , \\text_out_reg[70] , \\text_out_reg[71] ,
    \\text_out_reg[50] , \\text_out_reg[59] , \\text_out_reg[91] ,
    \\text_out_reg[40] , \\text_out_reg[72] , \\u0_w_reg[0][4] ,
    \\u0_w_reg[1][4] , \\u0_w_reg[3][4] , \\text_out_reg[9] ,
    \\text_out_reg[31] , \\text_out_reg[102] , \\text_out_reg[55] ,
    \\text_out_reg[54] , \\text_out_reg[90] , \\text_out_reg[119] ,
    \\text_out_reg[22] , \\text_out_reg[103] , \\text_out_reg[15] ,
    \\text_out_reg[14] , \\text_out_reg[92] , \\text_out_reg[116] ,
    \\text_out_reg[66] , \\text_out_reg[11] , \\text_out_reg[34] ,
    \\text_out_reg[27] , \\text_out_reg[2] , \\text_out_reg[28] ,
    \\text_out_reg[25] , \\u0_w_reg[3][7] , \\text_out_reg[58] ,
    \\text_out_reg[122] , \\text_out_reg[3] , \\u0_w_reg[1][18] ,
    \\text_out_reg[65] , \\u0_w_reg[1][7] , \\u0_w_reg[0][2] ,
    \\u0_w_reg[1][2] , \\u0_w_reg[3][18] , \\u0_w_reg[3][2] ,
    \\u0_w_reg[0][23] , \\u0_w_reg[3][23] , \\text_out_reg[107] ,
    \\u0_w_reg[0][20] , \\u0_w_reg[1][20] , \\u0_w_reg[3][20] ,
    \\text_out_reg[97] , \\text_out_reg[63] , \\text_out_reg[96] ,
    \\text_out_reg[113] , \\text_out_reg[127] , \\text_out_reg[118] ,
    \\text_out_reg[26] , \\text_out_reg[98] , \\text_out_reg[52] ,
    \\text_out_reg[84] , \\text_out_reg[95] , \\u0_w_reg[0][7] ,
    \\u0_w_reg[0][18] , \\u0_w_reg[3][1] , \\u0_w_reg[1][1] ,
    \\text_out_reg[20] , \\u0_w_reg[1][23] , \\u0_w_reg[0][1] ,
    \\text_out_reg[86] , \\text_out_reg[81] , \\text_out_reg[99] ,
    \\text_out_reg[87] , \\text_out_reg[17] , \\text_out_reg[49] ,
    \\text_out_reg[8] , \\u0_r0_out_reg[28] , \\u0_r0_out_reg[26] ,
    \\u0_r0_out_reg[27] , \\dcnt_reg[3] , \\u0_r0_out_reg[29] ,
    \\u0_r0_out_reg[25] , \\dcnt_reg[2] , \\u0_r0_out_reg[30] ,
    \\u0_r0_out_reg[31] , \\dcnt_reg[1] , \\u0_r0_out_reg[24] ,
    \\dcnt_reg[0] , \\u0_r0_rcnt_reg[3] , done_reg, \\text_in_r_reg[116] ,
    \\text_in_r_reg[111] , \\text_in_r_reg[37] , \\text_in_r_reg[14] ,
    \\text_in_r_reg[67] , \\text_in_r_reg[47] , \\text_in_r_reg[18] ,
    \\text_in_r_reg[0] , \\text_in_r_reg[68] , \\text_in_r_reg[49] ,
    \\text_in_r_reg[42] , \\text_in_r_reg[127] , \\text_in_r_reg[64] ,
    \\text_in_r_reg[54] , \\text_in_r_reg[35] , \\text_in_r_reg[6] ,
    \\text_in_r_reg[17] , \\text_in_r_reg[108] , \\text_in_r_reg[11] ,
    \\text_in_r_reg[123] , \\text_in_r_reg[24] , \\text_in_r_reg[26] ,
    \\text_in_r_reg[29] , \\text_in_r_reg[46] , \\text_in_r_reg[55] ,
    \\text_in_r_reg[61] , \\text_in_r_reg[63] , \\text_in_r_reg[78] ,
    \\text_in_r_reg[81] , \\text_in_r_reg[86] , \\text_in_r_reg[8] ,
    \\text_in_r_reg[99] , \\text_in_r_reg[91] , \\text_in_r_reg[39] ,
    \\text_in_r_reg[60] , \\text_in_r_reg[103] , \\text_in_r_reg[23] ,
    \\text_in_r_reg[58] , \\text_in_r_reg[3] , \\text_in_r_reg[118] ,
    \\text_in_r_reg[59] , \\text_in_r_reg[96] , \\text_in_r_reg[70] ,
    \\text_in_r_reg[51] , \\text_in_r_reg[92] , \\text_in_r_reg[107] ,
    \\text_in_r_reg[28] , \\text_in_r_reg[77] , \\text_in_r_reg[1] ,
    \\text_in_r_reg[19] , \\text_in_r_reg[56] , \\text_in_r_reg[90] ,
    \\text_in_r_reg[69] , \\text_in_r_reg[12] , \\text_in_r_reg[85] ,
    \\text_in_r_reg[80] , \\text_in_r_reg[66] , \\text_in_r_reg[9] ,
    \\text_in_r_reg[53] , \\text_in_r_reg[45] , \\text_in_r_reg[52] ,
    \\text_in_r_reg[97] , \\text_in_r_reg[10] , \\text_in_r_reg[34] ,
    \\text_in_r_reg[110] , \\text_in_r_reg[30] , \\text_in_r_reg[104] ,
    \\text_in_r_reg[65] , \\text_in_r_reg[79] , \\text_in_r_reg[7] ,
    \\text_in_r_reg[82] , \\text_in_r_reg[126] , \\text_in_r_reg[105] ,
    \\text_in_r_reg[13] , \\text_in_r_reg[120] , \\text_in_r_reg[84] ,
    \\text_in_r_reg[74] , \\text_in_r_reg[16] , \\text_in_r_reg[40] ,
    \\text_in_r_reg[15] , \\text_in_r_reg[121] , \\text_in_r_reg[41] ,
    \\text_in_r_reg[36] , \\text_in_r_reg[20] , \\u0_r0_rcnt_reg[2] ,
    \\text_in_r_reg[32] , \\text_in_r_reg[75] , \\text_in_r_reg[88] ,
    \\text_in_r_reg[33] , \\u0_r0_rcnt_reg[1] , \\text_in_r_reg[125] ,
    \\text_in_r_reg[2] , \\text_in_r_reg[44] , \\text_in_r_reg[72] ,
    \\text_in_r_reg[101] , \\text_in_r_reg[106] , \\text_in_r_reg[4] ,
    \\text_in_r_reg[43] , \\text_in_r_reg[112] , \\text_in_r_reg[93] ,
    \\text_in_r_reg[73] , \\text_in_r_reg[50] , \\text_in_r_reg[100] ,
    \\text_in_r_reg[114] , \\text_in_r_reg[25] , \\text_in_r_reg[57] ,
    \\text_in_r_reg[95] , \\text_in_r_reg[124] , \\text_in_r_reg[115] ,
    \\text_in_r_reg[98] , \\text_in_r_reg[31] , \\text_in_r_reg[122] ,
    \\text_in_r_reg[119] , \\text_in_r_reg[102] , \\text_in_r_reg[76] ,
    \\text_in_r_reg[113] , \\text_in_r_reg[94] , \\text_in_r_reg[62] ,
    \\text_in_r_reg[48] , \\text_in_r_reg[27] , \\text_in_r_reg[109] ,
    \\text_in_r_reg[117] , \\u0_r0_rcnt_reg[0] , \\text_in_r_reg[21] ,
    \\text_in_r_reg[5] , \\text_in_r_reg[22] , \\text_in_r_reg[83] ,
    \\text_in_r_reg[38] , \\text_in_r_reg[71] , \\text_in_r_reg[89] ,
    \\text_in_r_reg[87] , ld_r_reg;
  wire \new_[920]_ , \new_[921]_ , \new_[922]_ , \new_[923]_ , \new_[924]_ ,
    \new_[925]_ , \new_[926]_ , \new_[927]_ , \new_[928]_ , \new_[929]_ ,
    \new_[930]_ , \new_[931]_ , \new_[932]_ , \new_[933]_ , \new_[934]_ ,
    \new_[935]_ , \new_[936]_ , \new_[937]_ , \new_[938]_ , \new_[939]_ ,
    \new_[940]_ , \new_[941]_ , \new_[942]_ , \new_[943]_ , \new_[944]_ ,
    \new_[945]_ , \new_[946]_ , \new_[947]_ , \new_[948]_ , \new_[949]_ ,
    \new_[950]_ , \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[954]_ ,
    \new_[955]_ , \new_[956]_ , \new_[957]_ , \new_[958]_ , \new_[959]_ ,
    \new_[960]_ , \new_[961]_ , \new_[962]_ , \new_[963]_ , \new_[964]_ ,
    \new_[965]_ , \new_[970]_ , \new_[972]_ , \new_[973]_ , \new_[974]_ ,
    \new_[975]_ , \new_[976]_ , \new_[977]_ , \new_[979]_ , \new_[980]_ ,
    \new_[981]_ , \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ ,
    \new_[986]_ , \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ ,
    \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ ,
    \new_[996]_ , \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ ,
    \new_[1001]_ , \new_[1002]_ , \new_[1003]_ , \new_[1004]_ ,
    \new_[1005]_ , \new_[1006]_ , \new_[1007]_ , \new_[1008]_ ,
    \new_[1009]_ , \new_[1021]_ , \new_[1022]_ , \new_[1023]_ ,
    \new_[1024]_ , \new_[1025]_ , \new_[1026]_ , \new_[1027]_ ,
    \new_[1028]_ , \new_[1029]_ , \new_[1030]_ , \new_[1031]_ ,
    \new_[1032]_ , \new_[1033]_ , \new_[1034]_ , \new_[1035]_ ,
    \new_[1036]_ , \new_[1037]_ , \new_[1038]_ , \new_[1039]_ ,
    \new_[1040]_ , \new_[1041]_ , \new_[1042]_ , \new_[1043]_ ,
    \new_[1044]_ , \new_[1045]_ , \new_[1046]_ , \new_[1047]_ ,
    \new_[1078]_ , \new_[1079]_ , \new_[1080]_ , \new_[1081]_ ,
    \new_[1082]_ , \new_[1083]_ , \new_[1084]_ , \new_[1085]_ ,
    \new_[1086]_ , \new_[1087]_ , \new_[1088]_ , \new_[1089]_ ,
    \new_[1091]_ , \new_[1110]_ , \new_[1113]_ , \new_[1114]_ ,
    \new_[1130]_ , \new_[1133]_ , \new_[1134]_ , \new_[1135]_ ,
    \new_[1136]_ , \new_[1137]_ , \new_[1138]_ , \new_[1139]_ ,
    \new_[1140]_ , \new_[1141]_ , \new_[1142]_ , \new_[1143]_ ,
    \new_[1163]_ , \new_[1166]_ , \new_[1168]_ , \new_[1169]_ ,
    \new_[1170]_ , \new_[1171]_ , \new_[1172]_ , \new_[1173]_ ,
    \new_[1174]_ , \new_[1175]_ , \new_[1178]_ , \new_[1181]_ ,
    \new_[1182]_ , \new_[1184]_ , \new_[1185]_ , \new_[1186]_ ,
    \new_[1187]_ , \new_[1188]_ , \new_[1189]_ , \new_[1190]_ ,
    \new_[1191]_ , \new_[1192]_ , \new_[1193]_ , \new_[1194]_ ,
    \new_[1195]_ , \new_[1196]_ , \new_[1197]_ , \new_[1198]_ ,
    \new_[1199]_ , \new_[1201]_ , \new_[1202]_ , \new_[1203]_ ,
    \new_[1204]_ , \new_[1205]_ , \new_[1206]_ , \new_[1207]_ ,
    \new_[1208]_ , \new_[1213]_ , \new_[1214]_ , \new_[1215]_ ,
    \new_[1216]_ , \new_[1217]_ , \new_[1218]_ , \new_[1219]_ ,
    \new_[1220]_ , \new_[1222]_ , \new_[1225]_ , \new_[1226]_ ,
    \new_[1227]_ , \new_[1228]_ , \new_[1229]_ , \new_[1230]_ ,
    \new_[1231]_ , \new_[1233]_ , \new_[1234]_ , \new_[1235]_ ,
    \new_[1236]_ , \new_[1237]_ , \new_[1238]_ , \new_[1239]_ ,
    \new_[1240]_ , \new_[1241]_ , \new_[1242]_ , \new_[1243]_ ,
    \new_[1244]_ , \new_[1245]_ , \new_[1246]_ , \new_[1247]_ ,
    \new_[1248]_ , \new_[1249]_ , \new_[1250]_ , \new_[1251]_ ,
    \new_[1252]_ , \new_[1253]_ , \new_[1254]_ , \new_[1257]_ ,
    \new_[1258]_ , \new_[1259]_ , \new_[1261]_ , \new_[1262]_ ,
    \new_[1263]_ , \new_[1265]_ , \new_[1268]_ , \new_[1269]_ ,
    \new_[1270]_ , \new_[1271]_ , \new_[1272]_ , \new_[1273]_ ,
    \new_[1274]_ , \new_[1275]_ , \new_[1276]_ , \new_[1277]_ ,
    \new_[1278]_ , \new_[1279]_ , \new_[1280]_ , \new_[1281]_ ,
    \new_[1282]_ , \new_[1283]_ , \new_[1284]_ , \new_[1286]_ ,
    \new_[1287]_ , \new_[1288]_ , \new_[1289]_ , \new_[1290]_ ,
    \new_[1291]_ , \new_[1292]_ , \new_[1293]_ , \new_[1294]_ ,
    \new_[1295]_ , \new_[1296]_ , \new_[1299]_ , \new_[1301]_ ,
    \new_[1302]_ , \new_[1303]_ , \new_[1304]_ , \new_[1305]_ ,
    \new_[1306]_ , \new_[1307]_ , \new_[1308]_ , \new_[1309]_ ,
    \new_[1310]_ , \new_[1311]_ , \new_[1312]_ , \new_[1313]_ ,
    \new_[1314]_ , \new_[1315]_ , \new_[1316]_ , \new_[1317]_ ,
    \new_[1318]_ , \new_[1319]_ , \new_[1320]_ , \new_[1321]_ ,
    \new_[1322]_ , \new_[1323]_ , \new_[1324]_ , \new_[1325]_ ,
    \new_[1326]_ , \new_[1327]_ , \new_[1328]_ , \new_[1329]_ ,
    \new_[1330]_ , \new_[1331]_ , \new_[1332]_ , \new_[1333]_ ,
    \new_[1334]_ , \new_[1335]_ , \new_[1336]_ , \new_[1337]_ ,
    \new_[1338]_ , \new_[1339]_ , \new_[1341]_ , \new_[1342]_ ,
    \new_[1343]_ , \new_[1344]_ , \new_[1345]_ , \new_[1346]_ ,
    \new_[1347]_ , \new_[1348]_ , \new_[1349]_ , \new_[1350]_ ,
    \new_[1351]_ , \new_[1352]_ , \new_[1353]_ , \new_[1354]_ ,
    \new_[1361]_ , \new_[1362]_ , \new_[1364]_ , \new_[1365]_ ,
    \new_[1366]_ , \new_[1367]_ , \new_[1368]_ , \new_[1369]_ ,
    \new_[1370]_ , \new_[1371]_ , \new_[1372]_ , \new_[1373]_ ,
    \new_[1374]_ , \new_[1375]_ , \new_[1376]_ , \new_[1377]_ ,
    \new_[1378]_ , \new_[1379]_ , \new_[1380]_ , \new_[1381]_ ,
    \new_[1382]_ , \new_[1383]_ , \new_[1384]_ , \new_[1385]_ ,
    \new_[1386]_ , \new_[1387]_ , \new_[1388]_ , \new_[1389]_ ,
    \new_[1390]_ , \new_[1391]_ , \new_[1392]_ , \new_[1393]_ ,
    \new_[1394]_ , \new_[1395]_ , \new_[1396]_ , \new_[1397]_ ,
    \new_[1398]_ , \new_[1399]_ , \new_[1400]_ , \new_[1401]_ ,
    \new_[1402]_ , \new_[1403]_ , \new_[1404]_ , \new_[1405]_ ,
    \new_[1406]_ , \new_[1407]_ , \new_[1408]_ , \new_[1409]_ ,
    \new_[1410]_ , \new_[1411]_ , \new_[1412]_ , \new_[1414]_ ,
    \new_[1417]_ , \new_[1418]_ , \new_[1419]_ , \new_[1420]_ ,
    \new_[1421]_ , \new_[1422]_ , \new_[1423]_ , \new_[1424]_ ,
    \new_[1425]_ , \new_[1426]_ , \new_[1427]_ , \new_[1428]_ ,
    \new_[1429]_ , \new_[1430]_ , \new_[1431]_ , \new_[1432]_ ,
    \new_[1433]_ , \new_[1434]_ , \new_[1437]_ , \new_[1439]_ ,
    \new_[1440]_ , \new_[1441]_ , \new_[1442]_ , \new_[1443]_ ,
    \new_[1444]_ , \new_[1445]_ , \new_[1446]_ , \new_[1447]_ ,
    \new_[1448]_ , \new_[1449]_ , \new_[1450]_ , \new_[1451]_ ,
    \new_[1452]_ , \new_[1453]_ , \new_[1454]_ , \new_[1455]_ ,
    \new_[1456]_ , \new_[1457]_ , \new_[1458]_ , \new_[1459]_ ,
    \new_[1460]_ , \new_[1461]_ , \new_[1462]_ , \new_[1463]_ ,
    \new_[1464]_ , \new_[1465]_ , \new_[1466]_ , \new_[1467]_ ,
    \new_[1468]_ , \new_[1469]_ , \new_[1470]_ , \new_[1471]_ ,
    \new_[1472]_ , \new_[1473]_ , \new_[1474]_ , \new_[1475]_ ,
    \new_[1476]_ , \new_[1477]_ , \new_[1478]_ , \new_[1479]_ ,
    \new_[1480]_ , \new_[1481]_ , \new_[1482]_ , \new_[1483]_ ,
    \new_[1484]_ , \new_[1485]_ , \new_[1486]_ , \new_[1487]_ ,
    \new_[1488]_ , \new_[1489]_ , \new_[1490]_ , \new_[1491]_ ,
    \new_[1492]_ , \new_[1493]_ , \new_[1494]_ , \new_[1495]_ ,
    \new_[1496]_ , \new_[1497]_ , \new_[1498]_ , \new_[1499]_ ,
    \new_[1500]_ , \new_[1501]_ , \new_[1502]_ , \new_[1503]_ ,
    \new_[1504]_ , \new_[1506]_ , \new_[1507]_ , \new_[1508]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1513]_ ,
    \new_[1515]_ , \new_[1516]_ , \new_[1517]_ , \new_[1518]_ ,
    \new_[1519]_ , \new_[1533]_ , \new_[1536]_ , \new_[1542]_ ,
    \new_[1543]_ , \new_[1544]_ , \new_[1545]_ , \new_[1549]_ ,
    \new_[1551]_ , \new_[1552]_ , \new_[1553]_ , \new_[1556]_ ,
    \new_[1557]_ , \new_[1558]_ , \new_[1559]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1562]_ , \new_[1563]_ , \new_[1564]_ ,
    \new_[1565]_ , \new_[1566]_ , \new_[1567]_ , \new_[1568]_ ,
    \new_[1569]_ , \new_[1570]_ , \new_[1571]_ , \new_[1572]_ ,
    \new_[1573]_ , \new_[1574]_ , \new_[1575]_ , \new_[1576]_ ,
    \new_[1577]_ , \new_[1578]_ , \new_[1579]_ , \new_[1580]_ ,
    \new_[1581]_ , \new_[1582]_ , \new_[1583]_ , \new_[1584]_ ,
    \new_[1585]_ , \new_[1586]_ , \new_[1587]_ , \new_[1588]_ ,
    \new_[1589]_ , \new_[1590]_ , \new_[1591]_ , \new_[1592]_ ,
    \new_[1593]_ , \new_[1594]_ , \new_[1595]_ , \new_[1596]_ ,
    \new_[1597]_ , \new_[1598]_ , \new_[1599]_ , \new_[1600]_ ,
    \new_[1601]_ , \new_[1602]_ , \new_[1603]_ , \new_[1604]_ ,
    \new_[1605]_ , \new_[1606]_ , \new_[1607]_ , \new_[1608]_ ,
    \new_[1609]_ , \new_[1610]_ , \new_[1611]_ , \new_[1612]_ ,
    \new_[1613]_ , \new_[1614]_ , \new_[1615]_ , \new_[1616]_ ,
    \new_[1617]_ , \new_[1618]_ , \new_[1619]_ , \new_[1620]_ ,
    \new_[1621]_ , \new_[1622]_ , \new_[1623]_ , \new_[1624]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1627]_ , \new_[1628]_ ,
    \new_[1629]_ , \new_[1630]_ , \new_[1631]_ , \new_[1632]_ ,
    \new_[1633]_ , \new_[1634]_ , \new_[1635]_ , \new_[1636]_ ,
    \new_[1637]_ , \new_[1638]_ , \new_[1639]_ , \new_[1640]_ ,
    \new_[1641]_ , \new_[1642]_ , \new_[1643]_ , \new_[1644]_ ,
    \new_[1645]_ , \new_[1646]_ , \new_[1647]_ , \new_[1648]_ ,
    \new_[1649]_ , \new_[1650]_ , \new_[1651]_ , \new_[1656]_ ,
    \new_[1658]_ , \new_[1659]_ , \new_[1660]_ , \new_[1661]_ ,
    \new_[1662]_ , \new_[1663]_ , \new_[1664]_ , \new_[1665]_ ,
    \new_[1666]_ , \new_[1667]_ , \new_[1668]_ , \new_[1669]_ ,
    \new_[1670]_ , \new_[1671]_ , \new_[1672]_ , \new_[1673]_ ,
    \new_[1674]_ , \new_[1675]_ , \new_[1696]_ , \new_[1699]_ ,
    \new_[1705]_ , \new_[1706]_ , \new_[1707]_ , \new_[1711]_ ,
    \new_[1712]_ , \new_[1715]_ , \new_[1716]_ , \new_[1718]_ ,
    \new_[1719]_ , \new_[1720]_ , \new_[1721]_ , \new_[1722]_ ,
    \new_[1723]_ , \new_[1724]_ , \new_[1725]_ , \new_[1726]_ ,
    \new_[1727]_ , \new_[1728]_ , \new_[1729]_ , \new_[1730]_ ,
    \new_[1731]_ , \new_[1732]_ , \new_[1733]_ , \new_[1734]_ ,
    \new_[1735]_ , \new_[1736]_ , \new_[1737]_ , \new_[1738]_ ,
    \new_[1739]_ , \new_[1740]_ , \new_[1744]_ , \new_[1745]_ ,
    \new_[1746]_ , \new_[1747]_ , \new_[1748]_ , \new_[1751]_ ,
    \new_[1752]_ , \new_[1753]_ , \new_[1754]_ , \new_[1755]_ ,
    \new_[1756]_ , \new_[1757]_ , \new_[1758]_ , \new_[1759]_ ,
    \new_[1760]_ , \new_[1761]_ , \new_[1762]_ , \new_[1763]_ ,
    \new_[1764]_ , \new_[1765]_ , \new_[1766]_ , \new_[1767]_ ,
    \new_[1768]_ , \new_[1769]_ , \new_[1770]_ , \new_[1771]_ ,
    \new_[1773]_ , \new_[1774]_ , \new_[1775]_ , \new_[1776]_ ,
    \new_[1777]_ , \new_[1778]_ , \new_[1779]_ , \new_[1780]_ ,
    \new_[1781]_ , \new_[1782]_ , \new_[1783]_ , \new_[1784]_ ,
    \new_[1785]_ , \new_[1786]_ , \new_[1787]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1791]_ , \new_[1792]_ ,
    \new_[1793]_ , \new_[1794]_ , \new_[1795]_ , \new_[1796]_ ,
    \new_[1797]_ , \new_[1798]_ , \new_[1799]_ , \new_[1800]_ ,
    \new_[1801]_ , \new_[1803]_ , \new_[1804]_ , \new_[1805]_ ,
    \new_[1806]_ , \new_[1807]_ , \new_[1808]_ , \new_[1809]_ ,
    \new_[1810]_ , \new_[1811]_ , \new_[1812]_ , \new_[1813]_ ,
    \new_[1814]_ , \new_[1815]_ , \new_[1816]_ , \new_[1817]_ ,
    \new_[1818]_ , \new_[1819]_ , \new_[1820]_ , \new_[1821]_ ,
    \new_[1822]_ , \new_[1823]_ , \new_[1825]_ , \new_[1826]_ ,
    \new_[1827]_ , \new_[1828]_ , \new_[1829]_ , \new_[1830]_ ,
    \new_[1831]_ , \new_[1832]_ , \new_[1833]_ , \new_[1834]_ ,
    \new_[1835]_ , \new_[1836]_ , \new_[1837]_ , \new_[1838]_ ,
    \new_[1839]_ , \new_[1840]_ , \new_[1842]_ , \new_[1843]_ ,
    \new_[1844]_ , \new_[1845]_ , \new_[1847]_ , \new_[1848]_ ,
    \new_[1849]_ , \new_[1850]_ , \new_[1851]_ , \new_[1852]_ ,
    \new_[1853]_ , \new_[1854]_ , \new_[1855]_ , \new_[1861]_ ,
    \new_[1862]_ , \new_[1863]_ , \new_[1864]_ , \new_[1865]_ ,
    \new_[1866]_ , \new_[1867]_ , \new_[1868]_ , \new_[1869]_ ,
    \new_[1870]_ , \new_[1872]_ , \new_[1874]_ , \new_[1875]_ ,
    \new_[1877]_ , \new_[1878]_ , \new_[1879]_ , \new_[1903]_ ,
    \new_[1905]_ , \new_[1906]_ , \new_[1907]_ , \new_[1908]_ ,
    \new_[1909]_ , \new_[1912]_ , \new_[1914]_ , \new_[1915]_ ,
    \new_[1916]_ , \new_[1917]_ , \new_[1918]_ , \new_[1919]_ ,
    \new_[1920]_ , \new_[1921]_ , \new_[1922]_ , \new_[1923]_ ,
    \new_[1927]_ , \new_[1928]_ , \new_[1929]_ , \new_[1930]_ ,
    \new_[1931]_ , \new_[1932]_ , \new_[1933]_ , \new_[1934]_ ,
    \new_[1935]_ , \new_[1936]_ , \new_[1937]_ , \new_[1938]_ ,
    \new_[1939]_ , \new_[1940]_ , \new_[1941]_ , \new_[1942]_ ,
    \new_[1943]_ , \new_[1947]_ , \new_[1948]_ , \new_[1949]_ ,
    \new_[1950]_ , \new_[1951]_ , \new_[1952]_ , \new_[1953]_ ,
    \new_[1954]_ , \new_[1955]_ , \new_[1956]_ , \new_[1957]_ ,
    \new_[1958]_ , \new_[1959]_ , \new_[1960]_ , \new_[1964]_ ,
    \new_[1966]_ , \new_[1969]_ , \new_[1971]_ , \new_[1972]_ ,
    \new_[1973]_ , \new_[1974]_ , \new_[1975]_ , \new_[1976]_ ,
    \new_[1977]_ , \new_[1978]_ , \new_[1979]_ , \new_[1980]_ ,
    \new_[1981]_ , \new_[1984]_ , \new_[1985]_ , \new_[1986]_ ,
    \new_[1987]_ , \new_[1988]_ , \new_[1989]_ , \new_[1990]_ ,
    \new_[1991]_ , \new_[1992]_ , \new_[1993]_ , \new_[1994]_ ,
    \new_[1995]_ , \new_[1996]_ , \new_[1997]_ , \new_[1998]_ ,
    \new_[1999]_ , \new_[2000]_ , \new_[2001]_ , \new_[2002]_ ,
    \new_[2003]_ , \new_[2004]_ , \new_[2005]_ , \new_[2006]_ ,
    \new_[2008]_ , \new_[2009]_ , \new_[2010]_ , \new_[2011]_ ,
    \new_[2014]_ , \new_[2015]_ , \new_[2016]_ , \new_[2017]_ ,
    \new_[2018]_ , \new_[2019]_ , \new_[2020]_ , \new_[2021]_ ,
    \new_[2022]_ , \new_[2023]_ , \new_[2024]_ , \new_[2025]_ ,
    \new_[2026]_ , \new_[2027]_ , \new_[2028]_ , \new_[2029]_ ,
    \new_[2030]_ , \new_[2031]_ , \new_[2032]_ , \new_[2033]_ ,
    \new_[2034]_ , \new_[2035]_ , \new_[2038]_ , \new_[2039]_ ,
    \new_[2040]_ , \new_[2041]_ , \new_[2042]_ , \new_[2043]_ ,
    \new_[2044]_ , \new_[2045]_ , \new_[2046]_ , \new_[2047]_ ,
    \new_[2048]_ , \new_[2049]_ , \new_[2050]_ , \new_[2051]_ ,
    \new_[2052]_ , \new_[2055]_ , \new_[2056]_ , \new_[2057]_ ,
    \new_[2058]_ , \new_[2060]_ , \new_[2061]_ , \new_[2068]_ ,
    \new_[2072]_ , \new_[2078]_ , \new_[2079]_ , \new_[2080]_ ,
    \new_[2095]_ , \new_[2096]_ , \new_[2101]_ , \new_[2102]_ ,
    \new_[2103]_ , \new_[2104]_ , \new_[2106]_ , \new_[2107]_ ,
    \new_[2110]_ , \new_[2111]_ , \new_[2112]_ , \new_[2115]_ ,
    \new_[2118]_ , \new_[2119]_ , \new_[2120]_ , \new_[2121]_ ,
    \new_[2122]_ , \new_[2123]_ , \new_[2124]_ , \new_[2125]_ ,
    \new_[2133]_ , \new_[2134]_ , \new_[2135]_ , \new_[2136]_ ,
    \new_[2137]_ , \new_[2142]_ , \new_[2143]_ , \new_[2145]_ ,
    \new_[2146]_ , \new_[2147]_ , \new_[2148]_ , \new_[2149]_ ,
    \new_[2150]_ , \new_[2151]_ , \new_[2152]_ , \new_[2153]_ ,
    \new_[2155]_ , \new_[2156]_ , \new_[2159]_ , \new_[2161]_ ,
    \new_[2164]_ , \new_[2166]_ , \new_[2167]_ , \new_[2176]_ ,
    \new_[2178]_ , \new_[2179]_ , \new_[2180]_ , \new_[2181]_ ,
    \new_[2182]_ , \new_[2183]_ , \new_[2184]_ , \new_[2185]_ ,
    \new_[2188]_ , \new_[2189]_ , \new_[2190]_ , \new_[2191]_ ,
    \new_[2193]_ , \new_[2194]_ , \new_[2195]_ , \new_[2196]_ ,
    \new_[2197]_ , \new_[2198]_ , \new_[2199]_ , \new_[2200]_ ,
    \new_[2201]_ , \new_[2202]_ , \new_[2203]_ , \new_[2204]_ ,
    \new_[2205]_ , \new_[2206]_ , \new_[2207]_ , \new_[2208]_ ,
    \new_[2209]_ , \new_[2211]_ , \new_[2212]_ , \new_[2213]_ ,
    \new_[2214]_ , \new_[2215]_ , \new_[2216]_ , \new_[2217]_ ,
    \new_[2218]_ , \new_[2219]_ , \new_[2220]_ , \new_[2221]_ ,
    \new_[2222]_ , \new_[2223]_ , \new_[2224]_ , \new_[2225]_ ,
    \new_[2226]_ , \new_[2229]_ , \new_[2230]_ , \new_[2231]_ ,
    \new_[2232]_ , \new_[2233]_ , \new_[2234]_ , \new_[2235]_ ,
    \new_[2236]_ , \new_[2239]_ , \new_[2241]_ , \new_[2243]_ ,
    \new_[2248]_ , \new_[2249]_ , \new_[2250]_ , \new_[2251]_ ,
    \new_[2252]_ , \new_[2253]_ , \new_[2254]_ , \new_[2255]_ ,
    \new_[2256]_ , \new_[2257]_ , \new_[2258]_ , \new_[2259]_ ,
    \new_[2260]_ , \new_[2261]_ , \new_[2262]_ , \new_[2263]_ ,
    \new_[2264]_ , \new_[2266]_ , \new_[2267]_ , \new_[2268]_ ,
    \new_[2269]_ , \new_[2270]_ , \new_[2272]_ , \new_[2273]_ ,
    \new_[2274]_ , \new_[2275]_ , \new_[2276]_ , \new_[2277]_ ,
    \new_[2278]_ , \new_[2279]_ , \new_[2280]_ , \new_[2281]_ ,
    \new_[2282]_ , \new_[2283]_ , \new_[2285]_ , \new_[2288]_ ,
    \new_[2289]_ , \new_[2291]_ , \new_[2292]_ , \new_[2293]_ ,
    \new_[2294]_ , \new_[2295]_ , \new_[2296]_ , \new_[2297]_ ,
    \new_[2298]_ , \new_[2300]_ , \new_[2301]_ , \new_[2302]_ ,
    \new_[2314]_ , \new_[2316]_ , \new_[2317]_ , \new_[2318]_ ,
    \new_[2319]_ , \new_[2320]_ , \new_[2321]_ , \new_[2323]_ ,
    \new_[2324]_ , \new_[2325]_ , \new_[2326]_ , \new_[2327]_ ,
    \new_[2328]_ , \new_[2330]_ , \new_[2334]_ , \new_[2335]_ ,
    \new_[2336]_ , \new_[2337]_ , \new_[2339]_ , \new_[2340]_ ,
    \new_[2341]_ , \new_[2343]_ , \new_[2344]_ , \new_[2345]_ ,
    \new_[2346]_ , \new_[2351]_ , \new_[2356]_ , \new_[2357]_ ,
    \new_[2358]_ , \new_[2359]_ , \new_[2360]_ , \new_[2361]_ ,
    \new_[2362]_ , \new_[2366]_ , \new_[2367]_ , \new_[2368]_ ,
    \new_[2369]_ , \new_[2370]_ , \new_[2371]_ , \new_[2372]_ ,
    \new_[2373]_ , \new_[2374]_ , \new_[2375]_ , \new_[2376]_ ,
    \new_[2377]_ , \new_[2385]_ , \new_[2386]_ , \new_[2387]_ ,
    \new_[2388]_ , \new_[2389]_ , \new_[2390]_ , \new_[2391]_ ,
    \new_[2392]_ , \new_[2393]_ , \new_[2394]_ , \new_[2395]_ ,
    \new_[2396]_ , \new_[2397]_ , \new_[2398]_ , \new_[2399]_ ,
    \new_[2400]_ , \new_[2401]_ , \new_[2402]_ , \new_[2403]_ ,
    \new_[2404]_ , \new_[2405]_ , \new_[2406]_ , \new_[2407]_ ,
    \new_[2408]_ , \new_[2409]_ , \new_[2410]_ , \new_[2411]_ ,
    \new_[2412]_ , \new_[2413]_ , \new_[2414]_ , \new_[2415]_ ,
    \new_[2416]_ , \new_[2417]_ , \new_[2418]_ , \new_[2419]_ ,
    \new_[2421]_ , \new_[2422]_ , \new_[2423]_ , \new_[2424]_ ,
    \new_[2425]_ , \new_[2426]_ , \new_[2427]_ , \new_[2428]_ ,
    \new_[2429]_ , \new_[2430]_ , \new_[2431]_ , \new_[2432]_ ,
    \new_[2433]_ , \new_[2434]_ , \new_[2435]_ , \new_[2436]_ ,
    \new_[2437]_ , \new_[2439]_ , \new_[2440]_ , \new_[2441]_ ,
    \new_[2442]_ , \new_[2443]_ , \new_[2444]_ , \new_[2445]_ ,
    \new_[2446]_ , \new_[2447]_ , \new_[2448]_ , \new_[2449]_ ,
    \new_[2454]_ , \new_[2455]_ , \new_[2456]_ , \new_[2457]_ ,
    \new_[2458]_ , \new_[2459]_ , \new_[2460]_ , \new_[2461]_ ,
    \new_[2462]_ , \new_[2469]_ , \new_[2471]_ , \new_[2473]_ ,
    \new_[2474]_ , \new_[2475]_ , \new_[2476]_ , \new_[2477]_ ,
    \new_[2478]_ , \new_[2481]_ , \new_[2482]_ , \new_[2483]_ ,
    \new_[2485]_ , \new_[2486]_ , \new_[2487]_ , \new_[2488]_ ,
    \new_[2489]_ , \new_[2490]_ , \new_[2491]_ , \new_[2492]_ ,
    \new_[2493]_ , \new_[2494]_ , \new_[2495]_ , \new_[2496]_ ,
    \new_[2497]_ , \new_[2498]_ , \new_[2499]_ , \new_[2500]_ ,
    \new_[2501]_ , \new_[2502]_ , \new_[2503]_ , \new_[2504]_ ,
    \new_[2505]_ , \new_[2506]_ , \new_[2507]_ , \new_[2508]_ ,
    \new_[2509]_ , \new_[2511]_ , \new_[2512]_ , \new_[2513]_ ,
    \new_[2514]_ , \new_[2515]_ , \new_[2516]_ , \new_[2517]_ ,
    \new_[2518]_ , \new_[2519]_ , \new_[2520]_ , \new_[2521]_ ,
    \new_[2522]_ , \new_[2523]_ , \new_[2524]_ , \new_[2525]_ ,
    \new_[2529]_ , \new_[2531]_ , \new_[2532]_ , \new_[2533]_ ,
    \new_[2534]_ , \new_[2535]_ , \new_[2536]_ , \new_[2537]_ ,
    \new_[2539]_ , \new_[2540]_ , \new_[2541]_ , \new_[2542]_ ,
    \new_[2543]_ , \new_[2544]_ , \new_[2545]_ , \new_[2546]_ ,
    \new_[2547]_ , \new_[2548]_ , \new_[2549]_ , \new_[2550]_ ,
    \new_[2551]_ , \new_[2552]_ , \new_[2553]_ , \new_[2554]_ ,
    \new_[2555]_ , \new_[2556]_ , \new_[2558]_ , \new_[2559]_ ,
    \new_[2560]_ , \new_[2561]_ , \new_[2562]_ , \new_[2563]_ ,
    \new_[2564]_ , \new_[2566]_ , \new_[2567]_ , \new_[2569]_ ,
    \new_[2570]_ , \new_[2571]_ , \new_[2572]_ , \new_[2573]_ ,
    \new_[2574]_ , \new_[2577]_ , \new_[2578]_ , \new_[2579]_ ,
    \new_[2580]_ , \new_[2581]_ , \new_[2582]_ , \new_[2583]_ ,
    \new_[2584]_ , \new_[2585]_ , \new_[2586]_ , \new_[2587]_ ,
    \new_[2589]_ , \new_[2590]_ , \new_[2591]_ , \new_[2592]_ ,
    \new_[2593]_ , \new_[2594]_ , \new_[2595]_ , \new_[2596]_ ,
    \new_[2597]_ , \new_[2599]_ , \new_[2600]_ , \new_[2601]_ ,
    \new_[2603]_ , \new_[2604]_ , \new_[2605]_ , \new_[2606]_ ,
    \new_[2607]_ , \new_[2611]_ , \new_[2617]_ , \new_[2618]_ ,
    \new_[2619]_ , \new_[2621]_ , \new_[2622]_ , \new_[2623]_ ,
    \new_[2624]_ , \new_[2625]_ , \new_[2626]_ , \new_[2627]_ ,
    \new_[2628]_ , \new_[2630]_ , \new_[2632]_ , \new_[2633]_ ,
    \new_[2634]_ , \new_[2637]_ , \new_[2638]_ , \new_[2639]_ ,
    \new_[2640]_ , \new_[2641]_ , \new_[2642]_ , \new_[2643]_ ,
    \new_[2644]_ , \new_[2645]_ , \new_[2646]_ , \new_[2647]_ ,
    \new_[2648]_ , \new_[2649]_ , \new_[2651]_ , \new_[2652]_ ,
    \new_[2653]_ , \new_[2654]_ , \new_[2655]_ , \new_[2657]_ ,
    \new_[2658]_ , \new_[2659]_ , \new_[2660]_ , \new_[2661]_ ,
    \new_[2662]_ , \new_[2663]_ , \new_[2664]_ , \new_[2665]_ ,
    \new_[2666]_ , \new_[2667]_ , \new_[2668]_ , \new_[2669]_ ,
    \new_[2670]_ , \new_[2671]_ , \new_[2672]_ , \new_[2673]_ ,
    \new_[2674]_ , \new_[2675]_ , \new_[2676]_ , \new_[2677]_ ,
    \new_[2678]_ , \new_[2679]_ , \new_[2680]_ , \new_[2681]_ ,
    \new_[2682]_ , \new_[2683]_ , \new_[2684]_ , \new_[2685]_ ,
    \new_[2686]_ , \new_[2687]_ , \new_[2688]_ , \new_[2689]_ ,
    \new_[2690]_ , \new_[2692]_ , \new_[2693]_ , \new_[2694]_ ,
    \new_[2695]_ , \new_[2696]_ , \new_[2697]_ , \new_[2699]_ ,
    \new_[2701]_ , \new_[2702]_ , \new_[2703]_ , \new_[2704]_ ,
    \new_[2705]_ , \new_[2706]_ , \new_[2707]_ , \new_[2708]_ ,
    \new_[2712]_ , \new_[2713]_ , \new_[2716]_ , \new_[2717]_ ,
    \new_[2718]_ , \new_[2719]_ , \new_[2720]_ , \new_[2722]_ ,
    \new_[2723]_ , \new_[2724]_ , \new_[2726]_ , \new_[2727]_ ,
    \new_[2728]_ , \new_[2729]_ , \new_[2730]_ , \new_[2731]_ ,
    \new_[2732]_ , \new_[2733]_ , \new_[2734]_ , \new_[2735]_ ,
    \new_[2736]_ , \new_[2738]_ , \new_[2739]_ , \new_[2740]_ ,
    \new_[2741]_ , \new_[2742]_ , \new_[2743]_ , \new_[2744]_ ,
    \new_[2745]_ , \new_[2746]_ , \new_[2747]_ , \new_[2748]_ ,
    \new_[2749]_ , \new_[2750]_ , \new_[2751]_ , \new_[2752]_ ,
    \new_[2754]_ , \new_[2755]_ , \new_[2759]_ , \new_[2760]_ ,
    \new_[2761]_ , \new_[2762]_ , \new_[2763]_ , \new_[2764]_ ,
    \new_[2765]_ , \new_[2766]_ , \new_[2767]_ , \new_[2768]_ ,
    \new_[2769]_ , \new_[2770]_ , \new_[2771]_ , \new_[2772]_ ,
    \new_[2773]_ , \new_[2774]_ , \new_[2775]_ , \new_[2777]_ ,
    \new_[2778]_ , \new_[2779]_ , \new_[2780]_ , \new_[2781]_ ,
    \new_[2783]_ , \new_[2785]_ , \new_[2787]_ , \new_[2788]_ ,
    \new_[2789]_ , \new_[2790]_ , \new_[2791]_ , \new_[2792]_ ,
    \new_[2793]_ , \new_[2794]_ , \new_[2795]_ , \new_[2797]_ ,
    \new_[2798]_ , \new_[2799]_ , \new_[2800]_ , \new_[2801]_ ,
    \new_[2802]_ , \new_[2803]_ , \new_[2804]_ , \new_[2805]_ ,
    \new_[2809]_ , \new_[2810]_ , \new_[2811]_ , \new_[2812]_ ,
    \new_[2813]_ , \new_[2814]_ , \new_[2815]_ , \new_[2816]_ ,
    \new_[2817]_ , \new_[2818]_ , \new_[2819]_ , \new_[2820]_ ,
    \new_[2821]_ , \new_[2822]_ , \new_[2823]_ , \new_[2824]_ ,
    \new_[2825]_ , \new_[2826]_ , \new_[2827]_ , \new_[2828]_ ,
    \new_[2829]_ , \new_[2830]_ , \new_[2831]_ , \new_[2832]_ ,
    \new_[2833]_ , \new_[2834]_ , \new_[2835]_ , \new_[2836]_ ,
    \new_[2837]_ , \new_[2838]_ , \new_[2839]_ , \new_[2840]_ ,
    \new_[2841]_ , \new_[2842]_ , \new_[2843]_ , \new_[2844]_ ,
    \new_[2845]_ , \new_[2846]_ , \new_[2847]_ , \new_[2848]_ ,
    \new_[2849]_ , \new_[2850]_ , \new_[2851]_ , \new_[2852]_ ,
    \new_[2853]_ , \new_[2854]_ , \new_[2855]_ , \new_[2856]_ ,
    \new_[2857]_ , \new_[2858]_ , \new_[2859]_ , \new_[2863]_ ,
    \new_[2864]_ , \new_[2865]_ , \new_[2866]_ , \new_[2867]_ ,
    \new_[2868]_ , \new_[2869]_ , \new_[2870]_ , \new_[2871]_ ,
    \new_[2872]_ , \new_[2875]_ , \new_[2876]_ , \new_[2877]_ ,
    \new_[2878]_ , \new_[2880]_ , \new_[2881]_ , \new_[2882]_ ,
    \new_[2883]_ , \new_[2884]_ , \new_[2885]_ , \new_[2886]_ ,
    \new_[2887]_ , \new_[2889]_ , \new_[2890]_ , \new_[2891]_ ,
    \new_[2896]_ , \new_[2897]_ , \new_[2898]_ , \new_[2899]_ ,
    \new_[2900]_ , \new_[2901]_ , \new_[2902]_ , \new_[2906]_ ,
    \new_[2913]_ , \new_[2914]_ , \new_[2915]_ , \new_[2916]_ ,
    \new_[2917]_ , \new_[2918]_ , \new_[2919]_ , \new_[2920]_ ,
    \new_[2921]_ , \new_[2925]_ , \new_[2926]_ , \new_[2927]_ ,
    \new_[2929]_ , \new_[2930]_ , \new_[2931]_ , \new_[2932]_ ,
    \new_[2933]_ , \new_[2934]_ , \new_[2935]_ , \new_[2936]_ ,
    \new_[2937]_ , \new_[2938]_ , \new_[2939]_ , \new_[2940]_ ,
    \new_[2941]_ , \new_[2943]_ , \new_[2944]_ , \new_[2945]_ ,
    \new_[2946]_ , \new_[2947]_ , \new_[2948]_ , \new_[2949]_ ,
    \new_[2950]_ , \new_[2951]_ , \new_[2952]_ , \new_[2954]_ ,
    \new_[2957]_ , \new_[2959]_ , \new_[2960]_ , \new_[2961]_ ,
    \new_[2962]_ , \new_[2963]_ , \new_[2964]_ , \new_[2965]_ ,
    \new_[2966]_ , \new_[2967]_ , \new_[2968]_ , \new_[2969]_ ,
    \new_[2970]_ , \new_[2971]_ , \new_[2972]_ , \new_[2973]_ ,
    \new_[2974]_ , \new_[2975]_ , \new_[2976]_ , \new_[2977]_ ,
    \new_[2978]_ , \new_[2979]_ , \new_[2980]_ , \new_[2981]_ ,
    \new_[2982]_ , \new_[2983]_ , \new_[2984]_ , \new_[2985]_ ,
    \new_[2986]_ , \new_[2987]_ , \new_[2988]_ , \new_[2989]_ ,
    \new_[2990]_ , \new_[2992]_ , \new_[2993]_ , \new_[2994]_ ,
    \new_[2995]_ , \new_[2996]_ , \new_[2997]_ , \new_[2998]_ ,
    \new_[2999]_ , \new_[3000]_ , \new_[3001]_ , \new_[3002]_ ,
    \new_[3003]_ , \new_[3004]_ , \new_[3005]_ , \new_[3006]_ ,
    \new_[3007]_ , \new_[3009]_ , \new_[3010]_ , \new_[3011]_ ,
    \new_[3012]_ , \new_[3013]_ , \new_[3014]_ , \new_[3015]_ ,
    \new_[3016]_ , \new_[3017]_ , \new_[3018]_ , \new_[3019]_ ,
    \new_[3020]_ , \new_[3021]_ , \new_[3022]_ , \new_[3023]_ ,
    \new_[3024]_ , \new_[3025]_ , \new_[3026]_ , \new_[3027]_ ,
    \new_[3028]_ , \new_[3029]_ , \new_[3030]_ , \new_[3031]_ ,
    \new_[3032]_ , \new_[3033]_ , \new_[3034]_ , \new_[3035]_ ,
    \new_[3036]_ , \new_[3037]_ , \new_[3038]_ , \new_[3039]_ ,
    \new_[3040]_ , \new_[3041]_ , \new_[3042]_ , \new_[3043]_ ,
    \new_[3044]_ , \new_[3045]_ , \new_[3046]_ , \new_[3047]_ ,
    \new_[3048]_ , \new_[3049]_ , \new_[3050]_ , \new_[3051]_ ,
    \new_[3052]_ , \new_[3053]_ , \new_[3054]_ , \new_[3055]_ ,
    \new_[3056]_ , \new_[3057]_ , \new_[3058]_ , \new_[3059]_ ,
    \new_[3060]_ , \new_[3061]_ , \new_[3062]_ , \new_[3063]_ ,
    \new_[3064]_ , \new_[3065]_ , \new_[3066]_ , \new_[3067]_ ,
    \new_[3068]_ , \new_[3069]_ , \new_[3070]_ , \new_[3071]_ ,
    \new_[3072]_ , \new_[3073]_ , \new_[3074]_ , \new_[3075]_ ,
    \new_[3076]_ , \new_[3077]_ , \new_[3078]_ , \new_[3079]_ ,
    \new_[3080]_ , \new_[3081]_ , \new_[3082]_ , \new_[3083]_ ,
    \new_[3084]_ , \new_[3085]_ , \new_[3086]_ , \new_[3087]_ ,
    \new_[3088]_ , \new_[3089]_ , \new_[3090]_ , \new_[3092]_ ,
    \new_[3093]_ , \new_[3094]_ , \new_[3095]_ , \new_[3096]_ ,
    \new_[3097]_ , \new_[3098]_ , \new_[3099]_ , \new_[3100]_ ,
    \new_[3101]_ , \new_[3102]_ , \new_[3103]_ , \new_[3104]_ ,
    \new_[3105]_ , \new_[3106]_ , \new_[3107]_ , \new_[3108]_ ,
    \new_[3109]_ , \new_[3110]_ , \new_[3111]_ , \new_[3112]_ ,
    \new_[3113]_ , \new_[3114]_ , \new_[3115]_ , \new_[3116]_ ,
    \new_[3117]_ , \new_[3118]_ , \new_[3119]_ , \new_[3120]_ ,
    \new_[3121]_ , \new_[3122]_ , \new_[3123]_ , \new_[3124]_ ,
    \new_[3125]_ , \new_[3126]_ , \new_[3127]_ , \new_[3128]_ ,
    \new_[3129]_ , \new_[3130]_ , \new_[3131]_ , \new_[3132]_ ,
    \new_[3133]_ , \new_[3134]_ , \new_[3135]_ , \new_[3136]_ ,
    \new_[3137]_ , \new_[3138]_ , \new_[3139]_ , \new_[3140]_ ,
    \new_[3141]_ , \new_[3142]_ , \new_[3143]_ , \new_[3144]_ ,
    \new_[3145]_ , \new_[3146]_ , \new_[3147]_ , \new_[3148]_ ,
    \new_[3149]_ , \new_[3150]_ , \new_[3151]_ , \new_[3152]_ ,
    \new_[3153]_ , \new_[3154]_ , \new_[3155]_ , \new_[3156]_ ,
    \new_[3157]_ , \new_[3158]_ , \new_[3159]_ , \new_[3160]_ ,
    \new_[3161]_ , \new_[3162]_ , \new_[3163]_ , \new_[3164]_ ,
    \new_[3165]_ , \new_[3166]_ , \new_[3167]_ , \new_[3168]_ ,
    \new_[3169]_ , \new_[3170]_ , \new_[3171]_ , \new_[3172]_ ,
    \new_[3173]_ , \new_[3174]_ , \new_[3175]_ , \new_[3176]_ ,
    \new_[3177]_ , \new_[3178]_ , \new_[3179]_ , \new_[3180]_ ,
    \new_[3181]_ , \new_[3182]_ , \new_[3183]_ , \new_[3184]_ ,
    \new_[3185]_ , \new_[3186]_ , \new_[3187]_ , \new_[3188]_ ,
    \new_[3189]_ , \new_[3190]_ , \new_[3191]_ , \new_[3192]_ ,
    \new_[3193]_ , \new_[3194]_ , \new_[3195]_ , \new_[3196]_ ,
    \new_[3197]_ , \new_[3198]_ , \new_[3199]_ , \new_[3200]_ ,
    \new_[3201]_ , \new_[3202]_ , \new_[3203]_ , \new_[3204]_ ,
    \new_[3205]_ , \new_[3206]_ , \new_[3207]_ , \new_[3208]_ ,
    \new_[3209]_ , \new_[3210]_ , \new_[3211]_ , \new_[3212]_ ,
    \new_[3213]_ , \new_[3214]_ , \new_[3215]_ , \new_[3216]_ ,
    \new_[3217]_ , \new_[3218]_ , \new_[3219]_ , \new_[3220]_ ,
    \new_[3223]_ , \new_[3224]_ , \new_[3225]_ , \new_[3226]_ ,
    \new_[3227]_ , \new_[3228]_ , \new_[3229]_ , \new_[3230]_ ,
    \new_[3231]_ , \new_[3232]_ , \new_[3233]_ , \new_[3234]_ ,
    \new_[3235]_ , \new_[3236]_ , \new_[3237]_ , \new_[3238]_ ,
    \new_[3239]_ , \new_[3240]_ , \new_[3241]_ , \new_[3242]_ ,
    \new_[3243]_ , \new_[3244]_ , \new_[3245]_ , \new_[3246]_ ,
    \new_[3247]_ , \new_[3248]_ , \new_[3249]_ , \new_[3250]_ ,
    \new_[3251]_ , \new_[3252]_ , \new_[3253]_ , \new_[3254]_ ,
    \new_[3255]_ , \new_[3256]_ , \new_[3257]_ , \new_[3258]_ ,
    \new_[3259]_ , \new_[3260]_ , \new_[3261]_ , \new_[3262]_ ,
    \new_[3263]_ , \new_[3264]_ , \new_[3265]_ , \new_[3266]_ ,
    \new_[3267]_ , \new_[3268]_ , \new_[3269]_ , \new_[3270]_ ,
    \new_[3271]_ , \new_[3272]_ , \new_[3273]_ , \new_[3274]_ ,
    \new_[3275]_ , \new_[3276]_ , \new_[3277]_ , \new_[3278]_ ,
    \new_[3279]_ , \new_[3280]_ , \new_[3282]_ , \new_[3283]_ ,
    \new_[3284]_ , \new_[3285]_ , \new_[3286]_ , \new_[3287]_ ,
    \new_[3288]_ , \new_[3289]_ , \new_[3290]_ , \new_[3291]_ ,
    \new_[3292]_ , \new_[3293]_ , \new_[3294]_ , \new_[3295]_ ,
    \new_[3296]_ , \new_[3297]_ , \new_[3298]_ , \new_[3299]_ ,
    \new_[3300]_ , \new_[3301]_ , \new_[3302]_ , \new_[3303]_ ,
    \new_[3304]_ , \new_[3305]_ , \new_[3306]_ , \new_[3307]_ ,
    \new_[3308]_ , \new_[3309]_ , \new_[3310]_ , \new_[3311]_ ,
    \new_[3312]_ , \new_[3313]_ , \new_[3314]_ , \new_[3315]_ ,
    \new_[3316]_ , \new_[3317]_ , \new_[3318]_ , \new_[3319]_ ,
    \new_[3320]_ , \new_[3321]_ , \new_[3322]_ , \new_[3323]_ ,
    \new_[3324]_ , \new_[3325]_ , \new_[3326]_ , \new_[3327]_ ,
    \new_[3328]_ , \new_[3329]_ , \new_[3330]_ , \new_[3331]_ ,
    \new_[3332]_ , \new_[3333]_ , \new_[3334]_ , \new_[3335]_ ,
    \new_[3336]_ , \new_[3337]_ , \new_[3338]_ , \new_[3339]_ ,
    \new_[3340]_ , \new_[3341]_ , \new_[3342]_ , \new_[3344]_ ,
    \new_[3345]_ , \new_[3346]_ , \new_[3347]_ , \new_[3348]_ ,
    \new_[3349]_ , \new_[3350]_ , \new_[3351]_ , \new_[3352]_ ,
    \new_[3353]_ , \new_[3354]_ , \new_[3355]_ , \new_[3356]_ ,
    \new_[3357]_ , \new_[3358]_ , \new_[3359]_ , \new_[3360]_ ,
    \new_[3361]_ , \new_[3362]_ , \new_[3363]_ , \new_[3364]_ ,
    \new_[3365]_ , \new_[3366]_ , \new_[3367]_ , \new_[3368]_ ,
    \new_[3369]_ , \new_[3370]_ , \new_[3371]_ , \new_[3372]_ ,
    \new_[3373]_ , \new_[3374]_ , \new_[3375]_ , \new_[3376]_ ,
    \new_[3377]_ , \new_[3378]_ , \new_[3379]_ , \new_[3380]_ ,
    \new_[3381]_ , \new_[3382]_ , \new_[3383]_ , \new_[3384]_ ,
    \new_[3385]_ , \new_[3386]_ , \new_[3387]_ , \new_[3388]_ ,
    \new_[3389]_ , \new_[3390]_ , \new_[3391]_ , \new_[3392]_ ,
    \new_[3393]_ , \new_[3394]_ , \new_[3395]_ , \new_[3396]_ ,
    \new_[3397]_ , \new_[3398]_ , \new_[3399]_ , \new_[3400]_ ,
    \new_[3401]_ , \new_[3402]_ , \new_[3403]_ , \new_[3404]_ ,
    \new_[3405]_ , \new_[3406]_ , \new_[3407]_ , \new_[3408]_ ,
    \new_[3409]_ , \new_[3410]_ , \new_[3411]_ , \new_[3412]_ ,
    \new_[3413]_ , \new_[3414]_ , \new_[3415]_ , \new_[3416]_ ,
    \new_[3417]_ , \new_[3418]_ , \new_[3419]_ , \new_[3420]_ ,
    \new_[3421]_ , \new_[3422]_ , \new_[3423]_ , \new_[3424]_ ,
    \new_[3425]_ , \new_[3426]_ , \new_[3427]_ , \new_[3428]_ ,
    \new_[3429]_ , \new_[3430]_ , \new_[3431]_ , \new_[3432]_ ,
    \new_[3433]_ , \new_[3434]_ , \new_[3435]_ , \new_[3436]_ ,
    \new_[3437]_ , \new_[3438]_ , \new_[3439]_ , \new_[3440]_ ,
    \new_[3441]_ , \new_[3442]_ , \new_[3443]_ , \new_[3444]_ ,
    \new_[3445]_ , \new_[3446]_ , \new_[3447]_ , \new_[3448]_ ,
    \new_[3449]_ , \new_[3450]_ , \new_[3451]_ , \new_[3452]_ ,
    \new_[3453]_ , \new_[3454]_ , \new_[3455]_ , \new_[3456]_ ,
    \new_[3457]_ , \new_[3458]_ , \new_[3459]_ , \new_[3460]_ ,
    \new_[3461]_ , \new_[3462]_ , \new_[3463]_ , \new_[3464]_ ,
    \new_[3465]_ , \new_[3466]_ , \new_[3467]_ , \new_[3468]_ ,
    \new_[3469]_ , \new_[3470]_ , \new_[3471]_ , \new_[3472]_ ,
    \new_[3473]_ , \new_[3474]_ , \new_[3475]_ , \new_[3476]_ ,
    \new_[3477]_ , \new_[3478]_ , \new_[3479]_ , \new_[3480]_ ,
    \new_[3481]_ , \new_[3482]_ , \new_[3483]_ , \new_[3484]_ ,
    \new_[3485]_ , \new_[3486]_ , \new_[3487]_ , \new_[3488]_ ,
    \new_[3489]_ , \new_[3490]_ , \new_[3491]_ , \new_[3492]_ ,
    \new_[3493]_ , \new_[3494]_ , \new_[3495]_ , \new_[3496]_ ,
    \new_[3497]_ , \new_[3498]_ , \new_[3499]_ , \new_[3500]_ ,
    \new_[3501]_ , \new_[3502]_ , \new_[3503]_ , \new_[3504]_ ,
    \new_[3505]_ , \new_[3506]_ , \new_[3507]_ , \new_[3508]_ ,
    \new_[3509]_ , \new_[3510]_ , \new_[3511]_ , \new_[3512]_ ,
    \new_[3513]_ , \new_[3514]_ , \new_[3515]_ , \new_[3516]_ ,
    \new_[3517]_ , \new_[3518]_ , \new_[3519]_ , \new_[3520]_ ,
    \new_[3521]_ , \new_[3522]_ , \new_[3523]_ , \new_[3524]_ ,
    \new_[3525]_ , \new_[3526]_ , \new_[3527]_ , \new_[3528]_ ,
    \new_[3529]_ , \new_[3530]_ , \new_[3531]_ , \new_[3532]_ ,
    \new_[3533]_ , \new_[3534]_ , \new_[3535]_ , \new_[3536]_ ,
    \new_[3537]_ , \new_[3538]_ , \new_[3539]_ , \new_[3540]_ ,
    \new_[3541]_ , \new_[3542]_ , \new_[3543]_ , \new_[3544]_ ,
    \new_[3545]_ , \new_[3546]_ , \new_[3547]_ , \new_[3548]_ ,
    \new_[3549]_ , \new_[3550]_ , \new_[3551]_ , \new_[3552]_ ,
    \new_[3553]_ , \new_[3554]_ , \new_[3555]_ , \new_[3556]_ ,
    \new_[3557]_ , \new_[3558]_ , \new_[3559]_ , \new_[3560]_ ,
    \new_[3561]_ , \new_[3562]_ , \new_[3563]_ , \new_[3564]_ ,
    \new_[3565]_ , \new_[3566]_ , \new_[3567]_ , \new_[3568]_ ,
    \new_[3569]_ , \new_[3570]_ , \new_[3571]_ , \new_[3572]_ ,
    \new_[3573]_ , \new_[3574]_ , \new_[3575]_ , \new_[3576]_ ,
    \new_[3577]_ , \new_[3578]_ , \new_[3579]_ , \new_[3580]_ ,
    \new_[3581]_ , \new_[3582]_ , \new_[3583]_ , \new_[3584]_ ,
    \new_[3585]_ , \new_[3586]_ , \new_[3587]_ , \new_[3588]_ ,
    \new_[3589]_ , \new_[3590]_ , \new_[3591]_ , \new_[3592]_ ,
    \new_[3593]_ , \new_[3594]_ , \new_[3595]_ , \new_[3596]_ ,
    \new_[3597]_ , \new_[3598]_ , \new_[3599]_ , \new_[3600]_ ,
    \new_[3601]_ , \new_[3602]_ , \new_[3603]_ , \new_[3604]_ ,
    \new_[3605]_ , \new_[3606]_ , \new_[3607]_ , \new_[3608]_ ,
    \new_[3609]_ , \new_[3610]_ , \new_[3611]_ , \new_[3612]_ ,
    \new_[3613]_ , \new_[3614]_ , \new_[3615]_ , \new_[3616]_ ,
    \new_[3617]_ , \new_[3618]_ , \new_[3619]_ , \new_[3620]_ ,
    \new_[3621]_ , \new_[3622]_ , \new_[3623]_ , \new_[3624]_ ,
    \new_[3625]_ , \new_[3626]_ , \new_[3627]_ , \new_[3628]_ ,
    \new_[3629]_ , \new_[3630]_ , \new_[3631]_ , \new_[3632]_ ,
    \new_[3633]_ , \new_[3634]_ , \new_[3635]_ , \new_[3636]_ ,
    \new_[3637]_ , \new_[3638]_ , \new_[3639]_ , \new_[3640]_ ,
    \new_[3641]_ , \new_[3642]_ , \new_[3643]_ , \new_[3644]_ ,
    \new_[3645]_ , \new_[3646]_ , \new_[3647]_ , \new_[3648]_ ,
    \new_[3649]_ , \new_[3650]_ , \new_[3651]_ , \new_[3652]_ ,
    \new_[3653]_ , \new_[3654]_ , \new_[3655]_ , \new_[3656]_ ,
    \new_[3657]_ , \new_[3658]_ , \new_[3659]_ , \new_[3660]_ ,
    \new_[3661]_ , \new_[3662]_ , \new_[3663]_ , \new_[3664]_ ,
    \new_[3665]_ , \new_[3666]_ , \new_[3667]_ , \new_[3668]_ ,
    \new_[3669]_ , \new_[3670]_ , \new_[3671]_ , \new_[3672]_ ,
    \new_[3673]_ , \new_[3674]_ , \new_[3675]_ , \new_[3676]_ ,
    \new_[3677]_ , \new_[3678]_ , \new_[3679]_ , \new_[3680]_ ,
    \new_[3681]_ , \new_[3682]_ , \new_[3683]_ , \new_[3684]_ ,
    \new_[3685]_ , \new_[3686]_ , \new_[3687]_ , \new_[3688]_ ,
    \new_[3689]_ , \new_[3690]_ , \new_[3691]_ , \new_[3692]_ ,
    \new_[3693]_ , \new_[3694]_ , \new_[3695]_ , \new_[3696]_ ,
    \new_[3697]_ , \new_[3698]_ , \new_[3699]_ , \new_[3700]_ ,
    \new_[3701]_ , \new_[3702]_ , \new_[3703]_ , \new_[3704]_ ,
    \new_[3705]_ , \new_[3706]_ , \new_[3707]_ , \new_[3708]_ ,
    \new_[3709]_ , \new_[3710]_ , \new_[3711]_ , \new_[3712]_ ,
    \new_[3713]_ , \new_[3714]_ , \new_[3715]_ , \new_[3716]_ ,
    \new_[3717]_ , \new_[3718]_ , \new_[3719]_ , \new_[3720]_ ,
    \new_[3721]_ , \new_[3722]_ , \new_[3723]_ , \new_[3724]_ ,
    \new_[3725]_ , \new_[3726]_ , \new_[3727]_ , \new_[3728]_ ,
    \new_[3729]_ , \new_[3730]_ , \new_[3731]_ , \new_[3732]_ ,
    \new_[3733]_ , \new_[3734]_ , \new_[3735]_ , \new_[3736]_ ,
    \new_[3737]_ , \new_[3738]_ , \new_[3739]_ , \new_[3740]_ ,
    \new_[3741]_ , \new_[3742]_ , \new_[3743]_ , \new_[3744]_ ,
    \new_[3745]_ , \new_[3746]_ , \new_[3747]_ , \new_[3748]_ ,
    \new_[3749]_ , \new_[3750]_ , \new_[3751]_ , \new_[3752]_ ,
    \new_[3753]_ , \new_[3754]_ , \new_[3755]_ , \new_[3756]_ ,
    \new_[3757]_ , \new_[3758]_ , \new_[3759]_ , \new_[3760]_ ,
    \new_[3761]_ , \new_[3762]_ , \new_[3763]_ , \new_[3764]_ ,
    \new_[3765]_ , \new_[3766]_ , \new_[3767]_ , \new_[3768]_ ,
    \new_[3769]_ , \new_[3770]_ , \new_[3771]_ , \new_[3772]_ ,
    \new_[3773]_ , \new_[3774]_ , \new_[3775]_ , \new_[3776]_ ,
    \new_[3777]_ , \new_[3778]_ , \new_[3779]_ , \new_[3780]_ ,
    \new_[3781]_ , \new_[3782]_ , \new_[3783]_ , \new_[3784]_ ,
    \new_[3785]_ , \new_[3786]_ , \new_[3787]_ , \new_[3788]_ ,
    \new_[3789]_ , \new_[3790]_ , \new_[3791]_ , \new_[3792]_ ,
    \new_[3793]_ , \new_[3794]_ , \new_[3795]_ , \new_[3796]_ ,
    \new_[3797]_ , \new_[3798]_ , \new_[3799]_ , \new_[3800]_ ,
    \new_[3801]_ , \new_[3802]_ , \new_[3803]_ , \new_[3804]_ ,
    \new_[3805]_ , \new_[3806]_ , \new_[3807]_ , \new_[3808]_ ,
    \new_[3809]_ , \new_[3810]_ , \new_[3811]_ , \new_[3812]_ ,
    \new_[3813]_ , \new_[3814]_ , \new_[3815]_ , \new_[3816]_ ,
    \new_[3817]_ , \new_[3818]_ , \new_[3819]_ , \new_[3820]_ ,
    \new_[3821]_ , \new_[3822]_ , \new_[3823]_ , \new_[3824]_ ,
    \new_[3825]_ , \new_[3826]_ , \new_[3827]_ , \new_[3828]_ ,
    \new_[3829]_ , \new_[3830]_ , \new_[3831]_ , \new_[3832]_ ,
    \new_[3833]_ , \new_[3834]_ , \new_[3835]_ , \new_[3836]_ ,
    \new_[3837]_ , \new_[3838]_ , \new_[3839]_ , \new_[3840]_ ,
    \new_[3841]_ , \new_[3842]_ , \new_[3843]_ , \new_[3844]_ ,
    \new_[3845]_ , \new_[3846]_ , \new_[3847]_ , \new_[3848]_ ,
    \new_[3849]_ , \new_[3850]_ , \new_[3851]_ , \new_[3852]_ ,
    \new_[3853]_ , \new_[3854]_ , \new_[3855]_ , \new_[3856]_ ,
    \new_[3857]_ , \new_[3858]_ , \new_[3859]_ , \new_[3860]_ ,
    \new_[3861]_ , \new_[3862]_ , \new_[3863]_ , \new_[3864]_ ,
    \new_[3865]_ , \new_[3866]_ , \new_[3867]_ , \new_[3868]_ ,
    \new_[3869]_ , \new_[3870]_ , \new_[3871]_ , \new_[3872]_ ,
    \new_[3873]_ , \new_[3874]_ , \new_[3875]_ , \new_[3876]_ ,
    \new_[3877]_ , \new_[3878]_ , \new_[3879]_ , \new_[3880]_ ,
    \new_[3881]_ , \new_[3882]_ , \new_[3883]_ , \new_[3884]_ ,
    \new_[3885]_ , \new_[3886]_ , \new_[3887]_ , \new_[3888]_ ,
    \new_[3889]_ , \new_[3890]_ , \new_[3891]_ , \new_[3892]_ ,
    \new_[3893]_ , \new_[3894]_ , \new_[3895]_ , \new_[3896]_ ,
    \new_[3897]_ , \new_[3898]_ , \new_[3899]_ , \new_[3900]_ ,
    \new_[3901]_ , \new_[3902]_ , \new_[3903]_ , \new_[3904]_ ,
    \new_[3905]_ , \new_[3906]_ , \new_[3907]_ , \new_[3908]_ ,
    \new_[3909]_ , \new_[3910]_ , \new_[3911]_ , \new_[3912]_ ,
    \new_[3913]_ , \new_[3914]_ , \new_[3915]_ , \new_[3916]_ ,
    \new_[3917]_ , \new_[3918]_ , \new_[3919]_ , \new_[3920]_ ,
    \new_[3921]_ , \new_[3922]_ , \new_[3923]_ , \new_[3924]_ ,
    \new_[3925]_ , \new_[3926]_ , \new_[3927]_ , \new_[3928]_ ,
    \new_[3929]_ , \new_[3930]_ , \new_[3931]_ , \new_[3932]_ ,
    \new_[3933]_ , \new_[3934]_ , \new_[3935]_ , \new_[3936]_ ,
    \new_[3937]_ , \new_[3938]_ , \new_[3939]_ , \new_[3940]_ ,
    \new_[3941]_ , \new_[3942]_ , \new_[3943]_ , \new_[3944]_ ,
    \new_[3945]_ , \new_[3946]_ , \new_[3947]_ , \new_[3948]_ ,
    \new_[3949]_ , \new_[3950]_ , \new_[3951]_ , \new_[3952]_ ,
    \new_[3953]_ , \new_[3954]_ , \new_[3955]_ , \new_[3956]_ ,
    \new_[3957]_ , \new_[3958]_ , \new_[3959]_ , \new_[3960]_ ,
    \new_[3961]_ , \new_[3962]_ , \new_[3963]_ , \new_[3964]_ ,
    \new_[3965]_ , \new_[3966]_ , \new_[3967]_ , \new_[3968]_ ,
    \new_[3969]_ , \new_[3970]_ , \new_[3971]_ , \new_[3972]_ ,
    \new_[3973]_ , \new_[3974]_ , \new_[3975]_ , \new_[3976]_ ,
    \new_[3977]_ , \new_[3978]_ , \new_[3979]_ , \new_[3980]_ ,
    \new_[3981]_ , \new_[3982]_ , \new_[3983]_ , \new_[3984]_ ,
    \new_[3985]_ , \new_[3986]_ , \new_[3987]_ , \new_[3988]_ ,
    \new_[3989]_ , \new_[3990]_ , \new_[3991]_ , \new_[3992]_ ,
    \new_[3993]_ , \new_[3994]_ , \new_[3995]_ , \new_[3996]_ ,
    \new_[3997]_ , \new_[3998]_ , \new_[3999]_ , \new_[4000]_ ,
    \new_[4001]_ , \new_[4002]_ , \new_[4003]_ , \new_[4004]_ ,
    \new_[4005]_ , \new_[4006]_ , \new_[4007]_ , \new_[4008]_ ,
    \new_[4009]_ , \new_[4010]_ , \new_[4011]_ , \new_[4012]_ ,
    \new_[4013]_ , \new_[4014]_ , \new_[4015]_ , \new_[4016]_ ,
    \new_[4017]_ , \new_[4018]_ , \new_[4019]_ , \new_[4020]_ ,
    \new_[4021]_ , \new_[4022]_ , \new_[4023]_ , \new_[4024]_ ,
    \new_[4025]_ , \new_[4026]_ , \new_[4027]_ , \new_[4028]_ ,
    \new_[4029]_ , \new_[4030]_ , \new_[4031]_ , \new_[4032]_ ,
    \new_[4033]_ , \new_[4034]_ , \new_[4035]_ , \new_[4036]_ ,
    \new_[4037]_ , \new_[4038]_ , \new_[4039]_ , \new_[4040]_ ,
    \new_[4041]_ , \new_[4042]_ , \new_[4043]_ , \new_[4044]_ ,
    \new_[4045]_ , \new_[4046]_ , \new_[4047]_ , \new_[4048]_ ,
    \new_[4049]_ , \new_[4050]_ , \new_[4051]_ , \new_[4052]_ ,
    \new_[4053]_ , \new_[4054]_ , \new_[4055]_ , \new_[4056]_ ,
    \new_[4057]_ , \new_[4058]_ , \new_[4059]_ , \new_[4060]_ ,
    \new_[4061]_ , \new_[4062]_ , \new_[4063]_ , \new_[4064]_ ,
    \new_[4065]_ , \new_[4066]_ , \new_[4067]_ , \new_[4068]_ ,
    \new_[4069]_ , \new_[4070]_ , \new_[4071]_ , \new_[4072]_ ,
    \new_[4073]_ , \new_[4074]_ , \new_[4075]_ , \new_[4076]_ ,
    \new_[4077]_ , \new_[4078]_ , \new_[4079]_ , \new_[4080]_ ,
    \new_[4081]_ , \new_[4082]_ , \new_[4083]_ , \new_[4084]_ ,
    \new_[4085]_ , \new_[4086]_ , \new_[4087]_ , \new_[4088]_ ,
    \new_[4089]_ , \new_[4090]_ , \new_[4091]_ , \new_[4092]_ ,
    \new_[4093]_ , \new_[4094]_ , \new_[4095]_ , \new_[4096]_ ,
    \new_[4097]_ , \new_[4098]_ , \new_[4099]_ , \new_[4100]_ ,
    \new_[4101]_ , \new_[4102]_ , \new_[4103]_ , \new_[4104]_ ,
    \new_[4105]_ , \new_[4106]_ , \new_[4107]_ , \new_[4108]_ ,
    \new_[4109]_ , \new_[4110]_ , \new_[4111]_ , \new_[4112]_ ,
    \new_[4113]_ , \new_[4114]_ , \new_[4115]_ , \new_[4116]_ ,
    \new_[4117]_ , \new_[4118]_ , \new_[4119]_ , \new_[4120]_ ,
    \new_[4121]_ , \new_[4122]_ , \new_[4123]_ , \new_[4124]_ ,
    \new_[4125]_ , \new_[4126]_ , \new_[4127]_ , \new_[4128]_ ,
    \new_[4129]_ , \new_[4130]_ , \new_[4131]_ , \new_[4132]_ ,
    \new_[4133]_ , \new_[4134]_ , \new_[4135]_ , \new_[4136]_ ,
    \new_[4137]_ , \new_[4138]_ , \new_[4139]_ , \new_[4140]_ ,
    \new_[4141]_ , \new_[4142]_ , \new_[4143]_ , \new_[4144]_ ,
    \new_[4145]_ , \new_[4146]_ , \new_[4147]_ , \new_[4148]_ ,
    \new_[4149]_ , \new_[4150]_ , \new_[4151]_ , \new_[4152]_ ,
    \new_[4153]_ , \new_[4154]_ , \new_[4155]_ , \new_[4156]_ ,
    \new_[4157]_ , \new_[4158]_ , \new_[4159]_ , \new_[4160]_ ,
    \new_[4161]_ , \new_[4162]_ , \new_[4163]_ , \new_[4164]_ ,
    \new_[4165]_ , \new_[4166]_ , \new_[4167]_ , \new_[4168]_ ,
    \new_[4169]_ , \new_[4170]_ , \new_[4171]_ , \new_[4172]_ ,
    \new_[4173]_ , \new_[4174]_ , \new_[4175]_ , \new_[4176]_ ,
    \new_[4177]_ , \new_[4178]_ , \new_[4179]_ , \new_[4180]_ ,
    \new_[4181]_ , \new_[4182]_ , \new_[4183]_ , \new_[4184]_ ,
    \new_[4185]_ , \new_[4186]_ , \new_[4187]_ , \new_[4188]_ ,
    \new_[4189]_ , \new_[4190]_ , \new_[4191]_ , \new_[4192]_ ,
    \new_[4193]_ , \new_[4194]_ , \new_[4195]_ , \new_[4196]_ ,
    \new_[4197]_ , \new_[4198]_ , \new_[4199]_ , \new_[4200]_ ,
    \new_[4201]_ , \new_[4202]_ , \new_[4203]_ , \new_[4204]_ ,
    \new_[4205]_ , \new_[4206]_ , \new_[4207]_ , \new_[4208]_ ,
    \new_[4209]_ , \new_[4210]_ , \new_[4211]_ , \new_[4212]_ ,
    \new_[4213]_ , \new_[4214]_ , \new_[4215]_ , \new_[4216]_ ,
    \new_[4217]_ , \new_[4218]_ , \new_[4219]_ , \new_[4220]_ ,
    \new_[4221]_ , \new_[4222]_ , \new_[4223]_ , \new_[4224]_ ,
    \new_[4225]_ , \new_[4226]_ , \new_[4227]_ , \new_[4228]_ ,
    \new_[4229]_ , \new_[4230]_ , \new_[4231]_ , \new_[4232]_ ,
    \new_[4233]_ , \new_[4234]_ , \new_[4235]_ , \new_[4236]_ ,
    \new_[4237]_ , \new_[4238]_ , \new_[4239]_ , \new_[4240]_ ,
    \new_[4241]_ , \new_[4242]_ , \new_[4243]_ , \new_[4244]_ ,
    \new_[4245]_ , \new_[4246]_ , \new_[4247]_ , \new_[4248]_ ,
    \new_[4249]_ , \new_[4250]_ , \new_[4251]_ , \new_[4252]_ ,
    \new_[4253]_ , \new_[4254]_ , \new_[4255]_ , \new_[4256]_ ,
    \new_[4257]_ , \new_[4258]_ , \new_[4259]_ , \new_[4260]_ ,
    \new_[4261]_ , \new_[4262]_ , \new_[4263]_ , \new_[4264]_ ,
    \new_[4265]_ , \new_[4266]_ , \new_[4267]_ , \new_[4268]_ ,
    \new_[4269]_ , \new_[4270]_ , \new_[4271]_ , \new_[4272]_ ,
    \new_[4273]_ , \new_[4274]_ , \new_[4275]_ , \new_[4276]_ ,
    \new_[4277]_ , \new_[4278]_ , \new_[4279]_ , \new_[4280]_ ,
    \new_[4281]_ , \new_[4282]_ , \new_[4283]_ , \new_[4284]_ ,
    \new_[4285]_ , \new_[4286]_ , \new_[4287]_ , \new_[4288]_ ,
    \new_[4289]_ , \new_[4290]_ , \new_[4291]_ , \new_[4292]_ ,
    \new_[4293]_ , \new_[4294]_ , \new_[4295]_ , \new_[4296]_ ,
    \new_[4297]_ , \new_[4298]_ , \new_[4299]_ , \new_[4300]_ ,
    \new_[4301]_ , \new_[4302]_ , \new_[4303]_ , \new_[4304]_ ,
    \new_[4305]_ , \new_[4306]_ , \new_[4307]_ , \new_[4308]_ ,
    \new_[4309]_ , \new_[4310]_ , \new_[4311]_ , \new_[4312]_ ,
    \new_[4313]_ , \new_[4314]_ , \new_[4315]_ , \new_[4316]_ ,
    \new_[4317]_ , \new_[4318]_ , \new_[4319]_ , \new_[4320]_ ,
    \new_[4321]_ , \new_[4322]_ , \new_[4323]_ , \new_[4324]_ ,
    \new_[4325]_ , \new_[4326]_ , \new_[4327]_ , \new_[4328]_ ,
    \new_[4329]_ , \new_[4330]_ , \new_[4331]_ , \new_[4332]_ ,
    \new_[4333]_ , \new_[4334]_ , \new_[4335]_ , \new_[4336]_ ,
    \new_[4337]_ , \new_[4338]_ , \new_[4339]_ , \new_[4340]_ ,
    \new_[4341]_ , \new_[4342]_ , \new_[4343]_ , \new_[4344]_ ,
    \new_[4345]_ , \new_[4346]_ , \new_[4347]_ , \new_[4348]_ ,
    \new_[4349]_ , \new_[4350]_ , \new_[4351]_ , \new_[4352]_ ,
    \new_[4353]_ , \new_[4354]_ , \new_[4355]_ , \new_[4356]_ ,
    \new_[4357]_ , \new_[4358]_ , \new_[4359]_ , \new_[4360]_ ,
    \new_[4361]_ , \new_[4362]_ , \new_[4363]_ , \new_[4364]_ ,
    \new_[4365]_ , \new_[4366]_ , \new_[4367]_ , \new_[4368]_ ,
    \new_[4369]_ , \new_[4370]_ , \new_[4371]_ , \new_[4372]_ ,
    \new_[4373]_ , \new_[4374]_ , \new_[4375]_ , \new_[4376]_ ,
    \new_[4377]_ , \new_[4378]_ , \new_[4379]_ , \new_[4380]_ ,
    \new_[4381]_ , \new_[4382]_ , \new_[4383]_ , \new_[4384]_ ,
    \new_[4385]_ , \new_[4386]_ , \new_[4387]_ , \new_[4388]_ ,
    \new_[4389]_ , \new_[4390]_ , \new_[4391]_ , \new_[4392]_ ,
    \new_[4393]_ , \new_[4394]_ , \new_[4395]_ , \new_[4396]_ ,
    \new_[4397]_ , \new_[4398]_ , \new_[4399]_ , \new_[4400]_ ,
    \new_[4401]_ , \new_[4402]_ , \new_[4403]_ , \new_[4404]_ ,
    \new_[4405]_ , \new_[4406]_ , \new_[4407]_ , \new_[4408]_ ,
    \new_[4409]_ , \new_[4410]_ , \new_[4411]_ , \new_[4412]_ ,
    \new_[4413]_ , \new_[4414]_ , \new_[4415]_ , \new_[4416]_ ,
    \new_[4417]_ , \new_[4418]_ , \new_[4419]_ , \new_[4420]_ ,
    \new_[4421]_ , \new_[4422]_ , \new_[4423]_ , \new_[4424]_ ,
    \new_[4425]_ , \new_[4426]_ , \new_[4427]_ , \new_[4428]_ ,
    \new_[4429]_ , \new_[4430]_ , \new_[4431]_ , \new_[4432]_ ,
    \new_[4433]_ , \new_[4434]_ , \new_[4435]_ , \new_[4436]_ ,
    \new_[4437]_ , \new_[4438]_ , \new_[4439]_ , \new_[4440]_ ,
    \new_[4441]_ , \new_[4442]_ , \new_[4443]_ , \new_[4444]_ ,
    \new_[4445]_ , \new_[4446]_ , \new_[4447]_ , \new_[4448]_ ,
    \new_[4449]_ , \new_[4450]_ , \new_[4451]_ , \new_[4452]_ ,
    \new_[4453]_ , \new_[4454]_ , \new_[4455]_ , \new_[4456]_ ,
    \new_[4457]_ , \new_[4458]_ , \new_[4459]_ , \new_[4460]_ ,
    \new_[4461]_ , \new_[4462]_ , \new_[4463]_ , \new_[4464]_ ,
    \new_[4465]_ , \new_[4466]_ , \new_[4467]_ , \new_[4468]_ ,
    \new_[4469]_ , \new_[4470]_ , \new_[4471]_ , \new_[4472]_ ,
    \new_[4473]_ , \new_[4474]_ , \new_[4475]_ , \new_[4476]_ ,
    \new_[4477]_ , \new_[4478]_ , \new_[4479]_ , \new_[4480]_ ,
    \new_[4481]_ , \new_[4482]_ , \new_[4483]_ , \new_[4484]_ ,
    \new_[4485]_ , \new_[4486]_ , \new_[4487]_ , \new_[4488]_ ,
    \new_[4489]_ , \new_[4490]_ , \new_[4491]_ , \new_[4492]_ ,
    \new_[4493]_ , \new_[4494]_ , \new_[4495]_ , \new_[4496]_ ,
    \new_[4497]_ , \new_[4498]_ , \new_[4499]_ , \new_[4500]_ ,
    \new_[4501]_ , \new_[4502]_ , \new_[4503]_ , \new_[4504]_ ,
    \new_[4505]_ , \new_[4506]_ , \new_[4507]_ , \new_[4508]_ ,
    \new_[4509]_ , \new_[4510]_ , \new_[4511]_ , \new_[4512]_ ,
    \new_[4513]_ , \new_[4514]_ , \new_[4515]_ , \new_[4516]_ ,
    \new_[4517]_ , \new_[4518]_ , \new_[4519]_ , \new_[4520]_ ,
    \new_[4521]_ , \new_[4522]_ , \new_[4523]_ , \new_[4524]_ ,
    \new_[4525]_ , \new_[4526]_ , \new_[4527]_ , \new_[4528]_ ,
    \new_[4529]_ , \new_[4530]_ , \new_[4531]_ , \new_[4532]_ ,
    \new_[4533]_ , \new_[4534]_ , \new_[4535]_ , \new_[4536]_ ,
    \new_[4537]_ , \new_[4538]_ , \new_[4539]_ , \new_[4540]_ ,
    \new_[4541]_ , \new_[4542]_ , \new_[4543]_ , \new_[4544]_ ,
    \new_[4545]_ , \new_[4546]_ , \new_[4547]_ , \new_[4548]_ ,
    \new_[4549]_ , \new_[4550]_ , \new_[4551]_ , \new_[4552]_ ,
    \new_[4553]_ , \new_[4554]_ , \new_[4555]_ , \new_[4556]_ ,
    \new_[4557]_ , \new_[4558]_ , \new_[4559]_ , \new_[4560]_ ,
    \new_[4561]_ , \new_[4562]_ , \new_[4563]_ , \new_[4564]_ ,
    \new_[4565]_ , \new_[4566]_ , \new_[4567]_ , \new_[4568]_ ,
    \new_[4569]_ , \new_[4570]_ , \new_[4571]_ , \new_[4572]_ ,
    \new_[4573]_ , \new_[4574]_ , \new_[4575]_ , \new_[4576]_ ,
    \new_[4577]_ , \new_[4578]_ , \new_[4579]_ , \new_[4580]_ ,
    \new_[4581]_ , \new_[4582]_ , \new_[4583]_ , \new_[4584]_ ,
    \new_[4585]_ , \new_[4586]_ , \new_[4587]_ , \new_[4588]_ ,
    \new_[4589]_ , \new_[4590]_ , \new_[4591]_ , \new_[4592]_ ,
    \new_[4593]_ , \new_[4594]_ , \new_[4595]_ , \new_[4596]_ ,
    \new_[4597]_ , \new_[4598]_ , \new_[4599]_ , \new_[4600]_ ,
    \new_[4601]_ , \new_[4602]_ , \new_[4603]_ , \new_[4604]_ ,
    \new_[4605]_ , \new_[4606]_ , \new_[4607]_ , \new_[4608]_ ,
    \new_[4609]_ , \new_[4610]_ , \new_[4611]_ , \new_[4612]_ ,
    \new_[4613]_ , \new_[4614]_ , \new_[4615]_ , \new_[4616]_ ,
    \new_[4617]_ , \new_[4618]_ , \new_[4619]_ , \new_[4620]_ ,
    \new_[4621]_ , \new_[4622]_ , \new_[4623]_ , \new_[4624]_ ,
    \new_[4625]_ , \new_[4626]_ , \new_[4627]_ , \new_[4628]_ ,
    \new_[4629]_ , \new_[4630]_ , \new_[4631]_ , \new_[4632]_ ,
    \new_[4633]_ , \new_[4634]_ , \new_[4635]_ , \new_[4636]_ ,
    \new_[4637]_ , \new_[4638]_ , \new_[4639]_ , \new_[4640]_ ,
    \new_[4641]_ , \new_[4642]_ , \new_[4643]_ , \new_[4644]_ ,
    \new_[4645]_ , \new_[4646]_ , \new_[4647]_ , \new_[4648]_ ,
    \new_[4649]_ , \new_[4650]_ , \new_[4651]_ , \new_[4652]_ ,
    \new_[4653]_ , \new_[4654]_ , \new_[4655]_ , \new_[4656]_ ,
    \new_[4657]_ , \new_[4658]_ , \new_[4659]_ , \new_[4660]_ ,
    \new_[4661]_ , \new_[4662]_ , \new_[4663]_ , \new_[4664]_ ,
    \new_[4665]_ , \new_[4666]_ , \new_[4667]_ , \new_[4668]_ ,
    \new_[4669]_ , \new_[4670]_ , \new_[4671]_ , \new_[4672]_ ,
    \new_[4673]_ , \new_[4674]_ , \new_[4675]_ , \new_[4676]_ ,
    \new_[4677]_ , \new_[4678]_ , \new_[4679]_ , \new_[4680]_ ,
    \new_[4681]_ , \new_[4682]_ , \new_[4683]_ , \new_[4684]_ ,
    \new_[4685]_ , \new_[4686]_ , \new_[4687]_ , \new_[4688]_ ,
    \new_[4689]_ , \new_[4690]_ , \new_[4691]_ , \new_[4692]_ ,
    \new_[4693]_ , \new_[4694]_ , \new_[4695]_ , \new_[4696]_ ,
    \new_[4697]_ , \new_[4698]_ , \new_[4699]_ , \new_[4700]_ ,
    \new_[4701]_ , \new_[4702]_ , \new_[4703]_ , \new_[4704]_ ,
    \new_[4705]_ , \new_[4706]_ , \new_[4707]_ , \new_[4708]_ ,
    \new_[4709]_ , \new_[4710]_ , \new_[4711]_ , \new_[4712]_ ,
    \new_[4713]_ , \new_[4714]_ , \new_[4715]_ , \new_[4716]_ ,
    \new_[4717]_ , \new_[4718]_ , \new_[4719]_ , \new_[4720]_ ,
    \new_[4721]_ , \new_[4722]_ , \new_[4723]_ , \new_[4724]_ ,
    \new_[4725]_ , \new_[4726]_ , \new_[4727]_ , \new_[4728]_ ,
    \new_[4729]_ , \new_[4730]_ , \new_[4731]_ , \new_[4732]_ ,
    \new_[4733]_ , \new_[4734]_ , \new_[4735]_ , \new_[4736]_ ,
    \new_[4737]_ , \new_[4738]_ , \new_[4739]_ , \new_[4740]_ ,
    \new_[4741]_ , \new_[4742]_ , \new_[4743]_ , \new_[4744]_ ,
    \new_[4745]_ , \new_[4746]_ , \new_[4747]_ , \new_[4748]_ ,
    \new_[4749]_ , \new_[4750]_ , \new_[4751]_ , \new_[4752]_ ,
    \new_[4753]_ , \new_[4754]_ , \new_[4755]_ , \new_[4756]_ ,
    \new_[4757]_ , \new_[4758]_ , \new_[4759]_ , \new_[4760]_ ,
    \new_[4761]_ , \new_[4762]_ , \new_[4763]_ , \new_[4764]_ ,
    \new_[4765]_ , \new_[4766]_ , \new_[4767]_ , \new_[4768]_ ,
    \new_[4769]_ , \new_[4770]_ , \new_[4771]_ , \new_[4772]_ ,
    \new_[4773]_ , \new_[4774]_ , \new_[4775]_ , \new_[4776]_ ,
    \new_[4777]_ , \new_[4778]_ , \new_[4779]_ , \new_[4780]_ ,
    \new_[4781]_ , \new_[4782]_ , \new_[4783]_ , \new_[4784]_ ,
    \new_[4785]_ , \new_[4786]_ , \new_[4787]_ , \new_[4788]_ ,
    \new_[4789]_ , \new_[4790]_ , \new_[4791]_ , \new_[4792]_ ,
    \new_[4793]_ , \new_[4794]_ , \new_[4795]_ , \new_[4796]_ ,
    \new_[4797]_ , \new_[4798]_ , \new_[4799]_ , \new_[4800]_ ,
    \new_[4801]_ , \new_[4802]_ , \new_[4803]_ , \new_[4804]_ ,
    \new_[4805]_ , \new_[4806]_ , \new_[4807]_ , \new_[4808]_ ,
    \new_[4809]_ , \new_[4810]_ , \new_[4811]_ , \new_[4812]_ ,
    \new_[4813]_ , \new_[4814]_ , \new_[4815]_ , \new_[4816]_ ,
    \new_[4817]_ , \new_[4818]_ , \new_[4819]_ , \new_[4820]_ ,
    \new_[4821]_ , \new_[4822]_ , \new_[4823]_ , \new_[4824]_ ,
    \new_[4825]_ , \new_[4826]_ , \new_[4827]_ , \new_[4828]_ ,
    \new_[4829]_ , \new_[4830]_ , \new_[4831]_ , \new_[4832]_ ,
    \new_[4833]_ , \new_[4834]_ , \new_[4835]_ , \new_[4836]_ ,
    \new_[4837]_ , \new_[4838]_ , \new_[4839]_ , \new_[4840]_ ,
    \new_[4841]_ , \new_[4842]_ , \new_[4843]_ , \new_[4844]_ ,
    \new_[4845]_ , \new_[4846]_ , \new_[4847]_ , \new_[4848]_ ,
    \new_[4849]_ , \new_[4850]_ , \new_[4851]_ , \new_[4852]_ ,
    \new_[4853]_ , \new_[4854]_ , \new_[4855]_ , \new_[4856]_ ,
    \new_[4857]_ , \new_[4858]_ , \new_[4859]_ , \new_[4860]_ ,
    \new_[4861]_ , \new_[4862]_ , \new_[4863]_ , \new_[4864]_ ,
    \new_[4865]_ , \new_[4866]_ , \new_[4867]_ , \new_[4868]_ ,
    \new_[4869]_ , \new_[4870]_ , \new_[4871]_ , \new_[4872]_ ,
    \new_[4873]_ , \new_[4874]_ , \new_[4875]_ , \new_[4876]_ ,
    \new_[4877]_ , \new_[4878]_ , \new_[4879]_ , \new_[4880]_ ,
    \new_[4881]_ , \new_[4882]_ , \new_[4883]_ , \new_[4884]_ ,
    \new_[4885]_ , \new_[4886]_ , \new_[4887]_ , \new_[4888]_ ,
    \new_[4889]_ , \new_[4890]_ , \new_[4891]_ , \new_[4892]_ ,
    \new_[4893]_ , \new_[4894]_ , \new_[4895]_ , \new_[4896]_ ,
    \new_[4897]_ , \new_[4898]_ , \new_[4899]_ , \new_[4900]_ ,
    \new_[4901]_ , \new_[4902]_ , \new_[4903]_ , \new_[4904]_ ,
    \new_[4905]_ , \new_[4906]_ , \new_[4907]_ , \new_[4908]_ ,
    \new_[4909]_ , \new_[4910]_ , \new_[4911]_ , \new_[4912]_ ,
    \new_[4913]_ , \new_[4914]_ , \new_[4915]_ , \new_[4916]_ ,
    \new_[4917]_ , \new_[4918]_ , \new_[4919]_ , \new_[4920]_ ,
    \new_[4921]_ , \new_[4922]_ , \new_[4923]_ , \new_[4924]_ ,
    \new_[4925]_ , \new_[4926]_ , \new_[4927]_ , \new_[4928]_ ,
    \new_[4929]_ , \new_[4930]_ , \new_[4931]_ , \new_[4932]_ ,
    \new_[4933]_ , \new_[4934]_ , \new_[4935]_ , \new_[4936]_ ,
    \new_[4937]_ , \new_[4938]_ , \new_[4939]_ , \new_[4940]_ ,
    \new_[4941]_ , \new_[4942]_ , \new_[4943]_ , \new_[4944]_ ,
    \new_[4945]_ , \new_[4946]_ , \new_[4947]_ , \new_[4948]_ ,
    \new_[4949]_ , \new_[4950]_ , \new_[4951]_ , \new_[4952]_ ,
    \new_[4953]_ , \new_[4954]_ , \new_[4955]_ , \new_[4956]_ ,
    \new_[4957]_ , \new_[4958]_ , \new_[4959]_ , \new_[4960]_ ,
    \new_[4961]_ , \new_[4962]_ , \new_[4963]_ , \new_[4964]_ ,
    \new_[4965]_ , \new_[4966]_ , \new_[4967]_ , \new_[4968]_ ,
    \new_[4969]_ , \new_[4970]_ , \new_[4971]_ , \new_[4972]_ ,
    \new_[4973]_ , \new_[4974]_ , \new_[4975]_ , \new_[4976]_ ,
    \new_[4977]_ , \new_[4978]_ , \new_[4979]_ , \new_[4980]_ ,
    \new_[4981]_ , \new_[4982]_ , \new_[4983]_ , \new_[4984]_ ,
    \new_[4985]_ , \new_[4986]_ , \new_[4987]_ , \new_[4988]_ ,
    \new_[4989]_ , \new_[4990]_ , \new_[4991]_ , \new_[4992]_ ,
    \new_[4993]_ , \new_[4994]_ , \new_[4995]_ , \new_[4996]_ ,
    \new_[4997]_ , \new_[4998]_ , \new_[4999]_ , \new_[5000]_ ,
    \new_[5001]_ , \new_[5002]_ , \new_[5003]_ , \new_[5004]_ ,
    \new_[5005]_ , \new_[5006]_ , \new_[5007]_ , \new_[5008]_ ,
    \new_[5009]_ , \new_[5010]_ , \new_[5011]_ , \new_[5012]_ ,
    \new_[5013]_ , \new_[5014]_ , \new_[5015]_ , \new_[5016]_ ,
    \new_[5017]_ , \new_[5018]_ , \new_[5019]_ , \new_[5020]_ ,
    \new_[5021]_ , \new_[5022]_ , \new_[5023]_ , \new_[5024]_ ,
    \new_[5025]_ , \new_[5026]_ , \new_[5027]_ , \new_[5028]_ ,
    \new_[5029]_ , \new_[5030]_ , \new_[5031]_ , \new_[5032]_ ,
    \new_[5033]_ , \new_[5034]_ , \new_[5035]_ , \new_[5036]_ ,
    \new_[5037]_ , \new_[5038]_ , \new_[5039]_ , \new_[5040]_ ,
    \new_[5041]_ , \new_[5042]_ , \new_[5043]_ , \new_[5044]_ ,
    \new_[5045]_ , \new_[5046]_ , \new_[5047]_ , \new_[5048]_ ,
    \new_[5049]_ , \new_[5050]_ , \new_[5051]_ , \new_[5052]_ ,
    \new_[5053]_ , \new_[5054]_ , \new_[5055]_ , \new_[5056]_ ,
    \new_[5057]_ , \new_[5058]_ , \new_[5059]_ , \new_[5060]_ ,
    \new_[5061]_ , \new_[5062]_ , \new_[5063]_ , \new_[5064]_ ,
    \new_[5065]_ , \new_[5066]_ , \new_[5067]_ , \new_[5068]_ ,
    \new_[5069]_ , \new_[5070]_ , \new_[5071]_ , \new_[5072]_ ,
    \new_[5073]_ , \new_[5074]_ , \new_[5075]_ , \new_[5076]_ ,
    \new_[5077]_ , \new_[5078]_ , \new_[5079]_ , \new_[5080]_ ,
    \new_[5081]_ , \new_[5082]_ , \new_[5083]_ , \new_[5084]_ ,
    \new_[5085]_ , \new_[5086]_ , \new_[5087]_ , \new_[5088]_ ,
    \new_[5089]_ , \new_[5090]_ , \new_[5091]_ , \new_[5092]_ ,
    \new_[5093]_ , \new_[5094]_ , \new_[5095]_ , \new_[5096]_ ,
    \new_[5097]_ , \new_[5098]_ , \new_[5099]_ , \new_[5100]_ ,
    \new_[5101]_ , \new_[5102]_ , \new_[5103]_ , \new_[5104]_ ,
    \new_[5105]_ , \new_[5106]_ , \new_[5107]_ , \new_[5108]_ ,
    \new_[5109]_ , \new_[5110]_ , \new_[5111]_ , \new_[5112]_ ,
    \new_[5113]_ , \new_[5114]_ , \new_[5115]_ , \new_[5116]_ ,
    \new_[5117]_ , \new_[5118]_ , \new_[5119]_ , \new_[5120]_ ,
    \new_[5121]_ , \new_[5122]_ , \new_[5123]_ , \new_[5124]_ ,
    \new_[5125]_ , \new_[5126]_ , \new_[5127]_ , \new_[5128]_ ,
    \new_[5129]_ , \new_[5130]_ , \new_[5131]_ , \new_[5132]_ ,
    \new_[5133]_ , \new_[5134]_ , \new_[5135]_ , \new_[5136]_ ,
    \new_[5137]_ , \new_[5138]_ , \new_[5139]_ , \new_[5140]_ ,
    \new_[5141]_ , \new_[5142]_ , \new_[5143]_ , \new_[5144]_ ,
    \new_[5145]_ , \new_[5146]_ , \new_[5147]_ , \new_[5148]_ ,
    \new_[5149]_ , \new_[5150]_ , \new_[5151]_ , \new_[5152]_ ,
    \new_[5153]_ , \new_[5154]_ , \new_[5155]_ , \new_[5156]_ ,
    \new_[5157]_ , \new_[5158]_ , \new_[5159]_ , \new_[5160]_ ,
    \new_[5161]_ , \new_[5162]_ , \new_[5163]_ , \new_[5164]_ ,
    \new_[5165]_ , \new_[5166]_ , \new_[5167]_ , \new_[5168]_ ,
    \new_[5169]_ , \new_[5170]_ , \new_[5171]_ , \new_[5172]_ ,
    \new_[5173]_ , \new_[5174]_ , \new_[5175]_ , \new_[5176]_ ,
    \new_[5177]_ , \new_[5178]_ , \new_[5179]_ , \new_[5180]_ ,
    \new_[5181]_ , \new_[5182]_ , \new_[5183]_ , \new_[5184]_ ,
    \new_[5185]_ , \new_[5186]_ , \new_[5187]_ , \new_[5188]_ ,
    \new_[5189]_ , \new_[5190]_ , \new_[5191]_ , \new_[5192]_ ,
    \new_[5193]_ , \new_[5194]_ , \new_[5195]_ , \new_[5196]_ ,
    \new_[5197]_ , \new_[5198]_ , \new_[5199]_ , \new_[5200]_ ,
    \new_[5201]_ , \new_[5202]_ , \new_[5203]_ , \new_[5204]_ ,
    \new_[5205]_ , \new_[5206]_ , \new_[5207]_ , \new_[5208]_ ,
    \new_[5209]_ , \new_[5210]_ , \new_[5211]_ , \new_[5212]_ ,
    \new_[5213]_ , \new_[5214]_ , \new_[5215]_ , \new_[5216]_ ,
    \new_[5217]_ , \new_[5218]_ , \new_[5219]_ , \new_[5220]_ ,
    \new_[5221]_ , \new_[5222]_ , \new_[5223]_ , \new_[5224]_ ,
    \new_[5225]_ , \new_[5226]_ , \new_[5227]_ , \new_[5228]_ ,
    \new_[5229]_ , \new_[5230]_ , \new_[5231]_ , \new_[5232]_ ,
    \new_[5233]_ , \new_[5234]_ , \new_[5235]_ , \new_[5236]_ ,
    \new_[5237]_ , \new_[5238]_ , \new_[5239]_ , \new_[5240]_ ,
    \new_[5241]_ , \new_[5242]_ , \new_[5243]_ , \new_[5244]_ ,
    \new_[5245]_ , \new_[5246]_ , \new_[5247]_ , \new_[5248]_ ,
    \new_[5249]_ , \new_[5250]_ , \new_[5251]_ , \new_[5252]_ ,
    \new_[5253]_ , \new_[5254]_ , \new_[5255]_ , \new_[5256]_ ,
    \new_[5257]_ , \new_[5258]_ , \new_[5259]_ , \new_[5260]_ ,
    \new_[5261]_ , \new_[5262]_ , \new_[5263]_ , \new_[5264]_ ,
    \new_[5265]_ , \new_[5266]_ , \new_[5267]_ , \new_[5268]_ ,
    \new_[5269]_ , \new_[5270]_ , \new_[5271]_ , \new_[5272]_ ,
    \new_[5273]_ , \new_[5274]_ , \new_[5275]_ , \new_[5276]_ ,
    \new_[5277]_ , \new_[5278]_ , \new_[5279]_ , \new_[5280]_ ,
    \new_[5281]_ , \new_[5282]_ , \new_[5283]_ , \new_[5284]_ ,
    \new_[5285]_ , \new_[5286]_ , \new_[5287]_ , \new_[5288]_ ,
    \new_[5289]_ , \new_[5290]_ , \new_[5291]_ , \new_[5292]_ ,
    \new_[5293]_ , \new_[5294]_ , \new_[5295]_ , \new_[5296]_ ,
    \new_[5297]_ , \new_[5298]_ , \new_[5299]_ , \new_[5300]_ ,
    \new_[5301]_ , \new_[5302]_ , \new_[5303]_ , \new_[5304]_ ,
    \new_[5305]_ , \new_[5306]_ , \new_[5307]_ , \new_[5308]_ ,
    \new_[5309]_ , \new_[5310]_ , \new_[5311]_ , \new_[5312]_ ,
    \new_[5313]_ , \new_[5314]_ , \new_[5315]_ , \new_[5316]_ ,
    \new_[5317]_ , \new_[5318]_ , \new_[5319]_ , \new_[5320]_ ,
    \new_[5321]_ , \new_[5322]_ , \new_[5323]_ , \new_[5324]_ ,
    \new_[5325]_ , \new_[5326]_ , \new_[5327]_ , \new_[5328]_ ,
    \new_[5329]_ , \new_[5330]_ , \new_[5331]_ , \new_[5332]_ ,
    \new_[5333]_ , \new_[5334]_ , \new_[5335]_ , \new_[5336]_ ,
    \new_[5337]_ , \new_[5338]_ , \new_[5339]_ , \new_[5340]_ ,
    \new_[5341]_ , \new_[5342]_ , \new_[5343]_ , \new_[5344]_ ,
    \new_[5345]_ , \new_[5346]_ , \new_[5347]_ , \new_[5348]_ ,
    \new_[5349]_ , \new_[5350]_ , \new_[5351]_ , \new_[5352]_ ,
    \new_[5353]_ , \new_[5354]_ , \new_[5355]_ , \new_[5356]_ ,
    \new_[5357]_ , \new_[5358]_ , \new_[5359]_ , \new_[5360]_ ,
    \new_[5361]_ , \new_[5362]_ , \new_[5363]_ , \new_[5364]_ ,
    \new_[5365]_ , \new_[5366]_ , \new_[5367]_ , \new_[5368]_ ,
    \new_[5369]_ , \new_[5370]_ , \new_[5371]_ , \new_[5372]_ ,
    \new_[5373]_ , \new_[5374]_ , \new_[5375]_ , \new_[5376]_ ,
    \new_[5377]_ , \new_[5378]_ , \new_[5379]_ , \new_[5380]_ ,
    \new_[5381]_ , \new_[5382]_ , \new_[5383]_ , \new_[5384]_ ,
    \new_[5385]_ , \new_[5386]_ , \new_[5387]_ , \new_[5388]_ ,
    \new_[5389]_ , \new_[5390]_ , \new_[5391]_ , \new_[5392]_ ,
    \new_[5393]_ , \new_[5394]_ , \new_[5395]_ , \new_[5396]_ ,
    \new_[5397]_ , \new_[5398]_ , \new_[5399]_ , \new_[5400]_ ,
    \new_[5401]_ , \new_[5402]_ , \new_[5403]_ , \new_[5404]_ ,
    \new_[5405]_ , \new_[5406]_ , \new_[5407]_ , \new_[5408]_ ,
    \new_[5409]_ , \new_[5410]_ , \new_[5411]_ , \new_[5412]_ ,
    \new_[5413]_ , \new_[5414]_ , \new_[5415]_ , \new_[5416]_ ,
    \new_[5417]_ , \new_[5418]_ , \new_[5419]_ , \new_[5420]_ ,
    \new_[5421]_ , \new_[5422]_ , \new_[5423]_ , \new_[5424]_ ,
    \new_[5425]_ , \new_[5426]_ , \new_[5427]_ , \new_[5428]_ ,
    \new_[5429]_ , \new_[5430]_ , \new_[5431]_ , \new_[5432]_ ,
    \new_[5433]_ , \new_[5434]_ , \new_[5435]_ , \new_[5436]_ ,
    \new_[5437]_ , \new_[5438]_ , \new_[5439]_ , \new_[5440]_ ,
    \new_[5441]_ , \new_[5442]_ , \new_[5443]_ , \new_[5444]_ ,
    \new_[5445]_ , \new_[5446]_ , \new_[5447]_ , \new_[5448]_ ,
    \new_[5449]_ , \new_[5450]_ , \new_[5451]_ , \new_[5452]_ ,
    \new_[5453]_ , \new_[5454]_ , \new_[5455]_ , \new_[5456]_ ,
    \new_[5457]_ , \new_[5458]_ , \new_[5459]_ , \new_[5460]_ ,
    \new_[5461]_ , \new_[5462]_ , \new_[5463]_ , \new_[5464]_ ,
    \new_[5465]_ , \new_[5466]_ , \new_[5467]_ , \new_[5468]_ ,
    \new_[5469]_ , \new_[5470]_ , \new_[5471]_ , \new_[5472]_ ,
    \new_[5473]_ , \new_[5474]_ , \new_[5475]_ , \new_[5476]_ ,
    \new_[5477]_ , \new_[5478]_ , \new_[5479]_ , \new_[5480]_ ,
    \new_[5481]_ , \new_[5482]_ , \new_[5483]_ , \new_[5484]_ ,
    \new_[5485]_ , \new_[5486]_ , \new_[5487]_ , \new_[5488]_ ,
    \new_[5489]_ , \new_[5490]_ , \new_[5491]_ , \new_[5492]_ ,
    \new_[5493]_ , \new_[5494]_ , \new_[5495]_ , \new_[5496]_ ,
    \new_[5497]_ , \new_[5498]_ , \new_[5499]_ , \new_[5500]_ ,
    \new_[5501]_ , \new_[5502]_ , \new_[5503]_ , \new_[5504]_ ,
    \new_[5505]_ , \new_[5506]_ , \new_[5507]_ , \new_[5508]_ ,
    \new_[5509]_ , \new_[5510]_ , \new_[5511]_ , \new_[5512]_ ,
    \new_[5513]_ , \new_[5514]_ , \new_[5515]_ , \new_[5516]_ ,
    \new_[5517]_ , \new_[5518]_ , \new_[5519]_ , \new_[5520]_ ,
    \new_[5521]_ , \new_[5522]_ , \new_[5523]_ , \new_[5524]_ ,
    \new_[5525]_ , \new_[5526]_ , \new_[5527]_ , \new_[5528]_ ,
    \new_[5529]_ , \new_[5530]_ , \new_[5531]_ , \new_[5532]_ ,
    \new_[5533]_ , \new_[5534]_ , \new_[5535]_ , \new_[5536]_ ,
    \new_[5537]_ , \new_[5538]_ , \new_[5539]_ , \new_[5540]_ ,
    \new_[5541]_ , \new_[5542]_ , \new_[5543]_ , \new_[5544]_ ,
    \new_[5545]_ , \new_[5546]_ , \new_[5547]_ , \new_[5548]_ ,
    \new_[5549]_ , \new_[5550]_ , \new_[5551]_ , \new_[5552]_ ,
    \new_[5553]_ , \new_[5554]_ , \new_[5555]_ , \new_[5556]_ ,
    \new_[5557]_ , \new_[5558]_ , \new_[5559]_ , \new_[5560]_ ,
    \new_[5561]_ , \new_[5562]_ , \new_[5563]_ , \new_[5564]_ ,
    \new_[5565]_ , \new_[5566]_ , \new_[5567]_ , \new_[5568]_ ,
    \new_[5569]_ , \new_[5570]_ , \new_[5571]_ , \new_[5572]_ ,
    \new_[5573]_ , \new_[5574]_ , \new_[5575]_ , \new_[5576]_ ,
    \new_[5577]_ , \new_[5578]_ , \new_[5579]_ , \new_[5580]_ ,
    \new_[5581]_ , \new_[5582]_ , \new_[5583]_ , \new_[5584]_ ,
    \new_[5585]_ , \new_[5586]_ , \new_[5587]_ , \new_[5588]_ ,
    \new_[5589]_ , \new_[5590]_ , \new_[5591]_ , \new_[5592]_ ,
    \new_[5593]_ , \new_[5594]_ , \new_[5595]_ , \new_[5596]_ ,
    \new_[5597]_ , \new_[5598]_ , \new_[5599]_ , \new_[5600]_ ,
    \new_[5601]_ , \new_[5602]_ , \new_[5603]_ , \new_[5604]_ ,
    \new_[5605]_ , \new_[5606]_ , \new_[5607]_ , \new_[5608]_ ,
    \new_[5609]_ , \new_[5610]_ , \new_[5611]_ , \new_[5612]_ ,
    \new_[5613]_ , \new_[5614]_ , \new_[5615]_ , \new_[5616]_ ,
    \new_[5617]_ , \new_[5618]_ , \new_[5619]_ , \new_[5620]_ ,
    \new_[5621]_ , \new_[5622]_ , \new_[5623]_ , \new_[5624]_ ,
    \new_[5625]_ , \new_[5626]_ , \new_[5627]_ , \new_[5628]_ ,
    \new_[5629]_ , \new_[5630]_ , \new_[5631]_ , \new_[5632]_ ,
    \new_[5633]_ , \new_[5634]_ , \new_[5635]_ , \new_[5636]_ ,
    \new_[5637]_ , \new_[5638]_ , \new_[5639]_ , \new_[5640]_ ,
    \new_[5641]_ , \new_[5642]_ , \new_[5643]_ , \new_[5644]_ ,
    \new_[5645]_ , \new_[5646]_ , \new_[5647]_ , \new_[5648]_ ,
    \new_[5649]_ , \new_[5650]_ , \new_[5651]_ , \new_[5652]_ ,
    \new_[5653]_ , \new_[5654]_ , \new_[5655]_ , \new_[5656]_ ,
    \new_[5657]_ , \new_[5658]_ , \new_[5659]_ , \new_[5660]_ ,
    \new_[5661]_ , \new_[5662]_ , \new_[5663]_ , \new_[5664]_ ,
    \new_[5665]_ , \new_[5666]_ , \new_[5667]_ , \new_[5668]_ ,
    \new_[5669]_ , \new_[5670]_ , \new_[5671]_ , \new_[5672]_ ,
    \new_[5673]_ , \new_[5674]_ , \new_[5675]_ , \new_[5676]_ ,
    \new_[5677]_ , \new_[5678]_ , \new_[5679]_ , \new_[5680]_ ,
    \new_[5681]_ , \new_[5682]_ , \new_[5683]_ , \new_[5684]_ ,
    \new_[5685]_ , \new_[5686]_ , \new_[5687]_ , \new_[5688]_ ,
    \new_[5689]_ , \new_[5690]_ , \new_[5691]_ , \new_[5692]_ ,
    \new_[5693]_ , \new_[5694]_ , \new_[5695]_ , \new_[5696]_ ,
    \new_[5697]_ , \new_[5698]_ , \new_[5699]_ , \new_[5700]_ ,
    \new_[5701]_ , \new_[5702]_ , \new_[5703]_ , \new_[5704]_ ,
    \new_[5705]_ , \new_[5706]_ , \new_[5707]_ , \new_[5708]_ ,
    \new_[5709]_ , \new_[5710]_ , \new_[5711]_ , \new_[5712]_ ,
    \new_[5713]_ , \new_[5714]_ , \new_[5715]_ , \new_[5716]_ ,
    \new_[5717]_ , \new_[5718]_ , \new_[5719]_ , \new_[5720]_ ,
    \new_[5721]_ , \new_[5722]_ , \new_[5723]_ , \new_[5724]_ ,
    \new_[5725]_ , \new_[5726]_ , \new_[5727]_ , \new_[5728]_ ,
    \new_[5729]_ , \new_[5730]_ , \new_[5731]_ , \new_[5732]_ ,
    \new_[5733]_ , \new_[5734]_ , \new_[5735]_ , \new_[5736]_ ,
    \new_[5737]_ , \new_[5738]_ , \new_[5739]_ , \new_[5740]_ ,
    \new_[5741]_ , \new_[5742]_ , \new_[5743]_ , \new_[5744]_ ,
    \new_[5745]_ , \new_[5746]_ , \new_[5747]_ , \new_[5748]_ ,
    \new_[5749]_ , \new_[5750]_ , \new_[5751]_ , \new_[5752]_ ,
    \new_[5753]_ , \new_[5754]_ , \new_[5755]_ , \new_[5756]_ ,
    \new_[5757]_ , \new_[5758]_ , \new_[5759]_ , \new_[5760]_ ,
    \new_[5761]_ , \new_[5762]_ , \new_[5763]_ , \new_[5764]_ ,
    \new_[5765]_ , \new_[5766]_ , \new_[5767]_ , \new_[5768]_ ,
    \new_[5769]_ , \new_[5770]_ , \new_[5771]_ , \new_[5772]_ ,
    \new_[5773]_ , \new_[5774]_ , \new_[5775]_ , \new_[5776]_ ,
    \new_[5777]_ , \new_[5778]_ , \new_[5779]_ , \new_[5780]_ ,
    \new_[5781]_ , \new_[5782]_ , \new_[5783]_ , \new_[5784]_ ,
    \new_[5785]_ , \new_[5786]_ , \new_[5787]_ , \new_[5788]_ ,
    \new_[5789]_ , \new_[5790]_ , \new_[5791]_ , \new_[5792]_ ,
    \new_[5793]_ , \new_[5794]_ , \new_[5795]_ , \new_[5796]_ ,
    \new_[5797]_ , \new_[5798]_ , \new_[5799]_ , \new_[5800]_ ,
    \new_[5801]_ , \new_[5802]_ , \new_[5803]_ , \new_[5804]_ ,
    \new_[5805]_ , \new_[5806]_ , \new_[5807]_ , \new_[5808]_ ,
    \new_[5809]_ , \new_[5810]_ , \new_[5811]_ , \new_[5812]_ ,
    \new_[5813]_ , \new_[5814]_ , \new_[5815]_ , \new_[5816]_ ,
    \new_[5817]_ , \new_[5818]_ , \new_[5819]_ , \new_[5820]_ ,
    \new_[5821]_ , \new_[5822]_ , \new_[5823]_ , \new_[5824]_ ,
    \new_[5825]_ , \new_[5826]_ , \new_[5827]_ , \new_[5828]_ ,
    \new_[5829]_ , \new_[5830]_ , \new_[5831]_ , \new_[5832]_ ,
    \new_[5833]_ , \new_[5834]_ , \new_[5835]_ , \new_[5836]_ ,
    \new_[5837]_ , \new_[5838]_ , \new_[5839]_ , \new_[5840]_ ,
    \new_[5841]_ , \new_[5842]_ , \new_[5843]_ , \new_[5844]_ ,
    \new_[5845]_ , \new_[5846]_ , \new_[5847]_ , \new_[5848]_ ,
    \new_[5849]_ , \new_[5850]_ , \new_[5851]_ , \new_[5852]_ ,
    \new_[5853]_ , \new_[5854]_ , \new_[5855]_ , \new_[5856]_ ,
    \new_[5857]_ , \new_[5858]_ , \new_[5859]_ , \new_[5860]_ ,
    \new_[5861]_ , \new_[5862]_ , \new_[5863]_ , \new_[5864]_ ,
    \new_[5865]_ , \new_[5866]_ , \new_[5867]_ , \new_[5868]_ ,
    \new_[5869]_ , \new_[5870]_ , \new_[5871]_ , \new_[5872]_ ,
    \new_[5873]_ , \new_[5874]_ , \new_[5875]_ , \new_[5876]_ ,
    \new_[5877]_ , \new_[5878]_ , \new_[5879]_ , \new_[5880]_ ,
    \new_[5881]_ , \new_[5882]_ , \new_[5883]_ , \new_[5884]_ ,
    \new_[5885]_ , \new_[5886]_ , \new_[5887]_ , \new_[5888]_ ,
    \new_[5889]_ , \new_[5890]_ , \new_[5891]_ , \new_[5892]_ ,
    \new_[5893]_ , \new_[5894]_ , \new_[5895]_ , \new_[5896]_ ,
    \new_[5897]_ , \new_[5898]_ , \new_[5899]_ , \new_[5900]_ ,
    \new_[5901]_ , \new_[5902]_ , \new_[5903]_ , \new_[5904]_ ,
    \new_[5905]_ , \new_[5906]_ , \new_[5907]_ , \new_[5908]_ ,
    \new_[5909]_ , \new_[5910]_ , \new_[5911]_ , \new_[5912]_ ,
    \new_[5913]_ , \new_[5914]_ , \new_[5915]_ , \new_[5916]_ ,
    \new_[5917]_ , \new_[5918]_ , \new_[5919]_ , \new_[5920]_ ,
    \new_[5921]_ , \new_[5922]_ , \new_[5923]_ , \new_[5924]_ ,
    \new_[5925]_ , \new_[5926]_ , \new_[5927]_ , \new_[5928]_ ,
    \new_[5929]_ , \new_[5930]_ , \new_[5931]_ , \new_[5932]_ ,
    \new_[5933]_ , \new_[5934]_ , \new_[5935]_ , \new_[5936]_ ,
    \new_[5937]_ , \new_[5938]_ , \new_[5939]_ , \new_[5940]_ ,
    \new_[5941]_ , \new_[5942]_ , \new_[5943]_ , \new_[5944]_ ,
    \new_[5945]_ , \new_[5946]_ , \new_[5947]_ , \new_[5948]_ ,
    \new_[5949]_ , \new_[5950]_ , \new_[5951]_ , \new_[5952]_ ,
    \new_[5953]_ , \new_[5954]_ , \new_[5955]_ , \new_[5956]_ ,
    \new_[5957]_ , \new_[5958]_ , \new_[5959]_ , \new_[5960]_ ,
    \new_[5961]_ , \new_[5962]_ , \new_[5963]_ , \new_[5964]_ ,
    \new_[5965]_ , \new_[5966]_ , \new_[5967]_ , \new_[5968]_ ,
    \new_[5969]_ , \new_[5970]_ , \new_[5971]_ , \new_[5972]_ ,
    \new_[5973]_ , \new_[5974]_ , \new_[5975]_ , \new_[5976]_ ,
    \new_[5977]_ , \new_[5978]_ , \new_[5979]_ , \new_[5980]_ ,
    \new_[5981]_ , \new_[5982]_ , \new_[5983]_ , \new_[5984]_ ,
    \new_[5985]_ , \new_[5986]_ , \new_[5987]_ , \new_[5988]_ ,
    \new_[5989]_ , \new_[5990]_ , \new_[5991]_ , \new_[5992]_ ,
    \new_[5993]_ , \new_[5994]_ , \new_[5995]_ , \new_[5996]_ ,
    \new_[5997]_ , \new_[5998]_ , \new_[5999]_ , \new_[6000]_ ,
    \new_[6001]_ , \new_[6002]_ , \new_[6003]_ , \new_[6004]_ ,
    \new_[6005]_ , \new_[6006]_ , \new_[6007]_ , \new_[6008]_ ,
    \new_[6009]_ , \new_[6010]_ , \new_[6011]_ , \new_[6012]_ ,
    \new_[6013]_ , \new_[6014]_ , \new_[6015]_ , \new_[6016]_ ,
    \new_[6017]_ , \new_[6018]_ , \new_[6019]_ , \new_[6020]_ ,
    \new_[6021]_ , \new_[6022]_ , \new_[6023]_ , \new_[6024]_ ,
    \new_[6025]_ , \new_[6026]_ , \new_[6027]_ , \new_[6028]_ ,
    \new_[6029]_ , \new_[6030]_ , \new_[6031]_ , \new_[6032]_ ,
    \new_[6033]_ , \new_[6034]_ , \new_[6035]_ , \new_[6036]_ ,
    \new_[6037]_ , \new_[6038]_ , \new_[6039]_ , \new_[6040]_ ,
    \new_[6041]_ , \new_[6042]_ , \new_[6043]_ , \new_[6044]_ ,
    \new_[6045]_ , \new_[6046]_ , \new_[6047]_ , \new_[6048]_ ,
    \new_[6049]_ , \new_[6050]_ , \new_[6051]_ , \new_[6052]_ ,
    \new_[6053]_ , \new_[6054]_ , \new_[6055]_ , \new_[6056]_ ,
    \new_[6057]_ , \new_[6058]_ , \new_[6059]_ , \new_[6060]_ ,
    \new_[6061]_ , \new_[6062]_ , \new_[6063]_ , \new_[6064]_ ,
    \new_[6065]_ , \new_[6066]_ , \new_[6067]_ , \new_[6068]_ ,
    \new_[6069]_ , \new_[6070]_ , \new_[6071]_ , \new_[6072]_ ,
    \new_[6073]_ , \new_[6074]_ , \new_[6075]_ , \new_[6076]_ ,
    \new_[6077]_ , \new_[6078]_ , \new_[6079]_ , \new_[6080]_ ,
    \new_[6081]_ , \new_[6082]_ , \new_[6083]_ , \new_[6084]_ ,
    \new_[6085]_ , \new_[6086]_ , \new_[6087]_ , \new_[6088]_ ,
    \new_[6089]_ , \new_[6090]_ , \new_[6091]_ , \new_[6092]_ ,
    \new_[6093]_ , \new_[6094]_ , \new_[6095]_ , \new_[6096]_ ,
    \new_[6097]_ , \new_[6098]_ , \new_[6099]_ , \new_[6100]_ ,
    \new_[6101]_ , \new_[6102]_ , \new_[6103]_ , \new_[6104]_ ,
    \new_[6105]_ , \new_[6106]_ , \new_[6107]_ , \new_[6108]_ ,
    \new_[6109]_ , \new_[6110]_ , \new_[6111]_ , \new_[6112]_ ,
    \new_[6113]_ , \new_[6114]_ , \new_[6115]_ , \new_[6116]_ ,
    \new_[6117]_ , \new_[6118]_ , \new_[6119]_ , \new_[6120]_ ,
    \new_[6121]_ , \new_[6122]_ , \new_[6123]_ , \new_[6124]_ ,
    \new_[6125]_ , \new_[6126]_ , \new_[6127]_ , \new_[6128]_ ,
    \new_[6129]_ , \new_[6130]_ , \new_[6131]_ , \new_[6132]_ ,
    \new_[6133]_ , \new_[6134]_ , \new_[6135]_ , \new_[6136]_ ,
    \new_[6137]_ , \new_[6138]_ , \new_[6139]_ , \new_[6140]_ ,
    \new_[6141]_ , \new_[6142]_ , \new_[6143]_ , \new_[6144]_ ,
    \new_[6145]_ , \new_[6146]_ , \new_[6147]_ , \new_[6148]_ ,
    \new_[6149]_ , \new_[6150]_ , \new_[6151]_ , \new_[6152]_ ,
    \new_[6153]_ , \new_[6154]_ , \new_[6155]_ , \new_[6156]_ ,
    \new_[6157]_ , \new_[6158]_ , \new_[6159]_ , \new_[6160]_ ,
    \new_[6161]_ , \new_[6162]_ , \new_[6163]_ , \new_[6164]_ ,
    \new_[6165]_ , \new_[6166]_ , \new_[6167]_ , \new_[6168]_ ,
    \new_[6169]_ , \new_[6170]_ , \new_[6171]_ , \new_[6172]_ ,
    \new_[6173]_ , \new_[6174]_ , \new_[6175]_ , \new_[6176]_ ,
    \new_[6177]_ , \new_[6178]_ , \new_[6179]_ , \new_[6180]_ ,
    \new_[6181]_ , \new_[6182]_ , \new_[6183]_ , \new_[6184]_ ,
    \new_[6185]_ , \new_[6186]_ , \new_[6187]_ , \new_[6188]_ ,
    \new_[6189]_ , \new_[6190]_ , \new_[6191]_ , \new_[6192]_ ,
    \new_[6193]_ , \new_[6194]_ , \new_[6195]_ , \new_[6196]_ ,
    \new_[6197]_ , \new_[6198]_ , \new_[6199]_ , \new_[6200]_ ,
    \new_[6201]_ , \new_[6202]_ , \new_[6203]_ , \new_[6204]_ ,
    \new_[6205]_ , \new_[6206]_ , \new_[6207]_ , \new_[6208]_ ,
    \new_[6209]_ , \new_[6210]_ , \new_[6211]_ , \new_[6212]_ ,
    \new_[6213]_ , \new_[6214]_ , \new_[6215]_ , \new_[6216]_ ,
    \new_[6217]_ , \new_[6218]_ , \new_[6219]_ , \new_[6220]_ ,
    \new_[6221]_ , \new_[6222]_ , \new_[6223]_ , \new_[6224]_ ,
    \new_[6225]_ , \new_[6226]_ , \new_[6227]_ , \new_[6228]_ ,
    \new_[6229]_ , \new_[6230]_ , \new_[6231]_ , \new_[6232]_ ,
    \new_[6233]_ , \new_[6234]_ , \new_[6235]_ , \new_[6236]_ ,
    \new_[6237]_ , \new_[6238]_ , \new_[6239]_ , \new_[6240]_ ,
    \new_[6241]_ , \new_[6242]_ , \new_[6243]_ , \new_[6244]_ ,
    \new_[6245]_ , \new_[6246]_ , \new_[6247]_ , \new_[6248]_ ,
    \new_[6249]_ , \new_[6250]_ , \new_[6251]_ , \new_[6252]_ ,
    \new_[6253]_ , \new_[6254]_ , \new_[6255]_ , \new_[6256]_ ,
    \new_[6257]_ , \new_[6258]_ , \new_[6259]_ , \new_[6260]_ ,
    \new_[6261]_ , \new_[6262]_ , \new_[6263]_ , \new_[6264]_ ,
    \new_[6265]_ , \new_[6266]_ , \new_[6267]_ , \new_[6268]_ ,
    \new_[6269]_ , \new_[6270]_ , \new_[6271]_ , \new_[6272]_ ,
    \new_[6273]_ , \new_[6274]_ , \new_[6275]_ , \new_[6276]_ ,
    \new_[6277]_ , \new_[6278]_ , \new_[6279]_ , \new_[6280]_ ,
    \new_[6281]_ , \new_[6282]_ , \new_[6283]_ , \new_[6284]_ ,
    \new_[6285]_ , \new_[6286]_ , \new_[6287]_ , \new_[6288]_ ,
    \new_[6289]_ , \new_[6290]_ , \new_[6291]_ , \new_[6292]_ ,
    \new_[6293]_ , \new_[6294]_ , \new_[6295]_ , \new_[6296]_ ,
    \new_[6297]_ , \new_[6298]_ , \new_[6299]_ , \new_[6300]_ ,
    \new_[6301]_ , \new_[6302]_ , \new_[6303]_ , \new_[6304]_ ,
    \new_[6305]_ , \new_[6306]_ , \new_[6307]_ , \new_[6308]_ ,
    \new_[6309]_ , \new_[6310]_ , \new_[6311]_ , \new_[6312]_ ,
    \new_[6313]_ , \new_[6314]_ , \new_[6315]_ , \new_[6316]_ ,
    \new_[6317]_ , \new_[6318]_ , \new_[6319]_ , \new_[6320]_ ,
    \new_[6321]_ , \new_[6322]_ , \new_[6323]_ , \new_[6324]_ ,
    \new_[6325]_ , \new_[6326]_ , \new_[6327]_ , \new_[6328]_ ,
    \new_[6329]_ , \new_[6330]_ , \new_[6331]_ , \new_[6332]_ ,
    \new_[6333]_ , \new_[6334]_ , \new_[6335]_ , \new_[6336]_ ,
    \new_[6337]_ , \new_[6338]_ , \new_[6339]_ , \new_[6340]_ ,
    \new_[6341]_ , \new_[6342]_ , \new_[6343]_ , \new_[6344]_ ,
    \new_[6345]_ , \new_[6346]_ , \new_[6347]_ , \new_[6348]_ ,
    \new_[6349]_ , \new_[6350]_ , \new_[6351]_ , \new_[6352]_ ,
    \new_[6353]_ , \new_[6354]_ , \new_[6355]_ , \new_[6356]_ ,
    \new_[6357]_ , \new_[6358]_ , \new_[6359]_ , \new_[6360]_ ,
    \new_[6361]_ , \new_[6362]_ , \new_[6363]_ , \new_[6364]_ ,
    \new_[6365]_ , \new_[6366]_ , \new_[6367]_ , \new_[6368]_ ,
    \new_[6369]_ , \new_[6370]_ , \new_[6371]_ , \new_[6372]_ ,
    \new_[6373]_ , \new_[6374]_ , \new_[6375]_ , \new_[6376]_ ,
    \new_[6377]_ , \new_[6378]_ , \new_[6379]_ , \new_[6380]_ ,
    \new_[6381]_ , \new_[6382]_ , \new_[6383]_ , \new_[6384]_ ,
    \new_[6385]_ , \new_[6386]_ , \new_[6387]_ , \new_[6388]_ ,
    \new_[6389]_ , \new_[6390]_ , \new_[6391]_ , \new_[6392]_ ,
    \new_[6393]_ , \new_[6394]_ , \new_[6395]_ , \new_[6396]_ ,
    \new_[6397]_ , \new_[6398]_ , \new_[6399]_ , \new_[6400]_ ,
    \new_[6401]_ , \new_[6402]_ , \new_[6403]_ , \new_[6404]_ ,
    \new_[6405]_ , \new_[6406]_ , \new_[6407]_ , \new_[6408]_ ,
    \new_[6409]_ , \new_[6410]_ , \new_[6411]_ , \new_[6412]_ ,
    \new_[6413]_ , \new_[6414]_ , \new_[6415]_ , \new_[6416]_ ,
    \new_[6417]_ , \new_[6418]_ , \new_[6419]_ , \new_[6420]_ ,
    \new_[6421]_ , \new_[6422]_ , \new_[6423]_ , \new_[6424]_ ,
    \new_[6425]_ , \new_[6426]_ , \new_[6427]_ , \new_[6428]_ ,
    \new_[6429]_ , \new_[6430]_ , \new_[6431]_ , \new_[6432]_ ,
    \new_[6433]_ , \new_[6434]_ , \new_[6435]_ , \new_[6436]_ ,
    \new_[6437]_ , \new_[6438]_ , \new_[6439]_ , \new_[6440]_ ,
    \new_[6441]_ , \new_[6442]_ , \new_[6443]_ , \new_[6444]_ ,
    \new_[6445]_ , \new_[6446]_ , \new_[6447]_ , \new_[6448]_ ,
    \new_[6449]_ , \new_[6450]_ , \new_[6451]_ , \new_[6452]_ ,
    \new_[6453]_ , \new_[6454]_ , \new_[6455]_ , \new_[6456]_ ,
    \new_[6457]_ , \new_[6458]_ , \new_[6459]_ , \new_[6460]_ ,
    \new_[6461]_ , \new_[6462]_ , \new_[6463]_ , \new_[6464]_ ,
    \new_[6465]_ , \new_[6466]_ , \new_[6467]_ , \new_[6468]_ ,
    \new_[6469]_ , \new_[6470]_ , \new_[6471]_ , \new_[6472]_ ,
    \new_[6473]_ , \new_[6474]_ , \new_[6475]_ , \new_[6476]_ ,
    \new_[6477]_ , \new_[6478]_ , \new_[6479]_ , \new_[6480]_ ,
    \new_[6481]_ , \new_[6482]_ , \new_[6483]_ , \new_[6484]_ ,
    \new_[6485]_ , \new_[6486]_ , \new_[6487]_ , \new_[6488]_ ,
    \new_[6489]_ , \new_[6490]_ , \new_[6491]_ , \new_[6492]_ ,
    \new_[6493]_ , \new_[6494]_ , \new_[6495]_ , \new_[6496]_ ,
    \new_[6497]_ , \new_[6498]_ , \new_[6499]_ , \new_[6500]_ ,
    \new_[6501]_ , \new_[6502]_ , \new_[6503]_ , \new_[6504]_ ,
    \new_[6505]_ , \new_[6506]_ , \new_[6507]_ , \new_[6508]_ ,
    \new_[6509]_ , \new_[6510]_ , \new_[6511]_ , \new_[6512]_ ,
    \new_[6513]_ , \new_[6514]_ , \new_[6515]_ , \new_[6516]_ ,
    \new_[6517]_ , \new_[6518]_ , \new_[6519]_ , \new_[6520]_ ,
    \new_[6521]_ , \new_[6522]_ , \new_[6523]_ , \new_[6524]_ ,
    \new_[6525]_ , \new_[6526]_ , \new_[6527]_ , \new_[6528]_ ,
    \new_[6529]_ , \new_[6530]_ , \new_[6531]_ , \new_[6532]_ ,
    \new_[6533]_ , \new_[6534]_ , \new_[6535]_ , \new_[6536]_ ,
    \new_[6537]_ , \new_[6538]_ , \new_[6539]_ , \new_[6540]_ ,
    \new_[6541]_ , \new_[6542]_ , \new_[6543]_ , \new_[6544]_ ,
    \new_[6545]_ , \new_[6546]_ , \new_[6547]_ , \new_[6548]_ ,
    \new_[6549]_ , \new_[6550]_ , \new_[6551]_ , \new_[6552]_ ,
    \new_[6553]_ , \new_[6554]_ , \new_[6555]_ , \new_[6556]_ ,
    \new_[6557]_ , \new_[6558]_ , \new_[6559]_ , \new_[6560]_ ,
    \new_[6561]_ , \new_[6562]_ , \new_[6563]_ , \new_[6564]_ ,
    \new_[6565]_ , \new_[6566]_ , \new_[6567]_ , \new_[6568]_ ,
    \new_[6569]_ , \new_[6570]_ , \new_[6571]_ , \new_[6572]_ ,
    \new_[6573]_ , \new_[6574]_ , \new_[6575]_ , \new_[6576]_ ,
    \new_[6577]_ , \new_[6578]_ , \new_[6579]_ , \new_[6580]_ ,
    \new_[6581]_ , \new_[6582]_ , \new_[6583]_ , \new_[6584]_ ,
    \new_[6585]_ , \new_[6586]_ , \new_[6587]_ , \new_[6588]_ ,
    \new_[6589]_ , \new_[6590]_ , \new_[6591]_ , \new_[6592]_ ,
    \new_[6593]_ , \new_[6594]_ , \new_[6595]_ , \new_[6596]_ ,
    \new_[6597]_ , \new_[6598]_ , \new_[6599]_ , \new_[6600]_ ,
    \new_[6601]_ , \new_[6602]_ , \new_[6603]_ , \new_[6604]_ ,
    \new_[6605]_ , \new_[6606]_ , \new_[6607]_ , \new_[6608]_ ,
    \new_[6609]_ , \new_[6610]_ , \new_[6611]_ , \new_[6612]_ ,
    \new_[6613]_ , \new_[6614]_ , \new_[6615]_ , \new_[6616]_ ,
    \new_[6617]_ , \new_[6618]_ , \new_[6619]_ , \new_[6620]_ ,
    \new_[6621]_ , \new_[6622]_ , \new_[6623]_ , \new_[6624]_ ,
    \new_[6625]_ , \new_[6626]_ , \new_[6627]_ , \new_[6628]_ ,
    \new_[6629]_ , \new_[6630]_ , \new_[6631]_ , \new_[6632]_ ,
    \new_[6633]_ , \new_[6634]_ , \new_[6635]_ , \new_[6636]_ ,
    \new_[6637]_ , \new_[6638]_ , \new_[6639]_ , \new_[6640]_ ,
    \new_[6641]_ , \new_[6642]_ , \new_[6643]_ , \new_[6644]_ ,
    \new_[6645]_ , \new_[6646]_ , \new_[6647]_ , \new_[6648]_ ,
    \new_[6649]_ , \new_[6650]_ , \new_[6651]_ , \new_[6652]_ ,
    \new_[6653]_ , \new_[6654]_ , \new_[6655]_ , \new_[6656]_ ,
    \new_[6657]_ , \new_[6658]_ , \new_[6659]_ , \new_[6660]_ ,
    \new_[6661]_ , \new_[6662]_ , \new_[6663]_ , \new_[6664]_ ,
    \new_[6665]_ , \new_[6666]_ , \new_[6667]_ , \new_[6668]_ ,
    \new_[6669]_ , \new_[6670]_ , \new_[6671]_ , \new_[6672]_ ,
    \new_[6673]_ , \new_[6674]_ , \new_[6675]_ , \new_[6676]_ ,
    \new_[6677]_ , \new_[6678]_ , \new_[6679]_ , \new_[6680]_ ,
    \new_[6681]_ , \new_[6682]_ , \new_[6683]_ , \new_[6684]_ ,
    \new_[6685]_ , \new_[6686]_ , \new_[6687]_ , \new_[6688]_ ,
    \new_[6689]_ , \new_[6690]_ , \new_[6691]_ , \new_[6692]_ ,
    \new_[6693]_ , \new_[6694]_ , \new_[6695]_ , \new_[6696]_ ,
    \new_[6697]_ , \new_[6698]_ , \new_[6699]_ , \new_[6700]_ ,
    \new_[6701]_ , \new_[6702]_ , \new_[6703]_ , \new_[6704]_ ,
    \new_[6705]_ , \new_[6706]_ , \new_[6707]_ , \new_[6708]_ ,
    \new_[6709]_ , \new_[6710]_ , \new_[6711]_ , \new_[6712]_ ,
    \new_[6713]_ , \new_[6714]_ , \new_[6715]_ , \new_[6716]_ ,
    \new_[6717]_ , \new_[6718]_ , \new_[6719]_ , \new_[6720]_ ,
    \new_[6721]_ , \new_[6722]_ , \new_[6723]_ , \new_[6724]_ ,
    \new_[6725]_ , \new_[6726]_ , \new_[6727]_ , \new_[6728]_ ,
    \new_[6729]_ , \new_[6730]_ , \new_[6731]_ , \new_[6732]_ ,
    \new_[6733]_ , \new_[6734]_ , \new_[6735]_ , \new_[6736]_ ,
    \new_[6737]_ , \new_[6738]_ , \new_[6739]_ , \new_[6740]_ ,
    \new_[6741]_ , \new_[6742]_ , \new_[6743]_ , \new_[6744]_ ,
    \new_[6745]_ , \new_[6746]_ , \new_[6747]_ , \new_[6748]_ ,
    \new_[6749]_ , \new_[6750]_ , \new_[6751]_ , \new_[6752]_ ,
    \new_[6753]_ , \new_[6754]_ , \new_[6755]_ , \new_[6756]_ ,
    \new_[6757]_ , \new_[6758]_ , \new_[6759]_ , \new_[6760]_ ,
    \new_[6761]_ , \new_[6762]_ , \new_[6763]_ , \new_[6764]_ ,
    \new_[6765]_ , \new_[6766]_ , \new_[6767]_ , \new_[6768]_ ,
    \new_[6769]_ , \new_[6770]_ , \new_[6771]_ , \new_[6772]_ ,
    \new_[6773]_ , \new_[6774]_ , \new_[6775]_ , \new_[6776]_ ,
    \new_[6777]_ , \new_[6778]_ , \new_[6779]_ , \new_[6780]_ ,
    \new_[6781]_ , \new_[6782]_ , \new_[6783]_ , \new_[6784]_ ,
    \new_[6785]_ , \new_[6786]_ , \new_[6787]_ , \new_[6788]_ ,
    \new_[6789]_ , \new_[6790]_ , \new_[6791]_ , \new_[6792]_ ,
    \new_[6793]_ , \new_[6794]_ , \new_[6795]_ , \new_[6796]_ ,
    \new_[6797]_ , \new_[6798]_ , \new_[6799]_ , \new_[6800]_ ,
    \new_[6801]_ , \new_[6802]_ , \new_[6803]_ , \new_[6804]_ ,
    \new_[6805]_ , \new_[6806]_ , \new_[6807]_ , \new_[6808]_ ,
    \new_[6809]_ , \new_[6810]_ , \new_[6811]_ , \new_[6812]_ ,
    \new_[6813]_ , \new_[6814]_ , \new_[6815]_ , \new_[6816]_ ,
    \new_[6817]_ , \new_[6818]_ , \new_[6819]_ , \new_[6820]_ ,
    \new_[6821]_ , \new_[6822]_ , \new_[6823]_ , \new_[6824]_ ,
    \new_[6825]_ , \new_[6826]_ , \new_[6827]_ , \new_[6828]_ ,
    \new_[6829]_ , \new_[6830]_ , \new_[6831]_ , \new_[6832]_ ,
    \new_[6833]_ , \new_[6834]_ , \new_[6835]_ , \new_[6836]_ ,
    \new_[6837]_ , \new_[6838]_ , \new_[6839]_ , \new_[6840]_ ,
    \new_[6841]_ , \new_[6842]_ , \new_[6843]_ , \new_[6844]_ ,
    \new_[6845]_ , \new_[6846]_ , \new_[6847]_ , \new_[6848]_ ,
    \new_[6849]_ , \new_[6850]_ , \new_[6851]_ , \new_[6852]_ ,
    \new_[6853]_ , \new_[6854]_ , \new_[6855]_ , \new_[6856]_ ,
    \new_[6857]_ , \new_[6858]_ , \new_[6859]_ , \new_[6860]_ ,
    \new_[6861]_ , \new_[6862]_ , \new_[6863]_ , \new_[6864]_ ,
    \new_[6865]_ , \new_[6866]_ , \new_[6867]_ , \new_[6868]_ ,
    \new_[6869]_ , \new_[6870]_ , \new_[6871]_ , \new_[6872]_ ,
    \new_[6873]_ , \new_[6874]_ , \new_[6875]_ , \new_[6876]_ ,
    \new_[6877]_ , \new_[6878]_ , \new_[6879]_ , \new_[6880]_ ,
    \new_[6881]_ , \new_[6882]_ , \new_[6883]_ , \new_[6884]_ ,
    \new_[6885]_ , \new_[6886]_ , \new_[6887]_ , \new_[6888]_ ,
    \new_[6889]_ , \new_[6890]_ , \new_[6891]_ , \new_[6892]_ ,
    \new_[6893]_ , \new_[6894]_ , \new_[6895]_ , \new_[6896]_ ,
    \new_[6897]_ , \new_[6898]_ , \new_[6899]_ , \new_[6900]_ ,
    \new_[6901]_ , \new_[6902]_ , \new_[6903]_ , \new_[6904]_ ,
    \new_[6905]_ , \new_[6906]_ , \new_[6907]_ , \new_[6908]_ ,
    \new_[6909]_ , \new_[6910]_ , \new_[6911]_ , \new_[6912]_ ,
    \new_[6913]_ , \new_[6914]_ , \new_[6915]_ , \new_[6916]_ ,
    \new_[6917]_ , \new_[6918]_ , \new_[6919]_ , \new_[6920]_ ,
    \new_[6921]_ , \new_[6922]_ , \new_[6923]_ , \new_[6924]_ ,
    \new_[6925]_ , \new_[6926]_ , \new_[6927]_ , \new_[6928]_ ,
    \new_[6929]_ , \new_[6930]_ , \new_[6931]_ , \new_[6932]_ ,
    \new_[6933]_ , \new_[6934]_ , \new_[6935]_ , \new_[6936]_ ,
    \new_[6937]_ , \new_[6938]_ , \new_[6939]_ , \new_[6940]_ ,
    \new_[6941]_ , \new_[6942]_ , \new_[6943]_ , \new_[6944]_ ,
    \new_[6945]_ , \new_[6946]_ , \new_[6947]_ , \new_[6948]_ ,
    \new_[6949]_ , \new_[6950]_ , \new_[6951]_ , \new_[6952]_ ,
    \new_[6953]_ , \new_[6954]_ , \new_[6955]_ , \new_[6956]_ ,
    \new_[6957]_ , \new_[6958]_ , \new_[6959]_ , \new_[6960]_ ,
    \new_[6961]_ , \new_[6962]_ , \new_[6963]_ , \new_[6964]_ ,
    \new_[6965]_ , \new_[6966]_ , \new_[6967]_ , \new_[6968]_ ,
    \new_[6969]_ , \new_[6970]_ , \new_[6971]_ , \new_[6972]_ ,
    \new_[6973]_ , \new_[6974]_ , \new_[6975]_ , \new_[6976]_ ,
    \new_[6977]_ , \new_[6978]_ , \new_[6979]_ , \new_[6980]_ ,
    \new_[6981]_ , \new_[6982]_ , \new_[6983]_ , \new_[6984]_ ,
    \new_[6985]_ , \new_[6986]_ , \new_[6987]_ , \new_[6988]_ ,
    \new_[6989]_ , \new_[6990]_ , \new_[6991]_ , \new_[6992]_ ,
    \new_[6993]_ , \new_[6994]_ , \new_[6995]_ , \new_[6996]_ ,
    \new_[6997]_ , \new_[6998]_ , \new_[6999]_ , \new_[7000]_ ,
    \new_[7001]_ , \new_[7002]_ , \new_[7003]_ , \new_[7004]_ ,
    \new_[7005]_ , \new_[7006]_ , \new_[7007]_ , \new_[7008]_ ,
    \new_[7009]_ , \new_[7010]_ , \new_[7011]_ , \new_[7012]_ ,
    \new_[7013]_ , \new_[7014]_ , \new_[7015]_ , \new_[7016]_ ,
    \new_[7017]_ , \new_[7018]_ , \new_[7019]_ , \new_[7020]_ ,
    \new_[7021]_ , \new_[7022]_ , \new_[7023]_ , \new_[7024]_ ,
    \new_[7025]_ , \new_[7026]_ , \new_[7027]_ , \new_[7028]_ ,
    \new_[7029]_ , \new_[7030]_ , \new_[7031]_ , \new_[7032]_ ,
    \new_[7033]_ , \new_[7034]_ , \new_[7035]_ , \new_[7036]_ ,
    \new_[7037]_ , \new_[7038]_ , \new_[7039]_ , \new_[7040]_ ,
    \new_[7041]_ , \new_[7042]_ , \new_[7043]_ , \new_[7044]_ ,
    \new_[7045]_ , \new_[7046]_ , \new_[7047]_ , \new_[7048]_ ,
    \new_[7049]_ , \new_[7050]_ , \new_[7051]_ , \new_[7052]_ ,
    \new_[7053]_ , \new_[7054]_ , \new_[7055]_ , \new_[7056]_ ,
    \new_[7057]_ , \new_[7058]_ , \new_[7059]_ , \new_[7060]_ ,
    \new_[7061]_ , \new_[7062]_ , \new_[7063]_ , \new_[7064]_ ,
    \new_[7065]_ , \new_[7066]_ , \new_[7067]_ , \new_[7068]_ ,
    \new_[7069]_ , \new_[7070]_ , \new_[7071]_ , \new_[7072]_ ,
    \new_[7073]_ , \new_[7074]_ , \new_[7075]_ , \new_[7076]_ ,
    \new_[7077]_ , \new_[7078]_ , \new_[7079]_ , \new_[7080]_ ,
    \new_[7081]_ , \new_[7082]_ , \new_[7083]_ , \new_[7084]_ ,
    \new_[7085]_ , \new_[7086]_ , \new_[7087]_ , \new_[7088]_ ,
    \new_[7089]_ , \new_[7090]_ , \new_[7091]_ , \new_[7092]_ ,
    \new_[7093]_ , \new_[7094]_ , \new_[7095]_ , \new_[7096]_ ,
    \new_[7097]_ , \new_[7098]_ , \new_[7099]_ , \new_[7100]_ ,
    \new_[7101]_ , \new_[7102]_ , \new_[7103]_ , \new_[7104]_ ,
    \new_[7105]_ , \new_[7106]_ , \new_[7107]_ , \new_[7108]_ ,
    \new_[7109]_ , \new_[7110]_ , \new_[7111]_ , \new_[7112]_ ,
    \new_[7113]_ , \new_[7114]_ , \new_[7115]_ , \new_[7116]_ ,
    \new_[7117]_ , \new_[7118]_ , \new_[7119]_ , \new_[7120]_ ,
    \new_[7121]_ , \new_[7122]_ , \new_[7123]_ , \new_[7124]_ ,
    \new_[7125]_ , \new_[7126]_ , \new_[7127]_ , \new_[7128]_ ,
    \new_[7129]_ , \new_[7130]_ , \new_[7131]_ , \new_[7132]_ ,
    \new_[7133]_ , \new_[7134]_ , \new_[7135]_ , \new_[7136]_ ,
    \new_[7137]_ , \new_[7138]_ , \new_[7139]_ , \new_[7140]_ ,
    \new_[7141]_ , \new_[7142]_ , \new_[7143]_ , \new_[7144]_ ,
    \new_[7145]_ , \new_[7146]_ , \new_[7147]_ , \new_[7148]_ ,
    \new_[7149]_ , \new_[7150]_ , \new_[7151]_ , \new_[7152]_ ,
    \new_[7153]_ , \new_[7154]_ , \new_[7155]_ , \new_[7156]_ ,
    \new_[7157]_ , \new_[7158]_ , \new_[7159]_ , \new_[7160]_ ,
    \new_[7161]_ , \new_[7162]_ , \new_[7163]_ , \new_[7164]_ ,
    \new_[7165]_ , \new_[7166]_ , \new_[7167]_ , \new_[7168]_ ,
    \new_[7169]_ , \new_[7170]_ , \new_[7171]_ , \new_[7172]_ ,
    \new_[7173]_ , \new_[7174]_ , \new_[7175]_ , \new_[7176]_ ,
    \new_[7177]_ , \new_[7178]_ , \new_[7179]_ , \new_[7180]_ ,
    \new_[7181]_ , \new_[7182]_ , \new_[7183]_ , \new_[7184]_ ,
    \new_[7185]_ , \new_[7186]_ , \new_[7187]_ , \new_[7188]_ ,
    \new_[7189]_ , \new_[7190]_ , \new_[7191]_ , \new_[7192]_ ,
    \new_[7193]_ , \new_[7194]_ , \new_[7195]_ , \new_[7196]_ ,
    \new_[7197]_ , \new_[7198]_ , \new_[7199]_ , \new_[7200]_ ,
    \new_[7201]_ , \new_[7202]_ , \new_[7203]_ , \new_[7204]_ ,
    \new_[7205]_ , \new_[7206]_ , \new_[7207]_ , \new_[7208]_ ,
    \new_[7209]_ , \new_[7210]_ , \new_[7211]_ , \new_[7212]_ ,
    \new_[7213]_ , \new_[7214]_ , \new_[7215]_ , \new_[7216]_ ,
    \new_[7217]_ , \new_[7218]_ , \new_[7219]_ , \new_[7220]_ ,
    \new_[7221]_ , \new_[7222]_ , \new_[7223]_ , \new_[7224]_ ,
    \new_[7225]_ , \new_[7226]_ , \new_[7227]_ , \new_[7228]_ ,
    \new_[7229]_ , \new_[7230]_ , \new_[7231]_ , \new_[7232]_ ,
    \new_[7233]_ , \new_[7234]_ , \new_[7235]_ , \new_[7236]_ ,
    \new_[7237]_ , \new_[7238]_ , \new_[7239]_ , \new_[7240]_ ,
    \new_[7241]_ , \new_[7242]_ , \new_[7243]_ , \new_[7244]_ ,
    \new_[7245]_ , \new_[7246]_ , \new_[7247]_ , \new_[7248]_ ,
    \new_[7249]_ , \new_[7250]_ , \new_[7251]_ , \new_[7252]_ ,
    \new_[7253]_ , \new_[7254]_ , \new_[7255]_ , \new_[7256]_ ,
    \new_[7257]_ , \new_[7258]_ , \new_[7259]_ , \new_[7260]_ ,
    \new_[7261]_ , \new_[7262]_ , \new_[7263]_ , \new_[7264]_ ,
    \new_[7265]_ , \new_[7266]_ , \new_[7267]_ , \new_[7268]_ ,
    \new_[7269]_ , \new_[7270]_ , \new_[7271]_ , \new_[7272]_ ,
    \new_[7273]_ , \new_[7274]_ , \new_[7275]_ , \new_[7276]_ ,
    \new_[7277]_ , \new_[7278]_ , \new_[7279]_ , \new_[7280]_ ,
    \new_[7281]_ , \new_[7282]_ , \new_[7283]_ , \new_[7284]_ ,
    \new_[7285]_ , \new_[7286]_ , \new_[7287]_ , \new_[7288]_ ,
    \new_[7289]_ , \new_[7290]_ , \new_[7291]_ , \new_[7292]_ ,
    \new_[7293]_ , \new_[7294]_ , \new_[7295]_ , \new_[7296]_ ,
    \new_[7297]_ , \new_[7298]_ , \new_[7299]_ , \new_[7300]_ ,
    \new_[7301]_ , \new_[7302]_ , \new_[7303]_ , \new_[7304]_ ,
    \new_[7305]_ , \new_[7306]_ , \new_[7307]_ , \new_[7308]_ ,
    \new_[7309]_ , \new_[7310]_ , \new_[7311]_ , \new_[7312]_ ,
    \new_[7313]_ , \new_[7314]_ , \new_[7315]_ , \new_[7316]_ ,
    \new_[7317]_ , \new_[7318]_ , \new_[7319]_ , \new_[7320]_ ,
    \new_[7321]_ , \new_[7322]_ , \new_[7323]_ , \new_[7324]_ ,
    \new_[7325]_ , \new_[7326]_ , \new_[7327]_ , \new_[7328]_ ,
    \new_[7329]_ , \new_[7330]_ , \new_[7331]_ , \new_[7332]_ ,
    \new_[7333]_ , \new_[7334]_ , \new_[7335]_ , \new_[7336]_ ,
    \new_[7337]_ , \new_[7338]_ , \new_[7339]_ , \new_[7340]_ ,
    \new_[7341]_ , \new_[7342]_ , \new_[7343]_ , \new_[7344]_ ,
    \new_[7345]_ , \new_[7346]_ , \new_[7347]_ , \new_[7348]_ ,
    \new_[7349]_ , \new_[7350]_ , \new_[7351]_ , \new_[7352]_ ,
    \new_[7353]_ , \new_[7354]_ , \new_[7355]_ , \new_[7356]_ ,
    \new_[7357]_ , \new_[7358]_ , \new_[7359]_ , \new_[7360]_ ,
    \new_[7361]_ , \new_[7362]_ , \new_[7363]_ , \new_[7364]_ ,
    \new_[7365]_ , \new_[7366]_ , \new_[7367]_ , \new_[7368]_ ,
    \new_[7369]_ , \new_[7370]_ , \new_[7371]_ , \new_[7372]_ ,
    \new_[7373]_ , \new_[7374]_ , \new_[7375]_ , \new_[7376]_ ,
    \new_[7377]_ , \new_[7378]_ , \new_[7379]_ , \new_[7380]_ ,
    \new_[7381]_ , \new_[7382]_ , \new_[7383]_ , \new_[7384]_ ,
    \new_[7385]_ , \new_[7386]_ , \new_[7387]_ , \new_[7388]_ ,
    \new_[7389]_ , \new_[7390]_ , \new_[7391]_ , \new_[7392]_ ,
    \new_[7393]_ , \new_[7394]_ , \new_[7395]_ , \new_[7396]_ ,
    \new_[7397]_ , \new_[7398]_ , \new_[7399]_ , \new_[7400]_ ,
    \new_[7401]_ , \new_[7402]_ , \new_[7403]_ , \new_[7404]_ ,
    \new_[7405]_ , \new_[7406]_ , \new_[7407]_ , \new_[7408]_ ,
    \new_[7409]_ , \new_[7410]_ , \new_[7411]_ , \new_[7412]_ ,
    \new_[7413]_ , \new_[7414]_ , \new_[7415]_ , \new_[7416]_ ,
    \new_[7417]_ , \new_[7418]_ , \new_[7419]_ , \new_[7420]_ ,
    \new_[7421]_ , \new_[7422]_ , \new_[7423]_ , \new_[7424]_ ,
    \new_[7425]_ , \new_[7426]_ , \new_[7427]_ , \new_[7428]_ ,
    \new_[7429]_ , \new_[7430]_ , \new_[7431]_ , \new_[7432]_ ,
    \new_[7433]_ , \new_[7434]_ , \new_[7435]_ , \new_[7436]_ ,
    \new_[7437]_ , \new_[7438]_ , \new_[7439]_ , \new_[7440]_ ,
    \new_[7441]_ , \new_[7442]_ , \new_[7443]_ , \new_[7444]_ ,
    \new_[7445]_ , \new_[7446]_ , \new_[7447]_ , \new_[7448]_ ,
    \new_[7449]_ , \new_[7450]_ , \new_[7451]_ , \new_[7452]_ ,
    \new_[7453]_ , \new_[7454]_ , \new_[7455]_ , \new_[7456]_ ,
    \new_[7457]_ , \new_[7458]_ , \new_[7459]_ , \new_[7460]_ ,
    \new_[7461]_ , \new_[7462]_ , \new_[7463]_ , \new_[7464]_ ,
    \new_[7465]_ , \new_[7466]_ , \new_[7467]_ , \new_[7468]_ ,
    \new_[7469]_ , \new_[7470]_ , \new_[7471]_ , \new_[7472]_ ,
    \new_[7473]_ , \new_[7474]_ , \new_[7475]_ , \new_[7476]_ ,
    \new_[7477]_ , \new_[7478]_ , \new_[7479]_ , \new_[7480]_ ,
    \new_[7481]_ , \new_[7482]_ , \new_[7483]_ , \new_[7484]_ ,
    \new_[7485]_ , \new_[7486]_ , \new_[7487]_ , \new_[7488]_ ,
    \new_[7489]_ , \new_[7490]_ , \new_[7491]_ , \new_[7492]_ ,
    \new_[7493]_ , \new_[7494]_ , \new_[7495]_ , \new_[7496]_ ,
    \new_[7497]_ , \new_[7498]_ , \new_[7499]_ , \new_[7500]_ ,
    \new_[7501]_ , \new_[7502]_ , \new_[7503]_ , \new_[7504]_ ,
    \new_[7505]_ , \new_[7506]_ , \new_[7507]_ , \new_[7508]_ ,
    \new_[7509]_ , \new_[7510]_ , \new_[7511]_ , \new_[7512]_ ,
    \new_[7513]_ , \new_[7514]_ , \new_[7515]_ , \new_[7516]_ ,
    \new_[7517]_ , \new_[7518]_ , \new_[7519]_ , \new_[7520]_ ,
    \new_[7521]_ , \new_[7522]_ , \new_[7523]_ , \new_[7524]_ ,
    \new_[7525]_ , \new_[7526]_ , \new_[7527]_ , \new_[7528]_ ,
    \new_[7529]_ , \new_[7530]_ , \new_[7531]_ , \new_[7532]_ ,
    \new_[7533]_ , \new_[7534]_ , \new_[7535]_ , \new_[7536]_ ,
    \new_[7537]_ , \new_[7538]_ , \new_[7539]_ , \new_[7540]_ ,
    \new_[7541]_ , \new_[7542]_ , \new_[7543]_ , \new_[7544]_ ,
    \new_[7545]_ , \new_[7546]_ , \new_[7547]_ , \new_[7548]_ ,
    \new_[7549]_ , \new_[7550]_ , \new_[7551]_ , \new_[7552]_ ,
    \new_[7553]_ , \new_[7554]_ , \new_[7555]_ , \new_[7556]_ ,
    \new_[7557]_ , \new_[7558]_ , \new_[7559]_ , \new_[7560]_ ,
    \new_[7561]_ , \new_[7562]_ , \new_[7563]_ , \new_[7564]_ ,
    \new_[7565]_ , \new_[7566]_ , \new_[7567]_ , \new_[7568]_ ,
    \new_[7569]_ , \new_[7570]_ , \new_[7571]_ , \new_[7572]_ ,
    \new_[7573]_ , \new_[7574]_ , \new_[7575]_ , \new_[7576]_ ,
    \new_[7577]_ , \new_[7578]_ , \new_[7579]_ , \new_[7580]_ ,
    \new_[7581]_ , \new_[7582]_ , \new_[7583]_ , \new_[7584]_ ,
    \new_[7585]_ , \new_[7586]_ , \new_[7587]_ , \new_[7588]_ ,
    \new_[7589]_ , \new_[7590]_ , \new_[7591]_ , \new_[7592]_ ,
    \new_[7593]_ , \new_[7594]_ , \new_[7595]_ , \new_[7596]_ ,
    \new_[7597]_ , \new_[7598]_ , \new_[7599]_ , \new_[7600]_ ,
    \new_[7601]_ , \new_[7602]_ , \new_[7603]_ , \new_[7604]_ ,
    \new_[7605]_ , \new_[7606]_ , \new_[7607]_ , \new_[7608]_ ,
    \new_[7609]_ , \new_[7610]_ , \new_[7611]_ , \new_[7612]_ ,
    \new_[7613]_ , \new_[7614]_ , \new_[7615]_ , \new_[7616]_ ,
    \new_[7617]_ , \new_[7618]_ , \new_[7619]_ , \new_[7620]_ ,
    \new_[7621]_ , \new_[7622]_ , \new_[7623]_ , \new_[7624]_ ,
    \new_[7625]_ , \new_[7626]_ , \new_[7627]_ , \new_[7628]_ ,
    \new_[7629]_ , \new_[7630]_ , \new_[7631]_ , \new_[7632]_ ,
    \new_[7633]_ , \new_[7634]_ , \new_[7635]_ , \new_[7636]_ ,
    \new_[7637]_ , \new_[7638]_ , \new_[7639]_ , \new_[7640]_ ,
    \new_[7641]_ , \new_[7642]_ , \new_[7643]_ , \new_[7644]_ ,
    \new_[7645]_ , \new_[7646]_ , \new_[7647]_ , \new_[7648]_ ,
    \new_[7649]_ , \new_[7650]_ , \new_[7651]_ , \new_[7652]_ ,
    \new_[7653]_ , \new_[7654]_ , \new_[7655]_ , \new_[7656]_ ,
    \new_[7657]_ , \new_[7658]_ , \new_[7659]_ , \new_[7660]_ ,
    \new_[7661]_ , \new_[7662]_ , \new_[7663]_ , \new_[7664]_ ,
    \new_[7665]_ , \new_[7666]_ , \new_[7667]_ , \new_[7668]_ ,
    \new_[7669]_ , \new_[7670]_ , \new_[7671]_ , \new_[7672]_ ,
    \new_[7673]_ , \new_[7674]_ , \new_[7675]_ , \new_[7676]_ ,
    \new_[7677]_ , \new_[7678]_ , \new_[7679]_ , \new_[7680]_ ,
    \new_[7681]_ , \new_[7682]_ , \new_[7683]_ , \new_[7684]_ ,
    \new_[7685]_ , \new_[7686]_ , \new_[7687]_ , \new_[7688]_ ,
    \new_[7689]_ , \new_[7690]_ , \new_[7691]_ , \new_[7692]_ ,
    \new_[7693]_ , \new_[7694]_ , \new_[7695]_ , \new_[7696]_ ,
    \new_[7697]_ , \new_[7698]_ , \new_[7699]_ , \new_[7700]_ ,
    \new_[7701]_ , \new_[7702]_ , \new_[7703]_ , \new_[7704]_ ,
    \new_[7705]_ , \new_[7706]_ , \new_[7707]_ , \new_[7708]_ ,
    \new_[7709]_ , \new_[7710]_ , \new_[7711]_ , \new_[7712]_ ,
    \new_[7713]_ , \new_[7714]_ , \new_[7715]_ , \new_[7716]_ ,
    \new_[7717]_ , \new_[7718]_ , \new_[7719]_ , \new_[7720]_ ,
    \new_[7721]_ , \new_[7722]_ , \new_[7723]_ , \new_[7724]_ ,
    \new_[7725]_ , \new_[7726]_ , \new_[7727]_ , \new_[7728]_ ,
    \new_[7729]_ , \new_[7730]_ , \new_[7731]_ , \new_[7732]_ ,
    \new_[7733]_ , \new_[7734]_ , \new_[7735]_ , \new_[7736]_ ,
    \new_[7737]_ , \new_[7738]_ , \new_[7739]_ , \new_[7740]_ ,
    \new_[7741]_ , \new_[7742]_ , \new_[7743]_ , \new_[7744]_ ,
    \new_[7745]_ , \new_[7746]_ , \new_[7747]_ , \new_[7748]_ ,
    \new_[7749]_ , \new_[7750]_ , \new_[7751]_ , \new_[7752]_ ,
    \new_[7753]_ , \new_[7754]_ , \new_[7755]_ , \new_[7756]_ ,
    \new_[7757]_ , \new_[7758]_ , \new_[7759]_ , \new_[7760]_ ,
    \new_[7761]_ , \new_[7762]_ , \new_[7763]_ , \new_[7764]_ ,
    \new_[7765]_ , \new_[7766]_ , \new_[7767]_ , \new_[7768]_ ,
    \new_[7769]_ , \new_[7770]_ , \new_[7771]_ , \new_[7772]_ ,
    \new_[7773]_ , \new_[7774]_ , \new_[7775]_ , \new_[7776]_ ,
    \new_[7777]_ , \new_[7778]_ , \new_[7779]_ , \new_[7780]_ ,
    \new_[7781]_ , \new_[7782]_ , \new_[7783]_ , \new_[7784]_ ,
    \new_[7785]_ , \new_[7786]_ , \new_[7787]_ , \new_[7788]_ ,
    \new_[7789]_ , \new_[7790]_ , \new_[7791]_ , \new_[7792]_ ,
    \new_[7793]_ , \new_[7794]_ , \new_[7795]_ , \new_[7796]_ ,
    \new_[7797]_ , \new_[7798]_ , \new_[7799]_ , \new_[7800]_ ,
    \new_[7801]_ , \new_[7802]_ , \new_[7803]_ , \new_[7804]_ ,
    \new_[7805]_ , \new_[7806]_ , \new_[7807]_ , \new_[7808]_ ,
    \new_[7809]_ , \new_[7810]_ , \new_[7811]_ , \new_[7812]_ ,
    \new_[7813]_ , \new_[7814]_ , \new_[7815]_ , \new_[7816]_ ,
    \new_[7817]_ , \new_[7818]_ , \new_[7819]_ , \new_[7820]_ ,
    \new_[7821]_ , \new_[7822]_ , \new_[7823]_ , \new_[7824]_ ,
    \new_[7825]_ , \new_[7826]_ , \new_[7827]_ , \new_[7828]_ ,
    \new_[7829]_ , \new_[7830]_ , \new_[7831]_ , \new_[7832]_ ,
    \new_[7833]_ , \new_[7834]_ , \new_[7835]_ , \new_[7836]_ ,
    \new_[7837]_ , \new_[7838]_ , \new_[7839]_ , \new_[7840]_ ,
    \new_[7841]_ , \new_[7842]_ , \new_[7843]_ , \new_[7844]_ ,
    \new_[7845]_ , \new_[7846]_ , \new_[7847]_ , \new_[7848]_ ,
    \new_[7849]_ , \new_[7850]_ , \new_[7851]_ , \new_[7852]_ ,
    \new_[7853]_ , \new_[7854]_ , \new_[7855]_ , \new_[7856]_ ,
    \new_[7857]_ , \new_[7858]_ , \new_[7859]_ , \new_[7860]_ ,
    \new_[7861]_ , \new_[7862]_ , \new_[7863]_ , \new_[7864]_ ,
    \new_[7865]_ , \new_[7866]_ , \new_[7867]_ , \new_[7868]_ ,
    \new_[7869]_ , \new_[7870]_ , \new_[7871]_ , \new_[7872]_ ,
    \new_[7873]_ , \new_[7874]_ , \new_[7875]_ , \new_[7876]_ ,
    \new_[7877]_ , \new_[7878]_ , \new_[7879]_ , \new_[7880]_ ,
    \new_[7881]_ , \new_[7882]_ , \new_[7883]_ , \new_[7884]_ ,
    \new_[7885]_ , \new_[7886]_ , \new_[7887]_ , \new_[7888]_ ,
    \new_[7889]_ , \new_[7890]_ , \new_[7891]_ , \new_[7892]_ ,
    \new_[7893]_ , \new_[7894]_ , \new_[7895]_ , \new_[7896]_ ,
    \new_[7897]_ , \new_[7898]_ , \new_[7899]_ , \new_[7900]_ ,
    \new_[7901]_ , \new_[7902]_ , \new_[7903]_ , \new_[7904]_ ,
    \new_[7905]_ , \new_[7906]_ , \new_[7907]_ , \new_[7908]_ ,
    \new_[7909]_ , \new_[7910]_ , \new_[7911]_ , \new_[7912]_ ,
    \new_[7913]_ , \new_[7914]_ , \new_[7915]_ , \new_[7916]_ ,
    \new_[7917]_ , \new_[7918]_ , \new_[7919]_ , \new_[7920]_ ,
    \new_[7921]_ , \new_[7922]_ , \new_[7923]_ , \new_[7924]_ ,
    \new_[7925]_ , \new_[7926]_ , \new_[7927]_ , \new_[7928]_ ,
    \new_[7929]_ , \new_[7930]_ , \new_[7931]_ , \new_[7932]_ ,
    \new_[7933]_ , \new_[7934]_ , \new_[7935]_ , \new_[7936]_ ,
    \new_[7937]_ , \new_[7938]_ , \new_[7939]_ , \new_[7940]_ ,
    \new_[7941]_ , \new_[7942]_ , \new_[7943]_ , \new_[7944]_ ,
    \new_[7945]_ , \new_[7946]_ , \new_[7947]_ , \new_[7948]_ ,
    \new_[7949]_ , \new_[7950]_ , \new_[7951]_ , \new_[7952]_ ,
    \new_[7953]_ , \new_[7954]_ , \new_[7955]_ , \new_[7956]_ ,
    \new_[7957]_ , \new_[7958]_ , \new_[7959]_ , \new_[7960]_ ,
    \new_[7961]_ , \new_[7962]_ , \new_[7963]_ , \new_[7964]_ ,
    \new_[7965]_ , \new_[7966]_ , \new_[7967]_ , \new_[7968]_ ,
    \new_[7969]_ , \new_[7970]_ , \new_[7971]_ , \new_[7972]_ ,
    \new_[7973]_ , \new_[7974]_ , \new_[7975]_ , \new_[7976]_ ,
    \new_[7977]_ , \new_[7978]_ , \new_[7979]_ , \new_[7980]_ ,
    \new_[7981]_ , \new_[7982]_ , \new_[7983]_ , \new_[7984]_ ,
    \new_[7985]_ , \new_[7986]_ , \new_[7987]_ , \new_[7988]_ ,
    \new_[7989]_ , \new_[7990]_ , \new_[7991]_ , \new_[7992]_ ,
    \new_[7993]_ , \new_[7994]_ , \new_[7995]_ , \new_[7996]_ ,
    \new_[7997]_ , \new_[7998]_ , \new_[7999]_ , \new_[8000]_ ,
    \new_[8001]_ , \new_[8002]_ , \new_[8003]_ , \new_[8004]_ ,
    \new_[8005]_ , \new_[8006]_ , \new_[8007]_ , \new_[8008]_ ,
    \new_[8009]_ , \new_[8010]_ , \new_[8011]_ , \new_[8012]_ ,
    \new_[8013]_ , \new_[8014]_ , \new_[8015]_ , \new_[8016]_ ,
    \new_[8017]_ , \new_[8018]_ , \new_[8019]_ , \new_[8020]_ ,
    \new_[8021]_ , \new_[8022]_ , \new_[8023]_ , \new_[8024]_ ,
    \new_[8025]_ , \new_[8026]_ , \new_[8027]_ , \new_[8028]_ ,
    \new_[8029]_ , \new_[8030]_ , \new_[8031]_ , \new_[8032]_ ,
    \new_[8033]_ , \new_[8034]_ , \new_[8035]_ , \new_[8036]_ ,
    \new_[8037]_ , \new_[8038]_ , \new_[8039]_ , \new_[8040]_ ,
    \new_[8041]_ , \new_[8043]_ , \new_[8044]_ , \new_[8045]_ ,
    \new_[8046]_ , \new_[8047]_ , \new_[8048]_ , \new_[8049]_ ,
    \new_[8050]_ , \new_[8051]_ , \new_[8052]_ , \new_[8053]_ ,
    \new_[8054]_ , \new_[8055]_ , \new_[8056]_ , \new_[8057]_ ,
    \new_[8058]_ , \new_[8059]_ , \new_[8060]_ , \new_[8061]_ ,
    \new_[8062]_ , \new_[8063]_ , \new_[8064]_ , \new_[8065]_ ,
    \new_[8066]_ , \new_[8067]_ , \new_[8068]_ , \new_[8069]_ ,
    \new_[8070]_ , \new_[8071]_ , \new_[8072]_ , \new_[8073]_ ,
    \new_[8074]_ , \new_[8075]_ , \new_[8076]_ , \new_[8077]_ ,
    \new_[8078]_ , \new_[8079]_ , \new_[8080]_ , \new_[8081]_ ,
    \new_[8082]_ , \new_[8083]_ , \new_[8084]_ , \new_[8085]_ ,
    \new_[8086]_ , \new_[8087]_ , \new_[8088]_ , \new_[8089]_ ,
    \new_[8090]_ , \new_[8091]_ , \new_[8092]_ , \new_[8093]_ ,
    \new_[8094]_ , \new_[8095]_ , \new_[8096]_ , \new_[8097]_ ,
    \new_[8098]_ , \new_[8099]_ , \new_[8100]_ , \new_[8101]_ ,
    \new_[8102]_ , \new_[8103]_ , \new_[8104]_ , \new_[8105]_ ,
    \new_[8106]_ , \new_[8107]_ , \new_[8108]_ , \new_[8109]_ ,
    \new_[8110]_ , \new_[8111]_ , \new_[8112]_ , \new_[8113]_ ,
    \new_[8114]_ , \new_[8115]_ , \new_[8116]_ , \new_[8119]_ ,
    \new_[8120]_ , \new_[8121]_ , \new_[8122]_ , \new_[8123]_ ,
    \new_[8124]_ , \new_[8125]_ , \new_[8126]_ , \new_[8127]_ ,
    \new_[8128]_ , \new_[8129]_ , \new_[8130]_ , \new_[8131]_ ,
    \new_[8132]_ , \new_[8133]_ , \new_[8134]_ , \new_[8135]_ ,
    \new_[8136]_ , \new_[8137]_ , \new_[8138]_ , \new_[8139]_ ,
    \new_[8140]_ , \new_[8141]_ , \new_[8142]_ , \new_[8143]_ ,
    \new_[8144]_ , \new_[8145]_ , \new_[8146]_ , \new_[8147]_ ,
    \new_[8148]_ , \new_[8149]_ , \new_[8150]_ , \new_[8151]_ ,
    \new_[8152]_ , \new_[8153]_ , \new_[8154]_ , \new_[8155]_ ,
    \new_[8156]_ , \new_[8157]_ , \new_[8158]_ , \new_[8159]_ ,
    \new_[8160]_ , \new_[8161]_ , \new_[8162]_ , \new_[8163]_ ,
    \new_[8164]_ , \new_[8165]_ , \new_[8166]_ , \new_[8167]_ ,
    \new_[8168]_ , \new_[8169]_ , \new_[8170]_ , \new_[8171]_ ,
    \new_[8172]_ , \new_[8173]_ , \new_[8174]_ , \new_[8175]_ ,
    \new_[8176]_ , \new_[8177]_ , \new_[8178]_ , \new_[8179]_ ,
    \new_[8180]_ , \new_[8181]_ , \new_[8182]_ , \new_[8183]_ ,
    \new_[8184]_ , \new_[8185]_ , \new_[8186]_ , \new_[8187]_ ,
    \new_[8188]_ , \new_[8189]_ , \new_[8190]_ , \new_[8191]_ ,
    \new_[8192]_ , \new_[8193]_ , \new_[8194]_ , \new_[8195]_ ,
    \new_[8196]_ , \new_[8197]_ , \new_[8198]_ , \new_[8199]_ ,
    \new_[8200]_ , \new_[8201]_ , \new_[8202]_ , \new_[8203]_ ,
    \new_[8204]_ , \new_[8205]_ , \new_[8206]_ , \new_[8207]_ ,
    \new_[8208]_ , \new_[8209]_ , \new_[8210]_ , \new_[8211]_ ,
    \new_[8212]_ , \new_[8213]_ , \new_[8214]_ , \new_[8215]_ ,
    \new_[8216]_ , \new_[8217]_ , \new_[8218]_ , \new_[8219]_ ,
    \new_[8220]_ , \new_[8221]_ , \new_[8222]_ , \new_[8223]_ ,
    \new_[8224]_ , \new_[8225]_ , \new_[8226]_ , \new_[8227]_ ,
    \new_[8228]_ , \new_[8229]_ , \new_[8230]_ , \new_[8231]_ ,
    \new_[8232]_ , \new_[8233]_ , \new_[8234]_ , \new_[8235]_ ,
    \new_[8236]_ , \new_[8237]_ , \new_[8238]_ , \new_[8239]_ ,
    \new_[8240]_ , \new_[8241]_ , \new_[8242]_ , \new_[8243]_ ,
    \new_[8244]_ , \new_[8245]_ , \new_[8246]_ , \new_[8247]_ ,
    \new_[8248]_ , \new_[8249]_ , \new_[8250]_ , \new_[8251]_ ,
    \new_[8252]_ , \new_[8253]_ , \new_[8254]_ , \new_[8255]_ ,
    \new_[8256]_ , \new_[8257]_ , \new_[8258]_ , \new_[8259]_ ,
    \new_[8260]_ , \new_[8261]_ , \new_[8262]_ , \new_[8263]_ ,
    \new_[8264]_ , \new_[8265]_ , \new_[8266]_ , \new_[8267]_ ,
    \new_[8268]_ , \new_[8269]_ , \new_[8270]_ , \new_[8271]_ ,
    \new_[8272]_ , \new_[8273]_ , \new_[8274]_ , \new_[8275]_ ,
    \new_[8276]_ , \new_[8277]_ , \new_[8278]_ , \new_[8279]_ ,
    \new_[8280]_ , \new_[8281]_ , \new_[8282]_ , \new_[8283]_ ,
    \new_[8284]_ , \new_[8285]_ , \new_[8286]_ , \new_[8287]_ ,
    \new_[8288]_ , \new_[8289]_ , \new_[8290]_ , \new_[8291]_ ,
    \new_[8292]_ , \new_[8293]_ , \new_[8294]_ , \new_[8295]_ ,
    \new_[8296]_ , \new_[8297]_ , \new_[8298]_ , \new_[8299]_ ,
    \new_[8300]_ , \new_[8301]_ , \new_[8302]_ , \new_[8303]_ ,
    \new_[8304]_ , \new_[8305]_ , \new_[8306]_ , \new_[8307]_ ,
    \new_[8308]_ , \new_[8309]_ , \new_[8310]_ , \new_[8311]_ ,
    \new_[8312]_ , \new_[8313]_ , \new_[8314]_ , \new_[8315]_ ,
    \new_[8316]_ , \new_[8317]_ , \new_[8318]_ , \new_[8319]_ ,
    \new_[8320]_ , \new_[8321]_ , \new_[8322]_ , \new_[8323]_ ,
    \new_[8324]_ , \new_[8325]_ , \new_[8326]_ , \new_[8327]_ ,
    \new_[8328]_ , \new_[8329]_ , \new_[8330]_ , \new_[8331]_ ,
    \new_[8332]_ , \new_[8333]_ , \new_[8334]_ , \new_[8335]_ ,
    \new_[8336]_ , \new_[8337]_ , \new_[8338]_ , \new_[8339]_ ,
    \new_[8340]_ , \new_[8341]_ , \new_[8342]_ , \new_[8343]_ ,
    \new_[8344]_ , \new_[8345]_ , \new_[8346]_ , \new_[8347]_ ,
    \new_[8348]_ , \new_[8349]_ , \new_[8350]_ , \new_[8351]_ ,
    \new_[8352]_ , \new_[8353]_ , \new_[8354]_ , \new_[8355]_ ,
    \new_[8356]_ , \new_[8357]_ , \new_[8358]_ , \new_[8359]_ ,
    \new_[8360]_ , \new_[8361]_ , \new_[8362]_ , \new_[8363]_ ,
    \new_[8364]_ , \new_[8365]_ , \new_[8366]_ , \new_[8367]_ ,
    \new_[8368]_ , \new_[8369]_ , \new_[8370]_ , \new_[8371]_ ,
    \new_[8372]_ , \new_[8373]_ , \new_[8374]_ , \new_[8375]_ ,
    \new_[8376]_ , \new_[8377]_ , \new_[8378]_ , \new_[8379]_ ,
    \new_[8380]_ , \new_[8381]_ , \new_[8382]_ , \new_[8383]_ ,
    \new_[8384]_ , \new_[8385]_ , \new_[8386]_ , \new_[8387]_ ,
    \new_[8388]_ , \new_[8389]_ , \new_[8390]_ , \new_[8391]_ ,
    \new_[8392]_ , \new_[8393]_ , \new_[8394]_ , \new_[8395]_ ,
    \new_[8396]_ , \new_[8397]_ , \new_[8398]_ , \new_[8399]_ ,
    \new_[8400]_ , \new_[8401]_ , \new_[8402]_ , \new_[8403]_ ,
    \new_[8404]_ , \new_[8405]_ , \new_[8406]_ , \new_[8407]_ ,
    \new_[8408]_ , \new_[8409]_ , \new_[8410]_ , \new_[8411]_ ,
    \new_[8412]_ , \new_[8413]_ , \new_[8414]_ , \new_[8415]_ ,
    \new_[8416]_ , \new_[8417]_ , \new_[8418]_ , \new_[8419]_ ,
    \new_[8420]_ , \new_[8421]_ , \new_[8422]_ , \new_[8423]_ ,
    \new_[8424]_ , \new_[8425]_ , \new_[8426]_ , \new_[8427]_ ,
    \new_[8428]_ , \new_[8429]_ , \new_[8430]_ , \new_[8431]_ ,
    \new_[8432]_ , \new_[8433]_ , \new_[8434]_ , \new_[8435]_ ,
    \new_[8436]_ , \new_[8437]_ , \new_[8438]_ , \new_[8439]_ ,
    \new_[8440]_ , \new_[8441]_ , \new_[8442]_ , \new_[8443]_ ,
    \new_[8444]_ , \new_[8445]_ , \new_[8446]_ , \new_[8447]_ ,
    \new_[8448]_ , \new_[8449]_ , \new_[8450]_ , \new_[8451]_ ,
    \new_[8452]_ , \new_[8453]_ , \new_[8454]_ , \new_[8455]_ ,
    \new_[8456]_ , \new_[8457]_ , \new_[8458]_ , \new_[8459]_ ,
    \new_[8460]_ , \new_[8461]_ , \new_[8462]_ , \new_[8463]_ ,
    \new_[8464]_ , \new_[8465]_ , \new_[8466]_ , \new_[8467]_ ,
    \new_[8468]_ , \new_[8469]_ , \new_[8470]_ , \new_[8471]_ ,
    \new_[8472]_ , \new_[8473]_ , \new_[8474]_ , \new_[8475]_ ,
    \new_[8476]_ , \new_[8477]_ , \new_[8478]_ , \new_[8479]_ ,
    \new_[8480]_ , \new_[8481]_ , \new_[8482]_ , \new_[8483]_ ,
    \new_[8484]_ , \new_[8485]_ , \new_[8486]_ , \new_[8487]_ ,
    \new_[8488]_ , \new_[8489]_ , \new_[8490]_ , \new_[8491]_ ,
    \new_[8492]_ , \new_[8493]_ , \new_[8494]_ , \new_[8495]_ ,
    \new_[8496]_ , \new_[8497]_ , \new_[8498]_ , \new_[8499]_ ,
    \new_[8500]_ , \new_[8501]_ , \new_[8502]_ , \new_[8503]_ ,
    \new_[8504]_ , \new_[8505]_ , \new_[8506]_ , \new_[8507]_ ,
    \new_[8509]_ , \new_[8510]_ , \new_[8511]_ , \new_[8512]_ ,
    \new_[8513]_ , \new_[8514]_ , \new_[8515]_ , \new_[8516]_ ,
    \new_[8517]_ , \new_[8518]_ , \new_[8519]_ , \new_[8520]_ ,
    \new_[8521]_ , \new_[8522]_ , \new_[8523]_ , \new_[8524]_ ,
    \new_[8525]_ , \new_[8526]_ , \new_[8527]_ , \new_[8528]_ ,
    \new_[8529]_ , \new_[8530]_ , \new_[8531]_ , \new_[8532]_ ,
    \new_[8533]_ , \new_[8534]_ , \new_[8535]_ , \new_[8536]_ ,
    \new_[8537]_ , \new_[8538]_ , \new_[8539]_ , \new_[8540]_ ,
    \new_[8541]_ , \new_[8542]_ , \new_[8543]_ , \new_[8544]_ ,
    \new_[8545]_ , \new_[8546]_ , \new_[8547]_ , \new_[8548]_ ,
    \new_[8549]_ , \new_[8550]_ , \new_[8551]_ , \new_[8552]_ ,
    \new_[8553]_ , \new_[8554]_ , \new_[8555]_ , \new_[8556]_ ,
    \new_[8557]_ , \new_[8558]_ , \new_[8559]_ , \new_[8560]_ ,
    \new_[8561]_ , \new_[8562]_ , \new_[8563]_ , \new_[8564]_ ,
    \new_[8565]_ , \new_[8566]_ , \new_[8567]_ , \new_[8568]_ ,
    \new_[8569]_ , \new_[8570]_ , \new_[8571]_ , \new_[8572]_ ,
    \new_[8573]_ , \new_[8574]_ , \new_[8575]_ , \new_[8576]_ ,
    \new_[8577]_ , \new_[8578]_ , \new_[8579]_ , \new_[8580]_ ,
    \new_[8581]_ , \new_[8582]_ , \new_[8583]_ , \new_[8584]_ ,
    \new_[8585]_ , \new_[8586]_ , \new_[8587]_ , \new_[8588]_ ,
    \new_[8589]_ , \new_[8590]_ , \new_[8591]_ , \new_[8592]_ ,
    \new_[8593]_ , \new_[8594]_ , \new_[8595]_ , \new_[8596]_ ,
    \new_[8597]_ , \new_[8598]_ , \new_[8599]_ , \new_[8600]_ ,
    \new_[8601]_ , \new_[8602]_ , \new_[8603]_ , \new_[8604]_ ,
    \new_[8605]_ , \new_[8606]_ , \new_[8607]_ , \new_[8608]_ ,
    \new_[8609]_ , \new_[8610]_ , \new_[8611]_ , \new_[8612]_ ,
    \new_[8613]_ , \new_[8614]_ , \new_[8615]_ , \new_[8616]_ ,
    \new_[8617]_ , \new_[8618]_ , \new_[8619]_ , \new_[8620]_ ,
    \new_[8621]_ , \new_[8622]_ , \new_[8623]_ , \new_[8624]_ ,
    \new_[8625]_ , \new_[8626]_ , \new_[8627]_ , \new_[8628]_ ,
    \new_[8629]_ , \new_[8630]_ , \new_[8631]_ , \new_[8632]_ ,
    \new_[8633]_ , \new_[8634]_ , \new_[8635]_ , \new_[8636]_ ,
    \new_[8637]_ , \new_[8638]_ , \new_[8639]_ , \new_[8640]_ ,
    \new_[8641]_ , \new_[8642]_ , \new_[8643]_ , \new_[8644]_ ,
    \new_[8645]_ , \new_[8646]_ , \new_[8647]_ , \new_[8648]_ ,
    \new_[8649]_ , \new_[8650]_ , \new_[8651]_ , \new_[8652]_ ,
    \new_[8653]_ , \new_[8654]_ , \new_[8655]_ , \new_[8656]_ ,
    \new_[8657]_ , \new_[8658]_ , \new_[8659]_ , \new_[8660]_ ,
    \new_[8661]_ , \new_[8662]_ , \new_[8663]_ , \new_[8664]_ ,
    \new_[8665]_ , \new_[8666]_ , \new_[8667]_ , \new_[8668]_ ,
    \new_[8669]_ , \new_[8670]_ , \new_[8671]_ , \new_[8672]_ ,
    \new_[8673]_ , \new_[8674]_ , \new_[8675]_ , \new_[8676]_ ,
    \new_[8677]_ , \new_[8678]_ , \new_[8679]_ , \new_[8680]_ ,
    \new_[8681]_ , \new_[8682]_ , \new_[8683]_ , \new_[8684]_ ,
    \new_[8685]_ , \new_[8686]_ , \new_[8687]_ , \new_[8688]_ ,
    \new_[8689]_ , \new_[8690]_ , \new_[8691]_ , \new_[8692]_ ,
    \new_[8693]_ , \new_[8694]_ , \new_[8695]_ , \new_[8696]_ ,
    \new_[8697]_ , \new_[8698]_ , \new_[8699]_ , \new_[8700]_ ,
    \new_[8701]_ , \new_[8702]_ , \new_[8703]_ , \new_[8704]_ ,
    \new_[8705]_ , \new_[8706]_ , \new_[8707]_ , \new_[8708]_ ,
    \new_[8709]_ , \new_[8710]_ , \new_[8711]_ , \new_[8712]_ ,
    \new_[8713]_ , \new_[8714]_ , \new_[8715]_ , \new_[8716]_ ,
    \new_[8717]_ , \new_[8718]_ , \new_[8719]_ , \new_[8720]_ ,
    \new_[8721]_ , \new_[8722]_ , \new_[8723]_ , \new_[8724]_ ,
    \new_[8725]_ , \new_[8726]_ , \new_[8727]_ , \new_[8728]_ ,
    \new_[8729]_ , \new_[8730]_ , \new_[8731]_ , \new_[8732]_ ,
    \new_[8733]_ , \new_[8734]_ , \new_[8735]_ , \new_[8736]_ ,
    \new_[8737]_ , \new_[8738]_ , \new_[8739]_ , \new_[8740]_ ,
    \new_[8741]_ , \new_[8742]_ , \new_[8743]_ , \new_[8744]_ ,
    \new_[8745]_ , \new_[8746]_ , \new_[8747]_ , \new_[8748]_ ,
    \new_[8749]_ , \new_[8750]_ , \new_[8751]_ , \new_[8752]_ ,
    \new_[8753]_ , \new_[8754]_ , \new_[8755]_ , \new_[8756]_ ,
    \new_[8757]_ , \new_[8758]_ , \new_[8759]_ , \new_[8760]_ ,
    \new_[8761]_ , \new_[8762]_ , \new_[8763]_ , \new_[8764]_ ,
    \new_[8765]_ , \new_[8766]_ , \new_[8767]_ , \new_[8768]_ ,
    \new_[8769]_ , \new_[8770]_ , \new_[8771]_ , \new_[8772]_ ,
    \new_[8773]_ , \new_[8774]_ , \new_[8775]_ , \new_[8776]_ ,
    \new_[8777]_ , \new_[8778]_ , \new_[8779]_ , \new_[8780]_ ,
    \new_[8781]_ , \new_[8782]_ , \new_[8783]_ , \new_[8784]_ ,
    \new_[8785]_ , \new_[8786]_ , \new_[8787]_ , \new_[8788]_ ,
    \new_[8789]_ , \new_[8790]_ , \new_[8791]_ , \new_[8792]_ ,
    \new_[8793]_ , \new_[8794]_ , \new_[8795]_ , \new_[8796]_ ,
    \new_[8797]_ , \new_[8798]_ , \new_[8799]_ , \new_[8800]_ ,
    \new_[8801]_ , \new_[8802]_ , \new_[8803]_ , \new_[8804]_ ,
    \new_[8805]_ , \new_[8806]_ , \new_[8807]_ , \new_[8808]_ ,
    \new_[8809]_ , \new_[8810]_ , \new_[8811]_ , \new_[8812]_ ,
    \new_[8813]_ , \new_[8814]_ , \new_[8815]_ , \new_[8816]_ ,
    \new_[8817]_ , \new_[8818]_ , \new_[8819]_ , \new_[8820]_ ,
    \new_[8821]_ , \new_[8822]_ , \new_[8823]_ , \new_[8824]_ ,
    \new_[8825]_ , \new_[8826]_ , \new_[8827]_ , \new_[8828]_ ,
    \new_[8829]_ , \new_[8830]_ , \new_[8831]_ , \new_[8832]_ ,
    \new_[8833]_ , \new_[8834]_ , \new_[8835]_ , \new_[8836]_ ,
    \new_[8837]_ , \new_[8838]_ , \new_[8839]_ , \new_[8840]_ ,
    \new_[8841]_ , \new_[8842]_ , \new_[8843]_ , \new_[8844]_ ,
    \new_[8845]_ , \new_[8846]_ , \new_[8847]_ , \new_[8848]_ ,
    \new_[8849]_ , \new_[8850]_ , \new_[8851]_ , \new_[8852]_ ,
    \new_[8853]_ , \new_[8854]_ , \new_[8855]_ , \new_[8856]_ ,
    \new_[8857]_ , \new_[8858]_ , \new_[8859]_ , \new_[8860]_ ,
    \new_[8861]_ , \new_[8862]_ , \new_[8863]_ , \new_[8864]_ ,
    \new_[8865]_ , \new_[8866]_ , \new_[8867]_ , \new_[8868]_ ,
    \new_[8869]_ , \new_[8870]_ , \new_[8871]_ , \new_[8872]_ ,
    \new_[8873]_ , \new_[8874]_ , \new_[8875]_ , \new_[8876]_ ,
    \new_[8877]_ , \new_[8878]_ , \new_[8879]_ , \new_[8880]_ ,
    \new_[8881]_ , \new_[8882]_ , \new_[8883]_ , \new_[8884]_ ,
    \new_[8885]_ , \new_[8886]_ , \new_[8887]_ , \new_[8888]_ ,
    \new_[8889]_ , \new_[8890]_ , \new_[8891]_ , \new_[8892]_ ,
    \new_[8893]_ , \new_[8894]_ , \new_[8895]_ , \new_[8896]_ ,
    \new_[8897]_ , \new_[8898]_ , \new_[8899]_ , \new_[8900]_ ,
    \new_[8901]_ , \new_[8902]_ , \new_[8903]_ , \new_[8904]_ ,
    \new_[8905]_ , \new_[8906]_ , \new_[8907]_ , \new_[8908]_ ,
    \new_[8909]_ , \new_[8910]_ , \new_[8911]_ , \new_[8912]_ ,
    \new_[8913]_ , \new_[8914]_ , \new_[8915]_ , \new_[8916]_ ,
    \new_[8917]_ , \new_[8918]_ , \new_[8919]_ , \new_[8920]_ ,
    \new_[8921]_ , \new_[8922]_ , \new_[8923]_ , \new_[8924]_ ,
    \new_[8925]_ , \new_[8926]_ , \new_[8927]_ , \new_[8928]_ ,
    \new_[8929]_ , \new_[8930]_ , \new_[8931]_ , \new_[8932]_ ,
    \new_[8933]_ , \new_[8934]_ , \new_[8935]_ , \new_[8936]_ ,
    \new_[8937]_ , \new_[8938]_ , \new_[8939]_ , \new_[8940]_ ,
    \new_[8941]_ , \new_[8942]_ , \new_[8943]_ , \new_[8944]_ ,
    \new_[8945]_ , \new_[8946]_ , \new_[8947]_ , \new_[8948]_ ,
    \new_[8949]_ , \new_[8950]_ , \new_[8951]_ , \new_[8952]_ ,
    \new_[8953]_ , \new_[8954]_ , \new_[8955]_ , \new_[8956]_ ,
    \new_[8957]_ , \new_[8958]_ , \new_[8959]_ , \new_[8960]_ ,
    \new_[8961]_ , \new_[8962]_ , \new_[8963]_ , \new_[8964]_ ,
    \new_[8965]_ , \new_[8966]_ , \new_[8967]_ , \new_[8968]_ ,
    \new_[8969]_ , \new_[8970]_ , \new_[8971]_ , \new_[8972]_ ,
    \new_[8973]_ , \new_[8974]_ , \new_[8975]_ , \new_[8976]_ ,
    \new_[8977]_ , \new_[8978]_ , \new_[8979]_ , \new_[8980]_ ,
    \new_[8981]_ , \new_[8982]_ , \new_[8983]_ , \new_[8984]_ ,
    \new_[8985]_ , \new_[8986]_ , \new_[8987]_ , \new_[8988]_ ,
    \new_[8989]_ , \new_[8990]_ , \new_[8991]_ , \new_[8992]_ ,
    \new_[8993]_ , \new_[8994]_ , \new_[8995]_ , \new_[8996]_ ,
    \new_[8997]_ , \new_[8998]_ , \new_[8999]_ , \new_[9000]_ ,
    \new_[9001]_ , \new_[9002]_ , \new_[9003]_ , \new_[9004]_ ,
    \new_[9005]_ , \new_[9006]_ , \new_[9007]_ , \new_[9008]_ ,
    \new_[9009]_ , \new_[9010]_ , \new_[9011]_ , \new_[9012]_ ,
    \new_[9013]_ , \new_[9014]_ , \new_[9015]_ , \new_[9016]_ ,
    \new_[9017]_ , \new_[9018]_ , \new_[9019]_ , \new_[9020]_ ,
    \new_[9021]_ , \new_[9022]_ , \new_[9023]_ , \new_[9024]_ ,
    \new_[9025]_ , \new_[9026]_ , \new_[9027]_ , \new_[9028]_ ,
    \new_[9029]_ , \new_[9030]_ , \new_[9031]_ , \new_[9032]_ ,
    \new_[9033]_ , \new_[9034]_ , \new_[9035]_ , \new_[9036]_ ,
    \new_[9037]_ , \new_[9038]_ , \new_[9039]_ , \new_[9040]_ ,
    \new_[9041]_ , \new_[9042]_ , \new_[9043]_ , \new_[9044]_ ,
    \new_[9045]_ , \new_[9046]_ , \new_[9047]_ , \new_[9048]_ ,
    \new_[9049]_ , \new_[9050]_ , \new_[9051]_ , \new_[9052]_ ,
    \new_[9053]_ , \new_[9054]_ , \new_[9055]_ , \new_[9056]_ ,
    \new_[9057]_ , \new_[9058]_ , \new_[9059]_ , \new_[9060]_ ,
    \new_[9061]_ , \new_[9062]_ , \new_[9063]_ , \new_[9064]_ ,
    \new_[9065]_ , \new_[9066]_ , \new_[9067]_ , \new_[9068]_ ,
    \new_[9069]_ , \new_[9070]_ , \new_[9071]_ , \new_[9072]_ ,
    \new_[9073]_ , \new_[9074]_ , \new_[9075]_ , \new_[9076]_ ,
    \new_[9077]_ , \new_[9078]_ , \new_[9079]_ , \new_[9080]_ ,
    \new_[9081]_ , \new_[9082]_ , \new_[9083]_ , \new_[9084]_ ,
    \new_[9085]_ , \new_[9086]_ , \new_[9087]_ , \new_[9088]_ ,
    \new_[9089]_ , \new_[9090]_ , \new_[9091]_ , \new_[9092]_ ,
    \new_[9093]_ , \new_[9094]_ , \new_[9095]_ , \new_[9096]_ ,
    \new_[9097]_ , \new_[9098]_ , \new_[9099]_ , \new_[9100]_ ,
    \new_[9101]_ , \new_[9102]_ , \new_[9103]_ , \new_[9104]_ ,
    \new_[9105]_ , \new_[9106]_ , \new_[9107]_ , \new_[9108]_ ,
    \new_[9109]_ , \new_[9110]_ , \new_[9111]_ , \new_[9112]_ ,
    \new_[9113]_ , \new_[9114]_ , \new_[9115]_ , \new_[9116]_ ,
    \new_[9117]_ , \new_[9118]_ , \new_[9119]_ , \new_[9120]_ ,
    \new_[9121]_ , \new_[9122]_ , \new_[9123]_ , \new_[9124]_ ,
    \new_[9125]_ , \new_[9126]_ , \new_[9127]_ , \new_[9128]_ ,
    \new_[9129]_ , \new_[9130]_ , \new_[9131]_ , \new_[9132]_ ,
    \new_[9133]_ , \new_[9134]_ , \new_[9135]_ , \new_[9136]_ ,
    \new_[9137]_ , \new_[9138]_ , \new_[9139]_ , \new_[9140]_ ,
    \new_[9141]_ , \new_[9142]_ , \new_[9143]_ , \new_[9144]_ ,
    \new_[9145]_ , \new_[9146]_ , \new_[9147]_ , \new_[9148]_ ,
    \new_[9149]_ , \new_[9150]_ , \new_[9151]_ , \new_[9152]_ ,
    \new_[9153]_ , \new_[9154]_ , \new_[9155]_ , \new_[9156]_ ,
    \new_[9157]_ , \new_[9158]_ , \new_[9159]_ , \new_[9160]_ ,
    \new_[9161]_ , \new_[9162]_ , \new_[9163]_ , \new_[9164]_ ,
    \new_[9165]_ , \new_[9166]_ , \new_[9167]_ , \new_[9168]_ ,
    \new_[9169]_ , \new_[9170]_ , \new_[9171]_ , \new_[9172]_ ,
    \new_[9173]_ , \new_[9174]_ , \new_[9175]_ , \new_[9176]_ ,
    \new_[9177]_ , \new_[9178]_ , \new_[9179]_ , \new_[9180]_ ,
    \new_[9181]_ , \new_[9182]_ , \new_[9183]_ , \new_[9184]_ ,
    \new_[9185]_ , \new_[9186]_ , \new_[9187]_ , \new_[9188]_ ,
    \new_[9189]_ , \new_[9190]_ , \new_[9191]_ , \new_[9192]_ ,
    \new_[9193]_ , \new_[9194]_ , \new_[9195]_ , \new_[9196]_ ,
    \new_[9197]_ , \new_[9198]_ , \new_[9199]_ , \new_[9200]_ ,
    \new_[9201]_ , \new_[9202]_ , \new_[9203]_ , \new_[9204]_ ,
    \new_[9205]_ , \new_[9206]_ , \new_[9207]_ , \new_[9208]_ ,
    \new_[9209]_ , \new_[9210]_ , \new_[9211]_ , \new_[9212]_ ,
    \new_[9213]_ , \new_[9214]_ , \new_[9215]_ , \new_[9216]_ ,
    \new_[9217]_ , \new_[9218]_ , \new_[9219]_ , \new_[9220]_ ,
    \new_[9221]_ , \new_[9222]_ , \new_[9223]_ , \new_[9224]_ ,
    \new_[9225]_ , \new_[9226]_ , \new_[9227]_ , \new_[9228]_ ,
    \new_[9229]_ , \new_[9230]_ , \new_[9231]_ , \new_[9232]_ ,
    \new_[9233]_ , \new_[9234]_ , \new_[9235]_ , \new_[9236]_ ,
    \new_[9237]_ , \new_[9238]_ , \new_[9239]_ , \new_[9240]_ ,
    \new_[9241]_ , \new_[9242]_ , \new_[9243]_ , \new_[9244]_ ,
    \new_[9245]_ , \new_[9246]_ , \new_[9247]_ , \new_[9248]_ ,
    \new_[9249]_ , \new_[9250]_ , \new_[9251]_ , \new_[9252]_ ,
    \new_[9253]_ , \new_[9254]_ , \new_[9255]_ , \new_[9256]_ ,
    \new_[9257]_ , \new_[9258]_ , \new_[9259]_ , \new_[9260]_ ,
    \new_[9261]_ , \new_[9262]_ , \new_[9263]_ , \new_[9264]_ ,
    \new_[9265]_ , \new_[9266]_ , \new_[9267]_ , \new_[9268]_ ,
    \new_[9269]_ , \new_[9270]_ , \new_[9271]_ , \new_[9272]_ ,
    \new_[9273]_ , \new_[9274]_ , \new_[9275]_ , \new_[9276]_ ,
    \new_[9277]_ , \new_[9278]_ , \new_[9279]_ , \new_[9280]_ ,
    \new_[9281]_ , \new_[9282]_ , \new_[9283]_ , \new_[9284]_ ,
    \new_[9285]_ , \new_[9286]_ , \new_[9287]_ , \new_[9288]_ ,
    \new_[9289]_ , \new_[9290]_ , \new_[9291]_ , \new_[9292]_ ,
    \new_[9293]_ , \new_[9294]_ , \new_[9295]_ , \new_[9296]_ ,
    \new_[9297]_ , \new_[9298]_ , \new_[9299]_ , \new_[9300]_ ,
    \new_[9301]_ , \new_[9302]_ , \new_[9303]_ , \new_[9304]_ ,
    \new_[9305]_ , \new_[9306]_ , \new_[9307]_ , \new_[9308]_ ,
    \new_[9309]_ , \new_[9310]_ , \new_[9311]_ , \new_[9312]_ ,
    \new_[9313]_ , \new_[9314]_ , \new_[9315]_ , \new_[9316]_ ,
    \new_[9317]_ , \new_[9318]_ , \new_[9319]_ , \new_[9320]_ ,
    \new_[9321]_ , \new_[9322]_ , \new_[9323]_ , \new_[9324]_ ,
    \new_[9325]_ , \new_[9326]_ , \new_[9327]_ , \new_[9328]_ ,
    \new_[9329]_ , \new_[9330]_ , \new_[9331]_ , \new_[9332]_ ,
    \new_[9333]_ , \new_[9334]_ , \new_[9335]_ , \new_[9336]_ ,
    \new_[9337]_ , \new_[9338]_ , \new_[9339]_ , \new_[9340]_ ,
    \new_[9341]_ , \new_[9342]_ , \new_[9343]_ , \new_[9344]_ ,
    \new_[9345]_ , \new_[9346]_ , \new_[9347]_ , \new_[9348]_ ,
    \new_[9349]_ , \new_[9350]_ , \new_[9351]_ , \new_[9352]_ ,
    \new_[9353]_ , \new_[9354]_ , \new_[9355]_ , \new_[9356]_ ,
    \new_[9357]_ , \new_[9358]_ , \new_[9359]_ , \new_[9360]_ ,
    \new_[9361]_ , \new_[9362]_ , \new_[9363]_ , \new_[9364]_ ,
    \new_[9365]_ , \new_[9366]_ , \new_[9367]_ , \new_[9368]_ ,
    \new_[9369]_ , \new_[9371]_ , \new_[9372]_ , \new_[9373]_ ,
    \new_[9374]_ , \new_[9375]_ , \new_[9376]_ , \new_[9377]_ ,
    \new_[9378]_ , \new_[9379]_ , \new_[9380]_ , \new_[9381]_ ,
    \new_[9382]_ , \new_[9383]_ , \new_[9384]_ , \new_[9385]_ ,
    \new_[9386]_ , \new_[9387]_ , \new_[9388]_ , \new_[9389]_ ,
    \new_[9390]_ , \new_[9391]_ , \new_[9392]_ , \new_[9393]_ ,
    \new_[9394]_ , \new_[9395]_ , \new_[9396]_ , \new_[9397]_ ,
    \new_[9398]_ , \new_[9399]_ , \new_[9400]_ , \new_[9401]_ ,
    \new_[9402]_ , \new_[9403]_ , \new_[9404]_ , \new_[9405]_ ,
    \new_[9406]_ , \new_[9407]_ , \new_[9408]_ , \new_[9409]_ ,
    \new_[9410]_ , \new_[9411]_ , \new_[9412]_ , \new_[9413]_ ,
    \new_[9414]_ , \new_[9415]_ , \new_[9416]_ , \new_[9417]_ ,
    \new_[9418]_ , \new_[9419]_ , \new_[9420]_ , \new_[9421]_ ,
    \new_[9422]_ , \new_[9423]_ , \new_[9424]_ , \new_[9425]_ ,
    \new_[9426]_ , \new_[9427]_ , \new_[9428]_ , \new_[9429]_ ,
    \new_[9430]_ , \new_[9431]_ , \new_[9432]_ , \new_[9433]_ ,
    \new_[9434]_ , \new_[9435]_ , \new_[9436]_ , \new_[9437]_ ,
    \new_[9438]_ , \new_[9439]_ , \new_[9440]_ , \new_[9441]_ ,
    \new_[9442]_ , \new_[9443]_ , \new_[9444]_ , \new_[9445]_ ,
    \new_[9446]_ , \new_[9447]_ , \new_[9448]_ , \new_[9449]_ ,
    \new_[9450]_ , \new_[9451]_ , \new_[9452]_ , \new_[9453]_ ,
    \new_[9454]_ , \new_[9455]_ , \new_[9456]_ , \new_[9457]_ ,
    \new_[9458]_ , \new_[9459]_ , \new_[9460]_ , \new_[9461]_ ,
    \new_[9462]_ , \new_[9463]_ , \new_[9464]_ , \new_[9465]_ ,
    \new_[9466]_ , \new_[9467]_ , \new_[9468]_ , \new_[9469]_ ,
    \new_[9470]_ , \new_[9471]_ , \new_[9472]_ , \new_[9473]_ ,
    \new_[9474]_ , \new_[9475]_ , \new_[9476]_ , \new_[9477]_ ,
    \new_[9478]_ , \new_[9479]_ , \new_[9480]_ , \new_[9481]_ ,
    \new_[9482]_ , \new_[9483]_ , \new_[9484]_ , \new_[9485]_ ,
    \new_[9486]_ , \new_[9487]_ , \new_[9488]_ , \new_[9489]_ ,
    \new_[9490]_ , \new_[9491]_ , \new_[9492]_ , \new_[9493]_ ,
    \new_[9494]_ , \new_[9495]_ , \new_[9496]_ , \new_[9497]_ ,
    \new_[9498]_ , \new_[9499]_ , \new_[9500]_ , \new_[9501]_ ,
    \new_[9502]_ , \new_[9503]_ , \new_[9504]_ , \new_[9505]_ ,
    \new_[9506]_ , \new_[9507]_ , \new_[9508]_ , \new_[9509]_ ,
    \new_[9510]_ , \new_[9511]_ , \new_[9512]_ , \new_[9513]_ ,
    \new_[9514]_ , \new_[9515]_ , \new_[9516]_ , \new_[9517]_ ,
    \new_[9518]_ , \new_[9519]_ , \new_[9520]_ , \new_[9521]_ ,
    \new_[9522]_ , \new_[9523]_ , \new_[9524]_ , \new_[9525]_ ,
    \new_[9526]_ , \new_[9527]_ , \new_[9528]_ , \new_[9529]_ ,
    \new_[9530]_ , \new_[9531]_ , \new_[9532]_ , \new_[9533]_ ,
    \new_[9534]_ , \new_[9535]_ , \new_[9536]_ , \new_[9537]_ ,
    \new_[9538]_ , \new_[9539]_ , \new_[9540]_ , \new_[9541]_ ,
    \new_[9542]_ , \new_[9543]_ , \new_[9544]_ , \new_[9545]_ ,
    \new_[9546]_ , \new_[9547]_ , \new_[9548]_ , \new_[9549]_ ,
    \new_[9550]_ , \new_[9551]_ , \new_[9552]_ , \new_[9553]_ ,
    \new_[9554]_ , \new_[9555]_ , \new_[9556]_ , \new_[9557]_ ,
    \new_[9558]_ , \new_[9559]_ , \new_[9560]_ , \new_[9561]_ ,
    \new_[9562]_ , \new_[9563]_ , \new_[9564]_ , \new_[9565]_ ,
    \new_[9566]_ , \new_[9567]_ , \new_[9568]_ , \new_[9569]_ ,
    \new_[9570]_ , \new_[9571]_ , \new_[9572]_ , \new_[9573]_ ,
    \new_[9574]_ , \new_[9575]_ , \new_[9576]_ , \new_[9577]_ ,
    \new_[9578]_ , \new_[9579]_ , \new_[9580]_ , \new_[9581]_ ,
    \new_[9582]_ , \new_[9583]_ , \new_[9584]_ , \new_[9585]_ ,
    \new_[9586]_ , \new_[9587]_ , \new_[9588]_ , \new_[9589]_ ,
    \new_[9590]_ , \new_[9591]_ , \new_[9592]_ , \new_[9593]_ ,
    \new_[9594]_ , \new_[9595]_ , \new_[9596]_ , \new_[9597]_ ,
    \new_[9598]_ , \new_[9599]_ , \new_[9600]_ , \new_[9601]_ ,
    \new_[9602]_ , \new_[9603]_ , \new_[9604]_ , \new_[9605]_ ,
    \new_[9606]_ , \new_[9607]_ , \new_[9608]_ , \new_[9609]_ ,
    \new_[9610]_ , \new_[9611]_ , \new_[9612]_ , \new_[9613]_ ,
    \new_[9614]_ , \new_[9615]_ , \new_[9616]_ , \new_[9617]_ ,
    \new_[9618]_ , \new_[9619]_ , \new_[9620]_ , \new_[9621]_ ,
    \new_[9622]_ , \new_[9623]_ , \new_[9624]_ , \new_[9625]_ ,
    \new_[9626]_ , \new_[9627]_ , \new_[9628]_ , \new_[9629]_ ,
    \new_[9630]_ , \new_[9631]_ , \new_[9632]_ , \new_[9633]_ ,
    \new_[9634]_ , \new_[9635]_ , \new_[9636]_ , \new_[9637]_ ,
    \new_[9638]_ , \new_[9639]_ , \new_[9640]_ , \new_[9641]_ ,
    \new_[9642]_ , \new_[9643]_ , \new_[9644]_ , \new_[9645]_ ,
    \new_[9646]_ , \new_[9647]_ , \new_[9648]_ , \new_[9649]_ ,
    \new_[9650]_ , \new_[9651]_ , \new_[9652]_ , \new_[9653]_ ,
    \new_[9654]_ , \new_[9655]_ , \new_[9656]_ , \new_[9657]_ ,
    \new_[9658]_ , \new_[9659]_ , \new_[9660]_ , \new_[9661]_ ,
    \new_[9662]_ , \new_[9663]_ , \new_[9664]_ , \new_[9665]_ ,
    \new_[9666]_ , \new_[9667]_ , \new_[9668]_ , \new_[9669]_ ,
    \new_[9670]_ , \new_[9671]_ , \new_[9672]_ , \new_[9673]_ ,
    \new_[9674]_ , \new_[9675]_ , \new_[9676]_ , \new_[9677]_ ,
    \new_[9678]_ , \new_[9679]_ , \new_[9680]_ , \new_[9681]_ ,
    \new_[9682]_ , \new_[9683]_ , \new_[9684]_ , \new_[9685]_ ,
    \new_[9686]_ , \new_[9687]_ , \new_[9688]_ , \new_[9689]_ ,
    \new_[9690]_ , \new_[9691]_ , \new_[9692]_ , \new_[9693]_ ,
    \new_[9694]_ , \new_[9695]_ , \new_[9696]_ , \new_[9697]_ ,
    \new_[9698]_ , \new_[9699]_ , \new_[9700]_ , \new_[9701]_ ,
    \new_[9702]_ , \new_[9703]_ , \new_[9704]_ , \new_[9705]_ ,
    \new_[9706]_ , \new_[9707]_ , \new_[9708]_ , \new_[9709]_ ,
    \new_[9710]_ , \new_[9711]_ , \new_[9712]_ , \new_[9713]_ ,
    \new_[9714]_ , \new_[9715]_ , \new_[9716]_ , \new_[9717]_ ,
    \new_[9718]_ , \new_[9719]_ , \new_[9720]_ , \new_[9721]_ ,
    \new_[9722]_ , \new_[9723]_ , \new_[9724]_ , \new_[9725]_ ,
    \new_[9726]_ , \new_[9727]_ , \new_[9728]_ , \new_[9729]_ ,
    \new_[9730]_ , \new_[9731]_ , \new_[9732]_ , \new_[9733]_ ,
    \new_[9734]_ , \new_[9735]_ , \new_[9736]_ , \new_[9737]_ ,
    \new_[9738]_ , \new_[9739]_ , \new_[9740]_ , \new_[9741]_ ,
    \new_[9742]_ , \new_[9743]_ , \new_[9744]_ , \new_[9745]_ ,
    \new_[9746]_ , \new_[9747]_ , \new_[9748]_ , \new_[9749]_ ,
    \new_[9750]_ , \new_[9751]_ , \new_[9752]_ , \new_[9753]_ ,
    \new_[9754]_ , \new_[9755]_ , \new_[9756]_ , \new_[9757]_ ,
    \new_[9758]_ , \new_[9759]_ , \new_[9760]_ , \new_[9761]_ ,
    \new_[9762]_ , \new_[9763]_ , \new_[9764]_ , \new_[9765]_ ,
    \new_[9766]_ , \new_[9767]_ , \new_[9768]_ , \new_[9769]_ ,
    \new_[9770]_ , \new_[9771]_ , \new_[9772]_ , \new_[9773]_ ,
    \new_[9774]_ , \new_[9775]_ , \new_[9776]_ , \new_[9777]_ ,
    \new_[9778]_ , \new_[9779]_ , \new_[9780]_ , \new_[9781]_ ,
    \new_[9782]_ , \new_[9783]_ , \new_[9784]_ , \new_[9785]_ ,
    \new_[9786]_ , \new_[9787]_ , \new_[9788]_ , \new_[9789]_ ,
    \new_[9790]_ , \new_[9791]_ , \new_[9792]_ , \new_[9793]_ ,
    \new_[9794]_ , \new_[9795]_ , \new_[9796]_ , \new_[9797]_ ,
    \new_[9798]_ , \new_[9799]_ , \new_[9800]_ , \new_[9801]_ ,
    \new_[9802]_ , \new_[9803]_ , \new_[9804]_ , \new_[9805]_ ,
    \new_[9806]_ , \new_[9807]_ , \new_[9808]_ , \new_[9809]_ ,
    \new_[9810]_ , \new_[9811]_ , \new_[9812]_ , \new_[9813]_ ,
    \new_[9814]_ , \new_[9815]_ , \new_[9816]_ , \new_[9817]_ ,
    \new_[9818]_ , \new_[9819]_ , \new_[9820]_ , \new_[9821]_ ,
    \new_[9822]_ , \new_[9823]_ , \new_[9824]_ , \new_[9825]_ ,
    \new_[9826]_ , \new_[9827]_ , \new_[9828]_ , \new_[9829]_ ,
    \new_[9830]_ , \new_[9831]_ , \new_[9832]_ , \new_[9833]_ ,
    \new_[9834]_ , \new_[9835]_ , \new_[9836]_ , \new_[9837]_ ,
    \new_[9838]_ , \new_[9839]_ , \new_[9840]_ , \new_[9841]_ ,
    \new_[9842]_ , \new_[9843]_ , \new_[9844]_ , \new_[9845]_ ,
    \new_[9846]_ , \new_[9847]_ , \new_[9848]_ , \new_[9849]_ ,
    \new_[9850]_ , \new_[9851]_ , \new_[9852]_ , \new_[9853]_ ,
    \new_[9854]_ , \new_[9855]_ , \new_[9856]_ , \new_[9857]_ ,
    \new_[9858]_ , \new_[9859]_ , \new_[9860]_ , \new_[9861]_ ,
    \new_[9862]_ , \new_[9863]_ , \new_[9864]_ , \new_[9865]_ ,
    \new_[9866]_ , \new_[9867]_ , \new_[9868]_ , \new_[9869]_ ,
    \new_[9870]_ , \new_[9871]_ , \new_[9872]_ , \new_[9873]_ ,
    \new_[9874]_ , \new_[9875]_ , \new_[9876]_ , \new_[9877]_ ,
    \new_[9878]_ , \new_[9879]_ , \new_[9880]_ , \new_[9881]_ ,
    \new_[9882]_ , \new_[9883]_ , \new_[9884]_ , \new_[9885]_ ,
    \new_[9886]_ , \new_[9887]_ , \new_[9888]_ , \new_[9889]_ ,
    \new_[9890]_ , \new_[9891]_ , \new_[9892]_ , \new_[9893]_ ,
    \new_[9894]_ , \new_[9895]_ , \new_[9896]_ , \new_[9897]_ ,
    \new_[9898]_ , \new_[9899]_ , \new_[9900]_ , \new_[9901]_ ,
    \new_[9902]_ , \new_[9903]_ , \new_[9904]_ , \new_[9905]_ ,
    \new_[9906]_ , \new_[9907]_ , \new_[9908]_ , \new_[9909]_ ,
    \new_[9910]_ , \new_[9911]_ , \new_[9912]_ , \new_[9913]_ ,
    \new_[9914]_ , \new_[9915]_ , \new_[9916]_ , \new_[9917]_ ,
    \new_[9918]_ , \new_[9919]_ , \new_[9920]_ , \new_[9921]_ ,
    \new_[9922]_ , \new_[9923]_ , \new_[9924]_ , \new_[9925]_ ,
    \new_[9926]_ , \new_[9927]_ , \new_[9928]_ , \new_[9929]_ ,
    \new_[9930]_ , \new_[9931]_ , \new_[9932]_ , \new_[9933]_ ,
    \new_[9934]_ , \new_[9935]_ , \new_[9936]_ , \new_[9937]_ ,
    \new_[9938]_ , \new_[9939]_ , \new_[9940]_ , \new_[9941]_ ,
    \new_[9942]_ , \new_[9943]_ , \new_[9944]_ , \new_[9945]_ ,
    \new_[9946]_ , \new_[9947]_ , \new_[9948]_ , \new_[9949]_ ,
    \new_[9950]_ , \new_[9951]_ , \new_[9952]_ , \new_[9953]_ ,
    \new_[9954]_ , \new_[9955]_ , \new_[9956]_ , \new_[9957]_ ,
    \new_[9958]_ , \new_[9959]_ , \new_[9960]_ , \new_[9961]_ ,
    \new_[9962]_ , \new_[9963]_ , \new_[9964]_ , \new_[9965]_ ,
    \new_[9966]_ , \new_[9967]_ , \new_[9968]_ , \new_[9969]_ ,
    \new_[9970]_ , \new_[9971]_ , \new_[9972]_ , \new_[9973]_ ,
    \new_[9974]_ , \new_[9975]_ , \new_[9976]_ , \new_[9977]_ ,
    \new_[9978]_ , \new_[9979]_ , \new_[9980]_ , \new_[9981]_ ,
    \new_[9982]_ , \new_[9983]_ , \new_[9984]_ , \new_[9985]_ ,
    \new_[9986]_ , \new_[9987]_ , \new_[9988]_ , \new_[9989]_ ,
    \new_[9990]_ , \new_[9991]_ , \new_[9992]_ , \new_[9993]_ ,
    \new_[9994]_ , \new_[9995]_ , \new_[9996]_ , \new_[9997]_ ,
    \new_[9998]_ , \new_[9999]_ , \new_[10000]_ , \new_[10001]_ ,
    \new_[10002]_ , \new_[10003]_ , \new_[10004]_ , \new_[10005]_ ,
    \new_[10006]_ , \new_[10007]_ , \new_[10008]_ , \new_[10009]_ ,
    \new_[10010]_ , \new_[10011]_ , \new_[10012]_ , \new_[10013]_ ,
    \new_[10014]_ , \new_[10015]_ , \new_[10016]_ , \new_[10017]_ ,
    \new_[10018]_ , \new_[10019]_ , \new_[10020]_ , \new_[10021]_ ,
    \new_[10022]_ , \new_[10023]_ , \new_[10024]_ , \new_[10025]_ ,
    \new_[10026]_ , \new_[10027]_ , \new_[10028]_ , \new_[10029]_ ,
    \new_[10030]_ , \new_[10031]_ , \new_[10032]_ , \new_[10033]_ ,
    \new_[10034]_ , \new_[10035]_ , \new_[10036]_ , \new_[10037]_ ,
    \new_[10038]_ , \new_[10039]_ , \new_[10040]_ , \new_[10041]_ ,
    \new_[10042]_ , \new_[10043]_ , \new_[10044]_ , \new_[10045]_ ,
    \new_[10046]_ , \new_[10047]_ , \new_[10048]_ , \new_[10049]_ ,
    \new_[10050]_ , \new_[10051]_ , \new_[10052]_ , \new_[10053]_ ,
    \new_[10054]_ , \new_[10055]_ , \new_[10056]_ , \new_[10057]_ ,
    \new_[10058]_ , \new_[10059]_ , \new_[10060]_ , \new_[10061]_ ,
    \new_[10062]_ , \new_[10063]_ , \new_[10064]_ , \new_[10065]_ ,
    \new_[10066]_ , \new_[10067]_ , \new_[10068]_ , \new_[10069]_ ,
    \new_[10070]_ , \new_[10071]_ , \new_[10072]_ , \new_[10073]_ ,
    \new_[10074]_ , \new_[10075]_ , \new_[10076]_ , \new_[10077]_ ,
    \new_[10078]_ , \new_[10079]_ , \new_[10080]_ , \new_[10081]_ ,
    \new_[10082]_ , \new_[10083]_ , \new_[10084]_ , \new_[10085]_ ,
    \new_[10086]_ , \new_[10087]_ , \new_[10088]_ , \new_[10089]_ ,
    \new_[10090]_ , \new_[10091]_ , \new_[10092]_ , \new_[10093]_ ,
    \new_[10094]_ , \new_[10095]_ , \new_[10096]_ , \new_[10097]_ ,
    \new_[10098]_ , \new_[10099]_ , \new_[10100]_ , \new_[10101]_ ,
    \new_[10102]_ , \new_[10103]_ , \new_[10104]_ , \new_[10105]_ ,
    \new_[10106]_ , \new_[10107]_ , \new_[10108]_ , \new_[10109]_ ,
    \new_[10110]_ , \new_[10111]_ , \new_[10112]_ , \new_[10113]_ ,
    \new_[10114]_ , \new_[10115]_ , \new_[10116]_ , \new_[10117]_ ,
    \new_[10118]_ , \new_[10119]_ , \new_[10120]_ , \new_[10121]_ ,
    \new_[10122]_ , \new_[10123]_ , \new_[10124]_ , \new_[10125]_ ,
    \new_[10126]_ , \new_[10127]_ , \new_[10128]_ , \new_[10129]_ ,
    \new_[10130]_ , \new_[10131]_ , \new_[10132]_ , \new_[10133]_ ,
    \new_[10134]_ , \new_[10135]_ , \new_[10136]_ , \new_[10137]_ ,
    \new_[10138]_ , \new_[10139]_ , \new_[10140]_ , \new_[10141]_ ,
    \new_[10142]_ , \new_[10143]_ , \new_[10144]_ , \new_[10145]_ ,
    \new_[10146]_ , \new_[10147]_ , \new_[10148]_ , \new_[10149]_ ,
    \new_[10150]_ , \new_[10151]_ , \new_[10152]_ , \new_[10153]_ ,
    \new_[10154]_ , \new_[10155]_ , \new_[10156]_ , \new_[10157]_ ,
    \new_[10158]_ , \new_[10159]_ , \new_[10160]_ , \new_[10161]_ ,
    \new_[10162]_ , \new_[10163]_ , \new_[10164]_ , \new_[10165]_ ,
    \new_[10166]_ , \new_[10167]_ , \new_[10168]_ , \new_[10169]_ ,
    \new_[10170]_ , \new_[10171]_ , \new_[10172]_ , \new_[10173]_ ,
    \new_[10174]_ , \new_[10175]_ , \new_[10176]_ , \new_[10177]_ ,
    \new_[10178]_ , \new_[10179]_ , \new_[10180]_ , \new_[10181]_ ,
    \new_[10182]_ , \new_[10183]_ , \new_[10184]_ , \new_[10185]_ ,
    \new_[10186]_ , \new_[10187]_ , \new_[10188]_ , \new_[10189]_ ,
    \new_[10190]_ , \new_[10191]_ , \new_[10192]_ , \new_[10193]_ ,
    \new_[10194]_ , \new_[10195]_ , \new_[10196]_ , \new_[10197]_ ,
    \new_[10198]_ , \new_[10199]_ , \new_[10200]_ , \new_[10201]_ ,
    \new_[10202]_ , \new_[10203]_ , \new_[10204]_ , \new_[10205]_ ,
    \new_[10206]_ , \new_[10207]_ , \new_[10208]_ , \new_[10209]_ ,
    \new_[10210]_ , \new_[10211]_ , \new_[10212]_ , \new_[10213]_ ,
    \new_[10214]_ , \new_[10215]_ , \new_[10216]_ , \new_[10217]_ ,
    \new_[10218]_ , \new_[10219]_ , \new_[10220]_ , \new_[10221]_ ,
    \new_[10222]_ , \new_[10223]_ , \new_[10224]_ , \new_[10225]_ ,
    \new_[10226]_ , \new_[10227]_ , \new_[10228]_ , \new_[10229]_ ,
    \new_[10230]_ , \new_[10231]_ , \new_[10232]_ , \new_[10233]_ ,
    \new_[10234]_ , \new_[10235]_ , \new_[10236]_ , \new_[10237]_ ,
    \new_[10238]_ , \new_[10239]_ , \new_[10240]_ , \new_[10241]_ ,
    \new_[10242]_ , \new_[10243]_ , \new_[10244]_ , \new_[10245]_ ,
    \new_[10246]_ , \new_[10247]_ , \new_[10248]_ , \new_[10249]_ ,
    \new_[10250]_ , \new_[10251]_ , \new_[10252]_ , \new_[10253]_ ,
    \new_[10254]_ , \new_[10255]_ , \new_[10256]_ , \new_[10257]_ ,
    \new_[10258]_ , \new_[10259]_ , \new_[10260]_ , \new_[10261]_ ,
    \new_[10262]_ , \new_[10263]_ , \new_[10264]_ , \new_[10265]_ ,
    \new_[10266]_ , \new_[10267]_ , \new_[10268]_ , \new_[10269]_ ,
    \new_[10270]_ , \new_[10271]_ , \new_[10272]_ , \new_[10273]_ ,
    \new_[10274]_ , \new_[10275]_ , \new_[10276]_ , \new_[10277]_ ,
    \new_[10278]_ , \new_[10279]_ , \new_[10280]_ , \new_[10281]_ ,
    \new_[10282]_ , \new_[10283]_ , \new_[10284]_ , \new_[10285]_ ,
    \new_[10286]_ , \new_[10287]_ , \new_[10288]_ , \new_[10289]_ ,
    \new_[10290]_ , \new_[10291]_ , \new_[10292]_ , \new_[10293]_ ,
    \new_[10294]_ , \new_[10295]_ , \new_[10296]_ , \new_[10297]_ ,
    \new_[10298]_ , \new_[10299]_ , \new_[10300]_ , \new_[10301]_ ,
    \new_[10302]_ , \new_[10303]_ , \new_[10304]_ , \new_[10305]_ ,
    \new_[10306]_ , \new_[10307]_ , \new_[10308]_ , \new_[10309]_ ,
    \new_[10310]_ , \new_[10311]_ , \new_[10312]_ , \new_[10313]_ ,
    \new_[10314]_ , \new_[10315]_ , \new_[10316]_ , \new_[10317]_ ,
    \new_[10318]_ , \new_[10319]_ , \new_[10320]_ , \new_[10321]_ ,
    \new_[10322]_ , \new_[10323]_ , \new_[10324]_ , \new_[10325]_ ,
    \new_[10326]_ , \new_[10327]_ , \new_[10328]_ , \new_[10329]_ ,
    \new_[10330]_ , \new_[10331]_ , \new_[10332]_ , \new_[10333]_ ,
    \new_[10334]_ , \new_[10335]_ , \new_[10336]_ , \new_[10337]_ ,
    \new_[10338]_ , \new_[10339]_ , \new_[10340]_ , \new_[10341]_ ,
    \new_[10342]_ , \new_[10343]_ , \new_[10344]_ , \new_[10345]_ ,
    \new_[10346]_ , \new_[10347]_ , \new_[10348]_ , \new_[10349]_ ,
    \new_[10350]_ , \new_[10351]_ , \new_[10352]_ , \new_[10353]_ ,
    \new_[10354]_ , \new_[10355]_ , \new_[10356]_ , \new_[10357]_ ,
    \new_[10358]_ , \new_[10359]_ , \new_[10360]_ , \new_[10361]_ ,
    \new_[10362]_ , \new_[10363]_ , \new_[10364]_ , \new_[10365]_ ,
    \new_[10366]_ , \new_[10367]_ , \new_[10368]_ , \new_[10369]_ ,
    \new_[10370]_ , \new_[10371]_ , \new_[10372]_ , \new_[10373]_ ,
    \new_[10374]_ , \new_[10375]_ , \new_[10376]_ , \new_[10377]_ ,
    \new_[10378]_ , \new_[10379]_ , \new_[10380]_ , \new_[10381]_ ,
    \new_[10382]_ , \new_[10383]_ , \new_[10384]_ , \new_[10385]_ ,
    \new_[10386]_ , \new_[10387]_ , \new_[10388]_ , \new_[10389]_ ,
    \new_[10390]_ , \new_[10391]_ , \new_[10392]_ , \new_[10393]_ ,
    \new_[10394]_ , \new_[10395]_ , \new_[10396]_ , \new_[10397]_ ,
    \new_[10398]_ , \new_[10399]_ , \new_[10400]_ , \new_[10401]_ ,
    \new_[10402]_ , \new_[10403]_ , \new_[10404]_ , \new_[10405]_ ,
    \new_[10406]_ , \new_[10407]_ , \new_[10408]_ , \new_[10409]_ ,
    \new_[10410]_ , \new_[10411]_ , \new_[10412]_ , \new_[10413]_ ,
    \new_[10414]_ , \new_[10415]_ , \new_[10416]_ , \new_[10417]_ ,
    \new_[10418]_ , \new_[10419]_ , \new_[10420]_ , \new_[10421]_ ,
    \new_[10422]_ , \new_[10423]_ , \new_[10424]_ , \new_[10425]_ ,
    \new_[10426]_ , \new_[10427]_ , \new_[10428]_ , \new_[10429]_ ,
    \new_[10430]_ , \new_[10431]_ , \new_[10432]_ , \new_[10433]_ ,
    \new_[10434]_ , \new_[10435]_ , \new_[10436]_ , \new_[10437]_ ,
    \new_[10438]_ , \new_[10439]_ , \new_[10440]_ , \new_[10441]_ ,
    \new_[10442]_ , \new_[10443]_ , \new_[10444]_ , \new_[10445]_ ,
    \new_[10446]_ , \new_[10447]_ , \new_[10448]_ , \new_[10449]_ ,
    \new_[10450]_ , \new_[10451]_ , \new_[10452]_ , \new_[10453]_ ,
    \new_[10454]_ , \new_[10455]_ , \new_[10456]_ , \new_[10457]_ ,
    \new_[10458]_ , \new_[10459]_ , \new_[10460]_ , \new_[10461]_ ,
    \new_[10462]_ , \new_[10463]_ , \new_[10464]_ , \new_[10465]_ ,
    \new_[10466]_ , \new_[10467]_ , \new_[10468]_ , \new_[10469]_ ,
    \new_[10470]_ , \new_[10471]_ , \new_[10472]_ , \new_[10473]_ ,
    \new_[10474]_ , \new_[10475]_ , \new_[10476]_ , \new_[10477]_ ,
    \new_[10478]_ , \new_[10479]_ , \new_[10480]_ , \new_[10481]_ ,
    \new_[10482]_ , \new_[10483]_ , \new_[10484]_ , \new_[10485]_ ,
    \new_[10486]_ , \new_[10487]_ , \new_[10488]_ , \new_[10489]_ ,
    \new_[10490]_ , \new_[10491]_ , \new_[10492]_ , \new_[10493]_ ,
    \new_[10494]_ , \new_[10495]_ , \new_[10496]_ , \new_[10497]_ ,
    \new_[10498]_ , \new_[10499]_ , \new_[10500]_ , \new_[10501]_ ,
    \new_[10502]_ , \new_[10503]_ , \new_[10504]_ , \new_[10505]_ ,
    \new_[10506]_ , \new_[10507]_ , \new_[10508]_ , \new_[10509]_ ,
    \new_[10510]_ , \new_[10511]_ , \new_[10512]_ , \new_[10513]_ ,
    \new_[10514]_ , \new_[10515]_ , \new_[10516]_ , \new_[10517]_ ,
    \new_[10518]_ , \new_[10519]_ , \new_[10520]_ , \new_[10521]_ ,
    \new_[10522]_ , \new_[10523]_ , \new_[10524]_ , \new_[10525]_ ,
    \new_[10526]_ , \new_[10527]_ , \new_[10528]_ , \new_[10529]_ ,
    \new_[10530]_ , \new_[10531]_ , \new_[10532]_ , \new_[10533]_ ,
    \new_[10534]_ , \new_[10535]_ , \new_[10536]_ , \new_[10537]_ ,
    \new_[10538]_ , \new_[10539]_ , \new_[10540]_ , \new_[10541]_ ,
    \new_[10542]_ , \new_[10543]_ , \new_[10544]_ , \new_[10545]_ ,
    \new_[10546]_ , \new_[10547]_ , \new_[10548]_ , \new_[10549]_ ,
    \new_[10550]_ , \new_[10551]_ , \new_[10552]_ , \new_[10553]_ ,
    \new_[10554]_ , \new_[10555]_ , \new_[10556]_ , \new_[10557]_ ,
    \new_[10558]_ , \new_[10559]_ , \new_[10560]_ , \new_[10561]_ ,
    \new_[10562]_ , \new_[10563]_ , \new_[10564]_ , \new_[10565]_ ,
    \new_[10566]_ , \new_[10567]_ , \new_[10568]_ , \new_[10569]_ ,
    \new_[10570]_ , \new_[10571]_ , \new_[10572]_ , \new_[10573]_ ,
    \new_[10574]_ , \new_[10575]_ , \new_[10576]_ , \new_[10577]_ ,
    \new_[10578]_ , \new_[10579]_ , \new_[10580]_ , \new_[10581]_ ,
    \new_[10582]_ , \new_[10583]_ , \new_[10584]_ , \new_[10585]_ ,
    \new_[10586]_ , \new_[10587]_ , \new_[10588]_ , \new_[10589]_ ,
    \new_[10590]_ , \new_[10591]_ , \new_[10592]_ , \new_[10593]_ ,
    \new_[10594]_ , \new_[10595]_ , \new_[10596]_ , \new_[10597]_ ,
    \new_[10598]_ , \new_[10599]_ , \new_[10600]_ , \new_[10601]_ ,
    \new_[10602]_ , \new_[10603]_ , \new_[10604]_ , \new_[10605]_ ,
    \new_[10606]_ , \new_[10607]_ , \new_[10608]_ , \new_[10609]_ ,
    \new_[10610]_ , \new_[10611]_ , \new_[10612]_ , \new_[10613]_ ,
    \new_[10614]_ , \new_[10615]_ , \new_[10616]_ , \new_[10617]_ ,
    \new_[10618]_ , \new_[10619]_ , \new_[10620]_ , \new_[10621]_ ,
    \new_[10622]_ , \new_[10623]_ , \new_[10624]_ , \new_[10625]_ ,
    \new_[10626]_ , \new_[10627]_ , \new_[10628]_ , \new_[10629]_ ,
    \new_[10630]_ , \new_[10631]_ , \new_[10632]_ , \new_[10633]_ ,
    \new_[10634]_ , \new_[10635]_ , \new_[10636]_ , \new_[10637]_ ,
    \new_[10638]_ , \new_[10639]_ , \new_[10640]_ , \new_[10641]_ ,
    \new_[10642]_ , \new_[10643]_ , \new_[10644]_ , \new_[10645]_ ,
    \new_[10646]_ , \new_[10647]_ , \new_[10648]_ , \new_[10649]_ ,
    \new_[10650]_ , \new_[10651]_ , \new_[10652]_ , \new_[10653]_ ,
    \new_[10654]_ , \new_[10655]_ , \new_[10656]_ , \new_[10657]_ ,
    \new_[10658]_ , \new_[10659]_ , \new_[10660]_ , \new_[10661]_ ,
    \new_[10662]_ , \new_[10663]_ , \new_[10664]_ , \new_[10665]_ ,
    \new_[10666]_ , \new_[10667]_ , \new_[10668]_ , \new_[10669]_ ,
    \new_[10670]_ , \new_[10671]_ , \new_[10672]_ , \new_[10673]_ ,
    \new_[10674]_ , \new_[10675]_ , \new_[10676]_ , \new_[10677]_ ,
    \new_[10678]_ , \new_[10679]_ , \new_[10680]_ , \new_[10681]_ ,
    \new_[10682]_ , \new_[10683]_ , \new_[10684]_ , \new_[10685]_ ,
    \new_[10686]_ , \new_[10687]_ , \new_[10688]_ , \new_[10689]_ ,
    \new_[10690]_ , \new_[10691]_ , \new_[10692]_ , \new_[10693]_ ,
    \new_[10694]_ , \new_[10695]_ , \new_[10696]_ , \new_[10697]_ ,
    \new_[10698]_ , \new_[10699]_ , \new_[10700]_ , \new_[10701]_ ,
    \new_[10702]_ , \new_[10703]_ , \new_[10704]_ , \new_[10705]_ ,
    \new_[10706]_ , \new_[10707]_ , \new_[10708]_ , \new_[10709]_ ,
    \new_[10710]_ , \new_[10711]_ , \new_[10712]_ , \new_[10713]_ ,
    \new_[10714]_ , \new_[10715]_ , \new_[10716]_ , \new_[10717]_ ,
    \new_[10718]_ , \new_[10719]_ , \new_[10720]_ , \new_[10721]_ ,
    \new_[10722]_ , \new_[10723]_ , \new_[10724]_ , \new_[10725]_ ,
    \new_[10726]_ , \new_[10727]_ , \new_[10728]_ , \new_[10729]_ ,
    \new_[10730]_ , \new_[10731]_ , \new_[10732]_ , \new_[10733]_ ,
    \new_[10734]_ , \new_[10735]_ , \new_[10736]_ , \new_[10737]_ ,
    \new_[10738]_ , \new_[10739]_ , \new_[10740]_ , \new_[10741]_ ,
    \new_[10742]_ , \new_[10743]_ , \new_[10744]_ , \new_[10745]_ ,
    \new_[10746]_ , \new_[10747]_ , \new_[10748]_ , \new_[10749]_ ,
    \new_[10750]_ , \new_[10751]_ , \new_[10752]_ , \new_[10753]_ ,
    \new_[10754]_ , \new_[10755]_ , \new_[10756]_ , \new_[10757]_ ,
    \new_[10758]_ , \new_[10759]_ , \new_[10760]_ , \new_[10761]_ ,
    \new_[10762]_ , \new_[10763]_ , \new_[10764]_ , \new_[10765]_ ,
    \new_[10766]_ , \new_[10767]_ , \new_[10768]_ , \new_[10769]_ ,
    \new_[10770]_ , \new_[10771]_ , \new_[10772]_ , \new_[10773]_ ,
    \new_[10774]_ , \new_[10775]_ , \new_[10776]_ , \new_[10777]_ ,
    \new_[10778]_ , \new_[10779]_ , \new_[10780]_ , \new_[10781]_ ,
    \new_[10782]_ , \new_[10783]_ , \new_[10784]_ , \new_[10785]_ ,
    \new_[10786]_ , \new_[10787]_ , \new_[10788]_ , \new_[10789]_ ,
    \new_[10790]_ , \new_[10791]_ , \new_[10792]_ , \new_[10793]_ ,
    \new_[10794]_ , \new_[10795]_ , \new_[10796]_ , \new_[10797]_ ,
    \new_[10798]_ , \new_[10799]_ , \new_[10800]_ , \new_[10801]_ ,
    \new_[10802]_ , \new_[10803]_ , \new_[10804]_ , \new_[10805]_ ,
    \new_[10806]_ , \new_[10807]_ , \new_[10808]_ , \new_[10809]_ ,
    \new_[10810]_ , \new_[10811]_ , \new_[10812]_ , \new_[10813]_ ,
    \new_[10814]_ , \new_[10815]_ , \new_[10816]_ , \new_[10817]_ ,
    \new_[10818]_ , \new_[10819]_ , \new_[10820]_ , \new_[10821]_ ,
    \new_[10822]_ , \new_[10823]_ , \new_[10824]_ , \new_[10825]_ ,
    \new_[10826]_ , \new_[10827]_ , \new_[10828]_ , \new_[10829]_ ,
    \new_[10830]_ , \new_[10831]_ , \new_[10832]_ , \new_[10833]_ ,
    \new_[10834]_ , \new_[10835]_ , \new_[10836]_ , \new_[10837]_ ,
    \new_[10838]_ , \new_[10839]_ , \new_[10840]_ , \new_[10841]_ ,
    \new_[10842]_ , \new_[10843]_ , \new_[10844]_ , \new_[10845]_ ,
    \new_[10846]_ , \new_[10847]_ , \new_[10848]_ , \new_[10849]_ ,
    \new_[10850]_ , \new_[10851]_ , \new_[10852]_ , \new_[10853]_ ,
    \new_[10854]_ , \new_[10855]_ , \new_[10856]_ , \new_[10857]_ ,
    \new_[10858]_ , \new_[10859]_ , \new_[10860]_ , \new_[10861]_ ,
    \new_[10862]_ , \new_[10863]_ , \new_[10864]_ , \new_[10865]_ ,
    \new_[10866]_ , \new_[10867]_ , \new_[10868]_ , \new_[10869]_ ,
    \new_[10870]_ , \new_[10871]_ , \new_[10872]_ , \new_[10873]_ ,
    \new_[10874]_ , \new_[10875]_ , \new_[10876]_ , \new_[10877]_ ,
    \new_[10878]_ , \new_[10879]_ , \new_[10880]_ , \new_[10881]_ ,
    \new_[10882]_ , \new_[10883]_ , \new_[10884]_ , \new_[10885]_ ,
    \new_[10886]_ , \new_[10887]_ , \new_[10888]_ , \new_[10889]_ ,
    \new_[10890]_ , \new_[10891]_ , \new_[10892]_ , \new_[10893]_ ,
    \new_[10894]_ , \new_[10895]_ , \new_[10896]_ , \new_[10897]_ ,
    \new_[10898]_ , \new_[10899]_ , \new_[10900]_ , \new_[10901]_ ,
    \new_[10902]_ , \new_[10903]_ , \new_[10904]_ , \new_[10905]_ ,
    \new_[10906]_ , \new_[10907]_ , \new_[10908]_ , \new_[10909]_ ,
    \new_[10910]_ , \new_[10911]_ , \new_[10912]_ , \new_[10913]_ ,
    \new_[10914]_ , \new_[10915]_ , \new_[10916]_ , \new_[10917]_ ,
    \new_[10918]_ , \new_[10919]_ , \new_[10920]_ , \new_[10921]_ ,
    \new_[10922]_ , \new_[10923]_ , \new_[10924]_ , \new_[10925]_ ,
    \new_[10926]_ , \new_[10927]_ , \new_[10928]_ , \new_[10929]_ ,
    \new_[10930]_ , \new_[10931]_ , \new_[10932]_ , \new_[10933]_ ,
    \new_[10934]_ , \new_[10935]_ , \new_[10936]_ , \new_[10937]_ ,
    \new_[10938]_ , \new_[10939]_ , \new_[10940]_ , \new_[10941]_ ,
    \new_[10942]_ , \new_[10943]_ , \new_[10944]_ , \new_[10945]_ ,
    \new_[10946]_ , \new_[10947]_ , \new_[10948]_ , \new_[10949]_ ,
    \new_[10950]_ , \new_[10951]_ , \new_[10952]_ , \new_[10953]_ ,
    \new_[10954]_ , \new_[10955]_ , \new_[10956]_ , \new_[10957]_ ,
    \new_[10958]_ , \new_[10959]_ , \new_[10960]_ , \new_[10961]_ ,
    \new_[10962]_ , \new_[10963]_ , \new_[10964]_ , \new_[10965]_ ,
    \new_[10966]_ , \new_[10967]_ , \new_[10968]_ , \new_[10969]_ ,
    \new_[10970]_ , \new_[10971]_ , \new_[10972]_ , \new_[10973]_ ,
    \new_[10974]_ , \new_[10975]_ , \new_[10976]_ , \new_[10977]_ ,
    \new_[10978]_ , \new_[10979]_ , \new_[10980]_ , \new_[10981]_ ,
    \new_[10982]_ , \new_[10983]_ , \new_[10984]_ , \new_[10985]_ ,
    \new_[10986]_ , \new_[10987]_ , \new_[10988]_ , \new_[10989]_ ,
    \new_[10990]_ , \new_[10991]_ , \new_[10992]_ , \new_[10993]_ ,
    \new_[10994]_ , \new_[10995]_ , \new_[10996]_ , \new_[10997]_ ,
    \new_[10998]_ , \new_[10999]_ , \new_[11000]_ , \new_[11001]_ ,
    \new_[11002]_ , \new_[11003]_ , \new_[11004]_ , \new_[11005]_ ,
    \new_[11006]_ , \new_[11007]_ , \new_[11008]_ , \new_[11009]_ ,
    \new_[11010]_ , \new_[11011]_ , \new_[11012]_ , \new_[11013]_ ,
    \new_[11014]_ , \new_[11015]_ , \new_[11016]_ , \new_[11017]_ ,
    \new_[11018]_ , \new_[11019]_ , \new_[11020]_ , \new_[11021]_ ,
    \new_[11022]_ , \new_[11023]_ , \new_[11024]_ , \new_[11025]_ ,
    \new_[11026]_ , \new_[11027]_ , \new_[11028]_ , \new_[11029]_ ,
    \new_[11030]_ , \new_[11031]_ , \new_[11032]_ , \new_[11033]_ ,
    \new_[11034]_ , \new_[11035]_ , \new_[11036]_ , \new_[11037]_ ,
    \new_[11038]_ , \new_[11039]_ , \new_[11040]_ , \new_[11041]_ ,
    \new_[11042]_ , \new_[11043]_ , \new_[11044]_ , \new_[11045]_ ,
    \new_[11046]_ , \new_[11047]_ , \new_[11048]_ , \new_[11049]_ ,
    \new_[11050]_ , \new_[11051]_ , \new_[11052]_ , \new_[11053]_ ,
    \new_[11054]_ , \new_[11055]_ , \new_[11056]_ , \new_[11057]_ ,
    \new_[11058]_ , \new_[11059]_ , \new_[11060]_ , \new_[11061]_ ,
    \new_[11062]_ , \new_[11063]_ , \new_[11064]_ , \new_[11065]_ ,
    \new_[11066]_ , \new_[11067]_ , \new_[11068]_ , \new_[11069]_ ,
    \new_[11070]_ , \new_[11071]_ , \new_[11072]_ , \new_[11073]_ ,
    \new_[11074]_ , \new_[11075]_ , \new_[11076]_ , \new_[11077]_ ,
    \new_[11078]_ , \new_[11079]_ , \new_[11080]_ , \new_[11081]_ ,
    \new_[11082]_ , \new_[11083]_ , \new_[11084]_ , \new_[11085]_ ,
    \new_[11086]_ , \new_[11087]_ , \new_[11088]_ , \new_[11089]_ ,
    \new_[11090]_ , \new_[11091]_ , \new_[11092]_ , \new_[11093]_ ,
    \new_[11094]_ , \new_[11095]_ , \new_[11096]_ , \new_[11097]_ ,
    \new_[11098]_ , \new_[11099]_ , \new_[11100]_ , \new_[11101]_ ,
    \new_[11102]_ , \new_[11103]_ , \new_[11104]_ , \new_[11105]_ ,
    \new_[11106]_ , \new_[11107]_ , \new_[11108]_ , \new_[11109]_ ,
    \new_[11110]_ , \new_[11111]_ , \new_[11112]_ , \new_[11113]_ ,
    \new_[11114]_ , \new_[11115]_ , \new_[11116]_ , \new_[11117]_ ,
    \new_[11118]_ , \new_[11119]_ , \new_[11120]_ , \new_[11121]_ ,
    \new_[11122]_ , \new_[11123]_ , \new_[11124]_ , \new_[11125]_ ,
    \new_[11126]_ , \new_[11127]_ , \new_[11128]_ , \new_[11129]_ ,
    \new_[11130]_ , \new_[11131]_ , \new_[11132]_ , \new_[11133]_ ,
    \new_[11134]_ , \new_[11135]_ , \new_[11136]_ , \new_[11137]_ ,
    \new_[11138]_ , \new_[11139]_ , \new_[11140]_ , \new_[11141]_ ,
    \new_[11142]_ , \new_[11143]_ , \new_[11144]_ , \new_[11145]_ ,
    \new_[11146]_ , \new_[11147]_ , \new_[11148]_ , \new_[11149]_ ,
    \new_[11150]_ , \new_[11151]_ , \new_[11152]_ , \new_[11153]_ ,
    \new_[11154]_ , \new_[11155]_ , \new_[11156]_ , \new_[11157]_ ,
    \new_[11158]_ , \new_[11159]_ , \new_[11160]_ , \new_[11161]_ ,
    \new_[11162]_ , \new_[11163]_ , \new_[11164]_ , \new_[11165]_ ,
    \new_[11166]_ , \new_[11167]_ , \new_[11168]_ , \new_[11169]_ ,
    \new_[11170]_ , \new_[11171]_ , \new_[11172]_ , \new_[11173]_ ,
    \new_[11174]_ , \new_[11175]_ , \new_[11176]_ , \new_[11177]_ ,
    \new_[11178]_ , \new_[11179]_ , \new_[11180]_ , \new_[11181]_ ,
    \new_[11182]_ , \new_[11183]_ , \new_[11184]_ , \new_[11185]_ ,
    \new_[11186]_ , \new_[11187]_ , \new_[11188]_ , \new_[11189]_ ,
    \new_[11190]_ , \new_[11191]_ , \new_[11192]_ , \new_[11193]_ ,
    \new_[11194]_ , \new_[11195]_ , \new_[11196]_ , \new_[11197]_ ,
    \new_[11198]_ , \new_[11199]_ , \new_[11200]_ , \new_[11201]_ ,
    \new_[11202]_ , \new_[11203]_ , \new_[11204]_ , \new_[11205]_ ,
    \new_[11206]_ , \new_[11207]_ , \new_[11208]_ , \new_[11209]_ ,
    \new_[11210]_ , \new_[11211]_ , \new_[11212]_ , \new_[11213]_ ,
    \new_[11214]_ , \new_[11215]_ , \new_[11216]_ , \new_[11217]_ ,
    \new_[11218]_ , \new_[11219]_ , \new_[11220]_ , \new_[11221]_ ,
    \new_[11222]_ , \new_[11223]_ , \new_[11224]_ , \new_[11225]_ ,
    \new_[11226]_ , \new_[11227]_ , \new_[11228]_ , \new_[11229]_ ,
    \new_[11231]_ , \new_[11232]_ , \new_[11233]_ , \new_[11234]_ ,
    \new_[11235]_ , \new_[11236]_ , \new_[11237]_ , \new_[11238]_ ,
    \new_[11239]_ , \new_[11240]_ , \new_[11241]_ , \new_[11242]_ ,
    \new_[11243]_ , \new_[11244]_ , \new_[11245]_ , \new_[11246]_ ,
    \new_[11247]_ , \new_[11248]_ , \new_[11249]_ , \new_[11250]_ ,
    \new_[11251]_ , \new_[11252]_ , \new_[11253]_ , \new_[11254]_ ,
    \new_[11255]_ , \new_[11256]_ , \new_[11257]_ , \new_[11258]_ ,
    \new_[11259]_ , \new_[11260]_ , \new_[11261]_ , \new_[11262]_ ,
    \new_[11263]_ , \new_[11264]_ , \new_[11265]_ , \new_[11266]_ ,
    \new_[11267]_ , \new_[11268]_ , \new_[11269]_ , \new_[11270]_ ,
    \new_[11271]_ , \new_[11272]_ , \new_[11273]_ , \new_[11274]_ ,
    \new_[11275]_ , \new_[11276]_ , \new_[11277]_ , \new_[11278]_ ,
    \new_[11279]_ , \new_[11280]_ , \new_[11281]_ , \new_[11282]_ ,
    \new_[11283]_ , \new_[11284]_ , \new_[11285]_ , \new_[11286]_ ,
    \new_[11287]_ , \new_[11288]_ , \new_[11289]_ , \new_[11290]_ ,
    \new_[11291]_ , \new_[11292]_ , \new_[11293]_ , \new_[11294]_ ,
    \new_[11295]_ , \new_[11296]_ , \new_[11297]_ , \new_[11298]_ ,
    \new_[11299]_ , \new_[11300]_ , \new_[11301]_ , \new_[11302]_ ,
    \new_[11303]_ , \new_[11304]_ , \new_[11305]_ , \new_[11306]_ ,
    \new_[11307]_ , \new_[11308]_ , \new_[11309]_ , \new_[11310]_ ,
    \new_[11311]_ , \new_[11312]_ , \new_[11313]_ , \new_[11314]_ ,
    \new_[11315]_ , \new_[11316]_ , \new_[11317]_ , \new_[11318]_ ,
    \new_[11319]_ , \new_[11320]_ , \new_[11321]_ , \new_[11322]_ ,
    \new_[11323]_ , \new_[11324]_ , \new_[11325]_ , \new_[11326]_ ,
    \new_[11327]_ , \new_[11328]_ , \new_[11329]_ , \new_[11330]_ ,
    \new_[11331]_ , \new_[11332]_ , \new_[11333]_ , \new_[11334]_ ,
    \new_[11335]_ , \new_[11336]_ , \new_[11337]_ , \new_[11338]_ ,
    \new_[11339]_ , \new_[11340]_ , \new_[11341]_ , \new_[11342]_ ,
    \new_[11343]_ , \new_[11344]_ , \new_[11345]_ , \new_[11346]_ ,
    \new_[11347]_ , \new_[11348]_ , \new_[11349]_ , \new_[11350]_ ,
    \new_[11351]_ , \new_[11352]_ , \new_[11353]_ , \new_[11354]_ ,
    \new_[11355]_ , \new_[11356]_ , \new_[11357]_ , \new_[11358]_ ,
    \new_[11359]_ , \new_[11360]_ , \new_[11361]_ , \new_[11362]_ ,
    \new_[11363]_ , \new_[11364]_ , \new_[11365]_ , \new_[11366]_ ,
    \new_[11367]_ , \new_[11368]_ , \new_[11369]_ , \new_[11370]_ ,
    \new_[11371]_ , \new_[11372]_ , \new_[11373]_ , \new_[11374]_ ,
    \new_[11375]_ , \new_[11376]_ , \new_[11377]_ , \new_[11378]_ ,
    \new_[11379]_ , \new_[11380]_ , \new_[11381]_ , \new_[11382]_ ,
    \new_[11383]_ , \new_[11384]_ , \new_[11385]_ , \new_[11386]_ ,
    \new_[11387]_ , \new_[11388]_ , \new_[11389]_ , \new_[11390]_ ,
    \new_[11391]_ , \new_[11392]_ , \new_[11393]_ , \new_[11394]_ ,
    \new_[11395]_ , \new_[11396]_ , \new_[11397]_ , \new_[11398]_ ,
    \new_[11399]_ , \new_[11400]_ , \new_[11401]_ , \new_[11402]_ ,
    \new_[11403]_ , \new_[11404]_ , \new_[11405]_ , \new_[11406]_ ,
    \new_[11407]_ , \new_[11408]_ , \new_[11409]_ , \new_[11410]_ ,
    \new_[11411]_ , \new_[11412]_ , \new_[11413]_ , \new_[11414]_ ,
    \new_[11415]_ , \new_[11416]_ , \new_[11417]_ , \new_[11418]_ ,
    \new_[11419]_ , \new_[11420]_ , \new_[11421]_ , \new_[11422]_ ,
    \new_[11423]_ , \new_[11424]_ , \new_[11425]_ , \new_[11426]_ ,
    \new_[11427]_ , \new_[11428]_ , \new_[11429]_ , \new_[11430]_ ,
    \new_[11431]_ , \new_[11432]_ , \new_[11433]_ , \new_[11434]_ ,
    \new_[11435]_ , \new_[11436]_ , \new_[11437]_ , \new_[11438]_ ,
    \new_[11439]_ , \new_[11440]_ , \new_[11441]_ , \new_[11442]_ ,
    \new_[11443]_ , \new_[11444]_ , \new_[11445]_ , \new_[11446]_ ,
    \new_[11447]_ , \new_[11448]_ , \new_[11449]_ , \new_[11450]_ ,
    \new_[11451]_ , \new_[11452]_ , \new_[11453]_ , \new_[11454]_ ,
    \new_[11455]_ , \new_[11456]_ , \new_[11457]_ , \new_[11458]_ ,
    \new_[11459]_ , \new_[11460]_ , \new_[11461]_ , \new_[11462]_ ,
    \new_[11463]_ , \new_[11464]_ , \new_[11465]_ , \new_[11466]_ ,
    \new_[11467]_ , \new_[11468]_ , \new_[11469]_ , \new_[11470]_ ,
    \new_[11471]_ , \new_[11472]_ , \new_[11473]_ , \new_[11474]_ ,
    \new_[11475]_ , \new_[11476]_ , \new_[11477]_ , \new_[11478]_ ,
    \new_[11479]_ , \new_[11480]_ , \new_[11481]_ , \new_[11482]_ ,
    \new_[11483]_ , \new_[11484]_ , \new_[11485]_ , \new_[11486]_ ,
    \new_[11487]_ , \new_[11488]_ , \new_[11489]_ , \new_[11490]_ ,
    \new_[11491]_ , \new_[11492]_ , \new_[11493]_ , \new_[11494]_ ,
    \new_[11495]_ , \new_[11496]_ , \new_[11497]_ , \new_[11498]_ ,
    \new_[11499]_ , \new_[11500]_ , \new_[11501]_ , \new_[11502]_ ,
    \new_[11503]_ , \new_[11504]_ , \new_[11505]_ , \new_[11506]_ ,
    \new_[11507]_ , \new_[11508]_ , \new_[11509]_ , \new_[11510]_ ,
    \new_[11511]_ , \new_[11512]_ , \new_[11513]_ , \new_[11514]_ ,
    \new_[11515]_ , \new_[11516]_ , \new_[11517]_ , \new_[11518]_ ,
    \new_[11519]_ , \new_[11520]_ , \new_[11521]_ , \new_[11522]_ ,
    \new_[11523]_ , \new_[11524]_ , \new_[11525]_ , \new_[11526]_ ,
    \new_[11527]_ , \new_[11528]_ , \new_[11529]_ , \new_[11530]_ ,
    \new_[11531]_ , \new_[11532]_ , \new_[11533]_ , \new_[11534]_ ,
    \new_[11535]_ , \new_[11536]_ , \new_[11537]_ , \new_[11538]_ ,
    \new_[11539]_ , \new_[11540]_ , \new_[11541]_ , \new_[11542]_ ,
    \new_[11543]_ , \new_[11544]_ , \new_[11545]_ , \new_[11546]_ ,
    \new_[11547]_ , \new_[11548]_ , \new_[11549]_ , \new_[11550]_ ,
    \new_[11551]_ , \new_[11552]_ , \new_[11553]_ , \new_[11554]_ ,
    \new_[11555]_ , \new_[11556]_ , \new_[11557]_ , \new_[11558]_ ,
    \new_[11559]_ , \new_[11560]_ , \new_[11561]_ , \new_[11562]_ ,
    \new_[11563]_ , \new_[11564]_ , \new_[11565]_ , \new_[11566]_ ,
    \new_[11567]_ , \new_[11568]_ , \new_[11569]_ , \new_[11570]_ ,
    \new_[11571]_ , \new_[11572]_ , \new_[11573]_ , \new_[11574]_ ,
    \new_[11575]_ , \new_[11576]_ , \new_[11577]_ , \new_[11578]_ ,
    \new_[11579]_ , \new_[11580]_ , \new_[11581]_ , \new_[11582]_ ,
    \new_[11583]_ , \new_[11584]_ , \new_[11585]_ , \new_[11586]_ ,
    \new_[11587]_ , \new_[11588]_ , \new_[11589]_ , \new_[11590]_ ,
    \new_[11591]_ , \new_[11592]_ , \new_[11593]_ , \new_[11594]_ ,
    \new_[11595]_ , \new_[11596]_ , \new_[11597]_ , \new_[11598]_ ,
    \new_[11599]_ , \new_[11600]_ , \new_[11601]_ , \new_[11602]_ ,
    \new_[11603]_ , \new_[11604]_ , \new_[11605]_ , \new_[11606]_ ,
    \new_[11607]_ , \new_[11608]_ , \new_[11609]_ , \new_[11610]_ ,
    \new_[11611]_ , \new_[11612]_ , \new_[11613]_ , \new_[11614]_ ,
    \new_[11615]_ , \new_[11616]_ , \new_[11617]_ , \new_[11618]_ ,
    \new_[11619]_ , \new_[11620]_ , \new_[11621]_ , \new_[11622]_ ,
    \new_[11623]_ , \new_[11624]_ , \new_[11625]_ , \new_[11626]_ ,
    \new_[11627]_ , \new_[11628]_ , \new_[11629]_ , \new_[11630]_ ,
    \new_[11631]_ , \new_[11632]_ , \new_[11633]_ , \new_[11634]_ ,
    \new_[11635]_ , \new_[11636]_ , \new_[11637]_ , \new_[11638]_ ,
    \new_[11639]_ , \new_[11640]_ , \new_[11641]_ , \new_[11642]_ ,
    \new_[11643]_ , \new_[11644]_ , \new_[11645]_ , \new_[11646]_ ,
    \new_[11647]_ , \new_[11648]_ , \new_[11649]_ , \new_[11650]_ ,
    \new_[11651]_ , \new_[11652]_ , \new_[11653]_ , \new_[11654]_ ,
    \new_[11655]_ , \new_[11656]_ , \new_[11657]_ , \new_[11658]_ ,
    \new_[11659]_ , \new_[11660]_ , \new_[11661]_ , \new_[11662]_ ,
    \new_[11663]_ , \new_[11664]_ , \new_[11665]_ , \new_[11666]_ ,
    \new_[11667]_ , \new_[11668]_ , \new_[11669]_ , \new_[11670]_ ,
    \new_[11671]_ , \new_[11672]_ , \new_[11673]_ , \new_[11674]_ ,
    \new_[11675]_ , \new_[11676]_ , \new_[11677]_ , \new_[11678]_ ,
    \new_[11679]_ , \new_[11680]_ , \new_[11681]_ , \new_[11682]_ ,
    \new_[11683]_ , \new_[11684]_ , \new_[11685]_ , \new_[11686]_ ,
    \new_[11687]_ , \new_[11688]_ , \new_[11689]_ , \new_[11690]_ ,
    \new_[11691]_ , \new_[11692]_ , \new_[11693]_ , \new_[11694]_ ,
    \new_[11695]_ , \new_[11696]_ , \new_[11697]_ , \new_[11698]_ ,
    \new_[11699]_ , \new_[11700]_ , \new_[11701]_ , \new_[11702]_ ,
    \new_[11703]_ , \new_[11704]_ , \new_[11705]_ , \new_[11706]_ ,
    \new_[11707]_ , \new_[11708]_ , \new_[11709]_ , \new_[11710]_ ,
    \new_[11711]_ , \new_[11712]_ , \new_[11713]_ , \new_[11714]_ ,
    \new_[11715]_ , \new_[11716]_ , \new_[11717]_ , \new_[11718]_ ,
    \new_[11719]_ , \new_[11720]_ , \new_[11721]_ , \new_[11722]_ ,
    \new_[11723]_ , \new_[11724]_ , \new_[11725]_ , \new_[11726]_ ,
    \new_[11727]_ , \new_[11728]_ , \new_[11729]_ , \new_[11730]_ ,
    \new_[11731]_ , \new_[11732]_ , \new_[11733]_ , \new_[11734]_ ,
    \new_[11735]_ , \new_[11736]_ , \new_[11737]_ , \new_[11738]_ ,
    \new_[11739]_ , \new_[11740]_ , \new_[11741]_ , \new_[11742]_ ,
    \new_[11743]_ , \new_[11744]_ , \new_[11745]_ , \new_[11746]_ ,
    \new_[11747]_ , \new_[11748]_ , \new_[11749]_ , \new_[11750]_ ,
    \new_[11751]_ , \new_[11752]_ , \new_[11753]_ , \new_[11754]_ ,
    \new_[11755]_ , \new_[11756]_ , \new_[11757]_ , \new_[11758]_ ,
    \new_[11759]_ , \new_[11760]_ , \new_[11761]_ , \new_[11762]_ ,
    \new_[11763]_ , \new_[11764]_ , \new_[11765]_ , \new_[11766]_ ,
    \new_[11767]_ , \new_[11768]_ , \new_[11769]_ , \new_[11770]_ ,
    \new_[11771]_ , \new_[11772]_ , \new_[11773]_ , \new_[11774]_ ,
    \new_[11775]_ , \new_[11776]_ , \new_[11777]_ , \new_[11778]_ ,
    \new_[11779]_ , \new_[11780]_ , \new_[11781]_ , \new_[11782]_ ,
    \new_[11783]_ , \new_[11784]_ , \new_[11785]_ , \new_[11786]_ ,
    \new_[11787]_ , \new_[11788]_ , \new_[11789]_ , \new_[11790]_ ,
    \new_[11791]_ , \new_[11792]_ , \new_[11793]_ , \new_[11794]_ ,
    \new_[11795]_ , \new_[11796]_ , \new_[11797]_ , \new_[11798]_ ,
    \new_[11799]_ , \new_[11800]_ , \new_[11801]_ , \new_[11802]_ ,
    \new_[11803]_ , \new_[11804]_ , \new_[11805]_ , \new_[11806]_ ,
    \new_[11807]_ , \new_[11808]_ , \new_[11809]_ , \new_[11810]_ ,
    \new_[11811]_ , \new_[11812]_ , \new_[11813]_ , \new_[11814]_ ,
    \new_[11815]_ , \new_[11816]_ , \new_[11817]_ , \new_[11818]_ ,
    \new_[11819]_ , \new_[11820]_ , \new_[11821]_ , \new_[11822]_ ,
    \new_[11823]_ , \new_[11824]_ , \new_[11825]_ , \new_[11826]_ ,
    \new_[11827]_ , \new_[11828]_ , \new_[11829]_ , \new_[11830]_ ,
    \new_[11831]_ , \new_[11832]_ , \new_[11833]_ , \new_[11834]_ ,
    \new_[11835]_ , \new_[11836]_ , \new_[11837]_ , \new_[11838]_ ,
    \new_[11839]_ , \new_[11840]_ , \new_[11841]_ , \new_[11842]_ ,
    \new_[11843]_ , \new_[11844]_ , \new_[11845]_ , \new_[11846]_ ,
    \new_[11847]_ , \new_[11848]_ , \new_[11849]_ , \new_[11850]_ ,
    \new_[11851]_ , \new_[11852]_ , \new_[11853]_ , \new_[11854]_ ,
    \new_[11855]_ , \new_[11856]_ , \new_[11857]_ , \new_[11858]_ ,
    \new_[11859]_ , \new_[11860]_ , \new_[11861]_ , \new_[11862]_ ,
    \new_[11863]_ , \new_[11864]_ , \new_[11865]_ , \new_[11866]_ ,
    \new_[11867]_ , \new_[11868]_ , \new_[11869]_ , \new_[11870]_ ,
    \new_[11871]_ , \new_[11872]_ , \new_[11873]_ , \new_[11874]_ ,
    \new_[11875]_ , \new_[11876]_ , \new_[11877]_ , \new_[11878]_ ,
    \new_[11879]_ , \new_[11880]_ , \new_[11881]_ , \new_[11882]_ ,
    \new_[11883]_ , \new_[11884]_ , \new_[11885]_ , \new_[11886]_ ,
    \new_[11887]_ , \new_[11888]_ , \new_[11889]_ , \new_[11890]_ ,
    \new_[11891]_ , \new_[11892]_ , \new_[11893]_ , \new_[11894]_ ,
    \new_[11895]_ , \new_[11896]_ , \new_[11897]_ , \new_[11898]_ ,
    \new_[11899]_ , \new_[11900]_ , \new_[11901]_ , \new_[11902]_ ,
    \new_[11903]_ , \new_[11904]_ , \new_[11905]_ , \new_[11906]_ ,
    \new_[11907]_ , \new_[11908]_ , \new_[11909]_ , \new_[11910]_ ,
    \new_[11911]_ , \new_[11912]_ , \new_[11913]_ , \new_[11914]_ ,
    \new_[11915]_ , \new_[11916]_ , \new_[11917]_ , \new_[11918]_ ,
    \new_[11919]_ , \new_[11920]_ , \new_[11921]_ , \new_[11922]_ ,
    \new_[11923]_ , \new_[11924]_ , \new_[11925]_ , \new_[11926]_ ,
    \new_[11927]_ , \new_[11928]_ , \new_[11929]_ , \new_[11930]_ ,
    \new_[11931]_ , \new_[11932]_ , \new_[11933]_ , \new_[11934]_ ,
    \new_[11935]_ , \new_[11936]_ , \new_[11937]_ , \new_[11938]_ ,
    \new_[11939]_ , \new_[11940]_ , \new_[11941]_ , \new_[11942]_ ,
    \new_[11943]_ , \new_[11944]_ , \new_[11945]_ , \new_[11946]_ ,
    \new_[11947]_ , \new_[11948]_ , \new_[11949]_ , \new_[11950]_ ,
    \new_[11951]_ , \new_[11952]_ , \new_[11953]_ , \new_[11954]_ ,
    \new_[11955]_ , \new_[11956]_ , \new_[11957]_ , \new_[11958]_ ,
    \new_[11959]_ , \new_[11960]_ , \new_[11961]_ , \new_[11962]_ ,
    \new_[11963]_ , \new_[11964]_ , \new_[11965]_ , \new_[11966]_ ,
    \new_[11967]_ , \new_[11968]_ , \new_[11969]_ , \new_[11970]_ ,
    \new_[11971]_ , \new_[11972]_ , \new_[11973]_ , \new_[11974]_ ,
    \new_[11975]_ , \new_[11976]_ , \new_[11977]_ , \new_[11978]_ ,
    \new_[11979]_ , \new_[11980]_ , \new_[11981]_ , \new_[11982]_ ,
    \new_[11983]_ , \new_[11984]_ , \new_[11985]_ , \new_[11986]_ ,
    \new_[11987]_ , \new_[11988]_ , \new_[11989]_ , \new_[11990]_ ,
    \new_[11991]_ , \new_[11992]_ , \new_[11993]_ , \new_[11994]_ ,
    \new_[11995]_ , \new_[11996]_ , \new_[11997]_ , \new_[11998]_ ,
    \new_[11999]_ , \new_[12000]_ , \new_[12001]_ , \new_[12002]_ ,
    \new_[12003]_ , \new_[12004]_ , \new_[12005]_ , \new_[12006]_ ,
    \new_[12007]_ , \new_[12008]_ , \new_[12009]_ , \new_[12010]_ ,
    \new_[12011]_ , \new_[12012]_ , \new_[12013]_ , \new_[12014]_ ,
    \new_[12015]_ , \new_[12016]_ , \new_[12017]_ , \new_[12018]_ ,
    \new_[12019]_ , \new_[12020]_ , \new_[12021]_ , \new_[12022]_ ,
    \new_[12023]_ , \new_[12024]_ , \new_[12025]_ , \new_[12026]_ ,
    \new_[12027]_ , \new_[12028]_ , \new_[12029]_ , \new_[12030]_ ,
    \new_[12031]_ , \new_[12032]_ , \new_[12033]_ , \new_[12034]_ ,
    \new_[12035]_ , \new_[12036]_ , \new_[12037]_ , \new_[12038]_ ,
    \new_[12039]_ , \new_[12040]_ , \new_[12041]_ , \new_[12042]_ ,
    \new_[12043]_ , \new_[12044]_ , \new_[12045]_ , \new_[12046]_ ,
    \new_[12047]_ , \new_[12048]_ , \new_[12049]_ , \new_[12050]_ ,
    \new_[12051]_ , \new_[12052]_ , \new_[12053]_ , \new_[12054]_ ,
    \new_[12055]_ , \new_[12056]_ , \new_[12057]_ , \new_[12058]_ ,
    \new_[12059]_ , \new_[12060]_ , \new_[12061]_ , \new_[12062]_ ,
    \new_[12063]_ , \new_[12064]_ , \new_[12065]_ , \new_[12066]_ ,
    \new_[12067]_ , \new_[12068]_ , \new_[12069]_ , \new_[12070]_ ,
    \new_[12071]_ , \new_[12072]_ , \new_[12073]_ , \new_[12074]_ ,
    \new_[12075]_ , \new_[12076]_ , \new_[12077]_ , \new_[12078]_ ,
    \new_[12079]_ , \new_[12080]_ , \new_[12081]_ , \new_[12082]_ ,
    \new_[12084]_ , \new_[12085]_ , \new_[12086]_ , \new_[12087]_ ,
    \new_[12088]_ , \new_[12089]_ , \new_[12090]_ , \new_[12091]_ ,
    \new_[12092]_ , \new_[12093]_ , \new_[12094]_ , \new_[12095]_ ,
    \new_[12096]_ , \new_[12097]_ , \new_[12098]_ , \new_[12099]_ ,
    \new_[12100]_ , \new_[12101]_ , \new_[12102]_ , \new_[12103]_ ,
    \new_[12104]_ , \new_[12105]_ , \new_[12106]_ , \new_[12107]_ ,
    \new_[12108]_ , \new_[12109]_ , \new_[12110]_ , \new_[12111]_ ,
    \new_[12112]_ , \new_[12113]_ , \new_[12114]_ , \new_[12115]_ ,
    \new_[12116]_ , \new_[12117]_ , \new_[12118]_ , \new_[12119]_ ,
    \new_[12120]_ , \new_[12121]_ , \new_[12122]_ , \new_[12123]_ ,
    \new_[12124]_ , \new_[12125]_ , \new_[12126]_ , \new_[12127]_ ,
    \new_[12128]_ , \new_[12129]_ , \new_[12130]_ , \new_[12131]_ ,
    \new_[12132]_ , \new_[12133]_ , \new_[12134]_ , \new_[12135]_ ,
    \new_[12136]_ , \new_[12137]_ , \new_[12138]_ , \new_[12139]_ ,
    \new_[12140]_ , \new_[12141]_ , \new_[12142]_ , \new_[12143]_ ,
    \new_[12144]_ , \new_[12145]_ , \new_[12146]_ , \new_[12147]_ ,
    \new_[12148]_ , \new_[12149]_ , \new_[12150]_ , \new_[12151]_ ,
    \new_[12152]_ , \new_[12153]_ , \new_[12154]_ , \new_[12155]_ ,
    \new_[12156]_ , \new_[12157]_ , \new_[12158]_ , \new_[12159]_ ,
    \new_[12160]_ , \new_[12161]_ , \new_[12162]_ , \new_[12163]_ ,
    \new_[12164]_ , \new_[12165]_ , \new_[12166]_ , \new_[12167]_ ,
    \new_[12168]_ , \new_[12169]_ , \new_[12170]_ , \new_[12171]_ ,
    \new_[12172]_ , \new_[12173]_ , \new_[12174]_ , \new_[12175]_ ,
    \new_[12176]_ , \new_[12177]_ , \new_[12178]_ , \new_[12179]_ ,
    \new_[12180]_ , \new_[12181]_ , \new_[12182]_ , \new_[12183]_ ,
    \new_[12184]_ , \new_[12185]_ , \new_[12186]_ , \new_[12187]_ ,
    \new_[12188]_ , \new_[12189]_ , \new_[12190]_ , \new_[12191]_ ,
    \new_[12192]_ , \new_[12193]_ , \new_[12194]_ , \new_[12195]_ ,
    \new_[12196]_ , \new_[12197]_ , \new_[12198]_ , \new_[12199]_ ,
    \new_[12200]_ , \new_[12201]_ , \new_[12202]_ , \new_[12203]_ ,
    \new_[12204]_ , \new_[12205]_ , \new_[12206]_ , \new_[12207]_ ,
    \new_[12208]_ , \new_[12209]_ , \new_[12210]_ , \new_[12211]_ ,
    \new_[12212]_ , \new_[12213]_ , \new_[12214]_ , \new_[12215]_ ,
    \new_[12216]_ , \new_[12217]_ , \new_[12218]_ , \new_[12219]_ ,
    \new_[12220]_ , \new_[12221]_ , \new_[12222]_ , \new_[12223]_ ,
    \new_[12224]_ , \new_[12225]_ , \new_[12226]_ , \new_[12227]_ ,
    \new_[12228]_ , \new_[12229]_ , \new_[12230]_ , \new_[12231]_ ,
    \new_[12232]_ , \new_[12233]_ , \new_[12234]_ , \new_[12235]_ ,
    \new_[12236]_ , \new_[12237]_ , \new_[12238]_ , \new_[12239]_ ,
    \new_[12240]_ , \new_[12241]_ , \new_[12242]_ , \new_[12243]_ ,
    \new_[12244]_ , \new_[12245]_ , \new_[12246]_ , \new_[12247]_ ,
    \new_[12248]_ , \new_[12249]_ , \new_[12250]_ , \new_[12251]_ ,
    \new_[12252]_ , \new_[12253]_ , \new_[12254]_ , \new_[12255]_ ,
    \new_[12256]_ , \new_[12257]_ , \new_[12258]_ , \new_[12259]_ ,
    \new_[12260]_ , \new_[12261]_ , \new_[12262]_ , \new_[12263]_ ,
    \new_[12264]_ , \new_[12265]_ , \new_[12266]_ , \new_[12267]_ ,
    \new_[12268]_ , \new_[12269]_ , \new_[12270]_ , \new_[12271]_ ,
    \new_[12272]_ , \new_[12273]_ , \new_[12274]_ , \new_[12275]_ ,
    \new_[12276]_ , \new_[12277]_ , \new_[12278]_ , \new_[12279]_ ,
    \new_[12280]_ , \new_[12281]_ , \new_[12282]_ , \new_[12283]_ ,
    \new_[12284]_ , \new_[12285]_ , \new_[12286]_ , \new_[12287]_ ,
    \new_[12288]_ , \new_[12289]_ , \new_[12290]_ , \new_[12291]_ ,
    \new_[12292]_ , \new_[12293]_ , \new_[12294]_ , \new_[12295]_ ,
    \new_[12296]_ , \new_[12297]_ , \new_[12298]_ , \new_[12299]_ ,
    \new_[12300]_ , \new_[12301]_ , \new_[12302]_ , \new_[12303]_ ,
    \new_[12304]_ , \new_[12305]_ , \new_[12306]_ , \new_[12307]_ ,
    \new_[12308]_ , \new_[12309]_ , \new_[12310]_ , \new_[12311]_ ,
    \new_[12312]_ , \new_[12313]_ , \new_[12314]_ , \new_[12315]_ ,
    \new_[12316]_ , \new_[12317]_ , \new_[12318]_ , \new_[12319]_ ,
    \new_[12320]_ , \new_[12321]_ , \new_[12322]_ , \new_[12323]_ ,
    \new_[12324]_ , \new_[12325]_ , \new_[12326]_ , \new_[12327]_ ,
    \new_[12328]_ , \new_[12329]_ , \new_[12330]_ , \new_[12331]_ ,
    \new_[12332]_ , \new_[12333]_ , \new_[12334]_ , \new_[12335]_ ,
    \new_[12336]_ , \new_[12337]_ , \new_[12338]_ , \new_[12339]_ ,
    \new_[12340]_ , \new_[12341]_ , \new_[12342]_ , \new_[12343]_ ,
    \new_[12344]_ , \new_[12345]_ , \new_[12346]_ , \new_[12347]_ ,
    \new_[12348]_ , \new_[12349]_ , \new_[12350]_ , \new_[12351]_ ,
    \new_[12352]_ , \new_[12353]_ , \new_[12354]_ , \new_[12355]_ ,
    \new_[12356]_ , \new_[12357]_ , \new_[12358]_ , \new_[12359]_ ,
    \new_[12360]_ , \new_[12361]_ , \new_[12362]_ , \new_[12363]_ ,
    \new_[12364]_ , \new_[12365]_ , \new_[12366]_ , \new_[12367]_ ,
    \new_[12368]_ , \new_[12369]_ , \new_[12370]_ , \new_[12371]_ ,
    \new_[12372]_ , \new_[12373]_ , \new_[12374]_ , \new_[12375]_ ,
    \new_[12376]_ , \new_[12377]_ , \new_[12378]_ , \new_[12379]_ ,
    \new_[12380]_ , \new_[12381]_ , \new_[12382]_ , \new_[12383]_ ,
    \new_[12384]_ , \new_[12385]_ , \new_[12386]_ , \new_[12387]_ ,
    \new_[12388]_ , \new_[12389]_ , \new_[12390]_ , \new_[12391]_ ,
    \new_[12392]_ , \new_[12393]_ , \new_[12394]_ , \new_[12395]_ ,
    \new_[12396]_ , \new_[12397]_ , \new_[12398]_ , \new_[12399]_ ,
    \new_[12400]_ , \new_[12401]_ , \new_[12402]_ , \new_[12403]_ ,
    \new_[12404]_ , \new_[12405]_ , \new_[12406]_ , \new_[12407]_ ,
    \new_[12409]_ , \new_[12410]_ , \new_[12411]_ , \new_[12412]_ ,
    \new_[12413]_ , \new_[12414]_ , \new_[12415]_ , \new_[12416]_ ,
    \new_[12417]_ , \new_[12418]_ , \new_[12419]_ , \new_[12420]_ ,
    \new_[12421]_ , \new_[12422]_ , \new_[12423]_ , \new_[12424]_ ,
    \new_[12425]_ , \new_[12426]_ , \new_[12427]_ , \new_[12428]_ ,
    \new_[12429]_ , \new_[12430]_ , \new_[12431]_ , \new_[12432]_ ,
    \new_[12433]_ , \new_[12434]_ , \new_[12435]_ , \new_[12436]_ ,
    \new_[12437]_ , \new_[12438]_ , \new_[12439]_ , \new_[12440]_ ,
    \new_[12441]_ , \new_[12442]_ , \new_[12443]_ , \new_[12444]_ ,
    \new_[12445]_ , \new_[12446]_ , \new_[12447]_ , \new_[12448]_ ,
    \new_[12449]_ , \new_[12450]_ , \new_[12451]_ , \new_[12452]_ ,
    \new_[12453]_ , \new_[12454]_ , \new_[12455]_ , \new_[12456]_ ,
    \new_[12457]_ , \new_[12458]_ , \new_[12459]_ , \new_[12460]_ ,
    \new_[12461]_ , \new_[12462]_ , \new_[12463]_ , \new_[12464]_ ,
    \new_[12465]_ , \new_[12466]_ , \new_[12467]_ , \new_[12468]_ ,
    \new_[12469]_ , \new_[12470]_ , \new_[12471]_ , \new_[12472]_ ,
    \new_[12473]_ , \new_[12474]_ , \new_[12475]_ , \new_[12476]_ ,
    \new_[12477]_ , \new_[12478]_ , \new_[12479]_ , \new_[12480]_ ,
    \new_[12481]_ , \new_[12482]_ , \new_[12483]_ , \new_[12484]_ ,
    \new_[12485]_ , \new_[12486]_ , \new_[12487]_ , \new_[12488]_ ,
    \new_[12489]_ , \new_[12490]_ , \new_[12491]_ , \new_[12492]_ ,
    \new_[12493]_ , \new_[12494]_ , \new_[12495]_ , \new_[12496]_ ,
    \new_[12497]_ , \new_[12498]_ , \new_[12499]_ , \new_[12500]_ ,
    \new_[12501]_ , \new_[12502]_ , \new_[12503]_ , \new_[12504]_ ,
    \new_[12505]_ , \new_[12506]_ , \new_[12507]_ , \new_[12508]_ ,
    \new_[12509]_ , \new_[12510]_ , \new_[12511]_ , \new_[12512]_ ,
    \new_[12513]_ , \new_[12514]_ , \new_[12515]_ , \new_[12516]_ ,
    \new_[12517]_ , \new_[12518]_ , \new_[12519]_ , \new_[12520]_ ,
    \new_[12521]_ , \new_[12522]_ , \new_[12523]_ , \new_[12524]_ ,
    \new_[12525]_ , \new_[12526]_ , \new_[12527]_ , \new_[12528]_ ,
    \new_[12529]_ , \new_[12530]_ , \new_[12531]_ , \new_[12532]_ ,
    \new_[12533]_ , \new_[12534]_ , \new_[12535]_ , \new_[12536]_ ,
    \new_[12537]_ , \new_[12538]_ , \new_[12539]_ , \new_[12540]_ ,
    \new_[12541]_ , \new_[12542]_ , \new_[12543]_ , \new_[12544]_ ,
    \new_[12545]_ , \new_[12546]_ , \new_[12547]_ , \new_[12548]_ ,
    \new_[12549]_ , \new_[12550]_ , \new_[12551]_ , \new_[12552]_ ,
    \new_[12553]_ , \new_[12554]_ , \new_[12555]_ , \new_[12556]_ ,
    \new_[12557]_ , \new_[12558]_ , \new_[12559]_ , \new_[12560]_ ,
    \new_[12561]_ , \new_[12562]_ , \new_[12563]_ , \new_[12564]_ ,
    \new_[12565]_ , \new_[12566]_ , \new_[12567]_ , \new_[12568]_ ,
    \new_[12569]_ , \new_[12570]_ , \new_[12571]_ , \new_[12572]_ ,
    \new_[12573]_ , \new_[12574]_ , \new_[12575]_ , \new_[12576]_ ,
    \new_[12577]_ , \new_[12578]_ , \new_[12579]_ , \new_[12580]_ ,
    \new_[12581]_ , \new_[12582]_ , \new_[12583]_ , \new_[12584]_ ,
    \new_[12585]_ , \new_[12586]_ , \new_[12587]_ , \new_[12588]_ ,
    \new_[12589]_ , \new_[12590]_ , \new_[12591]_ , \new_[12592]_ ,
    \new_[12593]_ , \new_[12594]_ , \new_[12595]_ , \new_[12596]_ ,
    \new_[12597]_ , \new_[12598]_ , \new_[12599]_ , \new_[12600]_ ,
    \new_[12601]_ , \new_[12602]_ , \new_[12603]_ , \new_[12604]_ ,
    \new_[12605]_ , \new_[12606]_ , \new_[12607]_ , \new_[12608]_ ,
    \new_[12609]_ , \new_[12610]_ , \new_[12611]_ , \new_[12612]_ ,
    \new_[12613]_ , \new_[12614]_ , \new_[12615]_ , \new_[12616]_ ,
    \new_[12617]_ , \new_[12618]_ , \new_[12619]_ , \new_[12620]_ ,
    \new_[12621]_ , \new_[12622]_ , \new_[12623]_ , \new_[12624]_ ,
    \new_[12625]_ , \new_[12626]_ , \new_[12627]_ , \new_[12628]_ ,
    \new_[12629]_ , \new_[12630]_ , \new_[12631]_ , \new_[12632]_ ,
    \new_[12633]_ , \new_[12634]_ , \new_[12635]_ , \new_[12636]_ ,
    \new_[12637]_ , \new_[12638]_ , \new_[12639]_ , \new_[12640]_ ,
    \new_[12641]_ , \new_[12642]_ , \new_[12643]_ , \new_[12644]_ ,
    \new_[12645]_ , \new_[12646]_ , \new_[12647]_ , \new_[12648]_ ,
    \new_[12649]_ , \new_[12650]_ , \new_[12651]_ , \new_[12652]_ ,
    \new_[12653]_ , \new_[12654]_ , \new_[12655]_ , \new_[12656]_ ,
    \new_[12657]_ , \new_[12658]_ , \new_[12659]_ , \new_[12660]_ ,
    \new_[12661]_ , \new_[12662]_ , \new_[12663]_ , \new_[12664]_ ,
    \new_[12665]_ , \new_[12666]_ , \new_[12667]_ , \new_[12668]_ ,
    \new_[12669]_ , \new_[12670]_ , \new_[12671]_ , \new_[12672]_ ,
    \new_[12673]_ , \new_[12674]_ , \new_[12675]_ , \new_[12676]_ ,
    \new_[12677]_ , \new_[12678]_ , \new_[12679]_ , \new_[12680]_ ,
    \new_[12681]_ , \new_[12682]_ , \new_[12683]_ , \new_[12684]_ ,
    \new_[12685]_ , \new_[12686]_ , \new_[12687]_ , \new_[12688]_ ,
    \new_[12689]_ , \new_[12690]_ , \new_[12691]_ , \new_[12692]_ ,
    \new_[12693]_ , \new_[12694]_ , \new_[12695]_ , \new_[12696]_ ,
    \new_[12697]_ , \new_[12698]_ , \new_[12699]_ , \new_[12700]_ ,
    \new_[12701]_ , \new_[12702]_ , \new_[12703]_ , \new_[12704]_ ,
    \new_[12705]_ , \new_[12706]_ , \new_[12707]_ , \new_[12708]_ ,
    \new_[12709]_ , \new_[12710]_ , \new_[12711]_ , \new_[12712]_ ,
    \new_[12713]_ , \new_[12714]_ , \new_[12715]_ , \new_[12716]_ ,
    \new_[12717]_ , \new_[12718]_ , \new_[12719]_ , \new_[12720]_ ,
    \new_[12721]_ , \new_[12722]_ , \new_[12723]_ , \new_[12724]_ ,
    \new_[12725]_ , \new_[12726]_ , \new_[12727]_ , \new_[12728]_ ,
    \new_[12729]_ , \new_[12730]_ , \new_[12731]_ , \new_[12732]_ ,
    \new_[12733]_ , \new_[12734]_ , \new_[12735]_ , \new_[12736]_ ,
    \new_[12737]_ , \new_[12738]_ , \new_[12739]_ , \new_[12740]_ ,
    \new_[12741]_ , \new_[12742]_ , \new_[12743]_ , \new_[12744]_ ,
    \new_[12745]_ , \new_[12746]_ , \new_[12747]_ , \new_[12748]_ ,
    \new_[12749]_ , \new_[12750]_ , \new_[12751]_ , \new_[12752]_ ,
    \new_[12753]_ , \new_[12754]_ , \new_[12755]_ , \new_[12756]_ ,
    \new_[12757]_ , \new_[12758]_ , \new_[12759]_ , \new_[12760]_ ,
    \new_[12761]_ , \new_[12762]_ , \new_[12763]_ , \new_[12764]_ ,
    \new_[12765]_ , \new_[12766]_ , \new_[12767]_ , \new_[12768]_ ,
    \new_[12769]_ , \new_[12770]_ , \new_[12771]_ , \new_[12772]_ ,
    \new_[12773]_ , \new_[12774]_ , \new_[12775]_ , \new_[12776]_ ,
    \new_[12777]_ , \new_[12778]_ , \new_[12779]_ , \new_[12780]_ ,
    \new_[12781]_ , \new_[12782]_ , \new_[12783]_ , \new_[12784]_ ,
    \new_[12785]_ , \new_[12786]_ , \new_[12787]_ , \new_[12788]_ ,
    \new_[12789]_ , \new_[12790]_ , \new_[12791]_ , \new_[12792]_ ,
    \new_[12793]_ , \new_[12794]_ , \new_[12795]_ , \new_[12796]_ ,
    \new_[12797]_ , \new_[12798]_ , \new_[12799]_ , \new_[12800]_ ,
    \new_[12801]_ , \new_[12802]_ , \new_[12803]_ , \new_[12804]_ ,
    \new_[12805]_ , \new_[12806]_ , \new_[12807]_ , \new_[12808]_ ,
    \new_[12809]_ , \new_[12810]_ , \new_[12811]_ , \new_[12812]_ ,
    \new_[12813]_ , \new_[12814]_ , \new_[12815]_ , \new_[12816]_ ,
    \new_[12817]_ , \new_[12818]_ , \new_[12819]_ , \new_[12820]_ ,
    \new_[12821]_ , \new_[12822]_ , \new_[12823]_ , \new_[12824]_ ,
    \new_[12825]_ , \new_[12826]_ , \new_[12827]_ , \new_[12828]_ ,
    \new_[12829]_ , \new_[12830]_ , \new_[12831]_ , \new_[12832]_ ,
    \new_[12833]_ , \new_[12834]_ , \new_[12835]_ , \new_[12836]_ ,
    \new_[12837]_ , \new_[12838]_ , \new_[12839]_ , \new_[12840]_ ,
    \new_[12841]_ , \new_[12842]_ , \new_[12843]_ , \new_[12844]_ ,
    \new_[12845]_ , \new_[12846]_ , \new_[12847]_ , \new_[12848]_ ,
    \new_[12849]_ , \new_[12850]_ , \new_[12851]_ , \new_[12852]_ ,
    \new_[12853]_ , \new_[12854]_ , \new_[12855]_ , \new_[12856]_ ,
    \new_[12857]_ , \new_[12858]_ , \new_[12859]_ , \new_[12860]_ ,
    \new_[12861]_ , \new_[12862]_ , \new_[12863]_ , \new_[12864]_ ,
    \new_[12865]_ , \new_[12866]_ , \new_[12867]_ , \new_[12868]_ ,
    \new_[12869]_ , \new_[12870]_ , \new_[12871]_ , \new_[12872]_ ,
    \new_[12873]_ , \new_[12874]_ , \new_[12875]_ , \new_[12876]_ ,
    \new_[12877]_ , \new_[12878]_ , \new_[12879]_ , \new_[12880]_ ,
    \new_[12881]_ , \new_[12882]_ , \new_[12883]_ , \new_[12884]_ ,
    \new_[12885]_ , \new_[12886]_ , \new_[12887]_ , \new_[12888]_ ,
    \new_[12889]_ , \new_[12890]_ , \new_[12891]_ , \new_[12892]_ ,
    \new_[12893]_ , \new_[12894]_ , \new_[12895]_ , \new_[12896]_ ,
    \new_[12897]_ , \new_[12898]_ , \new_[12899]_ , \new_[12900]_ ,
    \new_[12901]_ , \new_[12902]_ , \new_[12903]_ , \new_[12904]_ ,
    \new_[12905]_ , \new_[12906]_ , \new_[12907]_ , \new_[12908]_ ,
    \new_[12909]_ , \new_[12910]_ , \new_[12911]_ , \new_[12912]_ ,
    \new_[12913]_ , \new_[12914]_ , \new_[12915]_ , \new_[12916]_ ,
    \new_[12917]_ , \new_[12918]_ , \new_[12919]_ , \new_[12920]_ ,
    \new_[12921]_ , \new_[12922]_ , \new_[12923]_ , \new_[12924]_ ,
    \new_[12925]_ , \new_[12926]_ , \new_[12927]_ , \new_[12928]_ ,
    \new_[12929]_ , \new_[12930]_ , \new_[12931]_ , \new_[12932]_ ,
    \new_[12933]_ , \new_[12934]_ , \new_[12935]_ , \new_[12936]_ ,
    \new_[12937]_ , \new_[12938]_ , \new_[12939]_ , \new_[12940]_ ,
    \new_[12941]_ , \new_[12942]_ , \new_[12943]_ , \new_[12944]_ ,
    \new_[12945]_ , \new_[12946]_ , \new_[12947]_ , \new_[12948]_ ,
    \new_[12949]_ , \new_[12950]_ , \new_[12951]_ , \new_[12952]_ ,
    \new_[12953]_ , \new_[12954]_ , \new_[12955]_ , \new_[12956]_ ,
    \new_[12957]_ , \new_[12958]_ , \new_[12959]_ , \new_[12960]_ ,
    \new_[12961]_ , \new_[12962]_ , \new_[12963]_ , \new_[12964]_ ,
    \new_[12965]_ , \new_[12966]_ , \new_[12967]_ , \new_[12968]_ ,
    \new_[12969]_ , \new_[12970]_ , \new_[12971]_ , \new_[12972]_ ,
    \new_[12973]_ , \new_[12974]_ , \new_[12975]_ , \new_[12976]_ ,
    \new_[12977]_ , \new_[12978]_ , \new_[12979]_ , \new_[12980]_ ,
    \new_[12981]_ , \new_[12982]_ , \new_[12983]_ , \new_[12984]_ ,
    \new_[12985]_ , \new_[12986]_ , \new_[12987]_ , \new_[12988]_ ,
    \new_[12989]_ , \new_[12990]_ , \new_[12991]_ , \new_[12992]_ ,
    \new_[12993]_ , \new_[12994]_ , \new_[12995]_ , \new_[12996]_ ,
    \new_[12997]_ , \new_[12998]_ , \new_[12999]_ , \new_[13000]_ ,
    \new_[13001]_ , \new_[13002]_ , \new_[13003]_ , \new_[13004]_ ,
    \new_[13005]_ , \new_[13006]_ , \new_[13007]_ , \new_[13008]_ ,
    \new_[13009]_ , \new_[13010]_ , \new_[13011]_ , \new_[13012]_ ,
    \new_[13013]_ , \new_[13014]_ , \new_[13015]_ , \new_[13016]_ ,
    \new_[13017]_ , \new_[13018]_ , \new_[13019]_ , \new_[13020]_ ,
    \new_[13021]_ , \new_[13022]_ , \new_[13023]_ , \new_[13024]_ ,
    \new_[13025]_ , \new_[13026]_ , \new_[13027]_ , \new_[13028]_ ,
    \new_[13029]_ , \new_[13030]_ , \new_[13031]_ , \new_[13032]_ ,
    \new_[13033]_ , \new_[13034]_ , \new_[13035]_ , \new_[13036]_ ,
    \new_[13037]_ , \new_[13038]_ , \new_[13039]_ , \new_[13040]_ ,
    \new_[13041]_ , \new_[13042]_ , \new_[13043]_ , \new_[13044]_ ,
    \new_[13045]_ , \new_[13046]_ , \new_[13047]_ , \new_[13048]_ ,
    \new_[13049]_ , \new_[13050]_ , \new_[13051]_ , \new_[13052]_ ,
    \new_[13053]_ , \new_[13054]_ , \new_[13055]_ , \new_[13056]_ ,
    \new_[13057]_ , \new_[13058]_ , \new_[13059]_ , \new_[13060]_ ,
    \new_[13061]_ , \new_[13062]_ , \new_[13063]_ , \new_[13064]_ ,
    \new_[13065]_ , \new_[13066]_ , \new_[13067]_ , \new_[13068]_ ,
    \new_[13069]_ , \new_[13070]_ , \new_[13071]_ , \new_[13072]_ ,
    \new_[13073]_ , \new_[13074]_ , \new_[13075]_ , \new_[13076]_ ,
    \new_[13077]_ , \new_[13078]_ , \new_[13079]_ , \new_[13080]_ ,
    \new_[13081]_ , \new_[13082]_ , \new_[13083]_ , \new_[13084]_ ,
    \new_[13085]_ , \new_[13086]_ , \new_[13087]_ , \new_[13088]_ ,
    \new_[13089]_ , \new_[13090]_ , \new_[13091]_ , \new_[13092]_ ,
    \new_[13093]_ , \new_[13094]_ , \new_[13095]_ , \new_[13096]_ ,
    \new_[13097]_ , \new_[13098]_ , \new_[13099]_ , \new_[13100]_ ,
    \new_[13101]_ , \new_[13102]_ , \new_[13103]_ , \new_[13104]_ ,
    \new_[13105]_ , \new_[13106]_ , \new_[13107]_ , \new_[13108]_ ,
    \new_[13109]_ , \new_[13110]_ , \new_[13111]_ , \new_[13112]_ ,
    \new_[13113]_ , \new_[13114]_ , \new_[13115]_ , \new_[13116]_ ,
    \new_[13117]_ , \new_[13118]_ , \new_[13119]_ , \new_[13120]_ ,
    \new_[13121]_ , \new_[13122]_ , \new_[13123]_ , \new_[13124]_ ,
    \new_[13125]_ , \new_[13126]_ , \new_[13127]_ , \new_[13128]_ ,
    \new_[13129]_ , \new_[13130]_ , \new_[13131]_ , \new_[13132]_ ,
    \new_[13133]_ , \new_[13134]_ , \new_[13135]_ , \new_[13136]_ ,
    \new_[13137]_ , \new_[13138]_ , \new_[13139]_ , \new_[13140]_ ,
    \new_[13141]_ , \new_[13142]_ , \new_[13143]_ , \new_[13144]_ ,
    \new_[13145]_ , \new_[13146]_ , \new_[13147]_ , \new_[13148]_ ,
    \new_[13149]_ , \new_[13150]_ , \new_[13151]_ , \new_[13152]_ ,
    \new_[13153]_ , \new_[13154]_ , \new_[13155]_ , \new_[13156]_ ,
    \new_[13157]_ , \new_[13158]_ , \new_[13159]_ , \new_[13160]_ ,
    \new_[13161]_ , \new_[13162]_ , \new_[13163]_ , \new_[13164]_ ,
    \new_[13165]_ , \new_[13166]_ , \new_[13167]_ , \new_[13168]_ ,
    \new_[13169]_ , \new_[13170]_ , \new_[13171]_ , \new_[13172]_ ,
    \new_[13173]_ , \new_[13174]_ , \new_[13175]_ , \new_[13176]_ ,
    \new_[13177]_ , \new_[13178]_ , \new_[13179]_ , \new_[13180]_ ,
    \new_[13181]_ , \new_[13182]_ , \new_[13183]_ , \new_[13184]_ ,
    \new_[13185]_ , \new_[13186]_ , \new_[13187]_ , \new_[13188]_ ,
    \new_[13189]_ , \new_[13190]_ , \new_[13191]_ , \new_[13192]_ ,
    \new_[13193]_ , \new_[13194]_ , \new_[13195]_ , \new_[13196]_ ,
    \new_[13197]_ , \new_[13198]_ , \new_[13199]_ , \new_[13200]_ ,
    \new_[13201]_ , \new_[13202]_ , \new_[13203]_ , \new_[13204]_ ,
    \new_[13205]_ , \new_[13206]_ , \new_[13207]_ , \new_[13208]_ ,
    \new_[13209]_ , \new_[13210]_ , \new_[13211]_ , \new_[13212]_ ,
    \new_[13213]_ , \new_[13214]_ , \new_[13215]_ , \new_[13216]_ ,
    \new_[13217]_ , \new_[13218]_ , \new_[13219]_ , \new_[13220]_ ,
    \new_[13221]_ , \new_[13222]_ , \new_[13223]_ , \new_[13224]_ ,
    \new_[13225]_ , \new_[13226]_ , \new_[13227]_ , \new_[13228]_ ,
    \new_[13229]_ , \new_[13230]_ , \new_[13231]_ , \new_[13232]_ ,
    \new_[13233]_ , \new_[13234]_ , \new_[13235]_ , \new_[13236]_ ,
    \new_[13237]_ , \new_[13238]_ , \new_[13239]_ , \new_[13240]_ ,
    \new_[13241]_ , \new_[13242]_ , \new_[13243]_ , \new_[13244]_ ,
    \new_[13245]_ , \new_[13246]_ , \new_[13247]_ , \new_[13248]_ ,
    \new_[13249]_ , \new_[13250]_ , \new_[13251]_ , \new_[13252]_ ,
    \new_[13253]_ , \new_[13254]_ , \new_[13255]_ , \new_[13256]_ ,
    \new_[13257]_ , \new_[13258]_ , \new_[13259]_ , \new_[13260]_ ,
    \new_[13261]_ , \new_[13262]_ , \new_[13263]_ , \new_[13264]_ ,
    \new_[13265]_ , \new_[13266]_ , \new_[13267]_ , \new_[13268]_ ,
    \new_[13269]_ , \new_[13270]_ , \new_[13271]_ , \new_[13272]_ ,
    \new_[13273]_ , \new_[13274]_ , \new_[13275]_ , \new_[13276]_ ,
    \new_[13277]_ , \new_[13278]_ , \new_[13279]_ , \new_[13280]_ ,
    \new_[13281]_ , \new_[13282]_ , \new_[13283]_ , \new_[13284]_ ,
    \new_[13285]_ , \new_[13286]_ , \new_[13287]_ , \new_[13288]_ ,
    \new_[13289]_ , \new_[13290]_ , \new_[13291]_ , \new_[13292]_ ,
    \new_[13293]_ , \new_[13294]_ , \new_[13295]_ , \new_[13296]_ ,
    \new_[13297]_ , \new_[13298]_ , \new_[13299]_ , \new_[13300]_ ,
    \new_[13301]_ , \new_[13302]_ , \new_[13303]_ , \new_[13304]_ ,
    \new_[13305]_ , \new_[13306]_ , \new_[13307]_ , \new_[13308]_ ,
    \new_[13309]_ , \new_[13310]_ , \new_[13311]_ , \new_[13312]_ ,
    \new_[13313]_ , \new_[13314]_ , \new_[13315]_ , \new_[13316]_ ,
    \new_[13317]_ , \new_[13318]_ , \new_[13319]_ , \new_[13320]_ ,
    \new_[13321]_ , \new_[13322]_ , \new_[13323]_ , \new_[13324]_ ,
    \new_[13325]_ , \new_[13326]_ , \new_[13327]_ , \new_[13328]_ ,
    \new_[13329]_ , \new_[13330]_ , \new_[13331]_ , \new_[13332]_ ,
    \new_[13333]_ , \new_[13334]_ , \new_[13335]_ , \new_[13336]_ ,
    \new_[13337]_ , \new_[13338]_ , \new_[13339]_ , \new_[13340]_ ,
    \new_[13341]_ , \new_[13342]_ , \new_[13343]_ , \new_[13344]_ ,
    \new_[13345]_ , \new_[13346]_ , \new_[13347]_ , \new_[13348]_ ,
    \new_[13349]_ , \new_[13350]_ , \new_[13351]_ , \new_[13352]_ ,
    \new_[13353]_ , \new_[13354]_ , \new_[13355]_ , \new_[13356]_ ,
    \new_[13357]_ , \new_[13358]_ , \new_[13359]_ , \new_[13360]_ ,
    \new_[13361]_ , \new_[13362]_ , \new_[13363]_ , \new_[13364]_ ,
    \new_[13365]_ , \new_[13366]_ , \new_[13367]_ , \new_[13368]_ ,
    \new_[13369]_ , \new_[13370]_ , \new_[13371]_ , \new_[13372]_ ,
    \new_[13373]_ , \new_[13374]_ , \new_[13375]_ , \new_[13376]_ ,
    \new_[13377]_ , \new_[13378]_ , \new_[13379]_ , \new_[13380]_ ,
    \new_[13381]_ , \new_[13382]_ , \new_[13383]_ , \new_[13384]_ ,
    \new_[13385]_ , \new_[13386]_ , \new_[13387]_ , \new_[13388]_ ,
    \new_[13389]_ , \new_[13390]_ , \new_[13391]_ , \new_[13392]_ ,
    \new_[13393]_ , \new_[13394]_ , \new_[13395]_ , \new_[13396]_ ,
    \new_[13397]_ , \new_[13398]_ , \new_[13399]_ , \new_[13400]_ ,
    \new_[13401]_ , \new_[13402]_ , \new_[13403]_ , \new_[13404]_ ,
    \new_[13405]_ , \new_[13406]_ , \new_[13407]_ , \new_[13408]_ ,
    \new_[13409]_ , \new_[13410]_ , \new_[13411]_ , \new_[13412]_ ,
    \new_[13413]_ , \new_[13414]_ , \new_[13415]_ , \new_[13416]_ ,
    \new_[13417]_ , \new_[13418]_ , \new_[13419]_ , \new_[13420]_ ,
    \new_[13421]_ , \new_[13422]_ , \new_[13423]_ , \new_[13424]_ ,
    \new_[13425]_ , \new_[13426]_ , \new_[13427]_ , \new_[13428]_ ,
    \new_[13429]_ , \new_[13430]_ , \new_[13431]_ , \new_[13432]_ ,
    \new_[13433]_ , \new_[13434]_ , \new_[13435]_ , \new_[13436]_ ,
    \new_[13437]_ , \new_[13438]_ , \new_[13439]_ , \new_[13440]_ ,
    \new_[13441]_ , \new_[13442]_ , \new_[13443]_ , \new_[13444]_ ,
    \new_[13445]_ , \new_[13446]_ , \new_[13447]_ , \new_[13448]_ ,
    \new_[13449]_ , \new_[13450]_ , \new_[13451]_ , \new_[13452]_ ,
    \new_[13453]_ , \new_[13454]_ , \new_[13455]_ , \new_[13456]_ ,
    \new_[13457]_ , \new_[13458]_ , \new_[13459]_ , \new_[13460]_ ,
    \new_[13461]_ , \new_[13462]_ , \new_[13463]_ , \new_[13464]_ ,
    \new_[13465]_ , \new_[13466]_ , \new_[13467]_ , \new_[13468]_ ,
    \new_[13469]_ , \new_[13470]_ , \new_[13471]_ , \new_[13472]_ ,
    \new_[13473]_ , \new_[13474]_ , \new_[13475]_ , \new_[13477]_ ,
    \new_[13478]_ , \new_[13479]_ , \new_[13481]_ , \new_[13482]_ ,
    \new_[13483]_ , \new_[13484]_ , \new_[13485]_ , \new_[13486]_ ,
    \new_[13487]_ , \new_[13488]_ , \new_[13489]_ , \new_[13490]_ ,
    \new_[13491]_ , \new_[13492]_ , \new_[13493]_ , \new_[13494]_ ,
    \new_[13495]_ , \new_[13496]_ , \new_[13497]_ , \new_[13498]_ ,
    \new_[13499]_ , \new_[13500]_ , \new_[13501]_ , \new_[13502]_ ,
    \new_[13503]_ , \new_[13504]_ , \new_[13505]_ , \new_[13506]_ ,
    \new_[13507]_ , \new_[13508]_ , \new_[13509]_ , \new_[13510]_ ,
    \new_[13511]_ , \new_[13512]_ , \new_[13513]_ , \new_[13514]_ ,
    \new_[13516]_ , \new_[13517]_ , \new_[13518]_ , \new_[13520]_ ,
    \new_[13521]_ , \new_[13522]_ , \new_[13523]_ , \new_[13524]_ ,
    \new_[13525]_ , \new_[13526]_ , \new_[13527]_ , \new_[13528]_ ,
    \new_[13529]_ , \new_[13530]_ , \new_[13531]_ , \new_[13532]_ ,
    \new_[13533]_ , \new_[13534]_ , \new_[13535]_ , \new_[13536]_ ,
    \new_[13537]_ , \new_[13538]_ , \new_[13539]_ , \new_[13540]_ ,
    \new_[13541]_ , \new_[13542]_ , \new_[13543]_ , \new_[13544]_ ,
    \new_[13545]_ , \new_[13546]_ , \new_[13547]_ , \new_[13548]_ ,
    \new_[13549]_ , \new_[13550]_ , \new_[13551]_ , \new_[13552]_ ,
    \new_[13553]_ , \new_[13554]_ , \new_[13555]_ , \new_[13556]_ ,
    \new_[13557]_ , \new_[13558]_ , \new_[13559]_ , \new_[13560]_ ,
    \new_[13561]_ , \new_[13562]_ , \new_[13563]_ , \new_[13564]_ ,
    \new_[13565]_ , \new_[13566]_ , \new_[13567]_ , \new_[13568]_ ,
    \new_[13569]_ , \new_[13570]_ , \new_[13571]_ , \new_[13572]_ ,
    \new_[13573]_ , \new_[13574]_ , \new_[13575]_ , \new_[13576]_ ,
    \new_[13577]_ , \new_[13578]_ , \new_[13579]_ , \new_[13580]_ ,
    \new_[13581]_ , \new_[13582]_ , \new_[13583]_ , \new_[13584]_ ,
    \new_[13585]_ , \new_[13586]_ , \new_[13587]_ , \new_[13588]_ ,
    \new_[13589]_ , \new_[13590]_ , \new_[13591]_ , \new_[13592]_ ,
    \new_[13593]_ , \new_[13594]_ , \new_[13595]_ , \new_[13596]_ ,
    \new_[13598]_ , \new_[13599]_ , \new_[13600]_ , \new_[13601]_ ,
    \new_[13602]_ , \new_[13603]_ , \new_[13604]_ , \new_[13605]_ ,
    \new_[13606]_ , \new_[13607]_ , \new_[13608]_ , \new_[13609]_ ,
    \new_[13610]_ , \new_[13611]_ , \new_[13612]_ , \new_[13613]_ ,
    \new_[13614]_ , \new_[13615]_ , \new_[13616]_ , \new_[13617]_ ,
    \new_[13618]_ , \new_[13619]_ , \new_[13620]_ , \new_[13621]_ ,
    \new_[13622]_ , \new_[13623]_ , \new_[13624]_ , \new_[13625]_ ,
    \new_[13626]_ , \new_[13627]_ , \new_[13628]_ , \new_[13629]_ ,
    \new_[13630]_ , \new_[13631]_ , \new_[13632]_ , \new_[13633]_ ,
    \new_[13634]_ , \new_[13635]_ , \new_[13636]_ , \new_[13637]_ ,
    \new_[13638]_ , \new_[13639]_ , \new_[13640]_ , \new_[13641]_ ,
    \new_[13642]_ , \new_[13643]_ , \new_[13644]_ , \new_[13645]_ ,
    \new_[13646]_ , \new_[13647]_ , \new_[13648]_ , \new_[13649]_ ,
    \new_[13650]_ , \new_[13651]_ , \new_[13652]_ , \new_[13653]_ ,
    \new_[13654]_ , \new_[13655]_ , \new_[13656]_ , \new_[13657]_ ,
    \new_[13658]_ , \new_[13659]_ , \new_[13660]_ , \new_[13661]_ ,
    \new_[13662]_ , \new_[13663]_ , \new_[13664]_ , \new_[13665]_ ,
    \new_[13666]_ , \new_[13667]_ , \new_[13668]_ , \new_[13669]_ ,
    \new_[13670]_ , \new_[13671]_ , \new_[13672]_ , \new_[13673]_ ,
    \new_[13674]_ , \new_[13675]_ , \new_[13676]_ , \new_[13677]_ ,
    \new_[13678]_ , \new_[13679]_ , \new_[13680]_ , \new_[13681]_ ,
    \new_[13682]_ , \new_[13683]_ , \new_[13684]_ , \new_[13685]_ ,
    \new_[13686]_ , \new_[13687]_ , \new_[13688]_ , \new_[13689]_ ,
    \new_[13690]_ , \new_[13691]_ , \new_[13692]_ , \new_[13693]_ ,
    \new_[13694]_ , \new_[13695]_ , \new_[13696]_ , \new_[13697]_ ,
    \new_[13698]_ , \new_[13699]_ , \new_[13700]_ , \new_[13701]_ ,
    \new_[13702]_ , \new_[13703]_ , \new_[13704]_ , \new_[13705]_ ,
    \new_[13706]_ , \new_[13707]_ , \new_[13708]_ , \new_[13709]_ ,
    \new_[13710]_ , \new_[13711]_ , \new_[13712]_ , \new_[13713]_ ,
    \new_[13714]_ , \new_[13715]_ , \new_[13716]_ , \new_[13717]_ ,
    \new_[13718]_ , \new_[13719]_ , \new_[13720]_ , \new_[13721]_ ,
    \new_[13722]_ , \new_[13723]_ , \new_[13724]_ , \new_[13725]_ ,
    \new_[13726]_ , \new_[13727]_ , \new_[13728]_ , \new_[13729]_ ,
    \new_[13730]_ , \new_[13731]_ , \new_[13732]_ , \new_[13733]_ ,
    \new_[13734]_ , \new_[13735]_ , \new_[13736]_ , \new_[13737]_ ,
    \new_[13738]_ , \new_[13739]_ , \new_[13740]_ , \new_[13741]_ ,
    \new_[13742]_ , \new_[13743]_ , \new_[13744]_ , \new_[13745]_ ,
    \new_[13746]_ , \new_[13747]_ , \new_[13748]_ , \new_[13749]_ ,
    \new_[13750]_ , \new_[13751]_ , \new_[13752]_ , \new_[13753]_ ,
    \new_[13754]_ , \new_[13755]_ , \new_[13756]_ , \new_[13757]_ ,
    \new_[13758]_ , \new_[13759]_ , \new_[13760]_ , \new_[13761]_ ,
    \new_[13762]_ , \new_[13763]_ , \new_[13764]_ , \new_[13765]_ ,
    \new_[13766]_ , \new_[13767]_ , \new_[13768]_ , \new_[13769]_ ,
    \new_[13770]_ , \new_[13771]_ , \new_[13772]_ , \new_[13773]_ ,
    \new_[13774]_ , \new_[13775]_ , \new_[13776]_ , \new_[13777]_ ,
    \new_[13778]_ , \new_[13779]_ , \new_[13780]_ , \new_[13781]_ ,
    \new_[13782]_ , \new_[13783]_ , \new_[13784]_ , \new_[13785]_ ,
    \new_[13786]_ , \new_[13787]_ , \new_[13788]_ , \new_[13789]_ ,
    \new_[13790]_ , \new_[13791]_ , \new_[13792]_ , \new_[13793]_ ,
    \new_[13794]_ , \new_[13795]_ , \new_[13796]_ , \new_[13797]_ ,
    \new_[13798]_ , \new_[13799]_ , \new_[13800]_ , \new_[13801]_ ,
    \new_[13802]_ , \new_[13803]_ , \new_[13804]_ , \new_[13805]_ ,
    \new_[13806]_ , \new_[13807]_ , \new_[13808]_ , \new_[13809]_ ,
    \new_[13810]_ , \new_[13811]_ , \new_[13812]_ , \new_[13813]_ ,
    \new_[13814]_ , \new_[13815]_ , \new_[13816]_ , \new_[13817]_ ,
    \new_[13818]_ , \new_[13819]_ , \new_[13820]_ , \new_[13821]_ ,
    \new_[13822]_ , \new_[13823]_ , \new_[13824]_ , \new_[13825]_ ,
    \new_[13826]_ , \new_[13827]_ , \new_[13828]_ , \new_[13829]_ ,
    \new_[13830]_ , \new_[13831]_ , \new_[13832]_ , \new_[13833]_ ,
    \new_[13834]_ , \new_[13835]_ , \new_[13836]_ , \new_[13837]_ ,
    \new_[13838]_ , \new_[13839]_ , \new_[13840]_ , \new_[13841]_ ,
    \new_[13842]_ , \new_[13843]_ , \new_[13844]_ , \new_[13845]_ ,
    \new_[13846]_ , \new_[13847]_ , \new_[13848]_ , \new_[13849]_ ,
    \new_[13850]_ , \new_[13851]_ , \new_[13852]_ , \new_[13853]_ ,
    \new_[13854]_ , \new_[13855]_ , \new_[13856]_ , \new_[13857]_ ,
    \new_[13858]_ , \new_[13859]_ , \new_[13860]_ , \new_[13861]_ ,
    \new_[13862]_ , \new_[13863]_ , \new_[13864]_ , \new_[13865]_ ,
    \new_[13866]_ , \new_[13867]_ , \new_[13868]_ , \new_[13869]_ ,
    \new_[13870]_ , \new_[13871]_ , \new_[13872]_ , \new_[13873]_ ,
    \new_[13874]_ , \new_[13875]_ , \new_[13876]_ , \new_[13877]_ ,
    \new_[13878]_ , \new_[13879]_ , \new_[13880]_ , \new_[13881]_ ,
    \new_[13882]_ , \new_[13883]_ , \new_[13884]_ , \new_[13885]_ ,
    \new_[13886]_ , \new_[13887]_ , \new_[13888]_ , \new_[13889]_ ,
    \new_[13890]_ , \new_[13891]_ , \new_[13892]_ , \new_[13893]_ ,
    \new_[13894]_ , \new_[13895]_ , \new_[13896]_ , \new_[13897]_ ,
    \new_[13898]_ , \new_[13899]_ , \new_[13900]_ , \new_[13901]_ ,
    \new_[13902]_ , \new_[13903]_ , \new_[13904]_ , \new_[13905]_ ,
    \new_[13906]_ , \new_[13907]_ , \new_[13908]_ , \new_[13909]_ ,
    \new_[13910]_ , \new_[13911]_ , \new_[13912]_ , \new_[13913]_ ,
    \new_[13914]_ , \new_[13915]_ , \new_[13916]_ , \new_[13917]_ ,
    \new_[13918]_ , \new_[13919]_ , \new_[13920]_ , \new_[13921]_ ,
    \new_[13922]_ , \new_[13923]_ , \new_[13924]_ , \new_[13925]_ ,
    \new_[13926]_ , \new_[13927]_ , \new_[13928]_ , \new_[13929]_ ,
    \new_[13930]_ , \new_[13931]_ , \new_[13932]_ , \new_[13933]_ ,
    \new_[13934]_ , \new_[13935]_ , \new_[13936]_ , \new_[13937]_ ,
    \new_[13938]_ , \new_[13939]_ , \new_[13940]_ , \new_[13941]_ ,
    \new_[13942]_ , \new_[13943]_ , \new_[13944]_ , \new_[13945]_ ,
    \new_[13946]_ , \new_[13947]_ , \new_[13948]_ , \new_[13949]_ ,
    \new_[13950]_ , \new_[13951]_ , \new_[13952]_ , \new_[13953]_ ,
    \new_[13954]_ , \new_[13955]_ , \new_[13956]_ , \new_[13957]_ ,
    \new_[13958]_ , \new_[13959]_ , \new_[13960]_ , \new_[13961]_ ,
    \new_[13962]_ , \new_[13963]_ , \new_[13964]_ , \new_[13965]_ ,
    \new_[13966]_ , \new_[13967]_ , \new_[13968]_ , \new_[13969]_ ,
    \new_[13970]_ , \new_[13971]_ , \new_[13972]_ , \new_[13973]_ ,
    \new_[13974]_ , \new_[13975]_ , \new_[13976]_ , \new_[13977]_ ,
    \new_[13978]_ , \new_[13979]_ , \new_[13980]_ , \new_[13981]_ ,
    \new_[13982]_ , \new_[13983]_ , \new_[13984]_ , \new_[13985]_ ,
    \new_[13986]_ , \new_[13987]_ , \new_[13988]_ , \new_[13989]_ ,
    \new_[13990]_ , \new_[13991]_ , \new_[13992]_ , \new_[13993]_ ,
    \new_[13994]_ , \new_[13995]_ , \new_[13996]_ , \new_[13997]_ ,
    \new_[13998]_ , \new_[13999]_ , \new_[14000]_ , \new_[14001]_ ,
    \new_[14002]_ , \new_[14003]_ , \new_[14004]_ , \new_[14005]_ ,
    \new_[14006]_ , \new_[14007]_ , \new_[14008]_ , \new_[14009]_ ,
    \new_[14010]_ , \new_[14011]_ , \new_[14012]_ , \new_[14013]_ ,
    \new_[14014]_ , \new_[14015]_ , \new_[14016]_ , \new_[14017]_ ,
    \new_[14018]_ , \new_[14019]_ , \new_[14020]_ , \new_[14021]_ ,
    \new_[14022]_ , \new_[14023]_ , \new_[14024]_ , \new_[14025]_ ,
    \new_[14026]_ , \new_[14027]_ , \new_[14028]_ , \new_[14029]_ ,
    \new_[14030]_ , \new_[14031]_ , \new_[14032]_ , \new_[14033]_ ,
    \new_[14034]_ , \new_[14035]_ , \new_[14036]_ , \new_[14037]_ ,
    \new_[14038]_ , \new_[14039]_ , \new_[14040]_ , \new_[14041]_ ,
    \new_[14042]_ , \new_[14043]_ , \new_[14044]_ , \new_[14045]_ ,
    \new_[14046]_ , \new_[14047]_ , \new_[14048]_ , \new_[14049]_ ,
    \new_[14050]_ , \new_[14051]_ , \new_[14052]_ , \new_[14053]_ ,
    \new_[14054]_ , \new_[14055]_ , \new_[14056]_ , \new_[14057]_ ,
    \new_[14058]_ , \new_[14059]_ , \new_[14060]_ , \new_[14061]_ ,
    \new_[14062]_ , \new_[14063]_ , \new_[14064]_ , \new_[14065]_ ,
    \new_[14066]_ , \new_[14067]_ , \new_[14068]_ , \new_[14069]_ ,
    \new_[14070]_ , \new_[14071]_ , \new_[14072]_ , \new_[14073]_ ,
    \new_[14074]_ , \new_[14075]_ , \new_[14076]_ , \new_[14077]_ ,
    \new_[14078]_ , \new_[14079]_ , \new_[14080]_ , \new_[14081]_ ,
    \new_[14082]_ , \new_[14083]_ , \new_[14084]_ , \new_[14085]_ ,
    \new_[14086]_ , \new_[14087]_ , \new_[14088]_ , \new_[14089]_ ,
    \new_[14090]_ , \new_[14091]_ , \new_[14092]_ , \new_[14093]_ ,
    \new_[14094]_ , \new_[14095]_ , \new_[14096]_ , \new_[14097]_ ,
    \new_[14098]_ , \new_[14099]_ , \new_[14100]_ , \new_[14101]_ ,
    \new_[14102]_ , \new_[14103]_ , \new_[14104]_ , \new_[14105]_ ,
    \new_[14106]_ , \new_[14107]_ , \new_[14108]_ , \new_[14109]_ ,
    \new_[14110]_ , \new_[14111]_ , \new_[14112]_ , \new_[14113]_ ,
    \new_[14114]_ , \new_[14115]_ , \new_[14116]_ , \new_[14117]_ ,
    \new_[14118]_ , \new_[14119]_ , \new_[14120]_ , \new_[14121]_ ,
    \new_[14122]_ , \new_[14123]_ , \new_[14124]_ , \new_[14125]_ ,
    \new_[14126]_ , \new_[14127]_ , \new_[14128]_ , \new_[14129]_ ,
    \new_[14130]_ , \new_[14131]_ , \new_[14132]_ , \new_[14133]_ ,
    \new_[14134]_ , \new_[14135]_ , \new_[14136]_ , \new_[14137]_ ,
    \new_[14138]_ , \new_[14139]_ , \new_[14140]_ , \new_[14141]_ ,
    \new_[14142]_ , \new_[14143]_ , \new_[14144]_ , \new_[14145]_ ,
    \new_[14146]_ , \new_[14147]_ , \new_[14148]_ , \new_[14149]_ ,
    \new_[14150]_ , \new_[14151]_ , \new_[14152]_ , \new_[14153]_ ,
    \new_[14154]_ , \new_[14155]_ , \new_[14156]_ , \new_[14157]_ ,
    \new_[14158]_ , \new_[14159]_ , \new_[14160]_ , \new_[14161]_ ,
    \new_[14162]_ , \new_[14163]_ , \new_[14164]_ , \new_[14165]_ ,
    \new_[14166]_ , \new_[14167]_ , \new_[14168]_ , \new_[14169]_ ,
    \new_[14170]_ , \new_[14171]_ , \new_[14172]_ , \new_[14173]_ ,
    \new_[14174]_ , \new_[14175]_ , \new_[14176]_ , \new_[14177]_ ,
    \new_[14178]_ , \new_[14179]_ , \new_[14180]_ , \new_[14181]_ ,
    \new_[14182]_ , \new_[14183]_ , \new_[14184]_ , \new_[14185]_ ,
    \new_[14186]_ , \new_[14187]_ , \new_[14188]_ , \new_[14189]_ ,
    \new_[14190]_ , \new_[14191]_ , \new_[14192]_ , \new_[14193]_ ,
    \new_[14194]_ , \new_[14195]_ , \new_[14196]_ , \new_[14197]_ ,
    \new_[14198]_ , \new_[14199]_ , \new_[14200]_ , \new_[14201]_ ,
    \new_[14202]_ , \new_[14203]_ , \new_[14204]_ , \new_[14205]_ ,
    \new_[14206]_ , \new_[14207]_ , \new_[14208]_ , \new_[14209]_ ,
    \new_[14210]_ , \new_[14211]_ , \new_[14212]_ , \new_[14213]_ ,
    \new_[14214]_ , \new_[14215]_ , \new_[14216]_ , \new_[14217]_ ,
    \new_[14218]_ , \new_[14219]_ , \new_[14220]_ , \new_[14221]_ ,
    \new_[14222]_ , \new_[14223]_ , \new_[14224]_ , \new_[14225]_ ,
    \new_[14226]_ , \new_[14227]_ , \new_[14228]_ , \new_[14229]_ ,
    \new_[14230]_ , \new_[14231]_ , \new_[14232]_ , \new_[14233]_ ,
    \new_[14234]_ , \new_[14235]_ , \new_[14236]_ , \new_[14237]_ ,
    \new_[14238]_ , \new_[14239]_ , \new_[14240]_ , \new_[14241]_ ,
    \new_[14242]_ , \new_[14243]_ , \new_[14244]_ , \new_[14245]_ ,
    \new_[14246]_ , \new_[14247]_ , \new_[14248]_ , \new_[14249]_ ,
    \new_[14250]_ , \new_[14251]_ , \new_[14252]_ , \new_[14253]_ ,
    \new_[14254]_ , \new_[14255]_ , \new_[14256]_ , \new_[14257]_ ,
    \new_[14258]_ , \new_[14259]_ , \new_[14260]_ , \new_[14261]_ ,
    \new_[14262]_ , \new_[14263]_ , \new_[14264]_ , \new_[14265]_ ,
    \new_[14266]_ , \new_[14267]_ , \new_[14268]_ , \new_[14269]_ ,
    \new_[14270]_ , \new_[14271]_ , \new_[14272]_ , \new_[14273]_ ,
    \new_[14274]_ , \new_[14275]_ , \new_[14276]_ , \new_[14277]_ ,
    \new_[14278]_ , \new_[14279]_ , \new_[14280]_ , \new_[14281]_ ,
    \new_[14282]_ , \new_[14283]_ , \new_[14284]_ , \new_[14285]_ ,
    \new_[14286]_ , \new_[14287]_ , \new_[14288]_ , \new_[14289]_ ,
    \new_[14290]_ , \new_[14291]_ , \new_[14292]_ , \new_[14293]_ ,
    \new_[14294]_ , \new_[14295]_ , \new_[14296]_ , \new_[14297]_ ,
    \new_[14298]_ , \new_[14299]_ , \new_[14300]_ , \new_[14301]_ ,
    \new_[14302]_ , \new_[14303]_ , \new_[14304]_ , \new_[14305]_ ,
    \new_[14306]_ , \new_[14307]_ , \new_[14308]_ , \new_[14309]_ ,
    \new_[14310]_ , \new_[14311]_ , \new_[14312]_ , \new_[14313]_ ,
    \new_[14314]_ , \new_[14315]_ , \new_[14316]_ , \new_[14317]_ ,
    \new_[14318]_ , \new_[14319]_ , \new_[14320]_ , \new_[14321]_ ,
    \new_[14322]_ , \new_[14323]_ , \new_[14324]_ , \new_[14325]_ ,
    \new_[14326]_ , \new_[14327]_ , \new_[14328]_ , \new_[14329]_ ,
    \new_[14330]_ , \new_[14331]_ , \new_[14332]_ , \new_[14333]_ ,
    \new_[14334]_ , \new_[14335]_ , \new_[14336]_ , \new_[14337]_ ,
    \new_[14338]_ , \new_[14339]_ , \new_[14340]_ , \new_[14341]_ ,
    \new_[14342]_ , \new_[14343]_ , \new_[14344]_ , \new_[14345]_ ,
    \new_[14346]_ , \new_[14347]_ , \new_[14348]_ , \new_[14349]_ ,
    \new_[14350]_ , \new_[14351]_ , \new_[14352]_ , \new_[14353]_ ,
    \new_[14354]_ , \new_[14355]_ , \new_[14356]_ , \new_[14357]_ ,
    \new_[14358]_ , \new_[14359]_ , \new_[14360]_ , \new_[14361]_ ,
    \new_[14362]_ , \new_[14363]_ , \new_[14364]_ , \new_[14365]_ ,
    \new_[14366]_ , \new_[14367]_ , \new_[14368]_ , \new_[14369]_ ,
    \new_[14370]_ , \new_[14371]_ , \new_[14372]_ , \new_[14373]_ ,
    \new_[14374]_ , \new_[14375]_ , \new_[14376]_ , \new_[14377]_ ,
    \new_[14378]_ , \new_[14379]_ , \new_[14380]_ , \new_[14381]_ ,
    \new_[14382]_ , \new_[14383]_ , \new_[14384]_ , \new_[14385]_ ,
    \new_[14386]_ , \new_[14387]_ , \new_[14388]_ , \new_[14389]_ ,
    \new_[14390]_ , \new_[14391]_ , \new_[14392]_ , \new_[14393]_ ,
    \new_[14394]_ , \new_[14395]_ , \new_[14396]_ , \new_[14397]_ ,
    \new_[14398]_ , \new_[14399]_ , \new_[14400]_ , \new_[14401]_ ,
    \new_[14402]_ , \new_[14403]_ , \new_[14404]_ , \new_[14405]_ ,
    \new_[14406]_ , \new_[14407]_ , \new_[14408]_ , \new_[14409]_ ,
    \new_[14410]_ , \new_[14411]_ , \new_[14412]_ , \new_[14413]_ ,
    \new_[14414]_ , \new_[14415]_ , \new_[14416]_ , \new_[14417]_ ,
    \new_[14418]_ , \new_[14419]_ , \new_[14420]_ , \new_[14421]_ ,
    \new_[14422]_ , \new_[14423]_ , \new_[14424]_ , \new_[14425]_ ,
    \new_[14426]_ , \new_[14427]_ , \new_[14428]_ , \new_[14429]_ ,
    \new_[14430]_ , \new_[14431]_ , \new_[14432]_ , \new_[14433]_ ,
    \new_[14434]_ , \new_[14435]_ , \new_[14436]_ , \new_[14437]_ ,
    \new_[14438]_ , \new_[14439]_ , \new_[14440]_ , \new_[14441]_ ,
    \new_[14442]_ , \new_[14443]_ , \new_[14444]_ , \new_[14445]_ ,
    \new_[14446]_ , \new_[14447]_ , \new_[14448]_ , \new_[14449]_ ,
    \new_[14450]_ , \new_[14451]_ , \new_[14452]_ , \new_[14453]_ ,
    \new_[14454]_ , \new_[14455]_ , \new_[14456]_ , \new_[14457]_ ,
    \new_[14458]_ , \new_[14459]_ , \new_[14460]_ , \new_[14461]_ ,
    \new_[14462]_ , \new_[14463]_ , \new_[14464]_ , \new_[14465]_ ,
    \new_[14466]_ , \new_[14467]_ , \new_[14468]_ , \new_[14469]_ ,
    \new_[14470]_ , \new_[14471]_ , \new_[14472]_ , \new_[14473]_ ,
    \new_[14474]_ , \new_[14475]_ , \new_[14476]_ , \new_[14477]_ ,
    \new_[14478]_ , \new_[14479]_ , \new_[14480]_ , \new_[14481]_ ,
    \new_[14482]_ , \new_[14483]_ , \new_[14484]_ , \new_[14485]_ ,
    \new_[14486]_ , \new_[14487]_ , \new_[14488]_ , \new_[14489]_ ,
    \new_[14490]_ , \new_[14491]_ , \new_[14492]_ , \new_[14493]_ ,
    \new_[14494]_ , \new_[14495]_ , \new_[14496]_ , \new_[14497]_ ,
    \new_[14498]_ , \new_[14499]_ , \new_[14500]_ , \new_[14501]_ ,
    \new_[14502]_ , \new_[14503]_ , \new_[14504]_ , \new_[14505]_ ,
    \new_[14506]_ , \new_[14507]_ , \new_[14508]_ , \new_[14509]_ ,
    \new_[14510]_ , \new_[14511]_ , \new_[14512]_ , \new_[14513]_ ,
    \new_[14514]_ , \new_[14515]_ , \new_[14516]_ , \new_[14517]_ ,
    \new_[14518]_ , \new_[14519]_ , \new_[14520]_ , \new_[14521]_ ,
    \new_[14522]_ , \new_[14523]_ , \new_[14524]_ , \new_[14525]_ ,
    \new_[14526]_ , \new_[14527]_ , \new_[14528]_ , \new_[14529]_ ,
    \new_[14530]_ , \new_[14531]_ , \new_[14532]_ , \new_[14533]_ ,
    \new_[14534]_ , \new_[14535]_ , \new_[14536]_ , \new_[14537]_ ,
    \new_[14538]_ , \new_[14539]_ , \new_[14540]_ , \new_[14541]_ ,
    \new_[14542]_ , \new_[14543]_ , \new_[14544]_ , \new_[14545]_ ,
    \new_[14546]_ , \new_[14547]_ , \new_[14548]_ , \new_[14549]_ ,
    \new_[14550]_ , \new_[14551]_ , \new_[14552]_ , \new_[14553]_ ,
    \new_[14554]_ , \new_[14555]_ , \new_[14556]_ , \new_[14557]_ ,
    \new_[14558]_ , \new_[14559]_ , \new_[14560]_ , \new_[14561]_ ,
    \new_[14562]_ , \new_[14563]_ , \new_[14564]_ , \new_[14565]_ ,
    \new_[14566]_ , \new_[14567]_ , \new_[14568]_ , \new_[14569]_ ,
    \new_[14570]_ , \new_[14571]_ , \new_[14572]_ , \new_[14573]_ ,
    \new_[14574]_ , \new_[14575]_ , \new_[14576]_ , \new_[14577]_ ,
    \new_[14578]_ , \new_[14579]_ , \new_[14580]_ , \new_[14581]_ ,
    \new_[14582]_ , \new_[14583]_ , \new_[14584]_ , \new_[14585]_ ,
    \new_[14586]_ , \new_[14587]_ , \new_[14588]_ , \new_[14589]_ ,
    \new_[14590]_ , \new_[14591]_ , \new_[14592]_ , \new_[14593]_ ,
    \new_[14594]_ , \new_[14595]_ , \new_[14596]_ , \new_[14597]_ ,
    \new_[14598]_ , \new_[14599]_ , \new_[14600]_ , \new_[14601]_ ,
    \new_[14602]_ , \new_[14603]_ , \new_[14604]_ , \new_[14605]_ ,
    \new_[14606]_ , \new_[14607]_ , \new_[14608]_ , \new_[14609]_ ,
    \new_[14610]_ , \new_[14611]_ , \new_[14612]_ , \new_[14613]_ ,
    \new_[14614]_ , \new_[14615]_ , \new_[14616]_ , \new_[14617]_ ,
    \new_[14618]_ , \new_[14619]_ , \new_[14620]_ , \new_[14621]_ ,
    \new_[14622]_ , \new_[14623]_ , \new_[14624]_ , \new_[14625]_ ,
    \new_[14626]_ , \new_[14627]_ , \new_[14628]_ , \new_[14629]_ ,
    \new_[14630]_ , \new_[14631]_ , \new_[14632]_ , \new_[14633]_ ,
    \new_[14634]_ , \new_[14635]_ , \new_[14636]_ , \new_[14637]_ ,
    \new_[14638]_ , \new_[14639]_ , \new_[14640]_ , \new_[14642]_ ,
    \new_[14643]_ , \new_[14644]_ , \new_[14645]_ , \new_[14646]_ ,
    \new_[14647]_ , \new_[14648]_ , \new_[14649]_ , \new_[14650]_ ,
    \new_[14651]_ , \new_[14652]_ , \new_[14653]_ , \new_[14654]_ ,
    \new_[14655]_ , \new_[14656]_ , \new_[14657]_ , \new_[14658]_ ,
    \new_[14659]_ , \new_[14660]_ , \new_[14661]_ , \new_[14662]_ ,
    \new_[14663]_ , \new_[14664]_ , \new_[14665]_ , \new_[14666]_ ,
    \new_[14667]_ , \new_[14668]_ , \new_[14669]_ , \new_[14670]_ ,
    \new_[14671]_ , \new_[14672]_ , \new_[14673]_ , \new_[14674]_ ,
    \new_[14675]_ , \new_[14676]_ , \new_[14677]_ , \new_[14678]_ ,
    \new_[14679]_ , \new_[14680]_ , \new_[14681]_ , \new_[14682]_ ,
    \new_[14683]_ , \new_[14684]_ , \new_[14685]_ , \new_[14686]_ ,
    \new_[14687]_ , \new_[14688]_ , \new_[14689]_ , \new_[14690]_ ,
    \new_[14691]_ , \new_[14692]_ , \new_[14693]_ , \new_[14694]_ ,
    \new_[14695]_ , \new_[14696]_ , \new_[14697]_ , \new_[14698]_ ,
    \new_[14699]_ , \new_[14700]_ , \new_[14701]_ , \new_[14702]_ ,
    \new_[14703]_ , \new_[14704]_ , \new_[14705]_ , \new_[14706]_ ,
    \new_[14707]_ , \new_[14708]_ , \new_[14709]_ , \new_[14710]_ ,
    \new_[14711]_ , \new_[14712]_ , \new_[14713]_ , \new_[14714]_ ,
    \new_[14715]_ , \new_[14716]_ , \new_[14717]_ , \new_[14718]_ ,
    \new_[14719]_ , \new_[14720]_ , \new_[14721]_ , \new_[14722]_ ,
    \new_[14723]_ , \new_[14724]_ , \new_[14725]_ , \new_[14726]_ ,
    \new_[14727]_ , \new_[14728]_ , \new_[14729]_ , \new_[14730]_ ,
    \new_[14731]_ , \new_[14732]_ , \new_[14733]_ , \new_[14734]_ ,
    \new_[14735]_ , \new_[14736]_ , \new_[14737]_ , \new_[14738]_ ,
    \new_[14739]_ , \new_[14740]_ , \new_[14741]_ , \new_[14742]_ ,
    \new_[14743]_ , \new_[14744]_ , \new_[14745]_ , \new_[14746]_ ,
    \new_[14747]_ , \new_[14748]_ , \new_[14749]_ , \new_[14750]_ ,
    \new_[14751]_ , \new_[14752]_ , \new_[14753]_ , \new_[14754]_ ,
    \new_[14755]_ , \new_[14756]_ , \new_[14757]_ , \new_[14758]_ ,
    \new_[14759]_ , \new_[14760]_ , \new_[14761]_ , \new_[14762]_ ,
    \new_[14763]_ , \new_[14764]_ , \new_[14765]_ , \new_[14766]_ ,
    \new_[14767]_ , \new_[14768]_ , \new_[14769]_ , \new_[14770]_ ,
    \new_[14771]_ , \new_[14772]_ , \new_[14773]_ , \new_[14774]_ ,
    \new_[14775]_ , \new_[14776]_ , \new_[14777]_ , \new_[14778]_ ,
    \new_[14779]_ , \new_[14780]_ , \new_[14781]_ , \new_[14782]_ ,
    \new_[14783]_ , \new_[14784]_ , \new_[14785]_ , \new_[14786]_ ,
    \new_[14787]_ , \new_[14788]_ , \new_[14789]_ , \new_[14790]_ ,
    \new_[14791]_ , \new_[14792]_ , \new_[14793]_ , \new_[14794]_ ,
    \new_[14795]_ , \new_[14796]_ , \new_[14797]_ , \new_[14798]_ ,
    \new_[14799]_ , \new_[14800]_ , \new_[14801]_ , \new_[14802]_ ,
    \new_[14803]_ , \new_[14804]_ , \new_[14805]_ , \new_[14806]_ ,
    \new_[14807]_ , \new_[14808]_ , \new_[14809]_ , \new_[14810]_ ,
    \new_[14811]_ , \new_[14812]_ , \new_[14813]_ , \new_[14814]_ ,
    \new_[14815]_ , \new_[14816]_ , \new_[14817]_ , \new_[14818]_ ,
    \new_[14819]_ , \new_[14820]_ , \new_[14821]_ , \new_[14822]_ ,
    \new_[14823]_ , \new_[14824]_ , \new_[14825]_ , \new_[14826]_ ,
    \new_[14827]_ , \new_[14828]_ , \new_[14829]_ , \new_[14830]_ ,
    \new_[14831]_ , \new_[14832]_ , \new_[14833]_ , \new_[14834]_ ,
    \new_[14835]_ , \new_[14836]_ , \new_[14837]_ , \new_[14838]_ ,
    \new_[14839]_ , \new_[14840]_ , \new_[14841]_ , \new_[14842]_ ,
    \new_[14843]_ , \new_[14844]_ , \new_[14845]_ , \new_[14846]_ ,
    \new_[14847]_ , \new_[14848]_ , \new_[14849]_ , \new_[14850]_ ,
    \new_[14851]_ , \new_[14852]_ , \new_[14853]_ , \new_[14854]_ ,
    \new_[14855]_ , \new_[14856]_ , \new_[14857]_ , \new_[14858]_ ,
    \new_[14859]_ , \new_[14860]_ , \new_[14861]_ , \new_[14862]_ ,
    \new_[14863]_ , \new_[14864]_ , \new_[14865]_ , \new_[14866]_ ,
    \new_[14867]_ , \new_[14868]_ , \new_[14869]_ , \new_[14870]_ ,
    \new_[14871]_ , \new_[14872]_ , \new_[14873]_ , \new_[14874]_ ,
    \new_[14875]_ , \new_[14876]_ , \new_[14877]_ , \new_[14878]_ ,
    \new_[14879]_ , \new_[14880]_ , \new_[14881]_ , \new_[14882]_ ,
    \new_[14883]_ , \new_[14884]_ , \new_[14885]_ , \new_[14886]_ ,
    \new_[14887]_ , \new_[14888]_ , \new_[14889]_ , \new_[14890]_ ,
    \new_[14891]_ , \new_[14892]_ , \new_[14893]_ , \new_[14894]_ ,
    \new_[14895]_ , \new_[14896]_ , \new_[14897]_ , \new_[14898]_ ,
    \new_[14899]_ , \new_[14900]_ , \new_[14901]_ , \new_[14902]_ ,
    \new_[14903]_ , \new_[14904]_ , \new_[14905]_ , \new_[14906]_ ,
    \new_[14907]_ , \new_[14908]_ , \new_[14909]_ , \new_[14910]_ ,
    \new_[14911]_ , \new_[14912]_ , \new_[14913]_ , \new_[14914]_ ,
    \new_[14915]_ , \new_[14916]_ , \new_[14917]_ , \new_[14918]_ ,
    \new_[14919]_ , \new_[14920]_ , \new_[14921]_ , \new_[14922]_ ,
    \new_[14923]_ , \new_[14924]_ , \new_[14925]_ , \new_[14926]_ ,
    \new_[14927]_ , \new_[14928]_ , \new_[14929]_ , \new_[14930]_ ,
    \new_[14931]_ , \new_[14932]_ , \new_[14933]_ , \new_[14934]_ ,
    \new_[14935]_ , \new_[14936]_ , \new_[14937]_ , \new_[14938]_ ,
    \new_[14939]_ , \new_[14940]_ , \new_[14941]_ , \new_[14942]_ ,
    \new_[14943]_ , \new_[14944]_ , \new_[14945]_ , \new_[14946]_ ,
    \new_[14947]_ , \new_[14948]_ , \new_[14949]_ , \new_[14950]_ ,
    \new_[14951]_ , \new_[14952]_ , \new_[14953]_ , \new_[14954]_ ,
    \new_[14955]_ , \new_[14956]_ , \new_[14957]_ , \new_[14958]_ ,
    \new_[14959]_ , \new_[14960]_ , \new_[14961]_ , \new_[14962]_ ,
    \new_[14963]_ , \new_[14964]_ , \new_[14965]_ , \new_[14966]_ ,
    \new_[14967]_ , \new_[14968]_ , \new_[14969]_ , \new_[14970]_ ,
    \new_[14971]_ , \new_[14972]_ , \new_[14973]_ , \new_[14974]_ ,
    \new_[14975]_ , \new_[14976]_ , \new_[14977]_ , \new_[14978]_ ,
    \new_[14979]_ , \new_[14980]_ , \new_[14981]_ , \new_[14982]_ ,
    \new_[14983]_ , \new_[14984]_ , \new_[14985]_ , \new_[14986]_ ,
    \new_[14987]_ , \new_[14988]_ , \new_[14989]_ , \new_[14990]_ ,
    \new_[14991]_ , \new_[14992]_ , \new_[14993]_ , \new_[14994]_ ,
    \new_[14995]_ , \new_[14996]_ , \new_[14997]_ , \new_[14998]_ ,
    \new_[14999]_ , \new_[15000]_ , \new_[15001]_ , \new_[15002]_ ,
    \new_[15003]_ , \new_[15004]_ , \new_[15005]_ , \new_[15006]_ ,
    \new_[15007]_ , \new_[15008]_ , \new_[15009]_ , \new_[15010]_ ,
    \new_[15011]_ , \new_[15012]_ , \new_[15013]_ , \new_[15014]_ ,
    \new_[15015]_ , \new_[15016]_ , \new_[15017]_ , \new_[15018]_ ,
    \new_[15019]_ , \new_[15020]_ , \new_[15021]_ , \new_[15022]_ ,
    \new_[15023]_ , \new_[15024]_ , \new_[15025]_ , \new_[15026]_ ,
    \new_[15027]_ , \new_[15028]_ , \new_[15029]_ , \new_[15030]_ ,
    \new_[15031]_ , \new_[15032]_ , \new_[15033]_ , \new_[15034]_ ,
    \new_[15035]_ , \new_[15036]_ , \new_[15037]_ , \new_[15038]_ ,
    \new_[15039]_ , \new_[15040]_ , \new_[15041]_ , \new_[15042]_ ,
    \new_[15043]_ , \new_[15044]_ , \new_[15045]_ , \new_[15046]_ ,
    \new_[15047]_ , \new_[15048]_ , \new_[15049]_ , \new_[15050]_ ,
    \new_[15051]_ , \new_[15052]_ , \new_[15053]_ , \new_[15054]_ ,
    \new_[15055]_ , \new_[15056]_ , \new_[15057]_ , \new_[15058]_ ,
    \new_[15059]_ , \new_[15060]_ , \new_[15061]_ , \new_[15062]_ ,
    \new_[15063]_ , \new_[15064]_ , \new_[15065]_ , \new_[15066]_ ,
    \new_[15067]_ , \new_[15068]_ , \new_[15069]_ , \new_[15070]_ ,
    \new_[15071]_ , \new_[15072]_ , \new_[15073]_ , \new_[15074]_ ,
    \new_[15075]_ , \new_[15076]_ , \new_[15077]_ , \new_[15078]_ ,
    \new_[15079]_ , \new_[15080]_ , \new_[15081]_ , \new_[15082]_ ,
    \new_[15083]_ , \new_[15084]_ , \new_[15085]_ , \new_[15086]_ ,
    \new_[15087]_ , \new_[15088]_ , \new_[15089]_ , \new_[15090]_ ,
    \new_[15091]_ , \new_[15092]_ , \new_[15093]_ , \new_[15094]_ ,
    \new_[15095]_ , \new_[15096]_ , \new_[15097]_ , \new_[15098]_ ,
    \new_[15099]_ , \new_[15100]_ , \new_[15101]_ , \new_[15102]_ ,
    \new_[15103]_ , \new_[15104]_ , \new_[15105]_ , \new_[15106]_ ,
    \new_[15107]_ , \new_[15108]_ , \new_[15109]_ , \new_[15110]_ ,
    \new_[15111]_ , \new_[15112]_ , \new_[15113]_ , \new_[15114]_ ,
    \new_[15115]_ , \new_[15116]_ , \new_[15117]_ , \new_[15118]_ ,
    \new_[15119]_ , \new_[15120]_ , \new_[15121]_ , \new_[15122]_ ,
    \new_[15123]_ , \new_[15124]_ , \new_[15125]_ , \new_[15126]_ ,
    \new_[15127]_ , \new_[15128]_ , \new_[15129]_ , \new_[15130]_ ,
    \new_[15131]_ , \new_[15132]_ , \new_[15133]_ , \new_[15134]_ ,
    \new_[15135]_ , \new_[15136]_ , \new_[15137]_ , \new_[15138]_ ,
    \new_[15139]_ , \new_[15140]_ , \new_[15141]_ , \new_[15142]_ ,
    \new_[15143]_ , \new_[15144]_ , \new_[15145]_ , \new_[15146]_ ,
    \new_[15147]_ , \new_[15148]_ , \new_[15149]_ , \new_[15150]_ ,
    \new_[15151]_ , \new_[15152]_ , \new_[15153]_ , \new_[15154]_ ,
    \new_[15155]_ , \new_[15156]_ , \new_[15157]_ , \new_[15158]_ ,
    \new_[15159]_ , \new_[15160]_ , \new_[15161]_ , \new_[15162]_ ,
    \new_[15163]_ , \new_[15164]_ , \new_[15165]_ , \new_[15166]_ ,
    \new_[15167]_ , \new_[15168]_ , \new_[15169]_ , \new_[15170]_ ,
    \new_[15171]_ , \new_[15172]_ , \new_[15173]_ , \new_[15174]_ ,
    \new_[15175]_ , \new_[15176]_ , \new_[15177]_ , \new_[15178]_ ,
    \new_[15179]_ , \new_[15180]_ , \new_[15181]_ , \new_[15182]_ ,
    \new_[15183]_ , \new_[15184]_ , \new_[15185]_ , \new_[15186]_ ,
    \new_[15187]_ , \new_[15188]_ , \new_[15189]_ , \new_[15190]_ ,
    \new_[15191]_ , \new_[15192]_ , \new_[15193]_ , \new_[15194]_ ,
    \new_[15195]_ , \new_[15196]_ , \new_[15197]_ , \new_[15198]_ ,
    \new_[15199]_ , \new_[15200]_ , \new_[15201]_ , \new_[15202]_ ,
    \new_[15203]_ , \new_[15204]_ , \new_[15205]_ , \new_[15206]_ ,
    \new_[15207]_ , \new_[15208]_ , \new_[15209]_ , \new_[15210]_ ,
    \new_[15211]_ , \new_[15212]_ , \new_[15213]_ , \new_[15214]_ ,
    \new_[15215]_ , \new_[15216]_ , \new_[15217]_ , \new_[15218]_ ,
    \new_[15219]_ , \new_[15220]_ , \new_[15221]_ , \new_[15222]_ ,
    \new_[15223]_ , \new_[15224]_ , \new_[15225]_ , \new_[15226]_ ,
    \new_[15227]_ , \new_[15228]_ , \new_[15229]_ , \new_[15230]_ ,
    \new_[15231]_ , \new_[15232]_ , \new_[15233]_ , \new_[15234]_ ,
    \new_[15235]_ , \new_[15236]_ , \new_[15237]_ , \new_[15238]_ ,
    \new_[15239]_ , \new_[15240]_ , \new_[15241]_ , \new_[15242]_ ,
    \new_[15243]_ , \new_[15244]_ , \new_[15245]_ , \new_[15246]_ ,
    \new_[15247]_ , \new_[15248]_ , \new_[15249]_ , \new_[15250]_ ,
    \new_[15251]_ , \new_[15252]_ , \new_[15253]_ , \new_[15254]_ ,
    \new_[15255]_ , \new_[15256]_ , \new_[15257]_ , \new_[15258]_ ,
    \new_[15259]_ , \new_[15260]_ , \new_[15261]_ , \new_[15262]_ ,
    \new_[15263]_ , \new_[15264]_ , \new_[15265]_ , \new_[15266]_ ,
    \new_[15267]_ , \new_[15268]_ , \new_[15269]_ , \new_[15270]_ ,
    \new_[15271]_ , \new_[15272]_ , \new_[15273]_ , \new_[15274]_ ,
    \new_[15275]_ , \new_[15276]_ , \new_[15277]_ , \new_[15278]_ ,
    \new_[15279]_ , \new_[15280]_ , \new_[15281]_ , \new_[15282]_ ,
    \new_[15283]_ , \new_[15284]_ , \new_[15285]_ , \new_[15286]_ ,
    \new_[15287]_ , \new_[15288]_ , \new_[15289]_ , \new_[15290]_ ,
    \new_[15291]_ , \new_[15292]_ , \new_[15293]_ , \new_[15294]_ ,
    \new_[15295]_ , \new_[15296]_ , \new_[15297]_ , \new_[15298]_ ,
    \new_[15299]_ , \new_[15300]_ , \new_[15301]_ , \new_[15302]_ ,
    \new_[15303]_ , \new_[15304]_ , \new_[15305]_ , \new_[15306]_ ,
    \new_[15307]_ , \new_[15308]_ , \new_[15309]_ , \new_[15310]_ ,
    \new_[15311]_ , \new_[15312]_ , \new_[15313]_ , \new_[15314]_ ,
    \new_[15315]_ , \new_[15316]_ , \new_[15317]_ , \new_[15318]_ ,
    \new_[15319]_ , \new_[15320]_ , \new_[15321]_ , \new_[15322]_ ,
    \new_[15323]_ , \new_[15324]_ , \new_[15325]_ , \new_[15326]_ ,
    \new_[15327]_ , \new_[15328]_ , \new_[15329]_ , \new_[15330]_ ,
    \new_[15331]_ , \new_[15332]_ , \new_[15333]_ , \new_[15334]_ ,
    \new_[15335]_ , \new_[15336]_ , \new_[15337]_ , \new_[15338]_ ,
    \new_[15339]_ , \new_[15340]_ , \new_[15341]_ , \new_[15342]_ ,
    \new_[15343]_ , \new_[15344]_ , \new_[15345]_ , \new_[15346]_ ,
    \new_[15347]_ , \new_[15348]_ , \new_[15349]_ , \new_[15350]_ ,
    \new_[15351]_ , \new_[15352]_ , \new_[15353]_ , \new_[15354]_ ,
    \new_[15355]_ , \new_[15356]_ , \new_[15357]_ , \new_[15358]_ ,
    \new_[15359]_ , \new_[15360]_ , \new_[15361]_ , \new_[15362]_ ,
    \new_[15363]_ , \new_[15364]_ , \new_[15365]_ , \new_[15366]_ ,
    \new_[15367]_ , \new_[15368]_ , \new_[15369]_ , \new_[15370]_ ,
    \new_[15371]_ , \new_[15372]_ , \new_[15373]_ , \new_[15374]_ ,
    \new_[15375]_ , \new_[15376]_ , \new_[15377]_ , \new_[15378]_ ,
    \new_[15379]_ , \new_[15380]_ , \new_[15381]_ , \new_[15382]_ ,
    \new_[15383]_ , \new_[15384]_ , \new_[15385]_ , \new_[15386]_ ,
    \new_[15387]_ , \new_[15388]_ , \new_[15389]_ , \new_[15390]_ ,
    \new_[15391]_ , \new_[15392]_ , \new_[15393]_ , \new_[15394]_ ,
    \new_[15395]_ , \new_[15396]_ , \new_[15397]_ , \new_[15398]_ ,
    \new_[15399]_ , \new_[15400]_ , \new_[15401]_ , \new_[15402]_ ,
    \new_[15403]_ , \new_[15404]_ , \new_[15405]_ , \new_[15406]_ ,
    \new_[15407]_ , \new_[15408]_ , \new_[15409]_ , \new_[15410]_ ,
    \new_[15411]_ , \new_[15412]_ , \new_[15413]_ , \new_[15414]_ ,
    \new_[15415]_ , \new_[15416]_ , \new_[15417]_ , \new_[15418]_ ,
    \new_[15419]_ , \new_[15420]_ , \new_[15421]_ , \new_[15422]_ ,
    \new_[15423]_ , \new_[15424]_ , \new_[15425]_ , \new_[15426]_ ,
    \new_[15427]_ , \new_[15428]_ , \new_[15429]_ , \new_[15430]_ ,
    \new_[15431]_ , \new_[15432]_ , \new_[15433]_ , \new_[15434]_ ,
    \new_[15435]_ , \new_[15436]_ , \new_[15437]_ , \new_[15438]_ ,
    \new_[15439]_ , \new_[15440]_ , \new_[15441]_ , \new_[15442]_ ,
    \new_[15443]_ , \new_[15444]_ , \new_[15445]_ , \new_[15446]_ ,
    \new_[15447]_ , \new_[15448]_ , \new_[15449]_ , \new_[15450]_ ,
    \new_[15451]_ , \new_[15452]_ , \new_[15453]_ , \new_[15454]_ ,
    \new_[15455]_ , \new_[15456]_ , \new_[15457]_ , \new_[15458]_ ,
    \new_[15459]_ , \new_[15460]_ , \new_[15461]_ , \new_[15462]_ ,
    \new_[15463]_ , \new_[15464]_ , \new_[15465]_ , \new_[15466]_ ,
    \new_[15467]_ , \new_[15468]_ , \new_[15469]_ , \new_[15470]_ ,
    \new_[15471]_ , \new_[15472]_ , \new_[15473]_ , \new_[15474]_ ,
    \new_[15475]_ , \new_[15476]_ , \new_[15477]_ , \new_[15478]_ ,
    \new_[15479]_ , \new_[15480]_ , \new_[15481]_ , \new_[15482]_ ,
    \new_[15483]_ , \new_[15484]_ , \new_[15485]_ , \new_[15486]_ ,
    \new_[15487]_ , \new_[15488]_ , \new_[15489]_ , \new_[15490]_ ,
    \new_[15491]_ , \new_[15492]_ , \new_[15493]_ , \new_[15494]_ ,
    \new_[15495]_ , \new_[15496]_ , \new_[15497]_ , \new_[15498]_ ,
    \new_[15499]_ , \new_[15500]_ , \new_[15501]_ , \new_[15502]_ ,
    \new_[15503]_ , \new_[15504]_ , \new_[15505]_ , \new_[15506]_ ,
    \new_[15507]_ , \new_[15508]_ , \new_[15509]_ , \new_[15510]_ ,
    \new_[15511]_ , \new_[15512]_ , \new_[15513]_ , \new_[15514]_ ,
    \new_[15515]_ , \new_[15516]_ , \new_[15517]_ , \new_[15518]_ ,
    \new_[15519]_ , \new_[15520]_ , \new_[15521]_ , \new_[15522]_ ,
    \new_[15523]_ , \new_[15524]_ , \new_[15525]_ , \new_[15526]_ ,
    \new_[15527]_ , \new_[15528]_ , \new_[15529]_ , \new_[15530]_ ,
    \new_[15531]_ , \new_[15532]_ , \new_[15533]_ , \new_[15534]_ ,
    \new_[15535]_ , \new_[15536]_ , \new_[15537]_ , \new_[15538]_ ,
    \new_[15539]_ , \new_[15540]_ , \new_[15541]_ , \new_[15542]_ ,
    \new_[15543]_ , \new_[15544]_ , \new_[15545]_ , \new_[15546]_ ,
    \new_[15547]_ , \new_[15548]_ , \new_[15549]_ , \new_[15550]_ ,
    \new_[15551]_ , \new_[15552]_ , \new_[15553]_ , \new_[15554]_ ,
    \new_[15555]_ , \new_[15556]_ , \new_[15557]_ , \new_[15558]_ ,
    \new_[15559]_ , \new_[15560]_ , \new_[15561]_ , \new_[15562]_ ,
    \new_[15563]_ , \new_[15564]_ , \new_[15565]_ , \new_[15566]_ ,
    \new_[15567]_ , \new_[15568]_ , \new_[15569]_ , \new_[15570]_ ,
    \new_[15571]_ , \new_[15572]_ , \new_[15573]_ , \new_[15574]_ ,
    \new_[15575]_ , \new_[15576]_ , \new_[15577]_ , \new_[15578]_ ,
    \new_[15579]_ , \new_[15580]_ , \new_[15581]_ , \new_[15582]_ ,
    \new_[15583]_ , \new_[15584]_ , \new_[15585]_ , \new_[15586]_ ,
    \new_[15587]_ , \new_[15588]_ , \new_[15589]_ , \new_[15590]_ ,
    \new_[15591]_ , \new_[15592]_ , \new_[15593]_ , \new_[15594]_ ,
    \new_[15595]_ , \new_[15596]_ , \new_[15597]_ , \new_[15598]_ ,
    \new_[15599]_ , \new_[15600]_ , \new_[15601]_ , \new_[15602]_ ,
    \new_[15603]_ , \new_[15604]_ , \new_[15605]_ , \new_[15606]_ ,
    \new_[15607]_ , \new_[15608]_ , \new_[15609]_ , \new_[15610]_ ,
    \new_[15611]_ , \new_[15612]_ , \new_[15613]_ , \new_[15614]_ ,
    \new_[15615]_ , \new_[15616]_ , \new_[15617]_ , \new_[15618]_ ,
    \new_[15619]_ , \new_[15620]_ , \new_[15621]_ , \new_[15622]_ ,
    \new_[15623]_ , \new_[15624]_ , \new_[15625]_ , \new_[15626]_ ,
    \new_[15627]_ , \new_[15628]_ , \new_[15629]_ , \new_[15630]_ ,
    \new_[15631]_ , \new_[15632]_ , \new_[15633]_ , \new_[15634]_ ,
    \new_[15635]_ , \new_[15636]_ , \new_[15637]_ , \new_[15638]_ ,
    \new_[15639]_ , \new_[15640]_ , \new_[15641]_ , \new_[15642]_ ,
    \new_[15643]_ , \new_[15644]_ , \new_[15645]_ , \new_[15646]_ ,
    \new_[15647]_ , \new_[15648]_ , \new_[15649]_ , \new_[15650]_ ,
    \new_[15651]_ , \new_[15652]_ , \new_[15653]_ , \new_[15654]_ ,
    \new_[15655]_ , \new_[15656]_ , \new_[15657]_ , \new_[15658]_ ,
    \new_[15659]_ , \new_[15660]_ , \new_[15661]_ , \new_[15662]_ ,
    \new_[15663]_ , \new_[15664]_ , \new_[15665]_ , \new_[15666]_ ,
    \new_[15667]_ , \new_[15668]_ , \new_[15669]_ , \new_[15670]_ ,
    \new_[15671]_ , \new_[15672]_ , \new_[15673]_ , \new_[15674]_ ,
    \new_[15675]_ , \new_[15676]_ , \new_[15677]_ , \new_[15678]_ ,
    \new_[15679]_ , \new_[15680]_ , \new_[15681]_ , \new_[15682]_ ,
    \new_[15683]_ , \new_[15684]_ , \new_[15685]_ , \new_[15686]_ ,
    \new_[15687]_ , \new_[15688]_ , \new_[15689]_ , \new_[15690]_ ,
    \new_[15691]_ , \new_[15692]_ , \new_[15693]_ , \new_[15694]_ ,
    \new_[15695]_ , \new_[15696]_ , \new_[15697]_ , \new_[15698]_ ,
    \new_[15699]_ , \new_[15700]_ , \new_[15701]_ , \new_[15702]_ ,
    \new_[15703]_ , \new_[15704]_ , \new_[15705]_ , \new_[15706]_ ,
    \new_[15707]_ , \new_[15708]_ , \new_[15709]_ , \new_[15710]_ ,
    \new_[15711]_ , \new_[15712]_ , \new_[15713]_ , \new_[15714]_ ,
    \new_[15715]_ , \new_[15716]_ , \new_[15717]_ , \new_[15718]_ ,
    \new_[15719]_ , \new_[15720]_ , \new_[15721]_ , \new_[15722]_ ,
    \new_[15723]_ , \new_[15724]_ , \new_[15725]_ , \new_[15726]_ ,
    \new_[15727]_ , \new_[15728]_ , \new_[15729]_ , \new_[15730]_ ,
    \new_[15731]_ , \new_[15732]_ , \new_[15733]_ , \new_[15734]_ ,
    \new_[15735]_ , \new_[15736]_ , \new_[15737]_ , \new_[15738]_ ,
    \new_[15739]_ , \new_[15740]_ , \new_[15741]_ , \new_[15742]_ ,
    \new_[15743]_ , \new_[15744]_ , \new_[15745]_ , \new_[15746]_ ,
    \new_[15747]_ , \new_[15748]_ , \new_[15749]_ , \new_[15750]_ ,
    \new_[15751]_ , \new_[15752]_ , \new_[15753]_ , \new_[15754]_ ,
    \new_[15755]_ , \new_[15756]_ , \new_[15757]_ , \new_[15758]_ ,
    \new_[15759]_ , \new_[15760]_ , \new_[15761]_ , \new_[15762]_ ,
    \new_[15763]_ , \new_[15764]_ , \new_[15765]_ , \new_[15766]_ ,
    \new_[15767]_ , \new_[15768]_ , \new_[15769]_ , \new_[15770]_ ,
    \new_[15771]_ , \new_[15772]_ , \new_[15773]_ , \new_[15774]_ ,
    \new_[15775]_ , \new_[15776]_ , \new_[15777]_ , \new_[15778]_ ,
    \new_[15779]_ , \new_[15780]_ , \new_[15781]_ , \new_[15782]_ ,
    \new_[15783]_ , \new_[15784]_ , \new_[15785]_ , \new_[15786]_ ,
    \new_[15787]_ , \new_[15788]_ , \new_[15789]_ , \new_[15790]_ ,
    \new_[15791]_ , \new_[15792]_ , \new_[15793]_ , \new_[15794]_ ,
    \new_[15795]_ , \new_[15796]_ , \new_[15797]_ , \new_[15798]_ ,
    \new_[15799]_ , \new_[15800]_ , \new_[15801]_ , \new_[15802]_ ,
    \new_[15803]_ , \new_[15804]_ , \new_[15805]_ , \new_[15806]_ ,
    \new_[15807]_ , \new_[15808]_ , \new_[15809]_ , \new_[15810]_ ,
    \new_[15811]_ , \new_[15812]_ , \new_[15813]_ , \new_[15814]_ ,
    \new_[15815]_ , \new_[15816]_ , \new_[15817]_ , \new_[15818]_ ,
    \new_[15819]_ , \new_[15820]_ , \new_[15821]_ , \new_[15822]_ ,
    \new_[15823]_ , \new_[15824]_ , \new_[15825]_ , \new_[15826]_ ,
    \new_[15827]_ , \new_[15828]_ , \new_[15829]_ , \new_[15830]_ ,
    \new_[15831]_ , \new_[15832]_ , \new_[15833]_ , \new_[15834]_ ,
    \new_[15835]_ , \new_[15836]_ , \new_[15837]_ , \new_[15838]_ ,
    \new_[15839]_ , \new_[15840]_ , \new_[15841]_ , \new_[15842]_ ,
    \new_[15843]_ , \new_[15844]_ , \new_[15845]_ , \new_[15846]_ ,
    \new_[15847]_ , \new_[15848]_ , \new_[15849]_ , \new_[15850]_ ,
    \new_[15851]_ , \new_[15852]_ , \new_[15853]_ , \new_[15854]_ ,
    \new_[15855]_ , \new_[15856]_ , \new_[15857]_ , \new_[15858]_ ,
    \new_[15859]_ , \new_[15860]_ , \new_[15861]_ , \new_[15862]_ ,
    \new_[15863]_ , \new_[15864]_ , \new_[15865]_ , \new_[15866]_ ,
    \new_[15867]_ , \new_[15868]_ , \new_[15869]_ , \new_[15870]_ ,
    \new_[15871]_ , \new_[15872]_ , \new_[15873]_ , \new_[15874]_ ,
    \new_[15875]_ , \new_[15876]_ , \new_[15877]_ , \new_[15878]_ ,
    \new_[15879]_ , \new_[15880]_ , \new_[15881]_ , \new_[15882]_ ,
    \new_[15883]_ , \new_[15884]_ , \new_[15885]_ , \new_[15886]_ ,
    \new_[15887]_ , \new_[15888]_ , \new_[15889]_ , \new_[15890]_ ,
    \new_[15891]_ , \new_[15892]_ , \new_[15893]_ , \new_[15894]_ ,
    \new_[15895]_ , \new_[15896]_ , \new_[15897]_ , \new_[15898]_ ,
    \new_[15899]_ , \new_[15900]_ , \new_[15901]_ , \new_[15902]_ ,
    \new_[15903]_ , \new_[15904]_ , \new_[15905]_ , \new_[15906]_ ,
    \new_[15907]_ , \new_[15908]_ , \new_[15909]_ , \new_[15910]_ ,
    \new_[15911]_ , \new_[15912]_ , \new_[15913]_ , \new_[15914]_ ,
    \new_[15915]_ , \new_[15916]_ , \new_[15917]_ , \new_[15918]_ ,
    \new_[15919]_ , \new_[15920]_ , \new_[15921]_ , \new_[15922]_ ,
    \new_[15923]_ , \new_[15924]_ , \new_[15925]_ , \new_[15926]_ ,
    \new_[15927]_ , \new_[15928]_ , \new_[15929]_ , \new_[15930]_ ,
    \new_[15931]_ , \new_[15932]_ , \new_[15933]_ , \new_[15934]_ ,
    \new_[15935]_ , \new_[15936]_ , \new_[15937]_ , \new_[15938]_ ,
    \new_[15939]_ , \new_[15940]_ , \new_[15941]_ , \new_[15942]_ ,
    \new_[15943]_ , \new_[15944]_ , \new_[15945]_ , \new_[15946]_ ,
    \new_[15947]_ , \new_[15948]_ , \new_[15949]_ , \new_[15950]_ ,
    \new_[15951]_ , \new_[15952]_ , \new_[15953]_ , \new_[15954]_ ,
    \new_[15955]_ , \new_[15956]_ , \new_[15957]_ , \new_[15958]_ ,
    \new_[15959]_ , \new_[15960]_ , \new_[15961]_ , \new_[15962]_ ,
    \new_[15963]_ , \new_[15964]_ , \new_[15965]_ , \new_[15966]_ ,
    \new_[15967]_ , \new_[15968]_ , \new_[15969]_ , \new_[15970]_ ,
    \new_[15971]_ , \new_[15972]_ , \new_[15973]_ , \new_[15974]_ ,
    \new_[15975]_ , \new_[15976]_ , \new_[15977]_ , \new_[15978]_ ,
    \new_[15979]_ , \new_[15980]_ , \new_[15981]_ , \new_[15982]_ ,
    \new_[15983]_ , \new_[15984]_ , \new_[15985]_ , \new_[15986]_ ,
    \new_[15987]_ , \new_[15988]_ , \new_[15989]_ , \new_[15990]_ ,
    \new_[15991]_ , \new_[15992]_ , \new_[15993]_ , \new_[15994]_ ,
    \new_[15995]_ , \new_[15996]_ , \new_[15997]_ , \new_[15998]_ ,
    \new_[15999]_ , \new_[16000]_ , \new_[16001]_ , \new_[16002]_ ,
    \new_[16003]_ , \new_[16004]_ , \new_[16005]_ , \new_[16006]_ ,
    \new_[16007]_ , \new_[16008]_ , \new_[16009]_ , \new_[16010]_ ,
    \new_[16011]_ , \new_[16012]_ , \new_[16013]_ , \new_[16014]_ ,
    \new_[16015]_ , \new_[16016]_ , \new_[16017]_ , \new_[16018]_ ,
    \new_[16019]_ , \new_[16020]_ , \new_[16021]_ , \new_[16022]_ ,
    \new_[16023]_ , \new_[16024]_ , \new_[16025]_ , \new_[16026]_ ,
    \new_[16027]_ , \new_[16028]_ , \new_[16029]_ , \new_[16030]_ ,
    \new_[16031]_ , \new_[16032]_ , \new_[16033]_ , \new_[16034]_ ,
    \new_[16035]_ , \new_[16036]_ , \new_[16037]_ , \new_[16038]_ ,
    \new_[16039]_ , \new_[16040]_ , \new_[16041]_ , \new_[16042]_ ,
    \new_[16043]_ , \new_[16044]_ , \new_[16045]_ , \new_[16046]_ ,
    \new_[16047]_ , \new_[16048]_ , \new_[16049]_ , \new_[16050]_ ,
    \new_[16051]_ , \new_[16052]_ , \new_[16053]_ , \new_[16054]_ ,
    \new_[16055]_ , \new_[16056]_ , \new_[16057]_ , \new_[16058]_ ,
    \new_[16059]_ , \new_[16060]_ , \new_[16061]_ , \new_[16062]_ ,
    \new_[16063]_ , \new_[16064]_ , \new_[16065]_ , \new_[16066]_ ,
    \new_[16067]_ , \new_[16068]_ , \new_[16069]_ , \new_[16070]_ ,
    \new_[16071]_ , \new_[16072]_ , \new_[16073]_ , \new_[16074]_ ,
    \new_[16075]_ , \new_[16076]_ , \new_[16077]_ , \new_[16078]_ ,
    \new_[16079]_ , \new_[16080]_ , \new_[16081]_ , \new_[16082]_ ,
    \new_[16083]_ , \new_[16084]_ , \new_[16085]_ , \new_[16086]_ ,
    \new_[16087]_ , \new_[16088]_ , \new_[16089]_ , \new_[16090]_ ,
    \new_[16091]_ , \new_[16092]_ , \new_[16093]_ , \new_[16094]_ ,
    \new_[16095]_ , \new_[16096]_ , \new_[16097]_ , \new_[16098]_ ,
    \new_[16099]_ , \new_[16100]_ , \new_[16101]_ , \new_[16102]_ ,
    \new_[16103]_ , \new_[16104]_ , \new_[16105]_ , \new_[16106]_ ,
    \new_[16107]_ , \new_[16108]_ , \new_[16109]_ , \new_[16110]_ ,
    \new_[16111]_ , \new_[16112]_ , \new_[16113]_ , \new_[16114]_ ,
    \new_[16115]_ , \new_[16116]_ , \new_[16117]_ , \new_[16118]_ ,
    \new_[16119]_ , \new_[16120]_ , \new_[16121]_ , \new_[16122]_ ,
    \new_[16123]_ , \new_[16124]_ , \new_[16125]_ , \new_[16126]_ ,
    \new_[16127]_ , \new_[16128]_ , \new_[16129]_ , \new_[16130]_ ,
    \new_[16131]_ , \new_[16132]_ , \new_[16133]_ , \new_[16134]_ ,
    \new_[16135]_ , \new_[16136]_ , \new_[16137]_ , \new_[16138]_ ,
    \new_[16139]_ , \new_[16140]_ , \new_[16141]_ , \new_[16142]_ ,
    \new_[16143]_ , \new_[16144]_ , \new_[16145]_ , \new_[16146]_ ,
    \new_[16147]_ , \new_[16148]_ , \new_[16149]_ , \new_[16150]_ ,
    \new_[16151]_ , \new_[16152]_ , \new_[16153]_ , \new_[16154]_ ,
    \new_[16155]_ , \new_[16156]_ , \new_[16157]_ , \new_[16158]_ ,
    \new_[16159]_ , \new_[16160]_ , \new_[16161]_ , \new_[16162]_ ,
    \new_[16163]_ , \new_[16164]_ , \new_[16165]_ , \new_[16166]_ ,
    \new_[16167]_ , \new_[16168]_ , \new_[16169]_ , \new_[16170]_ ,
    \new_[16171]_ , \new_[16172]_ , \new_[16173]_ , \new_[16174]_ ,
    \new_[16175]_ , \new_[16176]_ , \new_[16177]_ , \new_[16178]_ ,
    \new_[16179]_ , \new_[16180]_ , \new_[16181]_ , \new_[16182]_ ,
    \new_[16183]_ , \new_[16184]_ , \new_[16185]_ , \new_[16186]_ ,
    \new_[16187]_ , \new_[16188]_ , \new_[16189]_ , \new_[16190]_ ,
    \new_[16191]_ , \new_[16192]_ , \new_[16193]_ , \new_[16194]_ ,
    \new_[16195]_ , \new_[16196]_ , \new_[16197]_ , \new_[16198]_ ,
    \new_[16199]_ , \new_[16200]_ , \new_[16201]_ , \new_[16202]_ ,
    \new_[16203]_ , \new_[16204]_ , \new_[16205]_ , \new_[16206]_ ,
    \new_[16207]_ , \new_[16208]_ , \new_[16209]_ , \new_[16210]_ ,
    \new_[16211]_ , \new_[16212]_ , \new_[16213]_ , \new_[16214]_ ,
    \new_[16215]_ , \new_[16216]_ , \new_[16217]_ , \new_[16218]_ ,
    \new_[16219]_ , \new_[16220]_ , \new_[16221]_ , \new_[16222]_ ,
    \new_[16223]_ , \new_[16224]_ , \new_[16225]_ , \new_[16226]_ ,
    \new_[16227]_ , \new_[16228]_ , \new_[16229]_ , \new_[16230]_ ,
    \new_[16231]_ , \new_[16232]_ , \new_[16233]_ , \new_[16234]_ ,
    \new_[16235]_ , \new_[16236]_ , \new_[16237]_ , \new_[16238]_ ,
    \new_[16239]_ , \new_[16240]_ , \new_[16241]_ , \new_[16242]_ ,
    \new_[16243]_ , \new_[16244]_ , \new_[16245]_ , \new_[16246]_ ,
    \new_[16247]_ , \new_[16249]_ , \new_[16250]_ , \new_[16251]_ ,
    \new_[16252]_ , \new_[16253]_ , \new_[16254]_ , \new_[16255]_ ,
    \new_[16256]_ , \new_[16257]_ , \new_[16258]_ , \new_[16259]_ ,
    \new_[16260]_ , \new_[16261]_ , \new_[16262]_ , \new_[16263]_ ,
    \new_[16264]_ , \new_[16265]_ , \new_[16266]_ , \new_[16267]_ ,
    \new_[16268]_ , \new_[16269]_ , \new_[16270]_ , \new_[16271]_ ,
    \new_[16272]_ , \new_[16273]_ , \new_[16274]_ , \new_[16275]_ ,
    \new_[16276]_ , \new_[16277]_ , \new_[16278]_ , \new_[16279]_ ,
    \new_[16280]_ , \new_[16281]_ , \new_[16282]_ , \new_[16283]_ ,
    \new_[16284]_ , \new_[16285]_ , \new_[16286]_ , \new_[16287]_ ,
    \new_[16288]_ , \new_[16289]_ , \new_[16290]_ , \new_[16291]_ ,
    \new_[16292]_ , \new_[16293]_ , \new_[16294]_ , \new_[16295]_ ,
    \new_[16296]_ , \new_[16297]_ , \new_[16298]_ , \new_[16299]_ ,
    \new_[16300]_ , \new_[16301]_ , \new_[16302]_ , \new_[16303]_ ,
    \new_[16304]_ , \new_[16305]_ , \new_[16306]_ , \new_[16307]_ ,
    \new_[16308]_ , \new_[16309]_ , \new_[16310]_ , \new_[16311]_ ,
    \new_[16312]_ , \new_[16313]_ , \new_[16314]_ , \new_[16315]_ ,
    \new_[16316]_ , \new_[16317]_ , \new_[16318]_ , \new_[16319]_ ,
    \new_[16320]_ , \new_[16321]_ , \new_[16322]_ , \new_[16323]_ ,
    \new_[16324]_ , \new_[16325]_ , \new_[16326]_ , \new_[16327]_ ,
    \new_[16328]_ , \new_[16329]_ , \new_[16330]_ , \new_[16331]_ ,
    \new_[16332]_ , \new_[16333]_ , \new_[16334]_ , \new_[16335]_ ,
    \new_[16336]_ , \new_[16337]_ , \new_[16338]_ , \new_[16339]_ ,
    \new_[16340]_ , \new_[16341]_ , \new_[16342]_ , \new_[16343]_ ,
    \new_[16344]_ , \new_[16345]_ , \new_[16346]_ , \new_[16347]_ ,
    \new_[16348]_ , \new_[16349]_ , \new_[16350]_ , \new_[16351]_ ,
    \new_[16352]_ , \new_[16353]_ , \new_[16354]_ , \new_[16355]_ ,
    \new_[16356]_ , \new_[16357]_ , \new_[16358]_ , \new_[16359]_ ,
    \new_[16360]_ , \new_[16361]_ , \new_[16362]_ , \new_[16363]_ ,
    \new_[16364]_ , \new_[16365]_ , \new_[16366]_ , \new_[16367]_ ,
    \new_[16368]_ , \new_[16369]_ , \new_[16370]_ , \new_[16371]_ ,
    \new_[16372]_ , \new_[16373]_ , \new_[16374]_ , \new_[16375]_ ,
    \new_[16376]_ , \new_[16377]_ , \new_[16378]_ , \new_[16379]_ ,
    \new_[16380]_ , \new_[16381]_ , \new_[16382]_ , \new_[16383]_ ,
    \new_[16384]_ , \new_[16385]_ , \new_[16386]_ , \new_[16387]_ ,
    \new_[16388]_ , \new_[16389]_ , \new_[16390]_ , \new_[16391]_ ,
    \new_[16392]_ , \new_[16393]_ , \new_[16394]_ , \new_[16395]_ ,
    \new_[16396]_ , \new_[16397]_ , \new_[16398]_ , \new_[16399]_ ,
    \new_[16400]_ , \new_[16401]_ , \new_[16402]_ , \new_[16403]_ ,
    \new_[16404]_ , \new_[16405]_ , \new_[16406]_ , \new_[16407]_ ,
    \new_[16408]_ , \new_[16409]_ , \new_[16410]_ , \new_[16411]_ ,
    \new_[16412]_ , \new_[16413]_ , \new_[16414]_ , \new_[16415]_ ,
    \new_[16416]_ , \new_[16417]_ , \new_[16418]_ , \new_[16419]_ ,
    \new_[16420]_ , \new_[16421]_ , \new_[16422]_ , \new_[16423]_ ,
    \new_[16424]_ , \new_[16425]_ , \new_[16426]_ , \new_[16427]_ ,
    \new_[16428]_ , \new_[16429]_ , \new_[16430]_ , \new_[16431]_ ,
    \new_[16432]_ , \new_[16433]_ , \new_[16434]_ , \new_[16435]_ ,
    \new_[16436]_ , \new_[16437]_ , \new_[16438]_ , \new_[16439]_ ,
    \new_[16440]_ , \new_[16441]_ , \new_[16442]_ , \new_[16443]_ ,
    \new_[16444]_ , \new_[16445]_ , \new_[16446]_ , \new_[16447]_ ,
    \new_[16448]_ , \new_[16449]_ , \new_[16450]_ , \new_[16451]_ ,
    \new_[16452]_ , \new_[16453]_ , \new_[16454]_ , \new_[16455]_ ,
    \new_[16456]_ , \new_[16457]_ , \new_[16458]_ , \new_[16459]_ ,
    \new_[16460]_ , \new_[16461]_ , \new_[16462]_ , \new_[16463]_ ,
    \new_[16464]_ , \new_[16465]_ , \new_[16466]_ , \new_[16467]_ ,
    \new_[16468]_ , \new_[16469]_ , \new_[16470]_ , \new_[16471]_ ,
    \new_[16472]_ , \new_[16473]_ , \new_[16474]_ , \new_[16475]_ ,
    \new_[16476]_ , \new_[16477]_ , \new_[16478]_ , \new_[16479]_ ,
    \new_[16480]_ , \new_[16481]_ , \new_[16482]_ , \new_[16483]_ ,
    \new_[16484]_ , \new_[16485]_ , \new_[16486]_ , \new_[16487]_ ,
    \new_[16488]_ , \new_[16489]_ , \new_[16490]_ , \new_[16491]_ ,
    \new_[16492]_ , \new_[16493]_ , \new_[16494]_ , \new_[16495]_ ,
    \new_[16496]_ , \new_[16497]_ , \new_[16498]_ , \new_[16499]_ ,
    \new_[16500]_ , \new_[16501]_ , \new_[16502]_ , \new_[16503]_ ,
    \new_[16504]_ , \new_[16505]_ , \new_[16506]_ , \new_[16507]_ ,
    \new_[16508]_ , \new_[16509]_ , \new_[16510]_ , \new_[16511]_ ,
    \new_[16512]_ , \new_[16513]_ , \new_[16514]_ , \new_[16515]_ ,
    \new_[16516]_ , \new_[16517]_ , \new_[16518]_ , \new_[16519]_ ,
    \new_[16520]_ , \new_[16521]_ , \new_[16522]_ , \new_[16523]_ ,
    \new_[16524]_ , \new_[16525]_ , \new_[16526]_ , \new_[16527]_ ,
    \new_[16528]_ , \new_[16529]_ , \new_[16530]_ , \new_[16531]_ ,
    \new_[16532]_ , \new_[16533]_ , \new_[16534]_ , \new_[16535]_ ,
    \new_[16536]_ , \new_[16537]_ , \new_[16538]_ , \new_[16539]_ ,
    \new_[16540]_ , \new_[16541]_ , \new_[16542]_ , \new_[16543]_ ,
    \new_[16544]_ , \new_[16545]_ , \new_[16546]_ , \new_[16547]_ ,
    \new_[16548]_ , \new_[16549]_ , \new_[16550]_ , \new_[16551]_ ,
    \new_[16552]_ , \new_[16553]_ , \new_[16554]_ , \new_[16555]_ ,
    \new_[16556]_ , \new_[16557]_ , \new_[16558]_ , \new_[16559]_ ,
    \new_[16560]_ , \new_[16561]_ , \new_[16562]_ , \new_[16563]_ ,
    \new_[16564]_ , \new_[16565]_ , \new_[16566]_ , \new_[16567]_ ,
    \new_[16568]_ , \new_[16569]_ , \new_[16570]_ , \new_[16571]_ ,
    \new_[16572]_ , \new_[16573]_ , \new_[16574]_ , \new_[16575]_ ,
    \new_[16576]_ , \new_[16577]_ , \new_[16578]_ , \new_[16579]_ ,
    \new_[16580]_ , \new_[16581]_ , \new_[16582]_ , \new_[16583]_ ,
    \new_[16584]_ , \new_[16585]_ , \new_[16586]_ , \new_[16587]_ ,
    \new_[16588]_ , \new_[16589]_ , \new_[16590]_ , \new_[16591]_ ,
    \new_[16592]_ , \new_[16593]_ , \new_[16594]_ , \new_[16595]_ ,
    \new_[16596]_ , \new_[16597]_ , \new_[16598]_ , \new_[16599]_ ,
    \new_[16600]_ , \new_[16601]_ , \new_[16602]_ , \new_[16603]_ ,
    \new_[16604]_ , \new_[16605]_ , \new_[16606]_ , \new_[16607]_ ,
    \new_[16608]_ , \new_[16609]_ , \new_[16610]_ , \new_[16611]_ ,
    \new_[16612]_ , \new_[16613]_ , \new_[16614]_ , \new_[16615]_ ,
    \new_[16616]_ , \new_[16617]_ , \new_[16618]_ , \new_[16619]_ ,
    \new_[16620]_ , \new_[16621]_ , \new_[16622]_ , \new_[16623]_ ,
    \new_[16624]_ , \new_[16625]_ , \new_[16626]_ , \new_[16627]_ ,
    \new_[16628]_ , \new_[16629]_ , \new_[16630]_ , \new_[16631]_ ,
    \new_[16632]_ , \new_[16633]_ , \new_[16634]_ , \new_[16635]_ ,
    \new_[16636]_ , \new_[16637]_ , \new_[16638]_ , \new_[16639]_ ,
    \new_[16640]_ , \new_[16641]_ , \new_[16642]_ , \new_[16643]_ ,
    \new_[16644]_ , \new_[16645]_ , \new_[16646]_ , \new_[16647]_ ,
    \new_[16648]_ , \new_[16649]_ , \new_[16650]_ , \new_[16651]_ ,
    \new_[16652]_ , \new_[16653]_ , \new_[16654]_ , \new_[16655]_ ,
    \new_[16656]_ , \new_[16657]_ , \new_[16658]_ , \new_[16659]_ ,
    \new_[16660]_ , \new_[16661]_ , \new_[16662]_ , \new_[16663]_ ,
    \new_[16664]_ , \new_[16665]_ , \new_[16666]_ , \new_[16667]_ ,
    \new_[16668]_ , \new_[16669]_ , \new_[16670]_ , \new_[16671]_ ,
    \new_[16672]_ , \new_[16673]_ , \new_[16674]_ , \new_[16675]_ ,
    \new_[16676]_ , \new_[16677]_ , \new_[16678]_ , \new_[16679]_ ,
    \new_[16680]_ , \new_[16681]_ , \new_[16682]_ , \new_[16683]_ ,
    \new_[16684]_ , \new_[16686]_ , \new_[16687]_ , \new_[16689]_ ,
    \new_[16690]_ , \new_[16691]_ , \new_[16692]_ , \new_[16693]_ ,
    \new_[16695]_ , \new_[16696]_ , \new_[16698]_ , \new_[16699]_ ,
    \new_[16700]_ , \new_[16701]_ , \new_[16702]_ , \new_[16703]_ ,
    \new_[16704]_ , \new_[16705]_ , \new_[16706]_ , \new_[16708]_ ,
    \new_[16709]_ , \new_[16710]_ , \new_[16711]_ , \new_[16712]_ ,
    \new_[16713]_ , \new_[16714]_ , \new_[16715]_ , \new_[16716]_ ,
    \new_[16718]_ , \new_[16719]_ , \new_[16720]_ , \new_[16721]_ ,
    \new_[16722]_ , \new_[16723]_ , \new_[16724]_ , \new_[16727]_ ,
    \new_[16728]_ , \new_[16729]_ , \new_[16730]_ , \new_[16731]_ ,
    \new_[16732]_ , \new_[16733]_ , \new_[16734]_ , \new_[16735]_ ,
    \new_[16737]_ , \new_[16738]_ , \new_[16739]_ , \new_[16740]_ ,
    \new_[16741]_ , \new_[16742]_ , \new_[16743]_ , \new_[16744]_ ,
    \new_[16745]_ , \new_[16746]_ , \new_[16747]_ , \new_[16748]_ ,
    \new_[16749]_ , \new_[16750]_ , \new_[16751]_ , \new_[16752]_ ,
    \new_[16753]_ , \new_[16754]_ , \new_[16755]_ , \new_[16756]_ ,
    \new_[16757]_ , \new_[16758]_ , \new_[16759]_ , \new_[16760]_ ,
    \new_[16762]_ , \new_[16763]_ , \new_[16764]_ , \new_[16765]_ ,
    \new_[16766]_ , \new_[16767]_ , \new_[16768]_ , \new_[16769]_ ,
    \new_[16770]_ , \new_[16771]_ , \new_[16772]_ , \new_[16773]_ ,
    \new_[16775]_ , \new_[16776]_ , \new_[16777]_ , \new_[16778]_ ,
    \new_[16780]_ , \new_[16781]_ , \new_[16782]_ , \new_[16783]_ ,
    \new_[16784]_ , \new_[16785]_ , \new_[16786]_ , \new_[16787]_ ,
    \new_[16788]_ , \new_[16789]_ , \new_[16790]_ , \new_[16791]_ ,
    \new_[16792]_ , \new_[16793]_ , \new_[16794]_ , \new_[16795]_ ,
    \new_[16796]_ , \new_[16797]_ , \new_[16798]_ , \new_[16799]_ ,
    \new_[16800]_ , \new_[16801]_ , \new_[16802]_ , \new_[16803]_ ,
    \new_[16804]_ , \new_[16805]_ , \new_[16806]_ , \new_[16807]_ ,
    \new_[16808]_ , \new_[16809]_ , \new_[16810]_ , \new_[16811]_ ,
    \new_[16812]_ , \new_[16813]_ , \new_[16814]_ , \new_[16815]_ ,
    \new_[16816]_ , \new_[16817]_ , \new_[16818]_ , \new_[16820]_ ,
    \new_[16821]_ , \new_[16823]_ , \new_[16824]_ , \new_[16825]_ ,
    \new_[16826]_ , \new_[16827]_ , \new_[16828]_ , \new_[16829]_ ,
    \new_[16830]_ , \new_[16831]_ , \new_[16832]_ , \new_[16833]_ ,
    \new_[16834]_ , \new_[16835]_ , \new_[16836]_ , \new_[16837]_ ,
    \new_[16838]_ , \new_[16839]_ , \new_[16840]_ , \new_[16842]_ ,
    \new_[16843]_ , \new_[16844]_ , \new_[16845]_ , \new_[16846]_ ,
    \new_[16847]_ , \new_[16848]_ , \new_[16849]_ , \new_[16850]_ ,
    \new_[16851]_ , \new_[16853]_ , \new_[16854]_ , \new_[16855]_ ,
    \new_[16857]_ , \new_[16858]_ , \new_[16859]_ , \new_[16860]_ ,
    \new_[16861]_ , \new_[16862]_ , \new_[16863]_ , \new_[16864]_ ,
    \new_[16865]_ , \new_[16866]_ , \new_[16867]_ , \new_[16869]_ ,
    \new_[16870]_ , \new_[16871]_ , \new_[16872]_ , \new_[16873]_ ,
    \new_[16874]_ , \new_[16875]_ , \new_[16876]_ , \new_[16877]_ ,
    \new_[16878]_ , \new_[16879]_ , \new_[16880]_ , \new_[16881]_ ,
    \new_[16882]_ , \new_[16883]_ , \new_[16884]_ , \new_[16885]_ ,
    \new_[16886]_ , \new_[16887]_ , \new_[16888]_ , \new_[16889]_ ,
    \new_[16890]_ , \new_[16891]_ , \new_[16892]_ , \new_[16893]_ ,
    \new_[16894]_ , \new_[16896]_ , \new_[16897]_ , \new_[16898]_ ,
    \new_[16899]_ , \new_[16900]_ , \new_[16901]_ , \new_[16902]_ ,
    \new_[16903]_ , \new_[16904]_ , \new_[16905]_ , \new_[16906]_ ,
    \new_[16907]_ , \new_[16908]_ , \new_[16909]_ , \new_[16910]_ ,
    \new_[16911]_ , \new_[16912]_ , \new_[16913]_ , \new_[16914]_ ,
    \new_[16915]_ , \new_[16916]_ , \new_[16918]_ , \new_[16919]_ ,
    \new_[16920]_ , \new_[16921]_ , \new_[16922]_ , \new_[16923]_ ,
    \new_[16924]_ , \new_[16925]_ , \new_[16926]_ , \new_[16927]_ ,
    \new_[16928]_ , \new_[16929]_ , \new_[16930]_ , \new_[16931]_ ,
    \new_[16932]_ , \new_[16933]_ , \new_[16934]_ , \new_[16935]_ ,
    \new_[16937]_ , \new_[16939]_ , \new_[16940]_ , \new_[16941]_ ,
    \new_[16942]_ , \new_[16943]_ , \new_[16945]_ , \new_[16946]_ ,
    \new_[16947]_ , \new_[16949]_ , \new_[16952]_ , \new_[16953]_ ,
    \new_[16954]_ , \new_[16955]_ , \new_[16956]_ , \new_[16958]_ ,
    \new_[16959]_ , \new_[16961]_ , \new_[16963]_ , \new_[16965]_ ,
    \new_[16967]_ , \new_[16969]_ , \new_[16970]_ , \new_[16972]_ ,
    \new_[16973]_ , \new_[16974]_ , \new_[16976]_ , \new_[16977]_ ,
    \new_[16978]_ , \new_[16979]_ , \new_[16980]_ , \new_[16981]_ ,
    \new_[16982]_ , \new_[16983]_ , \new_[16984]_ , \new_[16985]_ ,
    \new_[16986]_ , \new_[16987]_ , \new_[16988]_ , \new_[16990]_ ,
    \new_[16991]_ , \new_[16992]_ , \new_[16993]_ , \new_[16994]_ ,
    \new_[16995]_ , \new_[16996]_ , \new_[16997]_ , \new_[16998]_ ,
    \new_[16999]_ , \new_[17000]_ , \new_[17001]_ , \new_[17002]_ ,
    \new_[17003]_ , \new_[17004]_ , \new_[17005]_ , \new_[17006]_ ,
    \new_[17007]_ , \new_[17009]_ , \new_[17010]_ , \new_[17011]_ ,
    \new_[17012]_ , \new_[17013]_ , \new_[17014]_ , \new_[17015]_ ,
    \new_[17016]_ , \new_[17017]_ , \new_[17018]_ , \new_[17019]_ ,
    \new_[17020]_ , \new_[17023]_ , \new_[17024]_ , \new_[17025]_ ,
    \new_[17026]_ , \new_[17027]_ , \new_[17028]_ , \new_[17029]_ ,
    \new_[17030]_ , \new_[17031]_ , \new_[17032]_ , \new_[17033]_ ,
    \new_[17034]_ , \new_[17036]_ , \new_[17038]_ , \new_[17039]_ ,
    \new_[17040]_ , \new_[17041]_ , \new_[17042]_ , \new_[17043]_ ,
    \new_[17044]_ , \new_[17045]_ , \new_[17046]_ , \new_[17047]_ ,
    \new_[17048]_ , \new_[17049]_ , \new_[17051]_ , \new_[17052]_ ,
    \new_[17053]_ , \new_[17054]_ , \new_[17055]_ , \new_[17056]_ ,
    \new_[17057]_ , \new_[17058]_ , \new_[17060]_ , \new_[17061]_ ,
    \new_[17062]_ , \new_[17063]_ , \new_[17064]_ , \new_[17065]_ ,
    \new_[17066]_ , \new_[17067]_ , \new_[17068]_ , \new_[17070]_ ,
    \new_[17071]_ , \new_[17072]_ , \new_[17073]_ , \new_[17074]_ ,
    \new_[17075]_ , \new_[17076]_ , \new_[17077]_ , \new_[17079]_ ,
    \new_[17080]_ , \new_[17081]_ , \new_[17082]_ , \new_[17083]_ ,
    \new_[17084]_ , \new_[17085]_ , \new_[17086]_ , \new_[17087]_ ,
    \new_[17088]_ , \new_[17089]_ , \new_[17090]_ , \new_[17091]_ ,
    \new_[17092]_ , \new_[17093]_ , \new_[17094]_ , \new_[17095]_ ,
    \new_[17096]_ , \new_[17097]_ , \new_[17098]_ , \new_[17100]_ ,
    \new_[17101]_ , \new_[17102]_ , \new_[17104]_ , \new_[17105]_ ,
    \new_[17106]_ , \new_[17107]_ , \new_[17108]_ , \new_[17109]_ ,
    \new_[17110]_ , \new_[17112]_ , \new_[17113]_ , \new_[17114]_ ,
    \new_[17115]_ , \new_[17116]_ , \new_[17117]_ , \new_[17119]_ ,
    \new_[17121]_ , \new_[17123]_ , \new_[17125]_ , \new_[17129]_ ,
    \new_[17131]_ , \new_[17132]_ , \new_[17133]_ , \new_[17135]_ ,
    \new_[17137]_ , \new_[17138]_ , \new_[17139]_ , \new_[17141]_ ,
    \new_[17142]_ , \new_[17143]_ , \new_[17144]_ , \new_[17145]_ ,
    \new_[17146]_ , \new_[17147]_ , \new_[17148]_ , \new_[17149]_ ,
    \new_[17152]_ , \new_[17153]_ , \new_[17154]_ , \new_[17155]_ ,
    \new_[17156]_ , \new_[17158]_ , \new_[17159]_ , \new_[17162]_ ,
    \new_[17164]_ , \new_[17165]_ , \new_[17166]_ , \new_[17167]_ ,
    \new_[17168]_ , \new_[17169]_ , \new_[17170]_ , \new_[17171]_ ,
    \new_[17172]_ , \new_[17173]_ , \new_[17174]_ , \new_[17175]_ ,
    \new_[17176]_ , \new_[17178]_ , \new_[17179]_ , \new_[17180]_ ,
    \new_[17181]_ , \new_[17182]_ , \new_[17183]_ , \new_[17185]_ ,
    \new_[17186]_ , \new_[17188]_ , \new_[17189]_ , \new_[17190]_ ,
    \new_[17191]_ , \new_[17192]_ , \new_[17193]_ , \new_[17194]_ ,
    \new_[17195]_ , \new_[17196]_ , \new_[17197]_ , \new_[17199]_ ,
    \new_[17200]_ , \new_[17201]_ , \new_[17202]_ , \new_[17203]_ ,
    \new_[17204]_ , \new_[17205]_ , \new_[17206]_ , \new_[17207]_ ,
    \new_[17208]_ , \new_[17209]_ , \new_[17210]_ , \new_[17211]_ ,
    \new_[17212]_ , \new_[17213]_ , \new_[17214]_ , \new_[17215]_ ,
    \new_[17216]_ , \new_[17217]_ , \new_[17218]_ , \new_[17219]_ ,
    \new_[17220]_ , \new_[17221]_ , \new_[17222]_ , \new_[17223]_ ,
    \new_[17225]_ , \new_[17226]_ , \new_[17227]_ , \new_[17229]_ ,
    \new_[17230]_ , \new_[17231]_ , \new_[17233]_ , \new_[17235]_ ,
    \new_[17236]_ , \new_[17237]_ , \new_[17238]_ , \new_[17239]_ ,
    \new_[17240]_ , \new_[17241]_ , \new_[17242]_ , \new_[17243]_ ,
    \new_[17244]_ , \new_[17245]_ , \new_[17246]_ , \new_[17247]_ ,
    \new_[17248]_ , \new_[17249]_ , \new_[17250]_ , \new_[17251]_ ,
    \new_[17252]_ , \new_[17253]_ , \new_[17254]_ , \new_[17255]_ ,
    \new_[17256]_ , \new_[17257]_ , \new_[17258]_ , \new_[17259]_ ,
    \new_[17260]_ , \new_[17261]_ , \new_[17262]_ , \new_[17263]_ ,
    \new_[17264]_ , \new_[17265]_ , \new_[17266]_ , \new_[17267]_ ,
    \new_[17268]_ , \new_[17269]_ , \new_[17270]_ , \new_[17271]_ ,
    \new_[17273]_ , \new_[17274]_ , \new_[17275]_ , \new_[17277]_ ,
    \new_[17278]_ , \new_[17279]_ , \new_[17280]_ , \new_[17282]_ ,
    \new_[17283]_ , \new_[17284]_ , \new_[17285]_ , \new_[17287]_ ,
    \new_[17289]_ , \new_[17292]_ , \new_[17295]_ , \new_[17296]_ ,
    \new_[17298]_ , \new_[17300]_ , \new_[17301]_ , \new_[17302]_ ,
    \new_[17304]_ , \new_[17305]_ , \new_[17306]_ , \new_[17307]_ ,
    \new_[17308]_ , \new_[17309]_ , \new_[17310]_ , \new_[17311]_ ,
    \new_[17312]_ , \new_[17313]_ , \new_[17314]_ , \new_[17315]_ ,
    \new_[17316]_ , \new_[17317]_ , \new_[17318]_ , \new_[17319]_ ,
    \new_[17320]_ , \new_[17321]_ , \new_[17322]_ , \new_[17323]_ ,
    \new_[17324]_ , \new_[17325]_ , \new_[17326]_ , \new_[17327]_ ,
    \new_[17328]_ , \new_[17329]_ , \new_[17330]_ , \new_[17332]_ ,
    \new_[17333]_ , \new_[17334]_ , \new_[17335]_ , \new_[17336]_ ,
    \new_[17337]_ , \new_[17338]_ , \new_[17339]_ , \new_[17340]_ ,
    \new_[17341]_ , \new_[17342]_ , \new_[17343]_ , \new_[17344]_ ,
    \new_[17345]_ , \new_[17346]_ , \new_[17347]_ , \new_[17348]_ ,
    \new_[17349]_ , \new_[17350]_ , \new_[17351]_ , \new_[17352]_ ,
    \new_[17353]_ , \new_[17354]_ , \new_[17355]_ , \new_[17356]_ ,
    \new_[17357]_ , \new_[17358]_ , \new_[17359]_ , \new_[17360]_ ,
    \new_[17361]_ , \new_[17362]_ , \new_[17363]_ , \new_[17364]_ ,
    \new_[17365]_ , \new_[17366]_ , \new_[17367]_ , \new_[17368]_ ,
    \new_[17369]_ , \new_[17370]_ , \new_[17371]_ , \new_[17372]_ ,
    \new_[17373]_ , \new_[17375]_ , \new_[17376]_ , \new_[17377]_ ,
    \new_[17378]_ , \new_[17379]_ , \new_[17380]_ , \new_[17381]_ ,
    \new_[17382]_ , \new_[17383]_ , \new_[17384]_ , \new_[17385]_ ,
    \new_[17386]_ , \new_[17387]_ , \new_[17388]_ , \new_[17389]_ ,
    \new_[17390]_ , \new_[17391]_ , \new_[17392]_ , \new_[17393]_ ,
    \new_[17394]_ , \new_[17395]_ , \new_[17396]_ , \new_[17397]_ ,
    \new_[17399]_ , \new_[17400]_ , \new_[17401]_ , \new_[17402]_ ,
    \new_[17403]_ , \new_[17404]_ , \new_[17405]_ , \new_[17406]_ ,
    \new_[17407]_ , \new_[17408]_ , \new_[17409]_ , \new_[17410]_ ,
    \new_[17411]_ , \new_[17412]_ , \new_[17413]_ , \new_[17414]_ ,
    \new_[17415]_ , \new_[17416]_ , \new_[17417]_ , \new_[17418]_ ,
    \new_[17420]_ , \new_[17421]_ , \new_[17422]_ , \new_[17423]_ ,
    \new_[17424]_ , \new_[17425]_ , \new_[17426]_ , \new_[17427]_ ,
    \new_[17428]_ , \new_[17430]_ , \new_[17431]_ , \new_[17432]_ ,
    \new_[17433]_ , \new_[17434]_ , \new_[17435]_ , \new_[17436]_ ,
    \new_[17437]_ , \new_[17438]_ , \new_[17439]_ , \new_[17440]_ ,
    \new_[17441]_ , \new_[17443]_ , \new_[17444]_ , \new_[17445]_ ,
    \new_[17446]_ , \new_[17447]_ , \new_[17448]_ , \new_[17449]_ ,
    \new_[17450]_ , \new_[17451]_ , \new_[17452]_ , \new_[17453]_ ,
    \new_[17454]_ , \new_[17455]_ , \new_[17456]_ , \new_[17457]_ ,
    \new_[17458]_ , \new_[17459]_ , \new_[17460]_ , \new_[17461]_ ,
    \new_[17462]_ , \new_[17463]_ , \new_[17464]_ , \new_[17465]_ ,
    \new_[17466]_ , \new_[17467]_ , \new_[17468]_ , \new_[17469]_ ,
    \new_[17470]_ , \new_[17471]_ , \new_[17472]_ , \new_[17473]_ ,
    \new_[17474]_ , \new_[17475]_ , \new_[17476]_ , \new_[17477]_ ,
    \new_[17478]_ , \new_[17479]_ , \new_[17480]_ , \new_[17481]_ ,
    \new_[17482]_ , \new_[17483]_ , \new_[17484]_ , \new_[17485]_ ,
    \new_[17486]_ , \new_[17487]_ , \new_[17488]_ , \new_[17489]_ ,
    \new_[17490]_ , \new_[17491]_ , \new_[17492]_ , \new_[17493]_ ,
    \new_[17494]_ , \new_[17495]_ , \new_[17496]_ , \new_[17497]_ ,
    \new_[17498]_ , \new_[17499]_ , \new_[17500]_ , \new_[17501]_ ,
    \new_[17502]_ , \new_[17503]_ , \new_[17504]_ , \new_[17505]_ ,
    \new_[17506]_ , \new_[17507]_ , \new_[17508]_ , \new_[17509]_ ,
    \new_[17510]_ , \new_[17511]_ , \new_[17512]_ , \new_[17513]_ ,
    \new_[17514]_ , \new_[17515]_ , \new_[17516]_ , \new_[17517]_ ,
    \new_[17518]_ , \new_[17519]_ , \new_[17520]_ , \new_[17521]_ ,
    \new_[17522]_ , \new_[17523]_ , \new_[17524]_ , \new_[17525]_ ,
    \new_[17526]_ , \new_[17527]_ , \new_[17528]_ , \new_[17529]_ ,
    \new_[17530]_ , \new_[17531]_ , \new_[17532]_ , \new_[17533]_ ,
    \new_[17534]_ , \new_[17535]_ , \new_[17536]_ , \new_[17537]_ ,
    \new_[17538]_ , \new_[17539]_ , \new_[17540]_ , \new_[17541]_ ,
    \new_[17542]_ , \new_[17543]_ , \new_[17544]_ , \new_[17545]_ ,
    \new_[17546]_ , \new_[17547]_ , \new_[17548]_ , \new_[17549]_ ,
    \new_[17550]_ , \new_[17551]_ , \new_[17552]_ , \new_[17553]_ ,
    \new_[17554]_ , \new_[17555]_ , \new_[17556]_ , \new_[17557]_ ,
    \new_[17558]_ , \new_[17559]_ , \new_[17560]_ , \new_[17561]_ ,
    \new_[17562]_ , \new_[17563]_ , \new_[17564]_ , \new_[17565]_ ,
    \new_[17566]_ , \new_[17567]_ , \new_[17569]_ , \new_[17570]_ ,
    \new_[17571]_ , \new_[17572]_ , \new_[17573]_ , \new_[17574]_ ,
    \new_[17575]_ , \new_[17576]_ , \new_[17577]_ , \new_[17578]_ ,
    \new_[17579]_ , \new_[17580]_ , \new_[17581]_ , \new_[17582]_ ,
    \new_[17583]_ , \new_[17584]_ , \new_[17585]_ , \new_[17586]_ ,
    \new_[17587]_ , \new_[17588]_ , \new_[17589]_ , \new_[17590]_ ,
    \new_[17591]_ , \new_[17592]_ , \new_[17593]_ , \new_[17594]_ ,
    \new_[17595]_ , \new_[17596]_ , \new_[17597]_ , \new_[17598]_ ,
    \new_[17599]_ , \new_[17600]_ , \new_[17601]_ , \new_[17602]_ ,
    \new_[17603]_ , \new_[17604]_ , \new_[17605]_ , \new_[17606]_ ,
    \new_[17607]_ , \new_[17608]_ , \new_[17609]_ , \new_[17610]_ ,
    \new_[17611]_ , \new_[17612]_ , \new_[17613]_ , \new_[17614]_ ,
    \new_[17615]_ , \new_[17616]_ , \new_[17617]_ , \new_[17618]_ ,
    \new_[17619]_ , \new_[17620]_ , \new_[17621]_ , \new_[17622]_ ,
    \new_[17623]_ , \new_[17624]_ , \new_[17625]_ , \new_[17626]_ ,
    \new_[17627]_ , \new_[17628]_ , \new_[17629]_ , \new_[17630]_ ,
    \new_[17631]_ , \new_[17632]_ , \new_[17633]_ , \new_[17634]_ ,
    \new_[17635]_ , \new_[17636]_ , \new_[17637]_ , \new_[17638]_ ,
    \new_[17639]_ , \new_[17640]_ , \new_[17641]_ , \new_[17642]_ ,
    \new_[17643]_ , \new_[17644]_ , \new_[17645]_ , \new_[17646]_ ,
    \new_[17647]_ , \new_[17648]_ , \new_[17649]_ , \new_[17650]_ ,
    \new_[17651]_ , \new_[17652]_ , \new_[17653]_ , \new_[17654]_ ,
    \new_[17655]_ , \new_[17656]_ , \new_[17657]_ , \new_[17658]_ ,
    \new_[17659]_ , \new_[17660]_ , \new_[17661]_ , \new_[17662]_ ,
    \new_[17663]_ , \new_[17664]_ , \new_[17665]_ , \new_[17666]_ ,
    \new_[17667]_ , \new_[17668]_ , \new_[17669]_ , \new_[17670]_ ,
    \new_[17671]_ , \new_[17672]_ , \new_[17673]_ , \new_[17674]_ ,
    \new_[17675]_ , \new_[17676]_ , \new_[17677]_ , \new_[17678]_ ,
    \new_[17679]_ , \new_[17680]_ , \new_[17681]_ , \new_[17682]_ ,
    \new_[17683]_ , \new_[17684]_ , \new_[17685]_ , \new_[17686]_ ,
    \new_[17687]_ , \new_[17688]_ , \new_[17689]_ , \new_[17690]_ ,
    \new_[17691]_ , \new_[17692]_ , \new_[17693]_ , \new_[17694]_ ,
    \new_[17695]_ , \new_[17696]_ , \new_[17697]_ , \new_[17698]_ ,
    \new_[17699]_ , \new_[17700]_ , \new_[17701]_ , \new_[17702]_ ,
    \new_[17703]_ , \new_[17704]_ , \new_[17705]_ , \new_[17706]_ ,
    \new_[17707]_ , \new_[17708]_ , \new_[17709]_ , \new_[17710]_ ,
    \new_[17711]_ , \new_[17712]_ , \new_[17713]_ , \new_[17714]_ ,
    \new_[17715]_ , \new_[17716]_ , \new_[17717]_ , \new_[17718]_ ,
    \new_[17719]_ , \new_[17720]_ , \new_[17721]_ , \new_[17722]_ ,
    \new_[17723]_ , \new_[17724]_ , \new_[17725]_ , \new_[17726]_ ,
    \new_[17727]_ , \new_[17728]_ , \new_[17729]_ , \new_[17730]_ ,
    \new_[17731]_ , \new_[17732]_ , \new_[17733]_ , \new_[17734]_ ,
    \new_[17735]_ , \new_[17736]_ , \new_[17737]_ , \new_[17738]_ ,
    \new_[17739]_ , \new_[17740]_ , \new_[17741]_ , \new_[17742]_ ,
    \new_[17743]_ , \new_[17744]_ , \new_[17745]_ , \new_[17746]_ ,
    \new_[17747]_ , \new_[17748]_ , \new_[17749]_ , \new_[17750]_ ,
    \new_[17751]_ , \new_[17752]_ , \new_[17753]_ , \new_[17754]_ ,
    \new_[17755]_ , \new_[17756]_ , \new_[17757]_ , \new_[17758]_ ,
    \new_[17759]_ , \new_[17760]_ , \new_[17761]_ , \new_[17762]_ ,
    \new_[17763]_ , \new_[17764]_ , \new_[17765]_ , \new_[17766]_ ,
    \new_[17767]_ , \new_[17768]_ , \new_[17769]_ , \new_[17770]_ ,
    \new_[17771]_ , \new_[17772]_ , \new_[17773]_ , \new_[17774]_ ,
    \new_[17775]_ , \new_[17776]_ , \new_[17777]_ , \new_[17778]_ ,
    \new_[17779]_ , \new_[17780]_ , \new_[17781]_ , \new_[17782]_ ,
    \new_[17783]_ , \new_[17784]_ , \new_[17785]_ , \new_[17786]_ ,
    \new_[17787]_ , \new_[17788]_ , \new_[17789]_ , \new_[17790]_ ,
    \new_[17791]_ , \new_[17792]_ , \new_[17793]_ , \new_[17794]_ ,
    \new_[17795]_ , \new_[17796]_ , \new_[17797]_ , \new_[17798]_ ,
    \new_[17799]_ , \new_[17800]_ , \new_[17801]_ , \new_[17802]_ ,
    \new_[17803]_ , \new_[17804]_ , \new_[17805]_ , \new_[17806]_ ,
    \new_[17807]_ , \new_[17808]_ , \new_[17809]_ , \new_[17810]_ ,
    \new_[17811]_ , \new_[17812]_ , \new_[17813]_ , \new_[17814]_ ,
    \new_[17815]_ , \new_[17816]_ , \new_[17817]_ , \new_[17818]_ ,
    \new_[17819]_ , \new_[17820]_ , \new_[17821]_ , \new_[17822]_ ,
    \new_[17823]_ , \new_[17824]_ , \new_[17825]_ , \new_[17826]_ ,
    \new_[17827]_ , \new_[17828]_ , \new_[17829]_ , \new_[17830]_ ,
    \new_[17831]_ , \new_[17832]_ , \new_[17833]_ , \new_[17834]_ ,
    \new_[17835]_ , \new_[17836]_ , \new_[17837]_ , \new_[17838]_ ,
    \new_[17839]_ , \new_[17840]_ , \new_[17841]_ , \new_[17842]_ ,
    \new_[17843]_ , \new_[17844]_ , \new_[17845]_ , \new_[17846]_ ,
    \new_[17847]_ , \new_[17848]_ , \new_[17849]_ , \new_[17850]_ ,
    \new_[17851]_ , \new_[17852]_ , \new_[17853]_ , \new_[17854]_ ,
    \new_[17855]_ , \new_[17856]_ , \new_[17857]_ , \new_[17858]_ ,
    \new_[17859]_ , \new_[17860]_ , \new_[17861]_ , \new_[17862]_ ,
    \new_[17863]_ , \new_[17864]_ , \new_[17865]_ , \new_[17866]_ ,
    \new_[17867]_ , \new_[17868]_ , \new_[17869]_ , \new_[17870]_ ,
    \new_[17871]_ , \new_[17872]_ , \new_[17873]_ , \new_[17874]_ ,
    \new_[17875]_ , \new_[17876]_ , \new_[17877]_ , \new_[17878]_ ,
    \new_[17879]_ , \new_[17880]_ , \new_[17881]_ , \new_[17882]_ ,
    \new_[17883]_ , \new_[17884]_ , \new_[17885]_ , \new_[17886]_ ,
    \new_[17887]_ , \new_[17888]_ , \new_[17889]_ , \new_[17890]_ ,
    \new_[17891]_ , \new_[17892]_ , \new_[17893]_ , \new_[17894]_ ,
    \new_[17895]_ , \new_[17896]_ , \new_[17897]_ , \new_[17898]_ ,
    \new_[17899]_ , \new_[17900]_ , \new_[17901]_ , \new_[17902]_ ,
    \new_[17903]_ , \new_[17904]_ , \new_[17905]_ , \new_[17906]_ ,
    \new_[17907]_ , \new_[17908]_ , \new_[17909]_ , \new_[17910]_ ,
    \new_[17911]_ , \new_[17912]_ , \new_[17913]_ , \new_[17914]_ ,
    \new_[17915]_ , \new_[17916]_ , \new_[17917]_ , \new_[17918]_ ,
    \new_[17919]_ , \new_[17920]_ , \new_[17921]_ , \new_[17922]_ ,
    \new_[17923]_ , \new_[17924]_ , \new_[17925]_ , \new_[17926]_ ,
    \new_[17927]_ , \new_[17928]_ , \new_[17929]_ , \new_[17930]_ ,
    \new_[17931]_ , \new_[17932]_ , \new_[17933]_ , \new_[17934]_ ,
    \new_[17935]_ , \new_[17936]_ , \new_[17937]_ , \new_[17938]_ ,
    \new_[17939]_ , \new_[17940]_ , \new_[17941]_ , \new_[17942]_ ,
    \new_[17943]_ , \new_[17944]_ , \new_[17945]_ , \new_[17946]_ ,
    \new_[17947]_ , \new_[17948]_ , \new_[17949]_ , \new_[17950]_ ,
    \new_[17951]_ , \new_[17952]_ , \new_[17953]_ , \new_[17954]_ ,
    \new_[17955]_ , \new_[17956]_ , \new_[17957]_ , \new_[17958]_ ,
    \new_[17959]_ , \new_[17960]_ , \new_[17961]_ , \new_[17962]_ ,
    \new_[17963]_ , \new_[17964]_ , \new_[17965]_ , \new_[17966]_ ,
    \new_[17967]_ , \new_[17968]_ , \new_[17969]_ , \new_[17970]_ ,
    \new_[17971]_ , \new_[17972]_ , \new_[17973]_ , \new_[17974]_ ,
    \new_[17975]_ , \new_[17976]_ , \new_[17977]_ , \new_[17978]_ ,
    \new_[17979]_ , \new_[17980]_ , \new_[17981]_ , \new_[17982]_ ,
    \new_[17983]_ , \new_[17984]_ , \new_[17985]_ , \new_[17986]_ ,
    \new_[17987]_ , \new_[17988]_ , \new_[17989]_ , \new_[17990]_ ,
    \new_[17991]_ , \new_[17992]_ , \new_[17993]_ , \new_[17994]_ ,
    \new_[17995]_ , \new_[17996]_ , \new_[17997]_ , \new_[17998]_ ,
    \new_[17999]_ , \new_[18000]_ , \new_[18001]_ , \new_[18002]_ ,
    \new_[18003]_ , \new_[18004]_ , \new_[18005]_ , \new_[18006]_ ,
    \new_[18007]_ , \new_[18008]_ , \new_[18009]_ , \new_[18010]_ ,
    \new_[18011]_ , \new_[18012]_ , \new_[18013]_ , \new_[18014]_ ,
    \new_[18015]_ , \new_[18016]_ , \new_[18017]_ , \new_[18018]_ ,
    \new_[18019]_ , \new_[18020]_ , \new_[18021]_ , \new_[18022]_ ,
    \new_[18023]_ , \new_[18024]_ , \new_[18025]_ , \new_[18026]_ ,
    \new_[18028]_ , \new_[18030]_ , \new_[18031]_ , \new_[18032]_ ,
    \new_[18033]_ , \new_[18034]_ , \new_[18035]_ , \new_[18036]_ ,
    \new_[18037]_ , \new_[18038]_ , \new_[18039]_ , \new_[18040]_ ,
    \new_[18041]_ , \new_[18042]_ , \new_[18043]_ , \new_[18044]_ ,
    \new_[18045]_ , \new_[18046]_ , \new_[18048]_ , \new_[18049]_ ,
    \new_[18050]_ , \new_[18051]_ , \new_[18053]_ , \new_[18054]_ ,
    \new_[18055]_ , \new_[18056]_ , \new_[18057]_ , \new_[18058]_ ,
    \new_[18059]_ , \new_[18060]_ , \new_[18061]_ , \new_[18062]_ ,
    \new_[18063]_ , \new_[18064]_ , \new_[18065]_ , \new_[18066]_ ,
    \new_[18067]_ , \new_[18068]_ , \new_[18069]_ , \new_[18070]_ ,
    \new_[18071]_ , \new_[18073]_ , \new_[18074]_ , \new_[18075]_ ,
    \new_[18076]_ , \new_[18077]_ , \new_[18078]_ , \new_[18079]_ ,
    \new_[18080]_ , \new_[18081]_ , \new_[18082]_ , \new_[18083]_ ,
    \new_[18084]_ , \new_[18085]_ , \new_[18086]_ , \new_[18087]_ ,
    \new_[18088]_ , \new_[18089]_ , \new_[18090]_ , \new_[18091]_ ,
    \new_[18092]_ , \new_[18093]_ , \new_[18094]_ , \new_[18095]_ ,
    \new_[18096]_ , \new_[18097]_ , \new_[18098]_ , \new_[18099]_ ,
    \new_[18100]_ , \new_[18101]_ , \new_[18102]_ , \new_[18103]_ ,
    \new_[18104]_ , \new_[18105]_ , \new_[18106]_ , \new_[18107]_ ,
    \new_[18108]_ , \new_[18109]_ , \new_[18110]_ , \new_[18111]_ ,
    \new_[18112]_ , \new_[18113]_ , \new_[18115]_ , \new_[18116]_ ,
    \new_[18117]_ , \new_[18118]_ , \new_[18119]_ , \new_[18120]_ ,
    \new_[18121]_ , \new_[18122]_ , \new_[18123]_ , \new_[18124]_ ,
    \new_[18126]_ , \new_[18127]_ , \new_[18128]_ , \new_[18129]_ ,
    \new_[18130]_ , \new_[18131]_ , \new_[18132]_ , \new_[18133]_ ,
    \new_[18134]_ , \new_[18135]_ , \new_[18136]_ , \new_[18137]_ ,
    \new_[18138]_ , \new_[18139]_ , \new_[18140]_ , \new_[18141]_ ,
    \new_[18142]_ , \new_[18143]_ , \new_[18144]_ , \new_[18145]_ ,
    \new_[18146]_ , \new_[18148]_ , \new_[18149]_ , \new_[18150]_ ,
    \new_[18151]_ , \new_[18153]_ , \new_[18154]_ , \new_[18155]_ ,
    \new_[18156]_ , \new_[18157]_ , \new_[18158]_ , \new_[18159]_ ,
    \new_[18160]_ , \new_[18161]_ , \new_[18163]_ , \new_[18164]_ ,
    \new_[18165]_ , \new_[18166]_ , \new_[18167]_ , \new_[18168]_ ,
    \new_[18169]_ , \new_[18170]_ , \new_[18171]_ , \new_[18172]_ ,
    \new_[18173]_ , \new_[18174]_ , \new_[18175]_ , \new_[18176]_ ,
    \new_[18177]_ , \new_[18178]_ , \new_[18179]_ , \new_[18180]_ ,
    \new_[18181]_ , \new_[18182]_ , \new_[18183]_ , \new_[18184]_ ,
    \new_[18185]_ , \new_[18186]_ , \new_[18187]_ , \new_[18188]_ ,
    \new_[18189]_ , \new_[18190]_ , \new_[18191]_ , \new_[18192]_ ,
    \new_[18193]_ , \new_[18194]_ , \new_[18195]_ , \new_[18196]_ ,
    \new_[18197]_ , \new_[18198]_ , \new_[18199]_ , \new_[18200]_ ,
    \new_[18201]_ , \new_[18203]_ , \new_[18204]_ , \new_[18205]_ ,
    \new_[18206]_ , \new_[18207]_ , \new_[18208]_ , \new_[18209]_ ,
    \new_[18210]_ , \new_[18211]_ , \new_[18212]_ , \new_[18214]_ ,
    \new_[18215]_ , \new_[18216]_ , \new_[18217]_ , \new_[18218]_ ,
    \new_[18219]_ , \new_[18220]_ , \new_[18221]_ , \new_[18222]_ ,
    \new_[18223]_ , \new_[18224]_ , \new_[18226]_ , \new_[18227]_ ,
    \new_[18228]_ , \new_[18229]_ , \new_[18230]_ , \new_[18231]_ ,
    \new_[18232]_ , \new_[18233]_ , \new_[18234]_ , \new_[18235]_ ,
    \new_[18236]_ , \new_[18237]_ , \new_[18238]_ , \new_[18239]_ ,
    \new_[18240]_ , \new_[18241]_ , \new_[18242]_ , \new_[18243]_ ,
    \new_[18244]_ , \new_[18245]_ , \new_[18246]_ , \new_[18247]_ ,
    \new_[18248]_ , \new_[18249]_ , \new_[18250]_ , \new_[18251]_ ,
    \new_[18252]_ , \new_[18253]_ , \new_[18254]_ , \new_[18255]_ ,
    \new_[18256]_ , \new_[18257]_ , \new_[18259]_ , \new_[18260]_ ,
    \new_[18261]_ , \new_[18262]_ , \new_[18263]_ , \new_[18264]_ ,
    \new_[18266]_ , \new_[18269]_ , \new_[18270]_ , \new_[18271]_ ,
    \new_[18273]_ , \new_[18274]_ , \new_[18275]_ , \new_[18276]_ ,
    \new_[18277]_ , \new_[18278]_ , \new_[18279]_ , \new_[18280]_ ,
    \new_[18281]_ , \new_[18282]_ , \new_[18283]_ , \new_[18284]_ ,
    \new_[18285]_ , \new_[18286]_ , \new_[18287]_ , \new_[18288]_ ,
    \new_[18289]_ , \new_[18292]_ , \new_[18293]_ , \new_[18294]_ ,
    \new_[18295]_ , \new_[18296]_ , \new_[18297]_ , \new_[18299]_ ,
    \new_[18300]_ , \new_[18301]_ , \new_[18302]_ , \new_[18303]_ ,
    \new_[18304]_ , \new_[18305]_ , \new_[18306]_ , \new_[18307]_ ,
    \new_[18308]_ , \new_[18309]_ , \new_[18310]_ , \new_[18311]_ ,
    \new_[18312]_ , \new_[18313]_ , \new_[18314]_ , \new_[18316]_ ,
    \new_[18317]_ , \new_[18319]_ , \new_[18320]_ , \new_[18321]_ ,
    \new_[18322]_ , \new_[18323]_ , \new_[18325]_ , \new_[18326]_ ,
    \new_[18327]_ , \new_[18328]_ , \new_[18329]_ , \new_[18330]_ ,
    \new_[18331]_ , \new_[18332]_ , \new_[18334]_ , \new_[18335]_ ,
    \new_[18336]_ , \new_[18337]_ , \new_[18338]_ , \new_[18339]_ ,
    \new_[18340]_ , \new_[18341]_ , \new_[18342]_ , \new_[18343]_ ,
    \new_[18344]_ , \new_[18345]_ , \new_[18346]_ , \new_[18347]_ ,
    \new_[18348]_ , \new_[18349]_ , \new_[18350]_ , \new_[18351]_ ,
    \new_[18352]_ , \new_[18353]_ , \new_[18354]_ , \new_[18355]_ ,
    \new_[18356]_ , \new_[18358]_ , \new_[18359]_ , \new_[18360]_ ,
    \new_[18361]_ , \new_[18362]_ , \new_[18363]_ , \new_[18365]_ ,
    \new_[18366]_ , \new_[18367]_ , \new_[18368]_ , \new_[18369]_ ,
    \new_[18370]_ , \new_[18371]_ , \new_[18372]_ , \new_[18373]_ ,
    \new_[18374]_ , \new_[18375]_ , \new_[18376]_ , \new_[18377]_ ,
    \new_[18378]_ , \new_[18379]_ , \new_[18380]_ , \new_[18381]_ ,
    \new_[18382]_ , \new_[18385]_ , \new_[18386]_ , \new_[18387]_ ,
    \new_[18388]_ , \new_[18389]_ , \new_[18390]_ , \new_[18391]_ ,
    \new_[18392]_ , \new_[18393]_ , \new_[18394]_ , \new_[18395]_ ,
    \new_[18396]_ , \new_[18397]_ , \new_[18398]_ , \new_[18399]_ ,
    \new_[18400]_ , \new_[18401]_ , \new_[18402]_ , \new_[18403]_ ,
    \new_[18404]_ , \new_[18405]_ , \new_[18406]_ , \new_[18408]_ ,
    \new_[18409]_ , \new_[18410]_ , \new_[18411]_ , \new_[18412]_ ,
    \new_[18413]_ , \new_[18414]_ , \new_[18415]_ , \new_[18416]_ ,
    \new_[18417]_ , \new_[18418]_ , \new_[18419]_ , \new_[18420]_ ,
    \new_[18421]_ , \new_[18422]_ , \new_[18423]_ , \new_[18424]_ ,
    \new_[18425]_ , \new_[18426]_ , \new_[18427]_ , \new_[18428]_ ,
    \new_[18429]_ , \new_[18430]_ , \new_[18431]_ , \new_[18432]_ ,
    \new_[18433]_ , \new_[18434]_ , \new_[18435]_ , \new_[18436]_ ,
    \new_[18437]_ , \new_[18439]_ , \new_[18440]_ , \new_[18442]_ ,
    \new_[18443]_ , \new_[18445]_ , \new_[18446]_ , \new_[18447]_ ,
    \new_[18448]_ , \new_[18449]_ , \new_[18450]_ , \new_[18451]_ ,
    \new_[18452]_ , \new_[18453]_ , \new_[18454]_ , \new_[18455]_ ,
    \new_[18456]_ , \new_[18457]_ , \new_[18458]_ , \new_[18459]_ ,
    \new_[18460]_ , \new_[18461]_ , \new_[18462]_ , \new_[18463]_ ,
    \new_[18464]_ , \new_[18465]_ , \new_[18466]_ , \new_[18467]_ ,
    \new_[18468]_ , \new_[18469]_ , \new_[18470]_ , \new_[18471]_ ,
    \new_[18472]_ , \new_[18473]_ , \new_[18474]_ , \new_[18475]_ ,
    \new_[18476]_ , \new_[18477]_ , \new_[18478]_ , \new_[18479]_ ,
    \new_[18480]_ , \new_[18481]_ , \new_[18482]_ , \new_[18483]_ ,
    \new_[18484]_ , \new_[18485]_ , \new_[18486]_ , \new_[18487]_ ,
    \new_[18489]_ , \new_[18490]_ , \new_[18491]_ , \new_[18492]_ ,
    \new_[18493]_ , \new_[18494]_ , \new_[18496]_ , \new_[18497]_ ,
    \new_[18498]_ , \new_[18499]_ , \new_[18500]_ , \new_[18501]_ ,
    \new_[18502]_ , \new_[18503]_ , \new_[18504]_ , \new_[18505]_ ,
    \new_[18506]_ , \new_[18507]_ , \new_[18508]_ , \new_[18509]_ ,
    \new_[18510]_ , \new_[18511]_ , \new_[18513]_ , \new_[18514]_ ,
    \new_[18516]_ , \new_[18517]_ , \new_[18518]_ , \new_[18519]_ ,
    \new_[18520]_ , \new_[18521]_ , \new_[18522]_ , \new_[18523]_ ,
    \new_[18524]_ , \new_[18525]_ , \new_[18526]_ , \new_[18527]_ ,
    \new_[18528]_ , \new_[18529]_ , \new_[18530]_ , \new_[18532]_ ,
    \new_[18533]_ , \new_[18535]_ , \new_[18536]_ , \new_[18537]_ ,
    \new_[18538]_ , \new_[18539]_ , \new_[18540]_ , \new_[18541]_ ,
    \new_[18542]_ , \new_[18543]_ , \new_[18544]_ , \new_[18545]_ ,
    \new_[18546]_ , \new_[18547]_ , \new_[18548]_ , \new_[18549]_ ,
    \new_[18551]_ , \new_[18552]_ , \new_[18553]_ , \new_[18554]_ ,
    \new_[18555]_ , \new_[18556]_ , \new_[18557]_ , \new_[18558]_ ,
    \new_[18559]_ , \new_[18560]_ , \new_[18561]_ , \new_[18562]_ ,
    \new_[18563]_ , \new_[18564]_ , \new_[18565]_ , \new_[18566]_ ,
    \new_[18567]_ , \new_[18568]_ , \new_[18569]_ , \new_[18570]_ ,
    \new_[18571]_ , \new_[18572]_ , \new_[18573]_ , \new_[18574]_ ,
    \new_[18575]_ , \new_[18576]_ , \new_[18577]_ , \new_[18578]_ ,
    \new_[18579]_ , \new_[18580]_ , \new_[18582]_ , \new_[18583]_ ,
    \new_[18584]_ , \new_[18585]_ , \new_[18586]_ , \new_[18587]_ ,
    \new_[18588]_ , \new_[18589]_ , \new_[18590]_ , \new_[18591]_ ,
    \new_[18592]_ , \new_[18593]_ , \new_[18594]_ , \new_[18595]_ ,
    \new_[18596]_ , \new_[18597]_ , \new_[18598]_ , \new_[18599]_ ,
    \new_[18600]_ , \new_[18601]_ , \new_[18602]_ , \new_[18603]_ ,
    \new_[18604]_ , \new_[18605]_ , \new_[18606]_ , \new_[18607]_ ,
    \new_[18608]_ , \new_[18609]_ , \new_[18610]_ , \new_[18611]_ ,
    \new_[18612]_ , \new_[18613]_ , \new_[18614]_ , \new_[18615]_ ,
    \new_[18616]_ , \new_[18617]_ , \new_[18618]_ , \new_[18619]_ ,
    \new_[18620]_ , \new_[18621]_ , \new_[18622]_ , \new_[18623]_ ,
    \new_[18624]_ , \new_[18625]_ , \new_[18626]_ , \new_[18627]_ ,
    \new_[18628]_ , \new_[18629]_ , \new_[18630]_ , \new_[18631]_ ,
    \new_[18632]_ , \new_[18633]_ , \new_[18634]_ , \new_[18635]_ ,
    \new_[18636]_ , \new_[18637]_ , \new_[18638]_ , \new_[18639]_ ,
    \new_[18640]_ , \new_[18641]_ , \new_[18642]_ , \new_[18643]_ ,
    \new_[18644]_ , \new_[18645]_ , \new_[18646]_ , \new_[18647]_ ,
    \new_[18648]_ , \new_[18649]_ , \new_[18650]_ , \new_[18651]_ ,
    \new_[18652]_ , \new_[18653]_ , \new_[18654]_ , \new_[18655]_ ,
    \new_[18656]_ , \new_[18657]_ , \new_[18658]_ , \new_[18659]_ ,
    \new_[18660]_ , \new_[18661]_ , \new_[18662]_ , \new_[18663]_ ,
    \new_[18664]_ , \new_[18665]_ , \new_[18666]_ , \new_[18667]_ ,
    \new_[18668]_ , \new_[18669]_ , \new_[18670]_ , \new_[18671]_ ,
    \new_[18672]_ , \new_[18673]_ , \new_[18674]_ , \new_[18675]_ ,
    \new_[18676]_ , \new_[18677]_ , \new_[18678]_ , \new_[18679]_ ,
    \new_[18680]_ , \new_[18681]_ , \new_[18682]_ , \new_[18683]_ ,
    \new_[18684]_ , \new_[18685]_ , \new_[18686]_ , \new_[18687]_ ,
    \new_[18688]_ , \new_[18689]_ , \new_[18690]_ , \new_[18691]_ ,
    \new_[18692]_ , \new_[18693]_ , \new_[18694]_ , \new_[18695]_ ,
    \new_[18696]_ , \new_[18697]_ , \new_[18698]_ , \new_[18699]_ ,
    \new_[18700]_ , \new_[18701]_ , \new_[18702]_ , \new_[18703]_ ,
    \new_[18704]_ , \new_[18705]_ , \new_[18706]_ , \new_[18707]_ ,
    \new_[18708]_ , \new_[18709]_ , \new_[18710]_ , \new_[18711]_ ,
    \new_[18712]_ , \new_[18713]_ , \new_[18714]_ , \new_[18715]_ ,
    \new_[18716]_ , \new_[18717]_ , \new_[18718]_ , \new_[18719]_ ,
    \new_[18720]_ , \new_[18721]_ , \new_[18722]_ , \new_[18723]_ ,
    \new_[18724]_ , \new_[18725]_ , \new_[18726]_ , \new_[18727]_ ,
    \new_[18728]_ , \new_[18729]_ , \new_[18730]_ , \new_[18731]_ ,
    \new_[18732]_ , \new_[18733]_ , \new_[18734]_ , \new_[18735]_ ,
    \new_[18736]_ , \new_[18737]_ , \new_[18738]_ , \new_[18739]_ ,
    \new_[18740]_ , \new_[18741]_ , \new_[18742]_ , \new_[18743]_ ,
    \new_[18744]_ , \new_[18745]_ , \new_[18746]_ , \new_[18747]_ ,
    \new_[18748]_ , \new_[18749]_ , \new_[18750]_ , \new_[18751]_ ,
    \new_[18752]_ , \new_[18753]_ , \new_[18754]_ , \new_[18755]_ ,
    \new_[18756]_ , \new_[18757]_ , \new_[18758]_ , \new_[18759]_ ,
    \new_[18760]_ , \new_[18761]_ , \new_[18762]_ , \new_[18763]_ ,
    \new_[18764]_ , \new_[18765]_ , \new_[18766]_ , \new_[18767]_ ,
    \new_[18768]_ , \new_[18769]_ , \new_[18770]_ , \new_[18771]_ ,
    \new_[18772]_ , \new_[18773]_ , \new_[18774]_ , \new_[18775]_ ,
    \new_[18776]_ , \new_[18777]_ , \new_[18778]_ , \new_[18779]_ ,
    \new_[18780]_ , \new_[18781]_ , \new_[18782]_ , \new_[18783]_ ,
    \new_[18784]_ , \new_[18785]_ , \new_[18786]_ , \new_[18787]_ ,
    \new_[18788]_ , \new_[18789]_ , \new_[18790]_ , \new_[18791]_ ,
    \new_[18792]_ , \new_[18793]_ , \new_[18794]_ , \new_[18795]_ ,
    \new_[18796]_ , \new_[18797]_ , \new_[18798]_ , \new_[18799]_ ,
    \new_[18800]_ , \new_[18801]_ , \new_[18802]_ , \new_[18803]_ ,
    \new_[18804]_ , \new_[18805]_ , \new_[18806]_ , \new_[18807]_ ,
    \new_[18808]_ , \new_[18809]_ , \new_[18810]_ , \new_[18811]_ ,
    \new_[18812]_ , \new_[18813]_ , \new_[18814]_ , \new_[18815]_ ,
    \new_[18816]_ , \new_[18817]_ , \new_[18818]_ , \new_[18819]_ ,
    \new_[18820]_ , \new_[18821]_ , \new_[18822]_ , \new_[18823]_ ,
    \new_[18824]_ , \new_[18825]_ , \new_[18826]_ , \new_[18827]_ ,
    \new_[18828]_ , \new_[18829]_ , \new_[18830]_ , \new_[18831]_ ,
    \new_[18832]_ , \new_[18833]_ , \new_[18834]_ , \new_[18835]_ ,
    \new_[18836]_ , \new_[18837]_ , \new_[18838]_ , \new_[18839]_ ,
    \new_[18840]_ , \new_[18841]_ , \new_[18842]_ , \new_[18843]_ ,
    \new_[18844]_ , \new_[18845]_ , \new_[18846]_ , \new_[18847]_ ,
    \new_[18848]_ , \new_[18849]_ , \new_[18850]_ , \new_[18851]_ ,
    \new_[18852]_ , \new_[18853]_ , \new_[18854]_ , \new_[18855]_ ,
    \new_[18856]_ , \new_[18857]_ , \new_[18858]_ , \new_[18859]_ ,
    \new_[18860]_ , \new_[18861]_ , \new_[18862]_ , \new_[18863]_ ,
    \new_[18864]_ , \new_[18865]_ , \new_[18866]_ , \new_[18867]_ ,
    \new_[18868]_ , \new_[18869]_ , \new_[18870]_ , \new_[18871]_ ,
    \new_[18872]_ , \new_[18873]_ , \new_[18874]_ , \new_[18875]_ ,
    \new_[18876]_ , \new_[18877]_ , \new_[18878]_ , \new_[18879]_ ,
    \new_[18880]_ , \new_[18881]_ , \new_[18882]_ , \new_[18883]_ ,
    \new_[18884]_ , \new_[18885]_ , \new_[18886]_ , \new_[18887]_ ,
    \new_[18888]_ , \new_[18889]_ , \new_[18890]_ , \new_[18891]_ ,
    \new_[18892]_ , \new_[18893]_ , \new_[18894]_ , \new_[18895]_ ,
    \new_[18896]_ , \new_[18897]_ , \new_[18898]_ , \new_[18899]_ ,
    \new_[18900]_ , \new_[18901]_ , \new_[18902]_ , \new_[18903]_ ,
    \new_[18904]_ , \new_[18905]_ , \new_[18906]_ , \new_[18907]_ ,
    \new_[18908]_ , \new_[18909]_ , \new_[18910]_ , \new_[18911]_ ,
    \new_[18912]_ , \new_[18913]_ , \new_[18914]_ , \new_[18915]_ ,
    \new_[18916]_ , \new_[18917]_ , \new_[18918]_ , \new_[18919]_ ,
    \new_[18920]_ , \new_[18921]_ , \new_[18922]_ , \new_[18923]_ ,
    \new_[18924]_ , \new_[18925]_ , \new_[18926]_ , \new_[18927]_ ,
    \new_[18928]_ , \new_[18929]_ , \new_[18930]_ , \new_[18931]_ ,
    \new_[18932]_ , \new_[18933]_ , \new_[18934]_ , \new_[18935]_ ,
    \new_[18936]_ , \new_[18937]_ , \new_[18938]_ , \new_[18939]_ ,
    \new_[18940]_ , \new_[18941]_ , \new_[18942]_ , \new_[18943]_ ,
    \new_[18944]_ , \new_[18945]_ , \new_[18946]_ , \new_[18947]_ ,
    \new_[18948]_ , \new_[18949]_ , \new_[18950]_ , \new_[18951]_ ,
    \new_[18952]_ , \new_[18953]_ , \new_[18954]_ , \new_[18955]_ ,
    \new_[18956]_ , \new_[18957]_ , \new_[18958]_ , \new_[18959]_ ,
    \new_[18960]_ , \new_[18961]_ , \new_[18962]_ , \new_[18963]_ ,
    \new_[18964]_ , \new_[18965]_ , \new_[18966]_ , \new_[18967]_ ,
    \new_[18968]_ , \new_[18969]_ , \new_[18970]_ , \new_[18971]_ ,
    \new_[18972]_ , \new_[18973]_ , \new_[18974]_ , \new_[18975]_ ,
    \new_[18976]_ , \new_[18978]_ , \new_[18979]_ , \new_[18980]_ ,
    \new_[18981]_ , \new_[18982]_ , \new_[18983]_ , \new_[18984]_ ,
    \new_[18986]_ , \new_[18987]_ , \new_[18988]_ , \new_[18989]_ ,
    \new_[18990]_ , \new_[18991]_ , \new_[18992]_ , \new_[18993]_ ,
    \new_[18994]_ , \new_[18995]_ , \new_[18996]_ , \new_[18997]_ ,
    \new_[18998]_ , \new_[18999]_ , \new_[19000]_ , \new_[19001]_ ,
    \new_[19002]_ , \new_[19003]_ , \new_[19004]_ , \new_[19005]_ ,
    \new_[19006]_ , \new_[19007]_ , \new_[19008]_ , \new_[19009]_ ,
    \new_[19010]_ , \new_[19011]_ , \new_[19012]_ , \new_[19013]_ ,
    \new_[19014]_ , \new_[19015]_ , \new_[19016]_ , \new_[19017]_ ,
    \new_[19018]_ , \new_[19019]_ , \new_[19020]_ , \new_[19021]_ ,
    \new_[19022]_ , \new_[19023]_ , \new_[19024]_ , \new_[19025]_ ,
    \new_[19026]_ , \new_[19027]_ , \new_[19028]_ , \new_[19029]_ ,
    \new_[19030]_ , \new_[19031]_ , \new_[19032]_ , \new_[19033]_ ,
    \new_[19034]_ , \new_[19035]_ , \new_[19036]_ , \new_[19037]_ ,
    \new_[19038]_ , \new_[19039]_ , \new_[19040]_ , \new_[19041]_ ,
    \new_[19042]_ , \new_[19043]_ , \new_[19044]_ , \new_[19045]_ ,
    \new_[19046]_ , \new_[19047]_ , \new_[19048]_ , \new_[19049]_ ,
    \new_[19050]_ , \new_[19051]_ , \new_[19052]_ , \new_[19053]_ ,
    \new_[19054]_ , \new_[19055]_ , \new_[19056]_ , \new_[19057]_ ,
    \new_[19058]_ , \new_[19059]_ , \new_[19060]_ , \new_[19061]_ ,
    \new_[19062]_ , \new_[19063]_ , \new_[19064]_ , \new_[19065]_ ,
    \new_[19066]_ , \new_[19067]_ , \new_[19068]_ , \new_[19069]_ ,
    \new_[19070]_ , \new_[19071]_ , \new_[19072]_ , \new_[19073]_ ,
    \new_[19074]_ , \new_[19075]_ , \new_[19076]_ , \new_[19077]_ ,
    \new_[19078]_ , \new_[19079]_ , \new_[19080]_ , \new_[19081]_ ,
    \new_[19082]_ , \new_[19083]_ , \new_[19084]_ , \new_[19085]_ ,
    \new_[19086]_ , \new_[19087]_ , \new_[19088]_ , \new_[19089]_ ,
    \new_[19090]_ , \new_[19091]_ , \new_[19092]_ , \new_[19093]_ ,
    \new_[19094]_ , \new_[19095]_ , \new_[19096]_ , \new_[19097]_ ,
    \new_[19098]_ , \new_[19099]_ , \new_[19100]_ , \new_[19101]_ ,
    \new_[19102]_ , \new_[19103]_ , \new_[19104]_ , \new_[19105]_ ,
    \new_[19106]_ , \new_[19107]_ , \new_[19108]_ , \new_[19109]_ ,
    \new_[19110]_ , \new_[19111]_ , \new_[19112]_ , \new_[19113]_ ,
    \new_[19114]_ , \new_[19115]_ , \new_[19116]_ , \new_[19117]_ ,
    \new_[19118]_ , \new_[19119]_ , \new_[19120]_ , \new_[19121]_ ,
    \new_[19122]_ , \new_[19123]_ , \new_[19124]_ , \new_[19125]_ ,
    \new_[19126]_ , \new_[19127]_ , \new_[19128]_ , \new_[19129]_ ,
    \new_[19130]_ , \new_[19131]_ , \new_[19132]_ , \new_[19133]_ ,
    \new_[19134]_ , \new_[19135]_ , \new_[19136]_ , \new_[19137]_ ,
    \new_[19138]_ , \new_[19139]_ , \new_[19140]_ , \new_[19141]_ ,
    \new_[19142]_ , \new_[19143]_ , \new_[19144]_ , \new_[19145]_ ,
    \new_[19146]_ , \new_[19147]_ , \new_[19148]_ , \new_[19149]_ ,
    \new_[19150]_ , \new_[19151]_ , \new_[19152]_ , \new_[19153]_ ,
    \new_[19154]_ , \new_[19155]_ , \new_[19156]_ , \new_[19157]_ ,
    \new_[19158]_ , \new_[19159]_ , \new_[19160]_ , \new_[19161]_ ,
    \new_[19162]_ , \new_[19163]_ , \new_[19164]_ , \new_[19165]_ ,
    \new_[19166]_ , \new_[19167]_ , \new_[19168]_ , \new_[19169]_ ,
    \new_[19170]_ , \new_[19171]_ , \new_[19172]_ , \new_[19173]_ ,
    \new_[19174]_ , \new_[19175]_ , \new_[19176]_ , \new_[19177]_ ,
    \new_[19178]_ , \new_[19179]_ , \new_[19180]_ , \new_[19181]_ ,
    \new_[19182]_ , \new_[19183]_ , \new_[19184]_ , \new_[19185]_ ,
    \new_[19186]_ , \new_[19187]_ , \new_[19188]_ , \new_[19189]_ ,
    \new_[19190]_ , \new_[19191]_ , \new_[19192]_ , \new_[19193]_ ,
    \new_[19194]_ , \new_[19195]_ , \new_[19196]_ , \new_[19197]_ ,
    \new_[19198]_ , \new_[19199]_ , \new_[19200]_ , \new_[19201]_ ,
    \new_[19202]_ , \new_[19203]_ , \new_[19204]_ , \new_[19205]_ ,
    \new_[19206]_ , \new_[19207]_ , \new_[19208]_ , \new_[19209]_ ,
    \new_[19210]_ , \new_[19211]_ , \new_[19212]_ , \new_[19213]_ ,
    \new_[19214]_ , \new_[19215]_ , \new_[19216]_ , \new_[19217]_ ,
    \new_[19218]_ , \new_[19219]_ , \new_[19220]_ , \new_[19221]_ ,
    \new_[19222]_ , \new_[19223]_ , \new_[19224]_ , \new_[19225]_ ,
    \new_[19226]_ , \new_[19227]_ , \new_[19228]_ , \new_[19229]_ ,
    \new_[19230]_ , \new_[19231]_ , \new_[19232]_ , \new_[19233]_ ,
    \new_[19234]_ , \new_[19235]_ , \new_[19236]_ , \new_[19237]_ ,
    \new_[19238]_ , \new_[19239]_ , \new_[19240]_ , \new_[19241]_ ,
    \new_[19242]_ , \new_[19243]_ , \new_[19244]_ , \new_[19245]_ ,
    \new_[19246]_ , \new_[19247]_ , \new_[19248]_ , \new_[19249]_ ,
    \new_[19250]_ , \new_[19251]_ , \new_[19252]_ , \new_[19253]_ ,
    \new_[19254]_ , \new_[19255]_ , \new_[19256]_ , \new_[19257]_ ,
    \new_[19258]_ , \new_[19259]_ , \new_[19260]_ , \new_[19261]_ ,
    \new_[19262]_ , \new_[19263]_ , \new_[19264]_ , \new_[19265]_ ,
    \new_[19266]_ , \new_[19267]_ , \new_[19268]_ , \new_[19269]_ ,
    \new_[19270]_ , \new_[19271]_ , \new_[19272]_ , \new_[19273]_ ,
    \new_[19274]_ , \new_[19275]_ , \new_[19276]_ , \new_[19277]_ ,
    \new_[19278]_ , \new_[19279]_ , \new_[19280]_ , \new_[19281]_ ,
    \new_[19282]_ , \new_[19283]_ , \new_[19284]_ , \new_[19285]_ ,
    \new_[19286]_ , \new_[19287]_ , \new_[19288]_ , \new_[19289]_ ,
    \new_[19290]_ , \new_[19291]_ , \new_[19292]_ , \new_[19293]_ ,
    \new_[19294]_ , \new_[19295]_ , \new_[19296]_ , \new_[19297]_ ,
    \new_[19298]_ , \new_[19299]_ , \new_[19300]_ , \new_[19301]_ ,
    \new_[19302]_ , \new_[19303]_ , \new_[19304]_ , \new_[19305]_ ,
    \new_[19306]_ , \new_[19307]_ , \new_[19308]_ , \new_[19309]_ ,
    \new_[19310]_ , \new_[19311]_ , \new_[19312]_ , \new_[19313]_ ,
    \new_[19314]_ , \new_[19315]_ , \new_[19316]_ , \new_[19317]_ ,
    \new_[19318]_ , \new_[19319]_ , \new_[19320]_ , \new_[19321]_ ,
    \new_[19322]_ , \new_[19323]_ , \new_[19324]_ , \new_[19325]_ ,
    \new_[19326]_ , \new_[19327]_ , \new_[19328]_ , \new_[19329]_ ,
    \new_[19330]_ , \new_[19331]_ , \new_[19332]_ , \new_[19333]_ ,
    \new_[19334]_ , \new_[19335]_ , \new_[19336]_ , \new_[19337]_ ,
    \new_[19338]_ , \new_[19339]_ , \new_[19340]_ , \new_[19341]_ ,
    \new_[19342]_ , \new_[19343]_ , \new_[19344]_ , \new_[19345]_ ,
    \new_[19346]_ , \new_[19347]_ , \new_[19348]_ , \new_[19349]_ ,
    \new_[19350]_ , \new_[19351]_ , \new_[19352]_ , \new_[19353]_ ,
    \new_[19354]_ , \new_[19355]_ , \new_[19356]_ , \new_[19357]_ ,
    \new_[19358]_ , \new_[19359]_ , \new_[19360]_ , \new_[19361]_ ,
    \new_[19362]_ , \new_[19363]_ , \new_[19364]_ , \new_[19365]_ ,
    \new_[19366]_ , \new_[19367]_ , \new_[19368]_ , \new_[19369]_ ,
    \new_[19370]_ , \new_[19371]_ , \new_[19372]_ , \new_[19373]_ ,
    \new_[19374]_ , \new_[19375]_ , \new_[19376]_ , \new_[19377]_ ,
    \new_[19378]_ , \new_[19379]_ , \new_[19380]_ , \new_[19381]_ ,
    \new_[19382]_ , \new_[19383]_ , \new_[19384]_ , \new_[19385]_ ,
    \new_[19386]_ , \new_[19387]_ , \new_[19388]_ , \new_[19389]_ ,
    \new_[19390]_ , \new_[19391]_ , \new_[19392]_ , \new_[19393]_ ,
    \new_[19394]_ , \new_[19395]_ , \new_[19396]_ , \new_[19397]_ ,
    \new_[19398]_ , \new_[19399]_ , \new_[19400]_ , \new_[19401]_ ,
    \new_[19402]_ , \new_[19403]_ , \new_[19404]_ , \new_[19405]_ ,
    \new_[19406]_ , \new_[19407]_ , \new_[19408]_ , \new_[19409]_ ,
    \new_[19410]_ , \new_[19411]_ , \new_[19412]_ , \new_[19413]_ ,
    \new_[19414]_ , \new_[19415]_ , \new_[19416]_ , \new_[19417]_ ,
    \new_[19418]_ , \new_[19419]_ , \new_[19420]_ , \new_[19421]_ ,
    \new_[19422]_ , \new_[19423]_ , \new_[19424]_ , \new_[19425]_ ,
    \new_[19426]_ , \new_[19427]_ , \new_[19428]_ , \new_[19429]_ ,
    \new_[19430]_ , \new_[19431]_ , \new_[19432]_ , \new_[19433]_ ,
    \new_[19434]_ , \new_[19435]_ , \new_[19436]_ , \new_[19437]_ ,
    \new_[19438]_ , \new_[19439]_ , \new_[19440]_ , \new_[19441]_ ,
    \new_[19442]_ , \new_[19443]_ , \new_[19444]_ , \new_[19445]_ ,
    \new_[19446]_ , \new_[19447]_ , \new_[19448]_ , \new_[19449]_ ,
    \new_[19450]_ , \new_[19451]_ , \new_[19452]_ , \new_[19453]_ ,
    \new_[19454]_ , \new_[19455]_ , \new_[19456]_ , \new_[19457]_ ,
    \new_[19459]_ , \new_[19460]_ , \new_[19461]_ , \new_[19462]_ ,
    \new_[19463]_ , \new_[19464]_ , \new_[19465]_ , \new_[19466]_ ,
    \new_[19467]_ , \new_[19468]_ , \new_[19469]_ , \new_[19470]_ ,
    \new_[19471]_ , \new_[19472]_ , \new_[19473]_ , \new_[19474]_ ,
    \new_[19475]_ , \new_[19476]_ , \new_[19477]_ , \new_[19478]_ ,
    \new_[19479]_ , \new_[19480]_ , \new_[19481]_ , \new_[19482]_ ,
    \new_[19483]_ , \new_[19484]_ , \new_[19485]_ , \new_[19486]_ ,
    \new_[19487]_ , \new_[19488]_ , \new_[19489]_ , \new_[19490]_ ,
    \new_[19491]_ , \new_[19492]_ , \new_[19493]_ , \new_[19494]_ ,
    \new_[19495]_ , \new_[19496]_ , \new_[19497]_ , \new_[19498]_ ,
    \new_[19499]_ , \new_[19500]_ , \new_[19501]_ , \new_[19502]_ ,
    \new_[19503]_ , \new_[19504]_ , \new_[19505]_ , \new_[19506]_ ,
    \new_[19507]_ , \new_[19508]_ , \new_[19509]_ , \new_[19510]_ ,
    \new_[19511]_ , \new_[19512]_ , \new_[19513]_ , \new_[19514]_ ,
    \new_[19515]_ , \new_[19516]_ , \new_[19517]_ , \new_[19518]_ ,
    \new_[19519]_ , \new_[19520]_ , \new_[19521]_ , \new_[19522]_ ,
    \new_[19523]_ , \new_[19524]_ , \new_[19525]_ , \new_[19526]_ ,
    \new_[19527]_ , \new_[19528]_ , \new_[19529]_ , \new_[19530]_ ,
    \new_[19531]_ , \new_[19532]_ , \new_[19533]_ , \new_[19534]_ ,
    \new_[19535]_ , \new_[19536]_ , \new_[19537]_ , \new_[19538]_ ,
    \new_[19539]_ , \new_[19540]_ , \new_[19541]_ , \new_[19542]_ ,
    \new_[19543]_ , \new_[19544]_ , \new_[19545]_ , \new_[19546]_ ,
    \new_[19547]_ , \new_[19548]_ , \new_[19549]_ , \new_[19550]_ ,
    \new_[19551]_ , \new_[19552]_ , \new_[19553]_ , \new_[19554]_ ,
    \new_[19555]_ , \new_[19556]_ , \new_[19557]_ , \new_[19558]_ ,
    \new_[19559]_ , \new_[19560]_ , \new_[19561]_ , \new_[19562]_ ,
    \new_[19563]_ , \new_[19564]_ , \new_[19565]_ , \new_[19566]_ ,
    \new_[19567]_ , \new_[19568]_ , \new_[19569]_ , \new_[19570]_ ,
    \new_[19571]_ , \new_[19572]_ , \new_[19573]_ , \new_[19574]_ ,
    \new_[19575]_ , \new_[19576]_ , \new_[19577]_ , \new_[19578]_ ,
    \new_[19579]_ , \new_[19580]_ , \new_[19581]_ , \new_[19582]_ ,
    \new_[19583]_ , \new_[19584]_ , \new_[19585]_ , \new_[19586]_ ,
    \new_[19587]_ , \new_[19588]_ , \new_[19589]_ , \new_[19590]_ ,
    \new_[19591]_ , \new_[19592]_ , \new_[19593]_ , \new_[19594]_ ,
    \new_[19595]_ , \new_[19596]_ , \new_[19597]_ , \new_[19598]_ ,
    \new_[19599]_ , \new_[19600]_ , \new_[19601]_ , \new_[19602]_ ,
    \new_[19603]_ , \new_[19604]_ , \new_[19605]_ , \new_[19606]_ ,
    \new_[19607]_ , \new_[19608]_ , \new_[19609]_ , \new_[19610]_ ,
    \new_[19611]_ , \new_[19612]_ , \new_[19613]_ , \new_[19614]_ ,
    \new_[19615]_ , \new_[19616]_ , \new_[19617]_ , \new_[19618]_ ,
    \new_[19619]_ , \new_[19620]_ , \new_[19621]_ , \new_[19622]_ ,
    \new_[19623]_ , \new_[19624]_ , \new_[19625]_ , \new_[19626]_ ,
    \new_[19627]_ , \new_[19628]_ , \new_[19629]_ , \new_[19630]_ ,
    \new_[19631]_ , \new_[19632]_ , \new_[19633]_ , \new_[19634]_ ,
    \new_[19635]_ , \new_[19636]_ , \new_[19637]_ , \new_[19638]_ ,
    \new_[19639]_ , \new_[19640]_ , \new_[19641]_ , \new_[19642]_ ,
    \new_[19643]_ , \new_[19644]_ , \new_[19645]_ , \new_[19646]_ ,
    \new_[19647]_ , \new_[19648]_ , \new_[19649]_ , \new_[19650]_ ,
    \new_[19651]_ , \new_[19652]_ , \new_[19653]_ , \new_[19654]_ ,
    \new_[19655]_ , \new_[19656]_ , \new_[19657]_ , \new_[19658]_ ,
    \new_[19659]_ , \new_[19660]_ , \new_[19661]_ , \new_[19662]_ ,
    \new_[19663]_ , \new_[19664]_ , \new_[19665]_ , \new_[19666]_ ,
    \new_[19667]_ , \new_[19668]_ , \new_[19669]_ , \new_[19670]_ ,
    \new_[19671]_ , \new_[19672]_ , \new_[19673]_ , \new_[19674]_ ,
    \new_[19675]_ , \new_[19676]_ , \new_[19677]_ , \new_[19678]_ ,
    \new_[19679]_ , \new_[19680]_ , \new_[19681]_ , \new_[19682]_ ,
    \new_[19683]_ , \new_[19684]_ , \new_[19685]_ , \new_[19686]_ ,
    \new_[19687]_ , \new_[19688]_ , \new_[19689]_ , \new_[19690]_ ,
    \new_[19691]_ , \new_[19692]_ , \new_[19693]_ , \new_[19694]_ ,
    \new_[19695]_ , \new_[19696]_ , \new_[19697]_ , \new_[19698]_ ,
    \new_[19699]_ , \new_[19700]_ , \new_[19701]_ , \new_[19702]_ ,
    \new_[19703]_ , \new_[19704]_ , \new_[19705]_ , \new_[19706]_ ,
    \new_[19707]_ , \new_[19708]_ , \new_[19709]_ , \new_[19710]_ ,
    \new_[19711]_ , \new_[19712]_ , \new_[19713]_ , \new_[19714]_ ,
    \new_[19715]_ , \new_[19716]_ , \new_[19717]_ , \new_[19718]_ ,
    \new_[19719]_ , \new_[19720]_ , \new_[19721]_ , \new_[19722]_ ,
    \new_[19723]_ , \new_[19724]_ , \new_[19725]_ , \new_[19726]_ ,
    \new_[19727]_ , \new_[19728]_ , \new_[19729]_ , \new_[19730]_ ,
    \new_[19731]_ , \new_[19732]_ , \new_[19733]_ , \new_[19734]_ ,
    \new_[19735]_ , \new_[19736]_ , \new_[19737]_ , \new_[19738]_ ,
    \new_[19739]_ , \new_[19740]_ , \new_[19741]_ , \new_[19742]_ ,
    \new_[19743]_ , \new_[19744]_ , \new_[19745]_ , \new_[19746]_ ,
    \new_[19747]_ , \new_[19748]_ , \new_[19749]_ , \new_[19750]_ ,
    \new_[19751]_ , \new_[19752]_ , \new_[19753]_ , \new_[19754]_ ,
    \new_[19755]_ , \new_[19756]_ , \new_[19757]_ , \new_[19758]_ ,
    \new_[19759]_ , \new_[19760]_ , \new_[19761]_ , \new_[19762]_ ,
    \new_[19763]_ , \new_[19764]_ , \new_[19765]_ , \new_[19766]_ ,
    \new_[19767]_ , \new_[19768]_ , \new_[19769]_ , \new_[19770]_ ,
    \new_[19771]_ , \new_[19772]_ , \new_[19773]_ , \new_[19774]_ ,
    \new_[19775]_ , \new_[19776]_ , \new_[19777]_ , \new_[19778]_ ,
    \new_[19779]_ , \new_[19780]_ , \new_[19781]_ , \new_[19782]_ ,
    \new_[19783]_ , \new_[19784]_ , \new_[19785]_ , \new_[19786]_ ,
    \new_[19787]_ , \new_[19788]_ , \new_[19789]_ , \new_[19790]_ ,
    \new_[19791]_ , \new_[19792]_ , \new_[19793]_ , \new_[19794]_ ,
    \new_[19795]_ , \new_[19796]_ , \new_[19797]_ , \new_[19798]_ ,
    \new_[19799]_ , \new_[19800]_ , \new_[19801]_ , \new_[19802]_ ,
    \new_[19803]_ , \new_[19804]_ , \new_[19805]_ , \new_[19806]_ ,
    \new_[19807]_ , \new_[19808]_ , \new_[19809]_ , \new_[19810]_ ,
    \new_[19811]_ , \new_[19812]_ , \new_[19813]_ , \new_[19814]_ ,
    \new_[19815]_ , \new_[19816]_ , \new_[19817]_ , \new_[19818]_ ,
    \new_[19819]_ , \new_[19820]_ , \new_[19821]_ , \new_[19822]_ ,
    \new_[19823]_ , \new_[19824]_ , \new_[19825]_ , \new_[19826]_ ,
    \new_[19827]_ , \new_[19828]_ , \new_[19829]_ , \new_[19830]_ ,
    \new_[19831]_ , \new_[19832]_ , \new_[19833]_ , \new_[19834]_ ,
    \new_[19835]_ , \new_[19836]_ , \new_[19837]_ , \new_[19838]_ ,
    \new_[19839]_ , \new_[19840]_ , \new_[19841]_ , \new_[19842]_ ,
    \new_[19843]_ , \new_[19844]_ , \new_[19845]_ , \new_[19846]_ ,
    \new_[19847]_ , \new_[19848]_ , \new_[19849]_ , \new_[19850]_ ,
    \new_[19851]_ , \new_[19852]_ , \new_[19853]_ , \new_[19854]_ ,
    \new_[19855]_ , \new_[19856]_ , \new_[19857]_ , \new_[19858]_ ,
    \new_[19859]_ , \new_[19860]_ , \new_[19861]_ , \new_[19862]_ ,
    \new_[19863]_ , \new_[19864]_ , \new_[19865]_ , \new_[19866]_ ,
    \new_[19867]_ , \new_[19868]_ , \new_[19869]_ , \new_[19871]_ ,
    \new_[19872]_ , \new_[19873]_ , \new_[19874]_ , \new_[19875]_ ,
    \new_[19876]_ , \new_[19877]_ , \new_[19878]_ , \new_[19879]_ ,
    \new_[19880]_ , \new_[19881]_ , \new_[19882]_ , \new_[19883]_ ,
    \new_[19884]_ , \new_[19885]_ , \new_[19886]_ , \new_[19887]_ ,
    \new_[19888]_ , \new_[19889]_ , \new_[19890]_ , \new_[19891]_ ,
    \new_[19892]_ , \new_[19893]_ , \new_[19894]_ , \new_[19895]_ ,
    \new_[19896]_ , \new_[19897]_ , \new_[19898]_ , \new_[19899]_ ,
    \new_[19900]_ , \new_[19901]_ , \new_[19902]_ , \new_[19903]_ ,
    \new_[19904]_ , \new_[19905]_ , \new_[19906]_ , \new_[19907]_ ,
    \new_[19908]_ , \new_[19909]_ , \new_[19910]_ , \new_[19911]_ ,
    \new_[19912]_ , \new_[19913]_ , \new_[19914]_ , \new_[19915]_ ,
    \new_[19916]_ , \new_[19917]_ , \new_[19918]_ , \new_[19919]_ ,
    \new_[19920]_ , \new_[19921]_ , \new_[19922]_ , \new_[19923]_ ,
    \new_[19924]_ , \new_[19925]_ , \new_[19926]_ , \new_[19927]_ ,
    \new_[19928]_ , \new_[19929]_ , \new_[19930]_ , \new_[19931]_ ,
    \new_[19932]_ , \new_[19933]_ , \new_[19934]_ , \new_[19935]_ ,
    \new_[19936]_ , \new_[19937]_ , \new_[19938]_ , \new_[19939]_ ,
    \new_[19940]_ , \new_[19941]_ , \new_[19942]_ , \new_[19943]_ ,
    \new_[19944]_ , \new_[19945]_ , \new_[19946]_ , \new_[19947]_ ,
    \new_[19948]_ , \new_[19949]_ , \new_[19950]_ , \new_[19951]_ ,
    \new_[19952]_ , \new_[19953]_ , \new_[19954]_ , \new_[19955]_ ,
    \new_[19956]_ , \new_[19957]_ , \new_[19958]_ , \new_[19959]_ ,
    \new_[19960]_ , \new_[19961]_ , \new_[19962]_ , \new_[19963]_ ,
    \new_[19964]_ , \new_[19965]_ , \new_[19966]_ , \new_[19967]_ ,
    \new_[19968]_ , \new_[19969]_ , \new_[19970]_ , \new_[19971]_ ,
    \new_[19972]_ , \new_[19973]_ , \new_[19974]_ , \new_[19975]_ ,
    \new_[19976]_ , \new_[19977]_ , \new_[19978]_ , \new_[19979]_ ,
    \new_[19980]_ , \new_[19981]_ , \new_[19982]_ , \new_[19983]_ ,
    \new_[19984]_ , \new_[19985]_ , \new_[19986]_ , \new_[19987]_ ,
    \new_[19988]_ , \new_[19989]_ , \new_[19990]_ , \new_[19991]_ ,
    \new_[19992]_ , \new_[19993]_ , \new_[19994]_ , \new_[19995]_ ,
    \new_[19996]_ , \new_[19997]_ , \new_[19998]_ , \new_[19999]_ ,
    \new_[20000]_ , \new_[20001]_ , \new_[20002]_ , \new_[20003]_ ,
    \new_[20004]_ , \new_[20005]_ , \new_[20006]_ , \new_[20007]_ ,
    \new_[20008]_ , \new_[20009]_ , \new_[20010]_ , \new_[20011]_ ,
    \new_[20012]_ , \new_[20013]_ , \new_[20014]_ , \new_[20015]_ ,
    \new_[20016]_ , \new_[20017]_ , \new_[20018]_ , \new_[20019]_ ,
    \new_[20020]_ , \new_[20021]_ , \new_[20022]_ , \new_[20023]_ ,
    \new_[20024]_ , \new_[20025]_ , \new_[20026]_ , \new_[20027]_ ,
    \new_[20028]_ , \new_[20029]_ , \new_[20030]_ , \new_[20031]_ ,
    \new_[20032]_ , \new_[20033]_ , \new_[20034]_ , \new_[20035]_ ,
    \new_[20036]_ , \new_[20037]_ , \new_[20038]_ , \new_[20039]_ ,
    \new_[20040]_ , \new_[20041]_ , \new_[20042]_ , \new_[20043]_ ,
    \new_[20044]_ , \new_[20045]_ , \new_[20046]_ , \new_[20047]_ ,
    \new_[20048]_ , \new_[20049]_ , \new_[20050]_ , \new_[20051]_ ,
    \new_[20052]_ , \new_[20053]_ , \new_[20054]_ , \new_[20055]_ ,
    \new_[20056]_ , \new_[20057]_ , \new_[20058]_ , \new_[20059]_ ,
    \new_[20060]_ , \new_[20061]_ , \new_[20062]_ , \new_[20063]_ ,
    \new_[20064]_ , \new_[20065]_ , \new_[20066]_ , \new_[20067]_ ,
    \new_[20068]_ , \new_[20069]_ , \new_[20070]_ , \new_[20071]_ ,
    \new_[20072]_ , \new_[20073]_ , \new_[20074]_ , \new_[20075]_ ,
    \new_[20076]_ , \new_[20077]_ , \new_[20078]_ , \new_[20079]_ ,
    \new_[20080]_ , \new_[20081]_ , \new_[20082]_ , \new_[20083]_ ,
    \new_[20084]_ , \new_[20085]_ , \new_[20086]_ , \new_[20087]_ ,
    \new_[20088]_ , \new_[20089]_ , \new_[20090]_ , \new_[20091]_ ,
    \new_[20092]_ , \new_[20093]_ , \new_[20094]_ , \new_[20095]_ ,
    \new_[20096]_ , \new_[20097]_ , \new_[20098]_ , \new_[20099]_ ,
    \new_[20100]_ , \new_[20101]_ , \new_[20102]_ , \new_[20103]_ ,
    \new_[20104]_ , \new_[20105]_ , \new_[20106]_ , \new_[20107]_ ,
    \new_[20108]_ , \new_[20109]_ , \new_[20110]_ , \new_[20111]_ ,
    \new_[20112]_ , \new_[20113]_ , \new_[20114]_ , \new_[20115]_ ,
    \new_[20116]_ , \new_[20117]_ , \new_[20118]_ , \new_[20119]_ ,
    \new_[20120]_ , \new_[20121]_ , \new_[20122]_ , \new_[20123]_ ,
    \new_[20124]_ , \new_[20125]_ , \new_[20126]_ , \new_[20127]_ ,
    \new_[20128]_ , \new_[20129]_ , \new_[20130]_ , \new_[20131]_ ,
    \new_[20132]_ , \new_[20133]_ , \new_[20134]_ , \new_[20135]_ ,
    \new_[20136]_ , \new_[20137]_ , \new_[20138]_ , \new_[20139]_ ,
    \new_[20140]_ , \new_[20141]_ , \new_[20142]_ , \new_[20143]_ ,
    \new_[20144]_ , \new_[20145]_ , \new_[20146]_ , \new_[20147]_ ,
    \new_[20148]_ , \new_[20149]_ , \new_[20150]_ , \new_[20151]_ ,
    \new_[20152]_ , \new_[20153]_ , \new_[20154]_ , \new_[20155]_ ,
    \new_[20156]_ , \new_[20157]_ , \new_[20158]_ , \new_[20159]_ ,
    \new_[20160]_ , \new_[20161]_ , \new_[20162]_ , \new_[20163]_ ,
    \new_[20164]_ , \new_[20165]_ , \new_[20166]_ , \new_[20167]_ ,
    \new_[20168]_ , \new_[20169]_ , \new_[20170]_ , \new_[20171]_ ,
    \new_[20172]_ , \new_[20173]_ , \new_[20174]_ , \new_[20175]_ ,
    \new_[20176]_ , \new_[20177]_ , \new_[20178]_ , \new_[20179]_ ,
    \new_[20180]_ , \new_[20181]_ , \new_[20182]_ , \new_[20183]_ ,
    \new_[20184]_ , \new_[20185]_ , \new_[20186]_ , \new_[20187]_ ,
    \new_[20188]_ , \new_[20189]_ , \new_[20190]_ , \new_[20191]_ ,
    \new_[20192]_ , \new_[20193]_ , \new_[20194]_ , \new_[20195]_ ,
    \new_[20196]_ , \new_[20197]_ , \new_[20198]_ , \new_[20199]_ ,
    \new_[20200]_ , \new_[20201]_ , \new_[20202]_ , \new_[20203]_ ,
    \new_[20204]_ , \new_[20205]_ , \new_[20206]_ , \new_[20207]_ ,
    \new_[20208]_ , \new_[20209]_ , \new_[20210]_ , \new_[20211]_ ,
    \new_[20212]_ , \new_[20213]_ , \new_[20214]_ , \new_[20215]_ ,
    \new_[20216]_ , \new_[20217]_ , \new_[20218]_ , \new_[20219]_ ,
    \new_[20220]_ , \new_[20221]_ , \new_[20222]_ , \new_[20223]_ ,
    \new_[20224]_ , \new_[20225]_ , \new_[20226]_ , \new_[20227]_ ,
    \new_[20228]_ , \new_[20229]_ , \new_[20230]_ , \new_[20231]_ ,
    \new_[20232]_ , \new_[20233]_ , \new_[20234]_ , \new_[20235]_ ,
    \new_[20236]_ , \new_[20237]_ , \new_[20238]_ , \new_[20239]_ ,
    \new_[20240]_ , \new_[20241]_ , \new_[20242]_ , \new_[20243]_ ,
    \new_[20244]_ , \new_[20245]_ , \new_[20246]_ , \new_[20247]_ ,
    \new_[20248]_ , \new_[20249]_ , \new_[20250]_ , \new_[20251]_ ,
    \new_[20252]_ , \new_[20253]_ , \new_[20254]_ , \new_[20255]_ ,
    \new_[20256]_ , \new_[20257]_ , \new_[20258]_ , \new_[20259]_ ,
    \new_[20260]_ , \new_[20261]_ , \new_[20262]_ , \new_[20263]_ ,
    \new_[20264]_ , \new_[20265]_ , \new_[20266]_ , \new_[20267]_ ,
    \new_[20268]_ , \new_[20269]_ , \new_[20270]_ , \new_[20271]_ ,
    \new_[20272]_ , \new_[20273]_ , \new_[20274]_ , \new_[20275]_ ,
    \new_[20276]_ , \new_[20277]_ , \new_[20278]_ , \new_[20279]_ ,
    \new_[20280]_ , \new_[20281]_ , \new_[20282]_ , \new_[20283]_ ,
    \new_[20284]_ , \new_[20285]_ , \new_[20286]_ , \new_[20287]_ ,
    \new_[20288]_ , \new_[20289]_ , \new_[20290]_ , \new_[20291]_ ,
    \new_[20292]_ , \new_[20293]_ , \new_[20294]_ , \new_[20295]_ ,
    \new_[20296]_ , \new_[20297]_ , \new_[20298]_ , \new_[20299]_ ,
    \new_[20300]_ , \new_[20301]_ , \new_[20302]_ , \new_[20303]_ ,
    \new_[20304]_ , \new_[20305]_ , \new_[20306]_ , \new_[20307]_ ,
    \new_[20308]_ , \new_[20309]_ , \new_[20310]_ , \new_[20311]_ ,
    \new_[20312]_ , \new_[20313]_ , \new_[20314]_ , \new_[20315]_ ,
    \new_[20316]_ , \new_[20317]_ , \new_[20318]_ , \new_[20319]_ ,
    \new_[20320]_ , \new_[20321]_ , \new_[20322]_ , \new_[20323]_ ,
    \new_[20324]_ , \new_[20325]_ , \new_[20326]_ , \new_[20327]_ ,
    \new_[20328]_ , \new_[20329]_ , \new_[20330]_ , \new_[20331]_ ,
    \new_[20332]_ , \new_[20333]_ , \new_[20334]_ , \new_[20335]_ ,
    \new_[20336]_ , \new_[20337]_ , \new_[20338]_ , \new_[20339]_ ,
    \new_[20340]_ , \new_[20341]_ , \new_[20342]_ , \new_[20343]_ ,
    \new_[20344]_ , \new_[20345]_ , \new_[20346]_ , \new_[20347]_ ,
    \new_[20348]_ , \new_[20349]_ , \new_[20350]_ , \new_[20351]_ ,
    \new_[20352]_ , \new_[20353]_ , \new_[20354]_ , \new_[20355]_ ,
    \new_[20356]_ , \new_[20357]_ , \new_[20358]_ , \new_[20359]_ ,
    \new_[20360]_ , \new_[20361]_ , \new_[20362]_ , \new_[20363]_ ,
    \new_[20364]_ , \new_[20365]_ , \new_[20366]_ , \new_[20367]_ ,
    \new_[20368]_ , \new_[20369]_ , \new_[20370]_ , \new_[20371]_ ,
    \new_[20372]_ , \new_[20373]_ , \new_[20374]_ , \new_[20375]_ ,
    \new_[20376]_ , \new_[20377]_ , \new_[20378]_ , \new_[20379]_ ,
    \new_[20380]_ , \new_[20381]_ , \new_[20382]_ , \new_[20383]_ ,
    \new_[20384]_ , \new_[20385]_ , \new_[20386]_ , \new_[20387]_ ,
    \new_[20388]_ , \new_[20389]_ , \new_[20390]_ , \new_[20391]_ ,
    \new_[20392]_ , \new_[20393]_ , \new_[20394]_ , \new_[20395]_ ,
    \new_[20396]_ , \new_[20397]_ , \new_[20398]_ , \new_[20399]_ ,
    \new_[20400]_ , \new_[20401]_ , \new_[20402]_ , \new_[20403]_ ,
    \new_[20404]_ , \new_[20405]_ , \new_[20406]_ , \new_[20407]_ ,
    \new_[20408]_ , \new_[20409]_ , \new_[20410]_ , \new_[20411]_ ,
    \new_[20412]_ , \new_[20413]_ , \new_[20414]_ , \new_[20415]_ ,
    \new_[20416]_ , \new_[20417]_ , \new_[20418]_ , \new_[20419]_ ,
    \new_[20420]_ , \new_[20421]_ , \new_[20422]_ , \new_[20423]_ ,
    \new_[20424]_ , \new_[20425]_ , \new_[20426]_ , \new_[20427]_ ,
    \new_[20428]_ , \new_[20429]_ , \new_[20430]_ , \new_[20431]_ ,
    \new_[20432]_ , \new_[20433]_ , \new_[20434]_ , \new_[20435]_ ,
    \new_[20436]_ , \new_[20437]_ , \new_[20438]_ , \new_[20439]_ ,
    \new_[20440]_ , \new_[20441]_ , \new_[20442]_ , \new_[20443]_ ,
    \new_[20444]_ , \new_[20445]_ , \new_[20446]_ , \new_[20447]_ ,
    \new_[20448]_ , \new_[20449]_ , \new_[20450]_ , \new_[20451]_ ,
    \new_[20452]_ , \new_[20453]_ , \new_[20454]_ , \new_[20455]_ ,
    \new_[20456]_ , \new_[20457]_ , \new_[20458]_ , \new_[20459]_ ,
    \new_[20460]_ , \new_[20461]_ , \new_[20462]_ , \new_[20463]_ ,
    \new_[20464]_ , \new_[20465]_ , \new_[20466]_ , \new_[20467]_ ,
    \new_[20468]_ , \new_[20469]_ , \new_[20470]_ , \new_[20471]_ ,
    \new_[20472]_ , \new_[20473]_ , \new_[20474]_ , \new_[20475]_ ,
    \new_[20476]_ , \new_[20477]_ , \new_[20478]_ , \new_[20479]_ ,
    \new_[20480]_ , \new_[20481]_ , \new_[20482]_ , \new_[20483]_ ,
    \new_[20484]_ , \new_[20485]_ , \new_[20486]_ , \new_[20487]_ ,
    \new_[20488]_ , \new_[20489]_ , \new_[20490]_ , \new_[20491]_ ,
    \new_[20492]_ , \new_[20493]_ , \new_[20494]_ , \new_[20495]_ ,
    \new_[20496]_ , \new_[20497]_ , \new_[20498]_ , \new_[20499]_ ,
    \new_[20500]_ , \new_[20501]_ , \new_[20502]_ , \new_[20503]_ ,
    \new_[20504]_ , \new_[20505]_ , \new_[20506]_ , \new_[20507]_ ,
    \new_[20508]_ , \new_[20509]_ , \new_[20510]_ , \new_[20511]_ ,
    \new_[20512]_ , \new_[20513]_ , \new_[20514]_ , \new_[20515]_ ,
    \new_[20516]_ , \new_[20517]_ , \new_[20518]_ , \new_[20519]_ ,
    \new_[20520]_ , \new_[20521]_ , \new_[20522]_ , \new_[20523]_ ,
    \new_[20524]_ , \new_[20525]_ , \new_[20526]_ , \new_[20527]_ ,
    \new_[20528]_ , \new_[20529]_ , \new_[20530]_ , \new_[20531]_ ,
    \new_[20532]_ , \new_[20533]_ , \new_[20534]_ , \new_[20535]_ ,
    \new_[20536]_ , \new_[20537]_ , \new_[20538]_ , \new_[20539]_ ,
    \new_[20540]_ , \new_[20541]_ , \new_[20542]_ , \new_[20543]_ ,
    \new_[20544]_ , \new_[20545]_ , \new_[20546]_ , \new_[20547]_ ,
    \new_[20548]_ , \new_[20549]_ , \new_[20550]_ , \new_[20551]_ ,
    \new_[20552]_ , \new_[20553]_ , \new_[20554]_ , \new_[20555]_ ,
    \new_[20556]_ , \new_[20557]_ , \new_[20558]_ , \new_[20559]_ ,
    \new_[20560]_ , \new_[20561]_ , \new_[20562]_ , \new_[20563]_ ,
    \new_[20564]_ , \new_[20565]_ , \new_[20566]_ , \new_[20567]_ ,
    \new_[20568]_ , \new_[20569]_ , \new_[20570]_ , \new_[20571]_ ,
    \new_[20572]_ , \new_[20573]_ , \new_[20574]_ , \new_[20575]_ ,
    \new_[20576]_ , \new_[20577]_ , \new_[20578]_ , \new_[20579]_ ,
    \new_[20580]_ , \new_[20581]_ , \new_[20582]_ , \new_[20583]_ ,
    \new_[20584]_ , \new_[20585]_ , \new_[20586]_ , \new_[20587]_ ,
    \new_[20588]_ , \new_[20589]_ , \new_[20590]_ , \new_[20591]_ ,
    \new_[20592]_ , \new_[20593]_ , \new_[20594]_ , \new_[20595]_ ,
    \new_[20596]_ , \new_[20597]_ , \new_[20598]_ , \new_[20599]_ ,
    \new_[20600]_ , \new_[20601]_ , \new_[20602]_ , \new_[20603]_ ,
    \new_[20604]_ , \new_[20605]_ , \new_[20606]_ , \new_[20607]_ ,
    \new_[20608]_ , \new_[20609]_ , \new_[20610]_ , \new_[20611]_ ,
    \new_[20612]_ , \new_[20613]_ , \new_[20614]_ , \new_[20615]_ ,
    \new_[20616]_ , \new_[20617]_ , \new_[20618]_ , \new_[20619]_ ,
    \new_[20620]_ , \new_[20621]_ , \new_[20622]_ , \new_[20623]_ ,
    \new_[20624]_ , \new_[20625]_ , \new_[20626]_ , \new_[20627]_ ,
    \new_[20628]_ , \new_[20629]_ , \new_[20630]_ , \new_[20631]_ ,
    \new_[20632]_ , \new_[20633]_ , \new_[20634]_ , \new_[20635]_ ,
    \new_[20636]_ , \new_[20637]_ , \new_[20638]_ , \new_[20639]_ ,
    \new_[20640]_ , \new_[20641]_ , \new_[20642]_ , \new_[20643]_ ,
    \new_[20644]_ , \new_[20645]_ , \new_[20646]_ , \new_[20647]_ ,
    \new_[20648]_ , \new_[20649]_ , \new_[20650]_ , \new_[20651]_ ,
    \new_[20652]_ , \new_[20653]_ , \new_[20654]_ , \new_[20655]_ ,
    \new_[20656]_ , \new_[20657]_ , \new_[20658]_ , \new_[20659]_ ,
    \new_[20660]_ , \new_[20661]_ , \new_[20662]_ , \new_[20663]_ ,
    \new_[20664]_ , \new_[20665]_ , \new_[20666]_ , \new_[20667]_ ,
    \new_[20668]_ , \new_[20669]_ , \new_[20670]_ , \new_[20671]_ ,
    \new_[20672]_ , \new_[20673]_ , \new_[20674]_ , \new_[20675]_ ,
    \new_[20676]_ , \new_[20677]_ , \new_[20678]_ , \new_[20679]_ ,
    \new_[20680]_ , \new_[20681]_ , \new_[20682]_ , \new_[20683]_ ,
    \new_[20684]_ , \new_[20685]_ , \new_[20686]_ , \new_[20687]_ ,
    \new_[20688]_ , \new_[20689]_ , \new_[20690]_ , \new_[20691]_ ,
    \new_[20692]_ , \new_[20693]_ , \new_[20694]_ , \new_[20695]_ ,
    \new_[20696]_ , \new_[20697]_ , \new_[20698]_ , \new_[20699]_ ,
    \new_[20700]_ , \new_[20701]_ , \new_[20702]_ , \new_[20703]_ ,
    \new_[20704]_ , \new_[20705]_ , \new_[20706]_ , \new_[20707]_ ,
    \new_[20708]_ , \new_[20709]_ , \new_[20710]_ , \new_[20711]_ ,
    \new_[20712]_ , \new_[20713]_ , \new_[20714]_ , \new_[20715]_ ,
    \new_[20716]_ , \new_[20717]_ , \new_[20718]_ , \new_[20719]_ ,
    \new_[20720]_ , \new_[20721]_ , \new_[20722]_ , \new_[20723]_ ,
    \new_[20724]_ , \new_[20725]_ , \new_[20726]_ , \new_[20727]_ ,
    \new_[20728]_ , \new_[20729]_ , \new_[20730]_ , \new_[20731]_ ,
    \new_[20732]_ , \new_[20733]_ , \new_[20734]_ , \new_[20735]_ ,
    \new_[20736]_ , \new_[20737]_ , \new_[20738]_ , \new_[20739]_ ,
    \new_[20740]_ , \new_[20741]_ , \new_[20742]_ , \new_[20743]_ ,
    \new_[20744]_ , \new_[20745]_ , \new_[20746]_ , \new_[20747]_ ,
    \new_[20748]_ , \new_[20749]_ , \new_[20750]_ , \new_[20751]_ ,
    \new_[20752]_ , \new_[20753]_ , \new_[20754]_ , \new_[20755]_ ,
    \new_[20756]_ , \new_[20757]_ , \new_[20758]_ , \new_[20759]_ ,
    \new_[20760]_ , \new_[20761]_ , \new_[20762]_ , \new_[20763]_ ,
    \new_[20764]_ , \new_[20765]_ , \new_[20766]_ , \new_[20767]_ ,
    \new_[20768]_ , \new_[20769]_ , \new_[20770]_ , \new_[20771]_ ,
    \new_[20772]_ , \new_[20773]_ , \new_[20774]_ , \new_[20775]_ ,
    \new_[20776]_ , \new_[20777]_ , \new_[20778]_ , \new_[20779]_ ,
    \new_[20780]_ , \new_[20781]_ , \new_[20782]_ , \new_[20783]_ ,
    \new_[20784]_ , \new_[20785]_ , \new_[20786]_ , \new_[20787]_ ,
    \new_[20788]_ , \new_[20789]_ , \new_[20790]_ , \new_[20791]_ ,
    \new_[20792]_ , \new_[20793]_ , \new_[20794]_ , \new_[20795]_ ,
    \new_[20796]_ , \new_[20797]_ , \new_[20798]_ , \new_[20799]_ ,
    \new_[20800]_ , \new_[20801]_ , \new_[20802]_ , \new_[20803]_ ,
    \new_[20804]_ , \new_[20805]_ , \new_[20806]_ , \new_[20807]_ ,
    \new_[20808]_ , \new_[20809]_ , \new_[20810]_ , \new_[20811]_ ,
    \new_[20812]_ , \new_[20813]_ , \new_[20814]_ , \new_[20815]_ ,
    \new_[20816]_ , \new_[20817]_ , \new_[20818]_ , \new_[20819]_ ,
    \new_[20820]_ , \new_[20821]_ , \new_[20822]_ , \new_[20823]_ ,
    \new_[20824]_ , \new_[20825]_ , \new_[20826]_ , \new_[20827]_ ,
    \new_[20828]_ , \new_[20829]_ , \new_[20830]_ , \new_[20831]_ ,
    \new_[20832]_ , \new_[20833]_ , \new_[20834]_ , \new_[20835]_ ,
    \new_[20836]_ , \new_[20837]_ , \new_[20838]_ , \new_[20839]_ ,
    \new_[20840]_ , \new_[20841]_ , \new_[20842]_ , \new_[20843]_ ,
    \new_[20844]_ , \new_[20845]_ , \new_[20846]_ , \new_[20847]_ ,
    \new_[20848]_ , \new_[20849]_ , \new_[20850]_ , \new_[20851]_ ,
    \new_[20852]_ , \new_[20853]_ , \new_[20854]_ , \new_[20855]_ ,
    \new_[20856]_ , \new_[20857]_ , \new_[20858]_ , \new_[20859]_ ,
    \new_[20860]_ , \new_[20861]_ , \new_[20862]_ , \new_[20863]_ ,
    \new_[20864]_ , \new_[20865]_ , \new_[20866]_ , \new_[20867]_ ,
    \new_[20868]_ , \new_[20869]_ , \new_[20870]_ , \new_[20871]_ ,
    \new_[20872]_ , \new_[20873]_ , \new_[20874]_ , \new_[20875]_ ,
    \new_[20876]_ , \new_[20877]_ , \new_[20878]_ , \new_[20879]_ ,
    \new_[20880]_ , \new_[20881]_ , \new_[20882]_ , \new_[20883]_ ,
    \new_[20884]_ , \new_[20885]_ , \new_[20886]_ , \new_[20887]_ ,
    \new_[20888]_ , \new_[20889]_ , \new_[20890]_ , \new_[20891]_ ,
    \new_[20892]_ , \new_[20893]_ , \new_[20894]_ , \new_[20895]_ ,
    \new_[20896]_ , \new_[20897]_ , \new_[20898]_ , \new_[20899]_ ,
    \new_[20900]_ , \new_[20901]_ , \new_[20902]_ , \new_[20903]_ ,
    \new_[20904]_ , \new_[20905]_ , \new_[20906]_ , \new_[20907]_ ,
    \new_[20908]_ , \new_[20909]_ , \new_[20910]_ , \new_[20911]_ ,
    \new_[20912]_ , \new_[20913]_ , \new_[20914]_ , \new_[20915]_ ,
    \new_[20916]_ , \new_[20917]_ , \new_[20918]_ , \new_[20919]_ ,
    \new_[20920]_ , \new_[20921]_ , \new_[20922]_ , \new_[20923]_ ,
    \new_[20924]_ , \new_[20925]_ , \new_[20926]_ , \new_[20927]_ ,
    \new_[20928]_ , \new_[20929]_ , \new_[20930]_ , \new_[20931]_ ,
    \new_[20932]_ , \new_[20933]_ , \new_[20934]_ , \new_[20935]_ ,
    \new_[20936]_ , \new_[20937]_ , \new_[20938]_ , \new_[20939]_ ,
    \new_[20940]_ , \new_[20941]_ , \new_[20942]_ , \new_[20943]_ ,
    \new_[20944]_ , \new_[20945]_ , \new_[20946]_ , \new_[20947]_ ,
    \new_[20948]_ , \new_[20949]_ , \new_[20950]_ , \new_[20951]_ ,
    \new_[20952]_ , \new_[20953]_ , \new_[20954]_ , \new_[20955]_ ,
    \new_[20956]_ , \new_[20957]_ , \new_[20958]_ , \new_[20959]_ ,
    \new_[20960]_ , \new_[20961]_ , \new_[20962]_ , \new_[20963]_ ,
    \new_[20964]_ , \new_[20965]_ , \new_[20966]_ , \new_[20967]_ ,
    \new_[20968]_ , \new_[20969]_ , \new_[20970]_ , \new_[20971]_ ,
    \new_[20972]_ , \new_[20973]_ , \new_[20974]_ , \new_[20975]_ ,
    \new_[20976]_ , \new_[20977]_ , \new_[20978]_ , \new_[20979]_ ,
    \new_[20980]_ , \new_[20981]_ , \new_[20982]_ , \new_[20983]_ ,
    \new_[20984]_ , \new_[20985]_ , \new_[20986]_ , \new_[20987]_ ,
    \new_[20988]_ , \new_[20989]_ , \new_[20990]_ , \new_[20991]_ ,
    \new_[20992]_ , \new_[20993]_ , \new_[20994]_ , \new_[20995]_ ,
    \new_[20996]_ , \new_[20997]_ , \new_[20998]_ , \new_[20999]_ ,
    \new_[21000]_ , \new_[21001]_ , \new_[21002]_ , \new_[21003]_ ,
    \new_[21004]_ , \new_[21005]_ , \new_[21006]_ , \new_[21007]_ ,
    \new_[21008]_ , \new_[21009]_ , \new_[21010]_ , \new_[21011]_ ,
    \new_[21012]_ , \new_[21013]_ , \new_[21014]_ , \new_[21015]_ ,
    \new_[21016]_ , \new_[21017]_ , \new_[21018]_ , \new_[21019]_ ,
    \new_[21020]_ , \new_[21021]_ , \new_[21022]_ , \new_[21023]_ ,
    \new_[21024]_ , \new_[21025]_ , \new_[21026]_ , \new_[21027]_ ,
    \new_[21028]_ , \new_[21029]_ , \new_[21030]_ , \new_[21031]_ ,
    \new_[21032]_ , \new_[21033]_ , \new_[21034]_ , \new_[21035]_ ,
    \new_[21036]_ , \new_[21037]_ , \new_[21038]_ , \new_[21039]_ ,
    \new_[21040]_ , \new_[21041]_ , \new_[21042]_ , \new_[21043]_ ,
    \new_[21044]_ , \new_[21045]_ , \new_[21046]_ , \new_[21047]_ ,
    \new_[21048]_ , \new_[21049]_ , \new_[21050]_ , \new_[21051]_ ,
    \new_[21052]_ , \new_[21053]_ , \new_[21054]_ , \new_[21055]_ ,
    \new_[21056]_ , \new_[21057]_ , \new_[21058]_ , \new_[21059]_ ,
    \new_[21060]_ , \new_[21061]_ , \new_[21062]_ , \new_[21063]_ ,
    \new_[21064]_ , \new_[21065]_ , \new_[21066]_ , \new_[21067]_ ,
    \new_[21068]_ , \new_[21069]_ , \new_[21070]_ , \new_[21071]_ ,
    \new_[21072]_ , \new_[21073]_ , \new_[21074]_ , \new_[21075]_ ,
    \new_[21076]_ , \new_[21077]_ , \new_[21078]_ , \new_[21079]_ ,
    \new_[21080]_ , \new_[21081]_ , \new_[21082]_ , \new_[21083]_ ,
    \new_[21084]_ , \new_[21085]_ , \new_[21086]_ , \new_[21087]_ ,
    \new_[21088]_ , \new_[21089]_ , \new_[21090]_ , \new_[21091]_ ,
    \new_[21092]_ , \new_[21093]_ , \new_[21094]_ , \new_[21095]_ ,
    \new_[21096]_ , \new_[21097]_ , \new_[21098]_ , \new_[21099]_ ,
    \new_[21100]_ , \new_[21101]_ , \new_[21102]_ , \new_[21103]_ ,
    \new_[21104]_ , \new_[21105]_ , \new_[21106]_ , \new_[21107]_ ,
    \new_[21108]_ , \new_[21109]_ , \new_[21110]_ , \new_[21111]_ ,
    \new_[21112]_ , \new_[21113]_ , \new_[21114]_ , \new_[21115]_ ,
    \new_[21116]_ , \new_[21117]_ , \new_[21118]_ , \new_[21119]_ ,
    \new_[21120]_ , \new_[21121]_ , \new_[21122]_ , \new_[21123]_ ,
    \new_[21124]_ , \new_[21125]_ , \new_[21126]_ , \new_[21127]_ ,
    \new_[21128]_ , \new_[21129]_ , \new_[21130]_ , \new_[21131]_ ,
    \new_[21132]_ , \new_[21133]_ , \new_[21134]_ , \new_[21135]_ ,
    \new_[21136]_ , \new_[21137]_ , \new_[21138]_ , \new_[21139]_ ,
    \new_[21140]_ , \new_[21141]_ , \new_[21142]_ , \new_[21143]_ ,
    \new_[21144]_ , \new_[21145]_ , \new_[21146]_ , \new_[21147]_ ,
    \new_[21148]_ , \new_[21149]_ , \new_[21150]_ , \new_[21151]_ ,
    \new_[21152]_ , \new_[21153]_ , \new_[21154]_ , \new_[21155]_ ,
    \new_[21156]_ , \new_[21157]_ , \new_[21158]_ , \new_[21159]_ ,
    \new_[21160]_ , \new_[21161]_ , \new_[21162]_ , \new_[21163]_ ,
    \new_[21164]_ , \new_[21165]_ , \new_[21166]_ , \new_[21167]_ ,
    \new_[21168]_ , \new_[21169]_ , \new_[21170]_ , \new_[21171]_ ,
    \new_[21172]_ , \new_[21173]_ , \new_[21174]_ , \new_[21175]_ ,
    \new_[21176]_ , \new_[21177]_ , \new_[21178]_ , \new_[21179]_ ,
    \new_[21180]_ , \new_[21181]_ , \new_[21182]_ , \new_[21183]_ ,
    \new_[21184]_ , \new_[21185]_ , \new_[21186]_ , \new_[21187]_ ,
    \new_[21188]_ , \new_[21189]_ , \new_[21190]_ , \new_[21191]_ ,
    \new_[21192]_ , \new_[21193]_ , \new_[21194]_ , \new_[21195]_ ,
    \new_[21196]_ , \new_[21197]_ , \new_[21198]_ , \new_[21199]_ ,
    \new_[21200]_ , \new_[21201]_ , \new_[21202]_ , \new_[21203]_ ,
    \new_[21204]_ , \new_[21205]_ , \new_[21206]_ , \new_[21207]_ ,
    \new_[21208]_ , \new_[21209]_ , \new_[21210]_ , \new_[21211]_ ,
    \new_[21212]_ , \new_[21213]_ , \new_[21214]_ , \new_[21215]_ ,
    \new_[21216]_ , \new_[21217]_ , \new_[21218]_ , \new_[21219]_ ,
    \new_[21220]_ , \new_[21221]_ , \new_[21222]_ , \new_[21223]_ ,
    \new_[21224]_ , \new_[21225]_ , \new_[21226]_ , \new_[21227]_ ,
    \new_[21228]_ , \new_[21229]_ , \new_[21230]_ , \new_[21231]_ ,
    \new_[21232]_ , \new_[21233]_ , \new_[21234]_ , \new_[21235]_ ,
    \new_[21236]_ , \new_[21237]_ , \new_[21238]_ , \new_[21239]_ ,
    \new_[21240]_ , \new_[21241]_ , \new_[21242]_ , \new_[21244]_ ,
    \new_[21245]_ , \new_[21246]_ , \new_[21247]_ , \new_[21248]_ ,
    \new_[21249]_ , \new_[21250]_ , \new_[21251]_ , \new_[21252]_ ,
    \new_[21253]_ , \new_[21254]_ , \new_[21255]_ , \new_[21256]_ ,
    \new_[21257]_ , \new_[21258]_ , \new_[21259]_ , \new_[21260]_ ,
    \new_[21261]_ , \new_[21262]_ , \new_[21263]_ , \new_[21264]_ ,
    \new_[21265]_ , \new_[21266]_ , \new_[21267]_ , \new_[21268]_ ,
    \new_[21269]_ , \new_[21270]_ , \new_[21271]_ , \new_[21272]_ ,
    \new_[21273]_ , \new_[21274]_ , \new_[21275]_ , \new_[21276]_ ,
    \new_[21277]_ , \new_[21278]_ , \new_[21279]_ , \new_[21280]_ ,
    \new_[21281]_ , \new_[21282]_ , \new_[21283]_ , \new_[21284]_ ,
    \new_[21285]_ , \new_[21286]_ , \new_[21287]_ , \new_[21288]_ ,
    \new_[21289]_ , \new_[21290]_ , \new_[21291]_ , \new_[21292]_ ,
    \new_[21293]_ , \new_[21294]_ , \new_[21295]_ , \new_[21296]_ ,
    \new_[21297]_ , \new_[21298]_ , \new_[21299]_ , \new_[21300]_ ,
    \new_[21301]_ , \new_[21302]_ , \new_[21303]_ , \new_[21304]_ ,
    \new_[21305]_ , \new_[21306]_ , \new_[21307]_ , \new_[21308]_ ,
    \new_[21309]_ , \new_[21310]_ , \new_[21311]_ , \new_[21312]_ ,
    \new_[21313]_ , \new_[21314]_ , \new_[21315]_ , \new_[21316]_ ,
    \new_[21317]_ , \new_[21318]_ , \new_[21319]_ , \new_[21320]_ ,
    \new_[21321]_ , \new_[21322]_ , \new_[21323]_ , \new_[21324]_ ,
    \new_[21325]_ , \new_[21326]_ , \new_[21327]_ , \new_[21328]_ ,
    \new_[21329]_ , \new_[21330]_ , \new_[21331]_ , \new_[21332]_ ,
    \new_[21333]_ , \new_[21334]_ , \new_[21335]_ , \new_[21336]_ ,
    \new_[21337]_ , \new_[21338]_ , \new_[21339]_ , \new_[21340]_ ,
    \new_[21341]_ , \new_[21342]_ , \new_[21343]_ , \new_[21344]_ ,
    \new_[21345]_ , \new_[21346]_ , \new_[21347]_ , \new_[21348]_ ,
    \new_[21349]_ , \new_[21350]_ , \new_[21351]_ , \new_[21352]_ ,
    \new_[21353]_ , \new_[21354]_ , \new_[21355]_ , \new_[21356]_ ,
    \new_[21357]_ , \new_[21358]_ , \new_[21359]_ , \new_[21360]_ ,
    \new_[21361]_ , \new_[21362]_ , \new_[21363]_ , \new_[21364]_ ,
    \new_[21365]_ , \new_[21366]_ , \new_[21367]_ , \new_[21368]_ ,
    \new_[21369]_ , \new_[21370]_ , \new_[21371]_ , \new_[21372]_ ,
    \new_[21373]_ , \new_[21374]_ , \new_[21375]_ , \new_[21376]_ ,
    \new_[21377]_ , \new_[21378]_ , \new_[21379]_ , \new_[21380]_ ,
    \new_[21381]_ , \new_[21382]_ , \new_[21383]_ , \new_[21384]_ ,
    \new_[21385]_ , \new_[21386]_ , \new_[21387]_ , \new_[21388]_ ,
    \new_[21389]_ , \new_[21390]_ , \new_[21391]_ , \new_[21392]_ ,
    \new_[21393]_ , \new_[21394]_ , \new_[21395]_ , \new_[21396]_ ,
    \new_[21397]_ , \new_[21398]_ , \new_[21399]_ , \new_[21400]_ ,
    \new_[21401]_ , \new_[21402]_ , \new_[21403]_ , \new_[21404]_ ,
    \new_[21405]_ , \new_[21406]_ , \new_[21407]_ , \new_[21408]_ ,
    \new_[21409]_ , \new_[21410]_ , \new_[21411]_ , \new_[21412]_ ,
    \new_[21413]_ , \new_[21414]_ , \new_[21415]_ , \new_[21416]_ ,
    \new_[21417]_ , \new_[21418]_ , \new_[21419]_ , \new_[21420]_ ,
    \new_[21421]_ , \new_[21422]_ , \new_[21423]_ , \new_[21424]_ ,
    \new_[21425]_ , \new_[21426]_ , \new_[21427]_ , \new_[21428]_ ,
    \new_[21429]_ , \new_[21430]_ , \new_[21431]_ , \new_[21432]_ ,
    \new_[21433]_ , \new_[21434]_ , \new_[21435]_ , \new_[21436]_ ,
    \new_[21437]_ , \new_[21438]_ , \new_[21439]_ , \new_[21440]_ ,
    \new_[21441]_ , \new_[21442]_ , \new_[21443]_ , \new_[21444]_ ,
    \new_[21445]_ , \new_[21446]_ , \new_[21447]_ , \new_[21448]_ ,
    \new_[21449]_ , \new_[21450]_ , \new_[21451]_ , \new_[21452]_ ,
    \new_[21453]_ , \new_[21454]_ , \new_[21455]_ , \new_[21456]_ ,
    \new_[21457]_ , \new_[21458]_ , \new_[21459]_ , \new_[21460]_ ,
    \new_[21461]_ , \new_[21462]_ , \new_[21463]_ , \new_[21464]_ ,
    \new_[21465]_ , \new_[21466]_ , \new_[21467]_ , \new_[21468]_ ,
    \new_[21469]_ , \new_[21470]_ , \new_[21471]_ , \new_[21472]_ ,
    \new_[21473]_ , \new_[21474]_ , \new_[21475]_ , \new_[21476]_ ,
    \new_[21477]_ , \new_[21478]_ , \new_[21479]_ , \new_[21480]_ ,
    \new_[21481]_ , \new_[21482]_ , \new_[21483]_ , \new_[21484]_ ,
    \new_[21485]_ , \new_[21486]_ , \new_[21487]_ , \new_[21488]_ ,
    \new_[21489]_ , \new_[21490]_ , \new_[21491]_ , \new_[21492]_ ,
    \new_[21493]_ , \new_[21494]_ , \new_[21495]_ , \new_[21496]_ ,
    \new_[21497]_ , \new_[21498]_ , \new_[21499]_ , \new_[21500]_ ,
    \new_[21501]_ , \new_[21502]_ , \new_[21503]_ , \new_[21504]_ ,
    \new_[21505]_ , \new_[21506]_ , \new_[21507]_ , \new_[21508]_ ,
    \new_[21509]_ , \new_[21510]_ , \new_[21511]_ , \new_[21512]_ ,
    \new_[21513]_ , \new_[21514]_ , \new_[21515]_ , \new_[21516]_ ,
    \new_[21517]_ , \new_[21518]_ , \new_[21519]_ , \new_[21520]_ ,
    \new_[21521]_ , \new_[21522]_ , \new_[21523]_ , \new_[21524]_ ,
    \new_[21525]_ , \new_[21526]_ , \new_[21527]_ , \new_[21528]_ ,
    \new_[21529]_ , \new_[21530]_ , \new_[21531]_ , \new_[21532]_ ,
    \new_[21533]_ , \new_[21534]_ , \new_[21535]_ , \new_[21536]_ ,
    \new_[21537]_ , \new_[21538]_ , \new_[21539]_ , \new_[21540]_ ,
    \new_[21541]_ , \new_[21542]_ , \new_[21543]_ , \new_[21544]_ ,
    \new_[21545]_ , \new_[21546]_ , \new_[21547]_ , \new_[21548]_ ,
    \new_[21549]_ , \new_[21550]_ , \new_[21551]_ , \new_[21552]_ ,
    \new_[21553]_ , \new_[21554]_ , \new_[21555]_ , \new_[21556]_ ,
    \new_[21557]_ , \new_[21558]_ , \new_[21559]_ , \new_[21560]_ ,
    \new_[21561]_ , \new_[21562]_ , \new_[21563]_ , \new_[21564]_ ,
    \new_[21565]_ , \new_[21566]_ , \new_[21567]_ , \new_[21568]_ ,
    \new_[21569]_ , \new_[21570]_ , \new_[21571]_ , \new_[21572]_ ,
    \new_[21573]_ , \new_[21574]_ , \new_[21575]_ , \new_[21576]_ ,
    \new_[21577]_ , \new_[21578]_ , \new_[21579]_ , \new_[21580]_ ,
    \new_[21581]_ , \new_[21582]_ , \new_[21583]_ , \new_[21584]_ ,
    \new_[21585]_ , \new_[21586]_ , \new_[21587]_ , \new_[21588]_ ,
    \new_[21589]_ , \new_[21590]_ , \new_[21591]_ , \new_[21592]_ ,
    \new_[21593]_ , \new_[21594]_ , \new_[21595]_ , \new_[21596]_ ,
    \new_[21597]_ , \new_[21598]_ , \new_[21599]_ , \new_[21600]_ ,
    \new_[21601]_ , \new_[21602]_ , \new_[21603]_ , \new_[21604]_ ,
    \new_[21605]_ , \new_[21606]_ , \new_[21607]_ , \new_[21608]_ ,
    \new_[21609]_ , \new_[21610]_ , \new_[21611]_ , \new_[21612]_ ,
    \new_[21613]_ , \new_[21614]_ , \new_[21615]_ , \new_[21616]_ ,
    \new_[21617]_ , \new_[21618]_ , \new_[21619]_ , \new_[21620]_ ,
    \new_[21621]_ , \new_[21622]_ , \new_[21623]_ , \new_[21624]_ ,
    \new_[21625]_ , \new_[21626]_ , \new_[21627]_ , \new_[21628]_ ,
    \new_[21629]_ , \new_[21630]_ , \new_[21631]_ , \new_[21632]_ ,
    \new_[21633]_ , \new_[21634]_ , \new_[21635]_ , \new_[21636]_ ,
    \new_[21637]_ , \new_[21638]_ , \new_[21639]_ , \new_[21640]_ ,
    \new_[21641]_ , \new_[21642]_ , \new_[21643]_ , \new_[21644]_ ,
    \new_[21645]_ , \new_[21646]_ , \new_[21647]_ , \new_[21648]_ ,
    \new_[21649]_ , \new_[21650]_ , \new_[21651]_ , \new_[21652]_ ,
    \new_[21653]_ , \new_[21654]_ , \new_[21655]_ , \new_[21656]_ ,
    \new_[21657]_ , \new_[21658]_ , \new_[21659]_ , \new_[21660]_ ,
    \new_[21661]_ , \new_[21662]_ , \new_[21663]_ , \new_[21664]_ ,
    \new_[21665]_ , \new_[21666]_ , \new_[21667]_ , \new_[21668]_ ,
    \new_[21669]_ , \new_[21670]_ , \new_[21671]_ , \new_[21672]_ ,
    \new_[21673]_ , \new_[21674]_ , \new_[21675]_ , \new_[21676]_ ,
    \new_[21677]_ , \new_[21678]_ , \new_[21679]_ , \new_[21680]_ ,
    \new_[21681]_ , \new_[21682]_ , \new_[21683]_ , \new_[21684]_ ,
    \new_[21685]_ , \new_[21686]_ , \new_[21687]_ , \new_[21688]_ ,
    \new_[21689]_ , \new_[21690]_ , \new_[21691]_ , \new_[21692]_ ,
    \new_[21693]_ , \new_[21694]_ , \new_[21695]_ , \new_[21696]_ ,
    \new_[21697]_ , \new_[21698]_ , \new_[21699]_ , \new_[21700]_ ,
    \new_[21701]_ , \new_[21702]_ , \new_[21703]_ , \new_[21704]_ ,
    \new_[21705]_ , \new_[21706]_ , \new_[21707]_ , \new_[21708]_ ,
    \new_[21709]_ , \new_[21710]_ , \new_[21711]_ , \new_[21712]_ ,
    \new_[21713]_ , \new_[21714]_ , n778, n783, n788, n793, n798, n803,
    n808, n813, n818, n823, n828, n833, n838, n843, n848, n853, n858, n863,
    n868, n873, n878, n883, n888, n893, n898, n903, n908, n913, n918, n923,
    n928, n933, n938, n943, n948, n953, n958, n963, n968, n973, n978, n983,
    n988, n993, n998, n1003, n1008, n1013, n1018, n1023, n1028, n1033,
    n1038, n1043, n1048, n1053, n1058, n1063, n1068, n1073, n1078, n1083,
    n1088, n1093, n1098, n1103, n1108, n1113, n1118, n1123, n1128, n1133,
    n1138, n1143, n1148, n1153, n1158, n1163, n1168, n1173, n1178, n1183,
    n1188, n1193, n1198, n1203, n1208, n1213, n1218, n1223, n1228, n1233,
    n1238, n1243, n1248, n1253, n1258, n1263, n1268, n1273, n1278, n1283,
    n1288, n1293, n1298, n1303, n1308, n1313, n1318, n1323, n1328, n1333,
    n1338, n1343, n1348, n1353, n1358, n1363, n1368, n1373, n1378, n1383,
    n1388, n1393, n1398, n1403, n1408, n1413, n1418, n1423, n1428, n1433,
    n1438, n1443, n1448, n1453, n1458, n1463, n1468, n1473, n1478, n1483,
    n1488, n1493, n1498, n1503, n1508, n1513, n1518, n1523, n1528, n1533,
    n1538, n1543, n1548, n1553, n1558, n1563, n1568, n1573, n1578, n1583,
    n1588, n1593, n1598, n1603, n1608, n1613, n1618, n1623, n1628, n1633,
    n1638, n1643, n1648, n1653, n1658, n1663, n1668, n1673, n1678, n1683,
    n1688, n1693, n1698, n1703, n1708, n1713, n1718, n1723, n1728, n1733,
    n1738, n1743, n1748, n1753, n1758, n1763, n1768, n1773, n1778, n1783,
    n1788, n1793, n1798, n1803, n1808, n1813, n1818, n1823, n1828, n1833,
    n1838, n1843, n1848, n1853, n1858, n1863, n1868, n1873, n1878, n1883,
    n1888, n1893, n1898, n1903, n1908, n1913, n1918, n1923, n1928, n1933,
    n1938, n1943, n1948, n1953, n1958, n1963, n1968, n1973, n1978, n1983,
    n1988, n1993, n1998, n2003, n2008, n2013, n2018, n2023, n2028, n2033,
    n2038, n2043, n2048, n2053, n2058, n2063, n2068, n2073, n2078, n2083,
    n2088, n2093, n2098, n2103, n2108, n2113, n2118, n2123, n2128, n2133,
    n2138, n2143, n2148, n2153, n2158, n2163, n2168, n2173, n2178, n2183,
    n2188, n2193, n2198, n2203, n2208, n2213, n2218, n2223, n2228, n2233,
    n2238, n2243, n2248, n2253, n2258, n2263, n2268, n2273, n2278, n2283,
    n2288, n2293, n2298, n2303, n2308, n2313, n2318, n2323, n2328, n2333,
    n2338, n2343, n2348, n2353, n2358, n2363, n2368, n2373, n2378, n2383,
    n2388, n2393, n2398, n2403, n2408, n2413, n2418, n2423, n2428, n2433,
    n2438, n2443, n2448, n2453, n2458, n2463, n2468, n2473, n2478, n2483,
    n2488, n2493, n2498, n2503, n2508, n2513, n2518, n2523, n2528, n2533,
    n2538, n2543, n2548, n2553, n2558, n2563, n2568, n2573, n2578, n2583,
    n2588, n2593, n2598, n2603, n2608, n2613, n2618, n2623, n2628, n2633,
    n2638, n2643, n2648, n2653, n2658, n2663, n2668, n2673, n2678, n2683,
    n2688, n2693, n2698, n2703, n2708, n2713, n2718, n2723, n2728, n2733,
    n2738, n2743, n2748, n2753, n2758, n2763, n2768, n2773, n2778, n2783,
    n2788, n2793, n2798, n2803, n2808, n2813, n2818, n2823, n2828, n2833,
    n2838, n2843, n2848, n2853, n2858, n2863, n2868, n2873, n2878, n2883,
    n2888, n2893, n2898, n2903, n2908, n2913, n2918, n2923, n2928, n2933,
    n2938, n2943, n2948, n2953, n2958, n2963, n2968, n2973, n2978, n2983,
    n2988, n2993, n2998, n3003, n3008, n3013, n3018, n3023, n3028, n3033,
    n3038, n3043, n3048, n3053, n3058, n3063, n3068, n3073, n3078, n3083,
    n3088, n3093, n3098, n3103, n3108, n3113, n3118, n3123, n3128, n3133,
    n3138, n3143, n3148, n3153, n3158, n3163, n3168, n3173, n3178, n3183,
    n3188, n3193, n3198, n3203, n3208, n3213, n3218, n3223, n3228, n3233,
    n3238, n3243, n3248, n3253, n3258, n3263, n3268, n3273, n3278, n3283,
    n3288, n3293, n3298, n3303, n3308, n3313, n3318, n3323, n3328, n3333,
    n3338, n3343, n3348, n3353, n3358, n3363, n3368, n3373, n3378, n3383,
    n3388, n3393, n3398, n3403, n3408, n3413, n3418, n3423;
  assign \new_[920]_  = \\sa22_reg[4] ;
  assign \new_[921]_  = \\sa02_reg[1] ;
  assign \new_[922]_  = \\sa01_reg[1] ;
  assign \new_[923]_  = \\sa00_reg[1] ;
  assign \new_[924]_  = \\sa03_reg[4] ;
  assign \new_[925]_  = \\sa03_reg[3] ;
  assign \new_[926]_  = \\sa33_reg[0] ;
  assign \new_[927]_  = \\sa02_reg[4] ;
  assign \new_[928]_  = \\sa12_reg[3] ;
  assign \new_[929]_  = \\sa32_reg[3] ;
  assign \new_[930]_  = ~\\sa32_reg[0] ;
  assign \new_[931]_  = \\sa22_reg[3] ;
  assign \new_[932]_  = \\sa31_reg[0] ;
  assign \new_[933]_  = \\sa02_reg[3] ;
  assign \new_[934]_  = \\sa20_reg[3] ;
  assign \new_[935]_  = \\sa30_reg[0] ;
  assign \new_[936]_  = \\sa00_reg[4] ;
  assign \new_[937]_  = \\sa10_reg[0] ;
  assign \new_[938]_  = \\sa03_reg[0] ;
  assign \new_[939]_  = \\sa33_reg[3] ;
  assign \new_[940]_  = \\sa13_reg[0] ;
  assign \new_[941]_  = \\sa02_reg[6] ;
  assign \new_[942]_  = \\sa22_reg[5] ;
  assign \new_[943]_  = \\sa13_reg[4] ;
  assign \new_[944]_  = \\sa03_reg[1] ;
  assign \new_[945]_  = \\sa32_reg[5] ;
  assign \new_[946]_  = \\sa12_reg[1] ;
  assign \new_[947]_  = \\sa13_reg[3] ;
  assign \new_[948]_  = \\sa23_reg[3] ;
  assign \new_[949]_  = \\sa02_reg[0] ;
  assign \new_[950]_  = \\sa12_reg[0] ;
  assign \new_[951]_  = \\sa21_reg[4] ;
  assign \new_[952]_  = \\sa01_reg[4] ;
  assign \new_[953]_  = \\sa31_reg[5] ;
  assign \new_[954]_  = \\sa11_reg[1] ;
  assign \new_[955]_  = \\sa21_reg[3] ;
  assign \new_[956]_  = \\sa01_reg[0] ;
  assign \new_[957]_  = \\sa21_reg[5] ;
  assign \new_[958]_  = \\sa11_reg[0] ;
  assign \new_[959]_  = \\sa10_reg[1] ;
  assign \new_[960]_  = \\sa20_reg[1] ;
  assign \new_[961]_  = \\sa00_reg[5] ;
  assign \new_[962]_  = \\sa30_reg[6] ;
  assign \new_[963]_  = \\sa10_reg[3] ;
  assign \new_[964]_  = \\sa00_reg[0] ;
  assign \new_[965]_  = \\sa00_reg[7] ;
  assign n778 = ~\new_[13101]_  | (~\new_[1113]_  & ~\new_[15808]_ );
  assign n788 = ~\new_[12999]_  | (~\new_[1110]_  & ~\new_[14659]_ );
  assign n783 = ~\new_[12909]_  | (~\new_[1114]_  & ~\new_[13673]_ );
  assign n793 = ~\new_[12964]_  | (~\new_[1091]_  & ~\new_[15780]_ );
  assign \new_[970]_  = \\sa23_reg[6] ;
  assign n798 = ~\new_[8053]_  | (~\new_[1166]_  & ~\new_[14998]_ );
  assign \new_[972]_  = \\sa13_reg[6] ;
  assign \new_[973]_  = \\sa13_reg[1] ;
  assign \new_[974]_  = \\sa33_reg[4] ;
  assign \new_[975]_  = \\sa23_reg[7] ;
  assign \new_[976]_  = \\sa33_reg[7] ;
  assign \new_[977]_  = \\sa03_reg[6] ;
  assign n808 = ~\new_[12930]_  | (~\new_[1163]_  & ~\new_[17582]_ );
  assign \new_[979]_  = \\sa23_reg[0] ;
  assign \new_[980]_  = \\sa02_reg[5] ;
  assign \new_[981]_  = \\sa32_reg[6] ;
  assign \new_[982]_  = \\sa12_reg[6] ;
  assign \new_[983]_  = \\sa22_reg[6] ;
  assign \new_[984]_  = \\sa22_reg[1] ;
  assign \new_[985]_  = \\sa12_reg[4] ;
  assign \new_[986]_  = \\sa22_reg[0] ;
  assign \new_[987]_  = \\sa01_reg[6] ;
  assign \new_[988]_  = \\sa11_reg[6] ;
  assign \new_[989]_  = \\sa31_reg[6] ;
  assign \new_[990]_  = \\sa01_reg[5] ;
  assign \new_[991]_  = \\sa21_reg[1] ;
  assign \new_[992]_  = \\sa11_reg[3] ;
  assign \new_[993]_  = \\sa01_reg[3] ;
  assign \new_[994]_  = \\sa21_reg[0] ;
  assign \new_[995]_  = \\sa31_reg[3] ;
  assign \new_[996]_  = \\sa10_reg[5] ;
  assign \new_[997]_  = \\sa30_reg[5] ;
  assign \new_[998]_  = \\sa20_reg[5] ;
  assign \new_[999]_  = \\sa30_reg[1] ;
  assign \new_[1000]_  = \\sa00_reg[3] ;
  assign \new_[1001]_  = \\sa30_reg[4] ;
  assign \new_[1002]_  = \\sa10_reg[4] ;
  assign \new_[1003]_  = \\sa10_reg[6] ;
  assign \new_[1004]_  = \\sa20_reg[0] ;
  assign \new_[1005]_  = \\sa30_reg[3] ;
  assign \new_[1006]_  = \\sa30_reg[2] ;
  assign \new_[1007]_  = \\sa00_reg[6] ;
  assign \new_[1008]_  = \\sa20_reg[6] ;
  assign \new_[1009]_  = \\sa20_reg[2] ;
  assign n813 = ~\new_[12873]_  | (~\new_[1170]_  & ~\new_[15808]_ );
  assign n843 = ~\new_[13209]_  | (~\new_[1171]_  & ~\new_[15101]_ );
  assign n833 = ~\new_[12004]_  | (~\new_[1173]_  & ~\new_[14989]_ );
  assign n818 = ~\new_[13206]_  | (~\new_[1172]_  & ~\new_[15101]_ );
  assign n823 = ~\new_[11730]_  | (~\new_[1174]_  & ~\new_[13673]_ );
  assign n848 = ~\new_[12840]_  | (~\new_[1140]_  & ~\new_[15450]_ );
  assign n858 = ~\new_[11844]_  | (~\new_[1141]_  & ~\new_[15234]_ );
  assign n803 = ~\new_[5429]_  | (~\new_[1169]_  & ~\new_[15234]_ );
  assign n863 = ~\new_[13144]_  | (~\new_[1142]_  & ~\new_[15238]_ );
  assign n1003 = ~\new_[1133]_  | ~\new_[12517]_ ;
  assign n918 = ~\new_[6274]_  | (~\new_[1231]_  & ~\new_[15450]_ );
  assign \new_[1021]_  = \\sa03_reg[5] ;
  assign \new_[1022]_  = \\sa23_reg[4] ;
  assign \new_[1023]_  = \\sa33_reg[5] ;
  assign \new_[1024]_  = \\sa23_reg[5] ;
  assign \new_[1025]_  = \\sa33_reg[1] ;
  assign \new_[1026]_  = \\sa23_reg[1] ;
  assign \new_[1027]_  = \\sa33_reg[2] ;
  assign \new_[1028]_  = \\sa03_reg[2] ;
  assign \new_[1029]_  = \\sa23_reg[2] ;
  assign \new_[1030]_  = \\sa13_reg[7] ;
  assign \new_[1031]_  = \\sa03_reg[7] ;
  assign \new_[1032]_  = \\sa12_reg[5] ;
  assign \new_[1033]_  = \\sa32_reg[1] ;
  assign \new_[1034]_  = \\sa22_reg[7] ;
  assign \new_[1035]_  = \\sa02_reg[7] ;
  assign \new_[1036]_  = \\sa12_reg[7] ;
  assign \new_[1037]_  = \\sa21_reg[6] ;
  assign \new_[1038]_  = \\sa11_reg[5] ;
  assign \new_[1039]_  = \\sa31_reg[1] ;
  assign \new_[1040]_  = \\sa11_reg[4] ;
  assign \new_[1041]_  = \\sa31_reg[2] ;
  assign \new_[1042]_  = \\sa01_reg[7] ;
  assign \new_[1043]_  = \\sa21_reg[2] ;
  assign \new_[1044]_  = \\sa20_reg[4] ;
  assign \new_[1045]_  = \\sa20_reg[7] ;
  assign \new_[1046]_  = \\sa10_reg[7] ;
  assign \new_[1047]_  = \\sa30_reg[7] ;
  assign n963 = ~\new_[13288]_  | (~\new_[1208]_  & ~\new_[14998]_ );
  assign n888 = ~\new_[13300]_  | (~\new_[1217]_  & ~\new_[17582]_ );
  assign n893 = ~\new_[8097]_  | (~\new_[1222]_  & ~\new_[15235]_ );
  assign n938 = ~\new_[13262]_  | (~\new_[1215]_  & ~\new_[15779]_ );
  assign n943 = ~\new_[13320]_  | (~\new_[1214]_  & ~\new_[15779]_ );
  assign n933 = ~\new_[13201]_  | (~\new_[1213]_  & ~\new_[14659]_ );
  assign n873 = ~\new_[5409]_  | (~\new_[1199]_  & ~\new_[14924]_ );
  assign n948 = ~\new_[13134]_  | (~\new_[1216]_  & ~\new_[13518]_ );
  assign n868 = ~\new_[13258]_  | (~\new_[1195]_  & ~\new_[14924]_ );
  assign n953 = ~\new_[11753]_  | (~\new_[1218]_  & ~\new_[14924]_ );
  assign n903 = ~\new_[13042]_  | (~\new_[1225]_  & ~\new_[15808]_ );
  assign n878 = ~\new_[13264]_  | (~\new_[1198]_  & ~\new_[14657]_ );
  assign n908 = ~\new_[12456]_  | (~\new_[1226]_  & ~\new_[15101]_ );
  assign n968 = ~\new_[13243]_  | (~\new_[1219]_  & ~\new_[15233]_ );
  assign n958 = ~\new_[13079]_  | (~\new_[1220]_  & ~\new_[15239]_ );
  assign n923 = ~\new_[12902]_  | (~\new_[1230]_  & ~\new_[14989]_ );
  assign n928 = ~\new_[13255]_  | (~\new_[1229]_  & ~\new_[15233]_ );
  assign n983 = ~\new_[13011]_  | (~\new_[1182]_  & ~\new_[15239]_ );
  assign n898 = ~\new_[7042]_  | (~\new_[1227]_  & ~\new_[15234]_ );
  assign n988 = ~\new_[1175]_  | ~\new_[13050]_ ;
  assign n973 = ~\new_[13231]_  | (~\new_[1191]_  & ~\new_[15781]_ );
  assign n978 = ~\new_[13130]_  | (~\new_[1192]_  & ~\new_[15235]_ );
  assign n993 = ~\new_[12931]_  | (~\new_[1194]_  & ~\new_[15450]_ );
  assign n913 = ~\new_[5043]_  | (~\new_[1228]_  & ~\new_[15234]_ );
  assign n998 = ~\new_[13180]_  | (~\new_[1197]_  & ~\new_[15238]_ );
  assign n1183 = ~\new_[12974]_  | ~\new_[1189]_ ;
  assign n1178 = ~\new_[11816]_  | (~\new_[1252]_  & ~\new_[13533]_ );
  assign n1038 = ~\new_[9342]_  | ~\new_[1184]_ ;
  assign n828 = ~\new_[1130]_ ;
  assign n1188 = ~\new_[13481]_  | ~\new_[1190]_ ;
  assign \new_[1078]_  = \\sa13_reg[5] ;
  assign \new_[1079]_  = \\sa33_reg[6] ;
  assign \new_[1080]_  = \\sa32_reg[2] ;
  assign \new_[1081]_  = \\sa02_reg[2] ;
  assign \new_[1082]_  = \\sa12_reg[2] ;
  assign \new_[1083]_  = \\sa22_reg[2] ;
  assign \new_[1084]_  = \\sa01_reg[2] ;
  assign \new_[1085]_  = \\sa11_reg[2] ;
  assign \new_[1086]_  = \\sa11_reg[7] ;
  assign \new_[1087]_  = \\sa00_reg[2] ;
  assign \new_[1088]_  = \\u0_w_reg[2][19] ;
  assign \new_[1089]_  = \\sa10_reg[2] ;
  assign n1193 = ~\new_[13275]_  | (~\new_[1258]_  & ~\new_[13671]_ );
  assign \new_[1091]_  = \new_[1747]_  ? \new_[1263]_  : \new_[1931]_ ;
  assign n853 = ~\new_[1143]_ ;
  assign n1053 = ~\new_[1205]_  | ~\new_[12832]_ ;
  assign n1048 = ~\new_[13023]_  | (~\new_[1270]_  & ~\new_[14658]_ );
  assign n1098 = ~\new_[12149]_  | (~\new_[1265]_  & ~\new_[14658]_ );
  assign n1083 = ~\new_[1202]_  | ~\new_[13110]_ ;
  assign n1088 = ~\new_[1203]_  | ~\new_[13229]_ ;
  assign n1058 = ~\new_[12842]_  | ~\new_[1206]_ ;
  assign n1093 = ~\new_[1204]_  | ~\new_[12884]_ ;
  assign n1013 = ~\new_[1193]_  | ~\new_[9357]_ ;
  assign n1063 = ~\new_[12033]_  | ~\new_[1207]_ ;
  assign n1113 = ~\new_[13067]_  | (~\new_[1269]_  & ~\new_[15780]_ );
  assign n1068 = ~\new_[13295]_  | (~\new_[1275]_  & ~\new_[17582]_ );
  assign n1108 = ~\new_[12487]_  | (~\new_[1271]_  & ~\new_[14924]_ );
  assign n1073 = ~\new_[11247]_  | (~\new_[1278]_  & ~\new_[15808]_ );
  assign n1008 = ~\new_[1196]_  | ~\new_[9331]_ ;
  assign n1118 = ~\new_[11814]_  | (~\new_[1274]_  & ~\new_[15235]_ );
  assign n1123 = ~\new_[11834]_  | (~\new_[1273]_  & ~\new_[15782]_ );
  assign n1043 = ~\new_[12371]_  | (~\new_[1254]_  & ~\new_[13671]_ );
  assign \new_[1110]_  = \new_[1792]_  ? \new_[1262]_  : \new_[1972]_ ;
  assign n1078 = ~\new_[13109]_  | (~\new_[1283]_  & ~\new_[15233]_ );
  assign n838 = ~\new_[1168]_ ;
  assign \new_[1113]_  = \new_[1306]_  ? \new_[1823]_  : \new_[1259]_ ;
  assign \new_[1114]_  = \new_[1838]_  ? \new_[1261]_  : \new_[2038]_ ;
  assign n1033 = ~\new_[1181]_  | ~\new_[9297]_ ;
  assign n1028 = ~\new_[1201]_  | ~\new_[10636]_ ;
  assign n1023 = ~\new_[8103]_  | (~\new_[1281]_  & ~\new_[15238]_ );
  assign n1128 = ~\new_[12944]_  | (~\new_[1234]_  & ~\new_[15239]_ );
  assign n1138 = ~\new_[13010]_  | (~\new_[1235]_  & ~\new_[14998]_ );
  assign n1133 = ~\new_[12855]_  | (~\new_[1233]_  & ~\new_[15781]_ );
  assign n1143 = ~\new_[12998]_  | (~\new_[1246]_  & ~\new_[15781]_ );
  assign n1148 = ~\new_[12864]_  | (~\new_[1247]_  & ~\new_[15458]_ );
  assign n1153 = ~\new_[11962]_  | (~\new_[1248]_  & ~\new_[15780]_ );
  assign n1158 = ~\new_[13111]_  | (~\new_[1249]_  & ~\new_[15238]_ );
  assign n1018 = ~\new_[10687]_  | (~\new_[1282]_  & ~\new_[13533]_ );
  assign n1163 = ~\new_[1178]_  | ~\new_[12934]_ ;
  assign n1168 = ~\new_[11859]_  | (~\new_[1251]_  & ~\new_[14657]_ );
  assign n1173 = ~\new_[13305]_  | (~\new_[1250]_  & ~\new_[14657]_ );
  assign n1323 = ~\new_[1244]_  | ~\new_[13119]_ ;
  assign \new_[1130]_  = \new_[2844]_  ^ \new_[1313]_ ;
  assign n1318 = ~\new_[1245]_  | ~\new_[12965]_ ;
  assign n1328 = ~\new_[12147]_  | (~\new_[1301]_  & ~\new_[15450]_ );
  assign \new_[1133]_  = ~\new_[1253]_  | ~\new_[16131]_ ;
  assign \new_[1134]_  = \\sa13_reg[2] ;
  assign \new_[1135]_  = \\sa32_reg[7] ;
  assign \new_[1136]_  = \\sa32_reg[4] ;
  assign \new_[1137]_  = \\sa31_reg[7] ;
  assign \new_[1138]_  = \\sa31_reg[4] ;
  assign \new_[1139]_  = \\sa21_reg[7] ;
  assign \new_[1140]_  = \new_[1775]_  ? \new_[1315]_  : \new_[1947]_ ;
  assign \new_[1141]_  = \new_[21366]_  ? \new_[1746]_  : \new_[1309]_ ;
  assign \new_[1142]_  = \new_[2319]_  ? \new_[1311]_  : \new_[2571]_ ;
  assign \new_[1143]_  = \new_[2864]_  ^ \new_[1317]_ ;
  assign n1223 = ~\new_[10630]_  | (~\new_[1322]_  & ~\new_[15782]_ );
  assign n1208 = ~\new_[9313]_  | (~\new_[1333]_  & ~\new_[15782]_ );
  assign n1283 = ~\new_[13249]_  | (~\new_[1312]_  & ~\new_[15779]_ );
  assign n1278 = ~\new_[1257]_  | ~\new_[13290]_ ;
  assign n1253 = ~\new_[13191]_  | (~\new_[1326]_  & ~\new_[14658]_ );
  assign n1213 = ~\new_[9295]_  | (~\new_[1292]_  & ~\new_[14659]_ );
  assign n1233 = ~\new_[6319]_  | (~\new_[1286]_  & ~\new_[13671]_ );
  assign n1288 = ~\new_[13316]_  | (~\new_[1321]_  & ~\new_[17582]_ );
  assign n1293 = ~\new_[12793]_  | (~\new_[1323]_  & ~\new_[14998]_ );
  assign n1218 = ~\new_[11737]_  | (~\new_[1329]_  & ~\new_[15781]_ );
  assign n1298 = ~\new_[13043]_  | (~\new_[1325]_  & ~\new_[14659]_ );
  assign n1258 = ~\new_[12821]_  | (~\new_[1334]_  & ~\new_[13673]_ );
  assign n1248 = ~\new_[1277]_  | ~\new_[12034]_ ;
  assign n1203 = ~\new_[6392]_  | (~\new_[1332]_  & ~\new_[15458]_ );
  assign n1243 = ~\new_[1276]_  | ~\new_[9290]_ ;
  assign n1303 = ~\new_[1268]_  | ~\new_[13127]_ ;
  assign n1308 = ~\new_[13022]_  | (~\new_[1331]_  & ~\new_[15235]_ );
  assign n1263 = ~\new_[13301]_  | ~\new_[1272]_ ;
  assign n1238 = ~\new_[5382]_  | (~\new_[1293]_  & ~\new_[13671]_ );
  assign \new_[1163]_  = \new_[2556]_  ? \new_[1307]_  : \new_[2781]_ ;
  assign n1268 = ~\new_[13135]_  | ~\new_[1279]_ ;
  assign n1228 = ~\new_[6254]_  | (~\new_[1335]_  & ~\new_[15458]_ );
  assign \new_[1166]_  = \new_[1390]_  ? \new_[1536]_  : \new_[1310]_ ;
  assign n1273 = ~\new_[1280]_  | ~\new_[13001]_ ;
  assign \new_[1168]_  = \new_[2945]_  ^ \new_[1320]_ ;
  assign \new_[1169]_  = \new_[1610]_  ? \new_[1305]_  : \new_[1487]_ ;
  assign \new_[1170]_  = \new_[1387]_  ? \new_[2015]_  : \new_[1308]_ ;
  assign \new_[1171]_  = \new_[1780]_  ? \new_[1336]_  : \new_[1608]_ ;
  assign \new_[1172]_  = \new_[1738]_  ? \new_[1337]_  : \new_[1574]_ ;
  assign \new_[1173]_  = \new_[1316]_  ^ \new_[1836]_ ;
  assign \new_[1174]_  = \new_[1339]_  ? \new_[1463]_  : \new_[1284]_ ;
  assign \new_[1175]_  = ~\new_[1236]_  | ~\new_[16130]_ ;
  assign n1198 = ~\new_[10716]_  | (~\new_[1287]_  & ~\new_[15779]_ );
  assign n1313 = ~\new_[12024]_  | (~\new_[1294]_  & ~\new_[15458]_ );
  assign \new_[1178]_  = ~\new_[16130]_  | ~\new_[1296]_ ;
  assign n1378 = ~\new_[13013]_  | (~\new_[1365]_  & ~\new_[13533]_ );
  assign n1388 = ~\new_[12954]_  | (~\new_[1373]_  & ~\new_[13533]_ );
  assign \new_[1181]_  = ~\new_[1295]_  | ~\new_[19872]_ ;
  assign \new_[1182]_  = \new_[2627]_  ? \new_[1374]_  : \new_[2890]_ ;
  assign n1383 = \new_[1375]_  ? \new_[19371]_  : \key[51] ;
  assign \new_[1184]_  = ~\new_[1302]_  | ~\new_[16130]_ ;
  assign \new_[1185]_  = \\u0_w_reg[3][29] ;
  assign \new_[1186]_  = \\u0_w_reg[0][19] ;
  assign \new_[1187]_  = ~\\u0_w_reg[1][19] ;
  assign \new_[1188]_  = \\u0_w_reg[3][19] ;
  assign \new_[1189]_  = ~\new_[1304]_  | ~\new_[16131]_ ;
  assign \new_[1190]_  = ~\new_[1303]_  | ~\new_[15011]_ ;
  assign \new_[1191]_  = \new_[1448]_  ? \new_[1583]_  : \new_[1378]_ ;
  assign \new_[1192]_  = \new_[1976]_  ? \new_[1381]_  : \new_[2178]_ ;
  assign \new_[1193]_  = ~\new_[20592]_  | ~\new_[15011]_ ;
  assign \new_[1194]_  = \new_[1735]_  ^ \new_[1382]_ ;
  assign \new_[1195]_  = \new_[1800]_  ? \new_[1385]_  : \new_[1985]_ ;
  assign \new_[1196]_  = ~\new_[1299]_  | ~\new_[16131]_ ;
  assign \new_[1197]_  = \new_[2316]_  ? \new_[1391]_  : \new_[2567]_ ;
  assign \new_[1198]_  = \new_[1804]_  ? \new_[1386]_  : \new_[1986]_ ;
  assign \new_[1199]_  = \new_[1974]_  ? \new_[1398]_  : \new_[1794]_ ;
  assign n1333 = ~\new_[9301]_  | (~\new_[1361]_  & ~\new_[17582]_ );
  assign \new_[1201]_  = ~\new_[1338]_  | ~\new_[19872]_ ;
  assign \new_[1202]_  = ~\new_[1318]_  | ~\new_[16130]_ ;
  assign \new_[1203]_  = ~\new_[1319]_  | ~\new_[15011]_ ;
  assign \new_[1204]_  = ~\new_[1314]_  | ~\new_[16131]_ ;
  assign \new_[1205]_  = ~\new_[1327]_  | ~\new_[19872]_ ;
  assign \new_[1206]_  = ~\new_[1330]_  | ~\new_[15011]_ ;
  assign \new_[1207]_  = ~\new_[1328]_  | ~\new_[16130]_ ;
  assign \new_[1208]_  = \new_[1777]_  ? \new_[1371]_  : \new_[1949]_ ;
  assign n1363 = ~\new_[13063]_  | (~\new_[1403]_  & ~\new_[15239]_ );
  assign n1343 = ~\new_[13008]_  | (~\new_[1405]_  & ~\new_[15101]_ );
  assign n1368 = ~\new_[12844]_  | (~\new_[1404]_  & ~\new_[15233]_ );
  assign n1373 = ~\new_[1324]_  | ~\new_[10858]_ ;
  assign \new_[1213]_  = \new_[1457]_  ? \new_[1779]_  : \new_[1384]_ ;
  assign \new_[1214]_  = \new_[1783]_  ? \new_[1369]_  : \new_[1612]_ ;
  assign \new_[1215]_  = \new_[1459]_  ? \new_[1954]_  : \new_[1389]_ ;
  assign \new_[1216]_  = \new_[1379]_  ? \new_[1615]_  : \new_[1449]_ ;
  assign \new_[1217]_  = \new_[1814]_  ? \new_[1372]_  : \new_[1999]_ ;
  assign \new_[1218]_  = \new_[1399]_  ^ \new_[1791]_ ;
  assign \new_[1219]_  = \new_[1808]_  ? \new_[1392]_  : \new_[1991]_ ;
  assign \new_[1220]_  = \new_[1807]_  ? \new_[1395]_  : \new_[1988]_ ;
  assign n1348 = ~\new_[12896]_  | (~\new_[1407]_  & ~\new_[14989]_ );
  assign \new_[1222]_  = \new_[1456]_  ? \new_[1364]_  : \new_[1576]_ ;
  assign n1353 = ~\new_[12921]_  | (~\new_[1410]_  & ~\new_[14989]_ );
  assign n1358 = ~\new_[13095]_  | (~\new_[1408]_  & ~\new_[14658]_ );
  assign \new_[1225]_  = \new_[1825]_  ? \new_[1367]_  : \new_[1635]_ ;
  assign \new_[1226]_  = \new_[1380]_  ? \new_[1641]_  : \new_[1450]_ ;
  assign \new_[1227]_  = \new_[1914]_  ? \new_[1388]_  : \new_[2119]_ ;
  assign \new_[1228]_  = \new_[1383]_  ? \new_[1729]_  : \new_[1455]_ ;
  assign \new_[1229]_  = \new_[1647]_  ? \new_[1393]_  : \new_[1849]_ ;
  assign \new_[1230]_  = \new_[1651]_  ? \new_[1394]_  : \new_[1852]_ ;
  assign \new_[1231]_  = \new_[1919]_  ^ \new_[1396]_ ;
  assign n1338 = ~\new_[10701]_  | (~\new_[1362]_  & ~\new_[15782]_ );
  assign \new_[1233]_  = \new_[1932]_  ? \new_[1440]_  : \new_[1748]_ ;
  assign \new_[1234]_  = \new_[1543]_  ? \new_[1551]_  : \new_[1441]_ ;
  assign \new_[1235]_  = \new_[1716]_  ? \new_[1442]_  : \new_[1908]_ ;
  assign \new_[1236]_  = \new_[1623]_  ? \new_[1909]_  : \new_[1494]_ ;
  assign \new_[1237]_  = \\u0_w_reg[2][21] ;
  assign \new_[1238]_  = \\u0_w_reg[0][27] ;
  assign \new_[1239]_  = ~\\u0_w_reg[1][27] ;
  assign \new_[1240]_  = \\u0_w_reg[2][27] ;
  assign \new_[1241]_  = \\u0_w_reg[2][11] ;
  assign \new_[1242]_  = \\u0_w_reg[3][27] ;
  assign \new_[1243]_  = \\u0_w_reg[3][24] ;
  assign \new_[1244]_  = ~\new_[1376]_  | ~\new_[15011]_ ;
  assign \new_[1245]_  = ~\new_[1370]_  | ~\new_[16130]_ ;
  assign \new_[1246]_  = \new_[1582]_  ? \new_[1451]_  : \new_[1751]_ ;
  assign \new_[1247]_  = \new_[1569]_  ^ \new_[1485]_ ;
  assign \new_[1248]_  = \new_[2125]_  ? \new_[1458]_  : \new_[1920]_ ;
  assign \new_[1249]_  = \new_[1453]_  ? \new_[1462]_  : \new_[1571]_ ;
  assign \new_[1250]_  = \new_[1579]_  ? \new_[1465]_  : \new_[1460]_ ;
  assign \new_[1251]_  = \new_[2320]_  ? \new_[1464]_  : \new_[2573]_ ;
  assign \new_[1252]_  = \new_[1498]_  ? \new_[1796]_  : \new_[1628]_ ;
  assign \new_[1253]_  = ~\new_[1377]_  | (~\new_[1613]_  & ~\new_[21482]_ );
  assign \new_[1254]_  = \new_[1806]_  ? \new_[1493]_  : \new_[1990]_ ;
  assign n1398 = ~\new_[13153]_  | (~\new_[1482]_  & ~\new_[17582]_ );
  assign n1408 = ~\new_[11838]_  | (~\new_[1461]_  & ~\new_[17582]_ );
  assign \new_[1257]_  = ~\new_[1397]_  | ~\new_[16131]_ ;
  assign \new_[1258]_  = \new_[2241]_  ? \new_[1499]_  : \new_[2471]_ ;
  assign \new_[1259]_  = ~\new_[1306]_ ;
  assign n1418 = ~\new_[13112]_  | (~\new_[1483]_  & ~\new_[15780]_ );
  assign \new_[1261]_  = ~\new_[1400]_  | ~\new_[1471]_ ;
  assign \new_[1262]_  = ~\new_[1401]_  | ~\new_[1472]_ ;
  assign \new_[1263]_  = ~\new_[1402]_  | ~\new_[1473]_ ;
  assign n1413 = ~\new_[12914]_  | (~\new_[1481]_  & ~\new_[14659]_ );
  assign \new_[1265]_  = \new_[3120]_  ? \new_[1484]_  : \new_[2891]_ ;
  assign n1393 = ~\new_[5902]_  | (~\new_[1423]_  & ~\new_[14657]_ );
  assign n1403 = ~\new_[12827]_  | (~\new_[1497]_  & ~\new_[13673]_ );
  assign \new_[1268]_  = ~\new_[21238]_  | ~\new_[16130]_ ;
  assign \new_[1269]_  = \new_[1609]_  ? \new_[1491]_  : \new_[1486]_ ;
  assign \new_[1270]_  = \new_[2889]_  ? \new_[1500]_  : \new_[3119]_ ;
  assign \new_[1271]_  = \new_[1736]_  ? \new_[1492]_  : \new_[1572]_ ;
  assign \new_[1272]_  = ~\new_[1406]_  | ~\new_[16131]_ ;
  assign \new_[1273]_  = \new_[1626]_  ? \new_[1580]_  : \new_[1495]_ ;
  assign \new_[1274]_  = \new_[1809]_  ? \new_[1496]_  : \new_[1993]_ ;
  assign \new_[1275]_  = \new_[1638]_  ? \new_[1566]_  : \new_[1501]_ ;
  assign \new_[1276]_  = ~\new_[1368]_  | ~\new_[16130]_ ;
  assign \new_[1277]_  = ~\new_[1366]_  | ~\new_[16131]_ ;
  assign \new_[1278]_  = \new_[1454]_  ? \new_[1636]_  : \new_[1575]_ ;
  assign \new_[1279]_  = ~\new_[1409]_  | ~\new_[16131]_ ;
  assign \new_[1280]_  = ~\new_[1411]_  | ~\new_[15011]_ ;
  assign \new_[1281]_  = \new_[1923]_  ^ \new_[1446]_ ;
  assign \new_[1282]_  = \new_[1568]_  ? \new_[1915]_  : \new_[1452]_ ;
  assign \new_[1283]_  = \new_[1649]_  ? \new_[1414]_  : \new_[1850]_ ;
  assign \new_[1284]_  = ~\new_[1339]_ ;
  assign n1423 = ~\new_[18907]_  | ~\new_[1437]_ ;
  assign \new_[1286]_  = \new_[2754]_  ? \new_[1606]_  : \new_[2990]_ ;
  assign \new_[1287]_  = \new_[3122]_  ? \new_[1642]_  : \new_[21370]_ ;
  assign \new_[1288]_  = ~\\u0_w_reg[2][29] ;
  assign \new_[1289]_  = \\u0_w_reg[0][29] ;
  assign \new_[1290]_  = \\u0_w_reg[2][5] ;
  assign \new_[1291]_  = \\u0_w_reg[2][3] ;
  assign \new_[1292]_  = \new_[1829]_  ? \new_[1552]_  : \new_[2025]_ ;
  assign \new_[1293]_  = \new_[1977]_  ? \new_[1630]_  : \new_[2179]_ ;
  assign \new_[1294]_  = \new_[1776]_  ? \new_[1577]_  : \new_[1605]_ ;
  assign \new_[1295]_  = ~\new_[1447]_  | (~\new_[1782]_  & ~\new_[1834]_ );
  assign \new_[1296]_  = ~\new_[1439]_  | (~\new_[1981]_  & ~\new_[1752]_ );
  assign n1428 = \key[115]  ? \new_[19614]_  : \new_[1616]_ ;
  assign n1433 = \key[83]  ? \new_[19614]_  : \new_[1617]_ ;
  assign \new_[1299]_  = ~\new_[1444]_  | (~\new_[2035]_  & ~\new_[1842]_ );
  assign n1438 = \key[19]  ? \new_[19649]_  : \new_[1618]_ ;
  assign \new_[1301]_  = \new_[1785]_  ? \new_[1624]_  : \new_[1614]_ ;
  assign \new_[1302]_  = ~\new_[1443]_  | (~\new_[1844]_  & ~\new_[2190]_ );
  assign \new_[1303]_  = ~\new_[1445]_  | (~\new_[1973]_  & ~\new_[1835]_ );
  assign \new_[1304]_  = \new_[2193]_  ? \new_[1622]_  : \new_[2191]_ ;
  assign \new_[1305]_  = \new_[1634]_  ? \new_[2712]_  : \new_[1821]_ ;
  assign \new_[1306]_  = ~\new_[1602]_  | ~\new_[1480]_ ;
  assign \new_[1307]_  = ~\new_[1479]_  | ~\new_[1599]_ ;
  assign \new_[1308]_  = ~\new_[1387]_ ;
  assign \new_[1309]_  = ~\new_[21366]_ ;
  assign \new_[1310]_  = ~\new_[1390]_ ;
  assign \new_[1311]_  = ~\new_[1475]_  | ~\new_[1592]_ ;
  assign \new_[1312]_  = \new_[1711]_  ? \new_[1778]_  : \new_[1544]_ ;
  assign \new_[1313]_  = ~\new_[1470]_  | ~\new_[1587]_ ;
  assign \new_[1314]_  = \new_[1801]_  ? \new_[1950]_  : \new_[1625]_ ;
  assign \new_[1315]_  = ~\new_[1468]_  | ~\new_[1584]_ ;
  assign \new_[1316]_  = ~\new_[1469]_  | ~\new_[1586]_ ;
  assign \new_[1317]_  = ~\new_[1476]_  | ~\new_[1597]_ ;
  assign \new_[1318]_  = ~\new_[1466]_  | (~\new_[1952]_  & ~\new_[21479]_ );
  assign \new_[1319]_  = ~\new_[1467]_  | (~\new_[2149]_  & ~\new_[1753]_ );
  assign \new_[1320]_  = ~\new_[1478]_  | ~\new_[1598]_ ;
  assign \new_[1321]_  = \new_[1788]_  ? \new_[1567]_  : \new_[1964]_ ;
  assign \new_[1322]_  = \new_[1730]_  ? \new_[1549]_  : \new_[1918]_ ;
  assign \new_[1323]_  = \new_[1573]_  ? \new_[1611]_  : \new_[1737]_ ;
  assign \new_[1324]_  = ~\new_[1490]_  | ~\new_[15011]_ ;
  assign \new_[1325]_  = \new_[1629]_  ? \new_[1793]_  : \new_[1813]_ ;
  assign \new_[1326]_  = \new_[1712]_  ? \new_[1819]_  : \new_[1545]_ ;
  assign \new_[1327]_  = \new_[1797]_  ? \new_[1817]_  : \new_[1621]_ ;
  assign \new_[1328]_  = ~\new_[1489]_  | (~\new_[1837]_  & ~\new_[2219]_ );
  assign \new_[1329]_  = \new_[1650]_  ? \new_[1565]_  : \new_[1854]_ ;
  assign \new_[1330]_  = ~\new_[1488]_  | (~\new_[2221]_  & ~\new_[1754]_ );
  assign \new_[1331]_  = \new_[1987]_  ? \new_[1631]_  : \new_[1803]_ ;
  assign \new_[1332]_  = \new_[1578]_  ? \new_[1696]_  : \new_[1740]_ ;
  assign \new_[1333]_  = \new_[1699]_  ? \new_[1542]_  : \new_[1533]_ ;
  assign \new_[1334]_  = \new_[1830]_  ? \new_[1564]_  : \new_[2027]_ ;
  assign \new_[1335]_  = \new_[1627]_  ? \new_[1570]_  : \new_[1812]_ ;
  assign \new_[1336]_  = \new_[1632]_  ? \new_[2095]_  : \new_[1820]_ ;
  assign \new_[1337]_  = \new_[2011]_  ? \new_[2317]_  : \new_[1822]_ ;
  assign \new_[1338]_  = ~\new_[1412]_  | (~\new_[1784]_  & ~\new_[2134]_ );
  assign \new_[1339]_  = \new_[3063]_  ? \new_[1705]_  : \new_[2849]_ ;
  assign n1443 = \new_[1707]_  ? \new_[19371]_  : \key[53] ;
  assign \new_[1341]_  = \\u0_w_reg[1][29] ;
  assign \new_[1342]_  = \\u0_w_reg[0][30] ;
  assign \new_[1343]_  = ~\\u0_w_reg[1][30] ;
  assign \new_[1344]_  = \\u0_w_reg[3][30] ;
  assign \new_[1345]_  = \\u0_w_reg[0][21] ;
  assign \new_[1346]_  = ~\\u0_w_reg[1][21] ;
  assign \new_[1347]_  = \\u0_w_reg[2][0] ;
  assign \new_[1348]_  = \\u0_w_reg[2][10] ;
  assign \new_[1349]_  = \\u0_w_reg[2][14] ;
  assign \new_[1350]_  = \\u0_w_reg[2][30] ;
  assign \new_[1351]_  = \\u0_w_reg[2][16] ;
  assign \new_[1352]_  = \\u0_w_reg[2][8] ;
  assign \new_[1353]_  = \\u0_w_reg[2][15] ;
  assign \new_[1354]_  = \\u0_w_reg[3][21] ;
  assign \text_out[12]  = \\text_out_reg[12] ;
  assign n1448 = \new_[1731]_  ? \new_[19372]_  : \key[123] ;
  assign n1453 = \new_[1732]_  ? \new_[19372]_  : \key[91] ;
  assign n1458 = \new_[1733]_  ? \new_[19372]_  : \key[59] ;
  assign n1468 = \new_[1734]_  ? \new_[19415]_  : \key[27] ;
  assign n1463 = \new_[1745]_  ? \new_[19496]_  : \key[43] ;
  assign \new_[1361]_  = \new_[1907]_  ? \new_[2044]_  : \new_[1715]_ ;
  assign \new_[1362]_  = \new_[1798]_  ? \new_[2040]_  : \new_[1980]_ ;
  assign n1473 = ~\new_[18748]_  | ~\new_[1563]_ ;
  assign \new_[1364]_  = ~\new_[1556]_  | ~\new_[1718]_ ;
  assign \new_[1365]_  = \new_[2524]_  ? \new_[1781]_  : \new_[2523]_ ;
  assign \new_[1366]_  = \new_[2869]_  ? \new_[1790]_  : \new_[2868]_ ;
  assign \new_[1367]_  = ~\new_[1561]_  | ~\new_[1725]_ ;
  assign \new_[1368]_  = ~\new_[1553]_  | (~\new_[2164]_  & ~\new_[1992]_ );
  assign \new_[1369]_  = ~\new_[1562]_  | ~\new_[1728]_ ;
  assign \new_[1370]_  = ~\new_[1560]_  | (~\new_[1955]_  & ~\new_[2469]_ );
  assign \new_[1371]_  = ~\new_[1723]_  | ~\new_[1558]_ ;
  assign \new_[1372]_  = ~\new_[1724]_  | ~\new_[1559]_ ;
  assign \new_[1373]_  = \new_[1786]_  ? \new_[2043]_  : \new_[1958]_ ;
  assign \new_[1374]_  = \new_[2041]_  ? \new_[2166]_  : \new_[1840]_ ;
  assign \new_[1375]_  = \new_[18296]_  ^ \new_[1795]_ ;
  assign \new_[1376]_  = ~\new_[1557]_  | (~\new_[2031]_  & ~\new_[2194]_ );
  assign \new_[1377]_  = ~\new_[1613]_  | ~\new_[21482]_ ;
  assign \new_[1378]_  = ~\new_[1448]_ ;
  assign \new_[1379]_  = ~\new_[1449]_ ;
  assign \new_[1380]_  = ~\new_[1450]_ ;
  assign \new_[1381]_  = ~\new_[1771]_  | ~\new_[1604]_ ;
  assign \new_[1382]_  = ~\new_[1770]_  | ~\new_[1603]_ ;
  assign \new_[1383]_  = ~\new_[1455]_ ;
  assign \new_[1384]_  = ~\new_[1457]_ ;
  assign \new_[1385]_  = ~\new_[1600]_  | ~\new_[1766]_ ;
  assign \new_[1386]_  = ~\new_[1767]_  | ~\new_[1601]_ ;
  assign \new_[1387]_  = ~\new_[1588]_  | ~\new_[1759]_ ;
  assign \new_[1388]_  = ~\new_[1589]_  | ~\new_[1760]_ ;
  assign \new_[1389]_  = ~\new_[1459]_ ;
  assign \new_[1390]_  = ~\new_[1590]_  | ~\new_[1762]_ ;
  assign \new_[1391]_  = ~\new_[1591]_  | ~\new_[1757]_ ;
  assign \new_[1392]_  = ~\new_[1593]_  | ~\new_[1763]_ ;
  assign \new_[1393]_  = ~\new_[1594]_  | ~\new_[1764]_ ;
  assign \new_[1394]_  = ~\new_[1595]_  | ~\new_[1765]_ ;
  assign \new_[1395]_  = ~\new_[1596]_  | ~\new_[1758]_ ;
  assign \new_[1396]_  = \new_[2112]_  ? \new_[1833]_  : \new_[2341]_ ;
  assign \new_[1397]_  = ~\new_[1581]_  | (~\new_[2034]_  & ~\new_[2146]_ );
  assign \new_[1398]_  = \new_[2285]_  ? \new_[1833]_  : \new_[2533]_ ;
  assign \new_[1399]_  = ~\new_[1585]_  | ~\new_[1755]_ ;
  assign \new_[1400]_  = ~\new_[2449]_  | ~\new_[1502]_ ;
  assign \new_[1401]_  = ~\new_[2455]_  | ~\new_[1503]_ ;
  assign \new_[1402]_  = ~\new_[2230]_  | ~\new_[1504]_ ;
  assign \new_[1403]_  = \new_[2989]_  ? \new_[1799]_  : \new_[2988]_ ;
  assign \new_[1404]_  = \new_[1787]_  ? \new_[1805]_  : \new_[1959]_ ;
  assign \new_[1405]_  = \new_[1811]_  ? \new_[1839]_  : \new_[1998]_ ;
  assign \new_[1406]_  = ~\new_[1633]_  | (~\new_[1957]_  & ~\new_[2255]_ );
  assign \new_[1407]_  = \new_[2987]_  ? \new_[1845]_  : \new_[2986]_ ;
  assign \new_[1408]_  = \new_[1848]_  ? \new_[1815]_  : \new_[1643]_ ;
  assign \new_[1409]_  = ~\new_[1640]_  | (~\new_[1847]_  & ~\new_[21576]_ );
  assign \new_[1410]_  = \new_[1960]_  ? \new_[1644]_  : \new_[2156]_ ;
  assign \new_[1411]_  = ~\new_[1639]_  | (~\new_[2058]_  & ~\new_[1989]_ );
  assign \new_[1412]_  = ~\new_[1784]_  | ~\new_[2134]_ ;
  assign n1483 = \new_[1903]_  ? \new_[19372]_  : \key[125] ;
  assign \new_[1414]_  = \new_[2330]_  ? \new_[2024]_  : \new_[2599]_ ;
  assign n1478 = \new_[1905]_  ? \new_[19414]_  : \key[61] ;
  assign n1488 = \new_[1912]_  ? ld : \key[37] ;
  assign \new_[1417]_  = \\u0_w_reg[2][12] ;
  assign \new_[1418]_  = \\u0_w_reg[0][24] ;
  assign \new_[1419]_  = \\u0_w_reg[0][31] ;
  assign \new_[1420]_  = \\u0_w_reg[1][24] ;
  assign \new_[1421]_  = ~\\u0_w_reg[1][31] ;
  assign \new_[1422]_  = \\u0_w_reg[2][24] ;
  assign \new_[1423]_  = \new_[2142]_  ? \new_[1979]_  : \new_[1948]_ ;
  assign \new_[1424]_  = \\u0_w_reg[2][31] ;
  assign \new_[1425]_  = \\u0_w_reg[3][31] ;
  assign \new_[1426]_  = \\u0_w_reg[0][5] ;
  assign \new_[1427]_  = \\u0_w_reg[2][22] ;
  assign \new_[1428]_  = \\u0_w_reg[2][6] ;
  assign \new_[1429]_  = \\u0_w_reg[3][5] ;
  assign \new_[1430]_  = \\u0_w_reg[0][11] ;
  assign \new_[1431]_  = \\u0_w_reg[1][11] ;
  assign \new_[1432]_  = \\u0_w_reg[2][17] ;
  assign \new_[1433]_  = \\u0_w_reg[2][9] ;
  assign \new_[1434]_  = \\u0_w_reg[3][11] ;
  assign \text_out[125]  = \\text_out_reg[125] ;
  assign \text_out[44]  = \\text_out_reg[44] ;
  assign \new_[1437]_  = ~\new_[1706]_  | ~\new_[19649]_ ;
  assign n1493 = \new_[1930]_  ? \new_[19415]_  : \key[35] ;
  assign \new_[1439]_  = ~\new_[1981]_  | ~\new_[1752]_ ;
  assign \new_[1440]_  = ~\new_[1726]_  | ~\new_[1727]_ ;
  assign \new_[1441]_  = ~\new_[1543]_ ;
  assign \new_[1442]_  = ~\new_[1722]_  | ~\new_[1721]_ ;
  assign \new_[1443]_  = ~\new_[1844]_  | ~\new_[2661]_ ;
  assign \new_[1444]_  = ~\new_[2035]_  | ~\new_[1842]_ ;
  assign \new_[1445]_  = ~\new_[1973]_  | ~\new_[1835]_ ;
  assign \new_[1446]_  = \new_[2562]_  ? \new_[2014]_  : \new_[2792]_ ;
  assign \new_[1447]_  = ~\new_[1782]_  | ~\new_[1834]_ ;
  assign \new_[1448]_  = \new_[2266]_  ? \new_[20046]_  : \new_[2050]_ ;
  assign \new_[1449]_  = \new_[2267]_  ? \new_[2429]_  : \new_[2051]_ ;
  assign \new_[1450]_  = \new_[2268]_  ? \new_[2430]_  : \new_[2052]_ ;
  assign \new_[1451]_  = ~\new_[1774]_  | ~\new_[1773]_ ;
  assign \new_[1452]_  = ~\new_[1568]_ ;
  assign \new_[1453]_  = ~\new_[1571]_ ;
  assign \new_[1454]_  = ~\new_[1575]_ ;
  assign \new_[1455]_  = ~\new_[1936]_  | ~\new_[1768]_ ;
  assign \new_[1456]_  = ~\new_[1576]_ ;
  assign \new_[1457]_  = ~\new_[1937]_  | ~\new_[1769]_ ;
  assign \new_[1458]_  = \new_[2627]_  ? \new_[2016]_  : \new_[2890]_ ;
  assign \new_[1459]_  = ~\new_[1761]_  | ~\new_[1935]_ ;
  assign \new_[1460]_  = ~\new_[1579]_ ;
  assign \new_[1461]_  = \new_[2155]_  ^ \new_[1953]_ ;
  assign \new_[1462]_  = ~\new_[1756]_  | ~\new_[1934]_ ;
  assign \new_[1463]_  = \new_[2553]_  ? \new_[2026]_  : \new_[2780]_ ;
  assign \new_[1464]_  = \new_[1855]_  ? \new_[2020]_  : \new_[2072]_ ;
  assign \new_[1465]_  = \new_[2060]_  ? \new_[2021]_  : \new_[2279]_ ;
  assign \new_[1466]_  = ~\new_[21479]_  | ~\new_[1952]_ ;
  assign \new_[1467]_  = ~\new_[2149]_  | ~\new_[1753]_ ;
  assign \new_[1468]_  = ~\new_[2101]_  | ~\new_[1828]_ ;
  assign \new_[1469]_  = ~\new_[2325]_  | ~\new_[1831]_ ;
  assign \new_[1470]_  = ~\new_[2449]_  | ~\new_[1827]_ ;
  assign \new_[1471]_  = ~\new_[2448]_  | ~\new_[1645]_ ;
  assign \new_[1472]_  = ~\new_[2454]_  | ~\new_[1646]_ ;
  assign \new_[1473]_  = ~\new_[2229]_  | ~\new_[1648]_ ;
  assign \new_[1474]_  = ~\\u0_w_reg[1][5] ;
  assign \new_[1475]_  = ~\new_[2231]_  | ~\new_[1818]_ ;
  assign \new_[1476]_  = ~\new_[2230]_  | ~\new_[1826]_ ;
  assign \new_[1477]_  = \\u0_w_reg[2][13] ;
  assign \new_[1478]_  = ~\new_[2455]_  | ~\new_[1832]_ ;
  assign \new_[1479]_  = ~\new_[2458]_  | ~\new_[1816]_ ;
  assign \new_[1480]_  = ~\new_[1822]_  | ~\new_[3119]_ ;
  assign \new_[1481]_  = \new_[1927]_  ^ \new_[1971]_ ;
  assign \new_[1482]_  = \new_[2153]_  ^ \new_[2006]_ ;
  assign \new_[1483]_  = \new_[2176]_  ? \new_[1956]_  : \new_[1975]_ ;
  assign \new_[1484]_  = \new_[2249]_  ? \new_[2385]_  : \new_[2042]_ ;
  assign \new_[1485]_  = ~\new_[1810]_  | ~\new_[1995]_ ;
  assign \new_[1486]_  = ~\new_[1609]_ ;
  assign \new_[1487]_  = ~\new_[1610]_ ;
  assign \new_[1488]_  = ~\new_[2221]_  | ~\new_[1754]_ ;
  assign \new_[1489]_  = ~\new_[1837]_  | ~\new_[2219]_ ;
  assign \new_[1490]_  = ~\new_[1789]_  | (~\new_[2198]_  & ~\new_[2195]_ );
  assign \new_[1491]_  = \new_[2008]_  ? \new_[2208]_  : \new_[2223]_ ;
  assign \new_[1492]_  = \new_[2010]_  ? \new_[2422]_  : \new_[2225]_ ;
  assign \new_[1493]_  = \new_[2532]_  ? \new_[2029]_  : \new_[21538]_ ;
  assign \new_[1494]_  = ~\new_[1623]_ ;
  assign \new_[1495]_  = ~\new_[1626]_ ;
  assign \new_[1496]_  = \new_[2440]_  ? \new_[2022]_  : \new_[2701]_ ;
  assign \new_[1497]_  = \new_[1922]_  ^ \new_[2033]_ ;
  assign \new_[1498]_  = ~\new_[1628]_ ;
  assign \new_[1499]_  = ~\new_[1843]_  | ~\new_[2045]_ ;
  assign \new_[1500]_  = \new_[2248]_  ? \new_[2486]_  : \new_[2039]_ ;
  assign \new_[1501]_  = ~\new_[1638]_ ;
  assign \new_[1502]_  = ~\new_[1645]_ ;
  assign \new_[1503]_  = ~\new_[1646]_ ;
  assign \new_[1504]_  = ~\new_[1648]_ ;
  assign n1568 = \new_[19419]_  ^ \new_[2622]_ ;
  assign \new_[1506]_  = \\u0_w_reg[1][3] ;
  assign \new_[1507]_  = \\u0_w_reg[0][3] ;
  assign \new_[1508]_  = \\u0_w_reg[3][3] ;
  assign \new_[1509]_  = \\u0_w_reg[2][4] ;
  assign \new_[1510]_  = ~\\u0_w_reg[1][28] ;
  assign \new_[1511]_  = \\u0_w_reg[3][28] ;
  assign \text_out[93]  = \\text_out_reg[93] ;
  assign \new_[1513]_  = \\u0_w_reg[0][0] ;
  assign \text_out[61]  = \\text_out_reg[61] ;
  assign \new_[1515]_  = \\u0_w_reg[0][16] ;
  assign \new_[1516]_  = ~\\u0_w_reg[1][0] ;
  assign \new_[1517]_  = \\u0_w_reg[3][0] ;
  assign \new_[1518]_  = ~\\u0_w_reg[1][16] ;
  assign \new_[1519]_  = \\u0_w_reg[3][16] ;
  assign \text_out[101]  = \\text_out_reg[101] ;
  assign \text_out[108]  = \\text_out_reg[108] ;
  assign \text_out[43]  = \\text_out_reg[43] ;
  assign \text_out[109]  = \\text_out_reg[109] ;
  assign \text_out[117]  = \\text_out_reg[117] ;
  assign \text_out[76]  = \\text_out_reg[76] ;
  assign \text_out[111]  = \\text_out_reg[111] ;
  assign \text_out[48]  = \\text_out_reg[48] ;
  assign \text_out[80]  = \\text_out_reg[80] ;
  assign \text_out[112]  = \\text_out_reg[112] ;
  assign \text_out[46]  = \\text_out_reg[46] ;
  assign \text_out[126]  = \\text_out_reg[126] ;
  assign \text_out[10]  = \\text_out_reg[10] ;
  assign \new_[1533]_  = ~\new_[1699]_ ;
  assign n1503 = \new_[2143]_  ? \new_[19472]_  : \key[126] ;
  assign n1508 = \new_[2145]_  ? \new_[19496]_  : \key[94] ;
  assign \new_[1536]_  = \new_[2375]_  ^ \new_[2061]_ ;
  assign n1543 = \new_[2147]_  ? \new_[19451]_  : \key[62] ;
  assign n1513 = \new_[2148]_  ? \new_[19496]_  : \key[30] ;
  assign n1518 = \new_[2150]_  ? \new_[19496]_  : \key[117] ;
  assign n1523 = \new_[2151]_  ? \new_[19496]_  : \key[85] ;
  assign n1563 = \new_[2152]_  ? \new_[19338]_  : \key[21] ;
  assign \new_[1542]_  = ~\new_[1917]_  | ~\new_[2122]_ ;
  assign \new_[1543]_  = \new_[3241]_  ? \new_[2185]_  : \new_[21332]_ ;
  assign \new_[1544]_  = ~\new_[1711]_ ;
  assign \new_[1545]_  = ~\new_[1712]_ ;
  assign n1528 = \new_[2181]_  ? \new_[19414]_  : \key[32] ;
  assign n1533 = \new_[2180]_  ? \new_[19414]_  : \key[42] ;
  assign n1548 = \new_[2182]_  ? \new_[19414]_  : \key[48] ;
  assign \new_[1549]_  = ~\new_[1906]_  | ~\new_[2111]_ ;
  assign n1538 = \new_[2184]_  ? n3423 : \key[46] ;
  assign \new_[1551]_  = \new_[3277]_  ? \new_[2167]_  : \new_[3074]_ ;
  assign \new_[1552]_  = ~\new_[1916]_  | ~\new_[2121]_ ;
  assign \new_[1553]_  = ~\new_[2164]_  | ~\new_[1992]_ ;
  assign n1558 = \new_[2188]_  ? \new_[19414]_  : \key[47] ;
  assign n1553 = \new_[2189]_  ? \new_[19338]_  : \key[40] ;
  assign \new_[1556]_  = ~\new_[1853]_  | ~\new_[2376]_ ;
  assign \new_[1557]_  = ~\new_[2031]_  | ~\new_[2194]_ ;
  assign \new_[1558]_  = ~\new_[3242]_  | ~\new_[2399]_ ;
  assign \new_[1559]_  = ~\new_[3051]_  | ~\new_[1984]_ ;
  assign \new_[1560]_  = ~\new_[1955]_  | ~\new_[2469]_ ;
  assign \new_[1561]_  = ~\new_[20973]_  | ~\new_[3642]_ ;
  assign \new_[1562]_  = ~\new_[2399]_  | ~\new_[3687]_ ;
  assign \new_[1563]_  = ~\new_[1951]_  | ~\new_[19077]_ ;
  assign \new_[1564]_  = ~\new_[1938]_  | ~\new_[1939]_ ;
  assign \new_[1565]_  = ~\new_[1940]_  | ~\new_[1941]_ ;
  assign \new_[1566]_  = \new_[2987]_  ? \new_[2233]_  : \new_[2986]_ ;
  assign \new_[1567]_  = ~\new_[1942]_  | ~\new_[1943]_ ;
  assign \new_[1568]_  = \new_[2521]_  ? \new_[2685]_  : \new_[2269]_ ;
  assign \new_[1569]_  = \new_[2222]_  ^ \new_[2759]_ ;
  assign \new_[1570]_  = \new_[17475]_  ? \new_[2234]_  : \new_[18194]_ ;
  assign \new_[1571]_  = \new_[2687]_  ? \new_[2209]_  : \new_[2937]_ ;
  assign \new_[1572]_  = ~\new_[1736]_ ;
  assign \new_[1573]_  = ~\new_[1737]_ ;
  assign \new_[1574]_  = ~\new_[1738]_ ;
  assign \new_[1575]_  = \new_[2217]_  ? \new_[2211]_  : \new_[2431]_ ;
  assign \new_[1576]_  = \new_[2432]_  ? \new_[2212]_  : \new_[2690]_ ;
  assign \new_[1577]_  = \new_[2627]_  ? \new_[2224]_  : \new_[2890]_ ;
  assign \new_[1578]_  = ~\new_[1740]_ ;
  assign \new_[1579]_  = ~\new_[1933]_  | ~\new_[2133]_ ;
  assign \new_[1580]_  = \new_[2283]_  ? \new_[2235]_  : \new_[2555]_ ;
  assign \new_[1581]_  = ~\new_[2034]_  | ~\new_[2146]_ ;
  assign \new_[1582]_  = ~\new_[1751]_ ;
  assign \new_[1583]_  = \new_[3019]_  ? \new_[2243]_  : \new_[3227]_ ;
  assign \new_[1584]_  = ~\new_[2323]_  | ~\new_[2021]_ ;
  assign \new_[1585]_  = ~\new_[2324]_  | ~\new_[2023]_ ;
  assign \new_[1586]_  = ~\new_[2581]_  | ~\new_[2026]_ ;
  assign \new_[1587]_  = ~\new_[2448]_  | ~\new_[2019]_ ;
  assign \new_[1588]_  = ~\new_[2000]_  | ~\new_[2456]_ ;
  assign \new_[1589]_  = ~\new_[2458]_  | ~\new_[1851]_ ;
  assign \new_[1590]_  = ~\new_[2001]_  | ~\new_[2460]_ ;
  assign \new_[1591]_  = ~\new_[2017]_  | ~\new_[2772]_ ;
  assign \new_[1592]_  = ~\new_[2018]_  | ~\new_[2002]_ ;
  assign \new_[1593]_  = ~\new_[2003]_  | ~\new_[2232]_ ;
  assign \new_[1594]_  = ~\new_[2233]_  | ~\new_[2004]_ ;
  assign \new_[1595]_  = ~\new_[2019]_  | ~\new_[3007]_ ;
  assign \new_[1596]_  = ~\new_[2770]_  | ~\new_[2028]_ ;
  assign \new_[1597]_  = ~\new_[2229]_  | ~\new_[2017]_ ;
  assign \new_[1598]_  = ~\new_[2454]_  | ~\new_[2028]_ ;
  assign \new_[1599]_  = ~\new_[2457]_  | ~\new_[20411]_ ;
  assign \new_[1600]_  = ~\new_[20411]_  | ~\new_[2542]_ ;
  assign \new_[1601]_  = ~\new_[2005]_  | ~\new_[3163]_ ;
  assign \new_[1602]_  = ~\new_[2011]_  | ~\new_[2889]_ ;
  assign \new_[1603]_  = ~\new_[2009]_  | ~\new_[2992]_ ;
  assign \new_[1604]_  = ~\new_[2018]_  | ~\new_[2523]_ ;
  assign \new_[1605]_  = ~\new_[1776]_ ;
  assign \new_[1606]_  = \new_[2106]_  ? \new_[2540]_  : \new_[2334]_ ;
  assign \new_[1607]_  = \\u0_w_reg[3][26] ;
  assign \new_[1608]_  = ~\new_[1780]_ ;
  assign \new_[1609]_  = ~\new_[1996]_  | ~\new_[2206]_ ;
  assign \new_[1610]_  = ~\new_[1997]_  | ~\new_[2207]_ ;
  assign \new_[1611]_  = ~\new_[1969]_  | ~\new_[2161]_ ;
  assign \new_[1612]_  = ~\new_[1783]_ ;
  assign \new_[1613]_  = \new_[2056]_  ^ \new_[3080]_ ;
  assign \new_[1614]_  = ~\new_[1785]_ ;
  assign \new_[1615]_  = ~\new_[1978]_  | ~\new_[2183]_ ;
  assign \new_[1616]_  = \new_[1186]_  ^ \new_[2264]_ ;
  assign \new_[1617]_  = \new_[18334]_  ^ \new_[2264]_ ;
  assign \new_[1618]_  = \new_[5687]_  ^ \new_[2264]_ ;
  assign \new_[1619]_  = ~\\u0_w_reg[1][26] ;
  assign \new_[1620]_  = \\u0_w_reg[2][26] ;
  assign \new_[1621]_  = ~\new_[1797]_ ;
  assign \new_[1622]_  = \new_[2345]_  ? \new_[2570]_  : \new_[2120]_ ;
  assign \new_[1623]_  = ~\new_[2197]_  | ~\new_[1994]_ ;
  assign \new_[1624]_  = \new_[19560]_  ? \new_[2096]_  : \new_[2344]_ ;
  assign \new_[1625]_  = ~\new_[1801]_ ;
  assign \new_[1626]_  = \new_[3171]_  ? \new_[2220]_  : \new_[2947]_ ;
  assign \new_[1627]_  = ~\new_[1812]_ ;
  assign \new_[1628]_  = ~\new_[2049]_  | ~\new_[2262]_ ;
  assign \new_[1629]_  = ~\new_[1813]_ ;
  assign \new_[1630]_  = ~\new_[2048]_  | ~\new_[2261]_ ;
  assign \new_[1631]_  = ~\new_[2046]_  | ~\new_[2257]_ ;
  assign \new_[1632]_  = ~\new_[1820]_ ;
  assign \new_[1633]_  = ~\new_[1957]_  | ~\new_[2255]_ ;
  assign \new_[1634]_  = ~\new_[1821]_ ;
  assign \new_[1635]_  = ~\new_[1825]_ ;
  assign \new_[1636]_  = ~\new_[2032]_  | ~\new_[2239]_ ;
  assign \new_[1637]_  = \\u0_w_reg[0][26] ;
  assign \new_[1638]_  = ~\new_[2030]_  | ~\new_[2236]_ ;
  assign \new_[1639]_  = ~\new_[2058]_  | ~\new_[1989]_ ;
  assign \new_[1640]_  = ~\new_[1847]_  | ~\new_[21576]_ ;
  assign \new_[1641]_  = ~\new_[2047]_  | ~\new_[2260]_ ;
  assign \new_[1642]_  = \new_[2250]_  ^ \new_[2630]_ ;
  assign \new_[1643]_  = ~\new_[1848]_ ;
  assign \new_[1644]_  = \new_[21596]_  ? \new_[2327]_  : \new_[21597]_ ;
  assign \new_[1645]_  = ~\new_[2102]_  | (~\new_[2625]_  & ~\new_[3521]_ );
  assign \new_[1646]_  = ~\new_[2103]_  | (~\new_[2626]_  & ~\new_[20323]_ );
  assign \new_[1647]_  = ~\new_[1849]_ ;
  assign \new_[1648]_  = ~\new_[2104]_  | (~\new_[2624]_  & ~\new_[3519]_ );
  assign \new_[1649]_  = ~\new_[1850]_ ;
  assign \new_[1650]_  = ~\new_[1854]_ ;
  assign \new_[1651]_  = ~\new_[1852]_ ;
  assign \text_out[0]  = \\text_out_reg[0] ;
  assign \text_out[4]  = \\text_out_reg[4] ;
  assign \text_out[6]  = \\text_out_reg[6] ;
  assign \text_out[32]  = \\text_out_reg[32] ;
  assign \new_[1656]_  = \\u0_w_reg[3][14] ;
  assign \text_out[64]  = \\text_out_reg[64] ;
  assign \new_[1658]_  = \\u0_w_reg[2][18] ;
  assign \new_[1659]_  = \\u0_w_reg[2][2] ;
  assign \new_[1660]_  = \\u0_w_reg[2][23] ;
  assign \new_[1661]_  = \\u0_w_reg[2][20] ;
  assign \new_[1662]_  = \\u0_w_reg[2][28] ;
  assign \new_[1663]_  = \\u0_w_reg[0][10] ;
  assign \new_[1664]_  = \\u0_w_reg[0][13] ;
  assign \new_[1665]_  = \\u0_w_reg[0][15] ;
  assign \new_[1666]_  = \\u0_w_reg[0][8] ;
  assign \new_[1667]_  = ~\\u0_w_reg[1][13] ;
  assign \new_[1668]_  = \\u0_w_reg[1][14] ;
  assign \new_[1669]_  = \\u0_w_reg[1][15] ;
  assign \new_[1670]_  = \\u0_w_reg[1][10] ;
  assign \new_[1671]_  = \\u0_w_reg[1][8] ;
  assign \new_[1672]_  = \\u0_w_reg[3][10] ;
  assign \new_[1673]_  = \\u0_w_reg[3][13] ;
  assign \new_[1674]_  = \\u0_w_reg[3][15] ;
  assign \new_[1675]_  = \\u0_w_reg[3][8] ;
  assign \text_out[29]  = \\text_out_reg[29] ;
  assign \text_out[51]  = \\text_out_reg[51] ;
  assign \text_out[45]  = \\text_out_reg[45] ;
  assign \text_out[105]  = \\text_out_reg[105] ;
  assign \text_out[104]  = \\text_out_reg[104] ;
  assign \text_out[77]  = \\text_out_reg[77] ;
  assign \text_out[13]  = \\text_out_reg[13] ;
  assign \text_out[115]  = \\text_out_reg[115] ;
  assign \text_out[19]  = \\text_out_reg[19] ;
  assign \text_out[47]  = \\text_out_reg[47] ;
  assign \text_out[42]  = \\text_out_reg[42] ;
  assign \text_out[79]  = \\text_out_reg[79] ;
  assign \text_out[74]  = \\text_out_reg[74] ;
  assign \text_out[100]  = \\text_out_reg[100] ;
  assign \text_out[62]  = \\text_out_reg[62] ;
  assign \text_out[94]  = \\text_out_reg[94] ;
  assign \text_out[110]  = \\text_out_reg[110] ;
  assign \text_out[78]  = \\text_out_reg[78] ;
  assign \text_out[121]  = \\text_out_reg[121] ;
  assign \text_out[124]  = \\text_out_reg[124] ;
  assign \new_[1696]_  = \new_[2377]_  ^ \new_[2720]_ ;
  assign n1573 = \new_[2366]_  ? \new_[19496]_  : \key[44] ;
  assign n1578 = \new_[2367]_  ? \new_[19472]_  : \key[120] ;
  assign \new_[1699]_  = \new_[16682]_  ? \new_[2374]_  : \new_[19526]_ ;
  assign n1583 = \new_[2368]_  ? \new_[19383]_  : \key[127] ;
  assign n1593 = \new_[2369]_  ? \new_[19496]_  : \key[95] ;
  assign n1598 = \new_[2370]_  ? \new_[19451]_  : \key[56] ;
  assign n1603 = \new_[2371]_  ? \new_[19451]_  : \key[63] ;
  assign n1608 = \new_[2372]_  ? \new_[19496]_  : \key[31] ;
  assign \new_[1705]_  = ~\new_[2115]_  | ~\new_[2343]_ ;
  assign \new_[1706]_  = ~\new_[2123]_  | ~\new_[2124]_ ;
  assign \new_[1707]_  = \new_[18504]_  ^ \new_[2373]_ ;
  assign n1613 = \new_[2387]_  ? ld : \key[101] ;
  assign n1668 = \new_[2388]_  ? ld : \key[69] ;
  assign n1628 = \new_[2389]_  ? \new_[19371]_  : \key[5] ;
  assign \new_[1711]_  = \new_[3242]_  ? \new_[2393]_  : \new_[21618]_ ;
  assign \new_[1712]_  = \new_[3051]_  ? \new_[2395]_  : \new_[20655]_ ;
  assign n1618 = \new_[2391]_  ? \new_[19479]_  : \key[54] ;
  assign n1623 = \new_[2392]_  ? \new_[19479]_  : \key[38] ;
  assign \new_[1715]_  = ~\new_[1907]_ ;
  assign \new_[1716]_  = ~\new_[1908]_ ;
  assign n1673 = \new_[2397]_  ? \new_[19414]_  : \key[45] ;
  assign \new_[1718]_  = ~\new_[2057]_  | ~\new_[2645]_ ;
  assign \new_[1719]_  = \\u0_w_reg[0][28] ;
  assign \new_[1720]_  = \\u0_w_reg[0][14] ;
  assign \new_[1721]_  = ~\new_[3241]_  | ~\new_[2193]_ ;
  assign \new_[1722]_  = ~\new_[3052]_  | ~\new_[2191]_ ;
  assign \new_[1723]_  = ~\new_[3053]_  | ~\new_[21480]_ ;
  assign \new_[1724]_  = ~\new_[2837]_  | ~\new_[20974]_ ;
  assign \new_[1725]_  = ~\new_[20974]_  | ~\new_[3539]_ ;
  assign \new_[1726]_  = ~\new_[2193]_  | ~\new_[3541]_ ;
  assign \new_[1727]_  = ~\new_[2191]_  | ~\new_[3336]_ ;
  assign \new_[1728]_  = ~\new_[21480]_  | ~\new_[3645]_ ;
  assign \new_[1729]_  = \new_[2941]_  ? \new_[2716]_  : \new_[2689]_ ;
  assign \new_[1730]_  = ~\new_[1918]_ ;
  assign \new_[1731]_  = \new_[6250]_  ^ \new_[2433]_ ;
  assign \new_[1732]_  = \new_[18505]_  ^ \new_[2421]_ ;
  assign \new_[1733]_  = \new_[4985]_  ^ \new_[2436]_ ;
  assign \new_[1734]_  = \new_[6172]_  ^ \new_[2421]_ ;
  assign \new_[1735]_  = \new_[2424]_  ? \new_[2277]_  : \new_[2680]_ ;
  assign \new_[1736]_  = ~\new_[2135]_  | ~\new_[2359]_ ;
  assign \new_[1737]_  = \new_[2688]_  ? \new_[2425]_  : \new_[2939]_ ;
  assign \new_[1738]_  = ~\new_[2136]_  | ~\new_[2360]_ ;
  assign \new_[1739]_  = \\u0_w_reg[2][1] ;
  assign \new_[1740]_  = ~\new_[2361]_  | ~\new_[2137]_ ;
  assign n1633 = \key[107]  ? \new_[19649]_  : \new_[2439]_ ;
  assign n1638 = \key[75]  ? \new_[19614]_  : \new_[2441]_ ;
  assign n1653 = \key[11]  ? \new_[19649]_  : \new_[2443]_ ;
  assign \new_[1744]_  = \\u0_w_reg[2][7] ;
  assign \new_[1745]_  = \new_[18507]_  ^ \new_[2442]_ ;
  assign \new_[1746]_  = \new_[2281]_  ^ \new_[2705]_ ;
  assign \new_[1747]_  = ~\new_[1931]_ ;
  assign \new_[1748]_  = ~\new_[1932]_ ;
  assign n1643 = \new_[2481]_  ? \new_[19371]_  : \key[49] ;
  assign n1648 = \new_[2482]_  ? \new_[19414]_  : \key[41] ;
  assign \new_[1751]_  = \new_[3084]_  ? \new_[2478]_  : \new_[2865]_ ;
  assign \new_[1752]_  = \new_[3277]_  ^ \new_[2473]_ ;
  assign \new_[1753]_  = \new_[3075]_  ^ \new_[2475]_ ;
  assign \new_[1754]_  = \new_[3073]_  ^ \new_[2477]_ ;
  assign \new_[1755]_  = ~\new_[2580]_  | ~\new_[2235]_ ;
  assign \new_[1756]_  = ~\new_[2226]_  | ~\new_[2068]_ ;
  assign \new_[1757]_  = ~\new_[2494]_  | ~\new_[2771]_  | ~\new_[2495]_ ;
  assign \new_[1758]_  = ~\new_[2493]_  | ~\new_[3004]_  | ~\new_[2499]_ ;
  assign \new_[1759]_  = ~\new_[2213]_  | ~\new_[2717]_ ;
  assign \new_[1760]_  = ~\new_[2457]_  | ~\new_[2055]_ ;
  assign \new_[1761]_  = ~\new_[2214]_  | ~\new_[2459]_ ;
  assign \new_[1762]_  = ~\new_[2215]_  | ~\new_[20545]_ ;
  assign \new_[1763]_  = ~\new_[2461]_  | ~\new_[20321]_ ;
  assign \new_[1764]_  = ~\new_[2462]_  | ~\new_[2216]_ ;
  assign \new_[1765]_  = ~\new_[2498]_  | ~\new_[2775]_  | ~\new_[2497]_ ;
  assign \new_[1766]_  = ~\new_[20416]_  | ~\new_[2541]_  | ~\new_[20412]_ ;
  assign \new_[1767]_  = ~\new_[2218]_  | ~\new_[2930]_ ;
  assign \new_[1768]_  = ~\new_[2110]_  | ~\new_[2684]_ ;
  assign \new_[1769]_  = ~\new_[2225]_  | ~\new_[3310]_ ;
  assign \new_[1770]_  = ~\new_[2760]_  | ~\new_[2224]_ ;
  assign \new_[1771]_  = ~\new_[2231]_  | ~\new_[2524]_ ;
  assign \text_out[21]  = \\text_out_reg[21] ;
  assign \new_[1773]_  = ~\new_[2229]_  | ~\new_[2523]_ ;
  assign \new_[1774]_  = ~\new_[2230]_  | ~\new_[2524]_ ;
  assign \new_[1775]_  = ~\new_[1947]_ ;
  assign \new_[1776]_  = \new_[2994]_  ? \new_[2292]_  : \new_[2761]_ ;
  assign \new_[1777]_  = ~\new_[1949]_ ;
  assign \new_[1778]_  = \new_[3075]_  ? \new_[2386]_  : \new_[3278]_ ;
  assign \new_[1779]_  = \new_[2660]_  ^ \new_[2423]_ ;
  assign \new_[1780]_  = ~\new_[2205]_  | ~\new_[2415]_ ;
  assign \new_[1781]_  = \new_[3102]_  ? \new_[2275]_  : \new_[2875]_ ;
  assign \new_[1782]_  = ~\new_[2200]_  | ~\new_[2201]_ ;
  assign \new_[1783]_  = \new_[1474]_  ? \new_[2396]_  : \new_[19558]_ ;
  assign \new_[1784]_  = ~\new_[2202]_  | ~\new_[2203]_ ;
  assign \new_[1785]_  = ~\new_[2204]_  | ~\new_[2414]_ ;
  assign \new_[1786]_  = ~\new_[1958]_ ;
  assign \new_[1787]_  = ~\new_[1959]_ ;
  assign \new_[1788]_  = ~\new_[1964]_ ;
  assign \new_[1789]_  = ~\new_[2198]_  | ~\new_[2195]_ ;
  assign \new_[1790]_  = \new_[2339]_  ? \new_[2795]_  : \new_[2611]_ ;
  assign \new_[1791]_  = \new_[2699]_  ? \new_[2679]_  : \new_[2437]_ ;
  assign \new_[1792]_  = ~\new_[1972]_ ;
  assign \new_[1793]_  = \new_[2294]_  ? \new_[2427]_  : \new_[19747]_ ;
  assign \new_[1794]_  = ~\new_[1974]_ ;
  assign \new_[1795]_  = \new_[19124]_  ^ \new_[2518]_ ;
  assign \new_[1796]_  = \new_[2293]_  ? \new_[2314]_  : \new_[19591]_ ;
  assign \new_[1797]_  = ~\new_[2401]_  | ~\new_[2196]_ ;
  assign \new_[1798]_  = ~\new_[1980]_ ;
  assign \new_[1799]_  = \new_[2434]_  ? \new_[2274]_  : \new_[2694]_ ;
  assign \new_[1800]_  = ~\new_[1985]_ ;
  assign \new_[1801]_  = ~\new_[2405]_  | ~\new_[2199]_ ;
  assign n1658 = \new_[1289]_  ^ \new_[2515]_ ;
  assign \new_[1803]_  = ~\new_[1987]_ ;
  assign \new_[1804]_  = ~\new_[1986]_ ;
  assign \new_[1805]_  = \new_[3454]_  ? \new_[2435]_  : \new_[3286]_ ;
  assign \new_[1806]_  = ~\new_[1990]_ ;
  assign \new_[1807]_  = ~\new_[1988]_ ;
  assign \new_[1808]_  = ~\new_[1991]_ ;
  assign \new_[1809]_  = ~\new_[1993]_ ;
  assign \new_[1810]_  = ~\new_[2854]_  | ~\new_[2060]_ ;
  assign \new_[1811]_  = ~\new_[1998]_ ;
  assign \new_[1812]_  = ~\new_[2259]_  | ~\new_[2514]_ ;
  assign \new_[1813]_  = ~\new_[2263]_  | ~\new_[2517]_ ;
  assign \new_[1814]_  = ~\new_[1999]_ ;
  assign \new_[1815]_  = ~\new_[2258]_  | ~\new_[2512]_ ;
  assign \new_[1816]_  = ~\new_[20411]_ ;
  assign \new_[1817]_  = \new_[1428]_  ? \new_[2483]_  : \new_[19662]_ ;
  assign \new_[1818]_  = ~\new_[2002]_ ;
  assign \new_[1819]_  = \new_[3073]_  ? \new_[2489]_  : \new_[3275]_ ;
  assign \new_[1820]_  = ~\new_[2501]_  | ~\new_[2253]_ ;
  assign \new_[1821]_  = ~\new_[2502]_  | ~\new_[2254]_ ;
  assign \new_[1822]_  = ~\new_[2011]_ ;
  assign \new_[1823]_  = \new_[2525]_  ^ \new_[2318]_ ;
  assign n1663 = \new_[1417]_  ^ \new_[2837]_ ;
  assign \new_[1825]_  = \new_[19549]_  ? \new_[2519]_  : \new_[1290]_ ;
  assign \new_[1826]_  = ~\new_[2017]_ ;
  assign \new_[1827]_  = ~\new_[2019]_ ;
  assign \new_[1828]_  = ~\new_[2021]_ ;
  assign \new_[1829]_  = ~\new_[2025]_ ;
  assign \new_[1830]_  = ~\new_[2027]_ ;
  assign \new_[1831]_  = ~\new_[2026]_ ;
  assign \new_[1832]_  = ~\new_[2028]_ ;
  assign \new_[1833]_  = ~\new_[2256]_  | ~\new_[2506]_ ;
  assign \new_[1834]_  = \new_[14690]_  ^ \new_[2351]_ ;
  assign \new_[1835]_  = ~\new_[2251]_  | ~\new_[2487]_ ;
  assign \new_[1836]_  = \new_[2595]_  ? \new_[2569]_  : \new_[2328]_ ;
  assign \new_[1837]_  = ~\new_[2252]_  | ~\new_[2490]_ ;
  assign \new_[1838]_  = ~\new_[2038]_ ;
  assign \new_[1839]_  = \new_[1659]_  ? \new_[2321]_  : \new_[19792]_ ;
  assign \new_[1840]_  = ~\new_[2041]_ ;
  assign \text_out[120]  = \\text_out_reg[120] ;
  assign \new_[1842]_  = \new_[3167]_  ^ \new_[2358]_ ;
  assign \new_[1843]_  = ~\new_[2851]_  | ~\new_[2107]_ ;
  assign \new_[1844]_  = \new_[2356]_  ^ \new_[2618]_ ;
  assign \new_[1845]_  = \new_[2326]_  ? \new_[2273]_  : \new_[2590]_ ;
  assign \text_out[16]  = \\text_out_reg[16] ;
  assign \new_[1847]_  = \new_[3070]_  ^ \new_[2539]_ ;
  assign \new_[1848]_  = \new_[3434]_  ? \new_[2594]_  : \new_[3575]_ ;
  assign \new_[1849]_  = ~\new_[2278]_  | ~\new_[2551]_ ;
  assign \new_[1850]_  = ~\new_[2280]_  | ~\new_[2554]_ ;
  assign \new_[1851]_  = ~\new_[2055]_ ;
  assign \new_[1852]_  = ~\new_[2282]_  | ~\new_[2548]_ ;
  assign \new_[1853]_  = ~\new_[2057]_ ;
  assign \new_[1854]_  = \new_[3012]_  ? \new_[2638]_  : \new_[2785]_ ;
  assign \new_[1855]_  = ~\new_[2072]_ ;
  assign \text_out[5]  = \\text_out_reg[5] ;
  assign \text_out[37]  = \\text_out_reg[37] ;
  assign \text_out[35]  = \\text_out_reg[35] ;
  assign \text_out[69]  = \\text_out_reg[69] ;
  assign \text_out[67]  = \\text_out_reg[67] ;
  assign \new_[1861]_  = \\u0_w_reg[2][25] ;
  assign \new_[1862]_  = ~\\u0_w_reg[1][25] ;
  assign \new_[1863]_  = \\u0_w_reg[0][12] ;
  assign \new_[1864]_  = \\u0_w_reg[3][12] ;
  assign \new_[1865]_  = \\u0_w_reg[0][22] ;
  assign \new_[1866]_  = \\u0_w_reg[0][6] ;
  assign \new_[1867]_  = \\u0_w_reg[1][22] ;
  assign \new_[1868]_  = \\u0_w_reg[1][6] ;
  assign \new_[1869]_  = \\u0_w_reg[3][22] ;
  assign \new_[1870]_  = \\u0_w_reg[3][6] ;
  assign \text_out[56]  = \\text_out_reg[56] ;
  assign \new_[1872]_  = \\u0_w_reg[0][17] ;
  assign \text_out[88]  = \\text_out_reg[88] ;
  assign \new_[1874]_  = \\u0_w_reg[0][9] ;
  assign \new_[1875]_  = \\u0_w_reg[1][17] ;
  assign \text_out[53]  = \\text_out_reg[53] ;
  assign \new_[1877]_  = \\u0_w_reg[1][9] ;
  assign \new_[1878]_  = \\u0_w_reg[3][17] ;
  assign \new_[1879]_  = \\u0_w_reg[3][9] ;
  assign \text_out[85]  = \\text_out_reg[85] ;
  assign \text_out[83]  = \\text_out_reg[83] ;
  assign \text_out[24]  = \\text_out_reg[24] ;
  assign \text_out[75]  = \\text_out_reg[75] ;
  assign \text_out[123]  = \\text_out_reg[123] ;
  assign \text_out[73]  = \\text_out_reg[73] ;
  assign \text_out[106]  = \\text_out_reg[106] ;
  assign n1793 = \new_[1515]_  ^ \new_[2624]_ ;
  assign \text_out[82]  = \\text_out_reg[82] ;
  assign \text_out[30]  = \\text_out_reg[30] ;
  assign \text_out[23]  = \\text_out_reg[23] ;
  assign \text_out[18]  = \\text_out_reg[18] ;
  assign \text_out[114]  = \\text_out_reg[114] ;
  assign \text_out[57]  = \\text_out_reg[57] ;
  assign \text_out[89]  = \\text_out_reg[89] ;
  assign n1783 = \new_[1351]_  ^ \new_[2625]_ ;
  assign \text_out[60]  = \\text_out_reg[60] ;
  assign n1788 = \new_[19708]_  ^ \new_[2626]_ ;
  assign n1778 = \new_[1665]_  ^ \new_[2621]_ ;
  assign n1828 = \new_[2639]_  ? \new_[19472]_  : \key[122] ;
  assign n1818 = \new_[2640]_  ? \new_[19383]_  : \key[90] ;
  assign n1823 = \new_[2643]_  ? \new_[19451]_  : \key[58] ;
  assign n1813 = \new_[2644]_  ? \new_[19383]_  : \key[26] ;
  assign \new_[1903]_  = \new_[6995]_  ? \new_[2653]_  : \new_[6251]_ ;
  assign n1498 = \new_[2642]_  ? \new_[16274]_  : \new_[2641]_ ;
  assign \new_[1905]_  = \new_[5334]_  ? \new_[2652]_  : \new_[4986]_ ;
  assign \new_[1906]_  = ~\new_[2959]_  | ~\new_[2402]_ ;
  assign \new_[1907]_  = \new_[2883]_  ? \new_[2659]_  : \new_[2622]_ ;
  assign \new_[1908]_  = \new_[2884]_  ? \new_[2646]_  : \new_[3114]_ ;
  assign \new_[1909]_  = \new_[1866]_  ? \new_[2647]_  : \new_[19684]_ ;
  assign n1803 = \new_[1342]_  ^ \new_[2634]_ ;
  assign n1808 = \new_[19547]_  ^ \new_[3130]_ ;
  assign \new_[1912]_  = \new_[17745]_  ^ \new_[2654]_ ;
  assign n1798 = \new_[1349]_  ^ \new_[3123]_ ;
  assign \new_[1914]_  = ~\new_[2119]_ ;
  assign \new_[1915]_  = \new_[2531]_  ? \new_[2723]_  : \new_[2765]_ ;
  assign \new_[1916]_  = ~\new_[2883]_  | ~\new_[2398]_ ;
  assign \new_[1917]_  = ~\new_[2398]_  | ~\new_[3689]_ ;
  assign \new_[1918]_  = ~\new_[2637]_  | ~\new_[2362]_ ;
  assign \new_[1919]_  = \new_[2552]_  ^ \new_[2718]_ ;
  assign \new_[1920]_  = ~\new_[2125]_ ;
  assign \new_[1921]_  = \\u0_w_reg[1][12] ;
  assign \new_[1922]_  = \new_[3119]_  ? \new_[2717]_  : \new_[2889]_ ;
  assign \new_[1923]_  = \new_[21370]_  ? \new_[20545]_  : \new_[3122]_ ;
  assign n1683 = \key[99]  ? \new_[19649]_  : \new_[2693]_ ;
  assign n1678 = \key[67]  ? \new_[19649]_  : \new_[2692]_ ;
  assign n1688 = \key[3]  ? \new_[19649]_  : \new_[2696]_ ;
  assign \new_[1927]_  = \new_[3310]_  ? \new_[2719]_  : \new_[3120]_ ;
  assign \new_[1928]_  = \\u0_w_reg[3][25] ;
  assign \new_[1929]_  = \\u0_w_reg[0][25] ;
  assign \new_[1930]_  = \new_[18431]_  ^ \new_[2695]_ ;
  assign \new_[1931]_  = \new_[3226]_  ? \new_[2708]_  : \new_[3018]_ ;
  assign \new_[1932]_  = \new_[1426]_  ? \new_[2722]_  : \new_[19651]_ ;
  assign \new_[1933]_  = ~\new_[3086]_  | ~\new_[2445]_ ;
  assign \new_[1934]_  = ~\new_[2446]_  | ~\new_[2289]_ ;
  assign \new_[1935]_  = ~\new_[2428]_  | ~\new_[2719]_ ;
  assign \new_[1936]_  = ~\new_[2340]_  | ~\new_[2426]_ ;
  assign \new_[1937]_  = ~\new_[2444]_  | ~\new_[3121]_ ;
  assign \new_[1938]_  = ~\new_[2449]_  | ~\new_[2987]_ ;
  assign \new_[1939]_  = ~\new_[2448]_  | ~\new_[2986]_ ;
  assign \new_[1940]_  = ~\new_[2458]_  | ~\new_[2754]_ ;
  assign \new_[1941]_  = ~\new_[2457]_  | ~\new_[2990]_ ;
  assign \new_[1942]_  = ~\new_[2455]_  | ~\new_[2989]_ ;
  assign \new_[1943]_  = ~\new_[2454]_  | ~\new_[2988]_ ;
  assign n1693 = \new_[2529]_  ? n3423 : \key[36] ;
  assign n1698 = \key[92]  ? \new_[19649]_  : \new_[2534]_ ;
  assign n1703 = \key[28]  ? \new_[19649]_  : \new_[2535]_ ;
  assign \new_[1947]_  = ~\new_[2676]_  | ~\new_[2418]_ ;
  assign \new_[1948]_  = ~\new_[2142]_ ;
  assign \new_[1949]_  = \new_[3345]_  ? \new_[2648]_  : \new_[3545]_ ;
  assign \new_[1950]_  = \new_[1868]_  ? \new_[2649]_  : \new_[19575]_ ;
  assign \new_[1951]_  = ~\new_[2417]_  | ~\new_[2675]_ ;
  assign \new_[1952]_  = \new_[2617]_  ^ \new_[2913]_ ;
  assign \new_[1953]_  = \new_[2291]_  ? \new_[2651]_  : \new_[19590]_ ;
  assign \new_[1954]_  = \new_[2950]_  ^ \new_[2657]_ ;
  assign \new_[1955]_  = ~\new_[2409]_  | ~\new_[2411]_ ;
  assign \new_[1956]_  = ~\new_[2412]_  | ~\new_[2672]_ ;
  assign \new_[1957]_  = ~\new_[2673]_  | ~\new_[2413]_ ;
  assign \new_[1958]_  = \new_[3066]_  ? \new_[2549]_  : \new_[3266]_ ;
  assign \new_[1959]_  = \new_[3261]_  ? \new_[2550]_  : \new_[3409]_ ;
  assign \new_[1960]_  = ~\new_[2156]_ ;
  assign n1713 = \key[96]  ? \new_[19614]_  : \new_[2558]_ ;
  assign n1723 = \key[112]  ? \new_[19649]_  : \new_[2559]_ ;
  assign n1728 = \key[64]  ? \new_[19614]_  : \new_[2560]_ ;
  assign \new_[1964]_  = \new_[3169]_  ? \new_[2663]_  : \new_[2946]_ ;
  assign n1738 = \key[80]  ? \new_[19649]_  : \new_[2561]_ ;
  assign \new_[1966]_  = ~\new_[3344]_  | ~\new_[2400]_ ;
  assign n1733 = \key[0]  ? \new_[19614]_  : \new_[2563]_ ;
  assign n1743 = \key[16]  ? \new_[19614]_  : \new_[2564]_ ;
  assign \new_[1969]_  = ~\new_[2706]_  | ~\new_[2394]_ ;
  assign n1748 = \new_[1426]_  ^ \new_[3204]_ ;
  assign \new_[1971]_  = \new_[2948]_  ? \new_[2681]_  : \new_[2703]_ ;
  assign \new_[1972]_  = ~\new_[2390]_  | ~\new_[2655]_ ;
  assign \new_[1973]_  = \new_[3371]_  ? \new_[2574]_  : \new_[3204]_ ;
  assign \new_[1974]_  = \new_[3017]_  ? \new_[2536]_  : \new_[2788]_ ;
  assign \new_[1975]_  = ~\new_[2176]_ ;
  assign \new_[1976]_  = ~\new_[2178]_ ;
  assign \new_[1977]_  = ~\new_[2179]_ ;
  assign \new_[1978]_  = ~\new_[3160]_  | ~\new_[2474]_ ;
  assign \new_[1979]_  = \new_[3130]_  ? \new_[2547]_  : \new_[3329]_ ;
  assign \new_[1980]_  = ~\new_[2404]_  | ~\new_[2403]_ ;
  assign \new_[1981]_  = \new_[3317]_  ? \new_[2572]_  : \new_[3514]_ ;
  assign n1718 = \new_[19305]_  ^ \new_[21613]_ ;
  assign n1708 = \new_[1341]_  ^ \new_[2750]_ ;
  assign \new_[1984]_  = ~\new_[20974]_ ;
  assign \new_[1985]_  = ~\new_[2408]_  | ~\new_[2674]_ ;
  assign \new_[1986]_  = ~\new_[2416]_  | ~\new_[2677]_ ;
  assign \new_[1987]_  = \new_[3651]_  ? \new_[2697]_  : \new_[3690]_ ;
  assign \new_[1988]_  = ~\new_[2406]_  | ~\new_[2669]_ ;
  assign \new_[1989]_  = \new_[3123]_  ? \new_[2578]_  : \new_[3313]_ ;
  assign \new_[1990]_  = ~\new_[2419]_  | ~\new_[2678]_ ;
  assign \new_[1991]_  = ~\new_[2407]_  | ~\new_[2670]_ ;
  assign \new_[1992]_  = \new_[3513]_  ^ \new_[2579]_ ;
  assign \new_[1993]_  = ~\new_[2410]_  | ~\new_[2671]_ ;
  assign \new_[1994]_  = ~\new_[21481]_  | ~\new_[2515]_ ;
  assign \new_[1995]_  = ~\new_[2601]_  | ~\new_[2279]_ ;
  assign \new_[1996]_  = ~\new_[2603]_  | ~\new_[2283]_ ;
  assign \new_[1997]_  = ~\new_[2604]_  | ~\new_[2285]_ ;
  assign \new_[1998]_  = ~\new_[2513]_  | ~\new_[2748]_ ;
  assign \new_[1999]_  = \new_[3243]_  ? \new_[2735]_  : \new_[3396]_ ;
  assign \new_[2000]_  = ~\new_[2213]_ ;
  assign \new_[2001]_  = ~\new_[2215]_ ;
  assign \new_[2002]_  = ~\new_[2508]_  | (~\new_[20403]_  & ~\new_[3519]_ );
  assign \new_[2003]_  = ~\new_[20321]_ ;
  assign \new_[2004]_  = ~\new_[2216]_ ;
  assign \new_[2005]_  = ~\new_[2218]_ ;
  assign \new_[2006]_  = \new_[1744]_  ? \new_[2736]_  : \new_[19737]_ ;
  assign n1758 = \new_[1241]_  ^ \new_[2596]_ ;
  assign \new_[2008]_  = ~\new_[2223]_ ;
  assign \new_[2009]_  = ~\new_[2224]_ ;
  assign \new_[2010]_  = ~\new_[2225]_ ;
  assign \new_[2011]_  = ~\new_[2503]_  | ~\new_[2741]_ ;
  assign n1753 = \new_[1863]_  ^ \new_[3052]_ ;
  assign n1773 = \new_[1921]_  ^ \new_[3053]_ ;
  assign \new_[2014]_  = ~\new_[2507]_  | ~\new_[2747]_ ;
  assign \new_[2015]_  = \new_[2755]_  ^ \new_[2704]_ ;
  assign \new_[2016]_  = ~\new_[21367]_ ;
  assign \new_[2017]_  = ~\new_[2495]_  | ~\new_[2494]_ ;
  assign \new_[2018]_  = ~\new_[2496]_  & (~\new_[2878]_  | ~\new_[20052]_ );
  assign \new_[2019]_  = ~\new_[2497]_  | ~\new_[2498]_ ;
  assign \new_[2020]_  = \new_[2885]_  ? \new_[20403]_  : \new_[2624]_ ;
  assign \new_[2021]_  = ~\new_[2504]_  | ~\new_[2742]_ ;
  assign \new_[2022]_  = \new_[2887]_  ? \new_[20327]_  : \new_[2626]_ ;
  assign \new_[2023]_  = ~\new_[2235]_ ;
  assign \new_[2024]_  = \new_[2886]_  ? \new_[21121]_  : \new_[2625]_ ;
  assign \new_[2025]_  = \new_[20667]_  ? \new_[2633]_  : \new_[2995]_ ;
  assign \new_[2026]_  = ~\new_[2505]_  | ~\new_[2744]_ ;
  assign \new_[2027]_  = \new_[3062]_  ? \new_[2537]_  : \new_[2848]_ ;
  assign \new_[2028]_  = ~\new_[2499]_  | ~\new_[2493]_ ;
  assign \new_[2029]_  = \new_[2623]_  ? \new_[20646]_  : \new_[3116]_ ;
  assign \new_[2030]_  = ~\new_[2276]_  | ~\new_[3032]_ ;
  assign \new_[2031]_  = \new_[2878]_  ? \new_[3079]_  : \new_[2621]_ ;
  assign \new_[2032]_  = ~\new_[2447]_  | ~\new_[2270]_ ;
  assign \new_[2033]_  = \new_[2850]_  ? \new_[2566]_  : \new_[2597]_ ;
  assign \new_[2034]_  = ~\new_[2488]_  | ~\new_[2734]_ ;
  assign \new_[2035]_  = ~\new_[2491]_  | ~\new_[2492]_ ;
  assign n1763 = \new_[1664]_  ^ \new_[3074]_ ;
  assign n1768 = \new_[1345]_  ^ \new_[2589]_ ;
  assign \new_[2038]_  = ~\new_[2752]_  | ~\new_[2516]_ ;
  assign \new_[2039]_  = ~\new_[2248]_ ;
  assign \new_[2040]_  = \new_[19184]_  ? \new_[2628]_  : \new_[18519]_ ;
  assign \new_[2041]_  = ~\new_[2730]_  | ~\new_[2485]_ ;
  assign \new_[2042]_  = ~\new_[2249]_ ;
  assign \new_[2043]_  = \new_[3455]_  ? \new_[20331]_  : \new_[3287]_ ;
  assign \new_[2044]_  = \new_[3057]_  ? \new_[2632]_  : \new_[3251]_ ;
  assign \new_[2045]_  = ~\new_[3066]_  | ~\new_[2335]_ ;
  assign \new_[2046]_  = ~\new_[3409]_  | ~\new_[2336]_ ;
  assign \new_[2047]_  = ~\new_[2809]_  | ~\new_[2476]_ ;
  assign \new_[2048]_  = ~\new_[3297]_  | ~\new_[2337]_ ;
  assign \new_[2049]_  = ~\new_[2335]_  | ~\new_[3537]_ ;
  assign \new_[2050]_  = ~\new_[2266]_ ;
  assign \new_[2051]_  = ~\new_[2267]_ ;
  assign \new_[2052]_  = ~\new_[2268]_ ;
  assign \text_out[41]  = \\text_out_reg[41] ;
  assign n1848 = \new_[1347]_  ^ \new_[2835]_ ;
  assign \new_[2055]_  = ~\new_[2585]_  | (~\new_[3116]_  & ~\new_[3315]_ );
  assign \new_[2056]_  = ~\new_[2586]_  | (~\new_[3108]_  & ~\new_[20053]_ );
  assign \new_[2057]_  = ~\new_[2587]_  & (~\new_[21276]_  | ~\new_[19993]_ );
  assign \new_[2058]_  = \new_[3459]_  ? \new_[2852]_  : \new_[3288]_ ;
  assign n2018 = \new_[19025]_  ^ \new_[2884]_ ;
  assign \new_[2060]_  = ~\new_[2279]_ ;
  assign \new_[2061]_  = ~\new_[2584]_  & (~\new_[3634]_  | ~\new_[19993]_ );
  assign \text_out[1]  = \\text_out_reg[1] ;
  assign \text_out[7]  = \\text_out_reg[7] ;
  assign \text_out[38]  = \\text_out_reg[38] ;
  assign \text_out[36]  = \\text_out_reg[36] ;
  assign \text_out[33]  = \\text_out_reg[33] ;
  assign \text_out[39]  = \\text_out_reg[39] ;
  assign \new_[2068]_  = ~\new_[2289]_ ;
  assign \text_out[68]  = \\text_out_reg[68] ;
  assign \text_out[70]  = \\text_out_reg[70] ;
  assign \text_out[71]  = \\text_out_reg[71] ;
  assign \new_[2072]_  = ~\new_[2582]_  | ~\new_[2828]_ ;
  assign \text_out[50]  = \\text_out_reg[50] ;
  assign \text_out[59]  = \\text_out_reg[59] ;
  assign \text_out[91]  = \\text_out_reg[91] ;
  assign \text_out[40]  = \\text_out_reg[40] ;
  assign \text_out[72]  = \\text_out_reg[72] ;
  assign \new_[2078]_  = \\u0_w_reg[0][4] ;
  assign \new_[2079]_  = \\u0_w_reg[1][4] ;
  assign \new_[2080]_  = \\u0_w_reg[3][4] ;
  assign \text_out[9]  = \\text_out_reg[9] ;
  assign \text_out[31]  = \\text_out_reg[31] ;
  assign \text_out[102]  = \\text_out_reg[102] ;
  assign \text_out[55]  = \\text_out_reg[55] ;
  assign \text_out[54]  = \\text_out_reg[54] ;
  assign \text_out[90]  = \\text_out_reg[90] ;
  assign \text_out[119]  = \\text_out_reg[119] ;
  assign \text_out[22]  = \\text_out_reg[22] ;
  assign \text_out[103]  = \\text_out_reg[103] ;
  assign \text_out[15]  = \\text_out_reg[15] ;
  assign \text_out[14]  = \\text_out_reg[14] ;
  assign \text_out[92]  = \\text_out_reg[92] ;
  assign \text_out[116]  = \\text_out_reg[116] ;
  assign \text_out[66]  = \\text_out_reg[66] ;
  assign \new_[2095]_  = ~\new_[2583]_  | ~\new_[2831]_ ;
  assign \new_[2096]_  = ~\new_[2827]_  | (~\new_[3487]_  & ~\new_[2878]_ );
  assign n2003 = \new_[19700]_  ^ \new_[21595]_ ;
  assign n1998 = \new_[1353]_  ^ \new_[3288]_ ;
  assign n2013 = \new_[19761]_  ^ \new_[3286]_ ;
  assign n2008 = \new_[1669]_  ^ \new_[3291]_ ;
  assign \new_[2101]_  = ~\new_[2323]_ ;
  assign \new_[2102]_  = ~\new_[20888]_  | ~\new_[3626]_ ;
  assign \new_[2103]_  = ~\new_[3118]_  | ~\new_[3702]_ ;
  assign \new_[2104]_  = ~\new_[3117]_  | ~\new_[20053]_ ;
  assign n2068 = \new_[2906]_  ? \new_[19338]_  : \key[39] ;
  assign \new_[2106]_  = ~\new_[2334]_ ;
  assign \new_[2107]_  = ~\new_[2335]_ ;
  assign n1863 = \new_[2918]_  ? n3423 : \key[50] ;
  assign n1868 = \new_[2919]_  ? n3423 : \key[34] ;
  assign \new_[2110]_  = ~\new_[2340]_ ;
  assign \new_[2111]_  = ~\new_[2724]_  | ~\new_[2664]_ ;
  assign \new_[2112]_  = ~\new_[2341]_ ;
  assign n2023 = \new_[1350]_  ^ \new_[2896]_ ;
  assign n2028 = \new_[19121]_  ^ \new_[2897]_ ;
  assign \new_[2115]_  = ~\new_[20270]_  | ~\new_[3476]_ ;
  assign n2033 = \new_[18970]_  ^ \new_[3317]_ ;
  assign n2038 = \new_[1668]_  ^ \new_[3318]_ ;
  assign \new_[2118]_  = ~\new_[2876]_  | ~\new_[2619]_ ;
  assign \new_[2119]_  = \new_[3001]_  ? \new_[2957]_  : \new_[2764]_ ;
  assign \new_[2120]_  = ~\new_[2345]_ ;
  assign \new_[2121]_  = ~\new_[2661]_  | ~\new_[2622]_ ;
  assign \new_[2122]_  = ~\new_[2661]_  | ~\new_[3647]_ ;
  assign \new_[2123]_  = ~\new_[2642]_  | ~\new_[8023]_ ;
  assign \new_[2124]_  = ~\new_[2641]_  | ~\new_[9256]_ ;
  assign \new_[2125]_  = \new_[2867]_  ? \new_[2921]_  : \new_[3087]_ ;
  assign n1873 = \new_[2933]_  ? \new_[19479]_  : \key[55] ;
  assign n2043 = \new_[1929]_  ^ \new_[3334]_ ;
  assign \text_out[11]  = \\text_out_reg[11] ;
  assign \text_out[34]  = \\text_out_reg[34] ;
  assign n1843 = \new_[19184]_  ^ \new_[3347]_ ;
  assign n2063 = \new_[2960]_  ? ld : \key[33] ;
  assign n2048 = \new_[1719]_  ^ \new_[3336]_ ;
  assign \new_[2133]_  = ~\new_[2866]_  | ~\new_[2702]_ ;
  assign \new_[2134]_  = \new_[3170]_  ^ \new_[2801]_ ;
  assign \new_[2135]_  = ~\new_[2545]_  | ~\new_[2682]_ ;
  assign \new_[2136]_  = ~\new_[2546]_  | ~\new_[2683]_ ;
  assign \new_[2137]_  = ~\new_[2689]_  | ~\new_[21370]_ ;
  assign n1878 = \new_[2763]_  ? \new_[19472]_  : \key[52] ;
  assign \text_out[27]  = \\text_out_reg[27] ;
  assign n2053 = \new_[2766]_  ? \new_[19414]_  : \key[124] ;
  assign n1883 = \new_[2769]_  ? \new_[19371]_  : \key[60] ;
  assign \new_[2142]_  = \new_[3472]_  ? \new_[2779]_  : \new_[3297]_ ;
  assign \new_[2143]_  = \new_[10730]_  ^ \new_[2799]_ ;
  assign n1588 = \new_[17844]_  ^ \new_[2767]_ ;
  assign \new_[2145]_  = \new_[18471]_  ^ \new_[21668]_ ;
  assign \new_[2146]_  = \new_[3153]_  ^ \new_[2915]_ ;
  assign \new_[2147]_  = \new_[7053]_  ^ \new_[2802]_ ;
  assign \new_[2148]_  = \new_[9257]_  ^ \new_[21667]_ ;
  assign \new_[2149]_  = \new_[3318]_  ? \new_[2914]_  : \new_[3516]_ ;
  assign \new_[2150]_  = \new_[1345]_  ^ \new_[2985]_ ;
  assign \new_[2151]_  = \new_[17908]_  ^ \new_[2985]_ ;
  assign \new_[2152]_  = \new_[11488]_  ^ \new_[2985]_ ;
  assign \new_[2153]_  = \new_[3125]_  ? \new_[2775]_  : \new_[2896]_ ;
  assign n1838 = \new_[19114]_  ^ \new_[2762]_ ;
  assign \new_[2155]_  = \new_[3127]_  ? \new_[3004]_  : \new_[2897]_ ;
  assign \new_[2156]_  = \new_[3405]_  ? \new_[2778]_  : \new_[3570]_ ;
  assign n1888 = \key[106]  ? \new_[19614]_  : \new_[2787]_ ;
  assign n1923 = \key[74]  ? \new_[19649]_  : \new_[2789]_ ;
  assign \new_[2159]_  = ~\new_[3162]_  | ~\new_[2662]_ ;
  assign n1933 = \key[10]  ? \new_[19614]_  : \new_[2793]_ ;
  assign \new_[2161]_  = ~\new_[2951]_  | ~\new_[2658]_ ;
  assign n2058 = \key[110]  ? \new_[19649]_  : \new_[2797]_ ;
  assign n1913 = \key[78]  ? \new_[19649]_  : \new_[2804]_ ;
  assign \new_[2164]_  = \new_[3622]_  ? \new_[2798]_  : \new_[21276]_ ;
  assign n1853 = \key[14]  ? \new_[19649]_  : \new_[2803]_ ;
  assign \new_[2166]_  = ~\new_[2665]_  | (~\new_[3204]_  & ~\new_[19775]_ );
  assign \new_[2167]_  = ~\new_[2666]_  | (~\new_[3204]_  & ~\new_[19799]_ );
  assign n1893 = \key[109]  ? \new_[19649]_  : \new_[2810]_ ;
  assign n1898 = \key[111]  ? \new_[19649]_  : \new_[2811]_ ;
  assign n1903 = \key[104]  ? \new_[19614]_  : \new_[2812]_ ;
  assign n1908 = \key[77]  ? \new_[19614]_  : \new_[2813]_ ;
  assign n1918 = \key[79]  ? \new_[19614]_  : \new_[2815]_ ;
  assign n1928 = \key[72]  ? \new_[19614]_  : \new_[2816]_ ;
  assign n1938 = \key[13]  ? \new_[19614]_  : \new_[2819]_ ;
  assign n1943 = \key[15]  ? \new_[19649]_  : \new_[2820]_ ;
  assign \new_[2176]_  = \new_[3542]_  ? \new_[2944]_  : \new_[3341]_ ;
  assign n1948 = \key[8]  ? \new_[19614]_  : \new_[2821]_ ;
  assign \new_[2178]_  = ~\new_[2667]_  | ~\new_[2668]_ ;
  assign \new_[2179]_  = \new_[21487]_  ? \new_[2777]_  : \new_[21486]_ ;
  assign \new_[2180]_  = \new_[18305]_  ^ \new_[2790]_ ;
  assign \new_[2181]_  = \new_[19143]_  ^ \new_[2794]_ ;
  assign \new_[2182]_  = \new_[17732]_  ^ \new_[2791]_ ;
  assign \new_[2183]_  = ~\new_[2929]_  | ~\new_[2726]_ ;
  assign \new_[2184]_  = \new_[18426]_  ^ \new_[2800]_ ;
  assign \new_[2185]_  = \new_[3531]_  ? \new_[2984]_  : \new_[3632]_ ;
  assign n1953 = \new_[18390]_  ^ \new_[2982]_ ;
  assign n1833 = \new_[19340]_  ^ \new_[21708]_ ;
  assign \new_[2188]_  = \new_[18188]_  ^ \new_[2817]_ ;
  assign \new_[2189]_  = \new_[18696]_  ^ \new_[2818]_ ;
  assign \new_[2190]_  = ~\new_[2398]_ ;
  assign \new_[2191]_  = \new_[2840]_  ? \new_[2984]_  : \new_[20250]_ ;
  assign n1858 = \new_[19686]_  ^ \new_[21198]_ ;
  assign \new_[2193]_  = \new_[20250]_  ? \new_[2984]_  : \new_[2840]_ ;
  assign \new_[2194]_  = \new_[3317]_  ? \new_[2822]_  : \new_[3514]_ ;
  assign \new_[2195]_  = \new_[3318]_  ? \new_[2823]_  : \new_[3516]_ ;
  assign \new_[2196]_  = ~\new_[21577]_  | ~\new_[2749]_ ;
  assign \new_[2197]_  = ~\new_[2872]_  | ~\new_[2751]_ ;
  assign \new_[2198]_  = \new_[3465]_  ? \new_[2943]_  : \new_[3291]_ ;
  assign \new_[2199]_  = ~\new_[2871]_  | ~\new_[2750]_ ;
  assign \new_[2200]_  = ~\new_[3525]_  | ~\new_[2542]_ ;
  assign \new_[2201]_  = ~\new_[3323]_  | ~\new_[2541]_ ;
  assign \new_[2202]_  = ~\new_[3316]_  | ~\new_[2542]_ ;
  assign \new_[2203]_  = ~\new_[3513]_  | ~\new_[2541]_ ;
  assign \new_[2204]_  = ~\new_[2634]_  | ~\new_[2772]_ ;
  assign \new_[2205]_  = ~\new_[2855]_  | ~\new_[2553]_ ;
  assign \new_[2206]_  = ~\new_[2856]_  | ~\new_[2555]_ ;
  assign \new_[2207]_  = ~\new_[2857]_  | ~\new_[2533]_ ;
  assign \new_[2208]_  = ~\new_[2686]_  | ~\new_[2935]_ ;
  assign \new_[2209]_  = \new_[3541]_  ? \new_[2845]_  : \new_[3644]_ ;
  assign \text_out[2]  = \\text_out_reg[2] ;
  assign \new_[2211]_  = \new_[3642]_  ? \new_[2843]_  : \new_[3540]_ ;
  assign \new_[2212]_  = \new_[3689]_  ? \new_[3271]_  : \new_[21375]_ ;
  assign \new_[2213]_  = \new_[3672]_  ? \new_[2843]_  : \new_[3625]_ ;
  assign \new_[2214]_  = ~\new_[2428]_ ;
  assign \new_[2215]_  = \new_[3506]_  ? \new_[3271]_  : \new_[3507]_ ;
  assign \new_[2216]_  = ~\new_[2745]_  | (~\new_[21121]_  & ~\new_[3521]_ );
  assign \new_[2217]_  = ~\new_[2431]_ ;
  assign \new_[2218]_  = ~\new_[2746]_  | (~\new_[20646]_  & ~\new_[3315]_ );
  assign \new_[2219]_  = \new_[2972]_  ^ \new_[3016]_ ;
  assign \new_[2220]_  = ~\new_[2713]_  | ~\new_[2954]_ ;
  assign \new_[2221]_  = \new_[3123]_  ? \new_[2970]_  : \new_[3313]_ ;
  assign \new_[2222]_  = \new_[3408]_  ? \new_[2845]_  : \new_[19840]_ ;
  assign \new_[2223]_  = ~\new_[2738]_  | ~\new_[2739]_ ;
  assign \new_[2224]_  = ~\new_[2740]_  | ~\new_[2971]_ ;
  assign \new_[2225]_  = ~\new_[2444]_ ;
  assign \new_[2226]_  = ~\new_[2446]_ ;
  assign n1973 = \new_[1666]_  ^ \new_[20052]_ ;
  assign n2078 = \new_[1418]_  ^ \new_[20403]_ ;
  assign \new_[2229]_  = \new_[3585]_  ? \new_[20403]_  : \new_[3584]_ ;
  assign \new_[2230]_  = \new_[3584]_  ? \new_[20403]_  : \new_[3585]_ ;
  assign \new_[2231]_  = \new_[3108]_  ? \new_[20052]_  : \new_[3292]_ ;
  assign \new_[2232]_  = ~\new_[2461]_ ;
  assign \new_[2233]_  = ~\new_[2462]_ ;
  assign \new_[2234]_  = ~\new_[2733]_  | (~\new_[21487]_  & ~\new_[3130]_ );
  assign \new_[2235]_  = ~\new_[2743]_  | ~\new_[2974]_ ;
  assign \new_[2236]_  = ~\new_[2814]_  | ~\new_[2544]_ ;
  assign n1988 = \new_[1186]_  ^ \new_[2845]_ ;
  assign n1993 = \new_[19520]_  ^ \new_[3271]_ ;
  assign \new_[2239]_  = ~\new_[2707]_  | ~\new_[2522]_ ;
  assign n1958 = \new_[1088]_  ^ \new_[2843]_ ;
  assign \new_[2241]_  = ~\new_[2471]_ ;
  assign n1968 = \new_[19043]_  ^ \new_[2851]_ ;
  assign \new_[2243]_  = ~\new_[2964]_  | (~\new_[3266]_  & ~\new_[2878]_ );
  assign n1983 = \new_[18699]_  ^ \new_[2841]_ ;
  assign n2073 = \new_[19513]_  ^ \new_[3249]_ ;
  assign n1963 = \new_[1477]_  ^ \new_[3275]_ ;
  assign n1978 = \new_[19387]_  ^ \new_[3278]_ ;
  assign \new_[2248]_  = ~\new_[2729]_  | ~\new_[2961]_ ;
  assign \new_[2249]_  = ~\new_[2731]_  | ~\new_[2962]_ ;
  assign \new_[2250]_  = ~\new_[2963]_  | ~\new_[2732]_ ;
  assign \new_[2251]_  = ~\new_[3074]_  | ~\new_[21482]_ ;
  assign \new_[2252]_  = ~\new_[3275]_  | ~\new_[21577]_ ;
  assign \new_[2253]_  = ~\new_[3060]_  | ~\new_[20270]_ ;
  assign \new_[2254]_  = ~\new_[2600]_  | ~\new_[21474]_ ;
  assign \new_[2255]_  = \new_[3385]_  ^ \new_[2853]_ ;
  assign \new_[2256]_  = ~\new_[2600]_  | ~\new_[3273]_ ;
  assign \new_[2257]_  = ~\new_[3261]_  | ~\new_[2605]_ ;
  assign \new_[2258]_  = ~\new_[3570]_  | ~\new_[2606]_ ;
  assign \new_[2259]_  = ~\new_[2607]_  | ~\new_[3639]_ ;
  assign \new_[2260]_  = ~\new_[2577]_  | ~\new_[2727]_ ;
  assign \new_[2261]_  = ~\new_[3472]_  | ~\new_[2607]_ ;
  assign \new_[2262]_  = ~\new_[3111]_  | ~\new_[3334]_  | ~\new_[2882]_ ;
  assign \new_[2263]_  = ~\new_[2605]_  | ~\new_[3333]_ ;
  assign \new_[2264]_  = \new_[2518]_ ;
  assign \text_out[28]  = \\text_out_reg[28] ;
  assign \new_[2266]_  = ~\new_[2591]_  | (~\new_[3117]_  & ~\new_[3537]_ );
  assign \new_[2267]_  = ~\new_[2592]_  | (~\new_[3118]_  & ~\new_[3637]_ );
  assign \new_[2268]_  = ~\new_[2593]_  | (~\new_[20888]_  & ~\new_[3635]_ );
  assign \new_[2269]_  = ~\new_[2521]_ ;
  assign \new_[2270]_  = ~\new_[2522]_ ;
  assign \text_out[25]  = \\text_out_reg[25] ;
  assign \new_[2272]_  = \\u0_w_reg[3][7] ;
  assign \new_[2273]_  = (~\new_[3669]_  | ~\new_[21596]_ ) & (~\new_[3610]_  | ~\new_[21598]_ );
  assign \new_[2274]_  = (~\new_[3616]_  | ~\new_[3453]_ ) & (~\new_[3501]_  | ~\new_[3286]_ );
  assign \new_[2275]_  = ~\new_[2838]_  | ~\new_[2839]_ ;
  assign \new_[2276]_  = ~\new_[2544]_ ;
  assign \new_[2277]_  = ~\new_[2836]_  | ~\new_[3049]_ ;
  assign \new_[2278]_  = ~\new_[2835]_  | ~\new_[19618]_ ;
  assign \new_[2279]_  = ~\new_[2829]_  | ~\new_[3042]_ ;
  assign \new_[2280]_  = ~\new_[2835]_  | ~\new_[19593]_ ;
  assign \new_[2281]_  = ~\new_[2830]_  | (~\new_[3299]_  & ~\new_[19626]_ );
  assign \new_[2282]_  = ~\new_[2835]_  | ~\new_[19710]_ ;
  assign \new_[2283]_  = ~\new_[2555]_ ;
  assign \text_out[58]  = \\text_out_reg[58] ;
  assign \new_[2285]_  = ~\new_[2533]_ ;
  assign \text_out[122]  = \\text_out_reg[122] ;
  assign \text_out[3]  = \\text_out_reg[3] ;
  assign \new_[2288]_  = \\u0_w_reg[1][18] ;
  assign \new_[2289]_  = ~\new_[2832]_  | (~\new_[3300]_  & ~\new_[19720]_ );
  assign \text_out[65]  = \\text_out_reg[65] ;
  assign \new_[2291]_  = \\u0_w_reg[1][7] ;
  assign \new_[2292]_  = ~\new_[2833]_  | (~\new_[3300]_  & ~\new_[19793]_ );
  assign \new_[2293]_  = \\u0_w_reg[0][2] ;
  assign \new_[2294]_  = \\u0_w_reg[1][2] ;
  assign \new_[2295]_  = \\u0_w_reg[3][18] ;
  assign \new_[2296]_  = \\u0_w_reg[3][2] ;
  assign \new_[2297]_  = \\u0_w_reg[0][23] ;
  assign \new_[2298]_  = \\u0_w_reg[3][23] ;
  assign \text_out[107]  = \\text_out_reg[107] ;
  assign \new_[2300]_  = \\u0_w_reg[0][20] ;
  assign \new_[2301]_  = \\u0_w_reg[1][20] ;
  assign \new_[2302]_  = \\u0_w_reg[3][20] ;
  assign \text_out[97]  = \\text_out_reg[97] ;
  assign \text_out[63]  = \\text_out_reg[63] ;
  assign \text_out[96]  = \\text_out_reg[96] ;
  assign \text_out[113]  = \\text_out_reg[113] ;
  assign \text_out[127]  = \\text_out_reg[127] ;
  assign \text_out[118]  = \\text_out_reg[118] ;
  assign \text_out[26]  = \\text_out_reg[26] ;
  assign \text_out[98]  = \\text_out_reg[98] ;
  assign \text_out[52]  = \\text_out_reg[52] ;
  assign \text_out[84]  = \\text_out_reg[84] ;
  assign n2083 = \new_[19397]_  ^ \new_[3116]_ ;
  assign \new_[2314]_  = ~\new_[2826]_  | ~\new_[3041]_ ;
  assign n2098 = \new_[1291]_  ^ \new_[3092]_ ;
  assign \new_[2316]_  = ~\new_[2567]_ ;
  assign \new_[2317]_  = \new_[19571]_  ? \new_[3092]_  : \new_[1088]_ ;
  assign \new_[2318]_  = ~\new_[2834]_  & (~\new_[3589]_  | ~\new_[3285]_ );
  assign \new_[2319]_  = ~\new_[2571]_ ;
  assign \new_[2320]_  = ~\new_[2573]_ ;
  assign \new_[2321]_  = ~\new_[2825]_  | (~\new_[3575]_  & ~\new_[21597]_ );
  assign n2238 = \new_[1663]_  ^ \new_[3455]_ ;
  assign \new_[2323]_  = ~\new_[2824]_  & (~\new_[3292]_  | ~\new_[3455]_ );
  assign \new_[2324]_  = ~\new_[2580]_ ;
  assign \new_[2325]_  = ~\new_[2581]_ ;
  assign \new_[2326]_  = ~\new_[2590]_ ;
  assign \new_[2327]_  = ~\new_[2859]_  | (~\new_[3298]_  & ~\new_[19714]_ );
  assign \new_[2328]_  = ~\new_[2595]_ ;
  assign \text_out[95]  = \\text_out_reg[95] ;
  assign \new_[2330]_  = ~\new_[2599]_ ;
  assign n2263 = \new_[2346]_  ^ \new_[3518]_ ;
  assign n2258 = \new_[19507]_  ^ \new_[21588]_ ;
  assign n2243 = \new_[2288]_  ^ \new_[3501]_ ;
  assign \new_[2334]_  = (~\new_[21589]_  | ~\new_[3329]_ ) & (~\new_[21587]_  | ~\new_[3129]_ );
  assign \new_[2335]_  = ~\new_[2882]_  | ~\new_[3111]_ ;
  assign \new_[2336]_  = ~\new_[2605]_ ;
  assign \new_[2337]_  = ~\new_[2607]_ ;
  assign n2253 = \new_[19308]_  ^ \new_[3124]_ ;
  assign \new_[2339]_  = ~\new_[2611]_ ;
  assign \new_[2340]_  = ~\new_[2880]_  | (~\new_[3328]_  & ~\new_[3509]_ );
  assign \new_[2341]_  = ~\new_[2881]_  | (~\new_[3329]_  & ~\new_[21276]_ );
  assign n2248 = \new_[18378]_  ^ \new_[3126]_ ;
  assign \new_[2343]_  = ~\new_[2847]_  | ~\new_[3475]_ ;
  assign \new_[2344]_  = \\u0_w_reg[0][7] ;
  assign \new_[2345]_  = ~\new_[3103]_  | ~\new_[2877]_ ;
  assign \new_[2346]_  = \\u0_w_reg[0][18] ;
  assign n2293 = \new_[3154]_  ? \new_[19338]_  : \key[121] ;
  assign n2118 = \key[89]  ? \new_[19649]_  : \new_[3155]_ ;
  assign n2113 = \new_[3156]_  ? \new_[19479]_  : \key[57] ;
  assign n2288 = \key[25]  ? \new_[19649]_  : \new_[3157]_ ;
  assign \new_[2351]_  = ~\new_[2902]_  | (~\new_[3347]_  & ~\new_[21276]_ );
  assign n2268 = \new_[1861]_  ^ \new_[3132]_ ;
  assign n2273 = \new_[19699]_  ^ \new_[3535]_ ;
  assign n2088 = \new_[16682]_  ^ \new_[3167]_ ;
  assign n2278 = \new_[1662]_  ^ \new_[3539]_ ;
  assign \new_[2356]_  = ~\new_[2899]_  | (~\new_[3348]_  & ~\new_[18877]_ );
  assign \new_[2357]_  = ~\new_[2900]_  | (~\new_[3347]_  & ~\new_[18449]_ );
  assign \new_[2358]_  = ~\new_[2901]_  | (~\new_[3347]_  & ~\new_[18391]_ );
  assign \new_[2359]_  = ~\new_[2773]_  | ~\new_[2926]_ ;
  assign \new_[2360]_  = ~\new_[2774]_  | ~\new_[2927]_ ;
  assign \new_[2361]_  = ~\new_[2941]_  | ~\new_[3122]_ ;
  assign \new_[2362]_  = ~\new_[2931]_  | ~\new_[2990]_ ;
  assign n2123 = \new_[2997]_  ? \new_[18703]_  : \key[108] ;
  assign n2283 = \new_[2998]_  ? \new_[18703]_  : \key[76] ;
  assign n2128 = \new_[3000]_  ? ld : \key[12] ;
  assign \new_[2366]_  = \new_[17538]_  ^ \new_[2999]_ ;
  assign \new_[2367]_  = \new_[10857]_  ^ \new_[3015]_ ;
  assign \new_[2368]_  = \new_[10731]_  ^ \new_[3005]_ ;
  assign \new_[2369]_  = \new_[18532]_  ^ \new_[3003]_ ;
  assign \new_[2370]_  = \new_[8252]_  ^ \new_[3020]_ ;
  assign \new_[2371]_  = \new_[7056]_  ^ \new_[3006]_ ;
  assign \new_[2372]_  = \new_[11486]_  ^ \new_[3003]_ ;
  assign \new_[2373]_  = \new_[19325]_  ? \new_[3210]_  : \new_[1346]_ ;
  assign \new_[2374]_  = ~\new_[2925]_  | ~\new_[3159]_ ;
  assign \new_[2375]_  = ~\new_[3161]_  | ~\new_[2932]_ ;
  assign \new_[2376]_  = ~\new_[2645]_ ;
  assign \new_[2377]_  = ~\new_[3166]_  | ~\new_[2940]_ ;
  assign n2133 = \new_[3023]_  ? \new_[19383]_  : \key[118] ;
  assign n2138 = \key[102]  ? \new_[19649]_  : \new_[3024]_ ;
  assign n2143 = \key[86]  ? \new_[19649]_  : \new_[3025]_ ;
  assign n2148 = \key[70]  ? \new_[19614]_  : \new_[3026]_ ;
  assign n2153 = \key[22]  ? \new_[19649]_  : \new_[3028]_ ;
  assign n2158 = \key[6]  ? \new_[19614]_  : \new_[3029]_ ;
  assign n2103 = \new_[1474]_  ^ \new_[3153]_ ;
  assign \new_[2385]_  = ~\new_[2916]_  | (~\new_[3340]_  & ~\new_[19552]_ );
  assign \new_[2386]_  = ~\new_[2917]_  | (~\new_[3340]_  & ~\new_[1346]_ );
  assign \new_[2387]_  = \new_[1426]_  ^ \new_[3375]_ ;
  assign \new_[2388]_  = \new_[17883]_  ^ \new_[3375]_ ;
  assign \new_[2389]_  = \new_[10502]_  ^ \new_[3375]_ ;
  assign \new_[2390]_  = ~\new_[3342]_  | ~\new_[2952]_ ;
  assign \new_[2391]_  = \new_[18422]_  ^ \new_[3027]_ ;
  assign \new_[2392]_  = \new_[17890]_  ^ \new_[3022]_ ;
  assign \new_[2393]_  = \new_[3633]_  ? \new_[3207]_  : \new_[3681]_ ;
  assign \new_[2394]_  = ~\new_[2658]_ ;
  assign \new_[2395]_  = \new_[3631]_  ? \new_[21613]_  : \new_[19902]_ ;
  assign \new_[2396]_  = ~\new_[3152]_  | ~\new_[2920]_ ;
  assign \new_[2397]_  = \new_[18105]_  ^ \new_[3031]_ ;
  assign \new_[2398]_  = ~\new_[2661]_ ;
  assign \new_[2399]_  = \new_[20185]_  ? \new_[3207]_  : \new_[3248]_ ;
  assign \new_[2400]_  = ~\new_[2662]_ ;
  assign \new_[2401]_  = ~\new_[20993]_  | ~\new_[2981]_ ;
  assign \new_[2402]_  = ~\new_[2664]_ ;
  assign \new_[2403]_  = ~\new_[2869]_  | ~\new_[3372]_ ;
  assign \new_[2404]_  = ~\new_[2868]_  | ~\new_[3205]_ ;
  assign \new_[2405]_  = ~\new_[21240]_  | ~\new_[2983]_ ;
  assign \new_[2406]_  = ~\new_[21198]_  | ~\new_[19774]_ ;
  assign \new_[2407]_  = ~\new_[2938]_  | ~\new_[1518]_ ;
  assign \new_[2408]_  = ~\new_[21707]_  | ~\new_[18829]_ ;
  assign \new_[2409]_  = ~\new_[3317]_  | ~\new_[2772]_ ;
  assign \new_[2410]_  = ~\new_[2938]_  | ~\new_[19598]_ ;
  assign \new_[2411]_  = ~\new_[3514]_  | ~\new_[2771]_ ;
  assign \new_[2412]_  = ~\new_[2770]_  | ~\new_[3318]_ ;
  assign \new_[2413]_  = ~\new_[3313]_  | ~\new_[3220]_ ;
  assign \new_[2414]_  = ~\new_[2898]_  | ~\new_[2771]_ ;
  assign \new_[2415]_  = ~\new_[3076]_  | ~\new_[2780]_ ;
  assign \new_[2416]_  = ~\new_[21707]_  | ~\new_[19563]_ ;
  assign \new_[2417]_  = ~\new_[2768]_  | ~\new_[12484]_ ;
  assign \new_[2418]_  = ~\new_[2863]_  | ~\new_[3215]_ ;
  assign \new_[2419]_  = ~\new_[21709]_  | ~\new_[19718]_ ;
  assign n2108 = \new_[1506]_  ^ \new_[3180]_ ;
  assign \new_[2421]_  = \new_[6250]_  ^ \new_[3064]_ ;
  assign \new_[2422]_  = \new_[1187]_  ? \new_[3180]_  : \new_[19124]_ ;
  assign \new_[2423]_  = ~\new_[2936]_  & (~\new_[3653]_  | ~\new_[3354]_ );
  assign \new_[2424]_  = ~\new_[2680]_ ;
  assign \new_[2425]_  = \new_[3687]_  ? \new_[3068]_  : \new_[3646]_ ;
  assign \new_[2426]_  = ~\new_[2684]_ ;
  assign \new_[2427]_  = ~\new_[2934]_  | (~\new_[3690]_  & ~\new_[3286]_ );
  assign \new_[2428]_  = \new_[3701]_  ? \new_[3069]_  : \new_[20329]_ ;
  assign \new_[2429]_  = ~\new_[2976]_  | (~\new_[20559]_  & ~\new_[20323]_ );
  assign \new_[2430]_  = ~\new_[2977]_  | (~\new_[3521]_  & ~\new_[3255]_ );
  assign \new_[2431]_  = \new_[3674]_  ? \new_[20270]_  : \new_[3672]_ ;
  assign \new_[2432]_  = ~\new_[2690]_ ;
  assign \new_[2433]_  = \new_[1238]_  ^ \new_[3064]_ ;
  assign \new_[2434]_  = ~\new_[2694]_ ;
  assign \new_[2435]_  = ~\new_[2949]_  | (~\new_[3355]_  & ~\new_[19726]_ );
  assign \new_[2436]_  = \new_[19628]_  ^ \new_[3064]_ ;
  assign \new_[2437]_  = ~\new_[2699]_ ;
  assign n2223 = \new_[1431]_  ^ \new_[3071]_ ;
  assign \new_[2439]_  = \new_[1430]_  ^ \new_[3059]_ ;
  assign \new_[2440]_  = ~\new_[2701]_ ;
  assign \new_[2441]_  = \new_[17741]_  ^ \new_[3059]_ ;
  assign \new_[2442]_  = \new_[1431]_  ^ \new_[3059]_ ;
  assign \new_[2443]_  = \new_[6165]_  ^ \new_[3059]_ ;
  assign \new_[2444]_  = ~\new_[2973]_  | ~\new_[3189]_ ;
  assign \new_[2445]_  = ~\new_[2702]_ ;
  assign \new_[2446]_  = \new_[3292]_  ? \new_[21332]_  : \new_[3108]_ ;
  assign \new_[2447]_  = ~\new_[2707]_ ;
  assign \new_[2448]_  = \new_[3587]_  ? \new_[21121]_  : \new_[3467]_ ;
  assign \new_[2449]_  = \new_[3467]_  ? \new_[21121]_  : \new_[3587]_ ;
  assign n2228 = \new_[1238]_  ^ \new_[3065]_ ;
  assign n2218 = \new_[1243]_  ^ \new_[20646]_ ;
  assign n2163 = \new_[1422]_  ^ \new_[21121]_ ;
  assign n2173 = \new_[1420]_  ^ \new_[20328]_ ;
  assign \new_[2454]_  = \new_[3583]_  ? \new_[20327]_  : \new_[3456]_ ;
  assign \new_[2455]_  = \new_[3456]_  ? \new_[20327]_  : \new_[3583]_ ;
  assign \new_[2456]_  = ~\new_[2717]_ ;
  assign \new_[2457]_  = \new_[3461]_  ? \new_[20646]_  : \new_[3290]_ ;
  assign \new_[2458]_  = \new_[3290]_  ? \new_[20646]_  : \new_[3461]_ ;
  assign \new_[2459]_  = ~\new_[2719]_ ;
  assign \new_[2460]_  = ~\new_[20545]_ ;
  assign \new_[2461]_  = ~\new_[2967]_  & (~\new_[3465]_  | ~\new_[20559]_ );
  assign \new_[2462]_  = ~\new_[2968]_  & (~\new_[3459]_  | ~\new_[3255]_ );
  assign n2168 = \new_[3093]_  ? \new_[19415]_  : \key[113] ;
  assign n2178 = \key[105]  ? \new_[19649]_  : \new_[3094]_ ;
  assign n2183 = \new_[3095]_  ? ld : \key[81] ;
  assign n2193 = \key[73]  ? \new_[19614]_  : \new_[3096]_ ;
  assign n2198 = \new_[3099]_  ? ld : \key[17] ;
  assign n2203 = \key[9]  ? \new_[19614]_  : \new_[3100]_ ;
  assign \new_[2469]_  = \new_[3083]_  ^ \new_[3302]_ ;
  assign n2213 = \new_[19124]_  ^ \new_[3068]_ ;
  assign \new_[2471]_  = \new_[3485]_  ? \new_[3101]_  : \new_[3603]_ ;
  assign n2233 = \new_[1877]_  ^ \new_[3409]_ ;
  assign \new_[2473]_  = \new_[3128]_  ? \new_[20250]_  : \new_[3327]_ ;
  assign \new_[2474]_  = ~\new_[2726]_ ;
  assign \new_[2475]_  = \new_[3326]_  ? \new_[3055]_  : \new_[3527]_ ;
  assign \new_[2476]_  = ~\new_[2727]_ ;
  assign \new_[2477]_  = \new_[3322]_  ? \new_[19978]_  : \new_[3524]_ ;
  assign \new_[2478]_  = ~\new_[3183]_  | ~\new_[2965]_ ;
  assign n2188 = \new_[1237]_  ^ \new_[3054]_ ;
  assign n2208 = \new_[19325]_  ^ \new_[3055]_ ;
  assign \new_[2481]_  = \new_[18503]_  ^ \new_[3090]_ ;
  assign \new_[2482]_  = \new_[18212]_  ^ \new_[3098]_ ;
  assign \new_[2483]_  = ~\new_[2978]_  | ~\new_[2975]_ ;
  assign n2093 = \new_[19549]_  ^ \new_[3016]_ ;
  assign \new_[2485]_  = ~\new_[2840]_  | ~\new_[21176]_ ;
  assign \new_[2486]_  = ~\new_[2979]_  | (~\new_[3224]_  & ~\new_[1288]_ );
  assign \new_[2487]_  = ~\new_[3277]_  | ~\new_[2872]_ ;
  assign \new_[2488]_  = ~\new_[3278]_  | ~\new_[2870]_ ;
  assign \new_[2489]_  = ~\new_[2980]_  | (~\new_[3224]_  & ~\new_[19605]_ );
  assign \new_[2490]_  = ~\new_[3073]_  | ~\new_[20993]_ ;
  assign \new_[2491]_  = ~\new_[3251]_  | ~\new_[2869]_ ;
  assign \new_[2492]_  = ~\new_[3057]_  | ~\new_[2868]_ ;
  assign \new_[2493]_  = ~\new_[2887]_  | ~\new_[20559]_ ;
  assign \new_[2494]_  = ~\new_[2885]_  | ~\new_[20052]_ ;
  assign \new_[2495]_  = \new_[2885]_  | \new_[20052]_ ;
  assign \new_[2496]_  = ~\new_[3292]_  & ~\new_[20052]_ ;
  assign \new_[2497]_  = \new_[3255]_  | \new_[2886]_ ;
  assign \new_[2498]_  = ~\new_[2886]_  | ~\new_[3255]_ ;
  assign \new_[2499]_  = \new_[2887]_  | \new_[20559]_ ;
  assign \new_[2500]_  = \\u0_w_reg[3][1] ;
  assign \new_[2501]_  = ~\new_[2843]_  | ~\new_[2847]_ ;
  assign \new_[2502]_  = ~\new_[3271]_  | ~\new_[3416]_ ;
  assign \new_[2503]_  = ~\new_[21646]_  | ~\new_[2846]_ ;
  assign \new_[2504]_  = ~\new_[2845]_  | ~\new_[3263]_ ;
  assign \new_[2505]_  = ~\new_[2843]_  | ~\new_[3407]_ ;
  assign \new_[2506]_  = ~\new_[3271]_  | ~\new_[3417]_ ;
  assign \new_[2507]_  = ~\new_[2883]_  | ~\new_[3433]_ ;
  assign \new_[2508]_  = ~\new_[20403]_  | ~\new_[20053]_ ;
  assign \new_[2509]_  = \\u0_w_reg[1][1] ;
  assign \text_out[20]  = \\text_out_reg[20] ;
  assign \new_[2511]_  = \\u0_w_reg[1][23] ;
  assign \new_[2512]_  = ~\new_[3405]_  | ~\new_[2858]_ ;
  assign \new_[2513]_  = ~\new_[2858]_  | ~\new_[3331]_ ;
  assign \new_[2514]_  = ~\new_[3296]_  | ~\new_[3536]_  | ~\new_[3113]_ ;
  assign \new_[2515]_  = ~\new_[2751]_ ;
  assign \new_[2516]_  = ~\new_[2805]_  | ~\new_[3350]_ ;
  assign \new_[2517]_  = ~\new_[3294]_  | ~\new_[3133]_  | ~\new_[3112]_ ;
  assign \new_[2518]_  = ~\new_[3907]_  | ~\new_[6190]_  | ~\new_[3115]_  | ~\new_[6363]_ ;
  assign \new_[2519]_  = ~\new_[3097]_  | ~\new_[2783]_ ;
  assign \new_[2520]_  = \\u0_w_reg[0][1] ;
  assign \new_[2521]_  = ~\new_[2842]_  | (~\new_[3639]_  & ~\new_[20417]_ );
  assign \new_[2522]_  = ~\new_[3011]_  | (~\new_[3394]_  & ~\new_[19749]_ );
  assign \new_[2523]_  = \new_[3335]_  ? \new_[3474]_  : \new_[3537]_ ;
  assign \new_[2524]_  = \new_[3537]_  ? \new_[3474]_  : \new_[3334]_ ;
  assign \new_[2525]_  = ~\new_[3014]_  | ~\new_[3013]_ ;
  assign n2373 = \new_[3304]_  ? \new_[19415]_  : \key[100] ;
  assign n2378 = \new_[3305]_  ? \new_[19371]_  : \key[68] ;
  assign n2383 = \new_[3307]_  ? \new_[19371]_  : \key[4] ;
  assign \new_[2529]_  = \new_[18513]_  ^ \new_[3306]_ ;
  assign n2388 = \new_[19070]_  ^ \new_[3297]_ ;
  assign \new_[2531]_  = ~\new_[2765]_ ;
  assign \new_[2532]_  = ~\new_[21537]_ ;
  assign \new_[2533]_  = ~\new_[3236]_  | ~\new_[3044]_ ;
  assign \new_[2534]_  = \new_[17810]_  ^ \new_[3308]_ ;
  assign \new_[2535]_  = \new_[8020]_  ^ \new_[3308]_ ;
  assign \new_[2536]_  = ~\new_[3067]_  | ~\new_[3072]_ ;
  assign \new_[2537]_  = \new_[20004]_  ? \new_[20882]_  : \new_[3655]_ ;
  assign n2473 = \new_[17475]_  ^ \new_[3309]_ ;
  assign \new_[2539]_  = ~\new_[3045]_  | (~\new_[3460]_  & ~\new_[3626]_ );
  assign \new_[2540]_  = ~\new_[3240]_  | (~\new_[3309]_  & ~\new_[18998]_ );
  assign \new_[2541]_  = ~\new_[3046]_  | ~\new_[3047]_ ;
  assign \new_[2542]_  = \new_[3046]_  & \new_[3047]_ ;
  assign \new_[2543]_  = ~\new_[3048]_  | (~\new_[3466]_  & ~\new_[20323]_ );
  assign \new_[2544]_  = \new_[3658]_  ? \new_[20882]_  : \new_[3657]_ ;
  assign \new_[2545]_  = ~\new_[2773]_ ;
  assign \new_[2546]_  = ~\new_[2774]_ ;
  assign \new_[2547]_  = ~\new_[3247]_  | (~\new_[3309]_  & ~\new_[18187]_ );
  assign \new_[2548]_  = ~\new_[3050]_  | ~\new_[1422]_ ;
  assign \new_[2549]_  = \new_[3311]_  ? \new_[3473]_  : \new_[20873]_ ;
  assign \new_[2550]_  = \new_[3505]_  ? \new_[19818]_  : \new_[3314]_ ;
  assign \new_[2551]_  = ~\new_[3050]_  | ~\new_[1351]_ ;
  assign \new_[2552]_  = ~\new_[3058]_  | ~\new_[3258]_ ;
  assign \new_[2553]_  = ~\new_[2780]_ ;
  assign \new_[2554]_  = ~\new_[3050]_  | ~\new_[1352]_ ;
  assign \new_[2555]_  = ~\new_[3043]_  | ~\new_[3235]_ ;
  assign \new_[2556]_  = ~\new_[2781]_ ;
  assign \text_out[86]  = \\text_out_reg[86] ;
  assign \new_[2558]_  = \new_[1513]_  ^ \new_[3479]_ ;
  assign \new_[2559]_  = \new_[1515]_  ^ \new_[3301]_ ;
  assign \new_[2560]_  = \new_[18221]_  ^ \new_[3479]_ ;
  assign \new_[2561]_  = \new_[17508]_  ^ \new_[3301]_ ;
  assign \new_[2562]_  = ~\new_[2792]_ ;
  assign \new_[2563]_  = \new_[14965]_  ^ \new_[3479]_ ;
  assign \new_[2564]_  = \new_[14963]_  ^ \new_[3301]_ ;
  assign n2308 = \new_[14690]_  ^ \new_[3303]_ ;
  assign \new_[2566]_  = \new_[3284]_  ? \new_[20655]_  : \new_[3285]_ ;
  assign \new_[2567]_  = ~\new_[3033]_  | ~\new_[3229]_ ;
  assign n2398 = \new_[19684]_  ^ \new_[3302]_ ;
  assign \new_[2569]_  = \new_[19667]_  ? \new_[3285]_  : \new_[1241]_ ;
  assign \new_[2570]_  = ~\new_[3034]_  | (~\new_[3488]_  & ~\new_[19634]_ );
  assign \new_[2571]_  = ~\new_[3035]_  | ~\new_[3230]_ ;
  assign \new_[2572]_  = ~\new_[3036]_  | (~\new_[3488]_  & ~\new_[19646]_ );
  assign \new_[2573]_  = ~\new_[3037]_  | ~\new_[3231]_ ;
  assign \new_[2574]_  = ~\new_[3038]_  | (~\new_[3488]_  & ~\new_[19705]_ );
  assign n2393 = \new_[18025]_  ^ \new_[3289]_ ;
  assign n2323 = \new_[1739]_  ^ \new_[3575]_ ;
  assign \new_[2577]_  = ~\new_[2809]_ ;
  assign \new_[2578]_  = \new_[3467]_  ? \new_[3320]_  : \new_[3587]_ ;
  assign \new_[2579]_  = \new_[3290]_  ? \new_[19998]_  : \new_[3461]_ ;
  assign \new_[2580]_  = ~\new_[3039]_  & (~\new_[3465]_  | ~\new_[3454]_ );
  assign \new_[2581]_  = ~\new_[3040]_  & (~\new_[3459]_  | ~\new_[21599]_ );
  assign \new_[2582]_  = ~\new_[3108]_  | ~\new_[3630]_ ;
  assign \new_[2583]_  = ~\new_[3092]_  | ~\new_[19544]_ ;
  assign \new_[2584]_  = ~\new_[3634]_  & ~\new_[19993]_ ;
  assign \new_[2585]_  = ~\new_[3116]_  | ~\new_[3509]_ ;
  assign \new_[2586]_  = ~\new_[3108]_  | ~\new_[3623]_ ;
  assign \new_[2587]_  = ~\new_[21276]_  & ~\new_[19993]_ ;
  assign n2463 = \new_[1659]_  ^ \new_[3298]_ ;
  assign \new_[2589]_  = ~\new_[2840]_ ;
  assign \new_[2590]_  = ~\new_[3077]_  | (~\new_[3475]_  & ~\new_[19588]_ );
  assign \new_[2591]_  = ~\new_[3117]_  | ~\new_[3538]_ ;
  assign \new_[2592]_  = ~\new_[3118]_  | ~\new_[3638]_ ;
  assign \new_[2593]_  = ~\new_[20888]_  | ~\new_[3636]_ ;
  assign \new_[2594]_  = ~\new_[3085]_  | (~\new_[3475]_  & ~\new_[19700]_ );
  assign \new_[2595]_  = ~\new_[3088]_  | ~\new_[3089]_ ;
  assign \new_[2596]_  = ~\new_[2847]_ ;
  assign \new_[2597]_  = ~\new_[2850]_ ;
  assign n2328 = \new_[19737]_  ^ \new_[3589]_ ;
  assign \new_[2599]_  = ~\new_[3078]_  | ~\new_[3081]_ ;
  assign \new_[2600]_  = ~\new_[3271]_ ;
  assign \new_[2601]_  = ~\new_[2854]_ ;
  assign n2348 = \new_[1658]_  ^ \new_[3610]_ ;
  assign \new_[2603]_  = ~\new_[2856]_ ;
  assign \new_[2604]_  = ~\new_[2857]_ ;
  assign \new_[2605]_  = ~\new_[3112]_  | ~\new_[3294]_ ;
  assign \new_[2606]_  = ~\new_[2858]_ ;
  assign \new_[2607]_  = ~\new_[3113]_  | ~\new_[3296]_ ;
  assign n2418 = \new_[2297]_  ^ \new_[3624]_ ;
  assign n2433 = \new_[17553]_  ^ \new_[3622]_ ;
  assign n2403 = \new_[1660]_  ^ \new_[3319]_ ;
  assign \new_[2611]_  = ~\new_[3109]_  | ~\new_[3110]_ ;
  assign n2413 = \new_[19101]_  ^ \new_[3314]_ ;
  assign n2428 = \new_[19560]_  ^ \new_[3325]_ ;
  assign n2438 = \new_[18772]_  ^ \new_[3316]_ ;
  assign n2423 = \new_[17482]_  ^ \new_[3321]_ ;
  assign n2408 = \new_[1427]_  ^ \new_[3320]_ ;
  assign \new_[2617]_  = ~\new_[3104]_  | ~\new_[3107]_ ;
  assign \new_[2618]_  = ~\new_[3105]_  | ~\new_[3106]_ ;
  assign \new_[2619]_  = ~\new_[21003]_  | ~\new_[21187]_ ;
  assign \text_out[81]  = \\text_out_reg[81] ;
  assign \new_[2621]_  = ~\new_[2878]_ ;
  assign \new_[2622]_  = ~\new_[2883]_ ;
  assign \new_[2623]_  = ~\new_[20417]_ ;
  assign \new_[2624]_  = ~\new_[2885]_ ;
  assign \new_[2625]_  = ~\new_[2886]_ ;
  assign \new_[2626]_  = ~\new_[2887]_ ;
  assign \new_[2627]_  = \new_[3541]_  ? \new_[3632]_  : \new_[3644]_ ;
  assign \new_[2628]_  = ~\new_[3134]_  | ~\new_[3135]_ ;
  assign n2448 = \new_[2300]_  ^ \new_[3330]_ ;
  assign \new_[2630]_  = ~\new_[3136]_  | (~\new_[3346]_  & ~\new_[17484]_ );
  assign \text_out[99]  = \\text_out_reg[99] ;
  assign \new_[2632]_  = ~\new_[3137]_  | (~\new_[3346]_  & ~\new_[19123]_ );
  assign \new_[2633]_  = ~\new_[3138]_  | (~\new_[19882]_  & ~\new_[19603]_ );
  assign \new_[2634]_  = ~\new_[2898]_ ;
  assign n2478 = \new_[19166]_  ^ \new_[3647]_ ;
  assign n2443 = \new_[19306]_  ^ \new_[3645]_ ;
  assign \new_[2637]_  = ~\new_[3163]_  | ~\new_[3213]_ ;
  assign \new_[2638]_  = \new_[3593]_  ? \new_[3214]_  : \new_[3661]_ ;
  assign \new_[2639]_  = \new_[6249]_  ^ \new_[3223]_ ;
  assign \new_[2640]_  = \new_[18135]_  ^ \new_[3218]_ ;
  assign \new_[2641]_  = \new_[6251]_  ? \new_[3374]_  : \new_[6995]_ ;
  assign \new_[2642]_  = \new_[6995]_  ^ \new_[3374]_ ;
  assign \new_[2643]_  = \new_[4984]_  ^ \new_[3373]_ ;
  assign \new_[2644]_  = \new_[8022]_  ^ \new_[3218]_ ;
  assign \new_[2645]_  = ~\new_[3164]_  | (~\new_[20667]_  & ~\new_[18179]_ );
  assign \new_[2646]_  = ~\new_[3144]_  | (~\new_[20061]_  & ~\new_[19716]_ );
  assign \new_[2647]_  = ~\new_[3145]_  | ~\new_[3146]_ ;
  assign \new_[2648]_  = ~\new_[3139]_  | (~\new_[20474]_  & ~\new_[1667]_ );
  assign \new_[2649]_  = ~\new_[3140]_  | ~\new_[3141]_ ;
  assign n2338 = \new_[1868]_  ^ \new_[3341]_ ;
  assign \new_[2651]_  = ~\new_[3143]_  | ~\new_[3142]_ ;
  assign \new_[2652]_  = \new_[1341]_  ^ \new_[3374]_ ;
  assign \new_[2653]_  = \new_[1289]_  ^ \new_[3374]_ ;
  assign \new_[2654]_  = \new_[19558]_  ? \new_[3375]_  : \new_[1474]_ ;
  assign \new_[2655]_  = ~\new_[3158]_  | ~\new_[3177]_ ;
  assign n2333 = \new_[2079]_  ^ \new_[3345]_ ;
  assign \new_[2657]_  = ~\new_[3147]_  | ~\new_[3148]_ ;
  assign \new_[2658]_  = ~\new_[3149]_  | (~\new_[3544]_  & ~\new_[19733]_ );
  assign \new_[2659]_  = \new_[3634]_  ? \new_[3372]_  : \new_[21376]_ ;
  assign \new_[2660]_  = ~\new_[3150]_  | ~\new_[3151]_ ;
  assign \new_[2661]_  = \new_[3250]_  ? \new_[3372]_  : \new_[3399]_ ;
  assign \new_[2662]_  = \new_[3692]_  ? \new_[21198]_  : \new_[3691]_ ;
  assign \new_[2663]_  = \new_[20258]_  ? \new_[21198]_  : \new_[3572]_ ;
  assign \new_[2664]_  = \new_[3667]_  ? \new_[3214]_  : \new_[3605]_ ;
  assign \new_[2665]_  = ~\new_[20061]_  | ~\new_[19775]_ ;
  assign \new_[2666]_  = ~\new_[20061]_  | ~\new_[19799]_ ;
  assign \new_[2667]_  = ~\new_[2996]_  | ~\new_[3228]_ ;
  assign \new_[2668]_  = ~\new_[3021]_  | ~\new_[3332]_ ;
  assign \new_[2669]_  = ~\new_[3165]_  | ~\new_[1420]_ ;
  assign \new_[2670]_  = ~\new_[3165]_  | ~\new_[19708]_ ;
  assign \new_[2671]_  = ~\new_[3165]_  | ~\new_[1671]_ ;
  assign \new_[2672]_  = ~\new_[3516]_  | ~\new_[3004]_ ;
  assign \new_[2673]_  = ~\new_[3123]_  | ~\new_[3007]_ ;
  assign \new_[2674]_  = ~\new_[21710]_  | ~\new_[1243]_ ;
  assign \new_[2675]_  = ~\new_[3002]_  | ~\new_[13690]_ ;
  assign \new_[2676]_  = ~\new_[3082]_  | ~\new_[2993]_ ;
  assign \new_[2677]_  = ~\new_[21710]_  | ~\new_[19397]_ ;
  assign \new_[2678]_  = ~\new_[21710]_  | ~\new_[1675]_ ;
  assign \new_[2679]_  = \new_[19630]_  ? \new_[3354]_  : \new_[1431]_ ;
  assign \new_[2680]_  = ~\new_[3196]_  | ~\new_[3195]_ ;
  assign \new_[2681]_  = \new_[3353]_  ? \new_[21617]_  : \new_[3354]_ ;
  assign \new_[2682]_  = ~\new_[2926]_ ;
  assign \new_[2683]_  = ~\new_[2927]_ ;
  assign \new_[2684]_  = ~\new_[3200]_  | ~\new_[3368]_ ;
  assign \new_[2685]_  = ~\new_[3199]_  | (~\new_[19901]_  & ~\new_[3315]_ );
  assign \new_[2686]_  = ~\new_[3180]_  | ~\new_[1239]_ ;
  assign \new_[2687]_  = ~\new_[2937]_ ;
  assign \new_[2688]_  = ~\new_[2939]_ ;
  assign \new_[2689]_  = ~\new_[2941]_ ;
  assign \new_[2690]_  = ~\new_[3192]_  | ~\new_[3194]_ ;
  assign n2453 = \new_[2294]_  ^ \new_[3355]_ ;
  assign \new_[2692]_  = \new_[18040]_  ^ \new_[3264]_ ;
  assign \new_[2693]_  = \new_[1507]_  ^ \new_[3264]_ ;
  assign \new_[2694]_  = ~\new_[3172]_  | (~\new_[3557]_  & ~\new_[1619]_ );
  assign \new_[2695]_  = \new_[1506]_  ^ \new_[3264]_ ;
  assign \new_[2696]_  = \new_[5283]_  ^ \new_[3264]_ ;
  assign \new_[2697]_  = ~\new_[3176]_  | (~\new_[3557]_  & ~\new_[19761]_ );
  assign n2458 = \new_[18011]_  ^ \new_[3272]_ ;
  assign \new_[2699]_  = ~\new_[3178]_  | ~\new_[3179]_ ;
  assign n2343 = \new_[19590]_  ^ \new_[3653]_ ;
  assign \new_[2701]_  = ~\new_[3173]_  | ~\new_[3174]_ ;
  assign \new_[2702]_  = ~\new_[3190]_  | ~\new_[3191]_ ;
  assign \new_[2703]_  = ~\new_[2948]_ ;
  assign \new_[2704]_  = \new_[3631]_  ? \new_[20655]_  : \new_[3530]_ ;
  assign \new_[2705]_  = \new_[3531]_  ? \new_[21332]_  : \new_[3632]_ ;
  assign \new_[2706]_  = ~\new_[2951]_ ;
  assign \new_[2707]_  = \new_[3459]_  ? \new_[20655]_  : \new_[3460]_ ;
  assign \new_[2708]_  = ~\new_[3187]_  | (~\new_[19969]_  & ~\new_[3595]_ );
  assign n2468 = \new_[19408]_  ^ \new_[3273]_ ;
  assign n2363 = \new_[1352]_  ^ \new_[21619]_ ;
  assign n2353 = \new_[1240]_  ^ \new_[3259]_ ;
  assign \new_[2712]_  = ~\new_[3198]_  | ~\new_[3201]_ ;
  assign \new_[2713]_  = ~\new_[3071]_  | ~\new_[3558]_ ;
  assign n2368 = \new_[1671]_  ^ \new_[20559]_ ;
  assign n2358 = \new_[19628]_  ^ \new_[3270]_ ;
  assign \new_[2716]_  = ~\new_[3202]_  | ~\new_[3206]_ ;
  assign \new_[2717]_  = ~\new_[3184]_  | ~\new_[3357]_ ;
  assign \new_[2718]_  = ~\new_[3209]_  | ~\new_[3208]_ ;
  assign \new_[2719]_  = ~\new_[3186]_  | ~\new_[3358]_ ;
  assign \new_[2720]_  = ~\new_[3212]_  | ~\new_[3211]_ ;
  assign n2303 = \new_[2500]_  ^ \new_[21487]_ ;
  assign \new_[2722]_  = \new_[3277]_  ? \new_[3300]_  : \new_[21176]_ ;
  assign \new_[2723]_  = ~\new_[3359]_  | ~\new_[3188]_ ;
  assign \new_[2724]_  = ~\new_[2959]_ ;
  assign n2298 = \new_[1433]_  ^ \new_[3570]_ ;
  assign \new_[2726]_  = ~\new_[3181]_  | (~\new_[3409]_  & ~\new_[3465]_ );
  assign \new_[2727]_  = ~\new_[3182]_  | (~\new_[3570]_  & ~\new_[3459]_ );
  assign \new_[2728]_  = \new_[3525]_  ? \new_[3249]_  : \new_[3324]_ ;
  assign \new_[2729]_  = ~\new_[19978]_  | ~\new_[3276]_ ;
  assign \new_[2730]_  = ~\new_[20250]_  | ~\new_[3277]_ ;
  assign \new_[2731]_  = ~\new_[3055]_  | ~\new_[3279]_ ;
  assign \new_[2732]_  = ~\new_[3056]_  | ~\new_[20131]_ ;
  assign \new_[2733]_  = ~\new_[21487]_  | ~\new_[3131]_ ;
  assign \new_[2734]_  = ~\new_[3075]_  | ~\new_[21240]_ ;
  assign \new_[2735]_  = ~\new_[3203]_  | (~\new_[19853]_  & ~\new_[19760]_ );
  assign \new_[2736]_  = ~\new_[3193]_  | ~\new_[3197]_ ;
  assign n2313 = \new_[1428]_  ^ \new_[3225]_ ;
  assign \new_[2738]_  = ~\new_[3068]_  | ~\new_[3269]_ ;
  assign \new_[2739]_  = ~\new_[3267]_  | ~\new_[3071]_ ;
  assign \new_[2740]_  = ~\new_[3108]_  | ~\new_[3408]_ ;
  assign \new_[2741]_  = ~\new_[3458]_  | ~\new_[20270]_ ;
  assign \new_[2742]_  = ~\new_[3061]_  | ~\new_[3412]_ ;
  assign \new_[2743]_  = ~\new_[3069]_  | ~\new_[3415]_ ;
  assign \new_[2744]_  = ~\new_[3060]_  | ~\new_[20854]_ ;
  assign \new_[2745]_  = ~\new_[21121]_  | ~\new_[3626]_ ;
  assign \new_[2746]_  = ~\new_[20646]_  | ~\new_[3509]_ ;
  assign \new_[2747]_  = ~\new_[3431]_  | ~\new_[19993]_ ;
  assign \new_[2748]_  = ~\new_[3470]_  | ~\new_[3132]_  | ~\new_[3295]_ ;
  assign \new_[2749]_  = ~\new_[2981]_ ;
  assign \new_[2750]_  = ~\new_[2983]_ ;
  assign \new_[2751]_  = ~\new_[2984]_ ;
  assign \new_[2752]_  = ~\new_[3030]_  | ~\new_[3175]_ ;
  assign n2318 = \new_[1509]_  ^ \new_[3243]_ ;
  assign \new_[2754]_  = ~\new_[2990]_ ;
  assign \new_[2755]_  = ~\new_[3010]_  | ~\new_[3009]_ ;
  assign n2558 = \key[116]  ? \new_[19614]_  : \new_[3492]_ ;
  assign n2563 = \key[84]  ? \new_[19614]_  : \new_[3497]_ ;
  assign n2568 = \key[20]  ? \new_[19614]_  : \new_[3495]_ ;
  assign \new_[2759]_  = ~\new_[3244]_  | (~\new_[3591]_  & ~\new_[19766]_ );
  assign \new_[2760]_  = ~\new_[2992]_ ;
  assign \new_[2761]_  = ~\new_[2994]_ ;
  assign \new_[2762]_  = ~\new_[2995]_ ;
  assign \new_[2763]_  = \new_[18207]_  ^ \new_[3494]_ ;
  assign \new_[2764]_  = ~\new_[3001]_ ;
  assign \new_[2765]_  = ~\new_[3254]_  | (~\new_[3594]_  & ~\new_[21276]_ );
  assign \new_[2766]_  = \new_[6223]_  ^ \new_[3493]_ ;
  assign \new_[2767]_  = ~\new_[3002]_ ;
  assign \new_[2768]_  = ~\new_[3002]_ ;
  assign \new_[2769]_  = \new_[4974]_  ^ \new_[3496]_ ;
  assign \new_[2770]_  = ~\new_[3004]_ ;
  assign \new_[2771]_  = ~\new_[3239]_  | ~\new_[3237]_ ;
  assign \new_[2772]_  = \new_[3239]_  & \new_[3237]_ ;
  assign \new_[2773]_  = (~\new_[20323]_  | ~\new_[3453]_ ) & (~\new_[20329]_  | ~\new_[21676]_ );
  assign \new_[2774]_  = (~\new_[3626]_  | ~\new_[21599]_ ) & (~\new_[3674]_  | ~\new_[21426]_ );
  assign \new_[2775]_  = ~\new_[3007]_ ;
  assign n2588 = \new_[1872]_  ^ \new_[3474]_ ;
  assign \new_[2777]_  = ~\new_[3253]_  | (~\new_[20342]_  & ~\new_[19547]_ );
  assign \new_[2778]_  = \new_[3614]_  ? \new_[3662]_  : \new_[3500]_ ;
  assign \new_[2779]_  = \new_[3620]_  ? \new_[3664]_  : \new_[3511]_ ;
  assign \new_[2780]_  = ~\new_[3233]_  | ~\new_[3234]_ ;
  assign \new_[2781]_  = (~\new_[3489]_  & ~\new_[19765]_ ) | (~\new_[3606]_  & ~\new_[19340]_ );
  assign \text_out[87]  = \\text_out_reg[87] ;
  assign \new_[2783]_  = ~\new_[3276]_  | ~\new_[20578]_ ;
  assign \text_out[17]  = \\text_out_reg[17] ;
  assign \new_[2785]_  = ~\new_[3012]_ ;
  assign n2573 = \new_[19187]_  ^ \new_[3485]_ ;
  assign \new_[2787]_  = \new_[1663]_  ^ \new_[3469]_ ;
  assign \new_[2788]_  = ~\new_[3017]_ ;
  assign \new_[2789]_  = \new_[18463]_  ^ \new_[3469]_ ;
  assign \new_[2790]_  = \new_[1670]_  ^ \new_[3469]_ ;
  assign \new_[2791]_  = \new_[19708]_  ^ \new_[3482]_ ;
  assign \new_[2792]_  = ~\new_[3238]_  | ~\new_[3393]_ ;
  assign \new_[2793]_  = \new_[5287]_  ^ \new_[3469]_ ;
  assign \new_[2794]_  = \new_[19686]_  ? \new_[3479]_  : \new_[1516]_ ;
  assign \new_[2795]_  = ~\new_[3395]_  | ~\new_[3245]_ ;
  assign n2583 = \new_[1513]_  ^ \new_[3471]_ ;
  assign \new_[2797]_  = \new_[18970]_  ^ \new_[3481]_ ;
  assign \new_[2798]_  = ~\new_[3398]_  | ~\new_[3252]_ ;
  assign \new_[2799]_  = \new_[1342]_  ^ \new_[3484]_ ;
  assign \new_[2800]_  = \new_[1668]_  ^ \new_[3481]_ ;
  assign \new_[2801]_  = ~\new_[3411]_  | ~\new_[3260]_ ;
  assign \new_[2802]_  = \new_[19121]_  ^ \new_[3484]_ ;
  assign \new_[2803]_  = \new_[9253]_  ^ \new_[3481]_ ;
  assign \new_[2804]_  = \new_[18109]_  ^ \new_[3481]_ ;
  assign \new_[2805]_  = ~\new_[3030]_ ;
  assign n2593 = \new_[1419]_  ^ \new_[3463]_ ;
  assign n2578 = \new_[1424]_  ^ \new_[3468]_ ;
  assign n2623 = \new_[19698]_  ^ \new_[3457]_ ;
  assign \new_[2809]_  = ~\new_[3232]_  | (~\new_[3575]_  & ~\new_[19704]_ );
  assign \new_[2810]_  = \new_[1664]_  ^ \new_[3491]_ ;
  assign \new_[2811]_  = \new_[1665]_  ^ \new_[21154]_ ;
  assign \new_[2812]_  = \new_[1666]_  ^ \new_[3478]_ ;
  assign \new_[2813]_  = \new_[17524]_  ^ \new_[3491]_ ;
  assign \new_[2814]_  = ~\new_[3032]_ ;
  assign \new_[2815]_  = \new_[18419]_  ^ \new_[21154]_ ;
  assign \new_[2816]_  = \new_[17704]_  ^ \new_[3478]_ ;
  assign \new_[2817]_  = \new_[1669]_  ^ \new_[21154]_ ;
  assign \new_[2818]_  = \new_[1671]_  ^ \new_[3478]_ ;
  assign \new_[2819]_  = \new_[8024]_  ^ \new_[3491]_ ;
  assign \new_[2820]_  = \new_[10504]_  ^ \new_[21154]_ ;
  assign \new_[2821]_  = \new_[14967]_  ^ \new_[3478]_ ;
  assign \new_[2822]_  = \new_[3584]_  ? \new_[3522]_  : \new_[3585]_ ;
  assign \new_[2823]_  = \new_[3456]_  ? \new_[3629]_  : \new_[3583]_ ;
  assign \new_[2824]_  = ~\new_[3292]_  & ~\new_[3455]_ ;
  assign \new_[2825]_  = ~\new_[3575]_  | ~\new_[21597]_ ;
  assign \new_[2826]_  = ~\new_[3666]_  | ~\new_[20828]_ ;
  assign \new_[2827]_  = ~\new_[3487]_  | ~\new_[3292]_ ;
  assign \new_[2828]_  = ~\new_[3292]_  | ~\new_[3678]_ ;
  assign \new_[2829]_  = ~\new_[3584]_  | ~\new_[3312]_ ;
  assign \new_[2830]_  = ~\new_[3299]_  | ~\new_[19626]_ ;
  assign \new_[2831]_  = ~\new_[3284]_  | ~\new_[1240]_ ;
  assign \new_[2832]_  = ~\new_[3300]_  | ~\new_[19720]_ ;
  assign \new_[2833]_  = ~\new_[3299]_  | ~\new_[19793]_ ;
  assign \new_[2834]_  = ~\new_[3589]_  & ~\new_[3285]_ ;
  assign \new_[2835]_  = ~\new_[3050]_ ;
  assign \new_[2836]_  = ~\new_[3520]_  | ~\new_[20828]_ ;
  assign \new_[2837]_  = ~\new_[3051]_ ;
  assign \new_[2838]_  = ~\new_[3518]_  | ~\new_[3287]_ ;
  assign \new_[2839]_  = ~\new_[3621]_  | ~\new_[3455]_ ;
  assign \new_[2840]_  = ~\new_[20250]_ ;
  assign \new_[2841]_  = ~\new_[3057]_ ;
  assign \new_[2842]_  = ~\new_[20417]_  | ~\new_[3640]_ ;
  assign \new_[2843]_  = ~\new_[3060]_ ;
  assign \new_[2844]_  = \new_[3589]_  ? \new_[1347]_  : \new_[3659]_ ;
  assign \new_[2845]_  = ~\new_[3061]_ ;
  assign \new_[2846]_  = ~\new_[20270]_ ;
  assign \new_[2847]_  = ~\new_[20270]_ ;
  assign \new_[2848]_  = ~\new_[3062]_ ;
  assign \new_[2849]_  = ~\new_[3063]_ ;
  assign \new_[2850]_  = ~\new_[3423]_  | ~\new_[3280]_ ;
  assign \new_[2851]_  = ~\new_[3066]_ ;
  assign \new_[2852]_  = ~\new_[3430]_  | ~\new_[3282]_ ;
  assign \new_[2853]_  = ~\new_[3432]_  | ~\new_[3283]_ ;
  assign \new_[2854]_  = \new_[3624]_  ? \new_[3517]_  : \new_[20053]_ ;
  assign \new_[2855]_  = ~\new_[3076]_ ;
  assign \new_[2856]_  = \new_[3701]_  ? \new_[3503]_  : \new_[20329]_ ;
  assign \new_[2857]_  = \new_[3506]_  ? \new_[21586]_  : \new_[3507]_ ;
  assign \new_[2858]_  = ~\new_[3295]_  | ~\new_[3470]_ ;
  assign \new_[2859]_  = ~\new_[3298]_  | ~\new_[19714]_ ;
  assign n2498 = \new_[1637]_  ^ \new_[20872]_ ;
  assign n2603 = \new_[19532]_  ^ \new_[3510]_ ;
  assign n2493 = \new_[1620]_  ^ \new_[3499]_ ;
  assign \new_[2863]_  = ~\new_[3082]_ ;
  assign \new_[2864]_  = \new_[3630]_  ? \new_[1513]_  : \new_[3526]_ ;
  assign \new_[2865]_  = ~\new_[3084]_ ;
  assign \new_[2866]_  = ~\new_[3086]_ ;
  assign \new_[2867]_  = ~\new_[3087]_ ;
  assign \new_[2868]_  = \new_[19998]_  ? \new_[3525]_  : \new_[3523]_ ;
  assign \new_[2869]_  = \new_[3523]_  ? \new_[3525]_  : \new_[19998]_ ;
  assign \new_[2870]_  = ~\new_[21240]_ ;
  assign \new_[2871]_  = ~\new_[21240]_ ;
  assign \new_[2872]_  = \new_[20223]_  ? \new_[20054]_  : \new_[3628]_ ;
  assign n2598 = \new_[18961]_  ^ \new_[3522]_ ;
  assign n2608 = \new_[19591]_  ^ \new_[21624]_ ;
  assign \new_[2875]_  = ~\new_[3102]_ ;
  assign \new_[2876]_  = ~\new_[3320]_  | ~\new_[3313]_ ;
  assign \new_[2877]_  = ~\new_[3628]_  | ~\new_[20077]_ ;
  assign \new_[2878]_  = ~\new_[3108]_ ;
  assign \text_out[49]  = \\text_out_reg[49] ;
  assign \new_[2880]_  = ~\new_[3328]_  | ~\new_[3506]_ ;
  assign \new_[2881]_  = ~\new_[3329]_  | ~\new_[3706]_ ;
  assign \new_[2882]_  = ~\new_[3311]_  | ~\new_[3518]_ ;
  assign \new_[2883]_  = ~\new_[19993]_ ;
  assign \new_[2884]_  = ~\new_[3114]_ ;
  assign \new_[2885]_  = ~\new_[3117]_ ;
  assign \new_[2886]_  = ~\new_[20888]_ ;
  assign \new_[2887]_  = ~\new_[3118]_ ;
  assign n2483 = \new_[15893]_  ^ \new_[3536]_ ;
  assign \new_[2889]_  = ~\new_[3119]_ ;
  assign \new_[2890]_  = \new_[3644]_  ? \new_[3632]_  : \new_[3541]_ ;
  assign \new_[2891]_  = ~\new_[3120]_ ;
  assign n2648 = \new_[19373]_  ^ \new_[3533]_ ;
  assign n2613 = \new_[1661]_  ^ \new_[3530]_ ;
  assign n2618 = \new_[2301]_  ^ \new_[3532]_ ;
  assign \text_out[8]  = \\text_out_reg[8] ;
  assign \new_[2896]_  = ~\new_[3125]_ ;
  assign \new_[2897]_  = ~\new_[3127]_ ;
  assign \new_[2898]_  = ~\new_[3128]_ ;
  assign \new_[2899]_  = ~\new_[20623]_  | ~\new_[18877]_ ;
  assign \new_[2900]_  = ~\new_[3348]_  | ~\new_[18449]_ ;
  assign \new_[2901]_  = ~\new_[3348]_  | ~\new_[18391]_ ;
  assign \new_[2902]_  = ~\new_[3348]_  | ~\new_[3706]_ ;
  assign n2628 = \key[103]  ? \new_[19614]_  : \new_[3376]_ ;
  assign n2518 = \key[71]  ? \new_[19614]_  : \new_[3377]_ ;
  assign n2488 = \key[7]  ? \new_[19649]_  : \new_[3379]_ ;
  assign \new_[2906]_  = \new_[18354]_  ^ \new_[3378]_ ;
  assign n2633 = \key[114]  ? \new_[19614]_  : \new_[3381]_ ;
  assign n2523 = \key[98]  ? \new_[19614]_  : \new_[3382]_ ;
  assign n2508 = \key[82]  ? \new_[19649]_  : \new_[3388]_ ;
  assign n2528 = \key[66]  ? \new_[19614]_  : \new_[3383]_ ;
  assign n2533 = \key[18]  ? \new_[19614]_  : \new_[3386]_ ;
  assign n2538 = \key[2]  ? \new_[19614]_  : \new_[3387]_ ;
  assign \new_[2913]_  = ~\new_[3337]_  | (~\new_[3648]_  & ~\new_[1343]_ );
  assign \new_[2914]_  = ~\new_[3338]_  | (~\new_[3648]_  & ~\new_[19606]_ );
  assign \new_[2915]_  = ~\new_[3339]_  | (~\new_[3648]_  & ~\new_[19753]_ );
  assign \new_[2916]_  = ~\new_[3340]_  | ~\new_[19552]_ ;
  assign \new_[2917]_  = ~\new_[3340]_  | ~\new_[1346]_ ;
  assign \new_[2918]_  = \new_[17624]_  ^ \new_[3384]_ ;
  assign \new_[2919]_  = \new_[18388]_  ^ \new_[3380]_ ;
  assign \new_[2920]_  = ~\new_[3279]_  | ~\new_[3544]_ ;
  assign \new_[2921]_  = \new_[3660]_  ? \new_[21332]_  : \new_[21530]_ ;
  assign n2543 = \key[119]  ? \new_[19614]_  : \new_[3425]_ ;
  assign n2653 = \key[87]  ? \new_[19614]_  : \new_[3426]_ ;
  assign n2548 = \key[23]  ? \new_[19614]_  : \new_[3429]_ ;
  assign \new_[2925]_  = ~\new_[20131]_  | ~\new_[3216]_ ;
  assign \new_[2926]_  = ~\new_[3363]_  | ~\new_[3364]_ ;
  assign \new_[2927]_  = ~\new_[3365]_  | ~\new_[3366]_ ;
  assign n2513 = \new_[2509]_  ^ \new_[3690]_ ;
  assign \new_[2929]_  = ~\new_[3160]_ ;
  assign \new_[2930]_  = ~\new_[3163]_ ;
  assign \new_[2931]_  = ~\new_[3163]_ ;
  assign \new_[2932]_  = ~\new_[3217]_  | ~\new_[19166]_ ;
  assign \new_[2933]_  = \new_[18073]_  ^ \new_[3427]_ ;
  assign \new_[2934]_  = ~\new_[3690]_  | ~\new_[21676]_ ;
  assign \new_[2935]_  = ~\new_[3353]_  | ~\new_[19628]_ ;
  assign \new_[2936]_  = ~\new_[3653]_  & ~\new_[3354]_ ;
  assign \new_[2937]_  = \new_[20048]_  ? \new_[19840]_  : \new_[3623]_ ;
  assign \new_[2938]_  = ~\new_[3165]_ ;
  assign \new_[2939]_  = \new_[20329]_  ? \new_[20391]_  : \new_[3702]_ ;
  assign \new_[2940]_  = ~\new_[3217]_  | ~\new_[19419]_ ;
  assign \new_[2941]_  = ~\new_[3362]_  | ~\new_[3361]_ ;
  assign n2553 = \new_[1430]_  ^ \new_[19840]_ ;
  assign \new_[2943]_  = ~\new_[3549]_  | ~\new_[3349]_ ;
  assign \new_[2944]_  = ~\new_[3550]_  | ~\new_[3351]_ ;
  assign \new_[2945]_  = \new_[3653]_  ? \new_[19686]_  : \new_[3693]_ ;
  assign \new_[2946]_  = ~\new_[3169]_ ;
  assign \new_[2947]_  = ~\new_[3171]_ ;
  assign \new_[2948]_  = ~\new_[3555]_  | ~\new_[3352]_ ;
  assign \new_[2949]_  = ~\new_[3355]_  | ~\new_[19726]_ ;
  assign \new_[2950]_  = \new_[3633]_  ? \new_[21617]_  : \new_[3532]_ ;
  assign \new_[2951]_  = \new_[3465]_  ? \new_[21618]_  : \new_[3466]_ ;
  assign \new_[2952]_  = ~\new_[3177]_ ;
  assign n2503 = \new_[18773]_  ^ \new_[3433]_ ;
  assign \new_[2954]_  = ~\new_[3269]_  | ~\new_[3557]_ ;
  assign n2658 = \new_[3435]_  ? ld : \key[97] ;
  assign n2643 = \new_[3437]_  ? \new_[19415]_  : \key[65] ;
  assign \new_[2957]_  = ~\new_[3356]_  | ~\new_[3559]_ ;
  assign n2638 = \new_[3439]_  ? \new_[19415]_  : \key[1] ;
  assign \new_[2959]_  = ~\new_[3360]_  | (~\new_[21484]_  & ~\new_[19578]_ );
  assign \new_[2960]_  = \new_[18240]_  ^ \new_[3438]_ ;
  assign \new_[2961]_  = ~\new_[3246]_  | ~\new_[20523]_ ;
  assign \new_[2962]_  = ~\new_[3248]_  | ~\new_[20687]_ ;
  assign \new_[2963]_  = ~\new_[3249]_  | ~\new_[3400]_ ;
  assign \new_[2964]_  = ~\new_[3266]_  | ~\new_[3292]_ ;
  assign \new_[2965]_  = ~\new_[3265]_  | ~\new_[20352]_ ;
  assign \new_[2966]_  = ~\new_[3262]_  | ~\new_[19954]_ ;
  assign \new_[2967]_  = ~\new_[3464]_  & ~\new_[20559]_ ;
  assign \new_[2968]_  = ~\new_[3458]_  & ~\new_[3255]_ ;
  assign \new_[2969]_  = ~\new_[3367]_  | (~\new_[3562]_  & ~\new_[19569]_ );
  assign \new_[2970]_  = ~\new_[3369]_  | (~\new_[3562]_  & ~\new_[19781]_ );
  assign \new_[2971]_  = ~\new_[3293]_  | ~\new_[19840]_ ;
  assign \new_[2972]_  = ~\new_[3370]_  | (~\new_[3562]_  & ~\new_[19682]_ );
  assign \new_[2973]_  = ~\new_[20596]_  | ~\new_[3268]_ ;
  assign \new_[2974]_  = ~\new_[3267]_  | ~\new_[21027]_ ;
  assign \new_[2975]_  = ~\new_[3313]_  | ~\new_[19853]_ ;
  assign \new_[2976]_  = ~\new_[20559]_  | ~\new_[3701]_ ;
  assign \new_[2977]_  = ~\new_[3255]_  | ~\new_[3672]_ ;
  assign \new_[2978]_  = \new_[3313]_  | \new_[19853]_ ;
  assign \new_[2979]_  = ~\new_[3224]_  | ~\new_[1288]_ ;
  assign \new_[2980]_  = ~\new_[3224]_  | ~\new_[19605]_ ;
  assign \new_[2981]_  = ~\new_[21613]_ ;
  assign \new_[2982]_  = ~\new_[3205]_ ;
  assign \new_[2983]_  = ~\new_[3207]_ ;
  assign \new_[2984]_  = ~\new_[20445]_  | ~\new_[4201]_ ;
  assign \new_[2985]_  = \new_[3210]_ ;
  assign \new_[2986]_  = \new_[3534]_  ? \new_[3663]_  : \new_[3635]_ ;
  assign \new_[2987]_  = \new_[3635]_  ? \new_[3663]_  : \new_[3534]_ ;
  assign \new_[2988]_  = \new_[3535]_  ? \new_[19818]_  : \new_[3637]_ ;
  assign \new_[2989]_  = \new_[3637]_  ? \new_[19818]_  : \new_[3535]_ ;
  assign \new_[2990]_  = ~\new_[3213]_ ;
  assign n2673 = \new_[1507]_  ^ \new_[3591]_ ;
  assign \new_[2992]_  = ~\new_[3402]_  | (~\new_[21530]_  & ~\new_[19805]_ );
  assign \new_[2993]_  = ~\new_[3215]_ ;
  assign \new_[2994]_  = ~\new_[3403]_  | ~\new_[3404]_ ;
  assign \new_[2995]_  = ~\new_[20667]_ ;
  assign \new_[2996]_  = ~\new_[3332]_ ;
  assign \new_[2997]_  = \new_[1863]_  ^ \new_[3597]_ ;
  assign \new_[2998]_  = \new_[18342]_  ^ \new_[3597]_ ;
  assign \new_[2999]_  = \new_[1921]_  ^ \new_[3597]_ ;
  assign \new_[3000]_  = \new_[6170]_  ^ \new_[3597]_ ;
  assign \new_[3001]_  = ~\new_[3397]_  | ~\new_[3568]_ ;
  assign \new_[3002]_  = \new_[9673]_  ? \new_[3599]_  : \new_[10857]_ ;
  assign \new_[3003]_  = \new_[10731]_  ^ \new_[3592]_ ;
  assign \new_[3004]_  = ~\new_[3219]_ ;
  assign \new_[3005]_  = \new_[1419]_  ^ \new_[3592]_ ;
  assign \new_[3006]_  = \new_[19698]_  ^ \new_[3592]_ ;
  assign \new_[3007]_  = ~\new_[3220]_ ;
  assign n2668 = \new_[1875]_  ^ \new_[19817]_ ;
  assign \new_[3009]_  = ~\new_[3396]_  | ~\new_[1662]_ ;
  assign \new_[3010]_  = ~\new_[3394]_  | ~\new_[19633]_ ;
  assign \new_[3011]_  = ~\new_[3394]_  | ~\new_[19749]_ ;
  assign \new_[3012]_  = ~\new_[3389]_  | ~\new_[3565]_ ;
  assign \new_[3013]_  = ~\new_[3394]_  | ~\new_[19800]_ ;
  assign \new_[3014]_  = ~\new_[3396]_  | ~\new_[1417]_ ;
  assign \new_[3015]_  = \new_[1418]_  ? \new_[3599]_  : \new_[19784]_ ;
  assign \new_[3016]_  = ~\new_[3224]_ ;
  assign \new_[3017]_  = ~\new_[3391]_  | ~\new_[3567]_ ;
  assign \new_[3018]_  = ~\new_[3226]_ ;
  assign \new_[3019]_  = ~\new_[3227]_ ;
  assign \new_[3020]_  = \new_[1420]_  ? \new_[3599]_  : \new_[19774]_ ;
  assign \new_[3021]_  = ~\new_[3228]_ ;
  assign \new_[3022]_  = \new_[1868]_  ^ \new_[3602]_ ;
  assign \new_[3023]_  = \new_[18961]_  ^ \new_[3598]_ ;
  assign \new_[3024]_  = \new_[1866]_  ^ \new_[3602]_ ;
  assign \new_[3025]_  = \new_[18257]_  ^ \new_[3598]_ ;
  assign \new_[3026]_  = \new_[17899]_  ^ \new_[3602]_ ;
  assign \new_[3027]_  = \new_[1867]_  ^ \new_[3598]_ ;
  assign \new_[3028]_  = \new_[9258]_  ^ \new_[3598]_ ;
  assign \new_[3029]_  = \new_[12485]_  ^ \new_[3602]_ ;
  assign \new_[3030]_  = ~\new_[3390]_  | (~\new_[21699]_  & ~\new_[19783]_ );
  assign \new_[3031]_  = \new_[19387]_  ^ \new_[3609]_ ;
  assign \new_[3032]_  = ~\new_[3392]_  | (~\new_[21699]_  & ~\new_[19631]_ );
  assign \new_[3033]_  = ~\new_[3471]_  | ~\new_[19784]_ ;
  assign \new_[3034]_  = ~\new_[3486]_  | ~\new_[19634]_ ;
  assign \new_[3035]_  = ~\new_[3471]_  | ~\new_[19811]_ ;
  assign \new_[3036]_  = ~\new_[3486]_  | ~\new_[19646]_ ;
  assign \new_[3037]_  = ~\new_[3471]_  | ~\new_[19551]_ ;
  assign \new_[3038]_  = ~\new_[3486]_  | ~\new_[19705]_ ;
  assign \new_[3039]_  = ~\new_[3464]_  & ~\new_[3454]_ ;
  assign \new_[3040]_  = ~\new_[3458]_  & ~\new_[21599]_ ;
  assign \new_[3041]_  = ~\new_[3603]_  | ~\new_[3455]_ ;
  assign \new_[3042]_  = ~\new_[3585]_  | ~\new_[20873]_ ;
  assign \new_[3043]_  = ~\new_[20121]_  | ~\new_[3504]_ ;
  assign \new_[3044]_  = ~\new_[3462]_  | ~\new_[20629]_ ;
  assign \new_[3045]_  = ~\new_[3460]_  | ~\new_[3672]_ ;
  assign \new_[3046]_  = ~\new_[3506]_  | ~\new_[20546]_ ;
  assign \new_[3047]_  = ~\new_[3462]_  | ~\new_[20612]_ ;
  assign \new_[3048]_  = ~\new_[3466]_  | ~\new_[3701]_ ;
  assign \new_[3049]_  = ~\new_[3519]_  | ~\new_[3455]_ ;
  assign \new_[3050]_  = ~\new_[20882]_ ;
  assign \new_[3051]_  = ~\new_[20655]_ ;
  assign \new_[3052]_  = ~\new_[3241]_ ;
  assign \new_[3053]_  = ~\new_[3242]_ ;
  assign \new_[3054]_  = ~\new_[3246]_ ;
  assign \new_[3055]_  = ~\new_[3248]_ ;
  assign \new_[3056]_  = ~\new_[3249]_ ;
  assign \new_[3057]_  = ~\new_[3251]_ ;
  assign \new_[3058]_  = ~\new_[3667]_  | ~\new_[3498]_ ;
  assign \new_[3059]_  = ~\new_[3480]_  | ~\new_[3929]_ ;
  assign \new_[3060]_  = ~\new_[3256]_ ;
  assign \new_[3061]_  = ~\new_[3257]_ ;
  assign \new_[3062]_  = ~\new_[3419]_  | ~\new_[3420]_ ;
  assign \new_[3063]_  = ~\new_[3422]_  | ~\new_[3421]_ ;
  assign \new_[3064]_  = ~\new_[3483]_  | ~\new_[3756]_ ;
  assign \new_[3065]_  = ~\new_[3263]_ ;
  assign \new_[3066]_  = ~\new_[3266]_ ;
  assign \new_[3067]_  = ~\new_[21474]_  | ~\new_[3498]_ ;
  assign \new_[3068]_  = ~\new_[3267]_ ;
  assign \new_[3069]_  = ~\new_[3267]_ ;
  assign \new_[3070]_  = ~\new_[3424]_  | ~\new_[3428]_ ;
  assign \new_[3071]_  = ~\new_[3269]_ ;
  assign \new_[3072]_  = ~\new_[3416]_  | ~\new_[20342]_ ;
  assign \new_[3073]_  = ~\new_[3275]_ ;
  assign \new_[3074]_  = ~\new_[3277]_ ;
  assign \new_[3075]_  = ~\new_[3278]_ ;
  assign \new_[3076]_  = \new_[3672]_  ? \new_[3612]_  : \new_[3625]_ ;
  assign \new_[3077]_  = ~\new_[3475]_  | ~\new_[19588]_ ;
  assign \new_[3078]_  = ~\new_[3659]_  | ~\new_[3459]_ ;
  assign \new_[3079]_  = ~\new_[3441]_  | ~\new_[3442]_ ;
  assign \new_[3080]_  = ~\new_[3443]_  | ~\new_[3444]_ ;
  assign \new_[3081]_  = ~\new_[3588]_  | ~\new_[3460]_ ;
  assign \new_[3082]_  = ~\new_[3445]_  | ~\new_[3446]_ ;
  assign \new_[3083]_  = ~\new_[3447]_  | ~\new_[3448]_ ;
  assign \new_[3084]_  = ~\new_[3449]_  | ~\new_[3580]_ ;
  assign \new_[3085]_  = ~\new_[3475]_  | ~\new_[19700]_ ;
  assign \new_[3086]_  = ~\new_[3450]_  | ~\new_[3451]_ ;
  assign \new_[3087]_  = ~\new_[3452]_  | ~\new_[3581]_ ;
  assign \new_[3088]_  = ~\new_[3659]_  | ~\new_[3476]_ ;
  assign \new_[3089]_  = ~\new_[3588]_  | ~\new_[3475]_ ;
  assign \new_[3090]_  = \new_[1875]_  ^ \new_[3615]_ ;
  assign n2663 = \new_[1867]_  ^ \new_[3629]_ ;
  assign \new_[3092]_  = ~\new_[3284]_ ;
  assign \new_[3093]_  = \new_[1872]_  ^ \new_[3615]_ ;
  assign \new_[3094]_  = \new_[19043]_  ^ \new_[3618]_ ;
  assign \new_[3095]_  = \new_[17907]_  ^ \new_[3615]_ ;
  assign \new_[3096]_  = \new_[17897]_  ^ \new_[3618]_ ;
  assign \new_[3097]_  = ~\new_[20523]_  | ~\new_[20577]_ ;
  assign \new_[3098]_  = \new_[1877]_  ^ \new_[3618]_ ;
  assign \new_[3099]_  = \new_[11487]_  ^ \new_[3615]_ ;
  assign \new_[3100]_  = \new_[9254]_  ^ \new_[3618]_ ;
  assign \new_[3101]_  = ~\new_[3578]_  | ~\new_[3440]_ ;
  assign \new_[3102]_  = ~\new_[3579]_  | (~\new_[21625]_  & ~\new_[19810]_ );
  assign \new_[3103]_  = ~\new_[3522]_  | ~\new_[3515]_ ;
  assign \new_[3104]_  = ~\new_[3629]_  | ~\new_[3516]_ ;
  assign \new_[3105]_  = ~\new_[3512]_  | ~\new_[19998]_ ;
  assign \new_[3106]_  = ~\new_[3523]_  | ~\new_[19829]_ ;
  assign \new_[3107]_  = ~\new_[20119]_  | ~\new_[19943]_ ;
  assign \new_[3108]_  = ~\new_[3293]_ ;
  assign \new_[3109]_  = ~\new_[3507]_  | ~\new_[3706]_ ;
  assign \new_[3110]_  = ~\new_[3509]_  | ~\new_[21277]_ ;
  assign \new_[3111]_  = ~\new_[3621]_  | ~\new_[20873]_ ;
  assign \new_[3112]_  = ~\new_[3502]_  | ~\new_[3505]_ ;
  assign \new_[3113]_  = ~\new_[21586]_  | ~\new_[3620]_ ;
  assign \new_[3114]_  = ~\new_[3299]_ ;
  assign \new_[3115]_  = ~\new_[7356]_  & ~\new_[3529]_ ;
  assign \new_[3116]_  = \new_[20417]_ ;
  assign \new_[3117]_  = \new_[20735]_ ;
  assign \new_[3118]_  = \new_[20194]_ ;
  assign \new_[3119]_  = \new_[3686]_  ? \new_[19902]_  : \new_[3643]_ ;
  assign \new_[3120]_  = ~\new_[3310]_ ;
  assign \new_[3121]_  = ~\new_[3310]_ ;
  assign \new_[3122]_  = ~\new_[21370]_ ;
  assign \new_[3123]_  = ~\new_[3313]_ ;
  assign \new_[3124]_  = ~\new_[3315]_ ;
  assign \new_[3125]_  = ~\new_[3322]_ ;
  assign \new_[3126]_  = ~\new_[3323]_ ;
  assign \new_[3127]_  = ~\new_[3326]_ ;
  assign \new_[3128]_  = ~\new_[3327]_ ;
  assign \new_[3129]_  = ~\new_[3328]_ ;
  assign \new_[3130]_  = ~\new_[3329]_ ;
  assign \new_[3131]_  = ~\new_[3329]_ ;
  assign \new_[3132]_  = ~\new_[3331]_ ;
  assign \new_[3133]_  = ~\new_[3333]_ ;
  assign \new_[3134]_  = \new_[3512]_  | \new_[19882]_ ;
  assign \new_[3135]_  = ~\new_[3513]_  | ~\new_[19882]_ ;
  assign \new_[3136]_  = ~\new_[19882]_  | ~\new_[17484]_ ;
  assign \new_[3137]_  = ~\new_[19882]_  | ~\new_[19123]_ ;
  assign \new_[3138]_  = ~\new_[19882]_  | ~\new_[19603]_ ;
  assign \new_[3139]_  = ~\new_[20474]_  | ~\new_[1667]_ ;
  assign \new_[3140]_  = \new_[3516]_  | \new_[20474]_ ;
  assign \new_[3141]_  = ~\new_[3516]_  | ~\new_[20474]_ ;
  assign \new_[3142]_  = ~\new_[3542]_  | ~\new_[3466]_ ;
  assign \new_[3143]_  = ~\new_[3648]_  | ~\new_[3465]_ ;
  assign \new_[3144]_  = ~\new_[20061]_  | ~\new_[19716]_ ;
  assign \new_[3145]_  = \new_[3515]_  | \new_[20061]_ ;
  assign \new_[3146]_  = ~\new_[3514]_  | ~\new_[20061]_ ;
  assign \new_[3147]_  = ~\new_[3544]_  | ~\new_[1510]_ ;
  assign \new_[3148]_  = ~\new_[3545]_  | ~\new_[19306]_ ;
  assign \new_[3149]_  = ~\new_[3544]_  | ~\new_[19733]_ ;
  assign \new_[3150]_  = ~\new_[3544]_  | ~\new_[19732]_ ;
  assign \new_[3151]_  = ~\new_[3545]_  | ~\new_[1921]_ ;
  assign \new_[3152]_  = ~\new_[20687]_  | ~\new_[20173]_ ;
  assign \new_[3153]_  = ~\new_[3340]_ ;
  assign \new_[3154]_  = \new_[9330]_  ^ \new_[3576]_ ;
  assign \new_[3155]_  = \new_[17305]_  ^ \new_[3574]_ ;
  assign \new_[3156]_  = \new_[6245]_  ^ \new_[3577]_ ;
  assign \new_[3157]_  = \new_[8018]_  ^ \new_[3574]_ ;
  assign \new_[3158]_  = ~\new_[3342]_ ;
  assign \new_[3159]_  = ~\new_[3401]_  | ~\new_[20667]_ ;
  assign \new_[3160]_  = ~\new_[3543]_  | (~\new_[3690]_  & ~\new_[19796]_ );
  assign \new_[3161]_  = ~\new_[20667]_  | ~\new_[17578]_ ;
  assign \new_[3162]_  = ~\new_[3344]_ ;
  assign \new_[3163]_  = ~\new_[3561]_  | (~\new_[20413]_  & ~\new_[3706]_ );
  assign \new_[3164]_  = ~\new_[20667]_  | ~\new_[18179]_ ;
  assign \new_[3165]_  = ~\new_[21198]_ ;
  assign \new_[3166]_  = ~\new_[20667]_  | ~\new_[19098]_ ;
  assign \new_[3167]_  = ~\new_[3346]_ ;
  assign \new_[3168]_  = ~\new_[3547]_  | ~\new_[3548]_ ;
  assign \new_[3169]_  = ~\new_[3551]_  | ~\new_[3552]_ ;
  assign \new_[3170]_  = ~\new_[3347]_ ;
  assign \new_[3171]_  = ~\new_[3553]_  | ~\new_[3554]_ ;
  assign \new_[3172]_  = ~\new_[3557]_  | ~\new_[1619]_ ;
  assign \new_[3173]_  = ~\new_[3693]_  | ~\new_[3465]_ ;
  assign \new_[3174]_  = ~\new_[3652]_  | ~\new_[3466]_ ;
  assign \new_[3175]_  = ~\new_[3350]_ ;
  assign \new_[3176]_  = ~\new_[3557]_  | ~\new_[19761]_ ;
  assign \new_[3177]_  = ~\new_[3560]_  | (~\new_[20258]_  & ~\new_[19819]_ );
  assign \new_[3178]_  = ~\new_[3693]_  | ~\new_[3558]_ ;
  assign \new_[3179]_  = ~\new_[3652]_  | ~\new_[3557]_ ;
  assign \new_[3180]_  = ~\new_[3353]_ ;
  assign \new_[3181]_  = ~\new_[3410]_  | ~\new_[3464]_ ;
  assign \new_[3182]_  = ~\new_[3571]_  | ~\new_[3458]_ ;
  assign \new_[3183]_  = ~\new_[19969]_  | ~\new_[3590]_ ;
  assign \new_[3184]_  = ~\new_[21648]_  | ~\new_[3406]_ ;
  assign \new_[3185]_  = ~\new_[3585]_  | ~\new_[3412]_ ;
  assign \new_[3186]_  = ~\new_[20120]_  | ~\new_[3414]_ ;
  assign \new_[3187]_  = ~\new_[19969]_  | ~\new_[3595]_ ;
  assign \new_[3188]_  = ~\new_[21486]_  | ~\new_[19195]_ ;
  assign \new_[3189]_  = ~\new_[3464]_  | ~\new_[20391]_ ;
  assign \new_[3190]_  = ~\new_[19840]_  | ~\new_[21626]_ ;
  assign \new_[3191]_  = ~\new_[3408]_  | ~\new_[21627]_ ;
  assign \new_[3192]_  = \new_[3508]_  | \new_[21474]_ ;
  assign \new_[3193]_  = ~\new_[3562]_  | ~\new_[3459]_ ;
  assign \new_[3194]_  = ~\new_[3509]_  | ~\new_[21474]_ ;
  assign \new_[3195]_  = ~\new_[3621]_  | ~\new_[3412]_ ;
  assign \new_[3196]_  = \new_[3621]_  | \new_[3412]_ ;
  assign \new_[3197]_  = ~\new_[3385]_  | ~\new_[3460]_ ;
  assign \new_[3198]_  = ~\new_[3433]_  | ~\new_[19203]_ ;
  assign \new_[3199]_  = ~\new_[20413]_  | ~\new_[3506]_ ;
  assign \new_[3200]_  = ~\new_[21586]_  | ~\new_[3417]_ ;
  assign \new_[3201]_  = ~\new_[3431]_  | ~\new_[19408]_ ;
  assign \new_[3202]_  = ~\new_[3433]_  | ~\new_[18209]_ ;
  assign \new_[3203]_  = ~\new_[19853]_  | ~\new_[19760]_ ;
  assign \new_[3204]_  = ~\new_[3371]_ ;
  assign \new_[3205]_  = ~\new_[3372]_ ;
  assign \new_[3206]_  = ~\new_[3431]_  | ~\new_[19520]_ ;
  assign \new_[3207]_  = ~\new_[20309]_  | ~\new_[4420]_ ;
  assign \new_[3208]_  = ~\new_[3431]_  | ~\new_[18011]_ ;
  assign \new_[3209]_  = ~\new_[3433]_  | ~\new_[19156]_ ;
  assign \new_[3210]_  = \new_[3679]_  | \new_[3887]_  | \new_[7107]_  | \new_[9931]_ ;
  assign \new_[3211]_  = ~\new_[3606]_  | ~\new_[3433]_ ;
  assign \new_[3212]_  = ~\new_[3667]_  | ~\new_[3431]_ ;
  assign \new_[3213]_  = \new_[3640]_  ? \new_[20203]_  : \new_[3685]_ ;
  assign \new_[3214]_  = \new_[3723]_  | \new_[9894]_  | \new_[4104]_  | \new_[3933]_ ;
  assign \new_[3215]_  = ~\new_[3569]_  | (~\new_[21530]_  & ~\new_[19739]_ );
  assign \new_[3216]_  = ~\new_[20667]_ ;
  assign \new_[3217]_  = ~\new_[20667]_ ;
  assign \new_[3218]_  = \new_[6249]_  ^ \new_[3656]_ ;
  assign \new_[3219]_  = \new_[3703]_  ? \new_[20120]_  : \new_[20329]_ ;
  assign \new_[3220]_  = \new_[3708]_  ? \new_[21648]_  : \new_[3673]_ ;
  assign n2683 = \new_[19195]_  ^ \new_[3664]_ ;
  assign n2688 = \new_[1432]_  ^ \new_[3663]_ ;
  assign \new_[3223]_  = \new_[1637]_  ^ \new_[3656]_ ;
  assign \new_[3224]_  = \new_[19853]_ ;
  assign \new_[3225]_  = ~\new_[3385]_ ;
  assign \new_[3226]_  = ~\new_[3563]_  | (~\new_[21471]_  & ~\new_[19610]_ );
  assign \new_[3227]_  = ~\new_[3564]_  | (~\new_[3666]_  & ~\new_[19658]_ );
  assign \new_[3228]_  = ~\new_[3566]_  | (~\new_[21471]_  & ~\new_[19763]_ );
  assign \new_[3229]_  = ~\new_[3590]_  | ~\new_[1418]_ ;
  assign \new_[3230]_  = ~\new_[3590]_  | ~\new_[1515]_ ;
  assign \new_[3231]_  = ~\new_[3590]_  | ~\new_[1666]_ ;
  assign \new_[3232]_  = ~\new_[3575]_  | ~\new_[19704]_ ;
  assign \new_[3233]_  = ~\new_[21648]_  | ~\new_[3613]_ ;
  assign \new_[3234]_  = ~\new_[3586]_  | ~\new_[21085]_ ;
  assign \new_[3235]_  = ~\new_[3582]_  | ~\new_[21445]_ ;
  assign \new_[3236]_  = ~\new_[20546]_  | ~\new_[3619]_ ;
  assign \new_[3237]_  = ~\new_[3585]_  | ~\new_[20048]_ ;
  assign \new_[3238]_  = ~\new_[3607]_  | ~\new_[19114]_ ;
  assign \new_[3239]_  = ~\new_[19954]_  | ~\new_[3623]_ ;
  assign \new_[3240]_  = ~\new_[20342]_  | ~\new_[18998]_ ;
  assign \new_[3241]_  = ~\new_[21332]_ ;
  assign \new_[3242]_  = ~\new_[21618]_ ;
  assign \new_[3243]_  = ~\new_[3396]_ ;
  assign \new_[3244]_  = ~\new_[3591]_  | ~\new_[19766]_ ;
  assign \new_[3245]_  = ~\new_[3605]_  | ~\new_[18025]_ ;
  assign \new_[3246]_  = ~\new_[19978]_ ;
  assign \new_[3247]_  = ~\new_[20342]_  | ~\new_[18187]_ ;
  assign \new_[3248]_  = ~\new_[20185]_ ;
  assign \new_[3249]_  = \new_[3399]_ ;
  assign \new_[3250]_  = ~\new_[3399]_ ;
  assign \new_[3251]_  = ~\new_[3400]_ ;
  assign \new_[3252]_  = ~\new_[3605]_  | ~\new_[19308]_ ;
  assign \new_[3253]_  = ~\new_[20342]_  | ~\new_[19547]_ ;
  assign \new_[3254]_  = ~\new_[3594]_  | ~\new_[3706]_ ;
  assign \new_[3255]_  = ~\new_[3608]_  | ~\new_[5476]_ ;
  assign \new_[3256]_  = \new_[3716]_  | \new_[21377]_  | \new_[4671]_  | \new_[4128]_ ;
  assign \new_[3257]_  = \new_[20638]_  | \new_[3804]_  | \new_[4672]_  | \new_[4014]_ ;
  assign \new_[3258]_  = ~\new_[21285]_  | ~\new_[20342]_ ;
  assign \new_[3259]_  = ~\new_[3407]_ ;
  assign \new_[3260]_  = ~\new_[3605]_  | ~\new_[18765]_ ;
  assign \new_[3261]_  = ~\new_[3409]_ ;
  assign \new_[3262]_  = ~\new_[3412]_ ;
  assign \new_[3263]_  = ~\new_[3412]_ ;
  assign \new_[3264]_  = ~\new_[3601]_  | ~\new_[3861]_ ;
  assign \new_[3265]_  = ~\new_[19969]_ ;
  assign \new_[3266]_  = \new_[19969]_ ;
  assign \new_[3267]_  = ~\new_[3413]_ ;
  assign \new_[3268]_  = ~\new_[20391]_ ;
  assign \new_[3269]_  = ~\new_[20391]_ ;
  assign \new_[3270]_  = ~\new_[3415]_ ;
  assign \new_[3271]_  = \new_[3717]_  | \new_[21414]_  | \new_[4921]_  | \new_[4131]_ ;
  assign \new_[3272]_  = ~\new_[3416]_ ;
  assign \new_[3273]_  = ~\new_[3417]_ ;
  assign \new_[3274]_  = ~\new_[3605]_  | ~\new_[21277]_ ;
  assign \new_[3275]_  = \new_[20523]_ ;
  assign \new_[3276]_  = ~\new_[20523]_ ;
  assign \new_[3277]_  = ~\new_[21177]_ ;
  assign \new_[3278]_  = \new_[20687]_ ;
  assign \new_[3279]_  = ~\new_[20687]_ ;
  assign \new_[3280]_  = ~\new_[3588]_  | ~\new_[1509]_ ;
  assign n2678 = \new_[2511]_  ^ \new_[20322]_ ;
  assign \new_[3282]_  = ~\new_[3588]_  | ~\new_[1660]_ ;
  assign \new_[3283]_  = ~\new_[3588]_  | ~\new_[1353]_ ;
  assign \new_[3284]_  = ~\new_[3436]_ ;
  assign \new_[3285]_  = \new_[3436]_ ;
  assign \new_[3286]_  = ~\new_[3454]_ ;
  assign \new_[3287]_  = ~\new_[3455]_ ;
  assign \new_[3288]_  = ~\new_[3459]_ ;
  assign \new_[3289]_  = ~\new_[3461]_ ;
  assign \new_[3290]_  = ~\new_[3462]_ ;
  assign \new_[3291]_  = ~\new_[3465]_ ;
  assign \new_[3292]_  = ~\new_[20076]_ ;
  assign \new_[3293]_  = ~\new_[20068]_ ;
  assign \new_[3294]_  = ~\new_[3616]_  | ~\new_[21445]_ ;
  assign \new_[3295]_  = ~\new_[3611]_  | ~\new_[3614]_ ;
  assign \new_[3296]_  = ~\new_[21590]_  | ~\new_[20629]_ ;
  assign \new_[3297]_  = ~\new_[3472]_ ;
  assign \new_[3298]_  = ~\new_[3476]_ ;
  assign \new_[3299]_  = ~\new_[3477]_ ;
  assign \new_[3300]_  = ~\new_[3477]_ ;
  assign \new_[3301]_  = \new_[3482]_ ;
  assign \new_[3302]_  = ~\new_[3487]_ ;
  assign \new_[3303]_  = ~\new_[3489]_ ;
  assign \new_[3304]_  = \new_[19025]_  ^ \new_[21683]_ ;
  assign \new_[3305]_  = \new_[18205]_  ^ \new_[21683]_ ;
  assign \new_[3306]_  = \new_[2079]_  ^ \new_[3683]_ ;
  assign \new_[3307]_  = \new_[8021]_  ^ \new_[21683]_ ;
  assign \new_[3308]_  = ~\new_[3627]_  | (~\new_[3722]_  & ~\new_[6223]_ );
  assign \new_[3309]_  = ~\new_[3498]_ ;
  assign \new_[3310]_  = \new_[3730]_  ? \new_[3681]_  : \new_[3688]_ ;
  assign \new_[3311]_  = ~\new_[20873]_ ;
  assign \new_[3312]_  = ~\new_[20873]_ ;
  assign \new_[3313]_  = ~\new_[21187]_ ;
  assign \new_[3314]_  = ~\new_[3505]_ ;
  assign \new_[3315]_  = ~\new_[3507]_ ;
  assign \new_[3316]_  = ~\new_[3513]_ ;
  assign \new_[3317]_  = ~\new_[3514]_ ;
  assign \new_[3318]_  = ~\new_[3516]_ ;
  assign \new_[3319]_  = ~\new_[3521]_ ;
  assign \new_[3320]_  = ~\new_[21003]_ ;
  assign \new_[3321]_  = ~\new_[3523]_ ;
  assign \new_[3322]_  = ~\new_[3524]_ ;
  assign \new_[3323]_  = ~\new_[3525]_ ;
  assign \new_[3324]_  = ~\new_[3525]_ ;
  assign \new_[3325]_  = ~\new_[3526]_ ;
  assign \new_[3326]_  = ~\new_[3527]_ ;
  assign \new_[3327]_  = ~\new_[20054]_ ;
  assign \new_[3328]_  = ~\new_[3528]_ ;
  assign \new_[3329]_  = ~\new_[3528]_ ;
  assign \new_[3330]_  = ~\new_[3531]_ ;
  assign \new_[3331]_  = ~\new_[3534]_ ;
  assign \new_[3332]_  = \new_[3709]_  ? \new_[20352]_  : \new_[3677]_ ;
  assign \new_[3333]_  = ~\new_[3535]_ ;
  assign \new_[3334]_  = ~\new_[3537]_ ;
  assign \new_[3335]_  = ~\new_[3537]_ ;
  assign \new_[3336]_  = ~\new_[3541]_ ;
  assign \new_[3337]_  = ~\new_[3648]_  | ~\new_[1343]_ ;
  assign \new_[3338]_  = ~\new_[3648]_  | ~\new_[19606]_ ;
  assign \new_[3339]_  = ~\new_[3648]_  | ~\new_[19753]_ ;
  assign \new_[3340]_  = \new_[20474]_ ;
  assign \new_[3341]_  = ~\new_[3542]_ ;
  assign \new_[3342]_  = ~\new_[3649]_  | (~\new_[20567]_  & ~\new_[1862]_ );
  assign n2693 = \new_[1675]_  ^ \new_[19901]_ ;
  assign \new_[3344]_  = ~\new_[3650]_  | (~\new_[20567]_  & ~\new_[19731]_ );
  assign \new_[3345]_  = ~\new_[3545]_ ;
  assign \new_[3346]_  = \new_[19882]_ ;
  assign \new_[3347]_  = ~\new_[3546]_ ;
  assign \new_[3348]_  = ~\new_[3546]_ ;
  assign \new_[3349]_  = ~\new_[3652]_  | ~\new_[2511]_ ;
  assign \new_[3350]_  = ~\new_[3654]_  | (~\new_[20004]_  & ~\new_[3698]_ );
  assign \new_[3351]_  = ~\new_[3652]_  | ~\new_[1669]_ ;
  assign \new_[3352]_  = ~\new_[3652]_  | ~\new_[2079]_ ;
  assign \new_[3353]_  = ~\new_[3556]_ ;
  assign \new_[3354]_  = \new_[3556]_ ;
  assign \new_[3355]_  = ~\new_[3558]_ ;
  assign \new_[3356]_  = ~\new_[21485]_  | ~\new_[19561]_ ;
  assign \new_[3357]_  = ~\new_[3586]_  | ~\new_[20854]_ ;
  assign \new_[3358]_  = ~\new_[3582]_  | ~\new_[21027]_ ;
  assign \new_[3359]_  = ~\new_[21487]_  | ~\new_[18757]_ ;
  assign \new_[3360]_  = ~\new_[20101]_  | ~\new_[19578]_ ;
  assign \new_[3361]_  = ~\new_[3706]_  | ~\new_[21473]_ ;
  assign \new_[3362]_  = \new_[3707]_  | \new_[21473]_ ;
  assign \new_[3363]_  = \new_[3617]_  | \new_[21027]_ ;
  assign \new_[3364]_  = ~\new_[3616]_  | ~\new_[21027]_ ;
  assign \new_[3365]_  = \new_[3670]_  | \new_[20854]_ ;
  assign \new_[3366]_  = ~\new_[3669]_  | ~\new_[20854]_ ;
  assign \new_[3367]_  = ~\new_[3562]_  | ~\new_[19569]_ ;
  assign \new_[3368]_  = ~\new_[21590]_  | ~\new_[20550]_ ;
  assign \new_[3369]_  = ~\new_[3562]_  | ~\new_[19781]_ ;
  assign \new_[3370]_  = ~\new_[3562]_  | ~\new_[19682]_ ;
  assign \new_[3371]_  = ~\new_[20061]_ ;
  assign \new_[3372]_  = ~\new_[3573]_  | ~\new_[4988]_ ;
  assign \new_[3373]_  = \new_[19101]_  ^ \new_[3656]_ ;
  assign \new_[3374]_  = \new_[3712]_  | \new_[3980]_  | \new_[6377]_  | \new_[10943]_ ;
  assign \new_[3375]_  = \new_[3713]_  | \new_[3981]_  | \new_[6384]_  | \new_[10888]_ ;
  assign \new_[3376]_  = \new_[2344]_  ^ \new_[3697]_ ;
  assign \new_[3377]_  = \new_[17809]_  ^ \new_[3697]_ ;
  assign \new_[3378]_  = \new_[2291]_  ^ \new_[3697]_ ;
  assign \new_[3379]_  = \new_[10501]_  ^ \new_[3697]_ ;
  assign \new_[3380]_  = \new_[2294]_  ^ \new_[3695]_ ;
  assign \new_[3381]_  = \new_[2346]_  ^ \new_[21527]_ ;
  assign \new_[3382]_  = \new_[2293]_  ^ \new_[3695]_ ;
  assign \new_[3383]_  = \new_[17892]_  ^ \new_[3695]_ ;
  assign \new_[3384]_  = \new_[2288]_  ^ \new_[3694]_ ;
  assign \new_[3385]_  = ~\new_[3562]_ ;
  assign \new_[3386]_  = \new_[6947]_  ^ \new_[21527]_ ;
  assign \new_[3387]_  = \new_[6946]_  ^ \new_[3695]_ ;
  assign \new_[3388]_  = \new_[17604]_  ^ \new_[21527]_ ;
  assign \new_[3389]_  = ~\new_[3668]_  | ~\new_[16980]_ ;
  assign \new_[3390]_  = ~\new_[21699]_  | ~\new_[19783]_ ;
  assign \new_[3391]_  = ~\new_[3668]_  | ~\new_[18414]_ ;
  assign \new_[3392]_  = ~\new_[21700]_  | ~\new_[19631]_ ;
  assign \new_[3393]_  = ~\new_[21284]_  | ~\new_[18906]_ ;
  assign \new_[3394]_  = ~\new_[20577]_ ;
  assign \new_[3395]_  = ~\new_[3667]_  | ~\new_[18741]_ ;
  assign \new_[3396]_  = \new_[20577]_ ;
  assign \new_[3397]_  = ~\new_[20203]_  | ~\new_[3661]_ ;
  assign \new_[3398]_  = ~\new_[21284]_  | ~\new_[15923]_ ;
  assign \new_[3399]_  = ~\new_[7802]_  | ~\new_[7173]_  | ~\new_[3744]_  | ~\new_[3904]_ ;
  assign \new_[3400]_  = ~\new_[20131]_ ;
  assign \new_[3401]_  = ~\new_[20131]_ ;
  assign \new_[3402]_  = ~\new_[21530]_  | ~\new_[19805]_ ;
  assign \new_[3403]_  = ~\new_[3677]_  | ~\new_[21530]_ ;
  assign \new_[3404]_  = ~\new_[3660]_  | ~\new_[3709]_ ;
  assign \new_[3405]_  = ~\new_[3570]_ ;
  assign \new_[3406]_  = ~\new_[20854]_ ;
  assign \new_[3407]_  = ~\new_[20854]_ ;
  assign \new_[3408]_  = ~\new_[19842]_  & ~\new_[19847]_  & ~\new_[19852]_  & ~\new_[19850]_ ;
  assign \new_[3409]_  = ~\new_[3572]_ ;
  assign \new_[3410]_  = ~\new_[3572]_ ;
  assign \new_[3411]_  = ~\new_[21284]_  | ~\new_[18464]_ ;
  assign \new_[3412]_  = ~\new_[4415]_  | ~\new_[3789]_  | ~\new_[3739]_  | ~\new_[4129]_ ;
  assign \new_[3413]_  = \new_[20534]_  | \new_[3805]_  | \new_[4675]_  | \new_[4130]_ ;
  assign \new_[3414]_  = ~\new_[21027]_ ;
  assign \new_[3415]_  = ~\new_[21027]_ ;
  assign \new_[3416]_  = ~\new_[21473]_ ;
  assign \new_[3417]_  = ~\new_[20550]_ ;
  assign \new_[3418]_  = ~\new_[3891]_  & ~\new_[3665]_ ;
  assign \new_[3419]_  = ~\new_[3658]_  | ~\new_[19735]_ ;
  assign \new_[3420]_  = ~\new_[3657]_  | ~\new_[1739]_ ;
  assign \new_[3421]_  = ~\new_[3657]_  | ~\new_[1291]_ ;
  assign \new_[3422]_  = ~\new_[3658]_  | ~\new_[19579]_ ;
  assign \new_[3423]_  = ~\new_[3659]_  | ~\new_[19677]_ ;
  assign \new_[3424]_  = ~\new_[3659]_  | ~\new_[19595]_ ;
  assign \new_[3425]_  = \new_[2297]_  ^ \new_[3705]_ ;
  assign \new_[3426]_  = \new_[18556]_  ^ \new_[3705]_ ;
  assign \new_[3427]_  = \new_[2511]_  ^ \new_[3705]_ ;
  assign \new_[3428]_  = ~\new_[3657]_  | ~\new_[1424]_ ;
  assign \new_[3429]_  = \new_[9255]_  ^ \new_[3705]_ ;
  assign \new_[3430]_  = ~\new_[3659]_  | ~\new_[19814]_ ;
  assign \new_[3431]_  = ~\new_[20505]_  & ~\new_[20782]_  & ~\new_[4234]_  & ~\new_[5733]_ ;
  assign \new_[3432]_  = ~\new_[3659]_  | ~\new_[19776]_ ;
  assign \new_[3433]_  = \new_[20505]_  | \new_[20782]_  | \new_[4234]_  | \new_[5733]_ ;
  assign \new_[3434]_  = ~\new_[3575]_ ;
  assign \new_[3435]_  = \new_[19187]_  ^ \new_[3704]_ ;
  assign \new_[3436]_  = \new_[3738]_  | \new_[3923]_  | \new_[4230]_  | \new_[4976]_ ;
  assign \new_[3437]_  = \new_[17841]_  ^ \new_[3704]_ ;
  assign \new_[3438]_  = \new_[2509]_  ^ \new_[3704]_ ;
  assign \new_[3439]_  = \new_[10503]_  ^ \new_[3704]_ ;
  assign \new_[3440]_  = ~\new_[21626]_  | ~\new_[1663]_ ;
  assign \new_[3441]_  = ~\new_[3678]_  | ~\new_[19565]_ ;
  assign \new_[3442]_  = ~\new_[3675]_  | ~\new_[2297]_ ;
  assign \new_[3443]_  = ~\new_[3678]_  | ~\new_[19570]_ ;
  assign \new_[3444]_  = ~\new_[3675]_  | ~\new_[1419]_ ;
  assign \new_[3445]_  = ~\new_[3678]_  | ~\new_[21626]_ ;
  assign \new_[3446]_  = ~\new_[3676]_  | ~\new_[21627]_ ;
  assign \new_[3447]_  = ~\new_[3678]_  | ~\new_[19666]_ ;
  assign \new_[3448]_  = ~\new_[3675]_  | ~\new_[1665]_ ;
  assign \new_[3449]_  = ~\new_[3677]_  | ~\new_[2520]_ ;
  assign \new_[3450]_  = ~\new_[3678]_  | ~\new_[19768]_ ;
  assign \new_[3451]_  = ~\new_[3676]_  | ~\new_[1507]_ ;
  assign \new_[3452]_  = ~\new_[3677]_  | ~\new_[2078]_ ;
  assign \new_[3453]_  = ~\new_[21676]_ ;
  assign \new_[3454]_  = ~\new_[21677]_ ;
  assign \new_[3455]_  = ~\new_[20828]_ ;
  assign \new_[3456]_  = ~\new_[3582]_ ;
  assign \new_[3457]_  = ~\new_[3583]_ ;
  assign \new_[3458]_  = ~\new_[21646]_ ;
  assign \new_[3459]_  = ~\new_[21647]_ ;
  assign \new_[3460]_  = \new_[21647]_ ;
  assign \new_[3461]_  = ~\new_[20546]_ ;
  assign \new_[3462]_  = ~\new_[20546]_ ;
  assign \new_[3463]_  = ~\new_[3585]_ ;
  assign \new_[3464]_  = ~\new_[20596]_ ;
  assign \new_[3465]_  = ~\new_[20596]_ ;
  assign \new_[3466]_  = \new_[20596]_ ;
  assign \new_[3467]_  = ~\new_[3586]_ ;
  assign \new_[3468]_  = ~\new_[3587]_ ;
  assign \new_[3469]_  = ~\new_[9495]_  | ~\new_[4599]_  | ~\new_[6004]_  | ~\new_[3715]_ ;
  assign \new_[3470]_  = ~\new_[3669]_  | ~\new_[21085]_ ;
  assign \new_[3471]_  = ~\new_[3590]_ ;
  assign \new_[3472]_  = ~\new_[3594]_ ;
  assign \new_[3473]_  = ~\new_[3595]_ ;
  assign \new_[3474]_  = ~\new_[3595]_ ;
  assign \new_[3475]_  = ~\new_[21230]_ ;
  assign \new_[3476]_  = \new_[21230]_ ;
  assign \new_[3477]_  = ~\new_[3596]_ ;
  assign \new_[3478]_  = ~\new_[3780]_  | ~\new_[9390]_  | ~\new_[3751]_  | ~\new_[3914]_ ;
  assign \new_[3479]_  = ~\new_[3998]_  | ~\new_[5296]_  | ~\new_[8242]_  | ~\new_[3726]_ ;
  assign \new_[3480]_  = ~\new_[3680]_  & (~\new_[6478]_  | ~\new_[19780]_ );
  assign \new_[3481]_  = ~\new_[3953]_  | ~\new_[9345]_  | ~\new_[3725]_ ;
  assign \new_[3482]_  = ~\new_[3884]_  | ~\new_[8243]_  | ~\new_[3727]_ ;
  assign \new_[3483]_  = ~\new_[3600]_ ;
  assign \new_[3484]_  = ~\new_[3840]_  | ~\new_[3746]_  | ~\new_[6380]_  | ~\new_[3827]_ ;
  assign \new_[3485]_  = ~\new_[3603]_ ;
  assign \new_[3486]_  = ~\new_[3604]_ ;
  assign \new_[3487]_  = ~\new_[3604]_ ;
  assign \new_[3488]_  = ~\new_[3604]_ ;
  assign \new_[3489]_  = ~\new_[3606]_ ;
  assign \new_[3490]_  = ~\new_[3728]_  & ~\new_[4339]_  & ~\new_[4132]_ ;
  assign \new_[3491]_  = \new_[3609]_ ;
  assign \new_[3492]_  = \new_[2300]_  ^ \new_[3721]_ ;
  assign \new_[3493]_  = \new_[19626]_  ^ \new_[3722]_ ;
  assign \new_[3494]_  = \new_[2301]_  ^ \new_[3721]_ ;
  assign \new_[3495]_  = \new_[8019]_  ^ \new_[3721]_ ;
  assign \new_[3496]_  = \new_[1510]_  ^ \new_[3722]_ ;
  assign \new_[3497]_  = \new_[18057]_  ^ \new_[3721]_ ;
  assign \new_[3498]_  = ~\new_[20342]_ ;
  assign \new_[3499]_  = ~\new_[3614]_ ;
  assign \new_[3500]_  = ~\new_[3614]_ ;
  assign \new_[3501]_  = ~\new_[3616]_ ;
  assign \new_[3502]_  = ~\new_[3616]_ ;
  assign \new_[3503]_  = ~\new_[3617]_ ;
  assign \new_[3504]_  = ~\new_[21445]_ ;
  assign \new_[3505]_  = ~\new_[21445]_ ;
  assign \new_[3506]_  = ~\new_[20612]_ ;
  assign \new_[3507]_  = \new_[20612]_ ;
  assign \new_[3508]_  = ~\new_[20612]_ ;
  assign \new_[3509]_  = ~\new_[20612]_ ;
  assign \new_[3510]_  = ~\new_[3620]_ ;
  assign \new_[3511]_  = ~\new_[3620]_ ;
  assign \new_[3512]_  = ~\new_[19829]_ ;
  assign \new_[3513]_  = ~\new_[19829]_ ;
  assign \new_[3514]_  = ~\new_[20077]_ ;
  assign \new_[3515]_  = ~\new_[20077]_ ;
  assign \new_[3516]_  = ~\new_[19943]_ ;
  assign \new_[3517]_  = ~\new_[3621]_ ;
  assign \new_[3518]_  = ~\new_[3621]_ ;
  assign \new_[3519]_  = ~\new_[3624]_ ;
  assign \new_[3520]_  = ~\new_[20053]_ ;
  assign \new_[3521]_  = ~\new_[3625]_ ;
  assign \new_[3522]_  = ~\new_[3628]_ ;
  assign \new_[3523]_  = ~\new_[19998]_ ;
  assign \new_[3524]_  = ~\new_[21002]_ ;
  assign \new_[3525]_  = ~\new_[3682]_  | ~\new_[6696]_ ;
  assign \new_[3526]_  = ~\new_[3630]_ ;
  assign \new_[3527]_  = ~\new_[20114]_ ;
  assign \new_[3528]_  = ~\new_[21260]_ ;
  assign \new_[3529]_  = ~\new_[3875]_  | (~\new_[3731]_  & ~\new_[19693]_ );
  assign \new_[3530]_  = ~\new_[3631]_ ;
  assign \new_[3531]_  = ~\new_[3632]_ ;
  assign \new_[3532]_  = ~\new_[3633]_ ;
  assign \new_[3533]_  = ~\new_[3634]_ ;
  assign \new_[3534]_  = ~\new_[3635]_ ;
  assign \new_[3535]_  = ~\new_[3637]_ ;
  assign \new_[3536]_  = ~\new_[3639]_ ;
  assign \new_[3537]_  = ~\new_[3641]_ ;
  assign \new_[3538]_  = ~\new_[3641]_ ;
  assign \new_[3539]_  = ~\new_[3642]_ ;
  assign \new_[3540]_  = ~\new_[3642]_ ;
  assign \new_[3541]_  = ~\new_[3644]_ ;
  assign \new_[3542]_  = ~\new_[3648]_ ;
  assign \new_[3543]_  = ~\new_[3690]_  | ~\new_[19796]_ ;
  assign \new_[3544]_  = ~\new_[20173]_ ;
  assign \new_[3545]_  = \new_[20173]_ ;
  assign \new_[3546]_  = ~\new_[20623]_ ;
  assign \new_[3547]_  = ~\new_[3693]_  | ~\new_[1421]_ ;
  assign \new_[3548]_  = ~\new_[3691]_  | ~\new_[19698]_ ;
  assign \new_[3549]_  = ~\new_[3693]_  | ~\new_[19802]_ ;
  assign \new_[3550]_  = ~\new_[3693]_  | ~\new_[19690]_ ;
  assign \new_[3551]_  = ~\new_[3692]_  | ~\new_[19657]_ ;
  assign \new_[3552]_  = ~\new_[3691]_  | ~\new_[2509]_ ;
  assign \new_[3553]_  = ~\new_[3692]_  | ~\new_[19562]_ ;
  assign \new_[3554]_  = ~\new_[3691]_  | ~\new_[1506]_ ;
  assign \new_[3555]_  = ~\new_[3693]_  | ~\new_[19632]_ ;
  assign \new_[3556]_  = \new_[3758]_  | \new_[4010]_  | \new_[4233]_  | \new_[4981]_ ;
  assign \new_[3557]_  = ~\new_[20846]_ ;
  assign \new_[3558]_  = \new_[20846]_ ;
  assign \new_[3559]_  = ~\new_[21488]_  | ~\new_[15893]_ ;
  assign \new_[3560]_  = ~\new_[19820]_  | ~\new_[20258]_ ;
  assign \new_[3561]_  = ~\new_[20413]_  | ~\new_[3707]_ ;
  assign \new_[3562]_  = \new_[21456]_ ;
  assign \new_[3563]_  = ~\new_[21471]_  | ~\new_[19610]_ ;
  assign \new_[3564]_  = ~\new_[21472]_  | ~\new_[19658]_ ;
  assign \new_[3565]_  = ~\new_[21285]_  | ~\new_[2500]_ ;
  assign \new_[3566]_  = ~\new_[21472]_  | ~\new_[19763]_ ;
  assign \new_[3567]_  = ~\new_[21285]_  | ~\new_[18773]_ ;
  assign \new_[3568]_  = ~\new_[3700]_  | ~\new_[20603]_ ;
  assign \new_[3569]_  = ~\new_[21531]_  | ~\new_[19739]_ ;
  assign \new_[3570]_  = ~\new_[3655]_ ;
  assign \new_[3571]_  = ~\new_[3655]_ ;
  assign \new_[3572]_  = ~\new_[20259]_ ;
  assign \new_[3573]_  = ~\new_[3896]_  & ~\new_[21437]_ ;
  assign \new_[3574]_  = \new_[9330]_  ^ \new_[3736]_ ;
  assign \new_[3575]_  = \new_[21700]_ ;
  assign \new_[3576]_  = \new_[1929]_  ^ \new_[3736]_ ;
  assign \new_[3577]_  = \new_[19699]_  ^ \new_[3736]_ ;
  assign \new_[3578]_  = ~\new_[21627]_  | ~\new_[19797]_ ;
  assign \new_[3579]_  = ~\new_[21627]_  | ~\new_[19810]_ ;
  assign \new_[3580]_  = ~\new_[3709]_  | ~\new_[19616]_ ;
  assign \new_[3581]_  = ~\new_[3709]_  | ~\new_[19673]_ ;
  assign \new_[3582]_  = ~\new_[20121]_ ;
  assign \new_[3583]_  = ~\new_[20121]_ ;
  assign \new_[3584]_  = \new_[19955]_ ;
  assign \new_[3585]_  = ~\new_[19955]_ ;
  assign \new_[3586]_  = ~\new_[21649]_ ;
  assign \new_[3587]_  = ~\new_[21649]_ ;
  assign \new_[3588]_  = ~\new_[3658]_ ;
  assign \new_[3589]_  = ~\new_[3659]_ ;
  assign \new_[3590]_  = ~\new_[20352]_ ;
  assign \new_[3591]_  = ~\new_[3660]_ ;
  assign \new_[3592]_  = ~\new_[3745]_  | ~\new_[4289]_  | ~\new_[4013]_ ;
  assign \new_[3593]_  = ~\new_[3661]_ ;
  assign \new_[3594]_  = ~\new_[3661]_ ;
  assign \new_[3595]_  = ~\new_[20436]_ ;
  assign \new_[3596]_  = \new_[20145]_  | \new_[4127]_  | \new_[7757]_  | \new_[4244]_ ;
  assign \new_[3597]_  = ~\new_[3711]_  | ~\new_[5905]_ ;
  assign \new_[3598]_  = ~\new_[3888]_  | ~\new_[6394]_  | ~\new_[3741]_ ;
  assign \new_[3599]_  = ~\new_[3826]_  | ~\new_[8240]_  | ~\new_[3769]_  | ~\new_[3945]_ ;
  assign \new_[3600]_  = ~\new_[3876]_  | ~\new_[6957]_  | ~\new_[3737]_ ;
  assign \new_[3601]_  = ~\new_[3714]_  & (~\new_[8192]_  | ~\new_[18506]_ );
  assign \new_[3602]_  = ~\new_[3829]_  | ~\new_[3742]_  | ~\new_[7129]_ ;
  assign \new_[3603]_  = ~\new_[3666]_ ;
  assign \new_[3604]_  = ~\new_[19914]_ ;
  assign \new_[3605]_  = ~\new_[3668]_ ;
  assign \new_[3606]_  = ~\new_[21284]_ ;
  assign \new_[3607]_  = ~\new_[21284]_ ;
  assign \new_[3608]_  = ~\new_[3743]_  & ~\new_[4355]_  & ~\new_[4136]_ ;
  assign \new_[3609]_  = ~\new_[10787]_  | ~\new_[8288]_  | ~\new_[3720]_  | ~\new_[10911]_ ;
  assign \new_[3610]_  = ~\new_[3669]_ ;
  assign \new_[3611]_  = ~\new_[3669]_ ;
  assign \new_[3612]_  = ~\new_[3670]_ ;
  assign \new_[3613]_  = ~\new_[21085]_ ;
  assign \new_[3614]_  = ~\new_[21085]_ ;
  assign \new_[3615]_  = ~\new_[4098]_  | ~\new_[3719]_  | ~\new_[6360]_ ;
  assign \new_[3616]_  = ~\new_[20017]_ ;
  assign \new_[3617]_  = ~\new_[20017]_ ;
  assign \new_[3618]_  = ~\new_[3724]_  | ~\new_[3899]_ ;
  assign \new_[3619]_  = ~\new_[20629]_ ;
  assign \new_[3620]_  = ~\new_[20629]_ ;
  assign \new_[3621]_  = ~\new_[20539]_ ;
  assign \new_[3622]_  = ~\new_[21276]_ ;
  assign \new_[3623]_  = ~\new_[3671]_ ;
  assign \new_[3624]_  = \new_[3671]_ ;
  assign \new_[3625]_  = ~\new_[3673]_ ;
  assign \new_[3626]_  = ~\new_[3674]_ ;
  assign \new_[3627]_  = ~\new_[3722]_  | ~\new_[6223]_ ;
  assign \new_[3628]_  = ~\new_[20223]_ ;
  assign \new_[3629]_  = ~\new_[20119]_ ;
  assign \new_[3630]_  = ~\new_[3678]_ ;
  assign \new_[3631]_  = ~\new_[19902]_ ;
  assign \new_[3632]_  = ~\new_[3729]_  | ~\new_[3790]_ ;
  assign \new_[3633]_  = ~\new_[3681]_ ;
  assign \new_[3634]_  = ~\new_[21376]_ ;
  assign \new_[3635]_  = ~\new_[20943]_ ;
  assign \new_[3636]_  = ~\new_[20943]_ ;
  assign \new_[3637]_  = ~\new_[3684]_ ;
  assign \new_[3638]_  = ~\new_[3684]_ ;
  assign \new_[3639]_  = ~\new_[3685]_ ;
  assign \new_[3640]_  = ~\new_[3685]_ ;
  assign \new_[3641]_  = ~\new_[3733]_  | (~\new_[3822]_  & ~\new_[964]_ );
  assign \new_[3642]_  = ~\new_[3686]_ ;
  assign \new_[3643]_  = ~\new_[3686]_ ;
  assign \new_[3644]_  = ~\new_[3818]_  | ~\new_[3732]_ ;
  assign \new_[3645]_  = ~\new_[3687]_ ;
  assign \new_[3646]_  = ~\new_[3687]_ ;
  assign \new_[3647]_  = ~\new_[3689]_ ;
  assign \new_[3648]_  = \new_[20025]_ ;
  assign \new_[3649]_  = ~\new_[20568]_  | ~\new_[1862]_ ;
  assign \new_[3650]_  = ~\new_[20568]_  | ~\new_[19731]_ ;
  assign \new_[3651]_  = ~\new_[3690]_ ;
  assign \new_[3652]_  = ~\new_[3692]_ ;
  assign \new_[3653]_  = ~\new_[3693]_ ;
  assign \new_[3654]_  = ~\new_[20004]_  | ~\new_[3699]_ ;
  assign \new_[3655]_  = ~\new_[20005]_ ;
  assign \new_[3656]_  = ~\new_[3824]_  | ~\new_[3847]_  | ~\new_[5472]_  | ~\new_[4020]_ ;
  assign \new_[3657]_  = \new_[3696]_ ;
  assign \new_[3658]_  = ~\new_[3696]_ ;
  assign \new_[3659]_  = ~\new_[3696]_ ;
  assign \new_[3660]_  = ~\new_[21531]_ ;
  assign \new_[3661]_  = ~\new_[20603]_ ;
  assign \new_[3662]_  = ~\new_[3698]_ ;
  assign \new_[3663]_  = ~\new_[3698]_ ;
  assign \new_[3664]_  = ~\new_[3700]_ ;
  assign \new_[3665]_  = ~\new_[4085]_  | ~\new_[5426]_  | ~\new_[3799]_  | ~\new_[8607]_ ;
  assign \new_[3666]_  = \new_[21472]_ ;
  assign \new_[3667]_  = ~\new_[21285]_ ;
  assign \new_[3668]_  = ~\new_[21285]_ ;
  assign \new_[3669]_  = ~\new_[20952]_ ;
  assign \new_[3670]_  = ~\new_[20952]_ ;
  assign \new_[3671]_  = ~\new_[20049]_ ;
  assign \new_[3672]_  = ~\new_[3708]_ ;
  assign \new_[3673]_  = ~\new_[3708]_ ;
  assign \new_[3674]_  = \new_[3708]_ ;
  assign \new_[3675]_  = ~\new_[3709]_ ;
  assign \new_[3676]_  = ~\new_[3709]_ ;
  assign \new_[3677]_  = \new_[3710]_ ;
  assign \new_[3678]_  = ~\new_[3710]_ ;
  assign \new_[3679]_  = ~\new_[3750]_  | (~\new_[3844]_  & ~\new_[19391]_ );
  assign \new_[3680]_  = ~\new_[4045]_  | (~\new_[3776]_  & ~\new_[19661]_ );
  assign \new_[3681]_  = ~\new_[21639]_  | ~\new_[3833]_ ;
  assign \new_[3682]_  = ~\new_[3718]_ ;
  assign \new_[3683]_  = ~\new_[4054]_  | ~\new_[3835]_  | ~\new_[7123]_  | ~\new_[3915]_ ;
  assign \new_[3684]_  = ~\new_[3757]_  | (~\new_[3787]_  & ~\new_[18483]_ );
  assign \new_[3685]_  = ~\new_[20792]_  | ~\new_[3747]_ ;
  assign \new_[3686]_  = ~\new_[3755]_  | ~\new_[3871]_ ;
  assign \new_[3687]_  = ~\new_[3730]_ ;
  assign \new_[3688]_  = ~\new_[3730]_ ;
  assign \new_[3689]_  = ~\new_[21375]_ ;
  assign \new_[3690]_  = \new_[20568]_ ;
  assign \new_[3691]_  = \new_[3734]_ ;
  assign \new_[3692]_  = ~\new_[3734]_ ;
  assign \new_[3693]_  = ~\new_[3734]_ ;
  assign \new_[3694]_  = ~\new_[3880]_  | ~\new_[3846]_  | ~\new_[5054]_  | ~\new_[4019]_ ;
  assign \new_[3695]_  = ~\new_[3882]_  | ~\new_[3848]_  | ~\new_[6006]_  | ~\new_[4021]_ ;
  assign \new_[3696]_  = ~\new_[3735]_ ;
  assign \new_[3697]_  = ~\new_[3793]_  | ~\new_[4287]_  | ~\new_[4123]_ ;
  assign \new_[3698]_  = ~\new_[21006]_ ;
  assign \new_[3699]_  = ~\new_[21006]_ ;
  assign \new_[3700]_  = ~\new_[20203]_ ;
  assign \new_[3701]_  = ~\new_[20329]_ ;
  assign \new_[3702]_  = ~\new_[20329]_ ;
  assign \new_[3703]_  = ~\new_[20329]_ ;
  assign \new_[3704]_  = ~\new_[6364]_  | ~\new_[4099]_  | ~\new_[3768]_  | ~\new_[3878]_ ;
  assign \new_[3705]_  = ~\new_[4150]_  | ~\new_[3764]_  | ~\new_[4012]_ ;
  assign \new_[3706]_  = ~\new_[21278]_ ;
  assign \new_[3707]_  = ~\new_[21278]_ ;
  assign \new_[3708]_  = ~\new_[20752]_  | ~\new_[4004]_ ;
  assign \new_[3709]_  = \new_[20908]_ ;
  assign \new_[3710]_  = ~\new_[20908]_ ;
  assign \new_[3711]_  = ~\new_[3759]_  & (~\new_[4096]_  | ~\new_[19340]_ );
  assign \new_[3712]_  = ~\new_[3792]_  | ~\new_[3770]_ ;
  assign \new_[3713]_  = ~\new_[3771]_  | (~\new_[3845]_  & ~\new_[1243]_ );
  assign \new_[3714]_  = ~\new_[3941]_  | (~\new_[3803]_  & ~\new_[19672]_ );
  assign \new_[3715]_  = ~\new_[3777]_  & (~\new_[4746]_  | ~\new_[19780]_ );
  assign \new_[3716]_  = ~\new_[21008]_  & (~\new_[3820]_  | ~\new_[6296]_ );
  assign \new_[3717]_  = ~\new_[19017]_  & (~\new_[3821]_  | ~\new_[6303]_ );
  assign \new_[3718]_  = ~\new_[5013]_  | ~\new_[3902]_  | ~\new_[3832]_  | ~\new_[3898]_ ;
  assign \new_[3719]_  = ~\new_[3877]_  & (~\new_[3808]_  | ~\new_[19693]_ );
  assign \new_[3720]_  = ~\new_[3775]_  & (~\new_[3860]_  | ~\new_[19765]_ );
  assign \new_[3721]_  = ~\new_[3886]_  | ~\new_[3905]_  | ~\new_[6367]_  | ~\new_[3838]_ ;
  assign \new_[3722]_  = ~\new_[3890]_  | ~\new_[3906]_  | ~\new_[7115]_  | ~\new_[3992]_ ;
  assign \new_[3723]_  = ~\new_[3788]_  | ~\new_[11601]_ ;
  assign \new_[3724]_  = ~\new_[3772]_  & (~\new_[4251]_  | ~\new_[19340]_ );
  assign \new_[3725]_  = ~\new_[3765]_  & (~\new_[3989]_  | ~\new_[19396]_ );
  assign \new_[3726]_  = (~\new_[3816]_  | ~\new_[1243]_ ) & (~\new_[4429]_  | ~\new_[19452]_ );
  assign \new_[3727]_  = (~\new_[3817]_  | ~\new_[1675]_ ) & (~\new_[3983]_  | ~\new_[19693]_ );
  assign \new_[3728]_  = ~\new_[3825]_  | (~\new_[3810]_  & ~\new_[20310]_ );
  assign \new_[3729]_  = ~\new_[3748]_ ;
  assign \new_[3730]_  = ~\new_[3779]_  | ~\new_[3819]_ ;
  assign \new_[3731]_  = ~\new_[3754]_ ;
  assign \new_[3732]_  = ~\new_[3837]_  & (~\new_[20979]_  | ~\new_[20452]_ );
  assign \new_[3733]_  = ~\new_[19875]_  & (~\new_[3987]_  | ~\new_[964]_ );
  assign \new_[3734]_  = ~\new_[21350]_ ;
  assign \new_[3735]_  = ~\new_[3841]_  | ~\new_[4000]_  | ~\new_[4031]_ ;
  assign \new_[3736]_  = ~\new_[9352]_  | ~\new_[4241]_  | ~\new_[3798]_  | ~\new_[3879]_ ;
  assign \new_[3737]_  = ~\new_[1519]_  | (~\new_[3868]_  & ~\new_[5913]_ );
  assign \new_[3738]_  = ~\new_[19786]_  & (~\new_[3855]_  | ~\new_[6298]_ );
  assign \new_[3739]_  = ~\new_[964]_  | (~\new_[3870]_  & ~\new_[5878]_ );
  assign \new_[3740]_  = ~\new_[4226]_  | ~\new_[3797]_ ;
  assign \new_[3741]_  = ~\new_[3794]_  & (~\new_[4141]_  | ~\new_[19391]_ );
  assign \new_[3742]_  = ~\new_[3795]_  & (~\new_[4143]_  | ~\new_[1243]_ );
  assign \new_[3743]_  = ~\new_[3964]_  | (~\new_[3867]_  & ~\new_[19772]_ );
  assign \new_[3744]_  = ~\new_[3926]_  & (~\new_[3851]_  | ~\new_[21425]_ );
  assign \new_[3745]_  = (~\new_[3865]_  | ~\new_[1519]_ ) & (~\new_[4231]_  | ~\new_[19602]_ );
  assign \new_[3746]_  = ~\new_[5007]_  & ~\new_[3811]_ ;
  assign \new_[3747]_  = ~\new_[20772]_  | ~\new_[20295]_ ;
  assign \new_[3748]_  = ~\new_[4153]_  | ~\new_[3977]_  | ~\new_[3883]_  | ~\new_[5038]_ ;
  assign \new_[3749]_  = ~\new_[20418]_ ;
  assign \new_[3750]_  = ~\new_[3806]_  | ~\new_[1675]_ ;
  assign \new_[3751]_  = ~\new_[3812]_  | ~\new_[19396]_ ;
  assign \new_[3752]_  = ~\new_[3813]_  | ~\new_[937]_ ;
  assign \new_[3753]_  = (~\new_[21205]_  | ~\new_[3894]_ ) & (~\new_[4303]_  | ~\new_[19300]_ );
  assign \new_[3754]_  = ~\new_[3815]_  | ~\new_[5906]_ ;
  assign \new_[3755]_  = ~\new_[3976]_  & ~\new_[3836]_ ;
  assign \new_[3756]_  = ~\new_[3781]_ ;
  assign \new_[3757]_  = ~\new_[3839]_  & (~\new_[3986]_  | ~\new_[21452]_ );
  assign \new_[3758]_  = ~\new_[19564]_  & (~\new_[3857]_  | ~\new_[6300]_ );
  assign \new_[3759]_  = ~\new_[3843]_  | ~\new_[4211]_ ;
  assign \new_[3760]_  = ~\new_[19916]_  | (~\new_[20838]_  & ~\new_[5875]_ );
  assign \new_[3761]_  = ~\new_[994]_  | (~\new_[21018]_  & ~\new_[5881]_ );
  assign \new_[3762]_  = ~\new_[938]_  | (~\new_[3935]_  & ~\new_[6304]_ );
  assign \new_[3763]_  = ~\new_[19490]_  | (~\new_[20675]_  & ~\new_[11183]_ );
  assign \new_[3764]_  = ~\new_[3889]_  & (~\new_[4040]_  | ~\new_[19391]_ );
  assign \new_[3765]_  = ~\new_[3863]_  | (~\new_[7050]_  & ~\new_[17379]_ );
  assign \new_[3766]_  = ~\new_[20528]_  | (~\new_[3946]_  & ~\new_[10709]_ );
  assign \new_[3767]_  = ~\new_[19772]_  | (~\new_[3956]_  & ~\new_[6539]_ );
  assign \new_[3768]_  = ~\new_[19452]_  | (~\new_[3970]_  & ~\new_[7103]_ );
  assign \new_[3769]_  = ~\new_[3869]_  | ~\new_[19397]_ ;
  assign \new_[3770]_  = ~\new_[3852]_  | ~\new_[1519]_ ;
  assign \new_[3771]_  = ~\new_[3853]_  | ~\new_[19314]_ ;
  assign \new_[3772]_  = ~\new_[19340]_  & (~\new_[3971]_  | ~\new_[6391]_ );
  assign \new_[3773]_  = ~\new_[3866]_  | ~\new_[938]_ ;
  assign \new_[3774]_  = ~\new_[3858]_  | ~\new_[19807]_ ;
  assign \new_[3775]_  = ~\new_[4077]_  | (~\new_[3952]_  & ~\new_[19691]_ );
  assign \new_[3776]_  = ~\new_[3859]_  & (~\new_[9499]_  | ~\new_[19508]_ );
  assign \new_[3777]_  = ~\new_[3854]_  | ~\new_[4044]_ ;
  assign \new_[3778]_  = ~\new_[3901]_  | ~\new_[21205]_ ;
  assign \new_[3779]_  = ~\new_[3912]_  & ~\new_[3910]_ ;
  assign \new_[3780]_  = ~\new_[19691]_  | (~\new_[4003]_  & ~\new_[6153]_ );
  assign \new_[3781]_  = ~\new_[7365]_  | ~\new_[12116]_  | ~\new_[3908]_  | ~\new_[9812]_ ;
  assign \new_[3782]_  = ~\new_[8309]_  | ~\new_[4812]_  | ~\new_[4139]_  | ~\new_[7081]_ ;
  assign \new_[3783]_  = ~\new_[8422]_  & ~\new_[3909]_ ;
  assign \new_[3784]_  = ~\new_[7562]_  | ~\new_[4362]_  | ~\new_[4148]_  | ~\new_[7198]_ ;
  assign \new_[3785]_  = ~\new_[7591]_  | ~\new_[4363]_  | ~\new_[4149]_  | ~\new_[7209]_ ;
  assign \new_[3786]_  = ~\new_[3885]_  & (~\new_[4542]_  | ~\new_[19032]_ );
  assign \new_[3787]_  = ~\new_[4144]_  & ~\new_[3892]_ ;
  assign \new_[3788]_  = ~\new_[20783]_  | (~\new_[20088]_  & ~\new_[8971]_ );
  assign \new_[3789]_  = ~\new_[3920]_  | ~\new_[19807]_ ;
  assign \new_[3790]_  = ~\new_[6100]_  & (~\new_[4016]_  | ~\new_[958]_ );
  assign \new_[3791]_  = ~\new_[19470]_  | (~\new_[20332]_  & ~\new_[11371]_ );
  assign \new_[3792]_  = ~\new_[3924]_  | ~\new_[19602]_ ;
  assign \new_[3793]_  = (~\new_[4041]_  | ~\new_[19314]_ ) & (~\new_[4435]_  | ~\new_[19672]_ );
  assign \new_[3794]_  = ~\new_[3931]_  | (~\new_[6368]_  & ~\new_[18466]_ );
  assign \new_[3795]_  = ~\new_[3932]_  | (~\new_[7116]_  & ~\new_[18249]_ );
  assign \new_[3796]_  = ~\new_[21180]_  | (~\new_[4047]_  & ~\new_[11837]_ );
  assign \new_[3797]_  = ~\new_[19816]_  | (~\new_[4048]_  & ~\new_[7119]_ );
  assign \new_[3798]_  = ~\new_[19602]_  | (~\new_[4061]_  & ~\new_[7111]_ );
  assign \new_[3799]_  = ~\new_[3927]_  | ~\new_[20283]_ ;
  assign \new_[3800]_  = ~\new_[3937]_  | ~\new_[1004]_ ;
  assign \new_[3801]_  = ~\new_[3928]_  | ~\new_[20181]_ ;
  assign \new_[3802]_  = ~\new_[20914]_  | ~\new_[19273]_ ;
  assign \new_[3803]_  = ~\new_[3934]_  & (~\new_[8409]_  | ~\new_[19177]_ );
  assign \new_[3804]_  = ~\new_[19273]_  & (~\new_[4120]_  | ~\new_[4544]_ );
  assign \new_[3805]_  = ~\new_[19316]_  & (~\new_[21139]_  | ~\new_[4557]_ );
  assign \new_[3806]_  = ~\new_[8148]_  | ~\new_[4159]_  | ~\new_[4578]_  | ~\new_[7551]_ ;
  assign \new_[3807]_  = ~\new_[3966]_  | ~\new_[1004]_ ;
  assign \new_[3808]_  = \new_[4172]_  | \new_[7098]_  | \new_[6359]_  | \new_[9445]_ ;
  assign \new_[3809]_  = ~\new_[9473]_  & ~\new_[3974]_ ;
  assign \new_[3810]_  = ~\new_[9529]_  & ~\new_[3975]_ ;
  assign \new_[3811]_  = ~\new_[7196]_  | (~\new_[4075]_  & ~\new_[1519]_ );
  assign \new_[3812]_  = ~\new_[4281]_  | ~\new_[4912]_  | ~\new_[7573]_  | ~\new_[6338]_ ;
  assign \new_[3813]_  = ~\new_[8437]_  | ~\new_[4583]_  | ~\new_[4283]_  | ~\new_[7135]_ ;
  assign \new_[3814]_  = ~\new_[4284]_  | ~\new_[4815]_  | ~\new_[7434]_  | ~\new_[7140]_ ;
  assign \new_[3815]_  = ~\new_[3947]_  & (~\new_[5521]_  | ~\new_[19578]_ );
  assign \new_[3816]_  = ~\new_[4328]_  | ~\new_[4258]_  | ~\new_[9488]_  | ~\new_[9350]_ ;
  assign \new_[3817]_  = ~\new_[4329]_  | ~\new_[4261]_  | ~\new_[7405]_  | ~\new_[8112]_ ;
  assign \new_[3818]_  = ~\new_[5048]_  & (~\new_[4092]_  | ~\new_[964]_ );
  assign \new_[3819]_  = ~\new_[4707]_  & (~\new_[4093]_  | ~\new_[956]_ );
  assign \new_[3820]_  = ~\new_[3955]_  & (~\new_[4541]_  | ~\new_[18787]_ );
  assign \new_[3821]_  = ~\new_[3959]_  & (~\new_[20303]_  | ~\new_[19259]_ );
  assign \new_[3822]_  = ~\new_[4138]_  & ~\new_[3950]_ ;
  assign \new_[3823]_  = ~\new_[7924]_  | ~\new_[5005]_  | ~\new_[4266]_  | ~\new_[5731]_ ;
  assign \new_[3824]_  = ~\new_[3881]_ ;
  assign \new_[3825]_  = ~\new_[3984]_  | ~\new_[20310]_ ;
  assign \new_[3826]_  = ~\new_[19602]_  | (~\new_[4022]_  & ~\new_[5688]_ );
  assign \new_[3827]_  = \new_[4007]_  & \new_[12443]_ ;
  assign \new_[3828]_  = ~\new_[3985]_  | ~\new_[20452]_ ;
  assign \new_[3829]_  = \new_[4008]_  & \new_[12333]_ ;
  assign \new_[3830]_  = ~\new_[4009]_  | ~\new_[10638]_ ;
  assign \new_[3831]_  = ~\new_[4006]_  | ~\new_[20295]_ ;
  assign \new_[3832]_  = ~\new_[20794]_  | ~\new_[3995]_ ;
  assign \new_[3833]_  = ~\new_[5512]_  & (~\new_[4134]_  | ~\new_[950]_ );
  assign \new_[3834]_  = ~\new_[7748]_  & (~\new_[4135]_  | ~\new_[937]_ );
  assign \new_[3835]_  = ~\new_[3991]_  & (~\new_[4515]_  | ~\new_[18791]_ );
  assign \new_[3836]_  = ~\new_[3990]_  | ~\new_[4069]_ ;
  assign \new_[3837]_  = ~\new_[3993]_  | ~\new_[4070]_ ;
  assign \new_[3838]_  = ~\new_[4017]_  | ~\new_[1675]_ ;
  assign \new_[3839]_  = ~\new_[4942]_  | ~\new_[4029]_  | ~\new_[7377]_ ;
  assign \new_[3840]_  = ~\new_[4018]_  | ~\new_[1519]_ ;
  assign \new_[3841]_  = ~\new_[20361]_  | ~\new_[932]_ ;
  assign \new_[3842]_  = ~\new_[4042]_  | ~\new_[19316]_ ;
  assign \new_[3843]_  = ~\new_[4080]_  & (~\new_[4210]_  | ~\new_[19765]_ );
  assign \new_[3844]_  = ~\new_[4032]_  & ~\new_[6547]_ ;
  assign \new_[3845]_  = ~\new_[4033]_  & ~\new_[6551]_ ;
  assign \new_[3846]_  = ~\new_[4034]_  & (~\new_[4438]_  | ~\new_[19718]_ );
  assign \new_[3847]_  = ~\new_[4035]_  & (~\new_[4242]_  | ~\new_[19563]_ );
  assign \new_[3848]_  = ~\new_[4037]_  & (~\new_[4243]_  | ~\new_[19672]_ );
  assign \new_[3849]_  = ~\new_[4699]_  & ~\new_[4064]_ ;
  assign \new_[3850]_  = ~\new_[5266]_  | ~\new_[5955]_  | ~\new_[4704]_  | ~\new_[4484]_ ;
  assign \new_[3851]_  = ~\new_[5655]_  | ~\new_[6463]_  | ~\new_[4493]_  | ~\new_[5935]_ ;
  assign \new_[3852]_  = ~\new_[7118]_  | ~\new_[4311]_  | ~\new_[4813]_  | ~\new_[8442]_ ;
  assign \new_[3853]_  = ~\new_[8129]_  | ~\new_[4313]_  | ~\new_[4582]_  | ~\new_[8417]_ ;
  assign \new_[3854]_  = ~\new_[1517]_  | (~\new_[4217]_  & ~\new_[5143]_ );
  assign \new_[3855]_  = ~\new_[4052]_  & (~\new_[4497]_  | ~\new_[19002]_ );
  assign \new_[3856]_  = ~\new_[5460]_  | ~\new_[15028]_  | ~\new_[4073]_  | ~\new_[4793]_ ;
  assign \new_[3857]_  = ~\new_[4056]_  & (~\new_[4498]_  | ~\new_[19041]_ );
  assign \new_[3858]_  = ~\new_[4494]_  | ~\new_[6432]_  | ~\new_[5014]_  | ~\new_[6055]_ ;
  assign \new_[3859]_  = ~\new_[4471]_  | ~\new_[7049]_  | ~\new_[4450]_  | ~\new_[10768]_ ;
  assign \new_[3860]_  = ~\new_[13616]_  | ~\new_[13716]_  | ~\new_[4065]_  | ~\new_[5146]_ ;
  assign \new_[3861]_  = ~\new_[3930]_ ;
  assign \new_[3862]_  = ~\new_[7379]_  & ~\new_[4066]_ ;
  assign \new_[3863]_  = (~\new_[4218]_  | ~\new_[19691]_ ) & (~\new_[9494]_  | ~\new_[18594]_ );
  assign \new_[3864]_  = ~\new_[7004]_  | ~\new_[4430]_  | ~\new_[6188]_  | ~\new_[15497]_ ;
  assign \new_[3865]_  = ~\new_[5830]_  | ~\new_[4431]_  | ~\new_[5722]_  | ~\new_[17275]_ ;
  assign \new_[3866]_  = ~\new_[4483]_  | ~\new_[4814]_  | ~\new_[7447]_  | ~\new_[5924]_ ;
  assign \new_[3867]_  = ~\new_[6062]_  & ~\new_[4067]_ ;
  assign \new_[3868]_  = ~\new_[4478]_  | ~\new_[6372]_  | ~\new_[5058]_  | ~\new_[14291]_ ;
  assign \new_[3869]_  = ~\new_[4330]_  | ~\new_[4451]_  | ~\new_[7390]_  | ~\new_[7085]_ ;
  assign \new_[3870]_  = ~\new_[4481]_  | ~\new_[6171]_  | ~\new_[4516]_  | ~\new_[9284]_ ;
  assign \new_[3871]_  = ~\new_[5916]_  & (~\new_[949]_  | ~\new_[4228]_ );
  assign \new_[3872]_  = ~\new_[4050]_  & (~\new_[4558]_  | ~\new_[19051]_ );
  assign \new_[3873]_  = ~\new_[7797]_  | ~\new_[4463]_  | ~\new_[5390]_  | ~\new_[5570]_ ;
  assign \new_[3874]_  = ~\new_[21066]_  | (~\new_[4175]_  & ~\new_[4779]_ );
  assign \new_[3875]_  = ~\new_[4094]_  | ~\new_[19693]_ ;
  assign \new_[3876]_  = ~\new_[4095]_  | ~\new_[19563]_ ;
  assign \new_[3877]_  = ~\new_[19693]_  & (~\new_[4161]_  | ~\new_[5675]_ );
  assign \new_[3878]_  = ~\new_[1243]_  | (~\new_[4162]_  & ~\new_[5676]_ );
  assign \new_[3879]_  = ~\new_[1519]_  | (~\new_[4163]_  & ~\new_[5281]_ );
  assign \new_[3880]_  = ~\new_[3943]_ ;
  assign \new_[3881]_  = ~\new_[1878]_  & (~\new_[4160]_  | ~\new_[9540]_ );
  assign \new_[3882]_  = ~\new_[3944]_ ;
  assign \new_[3883]_  = ~\new_[20743]_  | (~\new_[4152]_  & ~\new_[13527]_ );
  assign \new_[3884]_  = \new_[4097]_  & \new_[5297]_ ;
  assign \new_[3885]_  = ~\new_[5285]_  | ~\new_[4277]_  | ~\new_[10680]_ ;
  assign \new_[3886]_  = ~\new_[4118]_  | ~\new_[19693]_ ;
  assign \new_[3887]_  = ~\new_[4100]_  | (~\new_[6791]_  & ~\new_[19578]_ );
  assign \new_[3888]_  = \new_[4106]_  & \new_[12311]_ ;
  assign \new_[3889]_  = ~\new_[1675]_  & (~\new_[4293]_  | ~\new_[4783]_ );
  assign \new_[3890]_  = ~\new_[4119]_  | ~\new_[19602]_ ;
  assign \new_[3891]_  = ~\new_[20950]_  & (~\new_[4155]_  | ~\new_[4344]_ );
  assign \new_[3892]_  = ~\new_[4371]_  | ~\new_[5438]_  | ~\new_[6024]_  | ~\new_[8313]_ ;
  assign \new_[3893]_  = ~\new_[5322]_  | ~\new_[4333]_  | ~\new_[4178]_  | ~\new_[5926]_ ;
  assign \new_[3894]_  = ~\new_[6902]_  | ~\new_[4352]_  | ~\new_[4904]_  | ~\new_[7171]_ ;
  assign \new_[3895]_  = ~\new_[4113]_  | ~\new_[12925]_ ;
  assign \new_[3896]_  = ~\new_[20295]_  & (~\new_[4156]_  | ~\new_[4353]_ );
  assign \new_[3897]_  = ~\new_[4115]_  | ~\new_[11943]_ ;
  assign \new_[3898]_  = \new_[4116]_  & \new_[10634]_ ;
  assign \new_[3899]_  = ~\new_[3967]_ ;
  assign \new_[3900]_  = ~\new_[6385]_  | ~\new_[4101]_ ;
  assign \new_[3901]_  = ~\new_[4121]_  | ~\new_[4350]_ ;
  assign \new_[3902]_  = ~\new_[5943]_  & (~\new_[4273]_  | ~\new_[19866]_ );
  assign \new_[3903]_  = ~\new_[5448]_  | (~\new_[4274]_  & ~\new_[956]_ );
  assign \new_[3904]_  = ~\new_[3973]_ ;
  assign \new_[3905]_  = ~\new_[4082]_  & (~\new_[4173]_  | ~\new_[18667]_ );
  assign \new_[3906]_  = ~\new_[4084]_  & (~\new_[4174]_  | ~\new_[19195]_ );
  assign \new_[3907]_  = (~\new_[4167]_  | ~\new_[19070]_ ) & (~\new_[14156]_  | ~\new_[18544]_ );
  assign \new_[3908]_  = (~\new_[4169]_  | ~\new_[1878]_ ) & (~\new_[16862]_  | ~\new_[11890]_ );
  assign \new_[3909]_  = ~\new_[8701]_  | ~\new_[5917]_  | ~\new_[4410]_  | ~\new_[4282]_ ;
  assign \new_[3910]_  = ~\new_[4088]_  | ~\new_[4071]_ ;
  assign \new_[3911]_  = ~\new_[4089]_  | ~\new_[4072]_ ;
  assign \new_[3912]_  = ~\new_[20140]_ ;
  assign \new_[3913]_  = ~\new_[3978]_ ;
  assign \new_[3914]_  = \new_[4151]_  & \new_[5719]_ ;
  assign \new_[3915]_  = ~\new_[4142]_  | ~\new_[1243]_ ;
  assign \new_[3916]_  = ~\new_[6716]_  | ~\new_[4666]_  | ~\new_[4028]_  | ~\new_[9973]_ ;
  assign \new_[3917]_  = ~\new_[950]_  | (~\new_[4193]_  & ~\new_[4940]_ );
  assign \new_[3918]_  = ~\new_[19816]_  & (~\new_[4194]_  | ~\new_[5236]_ );
  assign \new_[3919]_  = ~\new_[4319]_  | ~\new_[4140]_ ;
  assign \new_[3920]_  = ~\new_[4024]_  | (~\new_[4389]_  & ~\new_[18293]_ );
  assign \new_[3921]_  = ~\new_[4320]_  | ~\new_[4145]_ ;
  assign \new_[3922]_  = ~\new_[5571]_  | ~\new_[5313]_  | ~\new_[4417]_ ;
  assign \new_[3923]_  = ~\new_[19490]_  & (~\new_[4448]_  | ~\new_[4337]_ );
  assign \new_[3924]_  = ~\new_[5708]_  | ~\new_[4716]_  | ~\new_[6005]_  | ~\new_[5264]_ ;
  assign \new_[3925]_  = ~\new_[5984]_  | ~\new_[10505]_  | ~\new_[4214]_  | ~\new_[4800]_ ;
  assign \new_[3926]_  = ~\new_[19017]_  & (~\new_[4589]_  | ~\new_[4444]_ );
  assign \new_[3927]_  = ~\new_[5380]_  | ~\new_[6434]_  | ~\new_[4736]_  | ~\new_[6642]_ ;
  assign \new_[3928]_  = ~\new_[5012]_  | ~\new_[6427]_  | ~\new_[4744]_  | ~\new_[5490]_ ;
  assign \new_[3929]_  = ~\new_[4039]_ ;
  assign \new_[3930]_  = ~\new_[7358]_  | ~\new_[8277]_  | ~\new_[4212]_  | ~\new_[10927]_ ;
  assign \new_[3931]_  = (~\new_[4427]_  | ~\new_[19718]_ ) & (~\new_[7587]_  | ~\new_[1879]_ );
  assign \new_[3932]_  = (~\new_[4428]_  | ~\new_[19672]_ ) & (~\new_[8399]_  | ~\new_[19502]_ );
  assign \new_[3933]_  = \new_[4224]_  & \new_[930]_ ;
  assign \new_[3934]_  = ~\new_[4734]_  | ~\new_[7121]_  | ~\new_[5481]_  | ~\new_[15285]_ ;
  assign \new_[3935]_  = ~\new_[4742]_  | ~\new_[6175]_  | ~\new_[4326]_  | ~\new_[10697]_ ;
  assign \new_[3936]_  = ~\new_[7778]_  | ~\new_[4721]_  | ~\new_[5539]_  | ~\new_[5828]_ ;
  assign \new_[3937]_  = ~\new_[7776]_  | ~\new_[4722]_  | ~\new_[4409]_  | ~\new_[5025]_ ;
  assign \new_[3938]_  = ~\new_[7799]_  | ~\new_[4723]_  | ~\new_[4892]_  | ~\new_[6264]_ ;
  assign \new_[3939]_  = ~\new_[7824]_  | ~\new_[5598]_  | ~\new_[4725]_  | ~\new_[5392]_ ;
  assign \new_[3940]_  = ~\new_[4237]_  | ~\new_[20011]_ ;
  assign \new_[3941]_  = ~\new_[4232]_  | ~\new_[19672]_ ;
  assign \new_[3942]_  = ~\new_[4246]_  | ~\new_[19017]_ ;
  assign \new_[3943]_  = ~\new_[18667]_  & (~\new_[4307]_  | ~\new_[9518]_ );
  assign \new_[3944]_  = ~\new_[18791]_  & (~\new_[4312]_  | ~\new_[12131]_ );
  assign \new_[3945]_  = \new_[4240]_  & \new_[5303]_ ;
  assign \new_[3946]_  = ~\new_[6874]_  | ~\new_[4546]_  | ~\new_[5253]_  | ~\new_[8165]_ ;
  assign \new_[3947]_  = ~\new_[7102]_  | ~\new_[15262]_  | ~\new_[4474]_ ;
  assign \new_[3948]_  = ~\new_[4219]_  | ~\new_[20950]_ ;
  assign \new_[3949]_  = ~\new_[4220]_  | ~\new_[19816]_ ;
  assign \new_[3950]_  = ~\new_[4598]_  | ~\new_[5430]_  | ~\new_[5482]_  | ~\new_[7381]_ ;
  assign \new_[3951]_  = ~\new_[5349]_  | ~\new_[6186]_  | ~\new_[4454]_ ;
  assign \new_[3952]_  = ~\new_[4358]_  & ~\new_[4238]_ ;
  assign \new_[3953]_  = \new_[4252]_  & \new_[14946]_ ;
  assign \new_[3954]_  = ~\new_[5427]_  | ~\new_[4601]_  | ~\new_[8109]_  | ~\new_[4778]_ ;
  assign \new_[3955]_  = ~\new_[4472]_  | ~\new_[5686]_  | ~\new_[7966]_ ;
  assign \new_[3956]_  = ~\new_[6527]_  | ~\new_[6390]_  | ~\new_[4553]_  | ~\new_[9576]_ ;
  assign \new_[3957]_  = ~\new_[5363]_  | ~\new_[6199]_  | ~\new_[4457]_ ;
  assign \new_[3958]_  = ~\new_[4221]_  | ~\new_[21441]_ ;
  assign \new_[3959]_  = ~\new_[5691]_  | ~\new_[10400]_  | ~\new_[4486]_ ;
  assign \new_[3960]_  = ~\new_[5011]_  | ~\new_[13161]_  | ~\new_[4460]_ ;
  assign \new_[3961]_  = ~\new_[4255]_  | ~\new_[10708]_ ;
  assign \new_[3962]_  = ~\new_[6525]_  | ~\new_[5944]_  | ~\new_[4571]_  | ~\new_[7541]_ ;
  assign \new_[3963]_  = ~\new_[7285]_  | ~\new_[6442]_  | ~\new_[4573]_  | ~\new_[7565]_ ;
  assign \new_[3964]_  = ~\new_[4222]_  | ~\new_[19772]_ ;
  assign \new_[3965]_  = ~\new_[19017]_  | (~\new_[4301]_  & ~\new_[5291]_ );
  assign \new_[3966]_  = ~\new_[4955]_  | ~\new_[4646]_  | ~\new_[4453]_ ;
  assign \new_[3967]_  = ~\new_[4735]_  | ~\new_[4528]_  | ~\new_[9444]_  | ~\new_[12316]_ ;
  assign \new_[3968]_  = ~\new_[4687]_  | ~\new_[4408]_  | ~\new_[4456]_ ;
  assign \new_[3969]_  = ~\new_[5267]_  | ~\new_[4665]_  | ~\new_[4461]_ ;
  assign \new_[3970]_  = ~\new_[8712]_  | ~\new_[8264]_  | ~\new_[4321]_  | ~\new_[8292]_ ;
  assign \new_[3971]_  = ~\new_[4062]_ ;
  assign \new_[3972]_  = ~\new_[21205]_  & (~\new_[4300]_  | ~\new_[4681]_ );
  assign \new_[3973]_  = ~\new_[5824]_  | ~\new_[4604]_  | ~\new_[5871]_  | ~\new_[7513]_ ;
  assign \new_[3974]_  = ~\new_[8934]_  | ~\new_[6126]_  | ~\new_[7080]_  | ~\new_[4470]_ ;
  assign \new_[3975]_  = ~\new_[8635]_  | ~\new_[6433]_  | ~\new_[4649]_  | ~\new_[4476]_ ;
  assign \new_[3976]_  = ~\new_[4068]_ ;
  assign \new_[3977]_  = ~\new_[20645]_  | (~\new_[4346]_  & ~\new_[13527]_ );
  assign \new_[3978]_  = ~\new_[20295]_  | (~\new_[20551]_  & ~\new_[5990]_ );
  assign \new_[3979]_  = ~\new_[4076]_ ;
  assign \new_[3980]_  = ~\new_[5421]_  | ~\new_[4294]_  | ~\new_[8631]_ ;
  assign \new_[3981]_  = ~\new_[7024]_  | ~\new_[4295]_  | ~\new_[9768]_ ;
  assign \new_[3982]_  = ~\new_[5526]_  | ~\new_[4357]_  | ~\new_[6871]_ ;
  assign \new_[3983]_  = ~\new_[8239]_  | ~\new_[4682]_  | ~\new_[4971]_  | ~\new_[6129]_ ;
  assign \new_[3984]_  = ~\new_[5288]_  | ~\new_[6630]_  | ~\new_[4648]_  | ~\new_[5548]_ ;
  assign \new_[3985]_  = ~\new_[4652]_  | ~\new_[6032]_  | ~\new_[5289]_  | ~\new_[5559]_ ;
  assign \new_[3986]_  = ~\new_[4359]_  | ~\new_[5114]_  | ~\new_[6885]_ ;
  assign \new_[3987]_  = ~\new_[4364]_  | ~\new_[4632]_  | ~\new_[7983]_ ;
  assign \new_[3988]_  = ~\new_[4941]_  | ~\new_[7399]_  | ~\new_[4378]_ ;
  assign \new_[3989]_  = ~\new_[4168]_  | ~\new_[4935]_ ;
  assign \new_[3990]_  = ~\new_[4157]_  | ~\new_[18091]_ ;
  assign \new_[3991]_  = ~\new_[15893]_  & (~\new_[4388]_  | ~\new_[7432]_ );
  assign \new_[3992]_  = ~\new_[4279]_  | ~\new_[19397]_ ;
  assign \new_[3993]_  = ~\new_[20716]_  | ~\new_[17715]_ ;
  assign \new_[3994]_  = ~\new_[20743]_  | (~\new_[4356]_  & ~\new_[5135]_ );
  assign \new_[3995]_  = ~\new_[8456]_  | ~\new_[4906]_  | ~\new_[4189]_  | ~\new_[9903]_ ;
  assign \new_[3996]_  = ~\new_[7545]_  | ~\new_[4663]_  | ~\new_[4190]_  | ~\new_[9970]_ ;
  assign \new_[3997]_  = ~\new_[8434]_  | ~\new_[4644]_  | ~\new_[4187]_  | ~\new_[9803]_ ;
  assign \new_[3998]_  = ~\new_[4291]_  & (~\new_[5243]_  | ~\new_[15893]_ );
  assign \new_[3999]_  = ~\new_[20528]_  & (~\new_[4385]_  | ~\new_[5229]_ );
  assign \new_[4000]_  = ~\new_[4375]_  & ~\new_[4262]_ ;
  assign \new_[4001]_  = \new_[4288]_  & \new_[979]_ ;
  assign \new_[4002]_  = ~\new_[21180]_  & (~\new_[4384]_  | ~\new_[5237]_ );
  assign \new_[4003]_  = ~\new_[14024]_  | ~\new_[4679]_  | ~\new_[5562]_  | ~\new_[11459]_ ;
  assign \new_[4004]_  = ~\new_[4263]_  & (~\new_[4374]_  | ~\new_[19509]_ );
  assign \new_[4005]_  = ~\new_[4267]_  | (~\new_[5811]_  & ~\new_[19236]_ );
  assign \new_[4006]_  = ~\new_[4165]_  | (~\new_[4396]_  & ~\new_[18004]_ );
  assign \new_[4007]_  = (~\new_[4377]_  | ~\new_[19717]_ ) & (~\new_[10899]_  | ~\new_[19440]_ );
  assign \new_[4008]_  = (~\new_[4376]_  | ~\new_[18506]_ ) & (~\new_[9834]_  | ~\new_[19177]_ );
  assign \new_[4009]_  = (~\new_[4391]_  | ~\new_[19271]_ ) & (~\new_[10895]_  | ~\new_[19492]_ );
  assign \new_[4010]_  = ~\new_[19470]_  & (~\new_[4449]_  | ~\new_[4347]_ );
  assign \new_[4011]_  = (~\new_[4397]_  | ~\new_[19277]_ ) & (~\new_[11790]_  | ~\new_[18739]_ );
  assign \new_[4012]_  = ~\new_[19070]_  | (~\new_[4418]_  & ~\new_[4635]_ );
  assign \new_[4013]_  = ~\new_[19195]_  | (~\new_[4414]_  & ~\new_[4850]_ );
  assign \new_[4014]_  = ~\new_[4195]_  | ~\new_[9532]_ ;
  assign \new_[4015]_  = ~\new_[4196]_  & (~\new_[9246]_  | ~\new_[18752]_ );
  assign \new_[4016]_  = ~\new_[6653]_  | ~\new_[4197]_  | ~\new_[5239]_ ;
  assign \new_[4017]_  = ~\new_[6841]_  | ~\new_[9121]_  | ~\new_[4879]_  | ~\new_[4407]_ ;
  assign \new_[4018]_  = ~\new_[4191]_  | ~\new_[5227]_ ;
  assign \new_[4019]_  = ~\new_[4181]_  & (~\new_[9082]_  | ~\new_[17669]_ );
  assign \new_[4020]_  = ~\new_[4179]_  & (~\new_[7873]_  | ~\new_[18097]_ );
  assign \new_[4021]_  = ~\new_[8400]_  & ~\new_[4180]_ ;
  assign \new_[4022]_  = ~\new_[4677]_  | ~\new_[5552]_  | ~\new_[9393]_ ;
  assign \new_[4023]_  = ~\new_[9270]_  | ~\new_[4959]_  | ~\new_[5802]_  | ~\new_[8787]_ ;
  assign \new_[4024]_  = ~\new_[4164]_ ;
  assign \new_[4025]_  = ~\new_[5788]_  | (~\new_[4691]_  & ~\new_[19528]_ );
  assign \new_[4026]_  = ~\new_[19207]_  | (~\new_[4692]_  & ~\new_[10318]_ );
  assign \new_[4027]_  = ~\new_[19133]_  | (~\new_[4696]_  & ~\new_[8822]_ );
  assign \new_[4028]_  = ~\new_[4702]_  & ~\new_[6446]_  & ~\new_[13471]_ ;
  assign \new_[4029]_  = ~\new_[5470]_  & ~\new_[4405]_ ;
  assign \new_[4030]_  = ~\new_[5056]_  | ~\new_[11946]_  | ~\new_[12294]_  | ~\new_[11650]_ ;
  assign \new_[4031]_  = ~\new_[19786]_  | (~\new_[4533]_  & ~\new_[4654]_ );
  assign \new_[4032]_  = ~\new_[5263]_  | ~\new_[4422]_ ;
  assign \new_[4033]_  = ~\new_[4717]_  | ~\new_[5646]_  | ~\new_[8029]_ ;
  assign \new_[4034]_  = ~\new_[19718]_  & (~\new_[4708]_  | ~\new_[5547]_ );
  assign \new_[4035]_  = ~\new_[19563]_  & (~\new_[4710]_  | ~\new_[5157]_ );
  assign \new_[4036]_  = ~\new_[7257]_  | ~\new_[10521]_  | ~\new_[4426]_  | ~\new_[4785]_ ;
  assign \new_[4037]_  = ~\new_[19452]_  & (~\new_[4711]_  | ~\new_[5558]_ );
  assign \new_[4038]_  = ~\new_[7246]_  | ~\new_[12513]_  | ~\new_[4424]_  | ~\new_[4774]_ ;
  assign \new_[4039]_  = ~\new_[8266]_  | ~\new_[11037]_  | ~\new_[4423]_  | ~\new_[9444]_ ;
  assign \new_[4040]_  = ~\new_[5019]_  | ~\new_[5464]_  | ~\new_[6954]_  | ~\new_[15730]_ ;
  assign \new_[4041]_  = ~\new_[5831]_  | ~\new_[5052]_  | ~\new_[5716]_  | ~\new_[15593]_ ;
  assign \new_[4042]_  = ~\new_[7821]_  | ~\new_[5059]_  | ~\new_[4872]_  | ~\new_[5832]_ ;
  assign \new_[4043]_  = ~\new_[930]_  | (~\new_[4629]_  & ~\new_[5082]_ );
  assign \new_[4044]_  = ~\new_[4437]_  | ~\new_[19765]_ ;
  assign \new_[4045]_  = ~\new_[4442]_  | ~\new_[19661]_ ;
  assign \new_[4046]_  = ~\new_[19623]_  | (~\new_[4511]_  & ~\new_[12429]_ );
  assign \new_[4047]_  = ~\new_[6138]_  | ~\new_[4792]_  | ~\new_[4953]_  | ~\new_[8133]_ ;
  assign \new_[4048]_  = ~\new_[6897]_  | ~\new_[4802]_  | ~\new_[5258]_  | ~\new_[7159]_ ;
  assign \new_[4049]_  = ~\new_[5692]_  | ~\new_[11802]_  | ~\new_[4731]_ ;
  assign \new_[4050]_  = ~\new_[5290]_  | ~\new_[13283]_  | ~\new_[4738]_ ;
  assign \new_[4051]_  = ~\new_[4507]_  & ~\new_[7855]_  & ~\new_[4763]_ ;
  assign \new_[4052]_  = ~\new_[6168]_  | ~\new_[11082]_  | ~\new_[4728]_ ;
  assign \new_[4053]_  = ~\new_[9450]_  | ~\new_[5556]_  | ~\new_[4784]_  | ~\new_[8388]_ ;
  assign \new_[4054]_  = ~\new_[4447]_  | ~\new_[19452]_ ;
  assign \new_[4055]_  = ~\new_[10775]_  | ~\new_[4811]_  | ~\new_[5591]_  | ~\new_[8332]_ ;
  assign \new_[4056]_  = ~\new_[6173]_  | ~\new_[11152]_  | ~\new_[4737]_ ;
  assign \new_[4057]_  = ~\new_[8287]_  | ~\new_[5579]_  | ~\new_[4804]_  | ~\new_[7483]_ ;
  assign \new_[4058]_  = ~\new_[8289]_  | ~\new_[4806]_  | ~\new_[5583]_  | ~\new_[6043]_ ;
  assign \new_[4059]_  = ~\new_[5277]_  | ~\new_[4808]_  | ~\new_[6021]_  | ~\new_[5882]_ ;
  assign \new_[4060]_  = \new_[4446]_  & \new_[13166]_ ;
  assign \new_[4061]_  = ~\new_[8715]_  | ~\new_[8272]_  | ~\new_[7357]_  | ~\new_[4514]_ ;
  assign \new_[4062]_  = ~\new_[10874]_  | ~\new_[8288]_  | ~\new_[10768]_  | ~\new_[4513]_ ;
  assign \new_[4063]_  = ~\new_[926]_  & (~\new_[4508]_  | ~\new_[5080]_ );
  assign \new_[4064]_  = ~\new_[6421]_  | ~\new_[4441]_ ;
  assign \new_[4065]_  = (~\new_[4747]_  | ~\new_[2500]_ ) & (~\new_[6546]_  | ~\new_[17475]_ );
  assign \new_[4066]_  = ~\new_[9569]_  | ~\new_[4867]_  | ~\new_[6350]_  | ~\new_[4726]_ ;
  assign \new_[4067]_  = ~\new_[8696]_  | ~\new_[5196]_  | ~\new_[4745]_  | ~\new_[7201]_ ;
  assign \new_[4068]_  = ~\new_[20283]_  | (~\new_[4550]_  & ~\new_[5997]_ );
  assign \new_[4069]_  = ~\new_[19659]_  | (~\new_[4551]_  & ~\new_[9283]_ );
  assign \new_[4070]_  = ~\new_[19163]_  | (~\new_[4563]_  & ~\new_[9344]_ );
  assign \new_[4071]_  = ~\new_[19748]_  | (~\new_[4568]_  & ~\new_[20374]_ );
  assign \new_[4072]_  = ~\new_[18409]_  | (~\new_[4570]_  & ~\new_[8124]_ );
  assign \new_[4073]_  = ~\new_[4502]_  | ~\new_[19623]_ ;
  assign \new_[4074]_  = ~\new_[4491]_  | ~\new_[21267]_ ;
  assign \new_[4075]_  = ~\new_[4466]_  & ~\new_[5419]_ ;
  assign \new_[4076]_  = ~\new_[4890]_  | ~\new_[8222]_  | ~\new_[4602]_ ;
  assign \new_[4077]_  = ~\new_[4499]_  & ~\new_[6258]_ ;
  assign \new_[4078]_  = ~\new_[5166]_  | ~\new_[9467]_  | ~\new_[4972]_  | ~\new_[4653]_ ;
  assign \new_[4079]_  = ~\new_[20464]_  | (~\new_[4538]_  & ~\new_[5145]_ );
  assign \new_[4080]_  = \new_[4322]_  & \new_[19350]_ ;
  assign \new_[4081]_  = ~\new_[4577]_  & ~\new_[9078]_  & ~\new_[10075]_ ;
  assign \new_[4082]_  = ~\new_[18667]_  & (~\new_[4615]_  | ~\new_[8378]_ );
  assign \new_[4083]_  = ~\new_[18406]_  & (~\new_[4549]_  | ~\new_[6042]_ );
  assign \new_[4084]_  = ~\new_[18668]_  & (~\new_[4616]_  | ~\new_[8328]_ );
  assign \new_[4085]_  = ~\new_[19659]_  | (~\new_[4607]_  & ~\new_[5885]_ );
  assign \new_[4086]_  = ~\new_[4302]_  | ~\new_[984]_ ;
  assign \new_[4087]_  = ~\new_[19049]_  & (~\new_[4561]_  | ~\new_[7479]_ );
  assign \new_[4088]_  = ~\new_[4304]_  | ~\new_[19530]_ ;
  assign \new_[4089]_  = ~\new_[4305]_  | ~\new_[18583]_ ;
  assign \new_[4090]_  = ~\new_[19748]_  | (~\new_[4609]_  & ~\new_[5428]_ );
  assign \new_[4091]_  = ~\new_[19163]_  | (~\new_[4610]_  & ~\new_[5887]_ );
  assign \new_[4092]_  = ~\new_[4566]_  | ~\new_[5418]_  | ~\new_[4634]_ ;
  assign \new_[4093]_  = ~\new_[4569]_  | ~\new_[5035]_  | ~\new_[4842]_ ;
  assign \new_[4094]_  = ~\new_[12246]_  | ~\new_[4837]_  | ~\new_[4748]_  | ~\new_[5768]_ ;
  assign \new_[4095]_  = ~\new_[12209]_  | ~\new_[4838]_  | ~\new_[4750]_  | ~\new_[5339]_ ;
  assign \new_[4096]_  = ~\new_[9368]_  | ~\new_[14880]_  | ~\new_[4874]_  | ~\new_[4600]_ ;
  assign \new_[4097]_  = ~\new_[4500]_  & (~\new_[4945]_  | ~\new_[1879]_ );
  assign \new_[4098]_  = ~\new_[4473]_  & (~\new_[5629]_  | ~\new_[1879]_ );
  assign \new_[4099]_  = ~\new_[4475]_  & (~\new_[5246]_  | ~\new_[18791]_ );
  assign \new_[4100]_  = ~\new_[4501]_  & (~\new_[14246]_  | ~\new_[17669]_ );
  assign \new_[4101]_  = ~\new_[21008]_  | (~\new_[20758]_  & ~\new_[5073]_ );
  assign \new_[4102]_  = ~\new_[8286]_  | ~\new_[4863]_  | ~\new_[5442]_  | ~\new_[7478]_ ;
  assign \new_[4103]_  = ~\new_[21425]_  | (~\new_[4628]_  & ~\new_[5075]_ );
  assign \new_[4104]_  = ~\new_[4464]_  | ~\new_[5065]_ ;
  assign \new_[4105]_  = ~\new_[4455]_  | ~\new_[4956]_ ;
  assign \new_[4106]_  = (~\new_[4606]_  | ~\new_[19578]_ ) & (~\new_[12219]_  | ~\new_[19377]_ );
  assign \new_[4107]_  = ~\new_[4526]_  & ~\new_[7117]_  & ~\new_[5305]_ ;
  assign \new_[4108]_  = ~\new_[4527]_  & ~\new_[6379]_  & ~\new_[4978]_ ;
  assign \new_[4109]_  = ~\new_[4529]_  & ~\new_[5930]_  & ~\new_[5324]_ ;
  assign \new_[4110]_  = ~\new_[4697]_  & ~\new_[7168]_  & ~\new_[5326]_ ;
  assign \new_[4111]_  = ~\new_[4680]_  & ~\new_[5934]_  & ~\new_[4982]_ ;
  assign \new_[4112]_  = (~\new_[4619]_  | ~\new_[19049]_ ) & (~\new_[10938]_  | ~\new_[17796]_ );
  assign \new_[4113]_  = (~\new_[4620]_  | ~\new_[18942]_ ) & (~\new_[6854]_  | ~\new_[21630]_ );
  assign \new_[4114]_  = (~\new_[4621]_  | ~\new_[20513]_ ) & (~\new_[11003]_  | ~\new_[19798]_ );
  assign \new_[4115]_  = (~\new_[4622]_  | ~\new_[19257]_ ) & (~\new_[10983]_  | ~\new_[19491]_ );
  assign \new_[4116]_  = (~\new_[20381]_  | ~\new_[18004]_ ) & (~\new_[10644]_  | ~\new_[21559]_ );
  assign \new_[4117]_  = (~\new_[4623]_  | ~\new_[19748]_ ) & (~\new_[9298]_  | ~\new_[19243]_ );
  assign \new_[4118]_  = ~\new_[6139]_  | ~\new_[8115]_  | ~\new_[4338]_  | ~\new_[9828]_ ;
  assign \new_[4119]_  = ~\new_[5625]_  | ~\new_[8121]_  | ~\new_[4342]_  | ~\new_[10973]_ ;
  assign \new_[4120]_  = (~\new_[20706]_  | ~\new_[19246]_ ) & (~\new_[6581]_  | ~\new_[19276]_ );
  assign \new_[4121]_  = (~\new_[4608]_  | ~\new_[19300]_ ) & (~\new_[6587]_  | ~\new_[19236]_ );
  assign \new_[4122]_  = ~\new_[4260]_ ;
  assign \new_[4123]_  = ~\new_[15893]_  | (~\new_[5213]_  & ~\new_[4636]_ );
  assign \new_[4124]_  = ~\new_[6500]_  | ~\new_[4674]_  | ~\new_[6260]_ ;
  assign \new_[4125]_  = ~\new_[19751]_  & (~\new_[9077]_  | ~\new_[4660]_ );
  assign \new_[4126]_  = ~\new_[4367]_  | ~\new_[18198]_ ;
  assign \new_[4127]_  = ~\new_[4268]_ ;
  assign \new_[4128]_  = ~\new_[4386]_  | ~\new_[8499]_ ;
  assign \new_[4129]_  = ~\new_[4390]_  & (~\new_[6939]_  | ~\new_[18380]_ );
  assign \new_[4130]_  = ~\new_[21339]_  | ~\new_[8464]_ ;
  assign \new_[4131]_  = ~\new_[4395]_  | ~\new_[8517]_ ;
  assign \new_[4132]_  = \new_[4345]_  & \new_[19748]_ ;
  assign \new_[4133]_  = ~\new_[6620]_  | ~\new_[4401]_  | ~\new_[5238]_ ;
  assign \new_[4134]_  = ~\new_[6037]_  | ~\new_[4402]_  | ~\new_[5624]_ ;
  assign \new_[4135]_  = ~\new_[6044]_  | ~\new_[4403]_  | ~\new_[6910]_ ;
  assign \new_[4136]_  = ~\new_[4275]_ ;
  assign \new_[4137]_  = ~\new_[4524]_  & ~\new_[4404]_ ;
  assign \new_[4138]_  = ~\new_[4975]_  | ~\new_[4641]_  | ~\new_[8709]_ ;
  assign \new_[4139]_  = ~\new_[7837]_  & ~\new_[4327]_ ;
  assign \new_[4140]_  = ~\new_[4387]_  | ~\new_[18091]_ ;
  assign \new_[4141]_  = ~\new_[4379]_  | ~\new_[5618]_ ;
  assign \new_[4142]_  = ~\new_[8725]_  | ~\new_[11097]_  | ~\new_[5164]_  | ~\new_[4651]_ ;
  assign \new_[4143]_  = ~\new_[4380]_  | ~\new_[5228]_ ;
  assign \new_[4144]_  = ~\new_[4642]_  | ~\new_[5335]_  | ~\new_[8708]_ ;
  assign \new_[4145]_  = ~\new_[4393]_  | ~\new_[19530]_ ;
  assign \new_[4146]_  = ~\new_[5821]_  | (~\new_[4637]_  & ~\new_[954]_ );
  assign \new_[4147]_  = ~\new_[5385]_  | ~\new_[4373]_ ;
  assign \new_[4148]_  = ~\new_[8863]_  & ~\new_[4331]_ ;
  assign \new_[4149]_  = ~\new_[9062]_  & ~\new_[4332]_ ;
  assign \new_[4150]_  = ~\new_[4324]_  & (~\new_[10820]_  | ~\new_[18965]_ );
  assign \new_[4151]_  = ~\new_[4368]_  & (~\new_[4947]_  | ~\new_[19528]_ );
  assign \new_[4152]_  = ~\new_[6396]_  | ~\new_[4555]_  | ~\new_[5231]_ ;
  assign \new_[4153]_  = ~\new_[19512]_  | (~\new_[4854]_  & ~\new_[11063]_ );
  assign \new_[4154]_  = ~\new_[8993]_  & (~\new_[4951]_  | ~\new_[19787]_ );
  assign \new_[4155]_  = ~\new_[4530]_  & (~\new_[4943]_  | ~\new_[19659]_ );
  assign \new_[4156]_  = ~\new_[4531]_  & (~\new_[4944]_  | ~\new_[18004]_ );
  assign \new_[4157]_  = ~\new_[8900]_  | ~\new_[6647]_  | ~\new_[5358]_  | ~\new_[10016]_ ;
  assign \new_[4158]_  = (~\new_[4901]_  | ~\new_[19300]_ ) & (~\new_[11383]_  | ~\new_[15822]_ );
  assign \new_[4159]_  = ~\new_[8324]_  & ~\new_[4545]_ ;
  assign \new_[4160]_  = ~\new_[4525]_  & (~\new_[7670]_  | ~\new_[19507]_ );
  assign \new_[4161]_  = ~\new_[4594]_  & (~\new_[12577]_  | ~\new_[19377]_ );
  assign \new_[4162]_  = ~\new_[5401]_  | ~\new_[14195]_  | ~\new_[10093]_  | ~\new_[6159]_ ;
  assign \new_[4163]_  = ~\new_[5402]_  | ~\new_[13615]_  | ~\new_[10110]_  | ~\new_[5272]_ ;
  assign \new_[4164]_  = ~\new_[13265]_  | ~\new_[6224]_  | ~\new_[4686]_  | ~\new_[10149]_ ;
  assign \new_[4165]_  = ~\new_[4565]_  & (~\new_[6588]_  | ~\new_[19619]_ );
  assign \new_[4166]_  = ~\new_[13213]_  | ~\new_[7840]_  | ~\new_[5278]_  | ~\new_[5399]_ ;
  assign \new_[4167]_  = ~\new_[5410]_  | ~\new_[6629]_  | ~\new_[10639]_  | ~\new_[8749]_ ;
  assign \new_[4168]_  = (~\new_[4913]_  | ~\new_[19350]_ ) & (~\new_[5816]_  | ~\new_[19780]_ );
  assign \new_[4169]_  = ~\new_[5411]_  | ~\new_[7376]_  | ~\new_[12943]_  | ~\new_[9843]_ ;
  assign \new_[4170]_  = ~\new_[12743]_  | ~\new_[5663]_  | ~\new_[5031]_  | ~\new_[12391]_ ;
  assign \new_[4171]_  = ~\new_[6903]_  & ~\new_[4585]_ ;
  assign \new_[4172]_  = ~\new_[4809]_  | (~\new_[4915]_  & ~\new_[18988]_ );
  assign \new_[4173]_  = ~\new_[11107]_  | ~\new_[5388]_  | ~\new_[6631]_  | ~\new_[8874]_ ;
  assign \new_[4174]_  = ~\new_[10261]_  | ~\new_[5389]_  | ~\new_[7543]_  | ~\new_[7869]_ ;
  assign \new_[4175]_  = ~\new_[5252]_  | (~\new_[21169]_  & ~\new_[19504]_ );
  assign \new_[4176]_  = ~\new_[5441]_  | ~\new_[8774]_  | ~\new_[20781]_  | ~\new_[7675]_ ;
  assign \new_[4177]_  = ~\new_[5294]_  | (~\new_[4991]_  & ~\new_[19271]_ );
  assign \new_[4178]_  = ~\new_[4361]_ ;
  assign \new_[4179]_  = ~\new_[8639]_  | (~\new_[4998]_  & ~\new_[18757]_ );
  assign \new_[4180]_  = ~\new_[9717]_  | (~\new_[5000]_  & ~\new_[19561]_ );
  assign \new_[4181]_  = ~\new_[6782]_  | (~\new_[4996]_  & ~\new_[19578]_ );
  assign \new_[4182]_  = ~\new_[19133]_  | (~\new_[5027]_  & ~\new_[12750]_ );
  assign \new_[4183]_  = ~\new_[20941]_  | (~\new_[4987]_  & ~\new_[9138]_ );
  assign \new_[4184]_  = ~\new_[6556]_  | (~\new_[4992]_  & ~\new_[19509]_ );
  assign \new_[4185]_  = ~\new_[6568]_  | (~\new_[5003]_  & ~\new_[21417]_ );
  assign \new_[4186]_  = ~\new_[5474]_  | (~\new_[5004]_  & ~\new_[991]_ );
  assign \new_[4187]_  = ~\new_[5020]_  & ~\new_[7132]_  & ~\new_[13329]_ ;
  assign \new_[4188]_  = ~\new_[11636]_  | ~\new_[14892]_  | ~\new_[4966]_ ;
  assign \new_[4189]_  = ~\new_[5021]_  & ~\new_[7189]_  & ~\new_[12059]_ ;
  assign \new_[4190]_  = ~\new_[5023]_  & ~\new_[7195]_  & ~\new_[13333]_ ;
  assign \new_[4191]_  = ~\new_[4650]_  & (~\new_[5357]_  | ~\new_[19445]_ );
  assign \new_[4192]_  = ~\new_[20934]_  | (~\new_[6267]_  & ~\new_[19509]_ );
  assign \new_[4193]_  = ~\new_[4633]_  | (~\new_[5842]_  & ~\new_[19400]_ );
  assign \new_[4194]_  = (~\new_[5009]_  | ~\new_[1026]_ ) & (~\new_[6268]_  | ~\new_[19709]_ );
  assign \new_[4195]_  = (~\new_[20820]_  | ~\new_[19246]_ ) & (~\new_[12922]_  | ~\new_[17411]_ );
  assign \new_[4196]_  = ~\new_[7860]_  | ~\new_[4639]_ ;
  assign \new_[4197]_  = ~\new_[4963]_  & (~\new_[4990]_  | ~\new_[19334]_ );
  assign \new_[4198]_  = ~\new_[18808]_  | (~\new_[5039]_  & ~\new_[8307]_ );
  assign \new_[4199]_  = ~\new_[19246]_  | (~\new_[7554]_  & ~\new_[5042]_ );
  assign \new_[4200]_  = \new_[5047]_  & \new_[4693]_ ;
  assign \new_[4201]_  = ~\new_[4718]_  & ~\new_[6029]_ ;
  assign \new_[4202]_  = ~\new_[6504]_  | ~\new_[21408]_  | ~\new_[4713]_  | ~\new_[4797]_ ;
  assign \new_[4203]_  = ~\new_[7248]_  | ~\new_[11712]_  | ~\new_[4796]_  | ~\new_[4709]_ ;
  assign \new_[4204]_  = ~\new_[5707]_  | ~\new_[4957]_  | ~\new_[5063]_ ;
  assign \new_[4205]_  = ~\new_[5728]_  | ~\new_[5255]_  | ~\new_[5066]_ ;
  assign \new_[4206]_  = ~\new_[5734]_  | ~\new_[4960]_  | ~\new_[5067]_ ;
  assign \new_[4207]_  = ~\new_[6965]_  | ~\new_[5654]_  | ~\new_[5068]_ ;
  assign \new_[4208]_  = ~\new_[19002]_  | (~\new_[4756]_  & ~\new_[12760]_ );
  assign \new_[4209]_  = ~\new_[19041]_  | (~\new_[4757]_  & ~\new_[13345]_ );
  assign \new_[4210]_  = ~\new_[6914]_  | ~\new_[7012]_  | ~\new_[5071]_ ;
  assign \new_[4211]_  = ~\new_[19780]_  | (~\new_[4754]_  & ~\new_[7466]_ );
  assign \new_[4212]_  = (~\new_[4760]_  | ~\new_[18791]_ ) & (~\new_[16615]_  | ~\new_[11865]_ );
  assign \new_[4213]_  = ~\new_[19133]_  | (~\new_[4787]_  & ~\new_[8908]_ );
  assign \new_[4214]_  = ~\new_[19207]_  | (~\new_[4798]_  & ~\new_[8998]_ );
  assign \new_[4215]_  = ~\new_[19236]_  | (~\new_[4799]_  & ~\new_[10230]_ );
  assign \new_[4216]_  = \new_[4503]_  & \new_[19262]_ ;
  assign \new_[4217]_  = ~\new_[4719]_  | ~\new_[7010]_ ;
  assign \new_[4218]_  = ~\new_[7622]_  | ~\new_[5128]_  | ~\new_[7021]_  | ~\new_[5638]_ ;
  assign \new_[4219]_  = ~\new_[5137]_  | ~\new_[6616]_  | ~\new_[4865]_  | ~\new_[5282]_ ;
  assign \new_[4220]_  = ~\new_[5139]_  | ~\new_[7378]_  | ~\new_[6166]_  | ~\new_[5537]_ ;
  assign \new_[4221]_  = ~\new_[5175]_  | ~\new_[6655]_  | ~\new_[5689]_  | ~\new_[4893]_ ;
  assign \new_[4222]_  = ~\new_[5195]_  | ~\new_[7572]_  | ~\new_[5292]_  | ~\new_[5593]_ ;
  assign \new_[4223]_  = ~\new_[4509]_  | ~\new_[19442]_ ;
  assign \new_[4224]_  = ~\new_[5174]_  | ~\new_[5671]_  | ~\new_[5002]_  | ~\new_[10428]_ ;
  assign \new_[4225]_  = ~\new_[4505]_  | ~\new_[18612]_ ;
  assign \new_[4226]_  = ~\new_[4510]_  | ~\new_[19418]_ ;
  assign \new_[4227]_  = ~\new_[6014]_  | ~\new_[5182]_  | ~\new_[5275]_  | ~\new_[8058]_ ;
  assign \new_[4228]_  = ~\new_[4788]_  | ~\new_[5033]_  | ~\new_[5116]_ ;
  assign \new_[4229]_  = ~\new_[4810]_  | ~\new_[5036]_  | ~\new_[5119]_ ;
  assign \new_[4230]_  = ~\new_[4780]_  | ~\new_[5431]_  | ~\new_[7923]_ ;
  assign \new_[4231]_  = ~\new_[5709]_  | ~\new_[6151]_  | ~\new_[4554]_  | ~\new_[5307]_ ;
  assign \new_[4232]_  = ~\new_[10902]_  | ~\new_[5108]_  | ~\new_[5487]_  | ~\new_[5770]_ ;
  assign \new_[4233]_  = ~\new_[4794]_  | ~\new_[5440]_  | ~\new_[8974]_ ;
  assign \new_[4234]_  = ~\new_[4805]_  | ~\new_[6409]_  | ~\new_[9045]_ ;
  assign \new_[4235]_  = ~\new_[10766]_  | ~\new_[5125]_  | ~\new_[6354]_  | ~\new_[12135]_ ;
  assign \new_[4236]_  = ~\new_[9454]_  | ~\new_[5126]_  | ~\new_[5041]_  | ~\new_[12124]_ ;
  assign \new_[4237]_  = ~\new_[9440]_  | ~\new_[5127]_  | ~\new_[6356]_  | ~\new_[8345]_ ;
  assign \new_[4238]_  = ~\new_[8346]_  | ~\new_[5205]_  | ~\new_[8361]_  | ~\new_[7104]_ ;
  assign \new_[4239]_  = ~\new_[8267]_  | ~\new_[5129]_  | ~\new_[5446]_  | ~\new_[10811]_ ;
  assign \new_[4240]_  = ~\new_[4749]_  & (~\new_[4946]_  | ~\new_[18668]_ );
  assign \new_[4241]_  = ~\new_[4732]_  & (~\new_[5247]_  | ~\new_[1878]_ );
  assign \new_[4242]_  = ~\new_[5102]_  | ~\new_[9543]_  | ~\new_[9542]_  | ~\new_[12596]_ ;
  assign \new_[4243]_  = ~\new_[12133]_  | ~\new_[7202]_  | ~\new_[4831]_ ;
  assign \new_[4244]_  = ~\new_[19736]_  & (~\new_[4835]_  | ~\new_[5407]_ );
  assign \new_[4245]_  = ~\new_[9460]_  | ~\new_[5134]_  | ~\new_[5951]_  | ~\new_[6722]_ ;
  assign \new_[4246]_  = ~\new_[10771]_  | ~\new_[5131]_  | ~\new_[7162]_  | ~\new_[6665]_ ;
  assign \new_[4247]_  = ~\new_[8285]_  | ~\new_[7472]_  | ~\new_[5118]_  | ~\new_[10848]_ ;
  assign \new_[4248]_  = ~\new_[19812]_  | (~\new_[4836]_  & ~\new_[5074]_ );
  assign \new_[4249]_  = ~\new_[10773]_  | ~\new_[5132]_  | ~\new_[7192]_  | ~\new_[9665]_ ;
  assign \new_[4250]_  = ~\new_[8293]_  | ~\new_[5133]_  | ~\new_[6438]_  | ~\new_[6709]_ ;
  assign \new_[4251]_  = ~\new_[5564]_  | ~\new_[5403]_  | ~\new_[5678]_  | ~\new_[11159]_ ;
  assign \new_[4252]_  = (~\new_[4828]_  | ~\new_[19780]_ ) & (~\new_[9960]_  | ~\new_[17475]_ );
  assign \new_[4253]_  = (~\new_[4832]_  | ~\new_[19659]_ ) & (~\new_[11954]_  | ~\new_[19005]_ );
  assign \new_[4254]_  = (~\new_[4833]_  | ~\new_[20645]_ ) & (~\new_[10365]_  | ~\new_[19384]_ );
  assign \new_[4255]_  = (~\new_[4834]_  | ~\new_[19787]_ ) & (~\new_[11042]_  | ~\new_[17668]_ );
  assign \new_[4256]_  = ~\new_[4720]_  | ~\new_[5268]_ ;
  assign \new_[4257]_  = ~\new_[6471]_  & ~\new_[4536]_ ;
  assign \new_[4258]_  = ~\new_[9787]_  & ~\new_[4575]_ ;
  assign \new_[4259]_  = ~\new_[6480]_  & ~\new_[4539]_ ;
  assign \new_[4260]_  = ~\new_[5200]_  | ~\new_[5962]_  | ~\new_[5016]_ ;
  assign \new_[4261]_  = ~\new_[4576]_  & (~\new_[10707]_  | ~\new_[18965]_ );
  assign \new_[4262]_  = ~\new_[4920]_  | ~\new_[6759]_  | ~\new_[6003]_ ;
  assign \new_[4263]_  = ~\new_[6535]_  | ~\new_[4934]_  | ~\new_[5826]_ ;
  assign \new_[4264]_  = ~\new_[4596]_  | ~\new_[19599]_ ;
  assign \new_[4265]_  = ~\new_[4597]_  | ~\new_[19337]_ ;
  assign \new_[4266]_  = ~\new_[20789]_  | (~\new_[4896]_  & ~\new_[10241]_ );
  assign \new_[4267]_  = ~\new_[19236]_  | (~\new_[4897]_  & ~\new_[7925]_ );
  assign \new_[4268]_  = ~\new_[4574]_  | ~\new_[18612]_ ;
  assign \new_[4269]_  = ~\new_[19257]_  | (~\new_[4952]_  & ~\new_[10369]_ );
  assign \new_[4270]_  = ~\new_[19512]_  | (~\new_[4866]_  & ~\new_[5528]_ );
  assign \new_[4271]_  = ~\new_[19022]_  | (~\new_[4875]_  & ~\new_[5530]_ );
  assign \new_[4272]_  = ~\new_[4626]_  & ~\new_[4765]_ ;
  assign \new_[4273]_  = ~\new_[4840]_  | ~\new_[4766]_  | ~\new_[5221]_ ;
  assign \new_[4274]_  = ~\new_[4630]_  & ~\new_[4767]_ ;
  assign \new_[4275]_  = ~\new_[19032]_  | (~\new_[4929]_  & ~\new_[8294]_ );
  assign \new_[4276]_  = ~\new_[6745]_  | ~\new_[8849]_  | ~\new_[4645]_  | ~\new_[5295]_ ;
  assign \new_[4277]_  = ~\new_[960]_  | (~\new_[4878]_  & ~\new_[8931]_ );
  assign \new_[4278]_  = ~\new_[4883]_  & ~\new_[7023]_  & ~\new_[5271]_ ;
  assign \new_[4279]_  = ~\new_[8722]_  | ~\new_[8899]_  | ~\new_[5159]_  | ~\new_[4884]_ ;
  assign \new_[4280]_  = ~\new_[5820]_  | (~\new_[4849]_  & ~\new_[19442]_ );
  assign \new_[4281]_  = (~\new_[4887]_  | ~\new_[19780]_ ) & (~\new_[13503]_  | ~\new_[18076]_ );
  assign \new_[4282]_  = (~\new_[4889]_  | ~\new_[19277]_ ) & (~\new_[10721]_  | ~\new_[19625]_ );
  assign \new_[4283]_  = ~\new_[8940]_  & ~\new_[4522]_ ;
  assign \new_[4284]_  = ~\new_[10194]_  & ~\new_[4523]_ ;
  assign \new_[4285]_  = ~\new_[4900]_  & ~\new_[7025]_  & ~\new_[5664]_ ;
  assign \new_[4286]_  = ~\new_[5379]_  | ~\new_[10601]_  | ~\new_[11630]_  | ~\new_[5810]_ ;
  assign \new_[4287]_  = ~\new_[4518]_  & (~\new_[9582]_  | ~\new_[18998]_ );
  assign \new_[4288]_  = ~\new_[4895]_  | ~\new_[5034]_  | ~\new_[5273]_ ;
  assign \new_[4289]_  = ~\new_[4517]_  & (~\new_[8606]_  | ~\new_[18187]_ );
  assign \new_[4290]_  = ~\new_[5861]_  | ~\new_[13652]_  | ~\new_[4685]_  | ~\new_[4965]_ ;
  assign \new_[4291]_  = ~\new_[18791]_  & (~\new_[4871]_  | ~\new_[8264]_ );
  assign \new_[4292]_  = ~\new_[6952]_  | ~\new_[5300]_  | ~\new_[8902]_  | ~\new_[9817]_ ;
  assign \new_[4293]_  = ~\new_[4595]_  & ~\new_[5705]_ ;
  assign \new_[4294]_  = ~\new_[5794]_  & (~\new_[4917]_  | ~\new_[19717]_ );
  assign \new_[4295]_  = ~\new_[5359]_  & (~\new_[4918]_  | ~\new_[19561]_ );
  assign \new_[4296]_  = ~\new_[5726]_  | ~\new_[5727]_  | ~\new_[12977]_  | ~\new_[11056]_ ;
  assign \new_[4297]_  = ~\new_[6370]_  | ~\new_[4782]_  | ~\new_[5226]_ ;
  assign \new_[4298]_  = ~\new_[8879]_  & (~\new_[5244]_  | ~\new_[19271]_ );
  assign \new_[4299]_  = ~\new_[8834]_  & (~\new_[5245]_  | ~\new_[19257]_ );
  assign \new_[4300]_  = (~\new_[5219]_  | ~\new_[991]_ ) & (~\new_[5825]_  | ~\new_[21267]_ );
  assign \new_[4301]_  = ~\new_[7990]_  | ~\new_[5670]_  | ~\new_[5169]_  | ~\new_[8435]_ ;
  assign \new_[4302]_  = ~\new_[7976]_  | ~\new_[5795]_  | ~\new_[6644]_  | ~\new_[8948]_ ;
  assign \new_[4303]_  = ~\new_[6046]_  | ~\new_[5804]_  | ~\new_[6870]_  | ~\new_[8794]_ ;
  assign \new_[4304]_  = ~\new_[9074]_  | ~\new_[6048]_  | ~\new_[5805]_  | ~\new_[10139]_ ;
  assign \new_[4305]_  = ~\new_[8901]_  | ~\new_[5489]_  | ~\new_[5806]_  | ~\new_[8980]_ ;
  assign \new_[4306]_  = ~\new_[8037]_  | ~\new_[5639]_  | ~\new_[5784]_  | ~\new_[7777]_ ;
  assign \new_[4307]_  = ~\new_[4768]_  & (~\new_[7611]_  | ~\new_[19045]_ );
  assign \new_[4308]_  = ~\new_[12764]_  | ~\new_[6981]_  | ~\new_[5640]_  | ~\new_[14322]_ ;
  assign \new_[4309]_  = ~\new_[10523]_  | ~\new_[5641]_  | ~\new_[6982]_  | ~\new_[14173]_ ;
  assign \new_[4310]_  = ~\new_[8032]_  | ~\new_[5642]_  | ~\new_[5787]_  | ~\new_[8747]_ ;
  assign \new_[4311]_  = ~\new_[6701]_  & ~\new_[4786]_ ;
  assign \new_[4312]_  = ~\new_[4769]_  & (~\new_[7615]_  | ~\new_[19177]_ );
  assign \new_[4313]_  = ~\new_[7431]_  & ~\new_[4791]_ ;
  assign \new_[4314]_  = ~\new_[13888]_  | ~\new_[6998]_  | ~\new_[5648]_  | ~\new_[14251]_ ;
  assign \new_[4315]_  = ~\new_[9276]_  | ~\new_[5658]_  | ~\new_[6985]_  | ~\new_[13035]_ ;
  assign \new_[4316]_  = ~\new_[8036]_  | ~\new_[5649]_  | ~\new_[5798]_  | ~\new_[8768]_ ;
  assign \new_[4317]_  = ~\new_[11687]_  | ~\new_[6993]_  | ~\new_[5650]_  | ~\new_[15306]_ ;
  assign \new_[4318]_  = ~\new_[6997]_  | ~\new_[5657]_  | ~\new_[12770]_  | ~\new_[15195]_ ;
  assign \new_[4319]_  = ~\new_[5635]_  & ~\new_[4777]_ ;
  assign \new_[4320]_  = ~\new_[5257]_  & ~\new_[4801]_ ;
  assign \new_[4321]_  = (~\new_[5208]_  | ~\new_[19550]_ ) & (~\new_[5153]_  | ~\new_[15893]_ );
  assign \new_[4322]_  = ~\new_[11348]_  | ~\new_[5829]_  | ~\new_[8405]_  | ~\new_[11064]_ ;
  assign \new_[4323]_  = ~\new_[19659]_  | (~\new_[5343]_  & ~\new_[8930]_ );
  assign \new_[4324]_  = ~\new_[4997]_  | (~\new_[5302]_  & ~\new_[19070]_ );
  assign \new_[4325]_  = ~\new_[19748]_  | (~\new_[5345]_  & ~\new_[6894]_ );
  assign \new_[4326]_  = ~\new_[19170]_  | (~\new_[5346]_  & ~\new_[8898]_ );
  assign \new_[4327]_  = ~\new_[19334]_  & (~\new_[8613]_  | ~\new_[5408]_ );
  assign \new_[4328]_  = ~\new_[4519]_ ;
  assign \new_[4329]_  = ~\new_[4520]_ ;
  assign \new_[4330]_  = ~\new_[4521]_ ;
  assign \new_[4331]_  = ~\new_[19284]_  & (~\new_[9262]_  | ~\new_[5413]_ );
  assign \new_[4332]_  = ~\new_[19022]_  & (~\new_[9693]_  | ~\new_[5414]_ );
  assign \new_[4333]_  = ~\new_[5323]_  & ~\new_[9096]_  & ~\new_[9621]_ ;
  assign \new_[4334]_  = (~\new_[5330]_  | ~\new_[18798]_ ) & (~\new_[7949]_  | ~\new_[19559]_ );
  assign \new_[4335]_  = (~\new_[5331]_  | ~\new_[19102]_ ) & (~\new_[6905]_  | ~\new_[19382]_ );
  assign \new_[4336]_  = ~\new_[5900]_  | ~\new_[10887]_  | ~\new_[9437]_  | ~\new_[8033]_ ;
  assign \new_[4337]_  = ~\new_[4540]_ ;
  assign \new_[4338]_  = ~\new_[4880]_  | ~\new_[1879]_ ;
  assign \new_[4339]_  = ~\new_[19748]_  & (~\new_[5299]_  | ~\new_[9304]_ );
  assign \new_[4340]_  = ~\new_[8600]_  | ~\new_[5304]_  | ~\new_[6956]_ ;
  assign \new_[4341]_  = ~\new_[4885]_  | ~\new_[984]_ ;
  assign \new_[4342]_  = ~\new_[4888]_  | ~\new_[19195]_ ;
  assign \new_[4343]_  = ~\new_[5914]_  | ~\new_[9941]_  | ~\new_[5482]_  | ~\new_[7657]_ ;
  assign \new_[4344]_  = ~\new_[5310]_  & ~\new_[9152]_  & ~\new_[6832]_ ;
  assign \new_[4345]_  = ~\new_[5907]_  | ~\new_[9860]_  | ~\new_[6024]_  | ~\new_[7659]_ ;
  assign \new_[4346]_  = ~\new_[5312]_  | ~\new_[6960]_  | ~\new_[10884]_ ;
  assign \new_[4347]_  = ~\new_[4556]_ ;
  assign \new_[4348]_  = ~\new_[4894]_  | ~\new_[19418]_ ;
  assign \new_[4349]_  = ~\new_[5325]_  | ~\new_[8514]_  | ~\new_[6962]_ ;
  assign \new_[4350]_  = ~\new_[4562]_ ;
  assign \new_[4351]_  = ~\new_[5327]_  | ~\new_[7500]_  | ~\new_[6963]_ ;
  assign \new_[4352]_  = ~\new_[4905]_  | ~\new_[19300]_ ;
  assign \new_[4353]_  = ~\new_[5332]_  & ~\new_[21387]_  & ~\new_[7734]_ ;
  assign \new_[4354]_  = ~\new_[5018]_  | ~\new_[4930]_ ;
  assign \new_[4355]_  = ~\new_[19032]_  & (~\new_[5336]_  | ~\new_[21195]_ );
  assign \new_[4356]_  = ~\new_[4933]_  | ~\new_[5767]_ ;
  assign \new_[4357]_  = ~\new_[4844]_  & ~\new_[5400]_ ;
  assign \new_[4358]_  = ~\new_[7558]_  | (~\new_[5393]_  & ~\new_[19350]_ );
  assign \new_[4359]_  = ~\new_[4852]_  & ~\new_[5404]_ ;
  assign \new_[4360]_  = (~\new_[5365]_  | ~\new_[984]_ ) & (~\new_[6502]_  | ~\new_[15963]_ );
  assign \new_[4361]_  = ~\new_[7974]_  | (~\new_[5394]_  & ~\new_[19334]_ );
  assign \new_[4362]_  = ~\new_[4909]_  & (~\new_[11336]_  | ~\new_[17285]_ );
  assign \new_[4363]_  = ~\new_[4911]_  & (~\new_[10105]_  | ~\new_[17381]_ );
  assign \new_[4364]_  = ~\new_[4860]_  & ~\new_[5029]_ ;
  assign \new_[4365]_  = ~\new_[7913]_  | ~\new_[5865]_  | ~\new_[4961]_  | ~\new_[12469]_ ;
  assign \new_[4366]_  = ~\new_[7893]_  | ~\new_[5866]_  | ~\new_[4962]_  | ~\new_[21615]_ ;
  assign \new_[4367]_  = \new_[6002]_  | \new_[7847]_  | \new_[7868]_  | \new_[13061]_ ;
  assign \new_[4368]_  = ~\new_[2500]_  & (~\new_[5309]_  | ~\new_[8288]_ );
  assign \new_[4369]_  = ~\new_[4876]_  | ~\new_[19659]_ ;
  assign \new_[4370]_  = ~\new_[20941]_  | (~\new_[5396]_  & ~\new_[12530]_ );
  assign \new_[4371]_  = ~\new_[4891]_  | ~\new_[19748]_ ;
  assign \new_[4372]_  = ~\new_[19257]_  | (~\new_[5397]_  & ~\new_[13792]_ );
  assign \new_[4373]_  = ~\new_[18942]_  | (~\new_[5398]_  & ~\new_[13575]_ );
  assign \new_[4374]_  = ~\new_[4859]_  | (~\new_[5378]_  & ~\new_[19525]_ );
  assign \new_[4375]_  = ~\new_[5179]_  | ~\new_[4919]_ ;
  assign \new_[4376]_  = ~\new_[5859]_  | ~\new_[13847]_  | ~\new_[15668]_  | ~\new_[11097]_ ;
  assign \new_[4377]_  = ~\new_[12176]_  | ~\new_[5953]_  | ~\new_[6725]_  | ~\new_[15043]_ ;
  assign \new_[4378]_  = ~\new_[5455]_  & ~\new_[4845]_ ;
  assign \new_[4379]_  = \new_[5786]_  ? \new_[19578]_  : \new_[5356]_ ;
  assign \new_[4380]_  = \new_[5360]_  ? \new_[19561]_  : \new_[5375]_ ;
  assign \new_[4381]_  = ~\new_[4841]_  | (~\new_[5841]_  & ~\new_[19512]_ );
  assign \new_[4382]_  = (~\new_[5370]_  | ~\new_[19433]_ ) & (~\new_[7011]_  | ~\new_[19696]_ );
  assign \new_[4383]_  = (~\new_[5371]_  | ~\new_[1033]_ ) & (~\new_[7002]_  | ~\new_[19157]_ );
  assign \new_[4384]_  = (~\new_[5373]_  | ~\new_[18983]_ ) & (~\new_[5843]_  | ~\new_[19257]_ );
  assign \new_[4385]_  = (~\new_[5361]_  | ~\new_[960]_ ) & (~\new_[5395]_  | ~\new_[19271]_ );
  assign \new_[4386]_  = (~\new_[5416]_  | ~\new_[18649]_ ) & (~\new_[12851]_  | ~\new_[17470]_ );
  assign \new_[4387]_  = ~\new_[10941]_  | ~\new_[5908]_  | ~\new_[8375]_  | ~\new_[9823]_ ;
  assign \new_[4388]_  = ~\new_[4617]_ ;
  assign \new_[4389]_  = ~\new_[8419]_  & ~\new_[4886]_ ;
  assign \new_[4390]_  = ~\new_[7880]_  | ~\new_[4851]_ ;
  assign \new_[4391]_  = ~\new_[9930]_  | ~\new_[8531]_  | ~\new_[5867]_  | ~\new_[10513]_ ;
  assign \new_[4392]_  = ~\new_[7863]_  | ~\new_[4847]_ ;
  assign \new_[4393]_  = ~\new_[9918]_  | ~\new_[5925]_  | ~\new_[8483]_  | ~\new_[9869]_ ;
  assign \new_[4394]_  = ~\new_[7919]_  | ~\new_[4855]_ ;
  assign \new_[4395]_  = (~\new_[5415]_  | ~\new_[19433]_ ) & (~\new_[12841]_  | ~\new_[16632]_ );
  assign \new_[4396]_  = ~\new_[7494]_  & ~\new_[4902]_ ;
  assign \new_[4397]_  = ~\new_[5531]_  | ~\new_[7031]_  | ~\new_[8589]_  | ~\new_[11491]_ ;
  assign \new_[4398]_  = ~\new_[5214]_  & (~\new_[5457]_  | ~\new_[19032]_ );
  assign \new_[4399]_  = ~\new_[4923]_  & (~\new_[5991]_  | ~\new_[19236]_ );
  assign \new_[4400]_  = ~\new_[4924]_  & (~\new_[5467]_  | ~\new_[19051]_ );
  assign \new_[4401]_  = ~\new_[5270]_  & ~\new_[4882]_ ;
  assign \new_[4402]_  = ~\new_[5274]_  & ~\new_[4899]_ ;
  assign \new_[4403]_  = ~\new_[5276]_  & ~\new_[4903]_ ;
  assign \new_[4404]_  = ~\new_[5224]_  | (~\new_[5383]_  & ~\new_[19529]_ );
  assign \new_[4405]_  = ~\new_[5921]_  | ~\new_[5459]_  | ~\new_[5473]_ ;
  assign \new_[4406]_  = ~\new_[8116]_  & ~\new_[4977]_ ;
  assign \new_[4407]_  = ~\new_[4989]_  | ~\new_[19070]_ ;
  assign \new_[4408]_  = ~\new_[4655]_ ;
  assign \new_[4409]_  = ~\new_[5026]_  & ~\new_[14497]_ ;
  assign \new_[4410]_  = ~\new_[20982]_  | (~\new_[5432]_  & ~\new_[12579]_ );
  assign \new_[4411]_  = ~\new_[8853]_  | ~\new_[9284]_  | ~\new_[5941]_  | ~\new_[7534]_ ;
  assign \new_[4412]_  = ~\new_[18649]_  | (~\new_[7567]_  & ~\new_[5449]_ );
  assign \new_[4413]_  = ~\new_[5028]_  & ~\new_[14624]_ ;
  assign \new_[4414]_  = ~\new_[19507]_  & (~\new_[5471]_  | ~\new_[13909]_ );
  assign \new_[4415]_  = \new_[5912]_  & \new_[4979]_ ;
  assign \new_[4416]_  = ~\new_[8608]_  | ~\new_[5437]_  | ~\new_[8132]_ ;
  assign \new_[4417]_  = ~\new_[4980]_  & (~\new_[8966]_  | ~\new_[19448]_ );
  assign \new_[4418]_  = ~\new_[19045]_  & (~\new_[5468]_  | ~\new_[13886]_ );
  assign \new_[4419]_  = ~\new_[10323]_  | ~\new_[5507]_  | ~\new_[7530]_  | ~\new_[13245]_ ;
  assign \new_[4420]_  = ~\new_[5053]_  & ~\new_[6650]_ ;
  assign \new_[4421]_  = ~\new_[4698]_ ;
  assign \new_[4422]_  = (~\new_[5485]_  | ~\new_[1879]_ ) & (~\new_[9392]_  | ~\new_[19377]_ );
  assign \new_[4423]_  = (~\new_[5072]_  | ~\new_[19528]_ ) & (~\new_[17015]_  | ~\new_[11788]_ );
  assign \new_[4424]_  = ~\new_[5062]_  | ~\new_[19694]_ ;
  assign \new_[4425]_  = ~\new_[20941]_  | (~\new_[5083]_  & ~\new_[8843]_ );
  assign \new_[4426]_  = ~\new_[5070]_  | ~\new_[19051]_ ;
  assign \new_[4427]_  = ~\new_[7650]_  | ~\new_[6865]_  | ~\new_[7022]_  | ~\new_[5261]_ ;
  assign \new_[4428]_  = ~\new_[9767]_  | ~\new_[5534]_  | ~\new_[6278]_  | ~\new_[5262]_ ;
  assign \new_[4429]_  = ~\new_[8238]_  | ~\new_[5617]_  | ~\new_[5685]_  | ~\new_[6127]_ ;
  assign \new_[4430]_  = (~\new_[5084]_  | ~\new_[19780]_ ) & (~\new_[12425]_  | ~\new_[18076]_ );
  assign \new_[4431]_  = ~\new_[5060]_  & (~\new_[14261]_  | ~\new_[19115]_ );
  assign \new_[4432]_  = ~\new_[4753]_  | ~\new_[19157]_ ;
  assign \new_[4433]_  = \new_[4761]_  & \new_[18280]_ ;
  assign \new_[4434]_  = ~\new_[5599]_  | ~\new_[5667]_  | ~\new_[5015]_  | ~\new_[10407]_ ;
  assign \new_[4435]_  = ~\new_[5647]_  | ~\new_[4762]_  | ~\new_[5715]_ ;
  assign \new_[4436]_  = ~\new_[5089]_  & ~\new_[5443]_  & ~\new_[5744]_ ;
  assign \new_[4437]_  = ~\new_[8351]_  | ~\new_[8106]_  | ~\new_[5099]_ ;
  assign \new_[4438]_  = ~\new_[10799]_  | ~\new_[7207]_  | ~\new_[5101]_ ;
  assign \new_[4439]_  = ~\new_[10774]_  | ~\new_[5535]_  | ~\new_[6448]_  | ~\new_[9633]_ ;
  assign \new_[4440]_  = ~\new_[8283]_  | ~\new_[5527]_  | ~\new_[7157]_  | ~\new_[10846]_ ;
  assign \new_[4441]_  = ~\new_[20464]_  | (~\new_[5106]_  & ~\new_[5076]_ );
  assign \new_[4442]_  = ~\new_[10912]_  | ~\new_[6117]_  | ~\new_[4873]_  | ~\new_[5086]_ ;
  assign \new_[4443]_  = (~\new_[19640]_  | ~\new_[5103]_ ) & (~\new_[11973]_  | ~\new_[19237]_ );
  assign \new_[4444]_  = ~\new_[5077]_  & ~\new_[7174]_  & ~\new_[5743]_ ;
  assign \new_[4445]_  = ~\new_[9083]_  & (~\new_[5104]_  | ~\new_[21418]_ );
  assign \new_[4446]_  = (~\new_[5105]_  | ~\new_[19599]_ ) & (~\new_[10670]_  | ~\new_[20701]_ );
  assign \new_[4447]_  = ~\new_[6140]_  | ~\new_[8131]_  | ~\new_[4790]_  | ~\new_[9855]_ ;
  assign \new_[4448]_  = (~\new_[5096]_  | ~\new_[18763]_ ) & (~\new_[6578]_  | ~\new_[19740]_ );
  assign \new_[4449]_  = (~\new_[999]_  | ~\new_[5097]_ ) & (~\new_[6585]_  | ~\new_[19702]_ );
  assign \new_[4450]_  = ~\new_[4827]_  | ~\new_[19567]_ ;
  assign \new_[4451]_  = ~\new_[5156]_  & ~\new_[8735]_  & ~\new_[6757]_ ;
  assign \new_[4452]_  = ~\new_[4816]_  | ~\new_[20941]_ ;
  assign \new_[4453]_  = ~\new_[4817]_  | ~\new_[19271]_ ;
  assign \new_[4454]_  = ~\new_[19002]_  | (~\new_[5144]_  & ~\new_[10056]_ );
  assign \new_[4455]_  = ~\new_[4818]_  | ~\new_[19659]_ ;
  assign \new_[4456]_  = ~\new_[4822]_  | ~\new_[19709]_ ;
  assign \new_[4457]_  = ~\new_[19041]_  | (~\new_[5168]_  & ~\new_[10354]_ );
  assign \new_[4458]_  = ~\new_[4819]_  | ~\new_[19448]_ ;
  assign \new_[4459]_  = ~\new_[4820]_  | ~\new_[19170]_ ;
  assign \new_[4460]_  = ~\new_[4821]_  | ~\new_[19207]_ ;
  assign \new_[4461]_  = ~\new_[4823]_  | ~\new_[19257]_ ;
  assign \new_[4462]_  = ~\new_[4781]_  | ~\new_[19041]_ ;
  assign \new_[4463]_  = ~\new_[19170]_  | (~\new_[5249]_  & ~\new_[8959]_ );
  assign \new_[4464]_  = ~\new_[4795]_  | ~\new_[19157]_ ;
  assign \new_[4465]_  = ~\new_[19787]_  | (~\new_[5250]_  & ~\new_[9116]_ );
  assign \new_[4466]_  = ~\new_[4771]_  | (~\new_[6493]_  & ~\new_[1878]_ );
  assign \new_[4467]_  = ~\new_[5115]_  | ~\new_[8350]_  | ~\new_[7362]_ ;
  assign \new_[4468]_  = ~\new_[5117]_  | ~\new_[7552]_  | ~\new_[10765]_ ;
  assign \new_[4469]_  = ~\new_[19442]_  | (~\new_[5569]_  & ~\new_[5121]_ );
  assign \new_[4470]_  = (~\new_[5138]_  | ~\new_[19659]_ ) & (~\new_[10723]_  | ~\new_[18863]_ );
  assign \new_[4471]_  = ~\new_[4824]_  | ~\new_[19528]_ ;
  assign \new_[4472]_  = ~\new_[19284]_  | (~\new_[5149]_  & ~\new_[10078]_ );
  assign \new_[4473]_  = \new_[5353]_  | \new_[4825]_ ;
  assign \new_[4474]_  = ~\new_[18988]_  | (~\new_[5151]_  & ~\new_[12331]_ );
  assign \new_[4475]_  = \new_[5354]_  | \new_[4826]_ ;
  assign \new_[4476]_  = (~\new_[5154]_  | ~\new_[19748]_ ) & (~\new_[10727]_  | ~\new_[17960]_ );
  assign \new_[4477]_  = ~\new_[19318]_  | (~\new_[5215]_  & ~\new_[9420]_ );
  assign \new_[4478]_  = ~\new_[1878]_  | (~\new_[5158]_  & ~\new_[11173]_ );
  assign \new_[4479]_  = ~\new_[4829]_  | ~\new_[984]_ ;
  assign \new_[4480]_  = ~\new_[960]_  | (~\new_[5161]_  & ~\new_[6492]_ );
  assign \new_[4481]_  = ~\new_[19529]_  | (~\new_[5163]_  & ~\new_[10130]_ );
  assign \new_[4482]_  = ~\new_[19509]_  | (~\new_[5167]_  & ~\new_[7260]_ );
  assign \new_[4483]_  = ~\new_[8982]_  & ~\new_[4764]_ ;
  assign \new_[4484]_  = ~\new_[954]_  | (~\new_[5176]_  & ~\new_[7274]_ );
  assign \new_[4485]_  = ~\new_[18983]_  | (~\new_[5178]_  & ~\new_[8197]_ );
  assign \new_[4486]_  = ~\new_[959]_  | (~\new_[20898]_  & ~\new_[9048]_ );
  assign \new_[4487]_  = ~\new_[19467]_  | (~\new_[5181]_  & ~\new_[9384]_ );
  assign \new_[4488]_  = ~\new_[6087]_  | ~\new_[9126]_  | ~\new_[5183]_  | ~\new_[5328]_ ;
  assign \new_[4489]_  = ~\new_[1026]_  | (~\new_[5184]_  & ~\new_[7278]_ );
  assign \new_[4490]_  = ~\new_[5823]_  | (~\new_[5123]_  & ~\new_[19517]_ );
  assign \new_[4491]_  = ~\new_[5186]_  | ~\new_[6047]_  | ~\new_[5739]_ ;
  assign \new_[4492]_  = ~\new_[9747]_  | ~\new_[5234]_  | ~\new_[5740]_  | ~\new_[9020]_ ;
  assign \new_[4493]_  = ~\new_[959]_  | (~\new_[5187]_  & ~\new_[7279]_ );
  assign \new_[4494]_  = ~\new_[19529]_  | (~\new_[5191]_  & ~\new_[7283]_ );
  assign \new_[4495]_  = ~\new_[19318]_  | (~\new_[5150]_  & ~\new_[14168]_ );
  assign \new_[4496]_  = ~\new_[20152]_  & (~\new_[5225]_  | ~\new_[8602]_ );
  assign \new_[4497]_  = \new_[5862]_  | \new_[12876]_  | \new_[10070]_  | \new_[9288]_ ;
  assign \new_[4498]_  = \new_[5863]_  | \new_[13449]_  | \new_[10196]_  | \new_[21591]_ ;
  assign \new_[4499]_  = ~\new_[19528]_  & (~\new_[6317]_  | ~\new_[5206]_ );
  assign \new_[4500]_  = ~\new_[18667]_  & (~\new_[5148]_  | ~\new_[9439]_ );
  assign \new_[4501]_  = ~\new_[19070]_  & (~\new_[6336]_  | ~\new_[5209]_ );
  assign \new_[4502]_  = ~\new_[7792]_  | ~\new_[5679]_  | ~\new_[11926]_  | ~\new_[9882]_ ;
  assign \new_[4503]_  = ~\new_[6205]_  | ~\new_[6206]_  | ~\new_[10206]_  | ~\new_[9993]_ ;
  assign \new_[4504]_  = ~\new_[5090]_  | ~\new_[19003]_ ;
  assign \new_[4505]_  = ~\new_[6162]_  | ~\new_[13723]_  | ~\new_[6310]_  | ~\new_[14146]_ ;
  assign \new_[4506]_  = ~\new_[20844]_  | ~\new_[5109]_  | ~\new_[5610]_ ;
  assign \new_[4507]_  = ~\new_[8629]_  | ~\new_[7069]_  | ~\new_[6204]_  | ~\new_[6766]_ ;
  assign \new_[4508]_  = ~\new_[5217]_  & (~\new_[6136]_  | ~\new_[20152]_ );
  assign \new_[4509]_  = ~\new_[6873]_  | ~\new_[6239]_  | ~\new_[6638]_  | ~\new_[7972]_ ;
  assign \new_[4510]_  = ~\new_[6896]_  | ~\new_[6244]_  | ~\new_[5488]_  | ~\new_[8829]_ ;
  assign \new_[4511]_  = ~\new_[11702]_  | ~\new_[6155]_  | ~\new_[5809]_  | ~\new_[14158]_ ;
  assign \new_[4512]_  = ~\new_[4759]_ ;
  assign \new_[4513]_  = (~\new_[5607]_  | ~\new_[19780]_ ) & (~\new_[5563]_  | ~\new_[19350]_ );
  assign \new_[4514]_  = (~\new_[5604]_  | ~\new_[19717]_ ) & (~\new_[5555]_  | ~\new_[1878]_ );
  assign \new_[4515]_  = ~\new_[10390]_  | ~\new_[6263]_  | ~\new_[8414]_  | ~\new_[11122]_ ;
  assign \new_[4516]_  = ~\new_[19277]_  | (~\new_[5778]_  & ~\new_[6132]_ );
  assign \new_[4517]_  = ~\new_[5792]_  | (~\new_[5766]_  & ~\new_[1878]_ );
  assign \new_[4518]_  = ~\new_[5793]_  | (~\new_[5718]_  & ~\new_[18791]_ );
  assign \new_[4519]_  = ~\new_[18791]_  & (~\new_[5848]_  | ~\new_[7610]_ );
  assign \new_[4520]_  = ~\new_[1879]_  & (~\new_[5849]_  | ~\new_[7604]_ );
  assign \new_[4521]_  = ~\new_[19480]_  & (~\new_[5851]_  | ~\new_[8616]_ );
  assign \new_[4522]_  = ~\new_[959]_  & (~\new_[7608]_  | ~\new_[5855]_ );
  assign \new_[4523]_  = ~\new_[19457]_  & (~\new_[8619]_  | ~\new_[5856]_ );
  assign \new_[4524]_  = ~\new_[7066]_  | (~\new_[5760]_  & ~\new_[18739]_ );
  assign \new_[4525]_  = ~\new_[5210]_  | ~\new_[10942]_ ;
  assign \new_[4526]_  = ~\new_[6375]_  | ~\new_[7966]_  | ~\new_[8588]_  | ~\new_[10396]_ ;
  assign \new_[4527]_  = ~\new_[10047]_  | ~\new_[10680]_  | ~\new_[6378]_  | ~\new_[8597]_ ;
  assign \new_[4528]_  = ~\new_[5248]_  | ~\new_[19528]_ ;
  assign \new_[4529]_  = ~\new_[10347]_  | ~\new_[11802]_  | ~\new_[6407]_  | ~\new_[8509]_ ;
  assign \new_[4530]_  = ~\new_[6454]_  | ~\new_[11805]_  | ~\new_[11163]_  | ~\new_[7542]_ ;
  assign \new_[4531]_  = ~\new_[6423]_  | ~\new_[10697]_  | ~\new_[11277]_  | ~\new_[6691]_ ;
  assign \new_[4532]_  = (~\new_[5717]_  | ~\new_[18941]_ ) & (~\new_[7882]_  | ~\new_[19029]_ );
  assign \new_[4533]_  = ~\new_[8302]_  | ~\new_[5720]_  | ~\new_[5684]_ ;
  assign \new_[4534]_  = ~\new_[8301]_  | ~\new_[6215]_  | ~\new_[5681]_ ;
  assign \new_[4535]_  = ~\new_[8299]_  | ~\new_[5753]_  | ~\new_[5683]_ ;
  assign \new_[4536]_  = ~\new_[5817]_  | ~\new_[5201]_ ;
  assign \new_[4537]_  = ~\new_[6553]_  | ~\new_[5240]_ ;
  assign \new_[4538]_  = ~\new_[5203]_  | ~\new_[5700]_ ;
  assign \new_[4539]_  = ~\new_[5818]_  | ~\new_[5204]_ ;
  assign \new_[4540]_  = ~\new_[9827]_  | ~\new_[6483]_  | ~\new_[10073]_  | ~\new_[14025]_ ;
  assign \new_[4541]_  = ~\new_[9861]_  | ~\new_[11246]_  | ~\new_[5775]_ ;
  assign \new_[4542]_  = ~\new_[9809]_  | ~\new_[5776]_  | ~\new_[10085]_ ;
  assign \new_[4543]_  = ~\new_[5152]_  | ~\new_[19442]_ ;
  assign \new_[4544]_  = ~\new_[5769]_  & ~\new_[12337]_  & ~\new_[14396]_ ;
  assign \new_[4545]_  = ~\new_[11475]_  | ~\new_[11759]_  | ~\new_[5703]_ ;
  assign \new_[4546]_  = ~\new_[5155]_  | ~\new_[960]_ ;
  assign \new_[4547]_  = ~\new_[10000]_  | ~\new_[5712]_  | ~\new_[6955]_ ;
  assign \new_[4548]_  = ~\new_[9876]_  | ~\new_[10339]_  | ~\new_[5777]_ ;
  assign \new_[4549]_  = ~\new_[5790]_  & ~\new_[11183]_  & ~\new_[8890]_ ;
  assign \new_[4550]_  = ~\new_[8276]_  | ~\new_[6383]_  | ~\new_[7000]_  | ~\new_[6534]_ ;
  assign \new_[4551]_  = ~\new_[5711]_  | ~\new_[9991]_  | ~\new_[5710]_ ;
  assign \new_[4552]_  = ~\new_[6554]_  | ~\new_[5241]_ ;
  assign \new_[4553]_  = ~\new_[19442]_  | (~\new_[5721]_  & ~\new_[11758]_ );
  assign \new_[4554]_  = ~\new_[5162]_  | ~\new_[18668]_ ;
  assign \new_[4555]_  = ~\new_[5172]_  | ~\new_[19246]_ ;
  assign \new_[4556]_  = ~\new_[9893]_  | ~\new_[10201]_  | ~\new_[6501]_  | ~\new_[14230]_ ;
  assign \new_[4557]_  = ~\new_[20805]_  & ~\new_[12374]_  & ~\new_[15203]_ ;
  assign \new_[4558]_  = ~\new_[10974]_  | ~\new_[5782]_  | ~\new_[10240]_ ;
  assign \new_[4559]_  = ~\new_[6555]_  | ~\new_[5242]_ ;
  assign \new_[4560]_  = ~\new_[9959]_  | ~\new_[5732]_  | ~\new_[6961]_ ;
  assign \new_[4561]_  = ~\new_[5803]_  & ~\new_[11371]_  & ~\new_[9037]_ ;
  assign \new_[4562]_  = ~\new_[9942]_  | ~\new_[6515]_  | ~\new_[11287]_  | ~\new_[10696]_ ;
  assign \new_[4563]_  = ~\new_[5736]_  | ~\new_[9952]_  | ~\new_[5735]_ ;
  assign \new_[4564]_  = ~\new_[5180]_  | ~\new_[18997]_ ;
  assign \new_[4565]_  = ~\new_[9943]_  | ~\new_[6518]_  | ~\new_[20382]_  | ~\new_[10621]_ ;
  assign \new_[4566]_  = ~\new_[18895]_  | (~\new_[5737]_  & ~\new_[9286]_ );
  assign \new_[4567]_  = ~\new_[5738]_  | ~\new_[9889]_  | ~\new_[6964]_ ;
  assign \new_[4568]_  = ~\new_[6211]_  | ~\new_[9851]_  | ~\new_[5741]_ ;
  assign \new_[4569]_  = ~\new_[922]_  | (~\new_[5742]_  & ~\new_[8052]_ );
  assign \new_[4570]_  = ~\new_[5748]_  | ~\new_[9883]_  | ~\new_[5747]_ ;
  assign \new_[4571]_  = ~\new_[19418]_  | (~\new_[5755]_  & ~\new_[11931]_ );
  assign \new_[4572]_  = ~\new_[5386]_  | ~\new_[5223]_ ;
  assign \new_[4573]_  = ~\new_[18983]_  | (~\new_[5757]_  & ~\new_[10626]_ );
  assign \new_[4574]_  = ~\new_[8592]_  | ~\new_[6191]_  | ~\new_[5725]_ ;
  assign \new_[4575]_  = \new_[7617]_  | \new_[5142]_ ;
  assign \new_[4576]_  = \new_[7624]_  | \new_[5147]_ ;
  assign \new_[4577]_  = ~\new_[20152]_  & (~\new_[5674]_  | ~\new_[8188]_ );
  assign \new_[4578]_  = ~\new_[10089]_  & (~\new_[5834]_  | ~\new_[19578]_ );
  assign \new_[4579]_  = ~\new_[5107]_  | ~\new_[10039]_ ;
  assign \new_[4580]_  = ~\new_[7859]_  & (~\new_[5835]_  | ~\new_[20941]_ );
  assign \new_[4581]_  = ~\new_[5306]_  | (~\new_[5791]_  & ~\new_[19787]_ );
  assign \new_[4582]_  = ~\new_[11210]_  & (~\new_[5836]_  | ~\new_[19561]_ );
  assign \new_[4583]_  = (~\new_[5750]_  | ~\new_[17119]_ ) & (~\new_[11349]_  | ~\new_[17472]_ );
  assign \new_[4584]_  = ~\new_[5320]_  | (~\new_[5800]_  & ~\new_[19236]_ );
  assign \new_[4585]_  = ~\new_[10234]_  | ~\new_[6287]_  | ~\new_[5730]_  | ~\new_[20557]_ ;
  assign \new_[4586]_  = ~\new_[5110]_  | ~\new_[10203]_ ;
  assign \new_[4587]_  = ~\new_[7908]_  & (~\new_[5837]_  | ~\new_[19599]_ );
  assign \new_[4588]_  = ~\new_[7932]_  | (~\new_[5838]_  & ~\new_[1033]_ );
  assign \new_[4589]_  = ~\new_[9051]_  & (~\new_[5839]_  | ~\new_[19448]_ );
  assign \new_[4590]_  = ~\new_[6875]_  & (~\new_[5840]_  | ~\new_[19236]_ );
  assign \new_[4591]_  = ~\new_[10023]_  | ~\new_[6279]_  | ~\new_[5659]_  | ~\new_[11100]_ ;
  assign \new_[4592]_  = ~\new_[10115]_  | ~\new_[6282]_  | ~\new_[5661]_  | ~\new_[11356]_ ;
  assign \new_[4593]_  = ~\new_[10221]_  | ~\new_[6285]_  | ~\new_[5662]_  | ~\new_[7910]_ ;
  assign \new_[4594]_  = ~\new_[11952]_  | ~\new_[5269]_  | ~\new_[5847]_ ;
  assign \new_[4595]_  = ~\new_[6369]_  | ~\new_[10819]_  | ~\new_[8211]_  | ~\new_[10159]_ ;
  assign \new_[4596]_  = \new_[6544]_  | \new_[8856]_  | \new_[11360]_  | \new_[21341]_ ;
  assign \new_[4597]_  = \new_[6541]_  | \new_[21120]_  | \new_[8955]_  | \new_[13076]_ ;
  assign \new_[4598]_  = ~\new_[5140]_  | ~\new_[18293]_ ;
  assign \new_[4599]_  = (~\new_[5785]_  | ~\new_[19528]_ ) & (~\new_[16285]_  | ~\new_[12446]_ );
  assign \new_[4600]_  = (~\new_[5773]_  | ~\new_[19350]_ ) & (~\new_[9701]_  | ~\new_[18194]_ );
  assign \new_[4601]_  = ~\new_[5207]_  & (~\new_[10489]_  | ~\new_[19780]_ );
  assign \new_[4602]_  = ~\new_[19448]_  | (~\new_[5696]_  & ~\new_[10360]_ );
  assign \new_[4603]_  = ~\new_[18803]_  & (~\new_[5680]_  | ~\new_[12089]_ );
  assign \new_[4604]_  = ~\new_[19259]_  | (~\new_[5845]_  & ~\new_[11627]_ );
  assign \new_[4605]_  = ~\new_[6123]_  | (~\new_[5799]_  & ~\new_[18769]_ );
  assign \new_[4606]_  = ~\new_[6276]_  | ~\new_[12683]_  | ~\new_[14542]_  | ~\new_[9121]_ ;
  assign \new_[4607]_  = ~\new_[13775]_  | ~\new_[15177]_  | ~\new_[5669]_ ;
  assign \new_[4608]_  = ~\new_[9940]_  | ~\new_[8521]_  | ~\new_[6332]_  | ~\new_[9853]_ ;
  assign \new_[4609]_  = ~\new_[9281]_  | ~\new_[14991]_  | ~\new_[5672]_ ;
  assign \new_[4610]_  = ~\new_[8026]_  | ~\new_[14186]_  | ~\new_[5673]_ ;
  assign \new_[4611]_  = ~\new_[8752]_  | ~\new_[6318]_  | ~\new_[8465]_  | ~\new_[9811]_ ;
  assign \new_[4612]_  = ~\new_[11007]_  | ~\new_[6326]_  | ~\new_[9603]_  | ~\new_[10002]_ ;
  assign \new_[4613]_  = ~\new_[5111]_  | (~\new_[6259]_  & ~\new_[18763]_ );
  assign \new_[4614]_  = ~\new_[5113]_  | (~\new_[6262]_  & ~\new_[999]_ );
  assign \new_[4615]_  = ~\new_[4830]_ ;
  assign \new_[4616]_  = ~\new_[5160]_  & ~\new_[6164]_ ;
  assign \new_[4617]_  = ~\new_[8347]_  | ~\new_[5677]_  | ~\new_[5852]_ ;
  assign \new_[4618]_  = ~\new_[8819]_  | ~\new_[6295]_  | ~\new_[8578]_  | ~\new_[11524]_ ;
  assign \new_[4619]_  = ~\new_[8799]_  | ~\new_[6291]_  | ~\new_[9564]_  | ~\new_[11544]_ ;
  assign \new_[4620]_  = ~\new_[8758]_  | ~\new_[10183]_  | ~\new_[6292]_  | ~\new_[11287]_ ;
  assign \new_[4621]_  = ~\new_[11034]_  | ~\new_[6293]_  | ~\new_[8551]_  | ~\new_[11046]_ ;
  assign \new_[4622]_  = ~\new_[9988]_  | ~\new_[6294]_  | ~\new_[6694]_  | ~\new_[11608]_ ;
  assign \new_[4623]_  = ~\new_[6120]_  | ~\new_[7029]_  | ~\new_[6708]_  | ~\new_[11584]_ ;
  assign \new_[4624]_  = ~\new_[5615]_  & (~\new_[5992]_  | ~\new_[19257]_ );
  assign \new_[4625]_  = ~\new_[5608]_  & (~\new_[5812]_  | ~\new_[19653]_ );
  assign \new_[4626]_  = ~\new_[5202]_  | (~\new_[6255]_  & ~\new_[18641]_ );
  assign \new_[4627]_  = ~\new_[5613]_  & (~\new_[5813]_  | ~\new_[19049]_ );
  assign \new_[4628]_  = ~\new_[5218]_  | (~\new_[6257]_  & ~\new_[19433]_ );
  assign \new_[4629]_  = ~\new_[5616]_  | (~\new_[5814]_  & ~\new_[1033]_ );
  assign \new_[4630]_  = ~\new_[5222]_  | (~\new_[5815]_  & ~\new_[19530]_ );
  assign \new_[4631]_  = ~\new_[5366]_  | ~\new_[19120]_ ;
  assign \new_[4632]_  = ~\new_[19277]_  | (~\new_[21161]_  & ~\new_[6862]_ );
  assign \new_[4633]_  = ~\new_[19467]_  | (~\new_[6007]_  & ~\new_[7179]_ );
  assign \new_[4634]_  = ~\new_[19277]_  | (~\new_[5986]_  & ~\new_[8810]_ );
  assign \new_[4635]_  = ~\new_[18965]_  & (~\new_[9061]_  | ~\new_[5896]_ );
  assign \new_[4636]_  = ~\new_[18833]_  & (~\new_[6884]_  | ~\new_[5897]_ );
  assign \new_[4637]_  = ~\new_[5886]_  & ~\new_[11574]_  & ~\new_[14228]_ ;
  assign \new_[4638]_  = ~\new_[18280]_  & (~\new_[8977]_  | ~\new_[5898]_ );
  assign \new_[4639]_  = ~\new_[19322]_  | (~\new_[6410]_  & ~\new_[5987]_ );
  assign \new_[4640]_  = ~\new_[984]_  | (~\new_[6022]_  & ~\new_[10546]_ );
  assign \new_[4641]_  = ~\new_[5341]_  | ~\new_[18895]_ ;
  assign \new_[4642]_  = ~\new_[5344]_  | ~\new_[19530]_ ;
  assign \new_[4643]_  = ~\new_[5368]_  & (~\new_[15927]_  | ~\new_[18891]_ );
  assign \new_[4644]_  = ~\new_[5254]_  & (~\new_[12578]_  | ~\new_[17478]_ );
  assign \new_[4645]_  = ~\new_[4869]_ ;
  assign \new_[4646]_  = ~\new_[4870]_ ;
  assign \new_[4647]_  = ~\new_[5377]_  | ~\new_[18895]_ ;
  assign \new_[4648]_  = (~\new_[5972]_  | ~\new_[19748]_ ) & (~\new_[12946]_  | ~\new_[18021]_ );
  assign \new_[4649]_  = ~\new_[19243]_  | (~\new_[5911]_  & ~\new_[12635]_ );
  assign \new_[4650]_  = ~\new_[5376]_  & ~\new_[1878]_ ;
  assign \new_[4651]_  = ~\new_[5347]_  | ~\new_[19343]_ ;
  assign \new_[4652]_  = (~\new_[5977]_  | ~\new_[19277]_ ) & (~\new_[13028]_  | ~\new_[17977]_ );
  assign \new_[4653]_  = ~\new_[19457]_  | (~\new_[5949]_  & ~\new_[14164]_ );
  assign \new_[4654]_  = ~\new_[19740]_  & (~\new_[6065]_  | ~\new_[5954]_ );
  assign \new_[4655]_  = ~\new_[5918]_  | ~\new_[6882]_  | ~\new_[12897]_ ;
  assign \new_[4656]_  = ~\new_[19623]_  | (~\new_[6643]_  & ~\new_[5880]_ );
  assign \new_[4657]_  = ~\new_[5364]_  | ~\new_[19530]_ ;
  assign \new_[4658]_  = ~\new_[5319]_  | ~\new_[19300]_ ;
  assign \new_[4659]_  = ~\new_[5367]_  | ~\new_[18599]_ ;
  assign \new_[4660]_  = ~\new_[5870]_  & ~\new_[11146]_  & ~\new_[12272]_ ;
  assign \new_[4661]_  = ~\new_[19702]_  & (~\new_[8416]_  | ~\new_[5959]_ );
  assign \new_[4662]_  = ~\new_[19512]_  | (~\new_[5893]_  & ~\new_[12017]_ );
  assign \new_[4663]_  = ~\new_[5259]_  & (~\new_[10570]_  | ~\new_[18021]_ );
  assign \new_[4664]_  = ~\new_[19509]_  | (~\new_[5894]_  & ~\new_[13172]_ );
  assign \new_[4665]_  = ~\new_[4908]_ ;
  assign \new_[4666]_  = ~\new_[5260]_  & (~\new_[12502]_  | ~\new_[17977]_ );
  assign \new_[4667]_  = ~\new_[19400]_  | (~\new_[5895]_  & ~\new_[12151]_ );
  assign \new_[4668]_  = ~\new_[9801]_  | ~\new_[6996]_  | ~\new_[5901]_ ;
  assign \new_[4669]_  = ~\new_[11076]_  | ~\new_[10605]_  | ~\new_[5873]_ ;
  assign \new_[4670]_  = ~\new_[4914]_ ;
  assign \new_[4671]_  = ~\new_[10735]_  | ~\new_[5298]_  | ~\new_[6560]_ ;
  assign \new_[4672]_  = ~\new_[9353]_  | ~\new_[5301]_  | ~\new_[6010]_ ;
  assign \new_[4673]_  = ~\new_[10994]_  | ~\new_[10595]_  | ~\new_[5877]_ ;
  assign \new_[4674]_  = ~\new_[5314]_  | ~\new_[19448]_ ;
  assign \new_[4675]_  = ~\new_[9319]_  | ~\new_[5315]_  | ~\new_[6566]_ ;
  assign \new_[4676]_  = ~\new_[19326]_  | (~\new_[5947]_  & ~\new_[11883]_ );
  assign \new_[4677]_  = (~\new_[5973]_  | ~\new_[19803]_ ) & (~\new_[17255]_  | ~\new_[17488]_ );
  assign \new_[4678]_  = ~\new_[7425]_  | ~\new_[5308]_ ;
  assign \new_[4679]_  = (~\new_[5978]_  | ~\new_[19780]_ ) & (~\new_[14554]_  | ~\new_[17640]_ );
  assign \new_[4680]_  = ~\new_[6415]_  | ~\new_[13283]_  | ~\new_[10148]_  | ~\new_[8534]_ ;
  assign \new_[4681]_  = (~\new_[6008]_  | ~\new_[21630]_ ) & (~\new_[8951]_  | ~\new_[21634]_ );
  assign \new_[4682]_  = (~\new_[5970]_  | ~\new_[19578]_ ) & (~\new_[16445]_  | ~\new_[17761]_ );
  assign \new_[4683]_  = ~\new_[8832]_  | ~\new_[5279]_ ;
  assign \new_[4684]_  = ~\new_[10170]_  | ~\new_[5280]_ ;
  assign \new_[4685]_  = ~\new_[10280]_  & (~\new_[6016]_  | ~\new_[1025]_ );
  assign \new_[4686]_  = ~\new_[5477]_  | ~\new_[19163]_ ;
  assign \new_[4687]_  = ~\new_[5458]_  | ~\new_[19517]_ ;
  assign \new_[4688]_  = ~\new_[5465]_  | ~\new_[18803]_ ;
  assign \new_[4689]_  = ~\new_[20645]_  | (~\new_[5511]_  & ~\new_[6664]_ );
  assign \new_[4690]_  = ~\new_[5469]_  | ~\new_[20763]_ ;
  assign \new_[4691]_  = \new_[5435]_  & \new_[15325]_ ;
  assign \new_[4692]_  = ~\new_[5434]_  | ~\new_[7408]_ ;
  assign \new_[4693]_  = \new_[5466]_  & \new_[12089]_ ;
  assign \new_[4694]_  = ~\new_[5478]_  & ~\new_[19748]_ ;
  assign \new_[4695]_  = ~\new_[923]_  | (~\new_[7536]_  & ~\new_[6033]_ );
  assign \new_[4696]_  = ~\new_[5452]_  | ~\new_[7600]_ ;
  assign \new_[4697]_  = ~\new_[6411]_  | ~\new_[20702]_  | ~\new_[10049]_  | ~\new_[8529]_ ;
  assign \new_[4698]_  = ~\new_[17335]_  & (~\new_[5504]_  | ~\new_[15379]_ );
  assign \new_[4699]_  = ~\new_[17244]_  & (~\new_[5506]_  | ~\new_[13046]_ );
  assign \new_[4700]_  = ~\new_[15901]_  & (~\new_[5497]_  | ~\new_[13080]_ );
  assign \new_[4701]_  = \new_[5447]_  & \new_[18154]_ ;
  assign \new_[4702]_  = ~\new_[5450]_  | ~\new_[5950]_ ;
  assign \new_[4703]_  = ~\new_[5032]_ ;
  assign \new_[4704]_  = ~\new_[5045]_ ;
  assign \new_[4705]_  = ~\new_[19748]_  | (~\new_[5525]_  & ~\new_[7920]_ );
  assign \new_[4706]_  = ~\new_[5046]_ ;
  assign \new_[4707]_  = \new_[5088]_  & \new_[20486]_ ;
  assign \new_[4708]_  = ~\new_[6176]_  & (~\new_[5514]_  | ~\new_[19578]_ );
  assign \new_[4709]_  = ~\new_[5483]_  | ~\new_[19770]_ ;
  assign \new_[4710]_  = ~\new_[5695]_  & (~\new_[5515]_  | ~\new_[19323]_ );
  assign \new_[4711]_  = ~\new_[6179]_  & (~\new_[5516]_  | ~\new_[19561]_ );
  assign \new_[4712]_  = ~\new_[5484]_  | ~\new_[20789]_ ;
  assign \new_[4713]_  = ~\new_[19448]_  | (~\new_[5501]_  & ~\new_[8990]_ );
  assign \new_[4714]_  = ~\new_[19527]_  | (~\new_[5505]_  & ~\new_[10264]_ );
  assign \new_[4715]_  = ~\new_[5486]_  | ~\new_[19032]_ ;
  assign \new_[4716]_  = ~\new_[19480]_  | (~\new_[5523]_  & ~\new_[8191]_ );
  assign \new_[4717]_  = ~\new_[19405]_  | (~\new_[5524]_  & ~\new_[8193]_ );
  assign \new_[4718]_  = ~\new_[5482]_  | (~\new_[12816]_  & ~\new_[18739]_ );
  assign \new_[4719]_  = ~\new_[19780]_  | (~\new_[5540]_  & ~\new_[8859]_ );
  assign \new_[4720]_  = ~\new_[19483]_  | (~\new_[5595]_  & ~\new_[10380]_ );
  assign \new_[4721]_  = ~\new_[19748]_  | (~\new_[5628]_  & ~\new_[8906]_ );
  assign \new_[4722]_  = ~\new_[19271]_  | (~\new_[5634]_  & ~\new_[7852]_ );
  assign \new_[4723]_  = ~\new_[19448]_  | (~\new_[5630]_  & ~\new_[8965]_ );
  assign \new_[4724]_  = ~\new_[19163]_  | (~\new_[5631]_  & ~\new_[6909]_ );
  assign \new_[4725]_  = ~\new_[19659]_  | (~\new_[5633]_  & ~\new_[9162]_ );
  assign \new_[4726]_  = (~\new_[5538]_  | ~\new_[19242]_ ) & (~\new_[12045]_  | ~\new_[18937]_ );
  assign \new_[4727]_  = ~\new_[19536]_  | (~\new_[5602]_  & ~\new_[8253]_ );
  assign \new_[4728]_  = ~\new_[19453]_  | (~\new_[5543]_  & ~\new_[8872]_ );
  assign \new_[4729]_  = ~\new_[19378]_  | (~\new_[5549]_  & ~\new_[10097]_ );
  assign \new_[4730]_  = ~\new_[18997]_  | (~\new_[5553]_  & ~\new_[13055]_ );
  assign \new_[4731]_  = ~\new_[984]_  | (~\new_[5554]_  & ~\new_[9050]_ );
  assign \new_[4732]_  = \new_[5355]_  | \new_[5094]_ ;
  assign \new_[4733]_  = ~\new_[8641]_  | ~\new_[6193]_  | ~\new_[5230]_  | ~\new_[10055]_ ;
  assign \new_[4734]_  = ~\new_[19502]_  | (~\new_[5560]_  & ~\new_[13628]_ );
  assign \new_[4735]_  = ~\new_[7261]_  & ~\new_[5095]_ ;
  assign \new_[4736]_  = ~\new_[19378]_  | (~\new_[5565]_  & ~\new_[8194]_ );
  assign \new_[4737]_  = ~\new_[19441]_  | (~\new_[5572]_  & ~\new_[8968]_ );
  assign \new_[4738]_  = ~\new_[19517]_  | (~\new_[5574]_  & ~\new_[8986]_ );
  assign \new_[4739]_  = ~\new_[922]_  | (~\new_[5575]_  & ~\new_[8999]_ );
  assign \new_[4740]_  = ~\new_[19120]_  | (~\new_[5581]_  & ~\new_[9040]_ );
  assign \new_[4741]_  = ~\new_[9743]_  | ~\new_[6208]_  | ~\new_[5232]_  | ~\new_[11211]_ ;
  assign \new_[4742]_  = ~\new_[18583]_  | (~\new_[20211]_  & ~\new_[10106]_ );
  assign \new_[4743]_  = ~\new_[5093]_  | ~\new_[991]_ ;
  assign \new_[4744]_  = ~\new_[19530]_  | (~\new_[5587]_  & ~\new_[8202]_ );
  assign \new_[4745]_  = (~\new_[5594]_  | ~\new_[19271]_ ) & (~\new_[13351]_  | ~\new_[18941]_ );
  assign \new_[4746]_  = ~\new_[6236]_  | ~\new_[12190]_  | ~\new_[10786]_  | ~\new_[7033]_ ;
  assign \new_[4747]_  = \new_[5100]_  | \new_[9504]_ ;
  assign \new_[4748]_  = ~\new_[7961]_  & (~\new_[5623]_  | ~\new_[1879]_ );
  assign \new_[4749]_  = ~\new_[1878]_  & (~\new_[5566]_  | ~\new_[8272]_ );
  assign \new_[4750]_  = ~\new_[7874]_  & (~\new_[5627]_  | ~\new_[18668]_ );
  assign \new_[4751]_  = ~\new_[6934]_  | ~\new_[12513]_  | ~\new_[6308]_  | ~\new_[15264]_ ;
  assign \new_[4752]_  = ~\new_[6936]_  | ~\new_[11712]_  | ~\new_[6311]_  | ~\new_[14797]_ ;
  assign \new_[4753]_  = ~\new_[6937]_  | ~\new_[11675]_  | ~\new_[6312]_  | ~\new_[13184]_ ;
  assign \new_[4754]_  = ~\new_[9775]_  | ~\new_[9530]_  | ~\new_[5626]_  | ~\new_[9502]_ ;
  assign \new_[4755]_  = ~\new_[9060]_  | ~\new_[6994]_  | ~\new_[7498]_  | ~\new_[10202]_ ;
  assign \new_[4756]_  = ~\new_[11519]_  | ~\new_[6919]_  | ~\new_[6983]_  | ~\new_[13044]_ ;
  assign \new_[4757]_  = ~\new_[11590]_  | ~\new_[6922]_  | ~\new_[6991]_  | ~\new_[12850]_ ;
  assign \new_[4758]_  = ~\new_[9268]_  | ~\new_[6992]_  | ~\new_[6923]_  | ~\new_[12915]_ ;
  assign \new_[4759]_  = ~\new_[15165]_  | ~\new_[6974]_  | ~\new_[5636]_  | ~\new_[7965]_ ;
  assign \new_[4760]_  = ~\new_[7015]_  | ~\new_[8401]_  | ~\new_[13000]_  | ~\new_[11058]_ ;
  assign \new_[4761]_  = ~\new_[9976]_  | ~\new_[5529]_ ;
  assign \new_[4762]_  = ~\new_[5714]_  & (~\new_[6876]_  | ~\new_[19343]_ );
  assign \new_[4763]_  = ~\new_[1025]_  & (~\new_[6270]_  | ~\new_[9441]_ );
  assign \new_[4764]_  = ~\new_[18583]_  & (~\new_[9691]_  | ~\new_[6275]_ );
  assign \new_[4765]_  = ~\new_[7045]_  | (~\new_[6198]_  & ~\new_[19005]_ );
  assign \new_[4766]_  = ~\new_[6335]_  & (~\new_[6216]_  | ~\new_[21562]_ );
  assign \new_[4767]_  = ~\new_[7064]_  | (~\new_[6218]_  & ~\new_[1084]_ );
  assign \new_[4768]_  = ~\new_[5603]_  | ~\new_[10900]_ ;
  assign \new_[4769]_  = ~\new_[5605]_  | ~\new_[10929]_ ;
  assign \new_[4770]_  = ~\new_[10625]_  | ~\new_[6203]_  | ~\new_[8723]_ ;
  assign \new_[4771]_  = ~\new_[10144]_  & (~\new_[6181]_  | ~\new_[19239]_ );
  assign \new_[4772]_  = (~\new_[6213]_  | ~\new_[21631]_ ) & (~\new_[9085]_  | ~\new_[21630]_ );
  assign \new_[4773]_  = ~\new_[6156]_  | ~\new_[7077]_  | ~\new_[6466]_ ;
  assign \new_[4774]_  = ~\new_[19536]_  | (~\new_[10783]_  & ~\new_[6226]_ );
  assign \new_[4775]_  = ~\new_[19442]_  | (~\new_[6976]_  & ~\new_[6617]_ );
  assign \new_[4776]_  = ~\new_[18649]_  | (~\new_[6619]_  & ~\new_[6227]_ );
  assign \new_[4777]_  = ~\new_[8744]_  | ~\new_[7254]_  | ~\new_[7846]_  | ~\new_[13303]_ ;
  assign \new_[4778]_  = ~\new_[5542]_  | ~\new_[19528]_ ;
  assign \new_[4779]_  = ~\new_[10620]_  | ~\new_[7263]_  | ~\new_[10072]_  | ~\new_[11914]_ ;
  assign \new_[4780]_  = ~\new_[5544]_  | ~\new_[18763]_ ;
  assign \new_[4781]_  = ~\new_[6157]_  | ~\new_[7100]_  | ~\new_[6070]_ ;
  assign \new_[4782]_  = ~\new_[5550]_  | ~\new_[18649]_ ;
  assign \new_[4783]_  = ~\new_[5551]_  | ~\new_[19070]_ ;
  assign \new_[4784]_  = ~\new_[5557]_  | ~\new_[19453]_ ;
  assign \new_[4785]_  = ~\new_[19517]_  | (~\new_[6634]_  & ~\new_[6229]_ );
  assign \new_[4786]_  = ~\new_[12162]_  | ~\new_[14292]_  | ~\new_[6194]_ ;
  assign \new_[4787]_  = \new_[7258]_  | \new_[13650]_  | \new_[10670]_  | \new_[10949]_ ;
  assign \new_[4788]_  = ~\new_[921]_  | (~\new_[6219]_  & ~\new_[9300]_ );
  assign \new_[4789]_  = ~\new_[18808]_  | (~\new_[6639]_  & ~\new_[6230]_ );
  assign \new_[4790]_  = ~\new_[5561]_  | ~\new_[19502]_ ;
  assign \new_[4791]_  = ~\new_[13686]_  | ~\new_[14584]_  | ~\new_[6195]_ ;
  assign \new_[4792]_  = ~\new_[5567]_  | ~\new_[18983]_ ;
  assign \new_[4793]_  = ~\new_[18983]_  | (~\new_[6648]_  & ~\new_[6231]_ );
  assign \new_[4794]_  = ~\new_[5573]_  | ~\new_[999]_ ;
  assign \new_[4795]_  = ~\new_[6158]_  | ~\new_[7146]_  | ~\new_[6781]_ ;
  assign \new_[4796]_  = ~\new_[19318]_  | (~\new_[10803]_  & ~\new_[6228]_ );
  assign \new_[4797]_  = ~\new_[19433]_  | (~\new_[6232]_  & ~\new_[8472]_ );
  assign \new_[4798]_  = \new_[7271]_  | \new_[10365]_  | \new_[13646]_  | \new_[11008]_ ;
  assign \new_[4799]_  = ~\new_[10345]_  | ~\new_[7272]_  | ~\new_[7801]_  | ~\new_[8777]_ ;
  assign \new_[4800]_  = ~\new_[19246]_  | (~\new_[6658]_  & ~\new_[6233]_ );
  assign \new_[4801]_  = ~\new_[7803]_  | ~\new_[7273]_  | ~\new_[7918]_  | ~\new_[13216]_ ;
  assign \new_[4802]_  = ~\new_[5576]_  | ~\new_[1026]_ ;
  assign \new_[4803]_  = ~\new_[5577]_  | ~\new_[18808]_ ;
  assign \new_[4804]_  = ~\new_[5580]_  | ~\new_[19441]_ ;
  assign \new_[4805]_  = ~\new_[5582]_  | ~\new_[18619]_ ;
  assign \new_[4806]_  = ~\new_[5584]_  | ~\new_[19523]_ ;
  assign \new_[4807]_  = ~\new_[5586]_  | ~\new_[19433]_ ;
  assign \new_[4808]_  = ~\new_[991]_  | (~\new_[6209]_  & ~\new_[12953]_ );
  assign \new_[4809]_  = ~\new_[5545]_  | ~\new_[19070]_ ;
  assign \new_[4810]_  = ~\new_[18803]_  | (~\new_[6212]_  & ~\new_[9173]_ );
  assign \new_[4811]_  = ~\new_[5536]_  | ~\new_[19751]_ ;
  assign \new_[4812]_  = ~\new_[5541]_  & (~\new_[10052]_  | ~\new_[18498]_ );
  assign \new_[4813]_  = ~\new_[10113]_  & (~\new_[6266]_  | ~\new_[19803]_ );
  assign \new_[4814]_  = (~\new_[6201]_  | ~\new_[21561]_ ) & (~\new_[9033]_  | ~\new_[21562]_ );
  assign \new_[4815]_  = (~\new_[6202]_  | ~\new_[19382]_ ) & (~\new_[11251]_  | ~\new_[19587]_ );
  assign \new_[4816]_  = \new_[7292]_  | \new_[9167]_  | \new_[10042]_  | \new_[12851]_ ;
  assign \new_[4817]_  = \new_[7293]_  | \new_[8855]_  | \new_[11121]_  | \new_[15208]_ ;
  assign \new_[4818]_  = \new_[7294]_  | \new_[10098]_  | \new_[8831]_  | \new_[12495]_ ;
  assign \new_[4819]_  = \new_[7295]_  | \new_[11269]_  | \new_[9024]_  | \new_[12841]_ ;
  assign \new_[4820]_  = \new_[7296]_  | \new_[10250]_  | \new_[9117]_  | \new_[13251]_ ;
  assign \new_[4821]_  = \new_[7297]_  | \new_[9096]_  | \new_[11321]_  | \new_[12922]_ ;
  assign \new_[4822]_  = \new_[7300]_  | \new_[8923]_  | \new_[10346]_  | \new_[15257]_ ;
  assign \new_[4823]_  = \new_[7299]_  | \new_[9127]_  | \new_[10349]_  | \new_[12454]_ ;
  assign \new_[4824]_  = ~\new_[7193]_  | ~\new_[15325]_  | ~\new_[11176]_  | ~\new_[15225]_ ;
  assign \new_[4825]_  = ~\new_[6557]_  | (~\new_[6237]_  & ~\new_[1879]_ );
  assign \new_[4826]_  = ~\new_[6563]_  | (~\new_[6238]_  & ~\new_[19502]_ );
  assign \new_[4827]_  = ~\new_[7340]_  | ~\new_[10911]_  | ~\new_[10788]_  | ~\new_[15612]_ ;
  assign \new_[4828]_  = ~\new_[7019]_  | ~\new_[9125]_  | ~\new_[15612]_  | ~\new_[15095]_ ;
  assign \new_[4829]_  = ~\new_[9850]_  | ~\new_[7052]_  | ~\new_[8391]_  | ~\new_[9902]_ ;
  assign \new_[4830]_  = ~\new_[7303]_  | ~\new_[8786]_  | ~\new_[5850]_  | ~\new_[8364]_ ;
  assign \new_[4831]_  = (~\new_[6241]_  | ~\new_[19502]_ ) & (~\new_[11054]_  | ~\new_[19532]_ );
  assign \new_[4832]_  = ~\new_[7816]_  | ~\new_[7030]_  | ~\new_[6719]_  | ~\new_[11570]_ ;
  assign \new_[4833]_  = ~\new_[9954]_  | ~\new_[7027]_  | ~\new_[9655]_  | ~\new_[10559]_ ;
  assign \new_[4834]_  = ~\new_[8800]_  | ~\new_[7028]_  | ~\new_[8552]_  | ~\new_[11709]_ ;
  assign \new_[4835]_  = (~\new_[6234]_  | ~\new_[19339]_ ) & (~\new_[19483]_  | ~\new_[7130]_ );
  assign \new_[4836]_  = ~\new_[5614]_  | (~\new_[6256]_  & ~\new_[954]_ );
  assign \new_[4837]_  = ~\new_[5854]_  | ~\new_[19578]_ ;
  assign \new_[4838]_  = ~\new_[19717]_  | (~\new_[6346]_  & ~\new_[11380]_ );
  assign \new_[4839]_  = ~\new_[5807]_  | ~\new_[19751]_ ;
  assign \new_[4840]_  = ~\new_[19170]_  | (~\new_[6054]_  & ~\new_[7191]_ );
  assign \new_[4841]_  = ~\new_[19512]_  | (~\new_[9388]_  & ~\new_[6419]_ );
  assign \new_[4842]_  = ~\new_[19337]_  | (~\new_[6522]_  & ~\new_[8780]_ );
  assign \new_[4843]_  = ~\new_[17689]_  & (~\new_[8867]_  | ~\new_[6339]_ );
  assign \new_[4844]_  = ~\new_[7570]_  | ~\new_[11364]_  | ~\new_[6524]_ ;
  assign \new_[4845]_  = ~\new_[6357]_  | ~\new_[6558]_  | ~\new_[8184]_ ;
  assign \new_[4846]_  = ~\new_[17475]_  | (~\new_[10081]_  & ~\new_[6297]_ );
  assign \new_[4847]_  = ~\new_[921]_  | (~\new_[7105]_  & ~\new_[6487]_ );
  assign \new_[4848]_  = ~\new_[10359]_  | (~\new_[6321]_  & ~\new_[18789]_ );
  assign \new_[4849]_  = ~\new_[6309]_  & ~\new_[12574]_  & ~\new_[12154]_ ;
  assign \new_[4850]_  = ~\new_[19239]_  & (~\new_[7969]_  | ~\new_[6341]_ );
  assign \new_[4851]_  = ~\new_[923]_  | (~\new_[7126]_  & ~\new_[6497]_ );
  assign \new_[4852]_  = ~\new_[9580]_  | ~\new_[12306]_  | ~\new_[6468]_ ;
  assign \new_[4853]_  = ~\new_[21558]_  & (~\new_[8949]_  | ~\new_[6343]_ );
  assign \new_[4854]_  = ~\new_[8824]_  | (~\new_[6325]_  & ~\new_[17660]_ );
  assign \new_[4855]_  = ~\new_[922]_  | (~\new_[7155]_  & ~\new_[6507]_ );
  assign \new_[4856]_  = ~\new_[18942]_  & (~\new_[6604]_  | ~\new_[13741]_ );
  assign \new_[4857]_  = ~\new_[10322]_  | (~\new_[6333]_  & ~\new_[20903]_ );
  assign \new_[4858]_  = ~\new_[18650]_  & (~\new_[8925]_  | ~\new_[6345]_ );
  assign \new_[4859]_  = ~\new_[5765]_  | ~\new_[19237]_ ;
  assign \new_[4860]_  = ~\new_[9464]_  | ~\new_[20987]_  | ~\new_[6537]_ ;
  assign \new_[4861]_  = ~\new_[5774]_  | ~\new_[18091]_ ;
  assign \new_[4862]_  = ~\new_[5783]_  | ~\new_[19322]_ ;
  assign \new_[4863]_  = ~\new_[19322]_  | (~\new_[6331]_  & ~\new_[8667]_ );
  assign \new_[4864]_  = ~\new_[1025]_  | (~\new_[6337]_  & ~\new_[10871]_ );
  assign \new_[4865]_  = ~\new_[5827]_  | ~\new_[19378]_ ;
  assign \new_[4866]_  = ~\new_[17660]_  & (~\new_[6470]_  | ~\new_[13823]_ );
  assign \new_[4867]_  = ~\new_[18418]_  | (~\new_[6351]_  & ~\new_[12518]_ );
  assign \new_[4868]_  = ~\new_[19243]_  & (~\new_[6472]_  | ~\new_[8030]_ );
  assign \new_[4869]_  = ~\new_[19748]_  & (~\new_[9478]_  | ~\new_[6574]_ );
  assign \new_[4870]_  = ~\new_[6355]_  | ~\new_[7978]_  | ~\new_[10610]_ ;
  assign \new_[4871]_  = ~\new_[13553]_  & (~\new_[6456]_  | ~\new_[18998]_ );
  assign \new_[4872]_  = ~\new_[16418]_  & ~\new_[5844]_ ;
  assign \new_[4873]_  = \new_[5699]_  & \new_[9125]_ ;
  assign \new_[4874]_  = ~\new_[5693]_  & ~\new_[7963]_ ;
  assign \new_[4875]_  = ~\new_[18827]_  & (~\new_[6479]_  | ~\new_[11521]_ );
  assign \new_[4876]_  = ~\new_[10192]_  | ~\new_[12171]_  | ~\new_[6481]_ ;
  assign \new_[4877]_  = ~\new_[6358]_  | ~\new_[6904]_  | ~\new_[10694]_ ;
  assign \new_[4878]_  = ~\new_[10576]_  | ~\new_[13971]_  | ~\new_[7415]_  | ~\new_[11948]_ ;
  assign \new_[4879]_  = ~\new_[5694]_  & (~\new_[8114]_  | ~\new_[18965]_ );
  assign \new_[4880]_  = ~\new_[15080]_  | ~\new_[5771]_  | ~\new_[16077]_ ;
  assign \new_[4881]_  = ~\new_[19442]_  | (~\new_[8342]_  & ~\new_[6320]_ );
  assign \new_[4882]_  = ~\new_[18787]_  & (~\new_[6633]_  | ~\new_[6322]_ );
  assign \new_[4883]_  = ~\new_[19694]_  & (~\new_[8385]_  | ~\new_[6323]_ );
  assign \new_[4884]_  = ~\new_[5780]_  | ~\new_[19445]_ ;
  assign \new_[4885]_  = ~\new_[7369]_  | ~\new_[8395]_  | ~\new_[6469]_ ;
  assign \new_[4886]_  = ~\new_[5858]_  | ~\new_[10006]_ ;
  assign \new_[4887]_  = ~\new_[8621]_  | ~\new_[5853]_ ;
  assign \new_[4888]_  = ~\new_[12503]_  | ~\new_[5772]_  | ~\new_[13964]_ ;
  assign \new_[4889]_  = ~\new_[6389]_  | ~\new_[8692]_  | ~\new_[12308]_ ;
  assign \new_[4890]_  = ~\new_[19433]_  | (~\new_[9581]_  & ~\new_[6393]_ );
  assign \new_[4891]_  = ~\new_[10181]_  | ~\new_[10624]_  | ~\new_[6498]_ ;
  assign \new_[4892]_  = ~\new_[5173]_ ;
  assign \new_[4893]_  = ~\new_[944]_  | (~\new_[6398]_  & ~\new_[13096]_ );
  assign \new_[4894]_  = ~\new_[7370]_  | ~\new_[8474]_  | ~\new_[6503]_ ;
  assign \new_[4895]_  = ~\new_[19418]_  | (~\new_[7459]_  & ~\new_[6327]_ );
  assign \new_[4896]_  = ~\new_[9924]_  | ~\new_[6663]_  | ~\new_[9020]_  | ~\new_[11940]_ ;
  assign \new_[4897]_  = ~\new_[11015]_  | ~\new_[6666]_  | ~\new_[10677]_  | ~\new_[11272]_ ;
  assign \new_[4898]_  = ~\new_[12232]_  | ~\new_[8997]_  | ~\new_[5928]_  | ~\new_[10977]_ ;
  assign \new_[4899]_  = ~\new_[20537]_  & (~\new_[6036]_  | ~\new_[6329]_ );
  assign \new_[4900]_  = ~\new_[19770]_  & (~\new_[7475]_  | ~\new_[6330]_ );
  assign \new_[4901]_  = ~\new_[6613]_  | ~\new_[6041]_  | ~\new_[6516]_ ;
  assign \new_[4902]_  = ~\new_[5860]_  | ~\new_[9920]_ ;
  assign \new_[4903]_  = ~\new_[19259]_  & (~\new_[7505]_  | ~\new_[6334]_ );
  assign \new_[4904]_  = ~\new_[9874]_  & (~\new_[6520]_  | ~\new_[21267]_ );
  assign \new_[4905]_  = ~\new_[6344]_  | ~\new_[9068]_  | ~\new_[14299]_ ;
  assign \new_[4906]_  = ~\new_[9184]_  & (~\new_[6550]_  | ~\new_[19619]_ );
  assign \new_[4907]_  = ~\new_[5846]_  & ~\new_[12143]_ ;
  assign \new_[4908]_  = ~\new_[6437]_  | ~\new_[10356]_  | ~\new_[11926]_ ;
  assign \new_[4909]_  = ~\new_[21056]_  & (~\new_[6441]_  | ~\new_[21257]_ );
  assign \new_[4910]_  = ~\new_[5764]_  | ~\new_[19284]_ ;
  assign \new_[4911]_  = ~\new_[18606]_  & (~\new_[6453]_  | ~\new_[11585]_ );
  assign \new_[4912]_  = ~\new_[6770]_  & (~\new_[6444]_  | ~\new_[17475]_ );
  assign \new_[4913]_  = ~\new_[7306]_  | ~\new_[5701]_ ;
  assign \new_[4914]_  = ~\new_[19508]_  & (~\new_[6482]_  | ~\new_[12616]_ );
  assign \new_[4915]_  = ~\new_[7409]_  & ~\new_[5789]_ ;
  assign \new_[4916]_  = ~\new_[12217]_  | ~\new_[6760]_  | ~\new_[6376]_ ;
  assign \new_[4917]_  = ~\new_[5211]_ ;
  assign \new_[4918]_  = ~\new_[5212]_ ;
  assign \new_[4919]_  = ~\new_[5706]_  | ~\new_[17518]_ ;
  assign \new_[4920]_  = ~\new_[19002]_  | (~\new_[6436]_  & ~\new_[12828]_ );
  assign \new_[4921]_  = ~\new_[11933]_  | ~\new_[6207]_  | ~\new_[6570]_ ;
  assign \new_[4922]_  = ~\new_[5932]_  & (~\new_[6517]_  | ~\new_[21267]_ );
  assign \new_[4923]_  = ~\new_[19236]_  & (~\new_[6600]_  | ~\new_[8785]_ );
  assign \new_[4924]_  = ~\new_[19051]_  & (~\new_[6601]_  | ~\new_[9993]_ );
  assign \new_[4925]_  = ~\new_[5754]_  | ~\new_[17714]_ ;
  assign \new_[4926]_  = ~\new_[19041]_  | (~\new_[6430]_  & ~\new_[13121]_ );
  assign \new_[4927]_  = ~\new_[19051]_  | (~\new_[6435]_  & ~\new_[12911]_ );
  assign \new_[4928]_  = ~\new_[5756]_  | ~\new_[17697]_ ;
  assign \new_[4929]_  = ~\new_[8811]_  | ~\new_[6093]_  | ~\new_[6443]_ ;
  assign \new_[4930]_  = ~\new_[5758]_  | ~\new_[19257]_ ;
  assign \new_[4931]_  = ~\new_[19659]_  | (~\new_[6450]_  & ~\new_[15284]_ );
  assign \new_[4932]_  = ~\new_[5762]_  & (~\new_[11374]_  | ~\new_[19640]_ );
  assign \new_[4933]_  = ~\new_[20453]_  & (~\new_[11386]_  | ~\new_[20970]_ );
  assign \new_[4934]_  = ~\new_[20763]_  | (~\new_[6451]_  & ~\new_[15273]_ );
  assign \new_[4935]_  = (~\new_[6545]_  | ~\new_[17475]_ ) & (~\new_[11140]_  | ~\new_[19553]_ );
  assign \new_[4936]_  = ~\new_[7555]_  | ~\new_[5713]_ ;
  assign \new_[4937]_  = ~\new_[8284]_  & ~\new_[5637]_ ;
  assign \new_[4938]_  = ~\new_[7519]_  | ~\new_[5745]_ ;
  assign \new_[4939]_  = ~\new_[6689]_  | ~\new_[5746]_ ;
  assign \new_[4940]_  = ~\new_[7525]_  | ~\new_[5749]_ ;
  assign \new_[4941]_  = (~\new_[6596]_  | ~\new_[18786]_ ) & (~\new_[9308]_  | ~\new_[17544]_ );
  assign \new_[4942]_  = (~\new_[6592]_  | ~\new_[18154]_ ) & (~\new_[8063]_  | ~\new_[17939]_ );
  assign \new_[4943]_  = ~\new_[10378]_  | ~\new_[6819]_  | ~\new_[8425]_  | ~\new_[12035]_ ;
  assign \new_[4944]_  = ~\new_[13168]_  | ~\new_[6692]_  | ~\new_[6571]_ ;
  assign \new_[4945]_  = ~\new_[7341]_  | ~\new_[13496]_  | ~\new_[10040]_  | ~\new_[13558]_ ;
  assign \new_[4946]_  = ~\new_[7342]_  | ~\new_[14036]_  | ~\new_[12313]_  | ~\new_[12208]_ ;
  assign \new_[4947]_  = ~\new_[7343]_  | ~\new_[14880]_  | ~\new_[13560]_  | ~\new_[11181]_ ;
  assign \new_[4948]_  = ~\new_[8845]_  | (~\new_[6594]_  & ~\new_[18787]_ );
  assign \new_[4949]_  = ~\new_[8912]_  | (~\new_[6597]_  & ~\new_[20537]_ );
  assign \new_[4950]_  = ~\new_[8987]_  | (~\new_[6598]_  & ~\new_[20513]_ );
  assign \new_[4951]_  = ~\new_[13174]_  | ~\new_[8532]_  | ~\new_[6576]_ ;
  assign \new_[4952]_  = ~\new_[7344]_  | ~\new_[12003]_  | ~\new_[9142]_  | ~\new_[11546]_ ;
  assign \new_[4953]_  = ~\new_[19257]_  | (~\new_[10389]_  & ~\new_[6111]_ );
  assign \new_[4954]_  = ~\new_[5965]_  | ~\new_[19529]_ ;
  assign \new_[4955]_  = ~\new_[5966]_  | ~\new_[19442]_ ;
  assign \new_[4956]_  = ~\new_[5969]_  | ~\new_[921]_ ;
  assign \new_[4957]_  = ~\new_[19694]_  | (~\new_[10807]_  & ~\new_[6109]_ );
  assign \new_[4958]_  = ~\new_[5980]_  | ~\new_[922]_ ;
  assign \new_[4959]_  = ~\new_[21562]_  | (~\new_[6038]_  & ~\new_[20389]_ );
  assign \new_[4960]_  = ~\new_[19702]_  | (~\new_[9630]_  & ~\new_[6110]_ );
  assign \new_[4961]_  = ~\new_[20763]_  | (~\new_[6095]_  & ~\new_[8329]_ );
  assign \new_[4962]_  = ~\new_[21142]_  | (~\new_[6096]_  & ~\new_[8415]_ );
  assign \new_[4963]_  = ~\new_[19246]_  & (~\new_[6080]_  | ~\new_[20827]_ );
  assign \new_[4964]_  = ~\new_[19054]_  | (~\new_[6097]_  & ~\new_[8477]_ );
  assign \new_[4965]_  = ~\new_[19527]_  | (~\new_[6098]_  & ~\new_[9070]_ );
  assign \new_[4966]_  = ~\new_[21558]_  | (~\new_[6072]_  & ~\new_[15202]_ );
  assign \new_[4967]_  = ~\new_[5998]_  | ~\new_[19276]_ ;
  assign \new_[4968]_  = ~\new_[5999]_  | ~\new_[21142]_ ;
  assign \new_[4969]_  = ~\new_[19271]_  & (~\new_[7385]_  | ~\new_[6618]_ );
  assign \new_[4970]_  = ~\new_[18942]_  & (~\new_[9612]_  | ~\new_[6659]_ );
  assign \new_[4971]_  = ~\new_[5284]_ ;
  assign \new_[4972]_  = ~\new_[5920]_  | ~\new_[19102]_ ;
  assign \new_[4973]_  = ~\new_[5931]_  | ~\new_[19202]_ ;
  assign \new_[4974]_  = \new_[6223]_  ^ \new_[18602]_ ;
  assign \new_[4975]_  = ~\new_[6953]_  & (~\new_[8316]_  | ~\new_[18280]_ );
  assign \new_[4976]_  = ~\new_[5971]_  & ~\new_[19536]_ ;
  assign \new_[4977]_  = ~\new_[5910]_  | ~\new_[7644]_ ;
  assign \new_[4978]_  = ~\new_[19271]_  & (~\new_[6635]_  | ~\new_[7422]_ );
  assign \new_[4979]_  = ~\new_[5979]_  & ~\new_[11790]_ ;
  assign \new_[4980]_  = ~\new_[11103]_  | ~\new_[6027]_  | ~\new_[8653]_ ;
  assign \new_[4981]_  = ~\new_[5982]_  & ~\new_[19318]_ ;
  assign \new_[4982]_  = ~\new_[19709]_  & (~\new_[7507]_  | ~\new_[6045]_ );
  assign \new_[4983]_  = ~\new_[6053]_  & ~\new_[12798]_  & ~\new_[13314]_ ;
  assign \new_[4984]_  = \new_[6249]_  ^ \new_[18822]_ ;
  assign \new_[4985]_  = \new_[6250]_  ^ \new_[18723]_ ;
  assign \new_[4986]_  = ~\new_[5334]_ ;
  assign \new_[4987]_  = ~\new_[5948]_  | ~\new_[6710]_ ;
  assign \new_[4988]_  = ~\new_[5993]_  & ~\new_[6039]_ ;
  assign \new_[4989]_  = ~\new_[6753]_  | ~\new_[12948]_  | ~\new_[13620]_  | ~\new_[10040]_ ;
  assign \new_[4990]_  = ~\new_[11150]_  | ~\new_[5889]_  | ~\new_[11281]_ ;
  assign \new_[4991]_  = (~\new_[6660]_  | ~\new_[19088]_ ) & (~\new_[17373]_  | ~\new_[15461]_ );
  assign \new_[4992]_  = ~\new_[6621]_  & ~\new_[5874]_ ;
  assign \new_[4993]_  = ~\new_[5888]_  | ~\new_[18649]_ ;
  assign \new_[4994]_  = ~\new_[5351]_ ;
  assign \new_[4995]_  = ~\new_[5352]_ ;
  assign \new_[4996]_  = ~\new_[5983]_  & (~\new_[10923]_  | ~\new_[18965]_ );
  assign \new_[4997]_  = ~\new_[6000]_  & (~\new_[14775]_  | ~\new_[14984]_ );
  assign \new_[4998]_  = ~\new_[5975]_  & (~\new_[11060]_  | ~\new_[19239]_ );
  assign \new_[4999]_  = ~\new_[6637]_  & ~\new_[5879]_ ;
  assign \new_[5000]_  = ~\new_[5976]_  & (~\new_[10971]_  | ~\new_[18998]_ );
  assign \new_[5001]_  = ~\new_[7421]_  | (~\new_[6071]_  & ~\new_[17668]_ );
  assign \new_[5002]_  = ~\new_[5923]_  & ~\new_[10832]_ ;
  assign \new_[5003]_  = ~\new_[7453]_  & (~\new_[6082]_  | ~\new_[18077]_ );
  assign \new_[5004]_  = ~\new_[8481]_  & (~\new_[6083]_  | ~\new_[21638]_ );
  assign \new_[5005]_  = ~\new_[5890]_  | ~\new_[19120]_ ;
  assign \new_[5006]_  = ~\new_[5891]_  | ~\new_[21417]_ ;
  assign \new_[5007]_  = ~\new_[17688]_  & (~\new_[6074]_  | ~\new_[15224]_ );
  assign \new_[5008]_  = ~\new_[5372]_ ;
  assign \new_[5009]_  = ~\new_[6009]_  | ~\new_[6424]_ ;
  assign \new_[5010]_  = ~\new_[6017]_  & ~\new_[7223]_ ;
  assign \new_[5011]_  = ~\new_[5892]_  | ~\new_[19246]_ ;
  assign \new_[5012]_  = ~\new_[6018]_  & ~\new_[7224]_ ;
  assign \new_[5013]_  = ~\new_[5374]_ ;
  assign \new_[5014]_  = ~\new_[6019]_  & ~\new_[6464]_ ;
  assign \new_[5015]_  = ~\new_[5381]_ ;
  assign \new_[5016]_  = ~\new_[18525]_  | (~\new_[6641]_  & ~\new_[11755]_ );
  assign \new_[5017]_  = ~\new_[17629]_  | (~\new_[6056]_  & ~\new_[11784]_ );
  assign \new_[5018]_  = ~\new_[18300]_  | (~\new_[6061]_  & ~\new_[12956]_ );
  assign \new_[5019]_  = (~\new_[6094]_  | ~\new_[19070]_ ) & (~\new_[11345]_  | ~\new_[17669]_ );
  assign \new_[5020]_  = ~\new_[9375]_  | ~\new_[5899]_ ;
  assign \new_[5021]_  = ~\new_[6429]_  | ~\new_[5942]_ ;
  assign \new_[5022]_  = ~\new_[5883]_  & ~\new_[6654]_ ;
  assign \new_[5023]_  = ~\new_[5945]_  | ~\new_[5946]_ ;
  assign \new_[5024]_  = ~\new_[6714]_  & ~\new_[5884]_ ;
  assign \new_[5025]_  = ~\new_[7430]_  & ~\new_[5872]_ ;
  assign \new_[5026]_  = ~\new_[14119]_  | ~\new_[5960]_ ;
  assign \new_[5027]_  = ~\new_[13618]_  | (~\new_[6099]_  & ~\new_[18606]_ );
  assign \new_[5028]_  = ~\new_[13163]_  | ~\new_[5961]_ ;
  assign \new_[5029]_  = ~\new_[6872]_  | ~\new_[5864]_ ;
  assign \new_[5030]_  = (~\new_[6108]_  | ~\new_[19711]_ ) & (~\new_[12094]_  | ~\new_[19269]_ );
  assign \new_[5031]_  = (~\new_[6107]_  | ~\new_[21629]_ ) & (~\new_[13987]_  | ~\new_[19018]_ );
  assign \new_[5032]_  = ~\new_[5909]_  | ~\new_[6281]_ ;
  assign \new_[5033]_  = ~\new_[5915]_  & (~\new_[7424]_  | ~\new_[19204]_ );
  assign \new_[5034]_  = ~\new_[5417]_ ;
  assign \new_[5035]_  = ~\new_[5936]_  & (~\new_[6684]_  | ~\new_[21115]_ );
  assign \new_[5036]_  = ~\new_[5938]_  & (~\new_[7523]_  | ~\new_[21558]_ );
  assign \new_[5037]_  = \new_[5502]_  | \new_[19257]_ ;
  assign \new_[5038]_  = \new_[5499]_  | \new_[20645]_ ;
  assign \new_[5039]_  = ~\new_[6112]_  | ~\new_[9798]_  | ~\new_[12174]_ ;
  assign \new_[5040]_  = ~\new_[19659]_  | (~\new_[9152]_  & ~\new_[6122]_ );
  assign \new_[5041]_  = ~\new_[5433]_ ;
  assign \new_[5042]_  = ~\new_[6114]_  | ~\new_[8754]_  | ~\new_[12270]_ ;
  assign \new_[5043]_  = ~\new_[6023]_  | ~\new_[15777]_ ;
  assign \new_[5044]_  = ~\new_[5436]_ ;
  assign \new_[5045]_  = ~\new_[19436]_  & (~\new_[11258]_  | ~\new_[6149]_ );
  assign \new_[5046]_  = ~\new_[18606]_  & (~\new_[11290]_  | ~\new_[6147]_ );
  assign \new_[5047]_  = ~\new_[18409]_  | (~\new_[6118]_  & ~\new_[21387]_ );
  assign \new_[5048]_  = ~\new_[18973]_  & (~\new_[6119]_  | ~\new_[13875]_ );
  assign \new_[5049]_  = ~\new_[5509]_  | ~\new_[10509]_ ;
  assign \new_[5050]_  = ~\new_[6029]_  | ~\new_[19529]_ ;
  assign \new_[5051]_  = ~\new_[6028]_  | ~\new_[19277]_ ;
  assign \new_[5052]_  = (~\new_[6081]_  | ~\new_[19561]_ ) & (~\new_[12894]_  | ~\new_[18998]_ );
  assign \new_[5053]_  = ~\new_[6024]_  | (~\new_[9265]_  & ~\new_[19243]_ );
  assign \new_[5054]_  = ~\new_[6030]_  & (~\new_[11451]_  | ~\new_[19098]_ );
  assign \new_[5055]_  = ~\new_[17977]_  | (~\new_[6154]_  & ~\new_[11091]_ );
  assign \new_[5056]_  = ~\new_[5508]_  & (~\new_[13138]_  | ~\new_[18280]_ );
  assign \new_[5057]_  = ~\new_[7393]_  | ~\new_[6031]_ ;
  assign \new_[5058]_  = ~\new_[5522]_  | ~\new_[19323]_ ;
  assign \new_[5059]_  = ~\new_[19599]_  | (~\new_[6142]_  & ~\new_[8870]_ );
  assign \new_[5060]_  = ~\new_[19445]_  & (~\new_[6143]_  | ~\new_[11174]_ );
  assign \new_[5061]_  = ~\new_[19615]_  | (~\new_[6146]_  & ~\new_[10353]_ );
  assign \new_[5062]_  = ~\new_[9804]_  | ~\new_[6942]_  | ~\new_[15317]_  | ~\new_[9805]_ ;
  assign \new_[5063]_  = ~\new_[5517]_  | ~\new_[19536]_ ;
  assign \new_[5064]_  = ~\new_[10880]_  & ~\new_[5493]_ ;
  assign \new_[5065]_  = ~\new_[19523]_  | (~\new_[6131]_  & ~\new_[12825]_ );
  assign \new_[5066]_  = ~\new_[5518]_  | ~\new_[19339]_ ;
  assign \new_[5067]_  = ~\new_[5519]_  | ~\new_[19318]_ ;
  assign \new_[5068]_  = ~\new_[5520]_  | ~\new_[19120]_ ;
  assign \new_[5069]_  = ~\new_[18599]_  | (~\new_[6134]_  & ~\new_[7282]_ );
  assign \new_[5070]_  = ~\new_[7815]_  | ~\new_[6941]_  | ~\new_[12897]_  | ~\new_[9963]_ ;
  assign \new_[5071]_  = ~\new_[5496]_  & ~\new_[9961]_ ;
  assign \new_[5072]_  = ~\new_[8046]_  | ~\new_[8353]_  | ~\new_[13093]_  | ~\new_[10914]_ ;
  assign \new_[5073]_  = ~\new_[8087]_  | (~\new_[6959]_  & ~\new_[18789]_ );
  assign \new_[5074]_  = ~\new_[8084]_  | (~\new_[6969]_  & ~\new_[19384]_ );
  assign \new_[5075]_  = ~\new_[8085]_  | (~\new_[6970]_  & ~\new_[18769]_ );
  assign \new_[5076]_  = ~\new_[8086]_  | (~\new_[6971]_  & ~\new_[18827]_ );
  assign \new_[5077]_  = ~\new_[8151]_  | ~\new_[10400]_  | ~\new_[12396]_  | ~\new_[8543]_ ;
  assign \new_[5078]_  = ~\new_[6495]_  & (~\new_[6951]_  | ~\new_[18481]_ );
  assign \new_[5079]_  = ~\new_[6128]_  | ~\new_[15824]_ ;
  assign \new_[5080]_  = ~\new_[10734]_  & (~\new_[6966]_  | ~\new_[19145]_ );
  assign \new_[5081]_  = ~\new_[8201]_  & (~\new_[6967]_  | ~\new_[18124]_ );
  assign \new_[5082]_  = ~\new_[6125]_  | (~\new_[6690]_  & ~\new_[19357]_ );
  assign \new_[5083]_  = \new_[8185]_  | \new_[13672]_  | \new_[11973]_  | \new_[11039]_ ;
  assign \new_[5084]_  = ~\new_[8110]_  | ~\new_[13747]_  | ~\new_[10061]_  | ~\new_[10044]_ ;
  assign \new_[5085]_  = \new_[6130]_  & \new_[12204]_ ;
  assign \new_[5086]_  = ~\new_[6141]_  | ~\new_[19528]_ ;
  assign \new_[5087]_  = ~\new_[1033]_  | (~\new_[8466]_  & ~\new_[6978]_ );
  assign \new_[5088]_  = ~\new_[6116]_  | ~\new_[12595]_ ;
  assign \new_[5089]_  = ~\new_[8153]_  | ~\new_[11272]_  | ~\new_[21025]_  | ~\new_[7517]_ ;
  assign \new_[5090]_  = ~\new_[10918]_  | ~\new_[11820]_  | ~\new_[6926]_ ;
  assign \new_[5091]_  = ~\new_[6133]_  | ~\new_[15602]_ ;
  assign \new_[5092]_  = ~\new_[5510]_ ;
  assign \new_[5093]_  = ~\new_[8679]_  | ~\new_[9323]_  | ~\new_[6686]_  | ~\new_[6685]_ ;
  assign \new_[5094]_  = ~\new_[6561]_  | (~\new_[6986]_  & ~\new_[1878]_ );
  assign \new_[5095]_  = ~\new_[6572]_  | (~\new_[6990]_  & ~\new_[18594]_ );
  assign \new_[5096]_  = ~\new_[9826]_  | ~\new_[9552]_  | ~\new_[8079]_  | ~\new_[9806]_ ;
  assign \new_[5097]_  = ~\new_[9892]_  | ~\new_[9591]_  | ~\new_[8082]_  | ~\new_[9858]_ ;
  assign \new_[5098]_  = ~\new_[6160]_  & (~\new_[7008]_  | ~\new_[19751]_ );
  assign \new_[5099]_  = ~\new_[10772]_  & (~\new_[6999]_  | ~\new_[19439]_ );
  assign \new_[5100]_  = ~\new_[14619]_  | ~\new_[8071]_  | ~\new_[10792]_  | ~\new_[10917]_ ;
  assign \new_[5101]_  = (~\new_[6984]_  | ~\new_[19070]_ ) & (~\new_[8813]_  | ~\new_[19377]_ );
  assign \new_[5102]_  = (~\new_[6988]_  | ~\new_[1878]_ ) & (~\new_[10978]_  | ~\new_[19507]_ );
  assign \new_[5103]_  = ~\new_[9966]_  | ~\new_[8055]_  | ~\new_[8530]_  | ~\new_[11503]_ ;
  assign \new_[5104]_  = ~\new_[11030]_  | ~\new_[8059]_  | ~\new_[9654]_  | ~\new_[11004]_ ;
  assign \new_[5105]_  = ~\new_[7796]_  | ~\new_[9657]_  | ~\new_[8060]_  | ~\new_[20705]_ ;
  assign \new_[5106]_  = ~\new_[6137]_  | (~\new_[7001]_  & ~\new_[19022]_ );
  assign \new_[5107]_  = ~\new_[19740]_  | (~\new_[7566]_  & ~\new_[7226]_ );
  assign \new_[5108]_  = ~\new_[6273]_  | ~\new_[19561]_ ;
  assign \new_[5109]_  = ~\new_[19336]_  | (~\new_[7218]_  & ~\new_[9602]_ );
  assign \new_[5110]_  = ~\new_[19702]_  | (~\new_[7491]_  & ~\new_[7219]_ );
  assign \new_[5111]_  = ~\new_[1039]_  | (~\new_[7122]_  & ~\new_[8215]_ );
  assign \new_[5112]_  = ~\new_[19619]_  | (~\new_[7233]_  & ~\new_[9046]_ );
  assign \new_[5113]_  = ~\new_[19318]_  | (~\new_[8213]_  & ~\new_[7176]_ );
  assign \new_[5114]_  = ~\new_[19748]_  | (~\new_[7231]_  & ~\new_[6886]_ );
  assign \new_[5115]_  = ~\new_[19453]_  | (~\new_[7090]_  & ~\new_[9698]_ );
  assign \new_[5116]_  = ~\new_[19659]_  | (~\new_[7264]_  & ~\new_[8765]_ );
  assign \new_[5117]_  = ~\new_[19441]_  | (~\new_[7133]_  & ~\new_[10781]_ );
  assign \new_[5118]_  = ~\new_[19300]_  | (~\new_[7164]_  & ~\new_[9740]_ );
  assign \new_[5119]_  = ~\new_[19170]_  | (~\new_[7281]_  & ~\new_[9946]_ );
  assign \new_[5120]_  = \new_[6189]_  & \new_[7754]_ ;
  assign \new_[5121]_  = ~\new_[19088]_  & (~\new_[6883]_  | ~\new_[8090]_ );
  assign \new_[5122]_  = ~\new_[10392]_  | (~\new_[7059]_  & ~\new_[18827]_ );
  assign \new_[5123]_  = ~\new_[7038]_  & ~\new_[12538]_  & ~\new_[15218]_ ;
  assign \new_[5124]_  = ~\new_[19450]_  & (~\new_[6868]_  | ~\new_[7074]_ );
  assign \new_[5125]_  = ~\new_[973]_  | (~\new_[7046]_  & ~\new_[8625]_ );
  assign \new_[5126]_  = ~\new_[18895]_  | (~\new_[7047]_  & ~\new_[6817]_ );
  assign \new_[5127]_  = ~\new_[960]_  | (~\new_[7048]_  & ~\new_[7619]_ );
  assign \new_[5128]_  = ~\new_[6187]_  | ~\new_[18194]_ ;
  assign \new_[5129]_  = ~\new_[19378]_  | (~\new_[7051]_  & ~\new_[8634]_ );
  assign \new_[5130]_  = ~\new_[19530]_  | (~\new_[7055]_  & ~\new_[6777]_ );
  assign \new_[5131]_  = ~\new_[959]_  | (~\new_[7058]_  & ~\new_[9739]_ );
  assign \new_[5132]_  = ~\new_[19512]_  | (~\new_[7063]_  & ~\new_[7720]_ );
  assign \new_[5133]_  = ~\new_[18983]_  | (~\new_[7065]_  & ~\new_[9759]_ );
  assign \new_[5134]_  = ~\new_[1026]_  | (~\new_[7054]_  & ~\new_[7723]_ );
  assign \new_[5135]_  = ~\new_[19813]_  & (~\new_[8311]_  | ~\new_[7213]_ );
  assign \new_[5136]_  = ~\new_[9799]_  | ~\new_[8310]_  | ~\new_[11083]_  | ~\new_[8738]_ ;
  assign \new_[5137]_  = (~\new_[7244]_  | ~\new_[19659]_ ) & (~\new_[12837]_  | ~\new_[17478]_ );
  assign \new_[5138]_  = ~\new_[7082]_  | ~\new_[8611]_  | ~\new_[10290]_ ;
  assign \new_[5139]_  = (~\new_[7245]_  | ~\new_[19787]_ ) & (~\new_[13141]_  | ~\new_[17629]_ );
  assign \new_[5140]_  = ~\new_[10021]_  | ~\new_[12901]_  | ~\new_[7247]_ ;
  assign \new_[5141]_  = ~\new_[6235]_  | ~\new_[19284]_ ;
  assign \new_[5142]_  = ~\new_[18998]_  & (~\new_[7089]_  | ~\new_[13766]_ );
  assign \new_[5143]_  = ~\new_[12309]_  | ~\new_[6185]_  | ~\new_[10909]_ ;
  assign \new_[5144]_  = ~\new_[9926]_  | ~\new_[8487]_  | ~\new_[10055]_  | ~\new_[21547]_ ;
  assign \new_[5145]_  = ~\new_[19599]_  & (~\new_[8423]_  | ~\new_[7215]_ );
  assign \new_[5146]_  = ~\new_[8728]_  & (~\new_[7214]_  | ~\new_[19780]_ );
  assign \new_[5147]_  = ~\new_[19547]_  & (~\new_[7136]_  | ~\new_[13979]_ );
  assign \new_[5148]_  = ~\new_[13564]_  & (~\new_[7227]_  | ~\new_[18965]_ );
  assign \new_[5149]_  = ~\new_[13510]_  | ~\new_[12726]_  | ~\new_[8366]_  | ~\new_[13743]_ ;
  assign \new_[5150]_  = ~\new_[9865]_  | ~\new_[8430]_  | ~\new_[11178]_  | ~\new_[8761]_ ;
  assign \new_[5151]_  = ~\new_[7488]_  | ~\new_[15102]_  | ~\new_[12601]_  | ~\new_[11870]_ ;
  assign \new_[5152]_  = ~\new_[7368]_  | ~\new_[7458]_  | ~\new_[7252]_ ;
  assign \new_[5153]_  = ~\new_[8689]_  | ~\new_[8113]_  | ~\new_[12307]_  | ~\new_[14340]_ ;
  assign \new_[5154]_  = ~\new_[8615]_  | ~\new_[7108]_  | ~\new_[10142]_ ;
  assign \new_[5155]_  = ~\new_[7070]_  | ~\new_[9137]_  | ~\new_[14319]_ ;
  assign \new_[5156]_  = ~\new_[19115]_  & (~\new_[7194]_  | ~\new_[13763]_ );
  assign \new_[5157]_  = \new_[6192]_  & \new_[8389]_ ;
  assign \new_[5158]_  = ~\new_[8390]_  | ~\new_[15034]_  | ~\new_[12596]_  | ~\new_[14070]_ ;
  assign \new_[5159]_  = ~\new_[6178]_  & (~\new_[9354]_  | ~\new_[19239]_ );
  assign \new_[5160]_  = ~\new_[6272]_  | ~\new_[8387]_ ;
  assign \new_[5161]_  = ~\new_[7043]_  | ~\new_[10177]_  | ~\new_[6768]_ ;
  assign \new_[5162]_  = ~\new_[10573]_  | ~\new_[13615]_  | ~\new_[7225]_ ;
  assign \new_[5163]_  = ~\new_[12657]_  | ~\new_[10537]_  | ~\new_[8411]_  | ~\new_[10596]_ ;
  assign \new_[5164]_  = ~\new_[6180]_  & (~\new_[9360]_  | ~\new_[18998]_ );
  assign \new_[5165]_  = ~\new_[6242]_  | ~\new_[19022]_ ;
  assign \new_[5166]_  = (~\new_[7243]_  | ~\new_[19623]_ ) & (~\new_[14404]_  | ~\new_[18300]_ );
  assign \new_[5167]_  = ~\new_[9315]_  | ~\new_[11201]_  | ~\new_[6763]_ ;
  assign \new_[5168]_  = ~\new_[9975]_  | ~\new_[8312]_  | ~\new_[11211]_  | ~\new_[13361]_ ;
  assign \new_[5169]_  = ~\new_[18844]_  | (~\new_[7067]_  & ~\new_[13084]_ );
  assign \new_[5170]_  = ~\new_[19300]_  | (~\new_[7062]_  & ~\new_[10017]_ );
  assign \new_[5171]_  = ~\new_[11425]_  & ~\new_[6161]_ ;
  assign \new_[5172]_  = ~\new_[7035]_  | ~\new_[7897]_  | ~\new_[10613]_ ;
  assign \new_[5173]_  = ~\new_[7232]_  | ~\new_[15736]_  | ~\new_[11907]_ ;
  assign \new_[5174]_  = ~\new_[19523]_  | (~\new_[7057]_  & ~\new_[13049]_ );
  assign \new_[5175]_  = (~\new_[7269]_  | ~\new_[19170]_ ) & (~\new_[11918]_  | ~\new_[17663]_ );
  assign \new_[5176]_  = ~\new_[11260]_  | ~\new_[8072]_  | ~\new_[6784]_ ;
  assign \new_[5177]_  = ~\new_[6246]_  | ~\new_[21417]_ ;
  assign \new_[5178]_  = ~\new_[7044]_  | ~\new_[9030]_  | ~\new_[7685]_ ;
  assign \new_[5179]_  = ~\new_[6243]_  | ~\new_[18344]_ ;
  assign \new_[5180]_  = ~\new_[9369]_  | ~\new_[9634]_  | ~\new_[6798]_ ;
  assign \new_[5181]_  = ~\new_[8073]_  | ~\new_[11291]_  | ~\new_[6797]_ ;
  assign \new_[5182]_  = ~\new_[19523]_  | (~\new_[8527]_  & ~\new_[7061]_ );
  assign \new_[5183]_  = ~\new_[5585]_ ;
  assign \new_[5184]_  = ~\new_[8074]_  | ~\new_[9067]_  | ~\new_[6802]_ ;
  assign \new_[5185]_  = ~\new_[6248]_  | ~\new_[19504]_ ;
  assign \new_[5186]_  = ~\new_[21630]_  | (~\new_[9641]_  & ~\new_[7172]_ );
  assign \new_[5187]_  = ~\new_[9322]_  | ~\new_[10291]_  | ~\new_[6806]_ ;
  assign \new_[5188]_  = ~\new_[7234]_  & ~\new_[16334]_  & ~\new_[11912]_ ;
  assign \new_[5189]_  = ~\new_[6252]_  | ~\new_[19512]_ ;
  assign \new_[5190]_  = ~\new_[6253]_  | ~\new_[18538]_ ;
  assign \new_[5191]_  = ~\new_[8076]_  | ~\new_[10060]_  | ~\new_[6821]_ ;
  assign \new_[5192]_  = ~\new_[6225]_  | ~\new_[19424]_ ;
  assign \new_[5193]_  = ~\new_[5590]_ ;
  assign \new_[5194]_  = ~\new_[6277]_  | ~\new_[18341]_ ;
  assign \new_[5195]_  = (~\new_[7287]_  | ~\new_[19271]_ ) & (~\new_[13066]_  | ~\new_[18525]_ );
  assign \new_[5196]_  = ~\new_[19492]_  | (~\new_[7203]_  & ~\new_[11706]_ );
  assign \new_[5197]_  = ~\new_[5597]_ ;
  assign \new_[5198]_  = ~\new_[8651]_  & ~\new_[6200]_ ;
  assign \new_[5199]_  = ~\new_[7770]_  | ~\new_[9903]_  | ~\new_[10604]_  | ~\new_[7907]_ ;
  assign \new_[5200]_  = ~\new_[19032]_  | (~\new_[7096]_  & ~\new_[14377]_ );
  assign \new_[5201]_  = ~\new_[19179]_  | (~\new_[7084]_  & ~\new_[15223]_ );
  assign \new_[5202]_  = ~\new_[6182]_  | ~\new_[19378]_ ;
  assign \new_[5203]_  = ~\new_[21079]_  & (~\new_[11167]_  | ~\new_[19599]_ );
  assign \new_[5204]_  = ~\new_[19341]_  | (~\new_[7092]_  & ~\new_[15152]_ );
  assign \new_[5205]_  = ~\new_[9703]_  & (~\new_[7321]_  | ~\new_[2500]_ );
  assign \new_[5206]_  = ~\new_[14845]_  & (~\new_[7093]_  | ~\new_[17475]_ );
  assign \new_[5207]_  = ~\new_[8268]_  | ~\new_[8288]_  | ~\new_[10064]_  | ~\new_[12316]_ ;
  assign \new_[5208]_  = ~\new_[8295]_  | ~\new_[10092]_  | ~\new_[9523]_  | ~\new_[8577]_ ;
  assign \new_[5209]_  = ~\new_[13730]_  & (~\new_[7106]_  | ~\new_[19377]_ );
  assign \new_[5210]_  = (~\new_[7113]_  | ~\new_[18187]_ ) & (~\new_[16638]_  | ~\new_[19520]_ );
  assign \new_[5211]_  = ~\new_[13966]_  & (~\new_[7138]_  | ~\new_[19440]_ );
  assign \new_[5212]_  = ~\new_[15121]_  & (~\new_[7124]_  | ~\new_[17447]_ );
  assign \new_[5213]_  = ~\new_[19532]_  & (~\new_[7259]_  | ~\new_[16114]_ );
  assign \new_[5214]_  = ~\new_[19032]_  & (~\new_[7334]_  | ~\new_[9817]_ );
  assign \new_[5215]_  = ~\new_[9579]_  | ~\new_[7585]_  | ~\new_[8278]_  | ~\new_[15065]_ ;
  assign \new_[5216]_  = ~\new_[19170]_  | (~\new_[7142]_  & ~\new_[11906]_ );
  assign \new_[5217]_  = ~\new_[19483]_  & (~\new_[7336]_  | ~\new_[10964]_ );
  assign \new_[5218]_  = ~\new_[19433]_  | (~\new_[7338]_  & ~\new_[10985]_ );
  assign \new_[5219]_  = ~\new_[6549]_  | ~\new_[6214]_ ;
  assign \new_[5220]_  = ~\new_[19157]_  | (~\new_[7187]_  & ~\new_[15288]_ );
  assign \new_[5221]_  = ~\new_[18599]_  | (~\new_[7339]_  & ~\new_[10984]_ );
  assign \new_[5222]_  = ~\new_[6217]_  | ~\new_[922]_ ;
  assign \new_[5223]_  = ~\new_[6220]_  | ~\new_[18293]_ ;
  assign \new_[5224]_  = ~\new_[6221]_  | ~\new_[19529]_ ;
  assign \new_[5225]_  = ~\new_[11071]_  & ~\new_[6222]_ ;
  assign \new_[5226]_  = ~\new_[9453]_  & ~\new_[6148]_ ;
  assign \new_[5227]_  = (~\new_[7323]_  | ~\new_[19440]_ ) & (~\new_[10239]_  | ~\new_[19366]_ );
  assign \new_[5228]_  = (~\new_[7324]_  | ~\new_[19177]_ ) & (~\new_[10158]_  | ~\new_[18998]_ );
  assign \new_[5229]_  = (~\new_[7320]_  | ~\new_[19492]_ ) & (~\new_[7884]_  | ~\new_[19088]_ );
  assign \new_[5230]_  = ~\new_[5619]_ ;
  assign \new_[5231]_  = (~\new_[7267]_  | ~\new_[19179]_ ) & (~\new_[11190]_  | ~\new_[19687]_ );
  assign \new_[5232]_  = ~\new_[5620]_ ;
  assign \new_[5233]_  = ~\new_[9458]_  & ~\new_[6150]_ ;
  assign \new_[5234]_  = ~\new_[5621]_ ;
  assign \new_[5235]_  = ~\new_[7529]_  & (~\new_[7328]_  | ~\new_[20098]_ );
  assign \new_[5236]_  = (~\new_[7329]_  | ~\new_[17668]_ ) & (~\new_[10018]_  | ~\new_[19711]_ );
  assign \new_[5237]_  = (~\new_[7330]_  | ~\new_[19491]_ ) & (~\new_[7952]_  | ~\new_[19592]_ );
  assign \new_[5238]_  = ~\new_[9398]_  & (~\new_[7110]_  | ~\new_[18762]_ );
  assign \new_[5239]_  = ~\new_[9403]_  & (~\new_[7144]_  | ~\new_[19208]_ );
  assign \new_[5240]_  = ~\new_[6184]_  & (~\new_[15824]_  | ~\new_[11653]_ );
  assign \new_[5241]_  = ~\new_[6197]_  & (~\new_[15602]_  | ~\new_[11722]_ );
  assign \new_[5242]_  = (~\new_[7154]_  | ~\new_[17801]_ ) & (~\new_[15865]_  | ~\new_[11551]_ );
  assign \new_[5243]_  = ~\new_[8241]_  | ~\new_[14303]_  | ~\new_[10050]_  | ~\new_[13554]_ ;
  assign \new_[5244]_  = ~\new_[10654]_  | ~\new_[9551]_  | ~\new_[7315]_ ;
  assign \new_[5245]_  = ~\new_[12003]_  | ~\new_[8507]_  | ~\new_[7317]_ ;
  assign \new_[5246]_  = ~\new_[10929]_  | ~\new_[12355]_  | ~\new_[7253]_ ;
  assign \new_[5247]_  = ~\new_[10942]_  | ~\new_[12322]_  | ~\new_[7256]_ ;
  assign \new_[5248]_  = ~\new_[12190]_  | ~\new_[11117]_  | ~\new_[7262]_ ;
  assign \new_[5249]_  = ~\new_[8245]_  | ~\new_[13168]_  | ~\new_[8957]_  | ~\new_[15081]_ ;
  assign \new_[5250]_  = ~\new_[8248]_  | ~\new_[13174]_  | ~\new_[7958]_  | ~\new_[11623]_ ;
  assign \new_[5251]_  = ~\new_[6577]_  | ~\new_[19271]_ ;
  assign \new_[5252]_  = ~\new_[6580]_  | ~\new_[19504]_ ;
  assign \new_[5253]_  = ~\new_[19032]_  | (~\new_[8943]_  & ~\new_[6849]_ );
  assign \new_[5254]_  = ~\new_[18641]_  & (~\new_[7582]_  | ~\new_[7388]_ );
  assign \new_[5255]_  = ~\new_[6457]_  | ~\new_[19326]_ ;
  assign \new_[5256]_  = ~\new_[6586]_  | ~\new_[19787]_ ;
  assign \new_[5257]_  = ~\new_[19530]_  & (~\new_[10231]_  | ~\new_[7360]_ );
  assign \new_[5258]_  = ~\new_[19051]_  | (~\new_[9021]_  & ~\new_[6850]_ );
  assign \new_[5259]_  = ~\new_[922]_  & (~\new_[6704]_  | ~\new_[7546]_ );
  assign \new_[5260]_  = ~\new_[19529]_  & (~\new_[7394]_  | ~\new_[6717]_ );
  assign \new_[5261]_  = ~\new_[6536]_  | ~\new_[19578]_ ;
  assign \new_[5262]_  = ~\new_[6496]_  | ~\new_[19561]_ ;
  assign \new_[5263]_  = ~\new_[5643]_ ;
  assign \new_[5264]_  = ~\new_[5645]_ ;
  assign \new_[5265]_  = ~\new_[19271]_  | (~\new_[7597]_  & ~\new_[6847]_ );
  assign \new_[5266]_  = ~\new_[20641]_  | (~\new_[9613]_  & ~\new_[6848]_ );
  assign \new_[5267]_  = ~\new_[6528]_  | ~\new_[984]_ ;
  assign \new_[5268]_  = ~\new_[6531]_  | ~\new_[19424]_ ;
  assign \new_[5269]_  = ~\new_[19578]_  | (~\new_[6834]_  & ~\new_[9516]_ );
  assign \new_[5270]_  = ~\new_[18649]_  & (~\new_[6824]_  | ~\new_[11041]_ );
  assign \new_[5271]_  = ~\new_[19453]_  & (~\new_[6758]_  | ~\new_[9829]_ );
  assign \new_[5272]_  = ~\new_[19717]_  | (~\new_[6835]_  & ~\new_[10805]_ );
  assign \new_[5273]_  = ~\new_[19787]_  | (~\new_[6785]_  & ~\new_[8776]_ );
  assign \new_[5274]_  = ~\new_[946]_  & (~\new_[6788]_  | ~\new_[21349]_ );
  assign \new_[5275]_  = ~\new_[19600]_  | (~\new_[6799]_  & ~\new_[8790]_ );
  assign \new_[5276]_  = ~\new_[21417]_  & (~\new_[6803]_  | ~\new_[9938]_ );
  assign \new_[5277]_  = ~\new_[6413]_  | ~\new_[19236]_ ;
  assign \new_[5278]_  = ~\new_[19271]_  | (~\new_[6935]_  & ~\new_[6833]_ );
  assign \new_[5279]_  = ~\new_[6593]_  | ~\new_[1039]_ ;
  assign \new_[5280]_  = ~\new_[6595]_  | ~\new_[19318]_ ;
  assign \new_[5281]_  = ~\new_[18757]_  & (~\new_[6715]_  | ~\new_[8594]_ );
  assign \new_[5282]_  = ~\new_[6347]_  | ~\new_[19204]_ ;
  assign \new_[5283]_  = \new_[18749]_  ^ \new_[7337]_ ;
  assign \new_[5284]_  = ~\new_[19377]_  & (~\new_[7404]_  | ~\new_[12718]_ );
  assign \new_[5285]_  = ~\new_[6362]_  | ~\new_[19088]_ ;
  assign \new_[5286]_  = ~\new_[19072]_  | (~\new_[7417]_  & ~\new_[12813]_ );
  assign \new_[5287]_  = \new_[18835]_  ^ \new_[7347]_ ;
  assign \new_[5288]_  = ~\new_[6431]_  | ~\new_[17689]_ ;
  assign \new_[5289]_  = ~\new_[6386]_  | ~\new_[14951]_ ;
  assign \new_[5290]_  = ~\new_[6399]_  | ~\new_[18937]_ ;
  assign \new_[5291]_  = ~\new_[5690]_ ;
  assign \new_[5292]_  = ~\new_[6445]_  | ~\new_[18941]_ ;
  assign \new_[5293]_  = ~\new_[5698]_ ;
  assign \new_[5294]_  = \new_[6473]_  | \new_[20725]_ ;
  assign \new_[5295]_  = ~\new_[6475]_  & ~\new_[7389]_ ;
  assign \new_[5296]_  = ~\new_[6477]_  | ~\new_[18506]_ ;
  assign \new_[5297]_  = ~\new_[6484]_  | ~\new_[19578]_ ;
  assign \new_[5298]_  = ~\new_[19640]_  | (~\new_[7412]_  & ~\new_[7859]_ );
  assign \new_[5299]_  = ~\new_[5704]_ ;
  assign \new_[5300]_  = ~\new_[19029]_  | (~\new_[8381]_  & ~\new_[6786]_ );
  assign \new_[5301]_  = ~\new_[19813]_  | (~\new_[6912]_  & ~\new_[9533]_ );
  assign \new_[5302]_  = ~\new_[6371]_  & ~\new_[14330]_ ;
  assign \new_[5303]_  = \new_[6489]_  | \new_[18668]_ ;
  assign \new_[5304]_  = ~\new_[6490]_  | ~\new_[20679]_ ;
  assign \new_[5305]_  = ~\new_[20763]_  & (~\new_[6702]_  | ~\new_[8443]_ );
  assign \new_[5306]_  = \new_[6494]_  | \new_[20622]_ ;
  assign \new_[5307]_  = \new_[6529]_  & \new_[12339]_ ;
  assign \new_[5308]_  = ~\new_[6591]_  | ~\new_[19237]_ ;
  assign \new_[5309]_  = ~\new_[11128]_  & (~\new_[6739]_  | ~\new_[19553]_ );
  assign \new_[5310]_  = ~\new_[6584]_  & ~\new_[19659]_ ;
  assign \new_[5311]_  = ~\new_[6488]_  & ~\new_[11954]_ ;
  assign \new_[5312]_  = ~\new_[19384]_  | (~\new_[7442]_  & ~\new_[7669]_ );
  assign \new_[5313]_  = ~\new_[6652]_  & (~\new_[8457]_  | ~\new_[17472]_ );
  assign \new_[5314]_  = ~\new_[7443]_  | ~\new_[14163]_  | ~\new_[6892]_ ;
  assign \new_[5315]_  = ~\new_[19599]_  | (~\new_[7450]_  & ~\new_[7908]_ );
  assign \new_[5316]_  = ~\new_[6400]_  | ~\new_[17723]_ ;
  assign \new_[5317]_  = ~\new_[19787]_  | (~\new_[7451]_  & ~\new_[8993]_ );
  assign \new_[5318]_  = ~\new_[5729]_ ;
  assign \new_[5319]_  = ~\new_[7454]_  | ~\new_[9608]_  | ~\new_[8661]_ ;
  assign \new_[5320]_  = ~\new_[6506]_  | ~\new_[21273]_ ;
  assign \new_[5321]_  = ~\new_[6508]_  & ~\new_[9298]_ ;
  assign \new_[5322]_  = ~\new_[954]_  | (~\new_[6661]_  & ~\new_[9619]_ );
  assign \new_[5323]_  = ~\new_[6404]_  | ~\new_[7857]_ ;
  assign \new_[5324]_  = ~\new_[19257]_  & (~\new_[6671]_  | ~\new_[6672]_ );
  assign \new_[5325]_  = ~\new_[6512]_  | ~\new_[17796]_ ;
  assign \new_[5326]_  = ~\new_[19341]_  & (~\new_[6679]_  | ~\new_[7497]_ );
  assign \new_[5327]_  = ~\new_[6519]_  | ~\new_[20098]_ ;
  assign \new_[5328]_  = ~\new_[6521]_  & ~\new_[7514]_ ;
  assign \new_[5329]_  = ~\new_[6418]_  | ~\new_[17697]_ ;
  assign \new_[5330]_  = ~\new_[11991]_  | ~\new_[9090]_  | ~\new_[8057]_  | ~\new_[12047]_ ;
  assign \new_[5331]_  = ~\new_[10668]_  | ~\new_[11887]_  | ~\new_[7950]_  | ~\new_[13403]_ ;
  assign \new_[5332]_  = \new_[6589]_  & \new_[18803]_ ;
  assign \new_[5333]_  = ~\new_[6057]_  & (~\new_[8566]_  | ~\new_[18087]_ );
  assign \new_[5334]_  = \new_[6995]_  ^ \new_[18887]_ ;
  assign \new_[5335]_  = ~\new_[10581]_  & (~\new_[8445]_  | ~\new_[17689]_ );
  assign \new_[5336]_  = ~\new_[5759]_ ;
  assign \new_[5337]_  = ~\new_[6532]_  & ~\new_[6720]_ ;
  assign \new_[5338]_  = ~\new_[5761]_ ;
  assign \new_[5339]_  = ~\new_[6491]_  & (~\new_[12679]_  | ~\new_[18209]_ );
  assign \new_[5340]_  = ~\new_[6523]_  & ~\new_[6626]_ ;
  assign \new_[5341]_  = ~\new_[10655]_  | ~\new_[7083]_  | ~\new_[6866]_ ;
  assign \new_[5342]_  = ~\new_[7697]_  & ~\new_[6361]_ ;
  assign \new_[5343]_  = ~\new_[10424]_  | ~\new_[14333]_  | ~\new_[6776]_  | ~\new_[9803]_ ;
  assign \new_[5344]_  = ~\new_[12025]_  | ~\new_[7139]_  | ~\new_[6887]_ ;
  assign \new_[5345]_  = ~\new_[11421]_  | ~\new_[9970]_  | ~\new_[6783]_  | ~\new_[11885]_ ;
  assign \new_[5346]_  = ~\new_[10418]_  | ~\new_[9903]_  | ~\new_[13117]_  | ~\new_[6796]_ ;
  assign \new_[5347]_  = ~\new_[7651]_  | ~\new_[13239]_  | ~\new_[13630]_  | ~\new_[10050]_ ;
  assign \new_[5348]_  = ~\new_[8320]_  | (~\new_[7411]_  & ~\new_[19492]_ );
  assign \new_[5349]_  = ~\new_[6316]_  | ~\new_[1039]_ ;
  assign \new_[5350]_  = ~\new_[9266]_  | ~\new_[7403]_  | ~\new_[7402]_ ;
  assign \new_[5351]_  = ~\new_[9446]_  | ~\new_[6628]_  | ~\new_[6771]_ ;
  assign \new_[5352]_  = ~\new_[10341]_  | ~\new_[8365]_  | ~\new_[6748]_ ;
  assign \new_[5353]_  = ~\new_[18466]_  & (~\new_[6888]_  | ~\new_[11952]_ );
  assign \new_[5354]_  = ~\new_[18249]_  & (~\new_[6752]_  | ~\new_[14195]_ );
  assign \new_[5355]_  = ~\new_[17688]_  & (~\new_[6762]_  | ~\new_[13615]_ );
  assign \new_[5356]_  = ~\new_[6590]_  & (~\new_[13857]_  | ~\new_[19045]_ );
  assign \new_[5357]_  = ~\new_[7302]_  | ~\new_[6381]_ ;
  assign \new_[5358]_  = ~\new_[18863]_  | (~\new_[6795]_  & ~\new_[11745]_ );
  assign \new_[5359]_  = ~\new_[15893]_  & (~\new_[7653]_  | ~\new_[7428]_ );
  assign \new_[5360]_  = ~\new_[7308]_  & (~\new_[6828]_  | ~\new_[19177]_ );
  assign \new_[5361]_  = ~\new_[6552]_  | ~\new_[6387]_ ;
  assign \new_[5362]_  = ~\new_[6324]_  | ~\new_[18808]_ ;
  assign \new_[5363]_  = ~\new_[6328]_  | ~\new_[19318]_ ;
  assign \new_[5364]_  = ~\new_[9265]_  | ~\new_[7439]_  | ~\new_[7438]_ ;
  assign \new_[5365]_  = ~\new_[11929]_  | ~\new_[6314]_ ;
  assign \new_[5366]_  = ~\new_[11923]_  | ~\new_[6315]_ ;
  assign \new_[5367]_  = ~\new_[9273]_  | ~\new_[6674]_  | ~\new_[6673]_ ;
  assign \new_[5368]_  = ~\new_[6414]_  | ~\new_[8362]_ ;
  assign \new_[5369]_  = ~\new_[18473]_  & (~\new_[6805]_  | ~\new_[13723]_ );
  assign \new_[5370]_  = ~\new_[8330]_  | ~\new_[6420]_  | ~\new_[13949]_ ;
  assign \new_[5371]_  = ~\new_[8461]_  | ~\new_[6422]_  | ~\new_[12604]_ ;
  assign \new_[5372]_  = ~\new_[18393]_  & (~\new_[6815]_  | ~\new_[14192]_ );
  assign \new_[5373]_  = ~\new_[7452]_  | ~\new_[6426]_  | ~\new_[11509]_ ;
  assign \new_[5374]_  = ~\new_[18171]_  & (~\new_[6818]_  | ~\new_[12929]_ );
  assign \new_[5375]_  = ~\new_[6583]_  & (~\new_[13790]_  | ~\new_[19177]_ );
  assign \new_[5376]_  = ~\new_[6582]_  & (~\new_[12563]_  | ~\new_[18655]_ );
  assign \new_[5377]_  = ~\new_[12816]_  | ~\new_[7396]_  | ~\new_[7395]_ ;
  assign \new_[5378]_  = ~\new_[12806]_  & (~\new_[6730]_  | ~\new_[18714]_ );
  assign \new_[5379]_  = ~\new_[11723]_  & ~\new_[6307]_ ;
  assign \new_[5380]_  = ~\new_[6603]_  & ~\new_[7217]_ ;
  assign \new_[5381]_  = ~\new_[10107]_  | ~\new_[7599]_  | ~\new_[6831]_ ;
  assign \new_[5382]_  = ~\new_[6606]_  | ~\new_[15777]_ ;
  assign \new_[5383]_  = ~\new_[6063]_  & ~\new_[8161]_ ;
  assign \new_[5384]_  = ~\new_[17663]_  | (~\new_[7437]_  & ~\new_[11905]_ );
  assign \new_[5385]_  = ~\new_[15822]_  | (~\new_[6808]_  & ~\new_[14040]_ );
  assign \new_[5386]_  = ~\new_[6439]_  | ~\new_[17977]_ ;
  assign \new_[5387]_  = ~\new_[17478]_  | (~\new_[6723]_  & ~\new_[13254]_ );
  assign \new_[5388]_  = ~\new_[6366]_  & (~\new_[15737]_  | ~\new_[17292]_ );
  assign \new_[5389]_  = ~\new_[6374]_  & (~\new_[16545]_  | ~\new_[17792]_ );
  assign \new_[5390]_  = ~\new_[6649]_  & ~\new_[6299]_ ;
  assign \new_[5391]_  = ~\new_[6040]_  & ~\new_[6305]_ ;
  assign \new_[5392]_  = ~\new_[6721]_  & ~\new_[6306]_ ;
  assign \new_[5393]_  = ~\new_[5833]_ ;
  assign \new_[5394]_  = ~\new_[9618]_  & ~\new_[6458]_ ;
  assign \new_[5395]_  = ~\new_[9848]_  | ~\new_[13059]_  | ~\new_[10420]_  | ~\new_[6878]_ ;
  assign \new_[5396]_  = ~\new_[14232]_  | (~\new_[6836]_  & ~\new_[18569]_ );
  assign \new_[5397]_  = ~\new_[13165]_  | (~\new_[6839]_  & ~\new_[19247]_ );
  assign \new_[5398]_  = ~\new_[15329]_  | (~\new_[6840]_  & ~\new_[21629]_ );
  assign \new_[5399]_  = (~\new_[6842]_  | ~\new_[19088]_ ) & (~\new_[12749]_  | ~\new_[18166]_ );
  assign \new_[5400]_  = ~\new_[7946]_  | ~\new_[6280]_ ;
  assign \new_[5401]_  = (~\new_[6845]_  | ~\new_[19727]_ ) & (~\new_[13740]_  | ~\new_[19319]_ );
  assign \new_[5402]_  = (~\new_[6843]_  | ~\new_[19115]_ ) & (~\new_[16247]_  | ~\new_[18209]_ );
  assign \new_[5403]_  = (~\new_[6844]_  | ~\new_[18194]_ ) & (~\new_[16155]_  | ~\new_[18414]_ );
  assign \new_[5404]_  = ~\new_[7886]_  | ~\new_[6284]_ ;
  assign \new_[5405]_  = (~\new_[6846]_  | ~\new_[19247]_ ) & (~\new_[12667]_  | ~\new_[18692]_ );
  assign \new_[5406]_  = \new_[6052]_  | \new_[7186]_ ;
  assign \new_[5407]_  = \new_[6388]_  & \new_[8061]_ ;
  assign \new_[5408]_  = \new_[8850]_  & \new_[6352]_ ;
  assign \new_[5409]_  = ~\new_[6607]_  | ~\new_[14955]_ ;
  assign \new_[5410]_  = ~\new_[9800]_  & (~\new_[6740]_  | ~\new_[17734]_ );
  assign \new_[5411]_  = ~\new_[9968]_  & (~\new_[6764]_  | ~\new_[18332]_ );
  assign \new_[5412]_  = ~\new_[8969]_  | ~\new_[6397]_ ;
  assign \new_[5413]_  = \new_[10361]_  & \new_[6440]_ ;
  assign \new_[5414]_  = \new_[10399]_  & \new_[6452]_ ;
  assign \new_[5415]_  = ~\new_[9938]_  | ~\new_[6514]_  | ~\new_[8503]_ ;
  assign \new_[5416]_  = ~\new_[11041]_  | ~\new_[6486]_  | ~\new_[9486]_ ;
  assign \new_[5417]_  = ~\new_[6288]_  | ~\new_[6403]_ ;
  assign \new_[5418]_  = (~\new_[6680]_  | ~\new_[18280]_ ) & (~\new_[8250]_  | ~\new_[18739]_ );
  assign \new_[5419]_  = ~\new_[19323]_  & (~\new_[6765]_  | ~\new_[10875]_ );
  assign \new_[5420]_  = \new_[6076]_  | \new_[18787]_ ;
  assign \new_[5421]_  = \new_[6073]_  | \new_[19717]_ ;
  assign \new_[5422]_  = ~\new_[19032]_  & (~\new_[7888]_  | ~\new_[6877]_ );
  assign \new_[5423]_  = ~\new_[19436]_  | (~\new_[9029]_  & ~\new_[6898]_ );
  assign \new_[5424]_  = \new_[6104]_  | \new_[19748]_ ;
  assign \new_[5425]_  = \new_[6105]_  | \new_[18293]_ ;
  assign \new_[5426]_  = \new_[6106]_  | \new_[19659]_ ;
  assign \new_[5427]_  = ~\new_[6627]_  & (~\new_[17015]_  | ~\new_[15971]_ );
  assign \new_[5428]_  = ~\new_[17689]_  & (~\new_[6906]_  | ~\new_[12367]_ );
  assign \new_[5429]_  = ~\new_[6605]_  | ~\new_[15777]_ ;
  assign \new_[5430]_  = \new_[6349]_  | \new_[19529]_ ;
  assign \new_[5431]_  = ~\new_[6101]_  & ~\new_[10892]_ ;
  assign \new_[5432]_  = ~\new_[14005]_  | ~\new_[6853]_  | ~\new_[11207]_ ;
  assign \new_[5433]_  = ~\new_[6624]_  | ~\new_[12657]_ ;
  assign \new_[5434]_  = ~\new_[19072]_  | (~\new_[6927]_  & ~\new_[10599]_ );
  assign \new_[5435]_  = ~\new_[6627]_  & (~\new_[12705]_  | ~\new_[18194]_ );
  assign \new_[5436]_  = ~\new_[18569]_  & (~\new_[11222]_  | ~\new_[6915]_ );
  assign \new_[5437]_  = ~\new_[6067]_  | ~\new_[21631]_ ;
  assign \new_[5438]_  = \new_[6079]_  | \new_[922]_ ;
  assign \new_[5439]_  = ~\new_[5922]_ ;
  assign \new_[5440]_  = ~\new_[10938]_  & ~\new_[6102]_ ;
  assign \new_[5441]_  = ~\new_[21558]_  | (~\new_[6928]_  & ~\new_[10662]_ );
  assign \new_[5442]_  = ~\new_[5929]_ ;
  assign \new_[5443]_  = \new_[6086]_  & \new_[21638]_ ;
  assign \new_[5444]_  = \new_[6088]_  & \new_[19099]_ ;
  assign \new_[5445]_  = \new_[6090]_  | \new_[921]_ ;
  assign \new_[5446]_  = ~\new_[5940]_ ;
  assign \new_[5447]_  = ~\new_[6092]_  | ~\new_[14033]_ ;
  assign \new_[5448]_  = ~\new_[6650]_  | ~\new_[922]_ ;
  assign \new_[5449]_  = ~\new_[6860]_  | ~\new_[9980]_  | ~\new_[12283]_ ;
  assign \new_[5450]_  = ~\new_[6058]_  | ~\new_[19529]_ ;
  assign \new_[5451]_  = ~\new_[6626]_  | ~\new_[921]_ ;
  assign \new_[5452]_  = ~\new_[18361]_  | (~\new_[6929]_  & ~\new_[10642]_ );
  assign \new_[5453]_  = ~\new_[5952]_ ;
  assign \new_[5454]_  = ~\new_[5958]_ ;
  assign \new_[5455]_  = ~\new_[5968]_ ;
  assign \new_[5456]_  = ~\new_[6640]_  | ~\new_[18087]_ ;
  assign \new_[5457]_  = ~\new_[10603]_  | ~\new_[6075]_  | ~\new_[7794]_ ;
  assign \new_[5458]_  = ~\new_[9801]_  | ~\new_[14401]_  | ~\new_[6921]_ ;
  assign \new_[5459]_  = ~\new_[6050]_  | ~\new_[19748]_ ;
  assign \new_[5460]_  = ~\new_[6651]_  | ~\new_[19587]_ ;
  assign \new_[5461]_  = ~\new_[8455]_  & (~\new_[6933]_  | ~\new_[19243]_ );
  assign \new_[5462]_  = \new_[10829]_  | \new_[6611]_ ;
  assign \new_[5463]_  = ~\new_[8398]_  | ~\new_[6608]_ ;
  assign \new_[5464]_  = (~\new_[6769]_  | ~\new_[19578]_ ) & (~\new_[13006]_  | ~\new_[18965]_ );
  assign \new_[5465]_  = ~\new_[8774]_  | ~\new_[6920]_  | ~\new_[13246]_ ;
  assign \new_[5466]_  = ~\new_[5988]_ ;
  assign \new_[5467]_  = ~\new_[9343]_  | ~\new_[6814]_  | ~\new_[6856]_ ;
  assign \new_[5468]_  = \new_[6610]_  & \new_[13832]_ ;
  assign \new_[5469]_  = ~\new_[6059]_  | ~\new_[12898]_ ;
  assign \new_[5470]_  = ~\new_[5996]_ ;
  assign \new_[5471]_  = ~\new_[12778]_  & (~\new_[6881]_  | ~\new_[19520]_ );
  assign \new_[5472]_  = ~\new_[6615]_  & (~\new_[12472]_  | ~\new_[18179]_ );
  assign \new_[5473]_  = ~\new_[18021]_  | (~\new_[6925]_  & ~\new_[11217]_ );
  assign \new_[5474]_  = ~\new_[6069]_  | ~\new_[18701]_ ;
  assign \new_[5475]_  = ~\new_[10611]_  | ~\new_[6034]_ ;
  assign \new_[5476]_  = \new_[8814]_  ? \new_[18941]_  : \new_[12785]_ ;
  assign \new_[5477]_  = ~\new_[11328]_  | ~\new_[6901]_  | ~\new_[6916]_ ;
  assign \new_[5478]_  = ~\new_[6693]_  & ~\new_[6051]_ ;
  assign \new_[5479]_  = ~\new_[8475]_  & ~\new_[6657]_ ;
  assign \new_[5480]_  = ~\new_[20557]_  | ~\new_[12692]_  | ~\new_[7921]_ ;
  assign \new_[5481]_  = ~\new_[6115]_  | ~\new_[19550]_ ;
  assign \new_[5482]_  = ~\new_[6026]_ ;
  assign \new_[5483]_  = ~\new_[10935]_  | ~\new_[8014]_  | ~\new_[15214]_  | ~\new_[9842]_ ;
  assign \new_[5484]_  = ~\new_[9905]_  | ~\new_[8017]_  | ~\new_[14241]_  | ~\new_[9906]_ ;
  assign \new_[5485]_  = ~\new_[8048]_  | ~\new_[13576]_  | ~\new_[9380]_  | ~\new_[10366]_ ;
  assign \new_[5486]_  = ~\new_[7773]_  | ~\new_[8012]_  | ~\new_[10610]_  | ~\new_[9810]_ ;
  assign \new_[5487]_  = ~\new_[10126]_  & (~\new_[6913]_  | ~\new_[15893]_ );
  assign \new_[5488]_  = \new_[6856]_  & \new_[7783]_ ;
  assign \new_[5489]_  = ~\new_[8798]_  & ~\new_[9886]_ ;
  assign \new_[5490]_  = ~\new_[6945]_  | ~\new_[19337]_ ;
  assign \new_[5491]_  = ~\new_[6060]_ ;
  assign \new_[5492]_  = ~\new_[6911]_  | ~\new_[15963]_ ;
  assign \new_[5493]_  = ~\new_[991]_  & (~\new_[8618]_  | ~\new_[8051]_ );
  assign \new_[5494]_  = ~\new_[6064]_ ;
  assign \new_[5495]_  = ~\new_[923]_  | ~\new_[17522]_  | ~\new_[10561]_ ;
  assign \new_[5496]_  = ~\new_[19780]_  & (~\new_[10281]_  | ~\new_[8038]_ );
  assign \new_[5497]_  = ~\new_[6078]_ ;
  assign \new_[5498]_  = ~\new_[922]_  | ~\new_[17972]_  | ~\new_[10514]_ ;
  assign \new_[5499]_  = \new_[6890]_  & \new_[13585]_ ;
  assign \new_[5500]_  = \new_[6880]_  & \new_[12256]_ ;
  assign \new_[5501]_  = \new_[9382]_  | \new_[13487]_  | \new_[13118]_  | \new_[11006]_ ;
  assign \new_[5502]_  = ~\new_[6899]_  & (~\new_[11621]_  | ~\new_[19406]_ );
  assign \new_[5503]_  = ~\new_[6907]_  | ~\new_[13478]_ ;
  assign \new_[5504]_  = ~\new_[6084]_ ;
  assign \new_[5505]_  = \new_[9383]_  | \new_[11185]_  | \new_[14280]_  | \new_[12264]_ ;
  assign \new_[5506]_  = ~\new_[6089]_ ;
  assign \new_[5507]_  = ~\new_[6091]_ ;
  assign \new_[5508]_  = ~\new_[18280]_  & (~\new_[8025]_  | ~\new_[14683]_ );
  assign \new_[5509]_  = ~\new_[9011]_  & ~\new_[6953]_ ;
  assign \new_[5510]_  = ~\new_[10505]_  | (~\new_[10171]_  & ~\new_[18840]_ );
  assign \new_[5511]_  = ~\new_[6857]_  | ~\new_[10586]_ ;
  assign \new_[5512]_  = (~\new_[13342]_  & ~\new_[17980]_ ) | (~\new_[17666]_  & ~\new_[20809]_ );
  assign \new_[5513]_  = (~\new_[13607]_  & ~\new_[17132]_ ) | (~\new_[17512]_  & ~\new_[8041]_ );
  assign \new_[5514]_  = \new_[9386]_  | \new_[10083]_  | \new_[8880]_  | \new_[14156]_ ;
  assign \new_[5515]_  = ~\new_[14928]_  | ~\new_[15037]_  | ~\new_[6987]_  | ~\new_[10658]_ ;
  assign \new_[5516]_  = ~\new_[13464]_  | ~\new_[13848]_  | ~\new_[6989]_  | ~\new_[10643]_ ;
  assign \new_[5517]_  = ~\new_[9723]_  | ~\new_[9314]_  | ~\new_[7640]_  | ~\new_[8947]_ ;
  assign \new_[5518]_  = ~\new_[9730]_  | ~\new_[9318]_  | ~\new_[9598]_  | ~\new_[10216]_ ;
  assign \new_[5519]_  = ~\new_[9742]_  | ~\new_[9320]_  | ~\new_[7690]_  | ~\new_[9049]_ ;
  assign \new_[5520]_  = ~\new_[9722]_  | ~\new_[9321]_  | ~\new_[8677]_  | ~\new_[11303]_ ;
  assign \new_[5521]_  = ~\new_[9832]_  | ~\new_[14986]_  | ~\new_[6979]_  | ~\new_[14542]_ ;
  assign \new_[5522]_  = ~\new_[13603]_  | ~\new_[15130]_  | ~\new_[6980]_  | ~\new_[14485]_ ;
  assign \new_[5523]_  = ~\new_[16922]_  | ~\new_[9316]_  | ~\new_[10374]_  | ~\new_[10962]_ ;
  assign \new_[5524]_  = ~\new_[12227]_  | ~\new_[10371]_  | ~\new_[8047]_ ;
  assign \new_[5525]_  = ~\new_[9303]_  & ~\new_[21115]_ ;
  assign \new_[5526]_  = ~\new_[19659]_  | (~\new_[8175]_  & ~\new_[8862]_ );
  assign \new_[5527]_  = ~\new_[1033]_  | (~\new_[8142]_  & ~\new_[9736]_ );
  assign \new_[5528]_  = ~\new_[19208]_  & (~\new_[7835]_  | ~\new_[8088]_ );
  assign \new_[5529]_  = ~\new_[6121]_ ;
  assign \new_[5530]_  = ~\new_[18606]_  & (~\new_[7938]_  | ~\new_[8089]_ );
  assign \new_[5531]_  = ~\new_[6124]_ ;
  assign \new_[5532]_  = ~\new_[21635]_  & (~\new_[9005]_  | ~\new_[8067]_ );
  assign \new_[5533]_  = ~\new_[19215]_  & (~\new_[9135]_  | ~\new_[8099]_ );
  assign \new_[5534]_  = ~\new_[6958]_  | ~\new_[18998]_ ;
  assign \new_[5535]_  = ~\new_[946]_  | (~\new_[8078]_  & ~\new_[7668]_ );
  assign \new_[5536]_  = ~\new_[11333]_  | ~\new_[8098]_  | ~\new_[12890]_ ;
  assign \new_[5537]_  = ~\new_[7003]_  | ~\new_[19517]_ ;
  assign \new_[5538]_  = ~\new_[8102]_  | ~\new_[8612]_  | ~\new_[10024]_ ;
  assign \new_[5539]_  = ~\new_[8173]_  & ~\new_[15746]_  & ~\new_[11768]_ ;
  assign \new_[5540]_  = ~\new_[12269]_  | ~\new_[9492]_  | ~\new_[12900]_  | ~\new_[11126]_ ;
  assign \new_[5541]_  = ~\new_[19072]_  & (~\new_[8107]_  | ~\new_[12670]_ );
  assign \new_[5542]_  = ~\new_[15097]_  | ~\new_[15305]_  | ~\new_[8224]_ ;
  assign \new_[5543]_  = ~\new_[9509]_  | ~\new_[12811]_  | ~\new_[14598]_  | ~\new_[14087]_ ;
  assign \new_[5544]_  = ~\new_[9829]_  | ~\new_[7014]_  | ~\new_[9547]_ ;
  assign \new_[5545]_  = ~\new_[14079]_  | ~\new_[6977]_  | ~\new_[12329]_ ;
  assign \new_[5546]_  = ~\new_[19441]_  | (~\new_[8080]_  & ~\new_[11781]_ );
  assign \new_[5547]_  = \new_[6950]_  & \new_[7413]_ ;
  assign \new_[5548]_  = ~\new_[7005]_  | ~\new_[19530]_ ;
  assign \new_[5549]_  = ~\new_[9527]_  | ~\new_[12507]_  | ~\new_[12505]_  | ~\new_[21594]_ ;
  assign \new_[5550]_  = ~\new_[8062]_  | ~\new_[6908]_  | ~\new_[10699]_ ;
  assign \new_[5551]_  = ~\new_[12625]_  | ~\new_[11952]_  | ~\new_[8166]_ ;
  assign \new_[5552]_  = ~\new_[7006]_  | ~\new_[19195]_ ;
  assign \new_[5553]_  = ~\new_[8755]_  | ~\new_[9616]_  | ~\new_[11302]_  | ~\new_[14297]_ ;
  assign \new_[5554]_  = ~\new_[13698]_  | ~\new_[12550]_  | ~\new_[9535]_  | ~\new_[11887]_ ;
  assign \new_[5555]_  = ~\new_[8636]_  | ~\new_[9351]_  | ~\new_[11109]_  | ~\new_[14142]_ ;
  assign \new_[5556]_  = ~\new_[21620]_  & (~\new_[8189]_  | ~\new_[19740]_ );
  assign \new_[5557]_  = ~\new_[8091]_  | ~\new_[10109]_  | ~\new_[13466]_ ;
  assign \new_[5558]_  = \new_[8027]_  & \new_[6728]_ ;
  assign \new_[5559]_  = ~\new_[7007]_  | ~\new_[18895]_ ;
  assign \new_[5560]_  = ~\new_[8590]_  | ~\new_[15010]_  | ~\new_[13952]_  | ~\new_[13609]_ ;
  assign \new_[5561]_  = ~\new_[11700]_  | ~\new_[6975]_  | ~\new_[16173]_ ;
  assign \new_[5562]_  = ~\new_[7016]_  | ~\new_[19528]_ ;
  assign \new_[5563]_  = ~\new_[8700]_  | ~\new_[9362]_  | ~\new_[14672]_  | ~\new_[11149]_ ;
  assign \new_[5564]_  = ~\new_[14260]_  & (~\new_[8168]_  | ~\new_[19780]_ );
  assign \new_[5565]_  = ~\new_[9317]_  | ~\new_[9169]_  | ~\new_[7621]_ ;
  assign \new_[5566]_  = ~\new_[12207]_  & (~\new_[8169]_  | ~\new_[19366]_ );
  assign \new_[5567]_  = ~\new_[8092]_  | ~\new_[7895]_  | ~\new_[14051]_ ;
  assign \new_[5568]_  = ~\new_[21559]_  & (~\new_[8195]_  | ~\new_[11591]_ );
  assign \new_[5569]_  = ~\new_[19492]_  & (~\new_[8207]_  | ~\new_[11571]_ );
  assign \new_[5570]_  = ~\new_[8177]_  & ~\new_[16603]_  & ~\new_[13074]_ ;
  assign \new_[5571]_  = ~\new_[959]_  | (~\new_[10830]_  & ~\new_[8170]_ );
  assign \new_[5572]_  = ~\new_[9590]_  | ~\new_[12528]_  | ~\new_[11572]_  | ~\new_[15328]_ ;
  assign \new_[5573]_  = ~\new_[9898]_  | ~\new_[7017]_  | ~\new_[8595]_ ;
  assign \new_[5574]_  = ~\new_[9600]_  | ~\new_[11501]_  | ~\new_[12515]_  | ~\new_[11991]_ ;
  assign \new_[5575]_  = ~\new_[9609]_  | ~\new_[11573]_  | ~\new_[12738]_  | ~\new_[10659]_ ;
  assign \new_[5576]_  = ~\new_[8093]_  | ~\new_[9019]_  | ~\new_[13123]_ ;
  assign \new_[5577]_  = ~\new_[6895]_  | ~\new_[8065]_  | ~\new_[11896]_ ;
  assign \new_[5578]_  = ~\new_[18739]_  & (~\new_[8196]_  | ~\new_[9272]_ );
  assign \new_[5579]_  = ~\new_[12145]_  & (~\new_[8198]_  | ~\new_[19702]_ );
  assign \new_[5580]_  = ~\new_[8094]_  | ~\new_[10254]_  | ~\new_[13145]_ ;
  assign \new_[5581]_  = ~\new_[8511]_  | ~\new_[11701]_  | ~\new_[11605]_  | ~\new_[14109]_ ;
  assign \new_[5582]_  = ~\new_[7806]_  | ~\new_[7018]_  | ~\new_[20348]_ ;
  assign \new_[5583]_  = ~\new_[9899]_  & (~\new_[8199]_  | ~\new_[19600]_ );
  assign \new_[5584]_  = ~\new_[8095]_  | ~\new_[10275]_  | ~\new_[14020]_ ;
  assign \new_[5585]_  = ~\new_[19163]_  & (~\new_[7502]_  | ~\new_[8225]_ );
  assign \new_[5586]_  = ~\new_[8066]_  | ~\new_[7940]_  | ~\new_[8096]_ ;
  assign \new_[5587]_  = ~\new_[8075]_  | ~\new_[9101]_  | ~\new_[7699]_ ;
  assign \new_[5588]_  = ~\new_[21630]_  & (~\new_[8203]_  | ~\new_[12491]_ );
  assign \new_[5589]_  = ~\new_[17668]_  & (~\new_[8204]_  | ~\new_[10530]_ );
  assign \new_[5590]_  = ~\new_[16547]_  | ~\new_[8181]_  | ~\new_[13683]_ ;
  assign \new_[5591]_  = ~\new_[9873]_  & (~\new_[8208]_  | ~\new_[19615]_ );
  assign \new_[5592]_  = ~\new_[19491]_  & (~\new_[8206]_  | ~\new_[11560]_ );
  assign \new_[5593]_  = ~\new_[7009]_  | ~\new_[19442]_ ;
  assign \new_[5594]_  = ~\new_[8160]_  | ~\new_[9026]_  | ~\new_[9147]_ ;
  assign \new_[5595]_  = ~\new_[14863]_  | ~\new_[21132]_  | ~\new_[8584]_  | ~\new_[11363]_ ;
  assign \new_[5596]_  = ~\new_[19005]_  & (~\new_[8209]_  | ~\new_[13975]_ );
  assign \new_[5597]_  = ~\new_[19659]_  & (~\new_[7581]_  | ~\new_[8228]_ );
  assign \new_[5598]_  = ~\new_[8183]_  & ~\new_[15735]_  & ~\new_[12031]_ ;
  assign \new_[5599]_  = ~\new_[19453]_  | (~\new_[8077]_  & ~\new_[12023]_ );
  assign \new_[5600]_  = ~\new_[14194]_  | ~\new_[13723]_  | ~\new_[9548]_  | ~\new_[13561]_ ;
  assign \new_[5601]_  = ~\new_[11826]_  | ~\new_[10976]_  | ~\new_[7205]_  | ~\new_[9056]_ ;
  assign \new_[5602]_  = ~\new_[9497]_  | ~\new_[8583]_  | ~\new_[8265]_  | ~\new_[13793]_ ;
  assign \new_[5603]_  = (~\new_[8159]_  | ~\new_[18965]_ ) & (~\new_[16873]_  | ~\new_[19279]_ );
  assign \new_[5604]_  = ~\new_[9449]_  | ~\new_[10119]_  | ~\new_[7464]_  | ~\new_[9536]_ ;
  assign \new_[5605]_  = (~\new_[8128]_  | ~\new_[18998]_ ) & (~\new_[17509]_  | ~\new_[19408]_ );
  assign \new_[5606]_  = ~\new_[13920]_  | ~\new_[14198]_  | ~\new_[9503]_  | ~\new_[13891]_ ;
  assign \new_[5607]_  = ~\new_[9461]_  | ~\new_[11037]_  | ~\new_[8585]_  | ~\new_[9566]_ ;
  assign \new_[5608]_  = ~\new_[19653]_  & (~\new_[8232]_  | ~\new_[12233]_ );
  assign \new_[5609]_  = ~\new_[10987]_  | ~\new_[12882]_  | ~\new_[8064]_ ;
  assign \new_[5610]_  = ~\new_[6135]_ ;
  assign \new_[5611]_  = ~\new_[8494]_  | ~\new_[8495]_  | ~\new_[9456]_  | ~\new_[13821]_ ;
  assign \new_[5612]_  = ~\new_[15135]_  | ~\new_[20520]_  | ~\new_[8520]_  | ~\new_[16229]_ ;
  assign \new_[5613]_  = ~\new_[19702]_  & (~\new_[8234]_  | ~\new_[12229]_ );
  assign \new_[5614]_  = ~\new_[6968]_  | ~\new_[954]_ ;
  assign \new_[5615]_  = ~\new_[19257]_  & (~\new_[8235]_  | ~\new_[11056]_ );
  assign \new_[5616]_  = ~\new_[19537]_  | (~\new_[8237]_  & ~\new_[13593]_ );
  assign \new_[5617]_  = (~\new_[8186]_  | ~\new_[19550]_ ) & (~\new_[16376]_  | ~\new_[18262]_ );
  assign \new_[5618]_  = (~\new_[8229]_  | ~\new_[19045]_ ) & (~\new_[12422]_  | ~\new_[19547]_ );
  assign \new_[5619]_  = ~\new_[11082]_  | ~\new_[9670]_  | ~\new_[8155]_ ;
  assign \new_[5620]_  = ~\new_[11152]_  | ~\new_[9632]_  | ~\new_[8146]_ ;
  assign \new_[5621]_  = ~\new_[12153]_  | ~\new_[8538]_  | ~\new_[8150]_ ;
  assign \new_[5622]_  = (~\new_[8230]_  | ~\new_[20903]_ ) & (~\new_[11317]_  | ~\new_[17837]_ );
  assign \new_[5623]_  = ~\new_[8805]_  | ~\new_[10769]_  | ~\new_[8370]_  | ~\new_[9833]_ ;
  assign \new_[5624]_  = ~\new_[9404]_  & (~\new_[8144]_  | ~\new_[18606]_ );
  assign \new_[5625]_  = ~\new_[10152]_  & (~\new_[8190]_  | ~\new_[19717]_ );
  assign \new_[5626]_  = (~\new_[8139]_  | ~\new_[17475]_ ) & (~\new_[15353]_  | ~\new_[19508]_ );
  assign \new_[5627]_  = ~\new_[8756]_  | ~\new_[9429]_  | ~\new_[7548]_  | ~\new_[9846]_ ;
  assign \new_[5628]_  = ~\new_[9399]_  | ~\new_[13245]_  | ~\new_[10095]_  | ~\new_[11553]_ ;
  assign \new_[5629]_  = ~\new_[10900]_  | ~\new_[12351]_  | ~\new_[8210]_ ;
  assign \new_[5630]_  = ~\new_[9402]_  | ~\new_[14030]_  | ~\new_[8963]_  | ~\new_[11504]_ ;
  assign \new_[5631]_  = ~\new_[9407]_  | ~\new_[11946]_  | ~\new_[10340]_  | ~\new_[12777]_ ;
  assign \new_[5632]_  = ~\new_[9409]_  | ~\new_[11987]_  | ~\new_[9160]_  | ~\new_[11579]_ ;
  assign \new_[5633]_  = ~\new_[9408]_  | ~\new_[12035]_  | ~\new_[7975]_  | ~\new_[12799]_ ;
  assign \new_[5634]_  = ~\new_[9397]_  | ~\new_[10654]_  | ~\new_[8884]_  | ~\new_[11575]_ ;
  assign \new_[5635]_  = ~\new_[19378]_  & (~\new_[7858]_  | ~\new_[9447]_ );
  assign \new_[5636]_  = ~\new_[7331]_  | ~\new_[19623]_ ;
  assign \new_[5637]_  = ~\new_[946]_  & (~\new_[7848]_  | ~\new_[8732]_ );
  assign \new_[5638]_  = ~\new_[7249]_  | ~\new_[19780]_ ;
  assign \new_[5639]_  = ~\new_[18280]_  | (~\new_[8335]_  & ~\new_[12496]_ );
  assign \new_[5640]_  = ~\new_[17285]_  | (~\new_[8341]_  & ~\new_[13451]_ );
  assign \new_[5641]_  = ~\new_[19088]_  | (~\new_[8348]_  & ~\new_[11506]_ );
  assign \new_[5642]_  = ~\new_[18863]_  | (~\new_[8424]_  & ~\new_[13368]_ );
  assign \new_[5643]_  = ~\new_[1879]_  & (~\new_[8379]_  | ~\new_[7762]_ );
  assign \new_[5644]_  = ~\new_[20763]_  | (~\new_[10809]_  & ~\new_[7760]_ );
  assign \new_[5645]_  = ~\new_[19480]_  & (~\new_[7556]_  | ~\new_[10877]_ );
  assign \new_[5646]_  = ~\new_[6152]_ ;
  assign \new_[5647]_  = ~\new_[7333]_  & (~\new_[15888]_  | ~\new_[16932]_ );
  assign \new_[5648]_  = ~\new_[17381]_  | (~\new_[8431]_  & ~\new_[10565]_ );
  assign \new_[5649]_  = ~\new_[17689]_  | (~\new_[8454]_  & ~\new_[12654]_ );
  assign \new_[5650]_  = ~\new_[17837]_  | (~\new_[7467]_  & ~\new_[12698]_ );
  assign \new_[5651]_  = ~\new_[19257]_  | (~\new_[7469]_  & ~\new_[7763]_ );
  assign \new_[5652]_  = ~\new_[19341]_  | (~\new_[8525]_  & ~\new_[7764]_ );
  assign \new_[5653]_  = ~\new_[19787]_  | (~\new_[7503]_  & ~\new_[7765]_ );
  assign \new_[5654]_  = ~\new_[20513]_  | (~\new_[8536]_  & ~\new_[7766]_ );
  assign \new_[5655]_  = ~\new_[21422]_  | (~\new_[8541]_  & ~\new_[7761]_ );
  assign \new_[5656]_  = ~\new_[19236]_  | (~\new_[7515]_  & ~\new_[7767]_ );
  assign \new_[5657]_  = ~\new_[18498]_  | (~\new_[7538]_  & ~\new_[11641]_ );
  assign \new_[5658]_  = ~\new_[19711]_  | (~\new_[8429]_  & ~\new_[12790]_ );
  assign \new_[5659]_  = ~\new_[19694]_  | (~\new_[7740]_  & ~\new_[8318]_ );
  assign \new_[5660]_  = ~\new_[19271]_  | (~\new_[7632]_  & ~\new_[10991]_ );
  assign \new_[5661]_  = ~\new_[19702]_  | (~\new_[7741]_  & ~\new_[7561]_ );
  assign \new_[5662]_  = ~\new_[20789]_  | (~\new_[7744]_  & ~\new_[8468]_ );
  assign \new_[5663]_  = ~\new_[18942]_  | (~\new_[9610]_  & ~\new_[7745]_ );
  assign \new_[5664]_  = ~\new_[999]_  & (~\new_[7687]_  | ~\new_[9898]_ );
  assign \new_[5665]_  = ~\new_[19257]_  | (~\new_[7672]_  & ~\new_[7743]_ );
  assign \new_[5666]_  = ~\new_[19242]_  | (~\new_[7731]_  & ~\new_[8707]_ );
  assign \new_[5667]_  = ~\new_[7242]_  | ~\new_[19229]_ ;
  assign \new_[5668]_  = ~\new_[7250]_  | ~\new_[19702]_ ;
  assign \new_[5669]_  = ~\new_[18863]_  | (~\new_[7658]_  & ~\new_[15370]_ );
  assign \new_[5670]_  = ~\new_[7266]_  | ~\new_[21422]_ ;
  assign \new_[5671]_  = ~\new_[7268]_  | ~\new_[19157]_ ;
  assign \new_[5672]_  = ~\new_[17689]_  | (~\new_[7714]_  & ~\new_[13247]_ );
  assign \new_[5673]_  = ~\new_[19625]_  | (~\new_[7716]_  & ~\new_[15838]_ );
  assign \new_[5674]_  = ~\new_[8916]_  & (~\new_[8339]_  | ~\new_[18891]_ );
  assign \new_[5675]_  = ~\new_[7332]_  | ~\new_[19070]_ ;
  assign \new_[5676]_  = ~\new_[19561]_  & (~\new_[8438]_  | ~\new_[12129]_ );
  assign \new_[5677]_  = ~\new_[7304]_  & ~\new_[10888]_ ;
  assign \new_[5678]_  = ~\new_[7335]_  | ~\new_[19528]_ ;
  assign \new_[5679]_  = ~\new_[11225]_  & (~\new_[8450]_  | ~\new_[19215]_ );
  assign \new_[5680]_  = ~\new_[11265]_  & (~\new_[8491]_  | ~\new_[21557]_ );
  assign \new_[5681]_  = ~\new_[10761]_  & ~\new_[7185]_ ;
  assign \new_[5682]_  = ~\new_[10762]_  & ~\new_[7188]_ ;
  assign \new_[5683]_  = ~\new_[9433]_  & ~\new_[7190]_ ;
  assign \new_[5684]_  = ~\new_[9436]_  & ~\new_[7131]_ ;
  assign \new_[5685]_  = ~\new_[6167]_ ;
  assign \new_[5686]_  = ~\new_[7099]_  | ~\new_[21056]_ ;
  assign \new_[5687]_  = \new_[18630]_  ^ \new_[8244]_ ;
  assign \new_[5688]_  = ~\new_[19507]_  & (~\new_[8384]_  | ~\new_[12792]_ );
  assign \new_[5689]_  = ~\new_[7149]_  | ~\new_[21557]_ ;
  assign \new_[5690]_  = ~\new_[18077]_  | (~\new_[8436]_  & ~\new_[11692]_ );
  assign \new_[5691]_  = ~\new_[7166]_  | ~\new_[18077]_ ;
  assign \new_[5692]_  = ~\new_[7112]_  | ~\new_[19215]_ ;
  assign \new_[5693]_  = ~\new_[7309]_  | (~\new_[10412]_  & ~\new_[19528]_ );
  assign \new_[5694]_  = ~\new_[7312]_  | (~\new_[11397]_  & ~\new_[19070]_ );
  assign \new_[5695]_  = ~\new_[6177]_ ;
  assign \new_[5696]_  = ~\new_[7079]_  | ~\new_[8510]_ ;
  assign \new_[5697]_  = ~\new_[6183]_ ;
  assign \new_[5698]_  = ~\new_[10894]_  | ~\new_[8835]_  | ~\new_[7768]_ ;
  assign \new_[5699]_  = ~\new_[9824]_  & (~\new_[8356]_  | ~\new_[19553]_ );
  assign \new_[5700]_  = ~\new_[8357]_  & (~\new_[7518]_  | ~\new_[18361]_ );
  assign \new_[5701]_  = ~\new_[7094]_  | ~\new_[19508]_ ;
  assign \new_[5702]_  = ~\new_[19271]_  | (~\new_[8373]_  & ~\new_[8879]_ );
  assign \new_[5703]_  = ~\new_[7322]_  | ~\new_[18988]_ ;
  assign \new_[5704]_  = ~\new_[9970]_  | ~\new_[7967]_  | ~\new_[7771]_ ;
  assign \new_[5705]_  = ~\new_[9439]_  | ~\new_[10173]_  | ~\new_[8271]_ ;
  assign \new_[5706]_  = ~\new_[11197]_  | ~\new_[7075]_ ;
  assign \new_[5707]_  = ~\new_[7114]_  | ~\new_[19519]_ ;
  assign \new_[5708]_  = ~\new_[7325]_  | ~\new_[19507]_ ;
  assign \new_[5709]_  = ~\new_[7183]_  & ~\new_[9572]_ ;
  assign \new_[5710]_  = ~\new_[18650]_  | (~\new_[8408]_  & ~\new_[10551]_ );
  assign \new_[5711]_  = ~\new_[7284]_  | ~\new_[19404]_ ;
  assign \new_[5712]_  = ~\new_[19237]_  | (~\new_[8383]_  & ~\new_[7635]_ );
  assign \new_[5713]_  = ~\new_[20679]_  | (~\new_[8412]_  & ~\new_[9168]_ );
  assign \new_[5714]_  = ~\new_[8264]_  | ~\new_[12377]_  | ~\new_[9452]_ ;
  assign \new_[5715]_  = ~\new_[7125]_  & ~\new_[8432]_ ;
  assign \new_[5716]_  = \new_[7313]_  & \new_[12227]_ ;
  assign \new_[5717]_  = ~\new_[11948]_  | ~\new_[8917]_  | ~\new_[9305]_  | ~\new_[13322]_ ;
  assign \new_[5718]_  = ~\new_[7127]_  & ~\new_[16241]_ ;
  assign \new_[5719]_  = \new_[7265]_  | \new_[19528]_ ;
  assign \new_[5720]_  = ~\new_[6706]_  & (~\new_[9639]_  | ~\new_[18821]_ );
  assign \new_[5721]_  = ~\new_[7316]_  | ~\new_[10515]_ ;
  assign \new_[5722]_  = \new_[7314]_  & \new_[10962]_ ;
  assign \new_[5723]_  = ~\new_[10528]_  & (~\new_[7574]_  | ~\new_[18650]_ );
  assign \new_[5724]_  = ~\new_[19257]_  | (~\new_[8397]_  & ~\new_[8834]_ );
  assign \new_[5725]_  = ~\new_[19145]_  | (~\new_[8333]_  & ~\new_[13932]_ );
  assign \new_[5726]_  = ~\new_[19102]_  | (~\new_[8448]_  & ~\new_[10546]_ );
  assign \new_[5727]_  = ~\new_[19349]_  | (~\new_[8449]_  & ~\new_[7664]_ );
  assign \new_[5728]_  = ~\new_[7151]_  | ~\new_[20842]_ ;
  assign \new_[5729]_  = ~\new_[9914]_  | ~\new_[8779]_  | ~\new_[10235]_  | ~\new_[12251]_ ;
  assign \new_[5730]_  = ~\new_[7455]_  & (~\new_[8485]_  | ~\new_[18803]_ );
  assign \new_[5731]_  = \new_[7158]_  & \new_[8773]_ ;
  assign \new_[5732]_  = ~\new_[20701]_  | (~\new_[7471]_  & ~\new_[7684]_ );
  assign \new_[5733]_  = ~\new_[19523]_  & (~\new_[9628]_  | ~\new_[7932]_ );
  assign \new_[5734]_  = ~\new_[7167]_  | ~\new_[17796]_ ;
  assign \new_[5735]_  = ~\new_[19625]_  | (~\new_[7492]_  & ~\new_[11724]_ );
  assign \new_[5736]_  = ~\new_[18739]_  | (~\new_[9059]_  & ~\new_[7691]_ );
  assign \new_[5737]_  = ~\new_[14279]_  | ~\new_[6864]_  | ~\new_[8671]_ ;
  assign \new_[5738]_  = ~\new_[18769]_  | (~\new_[7504]_  & ~\new_[8673]_ );
  assign \new_[5739]_  = ~\new_[7220]_  | ~\new_[21638]_ ;
  assign \new_[5740]_  = ~\new_[19537]_  | (~\new_[7509]_  & ~\new_[8539]_ );
  assign \new_[5741]_  = ~\new_[17689]_  | (~\new_[8484]_  & ~\new_[10545]_ );
  assign \new_[5742]_  = ~\new_[14056]_  | ~\new_[7967]_  | ~\new_[7707]_ ;
  assign \new_[5743]_  = ~\new_[21422]_  & (~\new_[7511]_  | ~\new_[8542]_ );
  assign \new_[5744]_  = ~\new_[21267]_  & (~\new_[8545]_  | ~\new_[7516]_ );
  assign \new_[5745]_  = ~\new_[17796]_  | (~\new_[7521]_  & ~\new_[9140]_ );
  assign \new_[5746]_  = ~\new_[7326]_  | ~\new_[19384]_ ;
  assign \new_[5747]_  = ~\new_[21562]_  | (~\new_[7522]_  & ~\new_[10564]_ );
  assign \new_[5748]_  = ~\new_[7280]_  | ~\new_[21559]_ ;
  assign \new_[5749]_  = ~\new_[7327]_  | ~\new_[18399]_ ;
  assign \new_[5750]_  = ~\new_[7153]_  | ~\new_[13889]_ ;
  assign \new_[5751]_  = ~\new_[10079]_  | ~\new_[7072]_ ;
  assign \new_[5752]_  = ~\new_[6676]_  & (~\new_[8557]_  | ~\new_[21631]_ );
  assign \new_[5753]_  = ~\new_[6697]_  & (~\new_[9662]_  | ~\new_[19233]_ );
  assign \new_[5754]_  = ~\new_[11332]_  | ~\new_[7073]_ ;
  assign \new_[5755]_  = ~\new_[7318]_  | ~\new_[12768]_ ;
  assign \new_[5756]_  = ~\new_[9132]_  | ~\new_[7036]_ ;
  assign \new_[5757]_  = ~\new_[7319]_  | ~\new_[11612]_ ;
  assign \new_[5758]_  = ~\new_[7565]_  | ~\new_[13645]_  | ~\new_[7970]_ ;
  assign \new_[5759]_  = ~\new_[9987]_  | ~\new_[10377]_  | ~\new_[7772]_ ;
  assign \new_[5760]_  = ~\new_[7756]_  & ~\new_[12862]_  & ~\new_[12050]_ ;
  assign \new_[5761]_  = ~\new_[9973]_  | ~\new_[6864]_  | ~\new_[9784]_ ;
  assign \new_[5762]_  = ~\new_[11311]_  | ~\new_[7367]_  | ~\new_[8697]_ ;
  assign \new_[5763]_  = ~\new_[6729]_  & (~\new_[7589]_  | ~\new_[19013]_ );
  assign \new_[5764]_  = ~\new_[8603]_  | ~\new_[7228]_ ;
  assign \new_[5765]_  = ~\new_[9166]_  | ~\new_[7076]_ ;
  assign \new_[5766]_  = ~\new_[7208]_  & ~\new_[15279]_ ;
  assign \new_[5767]_  = ~\new_[8308]_  & (~\new_[7601]_  | ~\new_[19687]_ );
  assign \new_[5768]_  = ~\new_[7251]_  & (~\new_[13770]_  | ~\new_[19156]_ );
  assign \new_[5769]_  = ~\new_[7798]_  | ~\new_[7255]_ ;
  assign \new_[5770]_  = (~\new_[8410]_  | ~\new_[18833]_ ) & (~\new_[13736]_  | ~\new_[19203]_ );
  assign \new_[5771]_  = (~\new_[8376]_  | ~\new_[19547]_ ) & (~\new_[15892]_  | ~\new_[15586]_ );
  assign \new_[5772]_  = (~\new_[8403]_  | ~\new_[19206]_ ) & (~\new_[17488]_  | ~\new_[17017]_ );
  assign \new_[5773]_  = ~\new_[8628]_  | ~\new_[12994]_  | ~\new_[11181]_  | ~\new_[13667]_ ;
  assign \new_[5774]_  = ~\new_[11440]_  | ~\new_[7091]_  | ~\new_[7968]_ ;
  assign \new_[5775]_  = ~\new_[7625]_  & ~\new_[7097]_ ;
  assign \new_[5776]_  = ~\new_[7727]_  & ~\new_[7101]_ ;
  assign \new_[5777]_  = ~\new_[6756]_  & ~\new_[8119]_ ;
  assign \new_[5778]_  = ~\new_[10435]_  | ~\new_[9973]_  | ~\new_[11735]_  | ~\new_[7649]_ ;
  assign \new_[5779]_  = ~\new_[8649]_  | ~\new_[14116]_  | ~\new_[12368]_  | ~\new_[10235]_ ;
  assign \new_[5780]_  = ~\new_[8642]_  | ~\new_[14166]_  | ~\new_[13660]_  | ~\new_[12313]_ ;
  assign \new_[5781]_  = ~\new_[7673]_  & ~\new_[7147]_ ;
  assign \new_[5782]_  = ~\new_[7677]_  & ~\new_[7152]_ ;
  assign \new_[5783]_  = ~\new_[10663]_  | ~\new_[8141]_  | ~\new_[7922]_ ;
  assign \new_[5784]_  = ~\new_[18739]_  | (~\new_[7730]_  & ~\new_[14846]_ );
  assign \new_[5785]_  = ~\new_[13925]_  | ~\new_[7397]_  | ~\new_[8352]_ ;
  assign \new_[5786]_  = ~\new_[7301]_  & (~\new_[7662]_  | ~\new_[19045]_ );
  assign \new_[5787]_  = ~\new_[19005]_  | (~\new_[7620]_  & ~\new_[15284]_ );
  assign \new_[5788]_  = ~\new_[7290]_  & (~\new_[13474]_  | ~\new_[15005]_ );
  assign \new_[5789]_  = ~\new_[10274]_  | ~\new_[9574]_  | ~\new_[8275]_ ;
  assign \new_[5790]_  = ~\new_[6240]_ ;
  assign \new_[5791]_  = (~\new_[8406]_  | ~\new_[19450]_ ) & (~\new_[18157]_  | ~\new_[13344]_ );
  assign \new_[5792]_  = ~\new_[7288]_  & (~\new_[14855]_  | ~\new_[15064]_ );
  assign \new_[5793]_  = ~\new_[7289]_  & (~\new_[15829]_  | ~\new_[15332]_ );
  assign \new_[5794]_  = ~\new_[1878]_  & (~\new_[7629]_  | ~\new_[8426]_ );
  assign \new_[5795]_  = ~\new_[19102]_  | (~\new_[7993]_  & ~\new_[20087]_ );
  assign \new_[5796]_  = ~\new_[21629]_  | (~\new_[7663]_  & ~\new_[12591]_ );
  assign \new_[5797]_  = ~\new_[9879]_  | ~\new_[19838]_  | ~\new_[7769]_ ;
  assign \new_[5798]_  = ~\new_[19243]_  | (~\new_[7665]_  & ~\new_[15178]_ );
  assign \new_[5799]_  = ~\new_[16067]_  & (~\new_[8459]_  | ~\new_[18943]_ );
  assign \new_[5800]_  = (~\new_[8482]_  | ~\new_[21631]_ ) & (~\new_[16798]_  | ~\new_[18355]_ );
  assign \new_[5801]_  = ~\new_[13895]_  | (~\new_[7473]_  & ~\new_[21632]_ );
  assign \new_[5802]_  = ~\new_[21561]_  | (~\new_[7686]_  & ~\new_[11906]_ );
  assign \new_[5803]_  = ~\new_[6247]_ ;
  assign \new_[5804]_  = ~\new_[21629]_  | (~\new_[7700]_  & ~\new_[19837]_ );
  assign \new_[5805]_  = ~\new_[17689]_  | (~\new_[7704]_  & ~\new_[10635]_ );
  assign \new_[5806]_  = ~\new_[21562]_  | (~\new_[7710]_  & ~\new_[11776]_ );
  assign \new_[5807]_  = ~\new_[13195]_  | ~\new_[7041]_ ;
  assign \new_[5808]_  = ~\new_[16158]_  & (~\new_[7532]_  | ~\new_[18632]_ );
  assign \new_[5809]_  = ~\new_[19491]_  | (~\new_[7679]_  & ~\new_[13273]_ );
  assign \new_[5810]_  = ~\new_[7068]_  | ~\new_[20842]_ ;
  assign \new_[5811]_  = ~\new_[13999]_  & ~\new_[7275]_ ;
  assign \new_[5812]_  = ~\new_[8000]_  | ~\new_[9559]_  | ~\new_[8440]_ ;
  assign \new_[5813]_  = ~\new_[8004]_  | ~\new_[8547]_  | ~\new_[9651]_ ;
  assign \new_[5814]_  = ~\new_[9660]_  & ~\new_[7182]_ ;
  assign \new_[5815]_  = ~\new_[6707]_  & ~\new_[9374]_ ;
  assign \new_[5816]_  = ~\new_[12190]_  | ~\new_[7241]_  | ~\new_[12723]_ ;
  assign \new_[5817]_  = ~\new_[18522]_  | (~\new_[8321]_  & ~\new_[14017]_ );
  assign \new_[5818]_  = ~\new_[17323]_  | (~\new_[8363]_  & ~\new_[14365]_ );
  assign \new_[5819]_  = ~\new_[17470]_  | (~\new_[7643]_  & ~\new_[13181]_ );
  assign \new_[5820]_  = ~\new_[16811]_  | (~\new_[7645]_  & ~\new_[13284]_ );
  assign \new_[5821]_  = ~\new_[7160]_  | ~\new_[17411]_ ;
  assign \new_[5822]_  = ~\new_[21342]_  | (~\new_[7695]_  & ~\new_[12988]_ );
  assign \new_[5823]_  = ~\new_[17409]_  | (~\new_[7701]_  & ~\new_[15161]_ );
  assign \new_[5824]_  = ~\new_[7175]_  | ~\new_[16632]_ ;
  assign \new_[5825]_  = ~\new_[13317]_  | ~\new_[12274]_  | ~\new_[7948]_  | ~\new_[7994]_ ;
  assign \new_[5826]_  = ~\new_[16886]_  | (~\new_[7593]_  & ~\new_[13502]_ );
  assign \new_[5827]_  = ~\new_[8739]_  | ~\new_[14579]_  | ~\new_[12836]_  | ~\new_[12499]_ ;
  assign \new_[5828]_  = ~\new_[7391]_  & ~\new_[7032]_ ;
  assign \new_[5829]_  = (~\new_[7563]_  | ~\new_[18194]_ ) & (~\new_[15759]_  | ~\new_[16730]_ );
  assign \new_[5830]_  = (~\new_[7733]_  | ~\new_[19480]_ ) & (~\new_[11195]_  | ~\new_[18097]_ );
  assign \new_[5831]_  = ~\new_[9663]_  & (~\new_[7739]_  | ~\new_[19343]_ );
  assign \new_[5832]_  = ~\new_[8349]_  & ~\new_[7034]_ ;
  assign \new_[5833]_  = ~\new_[8718]_  | ~\new_[14059]_  | ~\new_[13805]_  | ~\new_[10549]_ ;
  assign \new_[5834]_  = ~\new_[8717]_  | ~\new_[14281]_  | ~\new_[10080]_  | ~\new_[15052]_ ;
  assign \new_[5835]_  = ~\new_[19939]_  | ~\new_[8506]_  | ~\new_[7751]_ ;
  assign \new_[5836]_  = ~\new_[8719]_  | ~\new_[14053]_  | ~\new_[10138]_  | ~\new_[15049]_ ;
  assign \new_[5837]_  = ~\new_[13208]_  | ~\new_[8526]_  | ~\new_[7752]_ ;
  assign \new_[5838]_  = ~\new_[9645]_  & ~\new_[7221]_ ;
  assign \new_[5839]_  = ~\new_[14030]_  | ~\new_[9646]_  | ~\new_[7753]_ ;
  assign \new_[5840]_  = ~\new_[20519]_  | ~\new_[6687]_  | ~\new_[8720]_ ;
  assign \new_[5841]_  = ~\new_[6917]_  & ~\new_[7307]_ ;
  assign \new_[5842]_  = ~\new_[6918]_  & ~\new_[8214]_ ;
  assign \new_[5843]_  = ~\new_[9929]_  | ~\new_[14376]_  | ~\new_[10423]_  | ~\new_[7953]_ ;
  assign \new_[5844]_  = ~\new_[11794]_  | ~\new_[7230]_ ;
  assign \new_[5845]_  = ~\new_[14307]_  | (~\new_[7749]_  & ~\new_[18077]_ );
  assign \new_[5846]_  = ~\new_[12561]_  | ~\new_[7238]_ ;
  assign \new_[5847]_  = (~\new_[7758]_  | ~\new_[18965]_ ) & (~\new_[16129]_  | ~\new_[19156]_ );
  assign \new_[5848]_  = (~\new_[7616]_  | ~\new_[19532]_ ) & (~\new_[18910]_  | ~\new_[15569]_ );
  assign \new_[5849]_  = (~\new_[7623]_  | ~\new_[19377]_ ) & (~\new_[17734]_  | ~\new_[12165]_ );
  assign \new_[5850]_  = ~\new_[10372]_  & (~\new_[8377]_  | ~\new_[19045]_ );
  assign \new_[5851]_  = (~\new_[7636]_  | ~\new_[18655]_ ) & (~\new_[18332]_  | ~\new_[15476]_ );
  assign \new_[5852]_  = ~\new_[10146]_  & (~\new_[8444]_  | ~\new_[17447]_ );
  assign \new_[5853]_  = \new_[11084]_  & \new_[7128]_ ;
  assign \new_[5854]_  = ~\new_[13968]_  | ~\new_[14966]_  | ~\new_[10879]_  | ~\new_[8371]_ ;
  assign \new_[5855]_  = ~\new_[11293]_  & ~\new_[7200]_ ;
  assign \new_[5856]_  = ~\new_[11244]_  & ~\new_[7150]_ ;
  assign \new_[5857]_  = ~\new_[7894]_  | ~\new_[7210]_ ;
  assign \new_[5858]_  = ~\new_[9841]_  & (~\new_[7661]_  | ~\new_[18739]_ );
  assign \new_[5859]_  = ~\new_[13599]_  & ~\new_[7216]_ ;
  assign \new_[5860]_  = ~\new_[9945]_  & (~\new_[7693]_  | ~\new_[21561]_ );
  assign \new_[5861]_  = ~\new_[11130]_  & (~\new_[7759]_  | ~\new_[19145]_ );
  assign \new_[5862]_  = ~\new_[11812]_  | ~\new_[10612]_  | ~\new_[8738]_  | ~\new_[15268]_ ;
  assign \new_[5863]_  = ~\new_[11909]_  | ~\new_[10666]_  | ~\new_[8761]_  | ~\new_[15258]_ ;
  assign \new_[5864]_  = ~\new_[18280]_  | (~\new_[8882]_  & ~\new_[7828]_ );
  assign \new_[5865]_  = ~\new_[21056]_  | (~\new_[8846]_  & ~\new_[7845]_ );
  assign \new_[5866]_  = ~\new_[18606]_  | (~\new_[8904]_  & ~\new_[7867]_ );
  assign \new_[5867]_  = ~\new_[18941]_  | (~\new_[7941]_  & ~\new_[13278]_ );
  assign \new_[5868]_  = \new_[6800]_  | \new_[20537]_ ;
  assign \new_[5869]_  = ~\new_[19262]_  & (~\new_[7943]_  | ~\new_[9066]_ );
  assign \new_[5870]_  = ~\new_[6290]_ ;
  assign \new_[5871]_  = \new_[6807]_  | \new_[21418]_ ;
  assign \new_[5872]_  = ~\new_[19271]_  & (~\new_[10674]_  | ~\new_[7779]_ );
  assign \new_[5873]_  = ~\new_[6677]_  | ~\new_[18288]_ ;
  assign \new_[5874]_  = \new_[7441]_  & \new_[21056]_ ;
  assign \new_[5875]_  = ~\new_[19021]_  & (~\new_[7782]_  | ~\new_[11708]_ );
  assign \new_[5876]_  = \new_[6754]_  | \new_[18941]_ ;
  assign \new_[5877]_  = ~\new_[6755]_  | ~\new_[18542]_ ;
  assign \new_[5878]_  = ~\new_[18280]_  & (~\new_[7787]_  | ~\new_[11491]_ );
  assign \new_[5879]_  = \new_[6773]_  & \new_[18606]_ ;
  assign \new_[5880]_  = \new_[6789]_  & \new_[19247]_ ;
  assign \new_[5881]_  = ~\new_[21638]_  & (~\new_[7790]_  | ~\new_[12818]_ );
  assign \new_[5882]_  = ~\new_[6804]_  | ~\new_[21638]_ ;
  assign \new_[5883]_  = ~\new_[19242]_  & (~\new_[12007]_  | ~\new_[7783]_ );
  assign \new_[5884]_  = ~\new_[19257]_  & (~\new_[12021]_  | ~\new_[7818]_ );
  assign \new_[5885]_  = ~\new_[18650]_  & (~\new_[7899]_  | ~\new_[12321]_ );
  assign \new_[5886]_  = ~\new_[19072]_  & (~\new_[7844]_  | ~\new_[12397]_ );
  assign \new_[5887]_  = ~\new_[18280]_  & (~\new_[7875]_  | ~\new_[12294]_ );
  assign \new_[5888]_  = ~\new_[7746]_  | ~\new_[6710]_ ;
  assign \new_[5889]_  = ~\new_[11921]_  & (~\new_[7901]_  | ~\new_[19208]_ );
  assign \new_[5890]_  = ~\new_[6837]_  | ~\new_[12139]_ ;
  assign \new_[5891]_  = ~\new_[6838]_  | ~\new_[8510]_ ;
  assign \new_[5892]_  = ~\new_[8716]_  | ~\new_[7408]_ ;
  assign \new_[5893]_  = ~\new_[15695]_  | ~\new_[15857]_  | ~\new_[7813]_ ;
  assign \new_[5894]_  = ~\new_[13430]_  | ~\new_[7817]_  | ~\new_[14601]_ ;
  assign \new_[5895]_  = ~\new_[16242]_  | ~\new_[15786]_  | ~\new_[7825]_ ;
  assign \new_[5896]_  = ~\new_[6340]_ ;
  assign \new_[5897]_  = ~\new_[6342]_ ;
  assign \new_[5898]_  = ~\new_[21166]_  | (~\new_[7876]_  & ~\new_[14887]_ );
  assign \new_[5899]_  = ~\new_[6774]_  | ~\new_[18786]_ ;
  assign \new_[5900]_  = ~\new_[18967]_  | (~\new_[7997]_  & ~\new_[10652]_ );
  assign \new_[5901]_  = ~\new_[19711]_  | (~\new_[7998]_  & ~\new_[10588]_ );
  assign \new_[5902]_  = ~\new_[7346]_  | ~\new_[16394]_ ;
  assign \new_[5903]_  = ~\new_[7354]_  | ~\new_[8839]_ ;
  assign \new_[5904]_  = ~\new_[17522]_  | (~\new_[7849]_  & ~\new_[12824]_ );
  assign \new_[5905]_  = ~\new_[18773]_  | (~\new_[7823]_  & ~\new_[15005]_ );
  assign \new_[5906]_  = ~\new_[7416]_  | ~\new_[19045]_ ;
  assign \new_[5907]_  = ~\new_[21115]_  | (~\new_[7999]_  & ~\new_[10698]_ );
  assign \new_[5908]_  = ~\new_[6365]_ ;
  assign \new_[5909]_  = ~\new_[19492]_  | (~\new_[7960]_  & ~\new_[11403]_ );
  assign \new_[5910]_  = ~\new_[6736]_  | ~\new_[20845]_ ;
  assign \new_[5911]_  = ~\new_[14037]_  | ~\new_[11366]_  | ~\new_[8764]_ ;
  assign \new_[5912]_  = ~\new_[19163]_  | (~\new_[7812]_  & ~\new_[7904]_ );
  assign \new_[5913]_  = ~\new_[18187]_  & (~\new_[7980]_  | ~\new_[15043]_ );
  assign \new_[5914]_  = ~\new_[18280]_  | (~\new_[8006]_  & ~\new_[20719]_ );
  assign \new_[5915]_  = ~\new_[19204]_  & (~\new_[10156]_  | ~\new_[7996]_ );
  assign \new_[5916]_  = \new_[6747]_  & \new_[21690]_ ;
  assign \new_[5917]_  = ~\new_[7407]_  | ~\new_[18895]_ ;
  assign \new_[5918]_  = ~\new_[18557]_  | (~\new_[7962]_  & ~\new_[12849]_ );
  assign \new_[5919]_  = \new_[6741]_  | \new_[18941]_ ;
  assign \new_[5920]_  = ~\new_[10508]_  | ~\new_[11543]_  | ~\new_[10041]_ ;
  assign \new_[5921]_  = ~\new_[6688]_  | ~\new_[16818]_ ;
  assign \new_[5922]_  = ~\new_[7435]_  | ~\new_[12738]_ ;
  assign \new_[5923]_  = ~\new_[6780]_  | ~\new_[10205]_ ;
  assign \new_[5924]_  = ~\new_[7448]_  | ~\new_[944]_ ;
  assign \new_[5925]_  = ~\new_[6401]_ ;
  assign \new_[5926]_  = \new_[6662]_  | \new_[19276]_ ;
  assign \new_[5927]_  = ~\new_[6742]_  | ~\new_[19491]_ ;
  assign \new_[5928]_  = ~\new_[6667]_  | ~\new_[17144]_ ;
  assign \new_[5929]_  = ~\new_[6670]_  | ~\new_[11721]_ ;
  assign \new_[5930]_  = ~\new_[6408]_ ;
  assign \new_[5931]_  = ~\new_[12747]_  | ~\new_[11607]_  | ~\new_[10200]_ ;
  assign \new_[5932]_  = ~\new_[7801]_  | ~\new_[8282]_  | ~\new_[9055]_ ;
  assign \new_[5933]_  = \new_[6743]_  | \new_[19450]_ ;
  assign \new_[5934]_  = ~\new_[6416]_ ;
  assign \new_[5935]_  = ~\new_[6417]_ ;
  assign \new_[5936]_  = ~\new_[17689]_  & (~\new_[7995]_  | ~\new_[10294]_ );
  assign \new_[5937]_  = \new_[6744]_  | \new_[21638]_ ;
  assign \new_[5938]_  = ~\new_[21562]_  & (~\new_[7989]_  | ~\new_[10134]_ );
  assign \new_[5939]_  = \new_[7345]_  | \new_[19215]_ ;
  assign \new_[5940]_  = ~\new_[7401]_  | ~\new_[12505]_ ;
  assign \new_[5941]_  = ~\new_[14951]_  | (~\new_[7836]_  & ~\new_[17245]_ );
  assign \new_[5942]_  = ~\new_[6779]_  | ~\new_[18752]_ ;
  assign \new_[5943]_  = ~\new_[6670]_  & ~\new_[18004]_ ;
  assign \new_[5944]_  = ~\new_[6822]_  & ~\new_[10031]_ ;
  assign \new_[5945]_  = ~\new_[7449]_  | ~\new_[19530]_ ;
  assign \new_[5946]_  = ~\new_[6823]_  | ~\new_[18154]_ ;
  assign \new_[5947]_  = ~\new_[6705]_  | ~\new_[10358]_ ;
  assign \new_[5948]_  = ~\new_[17874]_  | (~\new_[9358]_  & ~\new_[8005]_ );
  assign \new_[5949]_  = ~\new_[15219]_  | ~\new_[12716]_  | ~\new_[7826]_ ;
  assign \new_[5950]_  = ~\new_[6829]_  | ~\new_[18380]_ ;
  assign \new_[5951]_  = ~\new_[6447]_ ;
  assign \new_[5952]_  = ~\new_[13059]_  | ~\new_[12524]_  | ~\new_[6877]_  | ~\new_[9848]_ ;
  assign \new_[5953]_  = ~\new_[6772]_  & ~\new_[12320]_ ;
  assign \new_[5954]_  = ~\new_[14362]_  & ~\new_[7351]_ ;
  assign \new_[5955]_  = ~\new_[7456]_  & ~\new_[9012]_ ;
  assign \new_[5956]_  = ~\new_[6459]_ ;
  assign \new_[5957]_  = ~\new_[6461]_ ;
  assign \new_[5958]_  = ~\new_[9361]_  | ~\new_[12658]_  | ~\new_[10297]_  | ~\new_[12274]_ ;
  assign \new_[5959]_  = ~\new_[14162]_  & ~\new_[7350]_ ;
  assign \new_[5960]_  = ~\new_[6465]_ ;
  assign \new_[5961]_  = ~\new_[6467]_ ;
  assign \new_[5962]_  = ~\new_[19088]_  | (~\new_[7822]_  & ~\new_[10934]_ );
  assign \new_[5963]_  = ~\new_[7380]_  | ~\new_[19859]_ ;
  assign \new_[5964]_  = ~\new_[7383]_  | ~\new_[19088]_ ;
  assign \new_[5965]_  = ~\new_[9941]_  | ~\new_[9292]_  | ~\new_[7986]_ ;
  assign \new_[5966]_  = ~\new_[8811]_  | ~\new_[14786]_  | ~\new_[7987]_ ;
  assign \new_[5967]_  = ~\new_[8354]_  & (~\new_[8009]_  | ~\new_[18739]_ );
  assign \new_[5968]_  = ~\new_[7400]_  | ~\new_[17851]_ ;
  assign \new_[5969]_  = ~\new_[10887]_  | ~\new_[13104]_  | ~\new_[7988]_ ;
  assign \new_[5970]_  = ~\new_[14035]_  | (~\new_[7883]_  & ~\new_[19279]_ );
  assign \new_[5971]_  = \new_[7406]_  & \new_[10039]_ ;
  assign \new_[5972]_  = ~\new_[7419]_  | ~\new_[7900]_ ;
  assign \new_[5973]_  = ~\new_[14115]_  | (~\new_[7890]_  & ~\new_[19407]_ );
  assign \new_[5974]_  = ~\new_[7386]_  | ~\new_[20483]_ ;
  assign \new_[5975]_  = ~\new_[7427]_  | ~\new_[12669]_ ;
  assign \new_[5976]_  = ~\new_[7387]_  | ~\new_[12641]_ ;
  assign \new_[5977]_  = ~\new_[9560]_  | ~\new_[6879]_ ;
  assign \new_[5978]_  = ~\new_[7426]_  | ~\new_[14901]_ ;
  assign \new_[5979]_  = ~\new_[12292]_  | (~\new_[7833]_  & ~\new_[19625]_ );
  assign \new_[5980]_  = ~\new_[9860]_  | ~\new_[10661]_  | ~\new_[7991]_ ;
  assign \new_[5981]_  = ~\new_[7436]_  | ~\new_[21562]_ ;
  assign \new_[5982]_  = \new_[7445]_  & \new_[10203]_ ;
  assign \new_[5983]_  = \new_[7414]_  | \new_[12577]_ ;
  assign \new_[5984]_  = ~\new_[7457]_  | ~\new_[19208]_ ;
  assign \new_[5985]_  = ~\new_[6675]_  & (~\new_[8011]_  | ~\new_[21561]_ );
  assign \new_[5986]_  = ~\new_[13776]_  | ~\new_[11769]_  | ~\new_[6879]_  | ~\new_[15398]_ ;
  assign \new_[5987]_  = ~\new_[18923]_  & (~\new_[7854]_  | ~\new_[17376]_ );
  assign \new_[5988]_  = ~\new_[20802]_  | (~\new_[7921]_  & ~\new_[21557]_ );
  assign \new_[5989]_  = ~\new_[6681]_  & ~\new_[8270]_ ;
  assign \new_[5990]_  = ~\new_[9355]_  | ~\new_[7373]_ ;
  assign \new_[5991]_  = ~\new_[9341]_  | ~\new_[6811]_  | ~\new_[8794]_ ;
  assign \new_[5992]_  = ~\new_[11985]_  | ~\new_[6813]_  | ~\new_[7788]_ ;
  assign \new_[5993]_  = ~\new_[20781]_  | (~\new_[9273]_  & ~\new_[21561]_ );
  assign \new_[5994]_  = ~\new_[6700]_  & (~\new_[12470]_  | ~\new_[19384]_ );
  assign \new_[5995]_  = ~\new_[6703]_  | ~\new_[19450]_ ;
  assign \new_[5996]_  = ~\new_[7433]_  | ~\new_[17749]_ ;
  assign \new_[5997]_  = ~\new_[10587]_  | ~\new_[7374]_ ;
  assign \new_[5998]_  = ~\new_[6718]_  | ~\new_[14389]_ ;
  assign \new_[5999]_  = ~\new_[6726]_  | ~\new_[12161]_ ;
  assign \new_[6000]_  = ~\new_[17385]_  & (~\new_[7820]_  | ~\new_[14079]_ );
  assign \new_[6001]_  = \new_[9431]_  | \new_[7366]_ ;
  assign \new_[6002]_  = ~\new_[13285]_  | ~\new_[11566]_  | ~\new_[6858]_  | ~\new_[14279]_ ;
  assign \new_[6003]_  = ~\new_[7444]_  | ~\new_[17106]_ ;
  assign \new_[6004]_  = ~\new_[7398]_  & (~\new_[10477]_  | ~\new_[18906]_ );
  assign \new_[6005]_  = ~\new_[6548]_ ;
  assign \new_[6006]_  = ~\new_[7423]_  & (~\new_[11456]_  | ~\new_[17578]_ );
  assign \new_[6007]_  = ~\new_[14381]_  | ~\new_[10004]_  | ~\new_[12609]_ ;
  assign \new_[6008]_  = ~\new_[12658]_  | ~\new_[8960]_  | ~\new_[10232]_ ;
  assign \new_[6009]_  = ~\new_[10534]_  & ~\new_[7382]_ ;
  assign \new_[6010]_  = ~\new_[10180]_  & ~\new_[7361]_ ;
  assign \new_[6011]_  = \new_[7420]_  & \new_[8386]_ ;
  assign \new_[6012]_  = ~\new_[7229]_  | ~\new_[17663]_ ;
  assign \new_[6013]_  = \new_[6669]_  & \new_[7476]_ ;
  assign \new_[6014]_  = \new_[6678]_  & \new_[8528]_ ;
  assign \new_[6015]_  = ~\new_[20987]_  | ~\new_[13713]_  | ~\new_[7833]_ ;
  assign \new_[6016]_  = ~\new_[9949]_  | ~\new_[6683]_  | ~\new_[14806]_ ;
  assign \new_[6017]_  = ~\new_[8643]_  | ~\new_[7349]_ ;
  assign \new_[6018]_  = ~\new_[6826]_  | ~\new_[8258]_ ;
  assign \new_[6019]_  = ~\new_[6820]_  | ~\new_[8259]_ ;
  assign \new_[6020]_  = ~\new_[7375]_  | ~\new_[7429]_ ;
  assign \new_[6021]_  = \new_[8247]_  & \new_[7418]_ ;
  assign \new_[6022]_  = ~\new_[6711]_  | ~\new_[6712]_ ;
  assign \new_[6023]_  = \new_[14905]_  ^ \new_[19520]_ ;
  assign \new_[6024]_  = ~\new_[6609]_ ;
  assign \new_[6025]_  = ~\new_[6611]_ ;
  assign \new_[6026]_  = ~\new_[6853]_  & ~\new_[18280]_ ;
  assign \new_[6027]_  = ~\new_[6938]_  | ~\new_[21418]_ ;
  assign \new_[6028]_  = ~\new_[11735]_  | ~\new_[6853]_ ;
  assign \new_[6029]_  = ~\new_[6624]_ ;
  assign \new_[6030]_  = ~\new_[6629]_ ;
  assign \new_[6031]_  = ~\new_[6931]_  | ~\new_[19088]_ ;
  assign \new_[6032]_  = \new_[6932]_  | \new_[18280]_ ;
  assign \new_[6033]_  = ~\new_[14382]_  | ~\new_[6853]_ ;
  assign \new_[6034]_  = ~\new_[20620]_  | ~\new_[19711]_ ;
  assign \new_[6035]_  = ~\new_[7911]_  | ~\new_[12183]_ ;
  assign \new_[6036]_  = ~\new_[10334]_  & ~\new_[11078]_ ;
  assign \new_[6037]_  = \new_[7927]_  | \new_[18361]_ ;
  assign \new_[6038]_  = ~\new_[9883]_  | ~\new_[11811]_ ;
  assign \new_[6039]_  = ~\new_[6670]_ ;
  assign \new_[6040]_  = ~\new_[17866]_  & (~\new_[9349]_  | ~\new_[13340]_ );
  assign \new_[6041]_  = \new_[7926]_  & \new_[7786]_ ;
  assign \new_[6042]_  = ~\new_[11021]_  & ~\new_[7780]_ ;
  assign \new_[6043]_  = ~\new_[6682]_ ;
  assign \new_[6044]_  = \new_[7896]_  | \new_[17837]_ ;
  assign \new_[6045]_  = ~\new_[14272]_  & ~\new_[9802]_ ;
  assign \new_[6046]_  = \new_[11016]_  & \new_[7977]_ ;
  assign \new_[6047]_  = ~\new_[9928]_  & ~\new_[9874]_ ;
  assign \new_[6048]_  = ~\new_[7809]_  & ~\new_[11019]_ ;
  assign \new_[6049]_  = ~\new_[8015]_  | ~\new_[18409]_ ;
  assign \new_[6050]_  = ~\new_[11885]_  | ~\new_[8764]_ ;
  assign \new_[6051]_  = ~\new_[14149]_  | ~\new_[8764]_ ;
  assign \new_[6052]_  = ~\new_[7915]_  | ~\new_[10921]_ ;
  assign \new_[6053]_  = ~\new_[6695]_ ;
  assign \new_[6054]_  = ~\new_[7810]_  | ~\new_[10589]_ ;
  assign \new_[6055]_  = ~\new_[8016]_  | ~\new_[18293]_ ;
  assign \new_[6056]_  = ~\new_[11806]_  | ~\new_[7783]_ ;
  assign \new_[6057]_  = ~\new_[6705]_ ;
  assign \new_[6058]_  = ~\new_[7785]_  | ~\new_[14005]_ ;
  assign \new_[6059]_  = ~\new_[7944]_  | ~\new_[17469]_ ;
  assign \new_[6060]_  = ~\new_[7977]_  | ~\new_[12651]_ ;
  assign \new_[6061]_  = ~\new_[9359]_  | ~\new_[7818]_ ;
  assign \new_[6062]_  = ~\new_[7972]_  | ~\new_[12917]_ ;
  assign \new_[6063]_  = ~\new_[7807]_  | ~\new_[13252]_ ;
  assign \new_[6064]_  = ~\new_[19711]_  & (~\new_[9287]_  | ~\new_[15408]_ );
  assign \new_[6065]_  = ~\new_[6734]_ ;
  assign \new_[6066]_  = ~\new_[12513]_  | ~\new_[12295]_  | ~\new_[10531]_ ;
  assign \new_[6067]_  = ~\new_[8003]_  | ~\new_[10977]_ ;
  assign \new_[6068]_  = ~\new_[11712]_  | ~\new_[12406]_  | ~\new_[10532]_ ;
  assign \new_[6069]_  = ~\new_[12701]_  | ~\new_[10232]_  | ~\new_[11648]_ ;
  assign \new_[6070]_  = ~\new_[6749]_ ;
  assign \new_[6071]_  = ~\new_[8939]_  & ~\new_[10154]_ ;
  assign \new_[6072]_  = ~\new_[12585]_  | ~\new_[9883]_ ;
  assign \new_[6073]_  = ~\new_[10405]_  & (~\new_[14733]_  | ~\new_[19407]_ );
  assign \new_[6074]_  = ~\new_[13966]_  & (~\new_[11815]_  | ~\new_[19520]_ );
  assign \new_[6075]_  = ~\new_[7881]_  & ~\new_[10460]_ ;
  assign \new_[6076]_  = \new_[7887]_  & \new_[10071]_ ;
  assign \new_[6077]_  = \new_[7834]_  & \new_[13786]_ ;
  assign \new_[6078]_  = ~\new_[13725]_  | (~\new_[14259]_  & ~\new_[17469]_ );
  assign \new_[6079]_  = ~\new_[11818]_  & ~\new_[7793]_ ;
  assign \new_[6080]_  = ~\new_[6778]_ ;
  assign \new_[6081]_  = ~\new_[10711]_  | ~\new_[16124]_  | ~\new_[10033]_  | ~\new_[11334]_ ;
  assign \new_[6082]_  = ~\new_[7914]_  | ~\new_[13654]_ ;
  assign \new_[6083]_  = ~\new_[7964]_  | ~\new_[13648]_ ;
  assign \new_[6084]_  = ~\new_[21408]_  | (~\new_[14027]_  & ~\new_[18974]_ );
  assign \new_[6085]_  = \new_[9073]_  & \new_[7935]_ ;
  assign \new_[6086]_  = ~\new_[19236]_  & (~\new_[9365]_  | ~\new_[15897]_ );
  assign \new_[6087]_  = ~\new_[7947]_  | ~\new_[17522]_ ;
  assign \new_[6088]_  = ~\new_[7811]_  | ~\new_[12593]_ ;
  assign \new_[6089]_  = ~\new_[11669]_  | (~\new_[21678]_  & ~\new_[21495]_ );
  assign \new_[6090]_  = ~\new_[11851]_  & ~\new_[7781]_ ;
  assign \new_[6091]_  = ~\new_[17689]_  & (~\new_[9275]_  | ~\new_[13649]_ );
  assign \new_[6092]_  = ~\new_[9123]_  & ~\new_[10581]_ ;
  assign \new_[6093]_  = ~\new_[6827]_ ;
  assign \new_[6094]_  = ~\new_[11455]_  | ~\new_[7820]_ ;
  assign \new_[6095]_  = ~\new_[7775]_  | ~\new_[11763]_ ;
  assign \new_[6096]_  = ~\new_[7789]_  | ~\new_[11860]_ ;
  assign \new_[6097]_  = ~\new_[7800]_  | ~\new_[11855]_ ;
  assign \new_[6098]_  = ~\new_[11971]_  | ~\new_[7808]_ ;
  assign \new_[6099]_  = ~\new_[7939]_  & ~\new_[11219]_ ;
  assign \new_[6100]_  = ~\new_[12057]_  | (~\new_[18540]_  & ~\new_[9279]_ );
  assign \new_[6101]_  = ~\new_[10363]_  | ~\new_[7838]_ ;
  assign \new_[6102]_  = ~\new_[10204]_  | ~\new_[7871]_ ;
  assign \new_[6103]_  = ~\new_[7951]_  & (~\new_[12663]_  | ~\new_[18120]_ );
  assign \new_[6104]_  = ~\new_[7934]_  & (~\new_[11541]_  | ~\new_[17468]_ );
  assign \new_[6105]_  = ~\new_[7862]_  & (~\new_[12519]_  | ~\new_[17840]_ );
  assign \new_[6106]_  = ~\new_[7982]_  & (~\new_[11529]_  | ~\new_[17917]_ );
  assign \new_[6107]_  = ~\new_[7916]_  | ~\new_[10385]_ ;
  assign \new_[6108]_  = ~\new_[10520]_  | ~\new_[14664]_  | ~\new_[13359]_  | ~\new_[12768]_ ;
  assign \new_[6109]_  = ~\new_[7892]_  | ~\new_[12971]_ ;
  assign \new_[6110]_  = ~\new_[7909]_  | ~\new_[13193]_ ;
  assign \new_[6111]_  = ~\new_[10567]_  | ~\new_[7791]_ ;
  assign \new_[6112]_  = ~\new_[6851]_ ;
  assign \new_[6113]_  = ~\new_[20719]_  | ~\new_[19625]_ ;
  assign \new_[6114]_  = ~\new_[6852]_ ;
  assign \new_[6115]_  = ~\new_[9836]_  | ~\new_[16169]_  | ~\new_[8039]_  | ~\new_[15668]_ ;
  assign \new_[6116]_  = ~\new_[17689]_  | ~\new_[10514]_ ;
  assign \new_[6117]_  = ~\new_[8050]_  | ~\new_[19567]_ ;
  assign \new_[6118]_  = ~\new_[10403]_  & ~\new_[21562]_ ;
  assign \new_[6119]_  = ~\new_[18280]_  | ~\new_[10561]_ ;
  assign \new_[6120]_  = ~\new_[6859]_ ;
  assign \new_[6121]_  = ~\new_[10509]_  & ~\new_[18228]_ ;
  assign \new_[6122]_  = ~\new_[20660]_  & ~\new_[19204]_ ;
  assign \new_[6123]_  = \new_[8031]_  | \new_[18077]_ ;
  assign \new_[6124]_  = ~\new_[8070]_  & ~\new_[14951]_ ;
  assign \new_[6125]_  = ~\new_[8035]_  | ~\new_[19299]_ ;
  assign \new_[6126]_  = ~\new_[19404]_  | (~\new_[9337]_  & ~\new_[12733]_ );
  assign \new_[6127]_  = ~\new_[8044]_  | ~\new_[19502]_ ;
  assign \new_[6128]_  = ~\new_[18569]_  & ~\new_[8041]_ ;
  assign \new_[6129]_  = ~\new_[8049]_  | ~\new_[18667]_ ;
  assign \new_[6130]_  = \new_[10185]_  | \new_[21056]_ ;
  assign \new_[6131]_  = ~\new_[12242]_  | ~\new_[10834]_  | ~\new_[11242]_  | ~\new_[10993]_ ;
  assign \new_[6132]_  = ~\new_[8026]_  | ~\new_[16435]_ ;
  assign \new_[6133]_  = ~\new_[18606]_  & ~\new_[20809]_ ;
  assign \new_[6134]_  = ~\new_[9324]_  | ~\new_[9092]_  | ~\new_[8680]_ ;
  assign \new_[6135]_  = ~\new_[11363]_  | ~\new_[10838]_  | ~\new_[9367]_ ;
  assign \new_[6136]_  = \new_[9644]_  | \new_[11442]_  | \new_[20150]_  | \new_[13220]_ ;
  assign \new_[6137]_  = ~\new_[8034]_  | ~\new_[946]_ ;
  assign \new_[6138]_  = ~\new_[10626]_  | ~\new_[19102]_ ;
  assign \new_[6139]_  = ~\new_[10038]_  & (~\new_[9379]_  | ~\new_[19578]_ );
  assign \new_[6140]_  = ~\new_[10332]_  & (~\new_[9381]_  | ~\new_[19561]_ );
  assign \new_[6141]_  = ~\new_[10743]_  | ~\new_[9822]_  | ~\new_[16204]_  | ~\new_[9821]_ ;
  assign \new_[6142]_  = ~\new_[10747]_  | ~\new_[13208]_  | ~\new_[10054]_  | ~\new_[11505]_ ;
  assign \new_[6143]_  = ~\new_[8028]_  & (~\new_[17488]_  | ~\new_[16461]_ );
  assign \new_[6144]_  = ~\new_[11866]_  | ~\new_[15133]_  | ~\new_[10751]_  | ~\new_[11527]_ ;
  assign \new_[6145]_  = ~\new_[10749]_  | ~\new_[13921]_  | ~\new_[13217]_  | ~\new_[11646]_ ;
  assign \new_[6146]_  = ~\new_[10739]_  | ~\new_[13171]_  | ~\new_[12015]_  | ~\new_[13891]_ ;
  assign \new_[6147]_  = ~\new_[15479]_  & ~\new_[8043]_ ;
  assign \new_[6148]_  = ~\new_[19284]_  & (~\new_[8935]_  | ~\new_[8733]_ );
  assign \new_[6149]_  = ~\new_[14256]_  & ~\new_[8045]_ ;
  assign \new_[6150]_  = ~\new_[959]_  & (~\new_[10279]_  | ~\new_[8731]_ );
  assign \new_[6151]_  = ~\new_[8231]_  & (~\new_[15768]_  | ~\new_[15798]_ );
  assign \new_[6152]_  = ~\new_[19502]_  & (~\new_[10815]_  | ~\new_[8730]_ );
  assign \new_[6153]_  = ~\new_[19508]_  & (~\new_[8604]_  | ~\new_[16166]_ );
  assign \new_[6154]_  = ~\new_[11497]_  | ~\new_[8026]_ ;
  assign \new_[6155]_  = ~\new_[19587]_  | (~\new_[8575]_  & ~\new_[12674]_ );
  assign \new_[6156]_  = ~\new_[18481]_  | (~\new_[9507]_  & ~\new_[11538]_ );
  assign \new_[6157]_  = ~\new_[19233]_  | (~\new_[9519]_  & ~\new_[11699]_ );
  assign \new_[6158]_  = ~\new_[19357]_  | (~\new_[9594]_  & ~\new_[11611]_ );
  assign \new_[6159]_  = ~\new_[19550]_  | (~\new_[9773]_  & ~\new_[9525]_ );
  assign \new_[6160]_  = ~\new_[1025]_  & (~\new_[9526]_  | ~\new_[14386]_ );
  assign \new_[6161]_  = ~\new_[19300]_  & (~\new_[9615]_  | ~\new_[16210]_ );
  assign \new_[6162]_  = ~\new_[19021]_  | (~\new_[8659]_  & ~\new_[14321]_ );
  assign \new_[6163]_  = ~\new_[8070]_  | (~\new_[18442]_  & ~\new_[13397]_ );
  assign \new_[6164]_  = ~\new_[8587]_  | ~\new_[9845]_  | ~\new_[16212]_ ;
  assign \new_[6165]_  = \new_[18866]_  ^ \new_[9412]_ ;
  assign \new_[6166]_  = ~\new_[8100]_  | ~\new_[18798]_ ;
  assign \new_[6167]_  = ~\new_[19177]_  & (~\new_[9487]_  | ~\new_[12544]_ );
  assign \new_[6168]_  = ~\new_[8111]_  | ~\new_[19064]_ ;
  assign \new_[6169]_  = ~\new_[19381]_  | (~\new_[9571]_  & ~\new_[12598]_ );
  assign \new_[6170]_  = \new_[18897]_  ^ \new_[9400]_ ;
  assign \new_[6171]_  = ~\new_[18280]_  | (~\new_[8570]_  & ~\new_[12620]_ );
  assign \new_[6172]_  = \new_[18767]_  ^ \new_[9396]_ ;
  assign \new_[6173]_  = ~\new_[8136]_  | ~\new_[18795]_ ;
  assign \new_[6174]_  = ~\new_[17689]_  | (~\new_[9611]_  & ~\new_[12549]_ );
  assign \new_[6175]_  = ~\new_[21562]_  | (~\new_[8524]_  & ~\new_[12685]_ );
  assign \new_[6176]_  = ~\new_[6948]_ ;
  assign \new_[6177]_  = ~\new_[11396]_  & (~\new_[8686]_  | ~\new_[1878]_ );
  assign \new_[6178]_  = ~\new_[8217]_  | (~\new_[9187]_  & ~\new_[18668]_ );
  assign \new_[6179]_  = ~\new_[6949]_ ;
  assign \new_[6180]_  = ~\new_[8219]_  | (~\new_[9206]_  & ~\new_[19502]_ );
  assign \new_[6181]_  = ~\new_[13998]_  | ~\new_[10082]_  | ~\new_[14070]_  | ~\new_[14407]_ ;
  assign \new_[6182]_  = ~\new_[9605]_  | ~\new_[9991]_  | ~\new_[12199]_ ;
  assign \new_[6183]_  = ~\new_[9803]_  | ~\new_[7831]_  | ~\new_[9785]_ ;
  assign \new_[6184]_  = ~\new_[15901]_  & (~\new_[8623]_  | ~\new_[12469]_ );
  assign \new_[6185]_  = ~\new_[9961]_  & (~\new_[9493]_  | ~\new_[18750]_ );
  assign \new_[6186]_  = ~\new_[21620]_  & (~\new_[9599]_  | ~\new_[17983]_ );
  assign \new_[6187]_  = ~\new_[8221]_  | ~\new_[15225]_ ;
  assign \new_[6188]_  = \new_[8216]_  & \new_[10917]_ ;
  assign \new_[6189]_  = ~\new_[8187]_  | ~\new_[19003]_ ;
  assign \new_[6190]_  = ~\new_[19578]_  | (~\new_[9521]_  & ~\new_[10089]_ );
  assign \new_[6191]_  = ~\new_[21129]_  | ~\new_[19361]_ ;
  assign \new_[6192]_  = ~\new_[11204]_  & (~\new_[9541]_  | ~\new_[19228]_ );
  assign \new_[6193]_  = ~\new_[19453]_  | (~\new_[9470]_  & ~\new_[9545]_ );
  assign \new_[6194]_  = ~\new_[19480]_  | (~\new_[9549]_  & ~\new_[9531]_ );
  assign \new_[6195]_  = ~\new_[1928]_  | (~\new_[10810]_  & ~\new_[9562]_ );
  assign \new_[6196]_  = ~\new_[9563]_  | ~\new_[10000]_  | ~\new_[10968]_ ;
  assign \new_[6197]_  = ~\new_[17244]_  & (~\new_[8693]_  | ~\new_[21615]_ );
  assign \new_[6198]_  = ~\new_[8721]_  & ~\new_[13224]_  & ~\new_[12054]_ ;
  assign \new_[6199]_  = ~\new_[12145]_  & (~\new_[9466]_  | ~\new_[18909]_ );
  assign \new_[6200]_  = ~\new_[21629]_  & (~\new_[9584]_  | ~\new_[9585]_ );
  assign \new_[6201]_  = ~\new_[12771]_  | ~\new_[12918]_  | ~\new_[9900]_  | ~\new_[11375]_ ;
  assign \new_[6202]_  = ~\new_[9857]_  | ~\new_[13106]_  | ~\new_[13858]_  | ~\new_[10041]_ ;
  assign \new_[6203]_  = ~\new_[1025]_  | (~\new_[9604]_  & ~\new_[10842]_ );
  assign \new_[6204]_  = ~\new_[20842]_  | (~\new_[8581]_  & ~\new_[9506]_ );
  assign \new_[6205]_  = ~\new_[19711]_  | (~\new_[8496]_  & ~\new_[21623]_ );
  assign \new_[6206]_  = ~\new_[17668]_  | (~\new_[8497]_  & ~\new_[8664]_ );
  assign \new_[6207]_  = ~\new_[19448]_  | (~\new_[8518]_  & ~\new_[9051]_ );
  assign \new_[6208]_  = ~\new_[999]_  | (~\new_[8522]_  & ~\new_[8523]_ );
  assign \new_[6209]_  = ~\new_[15299]_  | ~\new_[13648]_  | ~\new_[8675]_ ;
  assign \new_[6210]_  = ~\new_[19361]_  | (~\new_[8535]_  & ~\new_[9069]_ );
  assign \new_[6211]_  = ~\new_[8200]_  | ~\new_[19243]_ ;
  assign \new_[6212]_  = ~\new_[14349]_  | ~\new_[7907]_  | ~\new_[9727]_ ;
  assign \new_[6213]_  = \new_[10309]_  | \new_[15184]_  | \new_[14254]_  | \new_[12058]_ ;
  assign \new_[6214]_  = ~\new_[21633]_  | (~\new_[8550]_  & ~\new_[21548]_ );
  assign \new_[6215]_  = ~\new_[7531]_  & (~\new_[9661]_  | ~\new_[20099]_ );
  assign \new_[6216]_  = ~\new_[20221]_  | ~\new_[10328]_  | ~\new_[10640]_  | ~\new_[13327]_ ;
  assign \new_[6217]_  = ~\new_[8567]_  | ~\new_[9851]_  | ~\new_[9971]_ ;
  assign \new_[6218]_  = ~\new_[8724]_  & ~\new_[13062]_  & ~\new_[12048]_ ;
  assign \new_[6219]_  = ~\new_[13687]_  | ~\new_[7832]_  | ~\new_[9263]_ ;
  assign \new_[6220]_  = ~\new_[8544]_  | ~\new_[16259]_  | ~\new_[9159]_ ;
  assign \new_[6221]_  = ~\new_[8586]_  | ~\new_[9952]_  | ~\new_[8816]_ ;
  assign \new_[6222]_  = ~\new_[9683]_  | ~\new_[15112]_  | ~\new_[8601]_ ;
  assign \new_[6223]_  = ~\\u0_r0_out_reg[28] ;
  assign \new_[6224]_  = (~\new_[8571]_  | ~\new_[19625]_ ) & (~\new_[12715]_  | ~\new_[18973]_ );
  assign \new_[6225]_  = ~\new_[7575]_  | ~\new_[8226]_ ;
  assign \new_[6226]_  = ~\new_[8622]_  | ~\new_[8101]_ ;
  assign \new_[6227]_  = ~\new_[8104]_  | (~\new_[10036]_  & ~\new_[19079]_ );
  assign \new_[6228]_  = ~\new_[8620]_  | ~\new_[8120]_ ;
  assign \new_[6229]_  = ~\new_[8684]_  | ~\new_[8125]_ ;
  assign \new_[6230]_  = ~\new_[8162]_  | (~\new_[10127]_  & ~\new_[18361]_ );
  assign \new_[6231]_  = ~\new_[8652]_  | ~\new_[8134]_ ;
  assign \new_[6232]_  = ~\new_[8137]_  | ~\new_[8658]_ ;
  assign \new_[6233]_  = ~\new_[8140]_  | (~\new_[10233]_  & ~\new_[19436]_ );
  assign \new_[6234]_  = ~\new_[9696]_  | ~\new_[14257]_  | ~\new_[11302]_  | ~\new_[13655]_ ;
  assign \new_[6235]_  = ~\new_[13727]_  | ~\new_[9485]_  | ~\new_[9484]_ ;
  assign \new_[6236]_  = (~\new_[9491]_  | ~\new_[18076]_ ) & (~\new_[17039]_  | ~\new_[18773]_ );
  assign \new_[6237]_  = ~\new_[7571]_  & (~\new_[9765]_  | ~\new_[18965]_ );
  assign \new_[6238]_  = ~\new_[8427]_  & (~\new_[9724]_  | ~\new_[18998]_ );
  assign \new_[6239]_  = ~\new_[18941]_  | (~\new_[9721]_  & ~\new_[21197]_ );
  assign \new_[6240]_  = ~\new_[19064]_  | (~\new_[8688]_  & ~\new_[21468]_ );
  assign \new_[6241]_  = ~\new_[11582]_  | ~\new_[10862]_  | ~\new_[9417]_ ;
  assign \new_[6242]_  = ~\new_[13669]_  | ~\new_[9568]_  | ~\new_[9567]_ ;
  assign \new_[6243]_  = ~\new_[15092]_  | (~\new_[9522]_  & ~\new_[18443]_ );
  assign \new_[6244]_  = ~\new_[18798]_  | (~\new_[8663]_  & ~\new_[19950]_ );
  assign \new_[6245]_  = \new_[9330]_  ^ \new_[18756]_ ;
  assign \new_[6246]_  = ~\new_[13590]_  | ~\new_[8501]_  | ~\new_[8500]_ ;
  assign \new_[6247]_  = ~\new_[18124]_  | (~\new_[8668]_  & ~\new_[14168]_ );
  assign \new_[6248]_  = ~\new_[11002]_  | ~\new_[12863]_  | ~\new_[9190]_  | ~\new_[8883]_ ;
  assign \new_[6249]_  = \\u0_r0_out_reg[26] ;
  assign \new_[6250]_  = \\u0_r0_out_reg[27] ;
  assign \new_[6251]_  = ~\new_[6995]_ ;
  assign \new_[6252]_  = ~\new_[13547]_  | ~\new_[8560]_  | ~\new_[8558]_ ;
  assign \new_[6253]_  = ~\new_[15115]_  | (~\new_[8561]_  & ~\new_[19217]_ );
  assign \new_[6254]_  = \new_[8255]_  | \new_[15530]_ ;
  assign \new_[6255]_  = ~\new_[9471]_  & ~\new_[8158]_ ;
  assign \new_[6256]_  = ~\new_[10852]_  & ~\new_[8154]_ ;
  assign \new_[6257]_  = ~\new_[7526]_  & ~\new_[9372]_ ;
  assign \new_[6258]_  = ~\new_[11412]_  | (~\new_[8632]_  & ~\new_[19780]_ );
  assign \new_[6259]_  = ~\new_[9194]_  & ~\new_[8218]_ ;
  assign \new_[6260]_  = ~\new_[8135]_  | ~\new_[17789]_ ;
  assign \new_[6261]_  = ~\new_[14822]_  | (~\new_[8669]_  & ~\new_[13391]_ );
  assign \new_[6262]_  = ~\new_[9205]_  & ~\new_[8220]_ ;
  assign \new_[6263]_  = ~\new_[8126]_  & (~\new_[16540]_  | ~\new_[18465]_ );
  assign \new_[6264]_  = (~\new_[8702]_  | ~\new_[19433]_ ) & (~\new_[8962]_  | ~\new_[17801]_ );
  assign \new_[6265]_  = ~\new_[7553]_  & ~\new_[8069]_ ;
  assign \new_[6266]_  = ~\new_[9776]_  | ~\new_[14125]_  | ~\new_[10112]_  | ~\new_[13957]_ ;
  assign \new_[6267]_  = ~\new_[7984]_  & ~\new_[8212]_ ;
  assign \new_[6268]_  = ~\new_[9948]_  | ~\new_[11966]_  | ~\new_[10439]_  | ~\new_[9091]_ ;
  assign \new_[6269]_  = ~\new_[17041]_  | (~\new_[8706]_  & ~\new_[12523]_ );
  assign \new_[6270]_  = ~\new_[7013]_ ;
  assign \new_[6271]_  = ~\new_[7870]_  | ~\new_[8108]_ ;
  assign \new_[6272]_  = ~\new_[10141]_  & ~\new_[8122]_ ;
  assign \new_[6273]_  = ~\new_[13950]_  | ~\new_[14715]_  | ~\new_[9792]_  | ~\new_[9556]_ ;
  assign \new_[6274]_  = ~\new_[8251]_  | ~\new_[16394]_ ;
  assign \new_[6275]_  = ~\new_[12375]_  & (~\new_[8655]_  | ~\new_[21559]_ );
  assign \new_[6276]_  = ~\new_[8172]_  & (~\new_[15323]_  | ~\new_[19377]_ );
  assign \new_[6277]_  = ~\new_[8205]_  | ~\new_[11691]_ ;
  assign \new_[6278]_  = ~\new_[11908]_  & (~\new_[8648]_  | ~\new_[19405]_ );
  assign \new_[6279]_  = ~\new_[18821]_  | (~\new_[8833]_  & ~\new_[11099]_ );
  assign \new_[6280]_  = ~\new_[19381]_  | (~\new_[10195]_  & ~\new_[9071]_ );
  assign \new_[6281]_  = ~\new_[7550]_  | ~\new_[19088]_ ;
  assign \new_[6282]_  = ~\new_[20341]_  | (~\new_[8897]_  & ~\new_[11370]_ );
  assign \new_[6283]_  = ~\new_[8439]_  | ~\new_[19102]_ ;
  assign \new_[6284]_  = ~\new_[17689]_  | (~\new_[10175]_  & ~\new_[8919]_ );
  assign \new_[6285]_  = ~\new_[18070]_  | (~\new_[8860]_  & ~\new_[8988]_ );
  assign \new_[6286]_  = ~\new_[18077]_  | (~\new_[8995]_  & ~\new_[9106]_ );
  assign \new_[6287]_  = ~\new_[21556]_  | (~\new_[9009]_  & ~\new_[11263]_ );
  assign \new_[6288]_  = ~\new_[7460]_  | ~\new_[19711]_ ;
  assign \new_[6289]_  = ~\new_[19179]_  & (~\new_[9023]_  | ~\new_[9010]_ );
  assign \new_[6290]_  = ~\new_[7512]_  | ~\new_[19145]_ ;
  assign \new_[6291]_  = ~\new_[19233]_  | (~\new_[9081]_  & ~\new_[13198]_ );
  assign \new_[6292]_  = ~\new_[21631]_  | (~\new_[9087]_  & ~\new_[10628]_ );
  assign \new_[6293]_  = ~\new_[19299]_  | (~\new_[8905]_  & ~\new_[13274]_ );
  assign \new_[6294]_  = ~\new_[19247]_  | (~\new_[9099]_  & ~\new_[13188]_ );
  assign \new_[6295]_  = ~\new_[19015]_  | (~\new_[8938]_  & ~\new_[13034]_ );
  assign \new_[6296]_  = \new_[7626]_  | \new_[17874]_ ;
  assign \new_[6297]_  = ~\new_[18773]_  & (~\new_[8868]_  | ~\new_[15635]_ );
  assign \new_[6298]_  = \new_[7627]_  | \new_[20680]_ ;
  assign \new_[6299]_  = ~\new_[19619]_  & (~\new_[11902]_  | ~\new_[8770]_ );
  assign \new_[6300]_  = \new_[7671]_  | \new_[18124]_ ;
  assign \new_[6301]_  = \new_[7678]_  | \new_[18798]_ ;
  assign \new_[6302]_  = \new_[7688]_  & \new_[18498]_ ;
  assign \new_[6303]_  = \new_[7680]_  | \new_[17837]_ ;
  assign \new_[6304]_  = ~\new_[21557]_  & (~\new_[8791]_  | ~\new_[20390]_ );
  assign \new_[6305]_  = ~\new_[19163]_  & (~\new_[11760]_  | ~\new_[8801]_ );
  assign \new_[6306]_  = ~\new_[19659]_  & (~\new_[13302]_  | ~\new_[8817]_ );
  assign \new_[6307]_  = \new_[7594]_  & \new_[19021]_ ;
  assign \new_[6308]_  = ~\new_[19519]_  | (~\new_[8895]_  & ~\new_[21612]_ );
  assign \new_[6309]_  = ~\new_[19612]_  & (~\new_[9027]_  | ~\new_[12301]_ );
  assign \new_[6310]_  = ~\new_[20842]_  | (~\new_[8996]_  & ~\new_[10300]_ );
  assign \new_[6311]_  = ~\new_[17796]_  | (~\new_[9057]_  & ~\new_[21592]_ );
  assign \new_[6312]_  = ~\new_[19798]_  | (~\new_[9075]_  & ~\new_[11248]_ );
  assign \new_[6313]_  = ~\new_[21557]_  & (~\new_[9094]_  | ~\new_[10236]_ );
  assign \new_[6314]_  = ~\new_[8469]_  | ~\new_[19247]_ ;
  assign \new_[6315]_  = ~\new_[19357]_  | (~\new_[8989]_  & ~\new_[10464]_ );
  assign \new_[6316]_  = ~\new_[7747]_  | ~\new_[10779]_ ;
  assign \new_[6317]_  = \new_[7618]_  & \new_[10793]_ ;
  assign \new_[6318]_  = ~\new_[8372]_  | ~\new_[19492]_ ;
  assign \new_[6319]_  = ~\new_[8236]_  | ~\new_[14955]_ ;
  assign \new_[6320]_  = ~\new_[7633]_  | ~\new_[12569]_ ;
  assign \new_[6321]_  = ~\new_[7655]_  & ~\new_[8809]_ ;
  assign \new_[6322]_  = ~\new_[13120]_  & (~\new_[8886]_  | ~\new_[17874]_ );
  assign \new_[6323]_  = ~\new_[13032]_  & (~\new_[8933]_  | ~\new_[19064]_ );
  assign \new_[6324]_  = ~\new_[8713]_  | ~\new_[7600]_ ;
  assign \new_[6325]_  = ~\new_[7667]_  & ~\new_[8763]_ ;
  assign \new_[6326]_  = ~\new_[8471]_  | ~\new_[19320]_ ;
  assign \new_[6327]_  = ~\new_[7683]_  | ~\new_[14332]_ ;
  assign \new_[6328]_  = ~\new_[7750]_  | ~\new_[10798]_ ;
  assign \new_[6329]_  = ~\new_[12834]_  & (~\new_[9031]_  | ~\new_[18361]_ );
  assign \new_[6330]_  = ~\new_[12846]_  & (~\new_[9120]_  | ~\new_[18795]_ );
  assign \new_[6331]_  = ~\new_[8256]_  | ~\new_[11595]_ ;
  assign \new_[6332]_  = ~\new_[7060]_ ;
  assign \new_[6333]_  = ~\new_[7696]_  & ~\new_[12230]_ ;
  assign \new_[6334]_  = ~\new_[15167]_  & (~\new_[9034]_  | ~\new_[17472]_ );
  assign \new_[6335]_  = ~\new_[21556]_  & (~\new_[10553]_  | ~\new_[20557]_ );
  assign \new_[6336]_  = \new_[7634]_  & \new_[10819]_ ;
  assign \new_[6337]_  = ~\new_[8260]_  | ~\new_[11666]_ ;
  assign \new_[6338]_  = ~\new_[19439]_  | (~\new_[9110]_  & ~\new_[15047]_ );
  assign \new_[6339]_  = ~\new_[19095]_  | (~\new_[9108]_  & ~\new_[14871]_ );
  assign \new_[6340]_  = \new_[8421]_  & \new_[19156]_ ;
  assign \new_[6341]_  = ~\new_[7071]_ ;
  assign \new_[6342]_  = \new_[8420]_  & \new_[19203]_ ;
  assign \new_[6343]_  = ~\new_[19275]_  | (~\new_[8950]_  & ~\new_[14080]_ );
  assign \new_[6344]_  = ~\new_[21631]_  | (~\new_[9185]_  & ~\new_[14833]_ );
  assign \new_[6345]_  = ~\new_[21695]_  | (~\new_[8875]_  & ~\new_[14874]_ );
  assign \new_[6346]_  = ~\new_[9795]_  | ~\new_[8392]_ ;
  assign \new_[6347]_  = ~\new_[12121]_  | ~\new_[11545]_  | ~\new_[11087]_ ;
  assign \new_[6348]_  = ~\new_[8314]_  | ~\new_[15763]_ ;
  assign \new_[6349]_  = ~\new_[11785]_  & ~\new_[7774]_ ;
  assign \new_[6350]_  = ~\new_[8315]_  | ~\new_[19517]_ ;
  assign \new_[6351]_  = ~\new_[12027]_  | ~\new_[11095]_  | ~\new_[8740]_ ;
  assign \new_[6352]_  = ~\new_[7086]_ ;
  assign \new_[6353]_  = \new_[8338]_  & \new_[18873]_ ;
  assign \new_[6354]_  = ~\new_[7087]_ ;
  assign \new_[6355]_  = ~\new_[18644]_  | (~\new_[9153]_  & ~\new_[13278]_ );
  assign \new_[6356]_  = ~\new_[7088]_ ;
  assign \new_[6357]_  = ~\new_[8433]_  | ~\new_[17770]_ ;
  assign \new_[6358]_  = ~\new_[17845]_  | (~\new_[9170]_  & ~\new_[12970]_ );
  assign \new_[6359]_  = ~\new_[8367]_  | ~\new_[14986]_ ;
  assign \new_[6360]_  = \new_[8269]_  & \new_[10173]_ ;
  assign \new_[6361]_  = ~\new_[11678]_  | ~\new_[8754]_  | ~\new_[11862]_ ;
  assign \new_[6362]_  = ~\new_[12572]_  | ~\new_[11644]_  | ~\new_[9144]_ ;
  assign \new_[6363]_  = \new_[8269]_  & \new_[10959]_ ;
  assign \new_[6364]_  = \new_[8277]_  & \new_[12377]_ ;
  assign \new_[6365]_  = ~\new_[19261]_  & (~\new_[8840]_  | ~\new_[16859]_ );
  assign \new_[6366]_  = \new_[8337]_  & \new_[19547]_ ;
  assign \new_[6367]_  = ~\new_[7630]_  | ~\new_[18011]_ ;
  assign \new_[6368]_  = \new_[7889]_  & \new_[14966]_ ;
  assign \new_[6369]_  = ~\new_[8382]_  & (~\new_[16198]_  | ~\new_[19547]_ );
  assign \new_[6370]_  = ~\new_[7109]_ ;
  assign \new_[6371]_  = \new_[11165]_  | \new_[8382]_ ;
  assign \new_[6372]_  = ~\new_[8273]_  & (~\new_[10176]_  | ~\new_[18187]_ );
  assign \new_[6373]_  = ~\new_[8274]_  | ~\new_[8837]_ ;
  assign \new_[6374]_  = \new_[8394]_  & \new_[19239]_ ;
  assign \new_[6375]_  = ~\new_[19079]_  | (~\new_[9039]_  & ~\new_[15579]_ );
  assign \new_[6376]_  = ~\new_[19215]_  | (~\new_[9213]_  & ~\new_[11873]_ );
  assign \new_[6377]_  = ~\new_[9542]_  | ~\new_[8272]_ ;
  assign \new_[6378]_  = ~\new_[19612]_  | (~\new_[8836]_  & ~\new_[16474]_ );
  assign \new_[6379]_  = ~\new_[7120]_ ;
  assign \new_[6380]_  = \new_[12208]_  & \new_[8392]_ ;
  assign \new_[6381]_  = ~\new_[7646]_  | ~\new_[19440]_ ;
  assign \new_[6382]_  = ~\new_[8881]_  | ~\new_[8334]_ ;
  assign \new_[6383]_  = ~\new_[7981]_  | ~\new_[19404]_ ;
  assign \new_[6384]_  = ~\new_[9550]_  | ~\new_[8264]_ ;
  assign \new_[6385]_  = ~\new_[7468]_  | ~\new_[18649]_ ;
  assign \new_[6386]_  = ~\new_[11554]_  | ~\new_[11565]_  | ~\new_[11207]_ ;
  assign \new_[6387]_  = ~\new_[7652]_  | ~\new_[19492]_ ;
  assign \new_[6388]_  = \new_[7721]_  | \new_[19145]_ ;
  assign \new_[6389]_  = ~\new_[7656]_  | ~\new_[20982]_ ;
  assign \new_[6390]_  = ~\new_[7728]_  & ~\new_[10032]_ ;
  assign \new_[6391]_  = ~\new_[8380]_  & ~\new_[14845]_ ;
  assign \new_[6392]_  = ~\new_[8233]_  | ~\new_[15777]_ ;
  assign \new_[6393]_  = ~\new_[8772]_  | ~\new_[11066]_  | ~\new_[9870]_ ;
  assign \new_[6394]_  = \new_[13558]_  & \new_[8371]_ ;
  assign \new_[6395]_  = ~\new_[17818]_  | (~\new_[8958]_  & ~\new_[12981]_ );
  assign \new_[6396]_  = ~\new_[7141]_ ;
  assign \new_[6397]_  = ~\new_[7143]_ ;
  assign \new_[6398]_  = ~\new_[14694]_  | ~\new_[12682]_  | ~\new_[8775]_ ;
  assign \new_[6399]_  = ~\new_[11533]_  | ~\new_[11500]_  | ~\new_[11095]_ ;
  assign \new_[6400]_  = ~\new_[8657]_  | ~\new_[7910]_ ;
  assign \new_[6401]_  = ~\new_[21115]_  & (~\new_[9006]_  | ~\new_[15053]_ );
  assign \new_[6402]_  = ~\new_[8489]_  | ~\new_[17549]_ ;
  assign \new_[6403]_  = ~\new_[18418]_  | (~\new_[9017]_  & ~\new_[11414]_ );
  assign \new_[6404]_  = ~\new_[19436]_  | (~\new_[9000]_  & ~\new_[16386]_ );
  assign \new_[6405]_  = ~\new_[7163]_ ;
  assign \new_[6406]_  = \new_[8458]_  & \new_[19241]_ ;
  assign \new_[6407]_  = ~\new_[19247]_  | (~\new_[8954]_  & ~\new_[13414]_ );
  assign \new_[6408]_  = ~\new_[19247]_  | ~\new_[984]_  | ~\new_[9174]_ ;
  assign \new_[6409]_  = ~\new_[7755]_  & ~\new_[11003]_ ;
  assign \new_[6410]_  = ~\new_[7481]_  | ~\new_[8792]_ ;
  assign \new_[6411]_  = ~\new_[18627]_  | (~\new_[8926]_  & ~\new_[15877]_ );
  assign \new_[6412]_  = ~\new_[7169]_ ;
  assign \new_[6413]_  = ~\new_[17757]_  | ~\new_[16210]_  | ~\new_[7786]_  | ~\new_[9200]_ ;
  assign \new_[6414]_  = ~\new_[7170]_ ;
  assign \new_[6415]_  = ~\new_[19266]_  | (~\new_[9111]_  & ~\new_[15627]_ );
  assign \new_[6416]_  = ~\new_[19450]_  | ~\new_[19517]_  | ~\new_[9172]_ ;
  assign \new_[6417]_  = ~\new_[18077]_  & (~\new_[8942]_  | ~\new_[9186]_ );
  assign \new_[6418]_  = ~\new_[7708]_  | ~\new_[13652]_ ;
  assign \new_[6419]_  = ~\new_[19687]_  & (~\new_[9072]_  | ~\new_[12249]_ );
  assign \new_[6420]_  = ~\new_[7178]_ ;
  assign \new_[6421]_  = ~\new_[8428]_  | ~\new_[946]_ ;
  assign \new_[6422]_  = ~\new_[7181]_ ;
  assign \new_[6423]_  = ~\new_[21562]_  | (~\new_[9015]_  & ~\new_[15958]_ );
  assign \new_[6424]_  = ~\new_[7713]_  | ~\new_[18418]_ ;
  assign \new_[6425]_  = ~\new_[7735]_  | ~\new_[19170]_ ;
  assign \new_[6426]_  = ~\new_[7184]_ ;
  assign \new_[6427]_  = ~\new_[7736]_  | ~\new_[19748]_ ;
  assign \new_[6428]_  = ~\new_[7955]_  | ~\new_[7486]_ ;
  assign \new_[6429]_  = ~\new_[8463]_  | ~\new_[944]_ ;
  assign \new_[6430]_  = ~\new_[9112]_  | ~\new_[7535]_ ;
  assign \new_[6431]_  = ~\new_[11578]_  | ~\new_[11516]_  | ~\new_[11366]_ ;
  assign \new_[6432]_  = ~\new_[7732]_  | ~\new_[18293]_ ;
  assign \new_[6433]_  = ~\new_[7540]_  | ~\new_[19530]_ ;
  assign \new_[6434]_  = ~\new_[7737]_  | ~\new_[19659]_ ;
  assign \new_[6435]_  = ~\new_[7959]_  | ~\new_[7541]_ ;
  assign \new_[6436]_  = ~\new_[9103]_  | ~\new_[7549]_ ;
  assign \new_[6437]_  = ~\new_[18086]_  | (~\new_[9133]_  & ~\new_[13188]_ );
  assign \new_[6438]_  = ~\new_[7197]_ ;
  assign \new_[6439]_  = ~\new_[8801]_  | ~\new_[10655]_  | ~\new_[12986]_ ;
  assign \new_[6440]_  = ~\new_[7199]_ ;
  assign \new_[6441]_  = ~\new_[11346]_  & ~\new_[7564]_ ;
  assign \new_[6442]_  = ~\new_[7725]_  & ~\new_[7906]_ ;
  assign \new_[6443]_  = ~\new_[19612]_  | (~\new_[9219]_  & ~\new_[10705]_ );
  assign \new_[6444]_  = ~\new_[13642]_  | ~\new_[8404]_  | ~\new_[12551]_ ;
  assign \new_[6445]_  = ~\new_[11681]_  | ~\new_[11644]_  | ~\new_[9144]_ ;
  assign \new_[6446]_  = ~\new_[19625]_  & (~\new_[9149]_  | ~\new_[12294]_ );
  assign \new_[6447]_  = ~\new_[7602]_  | ~\new_[12515]_ ;
  assign \new_[6448]_  = ~\new_[7204]_ ;
  assign \new_[6449]_  = ~\new_[7729]_  | ~\new_[14067]_ ;
  assign \new_[6450]_  = ~\new_[9141]_  | ~\new_[7584]_ ;
  assign \new_[6451]_  = ~\new_[9038]_  | ~\new_[7590]_ ;
  assign \new_[6452]_  = ~\new_[7211]_ ;
  assign \new_[6453]_  = ~\new_[11387]_  & ~\new_[7595]_ ;
  assign \new_[6454]_  = ~\new_[18967]_  | (~\new_[9136]_  & ~\new_[14795]_ );
  assign \new_[6455]_  = ~\new_[8393]_  & ~\new_[8913]_ ;
  assign \new_[6456]_  = \new_[7742]_  | \new_[12894]_ ;
  assign \new_[6457]_  = ~\new_[12237]_  | ~\new_[7905]_  | ~\new_[11243]_ ;
  assign \new_[6458]_  = ~\new_[10199]_  | ~\new_[11987]_  | ~\new_[9016]_ ;
  assign \new_[6459]_  = ~\new_[14376]_  | ~\new_[12691]_  | ~\new_[7928]_  | ~\new_[9929]_ ;
  assign \new_[6460]_  = ~\new_[7495]_  & ~\new_[10076]_ ;
  assign \new_[6461]_  = ~\new_[11966]_  | ~\new_[10538]_  | ~\new_[9066]_  | ~\new_[9948]_ ;
  assign \new_[6462]_  = ~\new_[12193]_  | ~\new_[11528]_  | ~\new_[7935]_  | ~\new_[12920]_ ;
  assign \new_[6463]_  = ~\new_[7222]_ ;
  assign \new_[6464]_  = ~\new_[9965]_  | ~\new_[7956]_  | ~\new_[8920]_ ;
  assign \new_[6465]_  = ~\new_[19612]_  & (~\new_[9209]_  | ~\new_[11523]_ );
  assign \new_[6466]_  = ~\new_[7078]_ ;
  assign \new_[6467]_  = ~\new_[19247]_  & (~\new_[9224]_  | ~\new_[12688]_ );
  assign \new_[6468]_  = ~\new_[7482]_  | ~\new_[19148]_ ;
  assign \new_[6469]_  = ~\new_[7642]_  | ~\new_[19222]_ ;
  assign \new_[6470]_  = ~\new_[19469]_  | (~\new_[9155]_  & ~\new_[15591]_ );
  assign \new_[6471]_  = \new_[8319]_  & \new_[19208]_ ;
  assign \new_[6472]_  = ~\new_[20486]_  | (~\new_[16965]_  & ~\new_[8838]_ );
  assign \new_[6473]_  = ~\new_[7945]_  & ~\new_[11758]_ ;
  assign \new_[6474]_  = ~\new_[8325]_  | ~\new_[18762]_ ;
  assign \new_[6475]_  = \new_[8322]_  & \new_[21115]_ ;
  assign \new_[6476]_  = ~\new_[8340]_  & (~\new_[10472]_  | ~\new_[19525]_ );
  assign \new_[6477]_  = ~\new_[8347]_  | (~\new_[15668]_  & ~\new_[18998]_ );
  assign \new_[6478]_  = ~\new_[7558]_  | (~\new_[13667]_  & ~\new_[18194]_ );
  assign \new_[6479]_  = ~\new_[21497]_  | (~\new_[16984]_  & ~\new_[9164]_ );
  assign \new_[6480]_  = \new_[8358]_  & \new_[18606]_ ;
  assign \new_[6481]_  = ~\new_[8360]_  | ~\new_[19204]_ ;
  assign \new_[6482]_  = ~\new_[15966]_  & (~\new_[8921]_  | ~\new_[19471]_ );
  assign \new_[6483]_  = ~\new_[20680]_  | (~\new_[21612]_  & ~\new_[12643]_ );
  assign \new_[6484]_  = ~\new_[8364]_  | (~\new_[14542]_  & ~\new_[18965]_ );
  assign \new_[6485]_  = ~\new_[8368]_  | ~\new_[17874]_ ;
  assign \new_[6486]_  = ~\new_[7614]_  | ~\new_[19260]_ ;
  assign \new_[6487]_  = ~\new_[18992]_  & (~\new_[8869]_  | ~\new_[17104]_ );
  assign \new_[6488]_  = ~\new_[10132]_  | (~\new_[8864]_  & ~\new_[18967]_ );
  assign \new_[6489]_  = \new_[11810]_  & \new_[8387]_ ;
  assign \new_[6490]_  = ~\new_[12885]_  | ~\new_[7866]_  | ~\new_[8891]_ ;
  assign \new_[6491]_  = ~\new_[19440]_  & (~\new_[10112]_  | ~\new_[12503]_ );
  assign \new_[6492]_  = ~\new_[8814]_  | ~\new_[10637]_  | ~\new_[10594]_ ;
  assign \new_[6493]_  = ~\new_[9586]_  & ~\new_[7647]_ ;
  assign \new_[6494]_  = ~\new_[7660]_  & ~\new_[11931]_ ;
  assign \new_[6495]_  = ~\new_[18481]_  & (~\new_[15577]_  | ~\new_[11100]_ );
  assign \new_[6496]_  = ~\new_[11189]_  | ~\new_[10462]_  | ~\new_[10972]_  | ~\new_[15254]_ ;
  assign \new_[6497]_  = ~\new_[18442]_  & (~\new_[9113]_  | ~\new_[14493]_ );
  assign \new_[6498]_  = ~\new_[8447]_  | ~\new_[18572]_ ;
  assign \new_[6499]_  = \new_[8452]_  & \new_[21556]_ ;
  assign \new_[6500]_  = ~\new_[8460]_  | ~\new_[17837]_ ;
  assign \new_[6501]_  = ~\new_[19233]_  | (~\new_[21592]_  & ~\new_[12671]_ );
  assign \new_[6502]_  = ~\new_[10876]_  | (~\new_[8985]_  & ~\new_[18692]_ );
  assign \new_[6503]_  = ~\new_[18270]_  | (~\new_[8991]_  & ~\new_[13588]_ );
  assign \new_[6504]_  = ~\new_[8473]_  | ~\new_[17472]_ ;
  assign \new_[6505]_  = ~\new_[8480]_  | ~\new_[21629]_ ;
  assign \new_[6506]_  = ~\new_[7681]_  | ~\new_[12743]_ ;
  assign \new_[6507]_  = ~\new_[18032]_  & (~\new_[9008]_  | ~\new_[14742]_ );
  assign \new_[6508]_  = ~\new_[10178]_  | (~\new_[8946]_  & ~\new_[21115]_ );
  assign \new_[6509]_  = ~\new_[8488]_  | ~\new_[19170]_ ;
  assign \new_[6510]_  = ~\new_[8490]_  | ~\new_[21558]_ ;
  assign \new_[6511]_  = ~\new_[7465]_  & (~\new_[10484]_  | ~\new_[18769]_ );
  assign \new_[6512]_  = ~\new_[15274]_  | ~\new_[7931]_  | ~\new_[9044]_ ;
  assign \new_[6513]_  = ~\new_[7484]_  | ~\new_[18070]_ ;
  assign \new_[6514]_  = ~\new_[7689]_  | ~\new_[18728]_ ;
  assign \new_[6515]_  = ~\new_[7490]_  | ~\new_[21631]_ ;
  assign \new_[6516]_  = ~\new_[18783]_  | (~\new_[8910]_  & ~\new_[20925]_ );
  assign \new_[6517]_  = ~\new_[7865]_  | (~\new_[13648]_  & ~\new_[21629]_ );
  assign \new_[6518]_  = ~\new_[7493]_  | ~\new_[21557]_ ;
  assign \new_[6519]_  = ~\new_[14347]_  | ~\new_[10277]_  | ~\new_[8825]_ ;
  assign \new_[6520]_  = ~\new_[11301]_  | ~\new_[8795]_  | ~\new_[10516]_ ;
  assign \new_[6521]_  = \new_[7510]_  & \new_[18280]_ ;
  assign \new_[6522]_  = ~\new_[13922]_  | ~\new_[11840]_  | ~\new_[7900]_  | ~\new_[15403]_ ;
  assign \new_[6523]_  = ~\new_[9437]_  | (~\new_[9266]_  & ~\new_[1081]_ );
  assign \new_[6524]_  = ~\new_[8355]_  | ~\new_[19378]_ ;
  assign \new_[6525]_  = ~\new_[7539]_  | ~\new_[18937]_ ;
  assign \new_[6526]_  = ~\new_[7544]_  | ~\new_[16879]_ ;
  assign \new_[6527]_  = ~\new_[7579]_  | ~\new_[19088]_ ;
  assign \new_[6528]_  = ~\new_[12217]_  | ~\new_[15358]_  | ~\new_[9176]_ ;
  assign \new_[6529]_  = ~\new_[8290]_  & ~\new_[9448]_ ;
  assign \new_[6530]_  = ~\new_[8402]_  & (~\new_[10482]_  | ~\new_[18827]_ );
  assign \new_[6531]_  = ~\new_[10933]_  | ~\new_[9207]_  | ~\new_[15371]_ ;
  assign \new_[6532]_  = \new_[7583]_  & \new_[18967]_ ;
  assign \new_[6533]_  = ~\new_[7586]_  | ~\new_[18650]_ ;
  assign \new_[6534]_  = ~\new_[8650]_  & (~\new_[9249]_  | ~\new_[19659]_ );
  assign \new_[6535]_  = ~\new_[7592]_  | ~\new_[17874]_ ;
  assign \new_[6536]_  = ~\new_[10286]_  | ~\new_[10469]_  | ~\new_[10963]_  | ~\new_[15375]_ ;
  assign \new_[6537]_  = ~\new_[7598]_  | ~\new_[19529]_ ;
  assign \new_[6538]_  = ~\new_[9428]_  | ~\new_[8296]_ ;
  assign \new_[6539]_  = \new_[9430]_  | \new_[8297]_ ;
  assign \new_[6540]_  = \new_[8261]_  | \new_[8300]_ ;
  assign \new_[6541]_  = ~\new_[11900]_  | ~\new_[12665]_  | ~\new_[7795]_  | ~\new_[14056]_ ;
  assign \new_[6542]_  = ~\new_[7533]_  | ~\new_[17585]_ ;
  assign \new_[6543]_  = ~\new_[7559]_  | ~\new_[17041]_ ;
  assign \new_[6544]_  = ~\new_[11770]_  | ~\new_[9994]_  | ~\new_[10572]_  | ~\new_[11736]_ ;
  assign \new_[6545]_  = ~\new_[10549]_  | ~\new_[13716]_  | ~\new_[12540]_  | ~\new_[16204]_ ;
  assign \new_[6546]_  = ~\new_[10368]_  | ~\new_[17785]_  | ~\new_[14076]_  | ~\new_[13794]_ ;
  assign \new_[6547]_  = ~\new_[9839]_  | ~\new_[13800]_  | ~\new_[11212]_  | ~\new_[14092]_ ;
  assign \new_[6548]_  = ~\new_[9813]_  | ~\new_[13936]_  | ~\new_[11388]_  | ~\new_[14176]_ ;
  assign \new_[6549]_  = ~\new_[12762]_  & ~\new_[8446]_ ;
  assign \new_[6550]_  = ~\new_[13281]_  | ~\new_[8407]_  | ~\new_[9989]_ ;
  assign \new_[6551]_  = ~\new_[9995]_  | ~\new_[13758]_  | ~\new_[12366]_  | ~\new_[15232]_ ;
  assign \new_[6552]_  = ~\new_[11577]_  & ~\new_[7576]_ ;
  assign \new_[6553]_  = ~\new_[19509]_  | ~\new_[8336]_  | ~\new_[18569]_ ;
  assign \new_[6554]_  = ~\new_[19467]_  | ~\new_[8418]_  | ~\new_[17381]_ ;
  assign \new_[6555]_  = ~\new_[19433]_  | ~\new_[8478]_  | ~\new_[18077]_ ;
  assign \new_[6556]_  = ~\new_[16886]_  | (~\new_[9208]_  & ~\new_[11112]_ );
  assign \new_[6557]_  = \new_[7605]_  | \new_[17385]_ ;
  assign \new_[6558]_  = ~\new_[17478]_  | (~\new_[9212]_  & ~\new_[11134]_ );
  assign \new_[6559]_  = ~\new_[7861]_  & ~\new_[8262]_ ;
  assign \new_[6560]_  = ~\new_[10084]_  & ~\new_[8263]_ ;
  assign \new_[6561]_  = \new_[7606]_  | \new_[18537]_ ;
  assign \new_[6562]_  = ~\new_[17323]_  | (~\new_[9226]_  & ~\new_[11219]_ );
  assign \new_[6563]_  = \new_[7607]_  | \new_[18373]_ ;
  assign \new_[6564]_  = ~\new_[18300]_  | (~\new_[9221]_  & ~\new_[10129]_ );
  assign \new_[6565]_  = ~\new_[8907]_  & ~\new_[8280]_ ;
  assign \new_[6566]_  = ~\new_[8984]_  & ~\new_[8291]_ ;
  assign \new_[6567]_  = ~\new_[7912]_  & ~\new_[9451]_ ;
  assign \new_[6568]_  = ~\new_[7609]_  | ~\new_[17789]_ ;
  assign \new_[6569]_  = ~\new_[7926]_  | (~\new_[11464]_  & ~\new_[17115]_ );
  assign \new_[6570]_  = ~\new_[10259]_  & ~\new_[8281]_ ;
  assign \new_[6571]_  = ~\new_[10316]_  & ~\new_[7712]_ ;
  assign \new_[6572]_  = \new_[17390]_  | \new_[7612]_ ;
  assign \new_[6573]_  = ~\new_[7596]_  | ~\new_[17323]_ ;
  assign \new_[6574]_  = (~\new_[9177]_  | ~\new_[17689]_ ) & (~\new_[17468]_  | ~\new_[15572]_ );
  assign \new_[6575]_  = (~\new_[9179]_  | ~\new_[21558]_ ) & (~\new_[18120]_  | ~\new_[15953]_ );
  assign \new_[6576]_  = ~\new_[10099]_  & ~\new_[8246]_ ;
  assign \new_[6577]_  = ~\new_[21196]_  | ~\new_[8854]_  | ~\new_[10414]_ ;
  assign \new_[6578]_  = ~\new_[21470]_  | ~\new_[7929]_  | ~\new_[9789]_ ;
  assign \new_[6579]_  = ~\new_[7885]_  | ~\new_[10133]_  | ~\new_[9790]_ ;
  assign \new_[6580]_  = ~\new_[10067]_  | ~\new_[9788]_  | ~\new_[7853]_ ;
  assign \new_[6581]_  = ~\new_[8893]_  | ~\new_[8953]_  | ~\new_[8734]_ ;
  assign \new_[6582]_  = ~\new_[12596]_  | ~\new_[9813]_  | ~\new_[10942]_  | ~\new_[14176]_ ;
  assign \new_[6583]_  = ~\new_[13952]_  | ~\new_[9995]_  | ~\new_[10929]_  | ~\new_[15232]_ ;
  assign \new_[6584]_  = ~\new_[7477]_  & ~\new_[9648]_ ;
  assign \new_[6585]_  = ~\new_[10198]_  | ~\new_[7902]_  | ~\new_[9793]_ ;
  assign \new_[6586]_  = ~\new_[19952]_  | ~\new_[7942]_  | ~\new_[9192]_ ;
  assign \new_[6587]_  = ~\new_[19836]_  | ~\new_[7937]_  | ~\new_[10882]_ ;
  assign \new_[6588]_  = ~\new_[10269]_  | ~\new_[10268]_  | ~\new_[9198]_ ;
  assign \new_[6589]_  = ~\new_[15289]_  | ~\new_[9900]_  | ~\new_[10403]_  | ~\new_[11375]_ ;
  assign \new_[6590]_  = ~\new_[12601]_  | ~\new_[9839]_  | ~\new_[10900]_  | ~\new_[14092]_ ;
  assign \new_[6591]_  = ~\new_[10519]_  | ~\new_[15830]_  | ~\new_[12310]_  | ~\new_[11656]_ ;
  assign \new_[6592]_  = ~\new_[12306]_  | ~\new_[12500]_  | ~\new_[8946]_ ;
  assign \new_[6593]_  = ~\new_[13802]_  | ~\new_[8317]_  | ~\new_[9806]_ ;
  assign \new_[6594]_  = ~\new_[8326]_  & ~\new_[8327]_ ;
  assign \new_[6595]_  = ~\new_[13719]_  | ~\new_[7569]_  | ~\new_[9858]_ ;
  assign \new_[6596]_  = ~\new_[11364]_  | ~\new_[12681]_  | ~\new_[8864]_ ;
  assign \new_[6597]_  = ~\new_[8413]_  & ~\new_[9558]_ ;
  assign \new_[6598]_  = ~\new_[8467]_  & ~\new_[9601]_ ;
  assign \new_[6599]_  = ~\new_[13714]_  | ~\new_[7462]_  | ~\new_[20714]_ ;
  assign \new_[6600]_  = ~\new_[11032]_  & ~\new_[7527]_ ;
  assign \new_[6601]_  = ~\new_[7528]_  & (~\new_[11567]_  | ~\new_[19107]_ );
  assign \new_[6602]_  = \new_[8441]_  & \new_[11658]_ ;
  assign \new_[6603]_  = ~\new_[8695]_  | ~\new_[8254]_ ;
  assign \new_[6604]_  = ~\new_[7474]_  & (~\new_[11009]_  | ~\new_[21638]_ );
  assign \new_[6605]_  = \new_[17116]_  ^ \new_[19408]_ ;
  assign \new_[6606]_  = \new_[15062]_  ^ \new_[19045]_ ;
  assign \new_[6607]_  = \new_[14782]_  ^ \new_[18773]_ ;
  assign \new_[6608]_  = ~\new_[7353]_ ;
  assign \new_[6609]_  = ~\new_[8764]_  & ~\new_[21115]_ ;
  assign \new_[6610]_  = \new_[7883]_  | \new_[19156]_ ;
  assign \new_[6611]_  = ~\new_[9857]_  & ~\new_[19102]_ ;
  assign \new_[6612]_  = ~\new_[7361]_ ;
  assign \new_[6613]_  = ~\new_[7371]_ ;
  assign \new_[6614]_  = ~\new_[11495]_  | ~\new_[12980]_  | ~\new_[10543]_  | ~\new_[11361]_ ;
  assign \new_[6615]_  = ~\new_[7376]_ ;
  assign \new_[6616]_  = \new_[8007]_  | \new_[18967]_ ;
  assign \new_[6617]_  = ~\new_[7839]_  | ~\new_[10594]_ ;
  assign \new_[6618]_  = ~\new_[7384]_ ;
  assign \new_[6619]_  = ~\new_[7930]_  | ~\new_[13313]_ ;
  assign \new_[6620]_  = \new_[7842]_  | \new_[19079]_ ;
  assign \new_[6621]_  = ~\new_[9861]_  | ~\new_[20940]_ ;
  assign \new_[6622]_  = ~\new_[7877]_  | ~\new_[10005]_ ;
  assign \new_[6623]_  = ~\new_[7843]_  | ~\new_[12282]_ ;
  assign \new_[6624]_  = ~\new_[7830]_  | ~\new_[17089]_ ;
  assign \new_[6625]_  = ~\new_[7851]_  | ~\new_[18380]_ ;
  assign \new_[6626]_  = ~\new_[7401]_ ;
  assign \new_[6627]_  = \new_[7864]_  & \new_[18194]_ ;
  assign \new_[6628]_  = ~\new_[7410]_ ;
  assign \new_[6629]_  = ~\new_[7856]_  | ~\new_[18965]_ ;
  assign \new_[6630]_  = \new_[8008]_  | \new_[21115]_ ;
  assign \new_[6631]_  = \new_[10963]_  & \new_[7820]_ ;
  assign \new_[6632]_  = ~\new_[7850]_  | ~\new_[18941]_ ;
  assign \new_[6633]_  = ~\new_[10282]_  & ~\new_[11351]_ ;
  assign \new_[6634]_  = ~\new_[7957]_  | ~\new_[10664]_ ;
  assign \new_[6635]_  = ~\new_[11102]_  & ~\new_[7971]_ ;
  assign \new_[6636]_  = ~\new_[11074]_  & ~\new_[12617]_ ;
  assign \new_[6637]_  = ~\new_[9985]_  | ~\new_[10004]_ ;
  assign \new_[6638]_  = \new_[7794]_  & \new_[7779]_ ;
  assign \new_[6639]_  = ~\new_[7891]_  | ~\new_[13272]_ ;
  assign \new_[6640]_  = ~\new_[14197]_  | ~\new_[9306]_  | ~\new_[21173]_ ;
  assign \new_[6641]_  = ~\new_[13270]_  | ~\new_[7779]_ ;
  assign \new_[6642]_  = ~\new_[8013]_  | ~\new_[19659]_ ;
  assign \new_[6643]_  = ~\new_[9876]_  | ~\new_[9857]_ ;
  assign \new_[6644]_  = \new_[7788]_  & \new_[7818]_ ;
  assign \new_[6645]_  = \new_[21298]_  | \new_[21631]_ ;
  assign \new_[6646]_  = ~\new_[7936]_  | ~\new_[19215]_ ;
  assign \new_[6647]_  = ~\new_[9896]_  & ~\new_[9996]_ ;
  assign \new_[6648]_  = ~\new_[7898]_  | ~\new_[11901]_ ;
  assign \new_[6649]_  = ~\new_[18171]_  & (~\new_[9289]_  | ~\new_[13339]_ );
  assign \new_[6650]_  = ~\new_[7435]_ ;
  assign \new_[6651]_  = ~\new_[10184]_  | ~\new_[10041]_ ;
  assign \new_[6652]_  = ~\new_[7443]_ ;
  assign \new_[6653]_  = ~\new_[7903]_  | ~\new_[19384]_ ;
  assign \new_[6654]_  = ~\new_[20622]_  & (~\new_[9325]_  | ~\new_[12069]_ );
  assign \new_[6655]_  = \new_[8010]_  | \new_[21558]_ ;
  assign \new_[6656]_  = \new_[8001]_  | \new_[19202]_ ;
  assign \new_[6657]_  = ~\new_[18077]_  & (~\new_[9291]_  | ~\new_[14964]_ );
  assign \new_[6658]_  = ~\new_[7917]_  | ~\new_[12856]_ ;
  assign \new_[6659]_  = \new_[7973]_  | \new_[21631]_ ;
  assign \new_[6660]_  = ~\new_[10517]_  | ~\new_[14215]_  | ~\new_[12524]_  | ~\new_[12424]_ ;
  assign \new_[6661]_  = ~\new_[11281]_  | ~\new_[11381]_ ;
  assign \new_[6662]_  = ~\new_[19687]_  | (~\new_[10678]_  & ~\new_[15430]_ );
  assign \new_[6663]_  = ~\new_[9183]_  & ~\new_[12957]_ ;
  assign \new_[6664]_  = ~\new_[10559]_  | ~\new_[9279]_  | ~\new_[15785]_ ;
  assign \new_[6665]_  = ~\new_[9236]_  | ~\new_[19054]_ ;
  assign \new_[6666]_  = ~\new_[7470]_ ;
  assign \new_[6667]_  = ~\new_[17172]_  | ~\new_[9302]_  | ~\new_[15142]_ ;
  assign \new_[6668]_  = ~\new_[8788]_  | ~\new_[12210]_ ;
  assign \new_[6669]_  = \new_[9036]_  | \new_[18795]_ ;
  assign \new_[6670]_  = ~\new_[8983]_  | ~\new_[21557]_ ;
  assign \new_[6671]_  = ~\new_[11218]_  & ~\new_[8851]_ ;
  assign \new_[6672]_  = ~\new_[14320]_  & ~\new_[10957]_ ;
  assign \new_[6673]_  = ~\new_[9237]_  | ~\new_[21556]_ ;
  assign \new_[6674]_  = ~\new_[11011]_  | ~\new_[21558]_ ;
  assign \new_[6675]_  = ~\new_[7481]_ ;
  assign \new_[6676]_  = ~\new_[7486]_ ;
  assign \new_[6677]_  = ~\new_[8828]_  | ~\new_[11094]_ ;
  assign \new_[6678]_  = ~\new_[7496]_ ;
  assign \new_[6679]_  = ~\new_[14191]_  & ~\new_[8821]_ ;
  assign \new_[6680]_  = ~\new_[10596]_  | ~\new_[10732]_  | ~\new_[10593]_ ;
  assign \new_[6681]_  = \new_[11185]_  & \new_[19145]_ ;
  assign \new_[6682]_  = ~\new_[19357]_  & (~\new_[10592]_  | ~\new_[13912]_ );
  assign \new_[6683]_  = ~\new_[7506]_ ;
  assign \new_[6684]_  = ~\new_[10659]_  | ~\new_[9304]_  | ~\new_[10627]_ ;
  assign \new_[6685]_  = ~\new_[15111]_  & ~\new_[21299]_ ;
  assign \new_[6686]_  = ~\new_[9079]_  & ~\new_[14312]_ ;
  assign \new_[6687]_  = ~\new_[12610]_  & ~\new_[9002]_ ;
  assign \new_[6688]_  = ~\new_[14037]_  | ~\new_[9303]_  | ~\new_[11764]_ ;
  assign \new_[6689]_  = ~\new_[8878]_  | ~\new_[19436]_ ;
  assign \new_[6690]_  = ~\new_[15488]_  & ~\new_[20435]_ ;
  assign \new_[6691]_  = \new_[10236]_  | \new_[21558]_ ;
  assign \new_[6692]_  = \new_[10236]_  & \new_[11594]_ ;
  assign \new_[6693]_  = ~\new_[9303]_  | ~\new_[11366]_ ;
  assign \new_[6694]_  = ~\new_[12150]_  & ~\new_[9130]_ ;
  assign \new_[6695]_  = ~\new_[9201]_  | ~\new_[21628]_ ;
  assign \new_[6696]_  = (~\new_[10582]_  | ~\new_[18175]_ ) & (~\new_[19199]_  | ~\new_[12729]_ );
  assign \new_[6697]_  = ~\new_[7535]_ ;
  assign \new_[6698]_  = ~\new_[9107]_  | ~\new_[17070]_ ;
  assign \new_[6699]_  = \new_[8920]_  | \new_[19163]_ ;
  assign \new_[6700]_  = ~\new_[20826]_ ;
  assign \new_[6701]_  = ~\new_[10112]_  & ~\new_[19115]_ ;
  assign \new_[6702]_  = ~\new_[14360]_  & ~\new_[20942]_ ;
  assign \new_[6703]_  = ~\new_[10897]_  | ~\new_[8783]_ ;
  assign \new_[6704]_  = ~\new_[7547]_ ;
  assign \new_[6705]_  = ~\new_[9122]_  | ~\new_[19145]_ ;
  assign \new_[6706]_  = ~\new_[7549]_ ;
  assign \new_[6707]_  = ~\new_[8796]_  | ~\new_[12991]_ ;
  assign \new_[6708]_  = ~\new_[15026]_  & ~\new_[9004]_ ;
  assign \new_[6709]_  = ~\new_[9238]_  | ~\new_[19257]_ ;
  assign \new_[6710]_  = ~\new_[9131]_  | ~\new_[19013]_ ;
  assign \new_[6711]_  = ~\new_[10996]_  | ~\new_[19247]_ ;
  assign \new_[6712]_  = ~\new_[9229]_  | ~\new_[19247]_ ;
  assign \new_[6713]_  = \new_[9054]_  | \new_[16889]_ ;
  assign \new_[6714]_  = ~\new_[16889]_  & (~\new_[10681]_  | ~\new_[12063]_ );
  assign \new_[6715]_  = ~\new_[11060]_  & ~\new_[12533]_ ;
  assign \new_[6716]_  = ~\new_[9151]_  | ~\new_[18280]_ ;
  assign \new_[6717]_  = ~\new_[7577]_ ;
  assign \new_[6718]_  = ~\new_[9155]_  | ~\new_[18621]_ ;
  assign \new_[6719]_  = ~\new_[15322]_  & ~\new_[8852]_ ;
  assign \new_[6720]_  = ~\new_[7584]_ ;
  assign \new_[6721]_  = ~\new_[18468]_  & (~\new_[10684]_  | ~\new_[13341]_ );
  assign \new_[6722]_  = ~\new_[9235]_  | ~\new_[19262]_ ;
  assign \new_[6723]_  = ~\new_[11836]_  | ~\new_[8817]_ ;
  assign \new_[6724]_  = \new_[9239]_  | \new_[19751]_ ;
  assign \new_[6725]_  = \new_[14485]_  & \new_[8899]_ ;
  assign \new_[6726]_  = ~\new_[9164]_  | ~\new_[21510]_ ;
  assign \new_[6727]_  = \new_[9240]_  | \new_[18606]_ ;
  assign \new_[6728]_  = ~\new_[9972]_  & ~\new_[8760]_ ;
  assign \new_[6729]_  = ~\new_[7590]_ ;
  assign \new_[6730]_  = ~\new_[14358]_  | ~\new_[16559]_  | ~\new_[12780]_ ;
  assign \new_[6731]_  = ~\new_[11381]_  | ~\new_[12758]_ ;
  assign \new_[6732]_  = ~\new_[9146]_  | ~\new_[15657]_ ;
  assign \new_[6733]_  = \new_[9241]_  | \new_[19021]_ ;
  assign \new_[6734]_  = ~\new_[11100]_  | ~\new_[11512]_ ;
  assign \new_[6735]_  = ~\new_[13786]_  | ~\new_[12301]_  | ~\new_[10510]_ ;
  assign \new_[6736]_  = ~\new_[9223]_  | ~\new_[10976]_ ;
  assign \new_[6737]_  = ~\new_[11675]_  | ~\new_[12378]_  | ~\new_[10554]_ ;
  assign \new_[6738]_  = ~\new_[10505]_  | ~\new_[12397]_  | ~\new_[10560]_ ;
  assign \new_[6739]_  = \new_[9216]_  | \new_[9961]_ ;
  assign \new_[6740]_  = \new_[8826]_  | \new_[16631]_ ;
  assign \new_[6741]_  = ~\new_[10120]_  & ~\new_[9178]_ ;
  assign \new_[6742]_  = ~\new_[14911]_  | ~\new_[11961]_  | ~\new_[11677]_  | ~\new_[16986]_ ;
  assign \new_[6743]_  = ~\new_[8823]_  & ~\new_[9182]_ ;
  assign \new_[6744]_  = ~\new_[8944]_  & ~\new_[9202]_ ;
  assign \new_[6745]_  = ~\new_[8941]_  | ~\new_[17818]_ ;
  assign \new_[6746]_  = \\dcnt_reg[3] ;
  assign \new_[6747]_  = ~\new_[8762]_  | ~\new_[12624]_ ;
  assign \new_[6748]_  = ~\new_[9064]_  | ~\new_[20341]_ ;
  assign \new_[6749]_  = ~\new_[19233]_  & (~\new_[10656]_  | ~\new_[17343]_ );
  assign \new_[6750]_  = ~\new_[7628]_ ;
  assign \new_[6751]_  = ~\new_[9269]_  & (~\new_[10641]_  | ~\new_[21567]_ );
  assign \new_[6752]_  = \new_[16139]_  & \new_[8928]_ ;
  assign \new_[6753]_  = ~\new_[7631]_ ;
  assign \new_[6754]_  = ~\new_[11506]_  & (~\new_[11882]_  | ~\new_[17051]_ );
  assign \new_[6755]_  = ~\new_[9143]_  | ~\new_[11353]_ ;
  assign \new_[6756]_  = \new_[8844]_  & \new_[19215]_ ;
  assign \new_[6757]_  = \new_[9114]_  & \new_[19206]_ ;
  assign \new_[6758]_  = ~\new_[11329]_  & ~\new_[9181]_ ;
  assign \new_[6759]_  = ~\new_[7637]_ ;
  assign \new_[6760]_  = ~\new_[7638]_ ;
  assign \new_[6761]_  = ~\new_[12674]_  & (~\new_[10715]_  | ~\new_[18982]_ );
  assign \new_[6762]_  = \new_[15291]_  & \new_[8892]_ ;
  assign \new_[6763]_  = ~\new_[7641]_ ;
  assign \new_[6764]_  = ~\new_[17242]_  | ~\new_[17143]_  | ~\new_[12947]_ ;
  assign \new_[6765]_  = ~\new_[11043]_  & (~\new_[14733]_  | ~\new_[19239]_ );
  assign \new_[6766]_  = \new_[8861]_  & \new_[14843]_ ;
  assign \new_[6767]_  = ~\new_[7648]_ ;
  assign \new_[6768]_  = ~\new_[7654]_ ;
  assign \new_[6769]_  = ~\new_[12010]_  | ~\new_[15103]_  | ~\new_[11235]_  | ~\new_[11340]_ ;
  assign \new_[6770]_  = \new_[8841]_  & \new_[18076]_ ;
  assign \new_[6771]_  = ~\new_[8932]_  | ~\new_[19145]_ ;
  assign \new_[6772]_  = ~\new_[8981]_  | ~\new_[11388]_ ;
  assign \new_[6773]_  = ~\new_[10163]_  | ~\new_[11984]_ ;
  assign \new_[6774]_  = ~\new_[9129]_  | ~\new_[9998]_ ;
  assign \new_[6775]_  = \new_[9329]_  | \new_[8781]_ ;
  assign \new_[6776]_  = ~\new_[8936]_  | ~\new_[18967]_ ;
  assign \new_[6777]_  = ~\new_[18572]_  & (~\new_[10627]_  | ~\new_[13366]_ );
  assign \new_[6778]_  = ~\new_[13871]_  | ~\new_[11990]_  | ~\new_[14389]_  | ~\new_[15385]_ ;
  assign \new_[6779]_  = ~\new_[9105]_  | ~\new_[9922]_ ;
  assign \new_[6780]_  = ~\new_[8972]_  | ~\new_[18070]_ ;
  assign \new_[6781]_  = \new_[8975]_  | \new_[19202]_ ;
  assign \new_[6782]_  = ~\new_[9007]_  | ~\new_[17669]_ ;
  assign \new_[6783]_  = ~\new_[9128]_  | ~\new_[21115]_ ;
  assign \new_[6784]_  = ~\new_[7682]_ ;
  assign \new_[6785]_  = ~\new_[9013]_  | ~\new_[9195]_ ;
  assign \new_[6786]_  = ~\new_[12566]_  | ~\new_[14215]_  | ~\new_[10585]_ ;
  assign \new_[6787]_  = ~\new_[8827]_  | ~\new_[15865]_ ;
  assign \new_[6788]_  = ~\new_[10246]_  & ~\new_[9180]_ ;
  assign \new_[6789]_  = ~\new_[8945]_  | ~\new_[12368]_ ;
  assign \new_[6790]_  = ~\new_[944]_  | ~\new_[18818]_  | ~\new_[21390]_ ;
  assign \new_[6791]_  = \new_[8842]_  & \new_[11212]_ ;
  assign \new_[6792]_  = ~\new_[19529]_  & (~\new_[13875]_  | ~\new_[10602]_ );
  assign \new_[6793]_  = ~\new_[8924]_  | ~\new_[21634]_ ;
  assign \new_[6794]_  = ~\new_[9335]_  | ~\new_[9969]_ ;
  assign \new_[6795]_  = ~\new_[9311]_  | ~\new_[9838]_ ;
  assign \new_[6796]_  = ~\new_[9058]_  | ~\new_[21556]_ ;
  assign \new_[6797]_  = ~\new_[7692]_ ;
  assign \new_[6798]_  = ~\new_[7694]_ ;
  assign \new_[6799]_  = ~\new_[13752]_  | ~\new_[11940]_  | ~\new_[11861]_  | ~\new_[15395]_ ;
  assign \new_[6800]_  = \new_[9063]_  & \new_[10077]_ ;
  assign \new_[6801]_  = \new_[9065]_  & \new_[11025]_ ;
  assign \new_[6802]_  = ~\new_[7698]_ ;
  assign \new_[6803]_  = ~\new_[11294]_  & ~\new_[9199]_ ;
  assign \new_[6804]_  = ~\new_[14296]_  | ~\new_[19838]_  | ~\new_[13108]_ ;
  assign \new_[6805]_  = ~\new_[7702]_ ;
  assign \new_[6806]_  = ~\new_[7706]_ ;
  assign \new_[6807]_  = \new_[10394]_  & \new_[9076]_ ;
  assign \new_[6808]_  = ~\new_[13945]_  | ~\new_[8785]_ ;
  assign \new_[6809]_  = ~\new_[7709]_ ;
  assign \new_[6810]_  = ~\new_[11672]_  | ~\new_[8771]_ ;
  assign \new_[6811]_  = ~\new_[9084]_  & ~\new_[9222]_ ;
  assign \new_[6812]_  = \new_[9086]_  & \new_[14926]_ ;
  assign \new_[6813]_  = ~\new_[9088]_  & ~\new_[11445]_ ;
  assign \new_[6814]_  = ~\new_[10310]_  & ~\new_[9214]_ ;
  assign \new_[6815]_  = \new_[9089]_  & \new_[11675]_ ;
  assign \new_[6816]_  = \new_[8894]_  & \new_[15028]_ ;
  assign \new_[6817]_  = ~\new_[17727]_  & (~\new_[10593]_  | ~\new_[12072]_ );
  assign \new_[6818]_  = \new_[8937]_  & \new_[11636]_ ;
  assign \new_[6819]_  = ~\new_[7717]_ ;
  assign \new_[6820]_  = ~\new_[7718]_ ;
  assign \new_[6821]_  = ~\new_[7719]_ ;
  assign \new_[6822]_  = ~\new_[18930]_  & (~\new_[10520]_  | ~\new_[13721]_ );
  assign \new_[6823]_  = ~\new_[9119]_  | ~\new_[9880]_ ;
  assign \new_[6824]_  = ~\new_[10104]_  & ~\new_[9197]_ ;
  assign \new_[6825]_  = ~\new_[7724]_ ;
  assign \new_[6826]_  = ~\new_[7726]_ ;
  assign \new_[6827]_  = ~\new_[19612]_  & (~\new_[10706]_  | ~\new_[15642]_ );
  assign \new_[6828]_  = ~\new_[15899]_  | ~\new_[8753]_  | ~\new_[14102]_ ;
  assign \new_[6829]_  = ~\new_[9148]_  | ~\new_[10896]_ ;
  assign \new_[6830]_  = ~\new_[9157]_  | ~\new_[17845]_ ;
  assign \new_[6831]_  = ~\new_[9171]_  | ~\new_[18288]_ ;
  assign \new_[6832]_  = \new_[9175]_  & \new_[17851]_ ;
  assign \new_[6833]_  = ~\new_[8742]_  | ~\new_[10689]_ ;
  assign \new_[6834]_  = ~\new_[8750]_  | ~\new_[12997]_ ;
  assign \new_[6835]_  = ~\new_[14105]_  | (~\new_[12947]_  & ~\new_[19520]_ );
  assign \new_[6836]_  = ~\new_[9035]_  & ~\new_[11112]_ ;
  assign \new_[6837]_  = \new_[15441]_  ? \new_[20100]_  : \new_[10722]_ ;
  assign \new_[6838]_  = ~\new_[14441]_  & ~\new_[9025]_ ;
  assign \new_[6839]_  = ~\new_[9047]_  & ~\new_[10129]_ ;
  assign \new_[6840]_  = ~\new_[9002]_  & (~\new_[10676]_  | ~\new_[17909]_ );
  assign \new_[6841]_  = ~\new_[9247]_  & (~\new_[17654]_  | ~\new_[15892]_ );
  assign \new_[6842]_  = ~\new_[11668]_  | ~\new_[13969]_  | ~\new_[12917]_  | ~\new_[10515]_ ;
  assign \new_[6843]_  = ~\new_[12678]_  | ~\new_[10325]_  | ~\new_[10573]_ ;
  assign \new_[6844]_  = ~\new_[13852]_  | ~\new_[14842]_  | ~\new_[15097]_  | ~\new_[15246]_ ;
  assign \new_[6845]_  = ~\new_[11582]_  | ~\new_[15661]_  | ~\new_[15175]_  | ~\new_[14995]_ ;
  assign \new_[6846]_  = ~\new_[11598]_  | ~\new_[13846]_  | ~\new_[11897]_  | ~\new_[11612]_ ;
  assign \new_[6847]_  = ~\new_[9154]_  | ~\new_[11928]_ ;
  assign \new_[6848]_  = ~\new_[9003]_  | ~\new_[13228]_ ;
  assign \new_[6849]_  = ~\new_[13954]_  | ~\new_[8782]_ ;
  assign \new_[6850]_  = ~\new_[12170]_  | ~\new_[8784]_ ;
  assign \new_[6851]_  = ~\new_[13356]_  & ~\new_[18361]_  & ~\new_[17552]_ ;
  assign \new_[6852]_  = ~\new_[10737]_  & ~\new_[19072]_  & ~\new_[17786]_ ;
  assign \new_[6853]_  = \new_[7785]_ ;
  assign \new_[6854]_  = ~\new_[7801]_ ;
  assign \new_[6855]_  = ~\new_[9363]_  | ~\new_[20491]_ ;
  assign \new_[6856]_  = ~\new_[7804]_ ;
  assign \new_[6857]_  = ~\new_[11941]_  | ~\new_[18840]_ ;
  assign \new_[6858]_  = ~\new_[9261]_  | ~\new_[14951]_ ;
  assign \new_[6859]_  = ~\new_[9293]_  & ~\new_[21115]_ ;
  assign \new_[6860]_  = ~\new_[7819]_ ;
  assign \new_[6861]_  = ~\new_[9277]_  | ~\new_[16840]_ ;
  assign \new_[6862]_  = ~\new_[11491]_  | ~\new_[9271]_ ;
  assign \new_[6863]_  = \new_[13586]_  | \new_[9309]_ ;
  assign \new_[6864]_  = ~\new_[7830]_ ;
  assign \new_[6865]_  = ~\new_[9260]_  | ~\new_[19547]_ ;
  assign \new_[6866]_  = ~\new_[7836]_ ;
  assign \new_[6867]_  = ~\new_[13053]_  & ~\new_[9344]_ ;
  assign \new_[6868]_  = \new_[12508]_  & \new_[11561]_ ;
  assign \new_[6869]_  = \new_[14029]_  | \new_[9282]_ ;
  assign \new_[6870]_  = \new_[12009]_  | \new_[21635]_ ;
  assign \new_[6871]_  = \new_[9266]_  | \new_[19204]_ ;
  assign \new_[6872]_  = ~\new_[11674]_  | ~\new_[18973]_ ;
  assign \new_[6873]_  = \new_[11266]_  | \new_[18941]_ ;
  assign \new_[6874]_  = ~\new_[11758]_  | ~\new_[18941]_ ;
  assign \new_[6875]_  = ~\new_[7865]_ ;
  assign \new_[6876]_  = ~\new_[16847]_  | ~\new_[10863]_  | ~\new_[14195]_  | ~\new_[11582]_ ;
  assign \new_[6877]_  = ~\new_[11705]_  | ~\new_[19088]_ ;
  assign \new_[6878]_  = ~\new_[7878]_ ;
  assign \new_[6879]_  = ~\new_[9259]_  | ~\new_[18280]_ ;
  assign \new_[6880]_  = \new_[11863]_  | \new_[17381]_ ;
  assign \new_[6881]_  = ~\new_[7890]_ ;
  assign \new_[6882]_  = ~\new_[12831]_  & ~\new_[7119]_ ;
  assign \new_[6883]_  = \new_[12566]_  & \new_[11663]_ ;
  assign \new_[6884]_  = \new_[15049]_  & \new_[13967]_ ;
  assign \new_[6885]_  = \new_[9265]_  | \new_[17689]_ ;
  assign \new_[6886]_  = ~\new_[11584]_  | ~\new_[11507]_ ;
  assign \new_[6887]_  = ~\new_[21112]_ ;
  assign \new_[6888]_  = \new_[16122]_  & \new_[8877]_ ;
  assign \new_[6889]_  = ~\new_[13266]_  & ~\new_[20374]_ ;
  assign \new_[6890]_  = \new_[11762]_  | \new_[19072]_ ;
  assign \new_[6891]_  = \new_[11600]_  | \new_[19215]_ ;
  assign \new_[6892]_  = ~\new_[9312]_  | ~\new_[17472]_ ;
  assign \new_[6893]_  = ~\new_[7906]_ ;
  assign \new_[6894]_  = ~\new_[9281]_  | ~\new_[14593]_ ;
  assign \new_[6895]_  = ~\new_[12690]_  & ~\new_[11689]_ ;
  assign \new_[6896]_  = \new_[11738]_  | \new_[18798]_ ;
  assign \new_[6897]_  = ~\new_[11931]_  | ~\new_[18798]_ ;
  assign \new_[6898]_  = ~\new_[15001]_  | ~\new_[9278]_ ;
  assign \new_[6899]_  = ~\new_[7928]_ ;
  assign \new_[6900]_  = \new_[12466]_  & \new_[9355]_ ;
  assign \new_[6901]_  = ~\new_[12774]_  & ~\new_[11502]_ ;
  assign \new_[6902]_  = ~\new_[11998]_  | ~\new_[21638]_ ;
  assign \new_[6903]_  = ~\new_[9273]_  & ~\new_[21557]_ ;
  assign \new_[6904]_  = ~\new_[12833]_  & ~\new_[9283]_ ;
  assign \new_[6905]_  = ~\new_[10876]_  | ~\new_[10508]_ ;
  assign \new_[6906]_  = ~\new_[9363]_  | ~\new_[16832]_ ;
  assign \new_[6907]_  = ~\new_[19208]_  & ~\new_[9280]_ ;
  assign \new_[6908]_  = ~\new_[12546]_  & ~\new_[11511]_ ;
  assign \new_[6909]_  = ~\new_[11989]_  | ~\new_[20720]_ ;
  assign \new_[6910]_  = ~\new_[9406]_  & (~\new_[10728]_  | ~\new_[18077]_ );
  assign \new_[6911]_  = ~\new_[15571]_  | ~\new_[13996]_ ;
  assign \new_[6912]_  = ~\new_[7974]_ ;
  assign \new_[6913]_  = ~\new_[12216]_  | ~\new_[8568]_  | ~\new_[10745]_ ;
  assign \new_[6914]_  = ~\new_[9378]_  | ~\new_[19567]_ ;
  assign \new_[6915]_  = ~\new_[12982]_  & ~\new_[9336]_ ;
  assign \new_[6916]_  = ~\new_[7992]_ ;
  assign \new_[6917]_  = ~\new_[19208]_  & (~\new_[16369]_  | ~\new_[10737]_ );
  assign \new_[6918]_  = ~\new_[16879]_  & (~\new_[15674]_  | ~\new_[13356]_ );
  assign \new_[6919]_  = ~\new_[18288]_  | (~\new_[10825]_  & ~\new_[10526]_ );
  assign \new_[6920]_  = ~\new_[9366]_  | ~\new_[21556]_ ;
  assign \new_[6921]_  = ~\new_[9364]_  | ~\new_[19711]_ ;
  assign \new_[6922]_  = ~\new_[19233]_  | (~\new_[10821]_  & ~\new_[12597]_ );
  assign \new_[6923]_  = ~\new_[18070]_  | (~\new_[9622]_  & ~\new_[10556]_ );
  assign \new_[6924]_  = ~\new_[10521]_  | ~\new_[12394]_  | ~\new_[11693]_ ;
  assign \new_[6925]_  = ~\new_[11550]_  | ~\new_[9281]_ ;
  assign \new_[6926]_  = ~\new_[19021]_  | (~\new_[10878]_  & ~\new_[13054]_ );
  assign \new_[6927]_  = ~\new_[9264]_  | ~\new_[15321]_ ;
  assign \new_[6928]_  = ~\new_[11613]_  | ~\new_[9356]_ ;
  assign \new_[6929]_  = ~\new_[9267]_  | ~\new_[20463]_ ;
  assign \new_[6930]_  = ~\new_[17583]_  & (~\new_[15894]_  | ~\new_[21651]_ );
  assign \new_[6931]_  = ~\new_[14633]_  | ~\new_[11663]_ ;
  assign \new_[6932]_  = ~\new_[9307]_  | ~\new_[18584]_ ;
  assign \new_[6933]_  = ~\new_[17993]_  & (~\new_[17485]_  | ~\new_[12757]_ );
  assign \new_[6934]_  = ~\new_[20680]_  | (~\new_[9749]_  & ~\new_[13040]_ );
  assign \new_[6935]_  = ~\new_[10513]_  | ~\new_[11703]_  | ~\new_[15738]_ ;
  assign \new_[6936]_  = ~\new_[18124]_  | (~\new_[9744]_  & ~\new_[14203]_ );
  assign \new_[6937]_  = ~\new_[19299]_  | (~\new_[9748]_  & ~\new_[11911]_ );
  assign \new_[6938]_  = ~\new_[9285]_  | ~\new_[14220]_ ;
  assign \new_[6939]_  = \new_[14555]_  | \new_[12862]_ ;
  assign \new_[6940]_  = \new_[13436]_  | \new_[13224]_ ;
  assign \new_[6941]_  = ~\new_[13665]_  & (~\new_[10785]_  | ~\new_[19450]_ );
  assign \new_[6942]_  = ~\new_[13608]_  & (~\new_[10782]_  | ~\new_[18821]_ );
  assign \new_[6943]_  = ~\new_[11825]_  | ~\new_[9293]_ ;
  assign \new_[6944]_  = \new_[13438]_  | \new_[13062]_ ;
  assign \new_[6945]_  = ~\new_[11821]_  | ~\new_[9294]_ ;
  assign \new_[6946]_  = \new_[18921]_  ^ \new_[10736]_ ;
  assign \new_[6947]_  = \new_[18760]_  ^ \new_[10742]_ ;
  assign \new_[6948]_  = ~\new_[11407]_  & (~\new_[9705]_  | ~\new_[19070]_ );
  assign \new_[6949]_  = ~\new_[11408]_  & (~\new_[9762]_  | ~\new_[1928]_ );
  assign \new_[6950]_  = ~\new_[11198]_  & (~\new_[10824]_  | ~\new_[18981]_ );
  assign \new_[6951]_  = ~\new_[12826]_  | ~\new_[14087]_  | ~\new_[11188]_  | ~\new_[12111]_ ;
  assign \new_[6952]_  = ~\new_[19612]_  | (~\new_[10802]_  & ~\new_[11645]_ );
  assign \new_[6953]_  = ~\new_[8026]_ ;
  assign \new_[6954]_  = \new_[9389]_  & \new_[13576]_ ;
  assign \new_[6955]_  = ~\new_[17285]_  | (~\new_[9669]_  & ~\new_[12532]_ );
  assign \new_[6956]_  = ~\new_[19064]_  | (~\new_[10806]_  & ~\new_[12581]_ );
  assign \new_[6957]_  = ~\new_[19717]_  | (~\new_[10859]_  & ~\new_[10113]_ );
  assign \new_[6958]_  = ~\new_[16217]_  | ~\new_[11180]_  | ~\new_[13609]_  | ~\new_[14410]_ ;
  assign \new_[6959]_  = ~\new_[9781]_  & ~\new_[15350]_  & ~\new_[13331]_ ;
  assign \new_[6960]_  = ~\new_[19072]_  | (~\new_[10828]_  & ~\new_[12709]_ );
  assign \new_[6961]_  = ~\new_[17381]_  | (~\new_[9624]_  & ~\new_[12442]_ );
  assign \new_[6962]_  = ~\new_[18795]_  | (~\new_[9627]_  & ~\new_[13828]_ );
  assign \new_[6963]_  = ~\new_[19202]_  | (~\new_[9637]_  & ~\new_[12814]_ );
  assign \new_[6964]_  = ~\new_[17837]_  | (~\new_[9638]_  & ~\new_[12697]_ );
  assign \new_[6965]_  = ~\new_[9371]_  | ~\new_[1080]_ ;
  assign \new_[6966]_  = ~\new_[12866]_  | ~\new_[11309]_  | ~\new_[15253]_  | ~\new_[12088]_ ;
  assign \new_[6967]_  = ~\new_[13238]_  | ~\new_[15328]_  | ~\new_[11314]_  | ~\new_[12056]_ ;
  assign \new_[6968]_  = ~\new_[9652]_  | ~\new_[10884]_  | ~\new_[10922]_ ;
  assign \new_[6969]_  = ~\new_[9778]_  & ~\new_[20967]_  & ~\new_[13330]_ ;
  assign \new_[6970]_  = ~\new_[9779]_  & ~\new_[20905]_  & ~\new_[13392]_ ;
  assign \new_[6971]_  = ~\new_[9780]_  & ~\new_[15228]_  & ~\new_[14411]_ ;
  assign \new_[6972]_  = (~\new_[10800]_  | ~\new_[19088]_ ) & (~\new_[12786]_  | ~\new_[18166]_ );
  assign \new_[6973]_  = (~\new_[10841]_  | ~\new_[19266]_ ) & (~\new_[12511]_  | ~\new_[18008]_ );
  assign \new_[6974]_  = (~\new_[10808]_  | ~\new_[19247]_ ) & (~\new_[12644]_  | ~\new_[18692]_ );
  assign \new_[6975]_  = (~\new_[10812]_  | ~\new_[19288]_ ) & (~\new_[18262]_  | ~\new_[16414]_ );
  assign \new_[6976]_  = ~\new_[9274]_  | ~\new_[9340]_ ;
  assign \new_[6977]_  = ~\new_[9725]_  & (~\new_[10822]_  | ~\new_[18965]_ );
  assign \new_[6978]_  = ~\new_[8656]_  | ~\new_[10726]_ ;
  assign \new_[6979]_  = ~\new_[9394]_  & ~\new_[9931]_ ;
  assign \new_[6980]_  = ~\new_[9395]_  & ~\new_[10943]_ ;
  assign \new_[6981]_  = ~\new_[18789]_  | (~\new_[9752]_  & ~\new_[15273]_ );
  assign \new_[6982]_  = ~\new_[19492]_  | (~\new_[9760]_  & ~\new_[14377]_ );
  assign \new_[6983]_  = ~\new_[9326]_  | ~\new_[20679]_ ;
  assign \new_[6984]_  = ~\new_[9327]_  | (~\new_[12430]_  & ~\new_[19547]_ );
  assign \new_[6985]_  = ~\new_[19320]_  | (~\new_[9766]_  & ~\new_[12911]_ );
  assign \new_[6986]_  = ~\new_[9477]_  & (~\new_[9711]_  | ~\new_[18187]_ );
  assign \new_[6987]_  = ~\new_[9387]_  & ~\new_[10116]_ ;
  assign \new_[6988]_  = ~\new_[10573]_  | ~\new_[8638]_  | ~\new_[10754]_ ;
  assign \new_[6989]_  = ~\new_[9385]_  & ~\new_[10329]_ ;
  assign \new_[6990]_  = ~\new_[9483]_  & (~\new_[9709]_  | ~\new_[19553]_ );
  assign \new_[6991]_  = ~\new_[9328]_  | ~\new_[17796]_ ;
  assign \new_[6992]_  = ~\new_[19798]_  | (~\new_[9737]_  & ~\new_[15288]_ );
  assign \new_[6993]_  = ~\new_[17119]_  | (~\new_[9738]_  & ~\new_[13024]_ );
  assign \new_[6994]_  = ~\new_[20099]_  | (~\new_[9745]_  & ~\new_[12825]_ );
  assign \new_[6995]_  = \\u0_r0_out_reg[29] ;
  assign \new_[6996]_  = ~\new_[8040]_ ;
  assign \new_[6997]_  = ~\new_[17660]_  | (~\new_[9754]_  & ~\new_[15223]_ );
  assign \new_[6998]_  = ~\new_[18827]_  | (~\new_[9770]_  & ~\new_[15152]_ );
  assign \new_[6999]_  = ~\new_[15097]_  | ~\new_[8627]_  | ~\new_[10758]_ ;
  assign \new_[7000]_  = ~\new_[8815]_  & (~\new_[9685]_  | ~\new_[17851]_ );
  assign \new_[7001]_  = ~\new_[9656]_  & ~\new_[9373]_ ;
  assign \new_[7002]_  = ~\new_[11605]_  | ~\new_[12193]_  | ~\new_[10438]_  | ~\new_[11168]_ ;
  assign \new_[7003]_  = ~\new_[10889]_  | ~\new_[14517]_  | ~\new_[14684]_  | ~\new_[12717]_ ;
  assign \new_[7004]_  = ~\new_[9480]_  & (~\new_[9772]_  | ~\new_[2500]_ );
  assign \new_[7005]_  = ~\new_[10960]_  | ~\new_[16495]_  | ~\new_[10685]_  | ~\new_[12627]_ ;
  assign \new_[7006]_  = ~\new_[17061]_  | ~\new_[17057]_  | ~\new_[8726]_  | ~\new_[14531]_ ;
  assign \new_[7007]_  = ~\new_[12215]_  | ~\new_[14565]_  | ~\new_[9339]_  | ~\new_[12612]_ ;
  assign \new_[7008]_  = ~\new_[14504]_  | ~\new_[10926]_  | ~\new_[15365]_  | ~\new_[16546]_ ;
  assign \new_[7009]_  = ~\new_[10998]_  | ~\new_[15640]_  | ~\new_[13276]_  | ~\new_[12785]_ ;
  assign \new_[7010]_  = ~\new_[11127]_  & (~\new_[9699]_  | ~\new_[19350]_ );
  assign \new_[7011]_  = ~\new_[10437]_  | ~\new_[14153]_  | ~\new_[12271]_  | ~\new_[10302]_ ;
  assign \new_[7012]_  = (~\new_[9786]_  | ~\new_[17475]_ ) & (~\new_[14260]_  | ~\new_[18076]_ );
  assign \new_[7013]_  = ~\new_[11116]_  | (~\new_[9751]_  & ~\new_[19249]_ );
  assign \new_[7014]_  = ~\new_[10776]_  & (~\new_[9704]_  | ~\new_[17944]_ );
  assign \new_[7015]_  = ~\new_[9852]_  & (~\new_[9719]_  | ~\new_[18910]_ );
  assign \new_[7016]_  = ~\new_[15181]_  | ~\new_[17785]_  | ~\new_[8727]_  | ~\new_[17616]_ ;
  assign \new_[7017]_  = ~\new_[12118]_  & (~\new_[9728]_  | ~\new_[18597]_ );
  assign \new_[7018]_  = ~\new_[10778]_  & (~\new_[9741]_  | ~\new_[17702]_ );
  assign \new_[7019]_  = ~\new_[10955]_  & ~\new_[9376]_ ;
  assign \new_[7020]_  = ~\new_[13194]_  | ~\new_[10993]_  | ~\new_[13192]_  | ~\new_[14099]_ ;
  assign \new_[7021]_  = ~\new_[9346]_  & (~\new_[9774]_  | ~\new_[19439]_ );
  assign \new_[7022]_  = ~\new_[9310]_  & (~\new_[9707]_  | ~\new_[1879]_ );
  assign \new_[7023]_  = ~\new_[8054]_ ;
  assign \new_[7024]_  = \new_[8694]_  | \new_[19561]_ ;
  assign \new_[7025]_  = ~\new_[8056]_ ;
  assign \new_[7026]_  = ~\new_[18942]_  & (~\new_[10301]_  | ~\new_[10297]_ );
  assign \new_[7027]_  = ~\new_[19436]_  | (~\new_[10296]_  & ~\new_[12847]_ );
  assign \new_[7028]_  = ~\new_[19711]_  | (~\new_[10320]_  & ~\new_[12849]_ );
  assign \new_[7029]_  = ~\new_[21115]_  | (~\new_[10348]_  & ~\new_[12981]_ );
  assign \new_[7030]_  = ~\new_[19261]_  | (~\new_[10382]_  & ~\new_[12970]_ );
  assign \new_[7031]_  = ~\new_[19625]_  | (~\new_[10384]_  & ~\new_[12824]_ );
  assign \new_[7032]_  = ~\new_[19748]_  & (~\new_[13143]_  | ~\new_[9932]_ );
  assign \new_[7033]_  = \new_[8626]_  | \new_[18194]_ ;
  assign \new_[7034]_  = ~\new_[20537]_  & (~\new_[9820]_  | ~\new_[11857]_ );
  assign \new_[7035]_  = ~\new_[19687]_  | (~\new_[10186]_  & ~\new_[13072]_ );
  assign \new_[7036]_  = ~\new_[18652]_  | (~\new_[10355]_  & ~\new_[14193]_ );
  assign \new_[7037]_  = ~\new_[20641]_  & (~\new_[10712]_  | ~\new_[9992]_ );
  assign \new_[7038]_  = ~\new_[19711]_  & (~\new_[10285]_  | ~\new_[12394]_ );
  assign \new_[7039]_  = ~\new_[19064]_  | (~\new_[10026]_  & ~\new_[10450]_ );
  assign \new_[7040]_  = ~\new_[18795]_  | (~\new_[10147]_  & ~\new_[10461]_ );
  assign \new_[7041]_  = ~\new_[19249]_  | (~\new_[10307]_  & ~\new_[10468]_ );
  assign \new_[7042]_  = \new_[9410]_  | \new_[19874]_ ;
  assign \new_[7043]_  = ~\new_[19088]_  | (~\new_[10121]_  & ~\new_[11552]_ );
  assign \new_[7044]_  = ~\new_[19592]_  | (~\new_[10247]_  & ~\new_[13843]_ );
  assign \new_[7045]_  = ~\new_[1081]_  | (~\new_[10506]_  & ~\new_[10381]_ );
  assign \new_[7046]_  = ~\new_[9413]_  | ~\new_[13746]_ ;
  assign \new_[7047]_  = ~\new_[9414]_  | ~\new_[13782]_ ;
  assign \new_[7048]_  = ~\new_[9415]_  | ~\new_[10515]_ ;
  assign \new_[7049]_  = ~\new_[11132]_  & (~\new_[10059]_  | ~\new_[18194]_ );
  assign \new_[7050]_  = ~\new_[8633]_  & ~\new_[14845]_ ;
  assign \new_[7051]_  = ~\new_[9419]_  | ~\new_[13454]_ ;
  assign \new_[7052]_  = ~\new_[9546]_  | ~\new_[19491]_ ;
  assign \new_[7053]_  = \new_[10730]_  ^ \new_[18758]_ ;
  assign \new_[7054]_  = ~\new_[9426]_  | ~\new_[12768]_ ;
  assign \new_[7055]_  = ~\new_[9421]_  | ~\new_[13831]_ ;
  assign \new_[7056]_  = \new_[10731]_  ^ \new_[18851]_ ;
  assign \new_[7057]_  = ~\new_[14648]_  | ~\new_[15751]_  | ~\new_[9897]_ ;
  assign \new_[7058]_  = ~\new_[9422]_  | ~\new_[13868]_ ;
  assign \new_[7059]_  = ~\new_[9797]_  & ~\new_[8665]_ ;
  assign \new_[7060]_  = ~\new_[21638]_  & (~\new_[10124]_  | ~\new_[15407]_ );
  assign \new_[7061]_  = ~\new_[8672]_  | ~\new_[11824]_ ;
  assign \new_[7062]_  = ~\new_[14499]_  | ~\new_[20926]_  | ~\new_[9977]_ ;
  assign \new_[7063]_  = ~\new_[9425]_  | ~\new_[12494]_ ;
  assign \new_[7064]_  = ~\new_[19243]_  | (~\new_[10540]_  & ~\new_[11110]_ );
  assign \new_[7065]_  = ~\new_[9427]_  | ~\new_[11612]_ ;
  assign \new_[7066]_  = ~\new_[18739]_  | (~\new_[10533]_  & ~\new_[20989]_ );
  assign \new_[7067]_  = ~\new_[12092]_  | ~\new_[14857]_  | ~\new_[9867]_ ;
  assign \new_[7068]_  = ~\new_[10128]_  | ~\new_[14198]_  | ~\new_[15723]_ ;
  assign \new_[7069]_  = ~\new_[19751]_  | (~\new_[10058]_  & ~\new_[12745]_ );
  assign \new_[7070]_  = ~\new_[19088]_  | (~\new_[10441]_  & ~\new_[11705]_ );
  assign \new_[7071]_  = \new_[9501]_  & \new_[18209]_ ;
  assign \new_[7072]_  = ~\new_[8555]_  | ~\new_[19085]_ ;
  assign \new_[7073]_  = ~\new_[21328]_  | (~\new_[12332]_  & ~\new_[10702]_ );
  assign \new_[7074]_  = ~\new_[17598]_  | (~\new_[10336]_  & ~\new_[13343]_ );
  assign \new_[7075]_  = ~\new_[18443]_  | (~\new_[12357]_  & ~\new_[10650]_ );
  assign \new_[7076]_  = ~\new_[8605]_  | ~\new_[16840]_ ;
  assign \new_[7077]_  = ~\new_[9469]_  & ~\new_[19860]_ ;
  assign \new_[7078]_  = ~\new_[18821]_  & (~\new_[10583]_  | ~\new_[14883]_ );
  assign \new_[7079]_  = ~\new_[8614]_  | ~\new_[17837]_ ;
  assign \new_[7080]_  = ~\new_[9474]_  | ~\new_[19378]_ ;
  assign \new_[7081]_  = ~\new_[19512]_  | (~\new_[10408]_  & ~\new_[21553]_ );
  assign \new_[7082]_  = ~\new_[9145]_  | ~\new_[19005]_ ;
  assign \new_[7083]_  = ~\new_[14951]_  | (~\new_[10498]_  & ~\new_[14433]_ );
  assign \new_[7084]_  = ~\new_[10030]_  | ~\new_[9468]_ ;
  assign \new_[7085]_  = ~\new_[19445]_  | (~\new_[12448]_  & ~\new_[12853]_ );
  assign \new_[7086]_  = ~\new_[8624]_  & ~\new_[19687]_ ;
  assign \new_[7087]_  = ~\new_[8504]_  | ~\new_[11670]_ ;
  assign \new_[7088]_  = ~\new_[9489]_  | ~\new_[10576]_ ;
  assign \new_[7089]_  = ~\new_[11310]_  & ~\new_[9490]_ ;
  assign \new_[7090]_  = ~\new_[9416]_  | ~\new_[11512]_ ;
  assign \new_[7091]_  = ~\new_[18863]_  | (~\new_[10499]_  & ~\new_[14444]_ );
  assign \new_[7092]_  = ~\new_[11227]_  | ~\new_[9500]_ ;
  assign \new_[7093]_  = ~\new_[10549]_  | ~\new_[12616]_  | ~\new_[10494]_ ;
  assign \new_[7094]_  = ~\new_[15342]_  | ~\new_[14717]_  | ~\new_[9837]_ ;
  assign \new_[7095]_  = ~\new_[11145]_  & ~\new_[9510]_ ;
  assign \new_[7096]_  = ~\new_[8871]_  | ~\new_[9576]_ ;
  assign \new_[7097]_  = ~\new_[9980]_  | ~\new_[11515]_  | ~\new_[10671]_ ;
  assign \new_[7098]_  = ~\new_[8711]_  | ~\new_[9439]_ ;
  assign \new_[7099]_  = ~\new_[19942]_  | ~\new_[12702]_  | ~\new_[12432]_ ;
  assign \new_[7100]_  = ~\new_[9517]_  & ~\new_[20482]_ ;
  assign \new_[7101]_  = ~\new_[9987]_  | ~\new_[12541]_  | ~\new_[12008]_ ;
  assign \new_[7102]_  = ~\new_[9445]_  & (~\new_[10087]_  | ~\new_[18965]_ );
  assign \new_[7103]_  = ~\new_[9524]_  | ~\new_[16169]_ ;
  assign \new_[7104]_  = ~\new_[19553]_  | (~\new_[14488]_  & ~\new_[10074]_ );
  assign \new_[7105]_  = ~\new_[9508]_  | ~\new_[9877]_ ;
  assign \new_[7106]_  = ~\new_[10080]_  | ~\new_[13886]_  | ~\new_[10496]_ ;
  assign \new_[7107]_  = ~\new_[8598]_  | ~\new_[9439]_ ;
  assign \new_[7108]_  = ~\new_[8690]_  | ~\new_[19243]_ ;
  assign \new_[7109]_  = ~\new_[18569]_  & (~\new_[10577]_  | ~\new_[10001]_ );
  assign \new_[7110]_  = ~\new_[9979]_  | ~\new_[13236]_  | ~\new_[13743]_ ;
  assign \new_[7111]_  = ~\new_[8587]_  | ~\new_[15130]_ ;
  assign \new_[7112]_  = ~\new_[10522]_  | ~\new_[11543]_  | ~\new_[10041]_ ;
  assign \new_[7113]_  = ~\new_[15256]_  | ~\new_[15043]_  | ~\new_[9964]_ ;
  assign \new_[7114]_  = ~\new_[10010]_  | ~\new_[8929]_  | ~\new_[14167]_ ;
  assign \new_[7115]_  = ~\new_[19520]_  | (~\new_[9863]_  & ~\new_[15064]_ );
  assign \new_[7116]_  = \new_[8647]_  & \new_[14715]_ ;
  assign \new_[7117]_  = ~\new_[8123]_ ;
  assign \new_[7118]_  = ~\new_[19366]_  | (~\new_[10034]_  & ~\new_[16744]_ );
  assign \new_[7119]_  = ~\new_[10206]_ ;
  assign \new_[7120]_  = ~\new_[18941]_  | ~\new_[960]_  | ~\new_[10406]_ ;
  assign \new_[7121]_  = ~\new_[9459]_  & (~\new_[10174]_  | ~\new_[18998]_ );
  assign \new_[7122]_  = ~\new_[18821]_  & (~\new_[10046]_  | ~\new_[12178]_ );
  assign \new_[7123]_  = ~\new_[8646]_  | ~\new_[19408]_ ;
  assign \new_[7124]_  = ~\new_[10138]_  | ~\new_[16114]_  | ~\new_[10497]_ ;
  assign \new_[7125]_  = \new_[13633]_  | \new_[9565]_ ;
  assign \new_[7126]_  = ~\new_[9496]_  | ~\new_[9982]_ ;
  assign \new_[7127]_  = \new_[12423]_  | \new_[9565]_ ;
  assign \new_[7128]_  = ~\new_[8127]_ ;
  assign \new_[7129]_  = \new_[13554]_  & \new_[9556]_ ;
  assign \new_[7130]_  = ~\new_[10409]_  | ~\new_[11040]_  | ~\new_[11343]_ ;
  assign \new_[7131]_  = ~\new_[8698]_  | ~\new_[12300]_ ;
  assign \new_[7132]_  = ~\new_[19261]_  & (~\new_[10228]_  | ~\new_[12321]_ );
  assign \new_[7133]_  = ~\new_[9411]_  | ~\new_[11684]_ ;
  assign \new_[7134]_  = ~\new_[10447]_  | ~\new_[12224]_  | ~\new_[10350]_ ;
  assign \new_[7135]_  = ~\new_[959]_  | (~\new_[10425]_  & ~\new_[15261]_ );
  assign \new_[7136]_  = ~\new_[11166]_  & ~\new_[9512]_ ;
  assign \new_[7137]_  = ~\new_[19300]_  | (~\new_[12450]_  & ~\new_[10628]_ );
  assign \new_[7138]_  = ~\new_[10112]_  | ~\new_[13909]_  | ~\new_[12478]_ ;
  assign \new_[7139]_  = ~\new_[17689]_  | (~\new_[10500]_  & ~\new_[14446]_ );
  assign \new_[7140]_  = ~\new_[19457]_  | (~\new_[10426]_  & ~\new_[13188]_ );
  assign \new_[7141]_  = ~\new_[19436]_  & (~\new_[11597]_  | ~\new_[9808]_ );
  assign \new_[7142]_  = ~\new_[8961]_  | ~\new_[9587]_ ;
  assign \new_[7143]_  = ~\new_[20100]_  & (~\new_[11604]_  | ~\new_[10197]_ );
  assign \new_[7144]_  = ~\new_[9868]_  | ~\new_[12014]_  | ~\new_[20966]_ ;
  assign \new_[7145]_  = ~\new_[8970]_  & ~\new_[9592]_ ;
  assign \new_[7146]_  = ~\new_[10833]_  & ~\new_[19888]_ ;
  assign \new_[7147]_  = ~\new_[9798]_  | ~\new_[10572]_  | ~\new_[11981]_ ;
  assign \new_[7148]_  = ~\new_[13744]_  | ~\new_[12803]_  | ~\new_[10402]_ ;
  assign \new_[7149]_  = ~\new_[10553]_  | ~\new_[11618]_  | ~\new_[11375]_ ;
  assign \new_[7150]_  = ~\new_[8654]_  & ~\new_[19587]_ ;
  assign \new_[7151]_  = ~\new_[17513]_  | ~\new_[9191]_  | ~\new_[11170]_ ;
  assign \new_[7152]_  = ~\new_[10894]_  | ~\new_[12631]_  | ~\new_[10609]_ ;
  assign \new_[7153]_  = ~\new_[11213]_  & ~\new_[9481]_ ;
  assign \new_[7154]_  = ~\new_[8660]_  | ~\new_[12156]_ ;
  assign \new_[7155]_  = ~\new_[9589]_  | ~\new_[9919]_ ;
  assign \new_[7156]_  = \new_[9617]_  | \new_[10318]_ ;
  assign \new_[7157]_  = \new_[9620]_  & \new_[11605]_ ;
  assign \new_[7158]_  = ~\new_[8492]_  | ~\new_[18855]_ ;
  assign \new_[7159]_  = ~\new_[17668]_  | (~\new_[11640]_  & ~\new_[9925]_ );
  assign \new_[7160]_  = ~\new_[10884]_  | ~\new_[14042]_  | ~\new_[13892]_ ;
  assign \new_[7161]_  = \new_[8498]_  & \new_[17767]_ ;
  assign \new_[7162]_  = ~\new_[8143]_ ;
  assign \new_[7163]_  = ~\new_[18606]_  & (~\new_[10558]_  | ~\new_[9866]_ );
  assign \new_[7164]_  = ~\new_[10757]_  | ~\new_[11714]_ ;
  assign \new_[7165]_  = ~\new_[8670]_  & ~\new_[11190]_ ;
  assign \new_[7166]_  = ~\new_[11510]_  | ~\new_[12779]_  | ~\new_[12168]_ ;
  assign \new_[7167]_  = ~\new_[10157]_  | ~\new_[9052]_  | ~\new_[13509]_ ;
  assign \new_[7168]_  = ~\new_[8147]_ ;
  assign \new_[7169]_  = ~\new_[18077]_  & (~\new_[10535]_  | ~\new_[12238]_ );
  assign \new_[7170]_  = ~\new_[19145]_  & (~\new_[10283]_  | ~\new_[13595]_ );
  assign \new_[7171]_  = ~\new_[21637]_  | (~\new_[11498]_  & ~\new_[9951]_ );
  assign \new_[7172]_  = ~\new_[13114]_  | ~\new_[13818]_  | ~\new_[9915]_ ;
  assign \new_[7173]_  = \new_[9134]_  & \new_[9623]_ ;
  assign \new_[7174]_  = ~\new_[8152]_ ;
  assign \new_[7175]_  = ~\new_[9889]_  | ~\new_[16235]_  | ~\new_[11695]_ ;
  assign \new_[7176]_  = ~\new_[20341]_  & (~\new_[10299]_  | ~\new_[13601]_ );
  assign \new_[7177]_  = ~\new_[8563]_  | ~\new_[954]_ ;
  assign \new_[7178]_  = ~\new_[18077]_  & (~\new_[10314]_  | ~\new_[13587]_ );
  assign \new_[7179]_  = ~\new_[16879]_  & (~\new_[10308]_  | ~\new_[12214]_ );
  assign \new_[7180]_  = ~\new_[17837]_  | ~\new_[18844]_  | ~\new_[12444]_ ;
  assign \new_[7181]_  = ~\new_[19299]_  & (~\new_[10117]_  | ~\new_[14875]_ );
  assign \new_[7182]_  = ~\new_[20432]_  | ~\new_[11431]_  | ~\new_[16128]_ ;
  assign \new_[7183]_  = \new_[13656]_  | \new_[9554]_ ;
  assign \new_[7184]_  = ~\new_[19587]_  & (~\new_[10401]_  | ~\new_[9881]_ );
  assign \new_[7185]_  = ~\new_[8681]_  | ~\new_[12382]_ ;
  assign \new_[7186]_  = \new_[8556]_  & \new_[16670]_ ;
  assign \new_[7187]_  = ~\new_[10304]_  | ~\new_[8553]_ ;
  assign \new_[7188]_  = ~\new_[8682]_  | ~\new_[11261]_ ;
  assign \new_[7189]_  = ~\new_[21562]_  & (~\new_[10191]_  | ~\new_[10236]_ );
  assign \new_[7190]_  = ~\new_[8683]_  | ~\new_[11209]_ ;
  assign \new_[7191]_  = ~\new_[13386]_  | ~\new_[9215]_  | ~\new_[20557]_ ;
  assign \new_[7192]_  = ~\new_[8157]_ ;
  assign \new_[7193]_  = ~\new_[8579]_  & ~\new_[15557]_ ;
  assign \new_[7194]_  = ~\new_[10094]_  & ~\new_[9534]_ ;
  assign \new_[7195]_  = ~\new_[21115]_  & (~\new_[10343]_  | ~\new_[12367]_ );
  assign \new_[7196]_  = \new_[9542]_  | \new_[19717]_ ;
  assign \new_[7197]_  = ~\new_[8572]_  | ~\new_[13698]_ ;
  assign \new_[7198]_  = ~\new_[973]_  | (~\new_[10444]_  & ~\new_[14157]_ );
  assign \new_[7199]_  = ~\new_[8691]_  & ~\new_[19327]_ ;
  assign \new_[7200]_  = ~\new_[8637]_  & ~\new_[18077]_ ;
  assign \new_[7201]_  = ~\new_[8580]_  | ~\new_[19442]_ ;
  assign \new_[7202]_  = \new_[9550]_  & \new_[13952]_ ;
  assign \new_[7203]_  = ~\new_[12895]_  | ~\new_[9144]_  | ~\new_[9984]_ ;
  assign \new_[7204]_  = ~\new_[9573]_  | ~\new_[13530]_ ;
  assign \new_[7205]_  = ~\new_[8593]_  | ~\new_[18643]_ ;
  assign \new_[7206]_  = ~\new_[8163]_ ;
  assign \new_[7207]_  = \new_[8598]_  & \new_[12601]_ ;
  assign \new_[7208]_  = \new_[12438]_  | \new_[9554]_ ;
  assign \new_[7209]_  = ~\new_[946]_  | (~\new_[10440]_  & ~\new_[13148]_ );
  assign \new_[7210]_  = ~\new_[8164]_ ;
  assign \new_[7211]_  = ~\new_[8699]_  & ~\new_[16879]_ ;
  assign \new_[7212]_  = ~\new_[11105]_  & ~\new_[8609]_ ;
  assign \new_[7213]_  = (~\new_[10015]_  | ~\new_[19208]_ ) & (~\new_[17113]_  | ~\new_[15566]_ );
  assign \new_[7214]_  = ~\new_[14946]_  | ~\new_[8729]_  | ~\new_[9822]_ ;
  assign \new_[7215]_  = (~\new_[10063]_  | ~\new_[20704]_ ) & (~\new_[16985]_  | ~\new_[15629]_ );
  assign \new_[7216]_  = ~\new_[12366]_  | ~\new_[12815]_  | ~\new_[10179]_ ;
  assign \new_[7217]_  = ~\new_[9856]_  | ~\new_[8914]_  | ~\new_[11255]_ ;
  assign \new_[7218]_  = ~\new_[11252]_  | ~\new_[13171]_  | ~\new_[10223]_ ;
  assign \new_[7219]_  = ~\new_[12347]_  | ~\new_[21321]_  | ~\new_[10262]_ ;
  assign \new_[7220]_  = ~\new_[10345]_  | ~\new_[13741]_  | ~\new_[11972]_ ;
  assign \new_[7221]_  = ~\new_[10289]_  | ~\new_[13921]_  | ~\new_[10288]_ ;
  assign \new_[7222]_  = ~\new_[14153]_  | ~\new_[14978]_  | ~\new_[9076]_  | ~\new_[12271]_ ;
  assign \new_[7223]_  = ~\new_[9989]_  | ~\new_[9095]_  | ~\new_[10319]_ ;
  assign \new_[7224]_  = ~\new_[9958]_  | ~\new_[9100]_  | ~\new_[11323]_ ;
  assign \new_[7225]_  = ~\new_[8644]_  & (~\new_[17488]_  | ~\new_[17460]_ );
  assign \new_[7226]_  = ~\new_[12343]_  | ~\new_[15133]_  | ~\new_[10393]_ ;
  assign \new_[7227]_  = ~\new_[9828]_  | ~\new_[14147]_  | ~\new_[15138]_ ;
  assign \new_[7228]_  = (~\new_[10069]_  | ~\new_[21056]_ ) & (~\new_[17581]_  | ~\new_[15720]_ );
  assign \new_[7229]_  = ~\new_[10465]_  | ~\new_[10236]_ ;
  assign \new_[7230]_  = ~\new_[8174]_ ;
  assign \new_[7231]_  = ~\new_[12005]_  | ~\new_[14524]_  | ~\new_[9872]_ ;
  assign \new_[7232]_  = \new_[9588]_  | \new_[18778]_ ;
  assign \new_[7233]_  = ~\new_[11953]_  | ~\new_[14831]_  | ~\new_[9921]_ ;
  assign \new_[7234]_  = ~\new_[17089]_  & (~\new_[10471]_  | ~\new_[13717]_ );
  assign \new_[7235]_  = ~\new_[8178]_ ;
  assign \new_[7236]_  = ~\new_[21632]_  | (~\new_[10467]_  & ~\new_[12590]_ );
  assign \new_[7237]_  = ~\new_[8179]_ ;
  assign \new_[7238]_  = ~\new_[8180]_ ;
  assign \new_[7239]_  = ~\new_[8182]_ ;
  assign \new_[7240]_  = \new_[8599]_  | \new_[21056]_ ;
  assign \new_[7241]_  = ~\new_[11326]_  & ~\new_[8728]_ ;
  assign \new_[7242]_  = ~\new_[9465]_  | ~\new_[14060]_ ;
  assign \new_[7243]_  = ~\new_[11872]_  | ~\new_[9577]_ ;
  assign \new_[7244]_  = ~\new_[9472]_  | ~\new_[10014]_ ;
  assign \new_[7245]_  = ~\new_[10657]_  | ~\new_[9475]_ ;
  assign \new_[7246]_  = ~\new_[8889]_  & (~\new_[13608]_  | ~\new_[18288]_ );
  assign \new_[7247]_  = ~\new_[9476]_  | ~\new_[17727]_ ;
  assign \new_[7248]_  = ~\new_[9118]_  & (~\new_[13614]_  | ~\new_[18542]_ );
  assign \new_[7249]_  = ~\new_[11289]_  | ~\new_[11443]_  | ~\new_[11064]_  | ~\new_[13881]_ ;
  assign \new_[7250]_  = ~\new_[8533]_  | ~\new_[14266]_ ;
  assign \new_[7251]_  = ~\new_[19377]_  & (~\new_[10080]_  | ~\new_[15080]_ );
  assign \new_[7252]_  = ~\new_[18898]_  | (~\new_[10335]_  & ~\new_[14477]_ );
  assign \new_[7253]_  = ~\new_[9528]_  & (~\new_[16509]_  | ~\new_[18910]_ );
  assign \new_[7254]_  = ~\new_[8548]_  | ~\new_[19204]_ ;
  assign \new_[7255]_  = ~\new_[8565]_  | ~\new_[19072]_ ;
  assign \new_[7256]_  = ~\new_[9538]_  & (~\new_[15549]_  | ~\new_[18332]_ );
  assign \new_[7257]_  = ~\new_[8569]_  | ~\new_[19711]_ ;
  assign \new_[7258]_  = \new_[9539]_  & \new_[18606]_ ;
  assign \new_[7259]_  = ~\new_[15096]_  & (~\new_[10243]_  | ~\new_[19408]_ );
  assign \new_[7260]_  = ~\new_[9981]_  | ~\new_[14259]_  | ~\new_[13313]_ ;
  assign \new_[7261]_  = ~\new_[17379]_  & (~\new_[10413]_  | ~\new_[10324]_ );
  assign \new_[7262]_  = ~\new_[9570]_  & (~\new_[18402]_  | ~\new_[14478]_ );
  assign \new_[7263]_  = ~\new_[9511]_  | ~\new_[19249]_ ;
  assign \new_[7264]_  = ~\new_[13826]_  | ~\new_[11924]_  | ~\new_[10014]_  | ~\new_[15433]_ ;
  assign \new_[7265]_  = \new_[13005]_  & \new_[9502]_ ;
  assign \new_[7266]_  = ~\new_[8591]_  | ~\new_[15189]_ ;
  assign \new_[7267]_  = ~\new_[9885]_  | ~\new_[8956]_  | ~\new_[12666]_ ;
  assign \new_[7268]_  = ~\new_[9593]_  | ~\new_[11861]_ ;
  assign \new_[7269]_  = ~\new_[9596]_  | ~\new_[10213]_ ;
  assign \new_[7270]_  = ~\new_[8973]_  & (~\new_[13641]_  | ~\new_[20099]_ );
  assign \new_[7271]_  = \new_[9606]_  & \new_[19687]_ ;
  assign \new_[7272]_  = ~\new_[9607]_  | ~\new_[21628]_ ;
  assign \new_[7273]_  = ~\new_[9614]_  | ~\new_[18572]_ ;
  assign \new_[7274]_  = ~\new_[9911]_  | ~\new_[10171]_  | ~\new_[12856]_ ;
  assign \new_[7275]_  = ~\new_[11184]_  | ~\new_[8608]_ ;
  assign \new_[7276]_  = ~\new_[21631]_  & (~\new_[12453]_  | ~\new_[10345]_ );
  assign \new_[7277]_  = ~\new_[8516]_  | ~\new_[17837]_ ;
  assign \new_[7278]_  = ~\new_[10897]_  | ~\new_[14829]_  | ~\new_[10664]_ ;
  assign \new_[7279]_  = ~\new_[9871]_  | ~\new_[14027]_  | ~\new_[12838]_ ;
  assign \new_[7280]_  = ~\new_[13077]_  | ~\new_[11594]_  | ~\new_[11313]_  | ~\new_[11308]_ ;
  assign \new_[7281]_  = ~\new_[12756]_  | ~\new_[12011]_  | ~\new_[10213]_  | ~\new_[14452]_ ;
  assign \new_[7282]_  = ~\new_[13582]_  | ~\new_[14275]_  | ~\new_[10663]_ ;
  assign \new_[7283]_  = ~\new_[9976]_  | ~\new_[21164]_  | ~\new_[10655]_ ;
  assign \new_[7284]_  = ~\new_[12451]_  | ~\new_[11292]_  | ~\new_[11586]_  | ~\new_[13490]_ ;
  assign \new_[7285]_  = ~\new_[8573]_  | ~\new_[19215]_ ;
  assign \new_[7286]_  = ~\new_[19491]_  & (~\new_[12253]_  | ~\new_[9878]_ );
  assign \new_[7287]_  = ~\new_[11945]_  | ~\new_[8576]_ ;
  assign \new_[7288]_  = ~\new_[18537]_  & (~\new_[9875]_  | ~\new_[14142]_ );
  assign \new_[7289]_  = ~\new_[18373]_  & (~\new_[9983]_  | ~\new_[14340]_ );
  assign \new_[7290]_  = ~\new_[17390]_  & (~\new_[12254]_  | ~\new_[14672]_ );
  assign \new_[7291]_  = \new_[9434]_  | \new_[9463]_ ;
  assign \new_[7292]_  = ~\new_[13268]_  | ~\new_[11515]_  | ~\new_[10907]_  | ~\new_[11319]_ ;
  assign \new_[7293]_  = ~\new_[12187]_  | ~\new_[12541]_  | ~\new_[11779]_  | ~\new_[12569]_ ;
  assign \new_[7294]_  = ~\new_[13177]_  | ~\new_[11547]_  | ~\new_[9904]_  | ~\new_[13687]_ ;
  assign \new_[7295]_  = ~\new_[11752]_  | ~\new_[21409]_  | ~\new_[11014]_  | ~\new_[14018]_ ;
  assign \new_[7296]_  = ~\new_[13226]_  | ~\new_[11643]_  | ~\new_[9935]_  | ~\new_[14349]_ ;
  assign \new_[7297]_  = ~\new_[11988]_  | ~\new_[11678]_  | ~\new_[9956]_  | ~\new_[10672]_ ;
  assign \new_[7298]_  = ~\new_[8562]_  | ~\new_[17252]_ ;
  assign \new_[7299]_  = ~\new_[11995]_  | ~\new_[11688]_  | ~\new_[11049]_  | ~\new_[14116]_ ;
  assign \new_[7300]_  = ~\new_[11773]_  | ~\new_[12631]_  | ~\new_[9859]_  | ~\new_[14332]_ ;
  assign \new_[7301]_  = \new_[12632]_  | \new_[9512]_ ;
  assign \new_[7302]_  = ~\new_[9534]_  & (~\new_[14636]_  | ~\new_[18332]_ );
  assign \new_[7303]_  = ~\new_[15340]_  & ~\new_[9515]_ ;
  assign \new_[7304]_  = ~\new_[17121]_  | ~\new_[9524]_ ;
  assign \new_[7305]_  = ~\new_[11002]_  | ~\new_[10217]_  | ~\new_[10212]_ ;
  assign \new_[7306]_  = ~\new_[9553]_  & (~\new_[15749]_  | ~\new_[18402]_ );
  assign \new_[7307]_  = ~\new_[15309]_  | ~\new_[9080]_  | ~\new_[12252]_ ;
  assign \new_[7308]_  = \new_[13885]_  | \new_[9490]_ ;
  assign \new_[7309]_  = ~\new_[10062]_  & (~\new_[10451]_  | ~\new_[19780]_ );
  assign \new_[7310]_  = ~\new_[9505]_  | ~\new_[18522]_ ;
  assign \new_[7311]_  = ~\new_[9438]_  | (~\new_[11187]_  & ~\new_[18414]_ );
  assign \new_[7312]_  = ~\new_[10249]_  & (~\new_[10455]_  | ~\new_[19578]_ );
  assign \new_[7313]_  = (~\new_[10456]_  | ~\new_[19532]_ ) & (~\new_[17193]_  | ~\new_[18849]_ );
  assign \new_[7314]_  = (~\new_[10457]_  | ~\new_[19440]_ ) & (~\new_[17194]_  | ~\new_[19228]_ );
  assign \new_[7315]_  = ~\new_[8903]_  & ~\new_[9401]_ ;
  assign \new_[7316]_  = ~\new_[14179]_  & ~\new_[9575]_ ;
  assign \new_[7317]_  = ~\new_[11278]_  & ~\new_[9405]_ ;
  assign \new_[7318]_  = ~\new_[12961]_  & ~\new_[8564]_ ;
  assign \new_[7319]_  = ~\new_[13310]_  & ~\new_[8574]_ ;
  assign \new_[7320]_  = ~\new_[10617]_  | ~\new_[8848]_  | ~\new_[12301]_ ;
  assign \new_[7321]_  = ~\new_[10925]_  | ~\new_[13667]_  | ~\new_[14062]_  | ~\new_[13642]_ ;
  assign \new_[7322]_  = ~\new_[13620]_  | ~\new_[10920]_  | ~\new_[12486]_  | ~\new_[12338]_ ;
  assign \new_[7323]_  = ~\new_[12503]_  | ~\new_[13936]_  | ~\new_[10112]_  | ~\new_[15347]_ ;
  assign \new_[7324]_  = ~\new_[11700]_  | ~\new_[13758]_  | ~\new_[10138]_  | ~\new_[11732]_ ;
  assign \new_[7325]_  = ~\new_[14961]_  | ~\new_[17061]_  | ~\new_[8915]_  | ~\new_[15544]_ ;
  assign \new_[7326]_  = ~\new_[11599]_  | ~\new_[15343]_  | ~\new_[12397]_  | ~\new_[20713]_ ;
  assign \new_[7327]_  = ~\new_[11620]_  | ~\new_[12800]_  | ~\new_[12369]_  | ~\new_[13644]_ ;
  assign \new_[7328]_  = ~\new_[11783]_  | ~\new_[10312]_  | ~\new_[12378]_ ;
  assign \new_[7329]_  = ~\new_[14379]_  | ~\new_[9093]_  | ~\new_[12394]_ ;
  assign \new_[7330]_  = ~\new_[15311]_  | ~\new_[9139]_  | ~\new_[12287]_ ;
  assign \new_[7331]_  = ~\new_[20085]_  | ~\new_[8918]_  | ~\new_[10445]_ ;
  assign \new_[7332]_  = ~\new_[13803]_  | ~\new_[12128]_  | ~\new_[9830]_ ;
  assign \new_[7333]_  = ~\new_[19405]_  & (~\new_[10490]_  | ~\new_[16266]_ );
  assign \new_[7334]_  = ~\new_[9583]_  & (~\new_[11508]_  | ~\new_[18941]_ );
  assign \new_[7335]_  = ~\new_[12553]_  | ~\new_[9629]_  | ~\new_[9821]_ ;
  assign \new_[7336]_  = ~\new_[11027]_  & ~\new_[8537]_ ;
  assign \new_[7337]_  = \new_[19768]_  ^ \new_[18414]_ ;
  assign \new_[7338]_  = ~\new_[11069]_  | ~\new_[8549]_ ;
  assign \new_[7339]_  = ~\new_[9864]_  | (~\new_[10470]_  & ~\new_[21562]_ );
  assign \new_[7340]_  = ~\new_[9498]_  & (~\new_[16730]_  | ~\new_[15926]_ );
  assign \new_[7341]_  = (~\new_[10013]_  | ~\new_[19377]_ ) & (~\new_[14330]_  | ~\new_[19547]_ );
  assign \new_[7342]_  = (~\new_[10136]_  | ~\new_[2295]_ ) & (~\new_[15279]_  | ~\new_[19366]_ );
  assign \new_[7343]_  = \new_[10368]_  ? \new_[18076]_  : \new_[15325]_ ;
  assign \new_[7344]_  = ~\new_[19102]_  | (~\new_[10704]_  & ~\new_[16470]_ );
  assign \new_[7345]_  = ~\new_[8249]_ ;
  assign \new_[7346]_  = \new_[14709]_  ^ \new_[19507]_ ;
  assign \new_[7347]_  = \new_[19797]_  ^ \new_[19547]_ ;
  assign \new_[7348]_  = ~\new_[9196]_  & ~\new_[19299]_ ;
  assign \new_[7349]_  = ~\new_[8257]_ ;
  assign \new_[7350]_  = \new_[9109]_  & \new_[18542]_ ;
  assign \new_[7351]_  = \new_[8865]_  & \new_[19064]_ ;
  assign \new_[7352]_  = \new_[9124]_  & \new_[19615]_ ;
  assign \new_[7353]_  = ~\new_[8740]_  & ~\new_[19711]_ ;
  assign \new_[7354]_  = ~\new_[8262]_ ;
  assign \new_[7355]_  = ~\new_[8263]_ ;
  assign \new_[7356]_  = ~\new_[8877]_  & ~\new_[19547]_ ;
  assign \new_[7357]_  = ~\new_[8273]_ ;
  assign \new_[7358]_  = \new_[8928]_  | \new_[18833]_ ;
  assign \new_[7359]_  = ~\new_[8280]_ ;
  assign \new_[7360]_  = ~\new_[9193]_  & (~\new_[13914]_  | ~\new_[17939]_ );
  assign \new_[7361]_  = ~\new_[8788]_  & ~\new_[19436]_ ;
  assign \new_[7362]_  = \new_[8746]_  | \new_[18481]_ ;
  assign \new_[7363]_  = ~\new_[8291]_ ;
  assign \new_[7364]_  = ~\new_[8294]_ ;
  assign \new_[7365]_  = \new_[8892]_  | \new_[19239]_ ;
  assign \new_[7366]_  = ~\new_[923]_  & (~\new_[12041]_  | ~\new_[10602]_ );
  assign \new_[7367]_  = ~\new_[9244]_  | ~\new_[19638]_ ;
  assign \new_[7368]_  = ~\new_[8304]_ ;
  assign \new_[7369]_  = ~\new_[8305]_ ;
  assign \new_[7370]_  = ~\new_[8306]_ ;
  assign \new_[7371]_  = ~\new_[21629]_  & (~\new_[15700]_  | ~\new_[13108]_ );
  assign \new_[7372]_  = ~\new_[9245]_  | ~\new_[19148]_ ;
  assign \new_[7373]_  = ~\new_[9250]_  | ~\new_[18599]_ ;
  assign \new_[7374]_  = ~\new_[9252]_  | ~\new_[19378]_ ;
  assign \new_[7375]_  = ~\new_[11074]_  | ~\new_[19711]_ ;
  assign \new_[7376]_  = ~\new_[8887]_  | ~\new_[18187]_ ;
  assign \new_[7377]_  = \new_[10178]_  & \new_[8849]_ ;
  assign \new_[7378]_  = \new_[9228]_  | \new_[19450]_ ;
  assign \new_[7379]_  = ~\new_[8829]_  | ~\new_[13359]_ ;
  assign \new_[7380]_  = \new_[9210]_  | \new_[18481]_ ;
  assign \new_[7381]_  = \new_[9211]_  | \new_[18280]_ ;
  assign \new_[7382]_  = ~\new_[8740]_  | ~\new_[12027]_ ;
  assign \new_[7383]_  = ~\new_[12303]_  | ~\new_[9144]_ ;
  assign \new_[7384]_  = ~\new_[19612]_  & (~\new_[10598]_  | ~\new_[14746]_ );
  assign \new_[7385]_  = \new_[9811]_  & \new_[11663]_ ;
  assign \new_[7386]_  = \new_[9225]_  | \new_[19233]_ ;
  assign \new_[7387]_  = ~\new_[19727]_  | (~\new_[14689]_  & ~\new_[13472]_ );
  assign \new_[7388]_  = ~\new_[8331]_ ;
  assign \new_[7389]_  = ~\new_[8334]_ ;
  assign \new_[7390]_  = ~\new_[8887]_  & ~\new_[12196]_ ;
  assign \new_[7391]_  = ~\new_[17996]_  & (~\new_[10714]_  | ~\new_[12066]_ );
  assign \new_[7392]_  = ~\new_[9022]_  | ~\new_[16875]_ ;
  assign \new_[7393]_  = ~\new_[10898]_  | ~\new_[19088]_ ;
  assign \new_[7394]_  = ~\new_[13856]_  & ~\new_[8743]_ ;
  assign \new_[7395]_  = ~\new_[9230]_  | ~\new_[17727]_ ;
  assign \new_[7396]_  = ~\new_[11077]_  | ~\new_[18280]_ ;
  assign \new_[7397]_  = ~\new_[10910]_  | ~\new_[18194]_ ;
  assign \new_[7398]_  = ~\new_[8353]_ ;
  assign \new_[7399]_  = \new_[10132]_  & \new_[9158]_ ;
  assign \new_[7400]_  = ~\new_[12556]_  | ~\new_[13490]_  | ~\new_[10579]_  | ~\new_[13306]_ ;
  assign \new_[7401]_  = ~\new_[21475]_  | ~\new_[19204]_ ;
  assign \new_[7402]_  = ~\new_[9233]_  | ~\new_[19204]_ ;
  assign \new_[7403]_  = ~\new_[10913]_  | ~\new_[18863]_ ;
  assign \new_[7404]_  = ~\new_[11166]_  & ~\new_[15088]_ ;
  assign \new_[7405]_  = \new_[8874]_  & \new_[17101]_ ;
  assign \new_[7406]_  = \new_[11094]_  | \new_[20680]_ ;
  assign \new_[7407]_  = ~\new_[10537]_  | ~\new_[11727]_  | ~\new_[15708]_ ;
  assign \new_[7408]_  = ~\new_[8876]_  | ~\new_[19687]_ ;
  assign \new_[7409]_  = ~\new_[12359]_  | ~\new_[8749]_ ;
  assign \new_[7410]_  = ~\new_[9231]_  & ~\new_[19145]_ ;
  assign \new_[7411]_  = ~\new_[10027]_  & ~\new_[11102]_ ;
  assign \new_[7412]_  = ~\new_[11300]_  & ~\new_[21056]_ ;
  assign \new_[7413]_  = ~\new_[9986]_  & ~\new_[8748]_ ;
  assign \new_[7414]_  = \new_[9232]_  & \new_[19547]_ ;
  assign \new_[7415]_  = ~\new_[8369]_ ;
  assign \new_[7416]_  = ~\new_[14391]_  | ~\new_[12683]_  | ~\new_[12993]_ ;
  assign \new_[7417]_  = ~\new_[11381]_  | ~\new_[12659]_ ;
  assign \new_[7418]_  = ~\new_[8374]_ ;
  assign \new_[7419]_  = ~\new_[8838]_  | ~\new_[18427]_ ;
  assign \new_[7420]_  = \new_[8888]_  | \new_[19064]_ ;
  assign \new_[7421]_  = \new_[10974]_  & \new_[8740]_ ;
  assign \new_[7422]_  = ~\new_[13280]_  & ~\new_[11055]_ ;
  assign \new_[7423]_  = ~\new_[8401]_ ;
  assign \new_[7424]_  = ~\new_[21594]_  | ~\new_[10590]_  | ~\new_[13311]_ ;
  assign \new_[7425]_  = ~\new_[9156]_  | ~\new_[19079]_ ;
  assign \new_[7426]_  = ~\new_[8921]_  | ~\new_[18414]_ ;
  assign \new_[7427]_  = ~\new_[19115]_  | (~\new_[16613]_  & ~\new_[12533]_ );
  assign \new_[7428]_  = ~\new_[8432]_ ;
  assign \new_[7429]_  = ~\new_[19450]_  | (~\new_[15760]_  & ~\new_[12617]_ );
  assign \new_[7430]_  = ~\new_[20725]_  & (~\new_[10615]_  | ~\new_[12065]_ );
  assign \new_[7431]_  = ~\new_[10138]_  & ~\new_[19288]_ ;
  assign \new_[7432]_  = \new_[9855]_  & \new_[10969]_ ;
  assign \new_[7433]_  = ~\new_[12736]_  | ~\new_[13543]_  | ~\new_[13703]_  | ~\new_[13225]_ ;
  assign \new_[7434]_  = \new_[8948]_  & \new_[11897]_ ;
  assign \new_[7435]_  = ~\new_[20484]_  | ~\new_[21115]_ ;
  assign \new_[7436]_  = ~\new_[13582]_  | ~\new_[8771]_ ;
  assign \new_[7437]_  = ~\new_[11904]_  | ~\new_[8770]_ ;
  assign \new_[7438]_  = ~\new_[9234]_  | ~\new_[17689]_ ;
  assign \new_[7439]_  = ~\new_[10975]_  | ~\new_[17689]_ ;
  assign \new_[7440]_  = ~\new_[8964]_  | ~\new_[18154]_ ;
  assign \new_[7441]_  = ~\new_[10037]_  | ~\new_[11300]_ ;
  assign \new_[7442]_  = ~\new_[8789]_  | ~\new_[10921]_ ;
  assign \new_[7443]_  = ~\new_[8967]_  | ~\new_[18077]_ ;
  assign \new_[7444]_  = ~\new_[12848]_  | ~\new_[8746]_  | ~\new_[14128]_ ;
  assign \new_[7445]_  = \new_[11353]_  | \new_[18124]_ ;
  assign \new_[7446]_  = \new_[8979]_  | \new_[19247]_ ;
  assign \new_[7447]_  = \new_[8980]_  & \new_[13638]_ ;
  assign \new_[7448]_  = ~\new_[20220]_  | ~\new_[14068]_  | ~\new_[15610]_ ;
  assign \new_[7449]_  = ~\new_[8764]_  | ~\new_[14037]_ ;
  assign \new_[7450]_  = ~\new_[11984]_  & ~\new_[18606]_ ;
  assign \new_[7451]_  = ~\new_[8927]_  & ~\new_[19450]_ ;
  assign \new_[7452]_  = ~\new_[8476]_ ;
  assign \new_[7453]_  = ~\new_[20306]_  | ~\new_[8793]_ ;
  assign \new_[7454]_  = ~\new_[9243]_  | ~\new_[21628]_ ;
  assign \new_[7455]_  = ~\new_[8486]_ ;
  assign \new_[7456]_  = ~\new_[9010]_  | ~\new_[12252]_ ;
  assign \new_[7457]_  = ~\new_[12390]_  | ~\new_[11381]_ ;
  assign \new_[7458]_  = \new_[8858]_  & \new_[12241]_ ;
  assign \new_[7459]_  = ~\new_[8927]_  | ~\new_[8835]_ ;
  assign \new_[7460]_  = ~\new_[11991]_  | ~\new_[19951]_  | ~\new_[11999]_ ;
  assign \new_[7461]_  = ~\new_[10088]_  & ~\new_[20725]_ ;
  assign \new_[7462]_  = ~\new_[8493]_ ;
  assign \new_[7463]_  = ~\new_[10140]_  & ~\new_[18412]_ ;
  assign \new_[7464]_  = \new_[10155]_  & \new_[9843]_ ;
  assign \new_[7465]_  = ~\new_[8503]_ ;
  assign \new_[7466]_  = \new_[12189]_  | \new_[9961]_ ;
  assign \new_[7467]_  = ~\new_[9889]_  | ~\new_[15374]_ ;
  assign \new_[7468]_  = ~\new_[8504]_ ;
  assign \new_[7469]_  = ~\new_[9978]_  | ~\new_[11943]_ ;
  assign \new_[7470]_  = ~\new_[13894]_  | ~\new_[15299]_  | ~\new_[11871]_ ;
  assign \new_[7471]_  = ~\new_[9985]_  | ~\new_[10005]_ ;
  assign \new_[7472]_  = ~\new_[9849]_  & ~\new_[12711]_ ;
  assign \new_[7473]_  = ~\new_[10248]_  & ~\new_[9928]_ ;
  assign \new_[7474]_  = \new_[10446]_  & \new_[21634]_ ;
  assign \new_[7475]_  = ~\new_[10370]_  & ~\new_[12315]_ ;
  assign \new_[7476]_  = \new_[10433]_  | \new_[18795]_ ;
  assign \new_[7477]_  = ~\new_[20660]_  | ~\new_[11087]_ ;
  assign \new_[7478]_  = ~\new_[19170]_  | (~\new_[14898]_  & ~\new_[11906]_ );
  assign \new_[7479]_  = ~\new_[11020]_  & ~\new_[9974]_ ;
  assign \new_[7480]_  = ~\new_[10252]_  | ~\new_[18752]_ ;
  assign \new_[7481]_  = ~\new_[10214]_  | ~\new_[21562]_ ;
  assign \new_[7482]_  = ~\new_[9869]_  | ~\new_[13724]_ ;
  assign \new_[7483]_  = ~\new_[8513]_ ;
  assign \new_[7484]_  = ~\new_[12378]_  | ~\new_[11657]_ ;
  assign \new_[7485]_  = ~\new_[10386]_  | ~\new_[18124]_ ;
  assign \new_[7486]_  = ~\new_[10326]_  | ~\new_[21636]_ ;
  assign \new_[7487]_  = ~\new_[10220]_  | ~\new_[17067]_ ;
  assign \new_[7488]_  = ~\new_[8519]_ ;
  assign \new_[7489]_  = ~\new_[10434]_  | ~\new_[12657]_ ;
  assign \new_[7490]_  = ~\new_[12727]_  | ~\new_[10232]_ ;
  assign \new_[7491]_  = ~\new_[12406]_  | ~\new_[15201]_ ;
  assign \new_[7492]_  = ~\new_[12213]_  | ~\new_[10021]_ ;
  assign \new_[7493]_  = ~\new_[10236]_  | ~\new_[11536]_ ;
  assign \new_[7494]_  = ~\new_[9944]_  | ~\new_[11919]_ ;
  assign \new_[7495]_  = ~\new_[10077]_  | ~\new_[12265]_ ;
  assign \new_[7496]_  = ~\new_[19299]_  & (~\new_[16924]_  | ~\new_[11783]_ );
  assign \new_[7497]_  = ~\new_[10334]_  & ~\new_[11387]_ ;
  assign \new_[7498]_  = \new_[12266]_  & \new_[9923]_ ;
  assign \new_[7499]_  = \new_[10215]_  | \new_[17244]_ ;
  assign \new_[7500]_  = ~\new_[9899]_  & ~\new_[13593]_ ;
  assign \new_[7501]_  = \new_[10466]_  | \new_[19145]_ ;
  assign \new_[7502]_  = ~\new_[20989]_  & ~\new_[15022]_ ;
  assign \new_[7503]_  = ~\new_[12247]_  | ~\new_[10708]_ ;
  assign \new_[7504]_  = ~\new_[20306]_  | ~\new_[12183]_ ;
  assign \new_[7505]_  = ~\new_[12417]_  & ~\new_[12444]_ ;
  assign \new_[7506]_  = ~\new_[19021]_  & (~\new_[11823]_  | ~\new_[16051]_ );
  assign \new_[7507]_  = ~\new_[10154]_  & ~\new_[10020]_ ;
  assign \new_[7508]_  = ~\new_[10225]_  & ~\new_[20622]_ ;
  assign \new_[7509]_  = ~\new_[12379]_  | ~\new_[10200]_ ;
  assign \new_[7510]_  = ~\new_[9953]_  | ~\new_[10509]_ ;
  assign \new_[7511]_  = ~\new_[14073]_  & ~\new_[9947]_ ;
  assign \new_[7512]_  = ~\new_[10295]_  | ~\new_[11666]_ ;
  assign \new_[7513]_  = \new_[10220]_  | \new_[17335]_ ;
  assign \new_[7514]_  = ~\new_[8544]_ ;
  assign \new_[7515]_  = ~\new_[9853]_  | ~\new_[12925]_ ;
  assign \new_[7516]_  = ~\new_[12263]_  & ~\new_[12392]_ ;
  assign \new_[7517]_  = \new_[10232]_  | \new_[21628]_ ;
  assign \new_[7518]_  = ~\new_[9959]_  | ~\new_[13046]_ ;
  assign \new_[7519]_  = ~\new_[18795]_  | (~\new_[13733]_  & ~\new_[14326]_ );
  assign \new_[7520]_  = ~\new_[10124]_  & ~\new_[21274]_ ;
  assign \new_[7521]_  = ~\new_[12406]_  | ~\new_[11955]_ ;
  assign \new_[7522]_  = ~\new_[12032]_  | ~\new_[10237]_ ;
  assign \new_[7523]_  = ~\new_[20221]_  | ~\new_[10604]_  | ~\new_[13089]_ ;
  assign \new_[7524]_  = \new_[10885]_  & \new_[21146]_ ;
  assign \new_[7525]_  = ~\new_[10245]_  | ~\new_[18361]_ ;
  assign \new_[7526]_  = ~\new_[11025]_  | ~\new_[10667]_ ;
  assign \new_[7527]_  = ~\new_[21638]_  & (~\new_[11534]_  | ~\new_[16229]_ );
  assign \new_[7528]_  = ~\new_[19266]_  & (~\new_[11549]_  | ~\new_[14052]_ );
  assign \new_[7529]_  = \new_[10311]_  & \new_[19357]_ ;
  assign \new_[7530]_  = \new_[12367]_  & \new_[12526]_ ;
  assign \new_[7531]_  = ~\new_[8553]_ ;
  assign \new_[7532]_  = ~\new_[16449]_  | ~\new_[10207]_ ;
  assign \new_[7533]_  = ~\new_[14243]_  | ~\new_[9923]_  | ~\new_[14316]_ ;
  assign \new_[7534]_  = \new_[12294]_  | \new_[19625]_ ;
  assign \new_[7535]_  = ~\new_[10189]_  | ~\new_[19059]_ ;
  assign \new_[7536]_  = ~\new_[10591]_  | ~\new_[11207]_ ;
  assign \new_[7537]_  = ~\new_[18292]_  & (~\new_[12000]_  | ~\new_[12068]_ );
  assign \new_[7538]_  = ~\new_[10884]_  | ~\new_[15312]_ ;
  assign \new_[7539]_  = ~\new_[9993]_  | ~\new_[12870]_ ;
  assign \new_[7540]_  = ~\new_[11573]_  | ~\new_[11841]_  | ~\new_[14784]_ ;
  assign \new_[7541]_  = ~\new_[10337]_  | ~\new_[19450]_ ;
  assign \new_[7542]_  = \new_[12321]_  | \new_[18967]_ ;
  assign \new_[7543]_  = \new_[11047]_  & \new_[9875]_ ;
  assign \new_[7544]_  = ~\new_[12399]_  | ~\new_[10402]_ ;
  assign \new_[7545]_  = ~\new_[10344]_  | ~\new_[21115]_ ;
  assign \new_[7546]_  = ~\new_[13914]_  & ~\new_[9884]_ ;
  assign \new_[7547]_  = ~\new_[9958]_  | ~\new_[14294]_ ;
  assign \new_[7548]_  = \new_[15347]_  & \new_[9990]_ ;
  assign \new_[7549]_  = ~\new_[10379]_  | ~\new_[19064]_ ;
  assign \new_[7550]_  = ~\new_[11948]_  | ~\new_[21195]_  | ~\new_[11756]_ ;
  assign \new_[7551]_  = ~\new_[16269]_  & ~\new_[10083]_ ;
  assign \new_[7552]_  = \new_[10474]_  | \new_[19441]_ ;
  assign \new_[7553]_  = ~\new_[18473]_  & (~\new_[11970]_  | ~\new_[14425]_ );
  assign \new_[7554]_  = ~\new_[11150]_  | ~\new_[9868]_ ;
  assign \new_[7555]_  = ~\new_[19064]_  | (~\new_[13697]_  & ~\new_[14154]_ );
  assign \new_[7556]_  = \new_[9846]_  & \new_[12443]_ ;
  assign \new_[7557]_  = \new_[10486]_  | \new_[21056]_ ;
  assign \new_[7558]_  = ~\new_[9824]_  | ~\new_[17475]_ ;
  assign \new_[7559]_  = ~\new_[10357]_  | ~\new_[11067]_ ;
  assign \new_[7560]_  = ~\new_[12432]_  | ~\new_[11671]_ ;
  assign \new_[7561]_  = ~\new_[11544]_  | ~\new_[13688]_  | ~\new_[16657]_ ;
  assign \new_[7562]_  = ~\new_[21251]_  & ~\new_[13016]_ ;
  assign \new_[7563]_  = ~\new_[9822]_  | ~\new_[13560]_ ;
  assign \new_[7564]_  = ~\new_[20940]_  | ~\new_[20938]_ ;
  assign \new_[7565]_  = ~\new_[10362]_  | ~\new_[19587]_ ;
  assign \new_[7566]_  = ~\new_[12295]_  | ~\new_[15638]_ ;
  assign \new_[7567]_  = ~\new_[10364]_  | ~\new_[9979]_ ;
  assign \new_[7568]_  = \new_[9981]_  | \new_[19079]_ ;
  assign \new_[7569]_  = \new_[10118]_  | \new_[18124]_ ;
  assign \new_[7570]_  = ~\new_[18786]_  | (~\new_[10864]_  & ~\new_[16317]_ );
  assign \new_[7571]_  = ~\new_[9832]_  | ~\new_[10920]_ ;
  assign \new_[7572]_  = \new_[10479]_  | \new_[19088]_ ;
  assign \new_[7573]_  = ~\new_[10057]_  & ~\new_[14039]_ ;
  assign \new_[7574]_  = ~\new_[10192]_  | ~\new_[11087]_ ;
  assign \new_[7575]_  = ~\new_[8582]_ ;
  assign \new_[7576]_  = ~\new_[9984]_  | ~\new_[12895]_ ;
  assign \new_[7577]_  = ~\new_[9965]_  | ~\new_[13689]_ ;
  assign \new_[7578]_  = ~\new_[18412]_  & (~\new_[13279]_  | ~\new_[12071]_ );
  assign \new_[7579]_  = ~\new_[9817]_  | ~\new_[14016]_ ;
  assign \new_[7580]_  = \new_[9911]_  | \new_[19072]_ ;
  assign \new_[7581]_  = ~\new_[10381]_  & ~\new_[13976]_ ;
  assign \new_[7582]_  = ~\new_[13702]_  & ~\new_[9825]_ ;
  assign \new_[7583]_  = ~\new_[9991]_  | ~\new_[14067]_ ;
  assign \new_[7584]_  = ~\new_[10051]_  | ~\new_[18967]_ ;
  assign \new_[7585]_  = ~\new_[10481]_  | ~\new_[19233]_ ;
  assign \new_[7586]_  = ~\new_[13604]_  | ~\new_[9997]_ ;
  assign \new_[7587]_  = ~\new_[8598]_ ;
  assign \new_[7588]_  = ~\new_[10402]_  | ~\new_[11718]_ ;
  assign \new_[7589]_  = ~\new_[10000]_  | ~\new_[13080]_ ;
  assign \new_[7590]_  = ~\new_[10391]_  | ~\new_[19079]_ ;
  assign \new_[7591]_  = ~\new_[11378]_  & ~\new_[12155]_ ;
  assign \new_[7592]_  = ~\new_[9981]_  | ~\new_[10001]_ ;
  assign \new_[7593]_  = ~\new_[12043]_  | ~\new_[9999]_ ;
  assign \new_[7594]_  = ~\new_[10397]_  | ~\new_[10965]_ ;
  assign \new_[7595]_  = ~\new_[10004]_  | ~\new_[14381]_ ;
  assign \new_[7596]_  = ~\new_[10005]_  | ~\new_[15592]_ ;
  assign \new_[7597]_  = ~\new_[12221]_  | ~\new_[10638]_ ;
  assign \new_[7598]_  = ~\new_[10006]_  | ~\new_[11569]_ ;
  assign \new_[7599]_  = ~\new_[8610]_ ;
  assign \new_[7600]_  = ~\new_[20703]_  | ~\new_[16879]_ ;
  assign \new_[7601]_  = ~\new_[10884]_  | ~\new_[12822]_ ;
  assign \new_[7602]_  = ~\new_[10029]_  | ~\new_[19711]_ ;
  assign \new_[7603]_  = ~\new_[11800]_  | ~\new_[21674]_  | ~\new_[15918]_ ;
  assign \new_[7604]_  = ~\new_[10065]_  & ~\new_[11526]_ ;
  assign \new_[7605]_  = \new_[10453]_  & \new_[10080]_ ;
  assign \new_[7606]_  = \new_[11432]_  & \new_[10112]_ ;
  assign \new_[7607]_  = \new_[10459]_  & \new_[10138]_ ;
  assign \new_[7608]_  = ~\new_[8617]_ ;
  assign \new_[7609]_  = ~\new_[21408]_  | ~\new_[10227]_  | ~\new_[11629]_ ;
  assign \new_[7610]_  = ~\new_[10102]_  & ~\new_[12649]_ ;
  assign \new_[7611]_  = ~\new_[10274]_  | (~\new_[18890]_  & ~\new_[19156]_ );
  assign \new_[7612]_  = \new_[11437]_  & \new_[10549]_ ;
  assign \new_[7613]_  = ~\new_[11830]_  | ~\new_[12810]_  | ~\new_[14732]_ ;
  assign \new_[7614]_  = ~\new_[16409]_  | ~\new_[16127]_  | ~\new_[14259]_ ;
  assign \new_[7615]_  = ~\new_[10092]_  | (~\new_[19263]_  & ~\new_[19203]_ );
  assign \new_[7616]_  = ~\new_[14063]_  | ~\new_[15104]_  | ~\new_[14993]_ ;
  assign \new_[7617]_  = ~\new_[19177]_  & (~\new_[15593]_  | ~\new_[13739]_ );
  assign \new_[7618]_  = ~\new_[10053]_  & (~\new_[14802]_  | ~\new_[18402]_ );
  assign \new_[7619]_  = ~\new_[19088]_  & (~\new_[11756]_  | ~\new_[15020]_ );
  assign \new_[7620]_  = ~\new_[10192]_  | (~\new_[16630]_  & ~\new_[21697]_ );
  assign \new_[7621]_  = ~\new_[8630]_ ;
  assign \new_[7622]_  = \new_[10160]_  | \new_[18194]_ ;
  assign \new_[7623]_  = ~\new_[11847]_  | ~\new_[15057]_  | ~\new_[16121]_ ;
  assign \new_[7624]_  = ~\new_[19377]_  & (~\new_[15730]_  | ~\new_[13927]_ );
  assign \new_[7625]_  = \new_[10143]_  & \new_[19079]_ ;
  assign \new_[7626]_  = ~\new_[10511]_  & (~\new_[11868]_  | ~\new_[20169]_ );
  assign \new_[7627]_  = ~\new_[10526]_  & (~\new_[11765]_  | ~\new_[18199]_ );
  assign \new_[7628]_  = \new_[10333]_  & \new_[18124]_ ;
  assign \new_[7629]_  = ~\new_[10116]_  & (~\new_[18332]_  | ~\new_[17860]_ );
  assign \new_[7630]_  = ~\new_[9816]_  | ~\new_[16556]_ ;
  assign \new_[7631]_  = \new_[10100]_  & \new_[18965]_ ;
  assign \new_[7632]_  = ~\new_[10153]_  | ~\new_[10419]_ ;
  assign \new_[7633]_  = ~\new_[10398]_  | ~\new_[19088]_ ;
  assign \new_[7634]_  = ~\new_[10083]_  & (~\new_[17734]_  | ~\new_[15536]_ );
  assign \new_[7635]_  = ~\new_[11513]_  | ~\new_[13693]_  | ~\new_[13073]_ ;
  assign \new_[7636]_  = ~\new_[14184]_  | ~\new_[15036]_  | ~\new_[13798]_ ;
  assign \new_[7637]_  = \new_[10035]_  & \new_[20680]_ ;
  assign \new_[7638]_  = ~\new_[19215]_  & (~\new_[13684]_  | ~\new_[12085]_ );
  assign \new_[7639]_  = \new_[10114]_  & \new_[10172]_ ;
  assign \new_[7640]_  = ~\new_[10166]_  & ~\new_[12932]_ ;
  assign \new_[7641]_  = ~\new_[18569]_  & (~\new_[16326]_  | ~\new_[13961]_ );
  assign \new_[7642]_  = ~\new_[13538]_  | ~\new_[16858]_  | ~\new_[14229]_ ;
  assign \new_[7643]_  = ~\new_[13839]_  | ~\new_[10000]_ ;
  assign \new_[7644]_  = \new_[10103]_  | \new_[19021]_ ;
  assign \new_[7645]_  = ~\new_[12575]_  | ~\new_[9817]_ ;
  assign \new_[7646]_  = \new_[10331]_  | \new_[10901]_ ;
  assign \new_[7647]_  = ~\new_[12606]_  | ~\new_[14345]_  | ~\new_[13615]_  | ~\new_[12868]_ ;
  assign \new_[7648]_  = ~\new_[12513]_  | (~\new_[13685]_  & ~\new_[19224]_ );
  assign \new_[7649]_  = ~\new_[10137]_  | ~\new_[19625]_ ;
  assign \new_[7650]_  = \new_[10169]_  | \new_[19547]_ ;
  assign \new_[7651]_  = ~\new_[8645]_ ;
  assign \new_[7652]_  = ~\new_[10090]_  | ~\new_[14852]_ ;
  assign \new_[7653]_  = ~\new_[10329]_  & (~\new_[18910]_  | ~\new_[17208]_ );
  assign \new_[7654]_  = ~\new_[19088]_  & (~\new_[14920]_  | ~\new_[11523]_ );
  assign \new_[7655]_  = ~\new_[10631]_  | ~\new_[12185]_ ;
  assign \new_[7656]_  = ~\new_[13173]_  | ~\new_[12789]_  | ~\new_[13717]_ ;
  assign \new_[7657]_  = \new_[10045]_  | \new_[14951]_ ;
  assign \new_[7658]_  = ~\new_[13955]_  | ~\new_[9991]_ ;
  assign \new_[7659]_  = \new_[10091]_  | \new_[21115]_ ;
  assign \new_[7660]_  = ~\new_[18984]_  & (~\new_[15123]_  | ~\new_[11561]_ );
  assign \new_[7661]_  = ~\new_[10168]_  | ~\new_[17225]_ ;
  assign \new_[7662]_  = \new_[10373]_  | \new_[9814]_ ;
  assign \new_[7663]_  = ~\new_[12293]_  | (~\new_[17172]_  & ~\new_[19018]_ );
  assign \new_[7664]_  = ~\new_[11493]_  | ~\new_[14247]_  | ~\new_[13068]_ ;
  assign \new_[7665]_  = ~\new_[10181]_  | (~\new_[17970]_  & ~\new_[18605]_ );
  assign \new_[7666]_  = \new_[10229]_  & \new_[10257]_ ;
  assign \new_[7667]_  = ~\new_[10600]_  | ~\new_[20712]_ ;
  assign \new_[7668]_  = ~\new_[18361]_  & (~\new_[11854]_  | ~\new_[16336]_ );
  assign \new_[7669]_  = ~\new_[11683]_  | ~\new_[15335]_  | ~\new_[12159]_ ;
  assign \new_[7670]_  = ~\new_[10119]_  | (~\new_[17108]_  & ~\new_[18938]_ );
  assign \new_[7671]_  = ~\new_[12597]_  & (~\new_[11916]_  | ~\new_[19136]_ );
  assign \new_[7672]_  = ~\new_[11608]_  | ~\new_[13846]_  | ~\new_[14622]_ ;
  assign \new_[7673]_  = \new_[10209]_  & \new_[18627]_ ;
  assign \new_[7674]_  = \new_[10210]_  & \new_[10212]_ ;
  assign \new_[7675]_  = \new_[10211]_  | \new_[21562]_ ;
  assign \new_[7676]_  = ~\new_[16660]_  | ~\new_[21680]_  | ~\new_[14714]_ ;
  assign \new_[7677]_  = \new_[10218]_  & \new_[19450]_ ;
  assign \new_[7678]_  = ~\new_[12790]_  & (~\new_[13102]_  | ~\new_[19180]_ );
  assign \new_[7679]_  = ~\new_[10184]_  | (~\new_[15831]_  & ~\new_[18325]_ );
  assign \new_[7680]_  = ~\new_[10557]_  & (~\new_[12172]_  | ~\new_[17135]_ );
  assign \new_[7681]_  = ~\new_[8662]_ ;
  assign \new_[7682]_  = ~\new_[19071]_  & (~\new_[15385]_  | ~\new_[13825]_ );
  assign \new_[7683]_  = ~\new_[10238]_  | ~\new_[18798]_ ;
  assign \new_[7684]_  = ~\new_[11679]_  | ~\new_[13610]_  | ~\new_[13204]_ ;
  assign \new_[7685]_  = ~\new_[8666]_ ;
  assign \new_[7686]_  = ~\new_[10237]_  | (~\new_[15636]_  & ~\new_[19275]_ );
  assign \new_[7687]_  = ~\new_[11276]_  & ~\new_[10432]_ ;
  assign \new_[7688]_  = ~\new_[10251]_  | ~\new_[11281]_ ;
  assign \new_[7689]_  = ~\new_[16084]_  | ~\new_[16802]_  | ~\new_[14027]_ ;
  assign \new_[7690]_  = ~\new_[10260]_  & ~\new_[13186]_ ;
  assign \new_[7691]_  = ~\new_[11650]_  | ~\new_[12980]_  | ~\new_[11989]_ ;
  assign \new_[7692]_  = ~\new_[18046]_  & (~\new_[16277]_  | ~\new_[11542]_ );
  assign \new_[7693]_  = ~\new_[10271]_  | ~\new_[14454]_ ;
  assign \new_[7694]_  = ~\new_[19145]_  & (~\new_[11809]_  | ~\new_[15447]_ );
  assign \new_[7695]_  = ~\new_[13913]_  | ~\new_[9959]_ ;
  assign \new_[7696]_  = ~\new_[10713]_  | ~\new_[20160]_ ;
  assign \new_[7697]_  = \new_[10086]_  & \new_[19687]_ ;
  assign \new_[7698]_  = ~\new_[19266]_  & (~\new_[14662]_  | ~\new_[11609]_ );
  assign \new_[7699]_  = ~\new_[8674]_ ;
  assign \new_[7700]_  = ~\new_[11969]_  | ~\new_[9853]_ ;
  assign \new_[7701]_  = ~\new_[11647]_  | ~\new_[9993]_ ;
  assign \new_[7702]_  = ~\new_[15383]_  | (~\new_[12095]_  & ~\new_[17979]_ );
  assign \new_[7703]_  = ~\new_[10539]_  | ~\new_[9939]_ ;
  assign \new_[7704]_  = ~\new_[10686]_  | ~\new_[9917]_ ;
  assign \new_[7705]_  = ~\new_[10556]_  & (~\new_[12087]_  | ~\new_[19014]_ );
  assign \new_[7706]_  = ~\new_[18077]_  & (~\new_[14443]_  | ~\new_[13681]_ );
  assign \new_[7707]_  = ~\new_[10293]_  | ~\new_[18847]_ ;
  assign \new_[7708]_  = ~\new_[8678]_ ;
  assign \new_[7709]_  = ~\new_[13977]_  | (~\new_[14305]_  & ~\new_[21328]_ );
  assign \new_[7710]_  = ~\new_[10619]_  | ~\new_[9944]_ ;
  assign \new_[7711]_  = \new_[10313]_  & \new_[10521]_ ;
  assign \new_[7712]_  = ~\new_[21558]_  & (~\new_[11555]_  | ~\new_[15600]_ );
  assign \new_[7713]_  = ~\new_[10317]_  | ~\new_[12182]_ ;
  assign \new_[7714]_  = ~\new_[13901]_  | ~\new_[9851]_ ;
  assign \new_[7715]_  = ~\new_[18803]_  & (~\new_[12593]_  | ~\new_[11797]_ );
  assign \new_[7716]_  = ~\new_[13812]_  | ~\new_[9952]_ ;
  assign \new_[7717]_  = ~\new_[18863]_  & (~\new_[11494]_  | ~\new_[21300]_ );
  assign \new_[7718]_  = ~\new_[14951]_  & (~\new_[14545]_  | ~\new_[12074]_ );
  assign \new_[7719]_  = ~\new_[18280]_  & (~\new_[15398]_  | ~\new_[13717]_ );
  assign \new_[7720]_  = ~\new_[19687]_  & (~\new_[12014]_  | ~\new_[15462]_ );
  assign \new_[7721]_  = ~\new_[8685]_ ;
  assign \new_[7722]_  = ~\new_[8687]_ ;
  assign \new_[7723]_  = ~\new_[19266]_  & (~\new_[11999]_  | ~\new_[16307]_ );
  assign \new_[7724]_  = \new_[10421]_  & \new_[19145]_ ;
  assign \new_[7725]_  = ~\new_[18731]_  & (~\new_[11598]_  | ~\new_[13943]_ );
  assign \new_[7726]_  = ~\new_[21115]_  & (~\new_[12016]_  | ~\new_[13347]_ );
  assign \new_[7727]_  = \new_[10208]_  & \new_[19612]_ ;
  assign \new_[7728]_  = ~\new_[19141]_  & (~\new_[11668]_  | ~\new_[13973]_ );
  assign \new_[7729]_  = ~\new_[10351]_  & ~\new_[10528]_ ;
  assign \new_[7730]_  = ~\new_[10021]_  | (~\new_[16553]_  & ~\new_[21166]_ );
  assign \new_[7731]_  = ~\new_[11709]_  | ~\new_[14664]_  | ~\new_[15729]_ ;
  assign \new_[7732]_  = ~\new_[11801]_  | ~\new_[9969]_ ;
  assign \new_[7733]_  = ~\new_[14334]_  | ~\new_[9875]_ ;
  assign \new_[7734]_  = ~\new_[18132]_  & (~\new_[12924]_  | ~\new_[14457]_ );
  assign \new_[7735]_  = ~\new_[13100]_  | ~\new_[9944]_ ;
  assign \new_[7736]_  = ~\new_[11748]_  | ~\new_[9917]_ ;
  assign \new_[7737]_  = ~\new_[11965]_  | ~\new_[9838]_ ;
  assign \new_[7738]_  = ~\new_[12038]_  | ~\new_[9999]_ ;
  assign \new_[7739]_  = ~\new_[12026]_  | ~\new_[9983]_ ;
  assign \new_[7740]_  = ~\new_[9807]_  | ~\new_[11792]_ ;
  assign \new_[7741]_  = ~\new_[9844]_  | ~\new_[11741]_ ;
  assign \new_[7742]_  = ~\new_[14878]_  | ~\new_[9855]_ ;
  assign \new_[7743]_  = ~\new_[9895]_  | ~\new_[11913]_ ;
  assign \new_[7744]_  = ~\new_[9908]_  | ~\new_[11922]_ ;
  assign \new_[7745]_  = ~\new_[11874]_  | ~\new_[9913]_ ;
  assign \new_[7746]_  = ~\new_[12878]_  & ~\new_[10043]_ ;
  assign \new_[7747]_  = ~\new_[12908]_  & (~\new_[12053]_  | ~\new_[19064]_ );
  assign \new_[7748]_  = (~\new_[14432]_  & ~\new_[18809]_ ) | (~\new_[17969]_  & ~\new_[14677]_ );
  assign \new_[7749]_  = ~\new_[10265]_  & ~\new_[11256]_ ;
  assign \new_[7750]_  = ~\new_[13185]_  & (~\new_[12098]_  | ~\new_[18542]_ );
  assign \new_[7751]_  = ~\new_[10190]_  & (~\new_[12730]_  | ~\new_[21056]_ );
  assign \new_[7752]_  = ~\new_[10066]_  & (~\new_[13212]_  | ~\new_[18046]_ );
  assign \new_[7753]_  = ~\new_[10305]_  & (~\new_[20163]_  | ~\new_[19094]_ );
  assign \new_[7754]_  = ~\new_[14280]_  & (~\new_[13528]_  | ~\new_[18643]_ );
  assign \new_[7755]_  = ~\new_[10263]_  | ~\new_[10222]_ ;
  assign \new_[7756]_  = ~\new_[12029]_  | (~\new_[10855]_  & ~\new_[19044]_ );
  assign \new_[7757]_  = ~\new_[10164]_  | ~\new_[11729]_ ;
  assign \new_[7758]_  = ~\new_[12625]_  | ~\new_[15017]_  | ~\new_[17101]_  | ~\new_[15046]_ ;
  assign \new_[7759]_  = ~\new_[11666]_  | ~\new_[11305]_  | ~\new_[16586]_ ;
  assign \new_[7760]_  = ~\new_[10161]_  | ~\new_[10649]_ ;
  assign \new_[7761]_  = ~\new_[10123]_  | ~\new_[10629]_ ;
  assign \new_[7762]_  = (~\new_[17405]_  | ~\new_[18981]_ ) & (~\new_[12165]_  | ~\new_[19156]_ );
  assign \new_[7763]_  = ~\new_[10244]_  | ~\new_[10679]_ ;
  assign \new_[7764]_  = ~\new_[10270]_  | ~\new_[10622]_ ;
  assign \new_[7765]_  = ~\new_[10338]_  | ~\new_[10683]_ ;
  assign \new_[7766]_  = ~\new_[10287]_  | ~\new_[13183]_ ;
  assign \new_[7767]_  = ~\new_[10122]_  | ~\new_[10688]_ ;
  assign \new_[7768]_  = \new_[11754]_  ? \new_[18937]_  : \new_[14052]_ ;
  assign \new_[7769]_  = \new_[11893]_  ? \new_[21629]_  : \new_[16229]_ ;
  assign \new_[7770]_  = ~\new_[10999]_  & (~\new_[11906]_  | ~\new_[21556]_ );
  assign \new_[7771]_  = \new_[12016]_  ? \new_[17960]_  : \new_[16195]_ ;
  assign \new_[7772]_  = \new_[11795]_  ? \new_[19088]_  : \new_[14897]_ ;
  assign \new_[7773]_  = ~\new_[8741]_ ;
  assign \new_[7774]_  = ~\new_[10596]_  & ~\new_[14951]_ ;
  assign \new_[7775]_  = ~\new_[12871]_  | ~\new_[17469]_ ;
  assign \new_[7776]_  = ~\new_[10705]_  | ~\new_[19088]_ ;
  assign \new_[7777]_  = ~\new_[8743]_ ;
  assign \new_[7778]_  = ~\new_[10698]_  | ~\new_[17689]_ ;
  assign \new_[7779]_  = ~\new_[8745]_ ;
  assign \new_[7780]_  = ~\new_[8746]_ ;
  assign \new_[7781]_  = ~\new_[21594]_  & ~\new_[18863]_ ;
  assign \new_[7782]_  = ~\new_[10633]_  | ~\new_[19728]_ ;
  assign \new_[7783]_  = ~\new_[8751]_ ;
  assign \new_[7784]_  = ~\new_[10632]_  | ~\new_[21307]_ ;
  assign \new_[7785]_  = \new_[13477]_  | \new_[18925]_  | \new_[19068]_  | \new_[19044]_ ;
  assign \new_[7786]_  = ~\new_[8757]_ ;
  assign \new_[7787]_  = ~\new_[10651]_  | ~\new_[16695]_ ;
  assign \new_[7788]_  = ~\new_[8759]_ ;
  assign \new_[7789]_  = ~\new_[21679]_  | ~\new_[21510]_ ;
  assign \new_[7790]_  = ~\new_[10676]_  | ~\new_[17115]_ ;
  assign \new_[7791]_  = ~\new_[10660]_  | ~\new_[19247]_ ;
  assign \new_[7792]_  = ~\new_[8766]_ ;
  assign \new_[7793]_  = ~\new_[10659]_  & ~\new_[17689]_ ;
  assign \new_[7794]_  = ~\new_[8767]_ ;
  assign \new_[7795]_  = ~\new_[10581]_  | ~\new_[21115]_ ;
  assign \new_[7796]_  = ~\new_[8769]_ ;
  assign \new_[7797]_  = ~\new_[10662]_  | ~\new_[21562]_ ;
  assign \new_[7798]_  = ~\new_[10578]_  | ~\new_[18840]_ ;
  assign \new_[7799]_  = ~\new_[10607]_  | ~\new_[17837]_ ;
  assign \new_[7800]_  = ~\new_[12869]_  | ~\new_[18974]_ ;
  assign \new_[7801]_  = ~\new_[8778]_ ;
  assign \new_[7802]_  = ~\new_[12697]_  | ~\new_[18077]_ ;
  assign \new_[7803]_  = ~\new_[10514]_  | ~\new_[18427]_ ;
  assign \new_[7804]_  = ~\new_[19711]_  & ~\new_[10530]_ ;
  assign \new_[7805]_  = ~\new_[10550]_  | ~\new_[19085]_ ;
  assign \new_[7806]_  = ~\new_[8790]_ ;
  assign \new_[7807]_  = \new_[12197]_  | \new_[18925]_  | \new_[19625]_  | \new_[21168]_ ;
  assign \new_[7808]_  = ~\new_[10738]_  | ~\new_[18652]_ ;
  assign \new_[7809]_  = ~\new_[8796]_ ;
  assign \new_[7810]_  = ~\new_[8798]_ ;
  assign \new_[7811]_  = ~\new_[21562]_  | ~\new_[21390]_ ;
  assign \new_[7812]_  = ~\new_[10591]_  & ~\new_[14951]_ ;
  assign \new_[7813]_  = ~\new_[8802]_ ;
  assign \new_[7814]_  = ~\new_[10588]_  | ~\new_[19450]_ ;
  assign \new_[7815]_  = ~\new_[8803]_ ;
  assign \new_[7816]_  = ~\new_[8806]_ ;
  assign \new_[7817]_  = ~\new_[8807]_ ;
  assign \new_[7818]_  = ~\new_[8808]_ ;
  assign \new_[7819]_  = ~\new_[13605]_  & ~\new_[19079]_  & ~\new_[16850]_ ;
  assign \new_[7820]_  = ~\new_[8813]_ ;
  assign \new_[7821]_  = ~\new_[10642]_  | ~\new_[18361]_ ;
  assign \new_[7822]_  = ~\new_[8814]_ ;
  assign \new_[7823]_  = \new_[12446]_  & \new_[18194]_ ;
  assign \new_[7824]_  = ~\new_[10652]_  | ~\new_[19381]_ ;
  assign \new_[7825]_  = ~\new_[8818]_ ;
  assign \new_[7826]_  = ~\new_[8820]_ ;
  assign \new_[7827]_  = ~\new_[8822]_ ;
  assign \new_[7828]_  = ~\new_[10566]_  | ~\new_[13539]_ ;
  assign \new_[7829]_  = ~\new_[10552]_  & ~\new_[12583]_ ;
  assign \new_[7830]_  = ~\new_[18973]_  & ~\new_[10682]_ ;
  assign \new_[7831]_  = ~\new_[21475]_ ;
  assign \new_[7832]_  = ~\new_[21476]_ ;
  assign \new_[7833]_  = ~\new_[8830]_ ;
  assign \new_[7834]_  = \new_[10637]_  | \new_[18166]_ ;
  assign \new_[7835]_  = ~\new_[12146]_  & ~\new_[15788]_ ;
  assign \new_[7836]_  = ~\new_[10593]_  | ~\new_[11650]_ ;
  assign \new_[7837]_  = \new_[10718]_  & \new_[19208]_ ;
  assign \new_[7838]_  = \new_[10605]_  | \new_[18288]_ ;
  assign \new_[7839]_  = ~\new_[8836]_ ;
  assign \new_[7840]_  = \new_[12158]_  | \new_[18941]_ ;
  assign \new_[7841]_  = \new_[10505]_  & \new_[15140]_ ;
  assign \new_[7842]_  = ~\new_[10700]_  & (~\new_[18370]_  | ~\new_[19081]_ );
  assign \new_[7843]_  = ~\new_[8843]_ ;
  assign \new_[7844]_  = ~\new_[10641]_  | ~\new_[17347]_ ;
  assign \new_[7845]_  = ~\new_[13962]_  | ~\new_[12780]_ ;
  assign \new_[7846]_  = ~\new_[8852]_ ;
  assign \new_[7847]_  = ~\new_[8853]_ ;
  assign \new_[7848]_  = ~\new_[13205]_  & ~\new_[14069]_ ;
  assign \new_[7849]_  = ~\new_[10566]_  | ~\new_[16769]_ ;
  assign \new_[7850]_  = ~\new_[20726]_ ;
  assign \new_[7851]_  = ~\new_[15480]_  | ~\new_[13173]_ ;
  assign \new_[7852]_  = ~\new_[10585]_  | ~\new_[11266]_ ;
  assign \new_[7853]_  = ~\new_[16284]_  & ~\new_[10552]_ ;
  assign \new_[7854]_  = ~\new_[13155]_  & ~\new_[15639]_ ;
  assign \new_[7855]_  = ~\new_[8873]_ ;
  assign \new_[7856]_  = ~\new_[8874]_ ;
  assign \new_[7857]_  = ~\new_[8876]_ ;
  assign \new_[7858]_  = ~\new_[10580]_  & ~\new_[14996]_ ;
  assign \new_[7859]_  = ~\new_[18233]_  & ~\new_[12780]_ ;
  assign \new_[7860]_  = ~\new_[17549]_  | ~\new_[13251]_ ;
  assign \new_[7861]_  = \new_[18644]_  & \new_[12744]_ ;
  assign \new_[7862]_  = ~\new_[10543]_  & ~\new_[18973]_ ;
  assign \new_[7863]_  = ~\new_[17770]_  | ~\new_[12495]_ ;
  assign \new_[7864]_  = ~\new_[10524]_  | ~\new_[14093]_ ;
  assign \new_[7865]_  = ~\new_[18403]_  | ~\new_[21662]_ ;
  assign \new_[7866]_  = ~\new_[8885]_ ;
  assign \new_[7867]_  = ~\new_[11520]_  | ~\new_[20809]_ ;
  assign \new_[7868]_  = ~\new_[12980]_  | ~\new_[15029]_ ;
  assign \new_[7869]_  = ~\new_[8887]_ ;
  assign \new_[7870]_  = ~\new_[18597]_  | ~\new_[10702]_ ;
  assign \new_[7871]_  = \new_[10595]_  | \new_[19233]_ ;
  assign \new_[7872]_  = \new_[12646]_  | \new_[18798]_ ;
  assign \new_[7873]_  = ~\new_[10733]_  | ~\new_[14184]_ ;
  assign \new_[7874]_  = ~\new_[8899]_ ;
  assign \new_[7875]_  = ~\new_[10651]_  | ~\new_[17359]_ ;
  assign \new_[7876]_  = ~\new_[10682]_  | ~\new_[17408]_ ;
  assign \new_[7877]_  = ~\new_[8908]_ ;
  assign \new_[7878]_  = ~\new_[14173]_  | ~\new_[12788]_ ;
  assign \new_[7879]_  = ~\new_[8916]_ ;
  assign \new_[7880]_  = ~\new_[15763]_  | ~\new_[13061]_ ;
  assign \new_[7881]_  = ~\new_[13213]_  | ~\new_[12424]_ ;
  assign \new_[7882]_  = ~\new_[13213]_  | ~\new_[11681]_ ;
  assign \new_[7883]_  = ~\new_[13770]_  & ~\new_[12904]_ ;
  assign \new_[7884]_  = ~\new_[13253]_  | ~\new_[12424]_ ;
  assign \new_[7885]_  = ~\new_[10544]_  & ~\new_[14031]_ ;
  assign \new_[7886]_  = ~\new_[12687]_  | ~\new_[18427]_ ;
  assign \new_[7887]_  = ~\new_[8922]_ ;
  assign \new_[7888]_  = \new_[12524]_  | \new_[18166]_ ;
  assign \new_[7889]_  = ~\new_[13730]_  & (~\new_[11963]_  | ~\new_[18011]_ );
  assign \new_[7890]_  = ~\new_[13624]_  & ~\new_[12164]_ ;
  assign \new_[7891]_  = ~\new_[8926]_ ;
  assign \new_[7892]_  = ~\new_[13047]_  | ~\new_[19036]_ ;
  assign \new_[7893]_  = ~\new_[12559]_  | ~\new_[21510]_ ;
  assign \new_[7894]_  = ~\new_[17944]_  | ~\new_[10650]_ ;
  assign \new_[7895]_  = ~\new_[12776]_  & ~\new_[11564]_ ;
  assign \new_[7896]_  = ~\new_[20163]_  & (~\new_[18276]_  | ~\new_[18861]_ );
  assign \new_[7897]_  = ~\new_[12766]_  & ~\new_[12393]_ ;
  assign \new_[7898]_  = ~\new_[8954]_ ;
  assign \new_[7899]_  = ~\new_[10632]_  | ~\new_[20661]_ ;
  assign \new_[7900]_  = ~\new_[9672]_  | ~\new_[21115]_ ;
  assign \new_[7901]_  = ~\new_[15656]_  | ~\new_[12877]_ ;
  assign \new_[7902]_  = ~\new_[10547]_  & ~\new_[11827]_ ;
  assign \new_[7903]_  = ~\new_[20713]_  | (~\new_[16062]_  & ~\new_[18717]_ );
  assign \new_[7904]_  = \new_[17840]_  & \new_[10561]_ ;
  assign \new_[7905]_  = ~\new_[8978]_ ;
  assign \new_[7906]_  = ~\new_[12691]_  & ~\new_[18731]_ ;
  assign \new_[7907]_  = ~\new_[8983]_ ;
  assign \new_[7908]_  = ~\new_[17742]_  & ~\new_[20809]_ ;
  assign \new_[7909]_  = ~\new_[13242]_  | ~\new_[19084]_ ;
  assign \new_[7910]_  = ~\new_[20435]_ ;
  assign \new_[7911]_  = ~\new_[8990]_ ;
  assign \new_[7912]_  = \new_[18557]_  & \new_[12617]_ ;
  assign \new_[7913]_  = ~\new_[12784]_  | ~\new_[18111]_ ;
  assign \new_[7914]_  = ~\new_[13990]_  & ~\new_[10647]_ ;
  assign \new_[7915]_  = ~\new_[8998]_ ;
  assign \new_[7916]_  = ~\new_[12798]_  & ~\new_[11587]_ ;
  assign \new_[7917]_  = ~\new_[9000]_ ;
  assign \new_[7918]_  = ~\new_[9004]_ ;
  assign \new_[7919]_  = ~\new_[16818]_  | ~\new_[13076]_ ;
  assign \new_[7920]_  = \new_[17468]_  & \new_[10514]_ ;
  assign \new_[7921]_  = ~\new_[9014]_ ;
  assign \new_[7922]_  = ~\new_[9015]_ ;
  assign \new_[7923]_  = ~\new_[19229]_  | ~\new_[21546]_  | ~\new_[20680]_ ;
  assign \new_[7924]_  = \new_[14241]_  & \new_[10555]_ ;
  assign \new_[7925]_  = ~\new_[12775]_  | ~\new_[13114]_ ;
  assign \new_[7926]_  = ~\new_[12534]_  | ~\new_[18355]_ ;
  assign \new_[7927]_  = ~\new_[13212]_  & (~\new_[16022]_  | ~\new_[19039]_ );
  assign \new_[7928]_  = ~\new_[12492]_  | ~\new_[19587]_ ;
  assign \new_[7929]_  = ~\new_[10527]_  & ~\new_[11746]_ ;
  assign \new_[7930]_  = ~\new_[9039]_ ;
  assign \new_[7931]_  = ~\new_[9043]_ ;
  assign \new_[7932]_  = ~\new_[17461]_  | ~\new_[10550]_ ;
  assign \new_[7933]_  = ~\new_[10518]_  & ~\new_[16181]_ ;
  assign \new_[7934]_  = ~\new_[13703]_  & ~\new_[18427]_ ;
  assign \new_[7935]_  = ~\new_[12362]_  | ~\new_[19299]_ ;
  assign \new_[7936]_  = ~\new_[9054]_ ;
  assign \new_[7937]_  = ~\new_[10562]_  & ~\new_[16244]_ ;
  assign \new_[7938]_  = ~\new_[10568]_  & ~\new_[15009]_ ;
  assign \new_[7939]_  = \new_[20698]_  & \new_[16827]_ ;
  assign \new_[7940]_  = ~\new_[10512]_  & ~\new_[12721]_ ;
  assign \new_[7941]_  = ~\new_[10576]_  | ~\new_[10515]_ ;
  assign \new_[7942]_  = ~\new_[10529]_  & ~\new_[14028]_ ;
  assign \new_[7943]_  = \new_[10538]_  | \new_[17598]_ ;
  assign \new_[7944]_  = ~\new_[12780]_  | ~\new_[14358]_ ;
  assign \new_[7945]_  = ~\new_[18166]_  & (~\new_[16296]_  | ~\new_[11663]_ );
  assign \new_[7946]_  = ~\new_[12244]_  | ~\new_[21689]_ ;
  assign \new_[7947]_  = ~\new_[10566]_  | ~\new_[13935]_ ;
  assign \new_[7948]_  = ~\new_[10710]_  & ~\new_[12711]_ ;
  assign \new_[7949]_  = ~\new_[12465]_  | ~\new_[11499]_ ;
  assign \new_[7950]_  = ~\new_[10660]_  | ~\new_[18982]_ ;
  assign \new_[7951]_  = ~\new_[10525]_  & ~\new_[18747]_ ;
  assign \new_[7952]_  = ~\new_[12326]_  | ~\new_[11849]_ ;
  assign \new_[7953]_  = ~\new_[9098]_ ;
  assign \new_[7954]_  = ~\new_[10592]_  | ~\new_[14231]_ ;
  assign \new_[7955]_  = ~\new_[10690]_  | ~\new_[21638]_ ;
  assign \new_[7956]_  = \new_[13689]_  & \new_[10543]_ ;
  assign \new_[7957]_  = ~\new_[9111]_ ;
  assign \new_[7958]_  = ~\new_[9115]_ ;
  assign \new_[7959]_  = ~\new_[10693]_  | ~\new_[18937]_ ;
  assign \new_[7960]_  = ~\new_[16356]_  | ~\new_[10617]_ ;
  assign \new_[7961]_  = ~\new_[9121]_ ;
  assign \new_[7962]_  = ~\new_[12537]_  | ~\new_[16972]_ ;
  assign \new_[7963]_  = ~\new_[9125]_ ;
  assign \new_[7964]_  = ~\new_[10675]_  & ~\new_[17131]_ ;
  assign \new_[7965]_  = ~\new_[9130]_ ;
  assign \new_[7966]_  = ~\new_[9131]_ ;
  assign \new_[7967]_  = ~\new_[20484]_ ;
  assign \new_[7968]_  = ~\new_[9136]_ ;
  assign \new_[7969]_  = ~\new_[14695]_  & ~\new_[12533]_ ;
  assign \new_[7970]_  = ~\new_[10692]_  | ~\new_[19587]_ ;
  assign \new_[7971]_  = ~\new_[9144]_ ;
  assign \new_[7972]_  = \new_[13468]_  | \new_[18166]_ ;
  assign \new_[7973]_  = ~\new_[10003]_  & ~\new_[14564]_ ;
  assign \new_[7974]_  = ~\new_[17113]_  | ~\new_[10578]_ ;
  assign \new_[7975]_  = ~\new_[9161]_ ;
  assign \new_[7976]_  = \new_[13395]_  | \new_[19102]_ ;
  assign \new_[7977]_  = ~\new_[9163]_ ;
  assign \new_[7978]_  = ~\new_[12019]_  & ~\new_[10709]_ ;
  assign \new_[7979]_  = ~\new_[13073]_  | ~\new_[10185]_ ;
  assign \new_[7980]_  = ~\new_[12853]_  & ~\new_[15476]_ ;
  assign \new_[7981]_  = ~\new_[10569]_  | ~\new_[9997]_ ;
  assign \new_[7982]_  = ~\new_[10579]_  & ~\new_[21693]_ ;
  assign \new_[7983]_  = \new_[12816]_  | \new_[18280]_ ;
  assign \new_[7984]_  = ~\new_[18762]_  & (~\new_[14890]_  | ~\new_[13605]_ );
  assign \new_[7985]_  = ~\new_[10653]_  | ~\new_[17041]_ ;
  assign \new_[7986]_  = ~\new_[10719]_  | ~\new_[14951]_ ;
  assign \new_[7987]_  = ~\new_[10725]_  | ~\new_[19088]_ ;
  assign \new_[7988]_  = ~\new_[10724]_  | ~\new_[19261]_ ;
  assign \new_[7989]_  = ~\new_[12093]_  & ~\new_[12433]_ ;
  assign \new_[7990]_  = ~\new_[10616]_  | ~\new_[17789]_ ;
  assign \new_[7991]_  = ~\new_[10720]_  | ~\new_[21115]_ ;
  assign \new_[7992]_  = ~\new_[14416]_  | (~\new_[12123]_  & ~\new_[19625]_ );
  assign \new_[7993]_  = ~\new_[13269]_  | ~\new_[9978]_ ;
  assign \new_[7994]_  = ~\new_[9203]_ ;
  assign \new_[7995]_  = ~\new_[15380]_  & ~\new_[10597]_ ;
  assign \new_[7996]_  = ~\new_[13465]_  & ~\new_[13289]_ ;
  assign \new_[7997]_  = ~\new_[12498]_  | ~\new_[10587]_ ;
  assign \new_[7998]_  = ~\new_[11698]_  | ~\new_[10206]_ ;
  assign \new_[7999]_  = ~\new_[10571]_  | ~\new_[20378]_ ;
  assign \new_[8000]_  = ~\new_[9217]_ ;
  assign \new_[8001]_  = ~\new_[10548]_  & (~\new_[18614]_  | ~\new_[17777]_ );
  assign \new_[8002]_  = ~\new_[12412]_  & (~\new_[15667]_  | ~\new_[19275]_ );
  assign \new_[8003]_  = ~\new_[11614]_  & ~\new_[10703]_ ;
  assign \new_[8004]_  = ~\new_[9220]_ ;
  assign \new_[8005]_  = ~\new_[10574]_  | ~\new_[14627]_ ;
  assign \new_[8006]_  = ~\new_[12573]_  | ~\new_[10695]_ ;
  assign \new_[8007]_  = ~\new_[18328]_  | (~\new_[14181]_  & ~\new_[21650]_ );
  assign \new_[8008]_  = ~\new_[17922]_  | (~\new_[16049]_  & ~\new_[12078]_ );
  assign \new_[8009]_  = ~\new_[18102]_  & (~\new_[18014]_  | ~\new_[12091]_ );
  assign \new_[8010]_  = ~\new_[18275]_  | (~\new_[17029]_  & ~\new_[12086]_ );
  assign \new_[8011]_  = \new_[10691]_  & \new_[19199]_ ;
  assign \new_[8012]_  = ~\new_[13675]_  & (~\new_[12120]_  | ~\new_[19088]_ );
  assign \new_[8013]_  = ~\new_[11986]_  | ~\new_[10836]_ ;
  assign \new_[8014]_  = ~\new_[13614]_  & (~\new_[10856]_  | ~\new_[19059]_ );
  assign \new_[8015]_  = ~\new_[10646]_  | ~\new_[10634]_ ;
  assign \new_[8016]_  = ~\new_[11743]_  | ~\new_[10648]_ ;
  assign \new_[8017]_  = ~\new_[13641]_  & (~\new_[12140]_  | ~\new_[20099]_ );
  assign \new_[8018]_  = \new_[18467]_  ^ \new_[10986]_ ;
  assign \new_[8019]_  = \new_[18611]_  ^ \new_[12113]_ ;
  assign \new_[8020]_  = \new_[18684]_  ^ \new_[12102]_ ;
  assign \new_[8021]_  = \new_[18820]_  ^ \new_[12100]_ ;
  assign \new_[8022]_  = \new_[18905]_  ^ \new_[12104]_ ;
  assign \new_[8023]_  = ~\new_[9256]_ ;
  assign \new_[8024]_  = \new_[18848]_  ^ \new_[12107]_ ;
  assign \new_[8025]_  = ~\new_[9259]_ ;
  assign \new_[8026]_  = ~\new_[9261]_ ;
  assign \new_[8027]_  = ~\new_[11355]_  & (~\new_[12132]_  | ~\new_[18849]_ );
  assign \new_[8028]_  = ~\new_[14125]_  | ~\new_[15042]_  | ~\new_[12105]_ ;
  assign \new_[8029]_  = ~\new_[10740]_  | ~\new_[19177]_ ;
  assign \new_[8030]_  = \new_[12757]_  | \new_[20492]_ ;
  assign \new_[8031]_  = ~\new_[11234]_  & (~\new_[12137]_  | ~\new_[18974]_ );
  assign \new_[8032]_  = \new_[14703]_  | \new_[21689]_ ;
  assign \new_[8033]_  = \new_[10012]_  | \new_[19204]_ ;
  assign \new_[8034]_  = ~\new_[10853]_  | ~\new_[9959]_  | ~\new_[11031]_ ;
  assign \new_[8035]_  = ~\new_[12879]_  | ~\new_[13357]_  | ~\new_[14109]_  | ~\new_[14455]_ ;
  assign \new_[8036]_  = \new_[15685]_  | \new_[18427]_ ;
  assign \new_[8037]_  = \new_[15710]_  | \new_[18973]_ ;
  assign \new_[8038]_  = (~\new_[12127]_  | ~\new_[19553]_ ) & (~\new_[15559]_  | ~\new_[17640]_ );
  assign \new_[8039]_  = ~\new_[10746]_  & ~\new_[10888]_ ;
  assign \new_[8040]_  = ~\new_[19711]_  & (~\new_[11734]_  | ~\new_[15499]_ );
  assign \new_[8041]_  = ~\new_[9277]_ ;
  assign n2698 = ~\new_[19363]_  & (~\new_[12084]_  | ~\new_[14785]_ );
  assign \new_[8043]_  = ~\new_[17552]_  & ~\new_[13356]_ ;
  assign \new_[8044]_  = ~\new_[17830]_  | ~\new_[15949]_  | ~\new_[9782]_  | ~\new_[14486]_ ;
  assign \new_[8045]_  = ~\new_[17786]_  & ~\new_[10737]_ ;
  assign \new_[8046]_  = ~\new_[9890]_  & (~\new_[12126]_  | ~\new_[18402]_ );
  assign \new_[8047]_  = (~\new_[10873]_  | ~\new_[19727]_ ) & (~\new_[18849]_  | ~\new_[18590]_ );
  assign \new_[8048]_  = (~\new_[10872]_  | ~\new_[18965]_ ) & (~\new_[18981]_  | ~\new_[17761]_ );
  assign \new_[8049]_  = ~\new_[17787]_  | ~\new_[16159]_  | ~\new_[9783]_  | ~\new_[14805]_ ;
  assign \new_[8050]_  = ~\new_[12734]_  | ~\new_[14949]_  | ~\new_[11398]_  | ~\new_[12125]_ ;
  assign \new_[8051]_  = ~\new_[11221]_  & (~\new_[12136]_  | ~\new_[21633]_ );
  assign \new_[8052]_  = ~\new_[9303]_ ;
  assign \new_[8053]_  = ~\new_[10744]_  | ~\new_[16394]_ ;
  assign \new_[8054]_  = ~\new_[19064]_  | (~\new_[11114]_  & ~\new_[21468]_ );
  assign \new_[8055]_  = ~\new_[18569]_  | (~\new_[11205]_  & ~\new_[14157]_ );
  assign \new_[8056]_  = ~\new_[19059]_  | (~\new_[11279]_  & ~\new_[14168]_ );
  assign \new_[8057]_  = ~\new_[13260]_  | ~\new_[19269]_ ;
  assign \new_[8058]_  = ~\new_[19202]_  | (~\new_[11136]_  & ~\new_[12825]_ );
  assign \new_[8059]_  = ~\new_[19094]_  | (~\new_[11324]_  & ~\new_[15261]_ );
  assign \new_[8060]_  = ~\new_[18046]_  | (~\new_[11231]_  & ~\new_[13148]_ );
  assign \new_[8061]_  = ~\new_[9674]_  | ~\new_[19021]_ ;
  assign \new_[8062]_  = ~\new_[19079]_  | (~\new_[11208]_  & ~\new_[14107]_ );
  assign \new_[8063]_  = ~\new_[21702]_  & ~\new_[19748]_ ;
  assign \new_[8064]_  = ~\new_[9731]_  | ~\new_[19299]_ ;
  assign \new_[8065]_  = ~\new_[18627]_  | (~\new_[11327]_  & ~\new_[14355]_ );
  assign \new_[8066]_  = ~\new_[18077]_  | (~\new_[11298]_  & ~\new_[14041]_ );
  assign \new_[8067]_  = ~\new_[19050]_  | (~\new_[11259]_  & ~\new_[15419]_ );
  assign \new_[8068]_  = ~\new_[19049]_  & (~\new_[11934]_  | ~\new_[11051]_ );
  assign \new_[8069]_  = ~\new_[19336]_  & (~\new_[13087]_  | ~\new_[11067]_ );
  assign \new_[8070]_  = ~\new_[9296]_ ;
  assign \new_[8071]_  = ~\new_[18194]_  | (~\new_[11123]_  & ~\new_[13915]_ );
  assign \new_[8072]_  = ~\new_[19244]_  | (~\new_[11262]_  & ~\new_[11667]_ );
  assign \new_[8073]_  = ~\new_[18046]_  | (~\new_[12403]_  & ~\new_[11531]_ );
  assign \new_[8074]_  = ~\new_[19266]_  | (~\new_[12407]_  & ~\new_[11662]_ );
  assign \new_[8075]_  = ~\new_[21115]_  | (~\new_[12411]_  & ~\new_[11664]_ );
  assign \new_[8076]_  = ~\new_[18280]_  | (~\new_[11120]_  & ~\new_[12529]_ );
  assign \new_[8077]_  = ~\new_[13606]_  | ~\new_[10883]_  | ~\new_[14904]_ ;
  assign \new_[8078]_  = ~\new_[10756]_  | ~\new_[13796]_ ;
  assign \new_[8079]_  = ~\new_[20686]_  | (~\new_[16297]_  & ~\new_[11147]_ );
  assign \new_[8080]_  = ~\new_[14505]_  | ~\new_[15911]_  | ~\new_[10932]_ ;
  assign \new_[8081]_  = ~\new_[9329]_ ;
  assign \new_[8082]_  = ~\new_[18137]_  | (~\new_[15969]_  & ~\new_[11237]_ );
  assign \new_[8083]_  = ~\new_[9332]_ ;
  assign \new_[8084]_  = ~\new_[19384]_  | (~\new_[13507]_  & ~\new_[11190]_ );
  assign \new_[8085]_  = ~\new_[9334]_ ;
  assign \new_[8086]_  = ~\new_[20701]_  | (~\new_[12802]_  & ~\new_[11191]_ );
  assign \new_[8087]_  = ~\new_[19237]_  | (~\new_[12755]_  & ~\new_[11377]_ );
  assign \new_[8088]_  = ~\new_[18840]_  | (~\new_[12297]_  & ~\new_[11767]_ );
  assign \new_[8089]_  = ~\new_[21508]_  | (~\new_[11089]_  & ~\new_[13020]_ );
  assign \new_[8090]_  = ~\new_[18166]_  | (~\new_[11115]_  & ~\new_[11154]_ );
  assign \new_[8091]_  = ~\new_[19240]_  | (~\new_[11426]_  & ~\new_[15669]_ );
  assign \new_[8092]_  = ~\new_[19592]_  | (~\new_[11169]_  & ~\new_[12492]_ );
  assign \new_[8093]_  = ~\new_[19266]_  | (~\new_[11402]_  & ~\new_[13711]_ );
  assign \new_[8094]_  = ~\new_[19233]_  | (~\new_[11415]_  & ~\new_[21094]_ );
  assign \new_[8095]_  = ~\new_[19202]_  | (~\new_[11416]_  & ~\new_[12362]_ );
  assign \new_[8096]_  = \new_[17997]_  | \new_[10729]_ ;
  assign \new_[8097]_  = ~\new_[10763]_  | ~\new_[16394]_ ;
  assign \new_[8098]_  = ~\new_[19249]_  | (~\new_[12611]_  & ~\new_[11423]_ );
  assign \new_[8099]_  = ~\new_[18692]_  | (~\new_[11796]_  & ~\new_[15074]_ );
  assign \new_[8100]_  = ~\new_[11499]_  | ~\new_[11500]_  | ~\new_[11095]_ ;
  assign \new_[8101]_  = ~\new_[18821]_  | (~\new_[11476]_  & ~\new_[15438]_ );
  assign \new_[8102]_  = ~\new_[9694]_  | ~\new_[19559]_ ;
  assign \new_[8103]_  = ~\new_[10753]_  | ~\new_[14955]_ ;
  assign \new_[8104]_  = ~\new_[18569]_  | (~\new_[11477]_  & ~\new_[14751]_ );
  assign \new_[8105]_  = ~\new_[9667]_  | ~\new_[14598]_ ;
  assign \new_[8106]_  = \new_[10787]_  & \new_[12723]_ ;
  assign \new_[8107]_  = ~\new_[10395]_  & ~\new_[10789]_ ;
  assign \new_[8108]_  = ~\new_[9347]_ ;
  assign \new_[8109]_  = \new_[10793]_  & \new_[11187]_ ;
  assign \new_[8110]_  = ~\new_[15044]_  & (~\new_[11142]_  | ~\new_[19553]_ );
  assign \new_[8111]_  = ~\new_[11525]_  | ~\new_[11725]_  | ~\new_[12305]_ ;
  assign \new_[8112]_  = ~\new_[19070]_  | (~\new_[12431]_  & ~\new_[14127]_ );
  assign \new_[8113]_  = ~\new_[19727]_  | (~\new_[11485]_  & ~\new_[17855]_ );
  assign \new_[8114]_  = ~\new_[13558]_  | ~\new_[15169]_  | ~\new_[11870]_ ;
  assign \new_[8115]_  = ~\new_[9706]_  | ~\new_[19377]_ ;
  assign \new_[8116]_  = ~\new_[10933]_  | (~\new_[10918]_  & ~\new_[18087]_ );
  assign n2703 = ~\new_[10752]_  & ~n3423;
  assign n2708 = ~\new_[10741]_  & ~n3423;
  assign \new_[8119]_  = ~\new_[12251]_  | ~\new_[11688]_  | ~\new_[11829]_ ;
  assign \new_[8120]_  = ~\new_[18542]_  | (~\new_[11481]_  & ~\new_[15170]_ );
  assign \new_[8121]_  = ~\new_[9716]_  | ~\new_[19507]_ ;
  assign \new_[8122]_  = ~\new_[19366]_  & (~\new_[11177]_  | ~\new_[13603]_ );
  assign \new_[8123]_  = ~\new_[19079]_  | ~\new_[973]_  | ~\new_[11390]_ ;
  assign \new_[8124]_  = ~\new_[9355]_ ;
  assign \new_[8125]_  = ~\new_[19266]_  | (~\new_[11479]_  & ~\new_[13348]_ );
  assign \new_[8126]_  = \new_[10817]_  & \new_[18833]_ ;
  assign \new_[8127]_  = ~\new_[18194]_  & (~\new_[11164]_  | ~\new_[13883]_ );
  assign \new_[8128]_  = ~\new_[13571]_  | ~\new_[13847]_  | ~\new_[10969]_ ;
  assign \new_[8129]_  = ~\new_[18998]_  | (~\new_[11111]_  & ~\new_[16346]_ );
  assign \new_[8130]_  = ~\new_[9679]_  | ~\new_[21095]_ ;
  assign \new_[8131]_  = ~\new_[9720]_  | ~\new_[17447]_ ;
  assign \new_[8132]_  = ~\new_[10823]_  | ~\new_[21630]_ ;
  assign \new_[8133]_  = ~\new_[19349]_  | (~\new_[11588]_  & ~\new_[10980]_ );
  assign \new_[8134]_  = ~\new_[19592]_  | (~\new_[11482]_  & ~\new_[13349]_ );
  assign \new_[8135]_  = ~\new_[13584]_  | ~\new_[12838]_  | ~\new_[11739]_ ;
  assign \new_[8136]_  = ~\new_[11602]_  | ~\new_[11568]_  | ~\new_[12386]_ ;
  assign \new_[8137]_  = ~\new_[19094]_  | (~\new_[11483]_  & ~\new_[14734]_ );
  assign \new_[8138]_  = \new_[12142]_  | \new_[10360]_ ;
  assign \new_[8139]_  = ~\new_[10966]_  | ~\new_[11751]_  | ~\new_[13805]_ ;
  assign \new_[8140]_  = ~\new_[18693]_  | (~\new_[11484]_  & ~\new_[15430]_ );
  assign \new_[8141]_  = ~\new_[21562]_  | (~\new_[11480]_  & ~\new_[13479]_ );
  assign \new_[8142]_  = ~\new_[10839]_  | ~\new_[20433]_ ;
  assign \new_[8143]_  = ~\new_[9623]_  | ~\new_[20906]_ ;
  assign \new_[8144]_  = ~\new_[10885]_  | ~\new_[11854]_  | ~\new_[14134]_ ;
  assign \new_[8145]_  = ~\new_[18818]_  | (~\new_[11280]_  & ~\new_[15194]_ );
  assign \new_[8146]_  = ~\new_[19233]_  | (~\new_[11080]_  & ~\new_[15514]_ );
  assign \new_[8147]_  = ~\new_[18046]_  | ~\new_[19022]_  | ~\new_[11391]_ ;
  assign \new_[8148]_  = ~\new_[18965]_  | (~\new_[11151]_  & ~\new_[15467]_ );
  assign \new_[8149]_  = ~\new_[9678]_  & ~\new_[19003]_ ;
  assign \new_[8150]_  = ~\new_[19357]_  | (~\new_[11250]_  & ~\new_[16597]_ );
  assign \new_[8151]_  = ~\new_[18778]_  | (~\new_[11254]_  & ~\new_[13506]_ );
  assign \new_[8152]_  = ~\new_[19094]_  | ~\new_[19433]_  | ~\new_[11392]_ ;
  assign \new_[8153]_  = ~\new_[21635]_  | (~\new_[13398]_  & ~\new_[11257]_ );
  assign \new_[8154]_  = ~\new_[11782]_  | ~\new_[11444]_  | ~\new_[12349]_ ;
  assign \new_[8155]_  = ~\new_[19064]_  | (~\new_[11096]_  & ~\new_[15554]_ );
  assign \new_[8156]_  = \new_[9620]_  | \new_[20513]_ ;
  assign \new_[8157]_  = ~\new_[9664]_  | ~\new_[20971]_ ;
  assign \new_[8158]_  = ~\new_[13306]_  | ~\new_[10449]_  | ~\new_[11364]_ ;
  assign \new_[8159]_  = ~\new_[14023]_  | ~\new_[12683]_  | ~\new_[13552]_ ;
  assign \new_[8160]_  = ~\new_[9763]_  | ~\new_[19492]_ ;
  assign \new_[8161]_  = ~\new_[11361]_  | ~\new_[12463]_  | ~\new_[20987]_ ;
  assign \new_[8162]_  = ~\new_[20704]_  | (~\new_[11478]_  & ~\new_[15463]_ );
  assign \new_[8163]_  = ~\new_[9678]_  | ~\new_[13820]_ ;
  assign \new_[8164]_  = ~\new_[19064]_  & (~\new_[11382]_  | ~\new_[12602]_ );
  assign \new_[8165]_  = ~\new_[19492]_  | (~\new_[12804]_  & ~\new_[10934]_ );
  assign \new_[8166]_  = ~\new_[9708]_  & (~\new_[15892]_  | ~\new_[16568]_ );
  assign \new_[8167]_  = ~\new_[12212]_  | ~\new_[12520]_  | ~\new_[10172]_  | ~\new_[13435]_ ;
  assign \new_[8168]_  = ~\new_[10954]_  | ~\new_[9684]_  | ~\new_[14138]_ ;
  assign \new_[8169]_  = ~\new_[10973]_  | ~\new_[12358]_  | ~\new_[13851]_ ;
  assign \new_[8170]_  = ~\new_[14012]_  | ~\new_[10760]_ ;
  assign \new_[8171]_  = ~\new_[13572]_  | ~\new_[15050]_  | ~\new_[10257]_  | ~\new_[13157]_ ;
  assign \new_[8172]_  = ~\new_[11212]_  | ~\new_[11193]_  | ~\new_[11344]_ ;
  assign \new_[8173]_  = ~\new_[17689]_  & (~\new_[11436]_  | ~\new_[12584]_ );
  assign \new_[8174]_  = ~\new_[18606]_  & (~\new_[11430]_  | ~\new_[11542]_ );
  assign \new_[8175]_  = ~\new_[11867]_  | ~\new_[14515]_  | ~\new_[10915]_ ;
  assign \new_[8176]_  = ~\new_[19064]_  & (~\new_[11441]_  | ~\new_[16675]_ );
  assign \new_[8177]_  = ~\new_[21558]_  & (~\new_[11438]_  | ~\new_[14629]_ );
  assign \new_[8178]_  = ~\new_[19006]_  & (~\new_[11446]_  | ~\new_[16101]_ );
  assign \new_[8179]_  = ~\new_[18795]_  & (~\new_[10952]_  | ~\new_[21622]_ );
  assign \new_[8180]_  = ~\new_[19266]_  & (~\new_[11439]_  | ~\new_[11609]_ );
  assign \new_[8181]_  = ~\new_[9377]_ ;
  assign \new_[8182]_  = ~\new_[19687]_  & (~\new_[11435]_  | ~\new_[13825]_ );
  assign \new_[8183]_  = ~\new_[19204]_  & (~\new_[11447]_  | ~\new_[13780]_ );
  assign \new_[8184]_  = ~\new_[10790]_  | ~\new_[19659]_ ;
  assign \new_[8185]_  = \new_[10784]_  & \new_[21056]_ ;
  assign \new_[8186]_  = ~\new_[15174]_  | (~\new_[11268]_  & ~\new_[19408]_ );
  assign \new_[8187]_  = ~\new_[10625]_  | (~\new_[13655]_  & ~\new_[19145]_ );
  assign \new_[8188]_  = ~\new_[10777]_  & ~\new_[9962]_ ;
  assign \new_[8189]_  = ~\new_[13569]_  | ~\new_[10108]_  | ~\new_[13784]_ ;
  assign \new_[8190]_  = ~\new_[13158]_  | ~\new_[13834]_  | ~\new_[9847]_  | ~\new_[15243]_ ;
  assign \new_[8191]_  = ~\new_[10939]_  | ~\new_[12947]_  | ~\new_[14142]_ ;
  assign \new_[8192]_  = ~\new_[10167]_  | (~\new_[13630]_  & ~\new_[18833]_ );
  assign \new_[8193]_  = ~\new_[10905]_  | ~\new_[14102]_  | ~\new_[14340]_ ;
  assign \new_[8194]_  = ~\new_[13604]_  | ~\new_[15310]_  | ~\new_[11440]_ ;
  assign \new_[8195]_  = ~\new_[19790]_  | (~\new_[17002]_  & ~\new_[11224]_ );
  assign \new_[8196]_  = ~\new_[21165]_  | (~\new_[16502]_  & ~\new_[11275]_ );
  assign \new_[8197]_  = ~\new_[12253]_  | ~\new_[14229]_  | ~\new_[11901]_ ;
  assign \new_[8198]_  = ~\new_[14335]_  | ~\new_[10253]_  | ~\new_[13900]_ ;
  assign \new_[8199]_  = ~\new_[13596]_  | ~\new_[10273]_  | ~\new_[13701]_ ;
  assign \new_[8200]_  = ~\new_[13237]_  | ~\new_[12526]_  | ~\new_[11307]_  | ~\new_[13543]_ ;
  assign \new_[8201]_  = ~\new_[18124]_  & (~\new_[16525]_  | ~\new_[11356]_ );
  assign \new_[8202]_  = ~\new_[10981]_  | ~\new_[11858]_  | ~\new_[12025]_ ;
  assign \new_[8203]_  = ~\new_[18656]_  | (~\new_[17350]_  & ~\new_[11090]_ );
  assign \new_[8204]_  = ~\new_[18224]_  | (~\new_[16735]_  & ~\new_[11093]_ );
  assign \new_[8205]_  = ~\new_[19499]_  | (~\new_[20586]_  & ~\new_[11206]_ );
  assign \new_[8206]_  = ~\new_[19406]_  | (~\new_[14838]_  & ~\new_[11365]_ );
  assign \new_[8207]_  = ~\new_[19281]_  | (~\new_[15666]_  & ~\new_[11354]_ );
  assign \new_[8208]_  = ~\new_[12640]_  | ~\new_[11199]_  | ~\new_[11061]_ ;
  assign \new_[8209]_  = ~\new_[21691]_  | (~\new_[17092]_  & ~\new_[11335]_ );
  assign \new_[8210]_  = ~\new_[10797]_  & (~\new_[14856]_  | ~\new_[17734]_ );
  assign \new_[8211]_  = (~\new_[11467]_  | ~\new_[19578]_ ) & (~\new_[15793]_  | ~\new_[18544]_ );
  assign \new_[8212]_  = ~\new_[14313]_  | ~\new_[10145]_  | ~\new_[12180]_ ;
  assign \new_[8213]_  = ~\new_[13159]_  | ~\new_[12739]_  | ~\new_[10994]_ ;
  assign \new_[8214]_  = ~\new_[15326]_  | ~\new_[10303]_  | ~\new_[12265]_ ;
  assign \new_[8215]_  = ~\new_[13149]_  | ~\new_[11637]_  | ~\new_[11076]_ ;
  assign \new_[8216]_  = ~\new_[10795]_  & (~\new_[15206]_  | ~\new_[18750]_ );
  assign \new_[8217]_  = ~\new_[10165]_  & (~\new_[11434]_  | ~\new_[19803]_ );
  assign \new_[8218]_  = ~\new_[12212]_  | ~\new_[11186]_  | ~\new_[14598]_ ;
  assign \new_[8219]_  = ~\new_[10096]_  & (~\new_[12464]_  | ~\new_[19561]_ );
  assign \new_[8220]_  = ~\new_[13572]_  | ~\new_[11304]_  | ~\new_[21095]_ ;
  assign \new_[8221]_  = ~\new_[9777]_  & (~\new_[18527]_  | ~\new_[15759]_ );
  assign \new_[8222]_  = ~\new_[9682]_  | ~\new_[17789]_ ;
  assign \new_[8223]_  = ~\new_[9671]_  | ~\new_[16886]_ ;
  assign \new_[8224]_  = ~\new_[10794]_  & (~\new_[17640]_  | ~\new_[17990]_ );
  assign \new_[8225]_  = (~\new_[11417]_  | ~\new_[19625]_ ) & (~\new_[17840]_  | ~\new_[15469]_ );
  assign \new_[8226]_  = ~\new_[14273]_  & ~\new_[9666]_ ;
  assign \new_[8227]_  = \new_[10981]_  ? \new_[17689]_  : \new_[12627]_ ;
  assign \new_[8228]_  = (~\new_[11410]_  | ~\new_[18863]_ ) & (~\new_[17917]_  | ~\new_[15628]_ );
  assign \new_[8229]_  = ~\new_[15080]_  | ~\new_[13800]_  | ~\new_[10080]_  | ~\new_[13256]_ ;
  assign \new_[8230]_  = ~\new_[20158]_  | ~\new_[10306]_  | ~\new_[12387]_ ;
  assign \new_[8231]_  = ~\new_[19480]_  & (~\new_[11466]_  | ~\new_[17146]_ );
  assign \new_[8232]_  = ~\new_[10951]_  & ~\new_[10813]_ ;
  assign \new_[8233]_  = \new_[14936]_  ^ \new_[19419]_ ;
  assign \new_[8234]_  = ~\new_[11029]_  & ~\new_[9649]_ ;
  assign \new_[8235]_  = ~\new_[9658]_  & (~\new_[11621]_  | ~\new_[19247]_ );
  assign \new_[8236]_  = \new_[14763]_  ^ \new_[19532]_ ;
  assign \new_[8237]_  = ~\new_[9955]_  | ~\new_[9659]_ ;
  assign \new_[8238]_  = ~\new_[13105]_  & (~\new_[11429]_  | ~\new_[17578]_ );
  assign \new_[8239]_  = ~\new_[11804]_  & (~\new_[11428]_  | ~\new_[19098]_ );
  assign \new_[8240]_  = \new_[10939]_  ? \new_[18187]_  : \new_[14531]_ ;
  assign \new_[8241]_  = (~\new_[11274]_  | ~\new_[17447]_ ) & (~\new_[16241]_  | ~\new_[19727]_ );
  assign \new_[8242]_  = \new_[10905]_  ? \new_[18998]_  : \new_[14486]_ ;
  assign \new_[8243]_  = \new_[13566]_  ? \new_[19547]_  : \new_[14805]_ ;
  assign \new_[8244]_  = \new_[19805]_  ^ \new_[18209]_ ;
  assign \new_[8245]_  = ~\new_[21557]_  | (~\new_[11786]_  & ~\new_[14597]_ );
  assign \new_[8246]_  = ~\new_[19107]_  & (~\new_[11530]_  | ~\new_[14811]_ );
  assign \new_[8247]_  = \new_[10436]_  | \new_[21638]_ ;
  assign \new_[8248]_  = ~\new_[19711]_  | (~\new_[11490]_  & ~\new_[16560]_ );
  assign \new_[8249]_  = ~\new_[13537]_  | ~\new_[13140]_  | ~\new_[16043]_  | ~\new_[14152]_ ;
  assign \new_[8250]_  = ~\new_[10410]_  | ~\new_[10272]_ ;
  assign \new_[8251]_  = \new_[14760]_  ^ \new_[18011]_ ;
  assign \new_[8252]_  = \new_[10857]_  ^ \new_[18679]_ ;
  assign \new_[8253]_  = ~\new_[10422]_  & ~\new_[18288]_ ;
  assign \new_[8254]_  = ~\new_[9418]_ ;
  assign \new_[8255]_  = \new_[16692]_  ^ \new_[18194]_ ;
  assign \new_[8256]_  = ~\new_[21557]_  | (~\new_[11997]_  & ~\new_[14506]_ );
  assign \new_[8257]_  = ~\new_[21557]_  & (~\new_[11968]_  | ~\new_[12588]_ );
  assign \new_[8258]_  = ~\new_[9423]_ ;
  assign \new_[8259]_  = ~\new_[9424]_ ;
  assign \new_[8260]_  = ~\new_[19249]_  | (~\new_[12036]_  & ~\new_[14736]_ );
  assign \new_[8261]_  = ~\new_[19517]_  & (~\new_[13406]_  | ~\new_[12027]_ );
  assign \new_[8262]_  = ~\new_[9809]_  & ~\new_[19088]_ ;
  assign \new_[8263]_  = ~\new_[9861]_  & ~\new_[21056]_ ;
  assign \new_[8264]_  = ~\new_[9442]_ ;
  assign \new_[8265]_  = ~\new_[9443]_ ;
  assign \new_[8266]_  = \new_[18194]_  | \new_[10324]_ ;
  assign \new_[8267]_  = \new_[15351]_  | \new_[18794]_  | \new_[19261]_  | \new_[21695]_ ;
  assign \new_[8268]_  = \new_[9821]_  | \new_[19553]_ ;
  assign \new_[8269]_  = \new_[9832]_  | \new_[19547]_ ;
  assign \new_[8270]_  = ~\new_[9446]_ ;
  assign \new_[8271]_  = \new_[9830]_  | \new_[18965]_ ;
  assign \new_[8272]_  = ~\new_[9448]_ ;
  assign \new_[8273]_  = \new_[10094]_  & \new_[19206]_ ;
  assign \new_[8274]_  = ~\new_[9451]_ ;
  assign \new_[8275]_  = ~\new_[9814]_  | ~\new_[18965]_ ;
  assign \new_[8276]_  = ~\new_[10381]_  | ~\new_[18863]_ ;
  assign \new_[8277]_  = \new_[9836]_  | \new_[18998]_ ;
  assign \new_[8278]_  = ~\new_[9455]_ ;
  assign \new_[8279]_  = \new_[13410]_  | \new_[20490]_  | \new_[18847]_  | \new_[19095]_ ;
  assign \new_[8280]_  = ~\new_[9876]_  & ~\new_[19592]_ ;
  assign \new_[8281]_  = ~\new_[20306]_  & ~\new_[18077]_ ;
  assign \new_[8282]_  = \new_[9915]_  | \new_[21629]_ ;
  assign \new_[8283]_  = \new_[9923]_  | \new_[19202]_ ;
  assign \new_[8284]_  = \new_[11191]_  & \new_[16879]_ ;
  assign \new_[8285]_  = ~\new_[9927]_  | ~\new_[21630]_ ;
  assign \new_[8286]_  = \new_[13378]_  | \new_[21394]_  | \new_[21557]_  | \new_[18747]_ ;
  assign \new_[8287]_  = ~\new_[12440]_  | ~\new_[19233]_ ;
  assign \new_[8288]_  = ~\new_[9457]_ ;
  assign \new_[8289]_  = ~\new_[19085]_  | ~\new_[19357]_  | ~\new_[11911]_ ;
  assign \new_[8290]_  = ~\new_[9990]_  & ~\new_[19206]_ ;
  assign \new_[8291]_  = ~\new_[9985]_  & ~\new_[18606]_ ;
  assign \new_[8292]_  = ~\new_[9459]_ ;
  assign \new_[8293]_  = \new_[13431]_  | \new_[18362]_  | \new_[19592]_  | \new_[18325]_ ;
  assign \new_[8294]_  = ~\new_[9984]_  & ~\new_[19088]_ ;
  assign \new_[8295]_  = ~\new_[9835]_  | ~\new_[19727]_ ;
  assign \new_[8296]_  = ~\new_[10488]_  | ~\new_[19748]_ ;
  assign \new_[8297]_  = ~\new_[960]_  & (~\new_[13984]_  | ~\new_[11975]_ );
  assign \new_[8298]_  = ~\new_[10491]_  | ~\new_[18942]_ ;
  assign \new_[8299]_  = ~\new_[10493]_  | ~\new_[19702]_ ;
  assign \new_[8300]_  = ~\new_[1026]_  & (~\new_[12923]_  | ~\new_[11807]_ );
  assign \new_[8301]_  = ~\new_[10492]_  | ~\new_[20789]_ ;
  assign \new_[8302]_  = ~\new_[10487]_  | ~\new_[19229]_ ;
  assign \new_[8303]_  = ~\new_[19378]_  & (~\new_[12039]_  | ~\new_[13299]_ );
  assign \new_[8304]_  = ~\new_[19088]_  & (~\new_[14823]_  | ~\new_[11948]_ );
  assign \new_[8305]_  = ~\new_[19587]_  & (~\new_[13439]_  | ~\new_[11887]_ );
  assign \new_[8306]_  = ~\new_[19711]_  & (~\new_[16440]_  | ~\new_[11991]_ );
  assign \new_[8307]_  = ~\new_[10007]_  | ~\new_[10885]_ ;
  assign \new_[8308]_  = ~\new_[9468]_ ;
  assign \new_[8309]_  = ~\new_[10009]_  & ~\new_[13052]_ ;
  assign \new_[8310]_  = \new_[10010]_  | \new_[20680]_ ;
  assign \new_[8311]_  = ~\new_[11190]_  & ~\new_[13700]_ ;
  assign \new_[8312]_  = ~\new_[10443]_  & ~\new_[12846]_ ;
  assign \new_[8313]_  = \new_[10463]_  | \new_[17689]_ ;
  assign \new_[8314]_  = ~\new_[14005]_  | ~\new_[10591]_  | ~\new_[14078]_ ;
  assign \new_[8315]_  = ~\new_[11501]_  | ~\new_[14010]_  | ~\new_[15535]_ ;
  assign \new_[8316]_  = ~\new_[10021]_  | ~\new_[11207]_ ;
  assign \new_[8317]_  = \new_[10022]_  | \new_[19240]_ ;
  assign \new_[8318]_  = ~\new_[11524]_  | ~\new_[13696]_  | ~\new_[15650]_ ;
  assign \new_[8319]_  = ~\new_[9911]_  | ~\new_[9808]_ ;
  assign \new_[8320]_  = \new_[9809]_  & \new_[9984]_ ;
  assign \new_[8321]_  = ~\new_[11798]_  | ~\new_[9992]_ ;
  assign \new_[8322]_  = ~\new_[9851]_  | ~\new_[14033]_ ;
  assign \new_[8323]_  = \new_[10452]_  | \new_[18941]_ ;
  assign \new_[8324]_  = ~\new_[10080]_  & ~\new_[19547]_ ;
  assign \new_[8325]_  = ~\new_[12304]_  | ~\new_[12432]_ ;
  assign \new_[8326]_  = ~\new_[21058]_  | ~\new_[16143]_ ;
  assign \new_[8327]_  = ~\new_[18762]_  & (~\new_[11774]_  | ~\new_[16281]_ );
  assign \new_[8328]_  = \new_[10973]_  & \new_[9964]_ ;
  assign \new_[8329]_  = ~\new_[11503]_  | ~\new_[12780]_  | ~\new_[14529]_ ;
  assign \new_[8330]_  = ~\new_[9481]_ ;
  assign \new_[8331]_  = ~\new_[9856]_  | ~\new_[13613]_ ;
  assign \new_[8332]_  = ~\new_[9482]_ ;
  assign \new_[8333]_  = ~\new_[10128]_  | ~\new_[12938]_ ;
  assign \new_[8334]_  = ~\new_[10008]_  | ~\new_[21115]_ ;
  assign \new_[8335]_  = ~\new_[9952]_  | ~\new_[10682]_ ;
  assign \new_[8336]_  = ~\new_[12680]_  | ~\new_[13693]_  | ~\new_[15830]_  | ~\new_[11342]_ ;
  assign \new_[8337]_  = ~\new_[9833]_  | ~\new_[13558]_ ;
  assign \new_[8338]_  = ~\new_[15448]_  | ~\new_[13017]_  | ~\new_[11697]_ ;
  assign \new_[8339]_  = ~\new_[12095]_  | ~\new_[14491]_  | ~\new_[16513]_ ;
  assign \new_[8340]_  = ~\new_[9486]_ ;
  assign \new_[8341]_  = ~\new_[10000]_  | ~\new_[14287]_ ;
  assign \new_[8342]_  = ~\new_[12302]_  | ~\new_[10377]_ ;
  assign \new_[8343]_  = ~\new_[10981]_  | ~\new_[9939]_ ;
  assign \new_[8344]_  = ~\new_[11842]_  | ~\new_[9932]_ ;
  assign \new_[8345]_  = ~\new_[10473]_  | ~\new_[19032]_ ;
  assign \new_[8346]_  = \new_[10549]_  | \new_[19553]_ ;
  assign \new_[8347]_  = ~\new_[9972]_  | ~\new_[19532]_ ;
  assign \new_[8348]_  = ~\new_[9818]_  | ~\new_[14002]_ ;
  assign \new_[8349]_  = ~\new_[17244]_  & (~\new_[14274]_  | ~\new_[12067]_ );
  assign \new_[8350]_  = \new_[10478]_  | \new_[19453]_ ;
  assign \new_[8351]_  = ~\new_[10475]_  | ~\new_[19780]_ ;
  assign \new_[8352]_  = ~\new_[10483]_  | ~\new_[18194]_ ;
  assign \new_[8353]_  = ~\new_[10057]_  | ~\new_[18194]_ ;
  assign \new_[8354]_  = ~\new_[9496]_ ;
  assign \new_[8355]_  = ~\new_[9823]_  | ~\new_[11710]_ ;
  assign \new_[8356]_  = ~\new_[12540]_  | ~\new_[10549]_ ;
  assign \new_[8357]_  = ~\new_[9500]_ ;
  assign \new_[8358]_  = ~\new_[12175]_  | ~\new_[9866]_ ;
  assign \new_[8359]_  = \new_[10454]_  | \new_[18650]_ ;
  assign \new_[8360]_  = ~\new_[21600]_  | ~\new_[9998]_ ;
  assign \new_[8361]_  = ~\new_[10053]_  & ~\new_[11132]_ ;
  assign \new_[8362]_  = ~\new_[9506]_ ;
  assign \new_[8363]_  = ~\new_[12955]_  | ~\new_[9820]_ ;
  assign \new_[8364]_  = ~\new_[9986]_  | ~\new_[19045]_ ;
  assign \new_[8365]_  = ~\new_[9513]_ ;
  assign \new_[8366]_  = ~\new_[9514]_ ;
  assign \new_[8367]_  = ~\new_[9515]_ ;
  assign \new_[8368]_  = ~\new_[12310]_  | ~\new_[10519]_ ;
  assign \new_[8369]_  = ~\new_[19612]_  & (~\new_[11898]_  | ~\new_[16493]_ );
  assign \new_[8370]_  = \new_[13256]_  & \new_[9831]_ ;
  assign \new_[8371]_  = ~\new_[9520]_ ;
  assign \new_[8372]_  = ~\new_[10088]_  | ~\new_[16270]_ ;
  assign \new_[8373]_  = ~\new_[12302]_  & ~\new_[19088]_ ;
  assign \new_[8374]_  = ~\new_[21631]_  & (~\new_[14559]_  | ~\new_[14208]_ );
  assign \new_[8375]_  = \new_[9838]_  & \new_[14004]_ ;
  assign \new_[8376]_  = ~\new_[13979]_  | ~\new_[12601]_  | ~\new_[12299]_ ;
  assign \new_[8377]_  = ~\new_[15052]_  | ~\new_[9832]_  | ~\new_[14353]_ ;
  assign \new_[8378]_  = \new_[9828]_  & \new_[13552]_ ;
  assign \new_[8379]_  = \new_[9833]_  & \new_[12311]_ ;
  assign \new_[8380]_  = ~\new_[9530]_ ;
  assign \new_[8381]_  = ~\new_[10706]_  | ~\new_[9809]_ ;
  assign \new_[8382]_  = \new_[10162]_  & \new_[18965]_ ;
  assign \new_[8383]_  = ~\new_[9862]_  | ~\new_[12282]_ ;
  assign \new_[8384]_  = ~\new_[10094]_  & ~\new_[12781]_ ;
  assign \new_[8385]_  = ~\new_[10019]_  & ~\new_[20864]_ ;
  assign \new_[8386]_  = \new_[10417]_  | \new_[19064]_ ;
  assign \new_[8387]_  = \new_[9815]_  | \new_[19206]_ ;
  assign \new_[8388]_  = ~\new_[9537]_ ;
  assign \new_[8389]_  = \new_[9815]_  & \new_[10973]_ ;
  assign \new_[8390]_  = ~\new_[9544]_ ;
  assign \new_[8391]_  = \new_[9978]_  & \new_[15311]_ ;
  assign \new_[8392]_  = ~\new_[10405]_  | ~\new_[19520]_ ;
  assign \new_[8393]_  = ~\new_[10071]_  | ~\new_[12180]_ ;
  assign \new_[8394]_  = ~\new_[9846]_  | ~\new_[12208]_ ;
  assign \new_[8395]_  = \new_[10375]_  & \new_[12224]_ ;
  assign \new_[8396]_  = \new_[21054]_  | \new_[15901]_ ;
  assign \new_[8397]_  = ~\new_[12368]_  & ~\new_[19592]_ ;
  assign \new_[8398]_  = \new_[9910]_  | \new_[19711]_ ;
  assign \new_[8399]_  = ~\new_[9550]_ ;
  assign \new_[8400]_  = ~\new_[18249]_  & (~\new_[12082]_  | ~\new_[14063]_ );
  assign \new_[8401]_  = ~\new_[10048]_  | ~\new_[19727]_ ;
  assign \new_[8402]_  = ~\new_[21348]_ ;
  assign \new_[8403]_  = ~\new_[13763]_  | ~\new_[12596]_  | ~\new_[12945]_ ;
  assign \new_[8404]_  = ~\new_[9553]_ ;
  assign \new_[8405]_  = ~\new_[11013]_  & ~\new_[10057]_ ;
  assign \new_[8406]_  = ~\new_[12652]_  | ~\new_[13094]_  | ~\new_[10538]_  | ~\new_[12859]_ ;
  assign \new_[8407]_  = ~\new_[20222]_  & ~\new_[9933]_ ;
  assign \new_[8408]_  = ~\new_[13240]_  | ~\new_[10192]_ ;
  assign \new_[8409]_  = ~\new_[14104]_  | ~\new_[13847]_  | ~\new_[14267]_ ;
  assign \new_[8410]_  = ~\new_[10138]_  | ~\new_[11700]_ ;
  assign \new_[8411]_  = ~\new_[9555]_ ;
  assign \new_[8412]_  = ~\new_[12295]_  | ~\new_[11828]_ ;
  assign \new_[8413]_  = ~\new_[21074]_  | ~\new_[13755]_ ;
  assign \new_[8414]_  = \new_[10972]_  & \new_[9983]_ ;
  assign \new_[8415]_  = ~\new_[20809]_  | ~\new_[20705]_  | ~\new_[16510]_ ;
  assign \new_[8416]_  = ~\new_[9561]_ ;
  assign \new_[8417]_  = ~\new_[16669]_  & ~\new_[10329]_ ;
  assign \new_[8418]_  = ~\new_[12636]_  | ~\new_[13610]_  | ~\new_[12800]_  | ~\new_[12820]_ ;
  assign \new_[8419]_  = ~\new_[9969]_  | ~\new_[14289]_ ;
  assign \new_[8420]_  = ~\new_[14549]_  | ~\new_[14104]_  | ~\new_[13571]_ ;
  assign \new_[8421]_  = ~\new_[15929]_  | ~\new_[14391]_  | ~\new_[14023]_ ;
  assign \new_[8422]_  = \new_[20723]_  | \new_[10717]_ ;
  assign \new_[8423]_  = ~\new_[11191]_  & ~\new_[15327]_ ;
  assign \new_[8424]_  = ~\new_[9991]_  | ~\new_[12028]_ ;
  assign \new_[8425]_  = \new_[12321]_  & \new_[11586]_ ;
  assign \new_[8426]_  = ~\new_[9572]_ ;
  assign \new_[8427]_  = ~\new_[9836]_  | ~\new_[10904]_ ;
  assign \new_[8428]_  = ~\new_[9573]_ ;
  assign \new_[8429]_  = ~\new_[9993]_  | ~\new_[12858]_ ;
  assign \new_[8430]_  = \new_[10157]_  | \new_[18542]_ ;
  assign \new_[8431]_  = ~\new_[9959]_  | ~\new_[14201]_ ;
  assign \new_[8432]_  = \new_[12226]_  & \new_[18833]_ ;
  assign \new_[8433]_  = ~\new_[14387]_  | ~\new_[20660]_  | ~\new_[13695]_ ;
  assign \new_[8434]_  = ~\new_[10383]_  | ~\new_[18967]_ ;
  assign \new_[8435]_  = \new_[10480]_  | \new_[18077]_ ;
  assign \new_[8436]_  = ~\new_[12168]_  | ~\new_[12796]_ ;
  assign \new_[8437]_  = \new_[10322]_  & \new_[13993]_ ;
  assign \new_[8438]_  = ~\new_[10971]_  & ~\new_[13472]_ ;
  assign \new_[8439]_  = ~\new_[11887]_  | ~\new_[20084]_  | ~\new_[14213]_ ;
  assign \new_[8440]_  = ~\new_[13697]_  & ~\new_[10025]_ ;
  assign \new_[8441]_  = \new_[9871]_  | \new_[17472]_ ;
  assign \new_[8442]_  = ~\new_[15330]_  & ~\new_[10116]_ ;
  assign \new_[8443]_  = ~\new_[10282]_  & ~\new_[11346]_ ;
  assign \new_[8444]_  = ~\new_[15049]_  | ~\new_[9836]_  | ~\new_[15267]_ ;
  assign \new_[8445]_  = ~\new_[10181]_  | ~\new_[11366]_ ;
  assign \new_[8446]_  = ~\new_[9585]_ ;
  assign \new_[8447]_  = ~\new_[11841]_  | ~\new_[9880]_ ;
  assign \new_[8448]_  = ~\new_[11894]_  | ~\new_[10184]_ ;
  assign \new_[8449]_  = ~\new_[13684]_  | ~\new_[9876]_ ;
  assign \new_[8450]_  = ~\new_[14308]_  | ~\new_[9881]_ ;
  assign \new_[8451]_  = ~\new_[20558]_  & ~\new_[10542]_ ;
  assign \new_[8452]_  = ~\new_[9883]_  | ~\new_[12929]_ ;
  assign \new_[8453]_  = ~\new_[9587]_ ;
  assign \new_[8454]_  = ~\new_[9851]_  | ~\new_[20488]_ ;
  assign \new_[8455]_  = ~\new_[9589]_ ;
  assign \new_[8456]_  = ~\new_[10193]_  | ~\new_[21557]_ ;
  assign \new_[8457]_  = ~\new_[9889]_  | ~\new_[15379]_ ;
  assign \new_[8458]_  = ~\new_[20036]_  | ~\new_[11951]_  | ~\new_[11520]_ ;
  assign \new_[8459]_  = ~\new_[13199]_  | ~\new_[16215]_  | ~\new_[14677]_ ;
  assign \new_[8460]_  = ~\new_[9871]_  | ~\new_[12238]_ ;
  assign \new_[8461]_  = ~\new_[9592]_ ;
  assign \new_[8462]_  = \new_[9902]_  & \new_[11325]_ ;
  assign \new_[8463]_  = ~\new_[9901]_  | ~\new_[12918]_ ;
  assign \new_[8464]_  = ~\new_[10495]_  | ~\new_[15657]_ ;
  assign \new_[8465]_  = \new_[12221]_  & \new_[10617]_ ;
  assign \new_[8466]_  = ~\new_[10219]_  | ~\new_[14243]_ ;
  assign \new_[8467]_  = ~\new_[9907]_  | ~\new_[13726]_ ;
  assign \new_[8468]_  = ~\new_[11610]_  | ~\new_[11046]_  | ~\new_[16459]_ ;
  assign \new_[8469]_  = ~\new_[12694]_  | ~\new_[14247]_  | ~\new_[12691]_  | ~\new_[11849]_ ;
  assign \new_[8470]_  = \new_[10222]_  & \new_[12382]_ ;
  assign \new_[8471]_  = ~\new_[10225]_  | ~\new_[13367]_ ;
  assign \new_[8472]_  = ~\new_[10226]_  | ~\new_[12838]_ ;
  assign \new_[8473]_  = ~\new_[12384]_  | ~\new_[12168]_ ;
  assign \new_[8474]_  = \new_[10404]_  & \new_[9909]_ ;
  assign \new_[8475]_  = ~\new_[20161]_  | ~\new_[13709]_ ;
  assign \new_[8476]_  = ~\new_[9857]_  | ~\new_[13106]_ ;
  assign \new_[8477]_  = ~\new_[11004]_  | ~\new_[14677]_  | ~\new_[14523]_ ;
  assign \new_[8478]_  = ~\new_[12699]_  | ~\new_[15237]_  | ~\new_[14978]_  | ~\new_[14240]_ ;
  assign \new_[8479]_  = ~\new_[10125]_  | ~\new_[20680]_ ;
  assign \new_[8480]_  = ~\new_[12293]_  | ~\new_[10345]_ ;
  assign \new_[8481]_  = ~\new_[11023]_  | ~\new_[9915]_ ;
  assign \new_[8482]_  = ~\new_[15118]_  | ~\new_[13114]_  | ~\new_[12018]_  | ~\new_[12658]_ ;
  assign \new_[8483]_  = \new_[9917]_  & \new_[14295]_ ;
  assign \new_[8484]_  = ~\new_[13009]_  | ~\new_[10182]_ ;
  assign \new_[8485]_  = ~\new_[9920]_  | ~\new_[13859]_ ;
  assign \new_[8486]_  = ~\new_[10276]_  | ~\new_[18752]_ ;
  assign \new_[8487]_  = ~\new_[10411]_  & ~\new_[13032]_ ;
  assign \new_[8488]_  = ~\new_[13117]_  | ~\new_[9900]_ ;
  assign \new_[8489]_  = ~\new_[12918]_  | ~\new_[10403]_  | ~\new_[14126]_ ;
  assign \new_[8490]_  = ~\new_[10237]_  | ~\new_[11375]_ ;
  assign \new_[8491]_  = ~\new_[14068]_  | ~\new_[9922]_ ;
  assign \new_[8492]_  = ~\new_[15445]_  | ~\new_[12022]_  | ~\new_[13874]_ ;
  assign \new_[8493]_  = ~\new_[19687]_  & (~\new_[13125]_  | ~\new_[15425]_ );
  assign \new_[8494]_  = ~\new_[11005]_  | ~\new_[18070]_ ;
  assign \new_[8495]_  = ~\new_[11450]_  | ~\new_[18070]_ ;
  assign \new_[8496]_  = ~\new_[11777]_  | ~\new_[12881]_ ;
  assign \new_[8497]_  = ~\new_[11734]_  | ~\new_[10974]_ ;
  assign \new_[8498]_  = ~\new_[15384]_  | ~\new_[14196]_  | ~\new_[12455]_ ;
  assign \new_[8499]_  = ~\new_[11468]_  | ~\new_[16875]_ ;
  assign \new_[8500]_  = ~\new_[11454]_  | ~\new_[17472]_ ;
  assign \new_[8501]_  = ~\new_[20162]_  | ~\new_[17472]_ ;
  assign \new_[8502]_  = ~\new_[11271]_  | ~\new_[17801]_ ;
  assign \new_[8503]_  = ~\new_[11320]_  | ~\new_[17472]_ ;
  assign \new_[8504]_  = ~\new_[11351]_  | ~\new_[19079]_ ;
  assign \new_[8505]_  = ~\new_[21274]_  & (~\new_[14723]_  | ~\new_[14839]_ );
  assign \new_[8506]_  = \new_[12310]_  & \new_[11513]_ ;
  assign \new_[8507]_  = \new_[12287]_  & \new_[11493]_ ;
  assign n2713 = ~\new_[18775]_  | (~\new_[12428]_  & ~\new_[19723]_ );
  assign \new_[8509]_  = ~\new_[9625]_ ;
  assign \new_[8510]_  = ~\new_[11384]_  | ~\new_[18077]_ ;
  assign \new_[8511]_  = ~\new_[9626]_ ;
  assign \new_[8512]_  = \new_[11175]_  | \new_[16889]_ ;
  assign \new_[8513]_  = ~\new_[19233]_  & (~\new_[13146]_  | ~\new_[13902]_ );
  assign \new_[8514]_  = \new_[13484]_  & \new_[12229]_ ;
  assign \new_[8515]_  = \new_[12260]_  & \new_[11783]_ ;
  assign \new_[8516]_  = ~\new_[12387]_  | ~\new_[11649]_ ;
  assign \new_[8517]_  = ~\new_[11474]_  | ~\new_[17801]_ ;
  assign \new_[8518]_  = ~\new_[13654]_  & ~\new_[18077]_ ;
  assign \new_[8519]_  = ~\new_[19742]_  & (~\new_[12958]_  | ~\new_[16003]_ );
  assign \new_[8520]_  = ~\new_[9631]_ ;
  assign \new_[8521]_  = ~\new_[13060]_  & ~\new_[11009]_ ;
  assign \new_[8522]_  = ~\new_[11353]_  | ~\new_[12386]_ ;
  assign \new_[8523]_  = ~\new_[11800]_  | ~\new_[10994]_ ;
  assign \new_[8524]_  = ~\new_[11375]_  | ~\new_[12552]_ ;
  assign \new_[8525]_  = ~\new_[10997]_  | ~\new_[13166]_ ;
  assign \new_[8526]_  = \new_[12369]_  & \new_[11679]_ ;
  assign \new_[8527]_  = ~\new_[12379]_  | ~\new_[11242]_ ;
  assign \new_[8528]_  = ~\new_[9635]_ ;
  assign \new_[8529]_  = ~\new_[9636]_ ;
  assign \new_[8530]_  = ~\new_[16533]_  & ~\new_[21383]_ ;
  assign \new_[8531]_  = ~\new_[15870]_  & ~\new_[11330]_ ;
  assign \new_[8532]_  = \new_[12394]_  & \new_[12508]_ ;
  assign \new_[8533]_  = ~\new_[11347]_  | ~\new_[19217]_ ;
  assign \new_[8534]_  = ~\new_[9640]_ ;
  assign \new_[8535]_  = ~\new_[15108]_  | ~\new_[12418]_ ;
  assign \new_[8536]_  = ~\new_[11848]_  | ~\new_[12260]_ ;
  assign \new_[8537]_  = ~\new_[19249]_  & (~\new_[12746]_  | ~\new_[14198]_ );
  assign \new_[8538]_  = ~\new_[9643]_ ;
  assign \new_[8539]_  = ~\new_[14227]_  | ~\new_[10987]_ ;
  assign \new_[8540]_  = ~\new_[11282]_  | ~\new_[17723]_ ;
  assign \new_[8541]_  = ~\new_[20160]_  | ~\new_[12835]_ ;
  assign \new_[8542]_  = ~\new_[12417]_  & ~\new_[11213]_ ;
  assign \new_[8543]_  = ~\new_[9647]_ ;
  assign \new_[8544]_  = ~\new_[11312]_  | ~\new_[18280]_ ;
  assign \new_[8545]_  = ~\new_[14366]_  & (~\new_[12711]_  | ~\new_[19018]_ );
  assign \new_[8546]_  = ~\new_[12771]_  | ~\new_[20218]_  | ~\new_[14284]_ ;
  assign \new_[8547]_  = ~\new_[9650]_ ;
  assign \new_[8548]_  = ~\new_[12321]_  | ~\new_[11558]_ ;
  assign \new_[8549]_  = ~\new_[9653]_ ;
  assign \new_[8550]_  = ~\new_[12248]_  | ~\new_[11876]_ ;
  assign \new_[8551]_  = ~\new_[15540]_  & ~\new_[11288]_ ;
  assign \new_[8552]_  = ~\new_[15903]_  & ~\new_[11253]_ ;
  assign \new_[8553]_  = ~\new_[11362]_  | ~\new_[20100]_ ;
  assign \new_[8554]_  = \new_[11323]_  | \new_[19748]_ ;
  assign \new_[8555]_  = ~\new_[17003]_  | ~\new_[13091]_  | ~\new_[14225]_ ;
  assign \new_[8556]_  = ~\new_[17185]_  | ~\new_[21554]_  | ~\new_[15001]_ ;
  assign \new_[8557]_  = ~\new_[11017]_  | ~\new_[14926]_ ;
  assign \new_[8558]_  = ~\new_[11458]_  | ~\new_[19687]_ ;
  assign \new_[8559]_  = ~\new_[11957]_  | ~\new_[11016]_ ;
  assign \new_[8560]_  = ~\new_[20709]_  | ~\new_[19436]_ ;
  assign \new_[8561]_  = ~\new_[17189]_  & ~\new_[11347]_ ;
  assign \new_[8562]_  = ~\new_[13292]_  | ~\new_[11051]_  | ~\new_[14338]_ ;
  assign \new_[8563]_  = ~\new_[9664]_ ;
  assign \new_[8564]_  = \new_[11404]_  & \new_[19266]_ ;
  assign \new_[8565]_  = ~\new_[12397]_  | ~\new_[11599]_ ;
  assign \new_[8566]_  = ~\new_[10964]_  | ~\new_[15383]_ ;
  assign \new_[8567]_  = ~\new_[9668]_ ;
  assign \new_[8568]_  = ~\new_[12830]_  & ~\new_[10971]_ ;
  assign \new_[8569]_  = ~\new_[12881]_  | ~\new_[11095]_ ;
  assign \new_[8570]_  = ~\new_[11207]_  | ~\new_[13953]_ ;
  assign \new_[8571]_  = ~\new_[12294]_  | ~\new_[11518]_ ;
  assign \new_[8572]_  = ~\new_[11264]_  | ~\new_[19587]_ ;
  assign \new_[8573]_  = ~\new_[11056]_  | ~\new_[14202]_ ;
  assign \new_[8574]_  = \new_[11424]_  & \new_[19247]_ ;
  assign \new_[8575]_  = ~\new_[11056]_  | ~\new_[14136]_ ;
  assign \new_[8576]_  = ~\new_[11354]_  | ~\new_[18166]_ ;
  assign \new_[8577]_  = \new_[12815]_  & \new_[10927]_ ;
  assign \new_[8578]_  = ~\new_[14525]_  & ~\new_[11148]_ ;
  assign \new_[8579]_  = ~\new_[19553]_  & (~\new_[12983]_  | ~\new_[18396]_ );
  assign \new_[8580]_  = ~\new_[13971]_  | ~\new_[14371]_  | ~\new_[16407]_ ;
  assign \new_[8581]_  = ~\new_[11630]_  | ~\new_[12324]_ ;
  assign \new_[8582]_  = ~\new_[13652]_  | ~\new_[11666]_ ;
  assign \new_[8583]_  = ~\new_[11449]_  | ~\new_[18821]_ ;
  assign \new_[8584]_  = ~\new_[11427]_  & ~\new_[13815]_ ;
  assign \new_[8585]_  = \new_[12309]_  & \new_[10914]_ ;
  assign \new_[8586]_  = ~\new_[9675]_ ;
  assign \new_[8587]_  = ~\new_[11179]_  | ~\new_[19239]_ ;
  assign \new_[8588]_  = ~\new_[9676]_ ;
  assign \new_[8589]_  = ~\new_[16731]_  & ~\new_[11196]_ ;
  assign \new_[8590]_  = ~\new_[9677]_ ;
  assign \new_[8591]_  = ~\new_[11079]_  | ~\new_[18974]_ ;
  assign \new_[8592]_  = \new_[10964]_  & \new_[10976]_ ;
  assign \new_[8593]_  = ~\new_[15413]_  | ~\new_[15048]_  | ~\new_[15298]_ ;
  assign \new_[8594]_  = ~\new_[11368]_  | ~\new_[19507]_ ;
  assign \new_[8595]_  = ~\new_[11371]_  | ~\new_[19233]_ ;
  assign \new_[8596]_  = \new_[11463]_  | \new_[19072]_ ;
  assign \new_[8597]_  = ~\new_[9680]_ ;
  assign \new_[8598]_  = ~\new_[11113]_  | ~\new_[18965]_ ;
  assign \new_[8599]_  = ~\new_[9681]_ ;
  assign \new_[8600]_  = \new_[13546]_  & \new_[12233]_ ;
  assign \new_[8601]_  = ~\new_[11026]_  | ~\new_[19145]_ ;
  assign \new_[8602]_  = \new_[11376]_  | \new_[18087]_ ;
  assign \new_[8603]_  = ~\new_[11377]_  & ~\new_[15000]_ ;
  assign \new_[8604]_  = ~\new_[11563]_  & ~\new_[12381]_ ;
  assign \new_[8605]_  = ~\new_[16943]_  | ~\new_[21706]_  | ~\new_[14287]_ ;
  assign \new_[8606]_  = ~\new_[10939]_  | ~\new_[12211]_ ;
  assign \new_[8607]_  = \new_[11255]_  | \new_[19659]_ ;
  assign \new_[8608]_  = ~\new_[21026]_  | ~\new_[21631]_ ;
  assign \new_[8609]_  = ~\new_[11076]_  | ~\new_[13149]_ ;
  assign \new_[8610]_  = ~\new_[11465]_  & ~\new_[19224]_ ;
  assign \new_[8611]_  = ~\new_[9687]_ ;
  assign \new_[8612]_  = ~\new_[12298]_  & ~\new_[11628]_ ;
  assign \new_[8613]_  = ~\new_[11104]_  & ~\new_[12761]_ ;
  assign \new_[8614]_  = ~\new_[20422]_  | ~\new_[11780]_  | ~\new_[12763]_ ;
  assign \new_[8615]_  = ~\new_[9688]_ ;
  assign \new_[8616]_  = ~\new_[11379]_  & ~\new_[13799]_ ;
  assign \new_[8617]_  = ~\new_[15196]_  | ~\new_[11581]_  | ~\new_[16481]_ ;
  assign \new_[8618]_  = ~\new_[12325]_  & ~\new_[11686]_ ;
  assign \new_[8619]_  = ~\new_[9689]_ ;
  assign \new_[8620]_  = ~\new_[9692]_ ;
  assign \new_[8621]_  = ~\new_[11331]_  & ~\new_[11517]_ ;
  assign \new_[8622]_  = ~\new_[10770]_ ;
  assign \new_[8623]_  = ~\new_[9695]_ ;
  assign \new_[8624]_  = ~\new_[9697]_ ;
  assign \new_[8625]_  = ~\new_[17874]_  & (~\new_[13236]_  | ~\new_[16314]_ );
  assign \new_[8626]_  = ~\new_[11125]_  & (~\new_[18600]_  | ~\new_[18773]_ );
  assign \new_[8627]_  = ~\new_[9700]_ ;
  assign \new_[8628]_  = ~\new_[9702]_ ;
  assign \new_[8629]_  = ~\new_[11137]_  | ~\new_[19249]_ ;
  assign \new_[8630]_  = ~\new_[18863]_  & (~\new_[15433]_  | ~\new_[13780]_ );
  assign \new_[8631]_  = ~\new_[1878]_  | ~\new_[17488]_  | ~\new_[15035]_ ;
  assign \new_[8632]_  = \new_[11215]_  & \new_[13616]_ ;
  assign \new_[8633]_  = ~\new_[14949]_  | (~\new_[15342]_  & ~\new_[18414]_ );
  assign \new_[8634]_  = ~\new_[19204]_  & (~\new_[13311]_  | ~\new_[15455]_ );
  assign \new_[8635]_  = ~\new_[11131]_  | ~\new_[21115]_ ;
  assign \new_[8636]_  = ~\new_[9710]_ ;
  assign \new_[8637]_  = ~\new_[9712]_ ;
  assign \new_[8638]_  = ~\new_[9713]_ ;
  assign \new_[8639]_  = ~\new_[19445]_  | ~\new_[19228]_  | ~\new_[12679]_ ;
  assign \new_[8640]_  = ~\new_[9714]_ ;
  assign \new_[8641]_  = ~\new_[18344]_  | (~\new_[13325]_  & ~\new_[15438]_ );
  assign \new_[8642]_  = ~\new_[9715]_ ;
  assign \new_[8643]_  = ~\new_[9718]_ ;
  assign \new_[8644]_  = \new_[11422]_  & \new_[18187]_ ;
  assign \new_[8645]_  = \new_[11352]_  & \new_[19636]_ ;
  assign \new_[8646]_  = ~\new_[10956]_  | ~\new_[16125]_ ;
  assign \new_[8647]_  = ~\new_[15121]_  & (~\new_[21705]_  | ~\new_[19408]_ );
  assign \new_[8648]_  = ~\new_[12262]_  | ~\new_[10969]_ ;
  assign \new_[8649]_  = ~\new_[11214]_  | ~\new_[19587]_ ;
  assign \new_[8650]_  = ~\new_[921]_  & (~\new_[12624]_  | ~\new_[13299]_ );
  assign \new_[8651]_  = \new_[11338]_  & \new_[21638]_ ;
  assign \new_[8652]_  = ~\new_[9726]_ ;
  assign \new_[8653]_  = ~\new_[11232]_  | ~\new_[18825]_ ;
  assign \new_[8654]_  = ~\new_[9729]_ ;
  assign \new_[8655]_  = ~\new_[12468]_  | ~\new_[12647]_  | ~\new_[14629]_ ;
  assign \new_[8656]_  = ~\new_[9732]_ ;
  assign \new_[8657]_  = ~\new_[18632]_  | (~\new_[16279]_  & ~\new_[12531]_ );
  assign \new_[8658]_  = ~\new_[9733]_ ;
  assign \new_[8659]_  = ~\new_[11676]_  | ~\new_[10964]_ ;
  assign \new_[8660]_  = ~\new_[9734]_ ;
  assign \new_[8661]_  = ~\new_[9735]_ ;
  assign \new_[8662]_  = ~\new_[17358]_  & (~\new_[12234]_  | ~\new_[15849]_ );
  assign \new_[8663]_  = ~\new_[11937]_  | ~\new_[12247]_ ;
  assign \new_[8664]_  = ~\new_[12508]_  | ~\new_[13094]_  | ~\new_[13200]_ ;
  assign \new_[8665]_  = ~\new_[11942]_  | ~\new_[10997]_ ;
  assign \new_[8666]_  = ~\new_[19247]_  & (~\new_[15432]_  | ~\new_[12688]_ );
  assign \new_[8667]_  = ~\new_[21558]_  & (~\new_[13089]_  | ~\new_[15394]_ );
  assign \new_[8668]_  = ~\new_[11992]_  | ~\new_[12239]_ ;
  assign \new_[8669]_  = ~\new_[12720]_  | ~\new_[11056]_ ;
  assign \new_[8670]_  = ~\new_[15767]_  & (~\new_[21670]_  | ~\new_[13714]_ );
  assign \new_[8671]_  = ~\new_[11138]_  | ~\new_[14951]_ ;
  assign \new_[8672]_  = ~\new_[11139]_  | ~\new_[19357]_ ;
  assign \new_[8673]_  = ~\new_[13785]_  | ~\new_[15237]_  | ~\new_[13083]_ ;
  assign \new_[8674]_  = ~\new_[17689]_  & (~\new_[15403]_  | ~\new_[12584]_ );
  assign \new_[8675]_  = ~\new_[11299]_  | ~\new_[21638]_ ;
  assign \new_[8676]_  = ~\new_[922]_  & (~\new_[12595]_  | ~\new_[13015]_ );
  assign \new_[8677]_  = ~\new_[11157]_  & ~\new_[12905]_ ;
  assign \new_[8678]_  = ~\new_[17979]_  & (~\new_[15841]_  | ~\new_[14806]_ );
  assign \new_[8679]_  = ~\new_[9750]_ ;
  assign \new_[8680]_  = ~\new_[9753]_ ;
  assign \new_[8681]_  = ~\new_[11341]_  | ~\new_[18957]_ ;
  assign \new_[8682]_  = ~\new_[11284]_  | ~\new_[18278]_ ;
  assign \new_[8683]_  = ~\new_[11200]_  | ~\new_[18909]_ ;
  assign \new_[8684]_  = ~\new_[9755]_ ;
  assign \new_[8685]_  = ~\new_[15660]_  | ~\new_[14293]_  | ~\new_[17301]_  | ~\new_[14150]_ ;
  assign \new_[8686]_  = ~\new_[9756]_ ;
  assign \new_[8687]_  = ~\new_[18066]_  & (~\new_[15048]_  | ~\new_[13781]_ );
  assign \new_[8688]_  = ~\new_[11835]_  | ~\new_[12206]_ ;
  assign \new_[8689]_  = ~\new_[9757]_ ;
  assign \new_[8690]_  = ~\new_[14346]_  | ~\new_[13737]_  | ~\new_[12584]_ ;
  assign \new_[8691]_  = ~\new_[9758]_ ;
  assign \new_[8692]_  = ~\new_[9746]_ ;
  assign \new_[8693]_  = ~\new_[9761]_ ;
  assign \new_[8694]_  = ~\new_[11216]_  & (~\new_[15477]_  | ~\new_[19408]_ );
  assign \new_[8695]_  = ~\new_[9764]_ ;
  assign \new_[8696]_  = ~\new_[11358]_  | ~\new_[19088]_ ;
  assign \new_[8697]_  = ~\new_[11389]_  | ~\new_[18873]_ ;
  assign \new_[8698]_  = ~\new_[11337]_  | ~\new_[17983]_ ;
  assign \new_[8699]_  = ~\new_[9769]_ ;
  assign \new_[8700]_  = ~\new_[9771]_ ;
  assign \new_[8701]_  = ~\new_[11108]_  | ~\new_[14951]_ ;
  assign \new_[8702]_  = ~\new_[11766]_  | ~\new_[13584]_ ;
  assign \new_[8703]_  = ~\new_[13048]_  | ~\new_[11016]_ ;
  assign \new_[8704]_  = \new_[11393]_  & \new_[17925]_ ;
  assign \new_[8705]_  = \new_[11394]_  & \new_[17749]_ ;
  assign \new_[8706]_  = ~\new_[11652]_  | ~\new_[12418]_ ;
  assign \new_[8707]_  = ~\new_[10946]_  | ~\new_[11793]_ ;
  assign \new_[8708]_  = ~\new_[18154]_  | (~\new_[17711]_  & ~\new_[13151]_ );
  assign \new_[8709]_  = ~\new_[18380]_  | (~\new_[17674]_  & ~\new_[13189]_ );
  assign \new_[8710]_  = ~\new_[18786]_  | (~\new_[17854]_  & ~\new_[13196]_ );
  assign \new_[8711]_  = ~\new_[11118]_  & (~\new_[18223]_  | ~\new_[15892]_ );
  assign \new_[8712]_  = ~\new_[11156]_  & (~\new_[18839]_  | ~\new_[18262]_ );
  assign \new_[8713]_  = ~\new_[13277]_  & ~\new_[11143]_ ;
  assign \new_[8714]_  = ~\new_[11241]_  | ~\new_[18752]_ ;
  assign \new_[8715]_  = ~\new_[11372]_  & (~\new_[18069]_  | ~\new_[17488]_ );
  assign \new_[8716]_  = \new_[14798]_  ? \new_[19687]_  : \new_[13332]_ ;
  assign \new_[8717]_  = \new_[14328]_  ? \new_[18965]_  : \new_[13256]_ ;
  assign \new_[8718]_  = \new_[12967]_  ? \new_[19553]_  : \new_[16204]_ ;
  assign \new_[8719]_  = ~\new_[12353]_  & (~\new_[12830]_  | ~\new_[18998]_ );
  assign \new_[8720]_  = ~\new_[11296]_  & (~\new_[13060]_  | ~\new_[21634]_ );
  assign \new_[8721]_  = ~\new_[11892]_  | (~\new_[12839]_  & ~\new_[18794]_ );
  assign \new_[8722]_  = ~\new_[11472]_  & (~\new_[18010]_  | ~\new_[17488]_ );
  assign \new_[8723]_  = ~\new_[18341]_  | (~\new_[13328]_  & ~\new_[15443]_ );
  assign \new_[8724]_  = ~\new_[12013]_  | (~\new_[13122]_  & ~\new_[20490]_ );
  assign \new_[8725]_  = ~\new_[11470]_  & (~\new_[18578]_  | ~\new_[18262]_ );
  assign \new_[8726]_  = ~\new_[10945]_  & (~\new_[18332]_  | ~\new_[18206]_ );
  assign \new_[8727]_  = ~\new_[10953]_  & (~\new_[21682]_  | ~\new_[18402]_ );
  assign \new_[8728]_  = ~\new_[10948]_  | ~\new_[13497]_ ;
  assign \new_[8729]_  = ~\new_[11135]_  & (~\new_[18003]_  | ~\new_[18750]_ );
  assign \new_[8730]_  = (~\new_[17855]_  | ~\new_[18849]_ ) & (~\new_[15569]_  | ~\new_[19319]_ );
  assign \new_[8731]_  = ~\new_[12571]_  & (~\new_[12829]_  | ~\new_[18778]_ );
  assign \new_[8732]_  = ~\new_[13985]_  & (~\new_[12155]_  | ~\new_[18046]_ );
  assign \new_[8733]_  = ~\new_[12787]_  & (~\new_[13016]_  | ~\new_[18569]_ );
  assign \new_[8734]_  = \new_[14399]_  & \new_[11819]_ ;
  assign \new_[8735]_  = \new_[11959]_  & \new_[19366]_ ;
  assign \new_[8736]_  = ~\new_[11950]_  & (~\new_[14512]_  | ~\new_[17461]_ );
  assign \new_[8737]_  = \new_[12062]_  & \new_[14848]_ ;
  assign \new_[8738]_  = \new_[18821]_  | \new_[11828]_ ;
  assign \new_[8739]_  = \new_[11586]_  | \new_[19261]_ ;
  assign \new_[8740]_  = ~\new_[9802]_ ;
  assign \new_[8741]_  = ~\new_[11948]_  & ~\new_[19088]_ ;
  assign \new_[8742]_  = ~\new_[10850]_  | ~\new_[18166]_ ;
  assign \new_[8743]_  = \new_[11839]_  & \new_[19625]_ ;
  assign \new_[8744]_  = ~\new_[11717]_  | ~\new_[21689]_ ;
  assign \new_[8745]_  = ~\new_[14375]_  & ~\new_[19474]_ ;
  assign \new_[8746]_  = ~\new_[9819]_ ;
  assign \new_[8747]_  = ~\new_[9825]_ ;
  assign \new_[8748]_  = ~\new_[9828]_ ;
  assign \new_[8749]_  = \new_[11870]_  | \new_[19547]_ ;
  assign \new_[8750]_  = ~\new_[11963]_  | ~\new_[19156]_ ;
  assign \new_[8751]_  = ~\new_[14424]_  & ~\new_[19269]_ ;
  assign \new_[8752]_  = ~\new_[10850]_  | ~\new_[19612]_ ;
  assign \new_[8753]_  = ~\new_[9835]_ ;
  assign \new_[8754]_  = ~\new_[9840]_ ;
  assign \new_[8755]_  = ~\new_[11883]_  | ~\new_[19021]_ ;
  assign \new_[8756]_  = ~\new_[11815]_  | ~\new_[18187]_ ;
  assign \new_[8757]_  = ~\new_[21635]_  & ~\new_[13897]_ ;
  assign \new_[8758]_  = ~\new_[9854]_ ;
  assign \new_[8759]_  = ~\new_[19592]_  & ~\new_[11560]_ ;
  assign \new_[8760]_  = ~\new_[9855]_ ;
  assign \new_[8761]_  = \new_[11956]_  | \new_[19161]_ ;
  assign \new_[8762]_  = ~\new_[19204]_  | ~\new_[11717]_ ;
  assign \new_[8763]_  = ~\new_[9868]_ ;
  assign \new_[8764]_  = \new_[16041]_  | \new_[21515]_  | \new_[18427]_  | \new_[18810]_ ;
  assign \new_[8765]_  = ~\new_[9877]_ ;
  assign \new_[8766]_  = ~\new_[11887]_  & ~\new_[19102]_ ;
  assign \new_[8767]_  = ~\new_[19088]_  & ~\new_[11571]_ ;
  assign \new_[8768]_  = ~\new_[9884]_ ;
  assign \new_[8769]_  = ~\new_[11877]_  & ~\new_[18046]_ ;
  assign \new_[8770]_  = ~\new_[9886]_ ;
  assign \new_[8771]_  = ~\new_[9888]_ ;
  assign \new_[8772]_  = ~\new_[9891]_ ;
  assign \new_[8773]_  = ~\new_[9899]_ ;
  assign \new_[8774]_  = ~\new_[14718]_  | ~\new_[21558]_  | ~\new_[18275]_ ;
  assign \new_[8775]_  = \new_[11594]_  | \new_[21562]_ ;
  assign \new_[8776]_  = ~\new_[9909]_ ;
  assign \new_[8777]_  = ~\new_[9912]_ ;
  assign \new_[8778]_  = ~\new_[11843]_  & ~\new_[19018]_ ;
  assign \new_[8779]_  = \new_[11961]_  | \new_[19587]_ ;
  assign \new_[8780]_  = ~\new_[9919]_ ;
  assign \new_[8781]_  = ~\new_[20221]_  & ~\new_[21563]_ ;
  assign \new_[8782]_  = ~\new_[11799]_  | ~\new_[18941]_ ;
  assign \new_[8783]_  = ~\new_[9925]_ ;
  assign \new_[8784]_  = ~\new_[11747]_  | ~\new_[19107]_ ;
  assign \new_[8785]_  = ~\new_[9928]_ ;
  assign \new_[8786]_  = ~\new_[9931]_ ;
  assign \new_[8787]_  = ~\new_[9933]_ ;
  assign \new_[8788]_  = ~\new_[9934]_ ;
  assign \new_[8789]_  = ~\new_[9934]_ ;
  assign \new_[8790]_  = ~\new_[13873]_  & ~\new_[19202]_ ;
  assign \new_[8791]_  = ~\new_[11960]_  | ~\new_[21395]_ ;
  assign \new_[8792]_  = ~\new_[9946]_ ;
  assign \new_[8793]_  = ~\new_[9947]_ ;
  assign \new_[8794]_  = ~\new_[9950]_ ;
  assign \new_[8795]_  = ~\new_[11587]_  | ~\new_[21629]_ ;
  assign \new_[8796]_  = \new_[16041]_  | \new_[21515]_  | \new_[21115]_  | \new_[18605]_ ;
  assign \new_[8797]_  = ~\new_[11536]_  & ~\new_[19619]_ ;
  assign \new_[8798]_  = ~\new_[21563]_  & ~\new_[11591]_ ;
  assign \new_[8799]_  = \new_[11949]_  | \new_[18542]_ ;
  assign \new_[8800]_  = ~\new_[9957]_ ;
  assign \new_[8801]_  = ~\new_[9967]_ ;
  assign \new_[8802]_  = ~\new_[11683]_  & ~\new_[19436]_ ;
  assign \new_[8803]_  = ~\new_[11991]_  & ~\new_[19266]_ ;
  assign \new_[8804]_  = ~\new_[12099]_  | ~\new_[20845]_ ;
  assign \new_[8805]_  = ~\new_[11963]_  | ~\new_[18965]_ ;
  assign \new_[8806]_  = ~\new_[11757]_  & ~\new_[19261]_ ;
  assign \new_[8807]_  = ~\new_[11513]_  & ~\new_[19079]_ ;
  assign \new_[8808]_  = ~\new_[13996]_  & ~\new_[18692]_ ;
  assign \new_[8809]_  = ~\new_[9979]_ ;
  assign \new_[8810]_  = ~\new_[9982]_ ;
  assign \new_[8811]_  = ~\new_[21550]_  | ~\new_[19612]_  | ~\new_[17626]_ ;
  assign \new_[8812]_  = ~\new_[11873]_  | ~\new_[19592]_ ;
  assign \new_[8813]_  = ~\new_[11847]_  & ~\new_[19156]_ ;
  assign \new_[8814]_  = ~\new_[11935]_  | ~\new_[19446]_ ;
  assign \new_[8815]_  = ~\new_[11558]_  & ~\new_[19659]_ ;
  assign \new_[8816]_  = ~\new_[11596]_  | ~\new_[14951]_ ;
  assign \new_[8817]_  = ~\new_[9996]_ ;
  assign \new_[8818]_  = ~\new_[11679]_  & ~\new_[18627]_ ;
  assign \new_[8819]_  = \new_[11895]_  | \new_[19015]_ ;
  assign \new_[8820]_  = ~\new_[11493]_  & ~\new_[19215]_ ;
  assign \new_[8821]_  = ~\new_[10004]_ ;
  assign \new_[8822]_  = ~\new_[18734]_  & ~\new_[11520]_ ;
  assign \new_[8823]_  = ~\new_[11660]_  | ~\new_[16312]_ ;
  assign \new_[8824]_  = ~\new_[10009]_ ;
  assign \new_[8825]_  = ~\new_[10011]_ ;
  assign \new_[8826]_  = \new_[11963]_  | \new_[16873]_ ;
  assign \new_[8827]_  = ~\new_[18077]_  & ~\new_[14677]_ ;
  assign \new_[8828]_  = \new_[11808]_  & \new_[13149]_ ;
  assign \new_[8829]_  = \new_[13715]_  | \new_[17598]_ ;
  assign \new_[8830]_  = ~\new_[11569]_  & ~\new_[18423]_ ;
  assign \new_[8831]_  = ~\new_[13490]_  | ~\new_[12560]_ ;
  assign \new_[8832]_  = \new_[13793]_  | \new_[19064]_ ;
  assign \new_[8833]_  = ~\new_[15485]_  | ~\new_[11512]_ ;
  assign \new_[8834]_  = ~\new_[18117]_  & ~\new_[13846]_ ;
  assign \new_[8835]_  = ~\new_[10029]_ ;
  assign \new_[8836]_  = ~\new_[11756]_  | ~\new_[12566]_ ;
  assign \new_[8837]_  = ~\new_[10031]_ ;
  assign \new_[8838]_  = ~\new_[11507]_  | ~\new_[14304]_ ;
  assign \new_[8839]_  = ~\new_[10032]_ ;
  assign \new_[8840]_  = ~\new_[11529]_  | ~\new_[21686]_ ;
  assign \new_[8841]_  = ~\new_[15497]_  | ~\new_[14414]_ ;
  assign \new_[8842]_  = \new_[13800]_  | \new_[19156]_ ;
  assign \new_[8843]_  = ~\new_[14155]_  & ~\new_[18569]_ ;
  assign \new_[8844]_  = ~\new_[11600]_  | ~\new_[13636]_ ;
  assign \new_[8845]_  = \new_[13727]_  | \new_[19079]_ ;
  assign \new_[8846]_  = ~\new_[14155]_  | ~\new_[13746]_ ;
  assign \new_[8847]_  = ~\new_[11496]_  | ~\new_[17544]_ ;
  assign \new_[8848]_  = ~\new_[11661]_  & ~\new_[11508]_ ;
  assign \new_[8849]_  = ~\new_[12506]_  | ~\new_[17818]_ ;
  assign \new_[8850]_  = ~\new_[20825]_  | ~\new_[14212]_ ;
  assign \new_[8851]_  = ~\new_[10041]_ ;
  assign \new_[8852]_  = ~\new_[19261]_  & ~\new_[13816]_ ;
  assign \new_[8853]_  = ~\new_[15838]_  | ~\new_[14951]_ ;
  assign \new_[8854]_  = ~\new_[11532]_  & ~\new_[15164]_ ;
  assign \new_[8855]_  = ~\new_[10047]_ ;
  assign \new_[8856]_  = ~\new_[10049]_ ;
  assign \new_[8857]_  = ~\new_[14580]_  | ~\new_[14375]_ ;
  assign \new_[8858]_  = ~\new_[11706]_  | ~\new_[17373]_ ;
  assign \new_[8859]_  = \new_[11517]_  | \new_[15353]_ ;
  assign \new_[8860]_  = ~\new_[16151]_  | ~\new_[20433]_ ;
  assign \new_[8861]_  = ~\new_[19021]_  | (~\new_[13381]_  & ~\new_[14736]_ );
  assign \new_[8862]_  = \new_[13368]_  | \new_[11717]_ ;
  assign \new_[8863]_  = \new_[12060]_  & \new_[19013]_ ;
  assign \new_[8864]_  = \new_[11710]_  | \new_[21686]_ ;
  assign \new_[8865]_  = ~\new_[15802]_  | ~\new_[11808]_ ;
  assign \new_[8866]_  = ~\new_[13820]_  | ~\new_[15253]_ ;
  assign \new_[8867]_  = \new_[12526]_  & \new_[13724]_ ;
  assign \new_[8868]_  = ~\new_[14290]_  & ~\new_[14094]_ ;
  assign \new_[8869]_  = ~\new_[13602]_  & ~\new_[15874]_ ;
  assign \new_[8870]_  = ~\new_[13204]_  | ~\new_[11863]_ ;
  assign \new_[8871]_  = ~\new_[11775]_  | ~\new_[18941]_ ;
  assign \new_[8872]_  = ~\new_[11527]_  | ~\new_[11731]_ ;
  assign \new_[8873]_  = \new_[11630]_  | \new_[18709]_ ;
  assign \new_[8874]_  = \new_[13979]_  | \new_[19156]_ ;
  assign \new_[8875]_  = ~\new_[12028]_  | ~\new_[16899]_ ;
  assign \new_[8876]_  = ~\new_[14058]_  & ~\new_[18621]_ ;
  assign \new_[8877]_  = \new_[13803]_  | \new_[19156]_ ;
  assign \new_[8878]_  = ~\new_[15367]_  | ~\new_[11782]_ ;
  assign \new_[8879]_  = ~\new_[18657]_  & ~\new_[11703]_ ;
  assign \new_[8880]_  = \new_[13540]_  | \new_[11526]_ ;
  assign \new_[8881]_  = ~\new_[11845]_  | ~\new_[21115]_ ;
  assign \new_[8882]_  = ~\new_[10855]_  | ~\new_[13782]_ ;
  assign \new_[8883]_  = ~\new_[11771]_  & ~\new_[12611]_ ;
  assign \new_[8884]_  = ~\new_[10101]_ ;
  assign \new_[8885]_  = ~\new_[14288]_  & (~\new_[16673]_  | ~\new_[17521]_ );
  assign \new_[8886]_  = ~\new_[16127]_  | ~\new_[21706]_ ;
  assign \new_[8887]_  = ~\new_[13763]_  & ~\new_[18209]_ ;
  assign \new_[8888]_  = \new_[15671]_  & \new_[11828]_ ;
  assign \new_[8889]_  = ~\new_[10107]_ ;
  assign \new_[8890]_  = ~\new_[20232]_  & ~\new_[19015]_ ;
  assign \new_[8891]_  = ~\new_[10111]_ ;
  assign \new_[8892]_  = \new_[13729]_  | \new_[18938]_ ;
  assign \new_[8893]_  = ~\new_[21043]_  | ~\new_[17758]_ ;
  assign \new_[8894]_  = \new_[14229]_  | \new_[18692]_ ;
  assign \new_[8895]_  = \new_[11765]_  & \new_[16619]_ ;
  assign \new_[8896]_  = \new_[13590]_  | \new_[18077]_ ;
  assign \new_[8897]_  = ~\new_[15016]_  | ~\new_[11684]_ ;
  assign \new_[8898]_  = ~\new_[11636]_  | ~\new_[20388]_ ;
  assign \new_[8899]_  = \new_[18187]_  | \new_[14117]_ ;
  assign \new_[8900]_  = \new_[11983]_  | \new_[18650]_ ;
  assign \new_[8901]_  = \new_[11903]_  | \new_[21563]_ ;
  assign \new_[8902]_  = ~\new_[10709]_ ;
  assign \new_[8903]_  = \new_[13668]_  & \new_[19088]_ ;
  assign \new_[8904]_  = ~\new_[12042]_  | ~\new_[13796]_ ;
  assign \new_[8905]_  = ~\new_[13873]_  | ~\new_[11562]_ ;
  assign \new_[8906]_  = ~\new_[13237]_  | ~\new_[11996]_ ;
  assign \new_[8907]_  = ~\new_[18731]_  & ~\new_[11325]_ ;
  assign \new_[8908]_  = ~\new_[12042]_  & ~\new_[16879]_ ;
  assign \new_[8909]_  = ~\new_[20218]_  | ~\new_[11595]_ ;
  assign \new_[8910]_  = ~\new_[16837]_  | ~\new_[11876]_ ;
  assign \new_[8911]_  = ~\new_[10131]_ ;
  assign \new_[8912]_  = \new_[13669]_  | \new_[18361]_ ;
  assign \new_[8913]_  = ~\new_[14313]_  | ~\new_[15830]_ ;
  assign \new_[8914]_  = ~\new_[13286]_  & ~\new_[12795]_ ;
  assign \new_[8915]_  = ~\new_[10136]_ ;
  assign \new_[8916]_  = ~\new_[11630]_  & ~\new_[17926]_ ;
  assign \new_[8917]_  = ~\new_[11799]_  | ~\new_[19127]_ ;
  assign \new_[8918]_  = ~\new_[11514]_  & ~\new_[15265]_ ;
  assign \new_[8919]_  = ~\new_[11619]_  | ~\new_[11507]_ ;
  assign \new_[8920]_  = ~\new_[11589]_  | ~\new_[14951]_ ;
  assign \new_[8921]_  = ~\new_[14412]_  | ~\new_[13852]_ ;
  assign \new_[8922]_  = ~\new_[15830]_  & ~\new_[18111]_ ;
  assign \new_[8923]_  = ~\new_[10148]_ ;
  assign \new_[8924]_  = ~\new_[11932]_  | ~\new_[14997]_ ;
  assign \new_[8925]_  = \new_[11586]_  & \new_[11710]_ ;
  assign \new_[8926]_  = ~\new_[11854]_  | ~\new_[11679]_ ;
  assign \new_[8927]_  = ~\new_[10154]_ ;
  assign \new_[8928]_  = \new_[13967]_  | \new_[19203]_ ;
  assign \new_[8929]_  = \new_[11492]_  & \new_[15094]_ ;
  assign \new_[8930]_  = ~\new_[13775]_  | ~\new_[16079]_ ;
  assign \new_[8931]_  = ~\new_[11575]_  | ~\new_[14897]_ ;
  assign \new_[8932]_  = ~\new_[16371]_  | ~\new_[11537]_ ;
  assign \new_[8933]_  = ~\new_[17366]_  | ~\new_[11875]_ ;
  assign \new_[8934]_  = ~\new_[11092]_  | ~\new_[19204]_ ;
  assign \new_[8935]_  = ~\new_[15030]_  & ~\new_[14397]_ ;
  assign \new_[8936]_  = ~\new_[11161]_  | ~\new_[13695]_ ;
  assign \new_[8937]_  = \new_[14275]_  | \new_[18747]_ ;
  assign \new_[8938]_  = ~\new_[14598]_  | ~\new_[11512]_ ;
  assign \new_[8939]_  = ~\new_[14183]_  | ~\new_[12027]_ ;
  assign \new_[8940]_  = \new_[12049]_  & \new_[19028]_ ;
  assign \new_[8941]_  = ~\new_[11619]_  | ~\new_[13731]_ ;
  assign \new_[8942]_  = ~\new_[11557]_  & ~\new_[17112]_ ;
  assign \new_[8943]_  = ~\new_[14170]_  | ~\new_[11975]_ ;
  assign \new_[8944]_  = ~\new_[11893]_  | ~\new_[17780]_ ;
  assign \new_[8945]_  = ~\new_[15364]_  & ~\new_[11927]_ ;
  assign \new_[8946]_  = \new_[13724]_  | \new_[19095]_ ;
  assign \new_[8947]_  = \new_[11492]_  & \new_[13793]_ ;
  assign \new_[8948]_  = \new_[11593]_  | \new_[18325]_ ;
  assign \new_[8949]_  = \new_[11594]_  & \new_[13859]_ ;
  assign \new_[8950]_  = ~\new_[11811]_  | ~\new_[17307]_ ;
  assign \new_[8951]_  = ~\new_[15277]_  | ~\new_[12018]_ ;
  assign \new_[8952]_  = ~\new_[13706]_  | ~\new_[13863]_ ;
  assign \new_[8953]_  = ~\new_[11592]_  & ~\new_[11726]_ ;
  assign \new_[8954]_  = ~\new_[14213]_  | ~\new_[11493]_ ;
  assign \new_[8955]_  = ~\new_[13543]_  | ~\new_[12555]_ ;
  assign \new_[8956]_  = ~\new_[15276]_  & ~\new_[14400]_ ;
  assign \new_[8957]_  = ~\new_[10188]_ ;
  assign \new_[8958]_  = ~\new_[11619]_  | ~\new_[15120]_ ;
  assign \new_[8959]_  = ~\new_[13077]_  | ~\new_[11903]_ ;
  assign \new_[8960]_  = \new_[12727]_  & \new_[14208]_ ;
  assign \new_[8961]_  = ~\new_[11742]_  | ~\new_[21558]_ ;
  assign \new_[8962]_  = ~\new_[17011]_  | ~\new_[14548]_  | ~\new_[16084]_  | ~\new_[17503]_ ;
  assign \new_[8963]_  = \new_[11510]_  | \new_[19028]_ ;
  assign \new_[8964]_  = ~\new_[13413]_  | ~\new_[14346]_ ;
  assign \new_[8965]_  = ~\new_[13083]_  | ~\new_[11780]_ ;
  assign \new_[8966]_  = ~\new_[14590]_  | ~\new_[11869]_ ;
  assign \new_[8967]_  = ~\new_[11581]_  | ~\new_[14014]_ ;
  assign \new_[8968]_  = ~\new_[21330]_  | ~\new_[14207]_ ;
  assign \new_[8969]_  = \new_[18335]_  | \new_[14225]_ ;
  assign \new_[8970]_  = ~\new_[10200]_ ;
  assign \new_[8971]_  = ~\new_[10202]_ ;
  assign \new_[8972]_  = ~\new_[15935]_  | ~\new_[11607]_ ;
  assign \new_[8973]_  = ~\new_[10205]_ ;
  assign \new_[8974]_  = ~\new_[19702]_  | ~\new_[14188]_  | ~\new_[18124]_ ;
  assign \new_[8975]_  = ~\new_[11626]_  & ~\new_[15540]_ ;
  assign \new_[8976]_  = \new_[11669]_  & \new_[15592]_ ;
  assign \new_[8977]_  = \new_[11650]_  & \new_[11569]_ ;
  assign \new_[8978]_  = ~\new_[12405]_  | ~\new_[21173]_ ;
  assign \new_[8979]_  = ~\new_[11778]_  & ~\new_[16294]_ ;
  assign \new_[8980]_  = ~\new_[10214]_ ;
  assign \new_[8981]_  = ~\new_[11694]_  | ~\new_[19115]_ ;
  assign \new_[8982]_  = \new_[12046]_  & \new_[21562]_ ;
  assign \new_[8983]_  = ~\new_[19462]_  & ~\new_[11811]_ ;
  assign \new_[8984]_  = ~\new_[18734]_  & ~\new_[13755]_ ;
  assign \new_[8985]_  = \new_[13358]_  & \new_[13860]_ ;
  assign \new_[8986]_  = ~\new_[11623]_  | ~\new_[14052]_ ;
  assign \new_[8987]_  = \new_[13821]_  | \new_[19202]_ ;
  assign \new_[8988]_  = ~\new_[13874]_  | ~\new_[11610]_ ;
  assign \new_[8989]_  = ~\new_[16128]_  | ~\new_[11528]_ ;
  assign \new_[8990]_  = ~\new_[17472]_  & ~\new_[13993]_ ;
  assign \new_[8991]_  = ~\new_[14829]_  | ~\new_[11980]_ ;
  assign \new_[8992]_  = ~\new_[11803]_  | ~\new_[17697]_ ;
  assign \new_[8993]_  = ~\new_[18914]_  & ~\new_[14664]_ ;
  assign \new_[8994]_  = ~\new_[13676]_  | ~\new_[17457]_ ;
  assign \new_[8995]_  = ~\new_[13993]_  | ~\new_[13868]_ ;
  assign \new_[8996]_  = ~\new_[18626]_  & ~\new_[11850]_ ;
  assign \new_[8997]_  = ~\new_[10230]_ ;
  assign \new_[8998]_  = ~\new_[14434]_  & ~\new_[19436]_ ;
  assign \new_[8999]_  = ~\new_[11553]_  | ~\new_[16195]_ ;
  assign \new_[9000]_  = ~\new_[12014]_  | ~\new_[11683]_ ;
  assign \new_[9001]_  = ~\new_[11659]_  | ~\new_[17939]_ ;
  assign \new_[9002]_  = ~\new_[10232]_ ;
  assign \new_[9003]_  = ~\new_[11767]_  | ~\new_[18621]_ ;
  assign \new_[9004]_  = ~\new_[18847]_  & ~\new_[14304]_ ;
  assign \new_[9005]_  = ~\new_[12610]_  & ~\new_[11632]_ ;
  assign \new_[9006]_  = ~\new_[11541]_  | ~\new_[18605]_ ;
  assign \new_[9007]_  = ~\new_[15017]_  & ~\new_[19156]_ ;
  assign \new_[9008]_  = ~\new_[13007]_  & ~\new_[14558]_ ;
  assign \new_[9009]_  = ~\new_[13638]_  | ~\new_[11595]_ ;
  assign \new_[9010]_  = ~\new_[21043]_  | ~\new_[18693]_ ;
  assign \new_[9011]_  = ~\new_[21164]_  & ~\new_[18973]_ ;
  assign \new_[9012]_  = ~\new_[15309]_  | ~\new_[11535]_ ;
  assign \new_[9013]_  = ~\new_[11889]_  & ~\new_[13369]_ ;
  assign \new_[9014]_  = ~\new_[13859]_  & ~\new_[18747]_ ;
  assign \new_[9015]_  = ~\new_[13089]_  | ~\new_[11594]_ ;
  assign \new_[9016]_  = ~\new_[20715]_  | ~\new_[19436]_ ;
  assign \new_[9017]_  = ~\new_[16485]_  | ~\new_[14379]_ ;
  assign \new_[9018]_  = ~\new_[13547]_  & ~\new_[19072]_ ;
  assign \new_[9019]_  = ~\new_[13748]_  & ~\new_[11625]_ ;
  assign \new_[9020]_  = ~\new_[11911]_  | ~\new_[20100]_ ;
  assign \new_[9021]_  = ~\new_[12935]_  | ~\new_[11807]_ ;
  assign \new_[9022]_  = ~\new_[14511]_  | ~\new_[14609]_ ;
  assign \new_[9023]_  = \new_[11535]_  | \new_[19151]_ ;
  assign \new_[9024]_  = ~\new_[15237]_  | ~\new_[11581]_ ;
  assign \new_[9025]_  = \new_[12051]_  & \new_[18778]_ ;
  assign \new_[9026]_  = ~\new_[11357]_  & ~\new_[12576]_ ;
  assign \new_[9027]_  = ~\new_[11882]_  | ~\new_[17710]_ ;
  assign \new_[9028]_  = ~\new_[13749]_  | ~\new_[15767]_ ;
  assign \new_[9029]_  = ~\new_[14434]_  | ~\new_[12494]_ ;
  assign \new_[9030]_  = \new_[11677]_  & \new_[11600]_ ;
  assign \new_[9031]_  = ~\new_[14714]_  | ~\new_[14159]_ ;
  assign \new_[9032]_  = ~\new_[12562]_  & ~\new_[11976]_ ;
  assign \new_[9033]_  = ~\new_[15726]_  | ~\new_[13863]_ ;
  assign \new_[9034]_  = ~\new_[16802]_  | ~\new_[14121]_ ;
  assign \new_[9035]_  = \new_[11868]_  & \new_[16595]_ ;
  assign \new_[9036]_  = \new_[17256]_  & \new_[11955]_ ;
  assign \new_[9037]_  = ~\new_[21329]_  & ~\new_[18542]_ ;
  assign \new_[9038]_  = ~\new_[11878]_  | ~\new_[18569]_ ;
  assign \new_[9039]_  = ~\new_[13236]_  | ~\new_[11513]_ ;
  assign \new_[9040]_  = ~\new_[11646]_  | ~\new_[16150]_ ;
  assign \new_[9041]_  = ~\new_[13478]_  | ~\new_[11522]_ ;
  assign \new_[9042]_  = ~\new_[11665]_  & ~\new_[15426]_ ;
  assign \new_[9043]_  = ~\new_[12076]_  & (~\new_[18609]_  | ~\new_[18901]_ );
  assign \new_[9044]_  = ~\new_[10256]_ ;
  assign \new_[9045]_  = \new_[18490]_  | \new_[11940]_ ;
  assign \new_[9046]_  = ~\new_[20390]_  | ~\new_[21389]_ ;
  assign \new_[9047]_  = ~\new_[17531]_  & (~\new_[15221]_  | ~\new_[14840]_ );
  assign \new_[9048]_  = ~\new_[11504]_  | ~\new_[14163]_ ;
  assign \new_[9049]_  = \new_[11616]_  & \new_[15065]_ ;
  assign \new_[9050]_  = ~\new_[11546]_  | ~\new_[13645]_ ;
  assign \new_[9051]_  = ~\new_[17997]_  & ~\new_[14677]_ ;
  assign \new_[9052]_  = \new_[11616]_  & \new_[15399]_ ;
  assign \new_[9053]_  = ~\new_[13108]_  | ~\new_[13897]_ ;
  assign \new_[9054]_  = \new_[13846]_  | \new_[18692]_ ;
  assign \new_[9055]_  = ~\new_[17144]_  | ~\new_[11632]_ ;
  assign \new_[9056]_  = ~\new_[10264]_ ;
  assign \new_[9057]_  = \new_[11916]_  & \new_[17948]_ ;
  assign \new_[9058]_  = ~\new_[10861]_  | ~\new_[14126]_ ;
  assign \new_[9059]_  = ~\new_[11880]_  | ~\new_[11735]_ ;
  assign \new_[9060]_  = \new_[11915]_  | \new_[20099]_ ;
  assign \new_[9061]_  = \new_[15052]_  & \new_[13803]_ ;
  assign \new_[9062]_  = \new_[12061]_  & \new_[16879]_ ;
  assign \new_[9063]_  = ~\new_[10278]_ ;
  assign \new_[9064]_  = ~\new_[16525]_  | ~\new_[11568]_ ;
  assign \new_[9065]_  = \new_[11780]_  | \new_[18077]_ ;
  assign \new_[9066]_  = ~\new_[13711]_  | ~\new_[18937]_ ;
  assign \new_[9067]_  = \new_[11660]_  & \new_[12646]_ ;
  assign \new_[9068]_  = ~\new_[15099]_  & ~\new_[11654]_ ;
  assign \new_[9069]_  = ~\new_[12567]_  | ~\new_[14150]_ ;
  assign \new_[9070]_  = ~\new_[13336]_  | ~\new_[11708]_ ;
  assign \new_[9071]_  = ~\new_[11624]_  | ~\new_[14642]_ ;
  assign \new_[9072]_  = ~\new_[11941]_  & ~\new_[16432]_ ;
  assign \new_[9073]_  = \new_[11528]_  | \new_[19085]_ ;
  assign \new_[9074]_  = \new_[11996]_  | \new_[17689]_ ;
  assign \new_[9075]_  = \new_[12087]_  & \new_[17942]_ ;
  assign \new_[9076]_  = ~\new_[20907]_  | ~\new_[17472]_ ;
  assign \new_[9077]_  = \new_[15663]_  & \new_[11708]_ ;
  assign \new_[9078]_  = ~\new_[11820]_  & ~\new_[18087]_ ;
  assign \new_[9079]_  = ~\new_[14189]_  | ~\new_[14997]_ ;
  assign \new_[9080]_  = ~\new_[10298]_ ;
  assign \new_[9081]_  = ~\new_[21095]_  | ~\new_[11684]_ ;
  assign \new_[9082]_  = ~\new_[12077]_  | ~\new_[11847]_ ;
  assign \new_[9083]_  = ~\new_[11933]_  & ~\new_[18077]_ ;
  assign \new_[9084]_  = ~\new_[12743]_  | ~\new_[12018]_ ;
  assign \new_[9085]_  = \new_[11998]_  | \new_[12591]_ ;
  assign \new_[9086]_  = \new_[11876]_  | \new_[17358]_ ;
  assign \new_[9087]_  = ~\new_[13897]_  | ~\new_[11714]_ ;
  assign \new_[9088]_  = ~\new_[10876]_  | ~\new_[11849]_ ;
  assign \new_[9089]_  = \new_[11791]_  | \new_[18969]_ ;
  assign \new_[9090]_  = ~\new_[11747]_  | ~\new_[19180]_ ;
  assign \new_[9091]_  = ~\new_[10315]_ ;
  assign \new_[9092]_  = \new_[12588]_  & \new_[10861]_ ;
  assign \new_[9093]_  = ~\new_[11625]_  & ~\new_[11567]_ ;
  assign \new_[9094]_  = ~\new_[11960]_  | ~\new_[17043]_ ;
  assign \new_[9095]_  = ~\new_[11936]_  & ~\new_[12562]_ ;
  assign \new_[9096]_  = ~\new_[10321]_ ;
  assign \new_[9097]_  = ~\new_[12990]_  | ~\new_[11915]_ ;
  assign \new_[9098]_  = ~\new_[14158]_  | ~\new_[13698]_ ;
  assign \new_[9099]_  = ~\new_[13698]_  | ~\new_[11612]_ ;
  assign \new_[9100]_  = ~\new_[13463]_  & ~\new_[12506]_ ;
  assign \new_[9101]_  = \new_[13939]_  & \new_[10903]_ ;
  assign \new_[9102]_  = ~\new_[15334]_  | ~\new_[12009]_ ;
  assign \new_[9103]_  = ~\new_[11831]_  | ~\new_[19240]_ ;
  assign \new_[9104]_  = ~\new_[13382]_  | ~\new_[14424]_ ;
  assign \new_[9105]_  = ~\new_[10327]_ ;
  assign \new_[9106]_  = ~\new_[15073]_  | ~\new_[14677]_ ;
  assign \new_[9107]_  = ~\new_[13441]_  | ~\new_[14042]_ ;
  assign \new_[9108]_  = ~\new_[20488]_  | ~\new_[16991]_ ;
  assign \new_[9109]_  = ~\new_[16955]_  | ~\new_[12030]_ ;
  assign \new_[9110]_  = ~\new_[15547]_  | ~\new_[14123]_ ;
  assign \new_[9111]_  = ~\new_[11999]_  | ~\new_[12509]_ ;
  assign \new_[9112]_  = ~\new_[11978]_  | ~\new_[18124]_ ;
  assign \new_[9113]_  = ~\new_[21163]_  & ~\new_[14311]_ ;
  assign \new_[9114]_  = ~\new_[17275]_  | ~\new_[13754]_ ;
  assign \new_[9115]_  = ~\new_[19450]_  & ~\new_[11533]_ ;
  assign \new_[9116]_  = ~\new_[13200]_  | ~\new_[11738]_ ;
  assign \new_[9117]_  = ~\new_[11308]_  | ~\new_[13862]_ ;
  assign \new_[9118]_  = ~\new_[10341]_ ;
  assign \new_[9119]_  = ~\new_[10342]_ ;
  assign \new_[9120]_  = ~\new_[16796]_  | ~\new_[12006]_ ;
  assign \new_[9121]_  = \new_[18965]_  | \new_[14050]_ ;
  assign \new_[9122]_  = ~\new_[11809]_  | ~\new_[12732]_ ;
  assign \new_[9123]_  = ~\new_[11858]_  & ~\new_[18605]_ ;
  assign \new_[9124]_  = ~\new_[14604]_  | ~\new_[11881]_ ;
  assign \new_[9125]_  = \new_[14412]_  | \new_[18076]_ ;
  assign \new_[9126]_  = ~\new_[11596]_  | ~\new_[17522]_ ;
  assign \new_[9127]_  = ~\new_[10347]_ ;
  assign \new_[9128]_  = ~\new_[10903]_  | ~\new_[11764]_ ;
  assign \new_[9129]_  = ~\new_[10352]_ ;
  assign \new_[9130]_  = ~\new_[19592]_  & ~\new_[14152]_ ;
  assign \new_[9131]_  = ~\new_[13663]_  & ~\new_[18083]_ ;
  assign \new_[9132]_  = ~\new_[13899]_  & ~\new_[13528]_ ;
  assign \new_[9133]_  = ~\new_[11598]_  | ~\new_[15405]_ ;
  assign \new_[9134]_  = ~\new_[10360]_ ;
  assign \new_[9135]_  = \new_[11493]_  & \new_[11325]_ ;
  assign \new_[9136]_  = ~\new_[13311]_  | ~\new_[11586]_ ;
  assign \new_[9137]_  = ~\new_[14571]_  & ~\new_[11661]_ ;
  assign \new_[9138]_  = ~\new_[19073]_  & ~\new_[11697]_ ;
  assign \new_[9139]_  = ~\new_[11564]_  & ~\new_[11621]_ ;
  assign \new_[9140]_  = ~\new_[11606]_  | ~\new_[15050]_ ;
  assign \new_[9141]_  = ~\new_[12037]_  | ~\new_[19204]_ ;
  assign \new_[9142]_  = ~\new_[10367]_ ;
  assign \new_[9143]_  = \new_[12030]_  & \new_[13159]_ ;
  assign \new_[9144]_  = ~\new_[11704]_  | ~\new_[18845]_ ;
  assign \new_[9145]_  = ~\new_[13294]_  | ~\new_[14666]_  | ~\new_[13780]_ ;
  assign \new_[9146]_  = ~\new_[15615]_  | ~\new_[13525]_ ;
  assign \new_[9147]_  = ~\new_[18898]_  | ~\new_[11154]_ ;
  assign \new_[9148]_  = ~\new_[10376]_ ;
  assign \new_[9149]_  = ~\new_[12554]_  & ~\new_[11596]_ ;
  assign \new_[9150]_  = ~\new_[12916]_  | ~\new_[20232]_ ;
  assign \new_[9151]_  = ~\new_[13813]_  | ~\new_[11361]_ ;
  assign \new_[9152]_  = \new_[17917]_  & \new_[11717]_ ;
  assign \new_[9153]_  = ~\new_[11668]_  | ~\new_[15396]_ ;
  assign \new_[9154]_  = ~\new_[11154]_  | ~\new_[18166]_ ;
  assign \new_[9155]_  = ~\new_[11711]_  | ~\new_[16243]_ ;
  assign \new_[9156]_  = ~\new_[14809]_  | ~\new_[11342]_ ;
  assign \new_[9157]_  = ~\new_[11624]_  | ~\new_[13882]_ ;
  assign \new_[9158]_  = ~\new_[12795]_  | ~\new_[17845]_ ;
  assign \new_[9159]_  = ~\new_[12012]_  | ~\new_[17089]_ ;
  assign \new_[9160]_  = ~\new_[10387]_ ;
  assign \new_[9161]_  = ~\new_[11715]_  & ~\new_[18863]_ ;
  assign \new_[9162]_  = ~\new_[12451]_  | ~\new_[11983]_ ;
  assign \new_[9163]_  = ~\new_[19018]_  & ~\new_[14615]_ ;
  assign \new_[9164]_  = ~\new_[20808]_  | ~\new_[15210]_ ;
  assign \new_[9165]_  = ~\new_[12159]_  | ~\new_[11762]_ ;
  assign \new_[9166]_  = \new_[11513]_  & \new_[16143]_ ;
  assign \new_[9167]_  = ~\new_[10396]_ ;
  assign \new_[9168]_  = ~\new_[11576]_  | ~\new_[12520]_ ;
  assign \new_[9169]_  = \new_[13795]_  & \new_[11161]_ ;
  assign \new_[9170]_  = ~\new_[11624]_  | ~\new_[16925]_ ;
  assign \new_[9171]_  = ~\new_[15577]_  | ~\new_[11725]_ ;
  assign \new_[9172]_  = ~\new_[13401]_  | ~\new_[13662]_  | ~\new_[15813]_ ;
  assign \new_[9173]_  = ~\new_[10403]_ ;
  assign \new_[9174]_  = ~\new_[15473]_  | ~\new_[14437]_  | ~\new_[15672]_ ;
  assign \new_[9175]_  = \new_[11856]_  | \new_[14444]_ ;
  assign \new_[9176]_  = ~\new_[12052]_  | ~\new_[19247]_ ;
  assign \new_[9177]_  = ~\new_[13388]_  | ~\new_[11764]_ ;
  assign \new_[9178]_  = ~\new_[11795]_  | (~\new_[16270]_  & ~\new_[18166]_ );
  assign \new_[9179]_  = ~\new_[12080]_  | ~\new_[14126]_ ;
  assign \new_[9180]_  = ~\new_[13896]_  | ~\new_[21347]_ ;
  assign \new_[9181]_  = ~\new_[12648]_  | ~\new_[21547]_ ;
  assign \new_[9182]_  = ~\new_[11754]_  | (~\new_[13367]_  & ~\new_[18984]_ );
  assign \new_[9183]_  = ~\new_[11939]_  | ~\new_[14099]_ ;
  assign \new_[9184]_  = \new_[11680]_  & \new_[17663]_ ;
  assign \new_[9185]_  = ~\new_[11925]_  | ~\new_[14615]_ ;
  assign \new_[9186]_  = ~\new_[13160]_  & ~\new_[11846]_ ;
  assign \new_[9187]_  = ~\new_[15434]_  & ~\new_[11890]_ ;
  assign \new_[9188]_  = ~\new_[15099]_  & ~\new_[11886]_ ;
  assign \new_[9189]_  = ~\new_[16117]_  | ~\new_[11701]_ ;
  assign \new_[9190]_  = ~\new_[10427]_ ;
  assign \new_[9191]_  = ~\new_[12020]_  & ~\new_[12686]_ ;
  assign \new_[9192]_  = ~\new_[10430]_ ;
  assign \new_[9193]_  = ~\new_[14418]_  | (~\new_[13370]_  & ~\new_[21115]_ );
  assign \new_[9194]_  = ~\new_[20680]_  & (~\new_[15116]_  | ~\new_[14825]_ );
  assign \new_[9195]_  = ~\new_[11622]_  & ~\new_[15257]_ ;
  assign \new_[9196]_  = ~\new_[11911]_  & (~\new_[18614]_  | ~\new_[18060]_ );
  assign \new_[9197]_  = ~\new_[13929]_  | ~\new_[11749]_ ;
  assign \new_[9198]_  = ~\new_[12582]_  & (~\new_[13440]_  | ~\new_[18120]_ );
  assign \new_[9199]_  = ~\new_[11655]_  | ~\new_[11744]_ ;
  assign \new_[9200]_  = ~\new_[11383]_  & (~\new_[17964]_  | ~\new_[21638]_ );
  assign \new_[9201]_  = ~\new_[11932]_  | ~\new_[14487]_ ;
  assign \new_[9202]_  = ~\new_[13928]_  | (~\new_[15407]_  & ~\new_[17358]_ );
  assign \new_[9203]_  = ~\new_[21635]_  & (~\new_[15784]_  | ~\new_[13447]_ );
  assign \new_[9204]_  = ~\new_[11884]_  | ~\new_[18522]_ ;
  assign \new_[9205]_  = ~\new_[18124]_  & (~\new_[15917]_  | ~\new_[15694]_ );
  assign \new_[9206]_  = ~\new_[11865]_  & (~\new_[18590]_  | ~\new_[19408]_ );
  assign \new_[9207]_  = ~\new_[12055]_  | ~\new_[19021]_ ;
  assign \new_[9208]_  = ~\new_[11720]_  | ~\new_[13725]_ ;
  assign \new_[9209]_  = ~\new_[13699]_  & ~\new_[11457]_ ;
  assign \new_[9210]_  = ~\new_[11548]_  & (~\new_[17147]_  | ~\new_[21542]_ );
  assign \new_[9211]_  = ~\new_[11707]_  & (~\new_[16323]_  | ~\new_[18973]_ );
  assign \new_[9212]_  = ~\new_[11685]_  | ~\new_[13775]_ ;
  assign \new_[9213]_  = ~\new_[11713]_  | ~\new_[12977]_ ;
  assign \new_[9214]_  = ~\new_[13783]_  | ~\new_[11817]_ ;
  assign \new_[9215]_  = ~\new_[10458]_ ;
  assign \new_[9216]_  = ~\new_[11690]_  | ~\new_[14086]_ ;
  assign \new_[9217]_  = ~\new_[14175]_  | ~\new_[11559]_ ;
  assign \new_[9218]_  = ~\new_[11580]_  & (~\new_[15828]_  | ~\new_[19275]_ );
  assign \new_[9219]_  = ~\new_[11639]_  | ~\new_[11229]_ ;
  assign \new_[9220]_  = ~\new_[15416]_  | ~\new_[11539]_ ;
  assign \new_[9221]_  = ~\new_[11583]_  | ~\new_[15028]_ ;
  assign \new_[9222]_  = ~\new_[13934]_  | ~\new_[11982]_ ;
  assign \new_[9223]_  = ~\new_[15032]_  & ~\new_[12099]_ ;
  assign \new_[9224]_  = ~\new_[13965]_  & ~\new_[11144]_ ;
  assign \new_[9225]_  = ~\new_[11642]_  & (~\new_[18543]_  | ~\new_[18045]_ );
  assign \new_[9226]_  = ~\new_[11617]_  | ~\new_[11669]_ ;
  assign \new_[9227]_  = ~\new_[17486]_  | (~\new_[16623]_  & ~\new_[13399]_ );
  assign \new_[9228]_  = ~\new_[18434]_  | (~\new_[17355]_  & ~\new_[13399]_ );
  assign \new_[9229]_  = ~\new_[11325]_  | (~\new_[17531]_  & ~\new_[17564]_ );
  assign \new_[9230]_  = ~\new_[15764]_  | ~\new_[11569]_ ;
  assign \new_[9231]_  = ~\new_[11761]_  | ~\new_[18115]_ ;
  assign \new_[9232]_  = ~\new_[13803]_  | (~\new_[18796]_  & ~\new_[17584]_ );
  assign \new_[9233]_  = ~\new_[15728]_  | ~\new_[11710]_ ;
  assign \new_[9234]_  = ~\new_[15739]_  | ~\new_[13724]_ ;
  assign \new_[9235]_  = ~\new_[14052]_  | (~\new_[18875]_  & ~\new_[17344]_ );
  assign \new_[9236]_  = ~\new_[14163]_  | (~\new_[17969]_  & ~\new_[16512]_ );
  assign \new_[9237]_  = ~\new_[15745]_  | ~\new_[13859]_ ;
  assign \new_[9238]_  = ~\new_[13645]_  | (~\new_[18711]_  & ~\new_[18309]_ );
  assign \new_[9239]_  = ~\new_[11883]_  & (~\new_[17471]_  | ~\new_[16958]_ );
  assign \new_[9240]_  = ~\new_[11899]_  | ~\new_[16022]_ ;
  assign \new_[9241]_  = ~\new_[18807]_  | (~\new_[17094]_  & ~\new_[16872]_ );
  assign \new_[9242]_  = ~\new_[11964]_  | ~\new_[11797]_ ;
  assign \new_[9243]_  = ~\new_[14864]_  | ~\new_[11633]_  | ~\new_[15897]_ ;
  assign \new_[9244]_  = ~\new_[12040]_  | ~\new_[13309]_ ;
  assign \new_[9245]_  = ~\new_[11944]_  | ~\new_[12665]_ ;
  assign \new_[9246]_  = ~\new_[15531]_  | ~\new_[20221]_ ;
  assign \new_[9247]_  = ~\new_[13496]_  | (~\new_[12280]_  & ~\new_[18846]_ );
  assign \new_[9248]_  = ~\new_[11958]_  | ~\new_[11566]_ ;
  assign \new_[9249]_  = ~\new_[11822]_  | ~\new_[11757]_ ;
  assign \new_[9250]_  = ~\new_[11977]_  | ~\new_[11643]_ ;
  assign \new_[9251]_  = ~\new_[11864]_  | ~\new_[11994]_ ;
  assign \new_[9252]_  = ~\new_[11853]_  | ~\new_[11547]_ ;
  assign \new_[9253]_  = \new_[18856]_  ^ \new_[13452]_ ;
  assign \new_[9254]_  = \new_[18712]_  ^ \new_[13456]_ ;
  assign \new_[9255]_  = \new_[18915]_  ^ \new_[12449]_ ;
  assign \new_[9256]_  = \new_[18880]_  ^ \new_[12693]_ ;
  assign \new_[9257]_  = \new_[18865]_  ^ \new_[13460]_ ;
  assign \new_[9258]_  = \new_[18918]_  ^ \new_[13459]_ ;
  assign \new_[9259]_  = ~\new_[12123]_  & ~\new_[18421]_ ;
  assign \new_[9260]_  = ~\new_[14913]_  | ~\new_[13627]_  | ~\new_[11870]_  | ~\new_[13326]_ ;
  assign \new_[9261]_  = ~\new_[10507]_ ;
  assign \new_[9262]_  = ~\new_[11350]_  & ~\new_[11696]_ ;
  assign \new_[9263]_  = ~\new_[11172]_  | ~\new_[19261]_ ;
  assign \new_[9264]_  = ~\new_[11993]_  | ~\new_[18621]_ ;
  assign \new_[9265]_  = ~\new_[10545]_ ;
  assign \new_[9266]_  = ~\new_[10551]_ ;
  assign \new_[9267]_  = ~\new_[14596]_  | ~\new_[21508]_ ;
  assign \new_[9268]_  = \new_[13498]_  | \new_[18682]_ ;
  assign \new_[9269]_  = ~\new_[10559]_ ;
  assign \new_[9270]_  = \new_[13594]_  | \new_[18747]_ ;
  assign \new_[9271]_  = ~\new_[10561]_ ;
  assign \new_[9272]_  = \new_[12091]_  | \new_[18973]_ ;
  assign \new_[9273]_  = ~\new_[10564]_ ;
  assign \new_[9274]_  = ~\new_[10563]_ ;
  assign \new_[9275]_  = ~\new_[9672]_ ;
  assign \new_[9276]_  = \new_[11980]_  | \new_[18984]_ ;
  assign \new_[9277]_  = ~\new_[12780]_ ;
  assign \new_[9278]_  = ~\new_[10578]_ ;
  assign \new_[9279]_  = ~\new_[10578]_ ;
  assign \new_[9280]_  = ~\new_[10578]_ ;
  assign \new_[9281]_  = ~\new_[10581]_ ;
  assign \new_[9282]_  = ~\new_[10583]_ ;
  assign \new_[9283]_  = ~\new_[10587]_ ;
  assign \new_[9284]_  = ~\new_[18584]_  | ~\new_[14665]_ ;
  assign \new_[9285]_  = ~\new_[12079]_  | ~\new_[18825]_ ;
  assign \new_[9286]_  = ~\new_[10591]_ ;
  assign \new_[9287]_  = ~\new_[14674]_  & ~\new_[12090]_ ;
  assign \new_[9288]_  = ~\new_[10605]_ ;
  assign \new_[9289]_  = \new_[13594]_  & \new_[15394]_ ;
  assign \new_[9290]_  = ~\new_[12106]_  | ~\new_[15523]_ ;
  assign \new_[9291]_  = ~\new_[16400]_  & ~\new_[14233]_ ;
  assign \new_[9292]_  = \new_[12074]_  | \new_[14951]_ ;
  assign \new_[9293]_  = ~\new_[10614]_ ;
  assign \new_[9294]_  = ~\new_[17468]_  | ~\new_[21703]_ ;
  assign \new_[9295]_  = \new_[12114]_  | \new_[15530]_ ;
  assign \new_[9296]_  = ~\new_[12074]_  & ~\new_[18423]_ ;
  assign \new_[9297]_  = ~\new_[12108]_  | ~\new_[15778]_ ;
  assign \new_[9298]_  = ~\new_[10624]_ ;
  assign \new_[9299]_  = ~\new_[13632]_  & ~\new_[19277]_ ;
  assign \new_[9300]_  = ~\new_[20660]_ ;
  assign \new_[9301]_  = ~\new_[11638]_  | ~\new_[14955]_ ;
  assign \new_[9302]_  = ~\new_[10628]_ ;
  assign \new_[9303]_  = ~\new_[21703]_  | ~\new_[16832]_ ;
  assign \new_[9304]_  = ~\new_[10635]_ ;
  assign \new_[9305]_  = ~\new_[14422]_  | ~\new_[18166]_ ;
  assign \new_[9306]_  = ~\new_[10645]_ ;
  assign \new_[9307]_  = ~\new_[14789]_  | ~\new_[12091]_ ;
  assign \new_[9308]_  = ~\new_[12075]_  & ~\new_[19659]_ ;
  assign \new_[9309]_  = ~\new_[10656]_ ;
  assign \new_[9310]_  = ~\new_[19578]_  & (~\new_[14451]_  | ~\new_[12436]_ );
  assign \new_[9311]_  = ~\new_[10665]_ ;
  assign \new_[9312]_  = ~\new_[10667]_ ;
  assign \new_[9313]_  = \new_[12110]_  | \new_[14826]_ ;
  assign \new_[9314]_  = ~\new_[19240]_  | (~\new_[12370]_  & ~\new_[13853]_ );
  assign \new_[9315]_  = ~\new_[21056]_  | (~\new_[12354]_  & ~\new_[12628]_ );
  assign \new_[9316]_  = ~\new_[18187]_  | (~\new_[12437]_  & ~\new_[13810]_ );
  assign \new_[9317]_  = ~\new_[19204]_  | (~\new_[12352]_  & ~\new_[13918]_ );
  assign \new_[9318]_  = ~\new_[19021]_  | (~\new_[12376]_  & ~\new_[15090]_ );
  assign \new_[9319]_  = ~\new_[10670]_ ;
  assign \new_[9320]_  = ~\new_[20341]_  | (~\new_[12402]_  & ~\new_[13708]_ );
  assign \new_[9321]_  = ~\new_[20100]_  | (~\new_[12410]_  & ~\new_[13808]_ );
  assign \new_[9322]_  = ~\new_[19094]_  | (~\new_[12319]_  & ~\new_[13759]_ );
  assign \new_[9323]_  = ~\new_[21635]_  | (~\new_[12416]_  & ~\new_[13931]_ );
  assign \new_[9324]_  = ~\new_[21558]_  | (~\new_[12419]_  & ~\new_[13773]_ );
  assign \new_[9325]_  = \new_[11980]_  & \new_[16307]_ ;
  assign \new_[9326]_  = ~\new_[12296]_  | ~\new_[14532]_  | ~\new_[15621]_ ;
  assign \new_[9327]_  = ~\new_[13830]_  & (~\new_[12434]_  | ~\new_[18965]_ );
  assign \new_[9328]_  = ~\new_[12314]_  | ~\new_[11891]_  | ~\new_[15717]_ ;
  assign \new_[9329]_  = ~\new_[21388]_  & ~\new_[13492]_ ;
  assign \new_[9330]_  = \\u0_r0_out_reg[25] ;
  assign \new_[9331]_  = ~\new_[12109]_  | ~\new_[15778]_ ;
  assign \new_[9332]_  = ~\new_[19202]_  & (~\new_[16664]_  | ~\new_[12400]_ );
  assign \new_[9333]_  = ~\new_[11651]_  & ~\new_[19170]_ ;
  assign \new_[9334]_  = ~\new_[19094]_  & (~\new_[12796]_  | ~\new_[12156]_ );
  assign \new_[9335]_  = \new_[12096]_  | \new_[18228]_ ;
  assign \new_[9336]_  = ~\new_[16850]_  & ~\new_[13605]_ ;
  assign \new_[9337]_  = ~\new_[14387]_  | ~\new_[11087]_  | ~\new_[13549]_ ;
  assign \new_[9338]_  = ~\new_[10732]_ ;
  assign \new_[9339]_  = \new_[12074]_  & \new_[12072]_ ;
  assign \new_[9340]_  = ~\new_[19088]_  | (~\new_[12479]_  & ~\new_[14456]_ );
  assign \new_[9341]_  = ~\new_[10690]_ ;
  assign \new_[9342]_  = ~\new_[12103]_  | ~\new_[15523]_ ;
  assign \new_[9343]_  = ~\new_[10693]_ ;
  assign \new_[9344]_  = ~\new_[10695]_ ;
  assign \new_[9345]_  = \new_[12125]_  & \new_[13560]_ ;
  assign \new_[9346]_  = ~\new_[19567]_  & (~\new_[12278]_  | ~\new_[13557]_ );
  assign \new_[9347]_  = ~\new_[18124]_  & (~\new_[12435]_  | ~\new_[12710]_ );
  assign \new_[9348]_  = ~\new_[10606]_ ;
  assign \new_[9349]_  = \new_[15710]_  & \new_[12072]_ ;
  assign \new_[9350]_  = ~\new_[19343]_  | (~\new_[12458]_  & ~\new_[13139]_ );
  assign \new_[9351]_  = ~\new_[19239]_  | (~\new_[12480]_  & ~\new_[16019]_ );
  assign \new_[9352]_  = \new_[12116]_  & \new_[12339]_ ;
  assign \new_[9353]_  = ~\new_[10365]_ ;
  assign \new_[9354]_  = ~\new_[12208]_  | ~\new_[14242]_  | ~\new_[14070]_ ;
  assign \new_[9355]_  = ~\new_[10267]_ ;
  assign \new_[9356]_  = ~\new_[10267]_ ;
  assign \new_[9357]_  = ~\new_[12112]_  | ~\new_[15523]_ ;
  assign \new_[9358]_  = ~\new_[10185]_ ;
  assign \new_[9359]_  = ~\new_[12073]_  | ~\new_[18692]_ ;
  assign \new_[9360]_  = ~\new_[13554]_  | ~\new_[16222]_  | ~\new_[13609]_ ;
  assign \new_[9361]_  = ~\new_[10710]_ ;
  assign \new_[9362]_  = ~\new_[19553]_  | (~\new_[12482]_  & ~\new_[18003]_ );
  assign \new_[9363]_  = ~\new_[14860]_  | ~\new_[12081]_ ;
  assign \new_[9364]_  = ~\new_[13417]_  | ~\new_[13640]_ ;
  assign \new_[9365]_  = ~\new_[17407]_  & ~\new_[13559]_ ;
  assign \new_[9366]_  = ~\new_[13469]_  | ~\new_[13594]_ ;
  assign \new_[9367]_  = ~\new_[19249]_  | (~\new_[12335]_  & ~\new_[15587]_ );
  assign \new_[9368]_  = ~\new_[12097]_  & (~\new_[16628]_  | ~\new_[15827]_ );
  assign \new_[9369]_  = ~\new_[19145]_  | (~\new_[12483]_  & ~\new_[15443]_ );
  assign n2718 = ~\new_[17681]_  & (~\new_[13475]_  | ~\new_[14785]_ );
  assign \new_[9371]_  = ~\new_[12152]_  | ~\new_[11162]_  | ~\new_[12939]_ ;
  assign \new_[9372]_  = ~\new_[13980]_  | ~\new_[14370]_  | ~\new_[12156]_  | ~\new_[14240]_ ;
  assign \new_[9373]_  = ~\new_[12820]_  | ~\new_[11433]_  | ~\new_[21616]_ ;
  assign \new_[9374]_  = ~\new_[13225]_  | ~\new_[12461]_  | ~\new_[12306]_ ;
  assign \new_[9375]_  = ~\new_[12119]_  | ~\new_[19378]_ ;
  assign \new_[9376]_  = ~\new_[13616]_  | ~\new_[11203]_  | ~\new_[13583]_ ;
  assign \new_[9377]_  = ~\new_[19145]_  & (~\new_[12467]_  | ~\new_[15003]_ );
  assign \new_[9378]_  = ~\new_[14130]_  | ~\new_[13751]_  | ~\new_[10916]_  | ~\new_[14066]_ ;
  assign \new_[9379]_  = ~\new_[14114]_  | ~\new_[16556]_  | ~\new_[10931]_  | ~\new_[16251]_ ;
  assign \new_[9380]_  = ~\new_[12130]_  & ~\new_[11963]_ ;
  assign \new_[9381]_  = ~\new_[14082]_  | ~\new_[16125]_  | ~\new_[10967]_  | ~\new_[16226]_ ;
  assign \new_[9382]_  = \new_[12141]_  & \new_[18077]_ ;
  assign \new_[9383]_  = \new_[10849]_  & \new_[19249]_ ;
  assign \new_[9384]_  = ~\new_[12175]_  | ~\new_[21678]_  | ~\new_[13272]_ ;
  assign \new_[9385]_  = ~\new_[15585]_  | ~\new_[16173]_  | ~\new_[12218]_  | ~\new_[13239]_ ;
  assign \new_[9386]_  = ~\new_[14177]_  | ~\new_[16077]_  | ~\new_[11036]_  | ~\new_[12948]_ ;
  assign \new_[9387]_  = ~\new_[14351]_  | ~\new_[13964]_  | ~\new_[11073]_  | ~\new_[14166]_ ;
  assign \new_[9388]_  = ~\new_[14106]_  | ~\new_[12592]_  | ~\new_[12210]_ ;
  assign \new_[9389]_  = (~\new_[12462]_  | ~\new_[19377]_ ) & (~\new_[16135]_  | ~\new_[18981]_ );
  assign \new_[9390]_  = \new_[12277]_  ? \new_[18194]_  : \new_[15181]_ ;
  assign \new_[9391]_  = \new_[12253]_  ? \new_[19102]_  : \new_[12716]_ ;
  assign \new_[9392]_  = ~\new_[13924]_  | ~\new_[17787]_  | ~\new_[11085]_  | ~\new_[15250]_ ;
  assign \new_[9393]_  = ~\new_[11852]_  & (~\new_[12460]_  | ~\new_[18179]_ );
  assign \new_[9394]_  = ~\new_[14218]_  | ~\new_[16077]_  | ~\new_[14832]_  | ~\new_[13496]_ ;
  assign \new_[9395]_  = ~\new_[16268]_  | ~\new_[13964]_  | ~\new_[13692]_  | ~\new_[14036]_ ;
  assign \new_[9396]_  = \new_[19766]_  ^ \new_[19203]_ ;
  assign \new_[9397]_  = ~\new_[19612]_  | (~\new_[13267]_  & ~\new_[16616]_ );
  assign \new_[9398]_  = ~\new_[17874]_  & (~\new_[13371]_  | ~\new_[14358]_ );
  assign \new_[9399]_  = ~\new_[21115]_  | (~\new_[12927]_  & ~\new_[16010]_ );
  assign \new_[9400]_  = \new_[19793]_  ^ \new_[19098]_ ;
  assign \new_[9401]_  = ~\new_[18941]_  & (~\new_[12633]_  | ~\new_[16263]_ );
  assign \new_[9402]_  = ~\new_[21413]_  | (~\new_[13082]_  & ~\new_[15992]_ );
  assign \new_[9403]_  = ~\new_[19072]_  & (~\new_[13387]_  | ~\new_[16243]_ );
  assign \new_[9404]_  = ~\new_[16879]_  & (~\new_[15718]_  | ~\new_[15210]_ );
  assign \new_[9405]_  = ~\new_[19247]_  & (~\new_[12773]_  | ~\new_[15599]_ );
  assign \new_[9406]_  = ~\new_[17472]_  & (~\new_[13423]_  | ~\new_[13199]_ );
  assign \new_[9407]_  = ~\new_[19625]_  | (~\new_[13248]_  & ~\new_[14608]_ );
  assign \new_[9408]_  = ~\new_[19261]_  | (~\new_[13128]_  & ~\new_[14498]_ );
  assign \new_[9409]_  = ~\new_[19244]_  | (~\new_[13307]_  & ~\new_[16432]_ );
  assign \new_[9410]_  = \new_[16854]_  ^ \new_[19561]_ ;
  assign \new_[9411]_  = ~\new_[19161]_  | (~\new_[13103]_  & ~\new_[15969]_ );
  assign \new_[9412]_  = \new_[19739]_  ^ \new_[19156]_ ;
  assign \new_[9413]_  = ~\new_[19079]_  | (~\new_[13039]_  & ~\new_[14724]_ );
  assign \new_[9414]_  = ~\new_[18280]_  | (~\new_[12942]_  & ~\new_[13412]_ );
  assign \new_[9415]_  = ~\new_[19088]_  | (~\new_[13126]_  & ~\new_[17394]_ );
  assign \new_[9416]_  = ~\new_[18821]_  | (~\new_[12323]_  & ~\new_[16297]_ );
  assign \new_[9417]_  = ~\new_[10755]_ ;
  assign \new_[9418]_  = ~\new_[19261]_  & (~\new_[13448]_  | ~\new_[13795]_ );
  assign \new_[9419]_  = ~\new_[19261]_  | (~\new_[13115]_  & ~\new_[13373]_ );
  assign \new_[9420]_  = ~\new_[11395]_  & ~\new_[18542]_ ;
  assign \new_[9421]_  = ~\new_[21115]_  | (~\new_[12888]_  & ~\new_[13372]_ );
  assign \new_[9422]_  = ~\new_[19094]_  | (~\new_[12865]_  & ~\new_[15512]_ );
  assign \new_[9423]_  = ~\new_[21115]_  & (~\new_[12952]_  | ~\new_[13939]_ );
  assign \new_[9424]_  = ~\new_[14951]_  & (~\new_[12421]_  | ~\new_[13951]_ );
  assign \new_[9425]_  = ~\new_[19687]_  | (~\new_[13244]_  & ~\new_[13580]_ );
  assign \new_[9426]_  = ~\new_[19450]_  | (~\new_[12144]_  & ~\new_[16387]_ );
  assign \new_[9427]_  = ~\new_[19592]_  | (~\new_[13182]_  & ~\new_[16640]_ );
  assign \new_[9428]_  = ~\new_[11141]_  | ~\new_[19748]_ ;
  assign \new_[9429]_  = ~\new_[10759]_ ;
  assign \new_[9430]_  = ~\new_[960]_  & (~\new_[14553]_  | ~\new_[12895]_ );
  assign \new_[9431]_  = \new_[11318]_  & \new_[19277]_ ;
  assign \new_[9432]_  = \new_[11322]_  & \new_[19006]_ ;
  assign \new_[9433]_  = ~\new_[999]_  & (~\new_[14562]_  | ~\new_[13159]_ );
  assign \new_[9434]_  = ~\new_[18983]_  & (~\new_[15624]_  | ~\new_[13106]_ );
  assign \new_[9435]_  = \new_[11367]_  & \new_[19659]_ ;
  assign \new_[9436]_  = ~\new_[1039]_  & (~\new_[13422]_  | ~\new_[13149]_ );
  assign \new_[9437]_  = ~\new_[10764]_ ;
  assign \new_[9438]_  = ~\new_[11045]_  | ~\new_[18194]_ ;
  assign \new_[9439]_  = \new_[10920]_  | \new_[19547]_ ;
  assign \new_[9440]_  = \new_[14476]_  | \new_[18496]_  | \new_[19612]_  | \new_[18166]_ ;
  assign \new_[9441]_  = ~\new_[10767]_ ;
  assign \new_[9442]_  = ~\new_[10904]_  & ~\new_[18998]_ ;
  assign \new_[9443]_  = ~\new_[11182]_  & ~\new_[18481]_ ;
  assign \new_[9444]_  = \new_[10966]_  | \new_[18194]_ ;
  assign \new_[9445]_  = \new_[11166]_  & \new_[18965]_ ;
  assign \new_[9446]_  = ~\new_[18652]_  | ~\new_[19145]_  | ~\new_[12611]_ ;
  assign \new_[9447]_  = ~\new_[11401]_  & (~\new_[13702]_  | ~\new_[17544]_ );
  assign \new_[9448]_  = ~\new_[10936]_  & ~\new_[19115]_ ;
  assign \new_[9449]_  = ~\new_[10901]_  | ~\new_[19366]_ ;
  assign \new_[9450]_  = ~\new_[18443]_  | ~\new_[20680]_  | ~\new_[13040]_ ;
  assign \new_[9451]_  = ~\new_[19450]_  & ~\new_[10974]_ ;
  assign \new_[9452]_  = ~\new_[10971]_  | ~\new_[19532]_ ;
  assign \new_[9453]_  = \new_[11377]_  & \new_[18569]_ ;
  assign \new_[9454]_  = \new_[14526]_  | \new_[17572]_  | \new_[19625]_  | \new_[18228]_ ;
  assign \new_[9455]_  = ~\new_[11369]_  & ~\new_[19233]_ ;
  assign \new_[9456]_  = \new_[11267]_  | \new_[18070]_ ;
  assign \new_[9457]_  = ~\new_[10925]_  & ~\new_[18076]_ ;
  assign \new_[9458]_  = \new_[11233]_  & \new_[17472]_ ;
  assign \new_[9459]_  = \new_[11310]_  & \new_[19288]_ ;
  assign \new_[9460]_  = \new_[14603]_  | \new_[19386]_  | \new_[19450]_  | \new_[18984]_ ;
  assign \new_[9461]_  = ~\new_[10930]_  | ~\new_[18076]_ ;
  assign \new_[9462]_  = ~\new_[1025]_  & (~\new_[13214]_  | ~\new_[13030]_ );
  assign \new_[9463]_  = ~\new_[18983]_  & (~\new_[14364]_  | ~\new_[12966]_ );
  assign \new_[9464]_  = ~\new_[18380]_  | (~\new_[12933]_  & ~\new_[16306]_ );
  assign \new_[9465]_  = ~\new_[11171]_  | ~\new_[20239]_ ;
  assign \new_[9466]_  = ~\new_[17182]_  | ~\new_[14367]_  | ~\new_[15137]_ ;
  assign \new_[9467]_  = \new_[11453]_  | \new_[19102]_ ;
  assign \new_[9468]_  = ~\new_[11081]_  | ~\new_[19071]_ ;
  assign \new_[9469]_  = ~\new_[10779]_ ;
  assign \new_[9470]_  = ~\new_[11094]_  | ~\new_[12305]_ ;
  assign \new_[9471]_  = ~\new_[10988]_  | ~\new_[12163]_ ;
  assign \new_[9472]_  = ~\new_[11335]_  | ~\new_[21686]_ ;
  assign \new_[9473]_  = \new_[11088]_  | \new_[11740]_ ;
  assign \new_[9474]_  = ~\new_[12507]_  | ~\new_[21600]_  | ~\new_[15570]_ ;
  assign \new_[9475]_  = ~\new_[11093]_  | ~\new_[18984]_ ;
  assign \new_[9476]_  = ~\new_[11727]_  | ~\new_[10896]_ ;
  assign \new_[9477]_  = ~\new_[13603]_  | ~\new_[10936]_ ;
  assign \new_[9478]_  = ~\new_[11110]_  & ~\new_[15060]_ ;
  assign \new_[9479]_  = ~\new_[19079]_  & (~\new_[13353]_  | ~\new_[15127]_ );
  assign \new_[9480]_  = ~\new_[17379]_  & (~\new_[13069]_  | ~\new_[13337]_ );
  assign \new_[9481]_  = ~\new_[11024]_  | ~\new_[11869]_ ;
  assign \new_[9482]_  = ~\new_[18087]_  & (~\new_[14089]_  | ~\new_[12639]_ );
  assign \new_[9483]_  = ~\new_[10925]_  | ~\new_[10966]_ ;
  assign \new_[9484]_  = ~\new_[11448]_  | ~\new_[17874]_ ;
  assign \new_[9485]_  = ~\new_[21060]_  | ~\new_[17874]_ ;
  assign \new_[9486]_  = ~\new_[21251]_  | ~\new_[19013]_ ;
  assign \new_[9487]_  = ~\new_[11310]_  & ~\new_[16120]_ ;
  assign \new_[9488]_  = \new_[11122]_  & \new_[15175]_ ;
  assign \new_[9489]_  = ~\new_[11359]_  | ~\new_[18941]_ ;
  assign \new_[9490]_  = ~\new_[10904]_  | ~\new_[16266]_ ;
  assign \new_[9491]_  = ~\new_[15095]_  | ~\new_[13557]_  | ~\new_[15860]_ ;
  assign \new_[9492]_  = ~\new_[11413]_  & ~\new_[14135]_ ;
  assign \new_[9493]_  = ~\new_[17353]_  | ~\new_[14123]_  | ~\new_[14842]_ ;
  assign \new_[9494]_  = ~\new_[10787]_ ;
  assign \new_[9495]_  = \new_[11406]_  | \new_[17379]_ ;
  assign \new_[9496]_  = ~\new_[20723]_  | ~\new_[17727]_ ;
  assign \new_[9497]_  = ~\new_[10893]_  | ~\new_[18288]_ ;
  assign \new_[9498]_  = ~\new_[13817]_  | ~\new_[14880]_  | ~\new_[12907]_ ;
  assign \new_[9499]_  = ~\new_[15211]_  | ~\new_[14123]_  | ~\new_[15095]_ ;
  assign \new_[9500]_  = ~\new_[11133]_  | ~\new_[18627]_ ;
  assign \new_[9501]_  = ~\new_[14533]_  | ~\new_[16353]_  | ~\new_[15256]_ ;
  assign \new_[9502]_  = \new_[10909]_  | \new_[18194]_ ;
  assign \new_[9503]_  = ~\new_[10791]_ ;
  assign \new_[9504]_  = ~\new_[13925]_  | ~\new_[14672]_  | ~\new_[15342]_ ;
  assign \new_[9505]_  = ~\new_[10921]_  | ~\new_[15140]_ ;
  assign \new_[9506]_  = ~\new_[10918]_  | ~\new_[11881]_ ;
  assign \new_[9507]_  = ~\new_[13546]_  | ~\new_[20232]_ ;
  assign \new_[9508]_  = ~\new_[11088]_  | ~\new_[19261]_ ;
  assign \new_[9509]_  = ~\new_[10796]_ ;
  assign \new_[9510]_  = ~\new_[10994]_  | ~\new_[13159]_ ;
  assign \new_[9511]_  = ~\new_[12418]_  | ~\new_[12567]_ ;
  assign \new_[9512]_  = ~\new_[10920]_  | ~\new_[14120]_ ;
  assign \new_[9513]_  = ~\new_[11461]_  & ~\new_[21328]_ ;
  assign \new_[9514]_  = ~\new_[18762]_  & (~\new_[14090]_  | ~\new_[13457]_ );
  assign \new_[9515]_  = \new_[11295]_  & \new_[18965]_ ;
  assign \new_[9516]_  = \new_[11473]_  | \new_[13770]_ ;
  assign \new_[9517]_  = ~\new_[10798]_ ;
  assign \new_[9518]_  = \new_[13979]_  & \new_[12436]_ ;
  assign \new_[9519]_  = ~\new_[13484]_  | ~\new_[21329]_ ;
  assign \new_[9520]_  = ~\new_[11212]_  & ~\new_[19156]_ ;
  assign \new_[9521]_  = ~\new_[13620]_  & ~\new_[19547]_ ;
  assign \new_[9522]_  = ~\new_[16728]_  & ~\new_[11171]_ ;
  assign \new_[9523]_  = \new_[12439]_  & \new_[11058]_ ;
  assign \new_[9524]_  = ~\new_[11155]_  | ~\new_[19727]_ ;
  assign \new_[9525]_  = \new_[11469]_  | \new_[13736]_ ;
  assign \new_[9526]_  = ~\new_[11206]_  | ~\new_[18709]_ ;
  assign \new_[9527]_  = ~\new_[10801]_ ;
  assign \new_[9528]_  = ~\new_[19177]_  & (~\new_[13758]_  | ~\new_[15498]_ );
  assign \new_[9529]_  = \new_[11192]_  | \new_[11938]_ ;
  assign \new_[9530]_  = ~\new_[11125]_  | ~\new_[19553]_ ;
  assign \new_[9531]_  = ~\new_[13660]_  | ~\new_[10937]_ ;
  assign \new_[9532]_  = ~\new_[11471]_  | ~\new_[17070]_ ;
  assign \new_[9533]_  = ~\new_[11281]_  & ~\new_[19436]_ ;
  assign \new_[9534]_  = ~\new_[10936]_  | ~\new_[17146]_ ;
  assign \new_[9535]_  = ~\new_[10804]_ ;
  assign \new_[9536]_  = ~\new_[12320]_  & ~\new_[10899]_ ;
  assign \new_[9537]_  = ~\new_[18481]_  & (~\new_[13129]_  | ~\new_[13838]_ );
  assign \new_[9538]_  = ~\new_[19440]_  & (~\new_[13936]_  | ~\new_[12868]_ );
  assign \new_[9539]_  = ~\new_[11951]_  | ~\new_[12214]_ ;
  assign \new_[9540]_  = \new_[13763]_  & \new_[13661]_ ;
  assign \new_[9541]_  = ~\new_[17102]_  | ~\new_[14420]_  | ~\new_[15038]_ ;
  assign \new_[9542]_  = ~\new_[11119]_  | ~\new_[18187]_ ;
  assign \new_[9543]_  = ~\new_[19717]_  | (~\new_[16593]_  & ~\new_[15279]_ );
  assign \new_[9544]_  = ~\new_[19239]_  & (~\new_[13298]_  | ~\new_[17692]_ );
  assign \new_[9545]_  = ~\new_[11830]_  | ~\new_[11076]_ ;
  assign \new_[9546]_  = ~\new_[11175]_  | ~\new_[16683]_ ;
  assign \new_[9547]_  = ~\new_[11183]_  | ~\new_[19015]_ ;
  assign \new_[9548]_  = ~\new_[11399]_  & ~\new_[13815]_ ;
  assign \new_[9549]_  = ~\new_[14262]_  | ~\new_[11158]_ ;
  assign \new_[9550]_  = ~\new_[11124]_  | ~\new_[18998]_ ;
  assign \new_[9551]_  = \new_[12301]_  & \new_[12566]_ ;
  assign \new_[9552]_  = \new_[12206]_  & \new_[11828]_ ;
  assign \new_[9553]_  = ~\new_[10925]_  | ~\new_[14380]_ ;
  assign \new_[9554]_  = \new_[11273]_  & \new_[19239]_ ;
  assign \new_[9555]_  = ~\new_[19625]_  & (~\new_[13037]_  | ~\new_[15537]_ );
  assign \new_[9556]_  = ~\new_[11216]_  | ~\new_[19408]_ ;
  assign \new_[9557]_  = ~\new_[10840]_ ;
  assign \new_[9558]_  = ~\new_[18606]_  & (~\new_[13033]_  | ~\new_[16310]_ );
  assign \new_[9559]_  = ~\new_[10814]_ ;
  assign \new_[9560]_  = ~\new_[11275]_  | ~\new_[18228]_ ;
  assign \new_[9561]_  = ~\new_[11356]_  | ~\new_[11684]_ ;
  assign \new_[9562]_  = ~\new_[13630]_  | ~\new_[10904]_ ;
  assign \new_[9563]_  = ~\new_[10816]_ ;
  assign \new_[9564]_  = ~\new_[16448]_  & ~\new_[11238]_ ;
  assign \new_[9565]_  = \new_[11286]_  & \new_[19636]_ ;
  assign \new_[9566]_  = ~\new_[12360]_  & ~\new_[11125]_ ;
  assign \new_[9567]_  = ~\new_[11460]_  | ~\new_[18361]_ ;
  assign \new_[9568]_  = ~\new_[21073]_  | ~\new_[18361]_ ;
  assign \new_[9569]_  = ~\new_[11101]_  | ~\new_[19711]_ ;
  assign \new_[9570]_  = \new_[11270]_  & \new_[18194]_ ;
  assign \new_[9571]_  = ~\new_[11087]_  | ~\new_[11715]_ ;
  assign \new_[9572]_  = \new_[11043]_  & \new_[19366]_ ;
  assign \new_[9573]_  = ~\new_[11078]_  | ~\new_[20704]_ ;
  assign \new_[9574]_  = \new_[11193]_  & \new_[10959]_ ;
  assign \new_[9575]_  = \new_[11411]_  & \new_[19612]_ ;
  assign \new_[9576]_  = ~\new_[11106]_  | ~\new_[18941]_ ;
  assign \new_[9577]_  = ~\new_[11365]_  | ~\new_[18285]_ ;
  assign \new_[9578]_  = \\dcnt_reg[2] ;
  assign \new_[9579]_  = ~\new_[10958]_  | ~\new_[20341]_ ;
  assign \new_[9580]_  = ~\new_[18154]_  | (~\new_[13092]_  & ~\new_[16189]_ );
  assign \new_[9581]_  = ~\new_[11373]_  | ~\new_[13574]_ ;
  assign \new_[9582]_  = ~\new_[10905]_  | ~\new_[12223]_ ;
  assign \new_[9583]_  = ~\new_[19612]_  & (~\new_[12642]_  | ~\new_[14897]_ );
  assign \new_[9584]_  = ~\new_[12534]_  & ~\new_[11086]_ ;
  assign \new_[9585]_  = \new_[11023]_  & \new_[16237]_ ;
  assign \new_[9586]_  = ~\new_[11047]_  | ~\new_[15193]_ ;
  assign \new_[9587]_  = ~\new_[11226]_  | ~\new_[21562]_ ;
  assign \new_[9588]_  = ~\new_[10827]_ ;
  assign \new_[9589]_  = ~\new_[11192]_  | ~\new_[21115]_ ;
  assign \new_[9590]_  = ~\new_[10831]_ ;
  assign \new_[9591]_  = \new_[12239]_  & \new_[11955]_ ;
  assign \new_[9592]_  = ~\new_[10987]_  | ~\new_[13906]_ ;
  assign \new_[9593]_  = ~\new_[11240]_  | ~\new_[18682]_ ;
  assign \new_[9594]_  = ~\new_[10992]_  | ~\new_[11915]_ ;
  assign \new_[9595]_  = ~\new_[10835]_ ;
  assign \new_[9596]_  = ~\new_[11224]_  | ~\new_[18747]_ ;
  assign \new_[9597]_  = ~\new_[12369]_  | ~\new_[11620]_ ;
  assign \new_[9598]_  = ~\new_[11245]_  & ~\new_[13589]_ ;
  assign \new_[9599]_  = ~\new_[16907]_  | ~\new_[14178]_  | ~\new_[21714]_ ;
  assign \new_[9600]_  = ~\new_[10837]_ ;
  assign \new_[9601]_  = ~\new_[18070]_  & (~\new_[12989]_  | ~\new_[16322]_ );
  assign \new_[9602]_  = ~\new_[21136]_  | ~\new_[12418]_ ;
  assign \new_[9603]_  = \new_[12247]_  & \new_[14379]_ ;
  assign \new_[9604]_  = ~\new_[14729]_  | ~\new_[10918]_ ;
  assign \new_[9605]_  = ~\new_[10843]_ ;
  assign \new_[9606]_  = ~\new_[21555]_  | ~\new_[12249]_ ;
  assign \new_[9607]_  = ~\new_[11843]_  | ~\new_[12248]_ ;
  assign \new_[9608]_  = ~\new_[14312]_  & ~\new_[11257]_ ;
  assign \new_[9609]_  = ~\new_[10845]_ ;
  assign \new_[9610]_  = ~\new_[12818]_  | ~\new_[21661]_  | ~\new_[16370]_ ;
  assign \new_[9611]_  = ~\new_[11366]_  | ~\new_[13822]_ ;
  assign \new_[9612]_  = ~\new_[11009]_  & ~\new_[11632]_ ;
  assign \new_[9613]_  = ~\new_[20712]_  | ~\new_[13116]_ ;
  assign \new_[9614]_  = ~\new_[12367]_  | ~\new_[11635]_ ;
  assign \new_[9615]_  = ~\new_[11090]_  | ~\new_[19750]_ ;
  assign \new_[9616]_  = \new_[11170]_  | \new_[19145]_ ;
  assign \new_[9617]_  = ~\new_[19072]_  & (~\new_[13354]_  | ~\new_[14990]_ );
  assign \new_[9618]_  = ~\new_[12397]_  | ~\new_[11683]_ ;
  assign \new_[9619]_  = ~\new_[14141]_  | ~\new_[12210]_ ;
  assign \new_[9620]_  = ~\new_[12373]_  | ~\new_[20100]_ ;
  assign \new_[9621]_  = ~\new_[12397]_  & ~\new_[19687]_ ;
  assign \new_[9622]_  = ~\new_[12255]_  | ~\new_[13091]_ ;
  assign \new_[9623]_  = ~\new_[12444]_  | ~\new_[17472]_ ;
  assign \new_[9624]_  = ~\new_[13241]_  | ~\new_[12399]_ ;
  assign \new_[9625]_  = ~\new_[12287]_  & ~\new_[19587]_ ;
  assign \new_[9626]_  = ~\new_[20100]_  & (~\new_[14480]_  | ~\new_[15991]_ );
  assign \new_[9627]_  = ~\new_[14269]_  | ~\new_[12314]_ ;
  assign \new_[9628]_  = \new_[12379]_  | \new_[19299]_ ;
  assign \new_[9629]_  = ~\new_[12441]_  | ~\new_[17475]_ ;
  assign \new_[9630]_  = ~\new_[12910]_  | ~\new_[12239]_ ;
  assign \new_[9631]_  = ~\new_[21629]_  & (~\new_[14148]_  | ~\new_[15505]_ );
  assign \new_[9632]_  = \new_[12406]_  | \new_[18542]_ ;
  assign \new_[9633]_  = ~\new_[21142]_  | (~\new_[13493]_  & ~\new_[15152]_ );
  assign \new_[9634]_  = ~\new_[13589]_  & ~\new_[12335]_ ;
  assign \new_[9635]_  = ~\new_[19299]_  & (~\new_[13598]_  | ~\new_[13694]_ );
  assign \new_[9636]_  = ~\new_[12369]_  & ~\new_[16879]_ ;
  assign \new_[9637]_  = ~\new_[16207]_  | ~\new_[12380]_ ;
  assign \new_[9638]_  = ~\new_[14342]_  | ~\new_[12384]_ ;
  assign \new_[9639]_  = ~\new_[12233]_  | ~\new_[12845]_ ;
  assign \new_[9640]_  = ~\new_[12394]_  & ~\new_[18937]_ ;
  assign \new_[9641]_  = ~\new_[15334]_  | ~\new_[12232]_ ;
  assign \new_[9642]_  = ~\new_[13837]_  | ~\new_[12738]_  | ~\new_[14301]_ ;
  assign \new_[9643]_  = ~\new_[12378]_  & ~\new_[19006]_ ;
  assign \new_[9644]_  = ~\new_[13652]_  | ~\new_[13321]_ ;
  assign \new_[9645]_  = ~\new_[12378]_  | ~\new_[14588]_ ;
  assign \new_[9646]_  = \new_[12387]_  & \new_[13785]_ ;
  assign \new_[9647]_  = ~\new_[12387]_  & ~\new_[19028]_ ;
  assign \new_[9648]_  = ~\new_[14000]_  | ~\new_[13549]_ ;
  assign \new_[9649]_  = ~\new_[19059]_  & (~\new_[13842]_  | ~\new_[14207]_ );
  assign \new_[9650]_  = ~\new_[12259]_  | ~\new_[13190]_ ;
  assign \new_[9651]_  = ~\new_[13733]_  & ~\new_[12440]_ ;
  assign \new_[9652]_  = ~\new_[10851]_ ;
  assign \new_[9653]_  = ~\new_[19094]_  & (~\new_[13988]_  | ~\new_[14163]_ );
  assign \new_[9654]_  = ~\new_[21407]_  & ~\new_[12401]_ ;
  assign \new_[9655]_  = ~\new_[16359]_  & ~\new_[12337]_ ;
  assign \new_[9656]_  = ~\new_[12256]_  | ~\new_[14952]_ ;
  assign \new_[9657]_  = ~\new_[15974]_  & ~\new_[12374]_ ;
  assign \new_[9658]_  = ~\new_[19592]_  & (~\new_[13827]_  | ~\new_[13645]_ );
  assign \new_[9659]_  = ~\new_[10854]_ ;
  assign \new_[9660]_  = ~\new_[12266]_  | ~\new_[14129]_ ;
  assign \new_[9661]_  = ~\new_[12255]_  | ~\new_[14192]_ ;
  assign \new_[9662]_  = ~\new_[12229]_  | ~\new_[12959]_ ;
  assign \new_[9663]_  = ~\new_[18249]_  & (~\new_[14670]_  | ~\new_[15381]_ );
  assign \new_[9664]_  = ~\new_[12328]_  | ~\new_[19208]_ ;
  assign \new_[9665]_  = \new_[12474]_  | \new_[19512]_ ;
  assign \new_[9666]_  = \new_[12452]_  & \new_[19021]_ ;
  assign \new_[9667]_  = ~\new_[20864]_  | ~\new_[18821]_ ;
  assign \new_[9668]_  = ~\new_[21115]_  & (~\new_[13956]_  | ~\new_[16195]_ );
  assign \new_[9669]_  = ~\new_[12963]_  | ~\new_[12304]_ ;
  assign \new_[9670]_  = \new_[12295]_  | \new_[19064]_ ;
  assign \new_[9671]_  = ~\new_[12282]_  | ~\new_[15714]_ ;
  assign \new_[9672]_  = ~\new_[13370]_  & ~\new_[18605]_ ;
  assign \new_[9673]_  = ~\new_[10857]_ ;
  assign \new_[9674]_  = ~\new_[15253]_  | ~\new_[14197]_  | ~\new_[15198]_ ;
  assign \new_[9675]_  = ~\new_[19625]_  & (~\new_[13974]_  | ~\new_[16259]_ );
  assign \new_[9676]_  = ~\new_[12310]_  & ~\new_[18569]_ ;
  assign \new_[9677]_  = ~\new_[19727]_  & (~\new_[14032]_  | ~\new_[15702]_ );
  assign \new_[9678]_  = ~\new_[12409]_  | ~\new_[19021]_ ;
  assign \new_[9679]_  = ~\new_[12315]_  | ~\new_[19233]_ ;
  assign \new_[9680]_  = ~\new_[12301]_  & ~\new_[18941]_ ;
  assign \new_[9681]_  = ~\new_[14809]_  | ~\new_[13961]_  | ~\new_[13982]_ ;
  assign \new_[9682]_  = ~\new_[12183]_  | ~\new_[21406]_ ;
  assign \new_[9683]_  = ~\new_[12475]_  | ~\new_[19145]_ ;
  assign \new_[9684]_  = ~\new_[12477]_  & ~\new_[12446]_ ;
  assign \new_[9685]_  = ~\new_[13910]_  | ~\new_[12505]_  | ~\new_[15071]_ ;
  assign \new_[9686]_  = ~\new_[18361]_  & (~\new_[14440]_  | ~\new_[15143]_ );
  assign \new_[9687]_  = ~\new_[14000]_  | ~\new_[12560]_  | ~\new_[15563]_ ;
  assign \new_[9688]_  = ~\new_[14149]_  | ~\new_[12555]_  | ~\new_[14792]_ ;
  assign \new_[9689]_  = ~\new_[15337]_  | ~\new_[12539]_  | ~\new_[16011]_ ;
  assign \new_[9690]_  = ~\new_[14227]_  | ~\new_[13923]_  | ~\new_[15986]_ ;
  assign \new_[9691]_  = ~\new_[10847]_ ;
  assign \new_[9692]_  = ~\new_[19161]_  & (~\new_[15452]_  | ~\new_[14083]_ );
  assign \new_[9693]_  = ~\new_[12388]_  & ~\new_[12809]_ ;
  assign \new_[9694]_  = ~\new_[14424]_  | ~\new_[13720]_  | ~\new_[13625]_ ;
  assign \new_[9695]_  = ~\new_[16840]_  & (~\new_[14916]_  | ~\new_[16143]_ );
  assign \new_[9696]_  = ~\new_[12356]_  | ~\new_[19145]_ ;
  assign \new_[9697]_  = ~\new_[14042]_  | ~\new_[14990]_  | ~\new_[13825]_ ;
  assign \new_[9698]_  = ~\new_[19240]_  & (~\new_[14007]_  | ~\new_[14693]_ );
  assign \new_[9699]_  = ~\new_[12318]_  | (~\new_[17785]_  & ~\new_[18076]_ );
  assign \new_[9700]_  = ~\new_[18194]_  & (~\new_[17616]_  | ~\new_[14315]_ );
  assign \new_[9701]_  = ~\new_[15225]_  | ~\new_[13560]_  | ~\new_[14315]_ ;
  assign \new_[9702]_  = \new_[12341]_  & \new_[18076]_ ;
  assign \new_[9703]_  = ~\new_[17064]_  & (~\new_[14131]_  | ~\new_[16507]_ );
  assign \new_[9704]_  = ~\new_[16145]_  | ~\new_[17366]_  | ~\new_[13685]_ ;
  assign \new_[9705]_  = ~\new_[10860]_ ;
  assign \new_[9706]_  = ~\new_[13728]_  | ~\new_[12181]_ ;
  assign \new_[9707]_  = ~\new_[12228]_  | ~\new_[13552]_ ;
  assign \new_[9708]_  = \new_[12459]_  & \new_[19547]_ ;
  assign \new_[9709]_  = ~\new_[15281]_  | ~\new_[13667]_  | ~\new_[14380]_ ;
  assign \new_[9710]_  = ~\new_[19239]_  & (~\new_[17097]_  | ~\new_[14591]_ );
  assign \new_[9711]_  = ~\new_[17146]_  | ~\new_[13660]_  | ~\new_[13705]_ ;
  assign \new_[9712]_  = ~\new_[16235]_  | ~\new_[15716]_  | ~\new_[13681]_ ;
  assign \new_[9713]_  = ~\new_[18187]_  & (~\new_[14242]_  | ~\new_[17057]_ );
  assign \new_[9714]_  = ~\new_[21328]_  & (~\new_[16703]_  | ~\new_[13719]_ );
  assign \new_[9715]_  = \new_[12364]_  & \new_[19366]_ ;
  assign \new_[9716]_  = ~\new_[15063]_  | ~\new_[12211]_ ;
  assign \new_[9717]_  = ~\new_[19502]_  | ~\new_[16646]_  | ~\new_[13736]_ ;
  assign \new_[9718]_  = ~\new_[21557]_  & (~\new_[13992]_  | ~\new_[15386]_ );
  assign \new_[9719]_  = ~\new_[18486]_  | ~\new_[17863]_  | ~\new_[14102]_ ;
  assign \new_[9720]_  = ~\new_[15066]_  | ~\new_[12223]_ ;
  assign \new_[9721]_  = ~\new_[12245]_  | ~\new_[12221]_ ;
  assign \new_[9722]_  = ~\new_[10865]_ ;
  assign \new_[9723]_  = ~\new_[10866]_ ;
  assign \new_[9724]_  = ~\new_[16266]_  | ~\new_[13630]_  | ~\new_[16192]_ ;
  assign \new_[9725]_  = ~\new_[18965]_  & (~\new_[16292]_  | ~\new_[14199]_ );
  assign \new_[9726]_  = ~\new_[19102]_  & (~\new_[15459]_  | ~\new_[14074]_ );
  assign \new_[9727]_  = ~\new_[12348]_  | ~\new_[21562]_ ;
  assign \new_[9728]_  = ~\new_[16796]_  | ~\new_[14582]_  | ~\new_[14305]_ ;
  assign \new_[9729]_  = ~\new_[13996]_  | ~\new_[13884]_  | ~\new_[14895]_ ;
  assign \new_[9730]_  = ~\new_[10867]_ ;
  assign \new_[9731]_  = ~\new_[13906]_  | ~\new_[12379]_  | ~\new_[14264]_ ;
  assign \new_[9732]_  = ~\new_[19006]_  & (~\new_[17173]_  | ~\new_[14244]_ );
  assign \new_[9733]_  = ~\new_[19028]_  & (~\new_[15437]_  | ~\new_[14014]_ );
  assign \new_[9734]_  = ~\new_[17457]_  & (~\new_[15390]_  | ~\new_[13709]_ );
  assign \new_[9735]_  = ~\new_[21638]_  & (~\new_[13494]_  | ~\new_[17083]_ );
  assign \new_[9736]_  = ~\new_[20099]_  & (~\new_[13682]_  | ~\new_[14876]_ );
  assign \new_[9737]_  = ~\new_[15520]_  | ~\new_[12380]_ ;
  assign \new_[9738]_  = ~\new_[15414]_  | ~\new_[12384]_ ;
  assign \new_[9739]_  = ~\new_[19094]_  & (~\new_[14161]_  | ~\new_[17503]_ );
  assign \new_[9740]_  = ~\new_[21631]_  & (~\new_[20926]_  | ~\new_[14296]_ );
  assign \new_[9741]_  = ~\new_[13498]_  | ~\new_[17231]_  | ~\new_[13963]_ ;
  assign \new_[9742]_  = ~\new_[10868]_ ;
  assign \new_[9743]_  = ~\new_[18538]_  | (~\new_[14408]_  & ~\new_[15170]_ );
  assign \new_[9744]_  = ~\new_[12603]_  | ~\new_[12229]_ ;
  assign \new_[9745]_  = ~\new_[13169]_  | ~\new_[12260]_ ;
  assign \new_[9746]_  = ~\new_[14382]_  | ~\new_[15029]_  | ~\new_[15598]_ ;
  assign \new_[9747]_  = ~\new_[18494]_  | (~\new_[14413]_  & ~\new_[15435]_ );
  assign \new_[9748]_  = ~\new_[13764]_  | ~\new_[12255]_ ;
  assign \new_[9749]_  = ~\new_[12819]_  | ~\new_[12233]_ ;
  assign \new_[9750]_  = ~\new_[21638]_  & (~\new_[17757]_  | ~\new_[13804]_ );
  assign \new_[9751]_  = ~\new_[10869]_ ;
  assign \new_[9752]_  = ~\new_[15551]_  | ~\new_[12304]_ ;
  assign \new_[9753]_  = ~\new_[21562]_  & (~\new_[14452]_  | ~\new_[14629]_ );
  assign \new_[9754]_  = ~\new_[15863]_  | ~\new_[12390]_ ;
  assign \new_[9755]_  = ~\new_[19266]_  & (~\new_[15393]_  | ~\new_[14165]_ );
  assign \new_[9756]_  = ~\new_[15301]_  & ~\new_[12207]_ ;
  assign \new_[9757]_  = ~\new_[19727]_  & (~\new_[17722]_  | ~\new_[14378]_ );
  assign \new_[9758]_  = ~\new_[14609]_  | ~\new_[15127]_  | ~\new_[13961]_ ;
  assign \new_[9759]_  = ~\new_[19587]_  & (~\new_[14213]_  | ~\new_[17068]_ );
  assign \new_[9760]_  = ~\new_[12303]_  | (~\new_[16642]_  & ~\new_[18166]_ );
  assign \new_[9761]_  = ~\new_[21513]_  & (~\new_[16298]_  | ~\new_[13755]_ );
  assign \new_[9762]_  = ~\new_[10870]_ ;
  assign \new_[9763]_  = ~\new_[14375]_  | ~\new_[13972]_  | ~\new_[13762]_ ;
  assign \new_[9764]_  = ~\new_[19261]_  & (~\new_[14003]_  | ~\new_[15409]_ );
  assign \new_[9765]_  = ~\new_[14120]_  | ~\new_[13620]_  | ~\new_[16256]_ ;
  assign \new_[9766]_  = ~\new_[12881]_  | (~\new_[15584]_  & ~\new_[18984]_ );
  assign \new_[9767]_  = \new_[12345]_  | \new_[18833]_ ;
  assign \new_[9768]_  = ~\new_[12288]_  | ~\new_[18262]_ ;
  assign \new_[9769]_  = ~\new_[15939]_  | ~\new_[15143]_  | ~\new_[13801]_ ;
  assign \new_[9770]_  = ~\new_[15597]_  | ~\new_[12399]_ ;
  assign \new_[9771]_  = ~\new_[19553]_  & (~\new_[14093]_  | ~\new_[16162]_ );
  assign \new_[9772]_  = ~\new_[14906]_  | ~\new_[12254]_ ;
  assign \new_[9773]_  = ~\new_[12962]_  | (~\new_[14102]_  & ~\new_[19408]_ );
  assign \new_[9774]_  = ~\new_[15187]_  | ~\new_[12317]_ ;
  assign \new_[9775]_  = ~\new_[12191]_  & (~\new_[17990]_  | ~\new_[18402]_ );
  assign \new_[9776]_  = \new_[14190]_  ? \new_[19206]_  : \new_[15347]_ ;
  assign \new_[9777]_  = ~\new_[13131]_  | (~\new_[15246]_  & ~\new_[18906]_ );
  assign \new_[9778]_  = ~\new_[15303]_  | (~\new_[14434]_  & ~\new_[21574]_ );
  assign \new_[9779]_  = ~\new_[13202]_  | (~\new_[13993]_  & ~\new_[18587]_ );
  assign \new_[9780]_  = ~\new_[15362]_  | (~\new_[14398]_  & ~\new_[18394]_ );
  assign \new_[9781]_  = ~\new_[14945]_  | (~\new_[14155]_  & ~\new_[17886]_ );
  assign \new_[9782]_  = ~\new_[12186]_  & (~\new_[18910]_  | ~\new_[18170]_ );
  assign \new_[9783]_  = ~\new_[12273]_  & (~\new_[17734]_  | ~\new_[18082]_ );
  assign \new_[9784]_  = \new_[14545]_  ? \new_[19625]_  : \new_[16259]_ ;
  assign \new_[9785]_  = \new_[14003]_  ? \new_[18863]_  : \new_[16671]_ ;
  assign \new_[9786]_  = ~\new_[12558]_  | (~\new_[14949]_  & ~\new_[19253]_ );
  assign \new_[9787]_  = \new_[12912]_  & \new_[19288]_ ;
  assign \new_[9788]_  = ~\new_[13335]_  & (~\new_[16931]_  | ~\new_[21483]_ );
  assign \new_[9789]_  = ~\new_[12893]_  & (~\new_[14560]_  | ~\new_[17954]_ );
  assign \new_[9790]_  = \new_[14640]_  & \new_[12996]_ ;
  assign \new_[9791]_  = ~\new_[13045]_  | ~\new_[19233]_ ;
  assign \new_[9792]_  = ~\new_[14139]_  & (~\new_[14563]_  | ~\new_[18262]_ );
  assign \new_[9793]_  = ~\new_[13086]_  & (~\new_[15697]_  | ~\new_[17536]_ );
  assign \new_[9794]_  = ~\new_[10881]_ ;
  assign \new_[9795]_  = ~\new_[12340]_  & (~\new_[13657]_  | ~\new_[17488]_ );
  assign \new_[9796]_  = ~\new_[13482]_  | ~\new_[19015]_ ;
  assign \new_[9797]_  = ~\new_[10885]_ ;
  assign \new_[9798]_  = ~\new_[10886]_ ;
  assign \new_[9799]_  = ~\new_[12828]_  | ~\new_[19015]_ ;
  assign \new_[9800]_  = ~\new_[12601]_  & ~\new_[19547]_ ;
  assign \new_[9801]_  = ~\new_[17349]_  | ~\new_[18596]_  | ~\new_[19266]_  | ~\new_[18434]_ ;
  assign \new_[9802]_  = ~\new_[12537]_  & ~\new_[18984]_ ;
  assign \new_[9803]_  = ~\new_[10890]_ ;
  assign \new_[9804]_  = ~\new_[10891]_ ;
  assign \new_[9805]_  = ~\new_[10892]_ ;
  assign \new_[9806]_  = ~\new_[10893]_ ;
  assign \new_[9807]_  = ~\new_[12932]_  | ~\new_[20239]_ ;
  assign \new_[9808]_  = \new_[12823]_  | \new_[19151]_ ;
  assign \new_[9809]_  = \new_[13282]_  | \new_[19474]_ ;
  assign \new_[9810]_  = ~\new_[10895]_ ;
  assign \new_[9811]_  = ~\new_[10898]_ ;
  assign \new_[9812]_  = ~\new_[10899]_ ;
  assign \new_[9813]_  = ~\new_[12533]_  | ~\new_[18187]_ ;
  assign \new_[9814]_  = \new_[12589]_  & \new_[18832]_ ;
  assign \new_[9815]_  = ~\new_[13362]_  | ~\new_[18209]_ ;
  assign \new_[9816]_  = ~\new_[19547]_  | ~\new_[13770]_ ;
  assign \new_[9817]_  = ~\new_[10906]_ ;
  assign \new_[9818]_  = ~\new_[10906]_ ;
  assign \new_[9819]_  = ~\new_[18443]_  & ~\new_[13041]_ ;
  assign \new_[9820]_  = ~\new_[10908]_ ;
  assign \new_[9821]_  = ~\new_[10910]_ ;
  assign \new_[9822]_  = ~\new_[12899]_  | ~\new_[18414]_ ;
  assign \new_[9823]_  = ~\new_[10913]_ ;
  assign \new_[9824]_  = \new_[12446]_  & \new_[18414]_ ;
  assign \new_[9825]_  = \new_[13003]_  & \new_[19261]_ ;
  assign \new_[9826]_  = ~\new_[12932]_  | ~\new_[18288]_ ;
  assign \new_[9827]_  = ~\new_[12490]_  | ~\new_[18443]_ ;
  assign \new_[9828]_  = ~\new_[12867]_  | ~\new_[18832]_ ;
  assign \new_[9829]_  = ~\new_[10919]_ ;
  assign \new_[9830]_  = ~\new_[10923]_ ;
  assign \new_[9831]_  = ~\new_[10923]_ ;
  assign \new_[9832]_  = ~\new_[10924]_ ;
  assign \new_[9833]_  = ~\new_[12904]_  | ~\new_[18832]_ ;
  assign \new_[9834]_  = ~\new_[10927]_ ;
  assign \new_[9835]_  = \new_[13472]_  & \new_[19589]_ ;
  assign \new_[9836]_  = ~\new_[10928]_ ;
  assign \new_[9837]_  = ~\new_[10930]_ ;
  assign \new_[9838]_  = ~\new_[13289]_  | ~\new_[21689]_ ;
  assign \new_[9839]_  = ~\new_[12589]_  | ~\new_[19547]_ ;
  assign \new_[9840]_  = ~\new_[20713]_  & ~\new_[19208]_ ;
  assign \new_[9841]_  = \new_[21163]_  & \new_[18280]_ ;
  assign \new_[9842]_  = ~\new_[10938]_ ;
  assign \new_[9843]_  = ~\new_[10940]_ ;
  assign \new_[9844]_  = ~\new_[13186]_  | ~\new_[19217]_ ;
  assign \new_[9845]_  = ~\new_[10943]_ ;
  assign \new_[9846]_  = ~\new_[12164]_  | ~\new_[18209]_ ;
  assign \new_[9847]_  = ~\new_[12196]_  | ~\new_[19115]_ ;
  assign \new_[9848]_  = ~\new_[12744]_  | ~\new_[19088]_ ;
  assign \new_[9849]_  = ~\new_[10947]_ ;
  assign \new_[9850]_  = ~\new_[12167]_  | ~\new_[19102]_ ;
  assign \new_[9851]_  = ~\new_[10950]_ ;
  assign \new_[9852]_  = ~\new_[13952]_  & ~\new_[18998]_ ;
  assign \new_[9853]_  = ~\new_[18012]_  | ~\new_[19018]_  | ~\new_[16321]_ ;
  assign \new_[9854]_  = ~\new_[13187]_  & ~\new_[21638]_ ;
  assign \new_[9855]_  = ~\new_[12220]_  | ~\new_[19290]_ ;
  assign \new_[9856]_  = ~\new_[12791]_  | ~\new_[19381]_ ;
  assign \new_[9857]_  = ~\new_[10957]_ ;
  assign \new_[9858]_  = ~\new_[10958]_ ;
  assign \new_[9859]_  = ~\new_[12538]_  | ~\new_[19711]_ ;
  assign \new_[9860]_  = ~\new_[15209]_  | ~\new_[18847]_  | ~\new_[17922]_ ;
  assign \new_[9861]_  = ~\new_[10961]_ ;
  assign \new_[9862]_  = ~\new_[10961]_ ;
  assign \new_[9863]_  = \new_[19239]_  & \new_[12679]_ ;
  assign \new_[9864]_  = ~\new_[12562]_  | ~\new_[21558]_ ;
  assign \new_[9865]_  = ~\new_[13121]_  | ~\new_[19233]_ ;
  assign \new_[9866]_  = \new_[13046]_  | \new_[21513]_ ;
  assign \new_[9867]_  = ~\new_[10970]_ ;
  assign \new_[9868]_  = ~\new_[13791]_  | ~\new_[18621]_ ;
  assign \new_[9869]_  = ~\new_[10975]_ ;
  assign \new_[9870]_  = ~\new_[18974]_  | ~\new_[19094]_  | ~\new_[16168]_ ;
  assign \new_[9871]_  = ~\new_[15803]_  | ~\new_[19245]_  | ~\new_[18678]_  | ~\new_[18587]_ ;
  assign \new_[9872]_  = ~\new_[13007]_  | ~\new_[18605]_ ;
  assign \new_[9873]_  = ~\new_[10976]_ ;
  assign \new_[9874]_  = ~\new_[10977]_ ;
  assign \new_[9875]_  = ~\new_[10978]_ ;
  assign \new_[9876]_  = ~\new_[10979]_ ;
  assign \new_[9877]_  = \new_[12504]_  | \new_[19381]_ ;
  assign \new_[9878]_  = ~\new_[10980]_ ;
  assign \new_[9879]_  = ~\new_[10982]_ ;
  assign \new_[9880]_  = ~\new_[12527]_  | ~\new_[18427]_ ;
  assign \new_[9881]_  = ~\new_[18811]_  | ~\new_[18692]_  | ~\new_[15970]_ ;
  assign \new_[9882]_  = ~\new_[10983]_ ;
  assign \new_[9883]_  = ~\new_[10984]_ ;
  assign \new_[9884]_  = \new_[12361]_  & \new_[21115]_ ;
  assign \new_[9885]_  = ~\new_[13052]_  | ~\new_[19071]_ ;
  assign \new_[9886]_  = ~\new_[12468]_  & ~\new_[19275]_ ;
  assign \new_[9887]_  = ~\new_[15848]_  | ~\new_[18855]_ ;
  assign \new_[9888]_  = ~\new_[12929]_  & ~\new_[19275]_ ;
  assign \new_[9889]_  = ~\new_[10985]_ ;
  assign \new_[9890]_  = ~\new_[12723]_  & ~\new_[18076]_ ;
  assign \new_[9891]_  = ~\new_[14544]_  & ~\new_[19094]_  & ~\new_[17658]_ ;
  assign \new_[9892]_  = ~\new_[13186]_  | ~\new_[19233]_ ;
  assign \new_[9893]_  = ~\new_[12638]_  | ~\new_[19217]_ ;
  assign \new_[9894]_  = ~\new_[18770]_  & ~\new_[18060]_  & ~\new_[20099]_  & ~\new_[18501]_ ;
  assign \new_[9895]_  = ~\new_[12167]_  | ~\new_[18325]_ ;
  assign \new_[9896]_  = ~\new_[10988]_ ;
  assign \new_[9897]_  = ~\new_[10989]_ ;
  assign \new_[9898]_  = ~\new_[10990]_ ;
  assign \new_[9899]_  = ~\new_[10992]_ ;
  assign \new_[9900]_  = ~\new_[10995]_ ;
  assign \new_[9901]_  = ~\new_[10995]_ ;
  assign \new_[9902]_  = ~\new_[10996]_ ;
  assign \new_[9903]_  = ~\new_[11000]_ ;
  assign \new_[9904]_  = ~\new_[10528]_  | ~\new_[19204]_ ;
  assign \new_[9905]_  = ~\new_[11001]_ ;
  assign \new_[9906]_  = ~\new_[11003]_ ;
  assign \new_[9907]_  = ~\new_[11005]_ ;
  assign \new_[9908]_  = ~\new_[12905]_  | ~\new_[18969]_ ;
  assign \new_[9909]_  = \new_[12515]_  | \new_[19266]_ ;
  assign \new_[9910]_  = ~\new_[12522]_  & (~\new_[15836]_  | ~\new_[18984]_ );
  assign \new_[9911]_  = ~\new_[12891]_  | ~\new_[18840]_ ;
  assign \new_[9912]_  = ~\new_[13108]_  & ~\new_[21634]_ ;
  assign \new_[9913]_  = ~\new_[13364]_  | ~\new_[19018]_ ;
  assign \new_[9914]_  = ~\new_[13273]_  | ~\new_[19587]_ ;
  assign \new_[9915]_  = ~\new_[11010]_ ;
  assign \new_[9916]_  = ~\new_[11010]_ ;
  assign \new_[9917]_  = ~\new_[10597]_  | ~\new_[20485]_ ;
  assign \new_[9918]_  = ~\new_[13007]_  | ~\new_[18847]_ ;
  assign \new_[9919]_  = \new_[12737]_  | \new_[18847]_ ;
  assign \new_[9920]_  = ~\new_[11011]_ ;
  assign \new_[9921]_  = ~\new_[13155]_  | ~\new_[19275]_ ;
  assign \new_[9922]_  = ~\new_[21396]_  | ~\new_[19681]_  | ~\new_[16095]_ ;
  assign \new_[9923]_  = ~\new_[11012]_ ;
  assign \new_[9924]_  = ~\new_[12759]_  | ~\new_[19006]_ ;
  assign \new_[9925]_  = ~\new_[18984]_  & ~\new_[12870]_ ;
  assign \new_[9926]_  = ~\new_[12512]_  | ~\new_[20680]_ ;
  assign \new_[9927]_  = ~\new_[11016]_ ;
  assign \new_[9928]_  = ~\new_[11017]_ ;
  assign \new_[9929]_  = ~\new_[12420]_  | ~\new_[19215]_ ;
  assign \new_[9930]_  = ~\new_[11018]_ ;
  assign \new_[9931]_  = \new_[12577]_  & \new_[19153]_ ;
  assign \new_[9932]_  = ~\new_[11019]_ ;
  assign \new_[9933]_  = \new_[12412]_  & \new_[21558]_ ;
  assign \new_[9934]_  = ~\new_[12877]_  & ~\new_[18621]_ ;
  assign \new_[9935]_  = ~\new_[12706]_  | ~\new_[21558]_ ;
  assign \new_[9936]_  = ~\new_[12905]_  | ~\new_[19299]_ ;
  assign \new_[9937]_  = ~\new_[12493]_  | ~\new_[17457]_ ;
  assign \new_[9938]_  = \new_[20906]_  | \new_[18077]_ ;
  assign \new_[9939]_  = ~\new_[11022]_ ;
  assign \new_[9940]_  = ~\new_[13364]_  | ~\new_[21634]_ ;
  assign \new_[9941]_  = ~\new_[14665]_  | ~\new_[19625]_  | ~\new_[18584]_ ;
  assign \new_[9942]_  = ~\new_[21662]_  | ~\new_[17358]_ ;
  assign \new_[9943]_  = ~\new_[21390]_  | ~\new_[18747]_ ;
  assign \new_[9944]_  = ~\new_[12433]_  | ~\new_[19462]_ ;
  assign \new_[9945]_  = \new_[13155]_  & \new_[21562]_ ;
  assign \new_[9946]_  = ~\new_[20218]_  & ~\new_[21558]_ ;
  assign \new_[9947]_  = ~\new_[11024]_ ;
  assign \new_[9948]_  = ~\new_[12617]_  | ~\new_[19450]_ ;
  assign \new_[9949]_  = ~\new_[11026]_ ;
  assign \new_[9950]_  = ~\new_[12491]_  & ~\new_[21635]_ ;
  assign \new_[9951]_  = ~\new_[21297]_ ;
  assign \new_[9952]_  = ~\new_[11028]_ ;
  assign \new_[9953]_  = ~\new_[11028]_ ;
  assign \new_[9954]_  = ~\new_[11033]_ ;
  assign \new_[9955]_  = ~\new_[12570]_  | ~\new_[18994]_ ;
  assign \new_[9956]_  = ~\new_[12488]_  | ~\new_[19687]_ ;
  assign \new_[9957]_  = ~\new_[12935]_  & ~\new_[19450]_ ;
  assign \new_[9958]_  = ~\new_[12527]_  | ~\new_[21115]_ ;
  assign \new_[9959]_  = ~\new_[11035]_ ;
  assign \new_[9960]_  = ~\new_[11037]_ ;
  assign \new_[9961]_  = ~\new_[11038]_ ;
  assign \new_[9962]_  = ~\new_[11040]_ ;
  assign \new_[9963]_  = ~\new_[11042]_ ;
  assign \new_[9964]_  = ~\new_[11043]_ ;
  assign \new_[9965]_  = ~\new_[12626]_  | ~\new_[19625]_ ;
  assign \new_[9966]_  = ~\new_[11044]_ ;
  assign \new_[9967]_  = ~\new_[13173]_  & ~\new_[18421]_ ;
  assign \new_[9968]_  = ~\new_[12596]_  & ~\new_[18187]_ ;
  assign \new_[9969]_  = ~\new_[21601]_  | ~\new_[18228]_ ;
  assign \new_[9970]_  = ~\new_[11048]_ ;
  assign \new_[9971]_  = ~\new_[12506]_  | ~\new_[21115]_ ;
  assign \new_[9972]_  = \new_[12565]_  & \new_[19319]_ ;
  assign \new_[9973]_  = ~\new_[11050]_ ;
  assign \new_[9974]_  = ~\new_[11051]_ ;
  assign \new_[9975]_  = ~\new_[12794]_  | ~\new_[19161]_ ;
  assign \new_[9976]_  = ~\new_[13261]_  | ~\new_[18228]_ ;
  assign \new_[9977]_  = ~\new_[11052]_ ;
  assign \new_[9978]_  = ~\new_[13014]_  | ~\new_[18692]_ ;
  assign \new_[9979]_  = ~\new_[14679]_  | ~\new_[17469]_ ;
  assign \new_[9980]_  = ~\new_[11053]_ ;
  assign \new_[9981]_  = ~\new_[13263]_  | ~\new_[19265]_ ;
  assign \new_[9982]_  = \new_[12657]_  | \new_[14951]_ ;
  assign \new_[9983]_  = ~\new_[11054]_ ;
  assign \new_[9984]_  = ~\new_[11055]_ ;
  assign \new_[9985]_  = ~\new_[11057]_ ;
  assign \new_[9986]_  = \new_[12797]_  & \new_[19156]_ ;
  assign \new_[9987]_  = \new_[12941]_  | \new_[19088]_ ;
  assign \new_[9988]_  = ~\new_[11059]_ ;
  assign \new_[9989]_  = ~\new_[12661]_  | ~\new_[21562]_ ;
  assign \new_[9990]_  = ~\new_[11060]_ ;
  assign \new_[9991]_  = ~\new_[11062]_ ;
  assign \new_[9992]_  = ~\new_[11063]_ ;
  assign \new_[9993]_  = ~\new_[11065]_ ;
  assign \new_[9994]_  = ~\new_[12750]_  | ~\new_[18361]_ ;
  assign \new_[9995]_  = ~\new_[13472]_  | ~\new_[19288]_ ;
  assign \new_[9996]_  = ~\new_[13294]_  & ~\new_[21693]_ ;
  assign \new_[9997]_  = ~\new_[11068]_ ;
  assign \new_[9998]_  = ~\new_[12791]_  | ~\new_[21689]_ ;
  assign \new_[9999]_  = ~\new_[11070]_ ;
  assign \new_[10000]_  = ~\new_[11072]_ ;
  assign \new_[10001]_  = \new_[13080]_  | \new_[17469]_ ;
  assign \new_[10002]_  = ~\new_[11074]_ ;
  assign \new_[10003]_  = ~\new_[16309]_  | ~\new_[15758]_ ;
  assign \new_[10004]_  = ~\new_[11075]_ ;
  assign \new_[10005]_  = ~\new_[12655]_  | ~\new_[21508]_ ;
  assign \new_[10006]_  = ~\new_[11077]_ ;
  assign \new_[10007]_  = ~\new_[11078]_ ;
  assign \new_[10008]_  = ~\new_[12555]_  | ~\new_[13562]_ ;
  assign \new_[10009]_  = ~\new_[12670]_  & ~\new_[19151]_ ;
  assign \new_[10010]_  = ~\new_[15567]_  | ~\new_[19130]_ ;
  assign \new_[10011]_  = ~\new_[12990]_  | ~\new_[14588]_ ;
  assign \new_[10012]_  = ~\new_[12833]_  & ~\new_[15322]_ ;
  assign \new_[10013]_  = ~\new_[11085]_ ;
  assign \new_[10014]_  = ~\new_[12501]_  | ~\new_[18967]_ ;
  assign \new_[10015]_  = ~\new_[16521]_  | ~\new_[12975]_ ;
  assign \new_[10016]_  = ~\new_[11088]_ ;
  assign \new_[10017]_  = ~\new_[12735]_  | ~\new_[17780]_ ;
  assign \new_[10018]_  = ~\new_[15359]_  | ~\new_[12859]_ ;
  assign \new_[10019]_  = ~\new_[11094]_ ;
  assign \new_[10020]_  = ~\new_[11095]_ ;
  assign \new_[10021]_  = ~\new_[11098]_ ;
  assign \new_[10022]_  = ~\new_[13352]_  & ~\new_[15389]_ ;
  assign \new_[10023]_  = ~\new_[16174]_  | ~\new_[18443]_ ;
  assign \new_[10024]_  = ~\new_[18270]_  | ~\new_[13343]_ ;
  assign \new_[10025]_  = ~\new_[11100]_ ;
  assign \new_[10026]_  = ~\new_[14973]_  | ~\new_[12520]_ ;
  assign \new_[10027]_  = ~\new_[14015]_  | ~\new_[12895]_ ;
  assign \new_[10028]_  = ~\new_[11103]_ ;
  assign \new_[10029]_  = ~\new_[12858]_  & ~\new_[18008]_ ;
  assign \new_[10030]_  = ~\new_[12860]_  | ~\new_[18693]_ ;
  assign \new_[10031]_  = ~\new_[12622]_  & ~\new_[18930]_ ;
  assign \new_[10032]_  = ~\new_[12524]_  & ~\new_[19141]_ ;
  assign \new_[10033]_  = ~\new_[14204]_  & ~\new_[12894]_ ;
  assign \new_[10034]_  = ~\new_[11109]_ ;
  assign \new_[10035]_  = ~\new_[13129]_  | ~\new_[15377]_ ;
  assign \new_[10036]_  = ~\new_[17999]_  & ~\new_[12978]_ ;
  assign \new_[10037]_  = \new_[13057]_  & \new_[20938]_ ;
  assign \new_[10038]_  = \new_[13152]_  & \new_[19547]_ ;
  assign \new_[10039]_  = ~\new_[17954]_  | ~\new_[12490]_ ;
  assign \new_[10040]_  = ~\new_[11113]_ ;
  assign \new_[10041]_  = ~\new_[14974]_  | ~\new_[19082]_ ;
  assign \new_[10042]_  = ~\new_[13693]_  | ~\new_[12783]_ ;
  assign \new_[10043]_  = \new_[13324]_  & \new_[21056]_ ;
  assign \new_[10044]_  = \new_[12734]_  | \new_[19553]_ ;
  assign \new_[10045]_  = ~\new_[13053]_  & ~\new_[16731]_ ;
  assign \new_[10046]_  = ~\new_[12932]_  & ~\new_[20233]_ ;
  assign \new_[10047]_  = ~\new_[13284]_  | ~\new_[19612]_ ;
  assign \new_[10048]_  = ~\new_[11122]_ ;
  assign \new_[10049]_  = ~\new_[12988]_  | ~\new_[16879]_ ;
  assign \new_[10050]_  = ~\new_[11124]_ ;
  assign \new_[10051]_  = ~\new_[12560]_  | ~\new_[14392]_ ;
  assign \new_[10052]_  = \new_[20921]_  | \new_[15004]_ ;
  assign \new_[10053]_  = ~\new_[11126]_ ;
  assign \new_[10054]_  = ~\new_[11129]_ ;
  assign \new_[10055]_  = ~\new_[13040]_  | ~\new_[19064]_ ;
  assign \new_[10056]_  = ~\new_[12885]_  | ~\new_[12810]_ ;
  assign \new_[10057]_  = ~\new_[19253]_  & ~\new_[12551]_ ;
  assign \new_[10058]_  = ~\new_[15401]_  | ~\new_[15298]_ ;
  assign \new_[10059]_  = ~\new_[12734]_  | ~\new_[12618]_ ;
  assign \new_[10060]_  = \new_[13951]_  & \new_[12816]_ ;
  assign \new_[10061]_  = ~\new_[12852]_  & ~\new_[12425]_ ;
  assign \new_[10062]_  = ~\new_[17390]_  & ~\new_[12723]_ ;
  assign \new_[10063]_  = ~\new_[14704]_  | ~\new_[13211]_ ;
  assign \new_[10064]_  = ~\new_[13291]_  | ~\new_[19567]_ ;
  assign \new_[10065]_  = ~\new_[12486]_  | (~\new_[17573]_  & ~\new_[18699]_ );
  assign \new_[10066]_  = ~\new_[18606]_  & (~\new_[16313]_  | ~\new_[14585]_ );
  assign \new_[10067]_  = ~\new_[16958]_  | ~\new_[12611]_ ;
  assign \new_[10068]_  = ~\new_[14022]_  | ~\new_[13294]_ ;
  assign \new_[10069]_  = ~\new_[16031]_  | ~\new_[13057]_ ;
  assign \new_[10070]_  = ~\new_[12513]_  | ~\new_[14883]_ ;
  assign \new_[10071]_  = ~\new_[12753]_  | ~\new_[19013]_ ;
  assign \new_[10072]_  = ~\new_[11146]_ ;
  assign \new_[10073]_  = ~\new_[11148]_ ;
  assign \new_[10074]_  = ~\new_[11149]_ ;
  assign \new_[10075]_  = ~\new_[15816]_  & ~\new_[13293]_ ;
  assign \new_[10076]_  = ~\new_[15326]_  | ~\new_[12800]_ ;
  assign \new_[10077]_  = ~\new_[12724]_  | ~\new_[16879]_ ;
  assign \new_[10078]_  = ~\new_[19937]_  | ~\new_[16231]_ ;
  assign \new_[10079]_  = ~\new_[13029]_  & ~\new_[12531]_ ;
  assign \new_[10080]_  = ~\new_[15058]_  | ~\new_[18832]_ ;
  assign \new_[10081]_  = ~\new_[13805]_  | ~\new_[12553]_ ;
  assign \new_[10082]_  = ~\new_[11153]_ ;
  assign \new_[10083]_  = \new_[12992]_  & \new_[19742]_ ;
  assign \new_[10084]_  = \new_[18873]_  & \new_[14932]_ ;
  assign \new_[10085]_  = ~\new_[12574]_  & ~\new_[15870]_ ;
  assign \new_[10086]_  = ~\new_[13547]_  | ~\new_[12975]_ ;
  assign \new_[10087]_  = ~\new_[12718]_  | ~\new_[13968]_ ;
  assign \new_[10088]_  = ~\new_[12564]_  | ~\new_[18166]_ ;
  assign \new_[10089]_  = \new_[15892]_  & \new_[13770]_ ;
  assign \new_[10090]_  = \new_[13004]_  & \new_[15119]_ ;
  assign \new_[10091]_  = ~\new_[13266]_  & ~\new_[15026]_ ;
  assign \new_[10092]_  = ~\new_[11155]_ ;
  assign \new_[10093]_  = \new_[12641]_  | \new_[18998]_ ;
  assign \new_[10094]_  = ~\new_[11158]_ ;
  assign \new_[10095]_  = ~\new_[11160]_ ;
  assign \new_[10096]_  = ~\new_[13952]_  & ~\new_[18373]_ ;
  assign \new_[10097]_  = ~\new_[12799]_  | ~\new_[16671]_ ;
  assign \new_[10098]_  = ~\new_[11163]_ ;
  assign \new_[10099]_  = \new_[12857]_  & \new_[19266]_ ;
  assign \new_[10100]_  = \new_[16631]_  | \new_[12165]_ ;
  assign \new_[10101]_  = ~\new_[12572]_  & ~\new_[19088]_ ;
  assign \new_[10102]_  = ~\new_[13071]_  | (~\new_[18192]_  & ~\new_[18390]_ );
  assign \new_[10103]_  = ~\new_[16569]_  & (~\new_[18807]_  | ~\new_[14602]_ );
  assign \new_[10104]_  = ~\new_[12898]_  | ~\new_[16326]_ ;
  assign \new_[10105]_  = \new_[16418]_  | \new_[21075]_ ;
  assign \new_[10106]_  = ~\new_[15081]_  | ~\new_[15278]_ ;
  assign \new_[10107]_  = ~\new_[12812]_  | ~\new_[17944]_ ;
  assign \new_[10108]_  = ~\new_[13064]_  & ~\new_[14160]_ ;
  assign \new_[10109]_  = ~\new_[14205]_  & ~\new_[12643]_ ;
  assign \new_[10110]_  = \new_[12669]_  | \new_[19239]_ ;
  assign \new_[10111]_  = ~\new_[12916]_  | ~\new_[15638]_ ;
  assign \new_[10112]_  = ~\new_[15008]_  | ~\new_[19697]_ ;
  assign \new_[10113]_  = \new_[17488]_  & \new_[12679]_ ;
  assign \new_[10114]_  = \new_[12520]_  | \new_[18443]_ ;
  assign \new_[10115]_  = ~\new_[16563]_  | ~\new_[19217]_ ;
  assign \new_[10116]_  = \new_[15555]_  & \new_[18187]_ ;
  assign \new_[10117]_  = ~\new_[12906]_  & ~\new_[15915]_ ;
  assign \new_[10118]_  = ~\new_[13162]_  & ~\new_[15956]_ ;
  assign \new_[10119]_  = ~\new_[11179]_ ;
  assign \new_[10120]_  = ~\new_[12629]_  | ~\new_[17181]_ ;
  assign \new_[10121]_  = ~\new_[14652]_  | ~\new_[13253]_ ;
  assign \new_[10122]_  = ~\new_[15215]_  | ~\new_[19050]_ ;
  assign \new_[10123]_  = ~\new_[12985]_  | ~\new_[18017]_ ;
  assign \new_[10124]_  = ~\new_[15041]_  | ~\new_[20927]_ ;
  assign \new_[10125]_  = ~\new_[11182]_ ;
  assign \new_[10126]_  = ~\new_[11097]_ ;
  assign \new_[10127]_  = ~\new_[16288]_  & ~\new_[12913]_ ;
  assign \new_[10128]_  = ~\new_[11185]_ ;
  assign \new_[10129]_  = ~\new_[12287]_ ;
  assign \new_[10130]_  = ~\new_[12777]_  | ~\new_[16259]_ ;
  assign \new_[10131]_  = ~\new_[15142]_  & ~\new_[17812]_ ;
  assign \new_[10132]_  = ~\new_[17845]_  | ~\new_[14874]_ ;
  assign \new_[10133]_  = ~\new_[12754]_  | ~\new_[16782]_ ;
  assign \new_[10134]_  = ~\new_[13099]_  & (~\new_[16351]_  | ~\new_[21394]_ );
  assign \new_[10135]_  = ~\new_[12871]_  & ~\new_[13427]_ ;
  assign \new_[10136]_  = \new_[12853]_  & \new_[18209]_ ;
  assign \new_[10137]_  = ~\new_[12816]_  | ~\new_[14078]_ ;
  assign \new_[10138]_  = ~\new_[14994]_  | ~\new_[19319]_ ;
  assign \new_[10139]_  = ~\new_[11192]_ ;
  assign \new_[10140]_  = ~\new_[12689]_  | ~\new_[19367]_ ;
  assign \new_[10141]_  = ~\new_[14928]_  & ~\new_[19366]_ ;
  assign \new_[10142]_  = ~\new_[17559]_  | ~\new_[14871]_ ;
  assign \new_[10143]_  = ~\new_[13727]_  | ~\new_[13057]_ ;
  assign \new_[10144]_  = ~\new_[19366]_  & (~\new_[13615]_  | ~\new_[13960]_ );
  assign \new_[10145]_  = ~\new_[11194]_ ;
  assign \new_[10146]_  = ~\new_[13464]_  & ~\new_[18833]_ ;
  assign \new_[10147]_  = ~\new_[15693]_  | ~\new_[15050]_ ;
  assign \new_[10148]_  = ~\new_[15161]_  | ~\new_[19711]_ ;
  assign \new_[10149]_  = ~\new_[11196]_ ;
  assign \new_[10150]_  = \new_[13019]_  | \new_[19021]_ ;
  assign \new_[10151]_  = ~\new_[12454]_  | ~\new_[14822]_ ;
  assign \new_[10152]_  = \new_[13133]_  & \new_[19239]_ ;
  assign \new_[10153]_  = ~\new_[13132]_  & ~\new_[13623]_ ;
  assign \new_[10154]_  = ~\new_[11202]_ ;
  assign \new_[10155]_  = ~\new_[11204]_ ;
  assign \new_[10156]_  = ~\new_[12843]_  & (~\new_[17060]_  | ~\new_[18794]_ );
  assign \new_[10157]_  = ~\new_[15336]_  | ~\new_[21328]_ ;
  assign \new_[10158]_  = ~\new_[15231]_  | ~\new_[15498]_ ;
  assign \new_[10159]_  = ~\new_[12984]_  | ~\new_[19578]_ ;
  assign \new_[10160]_  = \new_[15305]_  & \new_[16166]_ ;
  assign \new_[10161]_  = ~\new_[14935]_  | ~\new_[18111]_ ;
  assign \new_[10162]_  = ~\new_[12568]_  | ~\new_[14199]_ ;
  assign \new_[10163]_  = \new_[13211]_  & \new_[14381]_ ;
  assign \new_[10164]_  = ~\new_[12801]_  | ~\new_[19021]_ ;
  assign \new_[10165]_  = ~\new_[12596]_  & ~\new_[18537]_ ;
  assign \new_[10166]_  = ~\new_[12848]_  | ~\new_[15377]_ ;
  assign \new_[10167]_  = ~\new_[11210]_ ;
  assign \new_[10168]_  = ~\new_[12519]_  | ~\new_[18228]_ ;
  assign \new_[10169]_  = ~\new_[13152]_  & ~\new_[15088]_ ;
  assign \new_[10170]_  = \new_[15065]_  | \new_[18795]_ ;
  assign \new_[10171]_  = ~\new_[11941]_ ;
  assign \new_[10172]_  = ~\new_[12812]_  | ~\new_[19015]_ ;
  assign \new_[10173]_  = ~\new_[15039]_  | ~\new_[18981]_ ;
  assign \new_[10174]_  = ~\new_[12544]_  | ~\new_[13950]_ ;
  assign \new_[10175]_  = ~\new_[13122]_  | ~\new_[13831]_ ;
  assign \new_[10176]_  = ~\new_[12792]_  | ~\new_[13941]_ ;
  assign \new_[10177]_  = \new_[12629]_  & \new_[12158]_ ;
  assign \new_[10178]_  = ~\new_[17972]_  | ~\new_[14871]_ ;
  assign \new_[10179]_  = ~\new_[12650]_  | ~\new_[18998]_ ;
  assign \new_[10180]_  = \new_[16670]_  & \new_[15788]_ ;
  assign \new_[10181]_  = ~\new_[11220]_ ;
  assign \new_[10182]_  = ~\new_[11220]_ ;
  assign \new_[10183]_  = \new_[15496]_  & \new_[12818]_ ;
  assign \new_[10184]_  = ~\new_[11225]_ ;
  assign \new_[10185]_  = ~\new_[13427]_  | ~\new_[18083]_ ;
  assign \new_[10186]_  = ~\new_[12670]_  | ~\new_[20971]_ ;
  assign \new_[10187]_  = ~\new_[13420]_  | ~\new_[12918]_ ;
  assign \new_[10188]_  = ~\new_[12552]_  & ~\new_[21562]_ ;
  assign \new_[10189]_  = ~\new_[21674]_  | ~\new_[14083]_ ;
  assign \new_[10190]_  = ~\new_[19079]_  & (~\new_[15896]_  | ~\new_[14503]_ );
  assign \new_[10191]_  = ~\new_[12580]_  & ~\new_[12562]_ ;
  assign \new_[10192]_  = ~\new_[11228]_ ;
  assign \new_[10193]_  = ~\new_[15185]_  | ~\new_[13386]_ ;
  assign \new_[10194]_  = \new_[13323]_  & \new_[19247]_ ;
  assign \new_[10195]_  = ~\new_[12839]_  | ~\new_[13454]_ ;
  assign \new_[10196]_  = ~\new_[13977]_  | ~\new_[17343]_ ;
  assign \new_[10197]_  = ~\new_[15357]_  & ~\new_[13088]_ ;
  assign \new_[10198]_  = ~\new_[17325]_  | ~\new_[21094]_ ;
  assign \new_[10199]_  = ~\new_[11236]_ ;
  assign \new_[10200]_  = ~\new_[12362]_  | ~\new_[19024]_ ;
  assign \new_[10201]_  = ~\new_[11238]_ ;
  assign \new_[10202]_  = ~\new_[11239]_ ;
  assign \new_[10203]_  = ~\new_[17536]_  | ~\new_[12638]_ ;
  assign \new_[10204]_  = ~\new_[18909]_  | ~\new_[12521]_ ;
  assign \new_[10205]_  = ~\new_[12362]_  | ~\new_[17702]_ ;
  assign \new_[10206]_  = ~\new_[17486]_  | ~\new_[13399]_ ;
  assign \new_[10207]_  = ~\new_[11240]_ ;
  assign \new_[10208]_  = ~\new_[12158]_  | ~\new_[14015]_ ;
  assign \new_[10209]_  = ~\new_[13669]_  | ~\new_[13211]_ ;
  assign \new_[10210]_  = \new_[15108]_  | \new_[17979]_ ;
  assign \new_[10211]_  = \new_[12466]_  & \new_[20388]_ ;
  assign \new_[10212]_  = ~\new_[12611]_  | ~\new_[19021]_ ;
  assign \new_[10213]_  = ~\new_[12607]_  | ~\new_[21560]_ ;
  assign \new_[10214]_  = ~\new_[19462]_  & ~\new_[12771]_ ;
  assign \new_[10215]_  = ~\new_[12586]_  | ~\new_[21496]_ ;
  assign \new_[10216]_  = ~\new_[12686]_  & ~\new_[13844]_ ;
  assign \new_[10217]_  = \new_[12863]_  & \new_[15108]_ ;
  assign \new_[10218]_  = ~\new_[12646]_  | ~\new_[14183]_ ;
  assign \new_[10219]_  = ~\new_[11250]_ ;
  assign \new_[10220]_  = ~\new_[15069]_  | ~\new_[18678]_ ;
  assign \new_[10221]_  = ~\new_[12672]_  | ~\new_[19085]_ ;
  assign \new_[10222]_  = \new_[12882]_  | \new_[18070]_ ;
  assign \new_[10223]_  = ~\new_[15825]_  | ~\new_[19021]_ ;
  assign \new_[10224]_  = ~\new_[11253]_ ;
  assign \new_[10225]_  = ~\new_[12675]_  | ~\new_[18984]_ ;
  assign \new_[10226]_  = ~\new_[11254]_ ;
  assign \new_[10227]_  = ~\new_[11256]_ ;
  assign \new_[10228]_  = ~\new_[12613]_  & ~\new_[12795]_ ;
  assign \new_[10229]_  = \new_[15050]_  | \new_[21328]_ ;
  assign \new_[10230]_  = ~\new_[12651]_  & ~\new_[21638]_ ;
  assign \new_[10231]_  = ~\new_[12615]_  & ~\new_[15302]_ ;
  assign \new_[10232]_  = ~\new_[15862]_  | ~\new_[19050]_ ;
  assign \new_[10233]_  = ~\new_[17473]_  & ~\new_[13058]_ ;
  assign \new_[10234]_  = ~\new_[15797]_  | ~\new_[19275]_ ;
  assign \new_[10235]_  = ~\new_[11264]_ ;
  assign \new_[10236]_  = ~\new_[14931]_  | ~\new_[19214]_ ;
  assign \new_[10237]_  = ~\new_[11265]_ ;
  assign \new_[10238]_  = ~\new_[15511]_  | ~\new_[14013]_ ;
  assign \new_[10239]_  = ~\new_[15212]_  | ~\new_[12868]_ ;
  assign \new_[10240]_  = ~\new_[12538]_  & ~\new_[15903]_ ;
  assign \new_[10241]_  = \new_[12473]_  | \new_[12751]_ ;
  assign \new_[10242]_  = ~\new_[11267]_ ;
  assign \new_[10243]_  = ~\new_[11268]_ ;
  assign \new_[10244]_  = ~\new_[15074]_  | ~\new_[18325]_ ;
  assign \new_[10245]_  = ~\new_[15051]_  | ~\new_[12820]_ ;
  assign \new_[10246]_  = ~\new_[12161]_  | ~\new_[16277]_ ;
  assign \new_[10247]_  = ~\new_[15776]_  | ~\new_[12326]_ ;
  assign \new_[10248]_  = ~\new_[14741]_  | ~\new_[12818]_ ;
  assign \new_[10249]_  = ~\new_[12601]_  & ~\new_[17385]_ ;
  assign \new_[10250]_  = ~\new_[11277]_ ;
  assign \new_[10251]_  = \new_[12975]_  & \new_[14106]_ ;
  assign \new_[10252]_  = ~\new_[13365]_  | ~\new_[12468]_ ;
  assign \new_[10253]_  = ~\new_[14133]_  & ~\new_[13142]_ ;
  assign \new_[10254]_  = ~\new_[16342]_  & ~\new_[12671]_ ;
  assign \new_[10255]_  = ~\new_[17367]_  | ~\new_[12362]_ ;
  assign \new_[10256]_  = ~\new_[13167]_  | ~\new_[15201]_ ;
  assign \new_[10257]_  = ~\new_[21094]_  | ~\new_[18542]_ ;
  assign \new_[10258]_  = ~\new_[20907]_  | ~\new_[17086]_ ;
  assign \new_[10259]_  = \new_[17767]_  & \new_[14979]_ ;
  assign \new_[10260]_  = ~\new_[13292]_  | ~\new_[15263]_ ;
  assign \new_[10261]_  = \new_[12358]_  | \new_[19115]_ ;
  assign \new_[10262]_  = ~\new_[13154]_  | ~\new_[20341]_ ;
  assign \new_[10263]_  = ~\new_[18855]_  | ~\new_[12531]_ ;
  assign \new_[10264]_  = ~\new_[14843]_  & ~\new_[19145]_ ;
  assign \new_[10265]_  = \new_[12172]_  & \new_[17395]_ ;
  assign \new_[10266]_  = ~\new_[11288]_ ;
  assign \new_[10267]_  = ~\new_[18815]_  & ~\new_[13411]_ ;
  assign \new_[10268]_  = \new_[12552]_  & \new_[12929]_ ;
  assign \new_[10269]_  = ~\new_[12805]_  | ~\new_[18175]_ ;
  assign \new_[10270]_  = ~\new_[13020]_  | ~\new_[21507]_ ;
  assign \new_[10271]_  = ~\new_[12663]_  | ~\new_[19275]_ ;
  assign \new_[10272]_  = ~\new_[13138]_  & (~\new_[17195]_  | ~\new_[17572]_ );
  assign \new_[10273]_  = ~\new_[15172]_  & ~\new_[12874]_ ;
  assign \new_[10274]_  = ~\new_[11295]_ ;
  assign \new_[10275]_  = ~\new_[15213]_  & ~\new_[12731]_ ;
  assign \new_[10276]_  = ~\new_[16349]_  | ~\new_[15406]_  | ~\new_[14821]_ ;
  assign \new_[10277]_  = ~\new_[11297]_ ;
  assign \new_[10278]_  = ~\new_[12800]_  & ~\new_[21513]_ ;
  assign \new_[10279]_  = ~\new_[16078]_  & ~\new_[13085]_ ;
  assign \new_[10280]_  = ~\new_[15112]_  & ~\new_[19145]_ ;
  assign \new_[10281]_  = \new_[13817]_  & \new_[12540]_ ;
  assign \new_[10282]_  = ~\new_[11300]_ ;
  assign \new_[10283]_  = ~\new_[13179]_  & ~\new_[17139]_ ;
  assign \new_[10284]_  = \new_[16224]_  & \new_[13321]_ ;
  assign \new_[10285]_  = ~\new_[13102]_  | ~\new_[17667]_ ;
  assign \new_[10286]_  = ~\new_[13152]_  & ~\new_[16182]_ ;
  assign \new_[10287]_  = ~\new_[15805]_  | ~\new_[19085]_ ;
  assign \new_[10288]_  = ~\new_[12892]_  | ~\new_[18994]_ ;
  assign \new_[10289]_  = ~\new_[11306]_ ;
  assign \new_[10290]_  = ~\new_[18635]_  | ~\new_[14874]_ ;
  assign \new_[10291]_  = \new_[12608]_  & \new_[13590]_ ;
  assign \new_[10292]_  = ~\new_[16025]_  & ~\new_[19145]_  & ~\new_[20768]_ ;
  assign \new_[10293]_  = ~\new_[14742]_  | ~\new_[14385]_ ;
  assign \new_[10294]_  = ~\new_[13175]_  & (~\new_[17330]_  | ~\new_[20490]_ );
  assign \new_[10295]_  = ~\new_[16240]_  & ~\new_[12611]_ ;
  assign \new_[10296]_  = ~\new_[20971]_  | ~\new_[12494]_ ;
  assign \new_[10297]_  = ~\new_[12711]_  | ~\new_[21631]_ ;
  assign \new_[10298]_  = ~\new_[15195]_  | ~\new_[20971]_ ;
  assign \new_[10299]_  = ~\new_[13186]_  & ~\new_[21331]_ ;
  assign \new_[10300]_  = ~\new_[12418]_ ;
  assign \new_[10301]_  = \new_[12658]_  | \new_[17358]_ ;
  assign \new_[10302]_  = ~\new_[11315]_ ;
  assign \new_[10303]_  = ~\new_[11316]_ ;
  assign \new_[10304]_  = ~\new_[13207]_  | ~\new_[19202]_ ;
  assign \new_[10305]_  = ~\new_[18077]_  & (~\new_[16401]_  | ~\new_[14285]_ );
  assign \new_[10306]_  = ~\new_[12721]_  & ~\new_[13707]_ ;
  assign \new_[10307]_  = ~\new_[21132]_  | ~\new_[13321]_ ;
  assign \new_[10308]_  = ~\new_[21681]_  & ~\new_[21398]_ ;
  assign \new_[10309]_  = ~\new_[12651]_  & ~\new_[18012]_ ;
  assign \new_[10310]_  = ~\new_[12465]_  | ~\new_[12859]_ ;
  assign \new_[10311]_  = ~\new_[16128]_  | ~\new_[15220]_ ;
  assign \new_[10312]_  = ~\new_[12731]_  & ~\new_[12570]_ ;
  assign \new_[10313]_  = \new_[14829]_  | \new_[17598]_ ;
  assign \new_[10314]_  = ~\new_[12869]_  & ~\new_[13565]_ ;
  assign \new_[10315]_  = ~\new_[13035]_  | ~\new_[12515]_ ;
  assign \new_[10316]_  = \new_[13099]_  & \new_[21558]_ ;
  assign \new_[10317]_  = \new_[14829]_  & \new_[15556]_ ;
  assign \new_[10318]_  = ~\new_[17452]_  & ~\new_[15001]_ ;
  assign \new_[10319]_  = ~\new_[12805]_  | ~\new_[21562]_ ;
  assign \new_[10320]_  = ~\new_[12515]_  | ~\new_[12769]_ ;
  assign \new_[10321]_  = ~\new_[17098]_  | ~\new_[19208]_ ;
  assign \new_[10322]_  = ~\new_[11320]_ ;
  assign \new_[10323]_  = ~\new_[13175]_  | ~\new_[17689]_ ;
  assign \new_[10324]_  = \new_[12553]_  | \new_[19253]_ ;
  assign \new_[10325]_  = ~\new_[12196]_  & ~\new_[16247]_ ;
  assign \new_[10326]_  = ~\new_[12775]_  | ~\new_[13494]_ ;
  assign \new_[10327]_  = ~\new_[14275]_  | ~\new_[15581]_ ;
  assign \new_[10328]_  = ~\new_[13124]_  | ~\new_[17797]_ ;
  assign \new_[10329]_  = \new_[15018]_  & \new_[19727]_ ;
  assign \new_[10330]_  = ~\new_[11330]_ ;
  assign \new_[10331]_  = ~\new_[12947]_  | ~\new_[15637]_ ;
  assign \new_[10332]_  = \new_[15260]_  & \new_[18833]_ ;
  assign \new_[10333]_  = ~\new_[13146]_  | ~\new_[15263]_ ;
  assign \new_[10334]_  = ~\new_[11984]_ ;
  assign \new_[10335]_  = ~\new_[13004]_  | ~\new_[13400]_ ;
  assign \new_[10336]_  = ~\new_[12858]_  | ~\new_[17218]_ ;
  assign \new_[10337]_  = ~\new_[12696]_  | ~\new_[14165]_ ;
  assign \new_[10338]_  = ~\new_[13343]_  | ~\new_[18984]_ ;
  assign \new_[10339]_  = ~\new_[13792]_  & ~\new_[12150]_ ;
  assign \new_[10340]_  = ~\new_[11339]_ ;
  assign \new_[10341]_  = ~\new_[21094]_  | ~\new_[18597]_ ;
  assign \new_[10342]_  = ~\new_[14687]_  | ~\new_[14869]_ ;
  assign \new_[10343]_  = ~\new_[12704]_  & ~\new_[12506]_ ;
  assign \new_[10344]_  = ~\new_[15093]_  | ~\new_[13225]_ ;
  assign \new_[10345]_  = ~\new_[11917]_ ;
  assign \new_[10346]_  = ~\new_[13094]_  | ~\new_[12696]_ ;
  assign \new_[10347]_  = ~\new_[13391]_  | ~\new_[19102]_ ;
  assign \new_[10348]_  = ~\new_[12737]_  | ~\new_[13831]_ ;
  assign \new_[10349]_  = ~\new_[14247]_  | ~\new_[12539]_ ;
  assign \new_[10350]_  = ~\new_[13038]_  & ~\new_[14448]_ ;
  assign \new_[10351]_  = ~\new_[15310]_  & ~\new_[21693]_ ;
  assign \new_[10352]_  = ~\new_[15310]_  | ~\new_[15526]_ ;
  assign \new_[10353]_  = ~\new_[13870]_  | ~\new_[13019]_ ;
  assign \new_[10354]_  = ~\new_[15274]_  | ~\new_[21675]_ ;
  assign \new_[10355]_  = ~\new_[17775]_  | ~\new_[13203]_ ;
  assign \new_[10356]_  = \new_[13684]_  & \new_[12977]_ ;
  assign \new_[10357]_  = ~\new_[13589]_  & (~\new_[14438]_  | ~\new_[18652]_ );
  assign \new_[10358]_  = ~\new_[13220]_  | ~\new_[19145]_ ;
  assign \new_[10359]_  = ~\new_[21251]_ ;
  assign \new_[10360]_  = ~\new_[18062]_  & ~\new_[12455]_ ;
  assign \new_[10361]_  = ~\new_[19260]_  | ~\new_[14935]_ ;
  assign \new_[10362]_  = ~\new_[12539]_  | ~\new_[14074]_ ;
  assign \new_[10363]_  = ~\new_[17983]_  | ~\new_[12587]_ ;
  assign \new_[10364]_  = ~\new_[11351]_ ;
  assign \new_[10365]_  = ~\new_[18180]_  & ~\new_[13222]_ ;
  assign \new_[10366]_  = ~\new_[12752]_  & ~\new_[12577]_ ;
  assign \new_[10367]_  = ~\new_[12543]_  & ~\new_[19215]_ ;
  assign \new_[10368]_  = ~\new_[14803]_  | ~\new_[19008]_ ;
  assign \new_[10369]_  = ~\new_[13068]_  | ~\new_[13395]_ ;
  assign \new_[10370]_  = ~\new_[11353]_ ;
  assign \new_[10371]_  = \new_[16141]_  & \new_[12641]_ ;
  assign \new_[10372]_  = ~\new_[12976]_  & ~\new_[19547]_ ;
  assign \new_[10373]_  = ~\new_[13170]_  | ~\new_[16745]_ ;
  assign \new_[10374]_  = \new_[14961]_  & \new_[12669]_ ;
  assign \new_[10375]_  = ~\new_[12429]_  | ~\new_[18322]_ ;
  assign \new_[10376]_  = ~\new_[21164]_  | ~\new_[15800]_ ;
  assign \new_[10377]_  = ~\new_[11359]_ ;
  assign \new_[10378]_  = ~\new_[12843]_  | ~\new_[18863]_ ;
  assign \new_[10379]_  = ~\new_[12810]_  | ~\new_[14009]_ ;
  assign \new_[10380]_  = ~\new_[12732]_  | ~\new_[13293]_ ;
  assign \new_[10381]_  = ~\new_[11364]_ ;
  assign \new_[10382]_  = ~\new_[12504]_  | ~\new_[13454]_ ;
  assign \new_[10383]_  = ~\new_[15290]_  | ~\new_[13306]_ ;
  assign \new_[10384]_  = ~\new_[12657]_  | ~\new_[13782]_ ;
  assign \new_[10385]_  = ~\new_[21662]_  & ~\new_[13987]_ ;
  assign \new_[10386]_  = ~\new_[11369]_ ;
  assign \new_[10387]_  = ~\new_[12659]_  & ~\new_[19072]_ ;
  assign \new_[10388]_  = ~\new_[16607]_  | ~\new_[14754]_  | ~\new_[16409]_  | ~\new_[16314]_ ;
  assign \new_[10389]_  = ~\new_[14283]_  | ~\new_[12966]_ ;
  assign \new_[10390]_  = ~\new_[12894]_  | ~\new_[19532]_ ;
  assign \new_[10391]_  = ~\new_[12783]_  | ~\new_[14113]_ ;
  assign \new_[10392]_  = ~\new_[11378]_ ;
  assign \new_[10393]_  = ~\new_[12312]_  | ~\new_[19015]_ ;
  assign \new_[10394]_  = \new_[14978]_  | \new_[17457]_ ;
  assign \new_[10395]_  = ~\new_[11381]_ ;
  assign \new_[10396]_  = ~\new_[13181]_  | ~\new_[19327]_ ;
  assign \new_[10397]_  = ~\new_[14193]_  & ~\new_[13462]_ ;
  assign \new_[10398]_  = ~\new_[15173]_  | ~\new_[13282]_ ;
  assign \new_[10399]_  = ~\new_[18037]_  | ~\new_[15761]_ ;
  assign \new_[10400]_  = ~\new_[11384]_ ;
  assign \new_[10401]_  = ~\new_[12725]_  & ~\new_[16470]_ ;
  assign \new_[10402]_  = ~\new_[11387]_ ;
  assign \new_[10403]_  = ~\new_[17043]_  | ~\new_[12729]_ ;
  assign \new_[10404]_  = ~\new_[12518]_  | ~\new_[18157]_ ;
  assign \new_[10405]_  = ~\new_[11388]_ ;
  assign \new_[10406]_  = ~\new_[14502]_  | ~\new_[15852]_  | ~\new_[15200]_ ;
  assign \new_[10407]_  = ~\new_[13210]_  | ~\new_[17106]_ ;
  assign \new_[10408]_  = ~\new_[15633]_  | ~\new_[20969]_ ;
  assign \new_[10409]_  = ~\new_[14828]_  & (~\new_[14482]_  | ~\new_[19249]_ );
  assign \new_[10410]_  = ~\new_[15144]_  & ~\new_[21601]_ ;
  assign \new_[10411]_  = ~\new_[12903]_  | ~\new_[15268]_ ;
  assign \new_[10412]_  = \new_[13360]_  & \new_[12900]_ ;
  assign \new_[10413]_  = ~\new_[14988]_  & ~\new_[14260]_ ;
  assign \new_[10414]_  = ~\new_[11400]_ ;
  assign \new_[10415]_  = ~\new_[12886]_  | ~\new_[17252]_ ;
  assign \new_[10416]_  = ~\new_[17027]_  | ~\new_[12528]_ ;
  assign \new_[10417]_  = ~\new_[15148]_  & (~\new_[16619]_  | ~\new_[21542]_ );
  assign \new_[10418]_  = ~\new_[12169]_  & ~\new_[12714]_ ;
  assign \new_[10419]_  = ~\new_[12514]_  & ~\new_[15208]_ ;
  assign \new_[10420]_  = ~\new_[11405]_ ;
  assign \new_[10421]_  = ~\new_[14089]_  | ~\new_[13233]_ ;
  assign \new_[10422]_  = ~\new_[13040]_  & (~\new_[17147]_  | ~\new_[21541]_ );
  assign \new_[10423]_  = ~\new_[11409]_ ;
  assign \new_[10424]_  = ~\new_[14265]_  & ~\new_[12600]_ ;
  assign \new_[10425]_  = ~\new_[15320]_  | ~\new_[20899]_ ;
  assign \new_[10426]_  = ~\new_[13384]_  | ~\new_[12550]_ ;
  assign \new_[10427]_  = ~\new_[19145]_  & (~\new_[16295]_  | ~\new_[16025]_ );
  assign \new_[10428]_  = ~\new_[13090]_  | ~\new_[17585]_ ;
  assign \new_[10429]_  = \new_[21138]_  | \new_[16569]_ ;
  assign \new_[10430]_  = ~\new_[14419]_  | (~\new_[14509]_  & ~\new_[19266]_ );
  assign \new_[10431]_  = ~\new_[13107]_  | ~\new_[17323]_ ;
  assign \new_[10432]_  = ~\new_[12713]_  | ~\new_[13361]_ ;
  assign \new_[10433]_  = ~\new_[15314]_  & (~\new_[17948]_  | ~\new_[18045]_ );
  assign \new_[10434]_  = ~\new_[12579]_  & (~\new_[16140]_  | ~\new_[18228]_ );
  assign \new_[10435]_  = ~\new_[14309]_  & ~\new_[12621]_ ;
  assign \new_[10436]_  = \new_[13405]_  & \new_[14210]_ ;
  assign \new_[10437]_  = ~\new_[11418]_ ;
  assign \new_[10438]_  = ~\new_[11419]_ ;
  assign \new_[10439]_  = ~\new_[11420]_ ;
  assign \new_[10440]_  = ~\new_[15691]_  | ~\new_[12807]_ ;
  assign \new_[10441]_  = ~\new_[12979]_  | ~\new_[13468]_ ;
  assign \new_[10442]_  = ~\new_[13312]_  | ~\new_[16886]_ ;
  assign \new_[10443]_  = ~\new_[13098]_  | ~\new_[15258]_ ;
  assign \new_[10444]_  = ~\new_[15460]_  | ~\new_[12726]_ ;
  assign \new_[10445]_  = ~\new_[12668]_  & (~\new_[16365]_  | ~\new_[17730]_ );
  assign \new_[10446]_  = ~\new_[13304]_  | ~\new_[12234]_ ;
  assign \new_[10447]_  = ~\new_[12525]_  & ~\new_[12454]_ ;
  assign \new_[10448]_  = ~\new_[16996]_  | ~\new_[12811]_ ;
  assign \new_[10449]_  = ~\new_[13136]_  & (~\new_[16408]_  | ~\new_[21693]_ );
  assign \new_[10450]_  = ~\new_[12548]_  | ~\new_[12885]_ ;
  assign \new_[10451]_  = ~\new_[12557]_  | ~\new_[14901]_ ;
  assign \new_[10452]_  = ~\new_[13467]_  & (~\new_[16035]_  | ~\new_[18166]_ );
  assign \new_[10453]_  = ~\new_[13730]_  & (~\new_[14501]_  | ~\new_[19156]_ );
  assign \new_[10454]_  = ~\new_[12510]_  & (~\new_[14676]_  | ~\new_[21697]_ );
  assign \new_[10455]_  = ~\new_[12703]_  | ~\new_[14035]_ ;
  assign \new_[10456]_  = ~\new_[12808]_  | ~\new_[15231]_ ;
  assign \new_[10457]_  = ~\new_[12653]_  | ~\new_[15212]_ ;
  assign \new_[10458]_  = ~\new_[13491]_  | ~\new_[13018]_ ;
  assign \new_[10459]_  = ~\new_[15121]_  & (~\new_[14592]_  | ~\new_[19290]_ );
  assign \new_[10460]_  = ~\new_[12634]_  | ~\new_[13012]_ ;
  assign \new_[10461]_  = ~\new_[12599]_  | ~\new_[15274]_ ;
  assign \new_[10462]_  = ~\new_[15373]_  & (~\new_[14519]_  | ~\new_[19589]_ );
  assign \new_[10463]_  = ~\new_[12545]_  & (~\new_[17042]_  | ~\new_[18427]_ );
  assign \new_[10464]_  = ~\new_[12695]_  | ~\new_[14347]_ ;
  assign \new_[10465]_  = ~\new_[12708]_  & ~\new_[12706]_ ;
  assign \new_[10466]_  = ~\new_[13738]_  & (~\new_[13485]_  | ~\new_[18652]_ );
  assign \new_[10467]_  = ~\new_[12535]_  | ~\new_[15277]_ ;
  assign \new_[10468]_  = ~\new_[13937]_  | ~\new_[15108]_ ;
  assign \new_[10469]_  = ~\new_[14034]_  & (~\new_[14484]_  | ~\new_[18832]_ );
  assign \new_[10470]_  = ~\new_[13867]_  & ~\new_[12637]_ ;
  assign \new_[10471]_  = ~\new_[13948]_  & ~\new_[12605]_ ;
  assign \new_[10472]_  = ~\new_[17696]_  & (~\new_[16012]_  | ~\new_[15545]_ );
  assign \new_[10473]_  = ~\new_[14897]_  | (~\new_[17615]_  & ~\new_[17592]_ );
  assign \new_[10474]_  = ~\new_[13121]_  & (~\new_[17325]_  | ~\new_[17709]_ );
  assign \new_[10475]_  = ~\new_[13444]_  | ~\new_[15325]_ ;
  assign \new_[10476]_  = \new_[13383]_  | \new_[14668]_ ;
  assign \new_[10477]_  = \new_[12972]_  & \new_[17640]_ ;
  assign \new_[10478]_  = ~\new_[12828]_  & (~\new_[17357]_  | ~\new_[17614]_ );
  assign \new_[10479]_  = ~\new_[17626]_  | (~\new_[17793]_  & ~\new_[14393]_ );
  assign \new_[10480]_  = ~\new_[13070]_  | ~\new_[18276]_ ;
  assign \new_[10481]_  = ~\new_[13338]_  | ~\new_[13719]_ ;
  assign \new_[10482]_  = ~\new_[18001]_  & (~\new_[21609]_  | ~\new_[14500]_ );
  assign \new_[10483]_  = ~\new_[16549]_  | ~\new_[12553]_ ;
  assign \new_[10484]_  = ~\new_[18564]_  & (~\new_[14663]_  | ~\new_[16515]_ );
  assign \new_[10485]_  = ~\new_[16998]_  | (~\new_[17368]_  & ~\new_[14393]_ );
  assign \new_[10486]_  = ~\new_[13234]_  | ~\new_[18370]_ ;
  assign \new_[10487]_  = \new_[13026]_  | \new_[14160]_ ;
  assign \new_[10488]_  = ~\new_[12995]_  | ~\new_[13015]_ ;
  assign \new_[10489]_  = ~\new_[13056]_  | ~\new_[14130]_ ;
  assign \new_[10490]_  = ~\new_[12940]_  & (~\new_[18849]_  | ~\new_[16414]_ );
  assign \new_[10491]_  = ~\new_[13612]_  | ~\new_[13164]_ ;
  assign \new_[10492]_  = \new_[14368]_  | \new_[12874]_ ;
  assign \new_[10493]_  = \new_[13227]_  | \new_[14133]_ ;
  assign \new_[10494]_  = ~\new_[18250]_  | (~\new_[15926]_  & ~\new_[16794]_ );
  assign \new_[10495]_  = ~\new_[13396]_  | ~\new_[14134]_ ;
  assign \new_[10496]_  = ~\new_[18319]_  | (~\new_[14501]_  & ~\new_[16871]_ );
  assign \new_[10497]_  = ~\new_[18323]_  | (~\new_[14592]_  & ~\new_[17296]_ );
  assign \new_[10498]_  = \new_[16378]_  & \new_[12960]_ ;
  assign \new_[10499]_  = \new_[16518]_  & \new_[13235]_ ;
  assign \new_[10500]_  = \new_[15623]_  & \new_[13156]_ ;
  assign \new_[10501]_  = \new_[18922]_  ^ \new_[13542]_ ;
  assign \new_[10502]_  = \new_[18892]_  ^ \new_[14653]_ ;
  assign \new_[10503]_  = \new_[18879]_  ^ \new_[14650]_ ;
  assign \new_[10504]_  = \new_[18828]_  ^ \new_[14649]_ ;
  assign \new_[10505]_  = ~\new_[11574]_ ;
  assign \new_[10506]_  = ~\new_[12121]_ ;
  assign \new_[10507]_  = ~\new_[12202]_  | ~\new_[21168]_ ;
  assign \new_[10508]_  = ~\new_[13349]_  | ~\new_[18285]_ ;
  assign \new_[10509]_  = ~\new_[11502]_ ;
  assign \new_[10510]_  = ~\new_[13429]_  | ~\new_[18166]_ ;
  assign \new_[10511]_  = ~\new_[11503]_ ;
  assign \new_[10512]_  = ~\new_[21409]_ ;
  assign \new_[10513]_  = ~\new_[11506]_ ;
  assign \new_[10514]_  = ~\new_[11507]_ ;
  assign \new_[10515]_  = ~\new_[12101]_ ;
  assign \new_[10516]_  = \new_[21631]_  | \new_[15849]_ ;
  assign \new_[10517]_  = ~\new_[13415]_  | ~\new_[18166]_ ;
  assign \new_[10518]_  = ~\new_[11510]_ ;
  assign \new_[10519]_  = ~\new_[11511]_ ;
  assign \new_[10520]_  = ~\new_[12094]_ ;
  assign \new_[10521]_  = ~\new_[12538]_ ;
  assign \new_[10522]_  = ~\new_[11514]_ ;
  assign \new_[10523]_  = \new_[13400]_  | \new_[18166]_ ;
  assign \new_[10524]_  = ~\new_[11517]_ ;
  assign \new_[10525]_  = ~\new_[12562]_ ;
  assign \new_[10526]_  = ~\new_[11524]_ ;
  assign \new_[10527]_  = ~\new_[11525]_ ;
  assign \new_[10528]_  = ~\new_[13775]_ ;
  assign \new_[10529]_  = ~\new_[11533]_ ;
  assign \new_[10530]_  = ~\new_[11540]_ ;
  assign \new_[10531]_  = ~\new_[13176]_  | ~\new_[18443]_ ;
  assign \new_[10532]_  = ~\new_[13374]_  | ~\new_[19217]_ ;
  assign \new_[10533]_  = ~\new_[11554]_ ;
  assign \new_[10534]_  = \new_[13334]_  & \new_[18270]_ ;
  assign \new_[10535]_  = ~\new_[13442]_  | ~\new_[18974]_ ;
  assign \new_[10536]_  = ~\new_[13394]_  | ~\new_[18973]_ ;
  assign \new_[10537]_  = ~\new_[12350]_  | ~\new_[19625]_ ;
  assign \new_[10538]_  = ~\new_[11567]_ ;
  assign \new_[10539]_  = ~\new_[13380]_  | ~\new_[18427]_ ;
  assign \new_[10540]_  = ~\new_[11578]_ ;
  assign \new_[10541]_  = ~\new_[11585]_ ;
  assign \new_[10542]_  = ~\new_[11595]_ ;
  assign \new_[10543]_  = ~\new_[11596]_ ;
  assign \new_[10544]_  = ~\new_[19942]_ ;
  assign \new_[10545]_  = ~\new_[10903]_ ;
  assign \new_[10546]_  = ~\new_[11600]_ ;
  assign \new_[10547]_  = ~\new_[11602]_ ;
  assign \new_[10548]_  = ~\new_[11604]_ ;
  assign \new_[10549]_  = ~\new_[15019]_  | ~\new_[19008]_ ;
  assign \new_[10550]_  = ~\new_[11610]_ ;
  assign \new_[10551]_  = ~\new_[11161]_ ;
  assign \new_[10552]_  = ~\new_[11615]_ ;
  assign \new_[10553]_  = ~\new_[13479]_  | ~\new_[19275]_ ;
  assign \new_[10554]_  = ~\new_[13424]_  | ~\new_[19085]_ ;
  assign \new_[10555]_  = ~\new_[11626]_ ;
  assign \new_[10556]_  = ~\new_[11046]_ ;
  assign \new_[10557]_  = ~\new_[11004]_ ;
  assign \new_[10558]_  = ~\new_[13426]_  | ~\new_[21499]_ ;
  assign \new_[10559]_  = ~\new_[11641]_ ;
  assign \new_[10560]_  = ~\new_[13418]_  | ~\new_[15767]_ ;
  assign \new_[10561]_  = ~\new_[13539]_ ;
  assign \new_[10562]_  = ~\new_[20522]_ ;
  assign \new_[10563]_  = ~\new_[19088]_  & (~\new_[16171]_  | ~\new_[14329]_ );
  assign \new_[10564]_  = ~\new_[10861]_ ;
  assign \new_[10565]_  = ~\new_[20705]_ ;
  assign \new_[10566]_  = ~\new_[11674]_ ;
  assign \new_[10567]_  = \new_[13358]_  | \new_[19102]_ ;
  assign \new_[10568]_  = ~\new_[11679]_ ;
  assign \new_[10569]_  = ~\new_[13416]_  | ~\new_[21697]_ ;
  assign \new_[10570]_  = \new_[17262]_  | \new_[13393]_ ;
  assign \new_[10571]_  = ~\new_[13393]_  | ~\new_[18427]_ ;
  assign \new_[10572]_  = ~\new_[11689]_ ;
  assign \new_[10573]_  = ~\new_[11694]_ ;
  assign \new_[10574]_  = ~\new_[14891]_  | ~\new_[18083]_ ;
  assign \new_[10575]_  = ~\new_[13437]_  | ~\new_[18569]_ ;
  assign \new_[10576]_  = ~\new_[11705]_ ;
  assign \new_[10577]_  = ~\new_[13390]_  | ~\new_[17469]_ ;
  assign \new_[10578]_  = ~\new_[11711]_ ;
  assign \new_[10579]_  = ~\new_[12795]_ ;
  assign \new_[10580]_  = ~\new_[11715]_ ;
  assign \new_[10581]_  = ~\new_[11716]_ ;
  assign \new_[10582]_  = ~\new_[11721]_ ;
  assign \new_[10583]_  = ~\new_[17147]_  | ~\new_[13176]_ ;
  assign \new_[10584]_  = ~\new_[20232]_ ;
  assign \new_[10585]_  = ~\new_[11733]_ ;
  assign \new_[10586]_  = ~\new_[15706]_  | ~\new_[19208]_ ;
  assign \new_[10587]_  = \new_[17583]_  | \new_[21651]_ ;
  assign \new_[10588]_  = ~\new_[11738]_ ;
  assign \new_[10589]_  = ~\new_[11742]_ ;
  assign \new_[10590]_  = ~\new_[11745]_ ;
  assign \new_[10591]_  = ~\new_[17359]_  | ~\new_[12342]_ ;
  assign \new_[10592]_  = \new_[18308]_  | \new_[15427]_ ;
  assign \new_[10593]_  = ~\new_[11750]_ ;
  assign \new_[10594]_  = ~\new_[11755]_ ;
  assign \new_[10595]_  = ~\new_[13375]_  | ~\new_[18023]_ ;
  assign \new_[10596]_  = ~\new_[12862]_ ;
  assign \new_[10597]_  = ~\new_[14304]_ ;
  assign \new_[10598]_  = ~\new_[17159]_  & ~\new_[15619]_ ;
  assign \new_[10599]_  = ~\new_[11762]_ ;
  assign \new_[10600]_  = \new_[13443]_  | \new_[18840]_ ;
  assign \new_[10601]_  = ~\new_[11771]_ ;
  assign \new_[10602]_  = ~\new_[11832]_ ;
  assign \new_[10603]_  = ~\new_[11775]_ ;
  assign \new_[10604]_  = ~\new_[11776]_ ;
  assign \new_[10605]_  = ~\new_[13176]_  | ~\new_[16797]_ ;
  assign \new_[10606]_  = ~\new_[13407]_  & ~\new_[18077]_ ;
  assign \new_[10607]_  = ~\new_[11780]_ ;
  assign \new_[10608]_  = ~\new_[11785]_ ;
  assign \new_[10609]_  = ~\new_[11789]_ ;
  assign \new_[10610]_  = ~\new_[18558]_  | ~\new_[21551]_ ;
  assign \new_[10611]_  = \new_[18930]_  | \new_[15123]_ ;
  assign \new_[10612]_  = \new_[17618]_  | \new_[14825]_ ;
  assign \new_[10613]_  = \new_[17628]_  | \new_[15568]_ ;
  assign \new_[10614]_  = ~\new_[18605]_  & ~\new_[13347]_ ;
  assign \new_[10615]_  = \new_[13400]_  & \new_[15020]_ ;
  assign \new_[10616]_  = ~\new_[13259]_  | ~\new_[20747]_ ;
  assign \new_[10617]_  = ~\new_[13668]_ ;
  assign \new_[10618]_  = \new_[18731]_  | \new_[13358]_ ;
  assign \new_[10619]_  = ~\new_[11813]_ ;
  assign \new_[10620]_  = ~\new_[15616]_  | ~\new_[17979]_ ;
  assign \new_[10621]_  = ~\new_[13363]_  | ~\new_[18818]_ ;
  assign \new_[10622]_  = ~\new_[15463]_  | ~\new_[19241]_ ;
  assign \new_[10623]_  = ~\new_[11818]_ ;
  assign \new_[10624]_  = ~\new_[17991]_  | ~\new_[13393]_ ;
  assign \new_[10625]_  = ~\new_[15616]_  | ~\new_[18167]_ ;
  assign \new_[10626]_  = ~\new_[10876]_ ;
  assign \new_[10627]_  = \new_[14742]_  | \new_[18637]_ ;
  assign \new_[10628]_  = ~\new_[11843]_ ;
  assign \new_[10629]_  = ~\new_[14734]_  | ~\new_[18825]_ ;
  assign \new_[10630]_  = \new_[12645]_  | \new_[15530]_ ;
  assign \new_[10631]_  = \new_[13377]_  | \new_[18111]_ ;
  assign \new_[10632]_  = ~\new_[15811]_  | ~\new_[14567]_ ;
  assign \new_[10633]_  = ~\new_[11850]_ ;
  assign \new_[10634]_  = ~\new_[18120]_  | ~\new_[12729]_ ;
  assign \new_[10635]_  = ~\new_[17993]_  & ~\new_[21701]_ ;
  assign \new_[10636]_  = ~\new_[13450]_  | ~\new_[15523]_ ;
  assign \new_[10637]_  = ~\new_[10850]_ ;
  assign \new_[10638]_  = ~\new_[18558]_  | ~\new_[15461]_ ;
  assign \new_[10639]_  = ~\new_[19098]_  | ~\new_[18981]_  | ~\new_[18310]_ ;
  assign \new_[10640]_  = ~\new_[15639]_  | ~\new_[19214]_ ;
  assign \new_[10641]_  = ~\new_[14221]_  | ~\new_[13222]_ ;
  assign \new_[10642]_  = ~\new_[11863]_ ;
  assign \new_[10643]_  = ~\new_[11865]_ ;
  assign \new_[10644]_  = ~\new_[12089]_ ;
  assign \new_[10645]_  = ~\new_[12250]_  & ~\new_[18709]_ ;
  assign \new_[10646]_  = ~\new_[13479]_  | ~\new_[18818]_ ;
  assign \new_[10647]_  = ~\new_[11869]_ ;
  assign \new_[10648]_  = ~\new_[17840]_  | ~\new_[12342]_ ;
  assign \new_[10649]_  = ~\new_[14751]_  | ~\new_[18873]_ ;
  assign \new_[10650]_  = ~\new_[11875]_ ;
  assign \new_[10651]_  = ~\new_[15711]_  | ~\new_[14607]_ ;
  assign \new_[10652]_  = ~\new_[11983]_ ;
  assign \new_[10653]_  = ~\new_[13432]_  | ~\new_[15594]_ ;
  assign \new_[10654]_  = ~\new_[21550]_  | ~\new_[18941]_ ;
  assign \new_[10655]_  = ~\new_[11888]_ ;
  assign \new_[10656]_  = ~\new_[18543]_  | ~\new_[13374]_ ;
  assign \new_[10657]_  = ~\new_[11889]_ ;
  assign \new_[10658]_  = ~\new_[11890]_ ;
  assign \new_[10659]_  = ~\new_[13062]_ ;
  assign \new_[10660]_  = ~\new_[11897]_ ;
  assign \new_[10661]_  = \new_[13347]_  | \new_[21115]_ ;
  assign \new_[10662]_  = ~\new_[11903]_ ;
  assign \new_[10663]_  = ~\new_[11905]_ ;
  assign \new_[10664]_  = ~\new_[11784]_ ;
  assign \new_[10665]_  = ~\new_[13461]_  & ~\new_[21686]_ ;
  assign \new_[10666]_  = \new_[18006]_  | \new_[15694]_ ;
  assign \new_[10667]_  = \new_[13376]_  | \new_[18766]_ ;
  assign \new_[10668]_  = ~\new_[13404]_  | ~\new_[18325]_ ;
  assign \new_[10669]_  = ~\new_[11915]_ ;
  assign \new_[10670]_  = ~\new_[17980]_  & ~\new_[13356]_ ;
  assign \new_[10671]_  = ~\new_[11920]_ ;
  assign \new_[10672]_  = ~\new_[11921]_ ;
  assign \new_[10673]_  = \new_[15820]_  | \new_[18930]_ ;
  assign \new_[10674]_  = ~\new_[18898]_  | ~\new_[13429]_ ;
  assign \new_[10675]_  = ~\new_[11932]_ ;
  assign \new_[10676]_  = ~\new_[13447]_  | ~\new_[15582]_ ;
  assign \new_[10677]_  = ~\new_[11383]_ ;
  assign \new_[10678]_  = ~\new_[13379]_  | ~\new_[16482]_ ;
  assign \new_[10679]_  = ~\new_[13349]_  | ~\new_[18086]_ ;
  assign \new_[10680]_  = ~\new_[17626]_  | ~\new_[21551]_ ;
  assign \new_[10681]_  = ~\new_[13404]_  & ~\new_[16202]_ ;
  assign \new_[10682]_  = ~\new_[13425]_  | ~\new_[19044]_ ;
  assign \new_[10683]_  = ~\new_[13348]_  | ~\new_[18557]_ ;
  assign \new_[10684]_  = \new_[14703]_  & \new_[15455]_ ;
  assign \new_[10685]_  = \new_[13347]_  & \new_[13366]_ ;
  assign \new_[10686]_  = ~\new_[11974]_ ;
  assign \new_[10687]_  = \new_[13453]_  | \new_[15530]_ ;
  assign \new_[10688]_  = ~\new_[14728]_  | ~\new_[18278]_ ;
  assign \new_[10689]_  = ~\new_[13428]_  | ~\new_[19088]_ ;
  assign \new_[10690]_  = ~\new_[19050]_  & ~\new_[15758]_ ;
  assign \new_[10691]_  = ~\new_[17338]_  | ~\new_[13411]_ ;
  assign \new_[10692]_  = ~\new_[11985]_ ;
  assign \new_[10693]_  = ~\new_[12177]_  & ~\new_[19269]_ ;
  assign \new_[10694]_  = ~\new_[11851]_ ;
  assign \new_[10695]_  = ~\new_[17807]_  | ~\new_[13483]_ ;
  assign \new_[10696]_  = \new_[13350]_  | \new_[17812]_ ;
  assign \new_[10697]_  = ~\new_[18275]_  | ~\new_[14718]_ ;
  assign \new_[10698]_  = ~\new_[11996]_ ;
  assign \new_[10699]_  = \new_[18233]_  | \new_[13457]_ ;
  assign \new_[10700]_  = ~\new_[11656]_ ;
  assign \new_[10701]_  = ~\new_[13458]_  | ~\new_[15777]_ ;
  assign \new_[10702]_  = ~\new_[12006]_ ;
  assign \new_[10703]_  = ~\new_[12009]_ ;
  assign \new_[10704]_  = ~\new_[13536]_  | ~\new_[12231]_ ;
  assign \new_[10705]_  = ~\new_[11266]_ ;
  assign \new_[10706]_  = ~\new_[12019]_ ;
  assign \new_[10707]_  = ~\new_[13419]_  | ~\new_[16807]_ ;
  assign \new_[10708]_  = ~\new_[18184]_  | ~\new_[13344]_ ;
  assign \new_[10709]_  = ~\new_[11229]_ ;
  assign \new_[10710]_  = ~\new_[18790]_  & ~\new_[13385]_ ;
  assign \new_[10711]_  = ~\new_[15182]_  & (~\new_[13659]_  | ~\new_[19288]_ );
  assign \new_[10712]_  = ~\new_[20825]_  | ~\new_[13418]_ ;
  assign \new_[10713]_  = \new_[13445]_  | \new_[17457]_ ;
  assign \new_[10714]_  = \new_[15685]_  & \new_[13366]_ ;
  assign \new_[10715]_  = ~\new_[15221]_  | ~\new_[14840]_ ;
  assign \new_[10716]_  = \new_[13455]_  | \new_[15530]_ ;
  assign \new_[10717]_  = ~\new_[10855]_ ;
  assign \new_[10718]_  = ~\new_[13421]_  | (~\new_[16979]_  & ~\new_[18840]_ );
  assign \new_[10719]_  = ~\new_[15692]_  | ~\new_[15710]_ ;
  assign \new_[10720]_  = ~\new_[15180]_  | ~\new_[15685]_ ;
  assign \new_[10721]_  = \new_[15665]_  | \new_[13412]_ ;
  assign \new_[10722]_  = ~\new_[15533]_  & (~\new_[17942]_  | ~\new_[18779]_ );
  assign \new_[10723]_  = \new_[13408]_  | \new_[13373]_ ;
  assign \new_[10724]_  = ~\new_[14800]_  | ~\new_[14703]_ ;
  assign \new_[10725]_  = ~\new_[15199]_  | ~\new_[14933]_ ;
  assign \new_[10726]_  = ~\new_[18994]_  | (~\new_[13513]_  & ~\new_[15435]_ );
  assign \new_[10727]_  = \new_[16053]_  | \new_[13372]_ ;
  assign \new_[10728]_  = ~\new_[13574]_  | ~\new_[14161]_  | ~\new_[20904]_ ;
  assign \new_[10729]_  = ~\new_[12079]_ ;
  assign \new_[10730]_  = \\u0_r0_out_reg[30] ;
  assign \new_[10731]_  = \\u0_r0_out_reg[31] ;
  assign \new_[10732]_  = ~\new_[17807]_  | ~\new_[12342]_ ;
  assign \new_[10733]_  = ~\new_[18209]_  | ~\new_[18179]_  | ~\new_[19308]_ ;
  assign \new_[10734]_  = ~\new_[19145]_  & (~\new_[16371]_  | ~\new_[13652]_ );
  assign \new_[10735]_  = ~\new_[11973]_ ;
  assign \new_[10736]_  = \new_[19591]_  ^ \new_[18194]_ ;
  assign \new_[10737]_  = ~\new_[11993]_ ;
  assign \new_[10738]_  = ~\new_[12095]_ ;
  assign \new_[10739]_  = ~\new_[19145]_  | (~\new_[14354]_  & ~\new_[16659]_ );
  assign \new_[10740]_  = ~\new_[16141]_  | ~\new_[17830]_  | ~\new_[12398]_  | ~\new_[13578]_ ;
  assign \new_[10741]_  = \new_[13517]_  ? \new_[17156]_  : \new_[14785]_ ;
  assign \new_[10742]_  = \new_[19175]_  ^ \new_[18187]_ ;
  assign \new_[10743]_  = \new_[13679]_  ? \new_[18076]_  : \new_[15342]_ ;
  assign \new_[10744]_  = \new_[14893]_  ^ \new_[19166]_ ;
  assign \new_[10745]_  = \new_[13521]_  ? \new_[18998]_  : \new_[14102]_ ;
  assign \new_[10746]_  = ~\new_[14927]_  | ~\new_[16173]_  | ~\new_[15607]_  | ~\new_[14303]_ ;
  assign \new_[10747]_  = ~\new_[20704]_  | (~\new_[14339]_  & ~\new_[21398]_ );
  assign \new_[10748]_  = ~\new_[18278]_  | ~\new_[18012]_  | ~\new_[14331]_ ;
  assign \new_[10749]_  = ~\new_[19006]_  | (~\new_[14048]_  & ~\new_[15915]_ );
  assign \new_[10750]_  = ~\new_[18542]_  | (~\new_[14143]_  & ~\new_[21331]_ );
  assign \new_[10751]_  = ~\new_[19064]_  | (~\new_[14098]_  & ~\new_[20233]_ );
  assign \new_[10752]_  = \new_[14785]_  ? \new_[17156]_  : \new_[13517]_ ;
  assign \new_[10753]_  = \new_[16752]_  ^ \new_[19114]_ ;
  assign \new_[10754]_  = ~\new_[12365]_  | ~\new_[19206]_ ;
  assign \new_[10755]_  = \new_[12426]_  & \new_[19727]_ ;
  assign \new_[10756]_  = ~\new_[18046]_  | (~\new_[14111]_  & ~\new_[15613]_ );
  assign \new_[10757]_  = ~\new_[21629]_  | (~\new_[14263]_  & ~\new_[13651]_ );
  assign \new_[10758]_  = ~\new_[18194]_  | (~\new_[14061]_  & ~\new_[17076]_ );
  assign \new_[10759]_  = ~\new_[19366]_  & (~\new_[14374]_  | ~\new_[16687]_ );
  assign \new_[10760]_  = ~\new_[12157]_  | ~\new_[18077]_ ;
  assign \new_[10761]_  = ~\new_[19537]_  & (~\new_[14521]_  | ~\new_[13906]_ );
  assign \new_[10762]_  = ~\new_[19300]_  & (~\new_[14481]_  | ~\new_[16237]_ );
  assign \new_[10763]_  = \new_[15850]_  ^ \new_[19373]_ ;
  assign \new_[10764]_  = ~\new_[13549]_  & ~\new_[18967]_ ;
  assign \new_[10765]_  = \new_[15632]_  | \new_[19444]_  | \new_[18795]_  | \new_[19217]_ ;
  assign \new_[10766]_  = \new_[17264]_  | \new_[17886]_  | \new_[19013]_  | \new_[16840]_ ;
  assign \new_[10767]_  = ~\new_[14729]_  | ~\new_[12732]_  | ~\new_[15524]_ ;
  assign \new_[10768]_  = ~\new_[12381]_  | ~\new_[19553]_ ;
  assign \new_[10769]_  = ~\new_[12115]_ ;
  assign \new_[10770]_  = ~\new_[20680]_  & (~\new_[15422]_  | ~\new_[14009]_ );
  assign \new_[10771]_  = \new_[15333]_  | \new_[17843]_  | \new_[18077]_  | \new_[18974]_ ;
  assign \new_[10772]_  = ~\new_[12254]_  & ~\new_[18194]_ ;
  assign \new_[10773]_  = \new_[15675]_  | \new_[21572]_  | \new_[18693]_  | \new_[18840]_ ;
  assign \new_[10774]_  = \new_[15561]_  | \new_[20699]_  | \new_[16879]_  | \new_[21508]_ ;
  assign \new_[10775]_  = ~\new_[12413]_  | ~\new_[19145]_ ;
  assign \new_[10776]_  = ~\new_[18288]_  & (~\new_[15468]_  | ~\new_[14087]_ );
  assign \new_[10777]_  = ~\new_[19021]_  & (~\new_[14884]_  | ~\new_[15253]_ );
  assign \new_[10778]_  = ~\new_[18070]_  & (~\new_[16390]_  | ~\new_[14109]_ );
  assign \new_[10779]_  = ~\new_[12290]_  | ~\new_[19064]_ ;
  assign \new_[10780]_  = \new_[12175]_  | \new_[18361]_ ;
  assign \new_[10781]_  = ~\new_[18124]_  & (~\new_[14182]_  | ~\new_[16704]_ );
  assign \new_[10782]_  = ~\new_[14178]_  | ~\new_[12178]_ ;
  assign \new_[10783]_  = ~\new_[15638]_  | ~\new_[12848]_  | ~\new_[14007]_ ;
  assign \new_[10784]_  = ~\new_[13017]_  | ~\new_[12276]_ ;
  assign \new_[10785]_  = ~\new_[14010]_  | ~\new_[12182]_ ;
  assign \new_[10786]_  = \new_[12317]_  & \new_[12551]_ ;
  assign \new_[10787]_  = ~\new_[12346]_  | ~\new_[18076]_ ;
  assign \new_[10788]_  = ~\new_[14845]_  & ~\new_[12225]_ ;
  assign \new_[10789]_  = ~\new_[12210]_  | ~\new_[14106]_ ;
  assign \new_[10790]_  = ~\new_[14333]_  | ~\new_[13549]_ ;
  assign \new_[10791]_  = ~\new_[19249]_  & (~\new_[14350]_  | ~\new_[15510]_ );
  assign \new_[10792]_  = \new_[13794]_  & \new_[12277]_ ;
  assign \new_[10793]_  = ~\new_[12189]_  | ~\new_[19553]_ ;
  assign \new_[10794]_  = \new_[12457]_  & \new_[18194]_ ;
  assign \new_[10795]_  = ~\new_[18194]_  & (~\new_[13765]_  | ~\new_[14680]_ );
  assign \new_[10796]_  = ~\new_[18821]_  & (~\new_[14071]_  | ~\new_[15315]_ );
  assign \new_[10797]_  = ~\new_[19377]_  & (~\new_[13800]_  | ~\new_[17158]_ );
  assign \new_[10798]_  = ~\new_[12330]_  | ~\new_[18795]_ ;
  assign \new_[10799]_  = ~\new_[19578]_  | (~\new_[15755]_  & ~\new_[14330]_ );
  assign \new_[10800]_  = ~\new_[12301]_  | ~\new_[12742]_ ;
  assign \new_[10801]_  = ~\new_[19261]_  & (~\new_[14639]_  | ~\new_[15652]_ );
  assign \new_[10802]_  = ~\new_[13021]_  | ~\new_[12303]_ ;
  assign \new_[10803]_  = ~\new_[15201]_  | ~\new_[13292]_  | ~\new_[14182]_ ;
  assign \new_[10804]_  = ~\new_[19215]_  & (~\new_[14118]_  | ~\new_[15959]_ );
  assign \new_[10805]_  = \new_[12476]_  | \new_[13624]_ ;
  assign \new_[10806]_  = ~\new_[14337]_  | ~\new_[12296]_ ;
  assign \new_[10807]_  = ~\new_[21466]_  | ~\new_[12206]_ ;
  assign \new_[10808]_  = ~\new_[12287]_  | ~\new_[12619]_ ;
  assign \new_[10809]_  = ~\new_[12185]_  | ~\new_[13078]_ ;
  assign \new_[10810]_  = ~\new_[13071]_  | ~\new_[13409]_ ;
  assign \new_[10811]_  = ~\new_[19659]_  | (~\new_[14647]_  & ~\new_[15284]_ );
  assign \new_[10812]_  = ~\new_[13766]_  | ~\new_[13952]_  | ~\new_[14222]_ ;
  assign \new_[10813]_  = ~\new_[18821]_  & (~\new_[13841]_  | ~\new_[14532]_ );
  assign \new_[10814]_  = ~\new_[12261]_  | ~\new_[12969]_ ;
  assign \new_[10815]_  = \new_[12216]_  & \new_[12333]_ ;
  assign \new_[10816]_  = ~\new_[19079]_  & (~\new_[13836]_  | ~\new_[16231]_ );
  assign \new_[10817]_  = ~\new_[12216]_  | ~\new_[13554]_ ;
  assign \new_[10818]_  = \\dcnt_reg[1] ;
  assign \new_[10819]_  = ~\new_[12179]_  | ~\new_[19547]_ ;
  assign \new_[10820]_  = ~\new_[13566]_  | ~\new_[12181]_ ;
  assign \new_[10821]_  = ~\new_[12229]_  | ~\new_[15354]_ ;
  assign \new_[10822]_  = ~\new_[12481]_  | ~\new_[16338]_ ;
  assign \new_[10823]_  = ~\new_[15496]_  | ~\new_[12232]_ ;
  assign \new_[10824]_  = ~\new_[16900]_  | ~\new_[12993]_  | ~\new_[15046]_ ;
  assign \new_[10825]_  = ~\new_[12233]_  | ~\new_[20866]_ ;
  assign \new_[10826]_  = ~\new_[19748]_  | (~\new_[14635]_  & ~\new_[15178]_ );
  assign \new_[10827]_  = ~\new_[14810]_  | ~\new_[13681]_  | ~\new_[13866]_ ;
  assign \new_[10828]_  = ~\new_[13081]_  | ~\new_[12390]_ ;
  assign \new_[10829]_  = ~\new_[19587]_  & (~\new_[14426]_  | ~\new_[13884]_ );
  assign \new_[10830]_  = ~\new_[12156]_  | ~\new_[13868]_ ;
  assign \new_[10831]_  = ~\new_[19059]_  & (~\new_[13995]_  | ~\new_[15466]_ );
  assign \new_[10832]_  = ~\new_[12471]_  & ~\new_[19085]_ ;
  assign \new_[10833]_  = ~\new_[12139]_ ;
  assign \new_[10834]_  = \new_[12152]_  | \new_[20100]_ ;
  assign \new_[10835]_  = ~\new_[16879]_  & (~\new_[14234]_  | ~\new_[15885]_ );
  assign \new_[10836]_  = ~\new_[17917]_  | ~\new_[20663]_ ;
  assign \new_[10837]_  = ~\new_[19711]_  & (~\new_[14245]_  | ~\new_[15622]_ );
  assign \new_[10838]_  = \new_[12418]_  | \new_[19021]_ ;
  assign \new_[10839]_  = ~\new_[19006]_  | (~\new_[14145]_  & ~\new_[15848]_ );
  assign \new_[10840]_  = ~\new_[18443]_  & (~\new_[16770]_  | ~\new_[13802]_ );
  assign \new_[10841]_  = ~\new_[12394]_  | ~\new_[12258]_ ;
  assign \new_[10842]_  = ~\new_[13655]_  | ~\new_[12324]_ ;
  assign \new_[10843]_  = ~\new_[19261]_  & (~\new_[13771]_  | ~\new_[16671]_ );
  assign \new_[10844]_  = ~\new_[21634]_  & (~\new_[14431]_  | ~\new_[14977]_ );
  assign \new_[10845]_  = ~\new_[21115]_  & (~\new_[14352]_  | ~\new_[14720]_ );
  assign \new_[10846]_  = ~\new_[19157]_  | (~\new_[15734]_  & ~\new_[15288]_ );
  assign \new_[10847]_  = ~\new_[15289]_  | ~\new_[13862]_  | ~\new_[16824]_ ;
  assign \new_[10848]_  = ~\new_[21267]_  | (~\new_[16541]_  & ~\new_[15270]_ );
  assign \new_[10849]_  = ~\new_[13595]_  | ~\new_[15298]_ ;
  assign \new_[10850]_  = ~\new_[13004]_ ;
  assign \new_[10851]_  = ~\new_[19687]_  & (~\new_[15113]_  | ~\new_[16218]_ );
  assign \new_[10852]_  = ~\new_[13585]_  | ~\new_[14019]_ ;
  assign \new_[10853]_  = ~\new_[12148]_ ;
  assign \new_[10854]_  = ~\new_[19299]_  & (~\new_[15014]_  | ~\new_[16150]_ );
  assign \new_[10855]_  = ~\new_[16092]_  | ~\new_[19068]_ ;
  assign \new_[10856]_  = ~\new_[14367]_  | ~\new_[13601]_ ;
  assign \new_[10857]_  = \\u0_r0_out_reg[24] ;
  assign \new_[10858]_  = ~\new_[18343]_  | ~\new_[13518]_ ;
  assign \new_[10859]_  = ~\new_[13660]_  & ~\new_[19239]_ ;
  assign \new_[10860]_  = ~\new_[16680]_  & ~\new_[13564]_ ;
  assign \new_[10861]_  = ~\new_[16095]_  | ~\new_[19181]_ ;
  assign \new_[10862]_  = ~\new_[12160]_ ;
  assign \new_[10863]_  = ~\new_[13674]_  | ~\new_[18998]_ ;
  assign \new_[10864]_  = \new_[15628]_  | \new_[14470]_ ;
  assign \new_[10865]_  = ~\new_[19202]_  & (~\new_[15395]_  | ~\new_[16101]_ );
  assign \new_[10866]_  = ~\new_[18821]_  & (~\new_[15454]_  | ~\new_[16675]_ );
  assign \new_[10867]_  = ~\new_[19249]_  & (~\new_[16178]_  | ~\new_[15003]_ );
  assign \new_[10868]_  = ~\new_[19059]_  & (~\new_[15440]_  | ~\new_[21622]_ );
  assign \new_[10869]_  = ~\new_[15003]_  | ~\new_[14992]_  | ~\new_[14819]_ ;
  assign \new_[10870]_  = ~\new_[16033]_  & ~\new_[13553]_ ;
  assign \new_[10871]_  = ~\new_[19145]_  & (~\new_[15198]_  | ~\new_[17180]_ );
  assign \new_[10872]_  = ~\new_[14919]_  | ~\new_[13835]_  | ~\new_[16014]_ ;
  assign \new_[10873]_  = ~\new_[15231]_  | ~\new_[15067]_  | ~\new_[15886]_ ;
  assign \new_[10874]_  = ~\new_[13670]_  & (~\new_[15827]_  | ~\new_[15654]_ );
  assign \new_[10875]_  = \new_[14108]_  & \new_[13661]_ ;
  assign \new_[10876]_  = ~\new_[17082]_  | ~\new_[15970]_ ;
  assign \new_[10877]_  = (~\new_[16019]_  | ~\new_[19228]_ ) & (~\new_[15476]_  | ~\new_[18938]_ );
  assign \new_[10878]_  = ~\new_[15307]_  | ~\new_[13655]_ ;
  assign \new_[10879]_  = ~\new_[14187]_  & (~\new_[15701]_  | ~\new_[15892]_ );
  assign \new_[10880]_  = \new_[14100]_  & \new_[21638]_ ;
  assign \new_[10881]_  = \new_[14348]_  & \new_[20100]_ ;
  assign \new_[10882]_  = \new_[14406]_  & \new_[15483]_ ;
  assign \new_[10883]_  = ~\new_[12173]_ ;
  assign \new_[10884]_  = \new_[18264]_  | \new_[16679]_  | \new_[19791]_  | \new_[21574]_ ;
  assign \new_[10885]_  = ~\new_[17651]_  | ~\new_[21580]_  | ~\new_[21508]_  | ~\new_[20699]_ ;
  assign \new_[10886]_  = ~\new_[13644]_  & ~\new_[18046]_ ;
  assign \new_[10887]_  = ~\new_[16601]_  | ~\new_[21658]_  | ~\new_[19261]_  | ~\new_[18328]_ ;
  assign \new_[10888]_  = \new_[13845]_  & \new_[19727]_ ;
  assign \new_[10889]_  = \new_[16088]_  | \new_[18567]_  | \new_[19266]_  | \new_[19269]_ ;
  assign \new_[10890]_  = ~\new_[14004]_  & ~\new_[19261]_ ;
  assign \new_[10891]_  = ~\new_[14087]_  & ~\new_[20680]_ ;
  assign \new_[10892]_  = ~\new_[14178]_  & ~\new_[19224]_ ;
  assign \new_[10893]_  = ~\new_[13989]_  & ~\new_[20865]_ ;
  assign \new_[10894]_  = \new_[14379]_  | \new_[19711]_ ;
  assign \new_[10895]_  = ~\new_[14371]_  & ~\new_[18166]_ ;
  assign \new_[10896]_  = ~\new_[19554]_  | ~\new_[19068]_  | ~\new_[16027]_ ;
  assign \new_[10897]_  = ~\new_[19386]_  | ~\new_[17598]_  | ~\new_[15521]_ ;
  assign \new_[10898]_  = ~\new_[13973]_  & ~\new_[18166]_ ;
  assign \new_[10899]_  = ~\new_[14420]_  & ~\new_[18209]_ ;
  assign \new_[10900]_  = ~\new_[13540]_  | ~\new_[19153]_ ;
  assign \new_[10901]_  = ~\new_[12184]_ ;
  assign \new_[10902]_  = \new_[13578]_  | \new_[19727]_ ;
  assign \new_[10903]_  = ~\new_[13489]_  | ~\new_[18893]_ ;
  assign \new_[10904]_  = ~\new_[12188]_ ;
  assign \new_[10905]_  = ~\new_[14001]_  | ~\new_[19290]_ ;
  assign \new_[10906]_  = ~\new_[13762]_  & ~\new_[19754]_ ;
  assign \new_[10907]_  = ~\new_[17490]_  | ~\new_[21056]_  | ~\new_[17886]_  | ~\new_[18111]_ ;
  assign \new_[10908]_  = ~\new_[13525]_  & ~\new_[21496]_ ;
  assign \new_[10909]_  = ~\new_[13742]_  | ~\new_[18414]_ ;
  assign \new_[10910]_  = ~\new_[14414]_  & ~\new_[19253]_ ;
  assign \new_[10911]_  = ~\new_[12191]_ ;
  assign \new_[10912]_  = \new_[14076]_  | \new_[19553]_ ;
  assign \new_[10913]_  = ~\new_[13882]_  & ~\new_[21695]_ ;
  assign \new_[10914]_  = ~\new_[12192]_ ;
  assign \new_[10915]_  = ~\new_[13602]_  | ~\new_[21686]_ ;
  assign \new_[10916]_  = ~\new_[14039]_  | ~\new_[18076]_ ;
  assign \new_[10917]_  = \new_[13883]_  | \new_[18194]_ ;
  assign \new_[10918]_  = ~\new_[12194]_ ;
  assign \new_[10919]_  = ~\new_[14598]_  & ~\new_[19064]_ ;
  assign \new_[10920]_  = ~\new_[12195]_ ;
  assign \new_[10921]_  = ~\new_[16608]_  | ~\new_[18264]_  | ~\new_[18621]_  | ~\new_[21574]_ ;
  assign \new_[10922]_  = ~\new_[13791]_  | ~\new_[19687]_ ;
  assign \new_[10923]_  = ~\new_[13927]_  & ~\new_[18832]_ ;
  assign \new_[10924]_  = ~\new_[14391]_  & ~\new_[18832]_ ;
  assign \new_[10925]_  = ~\new_[12198]_ ;
  assign \new_[10926]_  = ~\new_[12200]_ ;
  assign \new_[10927]_  = ~\new_[12201]_ ;
  assign \new_[10928]_  = ~\new_[14104]_  & ~\new_[19589]_ ;
  assign \new_[10929]_  = ~\new_[14661]_  | ~\new_[19288]_ ;
  assign \new_[10930]_  = \new_[13745]_  & \new_[19253]_ ;
  assign \new_[10931]_  = ~\new_[16104]_  | ~\new_[18965]_ ;
  assign \new_[10932]_  = ~\new_[12203]_ ;
  assign \new_[10933]_  = ~\new_[16799]_  | ~\new_[19249]_  | ~\new_[18115]_ ;
  assign \new_[10934]_  = ~\new_[14016]_  & ~\new_[18166]_ ;
  assign \new_[10935]_  = ~\new_[12205]_ ;
  assign \new_[10936]_  = ~\new_[21666]_ ;
  assign \new_[10937]_  = ~\new_[21665]_ ;
  assign \new_[10938]_  = ~\new_[14367]_  & ~\new_[19084]_ ;
  assign \new_[10939]_  = ~\new_[14026]_  | ~\new_[18938]_ ;
  assign \new_[10940]_  = ~\new_[14070]_  & ~\new_[19239]_ ;
  assign \new_[10941]_  = ~\new_[13602]_  | ~\new_[19261]_ ;
  assign \new_[10942]_  = ~\new_[14091]_  | ~\new_[18187]_ ;
  assign \new_[10943]_  = \new_[13643]_  & \new_[19239]_ ;
  assign \new_[10944]_  = ~\new_[14096]_  & (~\new_[16653]_  | ~\new_[19152]_ );
  assign \new_[10945]_  = ~\new_[13957]_  & ~\new_[19239]_ ;
  assign \new_[10946]_  = ~\new_[14112]_  | ~\new_[19269]_ ;
  assign \new_[10947]_  = ~\new_[14827]_  | ~\new_[21634]_  | ~\new_[18869]_ ;
  assign \new_[10948]_  = ~\new_[19553]_  | ~\new_[13745]_ ;
  assign \new_[10949]_  = ~\new_[14134]_  & ~\new_[18046]_ ;
  assign \new_[10950]_  = ~\new_[13797]_  & ~\new_[20492]_ ;
  assign \new_[10951]_  = \new_[13718]_  & \new_[19240]_ ;
  assign \new_[10952]_  = ~\new_[15056]_  & ~\new_[14326]_ ;
  assign \new_[10953]_  = ~\new_[13805]_  & ~\new_[18076]_ ;
  assign \new_[10954]_  = ~\new_[14327]_  | ~\new_[19253]_ ;
  assign \new_[10955]_  = ~\new_[14066]_  & ~\new_[18194]_ ;
  assign \new_[10956]_  = ~\new_[18833]_  | ~\new_[13736]_ ;
  assign \new_[10957]_  = ~\new_[19082]_  & ~\new_[13647]_ ;
  assign \new_[10958]_  = ~\new_[13769]_  & ~\new_[19084]_ ;
  assign \new_[10959]_  = ~\new_[12219]_ ;
  assign \new_[10960]_  = \new_[16186]_  | \new_[21515]_  | \new_[19154]_  | \new_[18637]_ ;
  assign \new_[10961]_  = ~\new_[21706]_  & ~\new_[18083]_ ;
  assign \new_[10962]_  = \new_[13798]_  | \new_[19115]_ ;
  assign \new_[10963]_  = \new_[19742]_  | \new_[13832]_ ;
  assign \new_[10964]_  = ~\new_[12222]_ ;
  assign \new_[10965]_  = ~\new_[12222]_ ;
  assign \new_[10966]_  = ~\new_[12225]_ ;
  assign \new_[10967]_  = ~\new_[14043]_  | ~\new_[19727]_ ;
  assign \new_[10968]_  = ~\new_[14679]_  | ~\new_[18569]_ ;
  assign \new_[10969]_  = ~\new_[12226]_ ;
  assign \new_[10970]_  = ~\new_[13785]_  & ~\new_[18778]_ ;
  assign \new_[10971]_  = ~\new_[13739]_  & ~\new_[19158]_ ;
  assign \new_[10972]_  = \new_[19727]_  | \new_[13890]_ ;
  assign \new_[10973]_  = ~\new_[14471]_  | ~\new_[18209]_ ;
  assign \new_[10974]_  = \new_[19269]_  | \new_[14013]_ ;
  assign \new_[10975]_  = ~\new_[13731]_  & ~\new_[18605]_ ;
  assign \new_[10976]_  = ~\new_[14193]_  | ~\new_[19268]_ ;
  assign \new_[10977]_  = ~\new_[14132]_  | ~\new_[19050]_ ;
  assign \new_[10978]_  = ~\new_[14184]_  & ~\new_[18938]_ ;
  assign \new_[10979]_  = ~\new_[14336]_  & ~\new_[18285]_ ;
  assign \new_[10980]_  = ~\new_[14202]_  & ~\new_[18285]_ ;
  assign \new_[10981]_  = ~\new_[18337]_  | ~\new_[19095]_  | ~\new_[15209]_ ;
  assign \new_[10982]_  = ~\new_[14208]_  & ~\new_[21631]_ ;
  assign \new_[10983]_  = ~\new_[14308]_  & ~\new_[18325]_ ;
  assign \new_[10984]_  = ~\new_[13861]_  & ~\new_[19181]_ ;
  assign \new_[10985]_  = ~\new_[13681]_  & ~\new_[18678]_ ;
  assign \new_[10986]_  = \new_[19610]_  ^ \new_[19561]_ ;
  assign \new_[10987]_  = ~\new_[12240]_ ;
  assign \new_[10988]_  = \new_[19381]_  | \new_[13975]_ ;
  assign \new_[10989]_  = ~\new_[14588]_  & ~\new_[19357]_ ;
  assign \new_[10990]_  = ~\new_[21095]_  & ~\new_[18124]_ ;
  assign \new_[10991]_  = ~\new_[12241]_ ;
  assign \new_[10992]_  = ~\new_[13880]_  | ~\new_[19085]_ ;
  assign \new_[10993]_  = \new_[19202]_  | \new_[14044]_ ;
  assign \new_[10994]_  = ~\new_[12243]_ ;
  assign \new_[10995]_  = ~\new_[13706]_  & ~\new_[19214]_ ;
  assign \new_[10996]_  = ~\new_[13943]_  & ~\new_[18285]_ ;
  assign \new_[10997]_  = ~\new_[14214]_  | ~\new_[21505]_ ;
  assign \new_[10998]_  = \new_[16017]_  | \new_[19398]_  | \new_[19612]_  | \new_[19446]_ ;
  assign \new_[10999]_  = ~\new_[13992]_  & ~\new_[21558]_ ;
  assign \new_[11000]_  = ~\new_[14239]_  & ~\new_[21562]_ ;
  assign \new_[11001]_  = ~\new_[14109]_  & ~\new_[19357]_ ;
  assign \new_[11002]_  = ~\new_[13528]_  | ~\new_[19021]_ ;
  assign \new_[11003]_  = ~\new_[13526]_  & ~\new_[18969]_ ;
  assign \new_[11004]_  = ~\new_[12698]_ ;
  assign \new_[11005]_  = ~\new_[13872]_  & ~\new_[19024]_ ;
  assign \new_[11006]_  = ~\new_[14248]_  & ~\new_[18778]_ ;
  assign \new_[11007]_  = ~\new_[14112]_  | ~\new_[18798]_ ;
  assign \new_[11008]_  = ~\new_[20966]_  & ~\new_[19687]_ ;
  assign \new_[11009]_  = ~\new_[13959]_  & ~\new_[19476]_ ;
  assign \new_[11010]_  = ~\new_[13579]_  & ~\new_[19050]_ ;
  assign \new_[11011]_  = ~\new_[13863]_  & ~\new_[19681]_ ;
  assign \new_[11012]_  = ~\new_[14226]_  & ~\new_[19196]_ ;
  assign \new_[11013]_  = ~\new_[12254]_ ;
  assign \new_[11014]_  = ~\new_[21412]_  | ~\new_[19094]_ ;
  assign \new_[11015]_  = ~\new_[13575]_  | ~\new_[21631]_ ;
  assign \new_[11016]_  = ~\new_[12257]_ ;
  assign \new_[11017]_  = \new_[13804]_  | \new_[19476]_ ;
  assign \new_[11018]_  = ~\new_[14170]_  & ~\new_[18941]_ ;
  assign \new_[11019]_  = ~\new_[19095]_  & ~\new_[14346]_ ;
  assign \new_[11020]_  = ~\new_[12259]_ ;
  assign \new_[11021]_  = ~\new_[12261]_ ;
  assign \new_[11022]_  = ~\new_[14033]_  & ~\new_[19095]_ ;
  assign \new_[11023]_  = ~\new_[12263]_ ;
  assign \new_[11024]_  = ~\new_[12267]_ ;
  assign \new_[11025]_  = ~\new_[12268]_ ;
  assign \new_[11026]_  = ~\new_[13781]_  & ~\new_[17979]_ ;
  assign \new_[11027]_  = \new_[13917]_  & \new_[19021]_ ;
  assign \new_[11028]_  = ~\new_[13717]_  & ~\new_[18973]_ ;
  assign \new_[11029]_  = \new_[13814]_  & \new_[19233]_ ;
  assign \new_[11030]_  = ~\new_[12275]_ ;
  assign \new_[11031]_  = ~\new_[13981]_  | ~\new_[18046]_ ;
  assign \new_[11032]_  = \new_[13664]_  & \new_[21634]_ ;
  assign \new_[11033]_  = ~\new_[14110]_  & ~\new_[19687]_ ;
  assign \new_[11034]_  = \new_[14038]_  | \new_[19299]_ ;
  assign \new_[11035]_  = ~\new_[13801]_  & ~\new_[21502]_ ;
  assign \new_[11036]_  = ~\new_[13730]_  | ~\new_[19547]_ ;
  assign \new_[11037]_  = \new_[14123]_  | \new_[18414]_ ;
  assign \new_[11038]_  = ~\new_[14290]_  | ~\new_[19253]_ ;
  assign \new_[11039]_  = ~\new_[13743]_  & ~\new_[21056]_ ;
  assign \new_[11040]_  = \new_[19249]_  | \new_[13820]_ ;
  assign \new_[11041]_  = \new_[13510]_  | \new_[19079]_ ;
  assign \new_[11042]_  = ~\new_[14010]_  & ~\new_[18008]_ ;
  assign \new_[11043]_  = ~\new_[13798]_  & ~\new_[19697]_ ;
  assign \new_[11044]_  = ~\new_[14238]_  & ~\new_[21056]_ ;
  assign \new_[11045]_  = ~\new_[12277]_ ;
  assign \new_[11046]_  = ~\new_[12279]_ ;
  assign \new_[11047]_  = \new_[19239]_  | \new_[13958]_ ;
  assign \new_[11048]_  = ~\new_[14295]_  & ~\new_[21115]_ ;
  assign \new_[11049]_  = ~\new_[13792]_  | ~\new_[19102]_ ;
  assign \new_[11050]_  = ~\new_[14289]_  & ~\new_[14951]_ ;
  assign \new_[11051]_  = ~\new_[12281]_ ;
  assign \new_[11052]_  = ~\new_[13818]_  & ~\new_[21635]_ ;
  assign \new_[11053]_  = ~\new_[13532]_  & ~\new_[19013]_ ;
  assign \new_[11054]_  = ~\new_[14063]_  & ~\new_[19319]_ ;
  assign \new_[11055]_  = ~\new_[13512]_  & ~\new_[18166]_ ;
  assign \new_[11056]_  = ~\new_[12284]_ ;
  assign \new_[11057]_  = ~\new_[14159]_  & ~\new_[21502]_ ;
  assign \new_[11058]_  = \new_[13609]_  | \new_[19288]_ ;
  assign \new_[11059]_  = ~\new_[14283]_  & ~\new_[19247]_ ;
  assign \new_[11060]_  = ~\new_[13754]_  & ~\new_[18209]_ ;
  assign \new_[11061]_  = ~\new_[13520]_  | ~\new_[19249]_ ;
  assign \new_[11062]_  = ~\new_[13780]_  & ~\new_[21692]_ ;
  assign \new_[11063]_  = ~\new_[14042]_  & ~\new_[18621]_ ;
  assign \new_[11064]_  = ~\new_[12285]_ ;
  assign \new_[11065]_  = ~\new_[13625]_  & ~\new_[18984]_ ;
  assign \new_[11066]_  = \new_[20158]_  | \new_[19028]_ ;
  assign \new_[11067]_  = ~\new_[12286]_ ;
  assign \new_[11068]_  = ~\new_[14067]_  & ~\new_[21689]_ ;
  assign \new_[11069]_  = ~\new_[13707]_  | ~\new_[19094]_ ;
  assign \new_[11070]_  = ~\new_[14609]_  & ~\new_[18083]_ ;
  assign \new_[11071]_  = ~\new_[13983]_  & ~\new_[19249]_ ;
  assign \new_[11072]_  = ~\new_[13961]_  & ~\new_[18083]_ ;
  assign \new_[11073]_  = ~\new_[13966]_  | ~\new_[18187]_ ;
  assign \new_[11074]_  = ~\new_[13721]_  & ~\new_[19269]_ ;
  assign \new_[11075]_  = ~\new_[13753]_  & ~\new_[21500]_ ;
  assign \new_[11076]_  = ~\new_[12289]_ ;
  assign \new_[11077]_  = ~\new_[13935]_  & ~\new_[19068]_ ;
  assign \new_[11078]_  = ~\new_[21502]_  & ~\new_[14201]_ ;
  assign \new_[11079]_  = ~\new_[14677]_  | ~\new_[16262]_ ;
  assign \new_[11080]_  = ~\new_[14182]_  | ~\new_[15201]_ ;
  assign \new_[11081]_  = ~\new_[13501]_  | ~\new_[14325]_ ;
  assign \new_[11082]_  = ~\new_[12290]_ ;
  assign \new_[11083]_  = ~\new_[20864]_ ;
  assign \new_[11084]_  = ~\new_[14094]_  | ~\new_[18402]_ ;
  assign \new_[11085]_  = ~\new_[14127]_  | ~\new_[19156]_ ;
  assign \new_[11086]_  = ~\new_[12293]_ ;
  assign \new_[11087]_  = ~\new_[13702]_  | ~\new_[21685]_ ;
  assign \new_[11088]_  = ~\new_[13910]_  & ~\new_[21688]_ ;
  assign \new_[11089]_  = ~\new_[14201]_  | ~\new_[17311]_ ;
  assign \new_[11090]_  = ~\new_[13855]_  | ~\new_[14210]_ ;
  assign \new_[11091]_  = ~\new_[12294]_ ;
  assign \new_[11092]_  = ~\new_[14630]_  | ~\new_[13882]_ ;
  assign \new_[11093]_  = ~\new_[14664]_  | ~\new_[16180]_ ;
  assign \new_[11094]_  = ~\new_[14006]_  | ~\new_[19224]_ ;
  assign \new_[11095]_  = ~\new_[13711]_  | ~\new_[19269]_ ;
  assign \new_[11096]_  = ~\new_[14007]_  | ~\new_[15638]_ ;
  assign \new_[11097]_  = \new_[19727]_  | \new_[13635]_ ;
  assign \new_[11098]_  = ~\new_[14268]_  & ~\new_[18421]_ ;
  assign \new_[11099]_  = ~\new_[21714]_  | ~\new_[13696]_ ;
  assign \new_[11100]_  = ~\new_[15252]_  | ~\new_[20239]_ ;
  assign \new_[11101]_  = ~\new_[14626]_  | ~\new_[13721]_ ;
  assign \new_[11102]_  = ~\new_[12302]_ ;
  assign \new_[11103]_  = ~\new_[13707]_  | ~\new_[18825]_ ;
  assign \new_[11104]_  = ~\new_[14605]_  | ~\new_[14141]_ ;
  assign \new_[11105]_  = ~\new_[12305]_ ;
  assign \new_[11106]_  = ~\new_[13787]_  | ~\new_[14329]_ ;
  assign \new_[11107]_  = \new_[14147]_  | \new_[19547]_ ;
  assign \new_[11108]_  = ~\new_[15744]_  | ~\new_[13935]_ ;
  assign \new_[11109]_  = \new_[14242]_  & \new_[13957]_ ;
  assign \new_[11110]_  = ~\new_[12306]_ ;
  assign \new_[11111]_  = ~\new_[12307]_ ;
  assign \new_[11112]_  = ~\new_[12310]_ ;
  assign \new_[11113]_  = ~\new_[14023]_  & ~\new_[19156]_ ;
  assign \new_[11114]_  = ~\new_[14007]_  | ~\new_[14087]_ ;
  assign \new_[11115]_  = ~\new_[14002]_  | ~\new_[17209]_ ;
  assign \new_[11116]_  = ~\new_[18891]_  | ~\new_[14314]_ ;
  assign \new_[11117]_  = ~\new_[15047]_  | ~\new_[18773]_ ;
  assign \new_[11118]_  = ~\new_[12311]_ ;
  assign \new_[11119]_  = ~\new_[12313]_ ;
  assign \new_[11120]_  = ~\new_[14942]_  | ~\new_[13813]_ ;
  assign \new_[11121]_  = ~\new_[14215]_  | ~\new_[13787]_ ;
  assign \new_[11122]_  = \new_[13766]_  | \new_[19290]_ ;
  assign \new_[11123]_  = ~\new_[14680]_  | ~\new_[16714]_ ;
  assign \new_[11124]_  = ~\new_[13571]_  & ~\new_[19319]_ ;
  assign \new_[11125]_  = ~\new_[14412]_  & ~\new_[19008]_ ;
  assign \new_[11126]_  = ~\new_[18194]_  | ~\new_[15900]_ ;
  assign \new_[11127]_  = ~\new_[17064]_  & (~\new_[16399]_  | ~\new_[16177]_ );
  assign \new_[11128]_  = ~\new_[12318]_ ;
  assign \new_[11129]_  = ~\new_[16879]_  & ~\new_[13744]_ ;
  assign \new_[11130]_  = \new_[13811]_  & \new_[17979]_ ;
  assign \new_[11131]_  = ~\new_[14634]_  | ~\new_[13731]_ ;
  assign \new_[11132]_  = ~\new_[14049]_  & ~\new_[19253]_ ;
  assign \new_[11133]_  = ~\new_[13986]_  | ~\new_[14054]_ ;
  assign \new_[11134]_  = ~\new_[12321]_ ;
  assign \new_[11135]_  = \new_[14094]_  & \new_[18414]_ ;
  assign \new_[11136]_  = ~\new_[13682]_  | ~\new_[14109]_ ;
  assign \new_[11137]_  = ~\new_[16547]_  | ~\new_[13781]_ ;
  assign \new_[11138]_  = ~\new_[14493]_  | ~\new_[14103]_ ;
  assign \new_[11139]_  = ~\new_[17231]_  | ~\new_[14225]_ ;
  assign \new_[11140]_  = ~\new_[14680]_  | ~\new_[14049]_ ;
  assign \new_[11141]_  = ~\new_[15705]_  | ~\new_[14037]_ ;
  assign \new_[11142]_  = ~\new_[17175]_  | ~\new_[16177]_  | ~\new_[14717]_ ;
  assign \new_[11143]_  = \new_[14409]_  & \new_[18606]_ ;
  assign \new_[11144]_  = ~\new_[12326]_ ;
  assign \new_[11145]_  = ~\new_[12386]_ ;
  assign \new_[11146]_  = ~\new_[14293]_  & ~\new_[19145]_ ;
  assign \new_[11147]_  = ~\new_[12327]_ ;
  assign \new_[11148]_  = ~\new_[19064]_  & ~\new_[16455]_ ;
  assign \new_[11149]_  = \new_[13805]_  & \new_[14315]_ ;
  assign \new_[11150]_  = ~\new_[12328]_ ;
  assign \new_[11151]_  = ~\new_[12329]_ ;
  assign \new_[11152]_  = ~\new_[12330]_ ;
  assign \new_[11153]_  = ~\new_[14271]_  & ~\new_[18179]_ ;
  assign \new_[11154]_  = ~\new_[13282]_ ;
  assign \new_[11155]_  = ~\new_[13635]_  & ~\new_[19290]_ ;
  assign \new_[11156]_  = ~\new_[12333]_ ;
  assign \new_[11157]_  = ~\new_[14243]_  | ~\new_[14231]_ ;
  assign \new_[11158]_  = ~\new_[14209]_  | ~\new_[18938]_ ;
  assign \new_[11159]_  = \new_[13925]_  | \new_[18194]_ ;
  assign \new_[11160]_  = ~\new_[13822]_  & ~\new_[17689]_ ;
  assign \new_[11161]_  = ~\new_[14616]_  | ~\new_[21684]_ ;
  assign \new_[11162]_  = \new_[13819]_  & \new_[15441]_ ;
  assign \new_[11163]_  = ~\new_[15370]_  | ~\new_[19204]_ ;
  assign \new_[11164]_  = ~\new_[12336]_ ;
  assign \new_[11165]_  = \new_[13516]_  & \new_[19547]_ ;
  assign \new_[11166]_  = ~\new_[12338]_ ;
  assign \new_[11167]_  = ~\new_[14985]_  | ~\new_[14381]_ ;
  assign \new_[11168]_  = ~\new_[13877]_  & ~\new_[14065]_ ;
  assign \new_[11169]_  = ~\new_[14217]_  | ~\new_[13858]_ ;
  assign \new_[11170]_  = ~\new_[16240]_  | ~\new_[19268]_ ;
  assign \new_[11171]_  = ~\new_[13696]_  | ~\new_[16455]_ ;
  assign \new_[11172]_  = ~\new_[17104]_  | ~\new_[13680]_ ;
  assign \new_[11173]_  = ~\new_[15042]_  | ~\new_[16188]_ ;
  assign \new_[11174]_  = ~\new_[13994]_  & ~\new_[14261]_ ;
  assign \new_[11175]_  = ~\new_[13879]_  | ~\new_[19410]_ ;
  assign \new_[11176]_  = ~\new_[13904]_  & ~\new_[15047]_ ;
  assign \new_[11177]_  = ~\new_[13994]_  & ~\new_[14695]_ ;
  assign \new_[11178]_  = ~\new_[12315]_ ;
  assign \new_[11179]_  = ~\new_[14117]_  & ~\new_[18209]_ ;
  assign \new_[11180]_  = ~\new_[12344]_ ;
  assign \new_[11181]_  = ~\new_[12346]_ ;
  assign \new_[11182]_  = \new_[13696]_  | \new_[20865]_ ;
  assign \new_[11183]_  = ~\new_[13938]_  & ~\new_[18443]_ ;
  assign \new_[11184]_  = ~\new_[14646]_  | ~\new_[21634]_ ;
  assign \new_[11185]_  = ~\new_[18972]_  & ~\new_[14293]_ ;
  assign \new_[11186]_  = ~\new_[14185]_  & ~\new_[14169]_ ;
  assign \new_[11187]_  = ~\new_[16069]_  | ~\new_[18076]_ ;
  assign \new_[11188]_  = ~\new_[13756]_  | ~\new_[18199]_ ;
  assign \new_[11189]_  = ~\new_[15260]_  & ~\new_[14001]_ ;
  assign \new_[11190]_  = ~\new_[12349]_ ;
  assign \new_[11191]_  = ~\new_[21615]_ ;
  assign \new_[11192]_  = ~\new_[13837]_  & ~\new_[20485]_ ;
  assign \new_[11193]_  = ~\new_[14127]_  | ~\new_[19742]_ ;
  assign \new_[11194]_  = ~\new_[14322]_  | ~\new_[13510]_ ;
  assign \new_[11195]_  = ~\new_[17057]_  | ~\new_[14423]_  | ~\new_[17242]_ ;
  assign \new_[11196]_  = ~\new_[19625]_  & ~\new_[14268]_ ;
  assign \new_[11197]_  = \new_[15638]_  & \new_[13802]_ ;
  assign \new_[11198]_  = ~\new_[12359]_ ;
  assign \new_[11199]_  = ~\new_[16098]_  & ~\new_[14174]_ ;
  assign \new_[11200]_  = ~\new_[15137]_  | ~\new_[13769]_ ;
  assign \new_[11201]_  = \new_[13850]_  & \new_[13727]_ ;
  assign \new_[11202]_  = ~\new_[14028]_  | ~\new_[19269]_ ;
  assign \new_[11203]_  = ~\new_[12360]_ ;
  assign \new_[11204]_  = ~\new_[14271]_  & ~\new_[19815]_ ;
  assign \new_[11205]_  = ~\new_[13510]_  | ~\new_[13746]_ ;
  assign \new_[11206]_  = ~\new_[16586]_  | ~\new_[14293]_ ;
  assign \new_[11207]_  = ~\new_[13856]_  | ~\new_[18421]_ ;
  assign \new_[11208]_  = ~\new_[21257]_  | ~\new_[13510]_ ;
  assign \new_[11209]_  = ~\new_[13814]_  | ~\new_[18909]_ ;
  assign \new_[11210]_  = \new_[18262]_  & \new_[13736]_ ;
  assign \new_[11211]_  = ~\new_[14203]_  | ~\new_[18124]_ ;
  assign \new_[11212]_  = ~\new_[15045]_  | ~\new_[19153]_ ;
  assign \new_[11213]_  = ~\new_[12168]_ ;
  assign \new_[11214]_  = ~\new_[16858]_  | ~\new_[14336]_ ;
  assign \new_[11215]_  = \new_[13716]_  | \new_[19253]_ ;
  assign \new_[11216]_  = ~\new_[12366]_ ;
  assign \new_[11217]_  = ~\new_[12367]_ ;
  assign \new_[11218]_  = ~\new_[12368]_ ;
  assign \new_[11219]_  = ~\new_[12369]_ ;
  assign \new_[11220]_  = ~\new_[14304]_  & ~\new_[18637]_ ;
  assign \new_[11221]_  = ~\new_[19258]_  & ~\new_[13579]_ ;
  assign \new_[11222]_  = \new_[13850]_  & \new_[16748]_ ;
  assign \new_[11223]_  = ~\new_[13911]_  | ~\new_[21634]_ ;
  assign \new_[11224]_  = ~\new_[21391]_  | ~\new_[14359]_ ;
  assign \new_[11225]_  = ~\new_[18325]_  & ~\new_[14152]_ ;
  assign \new_[11226]_  = ~\new_[13862]_  | ~\new_[14211]_ ;
  assign \new_[11227]_  = ~\new_[14075]_  | ~\new_[18606]_ ;
  assign \new_[11228]_  = ~\new_[13816]_  & ~\new_[21692]_ ;
  assign \new_[11229]_  = ~\new_[16998]_  | ~\new_[14393]_ ;
  assign n2728 = ~\new_[19363]_  & ~\new_[14095]_  & ~\new_[19723]_ ;
  assign \new_[11231]_  = ~\new_[13530]_  | ~\new_[13796]_ ;
  assign \new_[11232]_  = ~\new_[15073]_  | ~\new_[13849]_ ;
  assign \new_[11233]_  = ~\new_[12156]_ ;
  assign \new_[11234]_  = ~\new_[13785]_  | ~\new_[13709]_ ;
  assign \new_[11235]_  = \new_[14353]_  & \new_[14147]_ ;
  assign \new_[11236]_  = ~\new_[19687]_  & (~\new_[17317]_  | ~\new_[15609]_ );
  assign \new_[11237]_  = ~\new_[12372]_ ;
  assign \new_[11238]_  = ~\new_[18124]_  & ~\new_[14206]_ ;
  assign \new_[11239]_  = ~\new_[13905]_  & ~\new_[19085]_ ;
  assign \new_[11240]_  = ~\new_[13876]_  | ~\new_[16238]_ ;
  assign \new_[11241]_  = ~\new_[16283]_  | ~\new_[14211]_ ;
  assign \new_[11242]_  = ~\new_[12373]_ ;
  assign \new_[11243]_  = ~\new_[14314]_  | ~\new_[18709]_ ;
  assign \new_[11244]_  = ~\new_[18859]_  & ~\new_[14336]_ ;
  assign \new_[11245]_  = ~\new_[14617]_  | ~\new_[15112]_ ;
  assign \new_[11246]_  = \new_[13725]_  & \new_[15714]_ ;
  assign \new_[11247]_  = ~\new_[18042]_  | ~\new_[16394]_ ;
  assign \new_[11248]_  = ~\new_[12378]_ ;
  assign \new_[11249]_  = ~\new_[21076]_  | ~\new_[13753]_ ;
  assign \new_[11250]_  = ~\new_[13682]_  | ~\new_[14588]_ ;
  assign \new_[11251]_  = ~\new_[14873]_  | ~\new_[13943]_ ;
  assign \new_[11252]_  = ~\new_[12383]_ ;
  assign \new_[11253]_  = ~\new_[19711]_  & ~\new_[16180]_ ;
  assign \new_[11254]_  = ~\new_[14161]_  | ~\new_[13785]_ ;
  assign \new_[11255]_  = ~\new_[13702]_  | ~\new_[19381]_ ;
  assign \new_[11256]_  = ~\new_[12387]_ ;
  assign \new_[11257]_  = ~\new_[13818]_  | ~\new_[14296]_ ;
  assign \new_[11258]_  = ~\new_[13887]_  & ~\new_[15940]_ ;
  assign \new_[11259]_  = ~\new_[14741]_  | ~\new_[13579]_ ;
  assign \new_[11260]_  = \new_[14861]_  & \new_[13547]_ ;
  assign \new_[11261]_  = ~\new_[18278]_  | ~\new_[13664]_ ;
  assign \new_[11262]_  = ~\new_[14435]_  | ~\new_[15367]_ ;
  assign \new_[11263]_  = ~\new_[13706]_  | ~\new_[21391]_ ;
  assign \new_[11264]_  = ~\new_[14136]_  & ~\new_[18692]_ ;
  assign \new_[11265]_  = ~\new_[14359]_  & ~\new_[19681]_ ;
  assign \new_[11266]_  = ~\new_[16616]_  | ~\new_[19474]_ ;
  assign \new_[11267]_  = \new_[13876]_  | \new_[19024]_ ;
  assign \new_[11268]_  = \new_[15661]_  & \new_[13635]_ ;
  assign \new_[11269]_  = ~\new_[12396]_ ;
  assign \new_[11270]_  = ~\new_[14049]_  | ~\new_[13716]_ ;
  assign \new_[11271]_  = ~\new_[14547]_  | ~\new_[16235]_ ;
  assign \new_[11272]_  = ~\new_[21635]_  | ~\new_[14040]_ ;
  assign \new_[11273]_  = ~\new_[15037]_  | ~\new_[14591]_ ;
  assign \new_[11274]_  = ~\new_[12398]_ ;
  assign \new_[11275]_  = ~\new_[13539]_  | ~\new_[14268]_ ;
  assign \new_[11276]_  = ~\new_[14266]_  | ~\new_[15440]_ ;
  assign \new_[11277]_  = ~\new_[15202]_  | ~\new_[21562]_ ;
  assign \new_[11278]_  = \new_[13926]_  & \new_[19592]_ ;
  assign \new_[11279]_  = ~\new_[14182]_  | ~\new_[15328]_ ;
  assign \new_[11280]_  = ~\new_[13706]_  | ~\new_[16880]_ ;
  assign \new_[11281]_  = ~\new_[13991]_  | ~\new_[18621]_ ;
  assign \new_[11282]_  = ~\new_[12400]_ ;
  assign \new_[11283]_  = ~\new_[13590]_  | ~\new_[15282]_ ;
  assign \new_[11284]_  = ~\new_[15142]_  | ~\new_[13959]_ ;
  assign \new_[11285]_  = ~\new_[12401]_ ;
  assign \new_[11286]_  = ~\new_[13848]_  | ~\new_[14378]_ ;
  assign \new_[11287]_  = \new_[14210]_  | \new_[21629]_ ;
  assign \new_[11288]_  = ~\new_[19299]_  & ~\new_[13694]_ ;
  assign \new_[11289]_  = ~\new_[14260]_  & ~\new_[15179]_ ;
  assign \new_[11290]_  = \new_[13908]_  & \new_[17090]_ ;
  assign \new_[11291]_  = \new_[13908]_  & \new_[13669]_ ;
  assign \new_[11292]_  = ~\new_[12404]_ ;
  assign \new_[11293]_  = ~\new_[18246]_  & ~\new_[14121]_ ;
  assign \new_[11294]_  = ~\new_[15189]_  | ~\new_[14443]_ ;
  assign \new_[11295]_  = ~\new_[14050]_  & ~\new_[18832]_ ;
  assign \new_[11296]_  = ~\new_[21638]_  & (~\new_[17117]_  | ~\new_[14807]_ );
  assign \new_[11297]_  = ~\new_[13488]_  & (~\new_[18501]_  | ~\new_[18308]_ );
  assign \new_[11298]_  = ~\new_[13889]_  | ~\new_[20906]_ ;
  assign \new_[11299]_  = ~\new_[16837]_  | ~\new_[13579]_ ;
  assign \new_[11300]_  = ~\new_[14031]_  | ~\new_[19758]_ ;
  assign \new_[11301]_  = ~\new_[14306]_  & ~\new_[14282]_ ;
  assign \new_[11302]_  = ~\new_[12409]_ ;
  assign \new_[11303]_  = \new_[13819]_  & \new_[13821]_ ;
  assign \new_[11304]_  = ~\new_[14011]_  & ~\new_[13534]_ ;
  assign \new_[11305]_  = ~\new_[13520]_  & ~\new_[13811]_ ;
  assign \new_[11306]_  = ~\new_[19202]_  & (~\new_[15680]_  | ~\new_[17267]_ );
  assign \new_[11307]_  = ~\new_[12414]_ ;
  assign \new_[11308]_  = ~\new_[12412]_ ;
  assign \new_[11309]_  = ~\new_[13520]_  | ~\new_[18474]_ ;
  assign \new_[11310]_  = ~\new_[13409]_ ;
  assign \new_[11311]_  = ~\new_[14679]_  | ~\new_[18873]_ ;
  assign \new_[11312]_  = ~\new_[15029]_  | ~\new_[14310]_ ;
  assign \new_[11313]_  = ~\new_[14235]_  & ~\new_[13666]_ ;
  assign \new_[11314]_  = ~\new_[13768]_  | ~\new_[19136]_ ;
  assign \new_[11315]_  = ~\new_[15306]_  | ~\new_[20906]_ ;
  assign \new_[11316]_  = ~\new_[14251]_  | ~\new_[13530]_ ;
  assign \new_[11317]_  = ~\new_[14810]_  | ~\new_[14240]_ ;
  assign \new_[11318]_  = ~\new_[16678]_  | ~\new_[14005]_ ;
  assign \new_[11319]_  = ~\new_[13120]_ ;
  assign \new_[11320]_  = ~\new_[13889]_  & ~\new_[17457]_ ;
  assign \new_[11321]_  = ~\new_[15335]_  | ~\new_[13501]_ ;
  assign \new_[11322]_  = ~\new_[16499]_  | ~\new_[14264]_ ;
  assign \new_[11323]_  = ~\new_[13914]_  | ~\new_[18847]_ ;
  assign \new_[11324]_  = ~\new_[20906]_  | ~\new_[13868]_ ;
  assign \new_[11325]_  = ~\new_[12420]_ ;
  assign \new_[11326]_  = ~\new_[19553]_  & (~\new_[16319]_  | ~\new_[17316]_ );
  assign \new_[11327]_  = ~\new_[13854]_  | ~\new_[13530]_ ;
  assign \new_[11328]_  = ~\new_[13856]_  | ~\new_[16763]_ ;
  assign \new_[11329]_  = ~\new_[14060]_  | ~\new_[15454]_ ;
  assign \new_[11330]_  = ~\new_[19088]_  & ~\new_[14369]_ ;
  assign \new_[11331]_  = ~\new_[17056]_  | ~\new_[14062]_ ;
  assign \new_[11332]_  = \new_[15201]_  & \new_[13719]_ ;
  assign \new_[11333]_  = ~\new_[13772]_  & ~\new_[13815]_ ;
  assign \new_[11334]_  = \new_[13950]_  | \new_[19636]_ ;
  assign \new_[11335]_  = ~\new_[14642]_  | ~\new_[13816]_ ;
  assign \new_[11336]_  = \new_[19991]_  | \new_[14844]_ ;
  assign \new_[11337]_  = ~\new_[21714]_  | ~\new_[13989]_ ;
  assign \new_[11338]_  = ~\new_[21316]_  | ~\new_[13959]_ ;
  assign \new_[11339]_  = ~\new_[13953]_  & ~\new_[14951]_ ;
  assign \new_[11340]_  = \new_[13968]_  | \new_[18965]_ ;
  assign \new_[11341]_  = ~\new_[13874]_  | ~\new_[13872]_ ;
  assign \new_[11342]_  = ~\new_[13263]_ ;
  assign \new_[11343]_  = ~\new_[14870]_  & ~\new_[14172]_ ;
  assign \new_[11344]_  = ~\new_[13830]_  | ~\new_[19153]_ ;
  assign \new_[11345]_  = ~\new_[16159]_  | ~\new_[14421]_  | ~\new_[17576]_ ;
  assign \new_[11346]_  = ~\new_[12432]_ ;
  assign \new_[11347]_  = ~\new_[13688]_  | ~\new_[14206]_ ;
  assign \new_[11348]_  = \new_[14086]_  | \new_[19553]_ ;
  assign \new_[11349]_  = ~\new_[15736]_  | ~\new_[13849]_ ;
  assign \new_[11350]_  = ~\new_[14508]_  | ~\new_[14937]_ ;
  assign \new_[11351]_  = ~\new_[14287]_  & ~\new_[18083]_ ;
  assign \new_[11352]_  = ~\new_[17863]_  | ~\new_[14104]_ ;
  assign \new_[11353]_  = ~\new_[14101]_  | ~\new_[19084]_ ;
  assign \new_[11354]_  = ~\new_[13969]_  | ~\new_[16055]_ ;
  assign \new_[11355]_  = ~\new_[12439]_ ;
  assign \new_[11356]_  = ~\new_[12440]_ ;
  assign \new_[11357]_  = ~\new_[16478]_  | ~\new_[13622]_ ;
  assign \new_[11358]_  = ~\new_[15541]_  | ~\new_[13973]_ ;
  assign \new_[11359]_  = ~\new_[14002]_  & ~\new_[19474]_ ;
  assign \new_[11360]_  = ~\new_[13610]_  | ~\new_[13986]_ ;
  assign \new_[11361]_  = ~\new_[13261]_ ;
  assign \new_[11362]_  = ~\new_[13923]_  | ~\new_[14244]_ ;
  assign \new_[11363]_  = ~\new_[14321]_  | ~\new_[19249]_ ;
  assign \new_[11364]_  = ~\new_[15370]_  | ~\new_[21694]_ ;
  assign \new_[11365]_  = ~\new_[13846]_  | ~\new_[14152]_ ;
  assign \new_[11366]_  = ~\new_[13914]_  | ~\new_[18605]_ ;
  assign \new_[11367]_  = ~\new_[14572]_  | ~\new_[14387]_ ;
  assign \new_[11368]_  = ~\new_[13732]_  | ~\new_[15952]_ ;
  assign \new_[11369]_  = \new_[13688]_  | \new_[19217]_ ;
  assign \new_[11370]_  = ~\new_[15137]_  | ~\new_[13688]_ ;
  assign \new_[11371]_  = ~\new_[14430]_  & ~\new_[19217]_ ;
  assign \new_[11372]_  = ~\new_[12443]_ ;
  assign \new_[11373]_  = ~\new_[12444]_ ;
  assign \new_[11374]_  = ~\new_[14534]_  | ~\new_[20938]_ ;
  assign \new_[11375]_  = ~\new_[20222]_  | ~\new_[19428]_ ;
  assign \new_[11376]_  = ~\new_[14321]_  & (~\new_[16621]_  | ~\new_[18652]_ );
  assign \new_[11377]_  = ~\new_[12469]_ ;
  assign \new_[11378]_  = ~\new_[21507]_  & ~\new_[13854]_ ;
  assign \new_[11379]_  = ~\new_[14262]_  | (~\new_[18707]_  & ~\new_[19513]_ );
  assign \new_[11380]_  = ~\new_[13941]_  | ~\new_[15224]_ ;
  assign \new_[11381]_  = ~\new_[21043]_  | ~\new_[19409]_ ;
  assign \new_[11382]_  = ~\new_[15236]_  & ~\new_[15252]_ ;
  assign \new_[11383]_  = ~\new_[16665]_  & ~\new_[19050]_ ;
  assign \new_[11384]_  = ~\new_[14240]_  & ~\new_[18017]_ ;
  assign \new_[11385]_  = ~\new_[15001]_  | ~\new_[13750]_ ;
  assign \new_[11386]_  = ~\new_[15500]_  | ~\new_[14106]_ ;
  assign \new_[11387]_  = ~\new_[12447]_ ;
  assign \new_[11388]_  = ~\new_[14209]_  | ~\new_[19374]_ ;
  assign \new_[11389]_  = ~\new_[13962]_  | ~\new_[13893]_ ;
  assign \new_[11390]_  = ~\new_[15565]_  | ~\new_[16333]_  | ~\new_[16420]_ ;
  assign \new_[11391]_  = ~\new_[16974]_  | ~\new_[16591]_  | ~\new_[17188]_ ;
  assign \new_[11392]_  = ~\new_[15539]_  | ~\new_[16257]_  | ~\new_[16557]_ ;
  assign \new_[11393]_  = \new_[14324]_  | \new_[14433]_ ;
  assign \new_[11394]_  = \new_[13631]_  | \new_[14446]_ ;
  assign \new_[11395]_  = ~\new_[14203]_  & (~\new_[18543]_  | ~\new_[17155]_ );
  assign \new_[11396]_  = ~\new_[18836]_  & (~\new_[15688]_  | ~\new_[17242]_ );
  assign \new_[11397]_  = ~\new_[14156]_  & (~\new_[17761]_  | ~\new_[18011]_ );
  assign \new_[11398]_  = ~\new_[14415]_  & (~\new_[16628]_  | ~\new_[18601]_ );
  assign \new_[11399]_  = ~\new_[13637]_  | ~\new_[14297]_ ;
  assign \new_[11400]_  = ~\new_[14449]_  | (~\new_[14836]_  & ~\new_[19612]_ );
  assign \new_[11401]_  = ~\new_[14252]_  | (~\new_[15471]_  & ~\new_[19261]_ );
  assign \new_[11402]_  = ~\new_[15304]_  | ~\new_[13715]_ ;
  assign \new_[11403]_  = ~\new_[15474]_  | ~\new_[16055]_ ;
  assign \new_[11404]_  = ~\new_[13508]_  | ~\new_[14183]_ ;
  assign \new_[11405]_  = ~\new_[19088]_  & (~\new_[16654]_  | ~\new_[14757]_ );
  assign \new_[11406]_  = ~\new_[15900]_  & (~\new_[17451]_  | ~\new_[18935]_ );
  assign \new_[11407]_  = ~\new_[17927]_  & (~\new_[15646]_  | ~\new_[17576]_ );
  assign \new_[11408]_  = ~\new_[18033]_  & (~\new_[15686]_  | ~\new_[18486]_ );
  assign \new_[11409]_  = ~\new_[19592]_  & (~\new_[17216]_  | ~\new_[14840]_ );
  assign \new_[11410]_  = ~\new_[14539]_  | ~\new_[13695]_ ;
  assign \new_[11411]_  = ~\new_[15588]_  | ~\new_[14015]_ ;
  assign \new_[11412]_  = \new_[15835]_  | \new_[13883]_ ;
  assign \new_[11413]_  = ~\new_[14224]_  | ~\new_[13817]_ ;
  assign \new_[11414]_  = ~\new_[14573]_  | ~\new_[16180]_ ;
  assign \new_[11415]_  = ~\new_[14302]_  | ~\new_[14430]_ ;
  assign \new_[11416]_  = ~\new_[14046]_  | ~\new_[13905]_ ;
  assign \new_[11417]_  = ~\new_[14671]_  | ~\new_[14078]_ ;
  assign \new_[11418]_  = ~\new_[19094]_  & (~\new_[15834]_  | ~\new_[15608]_ );
  assign \new_[11419]_  = ~\new_[19006]_  & (~\new_[15132]_  | ~\new_[14865]_ );
  assign \new_[11420]_  = ~\new_[19711]_  & (~\new_[15799]_  | ~\new_[15560]_ );
  assign \new_[11421]_  = ~\new_[14255]_  & ~\new_[13864]_ ;
  assign \new_[11422]_  = ~\new_[16444]_  | ~\new_[13705]_ ;
  assign \new_[11423]_  = ~\new_[13581]_  | ~\new_[14180]_ ;
  assign \new_[11424]_  = ~\new_[14577]_  | ~\new_[13636]_ ;
  assign \new_[11425]_  = ~\new_[18416]_  & (~\new_[17246]_  | ~\new_[15505]_ );
  assign \new_[11426]_  = ~\new_[14249]_  | ~\new_[13938]_ ;
  assign \new_[11427]_  = ~\new_[14144]_  | ~\new_[14257]_ ;
  assign \new_[11428]_  = ~\new_[18846]_  & (~\new_[18349]_  | ~\new_[17646]_ );
  assign \new_[11429]_  = ~\new_[16997]_  & (~\new_[19248]_  | ~\new_[17690]_ );
  assign \new_[11430]_  = ~\new_[13903]_  & ~\new_[14236]_ ;
  assign \new_[11431]_  = ~\new_[13760]_  & (~\new_[16020]_  | ~\new_[19202]_ );
  assign \new_[11432]_  = ~\new_[13966]_  & (~\new_[15955]_  | ~\new_[18209]_ );
  assign \new_[11433]_  = ~\new_[14300]_  & (~\new_[15867]_  | ~\new_[21495]_ );
  assign \new_[11434]_  = ~\new_[16142]_  | ~\new_[14115]_ ;
  assign \new_[11435]_  = ~\new_[13807]_  & ~\new_[14372]_ ;
  assign \new_[11436]_  = ~\new_[13809]_  & ~\new_[13592]_ ;
  assign \new_[11437]_  = ~\new_[14845]_  & (~\new_[16794]_  | ~\new_[18414]_ );
  assign \new_[11438]_  = ~\new_[13865]_  & ~\new_[14055]_ ;
  assign \new_[11439]_  = ~\new_[13907]_  & ~\new_[14357]_ ;
  assign \new_[11440]_  = ~\new_[13254]_ ;
  assign \new_[11441]_  = ~\new_[13930]_  & ~\new_[14154]_ ;
  assign \new_[11442]_  = ~\new_[13933]_  | ~\new_[15204]_ ;
  assign \new_[11443]_  = ~\new_[15190]_  & (~\new_[15595]_  | ~\new_[18414]_ );
  assign \new_[11444]_  = ~\new_[15271]_  & (~\new_[14889]_  | ~\new_[19409]_ );
  assign \new_[11445]_  = ~\new_[13940]_  | ~\new_[14088]_ ;
  assign \new_[11446]_  = ~\new_[13944]_  & ~\new_[14124]_ ;
  assign \new_[11447]_  = ~\new_[13761]_  & ~\new_[14237]_ ;
  assign \new_[11448]_  = ~\new_[14625]_  | ~\new_[16143]_ ;
  assign \new_[11449]_  = ~\new_[14528]_  | ~\new_[13802]_ ;
  assign \new_[11450]_  = ~\new_[15742]_  | ~\new_[13726]_ ;
  assign \new_[11451]_  = \new_[14151]_  & \new_[15892]_ ;
  assign \new_[11452]_  = \new_[14794]_  | \new_[14390]_ ;
  assign \new_[11453]_  = ~\new_[17594]_  | (~\new_[17033]_  & ~\new_[16584]_ );
  assign \new_[11454]_  = ~\new_[15747]_  | ~\new_[13709]_ ;
  assign \new_[11455]_  = ~\new_[17734]_  | ~\new_[14501]_ ;
  assign \new_[11456]_  = \new_[14402]_  & \new_[18262]_ ;
  assign \new_[11457]_  = ~\new_[13253]_ ;
  assign \new_[11458]_  = ~\new_[14621]_  | ~\new_[13714]_ ;
  assign \new_[11459]_  = ~\new_[18906]_  | ~\new_[14276]_  | ~\new_[18750]_ ;
  assign \new_[11460]_  = ~\new_[15424]_  | ~\new_[13755]_ ;
  assign \new_[11461]_  = ~\new_[14403]_  | ~\new_[17382]_ ;
  assign \new_[11462]_  = ~\new_[18826]_  | (~\new_[17677]_  & ~\new_[16584]_ );
  assign \new_[11463]_  = ~\new_[14394]_  | ~\new_[18201]_ ;
  assign \new_[11464]_  = ~\new_[18403]_  | (~\new_[16622]_  & ~\new_[14827]_ );
  assign \new_[11465]_  = ~\new_[14405]_  | ~\new_[15792]_ ;
  assign \new_[11466]_  = ~\new_[14277]_  & (~\new_[19228]_  | ~\new_[17017]_ );
  assign \new_[11467]_  = ~\new_[14114]_  | (~\new_[18846]_  & ~\new_[16003]_ );
  assign \new_[11468]_  = ~\new_[14552]_  | ~\new_[13743]_ ;
  assign \new_[11469]_  = ~\new_[13847]_  | (~\new_[18913]_  & ~\new_[18665]_ );
  assign \new_[11470]_  = ~\new_[14303]_  | (~\new_[15832]_  & ~\new_[16997]_ );
  assign \new_[11471]_  = ~\new_[20966]_  | (~\new_[16062]_  & ~\new_[15999]_ );
  assign \new_[11472]_  = ~\new_[14036]_  | (~\new_[14730]_  & ~\new_[18123]_ );
  assign \new_[11473]_  = ~\new_[16364]_  | ~\new_[13878]_ ;
  assign \new_[11474]_  = ~\new_[14551]_  | ~\new_[20904]_ ;
  assign \new_[11475]_  = ~\new_[18304]_  | (~\new_[17405]_  & ~\new_[16472]_ );
  assign \new_[11476]_  = \new_[14472]_  & \new_[16246]_ ;
  assign \new_[11477]_  = \new_[16360]_  & \new_[14171]_ ;
  assign \new_[11478]_  = \new_[16463]_  & \new_[14286]_ ;
  assign \new_[11479]_  = \new_[16060]_  & \new_[14097]_ ;
  assign \new_[11480]_  = \new_[16677]_  & \new_[14673]_ ;
  assign \new_[11481]_  = \new_[14530]_  & \new_[16561]_ ;
  assign \new_[11482]_  = \new_[15670]_  & \new_[14216]_ ;
  assign \new_[11483]_  = \new_[16429]_  & \new_[14250]_ ;
  assign \new_[11484]_  = \new_[15733]_  & \new_[13499]_ ;
  assign \new_[11485]_  = \new_[14614]_  & \new_[16978]_ ;
  assign \new_[11486]_  = \new_[18453]_  ^ \new_[15774]_ ;
  assign \new_[11487]_  = \new_[18737]_  ^ \new_[14930]_ ;
  assign \new_[11488]_  = \new_[18830]_  ^ \new_[15766]_ ;
  assign \new_[11489]_  = ~\new_[14656]_  | ~\new_[17381]_ ;
  assign \new_[11490]_  = ~\new_[13640]_  | ~\new_[14835]_ ;
  assign \new_[11491]_  = ~\new_[12496]_ ;
  assign \new_[11492]_  = ~\new_[12497]_ ;
  assign \new_[11493]_  = ~\new_[13473]_ ;
  assign \new_[11494]_  = ~\new_[12501]_ ;
  assign \new_[11495]_  = ~\new_[14618]_  | ~\new_[18973]_ ;
  assign \new_[11496]_  = ~\new_[12505]_ ;
  assign \new_[11497]_  = ~\new_[16058]_  | ~\new_[18228]_ ;
  assign \new_[11498]_  = \new_[13529]_  & \new_[19018]_ ;
  assign \new_[11499]_  = ~\new_[15907]_  | ~\new_[18567]_  | ~\new_[18984]_  | ~\new_[19386]_ ;
  assign \new_[11500]_  = ~\new_[12516]_ ;
  assign \new_[11501]_  = ~\new_[15907]_  | ~\new_[17476]_  | ~\new_[19107]_  | ~\new_[18567]_ ;
  assign \new_[11502]_  = ~\new_[13634]_  & ~\new_[19097]_ ;
  assign \new_[11503]_  = ~\new_[13451]_ ;
  assign \new_[11504]_  = ~\new_[14489]_  | ~\new_[19028]_ ;
  assign \new_[11505]_  = ~\new_[14570]_  | ~\new_[17381]_ ;
  assign \new_[11506]_  = ~\new_[18575]_  & ~\new_[14652]_ ;
  assign \new_[11507]_  = ~\new_[14685]_  | ~\new_[18337]_ ;
  assign \new_[11508]_  = ~\new_[12524]_ ;
  assign \new_[11509]_  = \new_[14637]_  | \new_[18859]_ ;
  assign \new_[11510]_  = ~\new_[14233]_  | ~\new_[19538]_ ;
  assign \new_[11511]_  = ~\new_[14675]_  & ~\new_[19265]_ ;
  assign \new_[11512]_  = ~\new_[12536]_ ;
  assign \new_[11513]_  = ~\new_[12542]_ ;
  assign \new_[11514]_  = ~\new_[12543]_ ;
  assign \new_[11515]_  = ~\new_[12546]_ ;
  assign \new_[11516]_  = ~\new_[12549]_ ;
  assign \new_[11517]_  = \new_[14488]_  & \new_[19253]_ ;
  assign \new_[11518]_  = ~\new_[12554]_ ;
  assign \new_[11519]_  = \new_[16145]_  | \new_[18443]_ ;
  assign \new_[11520]_  = ~\new_[12559]_ ;
  assign \new_[11521]_  = \new_[14500]_  | \new_[21513]_ ;
  assign \new_[11522]_  = ~\new_[20969]_ ;
  assign \new_[11523]_  = ~\new_[12564]_ ;
  assign \new_[11524]_  = ~\new_[13355]_ ;
  assign \new_[11525]_  = ~\new_[14620]_  | ~\new_[18443]_ ;
  assign \new_[11526]_  = ~\new_[12568]_ ;
  assign \new_[11527]_  = ~\new_[13678]_  | ~\new_[18821]_ ;
  assign \new_[11528]_  = ~\new_[12570]_ ;
  assign \new_[11529]_  = ~\new_[13780]_ ;
  assign \new_[11530]_  = \new_[14509]_  | \new_[19269]_ ;
  assign \new_[11531]_  = \new_[14561]_  & \new_[21496]_ ;
  assign \new_[11532]_  = ~\new_[12572]_ ;
  assign \new_[11533]_  = ~\new_[13550]_  | ~\new_[18984]_ ;
  assign \new_[11534]_  = ~\new_[13651]_  | ~\new_[19050]_ ;
  assign \new_[11535]_  = ~\new_[13791]_ ;
  assign \new_[11536]_  = ~\new_[12580]_ ;
  assign \new_[11537]_  = ~\new_[12583]_ ;
  assign \new_[11538]_  = \new_[15962]_  & \new_[19036]_ ;
  assign \new_[11539]_  = ~\new_[14474]_  | ~\new_[19084]_ ;
  assign \new_[11540]_  = ~\new_[14516]_  & ~\new_[19269]_ ;
  assign \new_[11541]_  = ~\new_[12584]_ ;
  assign \new_[11542]_  = ~\new_[12586]_ ;
  assign \new_[11543]_  = ~\new_[12594]_ ;
  assign \new_[11544]_  = ~\new_[12597]_ ;
  assign \new_[11545]_  = ~\new_[12598]_ ;
  assign \new_[11546]_  = ~\new_[13555]_  | ~\new_[19102]_ ;
  assign \new_[11547]_  = ~\new_[12600]_ ;
  assign \new_[11548]_  = ~\new_[12602]_ ;
  assign \new_[11549]_  = ~\new_[14461]_  | ~\new_[18008]_ ;
  assign \new_[11550]_  = ~\new_[13567]_  | ~\new_[18427]_ ;
  assign \new_[11551]_  = ~\new_[20899]_ ;
  assign \new_[11552]_  = \new_[14477]_  & \new_[19754]_ ;
  assign \new_[11553]_  = ~\new_[14514]_  | ~\new_[21115]_ ;
  assign \new_[11554]_  = ~\new_[14433]_  | ~\new_[18228]_ ;
  assign \new_[11555]_  = ~\new_[12607]_ ;
  assign \new_[11556]_  = ~\new_[14688]_  | ~\new_[19208]_ ;
  assign \new_[11557]_  = ~\new_[12608]_ ;
  assign \new_[11558]_  = ~\new_[12613]_ ;
  assign \new_[11559]_  = ~\new_[14600]_  | ~\new_[19224]_ ;
  assign \new_[11560]_  = ~\new_[12614]_ ;
  assign \new_[11561]_  = ~\new_[12617]_ ;
  assign \new_[11562]_  = ~\new_[20434]_ ;
  assign \new_[11563]_  = ~\new_[12618]_ ;
  assign \new_[11564]_  = ~\new_[12619]_ ;
  assign \new_[11565]_  = ~\new_[12620]_ ;
  assign \new_[11566]_  = ~\new_[12621]_ ;
  assign \new_[11567]_  = ~\new_[12622]_ ;
  assign \new_[11568]_  = ~\new_[12623]_ ;
  assign \new_[11569]_  = ~\new_[12626]_ ;
  assign \new_[11570]_  = ~\new_[13368]_ ;
  assign \new_[11571]_  = ~\new_[12630]_ ;
  assign \new_[11572]_  = ~\new_[21094]_ ;
  assign \new_[11573]_  = ~\new_[21703]_  | ~\new_[19154]_ ;
  assign \new_[11574]_  = \new_[12488]_ ;
  assign \new_[11575]_  = ~\new_[14490]_  | ~\new_[19088]_ ;
  assign \new_[11576]_  = ~\new_[12643]_ ;
  assign \new_[11577]_  = \new_[14638]_  & \new_[18898]_ ;
  assign \new_[11578]_  = ~\new_[14446]_  | ~\new_[18605]_ ;
  assign \new_[11579]_  = ~\new_[14538]_  | ~\new_[19436]_ ;
  assign \new_[11580]_  = ~\new_[12647]_ ;
  assign \new_[11581]_  = ~\new_[13506]_  | ~\new_[18678]_ ;
  assign \new_[11582]_  = ~\new_[12650]_ ;
  assign \new_[11583]_  = ~\new_[14140]_  | ~\new_[18692]_ ;
  assign \new_[11584]_  = ~\new_[12654]_ ;
  assign \new_[11585]_  = ~\new_[12655]_ ;
  assign \new_[11586]_  = ~\new_[12445]_ ;
  assign \new_[11587]_  = ~\new_[12651]_ ;
  assign \new_[11588]_  = \new_[13523]_  & \new_[18285]_ ;
  assign \new_[11589]_  = ~\new_[12657]_ ;
  assign \new_[11590]_  = \new_[14582]_  | \new_[21328]_ ;
  assign \new_[11591]_  = ~\new_[12427]_ ;
  assign \new_[11592]_  = ~\new_[12659]_ ;
  assign \new_[11593]_  = ~\new_[12429]_ ;
  assign \new_[11594]_  = ~\new_[12660]_ ;
  assign \new_[11595]_  = ~\new_[12662]_ ;
  assign \new_[11596]_  = ~\new_[12664]_ ;
  assign \new_[11597]_  = ~\new_[14686]_  | ~\new_[18840]_ ;
  assign \new_[11598]_  = ~\new_[12667]_ ;
  assign \new_[11599]_  = ~\new_[12393]_ ;
  assign \new_[11600]_  = ~\new_[15970]_  | ~\new_[19729]_ ;
  assign \new_[11601]_  = ~\new_[14467]_  | ~\new_[17273]_ ;
  assign \new_[11602]_  = ~\new_[14594]_  | ~\new_[19217]_ ;
  assign \new_[11603]_  = ~\new_[12670]_ ;
  assign \new_[11604]_  = ~\new_[14442]_  | ~\new_[18682]_ ;
  assign \new_[11605]_  = ~\new_[12362]_ ;
  assign \new_[11606]_  = ~\new_[12671]_ ;
  assign \new_[11607]_  = ~\new_[12673]_ ;
  assign \new_[11608]_  = ~\new_[12674]_ ;
  assign \new_[11609]_  = ~\new_[12675]_ ;
  assign \new_[11610]_  = ~\new_[12676]_ ;
  assign \new_[11611]_  = \new_[14613]_  & \new_[18969]_ ;
  assign \new_[11612]_  = ~\new_[12677]_ ;
  assign \new_[11613]_  = ~\new_[21392]_  | ~\new_[19462]_ ;
  assign \new_[11614]_  = \new_[14611]_  & \new_[19476]_ ;
  assign \new_[11615]_  = ~\new_[14520]_  | ~\new_[18709]_ ;
  assign \new_[11616]_  = ~\new_[12684]_ ;
  assign \new_[11617]_  = ~\new_[14566]_  | ~\new_[21511]_ ;
  assign \new_[11618]_  = ~\new_[12685]_ ;
  assign \new_[11619]_  = ~\new_[12687]_ ;
  assign \new_[11620]_  = ~\new_[12690]_ ;
  assign \new_[11621]_  = ~\new_[12691]_ ;
  assign \new_[11622]_  = \new_[14475]_  & \new_[19266]_ ;
  assign \new_[11623]_  = ~\new_[14510]_  | ~\new_[19107]_ ;
  assign \new_[11624]_  = ~\new_[12244]_ ;
  assign \new_[11625]_  = ~\new_[12258]_ ;
  assign \new_[11626]_  = ~\new_[18501]_  & ~\new_[13488]_ ;
  assign \new_[11627]_  = ~\new_[21408]_ ;
  assign \new_[11628]_  = ~\new_[12696]_ ;
  assign \new_[11629]_  = ~\new_[13869]_  | ~\new_[17457]_ ;
  assign \new_[11630]_  = ~\new_[12700]_ ;
  assign \new_[11631]_  = ~\new_[14522]_  | ~\new_[20680]_ ;
  assign \new_[11632]_  = ~\new_[12234]_ ;
  assign \new_[11633]_  = ~\new_[12235]_ ;
  assign \new_[11634]_  = ~\new_[12702]_ ;
  assign \new_[11635]_  = ~\new_[12704]_ ;
  assign \new_[11636]_  = ~\new_[12706]_ ;
  assign \new_[11637]_  = ~\new_[14384]_  | ~\new_[17944]_ ;
  assign \new_[11638]_  = \new_[17201]_  ^ \new_[19513]_ ;
  assign \new_[11639]_  = ~\new_[13514]_  | ~\new_[18166]_ ;
  assign \new_[11640]_  = \new_[14535]_  & \new_[19269]_ ;
  assign \new_[11641]_  = ~\new_[21569]_  & ~\new_[14435]_ ;
  assign \new_[11642]_  = ~\new_[12710]_ ;
  assign \new_[11643]_  = ~\new_[12714]_ ;
  assign \new_[11644]_  = ~\new_[12166]_ ;
  assign \new_[11645]_  = ~\new_[12158]_ ;
  assign \new_[11646]_  = ~\new_[14576]_  | ~\new_[19202]_ ;
  assign \new_[11647]_  = ~\new_[14475]_  | ~\new_[17598]_ ;
  assign \new_[11648]_  = ~\new_[16273]_  | ~\new_[19018]_ ;
  assign \new_[11649]_  = ~\new_[12721]_ ;
  assign \new_[11650]_  = ~\new_[12722]_ ;
  assign \new_[11651]_  = ~\new_[12729]_ ;
  assign \new_[11652]_  = ~\new_[14602]_  | ~\new_[17979]_ ;
  assign \new_[11653]_  = ~\new_[12726]_ ;
  assign \new_[11654]_  = ~\new_[12727]_ ;
  assign \new_[11655]_  = ~\new_[14574]_  | ~\new_[18077]_ ;
  assign \new_[11656]_  = ~\new_[12730]_ ;
  assign \new_[11657]_  = ~\new_[12731]_ ;
  assign \new_[11658]_  = ~\new_[14578]_  | ~\new_[18077]_ ;
  assign \new_[11659]_  = ~\new_[12738]_ ;
  assign \new_[11660]_  = ~\new_[12740]_ ;
  assign \new_[11661]_  = ~\new_[12742]_ ;
  assign \new_[11662]_  = \new_[13588]_  & \new_[18008]_ ;
  assign \new_[11663]_  = ~\new_[12744]_ ;
  assign \new_[11664]_  = \new_[14610]_  & \new_[18605]_ ;
  assign \new_[11665]_  = ~\new_[12747]_ ;
  assign \new_[11666]_  = ~\new_[12748]_ ;
  assign \new_[11667]_  = \new_[13548]_  & \new_[19409]_ ;
  assign \new_[11668]_  = ~\new_[12749]_ ;
  assign \new_[11669]_  = ~\new_[12750]_ ;
  assign \new_[11670]_  = ~\new_[12753]_ ;
  assign \new_[11671]_  = ~\new_[12755]_ ;
  assign \new_[11672]_  = ~\new_[14537]_  | ~\new_[19462]_ ;
  assign \new_[11673]_  = \new_[18335]_  | \new_[13488]_ ;
  assign \new_[11674]_  = ~\new_[14691]_  & ~\new_[19554]_ ;
  assign \new_[11675]_  = ~\new_[12759]_ ;
  assign \new_[11676]_  = ~\new_[14482]_  | ~\new_[18652]_ ;
  assign \new_[11677]_  = ~\new_[12765]_ ;
  assign \new_[11678]_  = ~\new_[12766]_ ;
  assign \new_[11679]_  = ~\new_[12767]_ ;
  assign \new_[11680]_  = ~\new_[14536]_  | ~\new_[14837]_ ;
  assign \new_[11681]_  = ~\new_[14456]_  | ~\new_[18166]_ ;
  assign \new_[11682]_  = ~\new_[12771]_ ;
  assign \new_[11683]_  = ~\new_[12146]_ ;
  assign \new_[11684]_  = ~\new_[12772]_ ;
  assign \new_[11685]_  = ~\new_[14678]_  | ~\new_[21689]_ ;
  assign \new_[11686]_  = ~\new_[12775]_ ;
  assign \new_[11687]_  = \new_[16084]_  | \new_[17457]_ ;
  assign \new_[11688]_  = ~\new_[12776]_ ;
  assign \new_[11689]_  = ~\new_[18046]_  & ~\new_[15620]_ ;
  assign \new_[11690]_  = ~\new_[15926]_  | ~\new_[19008]_ ;
  assign \new_[11691]_  = \new_[16416]_  | \new_[17979]_ ;
  assign \new_[11692]_  = ~\new_[12779]_ ;
  assign \new_[11693]_  = ~\new_[14513]_  | ~\new_[17598]_ ;
  assign \new_[11694]_  = ~\new_[16590]_  & ~\new_[18209]_ ;
  assign \new_[11695]_  = ~\new_[14574]_  | ~\new_[17457]_ ;
  assign \new_[11696]_  = ~\new_[12783]_ ;
  assign \new_[11697]_  = ~\new_[12784]_ ;
  assign \new_[11698]_  = ~\new_[14543]_  | ~\new_[19269]_ ;
  assign \new_[11699]_  = \new_[14660]_  & \new_[19084]_ ;
  assign \new_[11700]_  = \new_[15899]_  | \new_[19290]_ ;
  assign \new_[11701]_  = ~\new_[14442]_  | ~\new_[19202]_ ;
  assign \new_[11702]_  = \new_[13538]_  | \new_[18285]_ ;
  assign \new_[11703]_  = ~\new_[12786]_ ;
  assign \new_[11704]_  = ~\new_[12788]_ ;
  assign \new_[11705]_  = ~\new_[12788]_ ;
  assign \new_[11706]_  = ~\new_[13468]_ ;
  assign \new_[11707]_  = ~\new_[12789]_ ;
  assign \new_[11708]_  = ~\new_[13462]_ ;
  assign \new_[11709]_  = ~\new_[12790]_ ;
  assign \new_[11710]_  = ~\new_[12791]_ ;
  assign \new_[11711]_  = ~\new_[14323]_  | ~\new_[21572]_ ;
  assign \new_[11712]_  = \new_[13977]_ ;
  assign \new_[11713]_  = ~\new_[13545]_  | ~\new_[18692]_ ;
  assign \new_[11714]_  = ~\new_[12798]_ ;
  assign \new_[11715]_  = ~\new_[14470]_  | ~\new_[21697]_ ;
  assign \new_[11716]_  = ~\new_[13600]_  | ~\new_[18605]_ ;
  assign \new_[11717]_  = ~\new_[14642]_ ;
  assign \new_[11718]_  = ~\new_[12802]_ ;
  assign \new_[11719]_  = ~\new_[12803]_ ;
  assign \new_[11720]_  = ~\new_[14595]_  | ~\new_[18111]_ ;
  assign \new_[11721]_  = ~\new_[12805]_ ;
  assign \new_[11722]_  = ~\new_[12807]_ ;
  assign \new_[11723]_  = ~\new_[14491]_  & ~\new_[17979]_ ;
  assign \new_[11724]_  = ~\new_[12816]_ ;
  assign \new_[11725]_  = ~\new_[12817]_ ;
  assign \new_[11726]_  = ~\new_[12822]_ ;
  assign \new_[11727]_  = ~\new_[12824]_ ;
  assign \new_[11728]_  = ~\new_[12825]_ ;
  assign \new_[11729]_  = ~\new_[14438]_  | ~\new_[18643]_ ;
  assign \new_[11730]_  = ~\new_[18044]_  | ~\new_[16394]_ ;
  assign \new_[11731]_  = ~\new_[12828]_ ;
  assign \new_[11732]_  = ~\new_[12830]_ ;
  assign \new_[11733]_  = ~\new_[14556]_  & ~\new_[19474]_ ;
  assign \new_[11734]_  = ~\new_[12831]_ ;
  assign \new_[11735]_  = ~\new_[18385]_  | ~\new_[16058]_ ;
  assign \new_[11736]_  = ~\new_[12834]_ ;
  assign \new_[11737]_  = \new_[14064]_  | \new_[14826]_ ;
  assign \new_[11738]_  = ~\new_[16560]_  | ~\new_[18008]_ ;
  assign \new_[11739]_  = ~\new_[13942]_  | ~\new_[17457]_ ;
  assign \new_[11740]_  = ~\new_[12839]_ ;
  assign \new_[11741]_  = ~\new_[16466]_  | ~\new_[18124]_ ;
  assign \new_[11742]_  = ~\new_[16349]_  & ~\new_[19275]_ ;
  assign \new_[11743]_  = ~\new_[14433]_  | ~\new_[17522]_ ;
  assign \new_[11744]_  = ~\new_[12841]_ ;
  assign \new_[11745]_  = ~\new_[17583]_  & ~\new_[20664]_ ;
  assign \new_[11746]_  = ~\new_[12845]_ ;
  assign \new_[11747]_  = ~\new_[13359]_ ;
  assign \new_[11748]_  = ~\new_[16832]_  | ~\new_[13567]_ ;
  assign \new_[11749]_  = ~\new_[12851]_ ;
  assign \new_[11750]_  = ~\new_[14493]_  & ~\new_[18228]_ ;
  assign \new_[11751]_  = ~\new_[12852]_ ;
  assign \new_[11752]_  = ~\new_[12854]_ ;
  assign \new_[11753]_  = ~\new_[17274]_  | ~\new_[16394]_ ;
  assign \new_[11754]_  = ~\new_[17667]_  | ~\new_[14543]_ ;
  assign \new_[11755]_  = ~\new_[14460]_  & ~\new_[18166]_ ;
  assign \new_[11756]_  = ~\new_[12861]_ ;
  assign \new_[11757]_  = ~\new_[13250]_ ;
  assign \new_[11758]_  = ~\new_[13213]_ ;
  assign \new_[11759]_  = ~\new_[19098]_  | ~\new_[14896]_  | ~\new_[18304]_ ;
  assign \new_[11760]_  = ~\new_[17664]_  | ~\new_[16058]_ ;
  assign \new_[11761]_  = ~\new_[17287]_  | ~\new_[16416]_ ;
  assign \new_[11762]_  = ~\new_[16432]_  | ~\new_[19151]_ ;
  assign \new_[11763]_  = ~\new_[16402]_  | ~\new_[19013]_ ;
  assign \new_[11764]_  = ~\new_[12872]_ ;
  assign \new_[11765]_  = ~\new_[14288]_  | ~\new_[14825]_ ;
  assign \new_[11766]_  = ~\new_[18728]_  | ~\new_[13869]_ ;
  assign \new_[11767]_  = ~\new_[12877]_ ;
  assign \new_[11768]_  = ~\new_[13649]_  & ~\new_[18153]_ ;
  assign \new_[11769]_  = ~\new_[13061]_ ;
  assign \new_[11770]_  = ~\new_[12880]_ ;
  assign \new_[11771]_  = ~\new_[16416]_  & ~\new_[19169]_ ;
  assign \new_[11772]_  = ~\new_[12882]_ ;
  assign \new_[11773]_  = ~\new_[12883]_ ;
  assign \new_[11774]_  = ~\new_[15720]_  & ~\new_[14546]_ ;
  assign \new_[11775]_  = ~\new_[14479]_  & ~\new_[18166]_ ;
  assign \new_[11776]_  = ~\new_[18815]_  & ~\new_[13712]_ ;
  assign \new_[11777]_  = ~\new_[14674]_  | ~\new_[18984]_ ;
  assign \new_[11778]_  = \new_[14465]_  | \new_[15765]_ ;
  assign \new_[11779]_  = ~\new_[12887]_ ;
  assign \new_[11780]_  = ~\new_[13565]_  | ~\new_[18678]_ ;
  assign \new_[11781]_  = \new_[16293]_  | \new_[16286]_ ;
  assign \new_[11782]_  = ~\new_[12891]_ ;
  assign \new_[11783]_  = ~\new_[12892]_ ;
  assign \new_[11784]_  = ~\new_[14428]_  & ~\new_[17598]_ ;
  assign \new_[11785]_  = \new_[17840]_  & \new_[14665]_ ;
  assign \new_[11786]_  = ~\new_[13594]_  | ~\new_[14881]_ ;
  assign \new_[11787]_  = \new_[14503]_  | \new_[19073]_ ;
  assign \new_[11788]_  = ~\new_[12900]_ ;
  assign \new_[11789]_  = ~\new_[16187]_  & ~\new_[19107]_ ;
  assign \new_[11790]_  = ~\new_[12901]_ ;
  assign \new_[11791]_  = ~\new_[12905]_ ;
  assign \new_[11792]_  = ~\new_[16579]_  | ~\new_[19064]_ ;
  assign \new_[11793]_  = ~\new_[16524]_  | ~\new_[19711]_ ;
  assign \new_[11794]_  = \new_[14585]_  | \new_[18734]_ ;
  assign \new_[11795]_  = ~\new_[17710]_  | ~\new_[13514]_ ;
  assign \new_[11796]_  = ~\new_[14136]_  | ~\new_[17236]_ ;
  assign \new_[11797]_  = \new_[13712]_  | \new_[21562]_ ;
  assign \new_[11798]_  = ~\new_[21671]_  | ~\new_[18840]_ ;
  assign \new_[11799]_  = ~\new_[12917]_ ;
  assign \new_[11800]_  = ~\new_[12919]_ ;
  assign \new_[11801]_  = ~\new_[17359]_  | ~\new_[16058]_ ;
  assign \new_[11802]_  = ~\new_[17594]_  | ~\new_[21606]_ ;
  assign \new_[11803]_  = ~\new_[12928]_ ;
  assign \new_[11804]_  = ~\new_[17191]_  & ~\new_[17385]_ ;
  assign \new_[11805]_  = ~\new_[18328]_  | ~\new_[13658]_ ;
  assign \new_[11806]_  = ~\new_[16324]_  | ~\new_[19269]_ ;
  assign \new_[11807]_  = \new_[14428]_  | \new_[19450]_ ;
  assign \new_[11808]_  = ~\new_[12936]_ ;
  assign \new_[11809]_  = ~\new_[14439]_  | ~\new_[18972]_ ;
  assign \new_[11810]_  = \new_[14485]_  | \new_[19115]_ ;
  assign \new_[11811]_  = ~\new_[13486]_  | ~\new_[18888]_ ;
  assign \new_[11812]_  = \new_[16160]_  | \new_[18821]_ ;
  assign \new_[11813]_  = ~\new_[14583]_  & ~\new_[19275]_ ;
  assign \new_[11814]_  = ~\new_[16860]_  | ~\new_[16394]_ ;
  assign \new_[11815]_  = ~\new_[12947]_ ;
  assign \new_[11816]_  = ~\new_[17903]_  | ~\new_[16394]_ ;
  assign \new_[11817]_  = ~\new_[14667]_  | ~\new_[19450]_ ;
  assign \new_[11818]_  = \new_[17468]_  & \new_[15209]_ ;
  assign \new_[11819]_  = ~\new_[12951]_ ;
  assign \new_[11820]_  = ~\new_[21138]_ ;
  assign \new_[11821]_  = ~\new_[14446]_  | ~\new_[17818]_ ;
  assign \new_[11822]_  = ~\new_[18635]_  | ~\new_[13658]_ ;
  assign \new_[11823]_  = ~\new_[17166]_  & ~\new_[14520]_ ;
  assign \new_[11824]_  = ~\new_[12957]_ ;
  assign \new_[11825]_  = ~\new_[17559]_  | ~\new_[15209]_ ;
  assign \new_[11826]_  = ~\new_[21130]_ ;
  assign \new_[11827]_  = ~\new_[12959]_ ;
  assign \new_[11828]_  = ~\new_[12312]_ ;
  assign \new_[11829]_  = \new_[14644]_  | \new_[19587]_ ;
  assign \new_[11830]_  = ~\new_[12968]_ ;
  assign \new_[11831]_  = ~\new_[12969]_ ;
  assign \new_[11832]_  = ~\new_[13632]_  & ~\new_[14951]_ ;
  assign \new_[11833]_  = \new_[19141]_  | \new_[16296]_ ;
  assign \new_[11834]_  = ~\new_[17900]_  | ~\new_[16394]_ ;
  assign \new_[11835]_  = ~\new_[12973]_ ;
  assign \new_[11836]_  = ~\new_[16335]_  | ~\new_[21689]_ ;
  assign \new_[11837]_  = ~\new_[12977]_ ;
  assign \new_[11838]_  = ~\new_[16732]_  | ~\new_[16394]_ ;
  assign \new_[11839]_  = ~\new_[12980]_ ;
  assign \new_[11840]_  = ~\new_[13076]_ ;
  assign \new_[11841]_  = ~\new_[12981]_ ;
  assign \new_[11842]_  = ~\new_[16236]_  | ~\new_[19095]_ ;
  assign \new_[11843]_  = ~\new_[12987]_ ;
  assign \new_[11844]_  = ~\new_[17653]_  | ~\new_[16394]_ ;
  assign \new_[11845]_  = ~\new_[12991]_ ;
  assign \new_[11846]_  = ~\new_[17658]_  & ~\new_[14544]_ ;
  assign \new_[11847]_  = ~\new_[12992]_ ;
  assign \new_[11848]_  = ~\new_[17461]_  | ~\new_[14442]_ ;
  assign \new_[11849]_  = ~\new_[21606]_  | ~\new_[18811]_ ;
  assign \new_[11850]_  = ~\new_[16870]_  & ~\new_[14602]_ ;
  assign \new_[11851]_  = \new_[17917]_  & \new_[13658]_ ;
  assign \new_[11852]_  = ~\new_[16590]_  & ~\new_[18537]_ ;
  assign \new_[11853]_  = ~\new_[17917]_  | ~\new_[15879]_ ;
  assign \new_[11854]_  = ~\new_[13002]_ ;
  assign \new_[11855]_  = ~\new_[16361]_  | ~\new_[18077]_ ;
  assign \new_[11856]_  = ~\new_[14492]_  | ~\new_[15644]_ ;
  assign \new_[11857]_  = ~\new_[18037]_  | ~\new_[14566]_ ;
  assign \new_[11858]_  = ~\new_[13007]_ ;
  assign \new_[11859]_  = ~\new_[18502]_  | ~\new_[16394]_ ;
  assign \new_[11860]_  = ~\new_[16234]_  | ~\new_[16879]_ ;
  assign \new_[11861]_  = ~\new_[14599]_  | ~\new_[18994]_ ;
  assign \new_[11862]_  = ~\new_[13025]_ ;
  assign \new_[11863]_  = ~\new_[21398]_  | ~\new_[21502]_ ;
  assign \new_[11864]_  = \new_[18923]_  | \new_[13492]_ ;
  assign \new_[11865]_  = ~\new_[14549]_  & ~\new_[19319]_ ;
  assign \new_[11866]_  = ~\new_[17954]_  | ~\new_[14620]_ ;
  assign \new_[11867]_  = ~\new_[16073]_  | ~\new_[19204]_ ;
  assign \new_[11868]_  = ~\new_[15442]_  | ~\new_[13605]_ ;
  assign \new_[11869]_  = ~\new_[13031]_ ;
  assign \new_[11870]_  = ~\new_[13036]_ ;
  assign \new_[11871]_  = ~\new_[13402]_ ;
  assign \new_[11872]_  = ~\new_[13038]_ ;
  assign \new_[11873]_  = ~\new_[13395]_ ;
  assign \new_[11874]_  = ~\new_[16271]_  | ~\new_[21638]_ ;
  assign \new_[11875]_  = ~\new_[13047]_ ;
  assign \new_[11876]_  = ~\new_[13364]_ ;
  assign \new_[11877]_  = ~\new_[13205]_ ;
  assign \new_[11878]_  = ~\new_[13051]_ ;
  assign \new_[11879]_  = ~\new_[16354]_  | ~\new_[18031]_ ;
  assign \new_[11880]_  = ~\new_[13053]_ ;
  assign \new_[11881]_  = ~\new_[13054]_ ;
  assign \new_[11882]_  = ~\new_[14587]_  | ~\new_[14757]_ ;
  assign \new_[11883]_  = ~\new_[14198]_ ;
  assign \new_[11884]_  = ~\new_[15504]_  | ~\new_[14507]_ ;
  assign \new_[11885]_  = ~\new_[17991]_  | ~\new_[13567]_ ;
  assign \new_[11886]_  = ~\new_[14606]_  & ~\new_[21635]_ ;
  assign \new_[11887]_  = ~\new_[13065]_ ;
  assign \new_[11888]_  = ~\new_[13632]_  & ~\new_[18228]_ ;
  assign \new_[11889]_  = ~\new_[14509]_  & ~\new_[18875]_ ;
  assign \new_[11890]_  = ~\new_[14533]_  & ~\new_[18938]_ ;
  assign \new_[11891]_  = ~\new_[13121]_ ;
  assign \new_[11892]_  = ~\new_[15874]_  | ~\new_[21689]_ ;
  assign \new_[11893]_  = ~\new_[17909]_  | ~\new_[14611]_ ;
  assign \new_[11894]_  = ~\new_[16580]_  | ~\new_[18325]_ ;
  assign \new_[11895]_  = ~\new_[13064]_ ;
  assign \new_[11896]_  = \new_[17742]_  | \new_[15885]_ ;
  assign \new_[11897]_  = ~\new_[21606]_  | ~\new_[19082]_ ;
  assign \new_[11898]_  = ~\new_[13570]_  & ~\new_[15704]_ ;
  assign \new_[11899]_  = ~\new_[17933]_  | ~\new_[14500]_ ;
  assign \new_[11900]_  = ~\new_[13075]_ ;
  assign \new_[11901]_  = ~\new_[12956]_ ;
  assign \new_[11902]_  = \new_[18923]_  | \new_[13504]_ ;
  assign \new_[11903]_  = ~\new_[14597]_  | ~\new_[19214]_ ;
  assign \new_[11904]_  = ~\new_[16023]_  | ~\new_[18747]_ ;
  assign \new_[11905]_  = ~\new_[16146]_  & ~\new_[19214]_ ;
  assign \new_[11906]_  = ~\new_[15278]_ ;
  assign \new_[11907]_  = \new_[14285]_  | \new_[18062]_ ;
  assign \new_[11908]_  = ~\new_[19550]_  & (~\new_[15249]_  | ~\new_[14915]_ );
  assign \new_[11909]_  = \new_[16626]_  | \new_[19161]_ ;
  assign \new_[11910]_  = ~\new_[13449]_ ;
  assign \new_[11911]_  = \new_[13088]_ ;
  assign \new_[11912]_  = ~\new_[14683]_  & ~\new_[18559]_ ;
  assign \new_[11913]_  = ~\new_[16588]_  | ~\new_[19247]_ ;
  assign \new_[11914]_  = \new_[18066]_  | \new_[16185]_ ;
  assign \new_[11915]_  = ~\new_[15915]_  | ~\new_[19196]_ ;
  assign \new_[11916]_  = ~\new_[14469]_  | ~\new_[15694]_ ;
  assign \new_[11917]_  = ~\new_[14210]_  & ~\new_[18126]_ ;
  assign \new_[11918]_  = \new_[14581]_  | \new_[15924]_ ;
  assign \new_[11919]_  = ~\new_[13099]_ ;
  assign \new_[11920]_  = ~\new_[16523]_  & ~\new_[21056]_ ;
  assign \new_[11921]_  = ~\new_[16032]_  & ~\new_[19244]_ ;
  assign \new_[11922]_  = ~\new_[16567]_  | ~\new_[19006]_ ;
  assign \new_[11923]_  = ~\new_[17367]_  | ~\new_[14442]_ ;
  assign \new_[11924]_  = ~\new_[12495]_ ;
  assign \new_[11925]_  = ~\new_[16115]_  | ~\new_[19476]_ ;
  assign \new_[11926]_  = ~\new_[17730]_  | ~\new_[21606]_ ;
  assign \new_[11927]_  = ~\new_[13106]_ ;
  assign \new_[11928]_  = ~\new_[14456]_  | ~\new_[18644]_ ;
  assign \new_[11929]_  = ~\new_[18322]_  | ~\new_[16119]_ ;
  assign \new_[11930]_  = \new_[16145]_  & \new_[14693]_ ;
  assign \new_[11931]_  = ~\new_[12465]_ ;
  assign \new_[11932]_  = ~\new_[13113]_ ;
  assign \new_[11933]_  = ~\new_[13118]_ ;
  assign \new_[11934]_  = \new_[19027]_  | \new_[14469]_ ;
  assign \new_[11935]_  = ~\new_[12424]_ ;
  assign \new_[11936]_  = ~\new_[13281]_ ;
  assign \new_[11937]_  = \new_[14628]_  | \new_[19269]_ ;
  assign \new_[11938]_  = ~\new_[13122]_ ;
  assign \new_[11939]_  = ~\new_[12395]_ ;
  assign \new_[11940]_  = ~\new_[12389]_ ;
  assign \new_[11941]_  = ~\new_[12363]_ ;
  assign \new_[11942]_  = \new_[14623]_  | \new_[21507]_ ;
  assign \new_[11943]_  = ~\new_[17730]_  | ~\new_[16119]_ ;
  assign \new_[11944]_  = ~\new_[17468]_  | ~\new_[15890]_ ;
  assign \new_[11945]_  = ~\new_[13132]_ ;
  assign \new_[11946]_  = ~\new_[14665]_  | ~\new_[19625]_ ;
  assign \new_[11947]_  = \new_[18106]_  | \new_[14288]_ ;
  assign \new_[11948]_  = ~\new_[13137]_ ;
  assign \new_[11949]_  = ~\new_[13142]_ ;
  assign \new_[11950]_  = ~\new_[13147]_ ;
  assign \new_[11951]_  = ~\new_[13148]_ ;
  assign \new_[11952]_  = ~\new_[13152]_ ;
  assign \new_[11953]_  = ~\new_[15978]_  | ~\new_[21557]_ ;
  assign \new_[11954]_  = ~\new_[12171]_ ;
  assign \new_[11955]_  = ~\new_[13154]_ ;
  assign \new_[11956]_  = ~\new_[13154]_ ;
  assign \new_[11957]_  = ~\new_[16153]_  | ~\new_[19018]_ ;
  assign \new_[11958]_  = ~\new_[17840]_  | ~\new_[16391]_ ;
  assign \new_[11959]_  = ~\new_[14586]_  | ~\new_[17887]_ ;
  assign \new_[11960]_  = ~\new_[13504]_  | ~\new_[14837]_ ;
  assign \new_[11961]_  = ~\new_[17082]_  | ~\new_[13545]_ ;
  assign \new_[11962]_  = ~\new_[17898]_  | ~\new_[16394]_ ;
  assign \new_[11963]_  = ~\new_[13170]_ ;
  assign \new_[11964]_  = \new_[20215]_  | \new_[19171]_ ;
  assign \new_[11965]_  = ~\new_[20661]_  | ~\new_[14678]_ ;
  assign \new_[11966]_  = ~\new_[18157]_  | ~\new_[13778]_ ;
  assign \new_[11967]_  = \new_[16270]_  | \new_[19141]_ ;
  assign \new_[11968]_  = \new_[15881]_  | \new_[19681]_ ;
  assign \new_[11969]_  = \new_[14459]_  | \new_[19018]_ ;
  assign \new_[11970]_  = \new_[13551]_  & \new_[17180]_ ;
  assign \new_[11971]_  = ~\new_[15936]_  | ~\new_[19021]_ ;
  assign \new_[11972]_  = ~\new_[14564]_  | ~\new_[19018]_ ;
  assign \new_[11973]_  = ~\new_[17132]_  & ~\new_[13605]_ ;
  assign \new_[11974]_  = ~\new_[14468]_  & ~\new_[18605]_ ;
  assign \new_[11975]_  = \new_[14460]_  | \new_[19612]_ ;
  assign \new_[11976]_  = ~\new_[13386]_ ;
  assign \new_[11977]_  = \new_[21388]_  | \new_[20215]_ ;
  assign \new_[11978]_  = ~\new_[13190]_ ;
  assign \new_[11979]_  = ~\new_[13346]_ ;
  assign \new_[11980]_  = ~\new_[13260]_ ;
  assign \new_[11981]_  = ~\new_[13197]_ ;
  assign \new_[11982]_  = ~\new_[14464]_  | ~\new_[21638]_ ;
  assign \new_[11983]_  = ~\new_[14498]_  | ~\new_[21693]_ ;
  assign \new_[11984]_  = ~\new_[14318]_  | ~\new_[21500]_ ;
  assign \new_[11985]_  = \new_[16452]_  | \new_[18926]_ ;
  assign \new_[11986]_  = ~\new_[14444]_  | ~\new_[17845]_ ;
  assign \new_[11987]_  = ~\new_[16570]_  | ~\new_[19687]_ ;
  assign \new_[11988]_  = ~\new_[12949]_ ;
  assign \new_[11989]_  = ~\new_[12950]_ ;
  assign \new_[11990]_  = ~\new_[12922]_ ;
  assign \new_[11991]_  = ~\new_[13215]_ ;
  assign \new_[11992]_  = ~\new_[13218]_ ;
  assign \new_[11993]_  = ~\new_[13222]_ ;
  assign \new_[11994]_  = ~\new_[13221]_ ;
  assign \new_[11995]_  = ~\new_[13223]_ ;
  assign \new_[11996]_  = ~\new_[16010]_  | ~\new_[18637]_ ;
  assign \new_[11997]_  = ~\new_[15406]_  | ~\new_[14454]_ ;
  assign \new_[11998]_  = ~\new_[12743]_ ;
  assign \new_[11999]_  = ~\new_[13230]_ ;
  assign \new_[12000]_  = \new_[16476]_  & \new_[16704]_ ;
  assign \new_[12001]_  = ~\new_[17551]_  | ~\new_[14594]_ ;
  assign \new_[12002]_  = \new_[13498]_  & \new_[14876]_ ;
  assign \new_[12003]_  = ~\new_[21606]_  | ~\new_[19587]_ ;
  assign \new_[12004]_  = ~\new_[18286]_  | ~\new_[16394]_ ;
  assign \new_[12005]_  = ~\new_[16070]_  | ~\new_[18572]_ ;
  assign \new_[12006]_  = ~\new_[13242]_ ;
  assign \new_[12007]_  = ~\new_[18270]_  | ~\new_[14513]_ ;
  assign \new_[12008]_  = ~\new_[12489]_ ;
  assign \new_[12009]_  = ~\new_[21548]_  | ~\new_[19050]_ ;
  assign \new_[12010]_  = ~\new_[15324]_  & (~\new_[14903]_  | ~\new_[19153]_ );
  assign \new_[12011]_  = ~\new_[13251]_ ;
  assign \new_[12012]_  = ~\new_[13252]_ ;
  assign \new_[12013]_  = ~\new_[14558]_  | ~\new_[18427]_ ;
  assign \new_[12014]_  = ~\new_[13257]_ ;
  assign \new_[12015]_  = ~\new_[18167]_  | ~\new_[14520]_ ;
  assign \new_[12016]_  = ~\new_[16832]_  | ~\new_[14685]_ ;
  assign \new_[12017]_  = \new_[15940]_  | \new_[14462]_ ;
  assign \new_[12018]_  = ~\new_[13271]_ ;
  assign \new_[12019]_  = ~\new_[18002]_  & ~\new_[14587]_ ;
  assign \new_[12020]_  = ~\new_[16185]_  & ~\new_[17979]_ ;
  assign \new_[12021]_  = ~\new_[19222]_  | ~\new_[14140]_ ;
  assign \new_[12022]_  = ~\new_[13274]_ ;
  assign \new_[12023]_  = \new_[15994]_  | \new_[14453]_ ;
  assign \new_[12024]_  = ~\new_[17759]_  | ~\new_[16394]_ ;
  assign \new_[12025]_  = ~\new_[13287]_ ;
  assign \new_[12026]_  = ~\new_[18910]_  | ~\new_[14592]_ ;
  assign \new_[12027]_  = ~\new_[12291]_ ;
  assign \new_[12028]_  = ~\new_[21652]_  | ~\new_[21306]_ ;
  assign \new_[12029]_  = ~\new_[14311]_  | ~\new_[18228]_ ;
  assign \new_[12030]_  = ~\new_[13297]_ ;
  assign \new_[12031]_  = ~\new_[21300]_  & ~\new_[18358]_ ;
  assign \new_[12032]_  = ~\new_[14496]_  | ~\new_[19462]_ ;
  assign \new_[12033]_  = ~\new_[18401]_  | ~\new_[13518]_ ;
  assign \new_[12034]_  = ~\new_[14654]_  | ~\new_[15778]_ ;
  assign \new_[12035]_  = ~\new_[13658]_  | ~\new_[19261]_ ;
  assign \new_[12036]_  = ~\new_[16290]_  | ~\new_[16185]_ ;
  assign \new_[12037]_  = ~\new_[12163]_ ;
  assign \new_[12038]_  = ~\new_[19260]_  | ~\new_[14595]_ ;
  assign \new_[12039]_  = ~\new_[15879]_  | ~\new_[17845]_ ;
  assign \new_[12040]_  = ~\new_[20164]_  | ~\new_[18873]_ ;
  assign \new_[12041]_  = ~\new_[16391]_  | ~\new_[17522]_ ;
  assign \new_[12042]_  = ~\new_[12155]_ ;
  assign \new_[12043]_  = ~\new_[16057]_  | ~\new_[16840]_ ;
  assign \new_[12044]_  = ~\new_[13317]_ ;
  assign \new_[12045]_  = \new_[14473]_  | \new_[16387]_ ;
  assign \new_[12046]_  = \new_[14557]_  | \new_[14506]_ ;
  assign \new_[12047]_  = \new_[17913]_  | \new_[14628]_ ;
  assign \new_[12048]_  = ~\new_[16700]_  & (~\new_[17354]_  | ~\new_[17485]_ );
  assign \new_[12049]_  = ~\new_[14655]_  | ~\new_[13556]_ ;
  assign \new_[12050]_  = ~\new_[17648]_  & (~\new_[14789]_  | ~\new_[18014]_ );
  assign \new_[12051]_  = ~\new_[16084]_  | (~\new_[17658]_  & ~\new_[18861]_ );
  assign \new_[12052]_  = ~\new_[14518]_  | ~\new_[13538]_ ;
  assign \new_[12053]_  = ~\new_[14589]_  | ~\new_[14643]_ ;
  assign \new_[12054]_  = ~\new_[17699]_  & (~\new_[14934]_  | ~\new_[15894]_ );
  assign \new_[12055]_  = ~\new_[17364]_  | ~\new_[13551]_ ;
  assign \new_[12056]_  = ~\new_[18920]_  | ~\new_[14632]_ ;
  assign \new_[12057]_  = \new_[14450]_  | \new_[18180]_ ;
  assign \new_[12058]_  = ~\new_[18048]_  & ~\new_[14459]_ ;
  assign \new_[12059]_  = ~\new_[17882]_  & (~\new_[17946]_  | ~\new_[15636]_ );
  assign \new_[12060]_  = ~\new_[14541]_  | (~\new_[16655]_  & ~\new_[18111]_ );
  assign \new_[12061]_  = ~\new_[14550]_  | (~\new_[17384]_  & ~\new_[21505]_ );
  assign \new_[12062]_  = ~\new_[14494]_  | ~\new_[17339]_ ;
  assign \new_[12063]_  = ~\new_[14540]_  & (~\new_[18577]_  | ~\new_[17528]_ );
  assign \new_[12064]_  = ~\new_[14427]_  & (~\new_[17529]_  | ~\new_[18814]_ );
  assign \new_[12065]_  = ~\new_[14575]_  & (~\new_[18575]_  | ~\new_[18365]_ );
  assign \new_[12066]_  = ~\new_[14682]_  & (~\new_[20490]_  | ~\new_[21533]_ );
  assign \new_[12067]_  = ~\new_[13541]_  & (~\new_[20699]_  | ~\new_[18782]_ );
  assign \new_[12068]_  = ~\new_[14429]_  & (~\new_[19444]_  | ~\new_[19389]_ );
  assign \new_[12069]_  = ~\new_[13626]_  & (~\new_[19386]_  | ~\new_[16740]_ );
  assign \new_[12070]_  = ~\new_[14612]_  & (~\new_[19379]_  | ~\new_[18779]_ );
  assign \new_[12071]_  = ~\new_[14568]_  & (~\new_[21572]_  | ~\new_[18717]_ );
  assign \new_[12072]_  = ~\new_[13568]_  | ~\new_[19426]_ ;
  assign \new_[12073]_  = ~\new_[13358]_ ;
  assign \new_[12074]_  = ~\new_[12202]_ ;
  assign \new_[12075]_  = ~\new_[20663]_ ;
  assign \new_[12076]_  = ~\new_[13374]_ ;
  assign \new_[12077]_  = ~\new_[19156]_  | ~\new_[19098]_  | ~\new_[17553]_ ;
  assign \new_[12078]_  = ~\new_[12757]_ ;
  assign \new_[12079]_  = ~\new_[21603]_ ;
  assign \new_[12080]_  = ~\new_[13389]_ ;
  assign \new_[12081]_  = ~\new_[13393]_ ;
  assign \new_[12082]_  = ~\new_[19203]_  | ~\new_[17578]_  | ~\new_[18025]_ ;
  assign n2723 = ~\new_[19363]_  & (~\new_[14972]_  | ~\new_[14785]_ );
  assign \new_[12084]_  = ~\new_[17156]_  | ~\new_[18715]_  | ~\new_[14787]_ ;
  assign \new_[12085]_  = ~\new_[12150]_ ;
  assign \new_[12086]_  = ~\new_[13411]_ ;
  assign \new_[12087]_  = ~\new_[17239]_  | ~\new_[14865]_ ;
  assign \new_[12088]_  = ~\new_[13591]_  | ~\new_[18115]_ ;
  assign \new_[12089]_  = ~\new_[17974]_  | ~\new_[21392]_ ;
  assign \new_[12090]_  = ~\new_[12177]_ ;
  assign \new_[12091]_  = ~\new_[13483]_ ;
  assign \new_[12092]_  = \new_[18246]_  | \new_[14663]_ ;
  assign \new_[12093]_  = ~\new_[13531]_  & ~\new_[21394]_ ;
  assign \new_[12094]_  = ~\new_[12537]_ ;
  assign \new_[12095]_  = ~\new_[13179]_ ;
  assign \new_[12096]_  = ~\new_[16600]_  & ~\new_[18523]_ ;
  assign \new_[12097]_  = ~\new_[18316]_  & ~\new_[14669]_ ;
  assign \new_[12098]_  = ~\new_[16467]_  | ~\new_[14582]_ ;
  assign \new_[12099]_  = ~\new_[13019]_ ;
  assign \new_[12100]_  = \new_[19673]_  ^ \new_[18906]_ ;
  assign \new_[12101]_  = ~\new_[14458]_  & ~\new_[18166]_ ;
  assign \new_[12102]_  = \new_[19626]_  ^ \new_[17578]_ ;
  assign \new_[12103]_  = \new_[15147]_  ^ \new_[18378]_ ;
  assign \new_[12104]_  = \new_[19810]_  ^ \new_[18998]_ ;
  assign \new_[12105]_  = ~\new_[19366]_  | (~\new_[15331]_  & ~\new_[16085]_ );
  assign \new_[12106]_  = \new_[14780]_  ^ \new_[19308]_ ;
  assign \new_[12107]_  = \new_[19716]_  ^ \new_[19603]_ ;
  assign \new_[12108]_  = \new_[15482]_  ^ \new_[18935]_ ;
  assign \new_[12109]_  = \new_[14700]_  ^ \new_[18772]_ ;
  assign \new_[12110]_  = \new_[17302]_  ^ \new_[16682]_ ;
  assign \new_[12111]_  = ~\new_[17574]_  | ~\new_[14436]_ ;
  assign \new_[12112]_  = \new_[17397]_  ^ \new_[17482]_ ;
  assign \new_[12113]_  = \new_[19720]_  ^ \new_[18179]_ ;
  assign \new_[12114]_  = \new_[15757]_  ^ \new_[19603]_ ;
  assign \new_[12115]_  = ~\new_[18965]_  & (~\new_[15294]_  | ~\new_[17062]_ );
  assign \new_[12116]_  = \new_[13603]_  | \new_[18187]_ ;
  assign \new_[12117]_  = \new_[16036]_  | \new_[19535]_  | \new_[19145]_  | \new_[18652]_ ;
  assign \new_[12118]_  = ~\new_[20341]_  & (~\new_[16487]_  | ~\new_[15328]_ );
  assign \new_[12119]_  = ~\new_[13549]_  | ~\new_[14387]_ ;
  assign \new_[12120]_  = ~\new_[14371]_  | ~\new_[14852]_ ;
  assign \new_[12121]_  = ~\new_[14444]_  | ~\new_[21688]_ ;
  assign \new_[12122]_  = ~\new_[13505]_  | ~\new_[16396]_ ;
  assign \new_[12123]_  = ~\new_[13470]_ ;
  assign \new_[12124]_  = ~\new_[19277]_  | (~\new_[15833]_  & ~\new_[14846]_ );
  assign \new_[12125]_  = \new_[13616]_  | \new_[18414]_ ;
  assign \new_[12126]_  = ~\new_[15342]_  | ~\new_[16177]_  | ~\new_[16775]_ ;
  assign \new_[12127]_  = ~\new_[14999]_  | ~\new_[14813]_  | ~\new_[15318]_ ;
  assign \new_[12128]_  = ~\new_[13619]_  | ~\new_[19377]_ ;
  assign \new_[12129]_  = ~\new_[13544]_  | ~\new_[17447]_ ;
  assign \new_[12130]_  = ~\new_[14079]_  | ~\new_[13566]_ ;
  assign \new_[12131]_  = \new_[13766]_  & \new_[14915]_ ;
  assign \new_[12132]_  = ~\new_[17445]_  | ~\new_[14267]_  | ~\new_[14995]_ ;
  assign \new_[12133]_  = ~\new_[19561]_  | (~\new_[15732]_  & ~\new_[16241]_ );
  assign \new_[12134]_  = \\dcnt_reg[0] ;
  assign \new_[12135]_  = ~\new_[20763]_  | (~\new_[15439]_  & ~\new_[15273]_ );
  assign \new_[12136]_  = ~\new_[14839]_  | ~\new_[13804]_  | ~\new_[14977]_ ;
  assign \new_[12137]_  = ~\new_[17266]_  | ~\new_[14121]_  | ~\new_[15374]_ ;
  assign \new_[12138]_  = \\u0_r0_rcnt_reg[3] ;
  assign \new_[12139]_  = ~\new_[13639]_  | ~\new_[19299]_ ;
  assign \new_[12140]_  = ~\new_[13526]_  | ~\new_[14875]_ ;
  assign \new_[12141]_  = ~\new_[14196]_  | ~\new_[13587]_ ;
  assign \new_[12142]_  = ~\new_[18077]_  & (~\new_[15387]_  | ~\new_[15716]_ );
  assign \new_[12143]_  = ~\new_[14626]_ ;
  assign \new_[12144]_  = ~\new_[15408]_  | ~\new_[15820]_ ;
  assign \new_[12145]_  = ~\new_[13484]_ ;
  assign \new_[12146]_  = ~\new_[19409]_  & ~\new_[14708]_ ;
  assign \new_[12147]_  = ~\new_[17487]_  | ~\new_[14955]_ ;
  assign \new_[12148]_  = ~\new_[20704]_  & (~\new_[16164]_  | ~\new_[16458]_ );
  assign \new_[12149]_  = ~\new_[17110]_  | ~\new_[14955]_ ;
  assign \new_[12150]_  = \new_[18826]_  & \new_[14783]_ ;
  assign \new_[12151]_  = \new_[16209]_  | \new_[15457]_ ;
  assign \new_[12152]_  = ~\new_[14796]_  | ~\new_[18979]_ ;
  assign \new_[12153]_  = ~\new_[13639]_ ;
  assign \new_[12154]_  = \new_[18644]_  & \new_[15666]_ ;
  assign \new_[12155]_  = ~\new_[14398]_ ;
  assign \new_[12156]_  = ~\new_[15280]_  | ~\new_[18678]_ ;
  assign \new_[12157]_  = ~\new_[17006]_  | ~\new_[15282]_ ;
  assign \new_[12158]_  = ~\new_[14847]_  | ~\new_[18166]_ ;
  assign \new_[12159]_  = ~\new_[14395]_ ;
  assign \new_[12160]_  = ~\new_[19727]_  & (~\new_[16222]_  | ~\new_[15949]_ );
  assign \new_[12161]_  = ~\new_[15715]_  | ~\new_[18627]_ ;
  assign \new_[12162]_  = ~\new_[18528]_  | (~\new_[16019]_  & ~\new_[16585]_ );
  assign \new_[12163]_  = \new_[15404]_  | \new_[21689]_ ;
  assign \new_[12164]_  = ~\new_[14117]_ ;
  assign \new_[12165]_  = ~\new_[14391]_ ;
  assign \new_[12166]_  = ~\new_[15396]_  & ~\new_[19446]_ ;
  assign \new_[12167]_  = ~\new_[14229]_ ;
  assign \new_[12168]_  = ~\new_[20907]_  | ~\new_[18616]_ ;
  assign \new_[12169]_  = ~\new_[17197]_  & ~\new_[21562]_ ;
  assign \new_[12170]_  = \new_[15123]_  | \new_[19107]_ ;
  assign \new_[12171]_  = ~\new_[17402]_  | ~\new_[15866]_ ;
  assign \new_[12172]_  = ~\new_[15575]_  | ~\new_[15608]_ ;
  assign \new_[12173]_  = ~\new_[15638]_  & ~\new_[18821]_ ;
  assign \new_[12174]_  = ~\new_[21495]_  | ~\new_[16879]_  | ~\new_[16288]_ ;
  assign \new_[12175]_  = ~\new_[16983]_  | ~\new_[21579]_  | ~\new_[21508]_  | ~\new_[20699]_ ;
  assign \new_[12176]_  = \new_[15243]_  | \new_[19239]_ ;
  assign \new_[12177]_  = ~\new_[13550]_ ;
  assign \new_[12178]_  = ~\new_[18533]_  | ~\new_[21521]_  | ~\new_[19130]_  | ~\new_[18035]_ ;
  assign \new_[12179]_  = ~\new_[13552]_ ;
  assign \new_[12180]_  = ~\new_[17425]_  | ~\new_[19035]_  | ~\new_[17886]_  | ~\new_[21056]_ ;
  assign \new_[12181]_  = \new_[14966]_  | \new_[19156]_ ;
  assign \new_[12182]_  = ~\new_[19454]_  | ~\new_[18008]_  | ~\new_[16007]_ ;
  assign \new_[12183]_  = ~\new_[16934]_  | ~\new_[18881]_  | ~\new_[18017]_  | ~\new_[18587]_ ;
  assign \new_[12184]_  = ~\new_[16877]_  | ~\new_[19123]_  | ~\new_[18209]_  | ~\new_[19675]_ ;
  assign \new_[12185]_  = ~\new_[15360]_  | ~\new_[18083]_ ;
  assign \new_[12186]_  = ~\new_[15049]_  & ~\new_[19288]_ ;
  assign \new_[12187]_  = ~\new_[16883]_  | ~\new_[18408]_  | ~\new_[19088]_  | ~\new_[18166]_ ;
  assign \new_[12188]_  = ~\new_[14995]_  & ~\new_[19319]_ ;
  assign \new_[12189]_  = ~\new_[13557]_ ;
  assign \new_[12190]_  = ~\new_[15353]_  | ~\new_[19553]_ ;
  assign \new_[12191]_  = \new_[15110]_  & \new_[19553]_ ;
  assign \new_[12192]_  = ~\new_[15225]_  & ~\new_[19553]_ ;
  assign \new_[12193]_  = ~\new_[16905]_  | ~\new_[19478]_  | ~\new_[18994]_  | ~\new_[19379]_ ;
  assign \new_[12194]_  = ~\new_[18972]_  & ~\new_[15048]_ ;
  assign \new_[12195]_  = ~\new_[15046]_  & ~\new_[18832]_ ;
  assign \new_[12196]_  = ~\new_[14271]_ ;
  assign \new_[12197]_  = ~\new_[13568]_ ;
  assign \new_[12198]_  = ~\new_[14842]_  & ~\new_[19008]_ ;
  assign \new_[12199]_  = ~\new_[20665]_  | ~\new_[21659]_  | ~\new_[19204]_  | ~\new_[18794]_ ;
  assign \new_[12200]_  = ~\new_[21136]_  & ~\new_[19021]_ ;
  assign \new_[12201]_  = ~\new_[14267]_  & ~\new_[19158]_ ;
  assign \new_[12202]_  = ~\new_[14447]_ ;
  assign \new_[12203]_  = ~\new_[15201]_  & ~\new_[19161]_ ;
  assign \new_[12204]_  = \new_[17391]_  | \new_[19035]_  | \new_[19941]_  | \new_[18083]_ ;
  assign \new_[12205]_  = ~\new_[15328]_  & ~\new_[19233]_ ;
  assign \new_[12206]_  = ~\new_[15148]_  | ~\new_[20865]_ ;
  assign \new_[12207]_  = \new_[15330]_  & \new_[19713]_ ;
  assign \new_[12208]_  = ~\new_[17422]_  | ~\new_[19123]_  | ~\new_[18209]_  | ~\new_[19675]_ ;
  assign \new_[12209]_  = \new_[15544]_  | \new_[19115]_ ;
  assign \new_[12210]_  = \new_[15002]_  | \new_[19409]_ ;
  assign \new_[12211]_  = \new_[15224]_  | \new_[18209]_ ;
  assign \new_[12212]_  = ~\new_[16851]_  | ~\new_[21520]_  | ~\new_[19064]_  | ~\new_[17529]_ ;
  assign \new_[12213]_  = ~\new_[15469]_  | ~\new_[18228]_ ;
  assign \new_[12214]_  = ~\new_[15009]_  | ~\new_[21498]_ ;
  assign \new_[12215]_  = \new_[17386]_  | \new_[18925]_  | \new_[19625]_  | \new_[19068]_ ;
  assign \new_[12216]_  = ~\new_[17746]_  | ~\new_[19319]_  | ~\new_[19335]_ ;
  assign \new_[12217]_  = ~\new_[17278]_  | ~\new_[18740]_  | ~\new_[19592]_  | ~\new_[17594]_ ;
  assign \new_[12218]_  = ~\new_[15121]_  | ~\new_[19288]_ ;
  assign \new_[12219]_  = ~\new_[15222]_  & ~\new_[18832]_ ;
  assign \new_[12220]_  = ~\new_[13571]_ ;
  assign \new_[12221]_  = ~\new_[15366]_  | ~\new_[18166]_ ;
  assign \new_[12222]_  = ~\new_[15003]_  & ~\new_[18972]_ ;
  assign \new_[12223]_  = \new_[14715]_  | \new_[19319]_ ;
  assign \new_[12224]_  = \new_[17564]_  | \new_[18026]_  | \new_[19592]_  | \new_[18811]_ ;
  assign \new_[12225]_  = ~\new_[15211]_  & ~\new_[18414]_ ;
  assign \new_[12226]_  = ~\new_[14993]_  & ~\new_[19158]_ ;
  assign \new_[12227]_  = \new_[14993]_  | \new_[19727]_ ;
  assign \new_[12228]_  = ~\new_[15039]_  | ~\new_[19547]_ ;
  assign \new_[12229]_  = ~\new_[13573]_ ;
  assign \new_[12230]_  = ~\new_[13574]_ ;
  assign \new_[12231]_  = ~\new_[14445]_ ;
  assign \new_[12232]_  = ~\new_[16935]_  | ~\new_[17532]_  | ~\new_[19018]_  | ~\new_[18012]_ ;
  assign \new_[12233]_  = ~\new_[13577]_ ;
  assign \new_[12234]_  = ~\new_[17277]_  | ~\new_[19096]_ ;
  assign \new_[12235]_  = ~\new_[15145]_  & ~\new_[19476]_ ;
  assign \new_[12236]_  = ~\new_[13584]_ ;
  assign \new_[12237]_  = ~\new_[15443]_  | ~\new_[18643]_ ;
  assign \new_[12238]_  = \new_[15379]_  | \new_[18017]_ ;
  assign \new_[12239]_  = ~\new_[15314]_  | ~\new_[19084]_ ;
  assign \new_[12240]_  = ~\new_[15086]_  & ~\new_[19024]_ ;
  assign \new_[12241]_  = \new_[16882]_  | \new_[19398]_  | \new_[18941]_  | \new_[18489]_ ;
  assign \new_[12242]_  = ~\new_[15288]_  | ~\new_[18070]_ ;
  assign \new_[12243]_  = ~\new_[15137]_  & ~\new_[19746]_ ;
  assign \new_[12244]_  = ~\new_[17162]_  & ~\new_[21306]_ ;
  assign \new_[12245]_  = \new_[15740]_  | \new_[18166]_ ;
  assign \new_[12246]_  = \new_[15250]_  | \new_[19547]_ ;
  assign \new_[12247]_  = ~\new_[15077]_  | ~\new_[18008]_ ;
  assign \new_[12248]_  = ~\new_[17556]_  | ~\new_[19047]_  | ~\new_[19750]_  | ~\new_[19096]_ ;
  assign \new_[12249]_  = ~\new_[15788]_  | ~\new_[19409]_ ;
  assign \new_[12250]_  = ~\new_[13591]_ ;
  assign \new_[12251]_  = \new_[15311]_  | \new_[19247]_ ;
  assign \new_[12252]_  = ~\new_[15788]_  | ~\new_[19436]_ ;
  assign \new_[12253]_  = ~\new_[17278]_  | ~\new_[18740]_  | ~\new_[18926]_  | ~\new_[18577]_ ;
  assign \new_[12254]_  = \new_[15227]_  | \new_[19008]_ ;
  assign \new_[12255]_  = ~\new_[13593]_ ;
  assign \new_[12256]_  = \new_[16916]_  | \new_[21580]_  | \new_[18046]_  | \new_[21505]_ ;
  assign \new_[12257]_  = ~\new_[19018]_  & ~\new_[14839]_ ;
  assign \new_[12258]_  = \new_[15556]_  | \new_[18008]_ ;
  assign \new_[12259]_  = \new_[18542]_  | \new_[15115]_ ;
  assign \new_[12260]_  = ~\new_[14968]_  | ~\new_[19196]_ ;
  assign \new_[12261]_  = \new_[19064]_  | \new_[15092]_ ;
  assign \new_[12262]_  = ~\new_[15477]_  | ~\new_[18998]_ ;
  assign \new_[12263]_  = ~\new_[15142]_  & ~\new_[19050]_ ;
  assign \new_[12264]_  = ~\new_[15253]_  & ~\new_[19249]_ ;
  assign \new_[12265]_  = ~\new_[15009]_  | ~\new_[16879]_ ;
  assign \new_[12266]_  = \new_[19202]_  | \new_[15106]_ ;
  assign \new_[12267]_  = ~\new_[15073]_  & ~\new_[17457]_ ;
  assign \new_[12268]_  = ~\new_[19094]_  & ~\new_[15084]_ ;
  assign \new_[12269]_  = ~\new_[14845]_  | ~\new_[18194]_ ;
  assign \new_[12270]_  = ~\new_[15223]_  | ~\new_[18693]_ ;
  assign \new_[12271]_  = ~\new_[14979]_  | ~\new_[18817]_ ;
  assign \new_[12272]_  = ~\new_[15348]_  & ~\new_[18087]_ ;
  assign \new_[12273]_  = ~\new_[15052]_  & ~\new_[18965]_ ;
  assign \new_[12274]_  = ~\new_[17556]_  | ~\new_[17532]_  | ~\new_[21635]_  | ~\new_[18012]_ ;
  assign \new_[12275]_  = ~\new_[14907]_  & ~\new_[18778]_ ;
  assign \new_[12276]_  = ~\new_[14932]_  | ~\new_[19758]_ ;
  assign \new_[12277]_  = ~\new_[15179]_  | ~\new_[19253]_ ;
  assign \new_[12278]_  = ~\new_[14980]_  | ~\new_[18076]_ ;
  assign \new_[12279]_  = ~\new_[15696]_  & ~\new_[18573]_ ;
  assign \new_[12280]_  = ~\new_[19098]_  | ~\new_[18391]_ ;
  assign \new_[12281]_  = ~\new_[15266]_  & ~\new_[19217]_ ;
  assign \new_[12282]_  = ~\new_[17348]_  | ~\new_[19035]_  | ~\new_[17886]_  | ~\new_[18111]_ ;
  assign \new_[12283]_  = ~\new_[15273]_  | ~\new_[19079]_ ;
  assign \new_[12284]_  = ~\new_[14895]_  & ~\new_[18325]_ ;
  assign \new_[12285]_  = ~\new_[15098]_  & ~\new_[19553]_ ;
  assign \new_[12286]_  = ~\new_[14819]_  & ~\new_[17979]_ ;
  assign \new_[12287]_  = ~\new_[15117]_  | ~\new_[19410]_ ;
  assign \new_[12288]_  = ~\new_[14993]_  & ~\new_[19561]_ ;
  assign \new_[12289]_  = ~\new_[20865]_  & ~\new_[21714]_ ;
  assign \new_[12290]_  = ~\new_[14973]_  & ~\new_[18443]_ ;
  assign \new_[12291]_  = ~\new_[15007]_  & ~\new_[19269]_ ;
  assign \new_[12292]_  = ~\new_[17522]_  | ~\new_[14887]_ ;
  assign \new_[12293]_  = ~\new_[14833]_  | ~\new_[19050]_ ;
  assign \new_[12294]_  = ~\new_[14739]_  | ~\new_[19188]_ ;
  assign \new_[12295]_  = ~\new_[20239]_  | ~\new_[15146]_ ;
  assign \new_[12296]_  = ~\new_[13608]_ ;
  assign \new_[12297]_  = ~\new_[15312]_  | ~\new_[17314]_ ;
  assign \new_[12298]_  = ~\new_[16201]_  | ~\new_[15316]_ ;
  assign \new_[12299]_  = ~\new_[15487]_  | ~\new_[18832]_ ;
  assign \new_[12300]_  = ~\new_[18148]_  | ~\new_[21520]_  | ~\new_[17983]_  | ~\new_[17529]_ ;
  assign \new_[12301]_  = ~\new_[15134]_  | ~\new_[18845]_ ;
  assign \new_[12302]_  = ~\new_[15164]_  | ~\new_[19474]_ ;
  assign \new_[12303]_  = ~\new_[13675]_ ;
  assign \new_[12304]_  = ~\new_[13672]_ ;
  assign \new_[12305]_  = ~\new_[15669]_  | ~\new_[19224]_ ;
  assign \new_[12306]_  = ~\new_[15352]_  | ~\new_[18637]_ ;
  assign \new_[12307]_  = \new_[16222]_  & \new_[15049]_ ;
  assign \new_[12308]_  = ~\new_[17664]_  | ~\new_[14887]_ ;
  assign \new_[12309]_  = \new_[15246]_  | \new_[19553]_ ;
  assign \new_[12310]_  = ~\new_[14844]_  | ~\new_[19265]_ ;
  assign \new_[12311]_  = \new_[15057]_  | \new_[19547]_ ;
  assign \new_[12312]_  = ~\new_[20865]_  & ~\new_[16713]_ ;
  assign \new_[12313]_  = \new_[15256]_  | \new_[18938]_ ;
  assign \new_[12314]_  = ~\new_[13614]_ ;
  assign \new_[12315]_  = ~\new_[19084]_  & ~\new_[15354]_ ;
  assign \new_[12316]_  = ~\new_[18750]_  | ~\new_[14980]_ ;
  assign \new_[12317]_  = \new_[15325]_  | \new_[19553]_ ;
  assign \new_[12318]_  = ~\new_[16730]_  | ~\new_[15179]_ ;
  assign \new_[12319]_  = ~\new_[15013]_  | ~\new_[14810]_ ;
  assign \new_[12320]_  = \new_[15162]_  & \new_[19713]_ ;
  assign \new_[12321]_  = ~\new_[15091]_  | ~\new_[21689]_ ;
  assign \new_[12322]_  = \new_[15034]_  | \new_[18938]_ ;
  assign \new_[12323]_  = ~\new_[15506]_  | ~\new_[16280]_ ;
  assign \new_[12324]_  = ~\new_[15150]_  | ~\new_[19568]_ ;
  assign \new_[12325]_  = ~\new_[17878]_  | ~\new_[14923]_ ;
  assign \new_[12326]_  = ~\new_[14838]_  | ~\new_[19729]_ ;
  assign \new_[12327]_  = ~\new_[15236]_  | ~\new_[19036]_ ;
  assign \new_[12328]_  = ~\new_[15312]_  & ~\new_[19151]_ ;
  assign \new_[12329]_  = \new_[15169]_  & \new_[15052]_ ;
  assign \new_[12330]_  = ~\new_[15693]_  & ~\new_[19217]_ ;
  assign \new_[12331]_  = ~\new_[15103]_  | ~\new_[15122]_ ;
  assign \new_[12332]_  = ~\new_[15354]_  | ~\new_[17652]_ ;
  assign \new_[12333]_  = \new_[15104]_  | \new_[19727]_ ;
  assign \new_[12334]_  = ~\new_[15208]_  | ~\new_[16811]_ ;
  assign \new_[12335]_  = ~\new_[21136]_  | ~\new_[15198]_ ;
  assign \new_[12336]_  = ~\new_[17265]_  | ~\new_[15227]_ ;
  assign \new_[12337]_  = ~\new_[19072]_  & ~\new_[16243]_ ;
  assign \new_[12338]_  = ~\new_[15045]_  | ~\new_[19738]_ ;
  assign \new_[12339]_  = ~\new_[14733]_  | ~\new_[19228]_ ;
  assign \new_[12340]_  = ~\new_[14373]_ ;
  assign \new_[12341]_  = ~\new_[16775]_  | ~\new_[15211]_ ;
  assign \new_[12342]_  = ~\new_[13632]_ ;
  assign \new_[12343]_  = ~\new_[13617]_ ;
  assign \new_[12344]_  = ~\new_[15175]_  & ~\new_[19335]_ ;
  assign \new_[12345]_  = ~\new_[15260]_  & ~\new_[16120]_ ;
  assign \new_[12346]_  = ~\new_[15860]_  & ~\new_[18414]_ ;
  assign \new_[12347]_  = ~\new_[13629]_ ;
  assign \new_[12348]_  = ~\new_[17376]_  | ~\new_[14925]_ ;
  assign \new_[12349]_  = ~\new_[17098]_  | ~\new_[19409]_ ;
  assign \new_[12350]_  = ~\new_[13632]_ ;
  assign \new_[12351]_  = \new_[15102]_  | \new_[19156]_ ;
  assign \new_[12352]_  = ~\new_[14727]_  | ~\new_[15290]_ ;
  assign \new_[12353]_  = ~\new_[18998]_  & (~\new_[16425]_  | ~\new_[17656]_ );
  assign \new_[12354]_  = ~\new_[15804]_  | ~\new_[14809]_ ;
  assign \new_[12355]_  = \new_[15010]_  | \new_[19203]_ ;
  assign \new_[12356]_  = ~\new_[16513]_  | ~\new_[14918]_ ;
  assign \new_[12357]_  = ~\new_[20866]_  | ~\new_[17298]_ ;
  assign \new_[12358]_  = ~\new_[14261]_ ;
  assign \new_[12359]_  = \new_[17101]_  | \new_[18965]_ ;
  assign \new_[12360]_  = \new_[14803]_  & \new_[19553]_ ;
  assign \new_[12361]_  = ~\new_[13543]_ ;
  assign \new_[12362]_  = ~\new_[13873]_ ;
  assign \new_[12363]_  = ~\new_[15543]_  | ~\new_[21568]_ ;
  assign \new_[12364]_  = ~\new_[17143]_  | ~\new_[16353]_ ;
  assign \new_[12365]_  = ~\new_[16687]_  | ~\new_[17887]_  | ~\new_[15952]_ ;
  assign \new_[12366]_  = ~\new_[14699]_  | ~\new_[19636]_ ;
  assign \new_[12367]_  = ~\new_[14987]_  | ~\new_[18427]_ ;
  assign \new_[12368]_  = ~\new_[15265]_  | ~\new_[19410]_ ;
  assign \new_[12369]_  = ~\new_[21075]_  | ~\new_[21505]_ ;
  assign \new_[12370]_  = ~\new_[15478]_  | ~\new_[15241]_ ;
  assign \new_[12371]_  = ~\new_[15769]_  | ~\new_[14955]_ ;
  assign \new_[12372]_  = ~\new_[21621]_  | ~\new_[19084]_ ;
  assign \new_[12373]_  = ~\new_[15287]_  & ~\new_[19085]_ ;
  assign \new_[12374]_  = ~\new_[18361]_  & ~\new_[15210]_ ;
  assign \new_[12375]_  = ~\new_[18923]_  & ~\new_[14925]_ ;
  assign \new_[12376]_  = ~\new_[16224]_  | ~\new_[14791]_ ;
  assign \new_[12377]_  = ~\new_[15477]_  | ~\new_[18849]_ ;
  assign \new_[12378]_  = ~\new_[14917]_  | ~\new_[18969]_ ;
  assign \new_[12379]_  = ~\new_[15426]_  | ~\new_[19024]_ ;
  assign \new_[12380]_  = ~\new_[13641]_ ;
  assign \new_[12381]_  = ~\new_[13642]_ ;
  assign \new_[12382]_  = ~\new_[16708]_  | ~\new_[19478]_  | ~\new_[18957]_  | ~\new_[19379]_ ;
  assign \new_[12383]_  = ~\new_[19021]_  & (~\new_[16368]_  | ~\new_[17827]_ );
  assign \new_[12384]_  = ~\new_[13487]_ ;
  assign \new_[12385]_  = ~\new_[15257]_  | ~\new_[17409]_ ;
  assign \new_[12386]_  = ~\new_[21094]_  | ~\new_[19084]_ ;
  assign \new_[12387]_  = ~\new_[15070]_  | ~\new_[18974]_ ;
  assign \new_[12388]_  = ~\new_[16352]_  | ~\new_[15436]_ ;
  assign \new_[12389]_  = ~\new_[17003]_  & ~\new_[19196]_ ;
  assign \new_[12390]_  = ~\new_[13646]_ ;
  assign \new_[12391]_  = \new_[14997]_  | \new_[21638]_ ;
  assign \new_[12392]_  = ~\new_[13648]_ ;
  assign \new_[12393]_  = ~\new_[14804]_  & ~\new_[18840]_ ;
  assign \new_[12394]_  = ~\new_[14983]_  | ~\new_[19269]_ ;
  assign \new_[12395]_  = ~\new_[14879]_  & ~\new_[20100]_ ;
  assign \new_[12396]_  = ~\new_[15280]_  | ~\new_[19028]_ ;
  assign \new_[12397]_  = ~\new_[15004]_  | ~\new_[19151]_ ;
  assign \new_[12398]_  = ~\new_[16037]_  | ~\new_[19319]_ ;
  assign \new_[12399]_  = ~\new_[13650]_ ;
  assign \new_[12400]_  = ~\new_[15357]_  | ~\new_[18682]_ ;
  assign \new_[12401]_  = ~\new_[19094]_  & ~\new_[16262]_ ;
  assign \new_[12402]_  = ~\new_[15166]_  | ~\new_[15168]_ ;
  assign \new_[12403]_  = ~\new_[15156]_  | ~\new_[15051]_ ;
  assign \new_[12404]_  = ~\new_[15811]_  & (~\new_[17583]_  | ~\new_[17707]_ );
  assign \new_[12405]_  = ~\new_[18167]_  | ~\new_[17171]_ ;
  assign \new_[12406]_  = ~\new_[15415]_  | ~\new_[19746]_ ;
  assign \new_[12407]_  = ~\new_[15449]_  | ~\new_[15359]_ ;
  assign n2743 = ~\new_[18775]_  | (~\new_[16329]_  & ~\new_[19723]_ );
  assign \new_[12409]_  = ~\new_[15411]_  & ~\new_[18709]_ ;
  assign \new_[12410]_  = ~\new_[15696]_  | ~\new_[15220]_ ;
  assign \new_[12411]_  = ~\new_[15495]_  | ~\new_[15093]_ ;
  assign \new_[12412]_  = ~\new_[14258]_ ;
  assign \new_[12413]_  = ~\new_[13652]_ ;
  assign \new_[12414]_  = ~\new_[14860]_  & (~\new_[17993]_  | ~\new_[18138]_ );
  assign \new_[12415]_  = ~\new_[13653]_ ;
  assign \new_[12416]_  = ~\new_[15277]_  | ~\new_[15355]_ ;
  assign \new_[12417]_  = ~\new_[13654]_ ;
  assign \new_[12418]_  = ~\new_[15021]_  | ~\new_[19568]_ ;
  assign \new_[12419]_  = ~\new_[15858]_  | ~\new_[15185]_ ;
  assign \new_[12420]_  = ~\new_[13860]_ ;
  assign \new_[12421]_  = \new_[17225]_  | \new_[18421]_ ;
  assign \new_[12422]_  = ~\new_[14919]_  | ~\new_[17158]_ ;
  assign \new_[12423]_  = ~\new_[15254]_  & ~\new_[19532]_ ;
  assign \new_[12424]_  = ~\new_[21551]_  | ~\new_[18615]_ ;
  assign \new_[12425]_  = ~\new_[14086]_ ;
  assign \new_[12426]_  = ~\new_[17465]_  | ~\new_[18469]_  | ~\new_[16040]_ ;
  assign \new_[12427]_  = ~\new_[19275]_  & ~\new_[15606]_ ;
  assign \new_[12428]_  = ~\new_[14749]_  & (~\new_[18813]_  | ~\new_[6746]_ );
  assign \new_[12429]_  = ~\new_[13858]_ ;
  assign \new_[12430]_  = \new_[15169]_  & \new_[16159]_ ;
  assign \new_[12431]_  = ~\new_[16427]_  | ~\new_[15102]_ ;
  assign \new_[12432]_  = ~\new_[14747]_  | ~\new_[19758]_ ;
  assign \new_[12433]_  = ~\new_[14359]_ ;
  assign \new_[12434]_  = ~\new_[17062]_  | ~\new_[16807]_  | ~\new_[16320]_ ;
  assign \new_[12435]_  = ~\new_[21621]_  & ~\new_[16227]_ ;
  assign \new_[12436]_  = \new_[15122]_  | \new_[19153]_ ;
  assign \new_[12437]_  = ~\new_[17207]_  | ~\new_[15212]_ ;
  assign \new_[12438]_  = ~\new_[15193]_  & ~\new_[19440]_ ;
  assign \new_[12439]_  = \new_[15175]_  | \new_[19727]_ ;
  assign \new_[12440]_  = ~\new_[13898]_ ;
  assign \new_[12441]_  = ~\new_[15905]_  | ~\new_[16940]_  | ~\new_[17179]_ ;
  assign \new_[12442]_  = ~\new_[13669]_ ;
  assign \new_[12443]_  = \new_[15036]_  | \new_[19239]_ ;
  assign \new_[12444]_  = ~\new_[15374]_  & ~\new_[18017]_ ;
  assign \new_[12445]_  = ~\new_[15493]_  & ~\new_[21684]_ ;
  assign \new_[12446]_  = ~\new_[13852]_ ;
  assign \new_[12447]_  = ~\new_[20291]_  | ~\new_[21506]_ ;
  assign \new_[12448]_  = ~\new_[16395]_  | ~\new_[15034]_ ;
  assign \new_[12449]_  = \new_[19565]_  ^ \new_[15923]_ ;
  assign \new_[12450]_  = ~\new_[15712]_  | ~\new_[15135]_ ;
  assign \new_[12451]_  = ~\new_[13677]_ ;
  assign \new_[12452]_  = ~\new_[15724]_  | ~\new_[15307]_ ;
  assign \new_[12453]_  = ~\new_[15589]_  & ~\new_[15270]_ ;
  assign \new_[12454]_  = ~\new_[17236]_  & ~\new_[19082]_ ;
  assign \new_[12455]_  = ~\new_[13676]_ ;
  assign \new_[12456]_  = \new_[18320]_  | \new_[19874]_ ;
  assign \new_[12457]_  = ~\new_[15281]_  | (~\new_[18316]_  & ~\new_[18906]_ );
  assign \new_[12458]_  = ~\new_[16450]_  | ~\new_[15010]_ ;
  assign \new_[12459]_  = ~\new_[15604]_  | ~\new_[16256]_ ;
  assign \new_[12460]_  = ~\new_[18123]_  & (~\new_[18613]_  | ~\new_[17876]_ );
  assign \new_[12461]_  = ~\new_[15183]_  & (~\new_[16564]_  | ~\new_[18637]_ );
  assign \new_[12462]_  = ~\new_[15012]_  | ~\new_[14919]_ ;
  assign \new_[12463]_  = ~\new_[15296]_  & (~\new_[16602]_  | ~\new_[19188]_ );
  assign \new_[12464]_  = ~\new_[15131]_  | ~\new_[15174]_ ;
  assign \new_[12465]_  = ~\new_[17832]_  | ~\new_[16007]_ ;
  assign \new_[12466]_  = ~\new_[14235]_ ;
  assign \new_[12467]_  = ~\new_[15125]_  & ~\new_[15643]_ ;
  assign \new_[12468]_  = ~\new_[15202]_ ;
  assign \new_[12469]_  = ~\new_[17217]_  | ~\new_[18083]_ ;
  assign \new_[12470]_  = ~\new_[18439]_  & (~\new_[17848]_  | ~\new_[16380]_ );
  assign \new_[12471]_  = ~\new_[17016]_  | (~\new_[18259]_  & ~\new_[16535]_ );
  assign \new_[12472]_  = \new_[15244]_  & \new_[17488]_ ;
  assign \new_[12473]_  = ~\new_[14347]_ ;
  assign \new_[12474]_  = ~\new_[15223]_  & (~\new_[17758]_  | ~\new_[16942]_ );
  assign \new_[12475]_  = ~\new_[15725]_  | ~\new_[14806]_ ;
  assign \new_[12476]_  = ~\new_[15043]_  | (~\new_[19255]_  & ~\new_[19223]_ );
  assign \new_[12477]_  = ~\new_[15095]_  | (~\new_[18962]_  & ~\new_[17502]_ );
  assign \new_[12478]_  = ~\new_[18222]_  | (~\new_[15955]_  & ~\new_[16462]_ );
  assign \new_[12479]_  = \new_[15538]_  & \new_[15157]_ ;
  assign \new_[12480]_  = \new_[15721]_  & \new_[16199]_ ;
  assign \new_[12481]_  = \new_[16712]_  ? \new_[19033]_  : \new_[17584]_ ;
  assign \new_[12482]_  = ~\new_[15762]_  & ~\new_[16008]_ ;
  assign \new_[12483]_  = \new_[16377]_  & \new_[15188]_ ;
  assign \new_[12484]_  = ~\new_[13690]_ ;
  assign \new_[12485]_  = \new_[18858]_  ^ \new_[16581]_ ;
  assign \new_[12486]_  = \new_[15492]_  | \new_[18832]_ ;
  assign \new_[12487]_  = ~\new_[17901]_  | ~\new_[14955]_ ;
  assign \new_[12488]_  = ~\new_[13840]_ ;
  assign \new_[12489]_  = ~\new_[16772]_  & ~\new_[19088]_ ;
  assign \new_[12490]_  = ~\new_[13696]_ ;
  assign \new_[12491]_  = ~\new_[14681]_ ;
  assign \new_[12492]_  = ~\new_[13698]_ ;
  assign \new_[12493]_  = ~\new_[14677]_ ;
  assign \new_[12494]_  = ~\new_[13700]_ ;
  assign \new_[12495]_  = ~\new_[16899]_  & ~\new_[21688]_ ;
  assign \new_[12496]_  = ~\new_[14942]_  & ~\new_[17572]_ ;
  assign \new_[12497]_  = ~\new_[15422]_  & ~\new_[20239]_ ;
  assign \new_[12498]_  = ~\new_[15866]_  | ~\new_[21693]_ ;
  assign \new_[12499]_  = \new_[15423]_  | \new_[18794]_ ;
  assign \new_[12500]_  = \new_[15392]_  | \new_[18427]_ ;
  assign \new_[12501]_  = ~\new_[15471]_  & ~\new_[21688]_ ;
  assign \new_[12502]_  = \new_[16849]_  | \new_[15690]_ ;
  assign \new_[12503]_  = \new_[15637]_  | \new_[18209]_ ;
  assign \new_[12504]_  = ~\new_[13702]_ ;
  assign \new_[12505]_  = ~\new_[13702]_ ;
  assign \new_[12506]_  = ~\new_[13703]_ ;
  assign \new_[12507]_  = ~\new_[20663]_  | ~\new_[19261]_ ;
  assign \new_[12508]_  = ~\new_[13704]_ ;
  assign \new_[12509]_  = ~\new_[13704]_ ;
  assign \new_[12510]_  = ~\new_[14666]_ ;
  assign \new_[12511]_  = ~\new_[14664]_ ;
  assign \new_[12512]_  = ~\new_[13710]_ ;
  assign \new_[12513]_  = \new_[13710]_ ;
  assign \new_[12514]_  = \new_[15662]_  & \new_[19088]_ ;
  assign \new_[12515]_  = ~\new_[13711]_ ;
  assign \new_[12516]_  = ~\new_[16972]_  & ~\new_[18008]_ ;
  assign \new_[12517]_  = ~\new_[18143]_  | ~\new_[15523]_ ;
  assign \new_[12518]_  = ~\new_[13715]_ ;
  assign \new_[12519]_  = ~\new_[13717]_ ;
  assign \new_[12520]_  = ~\new_[13718]_ ;
  assign \new_[12521]_  = ~\new_[13719]_ ;
  assign \new_[12522]_  = ~\new_[13720]_ ;
  assign \new_[12523]_  = ~\new_[13723]_ ;
  assign \new_[12524]_  = ~\new_[15461]_  | ~\new_[18575]_ ;
  assign \new_[12525]_  = \new_[15676]_  & \new_[19587]_ ;
  assign \new_[12526]_  = ~\new_[14645]_ ;
  assign \new_[12527]_  = ~\new_[13724]_ ;
  assign \new_[12528]_  = ~\new_[15417]_  | ~\new_[19161]_ ;
  assign \new_[12529]_  = \new_[14834]_  & \new_[18973]_ ;
  assign \new_[12530]_  = ~\new_[13725]_ ;
  assign \new_[12531]_  = ~\new_[13726]_ ;
  assign \new_[12532]_  = ~\new_[13727]_ ;
  assign \new_[12533]_  = ~\new_[13729]_ ;
  assign \new_[12534]_  = ~\new_[14615]_ ;
  assign \new_[12535]_  = ~\new_[15419]_  | ~\new_[19050]_ ;
  assign \new_[12536]_  = ~\new_[15509]_  & ~\new_[20865]_ ;
  assign \new_[12537]_  = ~\new_[13734]_ ;
  assign \new_[12538]_  = ~\new_[13735]_ ;
  assign \new_[12539]_  = ~\new_[15618]_  | ~\new_[18692]_ ;
  assign \new_[12540]_  = \new_[14717]_  | \new_[18414]_ ;
  assign \new_[12541]_  = ~\new_[14571]_ ;
  assign \new_[12542]_  = ~\new_[18083]_  & ~\new_[14862]_ ;
  assign \new_[12543]_  = ~\new_[15765]_  | ~\new_[19082]_ ;
  assign \new_[12544]_  = \new_[17445]_  | \new_[19290]_ ;
  assign \new_[12545]_  = ~\new_[13737]_ ;
  assign \new_[12546]_  = ~\new_[14862]_  & ~\new_[18569]_ ;
  assign \new_[12547]_  = ~\new_[13741]_ ;
  assign \new_[12548]_  = ~\new_[15515]_  | ~\new_[20239]_ ;
  assign \new_[12549]_  = ~\new_[15120]_  & ~\new_[18427]_ ;
  assign \new_[12550]_  = ~\new_[18244]_  | ~\new_[19174]_  | ~\new_[19102]_  | ~\new_[18026]_ ;
  assign \new_[12551]_  = ~\new_[13742]_ ;
  assign \new_[12552]_  = ~\new_[15550]_  | ~\new_[19275]_ ;
  assign \new_[12553]_  = ~\new_[13745]_ ;
  assign \new_[12554]_  = ~\new_[15800]_  & ~\new_[18973]_ ;
  assign \new_[12555]_  = ~\new_[15687]_  | ~\new_[18637]_ ;
  assign \new_[12556]_  = ~\new_[15617]_  | ~\new_[21689]_ ;
  assign \new_[12557]_  = ~\new_[14802]_  | ~\new_[18076]_ ;
  assign \new_[12558]_  = ~\new_[15206]_  | ~\new_[19253]_ ;
  assign \new_[12559]_  = ~\new_[13753]_ ;
  assign \new_[12560]_  = ~\new_[14795]_  | ~\new_[21684]_ ;
  assign \new_[12561]_  = \new_[14811]_  | \new_[18930]_ ;
  assign \new_[12562]_  = ~\new_[13757]_ ;
  assign \new_[12563]_  = ~\new_[16914]_  | ~\new_[17024]_ ;
  assign \new_[12564]_  = ~\new_[13762]_ ;
  assign \new_[12565]_  = ~\new_[13766]_ ;
  assign \new_[12566]_  = ~\new_[13767]_ ;
  assign \new_[12567]_  = ~\new_[13772]_ ;
  assign \new_[12568]_  = ~\new_[15467]_  | ~\new_[19738]_ ;
  assign \new_[12569]_  = ~\new_[13774]_ ;
  assign \new_[12570]_  = ~\new_[13779]_ ;
  assign \new_[12571]_  = ~\new_[15390]_  & ~\new_[19094]_ ;
  assign \new_[12572]_  = ~\new_[15619]_  | ~\new_[19754]_ ;
  assign \new_[12573]_  = ~\new_[15690]_  | ~\new_[18228]_ ;
  assign \new_[12574]_  = ~\new_[13786]_ ;
  assign \new_[12575]_  = ~\new_[15662]_  | ~\new_[18166]_ ;
  assign \new_[12576]_  = ~\new_[13787]_ ;
  assign \new_[12577]_  = ~\new_[13788]_ ;
  assign \new_[12578]_  = \new_[15810]_  | \new_[15866]_ ;
  assign \new_[12579]_  = ~\new_[13789]_ ;
  assign \new_[12580]_  = ~\new_[15581]_  & ~\new_[19181]_ ;
  assign \new_[12581]_  = ~\new_[13793]_ ;
  assign \new_[12582]_  = ~\new_[15683]_  & ~\new_[21562]_ ;
  assign \new_[12583]_  = ~\new_[15413]_  & ~\new_[19268]_ ;
  assign \new_[12584]_  = \new_[13797]_ ;
  assign \new_[12585]_  = ~\new_[15689]_  | ~\new_[19462]_ ;
  assign \new_[12586]_  = ~\new_[13801]_ ;
  assign \new_[12587]_  = ~\new_[13802]_ ;
  assign \new_[12588]_  = ~\new_[14253]_ ;
  assign \new_[12589]_  = ~\new_[13803]_ ;
  assign \new_[12590]_  = ~\new_[13804]_ ;
  assign \new_[12591]_  = \new_[14728]_  & \new_[19750]_ ;
  assign \new_[12592]_  = ~\new_[15361]_  | ~\new_[20825]_ ;
  assign \new_[12593]_  = \new_[14881]_  | \new_[21560]_ ;
  assign \new_[12594]_  = ~\new_[15405]_  & ~\new_[19082]_ ;
  assign \new_[12595]_  = \new_[15392]_  | \new_[21115]_ ;
  assign \new_[12596]_  = ~\new_[14209]_ ;
  assign \new_[12597]_  = ~\new_[15166]_  & ~\new_[19091]_ ;
  assign \new_[12598]_  = ~\new_[16925]_  & ~\new_[21689]_ ;
  assign \new_[12599]_  = ~\new_[14947]_  | ~\new_[19217]_ ;
  assign \new_[12600]_  = ~\new_[15421]_  & ~\new_[19381]_ ;
  assign \new_[12601]_  = ~\new_[15045]_ ;
  assign \new_[12602]_  = ~\new_[16720]_  | ~\new_[19224]_ ;
  assign \new_[12603]_  = ~\new_[14938]_  | ~\new_[19217]_ ;
  assign \new_[12604]_  = \new_[15748]_  | \new_[18335]_ ;
  assign \new_[12605]_  = ~\new_[13813]_ ;
  assign \new_[12606]_  = ~\new_[15678]_  | ~\new_[19697]_ ;
  assign \new_[12607]_  = ~\new_[15683]_  & ~\new_[19681]_ ;
  assign \new_[12608]_  = \new_[15437]_  | \new_[18766]_ ;
  assign \new_[12609]_  = ~\new_[15345]_  | ~\new_[18037]_ ;
  assign \new_[12610]_  = ~\new_[13818]_ ;
  assign \new_[12611]_  = ~\new_[13820]_ ;
  assign \new_[12612]_  = \new_[15410]_  | \new_[17572]_ ;
  assign \new_[12613]_  = ~\new_[15526]_  & ~\new_[21689]_ ;
  assign \new_[12614]_  = ~\new_[15699]_  & ~\new_[19082]_ ;
  assign \new_[12615]_  = ~\new_[13822]_ ;
  assign \new_[12616]_  = \new_[15553]_  | \new_[18414]_ ;
  assign \new_[12617]_  = ~\new_[13916]_ ;
  assign \new_[12618]_  = \new_[17353]_  | \new_[18414]_ ;
  assign \new_[12619]_  = \new_[14872]_  | \new_[18692]_ ;
  assign \new_[12620]_  = ~\new_[16769]_  & ~\new_[18228]_ ;
  assign \new_[12621]_  = ~\new_[15794]_  & ~\new_[19625]_ ;
  assign \new_[12622]_  = ~\new_[15141]_  | ~\new_[19801]_ ;
  assign \new_[12623]_  = ~\new_[17182]_  & ~\new_[21328]_ ;
  assign \new_[12624]_  = \new_[15453]_  | \new_[19261]_ ;
  assign \new_[12625]_  = ~\new_[13830]_ ;
  assign \new_[12626]_  = ~\new_[13829]_ ;
  assign \new_[12627]_  = \new_[15300]_  | \new_[20490]_ ;
  assign \new_[12628]_  = \new_[15486]_  & \new_[18083]_ ;
  assign \new_[12629]_  = ~\new_[13833]_ ;
  assign \new_[12630]_  = ~\new_[14712]_  & ~\new_[19474]_ ;
  assign \new_[12631]_  = ~\new_[13748]_ ;
  assign \new_[12632]_  = ~\new_[18436]_  & (~\new_[15930]_  | ~\new_[18890]_ );
  assign \new_[12633]_  = \new_[14836]_  | \new_[19474]_ ;
  assign \new_[12634]_  = ~\new_[15645]_  | ~\new_[18166]_ ;
  assign \new_[12635]_  = ~\new_[13837]_ ;
  assign \new_[12636]_  = ~\new_[15626]_  | ~\new_[21507]_ ;
  assign \new_[12637]_  = \new_[14710]_  & \new_[19181]_ ;
  assign \new_[12638]_  = ~\new_[13688]_ ;
  assign \new_[12639]_  = ~\new_[15501]_  | ~\new_[18709]_ ;
  assign \new_[12640]_  = \new_[15841]_  | \new_[19249]_ ;
  assign \new_[12641]_  = ~\new_[13845]_ ;
  assign \new_[12642]_  = ~\new_[15191]_  | ~\new_[19474]_ ;
  assign \new_[12643]_  = ~\new_[20234]_  & ~\new_[19036]_ ;
  assign \new_[12644]_  = ~\new_[13846]_ ;
  assign \new_[12645]_  = \new_[14948]_  ^ \new_[19578]_ ;
  assign \new_[12646]_  = ~\new_[16007]_  | ~\new_[18984]_ ;
  assign \new_[12647]_  = ~\new_[15391]_  | ~\new_[19181]_ ;
  assign \new_[12648]_  = ~\new_[15590]_  | ~\new_[19240]_ ;
  assign \new_[12649]_  = ~\new_[13848]_ ;
  assign \new_[12650]_  = ~\new_[17052]_  & ~\new_[19158]_ ;
  assign \new_[12651]_  = ~\new_[16501]_  | ~\new_[19018]_ ;
  assign \new_[12652]_  = ~\new_[15651]_  | ~\new_[18984]_ ;
  assign \new_[12653]_  = ~\new_[14849]_  | ~\new_[18938]_ ;
  assign \new_[12654]_  = ~\new_[15495]_  & ~\new_[20490]_ ;
  assign \new_[12655]_  = ~\new_[13854]_ ;
  assign \new_[12656]_  = \new_[15609]_  | \new_[17452]_ ;
  assign \new_[12657]_  = ~\new_[13856]_ ;
  assign \new_[12658]_  = ~\new_[13664]_ ;
  assign \new_[12659]_  = ~\new_[15625]_  | ~\new_[19409]_ ;
  assign \new_[12660]_  = ~\new_[17203]_  & ~\new_[19181]_ ;
  assign \new_[12661]_  = ~\new_[13859]_ ;
  assign \new_[12662]_  = ~\new_[15527]_  & ~\new_[19181]_ ;
  assign \new_[12663]_  = ~\new_[14629]_ ;
  assign \new_[12664]_  = ~\new_[14914]_  | ~\new_[19044]_ ;
  assign \new_[12665]_  = ~\new_[13864]_ ;
  assign \new_[12666]_  = \new_[21672]_  | \new_[19436]_ ;
  assign \new_[12667]_  = ~\new_[13647]_ ;
  assign \new_[12668]_  = ~\new_[15552]_  & ~\new_[19102]_ ;
  assign \new_[12669]_  = ~\new_[13643]_ ;
  assign \new_[12670]_  = ~\new_[14744]_  | ~\new_[21574]_ ;
  assign \new_[12671]_  = ~\new_[21326]_  & ~\new_[19084]_ ;
  assign \new_[12672]_  = ~\new_[13874]_ ;
  assign \new_[12673]_  = ~\new_[18979]_  & ~\new_[15445]_ ;
  assign \new_[12674]_  = ~\new_[15776]_  & ~\new_[18577]_ ;
  assign \new_[12675]_  = ~\new_[13625]_ ;
  assign \new_[12676]_  = ~\new_[13876]_ ;
  assign \new_[12677]_  = ~\new_[17036]_  & ~\new_[18692]_ ;
  assign \new_[12678]_  = ~\new_[13624]_ ;
  assign \new_[12679]_  = \new_[13624]_ ;
  assign \new_[12680]_  = ~\new_[15741]_  | ~\new_[16840]_ ;
  assign \new_[12681]_  = \new_[15453]_  | \new_[21689]_ ;
  assign \new_[12682]_  = \new_[15406]_  | \new_[21394]_ ;
  assign \new_[12683]_  = \new_[13878]_ ;
  assign \new_[12684]_  = ~\new_[15452]_  & ~\new_[19084]_ ;
  assign \new_[12685]_  = ~\new_[16880]_  & ~\new_[18747]_ ;
  assign \new_[12686]_  = ~\new_[15447]_  & ~\new_[18709]_ ;
  assign \new_[12687]_  = ~\new_[12757]_  & ~\new_[18337]_ ;
  assign \new_[12688]_  = ~\new_[13879]_ ;
  assign \new_[12689]_  = ~\new_[13825]_ ;
  assign \new_[12690]_  = ~\new_[14707]_  & ~\new_[21513]_ ;
  assign \new_[12691]_  = ~\new_[18811]_  | ~\new_[19174]_  | ~\new_[18244]_  | ~\new_[18026]_ ;
  assign \new_[12692]_  = \new_[14881]_  | \new_[19275]_ ;
  assign \new_[12693]_  = \new_[19775]_  ^ \new_[17484]_ ;
  assign \new_[12694]_  = ~\new_[14841]_  | ~\new_[18692]_ ;
  assign \new_[12695]_  = ~\new_[15754]_  | ~\new_[19024]_ ;
  assign \new_[12696]_  = ~\new_[15627]_  | ~\new_[18008]_ ;
  assign \new_[12697]_  = ~\new_[13590]_ ;
  assign \new_[12698]_  = ~\new_[15013]_  & ~\new_[18587]_ ;
  assign \new_[12699]_  = ~\new_[15484]_  | ~\new_[17457]_ ;
  assign \new_[12700]_  = ~\new_[13581]_ ;
  assign \new_[12701]_  = ~\new_[13575]_ ;
  assign \new_[12702]_  = \new_[15448]_  | \new_[18083]_ ;
  assign \new_[12703]_  = ~\new_[15536]_  | ~\new_[18965]_ ;
  assign \new_[12704]_  = ~\new_[14869]_  & ~\new_[18605]_ ;
  assign \new_[12705]_  = ~\new_[13881]_ ;
  assign \new_[12706]_  = ~\new_[13563]_ ;
  assign \new_[12707]_  = ~\new_[13889]_ ;
  assign \new_[12708]_  = \new_[14738]_  & \new_[19275]_ ;
  assign \new_[12709]_  = ~\new_[13547]_ ;
  assign \new_[12710]_  = ~\new_[17169]_  | ~\new_[19084]_ ;
  assign \new_[12711]_  = ~\new_[13897]_ ;
  assign \new_[12712]_  = ~\new_[13897]_ ;
  assign \new_[12713]_  = ~\new_[14938]_  | ~\new_[19059]_ ;
  assign \new_[12714]_  = ~\new_[17203]_  & ~\new_[21563]_ ;
  assign \new_[12715]_  = ~\new_[13539]_ ;
  assign \new_[12716]_  = \new_[15400]_  | \new_[18362]_ ;
  assign \new_[12717]_  = \new_[15408]_  | \new_[19386]_ ;
  assign \new_[12718]_  = \new_[16900]_  | \new_[18832]_ ;
  assign \new_[12719]_  = ~\new_[15472]_  | ~\new_[18840]_ ;
  assign \new_[12720]_  = ~\new_[15676]_  | ~\new_[18692]_ ;
  assign \new_[12721]_  = ~\new_[18678]_  & ~\new_[15516]_ ;
  assign \new_[12722]_  = ~\new_[15794]_  & ~\new_[19068]_ ;
  assign \new_[12723]_  = ~\new_[13904]_ ;
  assign \new_[12724]_  = ~\new_[13530]_ ;
  assign \new_[12725]_  = ~\new_[14229]_ ;
  assign \new_[12726]_  = ~\new_[17095]_  | ~\new_[19327]_ ;
  assign \new_[12727]_  = \new_[21549]_  | \new_[19050]_ ;
  assign \new_[12728]_  = ~\new_[13905]_ ;
  assign \new_[12729]_  = ~\new_[13712]_ ;
  assign \new_[12730]_  = ~\new_[13532]_ ;
  assign \new_[12731]_  = ~\new_[21593]_  & ~\new_[18682]_ ;
  assign \new_[12732]_  = ~\new_[15587]_  | ~\new_[18972]_ ;
  assign \new_[12733]_  = ~\new_[13910]_ ;
  assign \new_[12734]_  = ~\new_[14743]_  | ~\new_[19008]_ ;
  assign \new_[12735]_  = ~\new_[13911]_ ;
  assign \new_[12736]_  = ~\new_[15649]_  | ~\new_[20485]_ ;
  assign \new_[12737]_  = ~\new_[13914]_ ;
  assign \new_[12738]_  = ~\new_[13914]_ ;
  assign \new_[12739]_  = ~\new_[15339]_  | ~\new_[18597]_ ;
  assign \new_[12740]_  = ~\new_[15393]_  & ~\new_[18008]_ ;
  assign \new_[12741]_  = ~\new_[15647]_  | ~\new_[18124]_ ;
  assign \new_[12742]_  = \new_[15119]_  | \new_[19754]_ ;
  assign \new_[12743]_  = ~\new_[17909]_  | ~\new_[17277]_ ;
  assign \new_[12744]_  = ~\new_[13919]_ ;
  assign \new_[12745]_  = ~\new_[13920]_ ;
  assign \new_[12746]_  = ~\new_[15382]_  | ~\new_[19268]_ ;
  assign \new_[12747]_  = ~\new_[14731]_  | ~\new_[18682]_ ;
  assign \new_[12748]_  = ~\new_[15594]_  & ~\new_[18972]_ ;
  assign \new_[12749]_  = ~\new_[13512]_ ;
  assign \new_[12750]_  = ~\new_[13511]_ ;
  assign \new_[12751]_  = ~\new_[13923]_ ;
  assign \new_[12752]_  = ~\new_[13924]_ ;
  assign \new_[12753]_  = ~\new_[13510]_ ;
  assign \new_[12754]_  = ~\new_[13510]_ ;
  assign \new_[12755]_  = \new_[14751]_  & \new_[19052]_ ;
  assign \new_[12756]_  = ~\new_[15689]_  | ~\new_[21558]_ ;
  assign \new_[12757]_  = ~\new_[20489]_ ;
  assign \new_[12758]_  = ~\new_[13507]_ ;
  assign \new_[12759]_  = ~\new_[13505]_ ;
  assign \new_[12760]_  = ~\new_[13938]_ ;
  assign \new_[12761]_  = ~\new_[13501]_ ;
  assign \new_[12762]_  = \new_[15750]_  & \new_[18783]_ ;
  assign \new_[12763]_  = ~\new_[15864]_  | ~\new_[17457]_ ;
  assign \new_[12764]_  = \new_[16409]_  | \new_[18111]_ ;
  assign \new_[12765]_  = ~\new_[15459]_  & ~\new_[18926]_ ;
  assign \new_[12766]_  = ~\new_[14708]_  & ~\new_[19687]_ ;
  assign \new_[12767]_  = ~\new_[21507]_  & ~\new_[15620]_ ;
  assign \new_[12768]_  = ~\new_[13946]_ ;
  assign \new_[12769]_  = ~\new_[13946]_ ;
  assign \new_[12770]_  = \new_[15997]_  | \new_[15767]_ ;
  assign \new_[12771]_  = ~\new_[14738]_  | ~\new_[21394]_ ;
  assign \new_[12772]_  = ~\new_[21096]_  & ~\new_[19084]_ ;
  assign \new_[12773]_  = \new_[15552]_  | \new_[19082]_ ;
  assign \new_[12774]_  = ~\new_[13953]_ ;
  assign \new_[12775]_  = ~\new_[15558]_  | ~\new_[19750]_ ;
  assign \new_[12776]_  = ~\new_[21607]_  & ~\new_[19215]_ ;
  assign \new_[12777]_  = ~\new_[14921]_  | ~\new_[14951]_ ;
  assign \new_[12778]_  = ~\new_[13958]_ ;
  assign \new_[12779]_  = \new_[15384]_  | \new_[17457]_ ;
  assign \new_[12780]_  = ~\new_[14891]_  | ~\new_[17886]_ ;
  assign \new_[12781]_  = ~\new_[13960]_ ;
  assign \new_[12782]_  = ~\new_[21257]_ ;
  assign \new_[12783]_  = ~\new_[15579]_  | ~\new_[18448]_ ;
  assign \new_[12784]_  = ~\new_[13962]_ ;
  assign \new_[12785]_  = \new_[14746]_  | \new_[18496]_ ;
  assign \new_[12786]_  = ~\new_[13969]_ ;
  assign \new_[12787]_  = ~\new_[14916]_  & ~\new_[21056]_ ;
  assign \new_[12788]_  = ~\new_[13970]_ ;
  assign \new_[12789]_  = ~\new_[14914]_  | ~\new_[18973]_ ;
  assign \new_[12790]_  = ~\new_[15449]_  & ~\new_[19801]_ ;
  assign \new_[12791]_  = ~\new_[14651]_ ;
  assign \new_[12792]_  = \new_[17102]_  | \new_[18938]_ ;
  assign \new_[12793]_  = ~\new_[17813]_  | ~\new_[14955]_ ;
  assign \new_[12794]_  = ~\new_[13977]_ ;
  assign \new_[12795]_  = ~\new_[13978]_ ;
  assign \new_[12796]_  = ~\new_[14734]_  | ~\new_[18766]_ ;
  assign \new_[12797]_  = ~\new_[13979]_ ;
  assign \new_[12798]_  = ~\new_[20927]_  & ~\new_[14900]_ ;
  assign \new_[12799]_  = ~\new_[15773]_  | ~\new_[19204]_ ;
  assign \new_[12800]_  = ~\new_[13981]_ ;
  assign \new_[12801]_  = ~\new_[13983]_ ;
  assign \new_[12802]_  = \new_[15463]_  & \new_[21496]_ ;
  assign \new_[12803]_  = \new_[20036]_  | \new_[21499]_ ;
  assign \new_[12804]_  = \new_[15494]_  & \new_[18166]_ ;
  assign \new_[12805]_  = \new_[20222]_ ;
  assign \new_[12806]_  = ~\new_[15545]_  & ~\new_[16840]_ ;
  assign \new_[12807]_  = ~\new_[16891]_  | ~\new_[18046]_ ;
  assign \new_[12808]_  = ~\new_[15611]_  | ~\new_[19203]_ ;
  assign \new_[12809]_  = ~\new_[13986]_ ;
  assign \new_[12810]_  = ~\new_[15554]_  | ~\new_[19224]_ ;
  assign \new_[12811]_  = ~\new_[15412]_  | ~\new_[20680]_ ;
  assign \new_[12812]_  = ~\new_[14598]_ ;
  assign \new_[12813]_  = ~\new_[15814]_  & ~\new_[18840]_ ;
  assign \new_[12814]_  = ~\new_[13821]_ ;
  assign \new_[12815]_  = ~\new_[16037]_  | ~\new_[19288]_ ;
  assign \new_[12816]_  = ~\new_[16027]_  | ~\new_[18973]_ ;
  assign \new_[12817]_  = ~\new_[15418]_  & ~\new_[19036]_ ;
  assign \new_[12818]_  = \new_[19096]_  | \new_[15355]_ ;
  assign \new_[12819]_  = ~\new_[15590]_  | ~\new_[18443]_ ;
  assign \new_[12820]_  = ~\new_[16562]_  | ~\new_[18440]_ ;
  assign \new_[12821]_  = \new_[18215]_  | \new_[19874]_ ;
  assign \new_[12822]_  = ~\new_[13991]_ ;
  assign \new_[12823]_  = ~\new_[13991]_ ;
  assign \new_[12824]_  = ~\new_[19554]_  & ~\new_[15192]_ ;
  assign \new_[12825]_  = ~\new_[18501]_  & ~\new_[15427]_ ;
  assign \new_[12826]_  = ~\new_[15752]_  | ~\new_[19130]_ ;
  assign \new_[12827]_  = ~\new_[18185]_  | ~\new_[15777]_ ;
  assign \new_[12828]_  = ~\new_[14532]_ ;
  assign \new_[12829]_  = ~\new_[13993]_ ;
  assign \new_[12830]_  = ~\new_[15648]_  & ~\new_[19290]_ ;
  assign \new_[12831]_  = ~\new_[18446]_  & ~\new_[15664]_ ;
  assign \new_[12832]_  = \new_[18706]_  | \new_[14954]_ ;
  assign \new_[12833]_  = ~\new_[17583]_  & ~\new_[15811]_ ;
  assign \new_[12834]_  = ~\new_[16693]_  & ~\new_[17381]_ ;
  assign \new_[12835]_  = ~\new_[17339]_  | ~\new_[17145]_ ;
  assign \new_[12836]_  = \new_[15409]_  & \new_[15455]_ ;
  assign \new_[12837]_  = \new_[15562]_  | \new_[21565]_ ;
  assign \new_[12838]_  = ~\new_[13997]_ ;
  assign \new_[12839]_  = ~\new_[16076]_  | ~\new_[21693]_ ;
  assign \new_[12840]_  = ~\new_[17713]_  | ~\new_[15777]_ ;
  assign \new_[12841]_  = ~\new_[17266]_  & ~\new_[18766]_ ;
  assign \new_[12842]_  = ~\new_[18260]_  | ~\new_[15523]_ ;
  assign \new_[12843]_  = ~\new_[14004]_ ;
  assign \new_[12844]_  = ~\new_[18360]_  | ~\new_[14955]_ ;
  assign \new_[12845]_  = ~\new_[14006]_ ;
  assign \new_[12846]_  = ~\new_[15197]_  & ~\new_[19059]_ ;
  assign \new_[12847]_  = ~\new_[15709]_  & ~\new_[21570]_ ;
  assign \new_[12848]_  = ~\new_[14008]_ ;
  assign \new_[12849]_  = ~\new_[14010]_ ;
  assign \new_[12850]_  = ~\new_[14011]_ ;
  assign \new_[12851]_  = ~\new_[16943]_  & ~\new_[18966]_ ;
  assign \new_[12852]_  = ~\new_[15151]_  & ~\new_[18414]_ ;
  assign \new_[12853]_  = ~\new_[14420]_ ;
  assign \new_[12854]_  = ~\new_[15508]_  & ~\new_[18817]_ ;
  assign \new_[12855]_  = \new_[17893]_  | \new_[19874]_ ;
  assign \new_[12856]_  = ~\new_[14017]_ ;
  assign \new_[12857]_  = ~\new_[14379]_ ;
  assign \new_[12858]_  = ~\new_[15451]_  | ~\new_[19194]_ ;
  assign \new_[12859]_  = ~\new_[15521]_  | ~\new_[19801]_ ;
  assign \new_[12860]_  = ~\new_[14019]_ ;
  assign \new_[12861]_  = ~\new_[15173]_  & ~\new_[19754]_ ;
  assign \new_[12862]_  = ~\new_[14526]_  & ~\new_[18973]_ ;
  assign \new_[12863]_  = ~\new_[14745]_  | ~\new_[16958]_ ;
  assign \new_[12864]_  = ~\new_[17894]_  | ~\new_[14955]_ ;
  assign \new_[12865]_  = ~\new_[14964]_  | ~\new_[17067]_ ;
  assign \new_[12866]_  = ~\new_[15517]_  | ~\new_[19268]_ ;
  assign \new_[12867]_  = ~\new_[14023]_ ;
  assign \new_[12868]_  = ~\new_[14026]_ ;
  assign \new_[12869]_  = ~\new_[14027]_ ;
  assign \new_[12870]_  = ~\new_[14028]_ ;
  assign \new_[12871]_  = ~\new_[14259]_ ;
  assign \new_[12872]_  = ~\new_[15542]_  & ~\new_[18605]_ ;
  assign \new_[12873]_  = ~\new_[18470]_  | ~\new_[14955]_ ;
  assign \new_[12874]_  = ~\new_[15427]_  & ~\new_[19202]_ ;
  assign \new_[12875]_  = ~\new_[17298]_  & ~\new_[20239]_ ;
  assign \new_[12876]_  = ~\new_[18106]_  & ~\new_[21604]_ ;
  assign \new_[12877]_  = ~\new_[14212]_ ;
  assign \new_[12878]_  = ~\new_[16748]_  & ~\new_[18762]_ ;
  assign \new_[12879]_  = ~\new_[15533]_  | ~\new_[18979]_ ;
  assign \new_[12880]_  = ~\new_[15631]_  & ~\new_[17381]_ ;
  assign \new_[12881]_  = ~\new_[13665]_ ;
  assign \new_[12882]_  = ~\new_[18788]_  | ~\new_[16486]_ ;
  assign \new_[12883]_  = ~\new_[15806]_  & ~\new_[19266]_ ;
  assign \new_[12884]_  = \new_[17691]_  | \new_[14954]_ ;
  assign \new_[12885]_  = ~\new_[20867]_  | ~\new_[20865]_ ;
  assign \new_[12886]_  = ~\new_[16072]_  | ~\new_[21096]_ ;
  assign \new_[12887]_  = ~\new_[15513]_  & ~\new_[18941]_ ;
  assign \new_[12888]_  = ~\new_[15300]_  | ~\new_[15053]_ ;
  assign \new_[12889]_  = ~\new_[21549]_  | ~\new_[15849]_ ;
  assign \new_[12890]_  = \new_[18936]_  | \new_[15510]_ ;
  assign \new_[12891]_  = ~\new_[14058]_ ;
  assign \new_[12892]_  = ~\new_[14044]_ ;
  assign \new_[12893]_  = ~\new_[14045]_ ;
  assign \new_[12894]_  = \new_[16751]_  & \new_[19319]_ ;
  assign \new_[12895]_  = ~\new_[14047]_ ;
  assign \new_[12896]_  = ~\new_[18321]_  | ~\new_[14955]_ ;
  assign \new_[12897]_  = ~\new_[18184]_  | ~\new_[15521]_ ;
  assign \new_[12898]_  = ~\new_[15679]_  | ~\new_[19079]_ ;
  assign \new_[12899]_  = ~\new_[14412]_ ;
  assign \new_[12900]_  = \new_[15635]_  | \new_[18414]_ ;
  assign \new_[12901]_  = ~\new_[18385]_  | ~\new_[15690]_ ;
  assign \new_[12902]_  = \new_[17820]_  | \new_[15530]_ ;
  assign \new_[12903]_  = \new_[15490]_  | \new_[20680]_ ;
  assign \new_[12904]_  = ~\new_[14050]_ ;
  assign \new_[12905]_  = ~\new_[13963]_ ;
  assign \new_[12906]_  = ~\new_[13963]_ ;
  assign \new_[12907]_  = \new_[15503]_  | \new_[18076]_ ;
  assign \new_[12908]_  = ~\new_[15094]_  & ~\new_[19064]_ ;
  assign \new_[12909]_  = \new_[18904]_  | \new_[15530]_ ;
  assign \new_[12910]_  = ~\new_[17551]_  | ~\new_[15417]_ ;
  assign \new_[12911]_  = ~\new_[14052]_ ;
  assign \new_[12912]_  = ~\new_[15719]_  | ~\new_[18469]_ ;
  assign \new_[12913]_  = ~\new_[14054]_ ;
  assign \new_[12914]_  = ~\new_[18295]_  | ~\new_[14955]_ ;
  assign \new_[12915]_  = ~\new_[13877]_ ;
  assign \new_[12916]_  = ~\new_[14057]_ ;
  assign \new_[12917]_  = ~\new_[21550]_  | ~\new_[19754]_ ;
  assign \new_[12918]_  = ~\new_[13806]_ ;
  assign \new_[12919]_  = ~\new_[15197]_  & ~\new_[19084]_ ;
  assign \new_[12920]_  = ~\new_[14065]_ ;
  assign \new_[12921]_  = ~\new_[18074]_  | ~\new_[14955]_ ;
  assign \new_[12922]_  = ~\new_[17314]_  & ~\new_[19151]_ ;
  assign \new_[12923]_  = \new_[15622]_  | \new_[18930]_ ;
  assign \new_[12924]_  = ~\new_[15502]_  & (~\new_[17474]_  | ~\new_[21394]_ );
  assign \new_[12925]_  = ~\new_[18403]_  | ~\new_[16798]_ ;
  assign \new_[12926]_  = ~\new_[14069]_ ;
  assign \new_[12927]_  = ~\new_[15685]_  | ~\new_[15392]_ ;
  assign \new_[12928]_  = ~\new_[18369]_  | ~\new_[16799]_ ;
  assign \new_[12929]_  = ~\new_[14072]_ ;
  assign \new_[12930]_  = \new_[17129]_  | \new_[14826]_ ;
  assign \new_[12931]_  = ~\new_[17849]_  | ~\new_[14955]_ ;
  assign \new_[12932]_  = ~\new_[13685]_ ;
  assign \new_[12933]_  = \new_[15469]_  | \new_[16572]_ ;
  assign \new_[12934]_  = ~\new_[17817]_  | ~\new_[15523]_ ;
  assign \new_[12935]_  = ~\new_[14077]_ ;
  assign \new_[12936]_  = ~\new_[19224]_  & ~\new_[16814]_ ;
  assign \new_[12937]_  = ~\new_[21664]_  | ~\new_[19241]_ ;
  assign \new_[12938]_  = ~\new_[16903]_  | ~\new_[18652]_ ;
  assign \new_[12939]_  = ~\new_[14081]_ ;
  assign \new_[12940]_  = ~\new_[14082]_ ;
  assign \new_[12941]_  = ~\new_[13668]_ ;
  assign \new_[12942]_  = ~\new_[15410]_  | ~\new_[17225]_ ;
  assign \new_[12943]_  = ~\new_[18179]_  | ~\new_[19228]_  | ~\new_[17852]_ ;
  assign \new_[12944]_  = ~\new_[17517]_  | ~\new_[14955]_ ;
  assign \new_[12945]_  = ~\new_[15659]_  | ~\new_[19697]_ ;
  assign \new_[12946]_  = \new_[15673]_  | \new_[16087]_ ;
  assign \new_[12947]_  = ~\new_[15659]_  | ~\new_[19642]_ ;
  assign \new_[12948]_  = \new_[15492]_  | \new_[19742]_ ;
  assign \new_[12949]_  = ~\new_[15601]_  & ~\new_[19244]_ ;
  assign \new_[12950]_  = ~\new_[15713]_  & ~\new_[18228]_ ;
  assign \new_[12951]_  = ~\new_[21574]_  & ~\new_[19687]_  & ~\new_[17539]_ ;
  assign \new_[12952]_  = \new_[15053]_  | \new_[18637]_ ;
  assign \new_[12953]_  = \new_[18869]_  & \new_[14827]_ ;
  assign \new_[12954]_  = ~\new_[17320]_  | ~\new_[14955]_ ;
  assign \new_[12955]_  = ~\new_[15402]_  | ~\new_[21508]_ ;
  assign \new_[12956]_  = ~\new_[17164]_  & ~\new_[18926]_ ;
  assign \new_[12957]_  = ~\new_[17424]_  & ~\new_[20099]_ ;
  assign \new_[12958]_  = ~\new_[15487]_  & (~\new_[17463]_  | ~\new_[18832]_ );
  assign \new_[12959]_  = ~\new_[14101]_ ;
  assign \new_[12960]_  = \new_[15469]_  | \new_[19068]_ ;
  assign \new_[12961]_  = ~\new_[18914]_  & ~\new_[15614]_ ;
  assign \new_[12962]_  = ~\new_[15605]_  | ~\new_[18833]_ ;
  assign \new_[12963]_  = ~\new_[15720]_  | ~\new_[17469]_ ;
  assign \new_[12964]_  = \new_[17779]_  | \new_[19874]_ ;
  assign \new_[12965]_  = ~\new_[17905]_  | ~\new_[15778]_ ;
  assign \new_[12966]_  = \new_[17164]_  | \new_[19592]_ ;
  assign \new_[12967]_  = ~\new_[16949]_  & ~\new_[15206]_ ;
  assign \new_[12968]_  = ~\new_[15245]_  & ~\new_[20865]_ ;
  assign \new_[12969]_  = \new_[15722]_  | \new_[19224]_ ;
  assign \new_[12970]_  = ~\new_[18794]_  & ~\new_[16698]_ ;
  assign \new_[12971]_  = ~\new_[15438]_  | ~\new_[17983]_ ;
  assign \new_[12972]_  = ~\new_[18432]_  | ~\new_[17632]_ ;
  assign \new_[12973]_  = ~\new_[20239]_  & (~\new_[16617]_  | ~\new_[17773]_ );
  assign \new_[12974]_  = ~\new_[17555]_  | ~\new_[15778]_ ;
  assign \new_[12975]_  = \new_[15709]_  | \new_[19409]_ ;
  assign \new_[12976]_  = ~\new_[13540]_ ;
  assign \new_[12977]_  = ~\new_[16584]_  | ~\new_[18826]_ ;
  assign \new_[12978]_  = ~\new_[14113]_ ;
  assign \new_[12979]_  = ~\new_[15704]_  | ~\new_[19446]_ ;
  assign \new_[12980]_  = ~\new_[15655]_  | ~\new_[19188]_ ;
  assign \new_[12981]_  = ~\new_[15542]_  & ~\new_[18337]_ ;
  assign \new_[12982]_  = ~\new_[21055]_  & ~\new_[17469]_ ;
  assign \new_[12983]_  = ~\new_[15559]_  & (~\new_[17352]_  | ~\new_[19186]_ );
  assign \new_[12984]_  = ~\new_[14120]_ ;
  assign \new_[12985]_  = ~\new_[14121]_ ;
  assign \new_[12986]_  = ~\new_[17073]_  | ~\new_[21166]_ ;
  assign \new_[12987]_  = ~\new_[19096]_  & ~\new_[15753]_ ;
  assign \new_[12988]_  = ~\new_[13525]_ ;
  assign \new_[12989]_  = ~\new_[17816]_  & ~\new_[14731]_ ;
  assign \new_[12990]_  = ~\new_[13524]_ ;
  assign \new_[12991]_  = \new_[16816]_  | \new_[18427]_ ;
  assign \new_[12992]_  = ~\new_[17435]_  & ~\new_[19676]_ ;
  assign \new_[12993]_  = ~\new_[14127]_ ;
  assign \new_[12994]_  = ~\new_[14135]_ ;
  assign \new_[12995]_  = \new_[14720]_  | \new_[18153]_ ;
  assign \new_[12996]_  = ~\new_[13500]_ ;
  assign \new_[12997]_  = ~\new_[15630]_  | ~\new_[18965]_ ;
  assign \new_[12998]_  = \new_[18514]_  | \new_[19874]_ ;
  assign \new_[12999]_  = \new_[17023]_  | \new_[14826]_ ;
  assign \new_[13000]_  = ~\new_[17578]_  | ~\new_[16646]_  | ~\new_[18050]_ ;
  assign \new_[13001]_  = ~\new_[18387]_  | ~\new_[15523]_ ;
  assign \new_[13002]_  = ~\new_[14714]_  & ~\new_[21513]_ ;
  assign \new_[13003]_  = ~\new_[13490]_ ;
  assign \new_[13004]_  = ~\new_[15704]_  | ~\new_[19100]_ ;
  assign \new_[13005]_  = \new_[15612]_  | \new_[18076]_ ;
  assign \new_[13006]_  = ~\new_[14147]_ ;
  assign \new_[13007]_  = ~\new_[14687]_ ;
  assign \new_[13008]_  = \new_[18220]_  | \new_[19874]_ ;
  assign \new_[13009]_  = ~\new_[15572]_  | ~\new_[18427]_ ;
  assign \new_[13010]_  = \new_[18366]_  | \new_[15530]_ ;
  assign \new_[13011]_  = ~\new_[14939]_  | ~\new_[14955]_ ;
  assign \new_[13012]_  = ~\new_[15546]_  | ~\new_[19088]_ ;
  assign \new_[13013]_  = ~\new_[17815]_  | ~\new_[14955]_ ;
  assign \new_[13014]_  = ~\new_[14152]_ ;
  assign \new_[13015]_  = \new_[21701]_  | \new_[21115]_ ;
  assign \new_[13016]_  = ~\new_[14155]_ ;
  assign \new_[13017]_  = ~\new_[14157]_ ;
  assign \new_[13018]_  = ~\new_[15596]_  | ~\new_[21558]_ ;
  assign \new_[13019]_  = ~\new_[17139]_  | ~\new_[19268]_ ;
  assign \new_[13020]_  = ~\new_[14159]_ ;
  assign \new_[13021]_  = ~\new_[17159]_  | ~\new_[18166]_ ;
  assign \new_[13022]_  = ~\new_[17891]_  | ~\new_[15777]_ ;
  assign \new_[13023]_  = ~\new_[17310]_  | ~\new_[14955]_ ;
  assign \new_[13024]_  = ~\new_[14163]_ ;
  assign \new_[13025]_  = ~\new_[16760]_  & ~\new_[19072]_ ;
  assign \new_[13026]_  = ~\new_[15315]_  & ~\new_[18326]_ ;
  assign \new_[13027]_  = ~\new_[14168]_ ;
  assign \new_[13028]_  = \new_[15681]_  | \new_[16140]_ ;
  assign \new_[13029]_  = ~\new_[14588]_ ;
  assign \new_[13030]_  = ~\new_[14174]_ ;
  assign \new_[13031]_  = ~\new_[14854]_  & ~\new_[17457]_ ;
  assign \new_[13032]_  = ~\new_[15245]_  & ~\new_[19240]_ ;
  assign \new_[13033]_  = ~\new_[15629]_  & ~\new_[16410]_ ;
  assign \new_[13034]_  = ~\new_[14178]_ ;
  assign \new_[13035]_  = ~\new_[18270]_  | ~\new_[15451]_ ;
  assign \new_[13036]_  = ~\new_[17435]_  & ~\new_[19033]_ ;
  assign \new_[13037]_  = ~\new_[15856]_  & ~\new_[16140]_ ;
  assign \new_[13038]_  = ~\new_[15552]_  & ~\new_[18711]_ ;
  assign \new_[13039]_  = ~\new_[16281]_  | ~\new_[21055]_ ;
  assign \new_[13040]_  = \new_[15252]_ ;
  assign \new_[13041]_  = ~\new_[15252]_ ;
  assign \new_[13042]_  = \new_[17829]_  | \new_[15530]_ ;
  assign \new_[13043]_  = \new_[17833]_  | \new_[19874]_ ;
  assign \new_[13044]_  = ~\new_[14185]_ ;
  assign \new_[13045]_  = ~\new_[14812]_  | (~\new_[18382]_  & ~\new_[17155]_ );
  assign \new_[13046]_  = ~\new_[14318]_ ;
  assign \new_[13047]_  = ~\new_[15837]_  & ~\new_[18664]_ ;
  assign \new_[13048]_  = \new_[19258]_  | \new_[15582]_ ;
  assign \new_[13049]_  = ~\new_[15441]_  | ~\new_[14876]_ ;
  assign \new_[13050]_  = \new_[17720]_  | \new_[14954]_ ;
  assign \new_[13051]_  = \new_[15859]_  | \new_[18448]_ ;
  assign \new_[13052]_  = ~\new_[14434]_ ;
  assign \new_[13053]_  = ~\new_[18102]_  & ~\new_[15711]_ ;
  assign \new_[13054]_  = ~\new_[15489]_  & ~\new_[18972]_ ;
  assign \new_[13055]_  = ~\new_[14197]_ ;
  assign \new_[13056]_  = ~\new_[15559]_  | ~\new_[18750]_ ;
  assign \new_[13057]_  = ~\new_[14200]_ ;
  assign \new_[13058]_  = ~\new_[14325]_ ;
  assign \new_[13059]_  = ~\new_[17373]_  | ~\new_[14748]_ ;
  assign \new_[13060]_  = ~\new_[14208]_ ;
  assign \new_[13061]_  = ~\new_[17408]_  & ~\new_[18228]_ ;
  assign \new_[13062]_  = ~\new_[14705]_  & ~\new_[18605]_ ;
  assign \new_[13063]_  = ~\new_[17904]_  | ~\new_[15777]_ ;
  assign \new_[13064]_  = ~\new_[20239]_  & ~\new_[16893]_ ;
  assign \new_[13065]_  = ~\new_[13431]_  & ~\new_[19729]_ ;
  assign \new_[13066]_  = \new_[15920]_  | \new_[15704]_ ;
  assign \new_[13067]_  = ~\new_[18487]_  | ~\new_[15777]_ ;
  assign \new_[13068]_  = ~\new_[14463]_ ;
  assign \new_[13069]_  = \new_[16177]_  & \new_[17616]_ ;
  assign \new_[13070]_  = ~\new_[17295]_  | ~\new_[16515]_ ;
  assign \new_[13071]_  = \new_[15574]_  | \new_[19290]_ ;
  assign \new_[13072]_  = \new_[15543]_  & \new_[19151]_ ;
  assign \new_[13073]_  = ~\new_[14137]_ ;
  assign \new_[13074]_  = ~\new_[15600]_  & ~\new_[19171]_ ;
  assign \new_[13075]_  = ~\new_[15847]_  & ~\new_[19154]_ ;
  assign \new_[13076]_  = ~\new_[16991]_  & ~\new_[19095]_ ;
  assign \new_[13077]_  = ~\new_[14084]_ ;
  assign \new_[13078]_  = ~\new_[17581]_  | ~\new_[17095]_ ;
  assign \new_[13079]_  = \new_[17902]_  | \new_[14826]_ ;
  assign \new_[13080]_  = ~\new_[14031]_ ;
  assign \new_[13081]_  = ~\new_[15566]_  | ~\new_[18621]_ ;
  assign \new_[13082]_  = ~\new_[16084]_  | ~\new_[14737]_ ;
  assign \new_[13083]_  = ~\new_[14219]_ ;
  assign \new_[13084]_  = \new_[17112]_  | \new_[17074]_ ;
  assign \new_[13085]_  = ~\new_[14220]_ ;
  assign \new_[13086]_  = ~\new_[14223]_ ;
  assign \new_[13087]_  = \new_[19169]_  | \new_[14815]_ ;
  assign \new_[13088]_  = ~\new_[14226]_ ;
  assign \new_[13089]_  = \new_[17376]_  | \new_[19181]_ ;
  assign \new_[13090]_  = ~\new_[16969]_  | ~\new_[15677]_ ;
  assign \new_[13091]_  = ~\new_[13880]_ ;
  assign \new_[13092]_  = \new_[15572]_  | \new_[15968]_ ;
  assign \new_[13093]_  = ~\new_[18906]_  | ~\new_[18750]_  | ~\new_[17505]_ ;
  assign \new_[13094]_  = ~\new_[15451]_  | ~\new_[18008]_ ;
  assign \new_[13095]_  = ~\new_[18158]_  | ~\new_[14955]_ ;
  assign \new_[13096]_  = ~\new_[15386]_  | ~\new_[15394]_ ;
  assign \new_[13097]_  = ~\new_[13824]_ ;
  assign \new_[13098]_  = \new_[15024]_  | \new_[18542]_ ;
  assign \new_[13099]_  = ~\new_[14239]_ ;
  assign \new_[13100]_  = ~\new_[17043]_  | ~\new_[14738]_ ;
  assign \new_[13101]_  = ~\new_[17315]_  | ~\new_[14955]_ ;
  assign \new_[13102]_  = ~\new_[15664]_  | ~\new_[15560]_ ;
  assign \new_[13103]_  = ~\new_[14812]_  | ~\new_[16959]_ ;
  assign \new_[13104]_  = \new_[15409]_  | \new_[19261]_ ;
  assign \new_[13105]_  = ~\new_[17052]_  & ~\new_[18373]_ ;
  assign \new_[13106]_  = ~\new_[13691]_ ;
  assign \new_[13107]_  = ~\new_[15812]_  | ~\new_[15682]_ ;
  assign \new_[13108]_  = ~\new_[14254]_ ;
  assign \new_[13109]_  = ~\new_[18289]_  | ~\new_[15777]_ ;
  assign \new_[13110]_  = ~\new_[17781]_  | ~\new_[15523]_ ;
  assign \new_[13111]_  = ~\new_[17838]_  | ~\new_[14955]_ ;
  assign \new_[13112]_  = ~\new_[18435]_  | ~\new_[14955]_ ;
  assign \new_[13113]_  = ~\new_[20927]_  & ~\new_[15698]_ ;
  assign \new_[13114]_  = ~\new_[16929]_  | ~\new_[19018]_ ;
  assign \new_[13115]_  = ~\new_[15423]_  | ~\new_[16859]_ ;
  assign \new_[13116]_  = ~\new_[17113]_  | ~\new_[15388]_ ;
  assign \new_[13117]_  = ~\new_[13666]_ ;
  assign \new_[13118]_  = ~\new_[18809]_  & ~\new_[15608]_ ;
  assign \new_[13119]_  = ~\new_[17778]_  | ~\new_[15523]_ ;
  assign \new_[13120]_  = ~\new_[17205]_  & ~\new_[19013]_ ;
  assign \new_[13121]_  = ~\new_[14207]_ ;
  assign \new_[13122]_  = ~\new_[15209]_  | ~\new_[18637]_ ;
  assign \new_[13123]_  = \new_[18914]_  | \new_[15622]_ ;
  assign \new_[13124]_  = ~\new_[13638]_ ;
  assign \new_[13125]_  = ~\new_[15566]_  & ~\new_[15625]_ ;
  assign \new_[13126]_  = ~\new_[14746]_  | ~\new_[16270]_ ;
  assign \new_[13127]_  = ~\new_[17880]_  | ~\new_[15523]_ ;
  assign \new_[13128]_  = ~\new_[14703]_  | ~\new_[15453]_ ;
  assign \new_[13129]_  = ~\new_[16797]_  | ~\new_[15412]_ ;
  assign \new_[13130]_  = \new_[18214]_  | \new_[19874]_ ;
  assign \new_[13131]_  = ~\new_[17039]_  | ~\new_[19253]_ ;
  assign \new_[13132]_  = ~\new_[14836]_  & ~\new_[17615]_ ;
  assign \new_[13133]_  = ~\new_[13615]_ ;
  assign \new_[13134]_  = \new_[17725]_  | \new_[14826]_ ;
  assign \new_[13135]_  = ~\new_[18099]_  | ~\new_[15778]_ ;
  assign \new_[13136]_  = \new_[15810]_  & \new_[18967]_ ;
  assign \new_[13137]_  = ~\new_[19754]_  & ~\new_[16686]_ ;
  assign \new_[13138]_  = ~\new_[14289]_ ;
  assign \new_[13139]_  = ~\new_[14267]_ ;
  assign \new_[13140]_  = ~\new_[13926]_ ;
  assign \new_[13141]_  = \new_[15641]_  | \new_[16987]_ ;
  assign \new_[13142]_  = ~\new_[21328]_  & ~\new_[16947]_ ;
  assign \new_[13143]_  = \new_[18032]_  | \new_[14860]_ ;
  assign \new_[13144]_  = \new_[17570]_  | \new_[15530]_ ;
  assign \new_[13145]_  = \new_[18372]_  | \new_[15466]_ ;
  assign \new_[13146]_  = ~\new_[18023]_  | ~\new_[15417]_ ;
  assign \new_[13147]_  = \new_[15519]_  | \new_[19202]_ ;
  assign \new_[13148]_  = ~\new_[18440]_  & ~\new_[15428]_ ;
  assign \new_[13149]_  = ~\new_[14270]_ ;
  assign \new_[13150]_  = ~\new_[17325]_  | ~\new_[15417]_ ;
  assign \new_[13151]_  = ~\new_[13562]_ ;
  assign \new_[13152]_  = ~\new_[13522]_ ;
  assign \new_[13153]_  = ~\new_[17895]_  | ~\new_[14955]_ ;
  assign \new_[13154]_  = ~\new_[19431]_  & ~\new_[15475]_ ;
  assign \new_[13155]_  = ~\new_[14275]_ ;
  assign \new_[13156]_  = \new_[15572]_  | \new_[19095]_ ;
  assign \new_[13157]_  = ~\new_[13534]_ ;
  assign \new_[13158]_  = ~\new_[14277]_ ;
  assign \new_[13159]_  = ~\new_[14278]_ ;
  assign \new_[13160]_  = ~\new_[17067]_  & ~\new_[18974]_ ;
  assign \new_[13161]_  = ~\new_[13527]_ ;
  assign \new_[13162]_  = ~\new_[17329]_  | ~\new_[15573]_ ;
  assign \new_[13163]_  = \new_[15599]_  | \new_[18731]_ ;
  assign \new_[13164]_  = ~\new_[14282]_ ;
  assign \new_[13165]_  = ~\new_[18086]_  | ~\new_[14838]_ ;
  assign \new_[13166]_  = ~\new_[16985]_  | ~\new_[16891]_ ;
  assign \new_[13167]_  = ~\new_[21327]_ ;
  assign \new_[13168]_  = ~\new_[14718]_  | ~\new_[21558]_ ;
  assign \new_[13169]_  = ~\new_[13495]_ ;
  assign \new_[13170]_  = ~\new_[15487]_  | ~\new_[19098]_ ;
  assign \new_[13171]_  = ~\new_[16799]_  | ~\new_[19021]_ ;
  assign \new_[13172]_  = \new_[16161]_  | \new_[15420]_ ;
  assign \new_[13173]_  = ~\new_[15838]_ ;
  assign \new_[13174]_  = ~\new_[15521]_  | ~\new_[19107]_ ;
  assign \new_[13175]_  = ~\new_[14295]_ ;
  assign \new_[13176]_  = ~\new_[14288]_ ;
  assign \new_[13177]_  = ~\new_[14298]_ ;
  assign \new_[13178]_  = ~\new_[14627]_ ;
  assign \new_[13179]_  = ~\new_[14617]_ ;
  assign \new_[13180]_  = \new_[17784]_  | \new_[15530]_ ;
  assign \new_[13181]_  = ~\new_[14609]_ ;
  assign \new_[13182]_  = ~\new_[15400]_  | ~\new_[16683]_ ;
  assign \new_[13183]_  = ~\new_[15435]_  | ~\new_[18957]_ ;
  assign \new_[13184]_  = ~\new_[18855]_  | ~\new_[16894]_ ;
  assign \new_[13185]_  = ~\new_[15399]_  & ~\new_[18124]_ ;
  assign \new_[13186]_  = ~\new_[14305]_ ;
  assign \new_[13187]_  = ~\new_[14306]_ ;
  assign \new_[13188]_  = ~\new_[14308]_ ;
  assign \new_[13189]_  = ~\new_[14310]_ ;
  assign \new_[13190]_  = \new_[15573]_  | \new_[19084]_ ;
  assign \new_[13191]_  = ~\new_[18576]_  | ~\new_[14955]_ ;
  assign \new_[13192]_  = \new_[17754]_  | \new_[14865]_ ;
  assign \new_[13193]_  = ~\new_[15170]_  | ~\new_[18909]_ ;
  assign \new_[13194]_  = \new_[17341]_  | \new_[18994]_ ;
  assign \new_[13195]_  = ~\new_[16958]_  | ~\new_[17171]_ ;
  assign \new_[13196]_  = ~\new_[14392]_ ;
  assign \new_[13197]_  = ~\new_[16945]_  & ~\new_[18046]_ ;
  assign \new_[13198]_  = ~\new_[14367]_ ;
  assign \new_[13199]_  = ~\new_[14343]_ ;
  assign \new_[13200]_  = ~\new_[14021]_ ;
  assign \new_[13201]_  = ~\new_[17846]_  | ~\new_[14955]_ ;
  assign \new_[13202]_  = ~\new_[15491]_  | ~\new_[18616]_ ;
  assign \new_[13203]_  = ~\new_[14314]_ ;
  assign \new_[13204]_  = ~\new_[14317]_ ;
  assign \new_[13205]_  = ~\new_[15153]_  & ~\new_[21506]_ ;
  assign \new_[13206]_  = ~\new_[18574]_  | ~\new_[14955]_ ;
  assign \new_[13207]_  = ~\new_[14129]_ ;
  assign \new_[13208]_  = ~\new_[16562]_  | ~\new_[18046]_ ;
  assign \new_[13209]_  = ~\new_[18155]_  | ~\new_[14955]_ ;
  assign \new_[13210]_  = ~\new_[16532]_  | ~\new_[15509]_ ;
  assign \new_[13211]_  = \new_[15428]_  | \new_[21495]_ ;
  assign \new_[13212]_  = ~\new_[13644]_ ;
  assign \new_[13213]_  = ~\new_[17710]_  | ~\new_[14847]_ ;
  assign \new_[13214]_  = \new_[18066]_  | \new_[15510]_ ;
  assign \new_[13215]_  = ~\new_[16855]_  & ~\new_[18984]_ ;
  assign \new_[13216]_  = \new_[15053]_  | \new_[18153]_ ;
  assign \new_[13217]_  = ~\new_[17461]_  | ~\new_[14731]_ ;
  assign \new_[13218]_  = ~\new_[19431]_  & (~\new_[17955]_  | ~\new_[16093]_ );
  assign \new_[13219]_  = \new_[14807]_  | \new_[17812]_ ;
  assign \new_[13220]_  = ~\new_[15576]_  & ~\new_[18709]_ ;
  assign \new_[13221]_  = ~\new_[15386]_  & ~\new_[19214]_ ;
  assign \new_[13222]_  = ~\new_[14323]_ ;
  assign \new_[13223]_  = ~\new_[15580]_  & ~\new_[19247]_ ;
  assign \new_[13224]_  = ~\new_[15351]_  & ~\new_[21688]_ ;
  assign \new_[13225]_  = ~\new_[15209]_  | ~\new_[18337]_ ;
  assign \new_[13226]_  = ~\new_[13947]_ ;
  assign \new_[13227]_  = ~\new_[15466]_  & ~\new_[18948]_ ;
  assign \new_[13228]_  = ~\new_[15430]_  | ~\new_[18031]_ ;
  assign \new_[13229]_  = ~\new_[17889]_  | ~\new_[15523]_ ;
  assign \new_[13230]_  = ~\new_[15511]_  & ~\new_[18984]_ ;
  assign \new_[13231]_  = \new_[18058]_  | \new_[19874]_ ;
  assign \new_[13232]_  = \new_[17067]_  | \new_[18062]_ ;
  assign \new_[13233]_  = ~\new_[13844]_ ;
  assign \new_[13234]_  = ~\new_[16747]_  | ~\new_[15545]_ ;
  assign \new_[13235]_  = \new_[15628]_  | \new_[21686]_ ;
  assign \new_[13236]_  = ~\new_[14341]_ ;
  assign \new_[13237]_  = ~\new_[13777]_ ;
  assign \new_[13238]_  = ~\new_[14824]_  | ~\new_[21328]_ ;
  assign \new_[13239]_  = \new_[15574]_  | \new_[19636]_ ;
  assign \new_[13240]_  = ~\new_[15628]_  | ~\new_[21693]_ ;
  assign \new_[13241]_  = ~\new_[15629]_  | ~\new_[21513]_ ;
  assign \new_[13242]_  = ~\new_[15446]_  & ~\new_[19444]_ ;
  assign \new_[13243]_  = \new_[18064]_  | \new_[19874]_ ;
  assign \new_[13244]_  = ~\new_[15425]_  | ~\new_[16291]_ ;
  assign \new_[13245]_  = ~\new_[15209]_  | ~\new_[19154]_ ;
  assign \new_[13246]_  = \new_[15386]_  | \new_[21562]_ ;
  assign \new_[13247]_  = ~\new_[14346]_ ;
  assign \new_[13248]_  = ~\new_[15710]_  | ~\new_[16332]_ ;
  assign \new_[13249]_  = ~\new_[16812]_  | ~\new_[14955]_ ;
  assign \new_[13250]_  = ~\new_[15409]_  & ~\new_[21686]_ ;
  assign \new_[13251]_  = ~\new_[17307]_  & ~\new_[19428]_ ;
  assign \new_[13252]_  = \new_[17258]_  | \new_[19188]_ ;
  assign \new_[13253]_  = ~\new_[15666]_  | ~\new_[19474]_ ;
  assign \new_[13254]_  = ~\new_[21692]_  & ~\new_[12075]_ ;
  assign \new_[13255]_  = \new_[18677]_  | \new_[19874]_ ;
  assign \new_[13256]_  = \new_[15529]_  | \new_[19156]_ ;
  assign \new_[13257]_  = ~\new_[15656]_  & ~\new_[19409]_ ;
  assign \new_[13258]_  = \new_[15771]_  | \new_[15530]_ ;
  assign \new_[13259]_  = ~\new_[14706]_  | ~\new_[18017]_ ;
  assign \new_[13260]_  = ~\new_[13640]_ ;
  assign \new_[13261]_  = ~\new_[14356]_ ;
  assign \new_[13262]_  = ~\new_[17318]_  | ~\new_[15777]_ ;
  assign \new_[13263]_  = ~\new_[13663]_ ;
  assign \new_[13264]_  = \new_[16083]_  | \new_[19874]_ ;
  assign \new_[13265]_  = \new_[17225]_  | \new_[18559]_ ;
  assign \new_[13266]_  = ~\new_[17993]_  & ~\new_[14860]_ ;
  assign \new_[13267]_  = ~\new_[14933]_  | ~\new_[16296]_ ;
  assign \new_[13268]_  = ~\new_[14361]_ ;
  assign \new_[13269]_  = \new_[15727]_  | \new_[18285]_ ;
  assign \new_[13270]_  = ~\new_[17168]_  | ~\new_[18166]_ ;
  assign \new_[13271]_  = ~\new_[14363]_ ;
  assign \new_[13272]_  = ~\new_[14365]_ ;
  assign \new_[13273]_  = ~\new_[13645]_ ;
  assign \new_[13274]_  = ~\new_[13526]_ ;
  assign \new_[13275]_  = ~\new_[18178]_  | ~\new_[15777]_ ;
  assign \new_[13276]_  = \new_[17181]_  & \new_[15020]_ ;
  assign \new_[13277]_  = ~\new_[15153]_  & ~\new_[16879]_ ;
  assign \new_[13278]_  = ~\new_[14371]_ ;
  assign \new_[13279]_  = \new_[15997]_  & \new_[15462]_ ;
  assign \new_[13280]_  = ~\new_[13622]_ ;
  assign \new_[13281]_  = ~\new_[18175]_  | ~\new_[15502]_ ;
  assign \new_[13282]_  = ~\new_[13621]_ ;
  assign \new_[13283]_  = ~\new_[18434]_  | ~\new_[15521]_ ;
  assign \new_[13284]_  = ~\new_[14375]_ ;
  assign \new_[13285]_  = ~\new_[13611]_ ;
  assign \new_[13286]_  = ~\new_[13613]_ ;
  assign \new_[13287]_  = ~\new_[21701]_  & ~\new_[19095]_ ;
  assign \new_[13288]_  = \new_[17910]_  | \new_[19874]_ ;
  assign \new_[13289]_  = ~\new_[13816]_ ;
  assign \new_[13290]_  = ~\new_[17814]_  | ~\new_[15778]_ ;
  assign \new_[13291]_  = ~\new_[14380]_ ;
  assign \new_[13292]_  = ~\new_[14383]_ ;
  assign \new_[13293]_  = ~\new_[14172]_ ;
  assign \new_[13294]_  = ~\new_[15370]_ ;
  assign \new_[13295]_  = \new_[18437]_  | \new_[15530]_ ;
  assign \new_[13296]_  = ~\new_[15543]_  & ~\new_[16381]_ ;
  assign \new_[13297]_  = ~\new_[15787]_  & ~\new_[19084]_ ;
  assign \new_[13298]_  = ~\new_[15659]_  & (~\new_[17934]_  | ~\new_[19117]_ );
  assign \new_[13299]_  = \new_[20664]_  | \new_[19261]_ ;
  assign \new_[13300]_  = \new_[18359]_  | \new_[19874]_ ;
  assign \new_[13301]_  = ~\new_[18039]_  | ~\new_[15778]_ ;
  assign \new_[13302]_  = \new_[18992]_  | \new_[15811]_ ;
  assign \new_[13303]_  = \new_[16859]_  | \new_[18358]_ ;
  assign \new_[13304]_  = \new_[14864]_  | \new_[18012]_ ;
  assign \new_[13305]_  = ~\new_[17811]_  | ~\new_[14955]_ ;
  assign \new_[13306]_  = ~\new_[16076]_  | ~\new_[21306]_ ;
  assign \new_[13307]_  = ~\new_[16424]_  | ~\new_[21669]_ ;
  assign \new_[13308]_  = ~\new_[16409]_  | ~\new_[14916]_ ;
  assign \new_[13309]_  = ~\new_[14397]_ ;
  assign \new_[13310]_  = ~\new_[18117]_  & ~\new_[15464]_ ;
  assign \new_[13311]_  = \new_[17104]_  | \new_[21693]_ ;
  assign \new_[13312]_  = ~\new_[15089]_  | ~\new_[16828]_ ;
  assign \new_[13313]_  = ~\new_[13502]_ ;
  assign \new_[13314]_  = ~\new_[18751]_  & ~\new_[15145]_ ;
  assign \new_[13315]_  = ~\new_[14400]_ ;
  assign \new_[13316]_  = \new_[17500]_  | \new_[15530]_ ;
  assign \new_[13317]_  = ~\new_[18783]_  | ~\new_[16929]_ ;
  assign \new_[13318]_  = ~\new_[15743]_  | ~\new_[19021]_ ;
  assign \new_[13319]_  = ~\new_[17357]_  | ~\new_[15412]_ ;
  assign \new_[13320]_  = \new_[18395]_  | \new_[15530]_ ;
  assign \new_[13321]_  = ~\new_[16799]_  | ~\new_[19413]_ ;
  assign \new_[13322]_  = \new_[17327]_  | \new_[15740]_ ;
  assign \new_[13323]_  = \new_[15518]_  | \new_[16640]_ ;
  assign \new_[13324]_  = ~\new_[16409]_  | (~\new_[16850]_  & ~\new_[19081]_ );
  assign \new_[13325]_  = ~\new_[16520]_  | (~\new_[15977]_  & ~\new_[21520]_ );
  assign \new_[13326]_  = ~\new_[18133]_  | ~\new_[15737]_ ;
  assign \new_[13327]_  = ~\new_[18275]_  | ~\new_[15731]_ ;
  assign \new_[13328]_  = \new_[15528]_  | \new_[14745]_ ;
  assign \new_[13329]_  = ~\new_[18237]_  & (~\new_[16836]_  | ~\new_[16630]_ );
  assign \new_[13330]_  = ~\new_[17929]_  & (~\new_[16021]_  | ~\new_[17848]_ );
  assign \new_[13331]_  = ~\new_[17791]_  & (~\new_[16747]_  | ~\new_[16012]_ );
  assign \new_[13332]_  = ~\new_[14858]_  & (~\new_[17347]_  | ~\new_[18717]_ );
  assign \new_[13333]_  = ~\new_[17259]_  & (~\new_[17334]_  | ~\new_[17970]_ );
  assign \new_[13334]_  = ~\new_[15584]_  | (~\new_[19801]_  & ~\new_[18596]_ );
  assign \new_[13335]_  = ~\new_[18936]_  & (~\new_[21641]_  | ~\new_[17992]_ );
  assign \new_[13336]_  = ~\new_[15616]_  & (~\new_[18080]_  | ~\new_[17471]_ );
  assign \new_[13337]_  = ~\new_[15583]_  & (~\new_[19184]_  | ~\new_[18906]_ );
  assign \new_[13338]_  = ~\new_[17948]_  | ~\new_[17141]_ ;
  assign \new_[13339]_  = ~\new_[15507]_  & (~\new_[21396]_  | ~\new_[16690]_ );
  assign \new_[13340]_  = ~\new_[15707]_  & (~\new_[19044]_  | ~\new_[18477]_ );
  assign \new_[13341]_  = ~\new_[15465]_  & (~\new_[18794]_  | ~\new_[18327]_ );
  assign \new_[13342]_  = \new_[18151]_  | \new_[16879]_ ;
  assign \new_[13343]_  = ~\new_[14013]_ ;
  assign \new_[13344]_  = ~\new_[14428]_ ;
  assign \new_[13345]_  = ~\new_[14430]_ ;
  assign \new_[13346]_  = ~\new_[18335]_  & ~\new_[15653]_ ;
  assign \new_[13347]_  = ~\new_[13600]_ ;
  assign \new_[13348]_  = ~\new_[13662]_ ;
  assign \new_[13349]_  = ~\new_[14437]_ ;
  assign \new_[13350]_  = ~\new_[13651]_ ;
  assign \new_[13351]_  = \new_[14850]_  | \new_[17394]_ ;
  assign \new_[13352]_  = ~\new_[16741]_  | ~\new_[15722]_ ;
  assign \new_[13353]_  = ~\new_[15126]_  | ~\new_[18111]_ ;
  assign \new_[13354]_  = ~\new_[16636]_  | ~\new_[15767]_ ;
  assign \new_[13355]_  = ~\new_[20869]_  & ~\new_[15478]_ ;
  assign \new_[13356]_  = ~\new_[14596]_ ;
  assign \new_[13357]_  = ~\new_[15085]_  | ~\new_[19014]_ ;
  assign \new_[13358]_  = ~\new_[14445]_ ;
  assign \new_[13359]_  = ~\new_[15521]_  | ~\new_[18008]_ ;
  assign \new_[13360]_  = \new_[18128]_  | \new_[19253]_ ;
  assign \new_[13361]_  = ~\new_[14188]_ ;
  assign \new_[13362]_  = ~\new_[13763]_ ;
  assign \new_[13363]_  = ~\new_[14454]_ ;
  assign \new_[13364]_  = ~\new_[14189]_ ;
  assign \new_[13365]_  = ~\new_[14830]_  | ~\new_[18747]_ ;
  assign \new_[13366]_  = ~\new_[14953]_  | ~\new_[18605]_ ;
  assign \new_[13367]_  = ~\new_[14461]_ ;
  assign \new_[13368]_  = ~\new_[14727]_  & ~\new_[18794]_ ;
  assign \new_[13369]_  = ~\new_[14662]_ ;
  assign \new_[13370]_  = ~\new_[14466]_ ;
  assign \new_[13371]_  = \new_[16813]_  | \new_[17886]_ ;
  assign \new_[13372]_  = ~\new_[18605]_  & ~\new_[17354]_ ;
  assign \new_[13373]_  = ~\new_[14934]_  & ~\new_[21695]_ ;
  assign \new_[13374]_  = ~\new_[14469]_ ;
  assign \new_[13375]_  = ~\new_[14469]_ ;
  assign \new_[13376]_  = ~\new_[14233]_ ;
  assign \new_[13377]_  = ~\new_[16598]_  & ~\new_[15795]_ ;
  assign \new_[13378]_  = ~\new_[16095]_ ;
  assign \new_[13379]_  = ~\new_[14816]_  | ~\new_[21569]_ ;
  assign \new_[13380]_  = ~\new_[13649]_ ;
  assign \new_[13381]_  = ~\new_[14692]_  & ~\new_[18709]_ ;
  assign \new_[13382]_  = ~\new_[15809]_  | ~\new_[17598]_ ;
  assign \new_[13383]_  = ~\new_[15792]_  | ~\new_[18443]_ ;
  assign \new_[13384]_  = ~\new_[14783]_  | ~\new_[19102]_ ;
  assign \new_[13385]_  = ~\new_[13559]_ ;
  assign \new_[13386]_  = ~\new_[14718]_  | ~\new_[21396]_ ;
  assign \new_[13387]_  = \new_[15818]_  | \new_[21569]_ ;
  assign \new_[13388]_  = ~\new_[14495]_ ;
  assign \new_[13389]_  = ~\new_[15801]_  & ~\new_[18888]_ ;
  assign \new_[13390]_  = ~\new_[14503]_ ;
  assign \new_[13391]_  = ~\new_[13996]_ ;
  assign \new_[13392]_  = ~\new_[17862]_  & (~\new_[17295]_  | ~\new_[16604]_ );
  assign \new_[13393]_  = \new_[14685]_ ;
  assign \new_[13394]_  = ~\new_[14683]_ ;
  assign \new_[13395]_  = ~\new_[16470]_  | ~\new_[18926]_ ;
  assign \new_[13396]_  = \new_[17063]_  | \new_[18151]_ ;
  assign \new_[13397]_  = ~\new_[14665]_ ;
  assign \new_[13398]_  = ~\new_[14606]_ ;
  assign \new_[13399]_  = ~\new_[14516]_ ;
  assign \new_[13400]_  = ~\new_[14422]_ ;
  assign \new_[13401]_  = ~\new_[13778]_ ;
  assign \new_[13402]_  = ~\new_[15534]_  & ~\new_[21635]_ ;
  assign \new_[13403]_  = \new_[17123]_  | \new_[15727]_ ;
  assign \new_[13404]_  = ~\new_[13538]_ ;
  assign \new_[13405]_  = \new_[15826]_  | \new_[18012]_ ;
  assign \new_[13406]_  = ~\new_[15809]_  | ~\new_[19711]_ ;
  assign \new_[13407]_  = ~\new_[13506]_ ;
  assign \new_[13408]_  = ~\new_[15821]_  & ~\new_[21689]_ ;
  assign \new_[13409]_  = ~\new_[14699]_  | ~\new_[19589]_ ;
  assign \new_[13410]_  = ~\new_[13489]_ ;
  assign \new_[13411]_  = ~\new_[13486]_ ;
  assign \new_[13412]_  = ~\new_[14789]_  & ~\new_[18423]_ ;
  assign \new_[13413]_  = ~\new_[17345]_  | ~\new_[18427]_ ;
  assign \new_[13414]_  = ~\new_[14644]_ ;
  assign \new_[13415]_  = ~\new_[14556]_ ;
  assign \new_[13416]_  = ~\new_[21300]_ ;
  assign \new_[13417]_  = \new_[15796]_  | \new_[19270]_ ;
  assign \new_[13418]_  = ~\new_[14221]_ ;
  assign \new_[13419]_  = ~\new_[14716]_  | ~\new_[19098]_ ;
  assign \new_[13420]_  = ~\new_[14830]_  | ~\new_[21562]_ ;
  assign \new_[13421]_  = ~\new_[13580]_ ;
  assign \new_[13422]_  = ~\new_[21541]_  | ~\new_[19064]_  | ~\new_[17529]_ ;
  assign \new_[13423]_  = \new_[15124]_  | \new_[17843]_ ;
  assign \new_[13424]_  = ~\new_[13488]_ ;
  assign \new_[13425]_  = ~\new_[14691]_ ;
  assign \new_[13426]_  = ~\new_[14585]_ ;
  assign \new_[13427]_  = ~\new_[14675]_ ;
  assign \new_[13428]_  = ~\new_[14652]_ ;
  assign \new_[13429]_  = ~\new_[14587]_ ;
  assign \new_[13430]_  = ~\new_[19260]_  | ~\new_[15795]_ ;
  assign \new_[13431]_  = ~\new_[15970]_ ;
  assign \new_[13432]_  = ~\new_[17426]_  | ~\new_[18652]_ ;
  assign \new_[13433]_  = ~\new_[13548]_ ;
  assign \new_[13434]_  = ~\new_[17016]_  | ~\new_[19085]_ ;
  assign \new_[13435]_  = ~\new_[14169]_ ;
  assign \new_[13436]_  = ~\new_[17699]_  & ~\new_[17593]_ ;
  assign \new_[13437]_  = ~\new_[14601]_ ;
  assign \new_[13438]_  = ~\new_[16700]_  & ~\new_[17630]_ ;
  assign \new_[13439]_  = ~\new_[17594]_  | ~\new_[14783]_ ;
  assign \new_[13440]_  = ~\new_[18518]_  | ~\new_[17560]_ ;
  assign \new_[13441]_  = ~\new_[17380]_  | ~\new_[15767]_ ;
  assign \new_[13442]_  = ~\new_[14285]_ ;
  assign \new_[13443]_  = ~\new_[17361]_  & ~\new_[16976]_ ;
  assign \new_[13444]_  = ~\new_[16730]_  | ~\new_[16846]_ ;
  assign \new_[13445]_  = ~\new_[16596]_  & ~\new_[14940]_ ;
  assign \new_[13446]_  = ~\new_[17105]_  | (~\new_[17886]_  & ~\new_[18801]_ );
  assign \new_[13447]_  = ~\new_[14611]_ ;
  assign \new_[13448]_  = \new_[16859]_  | \new_[21688]_ ;
  assign \new_[13449]_  = ~\new_[19027]_  & ~\new_[15632]_ ;
  assign \new_[13450]_  = \new_[15842]_  ^ \new_[17553]_ ;
  assign \new_[13451]_  = ~\new_[17886]_  & ~\new_[15804]_ ;
  assign \new_[13452]_  = \new_[19705]_  ^ \new_[18391]_ ;
  assign \new_[13453]_  = \new_[14758]_  ^ \new_[18757]_ ;
  assign \new_[13454]_  = ~\new_[13976]_ ;
  assign \new_[13455]_  = \new_[14764]_  ^ \new_[17484]_ ;
  assign \new_[13456]_  = \new_[19763]_  ^ \new_[19578]_ ;
  assign \new_[13457]_  = ~\new_[20164]_ ;
  assign \new_[13458]_  = \new_[14756]_  ^ \new_[19184]_ ;
  assign \new_[13459]_  = \new_[19646]_  ^ \new_[18449]_ ;
  assign \new_[13460]_  = \new_[19634]_  ^ \new_[18877]_ ;
  assign \new_[13461]_  = ~\new_[21301]_  & ~\new_[16729]_ ;
  assign \new_[13462]_  = ~\new_[14791]_  & ~\new_[19535]_ ;
  assign \new_[13463]_  = ~\new_[14294]_ ;
  assign \new_[13464]_  = ~\new_[14661]_ ;
  assign \new_[13465]_  = ~\new_[14970]_  & ~\new_[18794]_ ;
  assign \new_[13466]_  = \new_[18208]_  | \new_[15315]_ ;
  assign \new_[13467]_  = ~\new_[13972]_ ;
  assign \new_[13468]_  = ~\new_[15775]_  | ~\new_[19100]_ ;
  assign \new_[13469]_  = \new_[15791]_  | \new_[21396]_ ;
  assign \new_[13470]_  = ~\new_[14859]_  & ~\new_[19019]_ ;
  assign \new_[13471]_  = ~\new_[17241]_  & (~\new_[16844]_  | ~\new_[16553]_ );
  assign \new_[13472]_  = ~\new_[13967]_ ;
  assign \new_[13473]_  = ~\new_[21607]_  & ~\new_[19082]_ ;
  assign \new_[13474]_  = \new_[19780]_  & \new_[18414]_ ;
  assign \new_[13475]_  = ~\new_[18715]_  | ~\new_[14787]_ ;
  assign n2738 = \new_[15807]_  & \new_[14787]_ ;
  assign \new_[13477]_  = ~\new_[13568]_ ;
  assign \new_[13478]_  = ~\new_[15767]_  & ~\new_[19179]_ ;
  assign \new_[13479]_  = ~\new_[14457]_ ;
  assign n2733 = \new_[16667]_  & \new_[14787]_ ;
  assign \new_[13481]_  = ~\new_[17642]_  | ~\new_[15523]_ ;
  assign \new_[13482]_  = ~\new_[15506]_  | (~\new_[15977]_  & ~\new_[21541]_ );
  assign \new_[13483]_  = ~\new_[14691]_ ;
  assign \new_[13484]_  = ~\new_[19444]_  | ~\new_[19084]_  | ~\new_[17271]_ ;
  assign \new_[13485]_  = ~\new_[14692]_ ;
  assign \new_[13486]_  = ~\new_[15606]_ ;
  assign \new_[13487]_  = ~\new_[16262]_  & ~\new_[18766]_ ;
  assign \new_[13488]_  = ~\new_[16486]_ ;
  assign \new_[13489]_  = ~\new_[14705]_ ;
  assign \new_[13490]_  = ~\new_[21652]_  | ~\new_[21685]_ ;
  assign \new_[13491]_  = ~\new_[16681]_  | ~\new_[19181]_ ;
  assign \new_[13492]_  = ~\new_[14718]_ ;
  assign \new_[13493]_  = ~\new_[17666]_  & ~\new_[17743]_ ;
  assign \new_[13494]_  = ~\new_[16321]_  | ~\new_[19018]_ ;
  assign \new_[13495]_  = ~\new_[19024]_  & (~\new_[17921]_  | ~\new_[18141]_ );
  assign \new_[13496]_  = ~\new_[18981]_  | ~\new_[16275]_ ;
  assign \new_[13497]_  = ~\new_[16730]_  | ~\new_[16045]_ ;
  assign \new_[13498]_  = ~\new_[15533]_ ;
  assign \new_[13499]_  = \new_[16249]_  | \new_[19409]_ ;
  assign \new_[13500]_  = ~\new_[17886]_  & ~\new_[19539]_  & ~\new_[17391]_ ;
  assign \new_[13501]_  = ~\new_[16386]_  | ~\new_[19409]_ ;
  assign \new_[13502]_  = ~\new_[17481]_  & ~\new_[18083]_ ;
  assign \new_[13503]_  = ~\new_[16853]_  | ~\new_[16468]_ ;
  assign \new_[13504]_  = ~\new_[14738]_ ;
  assign \new_[13505]_  = ~\new_[16325]_  | ~\new_[18979]_ ;
  assign \new_[13506]_  = ~\new_[15603]_ ;
  assign \new_[13507]_  = \new_[16005]_  & \new_[19409]_ ;
  assign \new_[13508]_  = ~\new_[14740]_ ;
  assign \new_[13509]_  = ~\new_[15226]_ ;
  assign \new_[13510]_  = ~\new_[14747]_ ;
  assign \new_[13511]_  = ~\new_[16209]_  | ~\new_[21506]_ ;
  assign \new_[13512]_  = ~\new_[15109]_ ;
  assign \new_[13513]_  = \new_[16498]_  & \new_[16272]_ ;
  assign \new_[13514]_  = ~\new_[14757]_ ;
  assign done = done_reg;
  assign \new_[13516]_  = ~\new_[15375]_ ;
  assign \new_[13517]_  = ~\new_[18307]_  | ~\new_[16610]_  | ~\new_[18113]_ ;
  assign \new_[13518]_  = ~\new_[15783]_ ;
  assign n2758 = ~\new_[16610]_  & ~n3423;
  assign \new_[13520]_  = ~\new_[14843]_ ;
  assign \new_[13521]_  = ~\new_[16696]_  & (~\new_[18323]_  | ~\new_[18144]_ );
  assign \new_[13522]_  = ~\new_[18319]_  | ~\new_[16661]_ ;
  assign \new_[13523]_  = ~\new_[15599]_ ;
  assign \new_[13524]_  = ~\new_[16490]_  & ~\new_[19196]_ ;
  assign \new_[13525]_  = ~\new_[17114]_ ;
  assign \new_[13526]_  = ~\new_[14796]_ ;
  assign \new_[13527]_  = ~\new_[15321]_ ;
  assign \new_[13528]_  = ~\new_[14806]_ ;
  assign \new_[13529]_  = ~\new_[14807]_ ;
  assign \new_[13530]_  = ~\new_[20291]_ ;
  assign \new_[13531]_  = ~\new_[17607]_  | ~\new_[18747]_ ;
  assign \new_[13532]_  = ~\new_[15344]_ ;
  assign \new_[13533]_  = ~\new_[14969]_ ;
  assign \new_[13534]_  = ~\new_[16620]_  & ~\new_[18006]_ ;
  assign \new_[13535]_  = ~\new_[18909]_  | ~\new_[17853]_ ;
  assign \new_[13536]_  = ~\new_[14818]_ ;
  assign \new_[13537]_  = ~\new_[17764]_  | ~\new_[18577]_ ;
  assign \new_[13538]_  = ~\new_[14818]_ ;
  assign \new_[13539]_  = ~\new_[16652]_  | ~\new_[19019]_ ;
  assign \new_[13540]_  = \new_[18245]_  & \new_[19033]_ ;
  assign \new_[13541]_  = ~\new_[16086]_  & ~\new_[21496]_ ;
  assign \new_[13542]_  = \new_[19560]_  ^ \new_[14690]_ ;
  assign \new_[13543]_  = ~\new_[20489]_  | ~\new_[18427]_ ;
  assign \new_[13544]_  = ~\new_[16923]_  | ~\new_[16040]_  | ~\new_[17543]_ ;
  assign \new_[13545]_  = ~\new_[14840]_ ;
  assign \new_[13546]_  = ~\new_[17529]_  | ~\new_[19036]_  | ~\new_[20867]_ ;
  assign \new_[13547]_  = ~\new_[16506]_  | ~\new_[19409]_ ;
  assign \new_[13548]_  = ~\new_[15656]_ ;
  assign \new_[13549]_  = \new_[17975]_  | \new_[21655]_  | \new_[21693]_  | \new_[19285]_ ;
  assign \new_[13550]_  = ~\new_[14853]_ ;
  assign \new_[13551]_  = ~\new_[15517]_ ;
  assign \new_[13552]_  = \new_[17774]_  | \new_[19603]_  | \new_[18832]_  | \new_[19676]_ ;
  assign \new_[13553]_  = \new_[16669]_  & \new_[19288]_ ;
  assign \new_[13554]_  = ~\new_[18730]_  | ~\new_[19685]_  | ~\new_[19589]_  | ~\new_[19655]_ ;
  assign \new_[13555]_  = ~\new_[15580]_ ;
  assign \new_[13556]_  = ~\new_[15512]_ ;
  assign \new_[13557]_  = \new_[17931]_  | \new_[19087]_  | \new_[19665]_  | \new_[19066]_ ;
  assign \new_[13558]_  = ~\new_[18838]_  | ~\new_[19603]_  | ~\new_[18832]_  | ~\new_[19098]_ ;
  assign \new_[13559]_  = ~\new_[16629]_  & ~\new_[19353]_ ;
  assign \new_[13560]_  = ~\new_[18601]_  | ~\new_[19087]_  | ~\new_[18414]_  | ~\new_[18906]_ ;
  assign \new_[13561]_  = ~\new_[21642]_  | ~\new_[18186]_  | ~\new_[19145]_  | ~\new_[18709]_ ;
  assign \new_[13562]_  = ~\new_[16205]_  | ~\new_[20492]_ ;
  assign \new_[13563]_  = ~\new_[19664]_  | ~\new_[17607]_  | ~\new_[17541]_  | ~\new_[19144]_ ;
  assign \new_[13564]_  = \new_[16269]_  & \new_[19742]_ ;
  assign \new_[13565]_  = ~\new_[15516]_ ;
  assign \new_[13566]_  = ~\new_[16182]_  | ~\new_[18832]_ ;
  assign \new_[13567]_  = ~\new_[14860]_ ;
  assign \new_[13568]_  = ~\new_[14859]_ ;
  assign \new_[13569]_  = ~\new_[18104]_  | ~\new_[21542]_  | ~\new_[20680]_  | ~\new_[19130]_ ;
  assign \new_[13570]_  = \new_[17546]_  & \new_[19754]_ ;
  assign \new_[13571]_  = ~\new_[16676]_  | ~\new_[19335]_ ;
  assign \new_[13572]_  = ~\new_[17765]_  | ~\new_[19116]_  | ~\new_[18542]_  | ~\new_[19444]_ ;
  assign \new_[13573]_  = ~\new_[21622]_  & ~\new_[19431]_ ;
  assign \new_[13574]_  = ~\new_[17686]_  | ~\new_[18881]_  | ~\new_[17457]_  | ~\new_[17843]_ ;
  assign \new_[13575]_  = ~\new_[14866]_ ;
  assign \new_[13576]_  = \new_[16121]_  | \new_[18965]_ ;
  assign \new_[13577]_  = ~\new_[16675]_  & ~\new_[20239]_ ;
  assign \new_[13578]_  = \new_[17465]_  | \new_[19319]_ ;
  assign \new_[13579]_  = ~\new_[15215]_ ;
  assign \new_[13580]_  = ~\new_[16021]_  & ~\new_[19367]_ ;
  assign \new_[13581]_  = ~\new_[20770]_  | ~\new_[19689]_ ;
  assign \new_[13582]_  = ~\new_[17611]_  | ~\new_[21491]_  | ~\new_[19214]_  | ~\new_[18888]_ ;
  assign \new_[13583]_  = ~\new_[15982]_  | ~\new_[18194]_ ;
  assign \new_[13584]_  = \new_[16235]_  | \new_[18766]_ ;
  assign \new_[13585]_  = \new_[17539]_  | \new_[18264]_  | \new_[19687]_  | \new_[19367]_ ;
  assign \new_[13586]_  = ~\new_[15214]_ ;
  assign \new_[13587]_  = ~\new_[16110]_  | ~\new_[19538]_ ;
  assign \new_[13588]_  = ~\new_[15511]_ ;
  assign \new_[13589]_  = ~\new_[16316]_  & ~\new_[18709]_ ;
  assign \new_[13590]_  = ~\new_[16004]_  | ~\new_[18616]_ ;
  assign \new_[13591]_  = ~\new_[17287]_  | ~\new_[16026]_ ;
  assign \new_[13592]_  = ~\new_[15093]_ ;
  assign \new_[13593]_  = ~\new_[16101]_  & ~\new_[18969]_ ;
  assign \new_[13594]_  = ~\new_[15639]_ ;
  assign \new_[13595]_  = ~\new_[19782]_  | ~\new_[19568]_  | ~\new_[17313]_ ;
  assign \new_[13596]_  = ~\new_[18398]_  | ~\new_[17777]_  | ~\new_[18994]_  | ~\new_[19196]_ ;
  assign n2748 = ~\new_[14882]_ ;
  assign \new_[13598]_  = ~\new_[17942]_  | ~\new_[17777]_ ;
  assign \new_[13599]_  = ~\new_[16226]_  & ~\new_[18833]_ ;
  assign \new_[13600]_  = ~\new_[15397]_ ;
  assign \new_[13601]_  = ~\new_[17968]_  | ~\new_[19116]_  | ~\new_[19084]_  | ~\new_[19091]_ ;
  assign \new_[13602]_  = ~\new_[15310]_ ;
  assign \new_[13603]_  = \new_[16353]_  | \new_[19697]_ ;
  assign \new_[13604]_  = ~\new_[17783]_  | ~\new_[21658]_  | ~\new_[21685]_  | ~\new_[21306]_ ;
  assign \new_[13605]_  = ~\new_[14891]_ ;
  assign \new_[13606]_  = \new_[18106]_  | \new_[16617]_ ;
  assign \new_[13607]_  = \new_[17534]_  | \new_[17874]_ ;
  assign \new_[13608]_  = ~\new_[16455]_  & ~\new_[19036]_ ;
  assign \new_[13609]_  = ~\new_[14894]_ ;
  assign \new_[13610]_  = ~\new_[15912]_  | ~\new_[21498]_ ;
  assign \new_[13611]_  = ~\new_[16063]_  & ~\new_[19625]_ ;
  assign \new_[13612]_  = ~\new_[16674]_  | ~\new_[18278]_ ;
  assign \new_[13613]_  = ~\new_[17544]_  | ~\new_[16477]_ ;
  assign \new_[13614]_  = ~\new_[16228]_  & ~\new_[19084]_ ;
  assign \new_[13615]_  = ~\new_[18222]_  | ~\new_[16488]_ ;
  assign \new_[13616]_  = ~\new_[17066]_  | ~\new_[18076]_ ;
  assign \new_[13617]_  = ~\new_[19015]_  & (~\new_[17010]_  | ~\new_[16920]_ );
  assign \new_[13618]_  = \new_[18734]_  | \new_[16406]_ ;
  assign \new_[13619]_  = ~\new_[17326]_  | ~\new_[16320]_  | ~\new_[16712]_ ;
  assign \new_[13620]_  = ~\new_[16198]_  | ~\new_[18832]_ ;
  assign \new_[13621]_  = ~\new_[16583]_  & ~\new_[18061]_ ;
  assign \new_[13622]_  = \new_[16100]_  | \new_[19754]_ ;
  assign \new_[13623]_  = ~\new_[14920]_ ;
  assign \new_[13624]_  = \new_[16462]_  & \new_[19642]_ ;
  assign \new_[13625]_  = ~\new_[14908]_ ;
  assign \new_[13626]_  = ~\new_[16088]_  & ~\new_[19269]_ ;
  assign \new_[13627]_  = ~\new_[16104]_  | ~\new_[19419]_ ;
  assign \new_[13628]_  = ~\new_[16124]_  | ~\new_[17138]_ ;
  assign \new_[13629]_  = ~\new_[18542]_  & (~\new_[16952]_  | ~\new_[17238]_ );
  assign \new_[13630]_  = ~\new_[16253]_  | ~\new_[19203]_ ;
  assign \new_[13631]_  = \new_[16437]_  | \new_[16637]_ ;
  assign \new_[13632]_  = ~\new_[14914]_ ;
  assign \new_[13633]_  = \new_[16253]_  & \new_[19636]_ ;
  assign \new_[13634]_  = ~\new_[14914]_ ;
  assign \new_[13635]_  = ~\new_[19655]_  | ~\new_[17746]_ ;
  assign \new_[13636]_  = ~\new_[15364]_ ;
  assign \new_[13637]_  = \new_[15998]_  | \new_[19145]_ ;
  assign \new_[13638]_  = ~\new_[15889]_  | ~\new_[19664]_ ;
  assign \new_[13639]_  = ~\new_[16128]_  & ~\new_[18682]_ ;
  assign \new_[13640]_  = ~\new_[15349]_ ;
  assign \new_[13641]_  = ~\new_[16238]_  & ~\new_[19024]_ ;
  assign \new_[13642]_  = ~\new_[17066]_  | ~\new_[19008]_ ;
  assign \new_[13643]_  = \new_[16488]_  & \new_[19117]_ ;
  assign \new_[13644]_  = ~\new_[15341]_ ;
  assign \new_[13645]_  = ~\new_[16134]_  | ~\new_[18692]_ ;
  assign \new_[13646]_  = ~\new_[16243]_  & ~\new_[19151]_ ;
  assign \new_[13647]_  = ~\new_[15082]_ ;
  assign \new_[13648]_  = ~\new_[16244]_  | ~\new_[19476]_ ;
  assign \new_[13649]_  = ~\new_[16049]_  | ~\new_[18947]_ ;
  assign \new_[13650]_  = ~\new_[16233]_  & ~\new_[21511]_ ;
  assign \new_[13651]_  = ~\new_[15407]_ ;
  assign \new_[13652]_  = ~\new_[15980]_  | ~\new_[18972]_ ;
  assign \new_[13653]_  = ~\new_[21483]_  | ~\new_[18186]_  | ~\new_[18643]_  | ~\new_[19535]_ ;
  assign \new_[13654]_  = ~\new_[16181]_  | ~\new_[18678]_ ;
  assign \new_[13655]_  = ~\new_[16284]_  | ~\new_[18972]_ ;
  assign \new_[13656]_  = \new_[15914]_  & \new_[19815]_ ;
  assign \new_[13657]_  = ~\new_[18672]_  | ~\new_[17747]_ ;
  assign \new_[13658]_  = ~\new_[15493]_ ;
  assign \new_[13659]_  = ~\new_[17756]_  | ~\new_[15899]_  | ~\new_[18486]_ ;
  assign \new_[13660]_  = ~\new_[15914]_  | ~\new_[18938]_ ;
  assign \new_[13661]_  = \new_[16188]_  | \new_[18187]_ ;
  assign \new_[13662]_  = ~\new_[16428]_  | ~\new_[19454]_ ;
  assign \new_[13663]_  = ~\new_[16423]_  | ~\new_[17886]_ ;
  assign \new_[13664]_  = ~\new_[15076]_ ;
  assign \new_[13665]_  = ~\new_[16180]_  & ~\new_[19269]_ ;
  assign \new_[13666]_  = ~\new_[18116]_  & ~\new_[16734]_ ;
  assign \new_[13667]_  = ~\new_[16069]_  | ~\new_[18414]_ ;
  assign \new_[13668]_  = ~\new_[19754]_  & ~\new_[16583]_ ;
  assign \new_[13669]_  = ~\new_[16372]_  | ~\new_[21500]_ ;
  assign \new_[13670]_  = ~\new_[14946]_ ;
  assign \new_[13671]_  = ~\new_[14954]_ ;
  assign \new_[13672]_  = ~\new_[16082]_  & ~\new_[18083]_ ;
  assign \new_[13673]_  = ~\new_[14969]_ ;
  assign \new_[13674]_  = ~\new_[16706]_  | ~\new_[16192]_ ;
  assign \new_[13675]_  = ~\new_[16055]_  & ~\new_[19446]_ ;
  assign \new_[13676]_  = ~\new_[15073]_ ;
  assign \new_[13677]_  = ~\new_[16587]_  & ~\new_[21693]_ ;
  assign \new_[13678]_  = ~\new_[15490]_ ;
  assign \new_[13679]_  = ~\new_[17076]_  & (~\new_[18250]_  | ~\new_[17655]_ );
  assign \new_[13680]_  = ~\new_[14874]_ ;
  assign \new_[13681]_  = ~\new_[15069]_ ;
  assign \new_[13682]_  = ~\new_[15363]_ ;
  assign \new_[13683]_  = \new_[16368]_  | \new_[18066]_ ;
  assign \new_[13684]_  = ~\new_[18826]_  | ~\new_[16355]_ ;
  assign \new_[13685]_  = ~\new_[16097]_  | ~\new_[17529]_ ;
  assign \new_[13686]_  = ~\new_[17924]_  | (~\new_[17855]_  & ~\new_[17213]_ );
  assign \new_[13687]_  = ~\new_[15297]_ ;
  assign \new_[13688]_  = ~\new_[16203]_  | ~\new_[19091]_ ;
  assign \new_[13689]_  = ~\new_[17337]_  | ~\new_[16417]_ ;
  assign \new_[13690]_  = \new_[17319]_  ^ \new_[18764]_ ;
  assign \new_[13691]_  = ~\new_[16574]_  & ~\new_[19410]_ ;
  assign \new_[13692]_  = ~\new_[17792]_  | ~\new_[16462]_ ;
  assign \new_[13693]_  = ~\new_[16662]_  | ~\new_[18966]_ ;
  assign \new_[13694]_  = ~\new_[14968]_ ;
  assign \new_[13695]_  = ~\new_[14971]_ ;
  assign \new_[13696]_  = ~\new_[15962]_  | ~\new_[18035]_ ;
  assign \new_[13697]_  = ~\new_[14973]_ ;
  assign \new_[13698]_  = ~\new_[14974]_ ;
  assign \new_[13699]_  = \new_[16571]_  & \new_[19474]_ ;
  assign \new_[13700]_  = ~\new_[21045]_  & ~\new_[19409]_ ;
  assign \new_[13701]_  = ~\new_[14975]_ ;
  assign \new_[13702]_  = \new_[14976]_ ;
  assign \new_[13703]_  = ~\new_[21704]_  | ~\new_[18810]_ ;
  assign \new_[13704]_  = ~\new_[15948]_  & ~\new_[18984]_ ;
  assign \new_[13705]_  = ~\new_[14958]_ ;
  assign \new_[13706]_  = ~\new_[15797]_ ;
  assign \new_[13707]_  = ~\new_[14978]_ ;
  assign \new_[13708]_  = \new_[16384]_  & \new_[19431]_ ;
  assign \new_[13709]_  = ~\new_[14979]_ ;
  assign \new_[13710]_  = ~\new_[15994]_  | ~\new_[19031]_ ;
  assign \new_[13711]_  = ~\new_[15790]_ ;
  assign \new_[13712]_  = ~\new_[15391]_ ;
  assign \new_[13713]_  = \new_[16332]_  | \new_[18973]_ ;
  assign \new_[13714]_  = ~\new_[15788]_ ;
  assign \new_[13715]_  = ~\new_[16411]_  | ~\new_[19270]_ ;
  assign \new_[13716]_  = ~\new_[14980]_ ;
  assign \new_[13717]_  = ~\new_[14981]_ ;
  assign \new_[13718]_  = ~\new_[14982]_ ;
  assign \new_[13719]_  = ~\new_[17235]_  | ~\new_[19091]_ ;
  assign \new_[13720]_  = ~\new_[18565]_  | ~\new_[17476]_  | ~\new_[18008]_  | ~\new_[18567]_ ;
  assign \new_[13721]_  = ~\new_[14983]_ ;
  assign \new_[13722]_  = ~\new_[18020]_  & ~\new_[16535]_ ;
  assign \new_[13723]_  = ~\new_[16328]_  | ~\new_[18652]_ ;
  assign \new_[13724]_  = ~\new_[15875]_  | ~\new_[19042]_ ;
  assign \new_[13725]_  = ~\new_[16161]_  | ~\new_[18111]_ ;
  assign \new_[13726]_  = ~\new_[15883]_  | ~\new_[19379]_ ;
  assign \new_[13727]_  = ~\new_[17871]_  | ~\new_[19758]_ ;
  assign \new_[13728]_  = ~\new_[16135]_  | ~\new_[19156]_ ;
  assign \new_[13729]_  = ~\new_[16488]_  | ~\new_[19192]_ ;
  assign \new_[13730]_  = ~\new_[14986]_ ;
  assign \new_[13731]_  = ~\new_[14987]_ ;
  assign \new_[13732]_  = ~\new_[17460]_  & ~\new_[16461]_ ;
  assign \new_[13733]_  = ~\new_[15693]_ ;
  assign \new_[13734]_  = ~\new_[16413]_  & ~\new_[19270]_ ;
  assign \new_[13735]_  = ~\new_[18565]_  | ~\new_[18461]_  | ~\new_[19548]_  | ~\new_[19270]_ ;
  assign \new_[13736]_  = ~\new_[15661]_ ;
  assign \new_[13737]_  = ~\new_[21703]_  | ~\new_[18893]_ ;
  assign \new_[13738]_  = ~\new_[14992]_ ;
  assign \new_[13739]_  = ~\new_[14994]_ ;
  assign \new_[13740]_  = ~\new_[14995]_ ;
  assign \new_[13741]_  = \new_[14997]_ ;
  assign \new_[13742]_  = ~\new_[14999]_ ;
  assign \new_[13743]_  = ~\new_[15350]_ ;
  assign \new_[13744]_  = ~\new_[16410]_  | ~\new_[21511]_ ;
  assign \new_[13745]_  = ~\new_[15564]_ ;
  assign \new_[13746]_  = ~\new_[15000]_ ;
  assign \new_[13747]_  = ~\new_[15557]_ ;
  assign \new_[13748]_  = ~\new_[15948]_  & ~\new_[19450]_ ;
  assign \new_[13749]_  = ~\new_[15001]_ ;
  assign \new_[13750]_  = ~\new_[15004]_ ;
  assign \new_[13751]_  = ~\new_[15005]_ ;
  assign \new_[13752]_  = ~\new_[16489]_  | ~\new_[19202]_ ;
  assign \new_[13753]_  = ~\new_[15006]_ ;
  assign \new_[13754]_  = ~\new_[15008]_ ;
  assign \new_[13755]_  = ~\new_[15009]_ ;
  assign \new_[13756]_  = ~\new_[15485]_ ;
  assign \new_[13757]_  = ~\new_[19061]_  | ~\new_[17607]_  | ~\new_[17541]_  | ~\new_[21492]_ ;
  assign \new_[13758]_  = ~\new_[15477]_ ;
  assign \new_[13759]_  = \new_[16464]_  & \new_[17457]_ ;
  assign \new_[13760]_  = \new_[16531]_  & \new_[19176]_ ;
  assign \new_[13761]_  = \new_[16080]_  & \new_[21697]_ ;
  assign \new_[13762]_  = ~\new_[15015]_ ;
  assign \new_[13763]_  = ~\new_[15951]_  | ~\new_[19192]_ ;
  assign \new_[13764]_  = ~\new_[16489]_  | ~\new_[19196]_ ;
  assign \new_[13765]_  = ~\new_[16647]_  | ~\new_[18414]_ ;
  assign \new_[13766]_  = ~\new_[15972]_  | ~\new_[19335]_ ;
  assign \new_[13767]_  = ~\new_[21552]_  & ~\new_[18166]_ ;
  assign \new_[13768]_  = ~\new_[15016]_ ;
  assign \new_[13769]_  = ~\new_[15415]_ ;
  assign \new_[13770]_  = ~\new_[15017]_ ;
  assign \new_[13771]_  = ~\new_[16172]_  | ~\new_[21684]_ ;
  assign \new_[13772]_  = ~\new_[16123]_  & ~\new_[19268]_ ;
  assign \new_[13773]_  = \new_[16624]_  & \new_[19275]_ ;
  assign \new_[13774]_  = ~\new_[16100]_  & ~\new_[18941]_ ;
  assign \new_[13775]_  = ~\new_[16305]_  | ~\new_[21697]_ ;
  assign \new_[13776]_  = ~\new_[16405]_  | ~\new_[14951]_ ;
  assign \new_[13777]_  = ~\new_[15895]_  & ~\new_[18637]_ ;
  assign \new_[13778]_  = ~\new_[16042]_  & ~\new_[19270]_ ;
  assign \new_[13779]_  = ~\new_[16016]_  | ~\new_[19212]_ ;
  assign \new_[13780]_  = ~\new_[15378]_ ;
  assign \new_[13781]_  = ~\new_[15021]_ ;
  assign \new_[13782]_  = ~\new_[15022]_ ;
  assign \new_[13783]_  = ~\new_[16102]_  | ~\new_[19269]_ ;
  assign \new_[13784]_  = ~\new_[15023]_ ;
  assign \new_[13785]_  = ~\new_[15025]_ ;
  assign \new_[13786]_  = ~\new_[16666]_  | ~\new_[18166]_ ;
  assign \new_[13787]_  = ~\new_[16474]_  | ~\new_[19754]_ ;
  assign \new_[13788]_  = ~\new_[16661]_  | ~\new_[18832]_ ;
  assign \new_[13789]_  = ~\new_[16058]_  | ~\new_[19044]_ ;
  assign \new_[13790]_  = ~\new_[17562]_  | ~\new_[17857]_ ;
  assign \new_[13791]_  = ~\new_[15343]_ ;
  assign \new_[13792]_  = ~\new_[15028]_ ;
  assign \new_[13793]_  = ~\new_[16575]_  | ~\new_[19031]_ ;
  assign \new_[13794]_  = \new_[16162]_  | \new_[19253]_ ;
  assign \new_[13795]_  = ~\new_[15031]_ ;
  assign \new_[13796]_  = ~\new_[15327]_ ;
  assign \new_[13797]_  = ~\new_[15033]_ ;
  assign \new_[13798]_  = ~\new_[15035]_ ;
  assign \new_[13799]_  = ~\new_[15037]_ ;
  assign \new_[13800]_  = ~\new_[15039]_ ;
  assign \new_[13801]_  = ~\new_[15040]_ ;
  assign \new_[13802]_  = ~\new_[16575]_  | ~\new_[20869]_ ;
  assign \new_[13803]_  = ~\new_[16661]_  | ~\new_[19676]_ ;
  assign \new_[13804]_  = ~\new_[15041]_ ;
  assign \new_[13805]_  = ~\new_[15295]_ ;
  assign \new_[13806]_  = ~\new_[15880]_  & ~\new_[19462]_ ;
  assign \new_[13807]_  = \new_[16090]_  & \new_[19409]_ ;
  assign \new_[13808]_  = \new_[16441]_  & \new_[19196]_ ;
  assign \new_[13809]_  = \new_[16643]_  & \new_[18637]_ ;
  assign \new_[13810]_  = \new_[16550]_  & \new_[19697]_ ;
  assign \new_[13811]_  = ~\new_[15048]_ ;
  assign \new_[13812]_  = ~\new_[16405]_  | ~\new_[18228]_ ;
  assign \new_[13813]_  = ~\new_[16502]_  | ~\new_[19426]_ ;
  assign \new_[13814]_  = ~\new_[15050]_ ;
  assign \new_[13815]_  = ~\new_[16382]_  & ~\new_[19145]_ ;
  assign \new_[13816]_  = ~\new_[19048]_  | ~\new_[17600]_ ;
  assign \new_[13817]_  = ~\new_[15149]_ ;
  assign \new_[13818]_  = ~\new_[15054]_ ;
  assign \new_[13819]_  = ~\new_[15055]_ ;
  assign \new_[13820]_  = ~\new_[15150]_ ;
  assign \new_[13821]_  = ~\new_[15883]_  | ~\new_[18979]_ ;
  assign \new_[13822]_  = ~\new_[15968]_  | ~\new_[18605]_ ;
  assign \new_[13823]_  = \new_[16380]_  | \new_[18840]_ ;
  assign \new_[13824]_  = ~\new_[20699]_  & ~\new_[20704]_  & ~\new_[16916]_ ;
  assign \new_[13825]_  = ~\new_[15087]_ ;
  assign \new_[13826]_  = ~\new_[15882]_  | ~\new_[19381]_ ;
  assign \new_[13827]_  = ~\new_[16276]_  | ~\new_[19082]_ ;
  assign \new_[13828]_  = ~\new_[15065]_ ;
  assign \new_[13829]_  = ~\new_[16027]_  | ~\new_[19044]_ ;
  assign \new_[13830]_  = ~\new_[17191]_  & ~\new_[19033]_ ;
  assign \new_[13831]_  = ~\new_[15060]_ ;
  assign \new_[13832]_  = ~\new_[15061]_ ;
  assign \new_[13833]_  = ~\new_[16171]_  & ~\new_[19474]_ ;
  assign \new_[13834]_  = ~\new_[15064]_ ;
  assign \new_[13835]_  = ~\new_[16631]_  | ~\new_[19156]_ ;
  assign \new_[13836]_  = ~\new_[21061]_  | ~\new_[18083]_ ;
  assign \new_[13837]_  = ~\new_[16000]_  | ~\new_[18810]_ ;
  assign \new_[13838]_  = ~\new_[16434]_  | ~\new_[20239]_ ;
  assign \new_[13839]_  = ~\new_[16500]_  | ~\new_[18111]_ ;
  assign \new_[13840]_  = ~\new_[16330]_  | ~\new_[19409]_ ;
  assign \new_[13841]_  = ~\new_[16157]_  | ~\new_[20239]_ ;
  assign \new_[13842]_  = ~\new_[15969]_  | ~\new_[19431]_ ;
  assign \new_[13843]_  = \new_[16009]_  & \new_[19082]_ ;
  assign \new_[13844]_  = ~\new_[19128]_  & ~\new_[16382]_ ;
  assign \new_[13845]_  = \new_[16651]_  & \new_[19298]_ ;
  assign \new_[13846]_  = ~\new_[16475]_  | ~\new_[18235]_ ;
  assign \new_[13847]_  = \new_[15886]_  | \new_[19655]_ ;
  assign \new_[13848]_  = ~\new_[16346]_  | ~\new_[19290]_ ;
  assign \new_[13849]_  = ~\new_[15070]_ ;
  assign \new_[13850]_  = ~\new_[15072]_ ;
  assign \new_[13851]_  = ~\new_[16462]_  | ~\new_[18938]_ ;
  assign \new_[13852]_  = ~\new_[15926]_  | ~\new_[18607]_ ;
  assign \new_[13853]_  = \new_[16447]_  & \new_[20865]_ ;
  assign \new_[13854]_  = ~\new_[16223]_  | ~\new_[18440]_ ;
  assign \new_[13855]_  = ~\new_[16551]_  | ~\new_[19096]_ ;
  assign \new_[13856]_  = \new_[15075]_ ;
  assign \new_[13857]_  = ~\new_[17038]_  | ~\new_[16460]_ ;
  assign \new_[13858]_  = ~\new_[16355]_  | ~\new_[18811]_ ;
  assign \new_[13859]_  = ~\new_[16095]_  | ~\new_[19144]_ ;
  assign \new_[13860]_  = ~\new_[15970]_  | ~\new_[18659]_ ;
  assign \new_[13861]_  = ~\new_[15078]_ ;
  assign \new_[13862]_  = ~\new_[15958]_  | ~\new_[19181]_ ;
  assign \new_[13863]_  = ~\new_[14931]_ ;
  assign \new_[13864]_  = ~\new_[16107]_  & ~\new_[21115]_ ;
  assign \new_[13865]_  = \new_[16148]_  & \new_[19181]_ ;
  assign \new_[13866]_  = ~\new_[16029]_  | ~\new_[18974]_ ;
  assign \new_[13867]_  = ~\new_[15278]_ ;
  assign \new_[13868]_  = ~\new_[15083]_ ;
  assign \new_[13869]_  = ~\new_[15575]_ ;
  assign \new_[13870]_  = ~\new_[21137]_ ;
  assign \new_[13871]_  = ~\new_[16442]_  | ~\new_[19687]_ ;
  assign \new_[13872]_  = ~\new_[14917]_ ;
  assign \new_[13873]_  = ~\new_[14910]_ ;
  assign \new_[13874]_  = \new_[15086]_ ;
  assign \new_[13875]_  = \new_[16332]_  | \new_[17089]_ ;
  assign \new_[13876]_  = ~\new_[16028]_  | ~\new_[18573]_ ;
  assign \new_[13877]_  = ~\new_[18335]_  & ~\new_[16491]_ ;
  assign \new_[13878]_  = \new_[16014]_  | \new_[19098]_ ;
  assign \new_[13879]_  = ~\new_[14895]_ ;
  assign \new_[13880]_  = ~\new_[15287]_ ;
  assign \new_[13881]_  = \new_[15905]_  | \new_[19253]_ ;
  assign \new_[13882]_  = ~\new_[15091]_ ;
  assign \new_[13883]_  = ~\new_[14888]_ ;
  assign \new_[13884]_  = ~\new_[16119]_  | ~\new_[19729]_ ;
  assign \new_[13885]_  = ~\new_[18430]_  & (~\new_[16831]_  | ~\new_[19263]_ );
  assign \new_[13886]_  = \new_[16422]_  | \new_[19156]_ ;
  assign \new_[13887]_  = ~\new_[14861]_ ;
  assign \new_[13888]_  = \new_[16660]_  | \new_[21508]_ ;
  assign \new_[13889]_  = ~\new_[16108]_  | ~\new_[18987]_ ;
  assign \new_[13890]_  = ~\new_[15096]_ ;
  assign \new_[13891]_  = ~\new_[15950]_  | ~\new_[19021]_ ;
  assign \new_[13892]_  = ~\new_[16442]_  | ~\new_[18840]_ ;
  assign \new_[13893]_  = ~\new_[14844]_ ;
  assign \new_[13894]_  = ~\new_[15099]_ ;
  assign \new_[13895]_  = \new_[20924]_  | \new_[19050]_ ;
  assign \new_[13896]_  = ~\new_[16362]_  | ~\new_[18046]_ ;
  assign \new_[13897]_  = ~\new_[14833]_ ;
  assign \new_[13898]_  = ~\new_[16227]_  | ~\new_[19084]_ ;
  assign \new_[13899]_  = ~\new_[21136]_ ;
  assign \new_[13900]_  = ~\new_[14820]_ ;
  assign \new_[13901]_  = ~\new_[16453]_  | ~\new_[18427]_ ;
  assign \new_[13902]_  = ~\new_[16483]_  | ~\new_[19217]_ ;
  assign \new_[13903]_  = \new_[16015]_  & \new_[21513]_ ;
  assign \new_[13904]_  = ~\new_[14813]_ ;
  assign \new_[13905]_  = ~\new_[16486]_  | ~\new_[19198]_ ;
  assign \new_[13906]_  = ~\new_[14801]_ ;
  assign \new_[13907]_  = \new_[16421]_  & \new_[18008]_ ;
  assign \new_[13908]_  = ~\new_[15105]_ ;
  assign \new_[13909]_  = \new_[16650]_  | \new_[18209]_ ;
  assign \new_[13910]_  = ~\new_[16635]_  | ~\new_[21306]_ ;
  assign \new_[13911]_  = ~\new_[16309]_  & ~\new_[19096]_ ;
  assign \new_[13912]_  = ~\new_[16341]_  | ~\new_[18969]_ ;
  assign \new_[13913]_  = ~\new_[16362]_  | ~\new_[21510]_ ;
  assign \new_[13914]_  = \new_[15107]_ ;
  assign \new_[13915]_  = \new_[16385]_  & \new_[18414]_ ;
  assign \new_[13916]_  = ~\new_[16007]_  | ~\new_[19194]_ ;
  assign \new_[13917]_  = ~\new_[15108]_ ;
  assign \new_[13918]_  = \new_[16191]_  & \new_[21685]_ ;
  assign \new_[13919]_  = ~\new_[16357]_  | ~\new_[18061]_ ;
  assign \new_[13920]_  = ~\new_[17171]_  | ~\new_[19021]_ ;
  assign \new_[13921]_  = ~\new_[16047]_  | ~\new_[19006]_ ;
  assign \new_[13922]_  = ~\new_[16453]_  | ~\new_[18847]_ ;
  assign \new_[13923]_  = ~\new_[16597]_  | ~\new_[19196]_ ;
  assign \new_[13924]_  = \new_[16292]_  | \new_[18832]_ ;
  assign \new_[13925]_  = ~\new_[15110]_ ;
  assign \new_[13926]_  = ~\new_[15311]_ ;
  assign \new_[13927]_  = ~\new_[15058]_ ;
  assign \new_[13928]_  = ~\new_[15111]_ ;
  assign \new_[13929]_  = ~\new_[16500]_  | ~\new_[19079]_ ;
  assign \new_[13930]_  = \new_[16555]_  & \new_[19031]_ ;
  assign \new_[13931]_  = \new_[16480]_  & \new_[20927]_ ;
  assign \new_[13932]_  = ~\new_[15112]_ ;
  assign \new_[13933]_  = ~\new_[16367]_  | ~\new_[18972]_ ;
  assign \new_[13934]_  = ~\new_[15868]_  | ~\new_[19018]_ ;
  assign \new_[13935]_  = ~\new_[14739]_ ;
  assign \new_[13936]_  = ~\new_[14733]_ ;
  assign \new_[13937]_  = ~\new_[16439]_  | ~\new_[18652]_ ;
  assign \new_[13938]_  = ~\new_[16530]_  | ~\new_[18903]_ ;
  assign \new_[13939]_  = ~\new_[15114]_ ;
  assign \new_[13940]_  = ~\new_[16375]_  | ~\new_[18926]_ ;
  assign \new_[13941]_  = ~\new_[16461]_  | ~\new_[18938]_ ;
  assign \new_[13942]_  = ~\new_[15390]_ ;
  assign \new_[13943]_  = ~\new_[15117]_ ;
  assign \new_[13944]_  = \new_[15873]_  & \new_[18979]_ ;
  assign \new_[13945]_  = ~\new_[17964]_  | ~\new_[17358]_ ;
  assign \new_[13946]_  = ~\new_[16348]_  & ~\new_[18984]_ ;
  assign \new_[13947]_  = ~\new_[16554]_  & ~\new_[21560]_ ;
  assign \new_[13948]_  = \new_[16536]_  & \new_[19068]_ ;
  assign \new_[13949]_  = \new_[16099]_  | \new_[18246]_ ;
  assign \new_[13950]_  = ~\new_[16430]_  | ~\new_[19290]_ ;
  assign \new_[13951]_  = ~\new_[14713]_ ;
  assign \new_[13952]_  = ~\new_[14699]_ ;
  assign \new_[13953]_  = ~\new_[16572]_  | ~\new_[19426]_ ;
  assign \new_[13954]_  = \new_[16296]_  | \new_[18941]_ ;
  assign \new_[13955]_  = ~\new_[15882]_  | ~\new_[21695]_ ;
  assign \new_[13956]_  = ~\new_[16137]_  | ~\new_[18605]_ ;
  assign \new_[13957]_  = ~\new_[14695]_ ;
  assign \new_[13958]_  = \new_[17876]_  | \new_[18209]_ ;
  assign \new_[13959]_  = ~\new_[15862]_ ;
  assign \new_[13960]_  = ~\new_[16019]_  | ~\new_[18938]_ ;
  assign \new_[13961]_  = ~\new_[15844]_ ;
  assign \new_[13962]_  = ~\new_[15128]_ ;
  assign \new_[13963]_  = ~\new_[16152]_  | ~\new_[19162]_ ;
  assign \new_[13964]_  = ~\new_[15129]_ ;
  assign \new_[13965]_  = \new_[15904]_  & \new_[19082]_ ;
  assign \new_[13966]_  = ~\new_[15130]_ ;
  assign \new_[13967]_  = ~\new_[19685]_  | ~\new_[19213]_  | ~\new_[18161]_ ;
  assign \new_[13968]_  = ~\new_[16565]_  | ~\new_[19738]_ ;
  assign \new_[13969]_  = ~\new_[16433]_  | ~\new_[19100]_ ;
  assign \new_[13970]_  = ~\new_[16301]_  & ~\new_[19023]_ ;
  assign \new_[13971]_  = ~\new_[18837]_  | ~\new_[18841]_  | ~\new_[19088]_  | ~\new_[19398]_ ;
  assign \new_[13972]_  = ~\new_[16645]_  | ~\new_[19446]_ ;
  assign \new_[13973]_  = ~\new_[15134]_ ;
  assign \new_[13974]_  = ~\new_[16300]_  | ~\new_[21168]_ ;
  assign \new_[13975]_  = ~\new_[15136]_ ;
  assign \new_[13976]_  = ~\new_[21564]_  & ~\new_[21697]_ ;
  assign \new_[13977]_  = ~\new_[16293]_  | ~\new_[19217]_ ;
  assign \new_[13978]_  = ~\new_[20663]_  | ~\new_[18852]_ ;
  assign \new_[13979]_  = ~\new_[16275]_  | ~\new_[19676]_ ;
  assign \new_[13980]_  = ~\new_[15925]_  | ~\new_[18678]_ ;
  assign \new_[13981]_  = ~\new_[15139]_ ;
  assign \new_[13982]_  = ~\new_[16469]_  | ~\new_[18083]_ ;
  assign \new_[13983]_  = \new_[16586]_  | \new_[18709]_ ;
  assign \new_[13984]_  = \new_[16493]_  | \new_[19141]_ ;
  assign \new_[13985]_  = ~\new_[16298]_  & ~\new_[18627]_ ;
  assign \new_[13986]_  = ~\new_[15877]_  | ~\new_[21505]_ ;
  assign \new_[13987]_  = ~\new_[15142]_ ;
  assign \new_[13988]_  = ~\new_[15919]_  | ~\new_[19538]_ ;
  assign \new_[13989]_  = ~\new_[15146]_ ;
  assign \new_[13990]_  = ~\new_[15282]_ ;
  assign \new_[13991]_  = ~\new_[16208]_  & ~\new_[21569]_ ;
  assign \new_[13992]_  = ~\new_[17043]_  | ~\new_[21392]_ ;
  assign \new_[13993]_  = ~\new_[21410]_  | ~\new_[18974]_ ;
  assign \new_[13994]_  = ~\new_[16094]_  & ~\new_[18209]_ ;
  assign \new_[13995]_  = ~\new_[16366]_  & ~\new_[15945]_ ;
  assign \new_[13996]_  = ~\new_[15532]_ ;
  assign \new_[13997]_  = ~\new_[16337]_  & ~\new_[18678]_ ;
  assign \new_[13998]_  = ~\new_[16638]_  | ~\new_[18209]_ ;
  assign \new_[13999]_  = ~\new_[17780]_  & ~\new_[21628]_ ;
  assign \new_[14000]_  = ~\new_[15155]_ ;
  assign \new_[14001]_  = ~\new_[15498]_ ;
  assign \new_[14002]_  = ~\new_[16504]_  | ~\new_[19023]_ ;
  assign \new_[14003]_  = ~\new_[20661]_  | ~\new_[15866]_ ;
  assign \new_[14004]_  = ~\new_[15444]_ ;
  assign \new_[14005]_  = ~\new_[15154]_ ;
  assign \new_[14006]_  = ~\new_[16068]_  & ~\new_[18664]_ ;
  assign \new_[14007]_  = ~\new_[15158]_ ;
  assign \new_[14008]_  = ~\new_[16068]_  & ~\new_[19130]_ ;
  assign \new_[14009]_  = ~\new_[16311]_  | ~\new_[19031]_ ;
  assign \new_[14010]_  = ~\new_[15159]_ ;
  assign \new_[14011]_  = ~\new_[19027]_  & ~\new_[15887]_ ;
  assign \new_[14012]_  = ~\new_[17339]_  | ~\new_[16400]_ ;
  assign \new_[14013]_  = ~\new_[15160]_ ;
  assign \new_[14014]_  = ~\new_[16211]_  | ~\new_[19538]_ ;
  assign \new_[14015]_  = ~\new_[15163]_ ;
  assign \new_[14016]_  = ~\new_[15164]_ ;
  assign \new_[14017]_  = ~\new_[16176]_  & ~\new_[19151]_ ;
  assign \new_[14018]_  = ~\new_[15167]_ ;
  assign \new_[14019]_  = \new_[16404]_  | \new_[19409]_ ;
  assign \new_[14020]_  = \new_[18022]_  | \new_[15991]_ ;
  assign \new_[14021]_  = ~\new_[15891]_  & ~\new_[18008]_ ;
  assign \new_[14022]_  = ~\new_[16605]_  | ~\new_[21688]_ ;
  assign \new_[14023]_  = ~\new_[16412]_  | ~\new_[19098]_ ;
  assign \new_[14024]_  = \new_[17390]_  | \new_[18396]_ ;
  assign \new_[14025]_  = ~\new_[16297]_  | ~\new_[17983]_ ;
  assign \new_[14026]_  = \new_[16457]_  & \new_[19675]_ ;
  assign \new_[14027]_  = ~\new_[16542]_  | ~\new_[19637]_ ;
  assign \new_[14028]_  = ~\new_[16175]_  & ~\new_[19454]_ ;
  assign \new_[14029]_  = ~\new_[15317]_ ;
  assign \new_[14030]_  = ~\new_[21410]_  | ~\new_[18817]_ ;
  assign \new_[14031]_  = ~\new_[19026]_  & ~\new_[17481]_ ;
  assign \new_[14032]_  = ~\new_[16503]_  & (~\new_[18196]_  | ~\new_[19425]_ );
  assign \new_[14033]_  = ~\new_[15302]_ ;
  assign \new_[14034]_  = \new_[16363]_  & \new_[19547]_ ;
  assign \new_[14035]_  = ~\new_[16436]_  | ~\new_[19153]_ ;
  assign \new_[14036]_  = ~\new_[19228]_  | ~\new_[15951]_ ;
  assign \new_[14037]_  = ~\new_[15171]_ ;
  assign \new_[14038]_  = ~\new_[15172]_ ;
  assign \new_[14039]_  = ~\new_[15246]_ ;
  assign \new_[14040]_  = ~\new_[14839]_ ;
  assign \new_[14041]_  = \new_[16542]_  & \new_[18616]_ ;
  assign \new_[14042]_  = ~\new_[17098]_ ;
  assign \new_[14043]_  = ~\new_[15175]_ ;
  assign \new_[14044]_  = ~\new_[15176]_ ;
  assign \new_[14045]_  = \new_[16446]_  | \new_[20680]_ ;
  assign \new_[14046]_  = ~\new_[16152]_  | ~\new_[19024]_ ;
  assign \new_[14047]_  = ~\new_[16573]_  & ~\new_[19474]_ ;
  assign \new_[14048]_  = ~\new_[15898]_  | ~\new_[17081]_ ;
  assign \new_[14049]_  = ~\new_[15179]_ ;
  assign \new_[14050]_  = ~\new_[19676]_  | ~\new_[17605]_ ;
  assign \new_[14051]_  = \new_[18117]_  | \new_[15959]_ ;
  assign \new_[14052]_  = ~\new_[16113]_  | ~\new_[18984]_ ;
  assign \new_[14053]_  = ~\new_[15182]_ ;
  assign \new_[14054]_  = ~\new_[16606]_  | ~\new_[21506]_ ;
  assign \new_[14055]_  = ~\new_[15185]_ ;
  assign \new_[14056]_  = ~\new_[15186]_ ;
  assign \new_[14057]_  = ~\new_[16668]_  & ~\new_[19130]_ ;
  assign \new_[14058]_  = ~\new_[16570]_  | ~\new_[21574]_ ;
  assign \new_[14059]_  = ~\new_[15044]_ ;
  assign \new_[14060]_  = ~\new_[15931]_  | ~\new_[19064]_ ;
  assign \new_[14061]_  = ~\new_[16468]_  | ~\new_[17179]_ ;
  assign \new_[14062]_  = \new_[16431]_  | \new_[18414]_ ;
  assign \new_[14063]_  = ~\new_[15018]_ ;
  assign \new_[14064]_  = \new_[14902]_  ^ \new_[16980]_ ;
  assign \new_[14065]_  = ~\new_[16397]_  & ~\new_[17754]_ ;
  assign \new_[14066]_  = \new_[17785]_  | \new_[19008]_ ;
  assign \new_[14067]_  = ~\new_[14996]_ ;
  assign \new_[14068]_  = ~\new_[15194]_ ;
  assign \new_[14069]_  = ~\new_[16039]_  & ~\new_[20704]_ ;
  assign \new_[14070]_  = ~\new_[15368]_ ;
  assign \new_[14071]_  = ~\new_[16393]_  & ~\new_[16097]_ ;
  assign \new_[14072]_  = ~\new_[16146]_  & ~\new_[19779]_ ;
  assign \new_[14073]_  = ~\new_[15196]_ ;
  assign \new_[14074]_  = ~\new_[16075]_  | ~\new_[18325]_ ;
  assign \new_[14075]_  = ~\new_[14952]_ ;
  assign \new_[14076]_  = \new_[15983]_  | \new_[19253]_ ;
  assign \new_[14077]_  = ~\new_[16312]_  & ~\new_[18008]_ ;
  assign \new_[14078]_  = ~\new_[15205]_ ;
  assign \new_[14079]_  = \new_[17822]_  | \new_[18832]_ ;
  assign \new_[14080]_  = ~\new_[14925]_ ;
  assign \new_[14081]_  = ~\new_[16664]_  & ~\new_[19085]_ ;
  assign \new_[14082]_  = \new_[17641]_  | \new_[19727]_ ;
  assign \new_[14083]_  = ~\new_[16656]_  | ~\new_[19217]_ ;
  assign \new_[14084]_  = ~\new_[16497]_  & ~\new_[19214]_ ;
  assign \new_[14085]_  = ~\new_[17983]_  | ~\new_[17501]_ ;
  assign \new_[14086]_  = ~\new_[15975]_  | ~\new_[19008]_ ;
  assign \new_[14087]_  = ~\new_[15207]_ ;
  assign \new_[14088]_  = ~\new_[16089]_  | ~\new_[19215]_ ;
  assign \new_[14089]_  = ~\new_[18080]_  | ~\new_[17171]_ ;
  assign \new_[14090]_  = ~\new_[16519]_  & ~\new_[15984]_ ;
  assign \new_[14091]_  = ~\new_[14928]_ ;
  assign \new_[14092]_  = ~\new_[17292]_  | ~\new_[16472]_ ;
  assign \new_[14093]_  = ~\new_[17726]_  | ~\new_[19186]_ ;
  assign \new_[14094]_  = ~\new_[15211]_ ;
  assign \new_[14095]_  = (~\new_[16705]_  | ~\new_[9578]_ ) & (~\new_[18555]_  | ~\new_[18411]_ );
  assign \new_[14096]_  = \new_[16109]_  & \new_[19327]_ ;
  assign \new_[14097]_  = \new_[16633]_  | \new_[18008]_ ;
  assign \new_[14098]_  = ~\new_[16145]_  | ~\new_[16770]_ ;
  assign \new_[14099]_  = ~\new_[15213]_ ;
  assign \new_[14100]_  = ~\new_[16374]_  | ~\new_[16074]_ ;
  assign \new_[14101]_  = ~\new_[19444]_  & ~\new_[16156]_ ;
  assign \new_[14102]_  = ~\new_[16503]_  | ~\new_[19335]_ ;
  assign \new_[14103]_  = ~\new_[14887]_ ;
  assign \new_[14104]_  = ~\new_[15569]_ ;
  assign \new_[14105]_  = ~\new_[16558]_  | ~\new_[19239]_ ;
  assign \new_[14106]_  = ~\new_[14868]_ ;
  assign \new_[14107]_  = \new_[15984]_  & \new_[19758]_ ;
  assign \new_[14108]_  = ~\new_[16308]_  | ~\new_[17488]_ ;
  assign \new_[14109]_  = ~\new_[15216]_ ;
  assign \new_[14110]_  = ~\new_[15276]_ ;
  assign \new_[14111]_  = ~\new_[16310]_  | ~\new_[17165]_ ;
  assign \new_[14112]_  = ~\new_[14829]_ ;
  assign \new_[14113]_  = ~\new_[16331]_  | ~\new_[18978]_ ;
  assign \new_[14114]_  = \new_[17822]_  | \new_[19742]_ ;
  assign \new_[14115]_  = ~\new_[16170]_  | ~\new_[19239]_ ;
  assign \new_[14116]_  = ~\new_[15217]_ ;
  assign \new_[14117]_  = ~\new_[19675]_  | ~\new_[16484]_ ;
  assign \new_[14118]_  = ~\new_[16443]_  & ~\new_[16126]_ ;
  assign \new_[14119]_  = \new_[16263]_  | \new_[19141]_ ;
  assign \new_[14120]_  = \new_[15878]_  | \new_[19156]_ ;
  assign \new_[14121]_  = ~\new_[14808]_ ;
  assign \new_[14122]_  = ~\new_[14808]_ ;
  assign \new_[14123]_  = ~\new_[14803]_ ;
  assign \new_[14124]_  = ~\new_[15220]_ ;
  assign \new_[14125]_  = ~\new_[16457]_  | ~\new_[19374]_ ;
  assign \new_[14126]_  = ~\new_[15229]_ ;
  assign \new_[14127]_  = ~\new_[15222]_ ;
  assign \new_[14128]_  = ~\new_[17501]_  | ~\new_[20239]_ ;
  assign \new_[14129]_  = \new_[16389]_  | \new_[19196]_ ;
  assign \new_[14130]_  = \new_[17850]_  | \new_[18076]_ ;
  assign \new_[14131]_  = ~\new_[16045]_  & ~\new_[18003]_ ;
  assign \new_[14132]_  = ~\new_[14741]_ ;
  assign \new_[14133]_  = ~\new_[16064]_  & ~\new_[19059]_ ;
  assign \new_[14134]_  = ~\new_[15228]_ ;
  assign \new_[14135]_  = ~\new_[16431]_  & ~\new_[19553]_ ;
  assign \new_[14136]_  = ~\new_[16584]_  | ~\new_[18811]_ ;
  assign \new_[14137]_  = ~\new_[16534]_  & ~\new_[18966]_ ;
  assign \new_[14138]_  = ~\new_[16514]_  | ~\new_[18194]_ ;
  assign \new_[14139]_  = ~\new_[14721]_ ;
  assign \new_[14140]_  = ~\new_[15221]_ ;
  assign \new_[14141]_  = \new_[16032]_  | \new_[19409]_ ;
  assign \new_[14142]_  = \new_[17569]_  | \new_[18209]_ ;
  assign \new_[14143]_  = ~\new_[16476]_  | ~\new_[16703]_ ;
  assign \new_[14144]_  = ~\new_[15230]_ ;
  assign \new_[14145]_  = ~\new_[15932]_  | ~\new_[16322]_ ;
  assign \new_[14146]_  = ~\new_[20586]_  | ~\new_[18643]_ ;
  assign \new_[14147]_  = ~\new_[15909]_  | ~\new_[18832]_ ;
  assign \new_[14148]_  = ~\new_[17847]_  & ~\new_[16674]_ ;
  assign \new_[14149]_  = ~\new_[15240]_ ;
  assign \new_[14150]_  = ~\new_[15825]_ ;
  assign \new_[14151]_  = \new_[18082]_  | \new_[16412]_ ;
  assign \new_[14152]_  = ~\new_[18659]_  | ~\new_[16075]_ ;
  assign \new_[14153]_  = ~\new_[17086]_  | ~\new_[16672]_ ;
  assign \new_[14154]_  = ~\new_[15241]_ ;
  assign \new_[14155]_  = ~\new_[16423]_  | ~\new_[18083]_ ;
  assign \new_[14156]_  = ~\new_[15929]_  & ~\new_[19156]_ ;
  assign \new_[14157]_  = ~\new_[16149]_  & ~\new_[17886]_ ;
  assign \new_[14158]_  = ~\new_[19222]_  | ~\new_[16584]_ ;
  assign \new_[14159]_  = ~\new_[15761]_ ;
  assign \new_[14160]_  = ~\new_[16183]_  & ~\new_[19240]_ ;
  assign \new_[14161]_  = ~\new_[15242]_ ;
  assign \new_[14162]_  = \new_[17536]_  & \new_[16594]_ ;
  assign \new_[14163]_  = ~\new_[16168]_  | ~\new_[18974]_ ;
  assign \new_[14164]_  = \new_[16194]_  | \new_[16202]_ ;
  assign \new_[14165]_  = ~\new_[17737]_  | ~\new_[19269]_ ;
  assign \new_[14166]_  = \new_[16508]_  | \new_[19456]_ ;
  assign \new_[14167]_  = ~\new_[15684]_ ;
  assign \new_[14168]_  = ~\new_[18609]_  & ~\new_[16064]_ ;
  assign \new_[14169]_  = ~\new_[16520]_  & ~\new_[17618]_ ;
  assign \new_[14170]_  = ~\new_[15247]_ ;
  assign \new_[14171]_  = \new_[15871]_  | \new_[19758]_ ;
  assign \new_[14172]_  = ~\new_[18709]_  & ~\new_[17775]_ ;
  assign \new_[14173]_  = ~\new_[18898]_  | ~\new_[16504]_ ;
  assign \new_[14174]_  = ~\new_[16316]_  & ~\new_[19021]_ ;
  assign \new_[14175]_  = ~\new_[15947]_  | ~\new_[19064]_ ;
  assign \new_[14176]_  = ~\new_[17792]_  | ~\new_[16585]_ ;
  assign \new_[14177]_  = \new_[16383]_  | \new_[19742]_ ;
  assign \new_[14178]_  = ~\new_[15567]_ ;
  assign \new_[14179]_  = ~\new_[18657]_  & ~\new_[16527]_ ;
  assign \new_[14180]_  = ~\new_[15957]_  | ~\new_[19568]_ ;
  assign \new_[14181]_  = ~\new_[14934]_ ;
  assign \new_[14182]_  = ~\new_[15578]_ ;
  assign \new_[14183]_  = ~\new_[15251]_ ;
  assign \new_[14184]_  = ~\new_[15555]_ ;
  assign \new_[14185]_  = ~\new_[18106]_  & ~\new_[16136]_ ;
  assign \new_[14186]_  = ~\new_[17522]_  | ~\new_[16502]_ ;
  assign \new_[14187]_  = ~\new_[15255]_ ;
  assign \new_[14188]_  = ~\new_[17652]_  & ~\new_[19431]_ ;
  assign \new_[14189]_  = ~\new_[16115]_  | ~\new_[19353]_ ;
  assign \new_[14190]_  = ~\new_[16170]_  & ~\new_[17194]_ ;
  assign \new_[14191]_  = ~\new_[15436]_ ;
  assign \new_[14192]_  = ~\new_[15426]_ ;
  assign \new_[14193]_  = ~\new_[15411]_ ;
  assign \new_[14194]_  = \new_[17926]_  | \new_[16025]_ ;
  assign \new_[14195]_  = ~\new_[15260]_ ;
  assign \new_[14196]_  = ~\new_[15261]_ ;
  assign \new_[14197]_  = ~\new_[18807]_  | ~\new_[17171]_ ;
  assign \new_[14198]_  = ~\new_[15913]_  | ~\new_[19568]_ ;
  assign \new_[14199]_  = ~\new_[17605]_  | ~\new_[19738]_ ;
  assign \new_[14200]_  = ~\new_[18083]_  & ~\new_[16149]_ ;
  assign \new_[14201]_  = ~\new_[15912]_  | ~\new_[20699]_ ;
  assign \new_[14202]_  = ~\new_[15265]_ ;
  assign \new_[14203]_  = ~\new_[15266]_ ;
  assign \new_[14204]_  = ~\new_[15267]_ ;
  assign \new_[14205]_  = ~\new_[15268]_ ;
  assign \new_[14206]_  = ~\new_[15314]_ ;
  assign \new_[14207]_  = ~\new_[15908]_  | ~\new_[19217]_ ;
  assign \new_[14208]_  = ~\new_[15283]_ ;
  assign \new_[14209]_  = ~\new_[16590]_  & ~\new_[19675]_ ;
  assign \new_[14210]_  = ~\new_[16321]_  | ~\new_[19617]_ ;
  assign \new_[14211]_  = ~\new_[16318]_  | ~\new_[19181]_ ;
  assign \new_[14212]_  = ~\new_[16232]_  & ~\new_[21571]_ ;
  assign \new_[14213]_  = ~\new_[15275]_ ;
  assign \new_[14214]_  = ~\new_[15210]_ ;
  assign \new_[14215]_  = ~\new_[16504]_  | ~\new_[19474]_ ;
  assign \new_[14216]_  = \new_[16580]_  | \new_[19082]_ ;
  assign \new_[14217]_  = ~\new_[16126]_  | ~\new_[19082]_ ;
  assign \new_[14218]_  = \new_[16529]_  | \new_[19153]_ ;
  assign \new_[14219]_  = ~\new_[16138]_  & ~\new_[18766]_ ;
  assign \new_[14220]_  = \new_[16337]_  | \new_[21413]_ ;
  assign \new_[14221]_  = ~\new_[14744]_ ;
  assign \new_[14222]_  = ~\new_[16503]_  | ~\new_[19158]_ ;
  assign \new_[14223]_  = \new_[16054]_  | \new_[19233]_ ;
  assign \new_[14224]_  = \new_[16197]_  | \new_[19553]_ ;
  assign \new_[14225]_  = ~\new_[15805]_ ;
  assign \new_[14226]_  = ~\new_[15100]_ ;
  assign \new_[14227]_  = ~\new_[15286]_ ;
  assign \new_[14228]_  = ~\new_[17452]_  & ~\new_[15987]_ ;
  assign \new_[14229]_  = ~\new_[16126]_  | ~\new_[18371]_ ;
  assign \new_[14230]_  = ~\new_[15969]_  | ~\new_[18909]_ ;
  assign \new_[14231]_  = ~\new_[18614]_  | ~\new_[16047]_ ;
  assign \new_[14232]_  = \new_[19073]_  | \new_[16559]_ ;
  assign \new_[14233]_  = ~\new_[15481]_ ;
  assign \new_[14234]_  = ~\new_[16091]_  & ~\new_[16052]_ ;
  assign \new_[14235]_  = ~\new_[18815]_  & ~\new_[16734]_ ;
  assign \new_[14236]_  = ~\new_[15051]_ ;
  assign \new_[14237]_  = ~\new_[15290]_ ;
  assign \new_[14238]_  = ~\new_[15030]_ ;
  assign \new_[14239]_  = ~\new_[15027]_ ;
  assign \new_[14240]_  = ~\new_[21410]_  | ~\new_[18987]_ ;
  assign \new_[14241]_  = ~\new_[17461]_  | ~\new_[16047]_ ;
  assign \new_[14242]_  = ~\new_[15292]_ ;
  assign \new_[14243]_  = ~\new_[15293]_ ;
  assign \new_[14244]_  = ~\new_[15941]_  | ~\new_[19024]_ ;
  assign \new_[14245]_  = ~\new_[16105]_  & ~\new_[16987]_ ;
  assign \new_[14246]_  = ~\new_[15294]_ ;
  assign \new_[14247]_  = ~\new_[16584]_  | ~\new_[18692]_ ;
  assign \new_[14248]_  = ~\new_[20905]_ ;
  assign \new_[14249]_  = ~\new_[16097]_  | ~\new_[19130]_ ;
  assign \new_[14250]_  = \new_[16400]_  | \new_[19538]_ ;
  assign \new_[14251]_  = ~\new_[18037]_  | ~\new_[15912]_ ;
  assign \new_[14252]_  = ~\new_[16538]_  | ~\new_[17917]_ ;
  assign \new_[14253]_  = ~\new_[16283]_  & ~\new_[19462]_ ;
  assign \new_[14254]_  = ~\new_[17906]_  & ~\new_[19476]_ ;
  assign \new_[14255]_  = ~\new_[21113]_  & ~\new_[19154]_ ;
  assign \new_[14256]_  = ~\new_[16291]_  & ~\new_[19151]_ ;
  assign \new_[14257]_  = ~\new_[14950]_ ;
  assign \new_[14258]_  = ~\new_[15872]_  | ~\new_[19681]_ ;
  assign \new_[14259]_  = ~\new_[15984]_  | ~\new_[19026]_ ;
  assign \new_[14260]_  = ~\new_[15305]_ ;
  assign \new_[14261]_  = \new_[16085]_  & \new_[18209]_ ;
  assign \new_[14262]_  = \new_[16508]_  | \new_[18209]_ ;
  assign \new_[14263]_  = ~\new_[16074]_  | ~\new_[16309]_ ;
  assign \new_[14264]_  = ~\new_[15308]_ ;
  assign \new_[14265]_  = ~\new_[16278]_  & ~\new_[19261]_ ;
  assign \new_[14266]_  = ~\new_[16419]_  | ~\new_[18542]_ ;
  assign \new_[14267]_  = ~\new_[16037]_ ;
  assign \new_[14268]_  = ~\new_[19097]_  | ~\new_[15944]_ ;
  assign \new_[14269]_  = ~\new_[16594]_  | ~\new_[21328]_ ;
  assign \new_[14270]_  = ~\new_[15990]_  & ~\new_[20239]_ ;
  assign \new_[14271]_  = ~\new_[17872]_  | ~\new_[19117]_ ;
  assign \new_[14272]_  = ~\new_[15316]_ ;
  assign \new_[14273]_  = ~\new_[16051]_  & ~\new_[18936]_ ;
  assign \new_[14274]_  = \new_[16660]_  & \new_[16336]_ ;
  assign \new_[14275]_  = ~\new_[15924]_  | ~\new_[19061]_ ;
  assign \new_[14276]_  = ~\new_[17867]_  | ~\new_[17632]_ ;
  assign \new_[14277]_  = ~\new_[17569]_  & ~\new_[19815]_ ;
  assign \new_[14278]_  = ~\new_[16641]_  & ~\new_[19746]_ ;
  assign \new_[14279]_  = ~\new_[15319]_ ;
  assign \new_[14280]_  = ~\new_[20768]_  & ~\new_[16025]_ ;
  assign \new_[14281]_  = ~\new_[15324]_ ;
  assign \new_[14282]_  = ~\new_[15943]_  & ~\new_[21635]_ ;
  assign \new_[14283]_  = ~\new_[14735]_ ;
  assign \new_[14284]_  = ~\new_[15924]_  | ~\new_[19428]_ ;
  assign \new_[14285]_  = ~\new_[16596]_  | ~\new_[18987]_ ;
  assign \new_[14286]_  = \new_[16265]_  | \new_[21502]_ ;
  assign \new_[14287]_  = ~\new_[16662]_  | ~\new_[21259]_ ;
  assign \new_[14288]_  = \new_[15837]_ ;
  assign \new_[14289]_  = ~\new_[15770]_ ;
  assign \new_[14290]_  = ~\new_[15860]_ ;
  assign \new_[14291]_  = ~\new_[15330]_ ;
  assign \new_[14292]_  = ~\new_[18179]_  | ~\new_[16876]_  | ~\new_[17792]_ ;
  assign \new_[14293]_  = ~\new_[16059]_  | ~\new_[19535]_ ;
  assign \new_[14294]_  = ~\new_[17939]_  | ~\new_[16637]_ ;
  assign \new_[14295]_  = ~\new_[15789]_ ;
  assign \new_[14296]_  = ~\new_[15772]_ ;
  assign \new_[14297]_  = ~\new_[18643]_  | ~\new_[16214]_ ;
  assign \new_[14298]_  = ~\new_[16576]_  & ~\new_[19261]_ ;
  assign \new_[14299]_  = ~\new_[18403]_  | ~\new_[16674]_ ;
  assign \new_[14300]_  = \new_[16473]_  & \new_[20704]_ ;
  assign \new_[14301]_  = ~\new_[16087]_  | ~\new_[19095]_ ;
  assign \new_[14302]_  = ~\new_[15945]_  | ~\new_[19084]_ ;
  assign \new_[14303]_  = ~\new_[18849]_  | ~\new_[15972]_ ;
  assign \new_[14304]_  = ~\new_[18947]_  | ~\new_[16205]_ ;
  assign \new_[14305]_  = ~\new_[15945]_  | ~\new_[19444]_ ;
  assign \new_[14306]_  = ~\new_[17780]_  & ~\new_[19018]_ ;
  assign \new_[14307]_  = \new_[18062]_  | \new_[16215]_ ;
  assign \new_[14308]_  = ~\new_[15522]_ ;
  assign \new_[14309]_  = ~\new_[17896]_  & ~\new_[14951]_ ;
  assign \new_[14310]_  = ~\new_[15944]_  | ~\new_[18973]_ ;
  assign \new_[14311]_  = ~\new_[15710]_ ;
  assign \new_[14312]_  = ~\new_[15943]_  & ~\new_[19018]_ ;
  assign \new_[14313]_  = ~\new_[16782]_  | ~\new_[16315]_ ;
  assign \new_[14314]_  = ~\new_[14918]_ ;
  assign \new_[14315]_  = ~\new_[15338]_ ;
  assign \new_[14316]_  = ~\new_[16279]_  | ~\new_[18682]_ ;
  assign \new_[14317]_  = ~\new_[16024]_  & ~\new_[21507]_ ;
  assign \new_[14318]_  = ~\new_[17694]_  & ~\new_[19182]_ ;
  assign \new_[14319]_  = \new_[18657]_  | \new_[16493]_ ;
  assign \new_[14320]_  = ~\new_[15337]_ ;
  assign \new_[14321]_  = ~\new_[14819]_ ;
  assign \new_[14322]_  = ~\new_[19260]_  | ~\new_[16662]_ ;
  assign \new_[14323]_  = ~\new_[15709]_ ;
  assign \new_[14324]_  = \new_[16258]_  | \new_[16417]_ ;
  assign \new_[14325]_  = ~\new_[16339]_  | ~\new_[19409]_ ;
  assign \new_[14326]_  = ~\new_[15168]_ ;
  assign \new_[14327]_  = ~\new_[15342]_ ;
  assign \new_[14328]_  = ~\new_[16436]_  & ~\new_[16135]_ ;
  assign \new_[14329]_  = ~\new_[16289]_  | ~\new_[18166]_ ;
  assign \new_[14330]_  = ~\new_[15122]_ ;
  assign \new_[14331]_  = ~\new_[17802]_  | ~\new_[15961]_ ;
  assign \new_[14332]_  = ~\new_[15346]_ ;
  assign \new_[14333]_  = ~\new_[17402]_  | ~\new_[16635]_ ;
  assign \new_[14334]_  = ~\new_[18332]_  | ~\new_[15955]_ ;
  assign \new_[14335]_  = ~\new_[18284]_  | ~\new_[18045]_  | ~\new_[18542]_  | ~\new_[19217]_ ;
  assign \new_[14336]_  = ~\new_[15074]_ ;
  assign \new_[14337]_  = ~\new_[16388]_  | ~\new_[19224]_ ;
  assign \new_[14338]_  = ~\new_[17853]_  | ~\new_[19217]_ ;
  assign \new_[14339]_  = ~\new_[16438]_  | ~\new_[16081]_ ;
  assign \new_[14340]_  = \new_[17641]_  | \new_[19158]_ ;
  assign \new_[14341]_  = ~\new_[16127]_  & ~\new_[18083]_ ;
  assign \new_[14342]_  = ~\new_[16400]_  | ~\new_[18017]_ ;
  assign \new_[14343]_  = ~\new_[16262]_ ;
  assign \new_[14344]_  = ~\new_[16341]_  | ~\new_[18957]_ ;
  assign \new_[14345]_  = ~\new_[16517]_  | ~\new_[19239]_ ;
  assign \new_[14346]_  = ~\new_[15352]_ ;
  assign \new_[14347]_  = ~\new_[16535]_  | ~\new_[19196]_ ;
  assign \new_[14348]_  = ~\new_[15932]_  | (~\new_[18182]_  & ~\new_[18060]_ );
  assign \new_[14349]_  = ~\new_[15356]_ ;
  assign \new_[14350]_  = ~\new_[17440]_  & ~\new_[15957]_ ;
  assign \new_[14351]_  = \new_[15916]_  | \new_[19374]_ ;
  assign \new_[14352]_  = ~\new_[16392]_  & ~\new_[16087]_ ;
  assign \new_[14353]_  = \new_[15993]_  | \new_[18832]_ ;
  assign \new_[14354]_  = ~\new_[15985]_  | ~\new_[16123]_ ;
  assign \new_[14355]_  = \new_[16052]_  & \new_[21513]_ ;
  assign \new_[14356]_  = ~\new_[16092]_  | ~\new_[19044]_ ;
  assign \new_[14357]_  = ~\new_[15359]_ ;
  assign \new_[14358]_  = ~\new_[15360]_ ;
  assign \new_[14359]_  = ~\new_[19779]_  | ~\new_[16318]_ ;
  assign \new_[14360]_  = ~\new_[14937]_ ;
  assign \new_[14361]_  = ~\new_[15928]_  & ~\new_[19013]_ ;
  assign \new_[14362]_  = \new_[17954]_  & \new_[16388]_ ;
  assign \new_[14363]_  = ~\new_[16501]_  | ~\new_[19096]_ ;
  assign \new_[14364]_  = \new_[15959]_  | \new_[18731]_ ;
  assign \new_[14365]_  = ~\new_[16039]_  & ~\new_[21513]_ ;
  assign \new_[14366]_  = ~\new_[14923]_ ;
  assign \new_[14367]_  = ~\new_[15336]_ ;
  assign \new_[14368]_  = ~\new_[15991]_  & ~\new_[18928]_ ;
  assign \new_[14369]_  = ~\new_[15366]_ ;
  assign \new_[14370]_  = ~\new_[16522]_  | ~\new_[18817]_ ;
  assign \new_[14371]_  = ~\new_[14959]_ ;
  assign \new_[14372]_  = ~\new_[15367]_ ;
  assign \new_[14373]_  = \new_[16537]_  | \new_[19815]_ ;
  assign \new_[14374]_  = ~\new_[18222]_  | ~\new_[16457]_ ;
  assign \new_[14375]_  = ~\new_[14929]_ ;
  assign \new_[14376]_  = ~\new_[18322]_  | ~\new_[16347]_ ;
  assign \new_[14377]_  = ~\new_[14897]_ ;
  assign \new_[14378]_  = ~\new_[17746]_  | ~\new_[19425]_ ;
  assign \new_[14379]_  = ~\new_[15313]_ ;
  assign \new_[14380]_  = \new_[15942]_  | \new_[18508]_ ;
  assign \new_[14381]_  = ~\new_[14886]_ ;
  assign \new_[14382]_  = ~\new_[14885]_ ;
  assign \new_[14383]_  = ~\new_[16156]_  & ~\new_[19084]_ ;
  assign \new_[14384]_  = ~\new_[17416]_  | (~\new_[17529]_  & ~\new_[21519]_ );
  assign \new_[14385]_  = ~\new_[14871]_ ;
  assign \new_[14386]_  = ~\new_[14870]_ ;
  assign \new_[14387]_  = ~\new_[15372]_ ;
  assign \new_[14388]_  = ~\new_[16243]_ ;
  assign \new_[14389]_  = ~\new_[16582]_  | ~\new_[19071]_ ;
  assign \new_[14390]_  = \new_[16093]_  & \new_[15887]_ ;
  assign \new_[14391]_  = ~\new_[14817]_ ;
  assign \new_[14392]_  = ~\new_[17600]_  | ~\new_[21695]_ ;
  assign \new_[14393]_  = ~\new_[14712]_ ;
  assign \new_[14394]_  = ~\new_[16021]_  | ~\new_[16380]_ ;
  assign \new_[14395]_  = ~\new_[16345]_  & ~\new_[19151]_ ;
  assign \new_[14396]_  = ~\new_[16291]_  & ~\new_[17452]_ ;
  assign \new_[14397]_  = ~\new_[17481]_  & ~\new_[21056]_ ;
  assign \new_[14398]_  = ~\new_[16562]_  | ~\new_[21507]_ ;
  assign \new_[14399]_  = ~\new_[16415]_  | ~\new_[17113]_ ;
  assign \new_[14400]_  = ~\new_[16176]_  & ~\new_[19687]_ ;
  assign \new_[14401]_  = \new_[16312]_  | \new_[19711]_ ;
  assign \new_[14402]_  = \new_[18170]_  | \new_[16676]_ ;
  assign \new_[14403]_  = ~\new_[17955]_  | ~\new_[15887]_ ;
  assign \new_[14404]_  = \new_[16167]_  | \new_[16126]_ ;
  assign \new_[14405]_  = ~\new_[17773]_  | ~\new_[16136]_ ;
  assign \new_[14406]_  = ~\new_[18403]_  | (~\new_[19234]_  & ~\new_[17556]_ );
  assign \new_[14407]_  = ~\new_[19155]_  | ~\new_[16545]_ ;
  assign \new_[14408]_  = ~\new_[16620]_  | (~\new_[18382]_  & ~\new_[19116]_ );
  assign \new_[14409]_  = ~\new_[16660]_  | (~\new_[17552]_  & ~\new_[19039]_ );
  assign \new_[14410]_  = ~\new_[18816]_  | ~\new_[16540]_ ;
  assign \new_[14411]_  = ~\new_[17063]_  & (~\new_[17933]_  | ~\new_[21609]_ );
  assign \new_[14412]_  = ~\new_[17726]_  | ~\new_[19555]_ ;
  assign \new_[14413]_  = ~\new_[16397]_  | (~\new_[18182]_  & ~\new_[19478]_ );
  assign \new_[14414]_  = ~\new_[15019]_ ;
  assign \new_[14415]_  = ~\new_[18460]_  & (~\new_[18128]_  | ~\new_[18283]_ );
  assign \new_[14416]_  = ~\new_[16479]_  | ~\new_[17840]_ ;
  assign \new_[14417]_  = ~\new_[16340]_  | ~\new_[16985]_ ;
  assign \new_[14418]_  = ~\new_[16494]_  | ~\new_[17468]_ ;
  assign \new_[14419]_  = ~\new_[16505]_  | ~\new_[18184]_ ;
  assign \new_[14420]_  = ~\new_[15162]_ ;
  assign \new_[14421]_  = ~\new_[16255]_  & (~\new_[19098]_  | ~\new_[18772]_ );
  assign \new_[14422]_  = ~\new_[14933]_ ;
  assign \new_[14423]_  = ~\new_[16006]_  & (~\new_[18179]_  | ~\new_[17482]_ );
  assign \new_[14424]_  = ~\new_[15161]_ ;
  assign \new_[14425]_  = ~\new_[16543]_  & (~\new_[19413]_  | ~\new_[18068]_ );
  assign \new_[14426]_  = ~\new_[15976]_  | ~\new_[18692]_ ;
  assign \new_[14427]_  = ~\new_[20242]_  & ~\new_[18443]_ ;
  assign \new_[14428]_  = ~\new_[15141]_ ;
  assign \new_[14429]_  = ~\new_[16048]_  & ~\new_[19217]_ ;
  assign \new_[14430]_  = ~\new_[16350]_  | ~\new_[19385]_ ;
  assign \new_[14431]_  = ~\new_[15938]_  | ~\new_[18012]_ ;
  assign \new_[14432]_  = \new_[18007]_  | \new_[17472]_ ;
  assign \new_[14433]_  = ~\new_[14957]_ ;
  assign \new_[14434]_  = ~\new_[16570]_  | ~\new_[19367]_ ;
  assign \new_[14435]_  = ~\new_[15706]_ ;
  assign \new_[14436]_  = ~\new_[17773]_  | ~\new_[16617]_ ;
  assign \new_[14437]_  = ~\new_[16627]_  | ~\new_[18371]_ ;
  assign \new_[14438]_  = ~\new_[15841]_ ;
  assign \new_[14439]_  = ~\new_[15413]_ ;
  assign \new_[14440]_  = ~\new_[16648]_  | ~\new_[21513]_ ;
  assign \new_[14441]_  = ~\new_[16213]_  & ~\new_[19094]_ ;
  assign \new_[14442]_  = ~\new_[15427]_ ;
  assign \new_[14443]_  = \new_[15876]_  | \new_[19538]_ ;
  assign \new_[14444]_  = ~\new_[15429]_ ;
  assign \new_[14445]_  = ~\new_[16426]_  & ~\new_[19053]_ ;
  assign \new_[14446]_  = ~\new_[15431]_ ;
  assign \new_[14447]_  = ~\new_[15996]_  | ~\new_[19741]_ ;
  assign \new_[14448]_  = ~\new_[15432]_ ;
  assign \new_[14449]_  = ~\new_[16304]_  | ~\new_[18558]_ ;
  assign \new_[14450]_  = \new_[15999]_  | \new_[19208]_ ;
  assign \new_[14451]_  = ~\new_[16282]_  | ~\new_[15892]_ ;
  assign \new_[14452]_  = ~\new_[15456]_ ;
  assign \new_[14453]_  = ~\new_[14693]_ ;
  assign \new_[14454]_  = ~\new_[14710]_ ;
  assign \new_[14455]_  = ~\new_[18598]_  | ~\new_[15989]_ ;
  assign \new_[14456]_  = ~\new_[15852]_ ;
  assign \new_[14457]_  = ~\new_[16577]_  | ~\new_[19434]_ ;
  assign \new_[14458]_  = ~\new_[15704]_ ;
  assign \new_[14459]_  = ~\new_[17137]_  & ~\new_[16622]_ ;
  assign \new_[14460]_  = ~\new_[15461]_ ;
  assign \new_[14461]_  = ~\new_[15820]_ ;
  assign \new_[14462]_  = ~\new_[15462]_ ;
  assign \new_[14463]_  = ~\new_[15979]_  & ~\new_[18926]_ ;
  assign \new_[14464]_  = ~\new_[15784]_ ;
  assign \new_[14465]_  = ~\new_[15464]_ ;
  assign \new_[14466]_  = ~\new_[16041]_  & ~\new_[18810]_ ;
  assign \new_[14467]_  = ~\new_[15751]_ ;
  assign \new_[14468]_  = ~\new_[16049]_  & ~\new_[17444]_ ;
  assign \new_[14469]_  = \new_[15446]_ ;
  assign \new_[14470]_  = ~\new_[15404]_ ;
  assign \new_[14471]_  = ~\new_[15256]_ ;
  assign \new_[14472]_  = ~\new_[17716]_  | ~\new_[19031]_ ;
  assign \new_[14473]_  = ~\new_[16578]_  & ~\new_[19269]_ ;
  assign \new_[14474]_  = ~\new_[15197]_ ;
  assign \new_[14475]_  = ~\new_[15007]_ ;
  assign \new_[14476]_  = ~\new_[14847]_ ;
  assign \new_[14477]_  = ~\new_[15173]_ ;
  assign \new_[14478]_  = ~\new_[15151]_ ;
  assign \new_[14479]_  = ~\new_[15619]_ ;
  assign \new_[14480]_  = ~\new_[15937]_  & ~\new_[16152]_ ;
  assign \new_[14481]_  = ~\new_[18012]_  | ~\new_[21631]_  | ~\new_[17387]_ ;
  assign \new_[14482]_  = ~\new_[15489]_ ;
  assign \new_[14483]_  = ~\new_[15024]_ ;
  assign \new_[14484]_  = ~\new_[15492]_ ;
  assign \new_[14485]_  = ~\new_[18938]_  | ~\new_[17852]_  | ~\new_[18179]_ ;
  assign \new_[14486]_  = \new_[18913]_  | \new_[17644]_ ;
  assign \new_[14487]_  = ~\new_[14726]_ ;
  assign \new_[14488]_  = ~\new_[15503]_ ;
  assign \new_[14489]_  = ~\new_[15508]_ ;
  assign \new_[14490]_  = ~\new_[15513]_ ;
  assign \new_[14491]_  = ~\new_[15517]_ ;
  assign \new_[14492]_  = ~\new_[15869]_  | ~\new_[18794]_ ;
  assign \new_[14493]_  = ~\new_[14834]_ ;
  assign \new_[14494]_  = ~\new_[15876]_  | ~\new_[17516]_ ;
  assign \new_[14495]_  = ~\new_[16013]_  & ~\new_[18810]_ ;
  assign \new_[14496]_  = ~\new_[14821]_ ;
  assign \new_[14497]_  = ~\new_[15541]_ ;
  assign \new_[14498]_  = ~\new_[15526]_ ;
  assign \new_[14499]_  = ~\new_[18783]_  | ~\new_[16622]_ ;
  assign \new_[14500]_  = ~\new_[14774]_ ;
  assign \new_[14501]_  = ~\new_[15529]_ ;
  assign \new_[14502]_  = ~\new_[14748]_ ;
  assign \new_[14503]_  = ~\new_[16598]_  | ~\new_[21259]_ ;
  assign \new_[14504]_  = \new_[19169]_  | \new_[16026]_ ;
  assign \new_[14505]_  = \new_[19027]_  | \new_[16093]_ ;
  assign \new_[14506]_  = ~\new_[15934]_  & ~\new_[19681]_ ;
  assign \new_[14507]_  = ~\new_[15543]_ ;
  assign \new_[14508]_  = ~\new_[17362]_  | ~\new_[17886]_ ;
  assign \new_[14509]_  = ~\new_[15548]_ ;
  assign \new_[14510]_  = ~\new_[15806]_ ;
  assign \new_[14511]_  = ~\new_[16002]_  | ~\new_[18111]_ ;
  assign \new_[14512]_  = ~\new_[18771]_  | ~\new_[17619]_ ;
  assign \new_[14513]_  = ~\new_[15664]_ ;
  assign \new_[14514]_  = ~\new_[15847]_ ;
  assign \new_[14515]_  = ~\new_[17402]_  | ~\new_[17499]_ ;
  assign \new_[14516]_  = ~\new_[15451]_ ;
  assign \new_[14517]_  = ~\new_[18270]_  | ~\new_[16623]_ ;
  assign \new_[14518]_  = \new_[16592]_  | \new_[18811]_ ;
  assign \new_[14519]_  = ~\new_[15574]_ ;
  assign \new_[14520]_  = ~\new_[15576]_ ;
  assign \new_[14521]_  = ~\new_[18060]_  | ~\new_[19357]_  | ~\new_[19379]_ ;
  assign \new_[14522]_  = ~\new_[14904]_ ;
  assign \new_[14523]_  = \new_[18809]_  | \new_[16512]_ ;
  assign \new_[14524]_  = ~\new_[17991]_  | ~\new_[17941]_ ;
  assign \new_[14525]_  = ~\new_[14883]_ ;
  assign \new_[14526]_  = ~\new_[16027]_ ;
  assign \new_[14527]_  = ~\new_[14862]_ ;
  assign \new_[14528]_  = ~\new_[16619]_  | ~\new_[16982]_ ;
  assign \new_[14529]_  = ~\new_[17588]_  | ~\new_[17671]_ ;
  assign \new_[14530]_  = ~\new_[17662]_  | ~\new_[19217]_ ;
  assign \new_[14531]_  = \new_[19255]_  | \new_[17747]_ ;
  assign \new_[14532]_  = ~\new_[16038]_  | ~\new_[20865]_ ;
  assign \new_[14533]_  = ~\new_[14849]_ ;
  assign \new_[14534]_  = ~\new_[16002]_  | ~\new_[21056]_ ;
  assign \new_[14535]_  = ~\new_[14811]_ ;
  assign \new_[14536]_  = ~\new_[15596]_ ;
  assign \new_[14537]_  = ~\new_[15600]_ ;
  assign \new_[14538]_  = ~\new_[15601]_ ;
  assign \new_[14539]_  = \new_[16046]_  | \new_[21306]_ ;
  assign \new_[14540]_  = ~\new_[17888]_  & ~\new_[18692]_ ;
  assign \new_[14541]_  = ~\new_[14724]_ ;
  assign \new_[14542]_  = ~\new_[19156]_  | ~\new_[18310]_  | ~\new_[19098]_ ;
  assign \new_[14543]_  = ~\new_[15560]_ ;
  assign \new_[14544]_  = ~\new_[15864]_ ;
  assign \new_[14545]_  = ~\new_[17359]_  | ~\new_[16652]_ ;
  assign \new_[14546]_  = ~\new_[15859]_ ;
  assign \new_[14547]_  = ~\new_[16618]_  | ~\new_[17457]_ ;
  assign \new_[14548]_  = \new_[16634]_  | \new_[19538]_ ;
  assign \new_[14549]_  = ~\new_[15611]_ ;
  assign \new_[14550]_  = ~\new_[15613]_ ;
  assign \new_[14551]_  = \new_[17862]_  | \new_[18007]_ ;
  assign \new_[14552]_  = \new_[17791]_  | \new_[17534]_ ;
  assign \new_[14553]_  = ~\new_[16611]_  | ~\new_[19088]_ ;
  assign \new_[14554]_  = \new_[17557]_  & \new_[16980]_ ;
  assign \new_[14555]_  = ~\new_[17648]_  & ~\new_[18424]_ ;
  assign \new_[14556]_  = ~\new_[17546]_  | ~\new_[18061]_ ;
  assign \new_[14557]_  = ~\new_[16644]_  & ~\new_[19681]_ ;
  assign \new_[14558]_  = ~\new_[15685]_ ;
  assign \new_[14559]_  = ~\new_[17919]_  | ~\new_[18012]_ ;
  assign \new_[14560]_  = ~\new_[19822]_  | ~\new_[17884]_ ;
  assign \new_[14561]_  = ~\new_[14714]_ ;
  assign \new_[14562]_  = ~\new_[17155]_  | ~\new_[18124]_  | ~\new_[19444]_ ;
  assign \new_[14563]_  = ~\new_[19016]_  | ~\new_[17644]_ ;
  assign \new_[14564]_  = ~\new_[15145]_ ;
  assign \new_[14565]_  = \new_[18442]_  | \new_[18014]_ ;
  assign \new_[14566]_  = ~\new_[15269]_ ;
  assign \new_[14567]_  = ~\new_[15866]_ ;
  assign \new_[14568]_  = ~\new_[16679]_  & ~\new_[18621]_ ;
  assign \new_[14569]_  = ~\new_[15758]_ ;
  assign \new_[14570]_  = ~\new_[15631]_ ;
  assign \new_[14571]_  = ~\new_[16791]_  & ~\new_[19088]_ ;
  assign \new_[14572]_  = ~\new_[16605]_  | ~\new_[18863]_ ;
  assign \new_[14573]_  = \new_[16649]_  | \new_[19386]_ ;
  assign \new_[14574]_  = ~\new_[14854]_ ;
  assign \new_[14575]_  = ~\new_[16017]_  & ~\new_[18166]_ ;
  assign \new_[14576]_  = ~\new_[14879]_ ;
  assign \new_[14577]_  = ~\new_[14867]_ ;
  assign \new_[14578]_  = ~\new_[14857]_ ;
  assign \new_[14579]_  = \new_[18992]_  | \new_[15894]_ ;
  assign \new_[14580]_  = ~\new_[16611]_  | ~\new_[18166]_ ;
  assign \new_[14581]_  = \new_[17776]_  & \new_[18747]_ ;
  assign \new_[14582]_  = ~\new_[14824]_ ;
  assign \new_[14583]_  = ~\new_[15731]_ ;
  assign \new_[14584]_  = ~\new_[17578]_  | ~\new_[16658]_  | ~\new_[18465]_ ;
  assign \new_[14585]_  = ~\new_[16018]_  | ~\new_[20699]_ ;
  assign \new_[14586]_  = ~\new_[15954]_  | ~\new_[18179]_ ;
  assign \new_[14587]_  = ~\new_[15775]_ ;
  assign \new_[14588]_  = ~\new_[15248]_ ;
  assign \new_[14589]_  = ~\new_[16619]_  | ~\new_[18814]_ ;
  assign \new_[14590]_  = ~\new_[16618]_  | ~\new_[18778]_ ;
  assign \new_[14591]_  = ~\new_[16484]_  | ~\new_[19117]_ ;
  assign \new_[14592]_  = ~\new_[15648]_ ;
  assign \new_[14593]_  = ~\new_[15026]_ ;
  assign \new_[14594]_  = ~\new_[15573]_ ;
  assign \new_[14595]_  = ~\new_[15442]_ ;
  assign \new_[14596]_  = ~\new_[15428]_ ;
  assign \new_[14597]_  = ~\new_[15581]_ ;
  assign \new_[14598]_  = ~\new_[15669]_ ;
  assign \new_[14599]_  = ~\new_[15680]_ ;
  assign \new_[14600]_  = ~\new_[15245]_ ;
  assign \new_[14601]_  = ~\new_[17588]_  | ~\new_[17425]_ ;
  assign \new_[14602]_  = ~\new_[14815]_ ;
  assign \new_[14603]_  = ~\new_[16007]_ ;
  assign \new_[14604]_  = ~\new_[16621]_  | ~\new_[19249]_ ;
  assign \new_[14605]_  = ~\new_[16599]_  | ~\new_[21574]_ ;
  assign \new_[14606]_  = ~\new_[15558]_ ;
  assign \new_[14607]_  = ~\new_[15690]_ ;
  assign \new_[14608]_  = ~\new_[15800]_ ;
  assign \new_[14609]_  = ~\new_[17217]_ ;
  assign \new_[14610]_  = ~\new_[14742]_ ;
  assign \new_[14611]_  = ~\new_[15753]_ ;
  assign \new_[14612]_  = ~\new_[17631]_  & ~\new_[19196]_ ;
  assign \new_[14613]_  = ~\new_[14865]_ ;
  assign \new_[14614]_  = ~\new_[17680]_  | ~\new_[19290]_ ;
  assign \new_[14615]_  = ~\new_[16273]_  | ~\new_[19096]_ ;
  assign \new_[14616]_  = ~\new_[15351]_ ;
  assign \new_[14617]_  = ~\new_[15957]_  | ~\new_[19689]_ ;
  assign \new_[14618]_  = ~\new_[15713]_ ;
  assign \new_[14619]_  = ~\new_[17557]_  | ~\new_[18750]_ ;
  assign \new_[14620]_  = ~\new_[15722]_ ;
  assign \new_[14621]_  = ~\new_[17347]_  | ~\new_[16608]_ ;
  assign \new_[14622]_  = ~\new_[15981]_  | ~\new_[17951]_ ;
  assign \new_[14623]_  = ~\new_[16018]_  & ~\new_[21608]_ ;
  assign \new_[14624]_  = ~\new_[14873]_ ;
  assign \new_[14625]_  = ~\new_[16595]_  | ~\new_[17348]_ ;
  assign \new_[14626]_  = ~\new_[17667]_  | ~\new_[16528]_ ;
  assign \new_[14627]_  = ~\new_[17428]_  | ~\new_[16662]_ ;
  assign \new_[14628]_  = ~\new_[17355]_  & ~\new_[16623]_ ;
  assign \new_[14629]_  = ~\new_[15078]_ ;
  assign \new_[14630]_  = ~\new_[15735]_ ;
  assign \new_[14631]_  = ~\new_[16619]_  | ~\new_[17614]_ ;
  assign \new_[14632]_  = ~\new_[17955]_  | ~\new_[16093]_ ;
  assign \new_[14633]_  = ~\new_[17710]_  | ~\new_[16625]_ ;
  assign \new_[14634]_  = ~\new_[15746]_ ;
  assign \new_[14635]_  = \new_[17939]_  & \new_[17941]_ ;
  assign \new_[14636]_  = ~\new_[18239]_  | (~\new_[18179]_  & ~\new_[19513]_ );
  assign \new_[14637]_  = ~\new_[16790]_  & ~\new_[16627]_ ;
  assign \new_[14638]_  = ~\new_[16642]_  | (~\new_[18575]_  & ~\new_[19647]_ );
  assign \new_[14639]_  = ~\new_[16492]_  & ~\new_[21565]_ ;
  assign \new_[14640]_  = ~\new_[17581]_  | (~\new_[18553]_  & ~\new_[17425]_ );
  assign n2753 = ~\new_[18775]_  | (~\new_[17309]_  & ~\new_[19723]_ );
  assign \new_[14642]_  = ~\new_[15866]_  | ~\new_[19048]_ ;
  assign \new_[14643]_  = ~\new_[15752]_ ;
  assign \new_[14644]_  = ~\new_[15618]_ ;
  assign \new_[14645]_  = ~\new_[16107]_  & ~\new_[19095]_ ;
  assign \new_[14646]_  = ~\new_[15902]_  | ~\new_[20924]_ ;
  assign \new_[14647]_  = \new_[17544]_  & \new_[17499]_ ;
  assign \new_[14648]_  = ~\new_[17702]_  | ~\new_[18020]_ ;
  assign \new_[14649]_  = \new_[19666]_  ^ \new_[18464]_ ;
  assign \new_[14650]_  = \new_[19616]_  ^ \new_[16980]_ ;
  assign \new_[14651]_  = ~\new_[16526]_  | ~\new_[21306]_ ;
  assign \new_[14652]_  = ~\new_[15658]_ ;
  assign \new_[14653]_  = \new_[19651]_  ^ \new_[16682]_ ;
  assign \new_[14654]_  = \new_[16995]_  ^ \new_[18025]_ ;
  assign \new_[14655]_  = \new_[16260]_  | \new_[18678]_ ;
  assign \new_[14656]_  = ~\new_[15786]_ ;
  assign \new_[14657]_  = ~\new_[14969]_ ;
  assign \new_[14658]_  = ~\new_[14969]_ ;
  assign \new_[14659]_  = ~\new_[15783]_ ;
  assign \new_[14660]_  = ~\new_[15694]_ ;
  assign \new_[14661]_  = \new_[16676]_  & \new_[19425]_ ;
  assign \new_[14662]_  = \new_[17550]_  | \new_[19269]_ ;
  assign \new_[14663]_  = ~\new_[14940]_ ;
  assign \new_[14664]_  = ~\new_[16451]_  | ~\new_[19801]_ ;
  assign \new_[14665]_  = ~\new_[15794]_ ;
  assign \new_[14666]_  = ~\new_[20663]_  | ~\new_[21686]_ ;
  assign \new_[14667]_  = ~\new_[15799]_ ;
  assign \new_[14668]_  = \new_[16617]_  & \new_[16136]_ ;
  assign \new_[14669]_  = ~\new_[15654]_ ;
  assign \new_[14670]_  = \new_[18486]_  & \new_[15949]_ ;
  assign \new_[14671]_  = \new_[16612]_  | \new_[19097]_ ;
  assign \new_[14672]_  = \new_[17850]_  | \new_[19253]_ ;
  assign \new_[14673]_  = \new_[15953]_  | \new_[19181]_ ;
  assign \new_[14674]_  = ~\new_[15614]_ ;
  assign \new_[14675]_  = ~\new_[15817]_ ;
  assign \new_[14676]_  = ~\new_[15821]_ ;
  assign \new_[14677]_  = ~\new_[16044]_  | ~\new_[18987]_ ;
  assign \new_[14678]_  = ~\new_[15811]_ ;
  assign \new_[14679]_  = ~\new_[15830]_ ;
  assign \new_[14680]_  = ~\new_[16589]_  | ~\new_[19665]_ ;
  assign \new_[14681]_  = ~\new_[15961]_  & ~\new_[19050]_ ;
  assign \new_[14682]_  = ~\new_[16186]_  & ~\new_[19095]_ ;
  assign \new_[14683]_  = ~\new_[16600]_  | ~\new_[19044]_ ;
  assign \new_[14684]_  = \new_[16312]_  & \new_[16307]_ ;
  assign \new_[14685]_  = ~\new_[15542]_ ;
  assign \new_[14686]_  = ~\new_[15609]_ ;
  assign \new_[14687]_  = ~\new_[16087]_  | ~\new_[18947]_ ;
  assign \new_[14688]_  = ~\new_[15857]_ ;
  assign \new_[14689]_  = ~\new_[18931]_  & ~\new_[17680]_ ;
  assign \new_[14690]_  = ~\new_[18935]_ ;
  assign \new_[14691]_  = ~\new_[15655]_ ;
  assign \new_[14692]_  = ~\new_[18140]_  | ~\new_[19535]_ ;
  assign \new_[14693]_  = ~\new_[17453]_  | ~\new_[20865]_ ;
  assign \new_[14694]_  = \new_[18923]_  | \new_[17338]_ ;
  assign \new_[14695]_  = ~\new_[16768]_  & ~\new_[19117]_ ;
  assign \new_[14696]_  = \\text_in_r_reg[116] ;
  assign \new_[14697]_  = \\text_in_r_reg[111] ;
  assign \new_[14698]_  = \\text_in_r_reg[37] ;
  assign \new_[14699]_  = ~\new_[17052]_  & ~\new_[19655]_ ;
  assign \new_[14700]_  = \\text_in_r_reg[14] ;
  assign \new_[14701]_  = \\text_in_r_reg[67] ;
  assign \new_[14702]_  = \\text_in_r_reg[47] ;
  assign \new_[14703]_  = ~\new_[15874]_ ;
  assign \new_[14704]_  = ~\new_[18585]_  | ~\new_[19039]_ ;
  assign \new_[14705]_  = ~\new_[15875]_ ;
  assign \new_[14706]_  = ~\new_[15876]_ ;
  assign \new_[14707]_  = ~\new_[21398]_ ;
  assign \new_[14708]_  = ~\new_[16570]_ ;
  assign \new_[14709]_  = \\text_in_r_reg[18] ;
  assign \new_[14710]_  = ~\new_[15881]_ ;
  assign \new_[14711]_  = \\text_in_r_reg[0] ;
  assign \new_[14712]_  = ~\new_[16504]_ ;
  assign \new_[14713]_  = ~\new_[17170]_  & ~\new_[19068]_ ;
  assign \new_[14714]_  = ~\new_[16983]_  | ~\new_[18968]_ ;
  assign \new_[14715]_  = ~\new_[16253]_ ;
  assign \new_[14716]_  = ~\new_[17553]_  & ~\new_[19156]_ ;
  assign \new_[14717]_  = ~\new_[15975]_ ;
  assign \new_[14718]_  = \new_[15889]_ ;
  assign \new_[14719]_  = \\text_in_r_reg[68] ;
  assign \new_[14720]_  = ~\new_[15890]_ ;
  assign \new_[14721]_  = \new_[17222]_  | \new_[19636]_ ;
  assign \new_[14722]_  = \\text_in_r_reg[49] ;
  assign \new_[14723]_  = ~\new_[17971]_  | ~\new_[17387]_ ;
  assign \new_[14724]_  = ~\new_[16747]_  & ~\new_[18966]_ ;
  assign \new_[14725]_  = \\text_in_r_reg[42] ;
  assign \new_[14726]_  = ~\new_[17289]_  & ~\new_[19096]_ ;
  assign \new_[14727]_  = ~\new_[16073]_ ;
  assign \new_[14728]_  = ~\new_[15897]_ ;
  assign \new_[14729]_  = \new_[17007]_  | \new_[18709]_ ;
  assign \new_[14730]_  = ~\new_[18179]_  | ~\new_[18449]_ ;
  assign \new_[14731]_  = ~\new_[16389]_ ;
  assign \new_[14732]_  = ~\new_[17574]_  | ~\new_[21520]_ ;
  assign \new_[14733]_  = \new_[17077]_  & \new_[19675]_ ;
  assign \new_[14734]_  = ~\new_[16257]_ ;
  assign \new_[14735]_  = ~\new_[16986]_  & ~\new_[18325]_ ;
  assign \new_[14736]_  = ~\new_[17287]_  & ~\new_[19268]_ ;
  assign \new_[14737]_  = ~\new_[16163]_ ;
  assign \new_[14738]_  = ~\new_[16734]_ ;
  assign \new_[14739]_  = ~\new_[19741]_  & ~\new_[16769]_ ;
  assign \new_[14740]_  = ~\new_[17371]_  & ~\new_[19801]_ ;
  assign \new_[14741]_  = ~\new_[16929]_  | ~\new_[19096]_ ;
  assign \new_[14742]_  = ~\new_[16792]_  | ~\new_[18810]_ ;
  assign \new_[14743]_  = ~\new_[15905]_ ;
  assign \new_[14744]_  = ~\new_[16232]_ ;
  assign \new_[14745]_  = ~\new_[17328]_  & ~\new_[17643]_ ;
  assign \new_[14746]_  = ~\new_[15906]_ ;
  assign \new_[14747]_  = ~\new_[19026]_  & ~\new_[16829]_ ;
  assign \new_[14748]_  = ~\new_[16788]_  & ~\new_[18408]_ ;
  assign \new_[14749]_  = ~\new_[18813]_  & ~\new_[17237]_ ;
  assign \new_[14750]_  = \\text_in_r_reg[127] ;
  assign \new_[14751]_  = ~\new_[16333]_ ;
  assign \new_[14752]_  = \\text_in_r_reg[64] ;
  assign \new_[14753]_  = \\text_in_r_reg[54] ;
  assign \new_[14754]_  = \new_[16902]_  | \new_[19265]_ ;
  assign \new_[14755]_  = \\text_in_r_reg[35] ;
  assign \new_[14756]_  = \\text_in_r_reg[6] ;
  assign \new_[14757]_  = ~\new_[16433]_ ;
  assign \new_[14758]_  = \\text_in_r_reg[17] ;
  assign \new_[14759]_  = \\text_in_r_reg[108] ;
  assign \new_[14760]_  = \\text_in_r_reg[11] ;
  assign \new_[14761]_  = \\text_in_r_reg[123] ;
  assign \new_[14762]_  = \\text_in_r_reg[24] ;
  assign \new_[14763]_  = \\text_in_r_reg[26] ;
  assign \new_[14764]_  = \\text_in_r_reg[29] ;
  assign \new_[14765]_  = \\text_in_r_reg[46] ;
  assign \new_[14766]_  = \\text_in_r_reg[55] ;
  assign \new_[14767]_  = \\text_in_r_reg[61] ;
  assign \new_[14768]_  = \\text_in_r_reg[63] ;
  assign \new_[14769]_  = \\text_in_r_reg[78] ;
  assign \new_[14770]_  = \\text_in_r_reg[81] ;
  assign \new_[14771]_  = \\text_in_r_reg[86] ;
  assign \new_[14772]_  = \\text_in_r_reg[8] ;
  assign \new_[14773]_  = \\text_in_r_reg[99] ;
  assign \new_[14774]_  = \new_[15912]_ ;
  assign \new_[14775]_  = \new_[19156]_  & \new_[19578]_ ;
  assign \new_[14776]_  = \\text_in_r_reg[91] ;
  assign \new_[14777]_  = \\text_in_r_reg[39] ;
  assign \new_[14778]_  = \\text_in_r_reg[60] ;
  assign \new_[14779]_  = \\text_in_r_reg[103] ;
  assign \new_[14780]_  = \\text_in_r_reg[23] ;
  assign \new_[14781]_  = \\text_in_r_reg[58] ;
  assign \new_[14782]_  = \\text_in_r_reg[3] ;
  assign \new_[14783]_  = ~\new_[16426]_ ;
  assign \new_[14784]_  = ~\new_[17438]_  | ~\new_[21115]_ ;
  assign \new_[14785]_  = ~\new_[18715]_  | ~\new_[17270]_  | ~\new_[18113]_ ;
  assign \new_[14786]_  = \new_[17181]_  | \new_[19088]_ ;
  assign \new_[14787]_  = ~\new_[17270]_  & ~\new_[18113]_ ;
  assign \new_[14788]_  = \\text_in_r_reg[118] ;
  assign \new_[14789]_  = ~\new_[16600]_ ;
  assign \new_[14790]_  = \\text_in_r_reg[59] ;
  assign \new_[14791]_  = ~\new_[15936]_ ;
  assign \new_[14792]_  = ~\new_[17324]_  | ~\new_[20490]_ ;
  assign \new_[14793]_  = \\text_in_r_reg[96] ;
  assign \new_[14794]_  = ~\new_[17382]_  | ~\new_[19217]_ ;
  assign \new_[14795]_  = ~\new_[16278]_ ;
  assign \new_[14796]_  = ~\new_[17142]_  & ~\new_[19198]_ ;
  assign \new_[14797]_  = ~\new_[18909]_  | ~\new_[17189]_ ;
  assign \new_[14798]_  = ~\new_[15940]_ ;
  assign \new_[14799]_  = \\text_in_r_reg[70] ;
  assign \new_[14800]_  = \new_[17340]_  | \new_[18794]_ ;
  assign \new_[14801]_  = ~\new_[16815]_  & ~\new_[19085]_ ;
  assign \new_[14802]_  = ~\new_[15942]_ ;
  assign \new_[14803]_  = ~\new_[17316]_  & ~\new_[19555]_ ;
  assign \new_[14804]_  = ~\new_[16432]_ ;
  assign \new_[14805]_  = ~\new_[18570]_  | ~\new_[18253]_ ;
  assign \new_[14806]_  = ~\new_[17313]_  | ~\new_[19782]_ ;
  assign \new_[14807]_  = ~\new_[17137]_  | ~\new_[19096]_ ;
  assign \new_[14808]_  = ~\new_[17251]_  & ~\new_[19637]_ ;
  assign \new_[14809]_  = ~\new_[16803]_  | ~\new_[19220]_ ;
  assign \new_[14810]_  = ~\new_[20494]_  | ~\new_[18974]_ ;
  assign \new_[14811]_  = ~\new_[17355]_  | ~\new_[19270]_ ;
  assign \new_[14812]_  = ~\new_[16496]_ ;
  assign \new_[14813]_  = ~\new_[17066]_ ;
  assign \new_[14814]_  = \\text_in_r_reg[51] ;
  assign \new_[14815]_  = ~\new_[16214]_ ;
  assign \new_[14816]_  = ~\new_[18264]_  & ~\new_[19151]_ ;
  assign \new_[14817]_  = ~\new_[16738]_  & ~\new_[19676]_ ;
  assign \new_[14818]_  = ~\new_[19053]_  & ~\new_[17417]_ ;
  assign \new_[14819]_  = ~\new_[15980]_ ;
  assign \new_[14820]_  = ~\new_[16703]_  & ~\new_[19161]_ ;
  assign \new_[14821]_  = ~\new_[15953]_ ;
  assign \new_[14822]_  = \new_[19215]_  & \new_[19623]_ ;
  assign \new_[14823]_  = \new_[17327]_  | \new_[18190]_ ;
  assign \new_[14824]_  = ~\new_[16476]_ ;
  assign \new_[14825]_  = ~\new_[15962]_ ;
  assign \new_[14826]_  = ~\new_[17582]_ ;
  assign \new_[14827]_  = ~\new_[15961]_ ;
  assign \new_[14828]_  = ~\new_[16178]_ ;
  assign \new_[14829]_  = ~\new_[16987]_  | ~\new_[19801]_ ;
  assign \new_[14830]_  = \new_[21396]_  & \new_[18485]_ ;
  assign \new_[14831]_  = ~\new_[17974]_  | ~\new_[17342]_ ;
  assign \new_[14832]_  = ~\new_[17292]_  | ~\new_[16871]_ ;
  assign \new_[14833]_  = ~\new_[18012]_  & ~\new_[16990]_ ;
  assign \new_[14834]_  = ~\new_[16379]_ ;
  assign \new_[14835]_  = ~\new_[16324]_ ;
  assign \new_[14836]_  = ~\new_[15965]_ ;
  assign \new_[14837]_  = ~\new_[21392]_ ;
  assign \new_[14838]_  = ~\new_[19459]_  & ~\new_[17351]_ ;
  assign \new_[14839]_  = ~\new_[16190]_ ;
  assign \new_[14840]_  = ~\new_[16475]_ ;
  assign \new_[14841]_  = ~\new_[15979]_ ;
  assign \new_[14842]_  = ~\new_[16155]_ ;
  assign \new_[14843]_  = ~\new_[16799]_  | ~\new_[19268]_ ;
  assign \new_[14844]_  = ~\new_[21259]_  & ~\new_[16765]_ ;
  assign \new_[14845]_  = \new_[17346]_  & \new_[19186]_ ;
  assign \new_[14846]_  = ~\new_[16259]_ ;
  assign \new_[14847]_  = \new_[16357]_ ;
  assign \new_[14848]_  = ~\new_[16250]_ ;
  assign \new_[14849]_  = \new_[19675]_  & \new_[16877]_ ;
  assign \new_[14850]_  = ~\new_[17045]_  & ~\new_[19446]_ ;
  assign \new_[14851]_  = \\text_in_r_reg[92] ;
  assign \new_[14852]_  = ~\new_[18459]_  | ~\new_[19398]_  | ~\new_[19446]_  | ~\new_[18857]_ ;
  assign \new_[14853]_  = ~\new_[16711]_  | ~\new_[19386]_ ;
  assign \new_[14854]_  = ~\new_[16994]_  | ~\new_[19251]_ ;
  assign \new_[14855]_  = \new_[18938]_  & \new_[19803]_ ;
  assign \new_[14856]_  = ~\new_[15993]_ ;
  assign \new_[14857]_  = ~\new_[19063]_  | ~\new_[17412]_ ;
  assign \new_[14858]_  = ~\new_[15997]_ ;
  assign \new_[14859]_  = ~\new_[15996]_ ;
  assign \new_[14860]_  = ~\new_[16000]_ ;
  assign \new_[14861]_  = \new_[16710]_  | \new_[18840]_ ;
  assign \new_[14862]_  = ~\new_[16423]_ ;
  assign \new_[14863]_  = ~\new_[21483]_  | ~\new_[19413]_  | ~\new_[19249]_  | ~\new_[17979]_ ;
  assign \new_[14864]_  = ~\new_[16935]_  | ~\new_[20927]_ ;
  assign \new_[14865]_  = ~\new_[16028]_ ;
  assign \new_[14866]_  = ~\new_[17446]_  | ~\new_[20927]_ ;
  assign \new_[14867]_  = ~\new_[16820]_  & ~\new_[18784]_ ;
  assign \new_[14868]_  = ~\new_[16909]_  & ~\new_[18621]_ ;
  assign \new_[14869]_  = ~\new_[16010]_ ;
  assign \new_[14870]_  = \new_[17263]_  & \new_[19145]_ ;
  assign \new_[14871]_  = ~\new_[17254]_  & ~\new_[20490]_ ;
  assign \new_[14872]_  = ~\new_[16470]_ ;
  assign \new_[14873]_  = ~\new_[17082]_  | ~\new_[17951]_ ;
  assign \new_[14874]_  = ~\new_[17396]_  & ~\new_[21306]_ ;
  assign \new_[14875]_  = ~\new_[18226]_  | ~\new_[19478]_  | ~\new_[19024]_  | ~\new_[19212]_ ;
  assign \new_[14876]_  = ~\new_[16708]_  | ~\new_[19024]_ ;
  assign \new_[14877]_  = \\text_in_r_reg[107] ;
  assign \new_[14878]_  = ~\new_[17296]_  | ~\new_[19319]_ ;
  assign \new_[14879]_  = ~\new_[16930]_  | ~\new_[19176]_ ;
  assign \new_[14880]_  = ~\new_[17200]_  | ~\new_[18750]_ ;
  assign \new_[14881]_  = ~\new_[16023]_ ;
  assign \new_[14882]_  = ~\new_[19371]_  & (~\new_[17566]_  | ~\new_[18113]_ );
  assign \new_[14883]_  = ~\new_[17147]_  | ~\new_[19062]_ ;
  assign \new_[14884]_  = ~\new_[18115]_  | ~\new_[16800]_ ;
  assign \new_[14885]_  = ~\new_[16993]_  & ~\new_[19426]_ ;
  assign \new_[14886]_  = ~\new_[17190]_  & ~\new_[21513]_ ;
  assign \new_[14887]_  = ~\new_[17269]_  & ~\new_[19044]_ ;
  assign \new_[14888]_  = ~\new_[17230]_  & ~\new_[18607]_ ;
  assign \new_[14889]_  = ~\new_[16032]_ ;
  assign \new_[14890]_  = ~\new_[16109]_ ;
  assign \new_[14891]_  = ~\new_[16149]_ ;
  assign \new_[14892]_  = ~\new_[18818]_  | ~\new_[17002]_ ;
  assign \new_[14893]_  = \\text_in_r_reg[28] ;
  assign \new_[14894]_  = ~\new_[16911]_  & ~\new_[19298]_ ;
  assign \new_[14895]_  = \new_[17071]_  | \new_[19189]_ ;
  assign \new_[14896]_  = ~\new_[19603]_  & ~\new_[19156]_ ;
  assign \new_[14897]_  = ~\new_[16825]_  | ~\new_[19754]_ ;
  assign \new_[14898]_  = \new_[18175]_  & \new_[17342]_ ;
  assign \new_[14899]_  = \\text_in_r_reg[77] ;
  assign \new_[14900]_  = ~\new_[16115]_ ;
  assign \new_[14901]_  = ~\new_[16949]_  | ~\new_[19553]_ ;
  assign \new_[14902]_  = \\text_in_r_reg[1] ;
  assign \new_[14903]_  = ~\new_[17772]_  | ~\new_[16745]_  | ~\new_[17576]_ ;
  assign \new_[14904]_  = ~\new_[16797]_  | ~\new_[16851]_ ;
  assign \new_[14905]_  = \\text_in_r_reg[19] ;
  assign \new_[14906]_  = ~\new_[16794]_  | ~\new_[18402]_ ;
  assign \new_[14907]_  = ~\new_[16078]_ ;
  assign \new_[14908]_  = ~\new_[17199]_  & ~\new_[19386]_ ;
  assign \new_[14909]_  = \\text_in_r_reg[56] ;
  assign \new_[14910]_  = ~\new_[18945]_  & ~\new_[16767]_ ;
  assign \new_[14911]_  = \new_[16683]_  | \new_[18285]_ ;
  assign \new_[14912]_  = \\text_in_r_reg[90] ;
  assign \new_[14913]_  = ~\new_[16873]_  | ~\new_[18832]_ ;
  assign \new_[14914]_  = ~\new_[15973]_ ;
  assign \new_[14915]_  = \new_[17138]_  | \new_[19727]_ ;
  assign \new_[14916]_  = ~\new_[16057]_ ;
  assign \new_[14917]_  = ~\new_[18945]_  & ~\new_[16784]_ ;
  assign \new_[14918]_  = \new_[19689]_  | \new_[20764]_ ;
  assign \new_[14919]_  = ~\new_[16867]_  | ~\new_[19156]_ ;
  assign \new_[14920]_  = \new_[18340]_  | \new_[18166]_ ;
  assign \new_[14921]_  = ~\new_[16063]_ ;
  assign \new_[14922]_  = \\text_in_r_reg[69] ;
  assign \new_[14923]_  = \new_[16719]_  | \new_[19476]_ ;
  assign \new_[14924]_  = ~\new_[16221]_ ;
  assign \new_[14925]_  = \new_[16734]_  | \new_[19061]_ ;
  assign \new_[14926]_  = ~\new_[16244]_ ;
  assign \new_[14927]_  = \new_[16937]_  | \new_[19636]_ ;
  assign \new_[14928]_  = ~\new_[17153]_  | ~\new_[19117]_ ;
  assign \new_[14929]_  = ~\new_[16686]_  & ~\new_[19100]_ ;
  assign \new_[14930]_  = \new_[19658]_  ^ \new_[18757]_ ;
  assign \new_[14931]_  = ~\new_[19150]_  & ~\new_[16880]_ ;
  assign \new_[14932]_  = ~\new_[16143]_ ;
  assign \new_[14933]_  = ~\new_[16230]_ ;
  assign \new_[14934]_  = ~\new_[21301]_ ;
  assign \new_[14935]_  = ~\new_[21256]_  & ~\new_[19026]_ ;
  assign \new_[14936]_  = \\text_in_r_reg[12] ;
  assign \new_[14937]_  = \new_[17205]_  | \new_[19758]_ ;
  assign \new_[14938]_  = ~\new_[16641]_ ;
  assign \new_[14939]_  = \new_[16684]_  ^ \new_[1289]_ ;
  assign \new_[14940]_  = ~\new_[16604]_ ;
  assign \new_[14941]_  = \\text_in_r_reg[85] ;
  assign \new_[14942]_  = ~\new_[16267]_ ;
  assign \new_[14943]_  = \\text_in_r_reg[80] ;
  assign \new_[14944]_  = \\text_in_r_reg[66] ;
  assign \new_[14945]_  = ~\new_[17257]_  | ~\new_[18083]_ ;
  assign \new_[14946]_  = \new_[17265]_  | \new_[19553]_ ;
  assign \new_[14947]_  = ~\new_[16639]_ ;
  assign \new_[14948]_  = \\text_in_r_reg[9] ;
  assign \new_[14949]_  = ~\new_[16069]_ ;
  assign \new_[14950]_  = ~\new_[17007]_  & ~\new_[19249]_ ;
  assign \new_[14951]_  = ~\new_[20982]_ ;
  assign \new_[14952]_  = \new_[17248]_  | \new_[21513]_ ;
  assign \new_[14953]_  = ~\new_[16041]_ ;
  assign \new_[14954]_  = ~\new_[17582]_ ;
  assign \new_[14955]_  = ~\new_[17005]_ ;
  assign \new_[14956]_  = \\text_in_r_reg[53] ;
  assign \new_[14957]_  = ~\new_[17282]_  | ~\new_[19097]_ ;
  assign \new_[14958]_  = ~\new_[17024]_  & ~\new_[19117]_ ;
  assign \new_[14959]_  = ~\new_[16757]_  & ~\new_[18615]_ ;
  assign \new_[14960]_  = \\text_in_r_reg[45] ;
  assign \new_[14961]_  = \new_[17097]_  | \new_[18938]_ ;
  assign \new_[14962]_  = \\text_in_r_reg[52] ;
  assign \new_[14963]_  = \new_[18608]_  ^ \new_[17721]_ ;
  assign \new_[14964]_  = ~\new_[16106]_ ;
  assign \new_[14965]_  = \new_[18917]_  ^ \new_[17989]_ ;
  assign \new_[14966]_  = ~\new_[16198]_ ;
  assign \new_[14967]_  = \new_[18658]_  ^ \new_[17823]_ ;
  assign \new_[14968]_  = ~\new_[16238]_ ;
  assign \new_[14969]_  = ~\new_[16220]_ ;
  assign \new_[14970]_  = ~\new_[19267]_  | ~\new_[21686]_ ;
  assign \new_[14971]_  = ~\new_[16698]_  & ~\new_[21686]_ ;
  assign \new_[14972]_  = ~\new_[16973]_  | ~\new_[18113]_ ;
  assign \new_[14973]_  = ~\new_[16845]_  | ~\new_[18035]_ ;
  assign \new_[14974]_  = ~\new_[19053]_  & ~\new_[17036]_ ;
  assign \new_[14975]_  = ~\new_[17081]_  & ~\new_[19357]_ ;
  assign \new_[14976]_  = ~\new_[21566]_  & ~\new_[18646]_ ;
  assign \new_[14977]_  = ~\new_[18271]_  | ~\new_[19168]_  | ~\new_[19750]_  | ~\new_[19047]_ ;
  assign \new_[14978]_  = ~\new_[18861]_  | ~\new_[19219]_  | ~\new_[18480]_  | ~\new_[19484]_ ;
  assign \new_[14979]_  = \new_[16110]_ ;
  assign \new_[14980]_  = \new_[17055]_  & \new_[18607]_ ;
  assign \new_[14981]_  = ~\new_[17088]_  & ~\new_[19741]_ ;
  assign \new_[14982]_  = ~\new_[16720]_  | ~\new_[18035]_ ;
  assign \new_[14983]_  = ~\new_[19801]_  & ~\new_[16972]_ ;
  assign \new_[14984]_  = ~\new_[16556]_ ;
  assign \new_[14985]_  = ~\new_[17336]_  | ~\new_[18627]_ ;
  assign \new_[14986]_  = ~\new_[18391]_  | ~\new_[18464]_  | ~\new_[19033]_  | ~\new_[19676]_ ;
  assign \new_[14987]_  = ~\new_[18959]_  & ~\new_[17072]_ ;
  assign \new_[14988]_  = ~\new_[17175]_  & ~\new_[19253]_ ;
  assign \new_[14989]_  = ~\new_[15922]_ ;
  assign \new_[14990]_  = ~\new_[18103]_  | ~\new_[19409]_  | ~\new_[18733]_  | ~\new_[18867]_ ;
  assign \new_[14991]_  = ~\new_[17972]_  | ~\new_[16965]_ ;
  assign \new_[14992]_  = ~\new_[17171]_  | ~\new_[19568]_ ;
  assign \new_[14993]_  = ~\new_[16465]_ ;
  assign \new_[14994]_  = ~\new_[19118]_  & ~\new_[17445]_ ;
  assign \new_[14995]_  = ~\new_[16116]_ ;
  assign \new_[14996]_  = ~\new_[20664]_  & ~\new_[18852]_ ;
  assign \new_[14997]_  = ~\new_[17277]_  | ~\new_[20927]_ ;
  assign \new_[14998]_  = ~\new_[16144]_ ;
  assign \new_[14999]_  = ~\new_[17200]_  | ~\new_[18607]_ ;
  assign \new_[15000]_  = ~\new_[16828]_  & ~\new_[18978]_ ;
  assign \new_[15001]_  = ~\new_[16398]_ ;
  assign \new_[15002]_  = ~\new_[16398]_ ;
  assign \new_[15003]_  = ~\new_[16118]_ ;
  assign \new_[15004]_  = ~\new_[21571]_  & ~\new_[17185]_ ;
  assign \new_[15005]_  = ~\new_[19553]_  & ~\new_[17175]_ ;
  assign \new_[15006]_  = ~\new_[16756]_  & ~\new_[19000]_ ;
  assign \new_[15007]_  = ~\new_[18450]_  | ~\new_[19454]_ ;
  assign \new_[15008]_  = ~\new_[19301]_  & ~\new_[17102]_ ;
  assign \new_[15009]_  = ~\new_[16373]_ ;
  assign \new_[15010]_  = ~\new_[17096]_  | ~\new_[19288]_ ;
  assign \new_[15011]_  = ~\new_[17582]_ ;
  assign \new_[15012]_  = ~\new_[16739]_  | ~\new_[19156]_ ;
  assign \new_[15013]_  = ~\new_[16361]_ ;
  assign \new_[15014]_  = ~\new_[17433]_  | ~\new_[19024]_ ;
  assign \new_[15015]_  = ~\new_[16791]_  & ~\new_[19100]_ ;
  assign \new_[15016]_  = ~\new_[17093]_  | ~\new_[19084]_ ;
  assign \new_[15017]_  = ~\new_[16871]_  | ~\new_[19098]_ ;
  assign \new_[15018]_  = ~\new_[16911]_  & ~\new_[19335]_ ;
  assign \new_[15019]_  = ~\new_[17353]_  & ~\new_[19066]_ ;
  assign \new_[15020]_  = ~\new_[16883]_  | ~\new_[18166]_ ;
  assign \new_[15021]_  = ~\new_[16786]_  & ~\new_[19719]_ ;
  assign \new_[15022]_  = ~\new_[17268]_  & ~\new_[19426]_ ;
  assign \new_[15023]_  = ~\new_[16770]_  & ~\new_[18821]_ ;
  assign \new_[15024]_  = ~\new_[18375]_  | ~\new_[19746]_ ;
  assign \new_[15025]_  = ~\new_[21411]_  & ~\new_[18974]_ ;
  assign \new_[15026]_  = \new_[18231]_  & \new_[17438]_ ;
  assign \new_[15027]_  = ~\new_[16734]_  & ~\new_[19664]_ ;
  assign \new_[15028]_  = ~\new_[18244]_  | ~\new_[19174]_  | ~\new_[19082]_  | ~\new_[19225]_ ;
  assign \new_[15029]_  = ~\new_[17245]_  | ~\new_[19426]_ ;
  assign \new_[15030]_  = ~\new_[16748]_  & ~\new_[19758]_ ;
  assign \new_[15031]_  = ~\new_[17080]_  & ~\new_[21692]_ ;
  assign \new_[15032]_  = \new_[16870]_  & \new_[19268]_ ;
  assign \new_[15033]_  = ~\new_[17048]_  & ~\new_[18947]_ ;
  assign \new_[15034]_  = ~\new_[17077]_  | ~\new_[19713]_ ;
  assign \new_[15035]_  = ~\new_[16768]_  & ~\new_[19675]_ ;
  assign \new_[15036]_  = ~\new_[17077]_  | ~\new_[18209]_ ;
  assign \new_[15037]_  = ~\new_[16744]_  | ~\new_[18209]_ ;
  assign \new_[15038]_  = ~\new_[16247]_ ;
  assign \new_[15039]_  = \new_[16906]_  & \new_[19098]_ ;
  assign \new_[15040]_  = ~\new_[17227]_  & ~\new_[18968]_ ;
  assign \new_[15041]_  = ~\new_[17247]_  & ~\new_[19617]_ ;
  assign \new_[15042]_  = ~\new_[16753]_  | ~\new_[19713]_ ;
  assign \new_[15043]_  = \new_[17207]_  | \new_[19675]_ ;
  assign \new_[15044]_  = \new_[17655]_  & \new_[19553]_ ;
  assign \new_[15045]_  = ~\new_[17191]_  & ~\new_[19098]_ ;
  assign \new_[15046]_  = ~\new_[16129]_ ;
  assign \new_[15047]_  = \new_[17055]_  & \new_[19553]_ ;
  assign \new_[15048]_  = ~\new_[16216]_ ;
  assign \new_[15049]_  = ~\new_[16132]_ ;
  assign \new_[15050]_  = ~\new_[17169]_  | ~\new_[19385]_ ;
  assign \new_[15051]_  = ~\new_[21500]_  | ~\new_[16984]_ ;
  assign \new_[15052]_  = ~\new_[16133]_ ;
  assign \new_[15053]_  = ~\new_[16137]_ ;
  assign \new_[15054]_  = ~\new_[16780]_  & ~\new_[19750]_ ;
  assign \new_[15055]_  = ~\new_[17173]_  & ~\new_[19176]_ ;
  assign \new_[15056]_  = \new_[16961]_  & \new_[19084]_ ;
  assign \new_[15057]_  = ~\new_[16906]_  | ~\new_[18832]_ ;
  assign \new_[15058]_  = ~\new_[19676]_  & ~\new_[16900]_ ;
  assign \new_[15059]_  = \\text_in_r_reg[97] ;
  assign \new_[15060]_  = ~\new_[17210]_  & ~\new_[18637]_ ;
  assign \new_[15061]_  = ~\new_[17646]_  & ~\new_[19033]_ ;
  assign \new_[15062]_  = \\text_in_r_reg[10] ;
  assign \new_[15063]_  = ~\new_[17194]_  | ~\new_[18209]_ ;
  assign \new_[15064]_  = ~\new_[16863]_  & ~\new_[19374]_ ;
  assign \new_[15065]_  = ~\new_[17235]_  | ~\new_[19217]_ ;
  assign \new_[15066]_  = ~\new_[17193]_  | ~\new_[19319]_ ;
  assign \new_[15067]_  = ~\new_[17280]_  | ~\new_[19589]_ ;
  assign \new_[15068]_  = \\text_in_r_reg[34] ;
  assign \new_[15069]_  = ~\new_[19679]_  & ~\new_[21411]_ ;
  assign \new_[15070]_  = ~\new_[19219]_  & ~\new_[17229]_ ;
  assign \new_[15071]_  = ~\new_[21565]_  | ~\new_[21693]_ ;
  assign \new_[15072]_  = ~\new_[17434]_  & ~\new_[18966]_ ;
  assign \new_[15073]_  = ~\new_[16065]_ ;
  assign \new_[15074]_  = ~\new_[16746]_  & ~\new_[18784]_ ;
  assign \new_[15075]_  = ~\new_[19097]_  & ~\new_[17268]_ ;
  assign \new_[15076]_  = ~\new_[16798]_  | ~\new_[18012]_ ;
  assign \new_[15077]_  = ~\new_[16180]_ ;
  assign \new_[15078]_  = ~\new_[17203]_  & ~\new_[19416]_ ;
  assign \new_[15079]_  = \\text_in_r_reg[110] ;
  assign \new_[15080]_  = \new_[16745]_  | \new_[19156]_ ;
  assign \new_[15081]_  = ~\new_[19681]_  | ~\new_[21563]_  | ~\new_[17611]_ ;
  assign \new_[15082]_  = ~\new_[16857]_  & ~\new_[19459]_ ;
  assign \new_[15083]_  = ~\new_[20747]_  & ~\new_[18974]_ ;
  assign \new_[15084]_  = ~\new_[16067]_ ;
  assign \new_[15085]_  = ~\new_[16151]_ ;
  assign \new_[15086]_  = ~\new_[16056]_ ;
  assign \new_[15087]_  = ~\new_[17306]_  & ~\new_[21575]_ ;
  assign \new_[15088]_  = \new_[17405]_  & \new_[19156]_ ;
  assign \new_[15089]_  = ~\new_[18553]_  | ~\new_[17469]_ ;
  assign \new_[15090]_  = \new_[16838]_  & \new_[17979]_ ;
  assign \new_[15091]_  = ~\new_[21306]_  & ~\new_[16925]_ ;
  assign \new_[15092]_  = ~\new_[16034]_ ;
  assign \new_[15093]_  = ~\new_[16965]_  | ~\new_[19095]_ ;
  assign \new_[15094]_  = ~\new_[15994]_ ;
  assign \new_[15095]_  = \new_[16714]_  | \new_[18906]_ ;
  assign \new_[15096]_  = ~\new_[17690]_  & ~\new_[19319]_ ;
  assign \new_[15097]_  = ~\new_[15982]_ ;
  assign \new_[15098]_  = ~\new_[15966]_ ;
  assign \new_[15099]_  = ~\new_[16780]_  & ~\new_[21638]_ ;
  assign \new_[15100]_  = ~\new_[18945]_  & ~\new_[16699]_ ;
  assign \new_[15101]_  = ~\new_[16144]_ ;
  assign \new_[15102]_  = ~\new_[16906]_  | ~\new_[18965]_ ;
  assign \new_[15103]_  = ~\new_[17214]_  | ~\new_[19742]_ ;
  assign \new_[15104]_  = ~\new_[17096]_  | ~\new_[19589]_ ;
  assign \new_[15105]_  = ~\new_[16919]_  & ~\new_[21498]_ ;
  assign \new_[15106]_  = ~\new_[16158]_ ;
  assign \new_[15107]_  = ~\new_[17210]_  & ~\new_[20490]_ ;
  assign \new_[15108]_  = ~\new_[16884]_  | ~\new_[19689]_ ;
  assign \new_[15109]_  = ~\new_[17009]_  & ~\new_[19100]_ ;
  assign \new_[15110]_  = \new_[16954]_  & \new_[19186]_ ;
  assign \new_[15111]_  = ~\new_[17083]_  & ~\new_[19050]_ ;
  assign \new_[15112]_  = ~\new_[17313]_  | ~\new_[17979]_ ;
  assign \new_[15113]_  = ~\new_[17100]_  | ~\new_[19367]_ ;
  assign \new_[15114]_  = ~\new_[16722]_  & ~\new_[18427]_ ;
  assign \new_[15115]_  = ~\new_[15884]_ ;
  assign \new_[15116]_  = ~\new_[15947]_ ;
  assign \new_[15117]_  = ~\new_[18784]_  & ~\new_[17040]_ ;
  assign \new_[15118]_  = ~\new_[16771]_  | ~\new_[19018]_ ;
  assign \new_[15119]_  = ~\new_[16616]_ ;
  assign \new_[15120]_  = ~\new_[16205]_ ;
  assign \new_[15121]_  = ~\new_[16169]_ ;
  assign \new_[15122]_  = ~\new_[17167]_  | ~\new_[18832]_ ;
  assign \new_[15123]_  = ~\new_[16324]_ ;
  assign \new_[15124]_  = ~\new_[18480]_  | ~\new_[18017]_ ;
  assign \new_[15125]_  = \new_[16913]_  & \new_[19268]_ ;
  assign \new_[15126]_  = ~\new_[16655]_ ;
  assign \new_[15127]_  = ~\new_[17095]_  | ~\new_[19758]_ ;
  assign \new_[15128]_  = ~\new_[17204]_  & ~\new_[21259]_ ;
  assign \new_[15129]_  = ~\new_[16768]_  & ~\new_[19713]_ ;
  assign \new_[15130]_  = ~\new_[18449]_  | ~\new_[15923]_  | ~\new_[19117]_  | ~\new_[19675]_ ;
  assign \new_[15131]_  = ~\new_[17208]_  | ~\new_[19727]_ ;
  assign \new_[15132]_  = ~\new_[16020]_ ;
  assign \new_[15133]_  = ~\new_[16890]_  | ~\new_[19064]_ ;
  assign \new_[15134]_  = ~\new_[18408]_  & ~\new_[16808]_ ;
  assign \new_[15135]_  = ~\new_[16798]_  | ~\new_[21638]_ ;
  assign \new_[15136]_  = ~\new_[17162]_  & ~\new_[21689]_ ;
  assign \new_[15137]_  = ~\new_[16563]_ ;
  assign \new_[15138]_  = ~\new_[16871]_  | ~\new_[19156]_ ;
  assign \new_[15139]_  = ~\new_[16891]_  | ~\new_[20699]_ ;
  assign \new_[15140]_  = ~\new_[16359]_ ;
  assign \new_[15141]_  = ~\new_[16175]_ ;
  assign \new_[15142]_  = ~\new_[16516]_ ;
  assign \new_[15143]_  = ~\new_[16891]_  | ~\new_[21501]_ ;
  assign \new_[15144]_  = ~\new_[17439]_  & ~\new_[17572]_ ;
  assign \new_[15145]_  = ~\new_[16165]_ ;
  assign \new_[15146]_  = ~\new_[18664]_  & ~\new_[16907]_ ;
  assign \new_[15147]_  = \\text_in_r_reg[30] ;
  assign \new_[15148]_  = ~\new_[16455]_ ;
  assign \new_[15149]_  = ~\new_[17230]_  & ~\new_[18194]_ ;
  assign \new_[15150]_  = ~\new_[19535]_  & ~\new_[16804]_ ;
  assign \new_[15151]_  = ~\new_[17352]_  | ~\new_[18607]_ ;
  assign \new_[15152]_  = ~\new_[16458]_ ;
  assign \new_[15153]_  = ~\new_[16209]_ ;
  assign \new_[15154]_  = ~\new_[17031]_  & ~\new_[19426]_ ;
  assign \new_[15155]_  = ~\new_[17211]_  & ~\new_[21689]_ ;
  assign \new_[15156]_  = ~\new_[16234]_ ;
  assign \new_[15157]_  = \new_[17159]_  | \new_[18845]_ ;
  assign \new_[15158]_  = ~\new_[17366]_  & ~\new_[20865]_ ;
  assign \new_[15159]_  = ~\new_[17226]_  & ~\new_[19454]_ ;
  assign \new_[15160]_  = ~\new_[16809]_  & ~\new_[19194]_ ;
  assign \new_[15161]_  = ~\new_[19801]_  & ~\new_[16855]_ ;
  assign \new_[15162]_  = ~\new_[17024]_  & ~\new_[19192]_ ;
  assign \new_[15163]_  = ~\new_[16757]_  & ~\new_[19754]_ ;
  assign \new_[15164]_  = ~\new_[17183]_  & ~\new_[18061]_ ;
  assign \new_[15165]_  = \new_[16683]_  | \new_[18731]_ ;
  assign \new_[15166]_  = ~\new_[16466]_ ;
  assign \new_[15167]_  = ~\new_[17372]_  & ~\new_[18817]_ ;
  assign \new_[15168]_  = ~\new_[17189]_  | ~\new_[19431]_ ;
  assign \new_[15169]_  = \new_[17012]_  | \new_[19156]_ ;
  assign \new_[15170]_  = ~\new_[16303]_ ;
  assign \new_[15171]_  = ~\new_[17283]_  & ~\new_[18637]_ ;
  assign \new_[15172]_  = ~\new_[16805]_  & ~\new_[18682]_ ;
  assign \new_[15173]_  = ~\new_[16999]_  | ~\new_[19104]_ ;
  assign \new_[15174]_  = ~\new_[16835]_  | ~\new_[19727]_ ;
  assign \new_[15175]_  = ~\new_[18144]_  | ~\new_[19425]_ ;
  assign \new_[15176]_  = ~\new_[17239]_  & ~\new_[18979]_ ;
  assign \new_[15177]_  = ~\new_[17845]_  | ~\new_[17092]_ ;
  assign \new_[15178]_  = ~\new_[16195]_ ;
  assign \new_[15179]_  = ~\new_[16196]_ ;
  assign \new_[15180]_  = \new_[16885]_  | \new_[20490]_ ;
  assign \new_[15181]_  = \new_[17179]_  | \new_[18906]_ ;
  assign \new_[15182]_  = \new_[18144]_  & \new_[19636]_ ;
  assign \new_[15183]_  = \new_[17262]_  & \new_[21115]_ ;
  assign \new_[15184]_  = \new_[20925]_  & \new_[19050]_ ;
  assign \new_[15185]_  = ~\new_[17002]_  | ~\new_[19275]_ ;
  assign \new_[15186]_  = ~\new_[17279]_  & ~\new_[19154]_ ;
  assign \new_[15187]_  = ~\new_[17076]_  | ~\new_[17640]_ ;
  assign \new_[15188]_  = \new_[16903]_  | \new_[19268]_ ;
  assign \new_[15189]_  = ~\new_[17206]_  | ~\new_[18077]_ ;
  assign \new_[15190]_  = \new_[17084]_  & \new_[19553]_ ;
  assign \new_[15191]_  = ~\new_[16270]_ ;
  assign \new_[15192]_  = ~\new_[16652]_ ;
  assign \new_[15193]_  = \new_[16869]_  | \new_[18938]_ ;
  assign \new_[15194]_  = ~\new_[21393]_  & ~\new_[18888]_ ;
  assign \new_[15195]_  = ~\new_[20825]_  | ~\new_[16810]_ ;
  assign \new_[15196]_  = \new_[17372]_  | \new_[18616]_ ;
  assign \new_[15197]_  = ~\new_[17141]_  | ~\new_[19785]_ ;
  assign \new_[15198]_  = ~\new_[15946]_ ;
  assign \new_[15199]_  = \new_[17383]_  | \new_[18408]_ ;
  assign \new_[15200]_  = ~\new_[17392]_  | ~\new_[18575]_ ;
  assign \new_[15201]_  = ~\new_[16200]_ ;
  assign \new_[15202]_  = ~\new_[16946]_  & ~\new_[19779]_ ;
  assign \new_[15203]_  = ~\new_[17165]_  & ~\new_[18734]_ ;
  assign \new_[15204]_  = ~\new_[17014]_  | ~\new_[19145]_ ;
  assign \new_[15205]_  = ~\new_[17449]_  & ~\new_[21168]_ ;
  assign \new_[15206]_  = \new_[17047]_  & \new_[19066]_ ;
  assign \new_[15207]_  = ~\new_[21604]_  & ~\new_[19130]_ ;
  assign \new_[15208]_  = ~\new_[17209]_  & ~\new_[18845]_ ;
  assign \new_[15209]_  = ~\new_[16107]_ ;
  assign \new_[15210]_  = \new_[16233]_ ;
  assign \new_[15211]_  = ~\new_[16050]_ ;
  assign \new_[15212]_  = ~\new_[17215]_  | ~\new_[19117]_ ;
  assign \new_[15213]_  = ~\new_[16762]_  & ~\new_[20100]_ ;
  assign \new_[15214]_  = ~\new_[17536]_  | ~\new_[17093]_ ;
  assign \new_[15215]_  = ~\new_[17219]_  & ~\new_[19096]_ ;
  assign \new_[15216]_  = ~\new_[16699]_  & ~\new_[19024]_ ;
  assign \new_[15217]_  = ~\new_[17025]_  & ~\new_[19247]_ ;
  assign \new_[15218]_  = \new_[18557]_  & \new_[16735]_ ;
  assign \new_[15219]_  = \new_[18859]_  | \new_[16776]_ ;
  assign \new_[15220]_  = ~\new_[16894]_  | ~\new_[19196]_ ;
  assign \new_[15221]_  = ~\new_[16355]_ ;
  assign \new_[15222]_  = ~\new_[15921]_ ;
  assign \new_[15223]_  = ~\new_[16218]_ ;
  assign \new_[15224]_  = ~\new_[15914]_ ;
  assign \new_[15225]_  = ~\new_[16219]_ ;
  assign \new_[15226]_  = ~\new_[17176]_  & ~\new_[19084]_ ;
  assign \new_[15227]_  = ~\new_[15900]_ ;
  assign \new_[15228]_  = ~\new_[21500]_  & ~\new_[17212]_ ;
  assign \new_[15229]_  = ~\new_[21393]_  & ~\new_[19664]_ ;
  assign \new_[15230]_  = ~\new_[16821]_  & ~\new_[19145]_ ;
  assign \new_[15231]_  = ~\new_[16912]_  | ~\new_[19425]_ ;
  assign \new_[15232]_  = ~\new_[18465]_  | ~\new_[17213]_ ;
  assign \new_[15233]_  = ~\new_[16144]_ ;
  assign \new_[15234]_  = ~\new_[16154]_ ;
  assign \new_[15235]_  = ~\new_[16144]_ ;
  assign \new_[15236]_  = ~\new_[16675]_ ;
  assign \new_[15237]_  = ~\new_[16718]_  | ~\new_[18678]_ ;
  assign \new_[15238]_  = ~\new_[16221]_ ;
  assign \new_[15239]_  = ~\new_[16221]_ ;
  assign \new_[15240]_  = ~\new_[17279]_  & ~\new_[18637]_ ;
  assign \new_[15241]_  = ~\new_[16728]_  | ~\new_[20239]_ ;
  assign \new_[15242]_  = ~\new_[16802]_  & ~\new_[19538]_ ;
  assign \new_[15243]_  = \new_[17061]_  | \new_[18209]_ ;
  assign \new_[15244]_  = \new_[18206]_  | \new_[17153]_ ;
  assign \new_[15245]_  = ~\new_[16982]_  | ~\new_[18664]_ ;
  assign \new_[15246]_  = ~\new_[17655]_  | ~\new_[19186]_ ;
  assign \new_[15247]_  = ~\new_[17181]_  & ~\new_[19446]_ ;
  assign \new_[15248]_  = ~\new_[17253]_  & ~\new_[19196]_ ;
  assign \new_[15249]_  = ~\new_[16696]_  | ~\new_[18262]_ ;
  assign \new_[15250]_  = \new_[17062]_  | \new_[19156]_ ;
  assign \new_[15251]_  = ~\new_[17226]_  & ~\new_[19548]_ ;
  assign \new_[15252]_  = ~\new_[20237]_  & ~\new_[21605]_ ;
  assign \new_[15253]_  = ~\new_[16225]_ ;
  assign \new_[15254]_  = \new_[16923]_  | \new_[19158]_ ;
  assign \new_[15255]_  = \new_[17223]_  | \new_[19153]_ ;
  assign \new_[15256]_  = ~\new_[17153]_  | ~\new_[19675]_ ;
  assign \new_[15257]_  = ~\new_[17218]_  & ~\new_[19269]_ ;
  assign \new_[15258]_  = ~\new_[16342]_ ;
  assign \new_[15259]_  = \\text_in_r_reg[104] ;
  assign \new_[15260]_  = ~\new_[18931]_  & ~\new_[16911]_ ;
  assign \new_[15261]_  = ~\new_[17456]_  & ~\new_[19637]_ ;
  assign \new_[15262]_  = ~\new_[16269]_ ;
  assign \new_[15263]_  = ~\new_[19076]_  | ~\new_[17093]_ ;
  assign \new_[15264]_  = ~\new_[17983]_  | ~\new_[16728]_ ;
  assign \new_[15265]_  = ~\new_[17164]_  & ~\new_[18659]_ ;
  assign \new_[15266]_  = ~\new_[16227]_ ;
  assign \new_[15267]_  = \new_[17250]_  | \new_[19203]_ ;
  assign \new_[15268]_  = ~\new_[16254]_ ;
  assign \new_[15269]_  = ~\new_[16223]_ ;
  assign \new_[15270]_  = ~\new_[16229]_ ;
  assign \new_[15271]_  = \new_[16928]_  & \new_[19687]_ ;
  assign \new_[15272]_  = \\text_in_r_reg[65] ;
  assign \new_[15273]_  = ~\new_[16231]_ ;
  assign \new_[15274]_  = ~\new_[17271]_  | ~\new_[19217]_ ;
  assign \new_[15275]_  = ~\new_[16858]_  & ~\new_[19729]_ ;
  assign \new_[15276]_  = ~\new_[17178]_  & ~\new_[18840]_ ;
  assign \new_[15277]_  = ~\new_[17350]_  | ~\new_[19476]_ ;
  assign \new_[15278]_  = ~\new_[17186]_  | ~\new_[19275]_ ;
  assign \new_[15279]_  = ~\new_[16188]_ ;
  assign \new_[15280]_  = ~\new_[16235]_ ;
  assign \new_[15281]_  = \new_[17316]_  | \new_[19008]_ ;
  assign \new_[15282]_  = \new_[17456]_  | \new_[18974]_ ;
  assign \new_[15283]_  = ~\new_[17219]_  & ~\new_[19476]_ ;
  assign \new_[15284]_  = ~\new_[16671]_ ;
  assign \new_[15285]_  = ~\new_[16669]_ ;
  assign \new_[15286]_  = ~\new_[17424]_  & ~\new_[19196]_ ;
  assign \new_[15287]_  = ~\new_[17377]_  | ~\new_[19162]_ ;
  assign \new_[15288]_  = ~\new_[16150]_ ;
  assign \new_[15289]_  = \new_[17001]_  | \new_[19462]_ ;
  assign \new_[15290]_  = ~\new_[17092]_  | ~\new_[21686]_ ;
  assign \new_[15291]_  = \new_[16863]_  | \new_[18209]_ ;
  assign \new_[15292]_  = ~\new_[17143]_  & ~\new_[18209]_ ;
  assign \new_[15293]_  = ~\new_[17079]_  & ~\new_[19024]_ ;
  assign \new_[15294]_  = ~\new_[18319]_  | ~\new_[18497]_ ;
  assign \new_[15295]_  = ~\new_[17230]_  & ~\new_[19008]_ ;
  assign \new_[15296]_  = \new_[16849]_  & \new_[14951]_ ;
  assign \new_[15297]_  = ~\new_[17211]_  & ~\new_[19261]_ ;
  assign \new_[15298]_  = ~\new_[16240]_ ;
  assign \new_[15299]_  = \new_[16719]_  | \new_[21635]_ ;
  assign \new_[15300]_  = ~\new_[16189]_ ;
  assign \new_[15301]_  = ~\new_[17061]_  & ~\new_[18187]_ ;
  assign \new_[15302]_  = ~\new_[17018]_  & ~\new_[18810]_ ;
  assign \new_[15303]_  = ~\new_[17174]_  | ~\new_[19409]_ ;
  assign \new_[15304]_  = ~\new_[16987]_  | ~\new_[19269]_ ;
  assign \new_[15305]_  = ~\new_[18250]_  | ~\new_[16954]_ ;
  assign \new_[15306]_  = ~\new_[18728]_  | ~\new_[16718]_ ;
  assign \new_[15307]_  = ~\new_[16245]_ ;
  assign \new_[15308]_  = ~\new_[17142]_  & ~\new_[18979]_ ;
  assign \new_[15309]_  = ~\new_[17758]_  | ~\new_[17414]_ ;
  assign \new_[15310]_  = ~\new_[21565]_  | ~\new_[19048]_ ;
  assign \new_[15311]_  = \new_[16746]_  | \new_[19674]_ ;
  assign \new_[15312]_  = ~\new_[16810]_  | ~\new_[21574]_ ;
  assign \new_[15313]_  = ~\new_[16809]_  & ~\new_[18984]_ ;
  assign \new_[15314]_  = ~\new_[16228]_ ;
  assign \new_[15315]_  = ~\new_[16239]_ ;
  assign \new_[15316]_  = \new_[16783]_  | \new_[18008]_ ;
  assign \new_[15317]_  = ~\new_[17954]_  | ~\new_[16890]_ ;
  assign \new_[15318]_  = ~\new_[16866]_  | ~\new_[19253]_ ;
  assign \new_[15319]_  = ~\new_[16993]_  & ~\new_[19625]_ ;
  assign \new_[15320]_  = ~\new_[18168]_  | ~\new_[18077]_ ;
  assign \new_[15321]_  = ~\new_[17856]_  | ~\new_[16810]_ ;
  assign \new_[15322]_  = ~\new_[16079]_ ;
  assign \new_[15323]_  = ~\new_[16251]_ ;
  assign \new_[15324]_  = \new_[18497]_  & \new_[19153]_ ;
  assign \new_[15325]_  = ~\new_[16778]_  | ~\new_[19253]_ ;
  assign \new_[15326]_  = ~\new_[16785]_  | ~\new_[17657]_ ;
  assign \new_[15327]_  = ~\new_[16750]_  & ~\new_[21496]_ ;
  assign \new_[15328]_  = ~\new_[16252]_ ;
  assign \new_[15329]_  = ~\new_[17350]_  | ~\new_[17144]_ ;
  assign \new_[15330]_  = ~\new_[18707]_  & ~\new_[16768]_ ;
  assign \new_[15331]_  = ~\new_[17242]_  | ~\new_[16863]_ ;
  assign \new_[15332]_  = ~\new_[16125]_ ;
  assign \new_[15333]_  = ~\new_[16004]_ ;
  assign \new_[15334]_  = ~\new_[16548]_ ;
  assign \new_[15335]_  = ~\new_[16810]_  | ~\new_[19367]_ ;
  assign \new_[15336]_  = ~\new_[17322]_  & ~\new_[19376]_ ;
  assign \new_[15337]_  = \new_[17025]_  | \new_[19729]_ ;
  assign \new_[15338]_  = ~\new_[16775]_  & ~\new_[19186]_ ;
  assign \new_[15339]_  = ~\new_[18038]_  | (~\new_[19444]_  & ~\new_[18799]_ );
  assign \new_[15340]_  = ~\new_[18436]_  & ~\new_[16712]_ ;
  assign \new_[15341]_  = ~\new_[21501]_  & ~\new_[17152]_ ;
  assign \new_[15342]_  = ~\new_[16866]_  | ~\new_[18906]_ ;
  assign \new_[15343]_  = ~\new_[16727]_  | ~\new_[21574]_ ;
  assign \new_[15344]_  = ~\new_[21252]_  & ~\new_[21256]_ ;
  assign \new_[15345]_  = ~\new_[16927]_  | (~\new_[20699]_  & ~\new_[21579]_ );
  assign \new_[15346]_  = ~\new_[16783]_  & ~\new_[19266]_ ;
  assign \new_[15347]_  = \new_[17515]_  | \new_[18209]_ ;
  assign \new_[15348]_  = ~\new_[16098]_ ;
  assign \new_[15349]_  = ~\new_[17221]_  & ~\new_[19270]_ ;
  assign \new_[15350]_  = ~\new_[18083]_  & ~\new_[17264]_ ;
  assign \new_[15351]_  = ~\new_[16526]_ ;
  assign \new_[15352]_  = ~\new_[18959]_  & ~\new_[16691]_ ;
  assign \new_[15353]_  = \new_[16874]_  & \new_[19186]_ ;
  assign \new_[15354]_  = ~\new_[17271]_  | ~\new_[19091]_ ;
  assign \new_[15355]_  = ~\new_[16271]_ ;
  assign \new_[15356]_  = ~\new_[17001]_  & ~\new_[21562]_ ;
  assign \new_[15357]_  = ~\new_[16101]_ ;
  assign \new_[15358]_  = \new_[16986]_  | \new_[19102]_ ;
  assign \new_[15359]_  = ~\new_[16735]_  | ~\new_[18008]_ ;
  assign \new_[15360]_  = ~\new_[16082]_ ;
  assign \new_[15361]_  = ~\new_[16963]_  | (~\new_[21574]_  & ~\new_[18009]_ );
  assign \new_[15362]_  = ~\new_[16702]_  | ~\new_[21513]_ ;
  assign \new_[15363]_  = ~\new_[17231]_  & ~\new_[18979]_ ;
  assign \new_[15364]_  = ~\new_[16817]_  & ~\new_[19674]_ ;
  assign \new_[15365]_  = \new_[17180]_  & \new_[17513]_ ;
  assign \new_[15366]_  = ~\new_[16055]_ ;
  assign \new_[15367]_  = ~\new_[17220]_  | ~\new_[19409]_ ;
  assign \new_[15368]_  = ~\new_[17240]_  & ~\new_[19117]_ ;
  assign \new_[15369]_  = \new_[17238]_  | \new_[18948]_ ;
  assign \new_[15370]_  = ~\new_[17154]_  & ~\new_[21306]_ ;
  assign \new_[15371]_  = \new_[17513]_  | \new_[19145]_ ;
  assign \new_[15372]_  = ~\new_[16733]_  & ~\new_[21688]_ ;
  assign \new_[15373]_  = \new_[16888]_  & \new_[19727]_ ;
  assign \new_[15374]_  = ~\new_[16718]_  | ~\new_[18987]_ ;
  assign \new_[15375]_  = \new_[17326]_  | \new_[18832]_ ;
  assign \new_[15376]_  = \new_[16920]_  | \new_[18326]_ ;
  assign \new_[15377]_  = ~\new_[18028]_  | ~\new_[16890]_ ;
  assign \new_[15378]_  = ~\new_[17034]_  & ~\new_[21306]_ ;
  assign \new_[15379]_  = ~\new_[16181]_ ;
  assign \new_[15380]_  = ~\new_[17308]_  & ~\new_[20490]_ ;
  assign \new_[15381]_  = ~\new_[17233]_  & (~\new_[17578]_  | ~\new_[18378]_ );
  assign \new_[15382]_  = ~\new_[16185]_ ;
  assign \new_[15383]_  = ~\new_[16284]_ ;
  assign \new_[15384]_  = ~\new_[16211]_ ;
  assign \new_[15385]_  = ~\new_[16179]_ ;
  assign \new_[15386]_  = ~\new_[17403]_  | ~\new_[19144]_ ;
  assign \new_[15387]_  = ~\new_[16864]_  | ~\new_[17457]_ ;
  assign \new_[15388]_  = ~\new_[16176]_ ;
  assign \new_[15389]_  = ~\new_[16280]_ ;
  assign \new_[15390]_  = ~\new_[16163]_ ;
  assign \new_[15391]_  = ~\new_[16146]_ ;
  assign \new_[15392]_  = ~\new_[16236]_ ;
  assign \new_[15393]_  = ~\new_[16113]_ ;
  assign \new_[15394]_  = ~\new_[17403]_  | ~\new_[19275]_ ;
  assign \new_[15395]_  = ~\new_[16287]_ ;
  assign \new_[15396]_  = ~\new_[16289]_ ;
  assign \new_[15397]_  = ~\new_[16898]_  | ~\new_[18947]_ ;
  assign \new_[15398]_  = ~\new_[16096]_ ;
  assign \new_[15399]_  = ~\new_[16293]_ ;
  assign \new_[15400]_  = ~\new_[16294]_ ;
  assign \new_[15401]_  = ~\new_[16800]_  | ~\new_[19249]_ ;
  assign \new_[15402]_  = ~\new_[16298]_ ;
  assign \new_[15403]_  = ~\new_[16299]_ ;
  assign \new_[15404]_  = ~\new_[16729]_  | ~\new_[21306]_ ;
  assign \new_[15405]_  = ~\new_[16075]_ ;
  assign \new_[15406]_  = ~\new_[16302]_ ;
  assign \new_[15407]_  = ~\new_[17415]_  | ~\new_[19353]_ ;
  assign \new_[15408]_  = ~\new_[16071]_ ;
  assign \new_[15409]_  = ~\new_[16305]_ ;
  assign \new_[15410]_  = ~\new_[16306]_ ;
  assign \new_[15411]_  = ~\new_[17094]_  | ~\new_[19719]_ ;
  assign \new_[15412]_  = ~\new_[16183]_ ;
  assign \new_[15413]_  = ~\new_[16059]_ ;
  assign \new_[15414]_  = \new_[21528]_  | \new_[18017]_ ;
  assign \new_[15415]_  = ~\new_[19444]_  & ~\new_[17182]_ ;
  assign \new_[15416]_  = ~\new_[16749]_  | ~\new_[18542]_ ;
  assign \new_[15417]_  = ~\new_[16064]_ ;
  assign \new_[15418]_  = ~\new_[16311]_ ;
  assign \new_[15419]_  = ~\new_[16665]_ ;
  assign \new_[15420]_  = ~\new_[16314]_ ;
  assign \new_[15421]_  = ~\new_[16076]_ ;
  assign \new_[15422]_  = ~\new_[16038]_ ;
  assign \new_[15423]_  = ~\new_[16317]_ ;
  assign \new_[15424]_  = ~\new_[16827]_  | ~\new_[17363]_ ;
  assign \new_[15425]_  = ~\new_[16193]_ ;
  assign \new_[15426]_  = ~\new_[17079]_  & ~\new_[19212]_ ;
  assign \new_[15427]_  = ~\new_[16016]_ ;
  assign \new_[15428]_  = ~\new_[16983]_  | ~\new_[21584]_ ;
  assign \new_[15429]_  = ~\new_[16709]_  | ~\new_[19342]_ ;
  assign \new_[15430]_  = \new_[16005]_ ;
  assign \new_[15431]_  = ~\new_[17399]_  | ~\new_[18810]_ ;
  assign \new_[15432]_  = \new_[17406]_  | \new_[19082]_ ;
  assign \new_[15433]_  = ~\new_[15988]_ ;
  assign \new_[15434]_  = ~\new_[18672]_  & ~\new_[18209]_ ;
  assign \new_[15435]_  = ~\new_[15960]_ ;
  assign \new_[15436]_  = \new_[16693]_  | \new_[21507]_ ;
  assign \new_[15437]_  = ~\new_[16168]_ ;
  assign \new_[15438]_  = ~\new_[15964]_ ;
  assign \new_[15439]_  = \new_[16782]_  & \new_[17671]_ ;
  assign \new_[15440]_  = \new_[17393]_  | \new_[19431]_ ;
  assign \new_[15441]_  = ~\new_[16325]_ ;
  assign \new_[15442]_  = ~\new_[21255]_ ;
  assign \new_[15443]_  = ~\new_[16327]_ ;
  assign \new_[15444]_  = ~\new_[17396]_  & ~\new_[21693]_ ;
  assign \new_[15445]_  = ~\new_[15941]_ ;
  assign \new_[15446]_  = ~\new_[16350]_ ;
  assign \new_[15447]_  = ~\new_[15913]_ ;
  assign \new_[15448]_  = ~\new_[16331]_ ;
  assign \new_[15449]_  = ~\new_[16524]_ ;
  assign \new_[15450]_  = ~\new_[16154]_ ;
  assign \new_[15451]_  = ~\new_[16413]_ ;
  assign \new_[15452]_  = ~\new_[15908]_ ;
  assign \new_[15453]_  = ~\new_[16335]_ ;
  assign \new_[15454]_  = \new_[19824]_  | \new_[20865]_ ;
  assign \new_[15455]_  = ~\new_[20665]_  | ~\new_[21688]_ ;
  assign \new_[15456]_  = ~\new_[18518]_  & ~\new_[19275]_ ;
  assign \new_[15457]_  = ~\new_[16336]_ ;
  assign \new_[15458]_  = ~\new_[16154]_ ;
  assign \new_[15459]_  = ~\new_[16134]_ ;
  assign \new_[15460]_  = ~\new_[18204]_  | ~\new_[19013]_ ;
  assign \new_[15461]_  = \new_[16645]_ ;
  assign \new_[15462]_  = ~\new_[18108]_  | ~\new_[18621]_ ;
  assign \new_[15463]_  = ~\new_[16591]_ ;
  assign \new_[15464]_  = ~\new_[16580]_ ;
  assign \new_[15465]_  = ~\new_[16970]_  & ~\new_[21688]_ ;
  assign \new_[15466]_  = ~\new_[16343]_ ;
  assign \new_[15467]_  = ~\new_[16529]_ ;
  assign \new_[15468]_  = ~\new_[17574]_  | ~\new_[18104]_ ;
  assign \new_[15469]_  = ~\new_[17044]_  & ~\new_[19097]_ ;
  assign \new_[15470]_  = \\text_in_r_reg[79] ;
  assign \new_[15471]_  = ~\new_[16344]_ ;
  assign \new_[15472]_  = ~\new_[16345]_ ;
  assign \new_[15473]_  = ~\new_[16347]_ ;
  assign \new_[15474]_  = \new_[17085]_  | \new_[18575]_ ;
  assign \new_[15475]_  = ~\new_[16350]_ ;
  assign \new_[15476]_  = ~\new_[16353]_ ;
  assign \new_[15477]_  = \new_[17096]_  & \new_[19655]_ ;
  assign \new_[15478]_  = ~\new_[16579]_ ;
  assign \new_[15479]_  = ~\new_[17165]_  & ~\new_[21499]_ ;
  assign \new_[15480]_  = ~\new_[17705]_  | ~\new_[18973]_ ;
  assign \new_[15481]_  = ~\new_[16977]_  | ~\new_[20495]_ ;
  assign \new_[15482]_  = \\text_in_r_reg[7] ;
  assign \new_[15483]_  = ~\new_[16992]_  | ~\new_[18454]_ ;
  assign \new_[15484]_  = ~\new_[16138]_ ;
  assign \new_[15485]_  = ~\new_[16890]_  | ~\new_[20865]_ ;
  assign \new_[15486]_  = ~\new_[16127]_ ;
  assign \new_[15487]_  = ~\new_[17191]_ ;
  assign \new_[15488]_  = ~\new_[15935]_ ;
  assign \new_[15489]_  = ~\new_[17426]_  | ~\new_[19719]_ ;
  assign \new_[15490]_  = ~\new_[20235]_  | ~\new_[20865]_ ;
  assign \new_[15491]_  = ~\new_[16084]_ ;
  assign \new_[15492]_  = ~\new_[17378]_  | ~\new_[19676]_ ;
  assign \new_[15493]_  = ~\new_[16076]_ ;
  assign \new_[15494]_  = ~\new_[16263]_ ;
  assign \new_[15495]_  = ~\new_[16070]_ ;
  assign \new_[15496]_  = ~\new_[17971]_  | ~\new_[17304]_ ;
  assign \new_[15497]_  = ~\new_[18250]_  | ~\new_[16846]_ ;
  assign \new_[15498]_  = ~\new_[18144]_  | ~\new_[19335]_ ;
  assign \new_[15499]_  = ~\new_[15903]_ ;
  assign \new_[15500]_  = ~\new_[17380]_  | ~\new_[19436]_ ;
  assign \new_[15501]_  = ~\new_[16368]_ ;
  assign \new_[15502]_  = ~\new_[17410]_  & ~\new_[18888]_ ;
  assign \new_[15503]_  = ~\new_[16846]_  | ~\new_[19066]_ ;
  assign \new_[15504]_  = ~\new_[18492]_  | ~\new_[18621]_ ;
  assign \new_[15505]_  = ~\new_[16115]_ ;
  assign \new_[15506]_  = ~\new_[16030]_ ;
  assign \new_[15507]_  = ~\new_[16910]_  & ~\new_[19428]_ ;
  assign \new_[15508]_  = ~\new_[16716]_  | ~\new_[19538]_ ;
  assign \new_[15509]_  = ~\new_[16097]_ ;
  assign \new_[15510]_  = ~\new_[16264]_ ;
  assign \new_[15511]_  = ~\new_[18243]_  | ~\new_[19386]_ ;
  assign \new_[15512]_  = ~\new_[17295]_  & ~\new_[18974]_ ;
  assign \new_[15513]_  = ~\new_[16999]_  | ~\new_[19754]_ ;
  assign \new_[15514]_  = ~\new_[16626]_ ;
  assign \new_[15515]_  = ~\new_[16668]_ ;
  assign \new_[15516]_  = ~\new_[15992]_ ;
  assign \new_[15517]_  = ~\new_[15985]_ ;
  assign \new_[15518]_  = ~\new_[16981]_  & ~\new_[19082]_ ;
  assign \new_[15519]_  = ~\new_[15967]_ ;
  assign \new_[15520]_  = \new_[21712]_  | \new_[19085]_ ;
  assign \new_[15521]_  = ~\new_[15948]_ ;
  assign \new_[15522]_  = ~\new_[16817]_  & ~\new_[18235]_ ;
  assign \new_[15523]_  = ~\new_[16742]_ ;
  assign \new_[15524]_  = \new_[18479]_  | \new_[17979]_ ;
  assign \new_[15525]_  = ~\new_[15928]_ ;
  assign \new_[15526]_  = ~\new_[15933]_ ;
  assign \new_[15527]_  = ~\new_[15924]_ ;
  assign \new_[15528]_  = \new_[16764]_  & \new_[19413]_ ;
  assign \new_[15529]_  = ~\new_[16275]_ ;
  assign \new_[15530]_  = ~\new_[16394]_ ;
  assign \new_[15531]_  = ~\new_[18275]_  | ~\new_[18107]_ ;
  assign \new_[15532]_  = ~\new_[17243]_  & ~\new_[19459]_ ;
  assign \new_[15533]_  = ~\new_[15898]_ ;
  assign \new_[15534]_  = ~\new_[20930]_  | ~\new_[19476]_ ;
  assign \new_[15535]_  = ~\new_[17312]_  | ~\new_[19266]_ ;
  assign \new_[15536]_  = ~\new_[15878]_ ;
  assign \new_[15537]_  = ~\new_[16391]_ ;
  assign \new_[15538]_  = ~\new_[16882]_  | ~\new_[18166]_ ;
  assign \new_[15539]_  = ~\new_[16672]_ ;
  assign \new_[15540]_  = ~\new_[16396]_ ;
  assign \new_[15541]_  = ~\new_[17710]_  | ~\new_[18425]_ ;
  assign \new_[15542]_  = ~\new_[16792]_  | ~\new_[21515]_ ;
  assign \new_[15543]_  = ~\new_[21045]_ ;
  assign \new_[15544]_  = \new_[16687]_  | \new_[18938]_ ;
  assign \new_[15545]_  = ~\new_[16662]_ ;
  assign \new_[15546]_  = ~\new_[16654]_ ;
  assign \new_[15547]_  = ~\new_[19553]_  | ~\new_[17505]_ ;
  assign \new_[15548]_  = ~\new_[17420]_  & ~\new_[19801]_ ;
  assign \new_[15549]_  = ~\new_[16094]_ ;
  assign \new_[15550]_  = ~\new_[16349]_ ;
  assign \new_[15551]_  = \new_[17105]_  | \new_[17469]_ ;
  assign \new_[15552]_  = ~\new_[16403]_ ;
  assign \new_[15553]_  = ~\new_[16589]_ ;
  assign \new_[15554]_  = ~\new_[16160]_ ;
  assign \new_[15555]_  = ~\new_[17240]_  & ~\new_[19192]_ ;
  assign \new_[15556]_  = ~\new_[16560]_ ;
  assign \new_[15557]_  = \new_[17109]_  & \new_[19553]_ ;
  assign \new_[15558]_  = ~\new_[15910]_ ;
  assign \new_[15559]_  = ~\new_[18432]_  & ~\new_[19555]_ ;
  assign \new_[15560]_  = ~\new_[16451]_ ;
  assign \new_[15561]_  = ~\new_[16372]_ ;
  assign \new_[15562]_  = \new_[18142]_  & \new_[21689]_ ;
  assign \new_[15563]_  = ~\new_[17356]_  | ~\new_[18794]_ ;
  assign \new_[15564]_  = ~\new_[16954]_  | ~\new_[19555]_ ;
  assign \new_[15565]_  = ~\new_[16315]_ ;
  assign \new_[15566]_  = \new_[16249]_ ;
  assign \new_[15567]_  = ~\new_[16814]_  & ~\new_[20869]_ ;
  assign \new_[15568]_  = ~\new_[16354]_ ;
  assign \new_[15569]_  = ~\new_[16737]_  & ~\new_[19118]_ ;
  assign \new_[15570]_  = ~\new_[18338]_  | ~\new_[19261]_ ;
  assign \new_[15571]_  = ~\new_[17300]_  | ~\new_[18692]_ ;
  assign \new_[15572]_  = ~\new_[17354]_  & ~\new_[18810]_ ;
  assign \new_[15573]_  = ~\new_[16897]_  | ~\new_[19624]_ ;
  assign \new_[15574]_  = ~\new_[16887]_  | ~\new_[19655]_ ;
  assign \new_[15575]_  = ~\new_[16108]_ ;
  assign \new_[15576]_  = ~\new_[16872]_  | ~\new_[19535]_ ;
  assign \new_[15577]_  = ~\new_[17676]_  | ~\new_[17147]_ ;
  assign \new_[15578]_  = ~\new_[16796]_  & ~\new_[19084]_ ;
  assign \new_[15579]_  = ~\new_[16523]_ ;
  assign \new_[15580]_  = ~\new_[17278]_  | ~\new_[19674]_ ;
  assign \new_[15581]_  = ~\new_[16261]_ ;
  assign \new_[15582]_  = ~\new_[16273]_ ;
  assign \new_[15583]_  = ~\new_[17931]_  & ~\new_[18414]_ ;
  assign \new_[15584]_  = ~\new_[16428]_ ;
  assign \new_[15585]_  = \new_[17437]_  | \new_[19727]_ ;
  assign \new_[15586]_  = ~\new_[16003]_ ;
  assign \new_[15587]_  = ~\new_[15998]_ ;
  assign \new_[15588]_  = ~\new_[16001]_ ;
  assign \new_[15589]_  = ~\new_[17436]_  & ~\new_[19476]_ ;
  assign \new_[15590]_  = ~\new_[15990]_ ;
  assign \new_[15591]_  = ~\new_[15987]_ ;
  assign \new_[15592]_  = ~\new_[15974]_ ;
  assign \new_[15593]_  = ~\new_[18323]_  | ~\new_[18455]_ ;
  assign \new_[15594]_  = ~\new_[15957]_ ;
  assign \new_[15595]_  = ~\new_[16431]_ ;
  assign \new_[15596]_  = ~\new_[17607]_  & ~\new_[19150]_  & ~\new_[19428]_ ;
  assign \new_[15597]_  = \new_[16927]_  | \new_[21513]_ ;
  assign \new_[15598]_  = ~\new_[17365]_  | ~\new_[19044]_ ;
  assign \new_[15599]_  = ~\new_[17033]_  | ~\new_[18811]_ ;
  assign \new_[15600]_  = ~\new_[17029]_  | ~\new_[19061]_ ;
  assign \new_[15601]_  = ~\new_[17454]_  | ~\new_[19367]_ ;
  assign \new_[15602]_  = ~\new_[21513]_  & ~\new_[21142]_ ;
  assign \new_[15603]_  = ~\new_[17260]_  | ~\new_[19679]_ ;
  assign \new_[15604]_  = \new_[17612]_  | \new_[19098]_ ;
  assign \new_[15605]_  = ~\new_[15886]_ ;
  assign \new_[15606]_  = ~\new_[15872]_ ;
  assign \new_[15607]_  = ~\new_[18465]_  | ~\new_[17296]_ ;
  assign \new_[15608]_  = ~\new_[16044]_ ;
  assign \new_[15609]_  = ~\new_[17361]_  | ~\new_[21569]_ ;
  assign \new_[15610]_  = ~\new_[18107]_  | ~\new_[21562]_ ;
  assign \new_[15611]_  = \new_[19655]_  & \new_[18161]_ ;
  assign \new_[15612]_  = ~\new_[17451]_  | ~\new_[17505]_ ;
  assign \new_[15613]_  = ~\new_[17933]_  & ~\new_[21513]_ ;
  assign \new_[15614]_  = ~\new_[16633]_ ;
  assign \new_[15615]_  = ~\new_[17336]_  | ~\new_[21513]_ ;
  assign \new_[15616]_  = ~\new_[16586]_ ;
  assign \new_[15617]_  = ~\new_[16587]_ ;
  assign \new_[15618]_  = ~\new_[16566]_ ;
  assign \new_[15619]_  = ~\new_[16358]_ ;
  assign \new_[15620]_  = ~\new_[16562]_ ;
  assign \new_[15621]_  = \new_[17416]_  | \new_[19036]_ ;
  assign \new_[15622]_  = ~\new_[16454]_ ;
  assign \new_[15623]_  = ~\new_[17981]_  | ~\new_[18605]_ ;
  assign \new_[15624]_  = ~\new_[17300]_  | ~\new_[19247]_ ;
  assign \new_[15625]_  = ~\new_[16404]_ ;
  assign \new_[15626]_  = ~\new_[16024]_ ;
  assign \new_[15627]_  = ~\new_[16187]_ ;
  assign \new_[15628]_  = ~\new_[19285]_  & ~\new_[21302]_ ;
  assign \new_[15629]_  = \new_[16265]_ ;
  assign \new_[15630]_  = ~\new_[16014]_ ;
  assign \new_[15631]_  = ~\new_[16983]_  | ~\new_[21513]_ ;
  assign \new_[15632]_  = ~\new_[17235]_ ;
  assign \new_[15633]_  = ~\new_[17455]_  | ~\new_[19208]_ ;
  assign \new_[15634]_  = \\text_in_r_reg[82] ;
  assign \new_[15635]_  = ~\new_[16647]_ ;
  assign \new_[15636]_  = ~\new_[16577]_ ;
  assign \new_[15637]_  = ~\new_[16085]_ ;
  assign \new_[15638]_  = ~\new_[16471]_ ;
  assign \new_[15639]_  = ~\new_[17418]_  & ~\new_[19150]_ ;
  assign \new_[15640]_  = ~\new_[18898]_  | ~\new_[17368]_ ;
  assign \new_[15641]_  = \new_[18450]_  & \new_[18984]_ ;
  assign \new_[15642]_  = ~\new_[15870]_ ;
  assign \new_[15643]_  = ~\new_[16224]_ ;
  assign \new_[15644]_  = ~\new_[16477]_ ;
  assign \new_[15645]_  = ~\new_[16100]_ ;
  assign \new_[15646]_  = ~\new_[19156]_  | ~\new_[19419]_  | ~\new_[18772]_ ;
  assign \new_[15647]_  = ~\new_[15911]_ ;
  assign \new_[15648]_  = ~\new_[15972]_ ;
  assign \new_[15649]_  = ~\new_[15895]_ ;
  assign \new_[15650]_  = ~\new_[16797]_  | ~\new_[17614]_ ;
  assign \new_[15651]_  = ~\new_[15891]_ ;
  assign \new_[15652]_  = ~\new_[15879]_ ;
  assign \new_[15653]_  = ~\new_[15883]_ ;
  assign \new_[15654]_  = ~\new_[18194]_  & ~\new_[19114]_ ;
  assign \new_[15655]_  = ~\new_[16843]_  & ~\new_[19197]_ ;
  assign \new_[15656]_  = ~\new_[17454]_  | ~\new_[21569]_ ;
  assign \new_[15657]_  = ~\new_[17244]_ ;
  assign \new_[15658]_  = ~\new_[16882]_  & ~\new_[19474]_ ;
  assign \new_[15659]_  = ~\new_[16590]_ ;
  assign \new_[15660]_  = ~\new_[18079]_  | ~\new_[18140]_ ;
  assign \new_[15661]_  = ~\new_[17296]_  | ~\new_[19655]_ ;
  assign \new_[15662]_  = ~\new_[16573]_ ;
  assign \new_[15663]_  = ~\new_[16569]_ ;
  assign \new_[15664]_  = ~\new_[16411]_ ;
  assign \new_[15665]_  = ~\new_[16881]_  & ~\new_[18228]_ ;
  assign \new_[15666]_  = ~\new_[17333]_  & ~\new_[19104]_ ;
  assign \new_[15667]_  = ~\new_[16497]_ ;
  assign \new_[15668]_  = ~\new_[19290]_  | ~\new_[18050]_  | ~\new_[17578]_ ;
  assign \new_[15669]_  = ~\new_[16865]_  & ~\new_[18640]_ ;
  assign \new_[15670]_  = ~\new_[17564]_  | ~\new_[18325]_ ;
  assign \new_[15671]_  = ~\new_[17574]_  | ~\new_[19256]_ ;
  assign \new_[15672]_  = ~\new_[16689]_  | ~\new_[18577]_ ;
  assign \new_[15673]_  = \new_[18314]_  & \new_[18637]_ ;
  assign \new_[15674]_  = ~\new_[16473]_ ;
  assign \new_[15675]_  = ~\new_[16506]_ ;
  assign \new_[15676]_  = ~\new_[16574]_ ;
  assign \new_[15677]_  = ~\new_[16152]_ ;
  assign \new_[15678]_  = ~\new_[16508]_ ;
  assign \new_[15679]_  = ~\new_[15896]_ ;
  assign \new_[15680]_  = ~\new_[18788]_  | ~\new_[16708]_ ;
  assign \new_[15681]_  = \new_[18256]_  & \new_[19068]_ ;
  assign \new_[15682]_  = ~\new_[16052]_ ;
  assign \new_[15683]_  = ~\new_[16147]_ ;
  assign \new_[15684]_  = ~\new_[17058]_  & ~\new_[19224]_ ;
  assign \new_[15685]_  = ~\new_[16456]_ ;
  assign \new_[15686]_  = ~\new_[19203]_  | ~\new_[19166]_  | ~\new_[18378]_ ;
  assign \new_[15687]_  = ~\new_[21113]_ ;
  assign \new_[15688]_  = ~\new_[18938]_  | ~\new_[19373]_  | ~\new_[17482]_ ;
  assign \new_[15689]_  = ~\new_[15880]_ ;
  assign \new_[15690]_  = \new_[16652]_ ;
  assign \new_[15691]_  = ~\new_[17698]_  | ~\new_[16879]_ ;
  assign \new_[15692]_  = \new_[17360]_  | \new_[19044]_ ;
  assign \new_[15693]_  = ~\new_[17093]_  | ~\new_[19091]_ ;
  assign \new_[15694]_  = ~\new_[16203]_ ;
  assign \new_[15695]_  = ~\new_[20825]_  | ~\new_[16976]_ ;
  assign \new_[15696]_  = ~\new_[16567]_ ;
  assign \new_[15697]_  = ~\new_[17393]_  | ~\new_[17401]_ ;
  assign \new_[15698]_  = ~\new_[16551]_ ;
  assign \new_[15699]_  = ~\new_[16584]_ ;
  assign \new_[15700]_  = ~\new_[18869]_  | ~\new_[17304]_ ;
  assign \new_[15701]_  = ~\new_[18484]_  | ~\new_[18735]_ ;
  assign \new_[15702]_  = ~\new_[16414]_ ;
  assign \new_[15703]_  = \\text_in_r_reg[126] ;
  assign \new_[15704]_  = ~\new_[16301]_ ;
  assign \new_[15705]_  = ~\new_[17345]_  | ~\new_[21115]_ ;
  assign \new_[15706]_  = ~\new_[17431]_  & ~\new_[19409]_ ;
  assign \new_[15707]_  = ~\new_[17386]_  & ~\new_[18421]_ ;
  assign \new_[15708]_  = ~\new_[18732]_  | ~\new_[14951]_ ;
  assign \new_[15709]_  = ~\new_[18867]_  | ~\new_[17454]_ ;
  assign \new_[15710]_  = ~\new_[15995]_ ;
  assign \new_[15711]_  = ~\new_[16058]_ ;
  assign \new_[15712]_  = ~\new_[21631]_  | ~\new_[17304]_ ;
  assign \new_[15713]_  = ~\new_[16833]_  | ~\new_[19019]_ ;
  assign \new_[15714]_  = ~\new_[16533]_ ;
  assign \new_[15715]_  = ~\new_[16313]_ ;
  assign \new_[15716]_  = ~\new_[17145]_  | ~\new_[18974]_ ;
  assign \new_[15717]_  = \new_[18038]_  | \new_[19084]_ ;
  assign \new_[15718]_  = \new_[16755]_  | \new_[20699]_ ;
  assign \new_[15719]_  = ~\new_[17375]_  | ~\new_[17578]_ ;
  assign \new_[15720]_  = \new_[15871]_ ;
  assign \new_[15721]_  = ~\new_[18134]_  | ~\new_[19117]_ ;
  assign \new_[15722]_  = ~\new_[16901]_  | ~\new_[18640]_ ;
  assign \new_[15723]_  = \new_[16988]_  | \new_[18709]_ ;
  assign \new_[15724]_  = ~\new_[16539]_ ;
  assign \new_[15725]_  = ~\new_[18369]_  | ~\new_[17054]_ ;
  assign \new_[15726]_  = ~\new_[16603]_ ;
  assign \new_[15727]_  = ~\new_[17033]_  & ~\new_[17677]_ ;
  assign \new_[15728]_  = ~\new_[20661]_  | ~\new_[17332]_ ;
  assign \new_[15729]_  = \new_[17427]_  | \new_[17344]_ ;
  assign \new_[15730]_  = ~\new_[18319]_  | ~\new_[17597]_ ;
  assign \new_[15731]_  = ~\new_[17504]_  | ~\new_[17338]_ ;
  assign \new_[15732]_  = \new_[18465]_  & \new_[18455]_ ;
  assign \new_[15733]_  = ~\new_[17431]_  | ~\new_[19151]_ ;
  assign \new_[15734]_  = \new_[17367]_  & \new_[18173]_ ;
  assign \new_[15735]_  = ~\new_[20662]_  & ~\new_[16759]_ ;
  assign \new_[15736]_  = ~\new_[17395]_  | ~\new_[17260]_ ;
  assign \new_[15737]_  = ~\new_[18349]_  | ~\new_[18812]_ ;
  assign \new_[15738]_  = \new_[17423]_  | \new_[17592]_ ;
  assign \new_[15739]_  = ~\new_[16832]_  | ~\new_[17369]_ ;
  assign \new_[15740]_  = ~\new_[17793]_  & ~\new_[17368]_ ;
  assign \new_[15741]_  = ~\new_[16534]_ ;
  assign \new_[15742]_  = ~\new_[17942]_  | ~\new_[17388]_ ;
  assign \new_[15743]_  = ~\new_[16546]_ ;
  assign \new_[15744]_  = ~\new_[16334]_ ;
  assign \new_[15745]_  = ~\new_[17043]_  | ~\new_[17065]_ ;
  assign \new_[15746]_  = ~\new_[17554]_  & ~\new_[18509]_ ;
  assign \new_[15747]_  = ~\new_[17395]_  | ~\new_[16934]_ ;
  assign \new_[15748]_  = ~\new_[17370]_  & ~\new_[21711]_ ;
  assign \new_[15749]_  = ~\new_[18299]_  | (~\new_[19526]_  & ~\new_[18906]_ );
  assign \new_[15750]_  = ~\new_[17436]_  | (~\new_[18096]_  & ~\new_[19096]_ );
  assign \new_[15751]_  = ~\new_[18788]_  | ~\new_[16905]_ ;
  assign \new_[15752]_  = ~\new_[16145]_ ;
  assign \new_[15753]_  = ~\new_[16551]_ ;
  assign \new_[15754]_  = ~\new_[16490]_ ;
  assign \new_[15755]_  = \new_[17292]_  & \new_[17597]_ ;
  assign \new_[15756]_  = \\text_in_r_reg[105] ;
  assign \new_[15757]_  = \\text_in_r_reg[13] ;
  assign \new_[15758]_  = ~\new_[16933]_  | ~\new_[19353]_ ;
  assign \new_[15759]_  = ~\new_[18432]_  | ~\new_[17867]_ ;
  assign \new_[15760]_  = \new_[17667]_  & \new_[16908]_ ;
  assign \new_[15761]_  = ~\new_[19182]_  & ~\new_[17152]_ ;
  assign \new_[15762]_  = \new_[18301]_  & \new_[19665]_ ;
  assign \new_[15763]_  = \new_[14951]_  & \new_[19277]_ ;
  assign \new_[15764]_  = ~\new_[17359]_  | ~\new_[17389]_ ;
  assign \new_[15765]_  = ~\new_[16452]_ ;
  assign \new_[15766]_  = \new_[19799]_  ^ \new_[19123]_ ;
  assign \new_[15767]_  = ~\new_[19469]_ ;
  assign \new_[15768]_  = \new_[19115]_  & \new_[18179]_ ;
  assign \new_[15769]_  = \new_[14772]_  ^ \new_[1675]_ ;
  assign \new_[15770]_  = ~\new_[17269]_  & ~\new_[21166]_ ;
  assign \new_[15771]_  = \new_[14762]_  ^ \new_[18829]_ ;
  assign \new_[15772]_  = ~\new_[16837]_  & ~\new_[20927]_ ;
  assign \new_[15773]_  = ~\new_[16576]_ ;
  assign \new_[15774]_  = \new_[19570]_  ^ \new_[18741]_ ;
  assign \new_[15775]_  = ~\new_[16583]_ ;
  assign \new_[15776]_  = ~\new_[16588]_ ;
  assign \new_[15777]_  = ~\new_[16742]_ ;
  assign \new_[15778]_  = ~\new_[16742]_ ;
  assign \new_[15779]_  = ~\new_[16154]_ ;
  assign \new_[15780]_  = ~\new_[16221]_ ;
  assign \new_[15781]_  = ~\new_[15922]_ ;
  assign \new_[15782]_  = ~\new_[15922]_ ;
  assign \new_[15783]_  = ~\new_[16103]_ ;
  assign \new_[15784]_  = ~\new_[18392]_  | ~\new_[17387]_ ;
  assign \new_[15785]_  = ~\new_[17525]_  | ~\new_[16942]_ ;
  assign \new_[15786]_  = ~\new_[18585]_  | ~\new_[18176]_ ;
  assign \new_[15787]_  = ~\new_[16203]_ ;
  assign \new_[15788]_  = ~\new_[16112]_ ;
  assign \new_[15789]_  = ~\new_[17254]_  & ~\new_[18427]_ ;
  assign \new_[15790]_  = ~\new_[16111]_ ;
  assign \new_[15791]_  = ~\new_[16690]_  | ~\new_[19428]_ ;
  assign \new_[15792]_  = ~\new_[19064]_  & ~\new_[18199]_ ;
  assign \new_[15793]_  = \new_[19098]_  & \new_[17553]_ ;
  assign \new_[15794]_  = ~\new_[16092]_ ;
  assign \new_[15795]_  = ~\new_[16012]_ ;
  assign \new_[15796]_  = ~\new_[16740]_  | ~\new_[19548]_ ;
  assign \new_[15797]_  = ~\new_[16915]_  & ~\new_[19434]_ ;
  assign \new_[15798]_  = \new_[19308]_  & \new_[19717]_ ;
  assign \new_[15799]_  = \new_[17028]_  | \new_[19386]_ ;
  assign \new_[15800]_  = ~\new_[16614]_ ;
  assign \new_[15801]_  = ~\new_[16351]_ ;
  assign \new_[15802]_  = ~\new_[16797]_  | ~\new_[19256]_ ;
  assign \new_[15803]_  = ~\new_[16634]_ ;
  assign \new_[15804]_  = ~\new_[16402]_ ;
  assign \new_[15805]_  = ~\new_[17239]_  & ~\new_[19162]_ ;
  assign \new_[15806]_  = ~\new_[17349]_  | ~\new_[19548]_ ;
  assign \new_[15807]_  = ~\new_[16830]_  & ~\new_[17156]_ ;
  assign \new_[15808]_  = ~\new_[15922]_ ;
  assign \new_[15809]_  = \new_[19801]_  & \new_[17032]_ ;
  assign \new_[15810]_  = ~\new_[19285]_  & ~\new_[16834]_ ;
  assign \new_[15811]_  = ~\new_[16635]_ ;
  assign \new_[15812]_  = ~\new_[18127]_  | ~\new_[21510]_ ;
  assign \new_[15813]_  = ~\new_[17413]_  | ~\new_[19386]_ ;
  assign \new_[15814]_  = ~\new_[16339]_ ;
  assign \new_[15815]_  = \\text_in_r_reg[120] ;
  assign \new_[15816]_  = ~\new_[19145]_  | ~\new_[19336]_ ;
  assign \new_[15817]_  = ~\new_[16902]_  & ~\new_[21259]_ ;
  assign \new_[15818]_  = ~\new_[18733]_  | ~\new_[19151]_ ;
  assign \new_[15819]_  = \\text_in_r_reg[84] ;
  assign \new_[15820]_  = ~\new_[16904]_  | ~\new_[19801]_ ;
  assign \new_[15821]_  = ~\new_[21306]_  | ~\new_[19267]_ ;
  assign \new_[15822]_  = \new_[18942]_  & \new_[21638]_ ;
  assign \new_[15823]_  = \\text_in_r_reg[74] ;
  assign \new_[15824]_  = ~\new_[18111]_  & ~\new_[20763]_ ;
  assign \new_[15825]_  = ~\new_[20764]_  & ~\new_[19568]_ ;
  assign \new_[15826]_  = ~\new_[15938]_ ;
  assign \new_[15827]_  = \new_[14690]_  & \new_[19253]_ ;
  assign \new_[15828]_  = ~\new_[16644]_ ;
  assign \new_[15829]_  = \new_[19203]_  & \new_[19550]_ ;
  assign \new_[15830]_  = ~\new_[17095]_  | ~\new_[19026]_ ;
  assign \new_[15831]_  = ~\new_[16627]_ ;
  assign \new_[15832]_  = ~\new_[17578]_  | ~\new_[18877]_ ;
  assign \new_[15833]_  = \new_[16763]_  & \new_[18927]_ ;
  assign \new_[15834]_  = ~\new_[16522]_ ;
  assign \new_[15835]_  = \new_[18460]_  | \new_[19780]_ ;
  assign \new_[15836]_  = ~\new_[16578]_ ;
  assign \new_[15837]_  = ~\new_[16530]_ ;
  assign \new_[15838]_  = ~\new_[16941]_  & ~\new_[19741]_ ;
  assign \new_[15839]_  = \\text_in_r_reg[16] ;
  assign \new_[15840]_  = \\text_in_r_reg[40] ;
  assign \new_[15841]_  = ~\new_[16659]_ ;
  assign \new_[15842]_  = \\text_in_r_reg[15] ;
  assign \new_[15843]_  = \\text_in_r_reg[121] ;
  assign \new_[15844]_  = ~\new_[19026]_  & ~\new_[16861]_ ;
  assign \new_[15845]_  = \\text_in_r_reg[41] ;
  assign \new_[15846]_  = \\text_in_r_reg[36] ;
  assign \new_[15847]_  = ~\new_[17019]_  | ~\new_[20487]_ ;
  assign \new_[15848]_  = ~\new_[16664]_ ;
  assign \new_[15849]_  = ~\new_[16153]_ ;
  assign \new_[15850]_  = \\text_in_r_reg[20] ;
  assign \new_[15851]_  = \\u0_r0_rcnt_reg[2] ;
  assign \new_[15852]_  = ~\new_[16781]_  | ~\new_[18408]_ ;
  assign \new_[15853]_  = \\text_in_r_reg[32] ;
  assign \new_[15854]_  = \\text_in_r_reg[75] ;
  assign \new_[15855]_  = \\text_in_r_reg[88] ;
  assign \new_[15856]_  = \new_[16833]_  & \new_[18423]_ ;
  assign \new_[15857]_  = ~\new_[17525]_  | ~\new_[18351]_ ;
  assign \new_[15858]_  = ~\new_[15978]_ ;
  assign \new_[15859]_  = ~\new_[20165]_  | ~\new_[17886]_ ;
  assign \new_[15860]_  = ~\new_[16874]_  | ~\new_[19066]_ ;
  assign \new_[15861]_  = \\text_in_r_reg[33] ;
  assign \new_[15862]_  = ~\new_[17172]_  & ~\new_[19096]_ ;
  assign \new_[15863]_  = \new_[16963]_  | \new_[18840]_ ;
  assign \new_[15864]_  = \new_[16044]_ ;
  assign \new_[15865]_  = ~\new_[17457]_  & ~\new_[19696]_ ;
  assign \new_[15866]_  = ~\new_[16698]_ ;
  assign \new_[15867]_  = ~\new_[16693]_ ;
  assign \new_[15868]_  = ~\new_[16719]_ ;
  assign \new_[15869]_  = ~\new_[21659]_  & ~\new_[21686]_ ;
  assign \new_[15870]_  = ~\new_[18002]_  & ~\new_[18190]_ ;
  assign \new_[15871]_  = ~\new_[17739]_  & ~\new_[17886]_ ;
  assign \new_[15872]_  = ~\new_[16915]_ ;
  assign \new_[15873]_  = ~\new_[17003]_ ;
  assign \new_[15874]_  = ~\new_[17953]_  & ~\new_[21306]_ ;
  assign \new_[15875]_  = ~\new_[16691]_ ;
  assign \new_[15876]_  = ~\new_[16994]_ ;
  assign \new_[15877]_  = ~\new_[16945]_ ;
  assign \new_[15878]_  = ~\new_[17761]_  | ~\new_[19098]_ ;
  assign \new_[15879]_  = ~\new_[17479]_  & ~\new_[21306]_ ;
  assign \new_[15880]_  = ~\new_[17776]_  | ~\new_[19150]_ ;
  assign \new_[15881]_  = ~\new_[17571]_  | ~\new_[19416]_ ;
  assign \new_[15882]_  = ~\new_[16733]_ ;
  assign \new_[15883]_  = ~\new_[16699]_ ;
  assign \new_[15884]_  = ~\new_[17480]_  & ~\new_[19431]_ ;
  assign \new_[15885]_  = ~\new_[21663]_ ;
  assign \new_[15886]_  = \new_[17680]_  | \new_[19589]_ ;
  assign \new_[15887]_  = ~\new_[17271]_ ;
  assign \new_[15888]_  = \new_[18998]_  & \new_[17578]_ ;
  assign \new_[15889]_  = ~\new_[17203]_ ;
  assign \new_[15890]_  = ~\new_[17485]_  & ~\new_[18959]_ ;
  assign \new_[15891]_  = ~\new_[18729]_  | ~\new_[19194]_ ;
  assign \new_[15892]_  = ~\new_[16724]_ ;
  assign \new_[15893]_  = ~\new_[19561]_ ;
  assign \new_[15894]_  = ~\new_[16729]_ ;
  assign \new_[15895]_  = ~\new_[17952]_  | ~\new_[18810]_ ;
  assign \new_[15896]_  = ~\new_[17588]_  | ~\new_[17490]_ ;
  assign \new_[15897]_  = ~\new_[17984]_  | ~\new_[19096]_ ;
  assign \new_[15898]_  = ~\new_[17202]_ ;
  assign \new_[15899]_  = ~\new_[16751]_ ;
  assign \new_[15900]_  = ~\new_[17881]_  & ~\new_[19066]_ ;
  assign \new_[15901]_  = ~\new_[16875]_ ;
  assign \new_[15902]_  = ~\new_[17909]_  | ~\new_[19321]_ ;
  assign \new_[15903]_  = ~\new_[18446]_  & ~\new_[17973]_ ;
  assign \new_[15904]_  = ~\new_[17236]_ ;
  assign \new_[15905]_  = ~\new_[21682]_  | ~\new_[19438]_ ;
  assign \new_[15906]_  = ~\new_[17533]_  & ~\new_[19446]_ ;
  assign \new_[15907]_  = ~\new_[16740]_ ;
  assign \new_[15908]_  = ~\new_[19785]_  & ~\new_[17467]_ ;
  assign \new_[15909]_  = ~\new_[16745]_ ;
  assign \new_[15910]_  = ~\new_[21654]_  | ~\new_[19353]_ ;
  assign \new_[15911]_  = ~\new_[18023]_  | ~\new_[17765]_ ;
  assign \new_[15912]_  = ~\new_[16756]_ ;
  assign \new_[15913]_  = ~\new_[17992]_  & ~\new_[19782]_ ;
  assign \new_[15914]_  = ~\new_[17569]_  & ~\new_[19301]_ ;
  assign \new_[15915]_  = ~\new_[17631]_  & ~\new_[19379]_ ;
  assign \new_[15916]_  = ~\new_[16753]_ ;
  assign \new_[15917]_  = ~\new_[16749]_ ;
  assign \new_[15918]_  = ~\new_[18920]_  | ~\new_[19116]_ ;
  assign \new_[15919]_  = ~\new_[17067]_ ;
  assign \new_[15920]_  = \new_[17684]_  & \new_[19754]_ ;
  assign \new_[15921]_  = ~\new_[17718]_  & ~\new_[19676]_ ;
  assign \new_[15922]_  = ~\new_[17026]_ ;
  assign \new_[15923]_  = ~\new_[19308]_ ;
  assign \new_[15924]_  = ~\new_[16766]_ ;
  assign \new_[15925]_  = ~\new_[17372]_ ;
  assign \new_[15926]_  = ~\new_[17316]_ ;
  assign \new_[15927]_  = \new_[17683]_  | \new_[17622]_ ;
  assign \new_[15928]_  = ~\new_[17661]_  | ~\new_[19052]_ ;
  assign \new_[15929]_  = ~\new_[16739]_ ;
  assign \new_[15930]_  = \new_[19098]_  | \new_[18699]_ ;
  assign \new_[15931]_  = ~\new_[17010]_ ;
  assign \new_[15932]_  = \new_[18648]_  | \new_[19085]_ ;
  assign \new_[15933]_  = ~\new_[17738]_  & ~\new_[21306]_ ;
  assign \new_[15934]_  = ~\new_[17029]_ ;
  assign \new_[15935]_  = ~\new_[21711]_  | ~\new_[18614]_ ;
  assign \new_[15936]_  = ~\new_[17957]_  & ~\new_[19568]_ ;
  assign \new_[15937]_  = \new_[17542]_  & \new_[19176]_ ;
  assign \new_[15938]_  = \new_[18271]_  & \new_[19476]_ ;
  assign \new_[15939]_  = ~\new_[17114]_ ;
  assign \new_[15940]_  = ~\new_[17178]_ ;
  assign \new_[15941]_  = ~\new_[16784]_ ;
  assign \new_[15942]_  = ~\new_[17557]_  | ~\new_[19066]_ ;
  assign \new_[15943]_  = ~\new_[16798]_ ;
  assign \new_[15944]_  = ~\new_[16769]_ ;
  assign \new_[15945]_  = ~\new_[21096]_ ;
  assign \new_[15946]_  = ~\new_[17558]_  & ~\new_[19268]_ ;
  assign \new_[15947]_  = ~\new_[17521]_  & ~\new_[21542]_ ;
  assign \new_[15948]_  = \new_[17199]_ ;
  assign \new_[15949]_  = ~\new_[17685]_  | ~\new_[19319]_ ;
  assign \new_[15950]_  = ~\new_[16821]_ ;
  assign \new_[15951]_  = ~\new_[17515]_ ;
  assign \new_[15952]_  = \new_[17747]_  | \new_[19117]_ ;
  assign \new_[15953]_  = ~\new_[17504]_  & ~\new_[19434]_ ;
  assign \new_[15954]_  = ~\new_[19308]_  & ~\new_[18209]_ ;
  assign \new_[15955]_  = ~\new_[17515]_ ;
  assign \new_[15956]_  = ~\new_[16959]_ ;
  assign \new_[15957]_  = ~\new_[16804]_ ;
  assign \new_[15958]_  = ~\new_[17197]_ ;
  assign \new_[15959]_  = ~\new_[16823]_ ;
  assign \new_[15960]_  = ~\new_[21713]_  | ~\new_[19198]_ ;
  assign \new_[15961]_  = ~\new_[16929]_ ;
  assign \new_[15962]_  = ~\new_[16814]_ ;
  assign \new_[15963]_  = ~\new_[16889]_ ;
  assign \new_[15964]_  = ~\new_[17676]_  | ~\new_[18903]_ ;
  assign \new_[15965]_  = ~\new_[17750]_  & ~\new_[18857]_ ;
  assign \new_[15966]_  = ~\new_[17632]_  & ~\new_[19186]_ ;
  assign \new_[15967]_  = ~\new_[17864]_  & ~\new_[18573]_ ;
  assign \new_[15968]_  = ~\new_[16816]_ ;
  assign \new_[15969]_  = ~\new_[17176]_ ;
  assign \new_[15970]_  = ~\new_[17243]_ ;
  assign \new_[15971]_  = \new_[18935]_  & \new_[18906]_ ;
  assign \new_[15972]_  = ~\new_[16737]_ ;
  assign \new_[15973]_  = ~\new_[17563]_  | ~\new_[19734]_ ;
  assign \new_[15974]_  = ~\new_[18001]_  & ~\new_[18151]_ ;
  assign \new_[15975]_  = ~\new_[17771]_  & ~\new_[19066]_ ;
  assign \new_[15976]_  = ~\new_[16981]_ ;
  assign \new_[15977]_  = ~\new_[17574]_ ;
  assign \new_[15978]_  = ~\new_[17821]_  & ~\new_[19681]_ ;
  assign \new_[15979]_  = ~\new_[17928]_  | ~\new_[18235]_ ;
  assign \new_[15980]_  = ~\new_[19782]_  & ~\new_[17865]_ ;
  assign \new_[15981]_  = ~\new_[18362]_  & ~\new_[18285]_ ;
  assign \new_[15982]_  = ~\new_[18396]_  & ~\new_[19253]_ ;
  assign \new_[15983]_  = ~\new_[17076]_ ;
  assign \new_[15984]_  = ~\new_[16828]_ ;
  assign \new_[15985]_  = ~\new_[17196]_ ;
  assign \new_[15986]_  = ~\new_[18598]_  | ~\new_[19478]_ ;
  assign \new_[15987]_  = ~\new_[17220]_ ;
  assign \new_[15988]_  = ~\new_[17665]_  & ~\new_[21688]_ ;
  assign \new_[15989]_  = \new_[18259]_  | \new_[18020]_ ;
  assign \new_[15990]_  = ~\new_[19823]_  | ~\new_[18664]_ ;
  assign \new_[15991]_  = ~\new_[16842]_ ;
  assign \new_[15992]_  = ~\new_[19251]_  & ~\new_[17649]_ ;
  assign \new_[15993]_  = ~\new_[17463]_  | ~\new_[19676]_ ;
  assign \new_[15994]_  = ~\new_[16893]_ ;
  assign \new_[15995]_  = ~\new_[19741]_  & ~\new_[17672]_ ;
  assign \new_[15996]_  = ~\new_[16843]_ ;
  assign \new_[15997]_  = ~\new_[17174]_ ;
  assign \new_[15998]_  = ~\new_[17547]_  | ~\new_[19782]_ ;
  assign \new_[15999]_  = ~\new_[17455]_ ;
  assign \new_[16000]_  = ~\new_[17254]_ ;
  assign \new_[16001]_  = ~\new_[17915]_  & ~\new_[18408]_ ;
  assign \new_[16002]_  = \new_[17886]_  & \new_[18663]_ ;
  assign \new_[16003]_  = \new_[18812]_  | \new_[19676]_ ;
  assign \new_[16004]_  = ~\new_[17249]_ ;
  assign \new_[16005]_  = \new_[17526]_  & \new_[21569]_ ;
  assign \new_[16006]_  = ~\new_[17736]_  & ~\new_[18938]_ ;
  assign \new_[16007]_  = ~\new_[16855]_ ;
  assign \new_[16008]_  = ~\new_[17990]_  & ~\new_[19186]_ ;
  assign \new_[16009]_  = ~\new_[16858]_ ;
  assign \new_[16010]_  = ~\new_[17923]_  & ~\new_[18947]_ ;
  assign \new_[16011]_  = ~\new_[17935]_  | ~\new_[18811]_ ;
  assign \new_[16012]_  = ~\new_[20165]_ ;
  assign \new_[16013]_  = ~\new_[17330]_ ;
  assign \new_[16014]_  = \new_[17584]_  | \new_[19738]_ ;
  assign \new_[16015]_  = ~\new_[17311]_ ;
  assign \new_[16016]_  = ~\new_[17079]_ ;
  assign \new_[16017]_  = ~\new_[16999]_ ;
  assign \new_[16018]_  = ~\new_[17933]_ ;
  assign \new_[16019]_  = \new_[17719]_  & \new_[19301]_ ;
  assign \new_[16020]_  = ~\new_[18308]_  & ~\new_[18842]_ ;
  assign \new_[16021]_  = ~\new_[17361]_ ;
  assign \new_[16022]_  = ~\new_[17063]_ ;
  assign \new_[16023]_  = ~\new_[17613]_  & ~\new_[19416]_ ;
  assign \new_[16024]_  = ~\new_[17621]_  | ~\new_[20699]_ ;
  assign \new_[16025]_  = ~\new_[16870]_ ;
  assign \new_[16026]_  = ~\new_[16872]_ ;
  assign \new_[16027]_  = ~\new_[16941]_ ;
  assign \new_[16028]_  = ~\new_[17142]_ ;
  assign \new_[16029]_  = ~\new_[17266]_ ;
  assign \new_[16030]_  = ~\new_[18885]_  & ~\new_[20865]_ ;
  assign \new_[16031]_  = ~\new_[17588]_  | ~\new_[19081]_ ;
  assign \new_[16032]_  = ~\new_[17937]_  | ~\new_[21572]_ ;
  assign \new_[16033]_  = ~\new_[17830]_  & ~\new_[18998]_ ;
  assign \new_[16034]_  = ~\new_[20868]_  & ~\new_[20239]_ ;
  assign \new_[16035]_  = ~\new_[17045]_ ;
  assign \new_[16036]_  = ~\new_[17313]_ ;
  assign \new_[16037]_  = ~\new_[17857]_  & ~\new_[19655]_ ;
  assign \new_[16038]_  = ~\new_[18964]_  & ~\new_[19824]_ ;
  assign \new_[16039]_  = ~\new_[16891]_ ;
  assign \new_[16040]_  = \new_[17644]_  | \new_[19298]_ ;
  assign \new_[16041]_  = ~\new_[16898]_ ;
  assign \new_[16042]_  = ~\new_[16904]_ ;
  assign \new_[16043]_  = \new_[17623]_  | \new_[18577]_ ;
  assign \new_[16044]_  = ~\new_[17456]_ ;
  assign \new_[16045]_  = ~\new_[17966]_  & ~\new_[18906]_ ;
  assign \new_[16046]_  = ~\new_[17060]_ ;
  assign \new_[16047]_  = ~\new_[16762]_ ;
  assign \new_[16048]_  = ~\new_[18375]_ ;
  assign \new_[16049]_  = ~\new_[17354]_ ;
  assign \new_[16050]_  = ~\new_[17670]_  & ~\new_[18607]_ ;
  assign \new_[16051]_  = ~\new_[16903]_ ;
  assign \new_[16052]_  = ~\new_[16750]_ ;
  assign \new_[16053]_  = ~\new_[17735]_  & ~\new_[19095]_ ;
  assign \new_[16054]_  = \new_[17548]_  | \new_[19444]_ ;
  assign \new_[16055]_  = ~\new_[18489]_  | ~\new_[17540]_ ;
  assign \new_[16056]_  = ~\new_[17870]_  & ~\new_[19162]_ ;
  assign \new_[16057]_  = ~\new_[17534]_  & ~\new_[21259]_ ;
  assign \new_[16058]_  = ~\new_[17269]_ ;
  assign \new_[16059]_  = ~\new_[16786]_ ;
  assign \new_[16060]_  = ~\new_[17695]_  | ~\new_[18984]_ ;
  assign \new_[16061]_  = \new_[17609]_  & \new_[19664]_ ;
  assign \new_[16062]_  = ~\new_[18201]_ ;
  assign \new_[16063]_  = ~\new_[17535]_  | ~\new_[19068]_ ;
  assign \new_[16064]_  = ~\new_[17169]_ ;
  assign \new_[16065]_  = ~\new_[19679]_  & ~\new_[17995]_ ;
  assign \new_[16066]_  = ~\new_[19096]_  & ~\new_[20931]_ ;
  assign \new_[16067]_  = ~\new_[17995]_  & ~\new_[18974]_ ;
  assign \new_[16068]_  = ~\new_[16720]_ ;
  assign \new_[16069]_  = ~\new_[17850]_  & ~\new_[18607]_ ;
  assign \new_[16070]_  = ~\new_[17981]_  & ~\new_[18605]_ ;
  assign \new_[16071]_  = ~\new_[17985]_  & ~\new_[18008]_ ;
  assign \new_[16072]_  = ~\new_[17956]_  | ~\new_[21328]_ ;
  assign \new_[16073]_  = ~\new_[17567]_  & ~\new_[21685]_ ;
  assign \new_[16074]_  = \new_[17802]_  | \new_[19018]_ ;
  assign \new_[16075]_  = ~\new_[17040]_ ;
  assign \new_[16076]_  = ~\new_[17034]_ ;
  assign \new_[16077]_  = \new_[17625]_  | \new_[19547]_ ;
  assign \new_[16078]_  = ~\new_[17492]_  & ~\new_[18616]_ ;
  assign \new_[16079]_  = \new_[17583]_  | \new_[17593]_ ;
  assign \new_[16080]_  = ~\new_[16899]_ ;
  assign \new_[16081]_  = ~\new_[17107]_ ;
  assign \new_[16082]_  = ~\new_[21259]_  | ~\new_[17752]_ ;
  assign \new_[16083]_  = \new_[15839]_  ^ \new_[19563]_ ;
  assign \new_[16084]_  = ~\new_[17192]_ ;
  assign \new_[16085]_  = ~\new_[17736]_  & ~\new_[19675]_ ;
  assign \new_[16086]_  = ~\new_[16983]_ ;
  assign \new_[16087]_  = ~\new_[17210]_ ;
  assign \new_[16088]_  = ~\new_[17349]_ ;
  assign \new_[16089]_  = ~\new_[17216]_ ;
  assign \new_[16090]_  = ~\new_[17314]_ ;
  assign \new_[16091]_  = \new_[17621]_  & \new_[21513]_ ;
  assign \new_[16092]_  = ~\new_[17088]_ ;
  assign \new_[16093]_  = ~\new_[16897]_ ;
  assign \new_[16094]_  = ~\new_[17934]_  | ~\new_[19675]_ ;
  assign \new_[16095]_  = ~\new_[16946]_ ;
  assign \new_[16096]_  = ~\new_[17965]_  & ~\new_[19426]_ ;
  assign \new_[16097]_  = ~\new_[16865]_ ;
  assign \new_[16098]_  = ~\new_[17513]_  & ~\new_[19268]_ ;
  assign \new_[16099]_  = ~\new_[18189]_  & ~\new_[21529]_ ;
  assign \new_[16100]_  = ~\new_[17606]_  | ~\new_[19023]_ ;
  assign \new_[16101]_  = ~\new_[16839]_ ;
  assign \new_[16102]_  = ~\new_[16783]_ ;
  assign \new_[16103]_  = ~\new_[19874]_ ;
  assign \new_[16104]_  = ~\new_[17101]_ ;
  assign \new_[16105]_  = \new_[18729]_  & \new_[18008]_ ;
  assign \new_[16106]_  = ~\new_[17516]_  & ~\new_[17457]_ ;
  assign \new_[16107]_  = \new_[17048]_ ;
  assign \new_[16108]_  = ~\new_[17251]_ ;
  assign \new_[16109]_  = ~\new_[17703]_  & ~\new_[17886]_ ;
  assign \new_[16110]_  = \new_[17599]_  & \new_[19637]_ ;
  assign \new_[16111]_  = ~\new_[17858]_  & ~\new_[19801]_ ;
  assign \new_[16112]_  = ~\new_[17788]_  | ~\new_[21570]_ ;
  assign \new_[16113]_  = ~\new_[17550]_  & ~\new_[19801]_ ;
  assign \new_[16114]_  = \new_[18018]_  | \new_[19203]_ ;
  assign \new_[16115]_  = ~\new_[16990]_ ;
  assign \new_[16116]_  = ~\new_[17690]_  & ~\new_[19335]_ ;
  assign \new_[16117]_  = ~\new_[18398]_  | ~\new_[19299]_ ;
  assign \new_[16118]_  = ~\new_[17706]_  & ~\new_[19782]_ ;
  assign \new_[16119]_  = ~\new_[17164]_ ;
  assign \new_[16120]_  = \new_[17855]_  & \new_[19589]_ ;
  assign \new_[16121]_  = \new_[17625]_  | \new_[19098]_ ;
  assign \new_[16122]_  = \new_[17772]_  | \new_[19156]_ ;
  assign \new_[16123]_  = ~\new_[17139]_ ;
  assign \new_[16124]_  = ~\new_[17620]_  | ~\new_[19727]_ ;
  assign \new_[16125]_  = \new_[17756]_  | \new_[19727]_ ;
  assign \new_[16126]_  = ~\new_[17036]_ ;
  assign \new_[16127]_  = ~\new_[17661]_  | ~\new_[19026]_ ;
  assign \new_[16128]_  = ~\new_[18842]_  | ~\new_[19198]_  | ~\new_[18398]_ ;
  assign \new_[16129]_  = ~\new_[17646]_  & ~\new_[19676]_ ;
  assign \new_[16130]_  = \new_[19874]_ ;
  assign \new_[16131]_  = \new_[19874]_ ;
  assign \new_[16132]_  = ~\new_[17914]_  & ~\new_[19319]_ ;
  assign \new_[16133]_  = ~\new_[17625]_  & ~\new_[19033]_ ;
  assign \new_[16134]_  = ~\new_[17637]_  & ~\new_[18784]_ ;
  assign \new_[16135]_  = \new_[17650]_  & \new_[19676]_ ;
  assign \new_[16136]_  = ~\new_[20867]_ ;
  assign \new_[16137]_  = ~\new_[17000]_ ;
  assign \new_[16138]_  = ~\new_[17687]_  | ~\new_[19219]_ ;
  assign \new_[16139]_  = \new_[17756]_  | \new_[19319]_ ;
  assign \new_[16140]_  = ~\new_[17268]_ ;
  assign \new_[16141]_  = \new_[17722]_  | \new_[19290]_ ;
  assign \new_[16142]_  = ~\new_[17860]_  | ~\new_[19115]_ ;
  assign \new_[16143]_  = ~\new_[17871]_  | ~\new_[21259]_ ;
  assign \new_[16144]_  = ~\new_[17026]_ ;
  assign \new_[16145]_  = ~\new_[17284]_ ;
  assign \new_[16146]_  = ~\new_[18785]_  | ~\new_[18036]_  | ~\new_[21490]_ ;
  assign \new_[16147]_  = ~\new_[17712]_  & ~\new_[19779]_ ;
  assign \new_[16148]_  = ~\new_[17307]_ ;
  assign \new_[16149]_  = ~\new_[17661]_  | ~\new_[19303]_ ;
  assign \new_[16150]_  = ~\new_[17877]_  | ~\new_[19176]_ ;
  assign \new_[16151]_  = ~\new_[18013]_  | ~\new_[19663]_ ;
  assign \new_[16152]_  = ~\new_[16767]_ ;
  assign \new_[16153]_  = ~\new_[17963]_  & ~\new_[19096]_ ;
  assign \new_[16154]_  = ~\new_[17026]_ ;
  assign \new_[16155]_  = ~\new_[17632]_  & ~\new_[19438]_ ;
  assign \new_[16156]_  = ~\new_[17169]_ ;
  assign \new_[16157]_  = ~\new_[17058]_ ;
  assign \new_[16158]_  = ~\new_[17870]_  & ~\new_[18979]_ ;
  assign \new_[16159]_  = ~\new_[18838]_  | ~\new_[18832]_ ;
  assign \new_[16160]_  = ~\new_[17912]_  | ~\new_[18664]_ ;
  assign \new_[16161]_  = ~\new_[16748]_ ;
  assign \new_[16162]_  = ~\new_[16778]_ ;
  assign \new_[16163]_  = ~\new_[18007]_  & ~\new_[19637]_ ;
  assign \new_[16164]_  = ~\new_[17717]_  | ~\new_[21502]_ ;
  assign \new_[16165]_  = ~\new_[17802]_  & ~\new_[19096]_ ;
  assign \new_[16166]_  = ~\new_[18003]_  | ~\new_[19253]_ ;
  assign \new_[16167]_  = \new_[17498]_  & \new_[19082]_ ;
  assign \new_[16168]_  = ~\new_[17466]_  & ~\new_[19637]_ ;
  assign \new_[16169]_  = ~\new_[18877]_  | ~\new_[18741]_  | ~\new_[19425]_  | ~\new_[19213]_ ;
  assign \new_[16170]_  = ~\new_[19255]_  & ~\new_[17673]_ ;
  assign \new_[16171]_  = ~\new_[16825]_ ;
  assign \new_[16172]_  = ~\new_[16859]_ ;
  assign \new_[16173]_  = \new_[17914]_  | \new_[19288]_ ;
  assign \new_[16174]_  = ~\new_[20868]_  & ~\new_[18964]_ ;
  assign \new_[16175]_  = ~\new_[17828]_  | ~\new_[18995]_ ;
  assign \new_[16176]_  = ~\new_[16727]_ ;
  assign \new_[16177]_  = ~\new_[17039]_ ;
  assign \new_[16178]_  = \new_[17992]_  | \new_[17979]_ ;
  assign \new_[16179]_  = ~\new_[18686]_  & ~\new_[19409]_ ;
  assign \new_[16180]_  = ~\new_[19801]_  | ~\new_[17737]_ ;
  assign \new_[16181]_  = ~\new_[18016]_  & ~\new_[19219]_ ;
  assign \new_[16182]_  = ~\new_[17158]_ ;
  assign \new_[16183]_  = ~\new_[16720]_ ;
  assign \new_[16184]_  = \new_[17687]_  & \new_[19538]_ ;
  assign \new_[16185]_  = ~\new_[17978]_  | ~\new_[18140]_ ;
  assign \new_[16186]_  = ~\new_[17019]_ ;
  assign \new_[16187]_  = ~\new_[18000]_  | ~\new_[19386]_ ;
  assign \new_[16188]_  = ~\new_[17645]_  | ~\new_[18209]_ ;
  assign \new_[16189]_  = ~\new_[17839]_  & ~\new_[18637]_ ;
  assign \new_[16190]_  = ~\new_[17906]_  & ~\new_[19353]_ ;
  assign \new_[16191]_  = ~\new_[17104]_ ;
  assign \new_[16192]_  = \new_[17857]_  | \new_[19290]_ ;
  assign \new_[16193]_  = ~\new_[17638]_  & ~\new_[19409]_ ;
  assign \new_[16194]_  = ~\new_[16986]_ ;
  assign \new_[16195]_  = ~\new_[17711]_  | ~\new_[20487]_ ;
  assign \new_[16196]_  = ~\new_[17655]_  | ~\new_[19555]_ ;
  assign \new_[16197]_  = ~\new_[17109]_ ;
  assign \new_[16198]_  = ~\new_[17822]_  & ~\new_[19676]_ ;
  assign \new_[16199]_  = \new_[17460]_  | \new_[18938]_ ;
  assign \new_[16200]_  = ~\new_[19084]_  & ~\new_[17804]_ ;
  assign \new_[16201]_  = ~\new_[17751]_  | ~\new_[19801]_ ;
  assign \new_[16202]_  = ~\new_[17068]_ ;
  assign \new_[16203]_  = ~\new_[17322]_ ;
  assign \new_[16204]_  = \new_[17670]_  | \new_[18414]_ ;
  assign \new_[16205]_  = ~\new_[17072]_ ;
  assign \new_[16206]_  = ~\new_[16750]_ ;
  assign \new_[16207]_  = ~\new_[17816]_  | ~\new_[18682]_ ;
  assign \new_[16208]_  = ~\new_[16727]_ ;
  assign \new_[16209]_  = ~\new_[17090]_ ;
  assign \new_[16210]_  = ~\new_[18454]_  | ~\new_[21631]_  | ~\new_[18392]_ ;
  assign \new_[16211]_  = ~\new_[17229]_ ;
  assign \new_[16212]_  = ~\new_[18332]_  | ~\new_[17460]_ ;
  assign \new_[16213]_  = ~\new_[17112]_ ;
  assign \new_[16214]_  = ~\new_[20764]_ ;
  assign \new_[16215]_  = ~\new_[20494]_ ;
  assign \new_[16216]_  = ~\new_[20298]_  & ~\new_[19782]_ ;
  assign \new_[16217]_  = ~\new_[17509]_  | ~\new_[19158]_ ;
  assign \new_[16218]_  = ~\new_[17473]_  | ~\new_[19409]_ ;
  assign \new_[16219]_  = ~\new_[17881]_  & ~\new_[19253]_ ;
  assign \new_[16220]_  = ~\new_[19874]_ ;
  assign \new_[16221]_  = ~\new_[17026]_ ;
  assign \new_[16222]_  = \new_[17863]_  | \new_[19319]_ ;
  assign \new_[16223]_  = ~\new_[17152]_ ;
  assign \new_[16224]_  = ~\new_[17979]_  | ~\new_[20586]_ ;
  assign \new_[16225]_  = ~\new_[17865]_  & ~\new_[19268]_ ;
  assign \new_[16226]_  = \new_[17830]_  | \new_[19290]_ ;
  assign \new_[16227]_  = ~\new_[19624]_  & ~\new_[17826]_ ;
  assign \new_[16228]_  = ~\new_[19444]_  | ~\new_[17994]_ ;
  assign \new_[16229]_  = ~\new_[17596]_  | ~\new_[19750]_ ;
  assign \new_[16230]_  = ~\new_[17510]_  & ~\new_[19023]_ ;
  assign \new_[16231]_  = ~\new_[17999]_  | ~\new_[19265]_ ;
  assign \new_[16232]_  = ~\new_[17937]_  | ~\new_[21049]_ ;
  assign \new_[16233]_  = ~\new_[18968]_  | ~\new_[21077]_ ;
  assign \new_[16234]_  = ~\new_[17762]_  & ~\new_[21506]_ ;
  assign \new_[16235]_  = ~\new_[17133]_ ;
  assign \new_[16236]_  = ~\new_[17630]_  & ~\new_[18959]_ ;
  assign \new_[16237]_  = ~\new_[17131]_ ;
  assign \new_[16238]_  = ~\new_[18945]_  | ~\new_[17808]_ ;
  assign \new_[16239]_  = ~\new_[17731]_  & ~\new_[18903]_ ;
  assign \new_[16240]_  = ~\new_[17834]_  & ~\new_[19719]_ ;
  assign \new_[16241]_  = ~\new_[17138]_ ;
  assign \new_[16242]_  = ~\new_[18037]_  | ~\new_[21608]_ ;
  assign \new_[16243]_  = ~\new_[21572]_  | ~\new_[17728]_ ;
  assign \new_[16244]_  = ~\new_[17755]_  & ~\new_[18012]_ ;
  assign \new_[16245]_  = ~\new_[17834]_  & ~\new_[17979]_ ;
  assign \new_[16246]_  = \new_[17693]_  | \new_[20239]_ ;
  assign \new_[16247]_  = ~\new_[17876]_  & ~\new_[19675]_ ;
  assign n2763 = ~\new_[16878]_ ;
  assign \new_[16249]_  = ~\new_[17805]_  & ~\new_[21574]_ ;
  assign \new_[16250]_  = ~\new_[18587]_  & ~\new_[19028]_  & ~\new_[18164]_ ;
  assign \new_[16251]_  = \new_[17787]_  | \new_[18832]_ ;
  assign \new_[16252]_  = ~\new_[17826]_  & ~\new_[19084]_ ;
  assign \new_[16253]_  = ~\new_[17641]_  & ~\new_[19655]_ ;
  assign \new_[16254]_  = ~\new_[17617]_  & ~\new_[19064]_ ;
  assign \new_[16255]_  = ~\new_[17774]_  & ~\new_[19156]_ ;
  assign \new_[16256]_  = \new_[17718]_  | \new_[18832]_ ;
  assign \new_[16257]_  = ~\new_[21529]_  | ~\new_[19219]_ ;
  assign \new_[16258]_  = \new_[17835]_  & \new_[19044]_ ;
  assign \new_[16259]_  = ~\new_[17674]_  | ~\new_[19068]_ ;
  assign \new_[16260]_  = ~\new_[16864]_ ;
  assign \new_[16261]_  = ~\new_[17782]_  & ~\new_[19779]_ ;
  assign \new_[16262]_  = ~\new_[19251]_  | ~\new_[17800]_ ;
  assign \new_[16263]_  = ~\new_[17793]_  | ~\new_[18496]_ ;
  assign \new_[16264]_  = ~\new_[17958]_  & ~\new_[19689]_ ;
  assign \new_[16265]_  = ~\new_[17933]_  & ~\new_[19182]_ ;
  assign \new_[16266]_  = \new_[17675]_  | \new_[19589]_ ;
  assign \new_[16267]_  = ~\new_[17511]_  & ~\new_[18973]_ ;
  assign \new_[16268]_  = \new_[17491]_  | \new_[19456]_ ;
  assign \new_[16269]_  = ~\new_[17573]_  & ~\new_[17625]_ ;
  assign \new_[16270]_  = ~\new_[17483]_  | ~\new_[18489]_ ;
  assign \new_[16271]_  = ~\new_[17733]_  & ~\new_[19750]_ ;
  assign \new_[16272]_  = \new_[17816]_  | \new_[19196]_ ;
  assign \new_[16273]_  = ~\new_[17219]_ ;
  assign \new_[16274]_  = \new_[19775]_  ^ \new_[19552]_ ;
  assign \new_[16275]_  = ~\new_[16738]_ ;
  assign \new_[16276]_  = ~\new_[16683]_ ;
  assign \new_[16277]_  = \new_[17565]_  | \new_[21511]_ ;
  assign \new_[16278]_  = ~\new_[17499]_  | ~\new_[21306]_ ;
  assign \new_[16279]_  = ~\new_[17081]_ ;
  assign \new_[16280]_  = \new_[17884]_  | \new_[19130]_ ;
  assign \new_[16281]_  = \new_[17988]_  | \new_[19052]_ ;
  assign \new_[16282]_  = ~\new_[17062]_ ;
  assign \new_[16283]_  = ~\new_[17186]_ ;
  assign \new_[16284]_  = ~\new_[17602]_  & ~\new_[19719]_ ;
  assign \new_[16285]_  = ~\new_[19112]_  & ~\new_[19780]_ ;
  assign \new_[16286]_  = ~\new_[16704]_ ;
  assign \new_[16287]_  = ~\new_[18771]_  & ~\new_[19024]_ ;
  assign \new_[16288]_  = ~\new_[16919]_ ;
  assign \new_[16289]_  = ~\new_[16808]_ ;
  assign \new_[16290]_  = ~\new_[17166]_ ;
  assign \new_[16291]_  = ~\new_[17100]_ ;
  assign \new_[16292]_  = ~\new_[17167]_ ;
  assign \new_[16293]_  = ~\new_[16947]_ ;
  assign \new_[16294]_  = ~\new_[18933]_  & ~\new_[19082]_ ;
  assign \new_[16295]_  = ~\new_[17014]_ ;
  assign \new_[16296]_  = ~\new_[17168]_ ;
  assign \new_[16297]_  = ~\new_[17058]_ ;
  assign \new_[16298]_  = ~\new_[17107]_ ;
  assign \new_[16299]_  = ~\new_[18015]_  & ~\new_[18605]_ ;
  assign \new_[16300]_  = ~\new_[17225]_ ;
  assign \new_[16301]_  = ~\new_[17450]_ ;
  assign \new_[16302]_  = ~\new_[17560]_  & ~\new_[19181]_ ;
  assign \new_[16303]_  = ~\new_[17873]_  | ~\new_[19385]_ ;
  assign \new_[16304]_  = ~\new_[18340]_  | ~\new_[18704]_ ;
  assign \new_[16305]_  = ~\new_[16956]_ ;
  assign \new_[16306]_  = ~\new_[17962]_  & ~\new_[19426]_ ;
  assign \new_[16307]_  = ~\new_[17828]_  | ~\new_[19269]_ ;
  assign \new_[16308]_  = ~\new_[16687]_ ;
  assign \new_[16309]_  = ~\new_[16921]_ ;
  assign \new_[16310]_  = \new_[17986]_  | \new_[21501]_ ;
  assign \new_[16311]_  = ~\new_[16907]_ ;
  assign \new_[16312]_  = ~\new_[17828]_  | ~\new_[19270]_ ;
  assign \new_[16313]_  = ~\new_[18585]_  | ~\new_[17651]_ ;
  assign \new_[16314]_  = ~\new_[17490]_  | ~\new_[18083]_ ;
  assign \new_[16315]_  = ~\new_[17987]_  & ~\new_[17886]_ ;
  assign \new_[16316]_  = ~\new_[17171]_ ;
  assign \new_[16317]_  = ~\new_[17950]_  & ~\new_[21695]_ ;
  assign \new_[16318]_  = ~\new_[16880]_ ;
  assign \new_[16319]_  = ~\new_[17084]_ ;
  assign \new_[16320]_  = \new_[18735]_  | \new_[19033]_ ;
  assign \new_[16321]_  = ~\new_[17172]_ ;
  assign \new_[16322]_  = \new_[17619]_  | \new_[19176]_ ;
  assign \new_[16323]_  = ~\new_[16881]_ ;
  assign \new_[16324]_  = ~\new_[17973]_  & ~\new_[19386]_ ;
  assign \new_[16325]_  = ~\new_[16805]_ ;
  assign \new_[16326]_  = \new_[18617]_  | \new_[19152]_ ;
  assign \new_[16327]_  = ~\new_[17622]_  | ~\new_[19782]_ ;
  assign \new_[16328]_  = ~\new_[17513]_ ;
  assign \new_[16329]_  = ~\new_[17920]_  & (~\new_[18813]_  | ~\new_[10818]_ );
  assign \new_[16330]_  = ~\new_[17178]_ ;
  assign \new_[16331]_  = ~\new_[16765]_ ;
  assign \new_[16332]_  = ~\new_[17073]_ ;
  assign \new_[16333]_  = ~\new_[17911]_  | ~\new_[21259]_ ;
  assign \new_[16334]_  = ~\new_[17932]_  & ~\new_[18121]_ ;
  assign \new_[16335]_  = ~\new_[17593]_  & ~\new_[21306]_ ;
  assign \new_[16336]_  = ~\new_[17651]_  | ~\new_[21513]_ ;
  assign \new_[16337]_  = ~\new_[17145]_ ;
  assign \new_[16338]_  = ~\new_[17405]_ ;
  assign \new_[16339]_  = ~\new_[17185]_ ;
  assign \new_[16340]_  = ~\new_[17565]_  | ~\new_[17986]_ ;
  assign \new_[16341]_  = ~\new_[17267]_ ;
  assign \new_[16342]_  = ~\new_[17804]_  & ~\new_[18542]_ ;
  assign \new_[16343]_  = ~\new_[17610]_  & ~\new_[19385]_ ;
  assign \new_[16344]_  = ~\new_[17975]_  & ~\new_[18852]_ ;
  assign \new_[16345]_  = ~\new_[17768]_  | ~\new_[21572]_ ;
  assign \new_[16346]_  = ~\new_[16937]_ ;
  assign \new_[16347]_  = ~\new_[17766]_  & ~\new_[18362]_ ;
  assign \new_[16348]_  = ~\new_[16987]_ ;
  assign \new_[16349]_  = ~\new_[17489]_  | ~\new_[19779]_ ;
  assign \new_[16350]_  = ~\new_[17049]_ ;
  assign \new_[16351]_  = ~\new_[17579]_  & ~\new_[19664]_ ;
  assign \new_[16352]_  = ~\new_[17591]_  | ~\new_[20699]_ ;
  assign \new_[16353]_  = \new_[17515]_  | \new_[19642]_ ;
  assign \new_[16354]_  = ~\new_[21571]_  & ~\new_[17848]_ ;
  assign \new_[16355]_  = ~\new_[16746]_ ;
  assign \new_[16356]_  = ~\new_[18078]_  | ~\new_[18496]_ ;
  assign \new_[16357]_  = ~\new_[16686]_ ;
  assign \new_[16358]_  = ~\new_[17938]_  | ~\new_[19104]_ ;
  assign \new_[16359]_  = ~\new_[18439]_  & ~\new_[18019]_ ;
  assign \new_[16360]_  = ~\new_[17587]_  | ~\new_[18966]_ ;
  assign \new_[16361]_  = ~\new_[17527]_  & ~\new_[18974]_ ;
  assign \new_[16362]_  = ~\new_[17190]_ ;
  assign \new_[16363]_  = ~\new_[17038]_ ;
  assign \new_[16364]_  = ~\new_[18570]_  | ~\new_[17597]_ ;
  assign \new_[16365]_  = \new_[17498]_  | \new_[18420]_ ;
  assign \new_[16366]_  = \new_[17916]_  & \new_[21328]_ ;
  assign \new_[16367]_  = ~\new_[17007]_ ;
  assign \new_[16368]_  = ~\new_[17825]_  | ~\new_[19719]_ ;
  assign \new_[16369]_  = ~\new_[16928]_ ;
  assign \new_[16370]_  = ~\new_[18392]_  | ~\new_[21653]_ ;
  assign \new_[16371]_  = ~\new_[17622]_  | ~\new_[18807]_ ;
  assign \new_[16372]_  = ~\new_[17212]_ ;
  assign \new_[16373]_  = ~\new_[17589]_  | ~\new_[19000]_ ;
  assign \new_[16374]_  = ~\new_[18869]_  | ~\new_[18271]_ ;
  assign \new_[16375]_  = ~\new_[17025]_ ;
  assign \new_[16376]_  = \new_[18590]_  & \new_[19550]_ ;
  assign \new_[16377]_  = ~\new_[17601]_  | ~\new_[18972]_ ;
  assign \new_[16378]_  = ~\new_[17511]_  | ~\new_[18421]_ ;
  assign \new_[16379]_  = ~\new_[17535]_  | ~\new_[19741]_ ;
  assign \new_[16380]_  = ~\new_[16810]_ ;
  assign \new_[16381]_  = \new_[17768]_  & \new_[19791]_ ;
  assign \new_[16382]_  = ~\new_[16799]_ ;
  assign \new_[16383]_  = ~\new_[17214]_ ;
  assign \new_[16384]_  = ~\new_[16796]_ ;
  assign \new_[16385]_  = ~\new_[16775]_ ;
  assign \new_[16386]_  = ~\new_[16760]_ ;
  assign \new_[16387]_  = ~\new_[17760]_  & ~\new_[18008]_ ;
  assign \new_[16388]_  = ~\new_[16741]_ ;
  assign \new_[16389]_  = ~\new_[17936]_  | ~\new_[18945]_ ;
  assign \new_[16390]_  = ~\new_[18598]_  | ~\new_[18398]_ ;
  assign \new_[16391]_  = ~\new_[18014]_  & ~\new_[19044]_ ;
  assign \new_[16392]_  = \new_[17952]_  & \new_[20487]_ ;
  assign \new_[16393]_  = \new_[17497]_  & \new_[20241]_ ;
  assign \new_[16394]_  = ~\new_[16742]_ ;
  assign \new_[16395]_  = ~\new_[17852]_  | ~\new_[18187]_ ;
  assign \new_[16396]_  = ~\new_[18614]_  | ~\new_[18398]_ ;
  assign \new_[16397]_  = ~\new_[17421]_ ;
  assign \new_[16398]_  = ~\new_[17708]_  & ~\new_[21574]_ ;
  assign \new_[16399]_  = ~\new_[18250]_  | ~\new_[19184]_ ;
  assign \new_[16400]_  = ~\new_[19637]_  & ~\new_[17918]_ ;
  assign \new_[16401]_  = ~\new_[17206]_ ;
  assign \new_[16402]_  = ~\new_[17587]_  & ~\new_[18083]_ ;
  assign \new_[16403]_  = ~\new_[17458]_  & ~\new_[18784]_ ;
  assign \new_[16404]_  = ~\new_[17803]_  | ~\new_[21574]_ ;
  assign \new_[16405]_  = ~\new_[17031]_ ;
  assign \new_[16406]_  = ~\new_[16984]_ ;
  assign \new_[16407]_  = ~\new_[18695]_  | ~\new_[19088]_ ;
  assign \new_[16408]_  = ~\new_[17211]_ ;
  assign \new_[16409]_  = ~\new_[17257]_ ;
  assign \new_[16410]_  = ~\new_[17248]_ ;
  assign \new_[16411]_  = ~\new_[16809]_ ;
  assign \new_[16412]_  = ~\new_[17646]_ ;
  assign \new_[16413]_  = ~\new_[17875]_  | ~\new_[18680]_ ;
  assign \new_[16414]_  = ~\new_[18864]_  & ~\new_[19655]_ ;
  assign \new_[16415]_  = ~\new_[18686]_  | ~\new_[17638]_ ;
  assign \new_[16416]_  = ~\new_[17094]_ ;
  assign \new_[16417]_  = ~\new_[17590]_  & ~\new_[19019]_ ;
  assign \new_[16418]_  = ~\new_[17552]_  & ~\new_[17743]_ ;
  assign \new_[16419]_  = ~\new_[16952]_ ;
  assign \new_[16420]_  = ~\new_[18112]_  | ~\new_[17886]_ ;
  assign \new_[16421]_  = ~\new_[17218]_ ;
  assign \new_[16422]_  = ~\new_[16867]_ ;
  assign \new_[16423]_  = ~\new_[16861]_ ;
  assign \new_[16424]_  = ~\new_[17174]_ ;
  assign \new_[16425]_  = ~\new_[16835]_ ;
  assign \new_[16426]_  = ~\new_[16787]_ ;
  assign \new_[16427]_  = ~\new_[18310]_  | ~\new_[18965]_ ;
  assign \new_[16428]_  = ~\new_[17221]_ ;
  assign \new_[16429]_  = ~\new_[17527]_  | ~\new_[18766]_ ;
  assign \new_[16430]_  = ~\new_[16923]_ ;
  assign \new_[16431]_  = ~\new_[17748]_  | ~\new_[19555]_ ;
  assign \new_[16432]_  = ~\new_[17530]_  & ~\new_[21570]_ ;
  assign \new_[16433]_  = ~\new_[16757]_ ;
  assign \new_[16434]_  = ~\new_[16920]_ ;
  assign \new_[16435]_  = ~\new_[16731]_ ;
  assign \new_[16436]_  = \new_[18570]_  & \new_[18838]_ ;
  assign \new_[16437]_  = \new_[17580]_  & \new_[18337]_ ;
  assign \new_[16438]_  = ~\new_[16702]_ ;
  assign \new_[16439]_  = ~\new_[16896]_ ;
  assign \new_[16440]_  = \new_[17913]_  | \new_[17973]_ ;
  assign \new_[16441]_  = ~\new_[17231]_ ;
  assign \new_[16442]_  = ~\new_[16909]_ ;
  assign \new_[16443]_  = \new_[17928]_  & \new_[19674]_ ;
  assign \new_[16444]_  = \new_[17795]_  | \new_[19675]_ ;
  assign \new_[16445]_  = \new_[17537]_  & \new_[19156]_ ;
  assign \new_[16446]_  = \new_[17519]_  | \new_[17529]_ ;
  assign \new_[16447]_  = ~\new_[17366]_ ;
  assign \new_[16448]_  = ~\new_[17343]_ ;
  assign \new_[16449]_  = ~\new_[16894]_ ;
  assign \new_[16450]_  = ~\new_[18050]_  | ~\new_[19727]_ ;
  assign \new_[16451]_  = ~\new_[17226]_ ;
  assign \new_[16452]_  = ~\new_[17507]_  | ~\new_[19459]_ ;
  assign \new_[16453]_  = ~\new_[17283]_ ;
  assign \new_[16454]_  = ~\new_[17477]_  & ~\new_[19386]_ ;
  assign \new_[16455]_  = ~\new_[20237]_  | ~\new_[17659]_ ;
  assign \new_[16456]_  = ~\new_[17970]_  & ~\new_[19042]_ ;
  assign \new_[16457]_  = ~\new_[16768]_ ;
  assign \new_[16458]_  = ~\new_[17577]_  | ~\new_[21501]_ ;
  assign \new_[16459]_  = ~\new_[18788]_  | ~\new_[18173]_ ;
  assign \new_[16460]_  = ~\new_[16871]_ ;
  assign \new_[16461]_  = ~\new_[16869]_ ;
  assign \new_[16462]_  = ~\new_[17024]_ ;
  assign \new_[16463]_  = ~\new_[17762]_  | ~\new_[21496]_ ;
  assign \new_[16464]_  = ~\new_[16802]_ ;
  assign \new_[16465]_  = ~\new_[17914]_  & ~\new_[19213]_ ;
  assign \new_[16466]_  = ~\new_[17662]_  & ~\new_[21328]_ ;
  assign \new_[16467]_  = ~\new_[17948]_  | ~\new_[19389]_ ;
  assign \new_[16468]_  = \new_[17867]_  | \new_[19186]_ ;
  assign \new_[16469]_  = ~\new_[16943]_ ;
  assign \new_[16470]_  = ~\new_[17888]_  & ~\new_[19459]_ ;
  assign \new_[16471]_  = ~\new_[17617]_  & ~\new_[20865]_ ;
  assign \new_[16472]_  = \new_[17654]_  & \new_[19603]_ ;
  assign \new_[16473]_  = ~\new_[17836]_  & ~\new_[18968]_ ;
  assign \new_[16474]_  = ~\new_[16772]_ ;
  assign \new_[16475]_  = ~\new_[16817]_ ;
  assign \new_[16476]_  = ~\new_[16806]_ ;
  assign \new_[16477]_  = ~\new_[17634]_  & ~\new_[19048]_ ;
  assign \new_[16478]_  = ~\new_[17930]_  | ~\new_[18496]_ ;
  assign \new_[16479]_  = ~\new_[17965]_  | ~\new_[17962]_ ;
  assign \new_[16480]_  = ~\new_[16837]_ ;
  assign \new_[16481]_  = ~\new_[17790]_  | ~\new_[18587]_ ;
  assign \new_[16482]_  = ~\new_[17414]_ ;
  assign \new_[16483]_  = ~\new_[17238]_ ;
  assign \new_[16484]_  = ~\new_[17102]_ ;
  assign \new_[16485]_  = ~\new_[17879]_  | ~\new_[19386]_ ;
  assign \new_[16486]_  = ~\new_[17239]_ ;
  assign \new_[16487]_  = ~\new_[18920]_  | ~\new_[18284]_ ;
  assign \new_[16488]_  = ~\new_[17240]_ ;
  assign \new_[16489]_  = ~\new_[16815]_ ;
  assign \new_[16490]_  = ~\new_[17542]_  | ~\new_[18945]_ ;
  assign \new_[16491]_  = ~\new_[17377]_ ;
  assign \new_[16492]_  = \new_[17885]_  & \new_[21685]_ ;
  assign \new_[16493]_  = ~\new_[16721]_ ;
  assign \new_[16494]_  = ~\new_[18015]_  | ~\new_[17839]_ ;
  assign \new_[16495]_  = \new_[18032]_  | \new_[17485]_ ;
  assign \new_[16496]_  = ~\new_[19084]_  & ~\new_[17955]_ ;
  assign \new_[16497]_  = ~\new_[17609]_  | ~\new_[19144]_ ;
  assign \new_[16498]_  = ~\new_[17520]_  | ~\new_[19176]_ ;
  assign \new_[16499]_  = ~\new_[18788]_  | ~\new_[19238]_ ;
  assign \new_[16500]_  = ~\new_[16789]_ ;
  assign \new_[16501]_  = ~\new_[16780]_ ;
  assign \new_[16502]_  = ~\new_[17462]_  & ~\new_[19741]_ ;
  assign \new_[16503]_  = ~\new_[17052]_ ;
  assign \new_[16504]_  = ~\new_[17009]_ ;
  assign \new_[16505]_  = ~\new_[17550]_  | ~\new_[17985]_ ;
  assign \new_[16506]_  = ~\new_[16773]_ ;
  assign \new_[16507]_  = ~\new_[18527]_  | ~\new_[19526]_ ;
  assign \new_[16508]_  = ~\new_[18806]_  | ~\new_[19675]_ ;
  assign \new_[16509]_  = ~\new_[17250]_ ;
  assign \new_[16510]_  = \new_[17980]_  | \new_[17743]_ ;
  assign \new_[16511]_  = \\u0_r0_rcnt_reg[1] ;
  assign \new_[16512]_  = ~\new_[17260]_ ;
  assign \new_[16513]_  = ~\new_[16838]_ ;
  assign \new_[16514]_  = ~\new_[16714]_ ;
  assign \new_[16515]_  = ~\new_[16718]_ ;
  assign \new_[16516]_  = ~\new_[17639]_  & ~\new_[19353]_ ;
  assign \new_[16517]_  = ~\new_[16914]_ ;
  assign \new_[16518]_  = ~\new_[17567]_  | ~\new_[21689]_ ;
  assign \new_[16519]_  = \new_[17740]_  & \new_[19758]_ ;
  assign \new_[16520]_  = \new_[17949]_  | \new_[17529]_ ;
  assign \new_[16521]_  = ~\new_[18708]_  | ~\new_[18103]_ ;
  assign \new_[16522]_  = ~\new_[17824]_  & ~\new_[19219]_ ;
  assign \new_[16523]_  = ~\new_[17671]_  | ~\new_[21259]_ ;
  assign \new_[16524]_  = ~\new_[17695]_  & ~\new_[19548]_ ;
  assign \new_[16525]_  = ~\new_[17873]_  | ~\new_[18543]_ ;
  assign \new_[16526]_  = ~\new_[17154]_ ;
  assign \new_[16527]_  = ~\new_[17159]_ ;
  assign \new_[16528]_  = ~\new_[17344]_ ;
  assign \new_[16529]_  = ~\new_[17597]_  | ~\new_[19676]_ ;
  assign \new_[16530]_  = ~\new_[16713]_ ;
  assign \new_[16531]_  = ~\new_[17424]_ ;
  assign \new_[16532]_  = ~\new_[19821]_  | ~\new_[19224]_ ;
  assign \new_[16533]_  = ~\new_[17696]_  & ~\new_[17534]_ ;
  assign \new_[16534]_  = ~\new_[17740]_  | ~\new_[19026]_ ;
  assign \new_[16535]_  = \new_[17377]_ ;
  assign \new_[16536]_  = ~\new_[17408]_ ;
  assign \new_[16537]_  = \new_[17673]_  | \new_[19642]_ ;
  assign \new_[16538]_  = ~\new_[17665]_  | ~\new_[17950]_ ;
  assign \new_[16539]_  = ~\new_[19782]_  & ~\new_[17943]_ ;
  assign \new_[16540]_  = ~\new_[19248]_  | ~\new_[18864]_ ;
  assign \new_[16541]_  = \new_[21653]_  & \new_[18355]_ ;
  assign \new_[16542]_  = ~\new_[20747]_ ;
  assign \new_[16543]_  = ~\new_[17608]_  & ~\new_[17979]_ ;
  assign \new_[16544]_  = \new_[17461]_  & \new_[17816]_ ;
  assign \new_[16545]_  = ~\new_[18613]_  | ~\new_[18721]_ ;
  assign \new_[16546]_  = ~\new_[17682]_  | ~\new_[17967]_ ;
  assign \new_[16547]_  = ~\new_[18369]_  | ~\new_[17471]_ ;
  assign \new_[16548]_  = ~\new_[17831]_  & ~\new_[19476]_ ;
  assign \new_[16549]_  = ~\new_[18250]_  | ~\new_[17748]_ ;
  assign \new_[16550]_  = ~\new_[17143]_ ;
  assign \new_[16551]_  = ~\new_[17261]_ ;
  assign \new_[16552]_  = ~\new_[17948]_  | ~\new_[17709]_ ;
  assign \new_[16553]_  = ~\new_[17282]_ ;
  assign \new_[16554]_  = ~\new_[17611]_  | ~\new_[19275]_ ;
  assign \new_[16555]_  = ~\new_[17298]_ ;
  assign \new_[16556]_  = \new_[17772]_  | \new_[19742]_ ;
  assign \new_[16557]_  = ~\new_[17982]_  | ~\new_[20749]_ ;
  assign \new_[16558]_  = ~\new_[17207]_ ;
  assign \new_[16559]_  = ~\new_[16803]_ ;
  assign \new_[16560]_  = ~\new_[17763]_  & ~\new_[19386]_ ;
  assign \new_[16561]_  = \new_[17799]_  | \new_[21328]_ ;
  assign \new_[16562]_  = ~\new_[17227]_ ;
  assign \new_[16563]_  = ~\new_[17480]_  & ~\new_[19785]_ ;
  assign \new_[16564]_  = ~\new_[17279]_ ;
  assign \new_[16565]_  = ~\new_[17326]_ ;
  assign \new_[16566]_  = ~\new_[17951]_  | ~\new_[19053]_ ;
  assign \new_[16567]_  = ~\new_[17520]_  & ~\new_[19176]_ ;
  assign \new_[16568]_  = ~\new_[16712]_ ;
  assign \new_[16569]_  = ~\new_[17679]_  & ~\new_[19128]_ ;
  assign \new_[16570]_  = ~\new_[17306]_ ;
  assign \new_[16571]_  = ~\new_[17209]_ ;
  assign \new_[16572]_  = ~\new_[17258]_ ;
  assign \new_[16573]_  = ~\new_[17684]_  | ~\new_[18615]_ ;
  assign \new_[16574]_  = ~\new_[17498]_  | ~\new_[18784]_ ;
  assign \new_[16575]_  = ~\new_[21604]_ ;
  assign \new_[16576]_  = ~\new_[17783]_  | ~\new_[21693]_ ;
  assign \new_[16577]_  = ~\new_[17418]_ ;
  assign \new_[16578]_  = ~\new_[19386]_  | ~\new_[17476]_ ;
  assign \new_[16579]_  = ~\new_[17716]_  & ~\new_[20241]_ ;
  assign \new_[16580]_  = ~\new_[19459]_  & ~\new_[17961]_ ;
  assign \new_[16581]_  = \new_[19684]_  ^ \new_[18519]_ ;
  assign \new_[16582]_  = ~\new_[17317]_ ;
  assign \new_[16583]_  = ~\new_[17606]_  | ~\new_[19788]_ ;
  assign \new_[16584]_  = ~\new_[16857]_ ;
  assign \new_[16585]_  = \new_[18010]_  & \new_[19123]_ ;
  assign \new_[16586]_  = ~\new_[17978]_  | ~\new_[18056]_ ;
  assign \new_[16587]_  = ~\new_[17885]_  | ~\new_[19285]_ ;
  assign \new_[16588]_  = ~\new_[17564]_  & ~\new_[19410]_ ;
  assign \new_[16589]_  = ~\new_[17806]_  & ~\new_[19555]_ ;
  assign \new_[16590]_  = ~\new_[17321]_ ;
  assign \new_[16591]_  = ~\new_[17701]_  | ~\new_[18968]_ ;
  assign \new_[16592]_  = ~\new_[17528]_  | ~\new_[19082]_ ;
  assign \new_[16593]_  = \new_[17792]_  & \new_[18676]_ ;
  assign \new_[16594]_  = ~\new_[17329]_ ;
  assign \new_[16595]_  = ~\new_[16850]_ ;
  assign \new_[16596]_  = ~\new_[17295]_ ;
  assign \new_[16597]_  = ~\new_[17341]_ ;
  assign \new_[16598]_  = ~\new_[16747]_ ;
  assign \new_[16599]_  = ~\new_[18009]_  & ~\new_[19409]_ ;
  assign \new_[16600]_  = ~\new_[17044]_ ;
  assign \new_[16601]_  = ~\new_[16970]_ ;
  assign \new_[16602]_  = ~\new_[16993]_ ;
  assign \new_[16603]_  = ~\new_[17947]_  & ~\new_[17700]_ ;
  assign \new_[16604]_  = ~\new_[16977]_ ;
  assign \new_[16605]_  = \new_[19048]_  & \new_[18660]_ ;
  assign \new_[16606]_  = ~\new_[20036]_ ;
  assign \new_[16607]_  = ~\new_[17886]_  | ~\new_[18651]_ ;
  assign \new_[16608]_  = ~\new_[17431]_ ;
  assign \new_[16609]_  = ~\new_[18019]_  & ~\new_[21569]_ ;
  assign \new_[16610]_  = ~\new_[17270]_ ;
  assign \new_[16611]_  = \new_[18575]_  & \new_[17459]_ ;
  assign \new_[16612]_  = ~\new_[17195]_ ;
  assign \new_[16613]_  = \new_[18222]_  & \new_[18806]_ ;
  assign \new_[16614]_  = ~\new_[17635]_  & ~\new_[19741]_ ;
  assign \new_[16615]_  = \new_[18833]_  & \new_[19550]_ ;
  assign \new_[16616]_  = ~\new_[17514]_  & ~\new_[19104]_ ;
  assign \new_[16617]_  = ~\new_[16901]_ ;
  assign \new_[16618]_  = \new_[20749]_  & \new_[17496]_ ;
  assign \new_[16619]_  = ~\new_[16793]_ ;
  assign \new_[16620]_  = \new_[17798]_  | \new_[19444]_ ;
  assign \new_[16621]_  = \new_[17643]_  & \new_[19535]_ ;
  assign \new_[16622]_  = \new_[16933]_ ;
  assign \new_[16623]_  = \new_[16711]_ ;
  assign \new_[16624]_  = ~\new_[17376]_ ;
  assign \new_[16625]_  = ~\new_[16882]_ ;
  assign \new_[16626]_  = ~\new_[17709]_  | ~\new_[19444]_ ;
  assign \new_[16627]_  = ~\new_[17417]_ ;
  assign \new_[16628]_  = ~\new_[19553]_  & ~\new_[18906]_ ;
  assign \new_[16629]_  = ~\new_[17415]_ ;
  assign \new_[16630]_  = ~\new_[16709]_ ;
  assign \new_[16631]_  = ~\new_[17012]_ ;
  assign \new_[16632]_  = \new_[19028]_  & \new_[21422]_ ;
  assign \new_[16633]_  = ~\new_[17760]_  & ~\new_[19386]_ ;
  assign \new_[16634]_  = ~\new_[16716]_ ;
  assign \new_[16635]_  = ~\new_[17396]_ ;
  assign \new_[16636]_  = ~\new_[16979]_ ;
  assign \new_[16637]_  = ~\new_[18005]_  & ~\new_[18810]_ ;
  assign \new_[16638]_  = ~\new_[17242]_ ;
  assign \new_[16639]_  = ~\new_[17916]_  | ~\new_[19091]_ ;
  assign \new_[16640]_  = ~\new_[17961]_  & ~\new_[18325]_ ;
  assign \new_[16641]_  = ~\new_[17956]_  | ~\new_[19444]_ ;
  assign \new_[16642]_  = ~\new_[16781]_ ;
  assign \new_[16643]_  = ~\new_[16991]_ ;
  assign \new_[16644]_  = ~\new_[18888]_  | ~\new_[17607]_ ;
  assign \new_[16645]_  = ~\new_[17183]_ ;
  assign \new_[16646]_  = ~\new_[16997]_ ;
  assign \new_[16647]_  = \new_[18980]_  & \new_[19555]_ ;
  assign \new_[16648]_  = ~\new_[17384]_ ;
  assign \new_[16649]_  = ~\new_[17476]_  | ~\new_[18008]_ ;
  assign \new_[16650]_  = ~\new_[17215]_ ;
  assign \new_[16651]_  = ~\new_[16911]_ ;
  assign \new_[16652]_  = ~\new_[17449]_ ;
  assign \new_[16653]_  = ~\new_[17205]_ ;
  assign \new_[16654]_  = \new_[17976]_  | \new_[19100]_ ;
  assign \new_[16655]_  = ~\new_[17886]_  | ~\new_[19147]_ ;
  assign \new_[16656]_  = ~\new_[17182]_ ;
  assign \new_[16657]_  = ~\new_[18023]_  | ~\new_[17709]_ ;
  assign \new_[16658]_  = ~\new_[17484]_  & ~\new_[19550]_ ;
  assign \new_[16659]_  = ~\new_[19719]_  & ~\new_[17679]_ ;
  assign \new_[16660]_  = ~\new_[16702]_ ;
  assign \new_[16661]_  = ~\new_[17435]_ ;
  assign \new_[16662]_  = ~\new_[17204]_ ;
  assign \new_[16663]_  = ~\new_[17942]_  | ~\new_[18173]_ ;
  assign \new_[16664]_  = ~\new_[17433]_ ;
  assign \new_[16665]_  = ~\new_[17556]_  | ~\new_[19096]_ ;
  assign \new_[16666]_  = ~\new_[17181]_ ;
  assign \new_[16667]_  = n3213 & \new_[17156]_ ;
  assign \new_[16668]_  = ~\new_[17497]_  | ~\new_[18903]_ ;
  assign \new_[16669]_  = ~\new_[18192]_  & ~\new_[17914]_ ;
  assign \new_[16670]_  = ~\new_[17452]_ ;
  assign \new_[16671]_  = ~\new_[17854]_  | ~\new_[21693]_ ;
  assign \new_[16672]_  = ~\new_[17744]_  & ~\new_[18987]_ ;
  assign \new_[16673]_  = ~\new_[17147]_ ;
  assign \new_[16674]_  = ~\new_[17633]_  & ~\new_[19353]_ ;
  assign \new_[16675]_  = ~\new_[17443]_ ;
  assign \new_[16676]_  = ~\new_[17690]_ ;
  assign \new_[16677]_  = ~\new_[17821]_  | ~\new_[19214]_ ;
  assign \new_[16678]_  = ~\new_[17705]_  | ~\new_[14951]_ ;
  assign \new_[16679]_  = ~\new_[17454]_ ;
  assign \new_[16680]_  = ~\new_[17787]_  & ~\new_[19547]_ ;
  assign \new_[16681]_  = ~\new_[17001]_ ;
  assign \new_[16682]_  = ~\new_[19526]_ ;
  assign \new_[16683]_  = ~\new_[18379]_  | ~\new_[19225]_ ;
  assign \new_[16684]_  = \\text_in_r_reg[125] ;
  assign n2973 = \new_[14793]_  ? \new_[19283]_  : \text_in[96] ;
  assign \new_[16686]_  = ~\new_[18100]_  | ~\new_[19788]_ ;
  assign \new_[16687]_  = ~\new_[18069]_  | ~\new_[19123]_ ;
  assign n3048 = \new_[14944]_  ? \new_[19283]_  : \text_in[66] ;
  assign \new_[16689]_  = ~\new_[18026]_  & ~\new_[19082]_ ;
  assign \new_[16690]_  = ~\new_[17541]_ ;
  assign \new_[16691]_  = ~\new_[18131]_  | ~\new_[21517]_ ;
  assign \new_[16692]_  = \\text_in_r_reg[2] ;
  assign \new_[16693]_  = ~\new_[18405]_  | ~\new_[19000]_ ;
  assign n2793 = \new_[14702]_  ? \new_[19497]_  : \text_in[47] ;
  assign \new_[16695]_  = ~\new_[17572]_ ;
  assign \new_[16696]_  = ~\new_[17465]_ ;
  assign n2833 = \new_[14753]_  ? \new_[19497]_  : \text_in[54] ;
  assign \new_[16698]_  = ~\new_[18217]_  | ~\new_[21659]_ ;
  assign \new_[16699]_  = ~\new_[18177]_  | ~\new_[19464]_ ;
  assign \new_[16700]_  = ~\new_[17922]_ ;
  assign \new_[16701]_  = \\text_in_r_reg[44] ;
  assign \new_[16702]_  = ~\new_[19000]_  & ~\new_[18200]_ ;
  assign \new_[16703]_  = ~\new_[17853]_ ;
  assign \new_[16704]_  = ~\new_[18149]_  | ~\new_[19746]_ ;
  assign \new_[16705]_  = ~\new_[18555]_  | ~\new_[19312]_ ;
  assign \new_[16706]_  = \new_[18347]_  | \new_[19335]_ ;
  assign n2943 = \new_[14779]_  ? ld : \text_in[103] ;
  assign \new_[16708]_  = ~\new_[17864]_ ;
  assign \new_[16709]_  = ~\new_[17953]_ ;
  assign \new_[16710]_  = ~\new_[17473]_ ;
  assign \new_[16711]_  = ~\new_[17477]_ ;
  assign \new_[16712]_  = \new_[18349]_  | \new_[19676]_ ;
  assign \new_[16713]_  = ~\new_[18381]_  | ~\new_[21521]_ ;
  assign \new_[16714]_  = \new_[18301]_  | \new_[19190]_ ;
  assign \new_[16715]_  = \\text_in_r_reg[72] ;
  assign \new_[16716]_  = ~\new_[17649]_ ;
  assign n2858 = \new_[14760]_  ? \new_[19497]_  : \text_in[11] ;
  assign \new_[16718]_  = ~\new_[17995]_ ;
  assign \new_[16719]_  = ~\new_[18350]_  | ~\new_[19617]_ ;
  assign \new_[16720]_  = ~\new_[17464]_ ;
  assign \new_[16721]_  = ~\new_[18331]_  & ~\new_[19100]_ ;
  assign \new_[16722]_  = ~\new_[17711]_ ;
  assign \new_[16723]_  = \\text_in_r_reg[101] ;
  assign \new_[16724]_  = ~\new_[19045]_  | ~\new_[19033]_ ;
  assign n2958 = \new_[14782]_  ? \new_[19283]_  : \text_in[3] ;
  assign n2998 = \new_[14893]_  ? \new_[19283]_  : \text_in[28] ;
  assign \new_[16727]_  = ~\new_[17493]_ ;
  assign \new_[16728]_  = ~\new_[19210]_  & ~\new_[18065]_ ;
  assign \new_[16729]_  = ~\new_[17479]_ ;
  assign \new_[16730]_  = ~\new_[17959]_ ;
  assign \new_[16731]_  = ~\new_[18102]_  & ~\new_[18424]_ ;
  assign \new_[16732]_  = \new_[17430]_  ^ \new_[2291]_ ;
  assign \new_[16733]_  = ~\new_[18142]_  | ~\new_[21306]_ ;
  assign \new_[16734]_  = ~\new_[18451]_  | ~\new_[21490]_ ;
  assign \new_[16735]_  = ~\new_[18524]_  & ~\new_[19386]_ ;
  assign n2868 = \new_[14762]_  ? \new_[19497]_  : \text_in[24] ;
  assign \new_[16737]_  = ~\new_[18266]_  | ~\new_[19685]_ ;
  assign \new_[16738]_  = ~\new_[18150]_  | ~\new_[19603]_ ;
  assign \new_[16739]_  = \new_[19098]_  & \new_[18253]_ ;
  assign \new_[16740]_  = ~\new_[18565]_ ;
  assign \new_[16741]_  = ~\new_[17693]_ ;
  assign \new_[16742]_  = ~\new_[17582]_ ;
  assign \new_[16743]_  = \\text_in_r_reg[106] ;
  assign \new_[16744]_  = ~\new_[17491]_ ;
  assign \new_[16745]_  = \new_[17774]_  | \new_[19676]_ ;
  assign \new_[16746]_  = ~\new_[18526]_  | ~\new_[18963]_ ;
  assign \new_[16747]_  = \new_[17739]_ ;
  assign \new_[16748]_  = ~\new_[18549]_  | ~\new_[21259]_ ;
  assign \new_[16749]_  = ~\new_[18901]_  & ~\new_[18045]_ ;
  assign \new_[16750]_  = ~\new_[20293]_ ;
  assign \new_[16751]_  = ~\new_[18238]_  & ~\new_[19655]_ ;
  assign \new_[16752]_  = \\text_in_r_reg[4] ;
  assign \new_[16753]_  = \new_[18024]_  & \new_[19697]_ ;
  assign \new_[16754]_  = \\text_in_r_reg[43] ;
  assign \new_[16755]_  = ~\new_[18975]_  | ~\new_[21495]_ ;
  assign \new_[16756]_  = ~\new_[18404]_  | ~\new_[21578]_ ;
  assign \new_[16757]_  = ~\new_[18433]_  | ~\new_[19788]_ ;
  assign \new_[16758]_  = \\text_in_r_reg[112] ;
  assign \new_[16759]_  = ~\new_[17499]_ ;
  assign \new_[16760]_  = ~\new_[18210]_  | ~\new_[21574]_ ;
  assign n2773 = \new_[14697]_  ? \new_[19283]_  : \text_in[111] ;
  assign \new_[16762]_  = ~\new_[18013]_ ;
  assign \new_[16763]_  = ~\new_[17495]_ ;
  assign \new_[16764]_  = ~\new_[19268]_  & ~\new_[18186]_ ;
  assign \new_[16765]_  = ~\new_[17752]_ ;
  assign \new_[16766]_  = ~\new_[18229]_  | ~\new_[21489]_ ;
  assign \new_[16767]_  = ~\new_[18248]_  | ~\new_[19463]_ ;
  assign \new_[16768]_  = ~\new_[17872]_ ;
  assign \new_[16769]_  = ~\new_[17506]_ ;
  assign \new_[16770]_  = ~\new_[17501]_ ;
  assign \new_[16771]_  = ~\new_[17831]_ ;
  assign \new_[16772]_  = ~\new_[18425]_  | ~\new_[19104]_ ;
  assign \new_[16773]_  = ~\new_[17788]_ ;
  assign n2788 = \new_[14701]_  ? \new_[19497]_  : \text_in[67] ;
  assign \new_[16775]_  = ~\new_[18353]_  | ~\new_[19438]_ ;
  assign \new_[16776]_  = ~\new_[17677]_ ;
  assign \new_[16777]_  = \\text_in_r_reg[93] ;
  assign \new_[16778]_  = ~\new_[18128]_  & ~\new_[19066]_ ;
  assign n3023 = \new_[14912]_  ? \new_[19283]_  : \text_in[90] ;
  assign \new_[16780]_  = ~\new_[17494]_ ;
  assign \new_[16781]_  = ~\new_[17510]_ ;
  assign \new_[16782]_  = ~\new_[17512]_ ;
  assign \new_[16783]_  = ~\new_[18345]_  | ~\new_[19801]_ ;
  assign \new_[16784]_  = ~\new_[17808]_ ;
  assign \new_[16785]_  = ~\new_[17666]_ ;
  assign \new_[16786]_  = ~\new_[17545]_ ;
  assign \new_[16787]_  = ~\new_[18094]_  & ~\new_[18963]_ ;
  assign \new_[16788]_  = ~\new_[17483]_ ;
  assign \new_[16789]_  = ~\new_[18553]_  | ~\new_[19026]_ ;
  assign \new_[16790]_  = ~\new_[18362]_  & ~\new_[18740]_ ;
  assign \new_[16791]_  = ~\new_[18433]_  | ~\new_[19647]_ ;
  assign \new_[16792]_  = ~\new_[17923]_ ;
  assign \new_[16793]_  = ~\new_[19139]_  | ~\new_[20239]_ ;
  assign \new_[16794]_  = ~\new_[17670]_ ;
  assign \new_[16795]_  = \\text_in_r_reg[73] ;
  assign \new_[16796]_  = ~\new_[18375]_  | ~\new_[19785]_ ;
  assign \new_[16797]_  = ~\new_[17521]_ ;
  assign \new_[16798]_  = ~\new_[17755]_ ;
  assign \new_[16799]_  = ~\new_[17706]_ ;
  assign \new_[16800]_  = ~\new_[17679]_ ;
  assign \new_[16801]_  = \\text_in_r_reg[50] ;
  assign \new_[16802]_  = ~\new_[18336]_  | ~\new_[20495]_ ;
  assign \new_[16803]_  = ~\new_[18145]_  & ~\new_[19026]_ ;
  assign \new_[16804]_  = ~\new_[18160]_  | ~\new_[18802]_ ;
  assign \new_[16805]_  = ~\new_[18541]_  | ~\new_[19379]_ ;
  assign \new_[16806]_  = ~\new_[18038]_  & ~\new_[19444]_ ;
  assign \new_[16807]_  = \new_[18349]_  | \new_[19156]_ ;
  assign \new_[16808]_  = ~\new_[17540]_ ;
  assign \new_[16809]_  = ~\new_[18345]_  | ~\new_[19200]_ ;
  assign \new_[16810]_  = ~\new_[17708]_ ;
  assign \new_[16811]_  = \new_[19088]_  & \new_[19271]_ ;
  assign \new_[16812]_  = \new_[14941]_  ^ \new_[19325]_ ;
  assign \new_[16813]_  = ~\new_[19147]_  | ~\new_[18111]_ ;
  assign \new_[16814]_  = ~\new_[20235]_  | ~\new_[21522]_ ;
  assign \new_[16815]_  = ~\new_[18067]_  | ~\new_[19379]_ ;
  assign \new_[16816]_  = ~\new_[18034]_  | ~\new_[18947]_ ;
  assign \new_[16817]_  = ~\new_[18146]_  | ~\new_[19132]_ ;
  assign \new_[16818]_  = \new_[21115]_  & \new_[19748]_ ;
  assign n2863 = \new_[14761]_  ? \new_[19414]_  : \text_in[123] ;
  assign \new_[16820]_  = ~\new_[17764]_ ;
  assign \new_[16821]_  = ~\new_[18056]_  | ~\new_[19568]_ ;
  assign n2978 = \new_[14799]_  ? \new_[19283]_  : \text_in[70] ;
  assign \new_[16823]_  = ~\new_[18475]_  & ~\new_[19459]_ ;
  assign \new_[16824]_  = ~\new_[18415]_  | ~\new_[21396]_ ;
  assign \new_[16825]_  = ~\new_[18340]_  & ~\new_[18489]_ ;
  assign \new_[16826]_  = \\text_in_r_reg[100] ;
  assign \new_[16827]_  = ~\new_[17552]_ ;
  assign \new_[16828]_  = ~\new_[17575]_ ;
  assign \new_[16829]_  = ~\new_[17575]_ ;
  assign \new_[16830]_  = ~n3213;
  assign \new_[16831]_  = \new_[19655]_  | \new_[18390]_ ;
  assign \new_[16832]_  = ~\new_[17554]_ ;
  assign \new_[16833]_  = ~\new_[17462]_ ;
  assign \new_[16834]_  = \new_[19267]_  | \new_[21685]_ ;
  assign \new_[16835]_  = ~\new_[18913]_  & ~\new_[18088]_ ;
  assign \new_[16836]_  = \new_[18794]_  | \new_[21658]_ ;
  assign \new_[16837]_  = ~\new_[20932]_  | ~\new_[19353]_ ;
  assign \new_[16838]_  = ~\new_[17558]_ ;
  assign \new_[16839]_  = ~\new_[18287]_  & ~\new_[19379]_ ;
  assign \new_[16840]_  = ~\new_[18714]_ ;
  assign n3058 = \new_[14956]_  ? ld : \text_in[53] ;
  assign \new_[16842]_  = ~\new_[18141]_  & ~\new_[18945]_ ;
  assign \new_[16843]_  = ~\new_[17563]_ ;
  assign \new_[16844]_  = \new_[19044]_  | \new_[18139]_ ;
  assign \new_[16845]_  = ~\new_[17617]_ ;
  assign \new_[16846]_  = ~\new_[17502]_ ;
  assign \new_[16847]_  = ~\new_[18262]_  | ~\new_[18363]_ ;
  assign \new_[16848]_  = \\text_in_r_reg[114] ;
  assign \new_[16849]_  = ~\new_[18445]_  & ~\new_[19097]_ ;
  assign \new_[16850]_  = ~\new_[21254]_  | ~\new_[19220]_ ;
  assign \new_[16851]_  = ~\new_[17884]_ ;
  assign n3193 = \new_[15853]_  ? \new_[19414]_  : \text_in[32] ;
  assign \new_[16853]_  = ~\new_[18527]_  | ~\new_[14690]_ ;
  assign \new_[16854]_  = \\text_in_r_reg[25] ;
  assign \new_[16855]_  = ~\new_[18263]_  | ~\new_[19092]_ ;
  assign n3108 = \new_[15470]_  ? \new_[19283]_  : \text_in[79] ;
  assign \new_[16857]_  = ~\new_[18376]_  | ~\new_[19146]_ ;
  assign \new_[16858]_  = ~\new_[18146]_  | ~\new_[19225]_ ;
  assign \new_[16859]_  = ~\new_[18098]_  | ~\new_[19342]_ ;
  assign \new_[16860]_  = \new_[16715]_  ^ \new_[1671]_ ;
  assign \new_[16861]_  = ~\new_[18329]_  | ~\new_[19395]_ ;
  assign \new_[16862]_  = \new_[19366]_  & \new_[19803]_ ;
  assign \new_[16863]_  = \new_[18472]_  | \new_[19642]_ ;
  assign \new_[16864]_  = \new_[20749]_  & \new_[18480]_ ;
  assign \new_[16865]_  = ~\new_[18163]_  | ~\new_[21524]_ ;
  assign \new_[16866]_  = ~\new_[18396]_ ;
  assign \new_[16867]_  = ~\new_[18059]_  & ~\new_[19676]_ ;
  assign n3008 = \new_[14902]_  ? \new_[19497]_  : \text_in[1] ;
  assign \new_[16869]_  = ~\new_[18206]_  | ~\new_[19192]_ ;
  assign \new_[16870]_  = ~\new_[17834]_ ;
  assign \new_[16871]_  = ~\new_[17718]_ ;
  assign \new_[16872]_  = ~\new_[17958]_ ;
  assign \new_[16873]_  = ~\new_[17576]_ ;
  assign \new_[16874]_  = ~\new_[17632]_ ;
  assign \new_[16875]_  = ~\new_[19079]_  & ~\new_[19638]_ ;
  assign \new_[16876]_  = ~\new_[19123]_  & ~\new_[19717]_ ;
  assign \new_[16877]_  = ~\new_[17747]_ ;
  assign \new_[16878]_  = ~\new_[19576]_  | ~\new_[19077]_  | ~\new_[19495]_  | ~\new_[12134]_ ;
  assign \new_[16879]_  = ~\new_[20701]_ ;
  assign \new_[16880]_  = ~\new_[17595]_ ;
  assign \new_[16881]_  = ~\new_[19097]_  | ~\new_[19159]_ ;
  assign \new_[16882]_  = ~\new_[17606]_ ;
  assign \new_[16883]_  = ~\new_[17750]_ ;
  assign \new_[16884]_  = ~\new_[17602]_ ;
  assign \new_[16885]_  = ~\new_[21533]_  | ~\new_[18893]_ ;
  assign \new_[16886]_  = ~\new_[19079]_  & ~\new_[973]_ ;
  assign \new_[16887]_  = ~\new_[17680]_ ;
  assign \new_[16888]_  = ~\new_[17562]_ ;
  assign \new_[16889]_  = \new_[19215]_  | \new_[19257]_ ;
  assign \new_[16890]_  = ~\new_[17617]_ ;
  assign \new_[16891]_  = ~\new_[17694]_ ;
  assign \new_[16892]_  = \\text_in_r_reg[57] ;
  assign \new_[16893]_  = ~\new_[18148]_  | ~\new_[19210]_ ;
  assign \new_[16894]_  = ~\new_[18520]_  & ~\new_[19597]_ ;
  assign n2853 = \new_[14759]_  ? \new_[19283]_  : \text_in[108] ;
  assign \new_[16896]_  = ~\new_[19689]_  | ~\new_[18317]_ ;
  assign \new_[16897]_  = ~\new_[17610]_ ;
  assign \new_[16898]_  = ~\new_[17678]_ ;
  assign \new_[16899]_  = ~\new_[21306]_  | ~\new_[18055]_ ;
  assign \new_[16900]_  = ~\new_[17605]_ ;
  assign \new_[16901]_  = ~\new_[17731]_ ;
  assign \new_[16902]_  = ~\new_[17661]_ ;
  assign \new_[16903]_  = ~\new_[18476]_  & ~\new_[19535]_ ;
  assign \new_[16904]_  = \new_[18461]_  & \new_[18995]_ ;
  assign \new_[16905]_  = ~\new_[17619]_ ;
  assign \new_[16906]_  = ~\new_[17822]_ ;
  assign \new_[16907]_  = ~\new_[17659]_ ;
  assign \new_[16908]_  = ~\new_[17695]_ ;
  assign \new_[16909]_  = ~\new_[18492]_  | ~\new_[21572]_ ;
  assign \new_[16910]_  = ~\new_[17611]_ ;
  assign \new_[16911]_  = ~\new_[18161]_  | ~\new_[19685]_ ;
  assign \new_[16912]_  = ~\new_[18018]_ ;
  assign \new_[16913]_  = ~\new_[17775]_ ;
  assign \new_[16914]_  = \new_[18499]_  | \new_[19675]_ ;
  assign \new_[16915]_  = ~\new_[18294]_  | ~\new_[21489]_ ;
  assign \new_[16916]_  = ~\new_[17651]_ ;
  assign n3083 = \new_[15068]_  ? \new_[19283]_  : \text_in[34] ;
  assign \new_[16918]_  = \\text_in_r_reg[95] ;
  assign \new_[16919]_  = ~\new_[17577]_ ;
  assign \new_[16920]_  = ~\new_[18119]_  | ~\new_[18640]_ ;
  assign \new_[16921]_  = ~\new_[18428]_  & ~\new_[19750]_ ;
  assign \new_[16922]_  = ~\new_[19228]_  | ~\new_[19250]_ ;
  assign \new_[16923]_  = ~\new_[18170]_  | ~\new_[19213]_ ;
  assign \new_[16924]_  = \new_[18182]_  | \new_[18779]_ ;
  assign \new_[16925]_  = ~\new_[17600]_ ;
  assign \new_[16926]_  = \\text_in_r_reg[124] ;
  assign \new_[16927]_  = ~\new_[17701]_ ;
  assign \new_[16928]_  = ~\new_[18273]_  & ~\new_[21572]_ ;
  assign \new_[16929]_  = ~\new_[17639]_ ;
  assign \new_[16930]_  = ~\new_[17631]_ ;
  assign \new_[16931]_  = ~\new_[19535]_  & ~\new_[19249]_ ;
  assign \new_[16932]_  = \new_[18025]_  & \new_[19550]_ ;
  assign \new_[16933]_  = ~\new_[17633]_ ;
  assign \new_[16934]_  = ~\new_[17527]_ ;
  assign \new_[16935]_  = ~\new_[17733]_ ;
  assign n3073 = \new_[15059]_  ? \new_[19283]_  : \text_in[97] ;
  assign \new_[16937]_  = ~\new_[18455]_  | ~\new_[19335]_ ;
  assign n2983 = \new_[14814]_  ? \new_[19414]_  : \text_in[51] ;
  assign \new_[16939]_  = ~\new_[20725]_ ;
  assign \new_[16940]_  = ~\new_[17990]_ ;
  assign \new_[16941]_  = ~\new_[18986]_  | ~\new_[19734]_ ;
  assign \new_[16942]_  = ~\new_[17998]_ ;
  assign \new_[16943]_  = ~\new_[19026]_  | ~\new_[18339]_ ;
  assign n3013 = \new_[14905]_  ? ld : \text_in[19] ;
  assign \new_[16945]_  = ~\new_[18254]_  | ~\new_[19000]_ ;
  assign \new_[16946]_  = ~\new_[19185]_  | ~\new_[21494]_ ;
  assign \new_[16947]_  = ~\new_[18149]_  | ~\new_[19624]_ ;
  assign n2903 = \new_[14769]_  ? \new_[19283]_  : \text_in[78] ;
  assign \new_[16949]_  = ~\new_[18962]_  & ~\new_[19172]_ ;
  assign n3053 = \new_[14948]_  ? \new_[18703]_  : \text_in[9] ;
  assign n3088 = \new_[15079]_  ? \new_[19497]_  : \text_in[110] ;
  assign \new_[16952]_  = ~\new_[19138]_  | ~\new_[18149]_ ;
  assign \new_[16953]_  = \\text_in_r_reg[115] ;
  assign \new_[16954]_  = ~\new_[17881]_ ;
  assign \new_[16955]_  = ~\new_[18023]_  | ~\new_[19111]_ ;
  assign \new_[16956]_  = ~\new_[20665]_  | ~\new_[19342]_ ;
  assign n3033 = \new_[14936]_  ? \new_[19283]_  : \text_in[12] ;
  assign \new_[16958]_  = ~\new_[17926]_ ;
  assign \new_[16959]_  = \new_[18547]_  | \new_[19084]_ ;
  assign n3118 = \new_[15634]_  ? \new_[19497]_  : \text_in[82] ;
  assign \new_[16961]_  = ~\new_[17652]_ ;
  assign n3098 = \new_[15259]_  ? ld : \text_in[104] ;
  assign \new_[16963]_  = ~\new_[17526]_ ;
  assign n2913 = \new_[14771]_  ? \new_[19414]_  : \text_in[86] ;
  assign \new_[16965]_  = ~\new_[18216]_  & ~\new_[18810]_ ;
  assign n2808 = \new_[14719]_  ? \new_[19497]_  : \text_in[68] ;
  assign \new_[16967]_  = \\text_in_r_reg[98] ;
  assign n2963 = \new_[14788]_  ? \new_[19283]_  : \text_in[118] ;
  assign \new_[16969]_  = ~\new_[18067]_  | ~\new_[18682]_ ;
  assign \new_[16970]_  = ~\new_[17783]_ ;
  assign n2838 = \new_[14755]_  ? \new_[19497]_  : \text_in[35] ;
  assign \new_[16972]_  = ~\new_[17737]_ ;
  assign \new_[16973]_  = ~\new_[18307]_  & ~\new_[17156]_ ;
  assign \new_[16974]_  = ~\new_[17657]_ ;
  assign n2993 = \new_[14877]_  ? \new_[19497]_  : \text_in[107] ;
  assign \new_[16976]_  = ~\new_[17848]_ ;
  assign \new_[16977]_  = ~\new_[17842]_ ;
  assign \new_[16978]_  = \new_[18363]_  | \new_[19298]_ ;
  assign \new_[16979]_  = ~\new_[21574]_  | ~\new_[18733]_ ;
  assign \new_[16980]_  = ~\new_[2500]_ ;
  assign \new_[16981]_  = ~\new_[19225]_  | ~\new_[19174]_ ;
  assign \new_[16982]_  = ~\new_[17716]_ ;
  assign \new_[16983]_  = ~\new_[21399]_ ;
  assign \new_[16984]_  = ~\new_[19000]_  & ~\new_[18389]_ ;
  assign \new_[16985]_  = ~\new_[17742]_ ;
  assign \new_[16986]_  = ~\new_[18376]_  | ~\new_[19053]_ ;
  assign \new_[16987]_  = ~\new_[17858]_ ;
  assign \new_[16988]_  = ~\new_[17622]_ ;
  assign n3158 = \new_[15840]_  ? \new_[19497]_  : \text_in[40] ;
  assign \new_[16990]_  = ~\new_[18350]_  | ~\new_[19324]_ ;
  assign \new_[16991]_  = ~\new_[18959]_  | ~\new_[18510]_ ;
  assign \new_[16992]_  = ~\new_[21634]_  & ~\new_[19096]_ ;
  assign \new_[16993]_  = ~\new_[18274]_  | ~\new_[19741]_ ;
  assign \new_[16994]_  = ~\new_[17466]_ ;
  assign \new_[16995]_  = \\text_in_r_reg[31] ;
  assign \new_[16996]_  = ~\new_[18104]_  | ~\new_[19064]_ ;
  assign \new_[16997]_  = ~\new_[18849]_ ;
  assign \new_[16998]_  = ~\new_[18002]_ ;
  assign \new_[16999]_  = ~\new_[17514]_ ;
  assign \new_[17000]_  = ~\new_[18219]_  | ~\new_[18947]_ ;
  assign \new_[17001]_  = ~\new_[18229]_  | ~\new_[19779]_ ;
  assign \new_[17002]_  = ~\new_[18165]_  & ~\new_[19779]_ ;
  assign \new_[17003]_  = ~\new_[19379]_  | ~\new_[18226]_ ;
  assign \new_[17004]_  = \\text_in_r_reg[122] ;
  assign \new_[17005]_  = ~\new_[17582]_ ;
  assign \new_[17006]_  = ~\new_[19063]_  | ~\new_[18861]_ ;
  assign \new_[17007]_  = ~\new_[20765]_  | ~\new_[19689]_ ;
  assign n2783 = \new_[14700]_  ? \new_[19414]_  : \text_in[14] ;
  assign \new_[17009]_  = ~\new_[18456]_  | ~\new_[19647]_ ;
  assign \new_[17010]_  = ~\new_[18093]_  | ~\new_[18148]_ ;
  assign \new_[17011]_  = ~\new_[20749]_  | ~\new_[18183]_ ;
  assign \new_[17012]_  = ~\new_[18793]_  | ~\new_[19676]_ ;
  assign \new_[17013]_  = \\text_in_r_reg[119] ;
  assign \new_[17014]_  = ~\new_[18252]_  & ~\new_[19268]_ ;
  assign \new_[17015]_  = \new_[19780]_  & \new_[18076]_ ;
  assign \new_[17016]_  = ~\new_[18994]_  & ~\new_[19014]_ ;
  assign \new_[17017]_  = ~\new_[17692]_ ;
  assign \new_[17018]_  = ~\new_[18172]_  | ~\new_[21517]_ ;
  assign \new_[17019]_  = ~\new_[17923]_ ;
  assign \new_[17020]_  = ~\new_[17715]_ ;
  assign n3188 = ~\new_[18113]_  & ~\new_[19363]_ ;
  assign n3018 = \new_[14909]_  ? \new_[19497]_  : \text_in[56] ;
  assign \new_[17023]_  = \new_[17432]_  ^ \new_[1862]_ ;
  assign \new_[17024]_  = ~\new_[18024]_  | ~\new_[19435]_ ;
  assign \new_[17025]_  = ~\new_[18526]_  | ~\new_[19189]_ ;
  assign \new_[17026]_  = \new_[17582]_ ;
  assign \new_[17027]_  = ~\new_[18284]_  | ~\new_[18795]_ ;
  assign \new_[17028]_  = \new_[18461]_  | \new_[18008]_ ;
  assign \new_[17029]_  = ~\new_[17504]_ ;
  assign \new_[17030]_  = \\text_in_r_reg[102] ;
  assign \new_[17031]_  = ~\new_[18256]_  | ~\new_[19741]_ ;
  assign \new_[17032]_  = ~\new_[17476]_ ;
  assign \new_[17033]_  = ~\new_[17961]_ ;
  assign \new_[17034]_  = ~\new_[18312]_  | ~\new_[21656]_ ;
  assign n3203 = \new_[15855]_  ? \new_[19497]_  : \text_in[88] ;
  assign \new_[17036]_  = ~\new_[17724]_ ;
  assign n2938 = \new_[14778]_  ? \new_[19497]_  : \text_in[60] ;
  assign \new_[17038]_  = \new_[18156]_  | \new_[19676]_ ;
  assign \new_[17039]_  = ~\new_[18299]_  & ~\new_[19555]_ ;
  assign \new_[17040]_  = ~\new_[17859]_ ;
  assign \new_[17041]_  = ~\new_[19145]_  & ~\new_[1025]_ ;
  assign \new_[17042]_  = ~\new_[17735]_ ;
  assign \new_[17043]_  = ~\new_[17947]_ ;
  assign \new_[17044]_  = ~\new_[18477]_  | ~\new_[19197]_ ;
  assign \new_[17045]_  = ~\new_[19100]_  | ~\new_[18841]_ ;
  assign \new_[17046]_  = \\text_in_r_reg[76] ;
  assign \new_[17047]_  = ~\new_[17867]_ ;
  assign \new_[17048]_  = ~\new_[18049]_  | ~\new_[21516]_ ;
  assign \new_[17049]_  = ~\new_[21098]_  | ~\new_[21100]_ ;
  assign n3063 = \new_[14960]_  ? \new_[19497]_  : \text_in[45] ;
  assign \new_[17051]_  = ~\new_[18496]_ ;
  assign \new_[17052]_  = ~\new_[17868]_ ;
  assign \new_[17053]_  = \\text_in_r_reg[113] ;
  assign \new_[17054]_  = ~\new_[17601]_ ;
  assign \new_[17055]_  = ~\new_[17850]_ ;
  assign \new_[17056]_  = ~\new_[18527]_  | ~\new_[19087]_ ;
  assign \new_[17057]_  = ~\new_[18681]_  | ~\new_[19117]_ ;
  assign \new_[17058]_  = ~\new_[18277]_  | ~\new_[20869]_ ;
  assign n2988 = \new_[14851]_  ? \new_[19497]_  : \text_in[92] ;
  assign \new_[17060]_  = ~\new_[18327]_  & ~\new_[21697]_ ;
  assign \new_[17061]_  = ~\new_[18681]_  | ~\new_[19675]_ ;
  assign \new_[17062]_  = ~\new_[18223]_  | ~\new_[19603]_ ;
  assign \new_[17063]_  = ~\new_[17769]_ ;
  assign \new_[17064]_  = ~\new_[2500]_  | ~\new_[18194]_ ;
  assign \new_[17065]_  = ~\new_[17821]_ ;
  assign \new_[17066]_  = ~\new_[18396]_  & ~\new_[19555]_ ;
  assign \new_[17067]_  = ~\new_[18582]_  | ~\new_[19679]_ ;
  assign \new_[17068]_  = ~\new_[18376]_  | ~\new_[18692]_ ;
  assign n2908 = \new_[14770]_  ? \new_[19283]_  : \text_in[81] ;
  assign \new_[17070]_  = ~\new_[18412]_ ;
  assign \new_[17071]_  = ~\new_[18146]_  | ~\new_[19146]_ ;
  assign \new_[17072]_  = ~\new_[17753]_ ;
  assign \new_[17073]_  = ~\new_[18424]_  & ~\new_[19741]_ ;
  assign \new_[17074]_  = ~\new_[17503]_ ;
  assign \new_[17075]_  = \\text_in_r_reg[94] ;
  assign \new_[17076]_  = \new_[18313]_  & \new_[19555]_ ;
  assign \new_[17077]_  = ~\new_[17569]_ ;
  assign n2888 = \new_[14766]_  ? \new_[19283]_  : \text_in[55] ;
  assign \new_[17079]_  = ~\new_[18541]_  | ~\new_[19478]_ ;
  assign \new_[17080]_  = ~\new_[17854]_ ;
  assign \new_[17081]_  = ~\new_[17729]_ ;
  assign \new_[17082]_  = ~\new_[17531]_ ;
  assign \new_[17083]_  = ~\new_[17596]_ ;
  assign \new_[17084]_  = ~\new_[18962]_  & ~\new_[14690]_ ;
  assign \new_[17085]_  = ~\new_[18841]_  | ~\new_[19754]_ ;
  assign \new_[17086]_  = ~\new_[17969]_ ;
  assign \new_[17087]_  = \\text_in_r_reg[62] ;
  assign \new_[17088]_  = ~\new_[18197]_  | ~\new_[19295]_ ;
  assign \new_[17089]_  = ~\new_[20982]_ ;
  assign \new_[17090]_  = ~\new_[18404]_  | ~\new_[18968]_ ;
  assign \new_[17091]_  = \\text_in_r_reg[48] ;
  assign \new_[17092]_  = ~\new_[18242]_  & ~\new_[19285]_ ;
  assign \new_[17093]_  = ~\new_[17804]_ ;
  assign \new_[17094]_  = ~\new_[20298]_ ;
  assign \new_[17095]_  = ~\new_[17481]_ ;
  assign \new_[17096]_  = ~\new_[17641]_ ;
  assign \new_[17097]_  = ~\new_[17645]_ ;
  assign \new_[17098]_  = ~\new_[18075]_  & ~\new_[21575]_ ;
  assign n2883 = \new_[14765]_  ? \new_[19497]_  : \text_in[46] ;
  assign \new_[17100]_  = ~\new_[17561]_ ;
  assign \new_[17101]_  = ~\new_[18497]_  | ~\new_[18832]_ ;
  assign \new_[17102]_  = ~\new_[17794]_ ;
  assign n2898 = \new_[14768]_  ? ld : \text_in[63] ;
  assign \new_[17104]_  = ~\new_[18217]_  | ~\new_[19342]_ ;
  assign \new_[17105]_  = ~\new_[17911]_ ;
  assign \new_[17106]_  = ~\new_[19064]_  & ~\new_[1039]_ ;
  assign \new_[17107]_  = ~\new_[18151]_  & ~\new_[19000]_ ;
  assign \new_[17108]_  = ~\new_[17719]_ ;
  assign \new_[17109]_  = \new_[18353]_  & \new_[19665]_ ;
  assign \new_[17110]_  = \new_[16777]_  ^ \new_[1341]_ ;
  assign n3148 = \new_[15823]_  ? \new_[19283]_  : \text_in[74] ;
  assign \new_[17112]_  = ~\new_[17492]_ ;
  assign \new_[17113]_  = ~\new_[17628]_ ;
  assign \new_[17114]_  = ~\new_[19000]_  & ~\new_[18397]_ ;
  assign \new_[17115]_  = ~\new_[18012]_ ;
  assign \new_[17116]_  = \\text_in_r_reg[27] ;
  assign \new_[17117]_  = ~\new_[18392]_  | ~\new_[18454]_ ;
  assign n2848 = \new_[14758]_  ? ld : \text_in[17] ;
  assign \new_[17119]_  = ~\new_[17472]_ ;
  assign n3183 = \new_[15850]_  ? \new_[19283]_  : \text_in[20] ;
  assign \new_[17121]_  = ~\new_[18910]_  | ~\new_[18363]_ ;
  assign n2928 = \new_[14776]_  ? \new_[19414]_  : \text_in[91] ;
  assign \new_[17123]_  = ~\new_[17594]_ ;
  assign n2878 = \new_[14764]_  ? \new_[19497]_  : \text_in[29] ;
  assign \new_[17125]_  = \\text_in_r_reg[109] ;
  assign n3028 = \new_[14922]_  ? \new_[19497]_  : \text_in[69] ;
  assign n3198 = \new_[15854]_  ? \new_[19497]_  : \text_in[75] ;
  assign n2968 = \new_[14790]_  ? \new_[19283]_  : \text_in[59] ;
  assign \new_[17129]_  = \new_[14711]_  ^ \new_[19765]_ ;
  assign n3043 = \new_[14943]_  ? ld : \text_in[80] ;
  assign \new_[17131]_  = ~\new_[18269]_  & ~\new_[19050]_ ;
  assign \new_[17132]_  = ~\new_[17588]_ ;
  assign \new_[17133]_  = ~\new_[18071]_  & ~\new_[19637]_ ;
  assign n3143 = \new_[15819]_  ? \new_[19414]_  : \text_in[84] ;
  assign \new_[17135]_  = ~\new_[17843]_ ;
  assign \new_[17137]_  = ~\new_[17802]_ ;
  assign \new_[17138]_  = ~\new_[18236]_  | ~\new_[19298]_ ;
  assign \new_[17139]_  = ~\new_[19782]_  & ~\new_[18118]_ ;
  assign n3128 = \new_[15756]_  ? ld : \text_in[105] ;
  assign \new_[17141]_  = ~\new_[17662]_ ;
  assign \new_[17142]_  = ~\new_[18521]_  | ~\new_[18960]_ ;
  assign \new_[17143]_  = ~\new_[18024]_  | ~\new_[19675]_ ;
  assign \new_[17144]_  = ~\new_[17812]_ ;
  assign \new_[17145]_  = ~\new_[18016]_ ;
  assign \new_[17146]_  = \new_[18181]_  | \new_[19697]_ ;
  assign \new_[17147]_  = ~\new_[17523]_ ;
  assign \new_[17148]_  = \\text_in_r_reg[117] ;
  assign \new_[17149]_  = ~\new_[18159]_  & ~\new_[19444]_ ;
  assign n3093 = \new_[15147]_  ? \new_[19283]_  : \text_in[30] ;
  assign n2923 = \new_[14773]_  ? \new_[19283]_  : \text_in[99] ;
  assign \new_[17152]_  = ~\new_[18405]_  | ~\new_[21584]_ ;
  assign \new_[17153]_  = ~\new_[17876]_ ;
  assign \new_[17154]_  = ~\new_[18255]_  | ~\new_[21657]_ ;
  assign \new_[17155]_  = ~\new_[18045]_ ;
  assign \new_[17156]_  = \\u0_r0_rcnt_reg[0] ;
  assign n2918 = \new_[14772]_  ? \new_[19497]_  : \text_in[8] ;
  assign \new_[17158]_  = ~\new_[18497]_  | ~\new_[19676]_ ;
  assign \new_[17159]_  = ~\new_[18458]_  & ~\new_[19104]_ ;
  assign n2873 = \new_[14763]_  ? \new_[19497]_  : \text_in[26] ;
  assign n3078 = \new_[15062]_  ? \new_[19283]_  : \text_in[10] ;
  assign \new_[17162]_  = ~\new_[20665]_  | ~\new_[21656]_ ;
  assign n3003 = \new_[14899]_  ? \new_[18703]_  : \text_in[77] ;
  assign \new_[17164]_  = ~\new_[18376]_  | ~\new_[19132]_ ;
  assign \new_[17165]_  = ~\new_[17717]_ ;
  assign \new_[17166]_  = ~\new_[19268]_  & ~\new_[21641]_ ;
  assign \new_[17167]_  = ~\new_[18484]_  & ~\new_[19098]_ ;
  assign \new_[17168]_  = ~\new_[19100]_  & ~\new_[18190]_ ;
  assign \new_[17169]_  = ~\new_[17647]_ ;
  assign \new_[17170]_  = ~\new_[17674]_ ;
  assign \new_[17171]_  = ~\new_[17602]_ ;
  assign \new_[17172]_  = ~\new_[17586]_ ;
  assign \new_[17173]_  = ~\new_[17877]_ ;
  assign \new_[17174]_  = ~\new_[18230]_  & ~\new_[21569]_ ;
  assign \new_[17175]_  = \new_[18447]_  | \new_[19066]_ ;
  assign \new_[17176]_  = ~\new_[18452]_  | ~\new_[19376]_ ;
  assign n2933 = \new_[14777]_  ? \new_[19497]_  : \text_in[39] ;
  assign \new_[17178]_  = ~\new_[18108]_  | ~\new_[21569]_ ;
  assign \new_[17179]_  = \new_[18283]_  | \new_[19253]_ ;
  assign \new_[17180]_  = ~\new_[21483]_  | ~\new_[19268]_ ;
  assign \new_[17181]_  = ~\new_[18456]_  | ~\new_[19023]_ ;
  assign \new_[17182]_  = ~\new_[17994]_ ;
  assign \new_[17183]_  = ~\new_[18456]_  | ~\new_[19788]_ ;
  assign n3113 = \new_[15482]_  ? ld : \text_in[7] ;
  assign \new_[17185]_  = ~\new_[17728]_ ;
  assign \new_[17186]_  = ~\new_[18518]_  & ~\new_[19434]_ ;
  assign n3168 = \new_[15843]_  ? \new_[18703]_  : \text_in[121] ;
  assign \new_[17188]_  = ~\new_[18110]_  | ~\new_[18394]_ ;
  assign \new_[17189]_  = ~\new_[19624]_  & ~\new_[18232]_ ;
  assign \new_[17190]_  = ~\new_[18127]_  | ~\new_[18968]_ ;
  assign \new_[17191]_  = ~\new_[17603]_ ;
  assign \new_[17192]_  = ~\new_[18282]_  & ~\new_[19679]_ ;
  assign \new_[17193]_  = ~\new_[17656]_ ;
  assign \new_[17194]_  = \new_[18297]_  & \new_[19675]_ ;
  assign \new_[17195]_  = ~\new_[18477]_  & ~\new_[18973]_ ;
  assign \new_[17196]_  = ~\new_[19413]_  & ~\new_[18053]_ ;
  assign \new_[17197]_  = ~\new_[18092]_  | ~\new_[19416]_ ;
  assign n2818 = \new_[14725]_  ? ld : \text_in[42] ;
  assign \new_[17199]_  = ~\new_[18243]_  | ~\new_[18680]_ ;
  assign \new_[17200]_  = ~\new_[17670]_ ;
  assign \new_[17201]_  = \\text_in_r_reg[21] ;
  assign \new_[17202]_  = ~\new_[18211]_  & ~\new_[19379]_ ;
  assign \new_[17203]_  = ~\new_[18251]_  | ~\new_[21489]_ ;
  assign \new_[17204]_  = ~\new_[18549]_  | ~\new_[19485]_ ;
  assign \new_[17205]_  = ~\new_[18281]_  | ~\new_[17886]_ ;
  assign \new_[17206]_  = ~\new_[18809]_  & ~\new_[18164]_ ;
  assign \new_[17207]_  = \new_[18134]_  | \new_[19697]_ ;
  assign \new_[17208]_  = ~\new_[17675]_ ;
  assign \new_[17209]_  = ~\new_[19100]_  | ~\new_[18459]_ ;
  assign \new_[17210]_  = ~\new_[18352]_  | ~\new_[21516]_ ;
  assign \new_[17211]_  = ~\new_[18571]_  | ~\new_[21306]_ ;
  assign \new_[17212]_  = ~\new_[17589]_ ;
  assign \new_[17213]_  = \new_[18578]_  & \new_[19685]_ ;
  assign \new_[17214]_  = \new_[18793]_  & \new_[19738]_ ;
  assign \new_[17215]_  = ~\new_[18478]_  & ~\new_[19675]_ ;
  assign \new_[17216]_  = \new_[18234]_  | \new_[18371]_ ;
  assign \new_[17217]_  = ~\new_[18400]_  & ~\new_[19026]_ ;
  assign \new_[17218]_  = ~\new_[19386]_  | ~\new_[18085]_ ;
  assign \new_[17219]_  = ~\new_[18350]_  | ~\new_[19354]_ ;
  assign \new_[17220]_  = ~\new_[21574]_  & ~\new_[18566]_ ;
  assign \new_[17221]_  = ~\new_[18565]_  | ~\new_[18995]_ ;
  assign \new_[17222]_  = \new_[18088]_  | \new_[19335]_ ;
  assign \new_[17223]_  = \new_[18374]_  | \new_[19098]_ ;
  assign n2948 = \new_[14780]_  ? \new_[19497]_  : \text_in[23] ;
  assign \new_[17225]_  = ~\new_[18330]_  | ~\new_[19554]_ ;
  assign \new_[17226]_  = ~\new_[18243]_  | ~\new_[19092]_ ;
  assign \new_[17227]_  = ~\new_[21578]_  | ~\new_[21400]_ ;
  assign n2953 = \new_[14781]_  ? \new_[19497]_  : \text_in[58] ;
  assign \new_[17229]_  = ~\new_[17800]_ ;
  assign \new_[17230]_  = ~\new_[17655]_ ;
  assign \new_[17231]_  = ~\new_[18521]_  | ~\new_[19597]_ ;
  assign n2843 = \new_[14756]_  ? \new_[19283]_  : \text_in[6] ;
  assign \new_[17233]_  = ~\new_[18238]_  & ~\new_[19203]_ ;
  assign n3133 = \new_[15757]_  ? \new_[19283]_  : \text_in[13] ;
  assign \new_[17235]_  = ~\new_[17826]_ ;
  assign \new_[17236]_  = ~\new_[19053]_  | ~\new_[18420]_ ;
  assign \new_[17237]_  = ~\new_[18813]_  & (~\new_[18589]_  | ~\new_[6746]_ );
  assign \new_[17238]_  = ~\new_[18195]_  | ~\new_[19444]_ ;
  assign \new_[17239]_  = ~\new_[18248]_  | ~\new_[18960]_ ;
  assign \new_[17240]_  = ~\new_[18169]_  | ~\new_[19435]_ ;
  assign \new_[17241]_  = \new_[18442]_  | \new_[19277]_ ;
  assign \new_[17242]_  = \new_[18239]_  | \new_[19642]_ ;
  assign \new_[17243]_  = ~\new_[19108]_  | ~\new_[19132]_ ;
  assign \new_[17244]_  = \new_[18046]_  | \new_[19599]_ ;
  assign \new_[17245]_  = ~\new_[17896]_ ;
  assign \new_[17246]_  = ~\new_[19234]_  | ~\new_[19750]_ ;
  assign \new_[17247]_  = ~\new_[17494]_ ;
  assign \new_[17248]_  = ~\new_[21611]_  | ~\new_[18968]_ ;
  assign \new_[17249]_  = ~\new_[17599]_ ;
  assign \new_[17250]_  = ~\new_[18196]_  | ~\new_[19655]_ ;
  assign \new_[17251]_  = ~\new_[18535]_  | ~\new_[20499]_ ;
  assign \new_[17252]_  = ~\new_[19059]_  & ~\new_[999]_ ;
  assign \new_[17253]_  = ~\new_[18013]_ ;
  assign \new_[17254]_  = ~\new_[18352]_  | ~\new_[21517]_ ;
  assign \new_[17255]_  = \new_[19250]_  & \new_[19717]_ ;
  assign \new_[17256]_  = \new_[18382]_  | \new_[19389]_ ;
  assign \new_[17257]_  = ~\new_[21259]_  & ~\new_[18516]_ ;
  assign \new_[17258]_  = ~\new_[18523]_  | ~\new_[19554]_ ;
  assign \new_[17259]_  = \new_[18032]_  | \new_[19337]_ ;
  assign \new_[17260]_  = ~\new_[17945]_ ;
  assign \new_[17261]_  = ~\new_[20932]_  | ~\new_[19670]_ ;
  assign \new_[17262]_  = ~\new_[18562]_  & ~\new_[18810]_ ;
  assign \new_[17263]_  = ~\new_[17827]_ ;
  assign \new_[17264]_  = ~\new_[17871]_ ;
  assign \new_[17265]_  = ~\new_[19503]_  | ~\new_[19654]_  | ~\new_[19253]_  | ~\new_[19087]_ ;
  assign \new_[17266]_  = ~\new_[20495]_  | ~\new_[18261]_ ;
  assign \new_[17267]_  = ~\new_[18259]_  | ~\new_[18945]_ ;
  assign \new_[17268]_  = ~\new_[18274]_  | ~\new_[19420]_ ;
  assign \new_[17269]_  = ~\new_[19254]_  | ~\new_[18274]_ ;
  assign \new_[17270]_  = \new_[12138]_  ^ \new_[18777]_ ;
  assign \new_[17271]_  = ~\new_[17480]_ ;
  assign n3038 = \new_[14941]_  ? \new_[19283]_  : \text_in[85] ;
  assign \new_[17273]_  = ~\new_[20098]_ ;
  assign \new_[17274]_  = \new_[15854]_  ^ \new_[1431]_ ;
  assign \new_[17275]_  = ~\new_[18222]_  | ~\new_[18676]_ ;
  assign n3163 = \new_[15842]_  ? \new_[19497]_  : \text_in[15] ;
  assign \new_[17277]_  = ~\new_[17906]_ ;
  assign \new_[17278]_  = ~\new_[17888]_ ;
  assign \new_[17279]_  = ~\new_[18352]_  | ~\new_[18947]_ ;
  assign \new_[17280]_  = ~\new_[17863]_ ;
  assign n3208 = \new_[15861]_  ? \new_[19497]_  : \text_in[33] ;
  assign \new_[17282]_  = ~\new_[17672]_ ;
  assign \new_[17283]_  = ~\new_[18314]_  | ~\new_[18959]_ ;
  assign \new_[17284]_  = ~\new_[18561]_  & ~\new_[18664]_ ;
  assign \new_[17285]_  = ~\new_[18789]_ ;
  assign n3178 = \new_[15846]_  ? \new_[19497]_  : \text_in[36] ;
  assign \new_[17287]_  = ~\new_[17825]_ ;
  assign n2803 = \new_[14711]_  ? \new_[19283]_  : \text_in[0] ;
  assign \new_[17289]_  = ~\new_[17919]_ ;
  assign n2828 = \new_[14752]_  ? \new_[19283]_  : \text_in[64] ;
  assign n2768 = \new_[14696]_  ? \new_[19283]_  : \text_in[116] ;
  assign \new_[17292]_  = ~\new_[17861]_ ;
  assign n3153 = \new_[15839]_  ? \new_[18703]_  : \text_in[16] ;
  assign n3138 = \new_[15815]_  ? ld : \text_in[120] ;
  assign \new_[17295]_  = \new_[17918]_ ;
  assign \new_[17296]_  = ~\new_[17857]_ ;
  assign n2813 = \new_[14722]_  ? \new_[19283]_  : \text_in[49] ;
  assign \new_[17298]_  = ~\new_[18964]_  | ~\new_[18533]_ ;
  assign n3123 = \new_[15703]_  ? \new_[19497]_  : \text_in[126] ;
  assign \new_[17300]_  = \new_[18577]_  & \new_[19328]_ ;
  assign \new_[17301]_  = ~\new_[18491]_  | ~\new_[19413]_ ;
  assign \new_[17302]_  = \\text_in_r_reg[5] ;
  assign n2778 = \new_[14698]_  ? \new_[19497]_  : \text_in[37] ;
  assign \new_[17304]_  = ~\new_[17963]_ ;
  assign \new_[17305]_  = \new_[19610]_  ^ \new_[1862]_ ;
  assign \new_[17306]_  = ~\new_[18580]_  | ~\new_[21046]_ ;
  assign \new_[17307]_  = ~\new_[19150]_  | ~\new_[18536]_ ;
  assign \new_[17308]_  = ~\new_[19165]_  | ~\new_[18605]_ ;
  assign \new_[17309]_  = \new_[12134]_  ^ \new_[18813]_ ;
  assign \new_[17310]_  = \new_[14767]_  ^ \new_[19305]_ ;
  assign \new_[17311]_  = ~\new_[19182]_  | ~\new_[18176]_ ;
  assign \new_[17312]_  = ~\new_[17973]_ ;
  assign \new_[17313]_  = ~\new_[17865]_ ;
  assign \new_[17314]_  = ~\new_[21570]_  | ~\new_[18351]_ ;
  assign \new_[17315]_  = \new_[16701]_  ^ \new_[1417]_ ;
  assign \new_[17316]_  = ~\new_[18462]_  | ~\new_[19503]_ ;
  assign \new_[17317]_  = ~\new_[18708]_  | ~\new_[18108]_ ;
  assign \new_[17318]_  = \new_[14851]_  ^ \new_[19306]_ ;
  assign \new_[17319]_  = \new_[19784]_  ^ \new_[18829]_ ;
  assign \new_[17320]_  = \new_[16848]_  ^ \new_[2346]_ ;
  assign \new_[17321]_  = ~\new_[19125]_  & ~\new_[19435]_ ;
  assign \new_[17322]_  = ~\new_[18368]_  | ~\new_[19412]_ ;
  assign \new_[17323]_  = ~\new_[18046]_  & ~\new_[946]_ ;
  assign \new_[17324]_  = ~\new_[21514]_  & ~\new_[18637]_ ;
  assign \new_[17325]_  = ~\new_[18006]_ ;
  assign \new_[17326]_  = ~\new_[18082]_  | ~\new_[19676]_ ;
  assign \new_[17327]_  = ~\new_[17626]_ ;
  assign \new_[17328]_  = ~\new_[17683]_ ;
  assign \new_[17329]_  = ~\new_[17799]_ ;
  assign \new_[17330]_  = ~\new_[21533]_  & ~\new_[18605]_ ;
  assign n2893 = \new_[14767]_  ? \new_[19414]_  : \text_in[61] ;
  assign \new_[17332]_  = ~\new_[17567]_ ;
  assign \new_[17333]_  = ~\new_[17546]_ ;
  assign \new_[17334]_  = \new_[20490]_  | \new_[21514]_ ;
  assign \new_[17335]_  = ~\new_[17801]_ ;
  assign \new_[17336]_  = \new_[18394]_  & \new_[19330]_ ;
  assign \new_[17337]_  = ~\new_[17495]_ ;
  assign \new_[17338]_  = ~\new_[17489]_ ;
  assign \new_[17339]_  = ~\new_[17997]_ ;
  assign \new_[17340]_  = ~\new_[18327]_  | ~\new_[21685]_ ;
  assign \new_[17341]_  = ~\new_[18173]_  | ~\new_[19379]_ ;
  assign \new_[17342]_  = ~\new_[17700]_ ;
  assign \new_[17343]_  = ~\new_[18543]_  | ~\new_[18284]_ ;
  assign \new_[17344]_  = ~\new_[18000]_ ;
  assign \new_[17345]_  = \new_[18337]_  & \new_[19368]_ ;
  assign \new_[17346]_  = ~\new_[17785]_ ;
  assign \new_[17347]_  = ~\new_[17786]_ ;
  assign \new_[17348]_  = ~\new_[17587]_ ;
  assign \new_[17349]_  = ~\new_[17763]_ ;
  assign \new_[17350]_  = ~\new_[18227]_  & ~\new_[19096]_ ;
  assign \new_[17351]_  = ~\new_[17928]_ ;
  assign \new_[17352]_  = ~\new_[17806]_ ;
  assign \new_[17353]_  = ~\new_[17726]_ ;
  assign \new_[17354]_  = ~\new_[21532]_  | ~\new_[21517]_ ;
  assign \new_[17355]_  = ~\new_[17760]_ ;
  assign \new_[17356]_  = ~\new_[21658]_  & ~\new_[21686]_ ;
  assign \new_[17357]_  = ~\new_[17618]_ ;
  assign \new_[17358]_  = ~\new_[18656]_ ;
  assign \new_[17359]_  = ~\new_[17932]_ ;
  assign \new_[17360]_  = ~\new_[18477]_  | ~\new_[18973]_ ;
  assign \new_[17361]_  = ~\new_[17805]_ ;
  assign \new_[17362]_  = ~\new_[18801]_  & ~\new_[18448]_ ;
  assign \new_[17363]_  = ~\new_[17762]_ ;
  assign \new_[17364]_  = \new_[18548]_  | \new_[19413]_ ;
  assign \new_[17365]_  = ~\new_[18139]_  & ~\new_[19426]_ ;
  assign \new_[17366]_  = ~\new_[20235]_  | ~\new_[20870]_ ;
  assign \new_[17367]_  = ~\new_[17754]_ ;
  assign \new_[17368]_  = \new_[17938]_ ;
  assign \new_[17369]_  = ~\new_[17981]_ ;
  assign \new_[17370]_  = ~\new_[18573]_  & ~\new_[19105]_ ;
  assign \new_[17371]_  = ~\new_[17879]_ ;
  assign \new_[17372]_  = ~\new_[18535]_  | ~\new_[19679]_ ;
  assign \new_[17373]_  = ~\new_[17615]_ ;
  assign n3173 = \new_[15845]_  ? \new_[19283]_  : \text_in[41] ;
  assign \new_[17375]_  = ~\new_[18025]_  & ~\new_[19203]_ ;
  assign \new_[17376]_  = ~\new_[18457]_  | ~\new_[21397]_ ;
  assign \new_[17377]_  = ~\new_[17870]_ ;
  assign \new_[17378]_  = ~\new_[17584]_ ;
  assign \new_[17379]_  = \new_[16980]_  | \new_[18194]_ ;
  assign \new_[17380]_  = \new_[21570]_  & \new_[19191]_ ;
  assign \new_[17381]_  = ~\new_[18827]_ ;
  assign \new_[17382]_  = ~\new_[18542]_  & ~\new_[19136]_ ;
  assign \new_[17383]_  = ~\new_[18365]_  | ~\new_[19474]_ ;
  assign \new_[17384]_  = ~\new_[20699]_  | ~\new_[18975]_ ;
  assign \new_[17385]_  = ~\new_[17537]_ ;
  assign \new_[17386]_  = ~\new_[17535]_ ;
  assign \new_[17387]_  = ~\new_[18271]_ ;
  assign \new_[17388]_  = ~\new_[17520]_ ;
  assign \new_[17389]_  = ~\new_[17511]_ ;
  assign \new_[17390]_  = \new_[2500]_  | \new_[19553]_ ;
  assign \new_[17391]_  = ~\new_[17490]_ ;
  assign \new_[17392]_  = ~\new_[19398]_  & ~\new_[19474]_ ;
  assign \new_[17393]_  = ~\new_[17956]_ ;
  assign \new_[17394]_  = ~\new_[18458]_  & ~\new_[19754]_ ;
  assign \new_[17395]_  = ~\new_[17658]_ ;
  assign \new_[17396]_  = ~\new_[18571]_  | ~\new_[21655]_ ;
  assign \new_[17397]_  = \\text_in_r_reg[22] ;
  assign n2798 = \new_[14709]_  ? ld : \text_in[18] ;
  assign \new_[17399]_  = ~\new_[17970]_ ;
  assign \new_[17400]_  = \\text_in_r_reg[83] ;
  assign \new_[17401]_  = ~\new_[17765]_ ;
  assign \new_[17402]_  = ~\new_[17707]_ ;
  assign \new_[17403]_  = ~\new_[17712]_ ;
  assign \new_[17404]_  = \\text_in_r_reg[38] ;
  assign \new_[17405]_  = \new_[18122]_  & \new_[19676]_ ;
  assign \new_[17406]_  = ~\new_[17498]_ ;
  assign \new_[17407]_  = ~\new_[18048]_  & ~\new_[19047]_ ;
  assign \new_[17408]_  = ~\new_[19741]_  | ~\new_[18546]_ ;
  assign \new_[17409]_  = \new_[19450]_  & \new_[19787]_ ;
  assign \new_[17410]_  = ~\new_[17571]_ ;
  assign \new_[17411]_  = \new_[19687]_  & \new_[19813]_ ;
  assign \new_[17412]_  = ~\new_[17516]_ ;
  assign \new_[17413]_  = ~\new_[18567]_  & ~\new_[19269]_ ;
  assign \new_[17414]_  = ~\new_[18054]_  & ~\new_[21570]_ ;
  assign \new_[17415]_  = \new_[18554]_  & \new_[19354]_ ;
  assign \new_[17416]_  = ~\new_[17676]_ ;
  assign \new_[17417]_  = ~\new_[18241]_  | ~\new_[19020]_ ;
  assign \new_[17418]_  = ~\new_[19227]_  | ~\new_[21494]_ ;
  assign n3068 = \new_[14962]_  ? \new_[19283]_  : \text_in[52] ;
  assign \new_[17420]_  = ~\new_[17828]_ ;
  assign \new_[17421]_  = ~\new_[18130]_  & ~\new_[19212]_ ;
  assign \new_[17422]_  = ~\new_[17673]_ ;
  assign \new_[17423]_  = \new_[19100]_  | \new_[19754]_ ;
  assign \new_[17424]_  = ~\new_[18248]_  | ~\new_[19379]_ ;
  assign \new_[17425]_  = ~\new_[17988]_ ;
  assign \new_[17426]_  = ~\new_[17992]_ ;
  assign \new_[17427]_  = \new_[19801]_  | \new_[18008]_ ;
  assign \new_[17428]_  = ~\new_[17696]_ ;
  assign n3103 = \new_[15272]_  ? \new_[19497]_  : \text_in[65] ;
  assign \new_[17430]_  = \\text_in_r_reg[71] ;
  assign \new_[17431]_  = ~\new_[17937]_ ;
  assign \new_[17432]_  = \\text_in_r_reg[89] ;
  assign \new_[17433]_  = ~\new_[17636]_ ;
  assign \new_[17434]_  = ~\new_[17999]_ ;
  assign \new_[17435]_  = ~\new_[19113]_  | ~\new_[19603]_ ;
  assign \new_[17436]_  = ~\new_[17984]_ ;
  assign \new_[17437]_  = ~\new_[17620]_ ;
  assign \new_[17438]_  = ~\new_[17630]_ ;
  assign \new_[17439]_  = ~\new_[19159]_  | ~\new_[18228]_ ;
  assign \new_[17440]_  = \new_[19568]_  & \new_[18317]_ ;
  assign \new_[17441]_  = ~\new_[18001]_ ;
  assign n2823 = \new_[14750]_  ? \new_[19283]_  : \text_in[127] ;
  assign \new_[17443]_  = ~\new_[18136]_  & ~\new_[18664]_ ;
  assign \new_[17444]_  = ~\new_[17485]_ ;
  assign \new_[17445]_  = ~\new_[17746]_ ;
  assign \new_[17446]_  = ~\new_[17780]_ ;
  assign \new_[17447]_  = ~\new_[19727]_ ;
  assign \new_[17448]_  = \\text_in_r_reg[87] ;
  assign \new_[17449]_  = ~\new_[18203]_  | ~\new_[19734]_ ;
  assign \new_[17450]_  = ~\new_[18302]_  & ~\new_[19788]_ ;
  assign \new_[17451]_  = \new_[18607]_  & \new_[18414]_ ;
  assign \new_[17452]_  = ~\new_[18031]_ ;
  assign \new_[17453]_  = ~\new_[17519]_ ;
  assign \new_[17454]_  = ~\new_[17530]_ ;
  assign \new_[17455]_  = ~\new_[18019]_ ;
  assign \new_[17456]_  = ~\new_[18336]_  | ~\new_[19484]_ ;
  assign \new_[17457]_  = ~\new_[18943]_ ;
  assign \new_[17458]_  = ~\new_[18376]_ ;
  assign \new_[17459]_  = ~\new_[18841]_ ;
  assign \new_[17460]_  = ~\new_[18613]_  & ~\new_[19301]_ ;
  assign \new_[17461]_  = ~\new_[18022]_ ;
  assign \new_[17462]_  = ~\new_[18850]_  | ~\new_[19420]_ ;
  assign \new_[17463]_  = ~\new_[18059]_ ;
  assign \new_[17464]_  = ~\new_[18720]_  | ~\new_[21522]_ ;
  assign \new_[17465]_  = ~\new_[18839]_  | ~\new_[19685]_ ;
  assign \new_[17466]_  = ~\new_[18552]_ ;
  assign \new_[17467]_  = ~\new_[18030]_ ;
  assign \new_[17468]_  = ~\new_[18568]_ ;
  assign \new_[17469]_  = ~\new_[18674]_ ;
  assign \new_[17470]_  = \new_[19013]_  & \new_[19638]_ ;
  assign \new_[17471]_  = ~\new_[18193]_ ;
  assign \new_[17472]_  = \new_[19094]_ ;
  assign \new_[17473]_  = ~\new_[18686]_  & ~\new_[21572]_ ;
  assign \new_[17474]_  = ~\new_[21492]_  & ~\new_[19462]_ ;
  assign \new_[17475]_  = ~\new_[18194]_ ;
  assign \new_[17476]_  = \new_[18461]_ ;
  assign \new_[17477]_  = ~\new_[18604]_  | ~\new_[18956]_ ;
  assign \new_[17478]_  = ~\new_[18863]_  & ~\new_[921]_ ;
  assign \new_[17479]_  = ~\new_[18660]_  | ~\new_[21657]_ ;
  assign \new_[17480]_  = ~\new_[18884]_  | ~\new_[19660]_ ;
  assign \new_[17481]_  = ~\new_[19596]_  | ~\new_[19173]_  | ~\new_[19140]_ ;
  assign \new_[17482]_  = ~\new_[18449]_ ;
  assign \new_[17483]_  = \new_[18841]_  & \new_[19398]_ ;
  assign \new_[17484]_  = ~\new_[18390]_ ;
  assign \new_[17485]_  = ~\new_[18034]_ ;
  assign \new_[17486]_  = ~\new_[18446]_ ;
  assign \new_[17487]_  = \new_[14779]_  ^ \new_[2344]_ ;
  assign \new_[17488]_  = ~\new_[18063]_ ;
  assign \new_[17489]_  = ~\new_[18051]_ ;
  assign \new_[17490]_  = \new_[18549]_ ;
  assign \new_[17491]_  = ~\new_[18676]_  | ~\new_[19675]_ ;
  assign \new_[17492]_  = ~\new_[18688]_  | ~\new_[20746]_ ;
  assign \new_[17493]_  = ~\new_[18900]_  | ~\new_[18939]_ ;
  assign \new_[17494]_  = ~\new_[19670]_  & ~\new_[20933]_ ;
  assign \new_[17495]_  = ~\new_[19625]_  | ~\new_[21165]_ ;
  assign \new_[17496]_  = ~\new_[18480]_ ;
  assign \new_[17497]_  = ~\new_[18065]_ ;
  assign \new_[17498]_  = \new_[18043]_ ;
  assign \new_[17499]_  = ~\new_[19344]_  & ~\new_[21660]_ ;
  assign \new_[17500]_  = \new_[15272]_  ^ \new_[19657]_ ;
  assign \new_[17501]_  = ~\new_[18698]_  & ~\new_[20237]_ ;
  assign \new_[17502]_  = ~\new_[19503]_  | ~\new_[18834]_ ;
  assign \new_[17503]_  = ~\new_[18688]_  | ~\new_[18974]_ ;
  assign \new_[17504]_  = ~\new_[18653]_  | ~\new_[21494]_ ;
  assign \new_[17505]_  = ~\new_[18447]_ ;
  assign \new_[17506]_  = ~\new_[18924]_  & ~\new_[19734]_ ;
  assign \new_[17507]_  = ~\new_[18475]_ ;
  assign \new_[17508]_  = \new_[19811]_  ^ \new_[1518]_ ;
  assign \new_[17509]_  = ~\new_[18486]_ ;
  assign \new_[17510]_  = ~\new_[18837]_  | ~\new_[19788]_ ;
  assign \new_[17511]_  = ~\new_[18274]_ ;
  assign \new_[17512]_  = ~\new_[19539]_  | ~\new_[18674]_ ;
  assign \new_[17513]_  = ~\new_[21483]_  | ~\new_[19413]_ ;
  assign \new_[17514]_  = ~\new_[18433]_ ;
  assign \new_[17515]_  = ~\new_[18806]_  | ~\new_[19435]_ ;
  assign \new_[17516]_  = ~\new_[18261]_ ;
  assign \new_[17517]_  = \new_[17148]_  ^ \new_[1345]_ ;
  assign \new_[17518]_  = ~\new_[18084]_ ;
  assign \new_[17519]_  = ~\new_[18148]_ ;
  assign \new_[17520]_  = ~\new_[18248]_ ;
  assign \new_[17521]_  = ~\new_[18093]_ ;
  assign \new_[17522]_  = ~\new_[18559]_ ;
  assign \new_[17523]_  = ~\new_[18028]_ ;
  assign \new_[17524]_  = \new_[19716]_  ^ \new_[1667]_ ;
  assign \new_[17525]_  = ~\new_[18180]_ ;
  assign \new_[17526]_  = ~\new_[18230]_ ;
  assign \new_[17527]_  = ~\new_[18535]_ ;
  assign \new_[17528]_  = ~\new_[18244]_ ;
  assign \new_[17529]_  = ~\new_[18199]_ ;
  assign \new_[17530]_  = ~\new_[18580]_ ;
  assign \new_[17531]_  = ~\new_[18797]_  | ~\new_[19674]_ ;
  assign \new_[17532]_  = ~\new_[18096]_ ;
  assign \new_[17533]_  = ~\new_[18459]_ ;
  assign \new_[17534]_  = ~\new_[18204]_ ;
  assign \new_[17535]_  = \new_[18203]_ ;
  assign \new_[17536]_  = ~\new_[18372]_ ;
  assign \new_[17537]_  = ~\new_[19547]_  & ~\new_[1879]_ ;
  assign \new_[17538]_  = \new_[19800]_  ^ \new_[19793]_ ;
  assign \new_[17539]_  = ~\new_[18108]_ ;
  assign \new_[17540]_  = ~\new_[18704]_  & ~\new_[19788]_ ;
  assign \new_[17541]_  = \new_[18036]_ ;
  assign \new_[17542]_  = ~\new_[18520]_ ;
  assign \new_[17543]_  = ~\new_[18363]_ ;
  assign \new_[17544]_  = ~\new_[18174]_ ;
  assign \new_[17545]_  = ~\new_[19055]_  & ~\new_[21640]_ ;
  assign \new_[17546]_  = ~\new_[18620]_  & ~\new_[19788]_ ;
  assign \new_[17547]_  = ~\new_[18193]_ ;
  assign \new_[17548]_  = ~\new_[18149]_ ;
  assign \new_[17549]_  = \new_[21560]_  & \new_[19170]_ ;
  assign \new_[17550]_  = ~\new_[18450]_ ;
  assign \new_[17551]_  = ~\new_[18372]_ ;
  assign \new_[17552]_  = ~\new_[18624]_  | ~\new_[21506]_ ;
  assign \new_[17553]_  = ~\new_[18464]_ ;
  assign \new_[17554]_  = ~\new_[18694]_  | ~\new_[19095]_ ;
  assign \new_[17555]_  = \new_[15703]_  ^ \new_[1342]_ ;
  assign \new_[17556]_  = ~\new_[18428]_ ;
  assign \new_[17557]_  = ~\new_[18128]_ ;
  assign \new_[17558]_  = ~\new_[18673]_  | ~\new_[19719]_ ;
  assign \new_[17559]_  = ~\new_[18032]_ ;
  assign \new_[17560]_  = ~\new_[18536]_ ;
  assign \new_[17561]_  = ~\new_[18862]_  | ~\new_[21575]_ ;
  assign \new_[17562]_  = \new_[18595]_  | \new_[19655]_ ;
  assign \new_[17563]_  = ~\new_[18041]_ ;
  assign \new_[17564]_  = ~\new_[18526]_ ;
  assign \new_[17565]_  = ~\new_[18127]_ ;
  assign \new_[17566]_  = \new_[18715]_  & \new_[17156]_ ;
  assign \new_[17567]_  = ~\new_[18571]_ ;
  assign n3213 = ~\new_[18715]_  & ~ld;
  assign \new_[17569]_  = ~\new_[18681]_  | ~\new_[19669]_ ;
  assign \new_[17570]_  = \new_[16758]_  ^ \new_[19811]_ ;
  assign \new_[17571]_  = \new_[18883]_  & \new_[21494]_ ;
  assign \new_[17572]_  = \new_[19554]_ ;
  assign \new_[17573]_  = ~\new_[18133]_ ;
  assign \new_[17574]_  = ~\new_[18603]_  & ~\new_[20241]_ ;
  assign \new_[17575]_  = ~\new_[19648]_  & ~\new_[21645]_ ;
  assign \new_[17576]_  = \new_[18890]_  | \new_[19676]_ ;
  assign \new_[17577]_  = ~\new_[18586]_  & ~\new_[18968]_ ;
  assign \new_[17578]_  = ~\new_[19166]_ ;
  assign \new_[17579]_  = ~\new_[18036]_ ;
  assign \new_[17580]_  = ~\new_[21515]_  & ~\new_[18893]_ ;
  assign \new_[17581]_  = ~\new_[18233]_ ;
  assign \new_[17582]_  = ld_r_reg;
  assign \new_[17583]_  = ~\new_[18646]_  | ~\new_[21693]_ ;
  assign \new_[17584]_  = ~\new_[18150]_ ;
  assign \new_[17585]_  = ~\new_[19299]_  & ~\new_[1033]_ ;
  assign \new_[17586]_  = ~\new_[18761]_  & ~\new_[19670]_ ;
  assign \new_[17587]_  = ~\new_[18281]_ ;
  assign \new_[17588]_  = ~\new_[21259]_  & ~\new_[19220]_ ;
  assign \new_[17589]_  = ~\new_[18397]_ ;
  assign \new_[17590]_  = ~\new_[18330]_ ;
  assign \new_[17591]_  = ~\new_[21579]_  & ~\new_[21513]_ ;
  assign \new_[17592]_  = ~\new_[18425]_ ;
  assign \new_[17593]_  = ~\new_[18338]_ ;
  assign \new_[17594]_  = ~\new_[18776]_  & ~\new_[19410]_ ;
  assign \new_[17595]_  = ~\new_[18724]_  & ~\new_[21494]_ ;
  assign \new_[17596]_  = ~\new_[18743]_  & ~\new_[19096]_ ;
  assign \new_[17597]_  = ~\new_[18303]_ ;
  assign \new_[17598]_  = ~\new_[18224]_ ;
  assign \new_[17599]_  = ~\new_[18071]_ ;
  assign \new_[17600]_  = ~\new_[18645]_  & ~\new_[21660]_ ;
  assign \new_[17601]_  = ~\new_[20765]_ ;
  assign \new_[17602]_  = ~\new_[20767]_  | ~\new_[19302]_  | ~\new_[18140]_ ;
  assign \new_[17603]_  = ~\new_[18932]_  & ~\new_[19603]_ ;
  assign \new_[17604]_  = \new_[19726]_  ^ \new_[19175]_ ;
  assign \new_[17605]_  = ~\new_[18735]_  & ~\new_[19603]_ ;
  assign \new_[17606]_  = ~\new_[18302]_ ;
  assign \new_[17607]_  = ~\new_[18485]_ ;
  assign \new_[17608]_  = ~\new_[18056]_ ;
  assign \new_[17609]_  = ~\new_[18165]_ ;
  assign \new_[17610]_  = ~\new_[18628]_  | ~\new_[19412]_ ;
  assign \new_[17611]_  = \new_[18457]_ ;
  assign \new_[17612]_  = \new_[18772]_  | \new_[19033]_ ;
  assign \new_[17613]_  = ~\new_[18107]_ ;
  assign \new_[17614]_  = ~\new_[18247]_ ;
  assign \new_[17615]_  = ~\new_[19695]_  | ~\new_[19281]_ ;
  assign \new_[17616]_  = ~\new_[18601]_  | ~\new_[19186]_ ;
  assign \new_[17617]_  = \new_[18136]_ ;
  assign \new_[17618]_  = ~\new_[20680]_  | ~\new_[19317]_ ;
  assign \new_[17619]_  = ~\new_[18226]_ ;
  assign \new_[17620]_  = \new_[18831]_  & \new_[19589]_ ;
  assign \new_[17621]_  = ~\new_[18389]_ ;
  assign \new_[17622]_  = ~\new_[18053]_ ;
  assign \new_[17623]_  = ~\new_[19174]_  | ~\new_[19729]_ ;
  assign \new_[17624]_  = \new_[19714]_  ^ \new_[19175]_ ;
  assign \new_[17625]_  = ~\new_[18497]_ ;
  assign \new_[17626]_  = ~\new_[18854]_  & ~\new_[18845]_ ;
  assign \new_[17627]_  = ~\new_[18685]_  & ~\new_[21657]_ ;
  assign \new_[17628]_  = ~\new_[19384]_  | ~\new_[19409]_ ;
  assign \new_[17629]_  = ~\new_[19450]_  & ~\new_[1026]_ ;
  assign \new_[17630]_  = ~\new_[18563]_ ;
  assign \new_[17631]_  = ~\new_[18521]_ ;
  assign \new_[17632]_  = ~\new_[18089]_ ;
  assign \new_[17633]_  = ~\new_[18727]_  | ~\new_[19670]_ ;
  assign \new_[17634]_  = ~\new_[18098]_ ;
  assign \new_[17635]_  = ~\new_[18203]_ ;
  assign \new_[17636]_  = ~\new_[18700]_  | ~\new_[19379]_ ;
  assign \new_[17637]_  = ~\new_[18043]_ ;
  assign \new_[17638]_  = ~\new_[18351]_ ;
  assign \new_[17639]_  = ~\new_[18661]_  | ~\new_[19417]_ ;
  assign \new_[17640]_  = ~\new_[18460]_ ;
  assign \new_[17641]_  = ~\new_[18730]_  | ~\new_[19685]_ ;
  assign \new_[17642]_  = \new_[15079]_  ^ \new_[18970]_ ;
  assign \new_[17643]_  = ~\new_[18140]_ ;
  assign \new_[17644]_  = ~\new_[18161]_ ;
  assign \new_[17645]_  = ~\new_[18672]_  & ~\new_[19675]_ ;
  assign \new_[17646]_  = ~\new_[18245]_ ;
  assign \new_[17647]_  = ~\new_[18884]_  | ~\new_[21100]_ ;
  assign \new_[17648]_  = ~\new_[18584]_ ;
  assign \new_[17649]_  = ~\new_[18336]_ ;
  assign \new_[17650]_  = ~\new_[18349]_ ;
  assign \new_[17651]_  = \new_[18404]_ ;
  assign \new_[17652]_  = ~\new_[19624]_  | ~\new_[18623]_ ;
  assign \new_[17653]_  = \new_[16926]_  ^ \new_[1719]_ ;
  assign \new_[17654]_  = ~\new_[19676]_  & ~\new_[18765]_ ;
  assign \new_[17655]_  = ~\new_[18780]_  & ~\new_[19205]_ ;
  assign \new_[17656]_  = ~\new_[18929]_  | ~\new_[19335]_ ;
  assign \new_[17657]_  = ~\new_[18639]_  & ~\new_[20699]_ ;
  assign \new_[17658]_  = ~\new_[18804]_  | ~\new_[18974]_ ;
  assign \new_[17659]_  = ~\new_[18713]_  & ~\new_[21525]_ ;
  assign \new_[17660]_  = ~\new_[18498]_ ;
  assign \new_[17661]_  = \new_[18329]_ ;
  assign \new_[17662]_  = ~\new_[21098]_ ;
  assign \new_[17663]_  = ~\new_[21558]_  & ~\new_[19322]_ ;
  assign \new_[17664]_  = ~\new_[18442]_ ;
  assign \new_[17665]_  = ~\new_[18142]_ ;
  assign \new_[17666]_  = ~\new_[20704]_  | ~\new_[21504]_ ;
  assign \new_[17667]_  = ~\new_[18539]_ ;
  assign \new_[17668]_  = ~\new_[19711]_ ;
  assign \new_[17669]_  = ~\new_[18466]_ ;
  assign \new_[17670]_  = ~\new_[18675]_  | ~\new_[19087]_ ;
  assign \new_[17671]_  = ~\new_[18500]_ ;
  assign \new_[17672]_  = ~\new_[18850]_  | ~\new_[19734]_ ;
  assign \new_[17673]_  = ~\new_[18681]_ ;
  assign \new_[17674]_  = ~\new_[18719]_  & ~\new_[19554]_ ;
  assign \new_[17675]_  = ~\new_[18590]_  | ~\new_[19655]_ ;
  assign \new_[17676]_  = ~\new_[18561]_ ;
  assign \new_[17677]_  = ~\new_[18475]_ ;
  assign \new_[17678]_  = ~\new_[18172]_ ;
  assign \new_[17679]_  = ~\new_[18511]_ ;
  assign \new_[17680]_  = ~\new_[18266]_ ;
  assign \new_[17681]_  = ~n3378;
  assign \new_[17682]_  = ~\new_[18972]_  & ~\new_[18647]_ ;
  assign \new_[17683]_  = ~\new_[19689]_  & ~\new_[18802]_ ;
  assign \new_[17684]_  = ~\new_[18340]_ ;
  assign \new_[17685]_  = ~\new_[18088]_ ;
  assign \new_[17686]_  = ~\new_[18164]_ ;
  assign \new_[17687]_  = ~\new_[20496]_ ;
  assign \new_[17688]_  = ~\new_[18097]_ ;
  assign \new_[17689]_  = ~\new_[19243]_ ;
  assign \new_[17690]_  = ~\new_[18482]_ ;
  assign \new_[17691]_  = \new_[14799]_  ^ \new_[19575]_ ;
  assign \new_[17692]_  = \new_[18721]_  | \new_[19192]_ ;
  assign \new_[17693]_  = ~\new_[18885]_  & ~\new_[18964]_ ;
  assign \new_[17694]_  = ~\new_[19577]_  | ~\new_[21585]_  | ~\new_[19039]_ ;
  assign \new_[17695]_  = ~\new_[18345]_ ;
  assign \new_[17696]_  = ~\new_[21259]_  | ~\new_[19758]_ ;
  assign \new_[17697]_  = ~\new_[18473]_ ;
  assign \new_[17698]_  = ~\new_[18151]_ ;
  assign \new_[17699]_  = ~\new_[18328]_ ;
  assign \new_[17700]_  = ~\new_[18092]_ ;
  assign \new_[17701]_  = ~\new_[18200]_ ;
  assign \new_[17702]_  = ~\new_[18335]_ ;
  assign \new_[17703]_  = ~\new_[18311]_ ;
  assign \new_[17704]_  = \new_[19551]_  ^ \new_[19598]_ ;
  assign \new_[17705]_  = \new_[19097]_  & \new_[18754]_ ;
  assign \new_[17706]_  = ~\new_[18745]_  | ~\new_[20301]_ ;
  assign \new_[17707]_  = \new_[18646]_  | \new_[21688]_ ;
  assign \new_[17708]_  = ~\new_[18900]_  | ~\new_[21046]_ ;
  assign \new_[17709]_  = ~\new_[18356]_ ;
  assign \new_[17710]_  = ~\new_[18191]_ ;
  assign \new_[17711]_  = ~\new_[18593]_  & ~\new_[18810]_ ;
  assign \new_[17712]_  = ~\new_[18294]_ ;
  assign \new_[17713]_  = \new_[14877]_  ^ \new_[1430]_ ;
  assign \new_[17714]_  = ~\new_[18292]_ ;
  assign \new_[17715]_  = ~\new_[18293]_ ;
  assign \new_[17716]_  = ~\new_[18163]_ ;
  assign \new_[17717]_  = ~\new_[18348]_ ;
  assign \new_[17718]_  = ~\new_[18793]_  | ~\new_[19603]_ ;
  assign \new_[17719]_  = ~\new_[18239]_ ;
  assign \new_[17720]_  = \new_[17030]_  ^ \new_[19684]_ ;
  assign \new_[17721]_  = \new_[19811]_  ^ \new_[19563]_ ;
  assign \new_[17722]_  = ~\new_[18236]_ ;
  assign \new_[17723]_  = ~\new_[18393]_ ;
  assign \new_[17724]_  = ~\new_[19348]_  & ~\new_[18746]_ ;
  assign \new_[17725]_  = \new_[14770]_  ^ \new_[19796]_ ;
  assign \new_[17726]_  = ~\new_[18283]_  & ~\new_[19205]_ ;
  assign \new_[17727]_  = ~\new_[20982]_ ;
  assign \new_[17728]_  = ~\new_[18824]_  & ~\new_[18939]_ ;
  assign \new_[17729]_  = ~\new_[18770]_  & ~\new_[19162]_ ;
  assign \new_[17730]_  = ~\new_[18117]_ ;
  assign \new_[17731]_  = ~\new_[21539]_  | ~\new_[21518]_ ;
  assign \new_[17732]_  = \new_[19811]_  ^ \new_[19618]_ ;
  assign \new_[17733]_  = ~\new_[18350]_ ;
  assign \new_[17734]_  = ~\new_[18436]_ ;
  assign \new_[17735]_  = ~\new_[20490]_  | ~\new_[19165]_ ;
  assign \new_[17736]_  = ~\new_[18024]_ ;
  assign \new_[17737]_  = ~\new_[18670]_  & ~\new_[19200]_ ;
  assign \new_[17738]_  = ~\new_[18217]_ ;
  assign \new_[17739]_  = ~\new_[18651]_  | ~\new_[19037]_ ;
  assign \new_[17740]_  = ~\new_[18145]_ ;
  assign \new_[17741]_  = \new_[19739]_  ^ \new_[19630]_ ;
  assign \new_[17742]_  = ~\new_[18827]_  | ~\new_[21506]_ ;
  assign \new_[17743]_  = ~\new_[18254]_ ;
  assign \new_[17744]_  = ~\new_[18582]_ ;
  assign \new_[17745]_  = \new_[19651]_  ^ \new_[19549]_ ;
  assign \new_[17746]_  = ~\new_[18916]_  & ~\new_[19309]_ ;
  assign \new_[17747]_  = ~\new_[18169]_ ;
  assign \new_[17748]_  = ~\new_[18301]_ ;
  assign \new_[17749]_  = \new_[17689]_  & \new_[922]_ ;
  assign \new_[17750]_  = ~\new_[18456]_ ;
  assign \new_[17751]_  = ~\new_[18596]_  & ~\new_[18008]_ ;
  assign \new_[17752]_  = ~\new_[20172]_  & ~\new_[18819]_ ;
  assign \new_[17753]_  = ~\new_[18792]_  & ~\new_[21517]_ ;
  assign \new_[17754]_  = ~\new_[20100]_  | ~\new_[19432]_ ;
  assign \new_[17755]_  = ~\new_[18661]_  | ~\new_[19354]_ ;
  assign \new_[17756]_  = \new_[18871]_  | \new_[19655]_ ;
  assign \new_[17757]_  = \new_[18743]_  | \new_[20927]_ ;
  assign \new_[17758]_  = ~\new_[18540]_ ;
  assign \new_[17759]_  = \new_[14759]_  ^ \new_[1863]_ ;
  assign \new_[17760]_  = ~\new_[19030]_  | ~\new_[18843]_ ;
  assign \new_[17761]_  = ~\new_[18484]_ ;
  assign \new_[17762]_  = ~\new_[18405]_ ;
  assign \new_[17763]_  = ~\new_[18243]_ ;
  assign \new_[17764]_  = ~\new_[18591]_  & ~\new_[19674]_ ;
  assign \new_[17765]_  = ~\new_[18547]_ ;
  assign \new_[17766]_  = ~\new_[18379]_ ;
  assign \new_[17767]_  = ~\new_[18062]_ ;
  assign \new_[17768]_  = ~\new_[18566]_ ;
  assign \new_[17769]_  = ~\new_[21078]_  & ~\new_[21502]_ ;
  assign \new_[17770]_  = \new_[19261]_  & \new_[19659]_ ;
  assign \new_[17771]_  = ~\new_[18353]_ ;
  assign \new_[17772]_  = \new_[18725]_  | \new_[19676]_ ;
  assign \new_[17773]_  = ~\new_[18119]_ ;
  assign \new_[17774]_  = ~\new_[18793]_ ;
  assign \new_[17775]_  = ~\new_[21643]_  | ~\new_[19689]_ ;
  assign \new_[17776]_  = ~\new_[18518]_ ;
  assign \new_[17777]_  = ~\new_[18060]_ ;
  assign \new_[17778]_  = \new_[17013]_  ^ \new_[2297]_ ;
  assign \new_[17779]_  = \new_[15843]_  ^ \new_[19610]_ ;
  assign \new_[17780]_  = ~\new_[18661]_  | ~\new_[19617]_ ;
  assign \new_[17781]_  = \new_[17075]_  ^ \new_[19121]_ ;
  assign \new_[17782]_  = ~\new_[18457]_ ;
  assign \new_[17783]_  = \new_[18217]_ ;
  assign \new_[17784]_  = \new_[15815]_  ^ \new_[19784]_ ;
  assign \new_[17785]_  = ~\new_[18601]_  | ~\new_[19438]_ ;
  assign \new_[17786]_  = ~\new_[21573]_  | ~\new_[19367]_ ;
  assign \new_[17787]_  = ~\new_[18838]_  | ~\new_[19676]_ ;
  assign \new_[17788]_  = ~\new_[18075]_ ;
  assign \new_[17789]_  = ~\new_[19094]_  & ~\new_[959]_ ;
  assign \new_[17790]_  = ~\new_[19245]_  & ~\new_[18616]_ ;
  assign \new_[17791]_  = ~\new_[18370]_ ;
  assign \new_[17792]_  = ~\new_[18545]_ ;
  assign \new_[17793]_  = ~\new_[18458]_ ;
  assign \new_[17794]_  = ~\new_[18669]_  & ~\new_[19721]_ ;
  assign \new_[17795]_  = \new_[18919]_  | \new_[19697]_ ;
  assign \new_[17796]_  = ~\new_[18542]_ ;
  assign \new_[17797]_  = ~\new_[21394]_ ;
  assign \new_[17798]_  = ~\new_[18452]_ ;
  assign \new_[17799]_  = ~\new_[18868]_  & ~\new_[19785]_ ;
  assign \new_[17800]_  = ~\new_[20751]_  & ~\new_[18633]_ ;
  assign \new_[17801]_  = ~\new_[19094]_  & ~\new_[19696]_ ;
  assign \new_[17802]_  = ~\new_[18993]_  | ~\new_[19321]_ ;
  assign \new_[17803]_  = ~\new_[18306]_ ;
  assign \new_[17804]_  = \new_[18159]_ ;
  assign \new_[17805]_  = ~\new_[18717]_  | ~\new_[18939]_ ;
  assign \new_[17806]_  = ~\new_[18902]_  | ~\new_[19654]_ ;
  assign \new_[17807]_  = ~\new_[18102]_ ;
  assign \new_[17808]_  = ~\new_[18960]_  & ~\new_[18774]_ ;
  assign \new_[17809]_  = \new_[19560]_  ^ \new_[19590]_ ;
  assign \new_[17810]_  = \new_[19626]_  ^ \new_[1510]_ ;
  assign \new_[17811]_  = \new_[14773]_  ^ \new_[1507]_ ;
  assign \new_[17812]_  = ~\new_[18278]_ ;
  assign \new_[17813]_  = \new_[15819]_  ^ \new_[2301]_ ;
  assign \new_[17814]_  = \new_[14769]_  ^ \new_[1668]_ ;
  assign \new_[17815]_  = \new_[17004]_  ^ \new_[1637]_ ;
  assign \new_[17816]_  = ~\new_[18648]_  & ~\new_[19379]_ ;
  assign \new_[17817]_  = \new_[14788]_  ^ \new_[18961]_ ;
  assign \new_[17818]_  = ~\new_[18153]_ ;
  assign \new_[17819]_  = \new_[16795]_  ^ \new_[19731]_ ;
  assign \new_[17820]_  = \new_[14909]_  ^ \new_[19710]_ ;
  assign \new_[17821]_  = ~\new_[18229]_ ;
  assign \new_[17822]_  = ~\new_[18838]_  | ~\new_[19603]_ ;
  assign \new_[17823]_  = \new_[19551]_  ^ \new_[19718]_ ;
  assign \new_[17824]_  = \new_[18634]_  | \new_[19538]_ ;
  assign \new_[17825]_  = ~\new_[18476]_ ;
  assign \new_[17826]_  = ~\new_[18623]_  | ~\new_[19412]_ ;
  assign \new_[17827]_  = ~\new_[20769]_  | ~\new_[21483]_ ;
  assign \new_[17828]_  = ~\new_[18090]_ ;
  assign \new_[17829]_  = \new_[14698]_  ^ \new_[19549]_ ;
  assign \new_[17830]_  = ~\new_[18730]_  | ~\new_[19655]_ ;
  assign \new_[17831]_  = ~\new_[18702]_  | ~\new_[19353]_ ;
  assign \new_[17832]_  = ~\new_[18539]_ ;
  assign \new_[17833]_  = \new_[14944]_  ^ \new_[19747]_ ;
  assign \new_[17834]_  = ~\new_[18673]_  | ~\new_[20767]_ ;
  assign \new_[17835]_  = ~\new_[18925]_  & ~\new_[18973]_ ;
  assign \new_[17836]_  = ~\new_[18429]_ ;
  assign \new_[17837]_  = ~\new_[20903]_ ;
  assign \new_[17838]_  = \new_[14696]_  ^ \new_[2300]_ ;
  assign \new_[17839]_  = ~\new_[18510]_ ;
  assign \new_[17840]_  = ~\new_[18530]_ ;
  assign \new_[17841]_  = \new_[19505]_  ^ \new_[19657]_ ;
  assign \new_[17842]_  = ~\new_[18882]_  | ~\new_[20751]_ ;
  assign \new_[17843]_  = \new_[20749]_ ;
  assign \new_[17844]_  = \new_[19784]_  ^ \new_[19774]_ ;
  assign \new_[17845]_  = ~\new_[18358]_ ;
  assign \new_[17846]_  = \new_[17046]_  ^ \new_[1921]_ ;
  assign \new_[17847]_  = \new_[18702]_  & \new_[20927]_ ;
  assign \new_[17848]_  = \new_[18306]_ ;
  assign \new_[17849]_  = \new_[16953]_  ^ \new_[1186]_ ;
  assign \new_[17850]_  = ~\new_[18601]_  | ~\new_[19087]_ ;
  assign \new_[17851]_  = \new_[18863]_  & \new_[921]_ ;
  assign \new_[17852]_  = ~\new_[18472]_ ;
  assign \new_[17853]_  = ~\new_[18683]_  & ~\new_[19444]_ ;
  assign \new_[17854]_  = ~\new_[18718]_  & ~\new_[19285]_ ;
  assign \new_[17855]_  = \new_[18618]_  & \new_[19213]_ ;
  assign \new_[17856]_  = ~\new_[18439]_ ;
  assign \new_[17857]_  = ~\new_[18831]_  | ~\new_[19309]_ ;
  assign \new_[17858]_  = \new_[18690]_  | \new_[19030]_ ;
  assign \new_[17859]_  = ~\new_[18933]_  & ~\new_[18963]_ ;
  assign \new_[17860]_  = ~\new_[18181]_ ;
  assign \new_[17861]_  = ~\new_[19547]_  | ~\new_[19279]_ ;
  assign \new_[17862]_  = ~\new_[18276]_ ;
  assign \new_[17863]_  = ~\new_[18831]_  | ~\new_[19213]_ ;
  assign \new_[17864]_  = ~\new_[18541]_ ;
  assign \new_[17865]_  = ~\new_[21643]_  | ~\new_[19055]_ ;
  assign \new_[17866]_  = ~\new_[18380]_ ;
  assign \new_[17867]_  = ~\new_[18462]_ ;
  assign \new_[17868]_  = ~\new_[18805]_  & ~\new_[19309]_ ;
  assign \new_[17869]_  = ~\new_[18564]_ ;
  assign \new_[17870]_  = ~\new_[18691]_  | ~\new_[19332]_ ;
  assign \new_[17871]_  = ~\new_[18400]_ ;
  assign \new_[17872]_  = ~\new_[18781]_  & ~\new_[19669]_ ;
  assign \new_[17873]_  = ~\new_[18038]_ ;
  assign \new_[17874]_  = ~\new_[19237]_ ;
  assign \new_[17875]_  = ~\new_[18090]_ ;
  assign \new_[17876]_  = ~\new_[18346]_ ;
  assign \new_[17877]_  = ~\new_[18771]_  & ~\new_[19597]_ ;
  assign \new_[17878]_  = ~\new_[18869]_  | ~\new_[19047]_ ;
  assign \new_[17879]_  = ~\new_[18843]_  & ~\new_[19548]_ ;
  assign \new_[17880]_  = \new_[16918]_  ^ \new_[19698]_ ;
  assign \new_[17881]_  = ~\new_[18980]_  | ~\new_[19205]_ ;
  assign \new_[17882]_  = \new_[18923]_  | \new_[19619]_ ;
  assign \new_[17883]_  = \new_[19651]_  ^ \new_[1474]_ ;
  assign \new_[17884]_  = ~\new_[18533]_ ;
  assign \new_[17885]_  = ~\new_[18242]_ ;
  assign \new_[17886]_  = ~\new_[20169]_ ;
  assign \new_[17887]_  = \new_[18613]_  | \new_[19117]_ ;
  assign \new_[17888]_  = ~\new_[18146]_ ;
  assign \new_[17889]_  = \new_[14771]_  ^ \new_[1867]_ ;
  assign \new_[17890]_  = \new_[19684]_  ^ \new_[19662]_ ;
  assign \new_[17891]_  = \new_[15823]_  ^ \new_[1670]_ ;
  assign \new_[17892]_  = \new_[19591]_  ^ \new_[19747]_ ;
  assign \new_[17893]_  = \new_[16723]_  ^ \new_[19651]_ ;
  assign \new_[17894]_  = \new_[14761]_  ^ \new_[1238]_ ;
  assign \new_[17895]_  = \new_[14777]_  ^ \new_[1744]_ ;
  assign \new_[17896]_  = ~\new_[18927]_  | ~\new_[19741]_ ;
  assign \new_[17897]_  = \new_[19287]_  ^ \new_[19731]_ ;
  assign \new_[17898]_  = \new_[16826]_  ^ \new_[19025]_ ;
  assign \new_[17899]_  = \new_[19684]_  ^ \new_[19575]_ ;
  assign \new_[17900]_  = \new_[14701]_  ^ \new_[1506]_ ;
  assign \new_[17901]_  = \new_[17400]_  ^ \new_[19124]_ ;
  assign \new_[17902]_  = \new_[15855]_  ^ \new_[19774]_ ;
  assign \new_[17903]_  = \new_[16967]_  ^ \new_[2293]_ ;
  assign \new_[17904]_  = \new_[14912]_  ^ \new_[19101]_ ;
  assign \new_[17905]_  = \new_[14697]_  ^ \new_[1665]_ ;
  assign \new_[17906]_  = ~\new_[18953]_  | ~\new_[19670]_ ;
  assign \new_[17907]_  = \new_[19658]_  ^ \new_[19796]_ ;
  assign \new_[17908]_  = \new_[19799]_  ^ \new_[1346]_ ;
  assign \new_[17909]_  = ~\new_[18517]_ ;
  assign \new_[17910]_  = \new_[14899]_  ^ \new_[1667]_ ;
  assign \new_[17911]_  = ~\new_[18516]_ ;
  assign \new_[17912]_  = ~\new_[18247]_ ;
  assign \new_[17913]_  = ~\new_[18434]_ ;
  assign \new_[17914]_  = ~\new_[18144]_ ;
  assign \new_[17915]_  = ~\new_[18078]_ ;
  assign \new_[17916]_  = ~\new_[18232]_ ;
  assign \new_[17917]_  = ~\new_[18551]_ ;
  assign \new_[17918]_  = ~\new_[18755]_  | ~\new_[20499]_ ;
  assign \new_[17919]_  = ~\new_[19321]_  & ~\new_[20927]_ ;
  assign \new_[17920]_  = ~\new_[18813]_  & ~\new_[18912]_ ;
  assign \new_[17921]_  = ~\new_[18259]_ ;
  assign \new_[17922]_  = ~\new_[19482]_  & ~\new_[18605]_ ;
  assign \new_[17923]_  = ~\new_[18049]_ ;
  assign \new_[17924]_  = ~\new_[18033]_ ;
  assign \new_[17925]_  = \new_[19625]_  & \new_[923]_ ;
  assign \new_[17926]_  = ~\new_[19499]_  | ~\new_[19145]_ ;
  assign \new_[17927]_  = ~\new_[18304]_ ;
  assign \new_[17928]_  = ~\new_[18823]_  & ~\new_[19132]_ ;
  assign \new_[17929]_  = ~\new_[18201]_ ;
  assign \new_[17930]_  = ~\new_[19647]_  & ~\new_[19474]_ ;
  assign \new_[17931]_  = ~\new_[18353]_ ;
  assign \new_[17932]_  = ~\new_[19510]_  | ~\new_[21168]_ ;
  assign \new_[17933]_  = ~\new_[18782]_  | ~\new_[21582]_ ;
  assign \new_[17934]_  = ~\new_[18478]_ ;
  assign \new_[17935]_  = ~\new_[18740]_  & ~\new_[19082]_ ;
  assign \new_[17936]_  = ~\new_[18141]_ ;
  assign \new_[17937]_  = ~\new_[21048]_ ;
  assign \new_[17938]_  = ~\new_[18331]_ ;
  assign \new_[17939]_  = ~\new_[18101]_ ;
  assign \new_[17940]_  = ~\new_[18494]_ ;
  assign \new_[17941]_  = ~\new_[18509]_ ;
  assign \new_[17942]_  = ~\new_[18410]_ ;
  assign \new_[17943]_  = ~\new_[18491]_ ;
  assign \new_[17944]_  = ~\new_[18106]_ ;
  assign \new_[17945]_  = ~\new_[18634]_  | ~\new_[20748]_ ;
  assign \new_[17946]_  = \new_[21396]_  | \new_[21491]_ ;
  assign \new_[17947]_  = ~\new_[21395]_  | ~\new_[19664]_ ;
  assign \new_[17948]_  = ~\new_[18529]_ ;
  assign \new_[17949]_  = ~\new_[18277]_ ;
  assign \new_[17950]_  = ~\new_[18055]_ ;
  assign \new_[17951]_  = ~\new_[18309]_ ;
  assign \new_[17952]_  = ~\new_[18216]_ ;
  assign \new_[17953]_  = ~\new_[21303]_  | ~\new_[21660]_ ;
  assign \new_[17954]_  = ~\new_[18208]_ ;
  assign \new_[17955]_  = ~\new_[18195]_ ;
  assign \new_[17956]_  = \new_[18030]_ ;
  assign \new_[17957]_  = ~\new_[18160]_ ;
  assign \new_[17958]_  = ~\new_[19522]_  | ~\new_[19055]_ ;
  assign \new_[17959]_  = ~\new_[18194]_  | ~\new_[18908]_ ;
  assign \new_[17960]_  = ~\new_[19243]_ ;
  assign \new_[17961]_  = ~\new_[18591]_  | ~\new_[19132]_ ;
  assign \new_[17962]_  = ~\new_[18546]_ ;
  assign \new_[17963]_  = ~\new_[18367]_ ;
  assign \new_[17964]_  = ~\new_[18269]_ ;
  assign \new_[17965]_  = ~\new_[18256]_ ;
  assign \new_[17966]_  = ~\new_[18313]_ ;
  assign \new_[17967]_  = ~\new_[18252]_ ;
  assign \new_[17968]_  = ~\new_[18547]_ ;
  assign \new_[17969]_  = ~\new_[18817]_  | ~\new_[19399]_ ;
  assign \new_[17970]_  = ~\new_[21534]_  | ~\new_[21517]_ ;
  assign \new_[17971]_  = \new_[19353]_  & \new_[19050]_ ;
  assign \new_[17972]_  = ~\new_[18153]_ ;
  assign \new_[17973]_  = ~\new_[18081]_ ;
  assign \new_[17974]_  = ~\new_[18116]_ ;
  assign \new_[17975]_  = ~\new_[20665]_ ;
  assign \new_[17976]_  = \new_[18841]_  | \new_[19754]_ ;
  assign \new_[17977]_  = ~\new_[14951]_  & ~\new_[923]_ ;
  assign \new_[17978]_  = ~\new_[18479]_ ;
  assign \new_[17979]_  = ~\new_[19499]_ ;
  assign \new_[17980]_  = ~\new_[18585]_ ;
  assign \new_[17981]_  = ~\new_[18352]_ ;
  assign \new_[17982]_  = ~\new_[18881]_  & ~\new_[18678]_ ;
  assign \new_[17983]_  = ~\new_[18326]_ ;
  assign \new_[17984]_  = ~\new_[18493]_ ;
  assign \new_[17985]_  = ~\new_[18085]_ ;
  assign \new_[17986]_  = ~\new_[18176]_ ;
  assign \new_[17987]_  = ~\new_[18129]_ ;
  assign \new_[17988]_  = ~\new_[18339]_ ;
  assign \new_[17989]_  = \new_[1513]_  ^ \new_[19340]_ ;
  assign \new_[17990]_  = ~\new_[18610]_  & ~\new_[19438]_ ;
  assign \new_[17991]_  = ~\new_[18138]_ ;
  assign \new_[17992]_  = ~\new_[18560]_ ;
  assign \new_[17993]_  = ~\new_[18231]_ ;
  assign \new_[17994]_  = ~\new_[19412]_  & ~\new_[18889]_ ;
  assign \new_[17995]_  = ~\new_[18377]_ ;
  assign \new_[17996]_  = ~\new_[18154]_ ;
  assign \new_[17997]_  = ~\new_[18886]_  | ~\new_[18974]_ ;
  assign \new_[17998]_  = ~\new_[18210]_ ;
  assign \new_[17999]_  = ~\new_[18617]_  & ~\new_[19026]_ ;
  assign \new_[18000]_  = ~\new_[18604]_  & ~\new_[19200]_ ;
  assign \new_[18001]_  = ~\new_[18968]_  | ~\new_[21513]_ ;
  assign \new_[18002]_  = ~\new_[18857]_  | ~\new_[18845]_ ;
  assign \new_[18003]_  = \new_[18600]_  & \new_[19438]_ ;
  assign \new_[18004]_  = ~\new_[19322]_ ;
  assign \new_[18005]_  = ~\new_[18219]_ ;
  assign \new_[18006]_  = ~\new_[18542]_  | ~\new_[19460]_ ;
  assign \new_[18007]_  = ~\new_[18168]_ ;
  assign \new_[18008]_  = ~\new_[19794]_ ;
  assign \new_[18009]_  = ~\new_[18264]_ ;
  assign \new_[18010]_  = ~\new_[19301]_  & ~\new_[19308]_ ;
  assign \new_[18011]_  = ~\new_[19156]_ ;
  assign \new_[18012]_  = ~\new_[19362]_ ;
  assign \new_[18013]_  = ~\new_[18287]_ ;
  assign \new_[18014]_  = ~\new_[18523]_ ;
  assign \new_[18015]_  = ~\new_[18314]_ ;
  assign \new_[18016]_  = ~\new_[18688]_  | ~\new_[20751]_ ;
  assign \new_[18017]_  = ~\new_[19149]_ ;
  assign \new_[18018]_  = \new_[18671]_  | \new_[19213]_ ;
  assign \new_[18019]_  = ~\new_[18579]_ ;
  assign \new_[18020]_  = ~\new_[18141]_ ;
  assign \new_[18021]_  = ~\new_[21115]_  & ~\new_[922]_ ;
  assign \new_[18022]_  = ~\new_[19531]_  | ~\new_[19024]_ ;
  assign \new_[18023]_  = ~\new_[18901]_ ;
  assign \new_[18024]_  = ~\new_[18781]_ ;
  assign \new_[18025]_  = ~\new_[18741]_ ;
  assign \new_[18026]_  = ~\new_[18740]_ ;
  assign n3388 = \new_[17302]_  ? \new_[19472]_  : \text_in[5] ;
  assign \new_[18028]_  = \new_[19210]_  & \new_[20865]_ ;
  assign n3273 = \new_[16801]_  ? \new_[19372]_  : \text_in[50] ;
  assign \new_[18030]_  = ~\new_[21100]_  & ~\new_[18951]_ ;
  assign \new_[18031]_  = ~\new_[19687]_  & ~\new_[19791]_ ;
  assign \new_[18032]_  = ~\new_[21115]_  | ~\new_[18605]_ ;
  assign \new_[18033]_  = ~\new_[19727]_  | ~\new_[1928]_ ;
  assign \new_[18034]_  = ~\new_[18710]_ ;
  assign \new_[18035]_  = ~\new_[18603]_ ;
  assign \new_[18036]_  = ~\new_[18653]_ ;
  assign \new_[18037]_  = \new_[20704]_  & \new_[21513]_ ;
  assign \new_[18038]_  = ~\new_[19111]_  | ~\new_[19412]_ ;
  assign \new_[18039]_  = \new_[14702]_  ^ \new_[1353]_ ;
  assign \new_[18040]_  = \new_[19768]_  ^ \new_[19562]_ ;
  assign \new_[18041]_  = ~\new_[19134]_  | ~\new_[19743]_ ;
  assign \new_[18042]_  = \new_[14962]_  ^ \new_[1661]_ ;
  assign \new_[18043]_  = ~\new_[19174]_  & ~\new_[18963]_ ;
  assign \new_[18044]_  = \new_[14755]_  ^ \new_[1291]_ ;
  assign \new_[18045]_  = ~\new_[18628]_ ;
  assign \new_[18046]_  = ~\new_[18827]_ ;
  assign n3223 = \new_[16692]_  ? \new_[19414]_  : \text_in[2] ;
  assign \new_[18048]_  = ~\new_[18869]_ ;
  assign \new_[18049]_  = ~\new_[18899]_ ;
  assign \new_[18050]_  = ~\new_[18871]_ ;
  assign \new_[18051]_  = ~\new_[19065]_  | ~\new_[21494]_ ;
  assign n3318 = \new_[16995]_  ? ld : \text_in[31] ;
  assign \new_[18053]_  = ~\new_[19302]_  | ~\new_[19055]_ ;
  assign \new_[18054]_  = ~\new_[18862]_ ;
  assign \new_[18055]_  = ~\new_[18645]_ ;
  assign \new_[18056]_  = \new_[18673]_ ;
  assign \new_[18057]_  = \new_[19720]_  ^ \new_[19733]_ ;
  assign \new_[18058]_  = \new_[17053]_  ^ \new_[19658]_ ;
  assign \new_[18059]_  = ~\new_[19355]_  | ~\new_[18699]_ ;
  assign \new_[18060]_  = ~\new_[18842]_ ;
  assign \new_[18061]_  = ~\new_[18854]_ ;
  assign \new_[18062]_  = ~\new_[18825]_ ;
  assign \new_[18063]_  = ~\new_[19507]_  | ~\new_[19117]_ ;
  assign \new_[18064]_  = \new_[14943]_  ^ \new_[1518]_ ;
  assign \new_[18065]_  = ~\new_[19712]_  | ~\new_[21523]_ ;
  assign \new_[18066]_  = ~\new_[18643]_ ;
  assign \new_[18067]_  = ~\new_[18771]_ ;
  assign \new_[18068]_  = ~\new_[18647]_ ;
  assign \new_[18069]_  = \new_[19301]_  & \new_[19771]_ ;
  assign \new_[18070]_  = ~\new_[19798]_ ;
  assign \new_[18071]_  = ~\new_[19060]_  | ~\new_[20751]_ ;
  assign n3363 = \new_[17116]_  ? \new_[19383]_  : \text_in[27] ;
  assign \new_[18073]_  = \new_[19814]_  ^ \new_[19565]_ ;
  assign \new_[18074]_  = \new_[16801]_  ^ \new_[1658]_ ;
  assign \new_[18075]_  = ~\new_[19004]_  | ~\new_[19582]_ ;
  assign \new_[18076]_  = ~\new_[19508]_ ;
  assign \new_[18077]_  = ~\new_[18769]_ ;
  assign \new_[18078]_  = ~\new_[18944]_  & ~\new_[19754]_ ;
  assign \new_[18079]_  = ~\new_[18626]_ ;
  assign \new_[18080]_  = ~\new_[20768]_ ;
  assign \new_[18081]_  = ~\new_[19201]_  & ~\new_[19030]_ ;
  assign \new_[18082]_  = ~\new_[18812]_ ;
  assign \new_[18083]_  = ~\new_[21258]_ ;
  assign \new_[18084]_  = \new_[19240]_  | \new_[19694]_ ;
  assign \new_[18085]_  = ~\new_[18670]_ ;
  assign \new_[18086]_  = ~\new_[18731]_ ;
  assign \new_[18087]_  = ~\new_[20842]_ ;
  assign \new_[18088]_  = ~\new_[18730]_ ;
  assign \new_[18089]_  = ~\new_[19172]_  & ~\new_[19622]_ ;
  assign \new_[18090]_  = ~\new_[19183]_  | ~\new_[19010]_ ;
  assign \new_[18091]_  = ~\new_[19659]_ ;
  assign \new_[18092]_  = ~\new_[19065]_  & ~\new_[21494]_ ;
  assign \new_[18093]_  = ~\new_[19210]_  & ~\new_[20865]_ ;
  assign \new_[18094]_  = ~\new_[18823]_ ;
  assign \new_[18095]_  = ~\new_[19218]_  | ~\new_[19417]_ ;
  assign \new_[18096]_  = ~\new_[19047]_ ;
  assign \new_[18097]_  = ~\new_[19366]_  & ~\new_[19717]_ ;
  assign \new_[18098]_  = \new_[19267]_  & \new_[21657]_ ;
  assign \new_[18099]_  = \new_[14768]_  ^ \new_[1424]_ ;
  assign \new_[18100]_  = ~\new_[18704]_ ;
  assign \new_[18101]_  = ~\new_[21115]_  | ~\new_[19106]_ ;
  assign \new_[18102]_  = ~\new_[19019]_  | ~\new_[21166]_ ;
  assign \new_[18103]_  = ~\new_[18717]_ ;
  assign \new_[18104]_  = ~\new_[18698]_ ;
  assign \new_[18105]_  = \new_[19760]_  ^ \new_[19716]_ ;
  assign \new_[18106]_  = ~\new_[20681]_  | ~\new_[20239]_ ;
  assign \new_[18107]_  = ~\new_[21494]_  & ~\new_[19227]_ ;
  assign \new_[18108]_  = \new_[18900]_ ;
  assign \new_[18109]_  = \new_[19345]_  ^ \new_[19753]_ ;
  assign \new_[18110]_  = ~\new_[21580]_  & ~\new_[21511]_ ;
  assign \new_[18111]_  = ~\new_[18714]_ ;
  assign \new_[18112]_  = ~\new_[19035]_  & ~\new_[19758]_ ;
  assign \new_[18113]_  = \new_[15851]_  ^ \new_[19515]_ ;
  assign n3258 = \new_[16758]_  ? \new_[19451]_  : \text_in[112] ;
  assign \new_[18115]_  = ~\new_[19481]_  & ~\new_[17979]_ ;
  assign \new_[18116]_  = \new_[21397]_  | \new_[19681]_ ;
  assign \new_[18117]_  = ~\new_[19349]_  | ~\new_[19082]_ ;
  assign \new_[18118]_  = ~\new_[18673]_ ;
  assign \new_[18119]_  = ~\new_[18885]_ ;
  assign \new_[18120]_  = ~\new_[21388]_ ;
  assign \new_[18121]_  = ~\new_[18927]_ ;
  assign \new_[18122]_  = ~\new_[18890]_ ;
  assign \new_[18123]_  = ~\new_[19228]_ ;
  assign \new_[18124]_  = ~\new_[17796]_ ;
  assign n3288 = \new_[16854]_  ? \new_[19383]_  : \text_in[25] ;
  assign \new_[18126]_  = ~\new_[18656]_ ;
  assign \new_[18127]_  = ~\new_[18586]_ ;
  assign \new_[18128]_  = \new_[19503]_  | \new_[19211]_ ;
  assign \new_[18129]_  = \new_[20166]_  & \new_[19596]_ ;
  assign \new_[18130]_  = ~\new_[18700]_ ;
  assign \new_[18131]_  = ~\new_[18792]_ ;
  assign \new_[18132]_  = ~\new_[18759]_ ;
  assign \new_[18133]_  = ~\new_[19419]_  & ~\new_[19738]_ ;
  assign \new_[18134]_  = ~\new_[18806]_ ;
  assign \new_[18135]_  = \new_[19810]_  ^ \new_[1619]_ ;
  assign \new_[18136]_  = ~\new_[19062]_  | ~\new_[21540]_ ;
  assign \new_[18137]_  = ~\new_[18795]_ ;
  assign \new_[18138]_  = \new_[20490]_  | \new_[18605]_ ;
  assign \new_[18139]_  = ~\new_[18925]_ ;
  assign \new_[18140]_  = ~\new_[19522]_ ;
  assign \new_[18141]_  = ~\new_[19226]_  | ~\new_[19464]_ ;
  assign \new_[18142]_  = ~\new_[18718]_ ;
  assign \new_[18143]_  = \new_[14750]_  ^ \new_[1419]_ ;
  assign \new_[18144]_  = ~\new_[19078]_  & ~\new_[19685]_ ;
  assign \new_[18145]_  = ~\new_[19140]_  | ~\new_[19395]_ ;
  assign \new_[18146]_  = ~\new_[18697]_ ;
  assign n3408 = \new_[17430]_  ? \new_[19372]_  : \text_in[71] ;
  assign \new_[18148]_  = \new_[18720]_ ;
  assign \new_[18149]_  = \new_[18884]_ ;
  assign \new_[18150]_  = ~\new_[18932]_ ;
  assign \new_[18151]_  = ~\new_[18654]_ ;
  assign n3308 = \new_[16953]_  ? \new_[19479]_  : \text_in[115] ;
  assign \new_[18153]_  = \new_[20487]_  | \new_[21115]_ ;
  assign \new_[18154]_  = ~\new_[21115]_  & ~\new_[19337]_ ;
  assign \new_[18155]_  = \new_[14790]_  ^ \new_[1240]_ ;
  assign \new_[18156]_  = \new_[19090]_  | \new_[19738]_ ;
  assign \new_[18157]_  = ~\new_[18875]_ ;
  assign \new_[18158]_  = \new_[14725]_  ^ \new_[1348]_ ;
  assign \new_[18159]_  = ~\new_[18950]_  | ~\new_[18951]_ ;
  assign \new_[18160]_  = ~\new_[20771]_ ;
  assign \new_[18161]_  = ~\new_[18916]_ ;
  assign n3218 = \new_[16684]_  ? \new_[19414]_  : \text_in[125] ;
  assign \new_[18163]_  = ~\new_[18768]_ ;
  assign \new_[18164]_  = ~\new_[18688]_ ;
  assign \new_[18165]_  = ~\new_[19227]_  | ~\new_[21489]_ ;
  assign \new_[18166]_  = ~\new_[19281]_ ;
  assign \new_[18167]_  = ~\new_[18936]_ ;
  assign \new_[18168]_  = ~\new_[18989]_  & ~\new_[20751]_ ;
  assign \new_[18169]_  = ~\new_[18669]_ ;
  assign \new_[18170]_  = ~\new_[18864]_ ;
  assign \new_[18171]_  = ~\new_[18752]_ ;
  assign \new_[18172]_  = ~\new_[18911]_ ;
  assign \new_[18173]_  = ~\new_[18722]_ ;
  assign \new_[18174]_  = ~\new_[19381]_  | ~\new_[21696]_ ;
  assign \new_[18175]_  = ~\new_[18744]_ ;
  assign \new_[18176]_  = ~\new_[20037]_ ;
  assign \new_[18177]_  = ~\new_[18774]_ ;
  assign \new_[18178]_  = \new_[16743]_  ^ \new_[1663]_ ;
  assign \new_[18179]_  = ~\new_[19373]_ ;
  assign \new_[18180]_  = ~\new_[18708]_ ;
  assign \new_[18181]_  = ~\new_[19250]_  | ~\new_[19675]_ ;
  assign \new_[18182]_  = ~\new_[18598]_ ;
  assign \new_[18183]_  = ~\new_[18861]_ ;
  assign \new_[18184]_  = ~\new_[18914]_ ;
  assign \new_[18185]_  = \new_[15846]_  ^ \new_[1509]_ ;
  assign \new_[18186]_  = ~\new_[18802]_ ;
  assign \new_[18187]_  = ~\new_[19507]_ ;
  assign \new_[18188]_  = \new_[19776]_  ^ \new_[19666]_ ;
  assign \new_[18189]_  = ~\new_[18987]_  & ~\new_[19245]_ ;
  assign \new_[18190]_  = ~\new_[18695]_ ;
  assign \new_[18191]_  = ~\new_[19390]_  | ~\new_[19754]_ ;
  assign \new_[18192]_  = ~\new_[18816]_ ;
  assign \new_[18193]_  = ~\new_[18140]_  | ~\new_[20301]_ ;
  assign \new_[18194]_  = ~\new_[19508]_ ;
  assign \new_[18195]_  = ~\new_[18868]_ ;
  assign \new_[18196]_  = ~\new_[18671]_ ;
  assign \new_[18197]_  = ~\new_[18705]_ ;
  assign \new_[18198]_  = ~\new_[18895]_ ;
  assign \new_[18199]_  = ~\new_[18664]_ ;
  assign \new_[18200]_  = ~\new_[19039]_  | ~\new_[21583]_ ;
  assign \new_[18201]_  = ~\new_[21573]_  & ~\new_[19151]_ ;
  assign n3278 = \new_[16826]_  ? ld : \text_in[100] ;
  assign \new_[18203]_  = ~\new_[18705]_ ;
  assign \new_[18204]_  = ~\new_[19140]_  & ~\new_[20172]_ ;
  assign \new_[18205]_  = \new_[19632]_  ^ \new_[19673]_ ;
  assign \new_[18206]_  = ~\new_[18721]_ ;
  assign \new_[18207]_  = \new_[19749]_  ^ \new_[19720]_ ;
  assign \new_[18208]_  = ~\new_[19519]_  | ~\new_[20865]_ ;
  assign \new_[18209]_  = ~\new_[19520]_ ;
  assign \new_[18210]_  = ~\new_[19191]_  & ~\new_[21049]_ ;
  assign \new_[18211]_  = ~\new_[19238]_  | ~\new_[19464]_ ;
  assign \new_[18212]_  = \new_[19631]_  ^ \new_[19287]_ ;
  assign n3243 = \new_[16743]_  ? \new_[19414]_  : \text_in[106] ;
  assign \new_[18214]_  = \new_[15756]_  ^ \new_[19287]_ ;
  assign \new_[18215]_  = \new_[15861]_  ^ \new_[19735]_ ;
  assign \new_[18216]_  = ~\new_[21534]_  | ~\new_[21516]_ ;
  assign \new_[18217]_  = ~\new_[18800]_ ;
  assign \new_[18218]_  = ~\new_[21478]_ ;
  assign \new_[18219]_  = \new_[19165]_  & \new_[21517]_ ;
  assign \new_[18220]_  = \new_[15068]_  ^ \new_[19792]_ ;
  assign \new_[18221]_  = \new_[1513]_  ^ \new_[19686]_ ;
  assign \new_[18222]_  = ~\new_[18753]_ ;
  assign \new_[18223]_  = \new_[19676]_  & \new_[19090]_ ;
  assign \new_[18224]_  = ~\new_[18008]_ ;
  assign n3328 = \new_[17013]_  ? \new_[19338]_  : \text_in[119] ;
  assign \new_[18226]_  = ~\new_[18774]_ ;
  assign \new_[18227]_  = ~\new_[18702]_ ;
  assign \new_[18228]_  = ~\new_[19388]_ ;
  assign \new_[18229]_  = ~\new_[18642]_ ;
  assign \new_[18230]_  = ~\new_[18991]_  | ~\new_[18939]_ ;
  assign \new_[18231]_  = \new_[18947]_  & \new_[20492]_ ;
  assign \new_[18232]_  = ~\new_[19764]_  | ~\new_[19660]_ ;
  assign \new_[18233]_  = ~\new_[19525]_  | ~\new_[19052]_ ;
  assign \new_[18234]_  = \new_[19174]_  | \new_[19674]_ ;
  assign \new_[18235]_  = ~\new_[18797]_ ;
  assign \new_[18236]_  = ~\new_[19016]_  & ~\new_[19213]_ ;
  assign \new_[18237]_  = \new_[18992]_  | \new_[19659]_ ;
  assign \new_[18238]_  = ~\new_[18831]_ ;
  assign \new_[18239]_  = ~\new_[19216]_  | ~\new_[19435]_ ;
  assign \new_[18240]_  = \new_[19735]_  ^ \new_[19505]_ ;
  assign \new_[18241]_  = ~\new_[18591]_ ;
  assign \new_[18242]_  = ~\new_[21303]_  | ~\new_[21656]_ ;
  assign \new_[18243]_  = ~\new_[18872]_ ;
  assign \new_[18244]_  = ~\new_[18591]_ ;
  assign \new_[18245]_  = ~\new_[19221]_  & ~\new_[19603]_ ;
  assign \new_[18246]_  = ~\new_[18728]_ ;
  assign \new_[18247]_  = ~\new_[21540]_  | ~\new_[21523]_ ;
  assign \new_[18248]_  = ~\new_[18738]_ ;
  assign \new_[18249]_  = \new_[19727]_  | \new_[19550]_ ;
  assign \new_[18250]_  = ~\new_[18636]_ ;
  assign \new_[18251]_  = ~\new_[18687]_ ;
  assign \new_[18252]_  = \new_[18140]_  | \new_[19689]_ ;
  assign \new_[18253]_  = ~\new_[18735]_ ;
  assign \new_[18254]_  = ~\new_[19330]_  & ~\new_[21581]_ ;
  assign \new_[18255]_  = ~\new_[18645]_ ;
  assign \new_[18256]_  = ~\new_[18719]_ ;
  assign \new_[18257]_  = \new_[19280]_  ^ \new_[19606]_ ;
  assign n3338 = \new_[17046]_  ? \new_[19451]_  : \text_in[76] ;
  assign \new_[18259]_  = ~\new_[18648]_ ;
  assign \new_[18260]_  = \new_[14753]_  ^ \new_[1427]_ ;
  assign \new_[18261]_  = ~\new_[18633]_ ;
  assign \new_[18262]_  = ~\new_[18631]_ ;
  assign \new_[18263]_  = ~\new_[18670]_ ;
  assign \new_[18264]_  = \new_[18867]_ ;
  assign n3418 = \new_[17448]_  ? ld : \text_in[87] ;
  assign \new_[18266]_  = ~\new_[18805]_ ;
  assign n3313 = \new_[16967]_  ? ld : \text_in[98] ;
  assign n3373 = \new_[17148]_  ? \new_[19479]_  : \text_in[117] ;
  assign \new_[18269]_  = ~\new_[19234]_  | ~\new_[19353]_ ;
  assign \new_[18270]_  = ~\new_[18588]_ ;
  assign \new_[18271]_  = ~\new_[18727]_ ;
  assign n3378 = ~\new_[17156]_  & ~ld;
  assign \new_[18273]_  = ~\new_[18592]_ ;
  assign \new_[18274]_  = ~\new_[18629]_ ;
  assign \new_[18275]_  = ~\new_[18940]_  & ~\new_[19181]_ ;
  assign \new_[18276]_  = ~\new_[19401]_  & ~\new_[18974]_ ;
  assign \new_[18277]_  = \new_[21543]_  & \new_[21521]_ ;
  assign \new_[18278]_  = ~\new_[21638]_  & ~\new_[19050]_ ;
  assign \new_[18279]_  = ~\new_[21522]_  & ~\new_[21543]_ ;
  assign \new_[18280]_  = ~\new_[18739]_ ;
  assign \new_[18281]_  = ~\new_[21644]_ ;
  assign \new_[18282]_  = ~\new_[19093]_  | ~\new_[20751]_ ;
  assign \new_[18283]_  = ~\new_[18980]_ ;
  assign \new_[18284]_  = ~\new_[18683]_ ;
  assign \new_[18285]_  = ~\new_[19423]_ ;
  assign \new_[18286]_  = \new_[16754]_  ^ \new_[1241]_ ;
  assign \new_[18287]_  = ~\new_[18976]_  | ~\new_[19274]_ ;
  assign \new_[18288]_  = ~\new_[19519]_ ;
  assign \new_[18289]_  = \new_[15840]_  ^ \new_[1352]_ ;
  assign n3398 = \new_[17400]_  ? \new_[19451]_  : \text_in[83] ;
  assign n3353 = \new_[17087]_  ? ld : \text_in[62] ;
  assign \new_[18292]_  = \new_[19059]_  | \new_[19770]_ ;
  assign \new_[18293]_  = ~\new_[18895]_ ;
  assign \new_[18294]_  = ~\new_[18736]_ ;
  assign \new_[18295]_  = \new_[14719]_  ^ \new_[2079]_ ;
  assign \new_[18296]_  = \new_[19571]_  ^ \new_[19805]_ ;
  assign \new_[18297]_  = ~\new_[18613]_ ;
  assign n3303 = \new_[16926]_  ? \new_[19414]_  : \text_in[124] ;
  assign \new_[18299]_  = ~\new_[18600]_ ;
  assign \new_[18300]_  = ~\new_[19587]_  & ~\new_[984]_ ;
  assign \new_[18301]_  = ~\new_[18675]_ ;
  assign \new_[18302]_  = ~\new_[19089]_  | ~\new_[19680]_ ;
  assign \new_[18303]_  = ~\new_[19090]_  | ~\new_[18699]_ ;
  assign \new_[18304]_  = \new_[19742]_  & \new_[1879]_ ;
  assign \new_[18305]_  = \new_[1348]_  ^ \new_[1663]_ ;
  assign \new_[18306]_  = ~\new_[19191]_  | ~\new_[19209]_ ;
  assign \new_[18307]_  = ~\new_[18715]_ ;
  assign \new_[18308]_  = ~\new_[18788]_ ;
  assign \new_[18309]_  = ~\new_[19174]_  | ~\new_[19146]_ ;
  assign \new_[18310]_  = ~\new_[18725]_ ;
  assign \new_[18311]_  = ~\new_[19147]_  & ~\new_[19650]_ ;
  assign \new_[18312]_  = ~\new_[18800]_ ;
  assign \new_[18313]_  = \new_[19503]_  & \new_[19087]_ ;
  assign \new_[18314]_  = ~\new_[18593]_ ;
  assign n3253 = \new_[16754]_  ? ld : \text_in[43] ;
  assign \new_[18316]_  = \new_[19184]_  | \new_[19665]_ ;
  assign \new_[18317]_  = ~\new_[20591]_ ;
  assign n3233 = \new_[16715]_  ? \new_[19472]_  : \text_in[72] ;
  assign \new_[18319]_  = ~\new_[18796]_ ;
  assign \new_[18320]_  = \new_[14722]_  ^ \new_[19704]_ ;
  assign \new_[18321]_  = \new_[14781]_  ^ \new_[1620]_ ;
  assign \new_[18322]_  = ~\new_[18711]_ ;
  assign \new_[18323]_  = ~\new_[18931]_ ;
  assign n3358 = \new_[17091]_  ? \new_[19372]_  : \text_in[48] ;
  assign \new_[18325]_  = ~\new_[19358]_ ;
  assign \new_[18326]_  = \new_[20681]_  | \new_[20241]_ ;
  assign \new_[18327]_  = ~\new_[21303]_ ;
  assign \new_[18328]_  = ~\new_[19122]_  & ~\new_[21685]_ ;
  assign \new_[18329]_  = ~\new_[18726]_ ;
  assign \new_[18330]_  = \new_[19231]_  & \new_[19734]_ ;
  assign \new_[18331]_  = ~\new_[19680]_  | ~\new_[19788]_ ;
  assign \new_[18332]_  = \new_[19815]_  & \new_[19697]_ ;
  assign n3248 = \new_[16752]_  ? \new_[19383]_  : \text_in[4] ;
  assign \new_[18334]_  = \new_[19805]_  ^ \new_[1187]_ ;
  assign \new_[18335]_  = ~\new_[20100]_  | ~\new_[18979]_ ;
  assign \new_[18336]_  = ~\new_[21477]_ ;
  assign \new_[18337]_  = ~\new_[18694]_ ;
  assign \new_[18338]_  = ~\new_[21303]_  & ~\new_[21657]_ ;
  assign \new_[18339]_  = ~\new_[18819]_ ;
  assign \new_[18340]_  = ~\new_[18638]_ ;
  assign \new_[18341]_  = \new_[19021]_  & \new_[1025]_ ;
  assign \new_[18342]_  = \new_[19793]_  ^ \new_[19732]_ ;
  assign \new_[18343]_  = \new_[17448]_  ^ \new_[2511]_ ;
  assign \new_[18344]_  = \new_[19015]_  & \new_[1039]_ ;
  assign \new_[18345]_  = ~\new_[18690]_ ;
  assign \new_[18346]_  = ~\new_[19235]_  & ~\new_[19669]_ ;
  assign \new_[18347]_  = \new_[19142]_  | \new_[19425]_ ;
  assign \new_[18348]_  = ~\new_[19135]_  | ~\new_[18968]_ ;
  assign \new_[18349]_  = ~\new_[18999]_  | ~\new_[19603]_ ;
  assign \new_[18350]_  = ~\new_[18716]_ ;
  assign \new_[18351]_  = ~\new_[18824]_ ;
  assign \new_[18352]_  = ~\new_[18742]_ ;
  assign \new_[18353]_  = ~\new_[18780]_ ;
  assign \new_[18354]_  = \new_[19560]_  ^ \new_[19737]_ ;
  assign \new_[18355]_  = ~\new_[18790]_ ;
  assign \new_[18356]_  = ~\new_[19069]_  | ~\new_[21097]_ ;
  assign n3293 = \new_[16892]_  ? ld : \text_in[57] ;
  assign \new_[18358]_  = \new_[19381]_  | \new_[21688]_ ;
  assign \new_[18359]_  = \new_[14960]_  ^ \new_[19760]_ ;
  assign \new_[18360]_  = \new_[15634]_  ^ \new_[2288]_ ;
  assign \new_[18361]_  = ~\new_[18827]_ ;
  assign \new_[18362]_  = ~\new_[18982]_ ;
  assign \new_[18363]_  = ~\new_[19248]_  & ~\new_[19213]_ ;
  assign n3348 = \new_[17075]_  ? ld : \text_in[94] ;
  assign \new_[18365]_  = ~\new_[18837]_ ;
  assign \new_[18366]_  = \new_[17125]_  ^ \new_[19716]_ ;
  assign \new_[18367]_  = ~\new_[19670]_  & ~\new_[19080]_ ;
  assign \new_[18368]_  = ~\new_[18870]_ ;
  assign \new_[18369]_  = ~\new_[18626]_ ;
  assign \new_[18370]_  = ~\new_[19293]_  & ~\new_[19758]_ ;
  assign \new_[18371]_  = ~\new_[18776]_ ;
  assign \new_[18372]_  = ~\new_[17796]_  | ~\new_[19084]_ ;
  assign \new_[18373]_  = \new_[19727]_  | \new_[1928]_ ;
  assign \new_[18374]_  = ~\new_[18838]_ ;
  assign \new_[18375]_  = ~\new_[18870]_ ;
  assign \new_[18376]_  = ~\new_[18878]_ ;
  assign \new_[18377]_  = ~\new_[19058]_  & ~\new_[20751]_ ;
  assign \new_[18378]_  = ~\new_[18877]_ ;
  assign \new_[18379]_  = \new_[19174]_  & \new_[19020]_ ;
  assign \new_[18380]_  = ~\new_[19625]_  & ~\new_[19277]_ ;
  assign \new_[18381]_  = ~\new_[18768]_ ;
  assign \new_[18382]_  = ~\new_[18920]_ ;
  assign n3368 = \new_[17125]_  ? \new_[19338]_  : \text_in[109] ;
  assign n3413 = \new_[17432]_  ? \new_[19383]_  : \text_in[89] ;
  assign \new_[18385]_  = ~\new_[19019]_  & ~\new_[19426]_ ;
  assign \new_[18386]_  = ~\new_[19318]_ ;
  assign \new_[18387]_  = \new_[14766]_  ^ \new_[1660]_ ;
  assign \new_[18388]_  = \new_[19591]_  ^ \new_[19792]_ ;
  assign \new_[18389]_  = ~\new_[19039]_  | ~\new_[21578]_ ;
  assign \new_[18390]_  = ~\new_[19685]_ ;
  assign \new_[18391]_  = ~\new_[18772]_ ;
  assign \new_[18392]_  = ~\new_[18012]_  & ~\new_[19050]_ ;
  assign \new_[18393]_  = \new_[19202]_  | \new_[19600]_ ;
  assign \new_[18394]_  = ~\new_[18624]_ ;
  assign \new_[18395]_  = \new_[14922]_  ^ \new_[1474]_ ;
  assign \new_[18396]_  = \new_[19046]_  | \new_[19205]_ ;
  assign \new_[18397]_  = ~\new_[20035]_  | ~\new_[21583]_ ;
  assign \new_[18398]_  = ~\new_[18770]_ ;
  assign \new_[18399]_  = ~\new_[18606]_ ;
  assign \new_[18400]_  = ~\new_[19126]_  | ~\new_[19596]_ ;
  assign \new_[18401]_  = \new_[14765]_  ^ \new_[1349]_ ;
  assign \new_[18402]_  = \new_[19553]_  & \new_[19190]_ ;
  assign \new_[18403]_  = ~\new_[18751]_ ;
  assign \new_[18404]_  = ~\new_[18689]_ ;
  assign \new_[18405]_  = ~\new_[20294]_ ;
  assign \new_[18406]_  = ~\new_[1039]_ ;
  assign n3383 = \new_[17201]_  ? \new_[19479]_  : \text_in[21] ;
  assign \new_[18408]_  = ~\new_[19127]_ ;
  assign \new_[18409]_  = ~\new_[18599]_ ;
  assign \new_[18410]_  = ~\new_[19014]_  | ~\new_[18979]_ ;
  assign \new_[18411]_  = ~\new_[18589]_ ;
  assign \new_[18412]_  = \new_[19244]_  | \new_[20641]_ ;
  assign \new_[18413]_  = \new_[17087]_  ^ \new_[1350]_ ;
  assign \new_[18414]_  = ~\new_[18773]_ ;
  assign \new_[18415]_  = ~\new_[21491]_  & ~\new_[19462]_ ;
  assign \new_[18416]_  = ~\new_[18701]_ ;
  assign \new_[18417]_  = ~\new_[18713]_ ;
  assign \new_[18418]_  = ~\new_[18798]_ ;
  assign \new_[18419]_  = \new_[19690]_  ^ \new_[19666]_ ;
  assign \new_[18420]_  = ~\new_[18933]_ ;
  assign \new_[18421]_  = ~\new_[19388]_ ;
  assign \new_[18422]_  = \new_[19781]_  ^ \new_[19280]_ ;
  assign \new_[18423]_  = ~\new_[21165]_ ;
  assign \new_[18424]_  = ~\new_[18732]_ ;
  assign \new_[18425]_  = ~\new_[19680]_  & ~\new_[19788]_ ;
  assign \new_[18426]_  = \new_[19682]_  ^ \new_[19345]_ ;
  assign \new_[18427]_  = ~\new_[20486]_ ;
  assign \new_[18428]_  = ~\new_[18953]_ ;
  assign \new_[18429]_  = ~\new_[18975]_  & ~\new_[21513]_ ;
  assign \new_[18430]_  = ~\new_[18910]_ ;
  assign \new_[18431]_  = \new_[19579]_  ^ \new_[19768]_ ;
  assign \new_[18432]_  = ~\new_[18935]_  | ~\new_[19211]_ ;
  assign \new_[18433]_  = ~\new_[18934]_ ;
  assign \new_[18434]_  = ~\new_[19356]_  & ~\new_[19548]_ ;
  assign \new_[18435]_  = \new_[15470]_  ^ \new_[1669]_ ;
  assign \new_[18436]_  = ~\new_[19742]_  | ~\new_[18832]_ ;
  assign \new_[18437]_  = \new_[15845]_  ^ \new_[19631]_ ;
  assign n3268 = \new_[16795]_  ? \new_[19372]_  : \text_in[73] ;
  assign \new_[18439]_  = ~\new_[21568]_  | ~\new_[19409]_ ;
  assign \new_[18440]_  = ~\new_[18896]_ ;
  assign n3298 = \new_[16918]_  ? \new_[19338]_  : \text_in[95] ;
  assign \new_[18442]_  = ~\new_[19625]_  | ~\new_[19188]_ ;
  assign \new_[18443]_  = ~\new_[20240]_ ;
  assign n3403 = \new_[17404]_  ? ld : \text_in[38] ;
  assign \new_[18445]_  = \new_[19159]_  | \new_[21166]_ ;
  assign \new_[18446]_  = ~\new_[19454]_  | ~\new_[18008]_ ;
  assign \new_[18447]_  = \new_[19211]_  | \new_[19654]_ ;
  assign \new_[18448]_  = ~\new_[18874]_ ;
  assign \new_[18449]_  = ~\new_[18919]_ ;
  assign \new_[18450]_  = ~\new_[19010]_  & ~\new_[19092]_ ;
  assign \new_[18451]_  = ~\new_[18642]_ ;
  assign \new_[18452]_  = \new_[19069]_  & \new_[19412]_ ;
  assign \new_[18453]_  = \new_[19595]_  ^ \new_[1421]_ ;
  assign \new_[18454]_  = \new_[18661]_ ;
  assign \new_[18455]_  = ~\new_[18665]_ ;
  assign \new_[18456]_  = ~\new_[18876]_ ;
  assign \new_[18457]_  = ~\new_[18687]_ ;
  assign \new_[18458]_  = ~\new_[18944]_  | ~\new_[19788]_ ;
  assign \new_[18459]_  = ~\new_[18704]_ ;
  assign \new_[18460]_  = ~\new_[19508]_  | ~\new_[19186]_ ;
  assign \new_[18461]_  = ~\new_[18604]_ ;
  assign \new_[18462]_  = ~\new_[18610]_ ;
  assign \new_[18463]_  = \new_[19797]_  ^ \new_[19761]_ ;
  assign \new_[18464]_  = ~\new_[18765]_ ;
  assign \new_[18465]_  = ~\new_[18622]_ ;
  assign \new_[18466]_  = \new_[19742]_  | \new_[19578]_ ;
  assign \new_[18467]_  = \new_[19783]_  ^ \new_[1862]_ ;
  assign \new_[18468]_  = ~\new_[18786]_ ;
  assign \new_[18469]_  = \new_[19248]_  | \new_[19298]_ ;
  assign \new_[18470]_  = \new_[14778]_  ^ \new_[1662]_ ;
  assign \new_[18471]_  = \new_[19634]_  ^ \new_[1343]_ ;
  assign \new_[18472]_  = \new_[19745]_  | \new_[19435]_ ;
  assign \new_[18473]_  = \new_[19145]_  | \new_[19336]_ ;
  assign \new_[18474]_  = ~\new_[19413]_ ;
  assign \new_[18475]_  = ~\new_[19132]_  | ~\new_[19328]_ ;
  assign \new_[18476]_  = ~\new_[18949]_  | ~\new_[19055]_ ;
  assign \new_[18477]_  = ~\new_[18850]_ ;
  assign \new_[18478]_  = ~\new_[19216]_  | ~\new_[19513]_ ;
  assign \new_[18479]_  = ~\new_[19689]_  | ~\new_[19055]_ ;
  assign \new_[18480]_  = \new_[18634]_ ;
  assign \new_[18481]_  = \new_[20680]_ ;
  assign \new_[18482]_  = ~\new_[19109]_  & ~\new_[19685]_ ;
  assign \new_[18483]_  = ~\new_[20310]_ ;
  assign \new_[18484]_  = \new_[19583]_  | \new_[19603]_ ;
  assign \new_[18485]_  = ~\new_[18785]_ ;
  assign \new_[18486]_  = \new_[19263]_  | \new_[19655]_ ;
  assign \new_[18487]_  = \new_[14776]_  ^ \new_[19628]_ ;
  assign n3323 = \new_[17004]_  ? \new_[19338]_  : \text_in[122] ;
  assign \new_[18489]_  = ~\new_[19127]_ ;
  assign \new_[18490]_  = ~\new_[19357]_  | ~\new_[19600]_ ;
  assign \new_[18491]_  = ~\new_[19568]_  & ~\new_[19272]_ ;
  assign \new_[18492]_  = ~\new_[18686]_ ;
  assign \new_[18493]_  = ~\new_[19354]_  | ~\new_[19168]_ ;
  assign \new_[18494]_  = \new_[20100]_  & \new_[1033]_ ;
  assign n3228 = \new_[16701]_  ? \new_[19472]_  : \text_in[44] ;
  assign \new_[18496]_  = ~\new_[19127]_ ;
  assign \new_[18497]_  = ~\new_[19012]_  & ~\new_[19603]_ ;
  assign \new_[18498]_  = ~\new_[19384]_ ;
  assign \new_[18499]_  = \new_[15923]_  | \new_[19697]_ ;
  assign \new_[18500]_  = ~\new_[19147]_  | ~\new_[19485]_ ;
  assign \new_[18501]_  = ~\new_[18614]_ ;
  assign \new_[18502]_  = \new_[15259]_  ^ \new_[1666]_ ;
  assign \new_[18503]_  = \new_[19704]_  ^ \new_[19658]_ ;
  assign \new_[18504]_  = \new_[19605]_  ^ \new_[19799]_ ;
  assign \new_[18505]_  = \new_[19766]_  ^ \new_[1239]_ ;
  assign \new_[18506]_  = ~\new_[18791]_ ;
  assign \new_[18507]_  = \new_[19667]_  ^ \new_[19739]_ ;
  assign \new_[18508]_  = ~\new_[18908]_ ;
  assign \new_[18509]_  = ~\new_[19165]_  | ~\new_[21516]_ ;
  assign \new_[18510]_  = ~\new_[18792]_ ;
  assign \new_[18511]_  = ~\new_[19302]_  & ~\new_[19055]_ ;
  assign n3283 = \new_[16848]_  ? \new_[19472]_  : \text_in[114] ;
  assign \new_[18513]_  = \new_[19677]_  ^ \new_[19673]_ ;
  assign \new_[18514]_  = \new_[15059]_  ^ \new_[19505]_ ;
  assign n3238 = \new_[16723]_  ? \new_[19451]_  : \text_in[101] ;
  assign \new_[18516]_  = ~\new_[19037]_  | ~\new_[19081]_ ;
  assign \new_[18517]_  = ~\new_[19645]_  | ~\new_[19050]_ ;
  assign \new_[18518]_  = ~\new_[18860]_ ;
  assign \new_[18519]_  = ~\new_[19184]_ ;
  assign \new_[18520]_  = ~\new_[19566]_  | ~\new_[19332]_ ;
  assign \new_[18521]_  = ~\new_[18894]_ ;
  assign \new_[18522]_  = ~\new_[19072]_  & ~\new_[954]_ ;
  assign \new_[18523]_  = ~\new_[18662]_ ;
  assign \new_[18524]_  = ~\new_[18729]_ ;
  assign \new_[18525]_  = ~\new_[18941]_  & ~\new_[960]_ ;
  assign \new_[18526]_  = ~\new_[18746]_ ;
  assign \new_[18527]_  = ~\new_[18955]_  & ~\new_[19008]_ ;
  assign \new_[18528]_  = ~\new_[18836]_ ;
  assign \new_[18529]_  = ~\new_[19493]_  | ~\new_[19431]_ ;
  assign \new_[18530]_  = ~\new_[1087]_  | ~\new_[19068]_ ;
  assign n3343 = \new_[17053]_  ? ld : \text_in[113] ;
  assign \new_[18532]_  = \new_[19570]_  ^ \new_[1421]_ ;
  assign \new_[18533]_  = ~\new_[18713]_ ;
  assign n3263 = \new_[16777]_  ? ld : \text_in[93] ;
  assign \new_[18535]_  = ~\new_[20750]_ ;
  assign \new_[18536]_  = ~\new_[18724]_ ;
  assign \new_[18537]_  = \new_[19713]_  | \new_[1878]_ ;
  assign \new_[18538]_  = \new_[18542]_  & \new_[999]_ ;
  assign \new_[18539]_  = ~\new_[19180]_  | ~\new_[18984]_ ;
  assign \new_[18540]_  = ~\new_[19687]_  | ~\new_[19040]_ ;
  assign \new_[18541]_  = \new_[18691]_ ;
  assign \new_[18542]_  = ~\new_[1006]_ ;
  assign \new_[18543]_  = ~\new_[18609]_ ;
  assign \new_[18544]_  = \new_[19153]_  & \new_[19578]_ ;
  assign \new_[18545]_  = ~\new_[19815]_  | ~\new_[19407]_ ;
  assign \new_[18546]_  = ~\new_[18924]_ ;
  assign \new_[18547]_  = ~\new_[18623]_ ;
  assign \new_[18548]_  = ~\new_[19268]_  | ~\new_[19272]_ ;
  assign \new_[18549]_  = ~\new_[18853]_ ;
  assign n3333 = \new_[17030]_  ? ld : \text_in[102] ;
  assign \new_[18551]_  = ~\new_[1081]_  | ~\new_[21686]_ ;
  assign \new_[18552]_  = ~\new_[19086]_  & ~\new_[20751]_ ;
  assign \new_[18553]_  = ~\new_[18617]_ ;
  assign \new_[18554]_  = ~\new_[18727]_ ;
  assign \new_[18555]_  = ~\new_[18813]_ ;
  assign \new_[18556]_  = \new_[19802]_  ^ \new_[19565]_ ;
  assign \new_[18557]_  = ~\new_[18930]_ ;
  assign \new_[18558]_  = ~\new_[18657]_ ;
  assign \new_[18559]_  = \new_[19625]_  | \new_[19068]_ ;
  assign \new_[18560]_  = ~\new_[18140]_  & ~\new_[20589]_ ;
  assign \new_[18561]_  = ~\new_[19256]_  | ~\new_[21521]_ ;
  assign \new_[18562]_  = \new_[19165]_  | \new_[20487]_ ;
  assign \new_[18563]_  = ~\new_[21534]_  & ~\new_[21517]_ ;
  assign \new_[18564]_  = ~\new_[18974]_  | ~\new_[19219]_ ;
  assign \new_[18565]_  = ~\new_[18843]_ ;
  assign \new_[18566]_  = ~\new_[18991]_  | ~\new_[19074]_ ;
  assign \new_[18567]_  = ~\new_[18596]_ ;
  assign \new_[18568]_  = ~\new_[1084]_  | ~\new_[18605]_ ;
  assign \new_[18569]_  = ~\new_[19525]_ ;
  assign \new_[18570]_  = ~\new_[19098]_  & ~\new_[18832]_ ;
  assign \new_[18571]_  = ~\new_[18685]_ ;
  assign \new_[18572]_  = ~\new_[19243]_ ;
  assign \new_[18573]_  = ~\new_[19500]_ ;
  assign \new_[18574]_  = \new_[14814]_  ^ \new_[1088]_ ;
  assign \new_[18575]_  = ~\new_[18854]_ ;
  assign \new_[18576]_  = \new_[14956]_  ^ \new_[1237]_ ;
  assign \new_[18577]_  = ~\new_[18982]_ ;
  assign \new_[18578]_  = ~\new_[19655]_  & ~\new_[19160]_ ;
  assign \new_[18579]_  = ~\new_[18991]_  & ~\new_[19209]_ ;
  assign \new_[18580]_  = ~\new_[18666]_ ;
  assign n3393 = \new_[17397]_  ? \new_[19479]_  : \text_in[22] ;
  assign \new_[18582]_  = \new_[19086]_  & \new_[20751]_ ;
  assign \new_[18583]_  = ~\new_[19619]_ ;
  assign \new_[18584]_  = ~\new_[19292]_  & ~\new_[18973]_ ;
  assign \new_[18585]_  = ~\new_[19000]_  & ~\new_[21513]_ ;
  assign \new_[18586]_  = ~\new_[19067]_ ;
  assign \new_[18587]_  = ~\new_[19009]_ ;
  assign \new_[18588]_  = ~\new_[19711]_  | ~\new_[18008]_ ;
  assign \new_[18589]_  = ~\new_[19312]_  | ~\new_[19759]_ ;
  assign \new_[18590]_  = ~\new_[19016]_ ;
  assign \new_[18591]_  = ~\new_[19056]_ ;
  assign \new_[18592]_  = ~\new_[19524]_  & ~\new_[19791]_ ;
  assign \new_[18593]_  = ~\new_[19252]_ ;
  assign \new_[18594]_  = ~\new_[19780]_ ;
  assign \new_[18595]_  = \new_[19393]_  | \new_[19425]_ ;
  assign \new_[18596]_  = ~\new_[18995]_ ;
  assign \new_[18597]_  = ~\new_[19027]_ ;
  assign \new_[18598]_  = ~\new_[19778]_  & ~\new_[19663]_ ;
  assign \new_[18599]_  = ~\new_[19170]_ ;
  assign \new_[18600]_  = \new_[19622]_  & \new_[19654]_ ;
  assign \new_[18601]_  = ~\new_[19172]_ ;
  assign \new_[18602]_  = \new_[19626]_  ^ \new_[19633]_ ;
  assign \new_[18603]_  = ~\new_[20237]_ ;
  assign \new_[18604]_  = ~\new_[19010]_ ;
  assign \new_[18605]_  = ~\new_[20486]_ ;
  assign \new_[18606]_  = \new_[20704]_ ;
  assign \new_[18607]_  = ~\new_[18955]_ ;
  assign \new_[18608]_  = \new_[19618]_  ^ \new_[1518]_ ;
  assign \new_[18609]_  = ~\new_[19076]_ ;
  assign \new_[18610]_  = ~\new_[19622]_  | ~\new_[19449]_ ;
  assign \new_[18611]_  = \new_[19733]_  ^ \new_[19749]_ ;
  assign \new_[18612]_  = ~\new_[18997]_ ;
  assign \new_[18613]_  = ~\new_[19461]_  | ~\new_[19435]_ ;
  assign \new_[18614]_  = \new_[19597]_  & \new_[19663]_ ;
  assign \new_[18615]_  = ~\new_[19390]_ ;
  assign \new_[18616]_  = ~\new_[19149]_ ;
  assign \new_[18617]_  = ~\new_[18990]_ ;
  assign \new_[18618]_  = ~\new_[19263]_ ;
  assign \new_[18619]_  = ~\new_[19157]_ ;
  assign \new_[18620]_  = ~\new_[19089]_ ;
  assign \new_[18621]_  = ~\new_[19469]_ ;
  assign \new_[18622]_  = ~\new_[19288]_  | ~\new_[19360]_ ;
  assign \new_[18623]_  = \new_[19230]_ ;
  assign \new_[18624]_  = ~\new_[20699]_ ;
  assign \new_[18625]_  = ~\new_[19330]_  | ~\new_[21585]_ ;
  assign \new_[18626]_  = ~\new_[19481]_  | ~\new_[19568]_ ;
  assign \new_[18627]_  = \new_[20704]_ ;
  assign \new_[18628]_  = ~\new_[19069]_ ;
  assign \new_[18629]_  = ~\new_[19411]_  | ~\new_[19402]_ ;
  assign \new_[18630]_  = \new_[19571]_  ^ \new_[1187]_ ;
  assign \new_[18631]_  = ~\new_[17447]_  | ~\new_[19290]_ ;
  assign \new_[18632]_  = ~\new_[19085]_ ;
  assign \new_[18633]_  = ~\new_[19060]_ ;
  assign \new_[18634]_  = \new_[19086]_ ;
  assign \new_[18635]_  = ~\new_[18992]_ ;
  assign \new_[18636]_  = ~\new_[19114]_  | ~\new_[19665]_ ;
  assign \new_[18637]_  = ~\new_[19007]_ ;
  assign \new_[18638]_  = ~\new_[19422]_  & ~\new_[19788]_ ;
  assign \new_[18639]_  = ~\new_[19135]_ ;
  assign \new_[18640]_  = ~\new_[19139]_ ;
  assign \new_[18641]_  = ~\new_[19659]_ ;
  assign \new_[18642]_  = ~\new_[19364]_  | ~\new_[19455]_ ;
  assign \new_[18643]_  = ~\new_[19178]_ ;
  assign \new_[18644]_  = ~\new_[19141]_ ;
  assign \new_[18645]_  = ~\new_[19232]_ ;
  assign \new_[18646]_  = ~\new_[19110]_ ;
  assign \new_[18647]_  = ~\new_[19272]_ ;
  assign \new_[18648]_  = ~\new_[19489]_  | ~\new_[19789]_ ;
  assign \new_[18649]_  = ~\new_[19638]_ ;
  assign \new_[18650]_  = ~\new_[1081]_ ;
  assign \new_[18651]_  = ~\new_[19081]_ ;
  assign \new_[18652]_  = ~\new_[19499]_ ;
  assign \new_[18653]_  = ~\new_[19227]_ ;
  assign \new_[18654]_  = ~\new_[19506]_  & ~\new_[21585]_ ;
  assign \new_[18655]_  = ~\new_[19366]_ ;
  assign \new_[18656]_  = ~\new_[19050]_ ;
  assign \new_[18657]_  = ~\new_[19029]_  | ~\new_[19754]_ ;
  assign \new_[18658]_  = \new_[19598]_  ^ \new_[19593]_ ;
  assign \new_[18659]_  = \new_[19189]_ ;
  assign \new_[18660]_  = ~\new_[19267]_ ;
  assign \new_[18661]_  = ~\new_[18958]_ ;
  assign \new_[18662]_  = ~\new_[19501]_  | ~\new_[19734]_ ;
  assign \new_[18663]_  = ~\new_[19147]_ ;
  assign \new_[18664]_  = ~\new_[19139]_ ;
  assign \new_[18665]_  = ~\new_[19393]_  | ~\new_[19611]_ ;
  assign \new_[18666]_  = ~\new_[19487]_  | ~\new_[19546]_ ;
  assign \new_[18667]_  = ~\new_[19578]_ ;
  assign \new_[18668]_  = ~\new_[19717]_ ;
  assign \new_[18669]_  = ~\new_[18954]_ ;
  assign \new_[18670]_  = ~\new_[18971]_ ;
  assign \new_[18671]_  = ~\new_[19315]_  | ~\new_[18390]_ ;
  assign \new_[18672]_  = ~\new_[19250]_ ;
  assign \new_[18673]_  = ~\new_[19264]_ ;
  assign \new_[18674]_  = ~\new_[19052]_ ;
  assign \new_[18675]_  = ~\new_[19046]_ ;
  assign \new_[18676]_  = ~\new_[19223]_ ;
  assign \new_[18677]_  = \new_[17091]_  ^ \new_[19618]_ ;
  assign \new_[18678]_  = ~\new_[19149]_ ;
  assign \new_[18679]_  = \new_[19784]_  ^ \new_[19710]_ ;
  assign \new_[18680]_  = ~\new_[18956]_ ;
  assign \new_[18681]_  = ~\new_[19235]_ ;
  assign \new_[18682]_  = ~\new_[19432]_ ;
  assign \new_[18683]_  = ~\new_[18950]_ ;
  assign \new_[18684]_  = \new_[19633]_  ^ \new_[1510]_ ;
  assign \new_[18685]_  = ~\new_[19494]_  | ~\new_[19344]_ ;
  assign \new_[18686]_  = ~\new_[19137]_ ;
  assign \new_[18687]_  = ~\new_[19365]_  | ~\new_[19572]_ ;
  assign \new_[18688]_  = ~\new_[19058]_ ;
  assign \new_[18689]_  = ~\new_[19506]_  | ~\new_[19692]_ ;
  assign \new_[18690]_  = ~\new_[19580]_  | ~\new_[19296]_ ;
  assign \new_[18691]_  = ~\new_[19038]_ ;
  assign \new_[18692]_  = ~\new_[19406]_ ;
  assign \new_[18693]_  = \new_[19687]_ ;
  assign \new_[18694]_  = ~\new_[18959]_ ;
  assign \new_[18695]_  = ~\new_[19437]_  & ~\new_[19788]_ ;
  assign \new_[18696]_  = \new_[19593]_  ^ \new_[19551]_ ;
  assign \new_[18697]_  = ~\new_[19542]_  | ~\new_[19629]_ ;
  assign \new_[18698]_  = ~\new_[19062]_ ;
  assign \new_[18699]_  = ~\new_[19603]_ ;
  assign \new_[18700]_  = \new_[19274]_  & \new_[19789]_ ;
  assign \new_[18701]_  = ~\new_[991]_  & ~\new_[21638]_ ;
  assign \new_[18702]_  = ~\new_[19670]_  & ~\new_[19321]_ ;
  assign \new_[18703]_  = ~\new_[19649]_ ;
  assign \new_[18704]_  = ~\new_[19164]_ ;
  assign \new_[18705]_  = ~\new_[19521]_  | ~\new_[19743]_ ;
  assign \new_[18706]_  = \new_[17404]_  ^ \new_[19662]_ ;
  assign \new_[18707]_  = ~\new_[19155]_ ;
  assign \new_[18708]_  = ~\new_[21571]_  & ~\new_[19409]_ ;
  assign \new_[18709]_  = ~\new_[19499]_ ;
  assign \new_[18710]_  = ~\new_[19368]_  | ~\new_[21517]_ ;
  assign \new_[18711]_  = ~\new_[19587]_  | ~\new_[19423]_ ;
  assign \new_[18712]_  = \new_[19731]_  ^ \new_[19631]_ ;
  assign \new_[18713]_  = ~\new_[19034]_ ;
  assign \new_[18714]_  = ~\new_[18978]_ ;
  assign \new_[18715]_  = \new_[16511]_  ^ \new_[19581]_ ;
  assign \new_[18716]_  = ~\new_[19533]_  | ~\new_[19586]_ ;
  assign \new_[18717]_  = ~\new_[18991]_ ;
  assign \new_[18718]_  = ~\new_[19131]_ ;
  assign \new_[18719]_  = ~\new_[19011]_ ;
  assign \new_[18720]_  = ~\new_[19001]_ ;
  assign \new_[18721]_  = ~\new_[19308]_  | ~\new_[19721]_ ;
  assign \new_[18722]_  = ~\new_[19274]_  | ~\new_[19463]_ ;
  assign \new_[18723]_  = \new_[19766]_  ^ \new_[19544]_ ;
  assign \new_[18724]_  = ~\new_[19185]_ ;
  assign \new_[18725]_  = \new_[19355]_  | \new_[19603]_ ;
  assign \new_[18726]_  = ~\new_[19311]_  | ~\new_[20167]_ ;
  assign \new_[18727]_  = ~\new_[19218]_ ;
  assign \new_[18728]_  = \new_[21413]_  & \new_[19538]_ ;
  assign \new_[18729]_  = ~\new_[19278]_  & ~\new_[19574]_ ;
  assign \new_[18730]_  = ~\new_[19109]_ ;
  assign \new_[18731]_  = \new_[19592]_  | \new_[19410]_ ;
  assign \new_[18732]_  = ~\new_[19411]_  & ~\new_[19734]_ ;
  assign \new_[18733]_  = ~\new_[19191]_ ;
  assign \new_[18734]_  = ~\new_[19241]_ ;
  assign \new_[18735]_  = ~\new_[19113]_ ;
  assign \new_[18736]_  = ~\new_[19364]_  | ~\new_[19514]_ ;
  assign \new_[18737]_  = \new_[19796]_  ^ \new_[19704]_ ;
  assign \new_[18738]_  = ~\new_[19566]_  | ~\new_[19346]_ ;
  assign \new_[18739]_  = ~\new_[19625]_ ;
  assign \new_[18740]_  = ~\new_[19020]_ ;
  assign \new_[18741]_  = ~\new_[19160]_ ;
  assign \new_[18742]_  = ~\new_[21536]_  | ~\new_[19286]_ ;
  assign \new_[18743]_  = ~\new_[19234]_ ;
  assign \new_[18744]_  = ~\new_[21562]_  | ~\new_[19403]_ ;
  assign \new_[18745]_  = ~\new_[19264]_ ;
  assign \new_[18746]_  = ~\new_[19518]_  | ~\new_[19430]_ ;
  assign \new_[18747]_  = ~\new_[19099]_ ;
  assign \new_[18748]_  = ~\key[24]  | ~\new_[19363]_ ;
  assign \new_[18749]_  = \new_[19562]_  ^ \new_[19579]_ ;
  assign \new_[18750]_  = ~\new_[19112]_ ;
  assign \new_[18751]_  = ~\new_[21632]_  | ~\new_[19476]_ ;
  assign \new_[18752]_  = ~\new_[21560]_  & ~\new_[19619]_ ;
  assign \new_[18753]_  = ~\new_[2302]_  | ~\new_[19697]_ ;
  assign \new_[18754]_  = ~\new_[19159]_ ;
  assign \new_[18755]_  = ~\new_[19093]_ ;
  assign \new_[18756]_  = \new_[19610]_  ^ \new_[19783]_ ;
  assign \new_[18757]_  = ~\new_[19195]_ ;
  assign \new_[18758]_  = \new_[19634]_  ^ \new_[19569]_ ;
  assign \new_[18759]_  = \new_[21557]_  & \new_[944]_ ;
  assign \new_[18760]_  = \new_[19726]_  ^ \new_[19714]_ ;
  assign \new_[18761]_  = ~\new_[18953]_ ;
  assign \new_[18762]_  = ~\new_[19237]_ ;
  assign \new_[18763]_  = ~\new_[19002]_ ;
  assign \new_[18764]_  = \new_[19710]_  ^ \new_[19774]_ ;
  assign \new_[18765]_  = ~\new_[19090]_ ;
  assign \new_[18766]_  = ~\new_[19149]_ ;
  assign \new_[18767]_  = \new_[19544]_  ^ \new_[1239]_ ;
  assign \new_[18768]_  = ~\new_[21544]_  | ~\new_[19712]_ ;
  assign \new_[18769]_  = ~\new_[21413]_ ;
  assign \new_[18770]_  = ~\new_[18976]_ ;
  assign \new_[18771]_  = ~\new_[19167]_ ;
  assign \new_[18772]_  = ~\new_[19355]_ ;
  assign \new_[18773]_  = ~\new_[19190]_ ;
  assign \new_[18774]_  = ~\new_[19119]_ ;
  assign \new_[18775]_  = ~rst | ~\new_[19415]_ ;
  assign \new_[18776]_  = ~\new_[19225]_ ;
  assign \new_[18777]_  = ~\new_[19515]_  & ~\new_[19635]_ ;
  assign \new_[18778]_  = \new_[21413]_ ;
  assign \new_[18779]_  = ~\new_[19238]_ ;
  assign \new_[18780]_  = ~\new_[19282]_  | ~\new_[19449]_ ;
  assign \new_[18781]_  = ~\new_[19461]_  | ~\new_[19608]_ ;
  assign \new_[18782]_  = ~\new_[19039]_ ;
  assign \new_[18783]_  = ~\new_[19258]_ ;
  assign \new_[18784]_  = ~\new_[18982]_ ;
  assign \new_[18785]_  = ~\new_[19065]_ ;
  assign \new_[18786]_  = ~\new_[19381]_  & ~\new_[19659]_ ;
  assign \new_[18787]_  = ~\new_[973]_ ;
  assign \new_[18788]_  = ~\new_[19597]_  & ~\new_[19663]_ ;
  assign \new_[18789]_  = ~\new_[19079]_ ;
  assign \new_[18790]_  = ~\new_[21631]_  | ~\new_[19333]_ ;
  assign \new_[18791]_  = ~\new_[19550]_ ;
  assign \new_[18792]_  = ~\new_[21308]_ ;
  assign \new_[18793]_  = ~\new_[19012]_ ;
  assign \new_[18794]_  = ~\new_[21307]_ ;
  assign \new_[18795]_  = \new_[18542]_ ;
  assign \new_[18796]_  = ~\new_[19419]_  | ~\new_[19738]_ ;
  assign \new_[18797]_  = ~\new_[19053]_ ;
  assign \new_[18798]_  = ~\new_[19559]_ ;
  assign \new_[18799]_  = ~\new_[19116]_ ;
  assign \new_[18800]_  = ~\new_[21304]_  | ~\new_[19683]_ ;
  assign \new_[18801]_  = ~\new_[19035]_ ;
  assign \new_[18802]_  = ~\new_[19055]_ ;
  assign \new_[18803]_  = ~\new_[19170]_ ;
  assign \new_[18804]_  = ~\new_[20749]_ ;
  assign \new_[18805]_  = ~\new_[19671]_  | ~\new_[19352]_ ;
  assign \new_[18806]_  = ~\new_[19125]_ ;
  assign \new_[18807]_  = ~\new_[19128]_ ;
  assign \new_[18808]_  = ~\new_[21142]_ ;
  assign \new_[18809]_  = ~\new_[19063]_ ;
  assign \new_[18810]_  = ~\new_[19482]_ ;
  assign \new_[18811]_  = \new_[19189]_ ;
  assign \new_[18812]_  = ~\new_[19468]_  | ~\new_[19603]_ ;
  assign \new_[18813]_  = \new_[19312]_  & \new_[19495]_ ;
  assign \new_[18814]_  = ~\new_[19256]_ ;
  assign \new_[18815]_  = ~\new_[19199]_ ;
  assign \new_[18816]_  = ~\new_[1511]_  & ~\new_[19589]_ ;
  assign \new_[18817]_  = ~\new_[20903]_ ;
  assign \new_[18818]_  = ~\new_[19171]_ ;
  assign \new_[18819]_  = ~\new_[19126]_ ;
  assign \new_[18820]_  = \new_[19632]_  ^ \new_[19677]_ ;
  assign \new_[18821]_  = ~\new_[20679]_ ;
  assign \new_[18822]_  = \new_[19810]_  ^ \new_[19588]_ ;
  assign \new_[18823]_  = ~\new_[19056]_ ;
  assign \new_[18824]_  = ~\new_[19004]_ ;
  assign \new_[18825]_  = ~\new_[21413]_  & ~\new_[19538]_ ;
  assign \new_[18826]_  = \new_[19459]_  & \new_[19674]_ ;
  assign \new_[18827]_  = ~\new_[20704]_ ;
  assign \new_[18828]_  = \new_[19776]_  ^ \new_[19690]_ ;
  assign \new_[18829]_  = ~\new_[1243]_ ;
  assign \new_[18830]_  = \new_[19605]_  ^ \new_[1346]_ ;
  assign \new_[18831]_  = ~\new_[19078]_ ;
  assign \new_[18832]_  = ~\new_[19279]_ ;
  assign \new_[18833]_  = ~\new_[19177]_ ;
  assign \new_[18834]_  = ~\new_[19205]_ ;
  assign \new_[18835]_  = \new_[19761]_  ^ \new_[19700]_ ;
  assign \new_[18836]_  = ~\new_[19366]_  | ~\new_[1878]_ ;
  assign \new_[18837]_  = ~\new_[18944]_ ;
  assign \new_[18838]_  = ~\new_[19221]_ ;
  assign \new_[18839]_  = \new_[19655]_  & \new_[19393]_ ;
  assign \new_[18840]_  = ~\new_[19469]_ ;
  assign \new_[18841]_  = ~\new_[19680]_ ;
  assign \new_[18842]_  = ~\new_[19226]_ ;
  assign \new_[18843]_  = ~\new_[19201]_ ;
  assign \new_[18844]_  = ~\new_[19448]_ ;
  assign \new_[18845]_  = ~\new_[19707]_ ;
  assign \new_[18846]_  = ~\new_[18981]_ ;
  assign \new_[18847]_  = ~\new_[19103]_ ;
  assign \new_[18848]_  = \new_[19760]_  ^ \new_[1667]_ ;
  assign \new_[18849]_  = ~\new_[19288]_  & ~\new_[19425]_ ;
  assign \new_[18850]_  = ~\new_[18946]_ ;
  assign \new_[18851]_  = \new_[19570]_  ^ \new_[19595]_ ;
  assign \new_[18852]_  = ~\new_[19122]_ ;
  assign \new_[18853]_  = ~\new_[19516]_  | ~\new_[20167]_ ;
  assign \new_[18854]_  = ~\new_[19023]_ ;
  assign \new_[18855]_  = \new_[18957]_ ;
  assign \new_[18856]_  = \new_[19753]_  ^ \new_[19682]_ ;
  assign \new_[18857]_  = \new_[19023]_ ;
  assign \new_[18858]_  = \new_[19575]_  ^ \new_[19662]_ ;
  assign \new_[18859]_  = ~\new_[19222]_ ;
  assign \new_[18860]_  = ~\new_[19514]_  & ~\new_[21494]_ ;
  assign \new_[18861]_  = \new_[19093]_ ;
  assign \new_[18862]_  = \new_[19524]_  & \new_[19582]_ ;
  assign \new_[18863]_  = ~\new_[19005]_ ;
  assign \new_[18864]_  = ~\new_[19291]_  | ~\new_[19685]_ ;
  assign \new_[18865]_  = \new_[19569]_  ^ \new_[1343]_ ;
  assign \new_[18866]_  = \new_[19630]_  ^ \new_[19667]_ ;
  assign \new_[18867]_  = ~\new_[19074]_ ;
  assign \new_[18868]_  = ~\new_[19389]_  | ~\new_[21100]_ ;
  assign \new_[18869]_  = ~\new_[19362]_  & ~\new_[20927]_ ;
  assign \new_[18870]_  = ~\new_[19389]_  | ~\new_[19777]_ ;
  assign \new_[18871]_  = \new_[19315]_  | \new_[19685]_ ;
  assign \new_[18872]_  = ~\new_[19347]_  | ~\new_[19604]_ ;
  assign \new_[18873]_  = ~\new_[19073]_ ;
  assign \new_[18874]_  = ~\new_[19265]_ ;
  assign \new_[18875]_  = ~\new_[19711]_  | ~\new_[19443]_ ;
  assign \new_[18876]_  = ~\new_[19437]_  | ~\new_[19701]_ ;
  assign \new_[18877]_  = ~\new_[19142]_ ;
  assign \new_[18878]_  = ~\new_[19518]_  | ~\new_[19629]_ ;
  assign \new_[18879]_  = \new_[19657]_  ^ \new_[19735]_ ;
  assign \new_[18880]_  = \new_[1288]_  ^ \new_[19552]_ ;
  assign \new_[18881]_  = ~\new_[19245]_ ;
  assign \new_[18882]_  = ~\new_[19086]_ ;
  assign \new_[18883]_  = ~\new_[19065]_ ;
  assign \new_[18884]_  = ~\new_[19193]_ ;
  assign \new_[18885]_  = ~\new_[19475]_  | ~\new_[21525]_ ;
  assign \new_[18886]_  = ~\new_[19094]_ ;
  assign \new_[18887]_  = \new_[19775]_  ^ \new_[1288]_ ;
  assign \new_[18888]_  = ~\new_[18940]_ ;
  assign \new_[18889]_  = ~\new_[19230]_ ;
  assign \new_[18890]_  = ~\new_[19355]_  | ~\new_[19603]_ ;
  assign \new_[18891]_  = ~\new_[19169]_ ;
  assign \new_[18892]_  = \new_[19549]_  ^ \new_[1474]_ ;
  assign \new_[18893]_  = ~\new_[19106]_ ;
  assign \new_[18894]_  = ~\new_[19668]_  | ~\new_[19489]_ ;
  assign \new_[18895]_  = ~\new_[19163]_ ;
  assign \new_[18896]_  = ~\new_[19182]_ ;
  assign \new_[18897]_  = \new_[19732]_  ^ \new_[19800]_ ;
  assign \new_[18898]_  = ~\new_[18996]_ ;
  assign \new_[18899]_  = ~\new_[21535]_  | ~\new_[19678]_ ;
  assign \new_[18900]_  = ~\new_[19057]_ ;
  assign \new_[18901]_  = ~\new_[19138]_ ;
  assign \new_[18902]_  = ~\new_[19087]_ ;
  assign \new_[18903]_  = \new_[20237]_ ;
  assign \new_[18904]_  = \new_[16892]_  ^ \new_[19783]_ ;
  assign \new_[18905]_  = \new_[19588]_  ^ \new_[1619]_ ;
  assign \new_[18906]_  = ~\new_[19114]_ ;
  assign \new_[18907]_  = ~\key[29]  | ~\new_[19363]_ ;
  assign \new_[18908]_  = ~\new_[19253]_ ;
  assign \new_[18909]_  = ~\new_[18948]_ ;
  assign \new_[18910]_  = \new_[19727]_  & \new_[19298]_ ;
  assign \new_[18911]_  = ~\new_[21536]_  | ~\new_[19678]_ ;
  assign \new_[18912]_  = ~\new_[19312]_  & (~\new_[12134]_  | ~\new_[10818]_ );
  assign \new_[18913]_  = \new_[19655]_  | \new_[19589]_ ;
  assign \new_[18914]_  = ~\new_[19559]_  | ~\new_[18008]_ ;
  assign \new_[18915]_  = \new_[19814]_  ^ \new_[19802]_ ;
  assign \new_[18916]_  = ~\new_[19075]_ ;
  assign \new_[18917]_  = \new_[1347]_  ^ \new_[19686]_ ;
  assign \new_[18918]_  = \new_[19606]_  ^ \new_[19781]_ ;
  assign \new_[18919]_  = ~\new_[19216]_ ;
  assign \new_[18920]_  = ~\new_[19493]_  & ~\new_[19431]_ ;
  assign \new_[18921]_  = \new_[19747]_  ^ \new_[19792]_ ;
  assign \new_[18922]_  = \new_[19590]_  ^ \new_[19737]_ ;
  assign \new_[18923]_  = ~\new_[21558]_  | ~\new_[19275]_ ;
  assign \new_[18924]_  = ~\new_[18986]_ ;
  assign \new_[18925]_  = \new_[19197]_ ;
  assign \new_[18926]_  = ~\new_[19083]_ ;
  assign \new_[18927]_  = ~\new_[19501]_  & ~\new_[19734]_ ;
  assign \new_[18928]_  = ~\new_[18957]_ ;
  assign \new_[18929]_  = ~\new_[19248]_ ;
  assign \new_[18930]_  = \new_[19711]_  | \new_[18008]_ ;
  assign \new_[18931]_  = ~\new_[19762]_  | ~\new_[19589]_ ;
  assign \new_[18932]_  = ~\new_[19557]_  | ~\new_[19468]_ ;
  assign \new_[18933]_  = ~\new_[19108]_ ;
  assign \new_[18934]_  = ~\new_[19466]_  | ~\new_[19701]_ ;
  assign \new_[18935]_  = ~\new_[19503]_ ;
  assign \new_[18936]_  = ~\new_[19568]_  | ~\new_[19361]_ ;
  assign \new_[18937]_  = ~\new_[19559]_ ;
  assign \new_[18938]_  = ~\new_[19407]_ ;
  assign \new_[18939]_  = ~\new_[19465]_ ;
  assign \new_[18940]_  = ~\new_[19434]_ ;
  assign \new_[18941]_  = ~\new_[19492]_ ;
  assign \new_[18942]_  = ~\new_[19300]_ ;
  assign \new_[18943]_  = ~\new_[19538]_ ;
  assign \new_[18944]_  = ~\new_[19437]_ ;
  assign \new_[18945]_  = ~\new_[19500]_ ;
  assign \new_[18946]_  = ~\new_[19411]_ ;
  assign \new_[18947]_  = ~\new_[19482]_ ;
  assign \new_[18948]_  = \new_[18542]_  | \new_[21328]_ ;
  assign \new_[18949]_  = ~\new_[19302]_ ;
  assign \new_[18950]_  = ~\new_[19764]_  & ~\new_[19613]_ ;
  assign \new_[18951]_  = ~\new_[19307]_ ;
  assign \new_[18952]_  = ~\new_[19487]_ ;
  assign \new_[18953]_  = ~\new_[19586]_  & ~\new_[19703]_ ;
  assign \new_[18954]_  = ~\new_[19745]_  & ~\new_[19608]_ ;
  assign \new_[18955]_  = ~\new_[19438]_ ;
  assign \new_[18956]_  = ~\new_[19534]_ ;
  assign \new_[18957]_  = ~\new_[19202]_  & ~\new_[19663]_ ;
  assign \new_[18958]_  = ~\new_[19703]_  | ~\new_[19586]_ ;
  assign \new_[18959]_  = ~\new_[20491]_ ;
  assign \new_[18960]_  = ~\new_[19332]_ ;
  assign \new_[18961]_  = ~\new_[19280]_ ;
  assign \new_[18962]_  = \new_[19555]_  | \new_[19767]_ ;
  assign \new_[18963]_  = ~\new_[19429]_ ;
  assign \new_[18964]_  = ~\new_[20238]_ ;
  assign \new_[18965]_  = ~\new_[19377]_ ;
  assign \new_[18966]_  = ~\new_[19369]_ ;
  assign \new_[18967]_  = ~\new_[1081]_ ;
  assign \new_[18968]_  = ~\new_[21078]_ ;
  assign \new_[18969]_  = ~\new_[19432]_ ;
  assign \new_[18970]_  = ~\new_[19345]_ ;
  assign \new_[18971]_  = ~\new_[19580]_  & ~\new_[19604]_ ;
  assign \new_[18972]_  = ~\new_[19499]_ ;
  assign \new_[18973]_  = ~\new_[21165]_ ;
  assign \new_[18974]_  = ~\new_[19399]_ ;
  assign \new_[18975]_  = ~\new_[19330]_ ;
  assign \new_[18976]_  = ~\new_[19566]_  & ~\new_[19769]_ ;
  assign \new_[18978]_  = ~\new_[19331]_ ;
  assign \new_[18979]_  = ~\new_[19432]_ ;
  assign \new_[18980]_  = ~\new_[19639]_  & ~\new_[19722]_ ;
  assign \new_[18981]_  = ~\new_[19724]_  & ~\new_[19738]_ ;
  assign \new_[18982]_  = \new_[19498]_ ;
  assign \new_[18983]_  = ~\new_[19257]_ ;
  assign \new_[18984]_  = ~\new_[19294]_ ;
  assign \new_[18986]_  = ~\new_[19756]_  & ~\new_[19806]_ ;
  assign \new_[18987]_  = ~\new_[19477]_ ;
  assign \new_[18988]_  = ~\new_[19578]_ ;
  assign \new_[18989]_  = ~\new_[20498]_ ;
  assign \new_[18990]_  = ~\new_[20167]_  & ~\new_[19648]_ ;
  assign \new_[18991]_  = ~\new_[19487]_ ;
  assign \new_[18992]_  = ~\new_[18967]_  | ~\new_[21697]_ ;
  assign \new_[18993]_  = ~\new_[19324]_ ;
  assign \new_[18994]_  = ~\new_[19531]_ ;
  assign \new_[18995]_  = ~\new_[19447]_ ;
  assign \new_[18996]_  = ~\new_[19612]_  | ~\new_[19754]_ ;
  assign \new_[18997]_  = ~\new_[19326]_ ;
  assign \new_[18998]_  = ~\new_[19532]_ ;
  assign \new_[18999]_  = ~\new_[19355]_ ;
  assign \new_[19000]_  = ~\new_[21402]_ ;
  assign \new_[19001]_  = ~\new_[19712]_  | ~\new_[21545]_ ;
  assign \new_[19002]_  = ~\new_[1039]_ ;
  assign \new_[19003]_  = ~\new_[19424]_ ;
  assign \new_[19004]_  = ~\new_[19688]_  & ~\new_[19730]_ ;
  assign \new_[19005]_  = ~\new_[18967]_ ;
  assign \new_[19006]_  = ~\new_[19798]_ ;
  assign \new_[19007]_  = \new_[20486]_ ;
  assign \new_[19008]_  = ~\new_[19511]_ ;
  assign \new_[19009]_  = ~\new_[19637]_ ;
  assign \new_[19010]_  = ~\new_[19296]_ ;
  assign \new_[19011]_  = ~\new_[19743]_  & ~\new_[19734]_ ;
  assign \new_[19012]_  = ~\new_[1656]_  | ~\new_[19583]_ ;
  assign \new_[19013]_  = \new_[19539]_ ;
  assign \new_[19014]_  = ~\new_[19379]_ ;
  assign \new_[19015]_  = ~\new_[19519]_ ;
  assign \new_[19016]_  = \new_[19808]_  | \new_[19685]_ ;
  assign \new_[19017]_  = ~\new_[937]_ ;
  assign \new_[19018]_  = ~\new_[19333]_ ;
  assign \new_[19019]_  = ~\new_[19292]_ ;
  assign \new_[19020]_  = \new_[19348]_ ;
  assign \new_[19021]_  = ~\new_[20842]_ ;
  assign \new_[19022]_  = ~\new_[21142]_ ;
  assign \new_[19023]_  = ~\new_[19390]_ ;
  assign \new_[19024]_  = ~\new_[19432]_ ;
  assign \new_[19025]_  = ~\new_[19673]_ ;
  assign \new_[19026]_  = ~\new_[19293]_ ;
  assign \new_[19027]_  = ~\new_[18542]_  | ~\new_[21328]_ ;
  assign \new_[19028]_  = ~\new_[20903]_ ;
  assign \new_[19029]_  = ~\new_[19695]_ ;
  assign \new_[19030]_  = ~\new_[19534]_ ;
  assign \new_[19031]_  = ~\new_[995]_ ;
  assign \new_[19032]_  = ~\new_[19442]_ ;
  assign \new_[19033]_  = ~\new_[19279]_ ;
  assign \new_[19034]_  = ~\new_[19712]_  & ~\new_[21545]_ ;
  assign \new_[19035]_  = \new_[19303]_ ;
  assign \new_[19036]_  = ~\new_[19375]_ ;
  assign \new_[19037]_  = ~\new_[19395]_ ;
  assign \new_[19038]_  = ~\new_[19668]_  | ~\new_[19566]_ ;
  assign \new_[19039]_  = ~\new_[21404]_ ;
  assign \new_[19040]_  = ~\new_[19367]_ ;
  assign \new_[19041]_  = ~\new_[999]_ ;
  assign \new_[19042]_  = ~\new_[20491]_ ;
  assign \new_[19043]_  = ~\new_[19287]_ ;
  assign \new_[19044]_  = ~\new_[19510]_ ;
  assign \new_[19045]_  = ~\new_[19547]_ ;
  assign \new_[19046]_  = ~\new_[19641]_  | ~\new_[19654]_ ;
  assign \new_[19047]_  = ~\new_[19324]_ ;
  assign \new_[19048]_  = \new_[19342]_ ;
  assign \new_[19049]_  = ~\new_[19318]_ ;
  assign \new_[19050]_  = ~\new_[19486]_ ;
  assign \new_[19051]_  = ~\new_[19418]_ ;
  assign \new_[19052]_  = ~\new_[19289]_ ;
  assign \new_[19053]_  = ~\new_[19392]_ ;
  assign \new_[19054]_  = ~\new_[19433]_ ;
  assign \new_[19055]_  = ~\new_[19310]_ ;
  assign \new_[19056]_  = ~\new_[19542]_ ;
  assign \new_[19057]_  = ~\new_[19688]_  | ~\new_[19730]_ ;
  assign \new_[19058]_  = ~\new_[20497]_  | ~\new_[19573]_ ;
  assign \new_[19059]_  = ~\new_[17796]_ ;
  assign \new_[19060]_  = ~\new_[20497]_  & ~\new_[19573]_ ;
  assign \new_[19061]_  = ~\new_[19297]_ ;
  assign \new_[19062]_  = ~\new_[19712]_  & ~\new_[21526]_ ;
  assign \new_[19063]_  = ~\new_[19637]_  & ~\new_[19621]_ ;
  assign \new_[19064]_  = ~\new_[20686]_ ;
  assign \new_[19065]_  = ~\new_[19514]_ ;
  assign \new_[19066]_  = ~\new_[19114]_ ;
  assign \new_[19067]_  = ~\new_[19692]_  & ~\new_[21583]_ ;
  assign \new_[19068]_  = ~\new_[21165]_ ;
  assign \new_[19069]_  = ~\new_[19307]_ ;
  assign \new_[19070]_  = ~\new_[19578]_ ;
  assign \new_[19071]_  = ~\new_[19384]_ ;
  assign \new_[19072]_  = ~\new_[19384]_ ;
  assign \new_[19073]_  = \new_[19941]_  | \new_[19758]_ ;
  assign \new_[19074]_  = \new_[19465]_ ;
  assign \new_[19075]_  = ~\new_[19671]_  & ~\new_[19808]_ ;
  assign \new_[19076]_  = \new_[19624]_  & \new_[19746]_ ;
  assign \new_[19077]_  = ~n3423;
  assign \new_[19078]_  = ~\new_[19757]_  | ~\new_[19609]_ ;
  assign \new_[19079]_  = ~\new_[1134]_ ;
  assign \new_[19080]_  = ~\new_[19321]_ ;
  assign \new_[19081]_  = \new_[19516]_ ;
  assign \new_[19082]_  = ~\new_[19423]_ ;
  assign \new_[19083]_  = ~\new_[19410]_ ;
  assign \new_[19084]_  = ~\new_[19460]_ ;
  assign \new_[19085]_  = ~\new_[19432]_ ;
  assign \new_[19086]_  = ~\new_[19488]_ ;
  assign \new_[19087]_  = ~\new_[19526]_ ;
  assign \new_[19088]_  = ~\new_[19029]_ ;
  assign \new_[19089]_  = ~\new_[19466]_ ;
  assign \new_[19090]_  = ~\new_[19468]_ ;
  assign \new_[19091]_  = ~\new_[19493]_ ;
  assign \new_[19092]_  = ~\new_[19534]_ ;
  assign \new_[19093]_  = ~\new_[20498]_ ;
  assign \new_[19094]_  = ~\new_[1089]_ ;
  assign \new_[19095]_  = ~\new_[20486]_ ;
  assign \new_[19096]_  = ~\new_[19362]_ ;
  assign \new_[19097]_  = ~\new_[19510]_ ;
  assign \new_[19098]_  = ~\new_[19419]_ ;
  assign \new_[19099]_  = ~\new_[19428]_ ;
  assign \new_[19100]_  = ~\new_[19390]_ ;
  assign \new_[19101]_  = ~\new_[1619]_ ;
  assign \new_[19102]_  = ~\new_[19491]_ ;
  assign \new_[19103]_  = ~\new_[21115]_ ;
  assign \new_[19104]_  = ~\new_[19390]_ ;
  assign \new_[19105]_  = ~\new_[19478]_ ;
  assign \new_[19106]_  = \new_[20486]_ ;
  assign \new_[19107]_  = ~\new_[19559]_ ;
  assign \new_[19108]_  = ~\new_[19744]_  & ~\new_[19629]_ ;
  assign \new_[19109]_  = ~\new_[19755]_  | ~\new_[19715]_ ;
  assign \new_[19110]_  = ~\new_[19285]_ ;
  assign \new_[19111]_  = ~\new_[19389]_ ;
  assign \new_[19112]_  = \new_[19553]_  | \new_[19665]_ ;
  assign \new_[19113]_  = ~\new_[19773]_  & ~\new_[19583]_ ;
  assign \new_[19114]_  = ~\new_[19555]_ ;
  assign \new_[19115]_  = ~\new_[2295]_ ;
  assign \new_[19116]_  = ~\new_[21097]_ ;
  assign \new_[19117]_  = ~\new_[19427]_ ;
  assign \new_[19118]_  = ~\new_[19394]_ ;
  assign \new_[19119]_  = ~\new_[19566]_  & ~\new_[19668]_ ;
  assign \new_[19120]_  = ~\new_[20513]_ ;
  assign \new_[19121]_  = ~\new_[1343]_ ;
  assign \new_[19122]_  = ~\new_[19342]_ ;
  assign \new_[19123]_  = ~\new_[19513]_ ;
  assign \new_[19124]_  = ~\new_[1187]_ ;
  assign \new_[19125]_  = ~\new_[19745]_  | ~\new_[2298]_ ;
  assign \new_[19126]_  = ~\new_[19706]_  & ~\new_[20167]_ ;
  assign \new_[19127]_  = \new_[19390]_ ;
  assign \new_[19128]_  = ~\new_[19689]_  | ~\new_[19568]_ ;
  assign \new_[19129]_  = ~\new_[20300]_  & ~\new_[19556]_ ;
  assign \new_[19130]_  = ~\new_[19317]_ ;
  assign \new_[19131]_  = ~\new_[19683]_  & ~\new_[21660]_ ;
  assign \new_[19132]_  = ~\new_[19429]_ ;
  assign \new_[19133]_  = ~\new_[19400]_ ;
  assign \new_[19134]_  = ~\new_[19521]_ ;
  assign \new_[19135]_  = \new_[19577]_  & \new_[21583]_ ;
  assign \new_[19136]_  = ~\new_[19444]_ ;
  assign \new_[19137]_  = ~\new_[19730]_  & ~\new_[19582]_ ;
  assign \new_[19138]_  = ~\new_[19376]_  & ~\new_[19746]_ ;
  assign \new_[19139]_  = ~\new_[20870]_ ;
  assign \new_[19140]_  = ~\new_[19311]_ ;
  assign \new_[19141]_  = \new_[19612]_  | \new_[19754]_ ;
  assign \new_[19142]_  = ~\new_[19315]_ ;
  assign \new_[19143]_  = \new_[1347]_  ^ \new_[1513]_ ;
  assign \new_[19144]_  = ~\new_[21395]_ ;
  assign \new_[19145]_  = ~\new_[20842]_ ;
  assign \new_[19146]_  = ~\new_[19348]_ ;
  assign \new_[19147]_  = ~\new_[20171]_ ;
  assign \new_[19148]_  = ~\new_[19337]_ ;
  assign \new_[19149]_  = ~\new_[19538]_ ;
  assign \new_[19150]_  = ~\new_[19421]_ ;
  assign \new_[19151]_  = ~\new_[19469]_ ;
  assign \new_[19152]_  = ~\new_[19331]_ ;
  assign \new_[19153]_  = ~\new_[19543]_ ;
  assign \new_[19154]_  = ~\new_[19351]_ ;
  assign \new_[19155]_  = ~\new_[2302]_  & ~\new_[19697]_ ;
  assign \new_[19156]_  = ~\new_[19279]_ ;
  assign \new_[19157]_  = ~\new_[19537]_ ;
  assign \new_[19158]_  = ~\new_[19408]_ ;
  assign \new_[19159]_  = ~\new_[19501]_ ;
  assign \new_[19160]_  = ~\new_[19393]_ ;
  assign \new_[19161]_  = ~\new_[1006]_ ;
  assign \new_[19162]_  = ~\new_[19500]_ ;
  assign \new_[19163]_  = ~\new_[19529]_ ;
  assign \new_[19164]_  = ~\new_[19601]_  & ~\new_[19701]_ ;
  assign \new_[19165]_  = ~\new_[19368]_ ;
  assign \new_[19166]_  = ~\new_[19335]_ ;
  assign \new_[19167]_  = ~\new_[19668]_  & ~\new_[19594]_ ;
  assign \new_[19168]_  = ~\new_[19321]_ ;
  assign \new_[19169]_  = ~\new_[19568]_  | ~\new_[20845]_ ;
  assign \new_[19170]_  = ~\new_[944]_ ;
  assign \new_[19171]_  = \new_[21560]_  | \new_[19664]_ ;
  assign \new_[19172]_  = ~\new_[19639]_  | ~\new_[19722]_ ;
  assign \new_[19173]_  = ~\new_[20171]_ ;
  assign \new_[19174]_  = ~\new_[19328]_ ;
  assign \new_[19175]_  = ~\new_[2346]_ ;
  assign \new_[19176]_  = ~\new_[19432]_ ;
  assign \new_[19177]_  = ~\new_[19288]_ ;
  assign \new_[19178]_  = \new_[19568]_  | \new_[20845]_ ;
  assign \new_[19179]_  = ~\new_[954]_ ;
  assign \new_[19180]_  = ~\new_[19386]_ ;
  assign \new_[19181]_  = ~\new_[19380]_ ;
  assign \new_[19182]_  = ~\new_[21402]_ ;
  assign \new_[19183]_  = ~\new_[19347]_ ;
  assign \new_[19184]_  = ~\new_[19654]_ ;
  assign \new_[19185]_  = ~\new_[19656]_  & ~\new_[19572]_ ;
  assign \new_[19186]_  = ~\new_[19511]_ ;
  assign \new_[19187]_  = ~\new_[19505]_ ;
  assign \new_[19188]_  = ~\new_[19388]_ ;
  assign \new_[19189]_  = ~\new_[19392]_ ;
  assign \new_[19190]_  = ~\new_[19471]_ ;
  assign \new_[19191]_  = ~\new_[19524]_ ;
  assign \new_[19192]_  = ~\new_[19373]_ ;
  assign \new_[19193]_  = ~\new_[19644]_  | ~\new_[19777]_ ;
  assign \new_[19194]_  = ~\new_[19356]_ ;
  assign \new_[19195]_  = ~\new_[19323]_ ;
  assign \new_[19196]_  = ~\new_[19432]_ ;
  assign \new_[19197]_  = ~\new_[19295]_ ;
  assign \new_[19198]_  = ~\new_[19778]_ ;
  assign \new_[19199]_  = \new_[19779]_  & \new_[19664]_ ;
  assign \new_[19200]_  = ~\new_[19447]_ ;
  assign \new_[19201]_  = ~\new_[19347]_ ;
  assign \new_[19202]_  = ~\new_[1080]_ ;
  assign \new_[19203]_  = ~\new_[19408]_ ;
  assign \new_[19204]_  = ~\new_[19404]_ ;
  assign \new_[19205]_  = ~\new_[19526]_ ;
  assign \new_[19206]_  = ~\new_[2295]_ ;
  assign \new_[19207]_  = ~\new_[19512]_ ;
  assign \new_[19208]_  = ~\new_[19384]_ ;
  assign \new_[19209]_  = ~\new_[19465]_ ;
  assign \new_[19210]_  = ~\new_[20238]_ ;
  assign \new_[19211]_  = ~\new_[19526]_ ;
  assign \new_[19212]_  = ~\new_[19778]_ ;
  assign \new_[19213]_  = ~\new_[19762]_ ;
  assign \new_[19214]_  = ~\new_[19403]_ ;
  assign \new_[19215]_  = ~\new_[19349]_ ;
  assign \new_[19216]_  = ~\new_[19461]_ ;
  assign \new_[19217]_  = ~\new_[19460]_ ;
  assign \new_[19218]_  = ~\new_[19533]_ ;
  assign \new_[19219]_  = ~\new_[19401]_ ;
  assign \new_[19220]_  = ~\new_[19331]_ ;
  assign \new_[19221]_  = ~\new_[19557]_  | ~\new_[19583]_ ;
  assign \new_[19222]_  = \new_[19620]_  & \new_[19674]_ ;
  assign \new_[19223]_  = ~\new_[19771]_  | ~\new_[1354]_ ;
  assign \new_[19224]_  = ~\new_[19375]_ ;
  assign \new_[19225]_  = ~\new_[19498]_ ;
  assign \new_[19226]_  = ~\new_[19274]_ ;
  assign \new_[19227]_  = ~\new_[19365]_ ;
  assign \new_[19228]_  = ~\new_[19456]_  & ~\new_[19697]_ ;
  assign \new_[19229]_  = ~\new_[1039]_ ;
  assign \new_[19230]_  = ~\new_[19764]_  & ~\new_[19777]_ ;
  assign \new_[19231]_  = ~\new_[19402]_ ;
  assign \new_[19232]_  = ~\new_[21305]_  & ~\new_[19809]_ ;
  assign \new_[19233]_  = ~\new_[1006]_ ;
  assign \new_[19234]_  = ~\new_[19584]_  & ~\new_[19670]_ ;
  assign \new_[19235]_  = ~\new_[19745]_  | ~\new_[19608]_ ;
  assign \new_[19236]_  = ~\new_[991]_ ;
  assign \new_[19237]_  = ~\new_[19327]_ ;
  assign \new_[19238]_  = ~\new_[19489]_ ;
  assign \new_[19239]_  = ~\new_[19440]_ ;
  assign \new_[19240]_  = ~\new_[19519]_ ;
  assign \new_[19241]_  = ~\new_[20704]_  & ~\new_[21513]_ ;
  assign \new_[19242]_  = ~\new_[1026]_ ;
  assign \new_[19243]_  = \new_[1084]_ ;
  assign \new_[19244]_  = ~\new_[19384]_ ;
  assign \new_[19245]_  = ~\new_[19484]_ ;
  assign \new_[19246]_  = ~\new_[19276]_ ;
  assign \new_[19247]_  = ~\new_[19491]_ ;
  assign \new_[19248]_  = ~\new_[19757]_  | ~\new_[19685]_ ;
  assign \new_[19249]_  = ~\new_[19361]_ ;
  assign \new_[19250]_  = ~\new_[19771]_  & ~\new_[19669]_ ;
  assign \new_[19251]_  = ~\new_[1002]_ ;
  assign \new_[19252]_  = ~\new_[19678]_  & ~\new_[21517]_ ;
  assign \new_[19253]_  = ~\new_[19471]_ ;
  assign \new_[19254]_  = ~\new_[19420]_ ;
  assign \new_[19255]_  = \new_[19301]_  | \new_[19697]_ ;
  assign \new_[19256]_  = ~\new_[19475]_ ;
  assign \new_[19257]_  = ~\new_[984]_ ;
  assign \new_[19258]_  = ~\new_[21635]_  | ~\new_[20927]_ ;
  assign \new_[19259]_  = ~\new_[959]_ ;
  assign \new_[19260]_  = \new_[19941]_  & \new_[19758]_ ;
  assign \new_[19261]_  = ~\new_[19404]_ ;
  assign \new_[19262]_  = ~\new_[19418]_ ;
  assign \new_[19263]_  = ~\new_[19671]_  | ~\new_[19685]_ ;
  assign \new_[19264]_  = ~\new_[20300]_  | ~\new_[1079]_ ;
  assign \new_[19265]_  = ~\new_[19289]_ ;
  assign \new_[19266]_  = ~\new_[19320]_ ;
  assign \new_[19267]_  = ~\new_[19344]_ ;
  assign \new_[19268]_  = ~\new_[19499]_ ;
  assign \new_[19269]_  = ~\new_[19443]_ ;
  assign \new_[19270]_  = ~\new_[19356]_ ;
  assign \new_[19271]_  = ~\new_[960]_ ;
  assign \new_[19272]_  = ~\new_[19302]_ ;
  assign \new_[19273]_  = ~\new_[20743]_ ;
  assign \new_[19274]_  = \new_[19668]_ ;
  assign \new_[19275]_  = ~\new_[19790]_ ;
  assign \new_[19276]_  = \new_[20970]_ ;
  assign \new_[19277]_  = ~\new_[923]_ ;
  assign \new_[19278]_  = ~\new_[19580]_ ;
  assign \new_[19279]_  = ~\new_[19738]_ ;
  assign \new_[19280]_  = \new_[19646]_ ;
  assign \new_[19281]_  = ~\new_[19754]_ ;
  assign \new_[19282]_  = ~\new_[19641]_ ;
  assign \new_[19283]_  = ~\new_[19649]_ ;
  assign \new_[19284]_  = ~\new_[19640]_ ;
  assign \new_[19285]_  = ~\new_[927]_ ;
  assign \new_[19286]_  = ~\new_[19678]_ ;
  assign \new_[19287]_  = \new_[19763]_ ;
  assign \new_[19288]_  = ~\new_[1607]_ ;
  assign \new_[19289]_  = ~\new_[19650]_ ;
  assign \new_[19290]_  = ~\new_[1242]_ ;
  assign \new_[19291]_  = ~\new_[19808]_ ;
  assign \new_[19292]_  = ~\new_[19741]_ ;
  assign \new_[19293]_  = ~\new_[20170]_ ;
  assign \new_[19294]_  = ~\new_[19548]_ ;
  assign \new_[19295]_  = ~\new_[19734]_ ;
  assign \new_[19296]_  = ~\new_[19604]_ ;
  assign \new_[19297]_  = ~\new_[19779]_ ;
  assign \new_[19298]_  = ~\new_[1242]_ ;
  assign \new_[19299]_  = ~\new_[19798]_ ;
  assign \new_[19300]_  = ~\new_[19236]_ ;
  assign \new_[19301]_  = ~\new_[2302]_ ;
  assign \new_[19302]_  = ~\new_[20590]_ ;
  assign \new_[19303]_  = \new_[19596]_ ;
  assign \new_[19304]_  = ~\new_[21205]_ ;
  assign \new_[19305]_  = ~\new_[1288]_ ;
  assign \new_[19306]_  = ~\new_[1510]_ ;
  assign \new_[19307]_  = ~\new_[19777]_ ;
  assign \new_[19308]_  = ~\new_[19771]_ ;
  assign \new_[19309]_  = ~\new_[19611]_ ;
  assign \new_[19310]_  = ~\new_[20589]_ ;
  assign \new_[19311]_  = ~\new_[19706]_ ;
  assign \new_[19312]_  = ~\new_[12134]_  & ~\new_[10818]_ ;
  assign \new_[19313]_  = ~\new_[19586]_ ;
  assign \new_[19314]_  = ~\new_[19672]_ ;
  assign \new_[19315]_  = ~\new_[19757]_ ;
  assign \new_[19316]_  = ~\new_[20464]_ ;
  assign \new_[19317]_  = ~\new_[20241]_ ;
  assign \new_[19318]_  = ~\new_[19702]_ ;
  assign \new_[19319]_  = ~\new_[1242]_ ;
  assign \new_[19320]_  = ~\new_[19711]_ ;
  assign \new_[19321]_  = ~\new_[19586]_ ;
  assign \new_[19322]_  = ~\new_[19619]_ ;
  assign \new_[19323]_  = ~\new_[1878]_ ;
  assign \new_[19324]_  = ~\new_[19670]_ ;
  assign \new_[19325]_  = ~\new_[1346]_ ;
  assign \new_[19326]_  = ~\new_[1025]_ ;
  assign \new_[19327]_  = ~\new_[1134]_ ;
  assign \new_[19328]_  = ~\new_[19629]_ ;
  assign \new_[19329]_  = ~\new_[19777]_ ;
  assign \new_[19330]_  = ~\new_[19577]_ ;
  assign \new_[19331]_  = ~\new_[19650]_ ;
  assign \new_[19332]_  = ~\new_[19594]_ ;
  assign \new_[19333]_  = ~\new_[19750]_ ;
  assign \new_[19334]_  = ~\new_[20645]_ ;
  assign \new_[19335]_  = ~\new_[19762]_ ;
  assign \new_[19336]_  = ~\new_[1025]_ ;
  assign \new_[19337]_  = ~\new_[922]_ ;
  assign \new_[19338]_  = ~\new_[19649]_ ;
  assign \new_[19339]_  = ~\new_[19615]_ ;
  assign \new_[19340]_  = ~\new_[19765]_ ;
  assign \new_[19341]_  = ~\new_[946]_ ;
  assign \new_[19342]_  = ~\new_[927]_ ;
  assign \new_[19343]_  = ~\new_[19561]_ ;
  assign \new_[19344]_  = ~\new_[19809]_ ;
  assign \new_[19345]_  = \new_[19705]_ ;
  assign \new_[19346]_  = ~\new_[19668]_ ;
  assign \new_[19347]_  = ~\new_[19580]_ ;
  assign \new_[19348]_  = \new_[19607]_ ;
  assign \new_[19349]_  = ~\new_[19620]_ ;
  assign \new_[19350]_  = ~\new_[19567]_ ;
  assign \new_[19351]_  = ~\new_[21115]_ ;
  assign \new_[19352]_  = ~\new_[19609]_ ;
  assign \new_[19353]_  = ~\new_[19645]_ ;
  assign \new_[19354]_  = \new_[19670]_ ;
  assign \new_[19355]_  = ~\new_[1656]_ ;
  assign \new_[19356]_  = ~\new_[19801]_ ;
  assign \new_[19357]_  = ~\new_[19798]_ ;
  assign \new_[19358]_  = ~\new_[19729]_ ;
  assign \new_[19359]_  = ~\new_[20751]_ ;
  assign \new_[19360]_  = ~\new_[19589]_ ;
  assign \new_[19361]_  = ~\new_[20845]_ ;
  assign \new_[19362]_  = ~\new_[19617]_ ;
  assign \new_[19363]_  = ~\new_[19649]_ ;
  assign \new_[19364]_  = \new_[19656]_ ;
  assign \new_[19365]_  = ~\new_[19656]_ ;
  assign \new_[19366]_  = ~\new_[2295]_ ;
  assign \new_[19367]_  = \new_[19791]_ ;
  assign \new_[19368]_  = ~\new_[19678]_ ;
  assign \new_[19369]_  = ~\new_[19758]_ ;
  assign \new_[19370]_  = ~\new_[20497]_ ;
  assign \new_[19371]_  = ~\new_[19649]_ ;
  assign \new_[19372]_  = ~\new_[19649]_ ;
  assign \new_[19373]_  = ~\new_[19675]_ ;
  assign \new_[19374]_  = ~\new_[2295]_ ;
  assign \new_[19375]_  = ~\new_[20865]_ ;
  assign \new_[19376]_  = ~\new_[1001]_ ;
  assign \new_[19377]_  = ~\new_[19547]_ ;
  assign \new_[19378]_  = ~\new_[19659]_ ;
  assign \new_[19379]_  = ~\new_[19778]_ ;
  assign \new_[19380]_  = ~\new_[19664]_ ;
  assign \new_[19381]_  = ~\new_[1081]_ ;
  assign \new_[19382]_  = ~\new_[19587]_ ;
  assign \new_[19383]_  = ~\new_[19649]_ ;
  assign \new_[19384]_  = ~\new_[19687]_ ;
  assign \new_[19385]_  = \new_[19376]_ ;
  assign \new_[19386]_  = ~\new_[19804]_ ;
  assign \new_[19387]_  = ~\new_[1667]_ ;
  assign \new_[19388]_  = ~\new_[21166]_ ;
  assign \new_[19389]_  = ~\new_[19764]_ ;
  assign \new_[19390]_  = ~\new_[19725]_ ;
  assign \new_[19391]_  = ~\new_[19718]_ ;
  assign \new_[19392]_  = ~\new_[19643]_ ;
  assign \new_[19393]_  = \new_[19609]_ ;
  assign \new_[19394]_  = ~\new_[19655]_ ;
  assign \new_[19395]_  = ~\new_[19648]_ ;
  assign \new_[19396]_  = ~\new_[19691]_ ;
  assign \new_[19397]_  = ~\new_[19563]_ ;
  assign \new_[19398]_  = ~\new_[19647]_ ;
  assign \new_[19399]_  = ~\new_[19621]_ ;
  assign \new_[19400]_  = \new_[946]_ ;
  assign \new_[19401]_  = ~\new_[20746]_ ;
  assign \new_[19402]_  = ~\new_[19743]_ ;
  assign \new_[19403]_  = ~\new_[19681]_ ;
  assign \new_[19404]_  = ~\new_[19381]_ ;
  assign \new_[19405]_  = ~\new_[19550]_ ;
  assign \new_[19406]_  = ~\new_[19674]_ ;
  assign \new_[19407]_  = ~\new_[19697]_ ;
  assign \new_[19408]_  = \new_[1242]_ ;
  assign \new_[19409]_  = ~\new_[19627]_ ;
  assign \new_[19410]_  = ~\new_[931]_ ;
  assign \new_[19411]_  = \new_[19756]_ ;
  assign \new_[19412]_  = ~\new_[19660]_ ;
  assign \new_[19413]_  = ~\new_[19728]_ ;
  assign \new_[19414]_  = ~\new_[19649]_ ;
  assign \new_[19415]_  = ~\new_[19649]_ ;
  assign \new_[19416]_  = ~\new_[924]_ ;
  assign \new_[19417]_  = ~\new_[19670]_ ;
  assign \new_[19418]_  = ~\new_[19709]_ ;
  assign \new_[19419]_  = ~\new_[19676]_ ;
  assign \new_[19420]_  = ~\new_[19734]_ ;
  assign \new_[19421]_  = ~\new_[21397]_ ;
  assign \new_[19422]_  = ~\new_[19680]_ ;
  assign \new_[19423]_  = ~\new_[19674]_ ;
  assign \new_[19424]_  = \new_[1025]_ ;
  assign \new_[19425]_  = ~\new_[1242]_ ;
  assign \new_[19426]_  = \new_[21166]_ ;
  assign \new_[19427]_  = ~\new_[19697]_ ;
  assign \new_[19428]_  = ~\new_[925]_ ;
  assign \new_[19429]_  = ~\new_[19607]_ ;
  assign \new_[19430]_  = ~\new_[19629]_ ;
  assign \new_[19431]_  = ~\new_[21325]_ ;
  assign \new_[19432]_  = ~\new_[19663]_ ;
  assign \new_[19433]_  = ~\new_[21422]_ ;
  assign \new_[19434]_  = ~\new_[924]_ ;
  assign \new_[19435]_  = ~\new_[1354]_ ;
  assign \new_[19436]_  = \new_[19687]_ ;
  assign \new_[19437]_  = \new_[19601]_ ;
  assign \new_[19438]_  = ~\new_[2080]_ ;
  assign \new_[19439]_  = ~\new_[19780]_ ;
  assign \new_[19440]_  = ~\new_[19815]_ ;
  assign \new_[19441]_  = ~\new_[19770]_ ;
  assign \new_[19442]_  = ~\new_[19271]_ ;
  assign \new_[19443]_  = \new_[19794]_ ;
  assign \new_[19444]_  = ~\new_[19545]_ ;
  assign \new_[19445]_  = ~\new_[19717]_ ;
  assign \new_[19446]_  = ~\new_[19707]_ ;
  assign \new_[19447]_  = ~\new_[19574]_ ;
  assign \new_[19448]_  = \new_[19696]_ ;
  assign \new_[19449]_  = ~\new_[19722]_ ;
  assign \new_[19450]_  = ~\new_[19559]_ ;
  assign \new_[19451]_  = ~\new_[19649]_ ;
  assign \new_[19452]_  = ~\new_[1243]_ ;
  assign \new_[19453]_  = ~\new_[19694]_ ;
  assign \new_[19454]_  = \new_[19801]_ ;
  assign \new_[19455]_  = ~\new_[19572]_ ;
  assign \new_[19456]_  = ~\new_[2295]_ ;
  assign \new_[19457]_  = ~\new_[19623]_ ;
  assign n3423 = ~\new_[19649]_ ;
  assign \new_[19459]_  = \new_[19643]_ ;
  assign \new_[19460]_  = ~\new_[19746]_ ;
  assign \new_[19461]_  = ~\new_[19745]_ ;
  assign \new_[19462]_  = \new_[19664]_ ;
  assign \new_[19463]_  = ~\new_[19789]_ ;
  assign \new_[19464]_  = \new_[19594]_ ;
  assign \new_[19465]_  = ~\new_[21047]_ ;
  assign \new_[19466]_  = ~\new_[19601]_ ;
  assign \new_[19467]_  = ~\new_[19599]_ ;
  assign \new_[19468]_  = ~\new_[19583]_ ;
  assign \new_[19469]_  = ~\new_[19791]_ ;
  assign \new_[19470]_  = ~\new_[19564]_ ;
  assign \new_[19471]_  = ~\new_[19767]_ ;
  assign \new_[19472]_  = ~\new_[19649]_ ;
  assign \new_[19473]_  = ~\new_[19692]_ ;
  assign \new_[19474]_  = ~\new_[19707]_ ;
  assign \new_[19475]_  = ~\new_[19712]_ ;
  assign \new_[19476]_  = \new_[19752]_ ;
  assign \new_[19477]_  = ~\new_[19679]_ ;
  assign \new_[19478]_  = \new_[19789]_ ;
  assign \new_[19479]_  = ~\new_[19649]_ ;
  assign \new_[19480]_  = ~\new_[19717]_ ;
  assign \new_[19481]_  = ~\new_[19782]_ ;
  assign \new_[19482]_  = ~\new_[20493]_ ;
  assign \new_[19483]_  = ~\new_[1025]_ ;
  assign \new_[19484]_  = \new_[20751]_ ;
  assign \new_[19485]_  = ~\new_[19596]_ ;
  assign \new_[19486]_  = ~\new_[19752]_ ;
  assign \new_[19487]_  = ~\new_[19688]_ ;
  assign \new_[19488]_  = ~\new_[19573]_ ;
  assign \new_[19489]_  = ~\new_[19566]_ ;
  assign \new_[19490]_  = ~\new_[19795]_ ;
  assign \new_[19491]_  = ~\new_[19592]_ ;
  assign \new_[19492]_  = ~\new_[19612]_ ;
  assign \new_[19493]_  = ~\new_[19376]_ ;
  assign \new_[19494]_  = \new_[21305]_ ;
  assign \new_[19495]_  = ~\new_[9578]_  & ~\new_[6746]_ ;
  assign \new_[19496]_  = ~\new_[19649]_ ;
  assign \new_[19497]_  = ~\new_[19649]_ ;
  assign \new_[19498]_  = ~\new_[19643]_ ;
  assign \new_[19499]_  = ~\new_[19568]_ ;
  assign \new_[19500]_  = ~\new_[19597]_ ;
  assign \new_[19501]_  = ~\new_[19743]_ ;
  assign \new_[19502]_  = ~\new_[19561]_ ;
  assign \new_[19503]_  = ~\new_[19641]_ ;
  assign \new_[19504]_  = ~\new_[19751]_ ;
  assign \new_[19505]_  = \new_[19616]_ ;
  assign \new_[19506]_  = \new_[21401]_ ;
  assign \new_[19507]_  = ~\new_[19713]_ ;
  assign \new_[19508]_  = ~\new_[19553]_ ;
  assign \new_[19509]_  = ~\new_[20941]_ ;
  assign \new_[19510]_  = ~\new_[19554]_ ;
  assign \new_[19511]_  = ~\new_[19665]_ ;
  assign \new_[19512]_  = ~\new_[19813]_ ;
  assign \new_[19513]_  = ~\new_[19721]_ ;
  assign \new_[19514]_  = \new_[19572]_ ;
  assign \new_[19515]_  = ~\new_[17156]_  | ~\new_[16511]_ ;
  assign \new_[19516]_  = \new_[19706]_ ;
  assign \new_[19517]_  = ~\new_[19787]_ ;
  assign \new_[19518]_  = \new_[19744]_ ;
  assign \new_[19519]_  = ~\new_[20681]_ ;
  assign \new_[19520]_  = ~\new_[19697]_ ;
  assign \new_[19521]_  = ~\new_[19756]_ ;
  assign \new_[19522]_  = ~\new_[20300]_ ;
  assign \new_[19523]_  = ~\new_[20513]_ ;
  assign \new_[19524]_  = \new_[19546]_ ;
  assign \new_[19525]_  = ~\new_[19941]_ ;
  assign \new_[19526]_  = ~\new_[19622]_ ;
  assign \new_[19527]_  = ~\new_[19751]_ ;
  assign \new_[19528]_  = ~\new_[19780]_ ;
  assign \new_[19529]_  = ~\new_[19277]_ ;
  assign \new_[19530]_  = ~\new_[19748]_ ;
  assign \new_[19531]_  = ~\new_[20100]_ ;
  assign \new_[19532]_  = ~\new_[19636]_ ;
  assign \new_[19533]_  = ~\new_[19584]_ ;
  assign \new_[19534]_  = ~\new_[19574]_ ;
  assign \new_[19535]_  = ~\new_[19728]_ ;
  assign \new_[19536]_  = ~\new_[19740]_ ;
  assign \new_[19537]_  = ~\new_[20789]_ ;
  assign \new_[19538]_  = ~\new_[19652]_ ;
  assign \new_[19539]_  = ~\new_[1134]_ ;
  assign \new_[19540]_  = ~\new_[20452]_ ;
  assign \new_[19541]_  = ~\new_[19730]_ ;
  assign \new_[19542]_  = ~\new_[19744]_ ;
  assign \new_[19543]_  = ~\new_[19742]_ ;
  assign \new_[19544]_  = ~\new_[1240]_ ;
  assign \new_[19545]_  = \new_[1001]_ ;
  assign \new_[19546]_  = ~\new_[1086]_ ;
  assign \new_[19547]_  = ~\new_[1672]_ ;
  assign \new_[19548]_  = ~\new_[948]_ ;
  assign \new_[19549]_  = ~\new_[1290]_ ;
  assign \new_[19550]_  = ~\new_[1928]_ ;
  assign \new_[19551]_  = ~\new_[1666]_ ;
  assign \new_[19552]_  = ~\new_[1341]_ ;
  assign \new_[19553]_  = ~\new_[2296]_ ;
  assign \new_[19554]_  = ~\new_[936]_ ;
  assign \new_[19555]_  = ~\new_[2080]_ ;
  assign \new_[19556]_  = ~\new_[1079]_ ;
  assign \new_[19557]_  = ~\new_[1656]_ ;
  assign \new_[19558]_  = ~\new_[1474]_ ;
  assign \new_[19559]_  = \new_[1029]_ ;
  assign \new_[19560]_  = ~\new_[2344]_ ;
  assign \new_[19561]_  = ~\new_[1928]_ ;
  assign \new_[19562]_  = ~\new_[1506]_ ;
  assign \new_[19563]_  = ~\new_[1519]_ ;
  assign \new_[19564]_  = ~\new_[935]_ ;
  assign \new_[19565]_  = ~\new_[2297]_ ;
  assign \new_[19566]_  = ~\new_[981]_ ;
  assign \new_[19567]_  = ~\new_[2500]_ ;
  assign \new_[19568]_  = ~\new_[939]_ ;
  assign \new_[19569]_  = ~\new_[1350]_ ;
  assign \new_[19570]_  = ~\new_[1419]_ ;
  assign \new_[19571]_  = ~\new_[1088]_ ;
  assign \new_[19572]_  = ~\new_[1031]_ ;
  assign \new_[19573]_  = ~\new_[1046]_ ;
  assign \new_[19574]_  = ~\new_[1024]_ ;
  assign \new_[19575]_  = ~\new_[1868]_ ;
  assign \new_[19576]_  = ~\new_[10818]_ ;
  assign \new_[19577]_  = ~\new_[1036]_ ;
  assign \new_[19578]_  = ~\new_[1879]_ ;
  assign \new_[19579]_  = ~\new_[1291]_ ;
  assign \new_[19580]_  = ~\new_[970]_ ;
  assign \new_[19581]_  = ~\new_[17156]_ ;
  assign \new_[19582]_  = ~\new_[1038]_ ;
  assign \new_[19583]_  = ~\new_[1674]_ ;
  assign \new_[19584]_  = ~\new_[1139]_ ;
  assign \new_[19585]_  = ~\new_[930]_ ;
  assign \new_[19586]_  = ~\new_[1037]_ ;
  assign \new_[19587]_  = ~\new_[1083]_ ;
  assign \new_[19588]_  = ~\new_[1620]_ ;
  assign \new_[19589]_  = ~\new_[1242]_ ;
  assign \new_[19590]_  = ~\new_[2291]_ ;
  assign \new_[19591]_  = ~\new_[2293]_ ;
  assign \new_[19592]_  = ~\new_[1083]_ ;
  assign \new_[19593]_  = ~\new_[1352]_ ;
  assign \new_[19594]_  = ~\new_[945]_ ;
  assign \new_[19595]_  = ~\new_[1424]_ ;
  assign \new_[19596]_  = ~\new_[1078]_ ;
  assign \new_[19597]_  = ~\new_[1136]_ ;
  assign \new_[19598]_  = ~\new_[1671]_ ;
  assign \new_[19599]_  = ~\new_[946]_ ;
  assign \new_[19600]_  = ~\new_[1033]_ ;
  assign \new_[19601]_  = ~\new_[1008]_ ;
  assign \new_[19602]_  = ~\new_[1519]_ ;
  assign \new_[19603]_  = ~\new_[1673]_ ;
  assign \new_[19604]_  = ~\new_[975]_ ;
  assign \new_[19605]_  = ~\new_[1237]_ ;
  assign \new_[19606]_  = ~\new_[1867]_ ;
  assign \new_[19607]_  = ~\new_[942]_ ;
  assign \new_[19608]_  = ~\new_[2298]_ ;
  assign \new_[19609]_  = ~\new_[1425]_ ;
  assign \new_[19610]_  = ~\new_[1929]_ ;
  assign \new_[19611]_  = \new_[1185]_ ;
  assign \new_[19612]_  = ~\new_[1009]_ ;
  assign \new_[19613]_  = ~\new_[997]_ ;
  assign \new_[19614]_  = ~ld;
  assign \new_[19615]_  = ~\new_[1025]_ ;
  assign \new_[19616]_  = ~\new_[2520]_ ;
  assign \new_[19617]_  = ~\new_[951]_ ;
  assign \new_[19618]_  = ~\new_[1351]_ ;
  assign \new_[19619]_  = ~\new_[944]_ ;
  assign \new_[19620]_  = ~\new_[1083]_ ;
  assign \new_[19621]_  = ~\new_[963]_ ;
  assign \new_[19622]_  = ~\new_[1429]_ ;
  assign \new_[19623]_  = ~\new_[984]_ ;
  assign \new_[19624]_  = ~\new_[1001]_ ;
  assign \new_[19625]_  = ~\new_[1087]_ ;
  assign \new_[19626]_  = ~\new_[1719]_ ;
  assign \new_[19627]_  = \new_[992]_ ;
  assign \new_[19628]_  = ~\new_[1239]_ ;
  assign \new_[19629]_  = ~\new_[1034]_ ;
  assign \new_[19630]_  = ~\new_[1431]_ ;
  assign \new_[19631]_  = ~\new_[1433]_ ;
  assign \new_[19632]_  = ~\new_[2079]_ ;
  assign \new_[19633]_  = ~\new_[1662]_ ;
  assign \new_[19634]_  = ~\new_[1342]_ ;
  assign \new_[19635]_  = ~\new_[15851]_ ;
  assign \new_[19636]_  = ~\new_[1607]_ ;
  assign \new_[19637]_  = ~\new_[1002]_ ;
  assign \new_[19638]_  = ~\new_[973]_ ;
  assign \new_[19639]_  = ~\new_[2272]_ ;
  assign \new_[19640]_  = ~\new_[973]_ ;
  assign \new_[19641]_  = \new_[2272]_ ;
  assign \new_[19642]_  = ~\new_[2302]_ ;
  assign \new_[19643]_  = ~\new_[920]_ ;
  assign \new_[19644]_  = ~\new_[962]_ ;
  assign \new_[19645]_  = \new_[951]_ ;
  assign \new_[19646]_  = ~\new_[1865]_ ;
  assign \new_[19647]_  = \new_[998]_ ;
  assign \new_[19648]_  = ~\new_[1078]_ ;
  assign \new_[19649]_  = ~ld;
  assign \new_[19650]_  = ~\new_[947]_ ;
  assign \new_[19651]_  = ~\new_[1426]_ ;
  assign \new_[19652]_  = \new_[963]_ ;
  assign \new_[19653]_  = ~\new_[1039]_ ;
  assign \new_[19654]_  = ~\new_[1870]_ ;
  assign \new_[19655]_  = ~\new_[1511]_ ;
  assign \new_[19656]_  = ~\new_[977]_ ;
  assign \new_[19657]_  = ~\new_[2509]_ ;
  assign \new_[19658]_  = ~\new_[1872]_ ;
  assign \new_[19659]_  = ~\new_[921]_ ;
  assign \new_[19660]_  = \new_[997]_ ;
  assign \new_[19661]_  = ~\new_[1517]_ ;
  assign \new_[19662]_  = ~\new_[1428]_ ;
  assign \new_[19663]_  = ~\new_[929]_ ;
  assign \new_[19664]_  = ~\new_[925]_ ;
  assign \new_[19665]_  = ~\new_[1508]_ ;
  assign \new_[19666]_  = ~\new_[1665]_ ;
  assign \new_[19667]_  = ~\new_[1241]_ ;
  assign \new_[19668]_  = ~\new_[1135]_ ;
  assign \new_[19669]_  = ~\new_[1354]_ ;
  assign \new_[19670]_  = ~\new_[957]_ ;
  assign \new_[19671]_  = ~\new_[1344]_ ;
  assign \new_[19672]_  = ~\new_[1243]_ ;
  assign \new_[19673]_  = ~\new_[2078]_ ;
  assign \new_[19674]_  = ~\new_[931]_ ;
  assign \new_[19675]_  = ~\new_[2302]_ ;
  assign \new_[19676]_  = ~\new_[1864]_ ;
  assign \new_[19677]_  = ~\new_[1509]_ ;
  assign \new_[19678]_  = ~\new_[1042]_ ;
  assign \new_[19679]_  = ~\new_[1002]_ ;
  assign \new_[19680]_  = \new_[1045]_ ;
  assign \new_[19681]_  = ~\new_[925]_ ;
  assign \new_[19682]_  = ~\new_[1349]_ ;
  assign \new_[19683]_  = ~\new_[1035]_ ;
  assign \new_[19684]_  = ~\new_[1866]_ ;
  assign \new_[19685]_  = ~\new_[1185]_ ;
  assign \new_[19686]_  = ~\new_[1516]_ ;
  assign \new_[19687]_  = ~\new_[1085]_ ;
  assign \new_[19688]_  = ~\new_[988]_ ;
  assign \new_[19689]_  = ~\new_[974]_ ;
  assign \new_[19690]_  = ~\new_[1669]_ ;
  assign \new_[19691]_  = ~\new_[1517]_ ;
  assign \new_[19692]_  = ~\new_[1036]_ ;
  assign \new_[19693]_  = ~\new_[1675]_ ;
  assign \new_[19694]_  = ~\new_[1039]_ ;
  assign \new_[19695]_  = ~\new_[1009]_ ;
  assign \new_[19696]_  = ~\new_[959]_ ;
  assign \new_[19697]_  = ~\new_[1188]_ ;
  assign \new_[19698]_  = ~\new_[1421]_ ;
  assign \new_[19699]_  = ~\new_[1862]_ ;
  assign \new_[19700]_  = ~\new_[1348]_ ;
  assign \new_[19701]_  = ~\new_[1045]_ ;
  assign \new_[19702]_  = ~\new_[999]_ ;
  assign \new_[19703]_  = ~\new_[1139]_ ;
  assign \new_[19704]_  = ~\new_[1432]_ ;
  assign \new_[19705]_  = ~\new_[1720]_ ;
  assign \new_[19706]_  = ~\new_[972]_ ;
  assign \new_[19707]_  = \new_[934]_ ;
  assign \new_[19708]_  = ~\new_[1518]_ ;
  assign \new_[19709]_  = ~\new_[1026]_ ;
  assign \new_[19710]_  = ~\new_[1422]_ ;
  assign \new_[19711]_  = ~\new_[1029]_ ;
  assign \new_[19712]_  = ~\new_[989]_ ;
  assign \new_[19713]_  = ~\new_[2295]_ ;
  assign \new_[19714]_  = ~\new_[1658]_ ;
  assign \new_[19715]_  = ~\new_[1425]_ ;
  assign \new_[19716]_  = ~\new_[1664]_ ;
  assign \new_[19717]_  = ~\new_[1878]_ ;
  assign \new_[19718]_  = ~\new_[1675]_ ;
  assign \new_[19719]_  = ~\new_[974]_ ;
  assign \new_[19720]_  = ~\new_[2300]_ ;
  assign \new_[19721]_  = ~\new_[1354]_ ;
  assign \new_[19722]_  = ~\new_[1870]_ ;
  assign \new_[19723]_  = ~rst;
  assign \new_[19724]_  = ~\new_[1672]_ ;
  assign \new_[19725]_  = ~\new_[1044]_ ;
  assign \new_[19726]_  = ~\new_[2288]_ ;
  assign \new_[19727]_  = ~\new_[1607]_ ;
  assign \new_[19728]_  = \new_[974]_ ;
  assign \new_[19729]_  = ~\new_[931]_ ;
  assign \new_[19730]_  = ~\new_[1086]_ ;
  assign \new_[19731]_  = ~\new_[1877]_ ;
  assign \new_[19732]_  = ~\new_[1921]_ ;
  assign \new_[19733]_  = ~\new_[2301]_ ;
  assign \new_[19734]_  = ~\new_[961]_ ;
  assign \new_[19735]_  = ~\new_[1739]_ ;
  assign \new_[19736]_  = ~\new_[926]_ ;
  assign \new_[19737]_  = ~\new_[1744]_ ;
  assign \new_[19738]_  = ~\new_[1434]_ ;
  assign \new_[19739]_  = ~\new_[1430]_ ;
  assign \new_[19740]_  = ~\new_[1039]_ ;
  assign \new_[19741]_  = ~\new_[936]_ ;
  assign \new_[19742]_  = ~\new_[1672]_ ;
  assign \new_[19743]_  = ~\new_[965]_ ;
  assign \new_[19744]_  = ~\new_[983]_ ;
  assign \new_[19745]_  = ~\new_[1869]_ ;
  assign \new_[19746]_  = ~\new_[1005]_ ;
  assign \new_[19747]_  = ~\new_[2294]_ ;
  assign \new_[19748]_  = ~\new_[922]_ ;
  assign \new_[19749]_  = ~\new_[1661]_ ;
  assign \new_[19750]_  = ~\new_[955]_ ;
  assign \new_[19751]_  = \new_[1025]_ ;
  assign \new_[19752]_  = ~\new_[955]_ ;
  assign \new_[19753]_  = ~\new_[1668]_ ;
  assign \new_[19754]_  = ~\new_[934]_ ;
  assign \new_[19755]_  = ~\new_[1344]_ ;
  assign \new_[19756]_  = ~\new_[1007]_ ;
  assign \new_[19757]_  = \new_[1344]_ ;
  assign \new_[19758]_  = ~\new_[947]_ ;
  assign \new_[19759]_  = ~\new_[9578]_ ;
  assign \new_[19760]_  = ~\new_[1477]_ ;
  assign \new_[19761]_  = ~\new_[1670]_ ;
  assign \new_[19762]_  = \new_[1511]_ ;
  assign \new_[19763]_  = ~\new_[1874]_ ;
  assign \new_[19764]_  = ~\new_[962]_ ;
  assign \new_[19765]_  = ~\new_[1517]_ ;
  assign \new_[19766]_  = ~\new_[1238]_ ;
  assign \new_[19767]_  = ~\new_[1508]_ ;
  assign \new_[19768]_  = ~\new_[1507]_ ;
  assign \new_[19769]_  = ~\new_[945]_ ;
  assign \new_[19770]_  = ~\new_[999]_ ;
  assign \new_[19771]_  = ~\new_[2298]_ ;
  assign \new_[19772]_  = ~\new_[1004]_ ;
  assign \new_[19773]_  = ~\new_[1656]_ ;
  assign \new_[19774]_  = ~\new_[1420]_ ;
  assign \new_[19775]_  = ~\new_[1289]_ ;
  assign \new_[19776]_  = ~\new_[1353]_ ;
  assign \new_[19777]_  = ~\new_[1047]_ ;
  assign \new_[19778]_  = \new_[1136]_ ;
  assign \new_[19779]_  = ~\new_[924]_ ;
  assign \new_[19780]_  = ~\new_[2500]_ ;
  assign \new_[19781]_  = ~\new_[1427]_ ;
  assign \new_[19782]_  = ~\new_[974]_ ;
  assign \new_[19783]_  = ~\new_[1861]_ ;
  assign \new_[19784]_  = ~\new_[1418]_ ;
  assign \new_[19785]_  = ~\new_[1001]_ ;
  assign \new_[19786]_  = ~\new_[932]_ ;
  assign \new_[19787]_  = ~\new_[1026]_ ;
  assign \new_[19788]_  = ~\new_[998]_ ;
  assign \new_[19789]_  = ~\new_[945]_ ;
  assign \new_[19790]_  = \new_[925]_ ;
  assign \new_[19791]_  = ~\new_[992]_ ;
  assign \new_[19792]_  = ~\new_[1659]_ ;
  assign \new_[19793]_  = ~\new_[1863]_ ;
  assign \new_[19794]_  = \new_[948]_ ;
  assign \new_[19795]_  = ~\new_[932]_ ;
  assign \new_[19796]_  = ~\new_[1875]_ ;
  assign \new_[19797]_  = ~\new_[1663]_ ;
  assign \new_[19798]_  = \new_[1080]_ ;
  assign \new_[19799]_  = ~\new_[1345]_ ;
  assign \new_[19800]_  = ~\new_[1417]_ ;
  assign \new_[19801]_  = ~\new_[1022]_ ;
  assign \new_[19802]_  = ~\new_[2511]_ ;
  assign \new_[19803]_  = ~\new_[1878]_ ;
  assign \new_[19804]_  = \new_[1022]_ ;
  assign \new_[19805]_  = ~\new_[1186]_ ;
  assign \new_[19806]_  = ~\new_[965]_ ;
  assign \new_[19807]_  = ~\new_[964]_ ;
  assign \new_[19808]_  = ~\new_[1425]_ ;
  assign \new_[19809]_  = ~\new_[1035]_ ;
  assign \new_[19810]_  = ~\new_[1637]_ ;
  assign \new_[19811]_  = ~\new_[1515]_ ;
  assign \new_[19812]_  = ~\new_[958]_ ;
  assign \new_[19813]_  = ~\new_[954]_ ;
  assign \new_[19814]_  = ~\new_[1660]_ ;
  assign \new_[19815]_  = ~\new_[2295]_ ;
  assign \new_[19816]_  = ~\new_[979]_ ;
  assign \new_[19817]_  = \new_[19818]_ ;
  assign \new_[19818]_  = \new_[21210]_ ;
  assign \new_[19819]_  = ~\new_[21210]_ ;
  assign \new_[19820]_  = ~\new_[21210]_ ;
  assign \new_[19821]_  = ~\new_[19822]_ ;
  assign \new_[19822]_  = \new_[19824]_ ;
  assign \new_[19823]_  = ~\new_[19824]_ ;
  assign \new_[19824]_  = ~\new_[18279]_ ;
  assign \new_[19825]_  = ~\new_[5192]_  | ~\new_[19826]_ ;
  assign \new_[19826]_  = ~\new_[9462]_  & ~\new_[7352]_ ;
  assign \new_[19827]_  = ~\new_[5333]_  | ~\new_[19828]_ ;
  assign \new_[19828]_  = \new_[7722]_  & \new_[13653]_ ;
  assign \new_[19829]_  = ~\new_[19833]_  | ~\new_[19830]_  | ~\new_[19831]_ ;
  assign \new_[19830]_  = ~\new_[3895]_  & ~\new_[3972]_ ;
  assign \new_[19831]_  = ~\new_[19832]_ ;
  assign \new_[19832]_  = ~\new_[994]_  & (~\new_[4399]_  | ~\new_[4772]_ );
  assign \new_[19833]_  = ~\new_[19834]_  & ~\new_[19839]_ ;
  assign \new_[19834]_  = ~\new_[19835]_  | (~\new_[10947]_  & ~\new_[21267]_ );
  assign \new_[19835]_  = \new_[19836]_  & \new_[19838]_ ;
  assign \new_[19836]_  = ~\new_[12712]_  | ~\new_[18355]_ ;
  assign \new_[19837]_  = ~\new_[19838]_ ;
  assign \new_[19838]_  = ~\new_[18454]_  | ~\new_[19018]_  | ~\new_[17532]_  | ~\new_[18012]_ ;
  assign \new_[19839]_  = ~\new_[21274]_  & (~\new_[6812]_  | ~\new_[12701]_ );
  assign \new_[19840]_  = ~\new_[19841]_  | ~\new_[19846]_ ;
  assign \new_[19841]_  = ~\new_[19842]_ ;
  assign \new_[19842]_  = ~\new_[21180]_  & (~\new_[19843]_  | ~\new_[19845]_ );
  assign \new_[19843]_  = ~\new_[19844]_  & ~\new_[4049]_ ;
  assign \new_[19844]_  = ~\new_[19587]_  & ~\new_[6761]_ ;
  assign \new_[19845]_  = ~\new_[4548]_  | ~\new_[19623]_ ;
  assign \new_[19846]_  = ~\new_[19847]_  & ~\new_[19848]_ ;
  assign \new_[19847]_  = ~\new_[986]_  & (~\new_[4512]_  | ~\new_[4479]_ );
  assign \new_[19848]_  = ~\new_[19849]_  | ~\new_[19851]_ ;
  assign \new_[19849]_  = ~\new_[19850]_ ;
  assign \new_[19850]_  = ~\new_[4341]_  | ~\new_[10151]_ ;
  assign \new_[19851]_  = ~\new_[19852]_ ;
  assign \new_[19852]_  = ~\new_[9882]_  | ~\new_[5724]_  | ~\new_[6565]_ ;
  assign \new_[19853]_  = ~\new_[19861]_  | ~\new_[19854]_  | ~\new_[19855]_ ;
  assign \new_[19854]_  = ~\new_[19795]_  | (~\new_[4204]_  & ~\new_[8167]_ );
  assign \new_[19855]_  = ~\new_[19856]_  & (~\new_[4751]_  | ~\new_[18406]_ );
  assign \new_[19856]_  = ~\new_[19859]_  | ~\new_[9667]_  | ~\new_[19857]_  | ~\new_[19858]_ ;
  assign \new_[19857]_  = \new_[19229]_  | \new_[7639]_ ;
  assign \new_[19858]_  = ~\new_[12876]_  & (~\new_[11147]_  | ~\new_[17518]_ );
  assign \new_[19859]_  = ~\new_[19860]_ ;
  assign \new_[19860]_  = ~\new_[11076]_  & ~\new_[19240]_ ;
  assign \new_[19861]_  = ~\new_[932]_  | (~\new_[4733]_  & ~\new_[4579]_ );
  assign \new_[19862]_  = \new_[6526]_  & \new_[11669]_ ;
  assign \new_[19863]_  = ~\new_[8822]_  & ~\new_[9686]_ ;
  assign \new_[19864]_  = ~\new_[7363]_  | ~\new_[21084]_ ;
  assign \new_[19865]_  = ~\new_[21357]_  | (~\new_[3873]_  & ~\new_[19866]_ );
  assign \new_[19866]_  = ~\new_[938]_ ;
  assign \new_[19867]_  = ~\new_[19869]_  & (~\new_[19868]_  | ~\new_[18583]_ );
  assign \new_[19868]_  = \new_[4853]_  | \new_[5568]_ ;
  assign \new_[19869]_  = ~\new_[5981]_  | ~\new_[5384]_  | ~\new_[5216]_ ;
  assign n883 = ~\new_[19871]_  | ~\new_[19873]_ ;
  assign \new_[19871]_  = ~\new_[20972]_  | ~\new_[19872]_ ;
  assign \new_[19872]_  = ~\new_[17582]_ ;
  assign \new_[19873]_  = ~\new_[18413]_  | ~\new_[15523]_ ;
  assign \new_[19874]_  = ~\new_[17582]_ ;
  assign \new_[19875]_  = ~\new_[19881]_  | ~\new_[5051]_  | ~\new_[19876]_  | ~\new_[19879]_ ;
  assign \new_[19876]_  = \new_[6348]_  & \new_[19877]_ ;
  assign \new_[19877]_  = ~\new_[19878]_  & (~\new_[6614]_  | ~\new_[17925]_ );
  assign \new_[19878]_  = ~\new_[12292]_  | ~\new_[9126]_ ;
  assign \new_[19879]_  = \new_[5055]_  & \new_[19880]_ ;
  assign \new_[19880]_  = ~\new_[9299]_  | ~\new_[16763]_ ;
  assign \new_[19881]_  = ~\new_[6015]_  | ~\new_[18380]_ ;
  assign \new_[19882]_  = ~\new_[4432]_  | ~\new_[19885]_  | ~\new_[19883]_  | ~\new_[19884]_ ;
  assign \new_[19883]_  = ~\new_[930]_  | (~\new_[4207]_  & ~\new_[6462]_ );
  assign \new_[19884]_  = ~\new_[20507]_  | (~\new_[4492]_  & ~\new_[4588]_ );
  assign \new_[19885]_  = ~\new_[19886]_  & ~\new_[19889]_ ;
  assign \new_[19886]_  = ~\new_[11979]_  | ~\new_[19887]_  | ~\new_[9620]_  | ~\new_[8540]_ ;
  assign \new_[19887]_  = ~\new_[19888]_ ;
  assign \new_[19888]_  = ~\new_[10987]_  & ~\new_[18070]_ ;
  assign \new_[19889]_  = ~\new_[19157]_  & ~\new_[6085]_ ;
  assign \new_[19890]_  = ~\new_[19891]_  & ~\new_[19892]_ ;
  assign \new_[19891]_  = ~\new_[6645]_  | ~\new_[11223]_ ;
  assign \new_[19892]_  = ~\new_[18942]_  & ~\new_[19893]_ ;
  assign \new_[19893]_  = ~\new_[12953]_  & ~\new_[5797]_ ;
  assign \new_[19894]_  = ~\new_[18942]_  | (~\new_[4416]_  & ~\new_[10131]_ );
  assign \new_[19895]_  = ~\new_[994]_  | (~\new_[19896]_  & ~\new_[19897]_ );
  assign \new_[19896]_  = ~\new_[5198]_  | ~\new_[5491]_ ;
  assign \new_[19897]_  = ~\new_[5064]_  | ~\new_[7137]_ ;
  assign \new_[19898]_  = ~\new_[21205]_  | (~\new_[19899]_  & ~\new_[19900]_ );
  assign \new_[19899]_  = ~\new_[5796]_  | ~\new_[5171]_ ;
  assign \new_[19900]_  = ~\new_[5170]_  | ~\new_[10748]_ ;
  assign \new_[19901]_  = \new_[20413]_ ;
  assign \new_[19902]_  = ~\new_[19909]_  | ~\new_[19907]_  | ~\new_[19904]_  | ~\new_[19903]_ ;
  assign \new_[19903]_  = ~\new_[4133]_  | ~\new_[940]_ ;
  assign \new_[19904]_  = \new_[19905]_  & \new_[19906]_ ;
  assign \new_[19905]_  = ~\new_[19509]_  | (~\new_[4848]_  & ~\new_[11070]_ );
  assign \new_[19906]_  = ~\new_[19640]_  | (~\new_[4547]_  & ~\new_[13178]_ );
  assign \new_[19907]_  = ~\new_[5513]_  & ~\new_[19908]_ ;
  assign \new_[19908]_  = ~\new_[19640]_  & ~\new_[5085]_ ;
  assign \new_[19909]_  = ~\new_[21386]_  | (~\new_[4297]_  & ~\new_[13178]_ );
  assign \new_[19910]_  = ~\new_[19911]_ ;
  assign \new_[19911]_  = ~\new_[18046]_  & (~\new_[10215]_  | ~\new_[17165]_ );
  assign \new_[19912]_  = ~\new_[21073]_  & (~\new_[21681]_  | ~\new_[18046]_ );
  assign \new_[19913]_  = ~\new_[16206]_  | ~\new_[19182]_ ;
  assign \new_[19914]_  = ~\new_[19924]_  | ~\new_[19915]_  | ~\new_[19923]_ ;
  assign \new_[19915]_  = ~\new_[19916]_  | ~\new_[19918]_ ;
  assign \new_[19916]_  = ~\new_[19917]_ ;
  assign \new_[19917]_  = ~\new_[926]_ ;
  assign \new_[19918]_  = ~\new_[19921]_  | ~\new_[5185]_  | ~\new_[19919]_ ;
  assign \new_[19919]_  = ~\new_[19920]_  | ~\new_[19424]_ ;
  assign \new_[19920]_  = ~\new_[4643]_ ;
  assign \new_[19921]_  = \new_[6210]_  & \new_[19922]_ ;
  assign \new_[19922]_  = \new_[19361]_  | \new_[10284]_ ;
  assign \new_[19923]_  = ~\new_[4063]_  & ~\new_[4125]_ ;
  assign \new_[19924]_  = \new_[19925]_  & \new_[19926]_ ;
  assign \new_[19925]_  = ~\new_[5369]_ ;
  assign \new_[19926]_  = ~\new_[19927]_  & ~\new_[19929]_ ;
  assign \new_[19927]_  = ~\new_[10067]_  | ~\new_[19928]_  | ~\new_[12405]_ ;
  assign \new_[19928]_  = ~\new_[10292]_ ;
  assign \new_[19929]_  = ~\new_[19930]_  | ~\new_[14197]_ ;
  assign \new_[19930]_  = ~\new_[8149]_ ;
  assign \new_[19931]_  = ~\new_[19932]_  | ~\new_[19938]_ ;
  assign \new_[19932]_  = ~\new_[19933]_  & ~\new_[19934]_ ;
  assign \new_[19933]_  = \new_[14527]_  & \new_[19327]_ ;
  assign \new_[19934]_  = ~\new_[19935]_  | ~\new_[19937]_ ;
  assign \new_[19935]_  = ~\new_[19936]_  | ~\new_[14546]_  | ~\new_[19152]_ ;
  assign \new_[19936]_  = ~\new_[21056]_ ;
  assign \new_[19937]_  = ~\new_[15525]_  | ~\new_[21056]_ ;
  assign \new_[19938]_  = ~\new_[18569]_  | (~\new_[13308]_  & ~\new_[13427]_ );
  assign \new_[19939]_  = ~\new_[19940]_ ;
  assign \new_[19940]_  = \new_[19327]_  & \new_[14527]_ ;
  assign \new_[19941]_  = ~\new_[1134]_ ;
  assign \new_[19942]_  = ~\new_[14546]_  | ~\new_[19152]_ ;
  assign \new_[19943]_  = ~\new_[19947]_  | ~\new_[19944]_  | ~\new_[19945]_ ;
  assign \new_[19944]_  = ~\new_[3961]_  & ~\new_[3918]_ ;
  assign \new_[19945]_  = ~\new_[19946]_ ;
  assign \new_[19946]_  = ~\new_[979]_  & (~\new_[4400]_  | ~\new_[4334]_ );
  assign \new_[19947]_  = ~\new_[19948]_  & ~\new_[19953]_ ;
  assign \new_[19948]_  = ~\new_[19949]_  | (~\new_[7602]_  & ~\new_[19262]_ );
  assign \new_[19949]_  = \new_[19951]_  & \new_[19952]_ ;
  assign \new_[19950]_  = ~\new_[19951]_ ;
  assign \new_[19951]_  = ~\new_[13344]_  | ~\new_[17486]_ ;
  assign \new_[19952]_  = ~\new_[13711]_  | ~\new_[18157]_ ;
  assign \new_[19953]_  = ~\new_[20622]_  & (~\new_[7711]_  | ~\new_[12870]_ );
  assign \new_[19954]_  = \new_[19955]_ ;
  assign \new_[19955]_  = ~\new_[19960]_  | ~\new_[19959]_  | ~\new_[19956]_  | ~\new_[19958]_ ;
  assign \new_[19956]_  = ~\new_[19957]_  | ~\new_[964]_ ;
  assign \new_[19957]_  = ~\new_[6113]_  | ~\new_[4724]_  | ~\new_[5391]_  | ~\new_[5188]_ ;
  assign \new_[19958]_  = ~\new_[19807]_  | (~\new_[4488]_  & ~\new_[6001]_ );
  assign \new_[19959]_  = ~\new_[4572]_  & ~\new_[4433]_ ;
  assign \new_[19960]_  = ~\new_[17715]_  | (~\new_[4638]_  & ~\new_[5578]_ );
  assign \new_[19961]_  = ~\new_[19962]_  & ~\new_[19963]_ ;
  assign \new_[19962]_  = ~\new_[6612]_  | ~\new_[20458]_ ;
  assign \new_[19963]_  = ~\new_[18412]_  & ~\new_[7165]_ ;
  assign \new_[19964]_  = ~\new_[18522]_  | ~\new_[6738]_ ;
  assign \new_[19965]_  = \new_[9041]_  & \new_[19966]_ ;
  assign \new_[19966]_  = ~\new_[19512]_  | ~\new_[19967]_  | ~\new_[19208]_ ;
  assign \new_[19967]_  = ~\new_[15335]_  | ~\new_[11535]_  | ~\new_[11782]_  | ~\new_[12719]_ ;
  assign \new_[19968]_  = ~\new_[19179]_  | (~\new_[6302]_  & ~\new_[6668]_ );
  assign \new_[19969]_  = ~\new_[4656]_  | ~\new_[19976]_  | ~\new_[19970]_  | ~\new_[19971]_ ;
  assign \new_[19970]_  = ~\new_[21180]_  | (~\new_[3856]_  & ~\new_[5462]_ );
  assign \new_[19971]_  = ~\new_[986]_  | ~\new_[19972]_ ;
  assign \new_[19972]_  = ~\new_[5665]_  | ~\new_[5405]_  | ~\new_[19973]_  | ~\new_[19975]_ ;
  assign \new_[19973]_  = ~\new_[19974]_ ;
  assign \new_[19974]_  = ~\new_[19257]_  & (~\new_[7446]_  | ~\new_[8462]_ );
  assign \new_[19975]_  = \new_[10876]_  & \new_[6891]_ ;
  assign \new_[19976]_  = ~\new_[19977]_ ;
  assign \new_[19977]_  = ~\new_[6893]_  | ~\new_[7359]_  | ~\new_[4360]_  | ~\new_[6564]_ ;
  assign \new_[19978]_  = ~\new_[19979]_  | ~\new_[19982]_ ;
  assign \new_[19979]_  = ~\new_[19981]_  & (~\new_[19980]_  | ~\new_[21386]_ );
  assign \new_[19980]_  = ~\new_[6455]_  | ~\new_[5644]_  | ~\new_[5044]_  | ~\new_[4482]_ ;
  assign \new_[19981]_  = ~\new_[21008]_  & (~\new_[4107]_  | ~\new_[4580]_ );
  assign \new_[19982]_  = ~\new_[19983]_  & ~\new_[19986]_ ;
  assign \new_[19983]_  = ~\new_[5819]_  | ~\new_[4370]_  | ~\new_[19984]_ ;
  assign \new_[19984]_  = ~\new_[19985]_  & (~\new_[18569]_  | ~\new_[12532]_ );
  assign \new_[19985]_  = ~\new_[21013]_  | ~\new_[8504]_ ;
  assign \new_[19986]_  = ~\new_[5420]_  | ~\new_[8396]_ ;
  assign \new_[19987]_  = ~\new_[19988]_  & (~\new_[7738]_  | ~\new_[19284]_ );
  assign \new_[19988]_  = ~\new_[11787]_  | ~\new_[7240]_ ;
  assign \new_[19989]_  = ~\new_[20941]_  | (~\new_[19931]_  & ~\new_[7979]_ );
  assign \new_[19990]_  = ~\new_[19991]_  & (~\new_[10388]_  | ~\new_[16875]_ );
  assign \new_[19991]_  = \new_[16595]_  & \new_[17671]_ ;
  assign \new_[19992]_  = ~\new_[9358]_  | ~\new_[17285]_ ;
  assign \new_[19993]_  = ~\new_[19994]_  | ~\new_[19996]_ ;
  assign \new_[19994]_  = \new_[3753]_  & \new_[19995]_ ;
  assign \new_[19995]_  = ~\new_[4059]_  | ~\new_[994]_ ;
  assign \new_[19996]_  = \new_[4074]_  & \new_[19997]_ ;
  assign \new_[19997]_  = (~\new_[16153]_  | ~\new_[17144]_ ) & (~\new_[21272]_  | ~\new_[21631]_ );
  assign \new_[19998]_  = ~\new_[4103]_  | ~\new_[4421]_  | ~\new_[19999]_  | ~\new_[20001]_ ;
  assign \new_[19999]_  = ~\new_[20000]_ ;
  assign \new_[20000]_  = ~\new_[19017]_  & (~\new_[4382]_  | ~\new_[5622]_ );
  assign \new_[20001]_  = ~\new_[20002]_  & ~\new_[20003]_ ;
  assign \new_[20002]_  = ~\new_[12835]_  | ~\new_[13574]_  | ~\new_[7180]_  | ~\new_[10258]_ ;
  assign \new_[20003]_  = ~\new_[4445]_ ;
  assign \new_[20004]_  = \new_[20005]_ ;
  assign \new_[20005]_  = ~\new_[20012]_  | ~\new_[20006]_  | ~\new_[20008]_  | ~\new_[20007]_ ;
  assign \new_[20006]_  = ~\new_[5903]_  & ~\new_[4177]_ ;
  assign \new_[20007]_  = ~\new_[1004]_  | (~\new_[4166]_  & ~\new_[4969]_ );
  assign \new_[20008]_  = ~\new_[20011]_  | (~\new_[20009]_  & ~\new_[20010]_ );
  assign \new_[20009]_  = ~\new_[7364]_  | ~\new_[4775]_  | ~\new_[8323]_ ;
  assign \new_[20010]_  = ~\new_[13786]_  | ~\new_[4715]_  | ~\new_[5964]_ ;
  assign \new_[20011]_  = ~\new_[1004]_ ;
  assign \new_[20012]_  = ~\new_[20013]_  & (~\new_[6735]_  | ~\new_[18525]_ );
  assign \new_[20013]_  = \new_[5348]_  & \new_[19032]_ ;
  assign \new_[20014]_  = \new_[17940]_  | \new_[5808]_ ;
  assign \new_[20015]_  = ~\new_[21218]_  | ~\new_[19585]_ ;
  assign \new_[20016]_  = ~\new_[930]_  | (~\new_[4534]_  & ~\new_[20428]_ );
  assign \new_[20017]_  = ~\new_[20024]_  | ~\new_[20018]_  | ~\new_[20022]_ ;
  assign \new_[20018]_  = ~\new_[950]_  | (~\new_[20019]_  & ~\new_[20020]_ );
  assign \new_[20019]_  = ~\new_[4264]_  | ~\new_[5362]_ ;
  assign \new_[20020]_  = ~\new_[20021]_  | ~\new_[20463]_ ;
  assign \new_[20021]_  = ~\new_[6406]_  & ~\new_[6622]_ ;
  assign \new_[20022]_  = ~\new_[20023]_  & (~\new_[21071]_  | ~\new_[4439]_ );
  assign \new_[20023]_  = ~\new_[6732]_  | ~\new_[6530]_  | ~\new_[5165]_  | ~\new_[5091]_ ;
  assign \new_[20024]_  = ~\new_[21142]_  | (~\new_[4314]_  & ~\new_[10541]_ );
  assign \new_[20025]_  = ~\new_[20026]_  | ~\new_[20027]_  | ~\new_[20029]_  | ~\new_[4112]_ ;
  assign \new_[20026]_  = ~\new_[19470]_  | (~\new_[4614]_  & ~\new_[4938]_ );
  assign \new_[20027]_  = ~\new_[20028]_ ;
  assign \new_[20028]_  = ~\new_[935]_  & (~\new_[4627]_  | ~\new_[5081]_ );
  assign \new_[20029]_  = \new_[20030]_  & \new_[20032]_ ;
  assign \new_[20030]_  = ~\new_[20031]_ ;
  assign \new_[20031]_  = ~\new_[18292]_  & (~\new_[6809]_  | ~\new_[12959]_ );
  assign \new_[20032]_  = ~\new_[20033]_  & ~\new_[20034]_ ;
  assign \new_[20033]_  = ~\new_[10198]_  | ~\new_[12910]_  | ~\new_[13027]_ ;
  assign \new_[20034]_  = ~\new_[19702]_  & ~\new_[9679]_ ;
  assign \new_[20035]_  = ~\new_[21401]_  & ~\new_[21403]_ ;
  assign \new_[20036]_  = ~\new_[21077]_ ;
  assign \new_[20037]_  = ~\new_[20035]_ ;
  assign \new_[20038]_  = ~\new_[19786]_  | (~\new_[4038]_  & ~\new_[5963]_ );
  assign \new_[20039]_  = ~\new_[20040]_  & (~\new_[4669]_  | ~\new_[19740]_ );
  assign \new_[20040]_  = ~\new_[19229]_  & (~\new_[7039]_  | ~\new_[13319]_ );
  assign \new_[20041]_  = ~\new_[932]_  | (~\new_[4683]_  & ~\new_[4591]_ );
  assign \new_[20042]_  = ~\new_[20043]_  & (~\new_[6066]_  | ~\new_[17106]_ );
  assign \new_[20043]_  = ~\new_[12300]_  | ~\new_[20044]_  | ~\new_[7838]_ ;
  assign \new_[20044]_  = ~\new_[20045]_ ;
  assign \new_[20045]_  = ~\new_[18084]_  & (~\new_[9557]_  | ~\new_[11100]_ );
  assign \new_[20046]_  = \new_[20047]_  ^ \new_[20051]_ ;
  assign \new_[20047]_  = \new_[20048]_ ;
  assign \new_[20048]_  = ~\new_[20049]_ ;
  assign \new_[20049]_  = ~\new_[20050]_ ;
  assign \new_[20050]_  = ~\new_[4270]_  | ~\new_[4257]_  | ~\new_[3994]_  | ~\new_[3802]_ ;
  assign \new_[20051]_  = ~\new_[21101]_  | ~\new_[9391]_ ;
  assign \new_[20052]_  = ~\new_[21101]_  | ~\new_[9391]_ ;
  assign \new_[20053]_  = ~\new_[20048]_ ;
  assign \new_[20054]_  = ~\new_[20059]_  | ~\new_[4011]_  | ~\new_[20055]_  | ~\new_[20056]_ ;
  assign \new_[20055]_  = ~\new_[19540]_  | ~\new_[3916]_ ;
  assign \new_[20056]_  = ~\new_[20057]_  & ~\new_[20058]_ ;
  assign \new_[20057]_  = ~\new_[5050]_ ;
  assign \new_[20058]_  = ~\new_[964]_  & ~\new_[4137]_ ;
  assign \new_[20059]_  = ~\new_[20060]_  & (~\new_[5049]_  | ~\new_[18380]_ );
  assign \new_[20060]_  = ~\new_[11328]_  | ~\new_[10648]_  | ~\new_[10732]_ ;
  assign \new_[20061]_  = ~\new_[20064]_  | ~\new_[20063]_  | ~\new_[20062]_  | ~\new_[4225]_ ;
  assign \new_[20062]_  = ~\new_[19917]_  | (~\new_[4205]_  & ~\new_[7305]_ );
  assign \new_[20063]_  = ~\new_[926]_  | (~\new_[4506]_  & ~\new_[4770]_ );
  assign \new_[20064]_  = ~\new_[20065]_  & ~\new_[20067]_ ;
  assign \new_[20065]_  = ~\new_[13561]_  | ~\new_[8992]_  | ~\new_[20066]_  | ~\new_[9678]_ ;
  assign \new_[20066]_  = \new_[10918]_  | \new_[19145]_ ;
  assign \new_[20067]_  = ~\new_[20152]_  & ~\new_[7674]_ ;
  assign \new_[20068]_  = ~\new_[20074]_  | ~\new_[20073]_  | ~\new_[20069]_  | ~\new_[20072]_ ;
  assign \new_[20069]_  = ~\new_[986]_  | (~\new_[20070]_  & ~\new_[20071]_ );
  assign \new_[20070]_  = ~\new_[4413]_ ;
  assign \new_[20071]_  = ~\new_[8812]_  | ~\new_[4269]_  | ~\new_[5024]_ ;
  assign \new_[20072]_  = ~\new_[21180]_  | (~\new_[3963]_  & ~\new_[7291]_ );
  assign \new_[20073]_  = ~\new_[7286]_  & ~\new_[4354]_ ;
  assign \new_[20074]_  = ~\new_[20075]_  | ~\new_[984]_ ;
  assign \new_[20075]_  = \new_[5533]_  | \new_[5592]_ ;
  assign \new_[20076]_  = \new_[20068]_ ;
  assign \new_[20077]_  = ~\new_[20081]_  | ~\new_[20078]_  | ~\new_[20079]_ ;
  assign \new_[20078]_  = ~\new_[4002]_  & ~\new_[3897]_ ;
  assign \new_[20079]_  = ~\new_[20080]_ ;
  assign \new_[20080]_  = ~\new_[986]_  & (~\new_[4624]_  | ~\new_[4335]_ );
  assign \new_[20081]_  = ~\new_[20082]_  & ~\new_[20086]_ ;
  assign \new_[20082]_  = ~\new_[20083]_  | (~\new_[19257]_  & ~\new_[8572]_ );
  assign \new_[20083]_  = \new_[20084]_  & \new_[20085]_ ;
  assign \new_[20084]_  = ~\new_[16119]_  | ~\new_[18826]_ ;
  assign \new_[20085]_  = ~\new_[18322]_  | ~\new_[12492]_ ;
  assign \new_[20086]_  = ~\new_[16889]_  & (~\new_[6816]_  | ~\new_[14202]_ );
  assign \new_[20087]_  = ~\new_[20084]_ ;
  assign \new_[20088]_  = ~\new_[20096]_  | ~\new_[20089]_  | ~\new_[20090]_ ;
  assign \new_[20089]_  = ~\new_[19157]_  | (~\new_[5412]_  & ~\new_[9690]_ );
  assign \new_[20090]_  = ~\new_[20091]_  & ~\new_[20094]_ ;
  assign \new_[20091]_  = ~\new_[16151]_  | ~\new_[9794]_  | ~\new_[20092]_ ;
  assign \new_[20092]_  = ~\new_[20093]_ ;
  assign \new_[20093]_  = ~\new_[1080]_  & (~\new_[16663]_  | ~\new_[13872]_ );
  assign \new_[20094]_  = ~\new_[19600]_  & ~\new_[20095]_ ;
  assign \new_[20095]_  = ~\new_[13274]_  & ~\new_[9189]_ ;
  assign \new_[20096]_  = ~\new_[20097]_  | ~\new_[20098]_ ;
  assign \new_[20097]_  = ~\new_[7145]_  | ~\new_[13905]_ ;
  assign \new_[20098]_  = ~\new_[20099]_ ;
  assign \new_[20099]_  = ~\new_[1080]_ ;
  assign \new_[20100]_  = ~\new_[1080]_ ;
  assign \new_[20101]_  = ~\new_[20110]_  | ~\new_[20109]_  | ~\new_[20106]_  | ~\new_[20102]_ ;
  assign \new_[20102]_  = ~\new_[930]_  | (~\new_[20103]_  & ~\new_[20105]_ );
  assign \new_[20103]_  = ~\new_[20104]_  | ~\new_[4712]_  | ~\new_[5087]_ ;
  assign \new_[20104]_  = \new_[7270]_  & \new_[11675]_ ;
  assign \new_[20105]_  = ~\new_[6656]_  | ~\new_[19887]_ ;
  assign \new_[20106]_  = ~\new_[20107]_  & ~\new_[20108]_ ;
  assign \new_[20107]_  = ~\new_[5316]_  | ~\new_[8470]_ ;
  assign \new_[20108]_  = ~\new_[4631]_ ;
  assign \new_[20109]_  = ~\new_[19585]_  | (~\new_[4593]_  & ~\new_[4950]_ );
  assign \new_[20110]_  = ~\new_[20111]_  & (~\new_[5609]_  | ~\new_[19157]_ );
  assign \new_[20111]_  = \new_[6737]_  & \new_[17585]_ ;
  assign \new_[20112]_  = ~\new_[7524]_  | ~\new_[3917]_  | ~\new_[3849]_  | ~\new_[4060]_ ;
  assign \new_[20113]_  = ~\new_[20112]_ ;
  assign \new_[20114]_  = ~\new_[20117]_  | ~\new_[4117]_  | ~\new_[20115]_  | ~\new_[20116]_ ;
  assign \new_[20115]_  = ~\new_[3903]_ ;
  assign \new_[20116]_  = ~\new_[3996]_  | ~\new_[956]_ ;
  assign \new_[20117]_  = ~\new_[20118]_  & ~\new_[4701]_ ;
  assign \new_[20118]_  = ~\new_[9304]_  | ~\new_[9001]_  | ~\new_[9294]_ ;
  assign \new_[20119]_  = ~\new_[20112]_ ;
  assign \new_[20120]_  = \new_[20121]_ ;
  assign \new_[20121]_  = ~\new_[20125]_  | ~\new_[20124]_  | ~\new_[20122]_  | ~\new_[20123]_ ;
  assign \new_[20122]_  = ~\new_[3936]_  | ~\new_[956]_ ;
  assign \new_[20123]_  = ~\new_[21453]_  | (~\new_[4276]_  & ~\new_[6538]_ );
  assign \new_[20124]_  = ~\new_[19530]_  | (~\new_[4868]_  & ~\new_[4843]_ );
  assign \new_[20125]_  = \new_[20126]_  & \new_[20127]_ ;
  assign \new_[20126]_  = ~\new_[19748]_  | (~\new_[6382]_  & ~\new_[15178]_ );
  assign \new_[20127]_  = ~\new_[20128]_  & (~\new_[8343]_  | ~\new_[17689]_ );
  assign \new_[20128]_  = ~\new_[20129]_  & ~\new_[20130]_ ;
  assign \new_[20129]_  = ~\new_[18021]_ ;
  assign \new_[20130]_  = ~\new_[13287]_  & ~\new_[8344]_ ;
  assign \new_[20131]_  = ~\new_[20136]_  | ~\new_[20132]_  | ~\new_[20134]_ ;
  assign \new_[20132]_  = ~\new_[20133]_ ;
  assign \new_[20133]_  = ~\new_[21205]_  & (~\new_[4436]_  | ~\new_[4590]_ );
  assign \new_[20134]_  = ~\new_[21205]_  | ~\new_[20135]_ ;
  assign \new_[20135]_  = ~\new_[5454]_  | ~\new_[5656]_  | ~\new_[4743]_  | ~\new_[5937]_ ;
  assign \new_[20136]_  = ~\new_[20137]_  & ~\new_[4147]_ ;
  assign \new_[20137]_  = ~\new_[10947]_  | ~\new_[8911]_  | ~\new_[20138]_  | ~\new_[20139]_ ;
  assign \new_[20138]_  = ~\new_[7026]_ ;
  assign \new_[20139]_  = ~\new_[7520]_  & (~\new_[21638]_  | ~\new_[12547]_ );
  assign \new_[20140]_  = ~\new_[21453]_  | (~\new_[20370]_  & ~\new_[20142]_ );
  assign \new_[20141]_  = ~\new_[8676]_ ;
  assign \new_[20142]_  = ~\new_[20143]_  | ~\new_[20144]_ ;
  assign \new_[20143]_  = ~\new_[9642]_  | ~\new_[17749]_ ;
  assign \new_[20144]_  = ~\new_[6943]_  | ~\new_[19337]_ ;
  assign \new_[20145]_  = ~\new_[20146]_  | ~\new_[20147]_ ;
  assign \new_[20146]_  = ~\new_[19736]_  | ~\new_[4055]_ ;
  assign \new_[20147]_  = ~\new_[20148]_  | ~\new_[1025]_ ;
  assign \new_[20148]_  = ~\new_[10150]_  | ~\new_[20149]_  | ~\new_[5456]_  | ~\new_[8873]_ ;
  assign \new_[20149]_  = ~\new_[20150]_  & ~\new_[20151]_ ;
  assign \new_[20150]_  = ~\new_[16416]_  & ~\new_[19178]_ ;
  assign \new_[20151]_  = ~\new_[11067]_ ;
  assign \new_[20152]_  = ~\new_[1025]_ ;
  assign \new_[20153]_  = ~\new_[7487]_  | ~\new_[18769]_ ;
  assign \new_[20154]_  = ~\new_[12869]_  | ~\new_[19094]_ ;
  assign \new_[20155]_  = ~\new_[20156]_  & ~\new_[20159]_ ;
  assign \new_[20156]_  = ~\new_[20157]_  | ~\new_[20158]_ ;
  assign \new_[20157]_  = \new_[18017]_  | \new_[13849]_ ;
  assign \new_[20158]_  = \new_[18974]_  | \new_[17251]_ ;
  assign \new_[20159]_  = ~\new_[20160]_ ;
  assign \new_[20160]_  = ~\new_[14343]_  | ~\new_[17457]_ ;
  assign \new_[20161]_  = ~\new_[20162]_ ;
  assign \new_[20162]_  = ~\new_[20157]_ ;
  assign \new_[20163]_  = ~\new_[20158]_ ;
  assign \new_[20164]_  = \new_[20165]_  & \new_[20169]_ ;
  assign \new_[20165]_  = ~\new_[20166]_  & ~\new_[20168]_ ;
  assign \new_[20166]_  = \new_[20167]_ ;
  assign \new_[20167]_  = ~\new_[1030]_ ;
  assign \new_[20168]_  = \new_[1078]_ ;
  assign \new_[20169]_  = \new_[943]_ ;
  assign \new_[20170]_  = ~\new_[943]_ ;
  assign \new_[20171]_  = ~\new_[20167]_ ;
  assign \new_[20172]_  = ~\new_[20168]_ ;
  assign \new_[20173]_  = ~\new_[20174]_ ;
  assign \new_[20174]_  = ~\new_[20180]_  | ~\new_[20178]_  | ~\new_[20175]_  | ~\new_[20177]_ ;
  assign \new_[20175]_  = ~\new_[20176]_  | ~\new_[19470]_ ;
  assign \new_[20176]_  = ~\new_[4285]_  | ~\new_[6013]_ ;
  assign \new_[20177]_  = ~\new_[4349]_  | ~\new_[18386]_ ;
  assign \new_[20178]_  = ~\new_[20179]_  & ~\new_[4087]_ ;
  assign \new_[20179]_  = ~\new_[7485]_  | ~\new_[13535]_ ;
  assign \new_[20180]_  = ~\new_[4057]_  | ~\new_[19564]_ ;
  assign \new_[20181]_  = ~\new_[956]_ ;
  assign \new_[20182]_  = ~\new_[10826]_  | ~\new_[8279]_  | ~\new_[5439]_  | ~\new_[5130]_ ;
  assign \new_[20183]_  = ~\new_[7440]_  | ~\new_[5498]_ ;
  assign \new_[20184]_  = ~\new_[4657]_  | ~\new_[5461]_ ;
  assign \new_[20185]_  = ~\new_[20186]_  | ~\new_[20189]_ ;
  assign \new_[20186]_  = ~\new_[20188]_  & (~\new_[20187]_  | ~\new_[20464]_ );
  assign \new_[20187]_  = ~\new_[6460]_  | ~\new_[5652]_  | ~\new_[4487]_  | ~\new_[4706]_ ;
  assign \new_[20188]_  = ~\new_[21071]_  & (~\new_[4110]_  | ~\new_[4587]_ );
  assign \new_[20189]_  = ~\new_[20190]_  & ~\new_[20193]_ ;
  assign \new_[20190]_  = ~\new_[5822]_  | ~\new_[5868]_  | ~\new_[20191]_ ;
  assign \new_[20191]_  = ~\new_[20192]_  & (~\new_[12442]_  | ~\new_[17381]_ );
  assign \new_[20192]_  = ~\new_[7827]_  | ~\new_[9573]_ ;
  assign \new_[20193]_  = ~\new_[4182]_  | ~\new_[7499]_ ;
  assign \new_[20194]_  = ~\new_[20199]_  | ~\new_[20195]_  | ~\new_[20196]_ ;
  assign \new_[20195]_  = ~\new_[19316]_  | ~\new_[3785]_ ;
  assign \new_[20196]_  = ~\new_[20197]_  & ~\new_[20198]_ ;
  assign \new_[20197]_  = ~\new_[6573]_  | ~\new_[10780]_  | ~\new_[11489]_ ;
  assign \new_[20198]_  = ~\new_[4027]_  | ~\new_[4198]_ ;
  assign \new_[20199]_  = ~\new_[21071]_  | (~\new_[20200]_  & ~\new_[20201]_ );
  assign \new_[20200]_  = ~\new_[10431]_  | ~\new_[4667]_  | ~\new_[6727]_ ;
  assign \new_[20201]_  = ~\new_[20202]_  | ~\new_[4968]_ ;
  assign \new_[20202]_  = ~\new_[18606]_  | (~\new_[7588]_  & ~\new_[11719]_ );
  assign \new_[20203]_  = ~\new_[20208]_  | ~\new_[20204]_  | ~\new_[20205]_ ;
  assign \new_[20204]_  = ~\new_[19017]_  | (~\new_[4202]_  & ~\new_[8138]_ );
  assign \new_[20205]_  = ~\new_[4559]_  & ~\new_[20206]_ ;
  assign \new_[20206]_  = \new_[20207]_  | \new_[4185]_ ;
  assign \new_[20207]_  = \new_[10028]_  | \new_[8281]_ ;
  assign \new_[20208]_  = ~\new_[937]_  | (~\new_[20209]_  & ~\new_[20210]_ );
  assign \new_[20209]_  = ~\new_[12156]_  | ~\new_[8994]_  | ~\new_[4964]_  | ~\new_[8896]_ ;
  assign \new_[20210]_  = ~\new_[6286]_  | (~\new_[5479]_  & ~\new_[19259]_ );
  assign \new_[20211]_  = ~\new_[20212]_  | ~\new_[20220]_ ;
  assign \new_[20212]_  = ~\new_[20216]_  & (~\new_[20213]_  | ~\new_[21559]_ );
  assign \new_[20213]_  = ~\new_[20214]_  | ~\new_[20215]_ ;
  assign \new_[20214]_  = ~\new_[15924]_  & ~\new_[16061]_ ;
  assign \new_[20215]_  = \new_[21396]_  | \new_[17338]_ ;
  assign \new_[20216]_  = ~\new_[20217]_  | ~\new_[20218]_ ;
  assign \new_[20217]_  = ~\new_[16095]_  | ~\new_[19403]_ ;
  assign \new_[20218]_  = ~\new_[20219]_  | ~\new_[19421]_ ;
  assign \new_[20219]_  = ~\new_[16766]_ ;
  assign \new_[20220]_  = ~\new_[15391]_  | ~\new_[21562]_ ;
  assign \new_[20221]_  = ~\new_[16095]_  | ~\new_[19403]_ ;
  assign \new_[20222]_  = ~\new_[20218]_ ;
  assign \new_[20223]_  = ~\new_[20228]_  | ~\new_[20226]_  | ~\new_[20224]_  | ~\new_[20225]_ ;
  assign \new_[20224]_  = \new_[4254]_  & \new_[4248]_ ;
  assign \new_[20225]_  = ~\new_[958]_  | (~\new_[4381]_  & ~\new_[4939]_ );
  assign \new_[20226]_  = ~\new_[20227]_  | ~\new_[17070]_ ;
  assign \new_[20227]_  = ~\new_[5092]_  | ~\new_[12822]_ ;
  assign \new_[20228]_  = ~\new_[20229]_ ;
  assign \new_[20229]_  = ~\new_[7177]_  | ~\new_[20230]_ ;
  assign \new_[20230]_  = ~\new_[20231]_ ;
  assign \new_[20231]_  = ~\new_[8893]_  | ~\new_[13116]_  | ~\new_[9868]_ ;
  assign \new_[20232]_  = ~\new_[20233]_  | ~\new_[20239]_ ;
  assign \new_[20233]_  = ~\new_[20234]_ ;
  assign \new_[20234]_  = ~\new_[20235]_  | ~\new_[18603]_ ;
  assign \new_[20235]_  = ~\new_[20236]_ ;
  assign \new_[20236]_  = ~\new_[21545]_  | ~\new_[19475]_ ;
  assign \new_[20237]_  = ~\new_[20238]_ ;
  assign \new_[20238]_  = ~\new_[20871]_ ;
  assign \new_[20239]_  = ~\new_[20240]_ ;
  assign \new_[20240]_  = \new_[995]_ ;
  assign \new_[20241]_  = ~\new_[995]_ ;
  assign \new_[20242]_  = ~\new_[20235]_ ;
  assign \new_[20243]_  = ~\new_[3997]_  | ~\new_[949]_ ;
  assign \new_[20244]_  = \new_[4253]_  & \new_[20245]_ ;
  assign \new_[20245]_  = ~\new_[20246]_  & (~\new_[6449]_  | ~\new_[18786]_ );
  assign \new_[20246]_  = ~\new_[10590]_  | ~\new_[10836]_ ;
  assign \new_[20247]_  = ~\new_[20248]_  & ~\new_[20249]_ ;
  assign \new_[20248]_  = ~\new_[5451]_  | ~\new_[8847]_ ;
  assign \new_[20249]_  = ~\new_[949]_  & ~\new_[4272]_ ;
  assign \new_[20250]_  = ~\new_[20257]_  | ~\new_[20256]_  | ~\new_[20251]_  | ~\new_[20252]_ ;
  assign \new_[20251]_  = ~\new_[3893]_  | ~\new_[958]_ ;
  assign \new_[20252]_  = ~\new_[4146]_  & ~\new_[20253]_ ;
  assign \new_[20253]_  = ~\new_[20254]_  | ~\new_[20255]_ ;
  assign \new_[20254]_  = ~\new_[6289]_ ;
  assign \new_[20255]_  = ~\new_[7463]_  & (~\new_[13749]_  | ~\new_[16670]_ );
  assign \new_[20256]_  = ~\new_[20743]_  | ~\new_[3850]_ ;
  assign \new_[20257]_  = (~\new_[12328]_  | ~\new_[19208]_ ) & (~\new_[19208]_  | ~\new_[12709]_ );
  assign \new_[20258]_  = \new_[20259]_ ;
  assign \new_[20259]_  = ~\new_[20260]_  | ~\new_[20268]_  | ~\new_[20269]_  | ~\new_[20263]_ ;
  assign \new_[20260]_  = ~\new_[20261]_  & (~\new_[5001]_  | ~\new_[19262]_ );
  assign \new_[20261]_  = ~\new_[20262]_ ;
  assign \new_[20262]_  = ~\new_[6373]_  & (~\new_[6924]_  | ~\new_[17629]_ );
  assign \new_[20263]_  = ~\new_[979]_  | ~\new_[20264]_ ;
  assign \new_[20264]_  = ~\new_[5666]_  | ~\new_[5030]_  | ~\new_[20265]_  | ~\new_[20267]_ ;
  assign \new_[20265]_  = ~\new_[20266]_ ;
  assign \new_[20266]_  = ~\new_[19787]_  & (~\new_[6636]_  | ~\new_[5494]_ );
  assign \new_[20267]_  = \new_[7872]_  & \new_[12465]_ ;
  assign \new_[20268]_  = ~\new_[4581]_ ;
  assign \new_[20269]_  = ~\new_[19816]_  | (~\new_[4036]_  & ~\new_[5463]_ );
  assign \new_[20270]_  = ~\new_[20271]_  | ~\new_[20274]_ ;
  assign \new_[20271]_  = ~\new_[20272]_  | ~\new_[20273]_ ;
  assign \new_[20272]_  = ~\new_[20011]_ ;
  assign \new_[20273]_  = ~\new_[3786]_  | ~\new_[5876]_ ;
  assign \new_[20274]_  = ~\new_[20275]_  & ~\new_[20277]_ ;
  assign \new_[20275]_  = ~\new_[20276]_  | ~\new_[6559]_  | ~\new_[4543]_  | ~\new_[5702]_ ;
  assign \new_[20276]_  = \new_[9810]_  & \new_[12334]_ ;
  assign \new_[20277]_  = ~\new_[1004]_  & (~\new_[20278]_  | ~\new_[20279]_ );
  assign \new_[20278]_  = ~\new_[4611]_  | ~\new_[19442]_ ;
  assign \new_[20279]_  = ~\new_[20280]_  & ~\new_[20281]_ ;
  assign \new_[20280]_  = ~\new_[10330]_  | ~\new_[11967]_  | ~\new_[6972]_ ;
  assign \new_[20281]_  = ~\new_[5251]_ ;
  assign \new_[20282]_  = ~\new_[20284]_  | (~\new_[3939]_  & ~\new_[20283]_ );
  assign \new_[20283]_  = ~\new_[949]_ ;
  assign \new_[20284]_  = ~\new_[20283]_  | ~\new_[5337]_  | ~\new_[20285]_  | ~\new_[5197]_ ;
  assign \new_[20285]_  = ~\new_[20286]_  & ~\new_[20287]_ ;
  assign \new_[20286]_  = ~\new_[9158]_  | ~\new_[6830]_ ;
  assign \new_[20287]_  = \new_[9435]_  | \new_[8303]_ ;
  assign \new_[20288]_  = ~\new_[20290]_  & (~\new_[20289]_  | ~\new_[921]_ );
  assign \new_[20289]_  = \new_[4858]_  | \new_[5596]_ ;
  assign \new_[20290]_  = ~\new_[6533]_  | ~\new_[4931]_  | ~\new_[5387]_ ;
  assign \new_[20291]_  = ~\new_[20292]_ ;
  assign \new_[20292]_  = ~\new_[20293]_  | ~\new_[21402]_ ;
  assign \new_[20293]_  = ~\new_[21583]_  & ~\new_[20294]_ ;
  assign \new_[20294]_  = ~\new_[19473]_  | ~\new_[19506]_ ;
  assign \new_[20295]_  = ~\new_[938]_ ;
  assign \new_[20296]_  = ~\new_[20297]_  | ~\new_[21365]_ ;
  assign \new_[20297]_  = ~\new_[9333]_  | ~\new_[18175]_ ;
  assign \new_[20298]_  = ~\new_[20299]_  | ~\new_[20301]_ ;
  assign \new_[20299]_  = ~\new_[1079]_  & ~\new_[19522]_ ;
  assign \new_[20300]_  = ~\new_[976]_ ;
  assign \new_[20301]_  = ~\new_[20589]_ ;
  assign \new_[20302]_  = ~\new_[1079]_ ;
  assign \new_[20303]_  = ~\new_[20308]_  | ~\new_[20304]_  | ~\new_[9348]_ ;
  assign \new_[20304]_  = ~\new_[21405]_  & ~\new_[20305]_ ;
  assign \new_[20305]_  = ~\new_[11066]_  | ~\new_[20306]_ ;
  assign \new_[20306]_  = ~\new_[20307]_ ;
  assign \new_[20307]_  = ~\new_[18678]_  & ~\new_[14122]_ ;
  assign \new_[20308]_  = ~\new_[11283]_  | ~\new_[18077]_ ;
  assign \new_[20309]_  = ~\new_[20317]_  & (~\new_[20311]_  | ~\new_[18483]_ );
  assign \new_[20310]_  = ~\new_[956]_ ;
  assign \new_[20311]_  = ~\new_[20314]_  | ~\new_[20312]_  | ~\new_[20313]_ ;
  assign \new_[20312]_  = ~\new_[4694]_  & (~\new_[4419]_  | ~\new_[19748]_ );
  assign \new_[20313]_  = ~\new_[21109]_ ;
  assign \new_[20314]_  = \new_[20315]_  & \new_[20316]_ ;
  assign \new_[20315]_  = ~\new_[8705]_ ;
  assign \new_[20316]_  = ~\new_[7920]_ ;
  assign \new_[20317]_  = ~\new_[4090]_  | ~\new_[3801]_  | ~\new_[20318]_ ;
  assign \new_[20318]_  = ~\new_[20319]_  & ~\new_[20320]_ ;
  assign \new_[20319]_  = ~\new_[8554]_ ;
  assign \new_[20320]_  = ~\new_[5424]_ ;
  assign \new_[20321]_  = \new_[20326]_  ^ \new_[20322]_ ;
  assign \new_[20322]_  = ~\new_[20323]_ ;
  assign \new_[20323]_  = \new_[20324]_ ;
  assign \new_[20324]_  = ~\new_[20325]_ ;
  assign \new_[20325]_  = ~\new_[4271]_  | ~\new_[4259]_  | ~\new_[3842]_  | ~\new_[4079]_ ;
  assign \new_[20326]_  = ~\new_[3490]_  | ~\new_[8227]_ ;
  assign \new_[20327]_  = ~\new_[3490]_  | ~\new_[8227]_ ;
  assign \new_[20328]_  = \new_[20327]_ ;
  assign \new_[20329]_  = ~\new_[20324]_ ;
  assign \new_[20330]_  = ~\new_[4983]_  | ~\new_[12743]_ ;
  assign \new_[20331]_  = \new_[2346]_  ^ \new_[21625]_ ;
  assign \new_[20332]_  = ~\new_[20340]_  | ~\new_[20339]_  | ~\new_[20333]_  | ~\new_[20334]_ ;
  assign \new_[20333]_  = ~\new_[19770]_  | (~\new_[6271]_  & ~\new_[7603]_ );
  assign \new_[20334]_  = ~\new_[20335]_  | ~\new_[20337]_ ;
  assign \new_[20335]_  = ~\new_[7095]_  | ~\new_[20336]_ ;
  assign \new_[20336]_  = \new_[14430]_  & \new_[17796]_ ;
  assign \new_[20337]_  = ~\new_[20338]_  | ~\new_[18542]_ ;
  assign \new_[20338]_  = \new_[16552]_  & \new_[13769]_ ;
  assign \new_[20339]_  = ~\new_[19441]_  | (~\new_[10416]_  & ~\new_[13198]_ );
  assign \new_[20340]_  = \new_[9791]_  & \new_[15016]_ ;
  assign \new_[20341]_  = ~\new_[1006]_ ;
  assign \new_[20342]_  = ~\new_[20343]_  | ~\new_[20349]_ ;
  assign \new_[20343]_  = ~\new_[20344]_  & (~\new_[20783]_  | ~\new_[3823]_ );
  assign \new_[20344]_  = ~\new_[20345]_  | ~\new_[20346]_ ;
  assign \new_[20345]_  = ~\new_[4440]_  | ~\new_[930]_ ;
  assign \new_[20346]_  = \new_[20347]_  & \new_[20348]_ ;
  assign \new_[20347]_  = \new_[13722]_  | \new_[13434]_ ;
  assign \new_[20348]_  = ~\new_[11239]_  | ~\new_[19299]_ ;
  assign \new_[20349]_  = \new_[20350]_  & \new_[20351]_ ;
  assign \new_[20350]_  = ~\new_[19157]_  | (~\new_[4758]_  & ~\new_[12728]_ );
  assign \new_[20351]_  = ~\new_[19120]_  | (~\new_[5611]_  & ~\new_[7348]_ );
  assign \new_[20352]_  = ~\new_[20353]_  | ~\new_[20358]_ ;
  assign \new_[20353]_  = ~\new_[20354]_  & ~\new_[20357]_ ;
  assign \new_[20354]_  = ~\new_[20355]_  | (~\new_[4406]_  & ~\new_[19751]_ );
  assign \new_[20355]_  = \new_[4730]_  & \new_[20356]_ ;
  assign \new_[20356]_  = \new_[19145]_  | \new_[19128]_  | \new_[17608]_  | \new_[18186]_ ;
  assign \new_[20357]_  = ~\new_[4051]_  & ~\new_[19917]_ ;
  assign \new_[20358]_  = ~\new_[20360]_  & (~\new_[20359]_  | ~\new_[21066]_ );
  assign \new_[20359]_  = ~\new_[7985]_  | ~\new_[4994]_  | ~\new_[5098]_ ;
  assign \new_[20360]_  = ~\new_[13318]_ ;
  assign \new_[20361]_  = ~\new_[20369]_  | ~\new_[20362]_  | ~\new_[20365]_ ;
  assign \new_[20362]_  = ~\new_[20364]_  & (~\new_[20363]_  | ~\new_[17518]_ );
  assign \new_[20363]_  = ~\new_[11930]_  | ~\new_[12064]_ ;
  assign \new_[20364]_  = ~\new_[19653]_  & (~\new_[8746]_  | ~\new_[11947]_ );
  assign \new_[20365]_  = ~\new_[20366]_  & ~\new_[8176]_ ;
  assign \new_[20366]_  = ~\new_[20367]_  | ~\new_[20368]_ ;
  assign \new_[20367]_  = ~\new_[10584]_  | ~\new_[18481]_ ;
  assign \new_[20368]_  = \new_[15376]_  & \new_[14631]_ ;
  assign \new_[20369]_  = ~\new_[19740]_  | (~\new_[6144]_  & ~\new_[9150]_ );
  assign \new_[20370]_  = ~\new_[20377]_  | ~\new_[20371]_  | ~\new_[20375]_ ;
  assign \new_[20371]_  = \new_[20141]_  & \new_[20372]_ ;
  assign \new_[20372]_  = ~\new_[20373]_  & ~\new_[20374]_ ;
  assign \new_[20373]_  = ~\new_[19337]_  & ~\new_[11635]_ ;
  assign \new_[20374]_  = ~\new_[17993]_  & ~\new_[12757]_ ;
  assign \new_[20375]_  = \new_[7372]_  & \new_[20376]_ ;
  assign \new_[20376]_  = ~\new_[17960]_  | ~\new_[11110]_ ;
  assign \new_[20377]_  = ~\new_[7703]_  | ~\new_[19103]_ ;
  assign \new_[20378]_  = ~\new_[20374]_ ;
  assign \new_[20379]_  = ~\new_[4928]_  | ~\new_[6825]_ ;
  assign \new_[20380]_  = ~\new_[6543]_  | ~\new_[4676]_  | ~\new_[5194]_ ;
  assign \new_[20381]_  = ~\new_[20386]_  | ~\new_[20385]_  | ~\new_[20382]_  | ~\new_[20384]_ ;
  assign \new_[20382]_  = ~\new_[20383]_ ;
  assign \new_[20383]_  = ~\new_[21563]_  & ~\new_[14359]_ ;
  assign \new_[20384]_  = ~\new_[13221]_  | ~\new_[21561]_ ;
  assign \new_[20385]_  = ~\new_[21557]_  | (~\new_[8909]_  & ~\new_[15194]_ );
  assign \new_[20386]_  = ~\new_[20387]_  & ~\new_[20389]_ ;
  assign \new_[20387]_  = ~\new_[20388]_ ;
  assign \new_[20388]_  = ~\new_[18107]_  | ~\new_[19199]_ ;
  assign \new_[20389]_  = ~\new_[15858]_  & ~\new_[21394]_ ;
  assign \new_[20390]_  = ~\new_[20389]_ ;
  assign \new_[20391]_  = ~\new_[20392]_  | ~\new_[20395]_ ;
  assign \new_[20392]_  = ~\new_[20393]_  | ~\new_[20394]_ ;
  assign \new_[20393]_  = ~\new_[19816]_ ;
  assign \new_[20394]_  = ~\new_[3872]_  | ~\new_[6301]_ ;
  assign \new_[20395]_  = ~\new_[20396]_  & ~\new_[20401]_ ;
  assign \new_[20396]_  = ~\new_[979]_  & (~\new_[20397]_  | ~\new_[20398]_ );
  assign \new_[20397]_  = ~\new_[19517]_  | ~\new_[4612]_ ;
  assign \new_[20398]_  = ~\new_[20399]_  & ~\new_[20400]_ ;
  assign \new_[20399]_  = ~\new_[10224]_  | ~\new_[10673]_  | ~\new_[6973]_ ;
  assign \new_[20400]_  = ~\new_[5256]_ ;
  assign \new_[20401]_  = ~\new_[20402]_  | ~\new_[6567]_  | ~\new_[4348]_  | ~\new_[5317]_ ;
  assign \new_[20402]_  = \new_[9963]_  & \new_[12385]_ ;
  assign \new_[20403]_  = ~\new_[20404]_  | ~\new_[20407]_ ;
  assign \new_[20404]_  = ~\new_[20405]_  & ~\new_[20406]_ ;
  assign \new_[20405]_  = ~\new_[3828]_ ;
  assign \new_[20406]_  = ~\new_[20452]_  & ~\new_[3783]_ ;
  assign \new_[20407]_  = ~\new_[20408]_  & (~\new_[4343]_  | ~\new_[18293]_ );
  assign \new_[20408]_  = ~\new_[20410]_  | (~\new_[20409]_  & ~\new_[18293]_ );
  assign \new_[20409]_  = \new_[5338]_  & \new_[10732]_ ;
  assign \new_[20410]_  = \new_[9976]_  ? \new_[18280]_  : \new_[12612]_ ;
  assign \new_[20411]_  = ~\new_[20412]_  | ~\new_[20416]_ ;
  assign \new_[20412]_  = \new_[20413]_  | \new_[20414]_ ;
  assign \new_[20413]_  = ~\new_[19898]_  | ~\new_[19895]_  | ~\new_[19890]_  | ~\new_[19894]_ ;
  assign \new_[20414]_  = ~\new_[20415]_ ;
  assign \new_[20415]_  = ~\new_[6602]_  | ~\new_[3965]_  | ~\new_[3752]_  | ~\new_[3979]_ ;
  assign \new_[20416]_  = ~\new_[20414]_  | ~\new_[20413]_ ;
  assign \new_[20417]_  = ~\new_[6602]_  | ~\new_[3965]_  | ~\new_[3979]_  | ~\new_[3752]_ ;
  assign \new_[20418]_  = ~\new_[20424]_  | ~\new_[20419]_  | ~\new_[20423]_ ;
  assign \new_[20419]_  = ~\new_[21425]_  | (~\new_[20420]_  & ~\new_[20421]_ );
  assign \new_[20420]_  = ~\new_[4807]_  | ~\new_[5233]_ ;
  assign \new_[20421]_  = ~\new_[6412]_  | ~\new_[20422]_ ;
  assign \new_[20422]_  = ~\new_[17869]_  | ~\new_[16718]_ ;
  assign \new_[20423]_  = ~\new_[18844]_  | (~\new_[4857]_  & ~\new_[12236]_ );
  assign \new_[20424]_  = ~\new_[20426]_  | (~\new_[4567]_  & ~\new_[20425]_ );
  assign \new_[20425]_  = ~\new_[20422]_  | ~\new_[19054]_ ;
  assign \new_[20426]_  = ~\new_[6801]_  | ~\new_[20427]_ ;
  assign \new_[20427]_  = ~\new_[19054]_ ;
  assign \new_[20428]_  = ~\new_[20513]_  & ~\new_[20429]_ ;
  assign \new_[20429]_  = ~\new_[16544]_  & ~\new_[20430]_ ;
  assign \new_[20430]_  = ~\new_[20433]_  | ~\new_[20431]_  | ~\new_[20432]_ ;
  assign \new_[20431]_  = ~\new_[9432]_ ;
  assign \new_[20432]_  = ~\new_[13088]_  | ~\new_[18979]_ ;
  assign \new_[20433]_  = ~\new_[20434]_ ;
  assign \new_[20434]_  = ~\new_[19196]_  & ~\new_[15677]_ ;
  assign \new_[20435]_  = ~\new_[20432]_ ;
  assign \new_[20436]_  = ~\new_[20444]_  | ~\new_[20439]_  | ~\new_[20437]_  | ~\new_[20438]_ ;
  assign \new_[20437]_  = ~\new_[19812]_  | (~\new_[3925]_  & ~\new_[7156]_ );
  assign \new_[20438]_  = \new_[19961]_  & \new_[19965]_ ;
  assign \new_[20439]_  = ~\new_[958]_  | (~\new_[20440]_  & ~\new_[20442]_ );
  assign \new_[20440]_  = ~\new_[20441]_  | ~\new_[4689]_  | ~\new_[5423]_ ;
  assign \new_[20441]_  = ~\new_[9018]_ ;
  assign \new_[20442]_  = ~\new_[12349]_  | ~\new_[20443]_  | ~\new_[9028]_ ;
  assign \new_[20443]_  = ~\new_[6599]_  | ~\new_[19334]_ ;
  assign \new_[20444]_  = \new_[19964]_  & \new_[19968]_ ;
  assign \new_[20445]_  = ~\new_[20450]_  & (~\new_[964]_  | ~\new_[20446]_ );
  assign \new_[20446]_  = ~\new_[20449]_  | ~\new_[20448]_  | ~\new_[4695]_  | ~\new_[20447]_ ;
  assign \new_[20447]_  = ~\new_[19163]_  | ~\new_[4030]_ ;
  assign \new_[20448]_  = ~\new_[4411]_ ;
  assign \new_[20449]_  = ~\new_[7904]_  & ~\new_[8704]_ ;
  assign \new_[20450]_  = ~\new_[20451]_  | ~\new_[3774]_  | ~\new_[4091]_ ;
  assign \new_[20451]_  = \new_[6699]_  & \new_[5425]_ ;
  assign \new_[20452]_  = ~\new_[964]_ ;
  assign \new_[20453]_  = ~\new_[20454]_  | ~\new_[20456]_ ;
  assign \new_[20454]_  = ~\new_[20455]_  | ~\new_[20645]_ ;
  assign \new_[20455]_  = ~\new_[11879]_  | ~\new_[13315]_ ;
  assign \new_[20456]_  = ~\new_[20457]_  & (~\new_[11385]_  | ~\new_[18031]_ );
  assign \new_[20457]_  = \new_[13791]_  & \new_[18031]_ ;
  assign \new_[20458]_  = ~\new_[20457]_ ;
  assign \new_[20459]_  = ~\new_[20468]_  | ~\new_[20467]_  | ~\new_[20465]_  | ~\new_[20460]_ ;
  assign \new_[20460]_  = ~\new_[20464]_  | (~\new_[20461]_  & ~\new_[20462]_ );
  assign \new_[20461]_  = ~\new_[4803]_  | ~\new_[4937]_ ;
  assign \new_[20462]_  = ~\new_[6405]_  | ~\new_[20463]_ ;
  assign \new_[20463]_  = ~\new_[14774]_  | ~\new_[17441]_ ;
  assign \new_[20464]_  = ~\new_[950]_ ;
  assign \new_[20465]_  = ~\new_[21142]_  | (~\new_[4560]_  & ~\new_[20466]_ );
  assign \new_[20466]_  = ~\new_[20463]_ ;
  assign \new_[20467]_  = ~\new_[19467]_  | (~\new_[5122]_  & ~\new_[10908]_ );
  assign \new_[20468]_  = ~\new_[20469]_ ;
  assign \new_[20469]_  = ~\new_[21142]_  & ~\new_[5500]_ ;
  assign \new_[20470]_  = ~\new_[6035]_ ;
  assign \new_[20471]_  = ~\new_[20472]_  & ~\new_[7161]_ ;
  assign \new_[20472]_  = ~\new_[20422]_ ;
  assign \new_[20473]_  = \new_[6511]_  & \new_[8502]_ ;
  assign \new_[20474]_  = ~\new_[20477]_  | ~\new_[20475]_  | ~\new_[20476]_ ;
  assign \new_[20475]_  = ~\new_[935]_  | (~\new_[4741]_  & ~\new_[4586]_ );
  assign \new_[20476]_  = ~\new_[19564]_  | (~\new_[4206]_  & ~\new_[8171]_ );
  assign \new_[20477]_  = ~\new_[20478]_  & (~\new_[4752]_  | ~\new_[19049]_ );
  assign \new_[20478]_  = ~\new_[11910]_  | ~\new_[20481]_  | ~\new_[20479]_  | ~\new_[9679]_ ;
  assign \new_[20479]_  = ~\new_[20480]_ ;
  assign \new_[20480]_  = ~\new_[19702]_  & ~\new_[7666]_ ;
  assign \new_[20481]_  = ~\new_[20482]_  & (~\new_[11237]_  | ~\new_[17714]_ );
  assign \new_[20482]_  = ~\new_[10994]_  & ~\new_[18124]_ ;
  assign \new_[20483]_  = ~\new_[20482]_ ;
  assign \new_[20484]_  = ~\new_[20485]_  & ~\new_[20488]_ ;
  assign \new_[20485]_  = ~\new_[20486]_ ;
  assign \new_[20486]_  = ~\new_[20487]_ ;
  assign \new_[20487]_  = ~\new_[993]_ ;
  assign \new_[20488]_  = ~\new_[20489]_  | ~\new_[20490]_ ;
  assign \new_[20489]_  = ~\new_[17678]_  & ~\new_[21517]_ ;
  assign \new_[20490]_  = ~\new_[20491]_ ;
  assign \new_[20491]_  = \new_[952]_ ;
  assign \new_[20492]_  = ~\new_[20486]_ ;
  assign \new_[20493]_  = ~\new_[952]_ ;
  assign \new_[20494]_  = ~\new_[20495]_  & ~\new_[20496]_ ;
  assign \new_[20495]_  = ~\new_[1002]_ ;
  assign \new_[20496]_  = ~\new_[20497]_  | ~\new_[996]_ ;
  assign \new_[20497]_  = ~\new_[1003]_ ;
  assign \new_[20498]_  = ~\new_[20497]_ ;
  assign \new_[20499]_  = \new_[20751]_ ;
  assign \new_[20500]_  = ~\new_[20501]_  & ~\new_[20504]_ ;
  assign \new_[20501]_  = ~\new_[20502]_  | ~\new_[20503]_ ;
  assign \new_[20502]_  = ~\new_[5751]_  | ~\new_[17723]_ ;
  assign \new_[20503]_  = ~\new_[7954]_  | ~\new_[19357]_ ;
  assign \new_[20504]_  = ~\new_[6542]_  | ~\new_[20014]_  | ~\new_[5220]_ ;
  assign \new_[20505]_  = ~\new_[20506]_ ;
  assign \new_[20506]_  = ~\new_[20507]_  | ~\new_[20508]_ ;
  assign \new_[20507]_  = ~\new_[930]_ ;
  assign \new_[20508]_  = ~\new_[4973]_  | ~\new_[20514]_  | ~\new_[20509]_  | ~\new_[4740]_ ;
  assign \new_[20509]_  = ~\new_[20510]_  | ~\new_[20513]_ ;
  assign \new_[20510]_  = ~\new_[20511]_  | ~\new_[20512]_ ;
  assign \new_[20511]_  = ~\new_[11772]_  & ~\new_[7020]_ ;
  assign \new_[20512]_  = ~\new_[12122]_  & ~\new_[13346]_ ;
  assign \new_[20513]_  = ~\new_[1033]_ ;
  assign \new_[20514]_  = ~\new_[20515]_  & ~\new_[20516]_ ;
  assign \new_[20515]_  = ~\new_[12153]_ ;
  assign \new_[20516]_  = ~\new_[17273]_  & ~\new_[7705]_ ;
  assign \new_[20517]_  = ~\new_[20521]_  | ~\new_[20520]_  | ~\new_[20518]_  | ~\new_[20519]_ ;
  assign \new_[20518]_  = ~\new_[21634]_  | (~\new_[12889]_  & ~\new_[20925]_ );
  assign \new_[20519]_  = ~\new_[16501]_  | ~\new_[21638]_ ;
  assign \new_[20520]_  = ~\new_[21635]_  | ~\new_[20930]_  | ~\new_[19476]_ ;
  assign \new_[20521]_  = ~\new_[14569]_  | ~\new_[21637]_  | ~\new_[19750]_ ;
  assign \new_[20522]_  = ~\new_[19750]_  | ~\new_[14569]_ ;
  assign \new_[20523]_  = ~\new_[20530]_  | ~\new_[20524]_  | ~\new_[20529]_ ;
  assign \new_[20524]_  = ~\new_[20525]_  | ~\new_[20526]_ ;
  assign \new_[20525]_  = ~\new_[1004]_  | ~\new_[4108]_  | ~\new_[4298]_ ;
  assign \new_[20526]_  = ~\new_[20528]_  | ~\new_[5265]_  | ~\new_[20527]_  | ~\new_[4480]_ ;
  assign \new_[20527]_  = \new_[5919]_  & \new_[5453]_ ;
  assign \new_[20528]_  = ~\new_[1004]_ ;
  assign \new_[20529]_  = ~\new_[4280]_ ;
  assign \new_[20530]_  = ~\new_[20531]_  & ~\new_[5422]_ ;
  assign \new_[20531]_  = ~\new_[20533]_  | ~\new_[9489]_  | ~\new_[7364]_  | ~\new_[20532]_ ;
  assign \new_[20532]_  = ~\new_[11645]_  | ~\new_[18941]_ ;
  assign \new_[20533]_  = ~\new_[7461]_ ;
  assign \new_[20534]_  = ~\new_[21071]_  & (~\new_[20538]_  | ~\new_[20535]_ );
  assign \new_[20535]_  = ~\new_[20536]_  | ~\new_[20537]_ ;
  assign \new_[20536]_  = ~\new_[9985]_  | ~\new_[5781]_  | ~\new_[8976]_ ;
  assign \new_[20537]_  = ~\new_[946]_ ;
  assign \new_[20538]_  = ~\new_[20696]_  & ~\new_[21038]_ ;
  assign \new_[20539]_  = ~\new_[20544]_  | ~\new_[20542]_  | ~\new_[20540]_  | ~\new_[20541]_ ;
  assign \new_[20540]_  = ~\new_[958]_  | (~\new_[3960]_  & ~\new_[5406]_ );
  assign \new_[20541]_  = ~\new_[20645]_  | (~\new_[4318]_  & ~\new_[11603]_ );
  assign \new_[20542]_  = ~\new_[20543]_  & (~\new_[4249]_  | ~\new_[20743]_ );
  assign \new_[20543]_  = ~\new_[5189]_  | ~\new_[5994]_ ;
  assign \new_[20544]_  = \new_[6698]_  & \new_[5503]_ ;
  assign \new_[20545]_  = \new_[3462]_  ? \new_[20547]_  : \new_[20546]_ ;
  assign \new_[20546]_  = ~\new_[19865]_  | ~\new_[19867]_ ;
  assign \new_[20547]_  = ~\new_[20548]_  & ~\new_[20549]_ ;
  assign \new_[20548]_  = ~\new_[3762]_  | ~\new_[3831]_ ;
  assign \new_[20549]_  = ~\new_[4015]_  | ~\new_[4200]_ ;
  assign \new_[20550]_  = ~\new_[3831]_  | ~\new_[3762]_  | ~\new_[4015]_  | ~\new_[4200]_ ;
  assign \new_[20551]_  = ~\new_[20554]_  | ~\new_[20552]_  | ~\new_[20553]_ ;
  assign \new_[20552]_  = ~\new_[7715]_  & (~\new_[8546]_  | ~\new_[18759]_ );
  assign \new_[20553]_  = ~\new_[6810]_  | ~\new_[21559]_ ;
  assign \new_[20554]_  = ~\new_[20555]_  & (~\new_[9251]_  | ~\new_[19619]_ );
  assign \new_[20555]_  = \new_[8797]_  | \new_[20556]_ ;
  assign \new_[20556]_  = ~\new_[20557]_  & ~\new_[21559]_ ;
  assign \new_[20557]_  = ~\new_[19462]_  | ~\new_[15202]_ ;
  assign \new_[20558]_  = ~\new_[20557]_ ;
  assign \new_[20559]_  = ~\new_[20560]_  | ~\new_[20564]_ ;
  assign \new_[20560]_  = ~\new_[20561]_  & ~\new_[20562]_ ;
  assign \new_[20561]_  = ~\new_[19816]_  & ~\new_[3862]_ ;
  assign \new_[20562]_  = ~\new_[3949]_  | ~\new_[20563]_ ;
  assign \new_[20563]_  = \new_[10897]_  ? \new_[19711]_  : \new_[12717]_ ;
  assign \new_[20564]_  = ~\new_[20566]_  & (~\new_[20565]_  | ~\new_[19262]_ );
  assign \new_[20565]_  = \new_[7353]_  | \new_[4668]_ ;
  assign \new_[20566]_  = ~\new_[19262]_  & (~\new_[5293]_  | ~\new_[19951]_ );
  assign \new_[20567]_  = \new_[20568]_ ;
  assign \new_[20568]_  = ~\new_[20574]_  | ~\new_[20571]_  | ~\new_[20569]_  | ~\new_[20570]_ ;
  assign \new_[20569]_  = ~\new_[935]_  | (~\new_[4592]_  & ~\new_[4684]_ );
  assign \new_[20570]_  = ~\new_[19564]_  | (~\new_[4203]_  & ~\new_[5974]_ );
  assign \new_[20571]_  = ~\new_[20572]_  & (~\new_[4673]_  | ~\new_[18386]_ );
  assign \new_[20572]_  = ~\new_[11209]_  | ~\new_[20573]_  | ~\new_[7871]_ ;
  assign \new_[20573]_  = ~\new_[17252]_  | ~\new_[6068]_ ;
  assign \new_[20574]_  = ~\new_[20575]_  & ~\new_[20576]_ ;
  assign \new_[20575]_  = ~\new_[18292]_  & (~\new_[11356]_  | ~\new_[8640]_ );
  assign \new_[20576]_  = ~\new_[19702]_  & (~\new_[7040]_  | ~\new_[13150]_ );
  assign \new_[20577]_  = ~\new_[20578]_ ;
  assign \new_[20578]_  = ~\new_[20579]_  | ~\new_[20584]_ ;
  assign \new_[20579]_  = ~\new_[20580]_  & ~\new_[20581]_ ;
  assign \new_[20580]_  = ~\new_[8479]_  | ~\new_[14085]_ ;
  assign \new_[20581]_  = ~\new_[20582]_  | ~\new_[20583]_ ;
  assign \new_[20582]_  = ~\new_[4340]_  | ~\new_[19740]_ ;
  assign \new_[20583]_  = ~\new_[4053]_  | ~\new_[19795]_ ;
  assign \new_[20584]_  = ~\new_[4083]_  & ~\new_[20585]_ ;
  assign \new_[20585]_  = ~\new_[19786]_  & (~\new_[6011]_  | ~\new_[4278]_ );
  assign \new_[20586]_  = ~\new_[19689]_  & ~\new_[20587]_ ;
  assign \new_[20587]_  = \new_[20588]_  | \new_[20590]_ ;
  assign \new_[20588]_  = \new_[20589]_ ;
  assign \new_[20589]_  = ~\new_[1023]_ ;
  assign \new_[20590]_  = \new_[1079]_ ;
  assign \new_[20591]_  = \new_[20588]_  | \new_[20590]_ ;
  assign \new_[20592]_  = ~\new_[20595]_  | (~\new_[20593]_  & ~\new_[20594]_ );
  assign \new_[20593]_  = \new_[3400]_  ^ \new_[2728]_ ;
  assign \new_[20594]_  = \new_[3316]_  ? \new_[2357]_  : \new_[3513]_ ;
  assign \new_[20595]_  = ~\new_[20594]_  | ~\new_[20593]_ ;
  assign \new_[20596]_  = ~\new_[20602]_  | ~\new_[20600]_  | ~\new_[20598]_  | ~\new_[20597]_ ;
  assign \new_[20597]_  = ~\new_[19816]_  | (~\new_[3962]_  & ~\new_[6540]_ );
  assign \new_[20598]_  = ~\new_[979]_  | ~\new_[20599]_ ;
  assign \new_[20599]_  = ~\new_[7814]_  | ~\new_[5022]_  | ~\new_[4907]_  | ~\new_[4465]_ ;
  assign \new_[20600]_  = ~\new_[20601]_ ;
  assign \new_[20601]_  = ~\new_[5017]_  | ~\new_[4927]_  | ~\new_[5995]_ ;
  assign \new_[20602]_  = ~\new_[19517]_  | (~\new_[5124]_  & ~\new_[5589]_ );
  assign \new_[20603]_  = ~\new_[20610]_  | ~\new_[20609]_  | ~\new_[20604]_  | ~\new_[20608]_ ;
  assign \new_[20604]_  = ~\new_[21205]_  | ~\new_[20605]_ ;
  assign \new_[20605]_  = ~\new_[20607]_  | ~\new_[20606]_  | ~\new_[4658]_  | ~\new_[4215]_ ;
  assign \new_[20606]_  = \new_[6505]_  & \new_[12701]_ ;
  assign \new_[20607]_  = ~\new_[10131]_  & ~\new_[10844]_ ;
  assign \new_[20608]_  = ~\new_[994]_  | (~\new_[4170]_  & ~\new_[4970]_ );
  assign \new_[20609]_  = ~\new_[4584]_ ;
  assign \new_[20610]_  = ~\new_[20611]_  & ~\new_[4186]_ ;
  assign \new_[20611]_  = ~\new_[8282]_  | ~\new_[11261]_ ;
  assign \new_[20612]_  = ~\new_[20614]_  | ~\new_[20613]_ ;
  assign \new_[20613]_  = (~\new_[937]_  | ~\new_[3938]_ ) & (~\new_[4605]_  | ~\new_[18844]_ );
  assign \new_[20614]_  = ~\new_[4124]_  & (~\new_[21425]_  | ~\new_[3922]_ );
  assign \new_[20615]_  = ~\new_[19787]_  | (~\new_[4315]_  & ~\new_[12518]_ );
  assign \new_[20616]_  = ~\new_[19517]_  | (~\new_[6020]_  & ~\new_[21623]_ );
  assign \new_[20617]_  = \new_[20618]_  & \new_[20619]_ ;
  assign \new_[20618]_  = ~\new_[9104]_  | ~\new_[20621]_ ;
  assign \new_[20619]_  = ~\new_[20620]_  | ~\new_[20621]_ ;
  assign \new_[20620]_  = ~\new_[17598]_  & ~\new_[14664]_ ;
  assign \new_[20621]_  = ~\new_[19242]_  & ~\new_[19450]_ ;
  assign \new_[20622]_  = ~\new_[20621]_ ;
  assign \new_[20623]_  = ~\new_[20627]_  | ~\new_[5008]_  | ~\new_[20624]_  | ~\new_[20626]_ ;
  assign \new_[20624]_  = ~\new_[20625]_ ;
  assign \new_[20625]_  = ~\new_[930]_  & (~\new_[4383]_  | ~\new_[5235]_ );
  assign \new_[20626]_  = \new_[4043]_  & \new_[4114]_ ;
  assign \new_[20627]_  = ~\new_[20628]_ ;
  assign \new_[20628]_  = ~\new_[10255]_  | ~\new_[11848]_  | ~\new_[8156]_  | ~\new_[11728]_ ;
  assign \new_[20629]_  = ~\new_[20635]_  | ~\new_[20634]_  | ~\new_[20630]_  | ~\new_[20633]_ ;
  assign \new_[20630]_  = ~\new_[20631]_  | ~\new_[938]_ ;
  assign \new_[20631]_  = ~\new_[6900]_  | ~\new_[20632]_  | ~\new_[4688]_  | ~\new_[4459]_ ;
  assign \new_[20632]_  = \new_[8081]_  & \new_[8145]_ ;
  assign \new_[20633]_  = ~\new_[21441]_  | ~\new_[4102]_ ;
  assign \new_[20634]_  = ~\new_[18409]_  | (~\new_[4023]_  & ~\new_[11682]_ );
  assign \new_[20635]_  = ~\new_[20636]_  & ~\new_[20637]_ ;
  assign \new_[20636]_  = ~\new_[4659]_  | ~\new_[6790]_ ;
  assign \new_[20637]_  = ~\new_[5985]_  | ~\new_[7480]_ ;
  assign \new_[20638]_  = ~\new_[19812]_  & (~\new_[20639]_  | ~\new_[20642]_ );
  assign \new_[20639]_  = ~\new_[20640]_  | ~\new_[20641]_ ;
  assign \new_[20640]_  = ~\new_[8788]_  | ~\new_[7841]_  | ~\new_[5342]_ ;
  assign \new_[20641]_  = ~\new_[954]_ ;
  assign \new_[20642]_  = ~\new_[20643]_  & ~\new_[20644]_ ;
  assign \new_[20643]_  = ~\new_[19072]_  & ~\new_[6751]_ ;
  assign \new_[20644]_  = ~\new_[7857]_  | ~\new_[20961]_  | ~\new_[5286]_ ;
  assign \new_[20645]_  = ~\new_[954]_ ;
  assign \new_[20646]_  = ~\new_[20647]_  | ~\new_[20648]_ ;
  assign \new_[20647]_  = \new_[3958]_  & \new_[3773]_ ;
  assign \new_[20648]_  = ~\new_[20649]_  & ~\new_[20652]_ ;
  assign \new_[20649]_  = ~\new_[20650]_ ;
  assign \new_[20650]_  = ~\new_[20651]_  & (~\new_[4176]_  | ~\new_[18409]_ );
  assign \new_[20651]_  = \new_[5199]_  & \new_[18583]_ ;
  assign \new_[20652]_  = ~\new_[20653]_  | (~\new_[13582]_  & ~\new_[21557]_ );
  assign \new_[20653]_  = ~\new_[21562]_  | ~\new_[20654]_ ;
  assign \new_[20654]_  = ~\new_[12682]_ ;
  assign \new_[20655]_  = ~\new_[20659]_  | ~\new_[3766]_  | ~\new_[20656]_  | ~\new_[4223]_ ;
  assign \new_[20656]_  = ~\new_[20657]_  & (~\new_[4292]_  | ~\new_[19032]_ );
  assign \new_[20657]_  = ~\new_[20528]_  & (~\new_[4703]_  | ~\new_[20658]_ );
  assign \new_[20658]_  = \new_[4881]_  & \new_[5660]_ ;
  assign \new_[20659]_  = \new_[6632]_  & \new_[11833]_ ;
  assign \new_[20660]_  = ~\new_[20661]_  | ~\new_[20663]_ ;
  assign \new_[20661]_  = ~\new_[20662]_ ;
  assign \new_[20662]_  = ~\new_[21307]_  | ~\new_[21686]_ ;
  assign \new_[20663]_  = ~\new_[20664]_ ;
  assign \new_[20664]_  = ~\new_[20665]_  | ~\new_[21657]_ ;
  assign \new_[20665]_  = ~\new_[20666]_ ;
  assign \new_[20666]_  = ~\new_[19494]_  | ~\new_[19683]_ ;
  assign \new_[20667]_  = ~\new_[20668]_  | ~\new_[20672]_ ;
  assign \new_[20668]_  = ~\new_[20669]_  & (~\new_[930]_  | ~\new_[4058]_ );
  assign \new_[20669]_  = ~\new_[20670]_  | ~\new_[20671]_ ;
  assign \new_[20670]_  = ~\new_[4755]_  | ~\new_[19523]_ ;
  assign \new_[20671]_  = (~\new_[16279]_  | ~\new_[18855]_ ) & (~\new_[10242]_  | ~\new_[17273]_ );
  assign \new_[20672]_  = (~\new_[19585]_  | ~\new_[4227]_ ) & (~\new_[4351]_  | ~\new_[19157]_ );
  assign \new_[20673]_  = ~\new_[19229]_  & ~\new_[9667]_ ;
  assign \new_[20674]_  = ~\new_[18084]_  & (~\new_[6767]_  | ~\new_[12845]_ );
  assign \new_[20675]_  = ~\new_[20685]_  | ~\new_[20676]_  | ~\new_[20677]_ ;
  assign \new_[20676]_  = ~\new_[19694]_  | (~\new_[5857]_  & ~\new_[7613]_ );
  assign \new_[20677]_  = ~\new_[20682]_  & (~\new_[20678]_  | ~\new_[20679]_ );
  assign \new_[20678]_  = ~\new_[7212]_  | ~\new_[13938]_ ;
  assign \new_[20679]_  = ~\new_[20680]_ ;
  assign \new_[20680]_  = \new_[20681]_ ;
  assign \new_[20681]_  = ~\new_[1041]_ ;
  assign \new_[20682]_  = ~\new_[15485]_  | ~\new_[20683]_  | ~\new_[9796]_ ;
  assign \new_[20683]_  = ~\new_[20684]_ ;
  assign \new_[20684]_  = ~\new_[20679]_  & (~\new_[14631]_  | ~\new_[13989]_ );
  assign \new_[20685]_  = ~\new_[19453]_  | (~\new_[10448]_  & ~\new_[13034]_ );
  assign \new_[20686]_  = ~\new_[20681]_ ;
  assign \new_[20687]_  = ~\new_[20693]_  | ~\new_[20692]_  | ~\new_[20688]_  | ~\new_[20690]_ ;
  assign \new_[20688]_  = ~\new_[20689]_  | ~\new_[979]_ ;
  assign \new_[20689]_  = ~\new_[4111]_  | ~\new_[4154]_ ;
  assign \new_[20690]_  = ~\new_[20691]_  | ~\new_[19816]_ ;
  assign \new_[20691]_  = ~\new_[5653]_  | ~\new_[5933]_  | ~\new_[4489]_  | ~\new_[5957]_ ;
  assign \new_[20692]_  = ~\new_[4490]_  & ~\new_[5869]_ ;
  assign \new_[20693]_  = ~\new_[20694]_ ;
  assign \new_[20694]_  = ~\new_[7602]_  | ~\new_[6608]_  | ~\new_[20695]_ ;
  assign \new_[20695]_  = ~\new_[7508]_  & (~\new_[21623]_  | ~\new_[19711]_ );
  assign \new_[20696]_  = ~\new_[20702]_  | (~\new_[20697]_  & ~\new_[16879]_ );
  assign \new_[20697]_  = ~\new_[20700]_  & (~\new_[20698]_  | ~\new_[18624]_ );
  assign \new_[20698]_  = ~\new_[13356]_  | ~\new_[15269]_ ;
  assign \new_[20699]_  = ~\new_[21402]_ ;
  assign \new_[20700]_  = ~\new_[20699]_  & ~\new_[15156]_ ;
  assign \new_[20701]_  = \new_[1082]_ ;
  assign \new_[20702]_  = ~\new_[20703]_ ;
  assign \new_[20703]_  = ~\new_[21498]_  & ~\new_[12820]_ ;
  assign \new_[20704]_  = ~\new_[1082]_ ;
  assign \new_[20705]_  = ~\new_[20700]_ ;
  assign \new_[20706]_  = ~\new_[20711]_  | ~\new_[20707]_  | ~\new_[20710]_ ;
  assign \new_[20707]_  = ~\new_[20708]_  & ~\new_[20709]_ ;
  assign \new_[20708]_  = ~\new_[18693]_  & (~\new_[10140]_  | ~\new_[16291]_ );
  assign \new_[20709]_  = ~\new_[13750]_  & ~\new_[19151]_ ;
  assign \new_[20710]_  = ~\new_[11941]_  | ~\new_[18693]_ ;
  assign \new_[20711]_  = \new_[20712]_  & \new_[20713]_ ;
  assign \new_[20712]_  = ~\new_[14388]_  | ~\new_[18840]_ ;
  assign \new_[20713]_  = \new_[19409]_  | \new_[16232]_ ;
  assign \new_[20714]_  = ~\new_[20709]_ ;
  assign \new_[20715]_  = ~\new_[20713]_ ;
  assign \new_[20716]_  = ~\new_[20718]_  | (~\new_[20717]_  & ~\new_[18739]_ );
  assign \new_[20717]_  = ~\new_[9338]_  & ~\new_[6794]_ ;
  assign \new_[20718]_  = ~\new_[20721]_  & (~\new_[20719]_  | ~\new_[18739]_ );
  assign \new_[20719]_  = ~\new_[20720]_ ;
  assign \new_[20720]_  = ~\new_[14608]_  | ~\new_[18423]_ ;
  assign \new_[20721]_  = ~\new_[8801]_  | ~\new_[20722]_  | ~\new_[7807]_ ;
  assign \new_[20722]_  = ~\new_[20723]_ ;
  assign \new_[20723]_  = ~\new_[18973]_  & ~\new_[13789]_ ;
  assign \new_[20724]_  = ~\new_[20725]_  & ~\new_[20726]_ ;
  assign \new_[20725]_  = \new_[19271]_  | \new_[18941]_ ;
  assign \new_[20726]_  = \new_[18166]_  | \new_[11703]_ ;
  assign \new_[20727]_  = ~\new_[20728]_  | ~\new_[20733]_  | ~\new_[20730]_  | ~\new_[20729]_ ;
  assign \new_[20728]_  = ~\new_[7537]_  & (~\new_[21324]_  | ~\new_[18124]_ );
  assign \new_[20729]_  = ~\new_[8068]_ ;
  assign \new_[20730]_  = ~\new_[20731]_ ;
  assign \new_[20731]_  = ~\new_[7237]_  | ~\new_[20732]_ ;
  assign \new_[20732]_  = \new_[15369]_  & \new_[16552]_ ;
  assign \new_[20733]_  = ~\new_[19702]_  | (~\new_[21319]_  & ~\new_[20734]_ );
  assign \new_[20734]_  = ~\new_[10750]_  | ~\new_[12001]_ ;
  assign \new_[20735]_  = ~\new_[20744]_  | ~\new_[20738]_  | ~\new_[20736]_  | ~\new_[20737]_ ;
  assign \new_[20736]_  = ~\new_[3782]_  | ~\new_[19273]_ ;
  assign \new_[20737]_  = \new_[4199]_  & \new_[4026]_ ;
  assign \new_[20738]_  = ~\new_[20743]_  | (~\new_[20739]_  & ~\new_[20741]_ );
  assign \new_[20739]_  = ~\new_[4662]_  | ~\new_[20740]_ ;
  assign \new_[20740]_  = \new_[9204]_  & \new_[8596]_ ;
  assign \new_[20741]_  = ~\new_[4967]_  | ~\new_[20742]_ ;
  assign \new_[20742]_  = ~\new_[19436]_  | (~\new_[6731]_  & ~\new_[12813]_ );
  assign \new_[20743]_  = ~\new_[958]_ ;
  assign \new_[20744]_  = ~\new_[20745]_ ;
  assign \new_[20745]_  = ~\new_[7310]_  | ~\new_[11556]_  | ~\new_[7580]_ ;
  assign \new_[20746]_  = ~\new_[1002]_ ;
  assign \new_[20747]_  = ~\new_[20497]_  | ~\new_[20748]_  | ~\new_[19488]_ ;
  assign \new_[20748]_  = \new_[996]_ ;
  assign \new_[20749]_  = \new_[20746]_ ;
  assign \new_[20750]_  = ~\new_[20497]_  | ~\new_[19488]_ ;
  assign \new_[20751]_  = ~\new_[996]_ ;
  assign \new_[20752]_  = ~\new_[20753]_  | ~\new_[20754]_ ;
  assign \new_[20753]_  = ~\new_[21386]_  | ~\new_[5763]_  | ~\new_[4932]_  | ~\new_[4910]_ ;
  assign \new_[20754]_  = ~\new_[19989]_  | ~\new_[20755]_  | ~\new_[19987]_ ;
  assign \new_[20755]_  = ~\new_[20756]_  & ~\new_[20757]_ ;
  assign \new_[20756]_  = ~\new_[19990]_  | ~\new_[940]_ ;
  assign \new_[20757]_  = ~\new_[19992]_ ;
  assign \new_[20758]_  = ~\new_[20759]_  | ~\new_[20760]_ ;
  assign \new_[20759]_  = ~\new_[6196]_  | ~\new_[973]_ ;
  assign \new_[20760]_  = ~\new_[20763]_  | (~\new_[20761]_  & ~\new_[20762]_ );
  assign \new_[20761]_  = ~\new_[12469]_  | ~\new_[11342]_  | ~\new_[12204]_ ;
  assign \new_[20762]_  = ~\new_[10944]_  | ~\new_[13051]_ ;
  assign \new_[20763]_  = ~\new_[973]_ ;
  assign \new_[20764]_  = ~\new_[20765]_  | ~\new_[20767]_ ;
  assign \new_[20765]_  = ~\new_[20766]_ ;
  assign \new_[20766]_  = ~\new_[19522]_  | ~\new_[20302]_ ;
  assign \new_[20767]_  = ~\new_[1023]_ ;
  assign \new_[20768]_  = ~\new_[20769]_ ;
  assign \new_[20769]_  = ~\new_[19568]_  & ~\new_[19689]_ ;
  assign \new_[20770]_  = ~\new_[20764]_ ;
  assign \new_[20771]_  = ~\new_[19522]_  | ~\new_[20302]_ ;
  assign \new_[20772]_  = ~\new_[20773]_  | ~\new_[20778]_ ;
  assign \new_[20773]_  = ~\new_[20774]_  & (~\new_[6775]_  | ~\new_[19170]_ );
  assign \new_[20774]_  = ~\new_[4862]_  | ~\new_[20775]_ ;
  assign \new_[20775]_  = ~\new_[20776]_  & ~\new_[20777]_ ;
  assign \new_[20776]_  = ~\new_[21562]_  & ~\new_[9900]_ ;
  assign \new_[20777]_  = ~\new_[8714]_  | ~\new_[11636]_ ;
  assign \new_[20778]_  = ~\new_[20779]_  & ~\new_[4603]_ ;
  assign \new_[20779]_  = ~\new_[6510]_  | ~\new_[20780]_ ;
  assign \new_[20780]_  = \new_[21562]_  | \new_[9218]_ ;
  assign \new_[20781]_  = ~\new_[20776]_ ;
  assign \new_[20782]_  = ~\new_[20783]_  & ~\new_[20784]_ ;
  assign \new_[20783]_  = ~\new_[930]_ ;
  assign \new_[20784]_  = ~\new_[20790]_  & (~\new_[20785]_  | ~\new_[20787]_ );
  assign \new_[20785]_  = ~\new_[8515]_  | ~\new_[9936]_  | ~\new_[20786]_  | ~\new_[8083]_ ;
  assign \new_[20786]_  = \new_[9907]_  & \new_[1033]_ ;
  assign \new_[20787]_  = ~\new_[20788]_  | ~\new_[9042]_  | ~\new_[8736]_ ;
  assign \new_[20788]_  = \new_[10255]_  & \new_[20789]_ ;
  assign \new_[20789]_  = ~\new_[1033]_ ;
  assign \new_[20790]_  = ~\new_[20791]_  | ~\new_[6513]_  | ~\new_[7805]_ ;
  assign \new_[20791]_  = \new_[9887]_  & \new_[10266]_ ;
  assign \new_[20792]_  = ~\new_[20795]_  & (~\new_[20793]_  | ~\new_[20794]_ );
  assign \new_[20793]_  = ~\new_[4171]_  | ~\new_[5112]_ ;
  assign \new_[20794]_  = ~\new_[20295]_ ;
  assign \new_[20795]_  = ~\new_[20803]_  | ~\new_[20796]_  | ~\new_[20800]_ ;
  assign \new_[20796]_  = ~\new_[20797]_  & ~\new_[20798]_ ;
  assign \new_[20797]_  = ~\new_[6402]_  | ~\new_[6509]_ ;
  assign \new_[20798]_  = ~\new_[20799]_  | ~\new_[6012]_ ;
  assign \new_[20799]_  = ~\new_[5480]_  | ~\new_[18752]_ ;
  assign \new_[20800]_  = ~\new_[20801]_  & ~\new_[20296]_ ;
  assign \new_[20801]_  = ~\new_[20802]_ ;
  assign \new_[20802]_  = ~\new_[18818]_  | ~\new_[14080]_ ;
  assign \new_[20803]_  = ~\new_[20804]_  | ~\new_[18759]_ ;
  assign \new_[20804]_  = ~\new_[9032]_  | ~\new_[8002]_ ;
  assign \new_[20805]_  = ~\new_[20806]_  | ~\new_[20807]_ ;
  assign \new_[20806]_  = ~\new_[9597]_  | ~\new_[18361]_ ;
  assign \new_[20807]_  = \new_[21504]_  | \new_[20808]_ ;
  assign \new_[20808]_  = ~\new_[14596]_  | ~\new_[18394]_ ;
  assign \new_[20809]_  = \new_[20808]_ ;
  assign \new_[20810]_  = ~\new_[20818]_  | ~\new_[20811]_  | ~\new_[20817]_ ;
  assign \new_[20811]_  = ~\new_[20812]_  | ~\new_[20815]_ ;
  assign \new_[20812]_  = ~\new_[20813]_  | ~\new_[20814]_ ;
  assign \new_[20813]_  = ~\new_[4256]_ ;
  assign \new_[20814]_  = ~\new_[19736]_  & ~\new_[5601]_ ;
  assign \new_[20815]_  = ~\new_[21066]_  | ~\new_[6724]_  | ~\new_[20816]_  | ~\new_[4864]_ ;
  assign \new_[20816]_  = \new_[7206]_  & \new_[12117]_ ;
  assign \new_[20817]_  = ~\new_[4286]_  | ~\new_[18612]_ ;
  assign \new_[20818]_  = ~\new_[20819]_  & ~\new_[4496]_ ;
  assign \new_[20819]_  = ~\new_[6733]_  | ~\new_[7879]_ ;
  assign \new_[20820]_  = ~\new_[20821]_  | ~\new_[20823]_ ;
  assign \new_[20821]_  = ~\new_[20822]_  & (~\new_[10009]_  | ~\new_[19208]_ );
  assign \new_[20822]_  = ~\new_[20971]_  & ~\new_[18693]_ ;
  assign \new_[20823]_  = ~\new_[20824]_  | ~\new_[20825]_ ;
  assign \new_[20824]_  = ~\new_[15997]_  | ~\new_[10171]_  | ~\new_[13433]_ ;
  assign \new_[20825]_  = \new_[19791]_  & \new_[19687]_ ;
  assign \new_[20826]_  = ~\new_[10009]_  | ~\new_[19208]_ ;
  assign \new_[20827]_  = ~\new_[20822]_ ;
  assign \new_[20828]_  = ~\new_[20829]_  & ~\new_[20832]_ ;
  assign \new_[20829]_  = ~\new_[20830]_  | ~\new_[20831]_ ;
  assign \new_[20830]_  = ~\new_[3969]_  | ~\new_[986]_ ;
  assign \new_[20831]_  = ~\new_[4250]_  | ~\new_[21180]_ ;
  assign \new_[20832]_  = ~\new_[6713]_  | ~\new_[20833]_  | ~\new_[4046]_ ;
  assign \new_[20833]_  = ~\new_[20834]_ ;
  assign \new_[20834]_  = ~\new_[5492]_  | ~\new_[4640]_  | ~\new_[20835]_ ;
  assign \new_[20835]_  = ~\new_[20836]_  & ~\new_[20837]_ ;
  assign \new_[20836]_  = ~\new_[18711]_  & ~\new_[13858]_ ;
  assign \new_[20837]_  = ~\new_[19215]_  & ~\new_[11462]_ ;
  assign \new_[20838]_  = ~\new_[20844]_  | ~\new_[20843]_  | ~\new_[20839]_  | ~\new_[20840]_ ;
  assign \new_[20839]_  = ~\new_[19527]_  | (~\new_[5600]_  & ~\new_[10429]_ );
  assign \new_[20840]_  = ~\new_[20841]_  | ~\new_[19145]_ ;
  assign \new_[20841]_  = ~\new_[7829]_  | ~\new_[12324]_ ;
  assign \new_[20842]_  = \new_[1027]_ ;
  assign \new_[20843]_  = ~\new_[19339]_  | (~\new_[5606]_  & ~\new_[8866]_ );
  assign \new_[20844]_  = ~\new_[16799]_  | ~\new_[18115]_ ;
  assign \new_[20845]_  = ~\new_[1027]_ ;
  assign \new_[20846]_  = ~\new_[20847]_  & ~\new_[20849]_ ;
  assign \new_[20847]_  = ~\new_[20848]_  | ~\new_[4209]_  | ~\new_[4477]_ ;
  assign \new_[20848]_  = \new_[11452]_  & \new_[8595]_ ;
  assign \new_[20849]_  = ~\new_[20850]_  & ~\new_[20852]_ ;
  assign \new_[20850]_  = ~\new_[4468]_  & ~\new_[20851]_ ;
  assign \new_[20851]_  = \new_[935]_  | \new_[8130]_ ;
  assign \new_[20852]_  = ~\new_[20853]_  & ~\new_[3957]_ ;
  assign \new_[20853]_  = \new_[19564]_  | \new_[6863]_ ;
  assign \new_[20854]_  = ~\new_[20859]_  | ~\new_[20855]_  | ~\new_[20858]_ ;
  assign \new_[20855]_  = ~\new_[4392]_  & ~\new_[20856]_ ;
  assign \new_[20856]_  = ~\new_[20857]_  | ~\new_[5040]_  | ~\new_[5311]_ ;
  assign \new_[20857]_  = ~\new_[6940]_  | ~\new_[18786]_ ;
  assign \new_[20858]_  = ~\new_[3919]_  | ~\new_[20283]_ ;
  assign \new_[20859]_  = ~\new_[20860]_  | ~\new_[949]_ ;
  assign \new_[20860]_  = ~\new_[11805]_  | ~\new_[4729]_  | ~\new_[20861]_  | ~\new_[4323]_ ;
  assign \new_[20861]_  = ~\new_[20862]_  & ~\new_[20863]_ ;
  assign \new_[20862]_  = ~\new_[18650]_  & (~\new_[7784]_  | ~\new_[11570]_ );
  assign \new_[20863]_  = ~\new_[6169]_ ;
  assign \new_[20864]_  = ~\new_[20865]_  & ~\new_[20866]_ ;
  assign \new_[20865]_  = ~\new_[995]_ ;
  assign \new_[20866]_  = ~\new_[20867]_  | ~\new_[20869]_ ;
  assign \new_[20867]_  = ~\new_[20868]_ ;
  assign \new_[20868]_  = ~\new_[21524]_  | ~\new_[18720]_ ;
  assign \new_[20869]_  = ~\new_[19139]_ ;
  assign \new_[20870]_  = \new_[20871]_ ;
  assign \new_[20871]_  = ~\new_[1138]_ ;
  assign \new_[20872]_  = \new_[20873]_ ;
  assign \new_[20873]_  = ~\new_[20876]_  | ~\new_[20874]_ ;
  assign \new_[20874]_  = ~\new_[20875]_  & (~\new_[4236]_  | ~\new_[19807]_ );
  assign \new_[20875]_  = ~\new_[6625]_  | ~\new_[5967]_  | ~\new_[4647]_  | ~\new_[5495]_ ;
  assign \new_[20876]_  = ~\new_[20879]_  & (~\new_[20877]_  | ~\new_[17020]_ );
  assign \new_[20877]_  = ~\new_[20878]_  | ~\new_[13789]_ ;
  assign \new_[20878]_  = ~\new_[4306]_ ;
  assign \new_[20879]_  = \new_[964]_  & \new_[20880]_ ;
  assign \new_[20880]_  = ~\new_[6867]_  | ~\new_[4954]_  | ~\new_[4126]_  | ~\new_[20881]_ ;
  assign \new_[20881]_  = \new_[5904]_  & \new_[10608]_ ;
  assign \new_[20882]_  = ~\new_[20885]_  | ~\new_[3763]_  | ~\new_[20883]_ ;
  assign \new_[20883]_  = (~\new_[19786]_  | ~\new_[4434]_ ) & (~\new_[20884]_  | ~\new_[19536]_ );
  assign \new_[20884]_  = \new_[21468]_  | \new_[5136]_ ;
  assign \new_[20885]_  = ~\new_[20886]_  & (~\new_[4773]_  | ~\new_[19002]_ );
  assign \new_[20886]_  = ~\new_[20887]_  | ~\new_[11631]_ ;
  assign \new_[20887]_  = \new_[16673]_  | \new_[21541]_  | \new_[18698]_  | \new_[18288]_ ;
  assign \new_[20888]_  = ~\new_[20893]_  | ~\new_[20892]_  | ~\new_[20889]_ ;
  assign \new_[20889]_  = ~\new_[20890]_  & ~\new_[20891]_ ;
  assign \new_[20890]_  = ~\new_[7568]_  | ~\new_[10575]_  | ~\new_[8223]_ ;
  assign \new_[20891]_  = ~\new_[4183]_  | ~\new_[4412]_ ;
  assign \new_[20892]_  = ~\new_[3784]_  | ~\new_[21385]_ ;
  assign \new_[20893]_  = ~\new_[21386]_  | (~\new_[20894]_  & ~\new_[20896]_ );
  assign \new_[20894]_  = ~\new_[20895]_  | ~\new_[4664]_ ;
  assign \new_[20895]_  = \new_[7557]_  & \new_[10442]_ ;
  assign \new_[20896]_  = ~\new_[4690]_  | ~\new_[20897]_ ;
  assign \new_[20897]_  = ~\new_[18569]_  | (~\new_[7560]_  & ~\new_[11634]_ );
  assign \new_[20898]_  = ~\new_[20906]_  | ~\new_[20904]_  | ~\new_[20899]_  | ~\new_[20900]_ ;
  assign \new_[20899]_  = ~\new_[17145]_  | ~\new_[19028]_ ;
  assign \new_[20900]_  = ~\new_[20901]_  | ~\new_[20903]_ ;
  assign \new_[20901]_  = ~\new_[21602]_  | ~\new_[20902]_ ;
  assign \new_[20902]_  = ~\new_[16542]_  & ~\new_[16184]_ ;
  assign \new_[20903]_  = \new_[1089]_ ;
  assign \new_[20904]_  = ~\new_[20905]_ ;
  assign \new_[20905]_  = ~\new_[18974]_  & ~\new_[17249]_ ;
  assign \new_[20906]_  = ~\new_[20907]_ ;
  assign \new_[20907]_  = ~\new_[20746]_  & ~\new_[20747]_ ;
  assign \new_[20908]_  = ~\new_[20911]_  | ~\new_[20910]_  | ~\new_[20909]_ ;
  assign \new_[20909]_  = ~\new_[19736]_  | (~\new_[19825]_  & ~\new_[19827]_ );
  assign \new_[20910]_  = ~\new_[20379]_  & ~\new_[20380]_ ;
  assign \new_[20911]_  = ~\new_[926]_  | (~\new_[20912]_  & ~\new_[20913]_ );
  assign \new_[20912]_  = ~\new_[5193]_  | ~\new_[5061]_ ;
  assign \new_[20913]_  = ~\new_[6265]_  | ~\new_[8804]_ ;
  assign \new_[20914]_  = ~\new_[20917]_  | ~\new_[20915]_  | ~\new_[20916]_ ;
  assign \new_[20915]_  = ~\new_[20970]_  | (~\new_[5632]_  & ~\new_[9165]_ );
  assign \new_[20916]_  = ~\new_[7037]_  & ~\new_[7578]_ ;
  assign \new_[20917]_  = \new_[20918]_  & \new_[7239]_ ;
  assign \new_[20918]_  = ~\new_[20919]_  & (~\new_[19072]_  | ~\new_[10599]_ );
  assign \new_[20919]_  = ~\new_[12656]_  | ~\new_[20920]_ ;
  assign \new_[20920]_  = ~\new_[20921]_ ;
  assign \new_[20921]_  = ~\new_[17786]_  & ~\new_[17998]_ ;
  assign \new_[20922]_  = ~\new_[20929]_  | ~\new_[20926]_  | ~\new_[20923]_  | ~\new_[20924]_ ;
  assign \new_[20923]_  = ~\new_[19321]_  | ~\new_[19096]_ ;
  assign \new_[20924]_  = ~\new_[20925]_ ;
  assign \new_[20925]_  = ~\new_[19096]_  & ~\new_[18493]_ ;
  assign \new_[20926]_  = ~\new_[18454]_  | ~\new_[20927]_ ;
  assign \new_[20927]_  = ~\new_[20928]_ ;
  assign \new_[20928]_  = \new_[955]_ ;
  assign \new_[20929]_  = ~\new_[20930]_  | ~\new_[20928]_ ;
  assign \new_[20930]_  = ~\new_[20931]_ ;
  assign \new_[20931]_  = ~\new_[20932]_ ;
  assign \new_[20932]_  = ~\new_[20933]_ ;
  assign \new_[20933]_  = ~\new_[19584]_  | ~\new_[19313]_ ;
  assign \new_[20934]_  = ~\new_[973]_  | (~\new_[20935]_  & ~\new_[20936]_ );
  assign \new_[20935]_  = ~\new_[18569]_  & (~\new_[12276]_  | ~\new_[10135]_ );
  assign \new_[20936]_  = ~\new_[20937]_  | ~\new_[20940]_  | ~\new_[20938]_ ;
  assign \new_[20937]_  = ~\new_[13446]_  | ~\new_[19260]_ ;
  assign \new_[20938]_  = ~\new_[20939]_ ;
  assign \new_[20939]_  = ~\new_[18978]_  & ~\new_[16789]_ ;
  assign \new_[20940]_  = \new_[19152]_  | \new_[13962]_ ;
  assign \new_[20941]_  = ~\new_[973]_ ;
  assign \new_[20942]_  = ~\new_[20940]_ ;
  assign \new_[20943]_  = ~\new_[20951]_  | ~\new_[20944]_  | ~\new_[20945]_ ;
  assign \new_[20944]_  = ~\new_[3982]_  | ~\new_[949]_ ;
  assign \new_[20945]_  = ~\new_[20950]_  | (~\new_[20946]_  & ~\new_[20948]_ );
  assign \new_[20946]_  = ~\new_[5445]_  | ~\new_[4369]_  | ~\new_[20947]_ ;
  assign \new_[20947]_  = \new_[5723]_  & \new_[8710]_ ;
  assign \new_[20948]_  = ~\new_[4861]_  | ~\new_[20949]_ ;
  assign \new_[20949]_  = \new_[8359]_  & \new_[9437]_ ;
  assign \new_[20950]_  = ~\new_[949]_ ;
  assign \new_[20951]_  = ~\new_[3988]_ ;
  assign \new_[20952]_  = ~\new_[20959]_  | ~\new_[20958]_  | ~\new_[20953]_  | ~\new_[20957]_ ;
  assign \new_[20953]_  = ~\new_[940]_  | (~\new_[20954]_  & ~\new_[20955]_ );
  assign \new_[20954]_  = ~\new_[4452]_  | ~\new_[4993]_ ;
  assign \new_[20955]_  = ~\new_[20956]_  | ~\new_[14627]_ ;
  assign \new_[20956]_  = ~\new_[6353]_  & ~\new_[6623]_ ;
  assign \new_[20957]_  = ~\new_[4235]_  | ~\new_[21008]_ ;
  assign \new_[20958]_  = ~\new_[19640]_  | (~\new_[4308]_  & ~\new_[12782]_ );
  assign \new_[20959]_  = ~\new_[20960]_ ;
  assign \new_[20960]_  = ~\new_[7392]_  | ~\new_[5141]_  | ~\new_[5079]_  | ~\new_[6476]_ ;
  assign \new_[20961]_  = ~\new_[20962]_  | ~\new_[954]_ ;
  assign \new_[20962]_  = ~\new_[20963]_  | ~\new_[20968]_ ;
  assign \new_[20963]_  = ~\new_[20964]_  & ~\new_[20965]_ ;
  assign \new_[20964]_  = ~\new_[19687]_  & (~\new_[13296]_  | ~\new_[15568]_ );
  assign \new_[20965]_  = ~\new_[20966]_  | ~\new_[16218]_  | ~\new_[11579]_ ;
  assign \new_[20966]_  = ~\new_[20967]_ ;
  assign \new_[20967]_  = ~\new_[19409]_  & ~\new_[16773]_ ;
  assign \new_[20968]_  = \new_[20969]_  & \new_[20971]_ ;
  assign \new_[20969]_  = ~\new_[15388]_  | ~\new_[19436]_ ;
  assign \new_[20970]_  = ~\new_[954]_ ;
  assign \new_[20971]_  = ~\new_[21043]_ ;
  assign \new_[20972]_  = \new_[20973]_  ^ \new_[20977]_ ;
  assign \new_[20973]_  = ~\new_[20974]_ ;
  assign \new_[20974]_  = ~\new_[20975]_  | ~\new_[20976]_ ;
  assign \new_[20975]_  = ~\new_[19978]_  | ~\new_[21614]_ ;
  assign \new_[20976]_  = \new_[19978]_  | \new_[21614]_ ;
  assign \new_[20977]_  = \new_[2969]_  ? \new_[2118]_  : \new_[20978]_ ;
  assign \new_[20978]_  = ~\new_[2969]_ ;
  assign \new_[20979]_  = ~\new_[20988]_  | ~\new_[20980]_  | ~\new_[20983]_ ;
  assign \new_[20980]_  = ~\new_[20981]_  | ~\new_[20982]_ ;
  assign \new_[20981]_  = ~\new_[5529]_  | ~\new_[10536]_ ;
  assign \new_[20982]_  = \new_[1087]_ ;
  assign \new_[20983]_  = ~\new_[20984]_  & (~\new_[7489]_  | ~\new_[17925]_ );
  assign \new_[20984]_  = ~\new_[20985]_  | ~\new_[20986]_ ;
  assign \new_[20985]_  = ~\new_[9344]_  & (~\new_[12554]_  | ~\new_[19529]_ );
  assign \new_[20986]_  = ~\new_[6792]_  & (~\new_[20989]_  | ~\new_[14951]_ );
  assign \new_[20987]_  = ~\new_[15838]_  | ~\new_[19068]_ ;
  assign \new_[20988]_  = (~\new_[18895]_  | ~\new_[9248]_ ) & (~\new_[6163]_  | ~\new_[18293]_ );
  assign \new_[20989]_  = ~\new_[20987]_ ;
  assign \new_[20990]_  = ~\new_[4504]_  | ~\new_[5329]_ ;
  assign \new_[20991]_  = ~\new_[20992]_  | ~\new_[4839]_  | ~\new_[6269]_ ;
  assign \new_[20992]_  = ~\new_[12415]_  & ~\new_[9078]_ ;
  assign \new_[20993]_  = \new_[20994]_  ? \new_[21002]_  : \new_[21001]_ ;
  assign \new_[20994]_  = ~\new_[21000]_  | ~\new_[20997]_  | ~\new_[20996]_  | ~\new_[20995]_ ;
  assign \new_[20995]_  = ~\new_[940]_  | (~\new_[4192]_  & ~\new_[4678]_ );
  assign \new_[20996]_  = ~\new_[3900]_ ;
  assign \new_[20997]_  = \new_[4443]_  & \new_[20998]_ ;
  assign \new_[20998]_  = ~\new_[20999]_ ;
  assign \new_[20999]_  = ~\new_[10133]_  | ~\new_[13078]_  | ~\new_[9979]_ ;
  assign \new_[21000]_  = ~\new_[4700]_ ;
  assign \new_[21001]_  = ~\new_[20994]_ ;
  assign \new_[21002]_  = ~\new_[20247]_  | ~\new_[20243]_  | ~\new_[20244]_ ;
  assign \new_[21003]_  = ~\new_[21004]_  & ~\new_[21005]_ ;
  assign \new_[21004]_  = ~\new_[20995]_ ;
  assign \new_[21005]_  = ~\new_[21000]_  | ~\new_[20996]_  | ~\new_[20997]_ ;
  assign \new_[21006]_  = ~\new_[21016]_  | ~\new_[21015]_  | ~\new_[21007]_  | ~\new_[21014]_ ;
  assign \new_[21007]_  = ~\new_[21008]_  | ~\new_[21009]_ ;
  assign \new_[21008]_  = ~\new_[940]_ ;
  assign \new_[21009]_  = ~\new_[4776]_  | ~\new_[4425]_  | ~\new_[21010]_ ;
  assign \new_[21010]_  = ~\new_[21011]_ ;
  assign \new_[21011]_  = ~\new_[21013]_  | ~\new_[13725]_  | ~\new_[21012]_  | ~\new_[6474]_ ;
  assign \new_[21012]_  = ~\new_[9479]_ ;
  assign \new_[21013]_  = ~\new_[9138]_ ;
  assign \new_[21014]_  = ~\new_[940]_  | (~\new_[4365]_  & ~\new_[4948]_ );
  assign \new_[21015]_  = ~\new_[4537]_ ;
  assign \new_[21016]_  = ~\new_[21017]_  & ~\new_[4184]_ ;
  assign \new_[21017]_  = ~\new_[7355]_  | ~\new_[11311]_ ;
  assign \new_[21018]_  = ~\new_[21025]_  | ~\new_[21024]_  | ~\new_[21019]_  | ~\new_[21023]_ ;
  assign \new_[21019]_  = ~\new_[19236]_  | (~\new_[21020]_  & ~\new_[21022]_ );
  assign \new_[21020]_  = ~\new_[9879]_  | ~\new_[6793]_  | ~\new_[21021]_ ;
  assign \new_[21021]_  = \new_[15496]_  & \new_[14866]_ ;
  assign \new_[21022]_  = ~\new_[9916]_  | ~\new_[9188]_ ;
  assign \new_[21023]_  = ~\new_[19300]_  | (~\new_[5612]_  & ~\new_[9053]_ );
  assign \new_[21024]_  = ~\new_[21631]_  | (~\new_[7663]_  & ~\new_[10562]_ );
  assign \new_[21025]_  = ~\new_[21026]_ ;
  assign \new_[21026]_  = ~\new_[14363]_  & ~\new_[19050]_ ;
  assign \new_[21027]_  = ~\new_[21033]_  | ~\new_[21028]_  | ~\new_[21032]_ ;
  assign \new_[21028]_  = ~\new_[4394]_  & ~\new_[21029]_ ;
  assign \new_[21029]_  = ~\new_[4705]_  | ~\new_[21030]_ ;
  assign \new_[21030]_  = ~\new_[21031]_  & (~\new_[6944]_  | ~\new_[18154]_ );
  assign \new_[21031]_  = ~\new_[5321]_ ;
  assign \new_[21032]_  = ~\new_[3921]_  | ~\new_[20181]_ ;
  assign \new_[21033]_  = ~\new_[21452]_  | ~\new_[21034]_ ;
  assign \new_[21034]_  = ~\new_[21118]_  | ~\new_[4739]_  | ~\new_[21035]_  | ~\new_[4325]_ ;
  assign \new_[21035]_  = ~\new_[21036]_  & ~\new_[21037]_ ;
  assign \new_[21036]_  = ~\new_[6174]_ ;
  assign \new_[21037]_  = ~\new_[17689]_  & (~\new_[6855]_  | ~\new_[11584]_ );
  assign \new_[21038]_  = ~\new_[21039]_  | ~\new_[21040]_ ;
  assign \new_[21039]_  = ~\new_[7148]_  | ~\new_[17381]_ ;
  assign \new_[21040]_  = ~\new_[946]_  | (~\new_[21041]_  & ~\new_[21042]_ );
  assign \new_[21041]_  = ~\new_[9595]_  | ~\new_[12807]_ ;
  assign \new_[21042]_  = ~\new_[16458]_  | ~\new_[13530]_  | ~\new_[14134]_  | ~\new_[11505]_ ;
  assign \new_[21043]_  = ~\new_[21044]_ ;
  assign \new_[21044]_  = \new_[21572]_  | \new_[21045]_ ;
  assign \new_[21045]_  = ~\new_[19541]_  | ~\new_[21046]_  | ~\new_[18952]_ ;
  assign \new_[21046]_  = ~\new_[21047]_ ;
  assign \new_[21047]_  = ~\new_[1038]_ ;
  assign \new_[21048]_  = ~\new_[18952]_  | ~\new_[19541]_ ;
  assign \new_[21049]_  = ~\new_[21046]_ ;
  assign \new_[21050]_  = ~\new_[21058]_  | ~\new_[21051]_  | ~\new_[21057]_ ;
  assign \new_[21051]_  = ~\new_[21052]_  & ~\new_[21053]_ ;
  assign \new_[21052]_  = ~\new_[11656]_  | ~\new_[12185]_ ;
  assign \new_[21053]_  = ~\new_[21056]_  & (~\new_[21054]_  | ~\new_[21055]_ );
  assign \new_[21054]_  = ~\new_[15844]_  | ~\new_[18966]_ ;
  assign \new_[21055]_  = ~\new_[18129]_  | ~\new_[19026]_ ;
  assign \new_[21056]_  = ~\new_[1134]_ ;
  assign \new_[21057]_  = ~\new_[12871]_  | ~\new_[19079]_ ;
  assign \new_[21058]_  = ~\new_[21059]_ ;
  assign \new_[21059]_  = ~\new_[17469]_  & ~\new_[13893]_ ;
  assign \new_[21060]_  = ~\new_[17469]_  & ~\new_[13893]_ ;
  assign \new_[21061]_  = ~\new_[21055]_ ;
  assign \new_[21062]_  = ~\new_[21066]_  | (~\new_[21063]_  & ~\new_[21065]_ );
  assign \new_[21063]_  = ~\new_[21064]_  | ~\new_[4714]_ ;
  assign \new_[21064]_  = \new_[5989]_  & \new_[13723]_ ;
  assign \new_[21065]_  = ~\new_[20066]_  | ~\new_[4564]_  | ~\new_[7501]_ ;
  assign \new_[21066]_  = ~\new_[926]_ ;
  assign \new_[21067]_  = ~\new_[19916]_  | ~\new_[4290]_ ;
  assign \new_[21068]_  = ~\new_[20990]_  & ~\new_[20991]_ ;
  assign \new_[21069]_  = ~\new_[4213]_  | ~\new_[4789]_ ;
  assign \new_[21070]_  = ~\new_[19862]_  | ~\new_[19863]_ ;
  assign \new_[21071]_  = ~\new_[950]_ ;
  assign \new_[21072]_  = ~\new_[4552]_ ;
  assign \new_[21073]_  = ~\new_[21074]_ ;
  assign \new_[21074]_  = ~\new_[21075]_  | ~\new_[21509]_ ;
  assign \new_[21075]_  = ~\new_[21076]_ ;
  assign \new_[21076]_  = ~\new_[21077]_  | ~\new_[21078]_ ;
  assign \new_[21077]_  = \new_[21578]_  & \new_[20035]_ ;
  assign \new_[21078]_  = \new_[985]_ ;
  assign \new_[21079]_  = ~\new_[21082]_  | ~\new_[21080]_ ;
  assign \new_[21080]_  = ~\new_[21081]_  & (~\new_[11249]_  | ~\new_[19241]_ );
  assign \new_[21081]_  = \new_[13981]_  & \new_[19241]_ ;
  assign \new_[21082]_  = ~\new_[21083]_  | ~\new_[21142]_ ;
  assign \new_[21083]_  = ~\new_[12937]_  | ~\new_[12926]_ ;
  assign \new_[21084]_  = ~\new_[21081]_ ;
  assign \new_[21085]_  = ~\new_[21089]_  | ~\new_[21088]_  | ~\new_[21086]_  | ~\new_[21087]_ ;
  assign \new_[21086]_  = ~\new_[20283]_  | ~\new_[4239]_ ;
  assign \new_[21087]_  = ~\new_[949]_  | (~\new_[4105]_  & ~\new_[4877]_ );
  assign \new_[21088]_  = ~\new_[19659]_  | (~\new_[4310]_  & ~\new_[12733]_ );
  assign \new_[21089]_  = ~\new_[21090]_ ;
  assign \new_[21090]_  = ~\new_[21093]_  | ~\new_[9508]_  | ~\new_[21091]_  | ~\new_[21092]_ ;
  assign \new_[21091]_  = ~\new_[5350]_  | ~\new_[18091]_ ;
  assign \new_[21092]_  = (~\new_[18786]_  | ~\new_[10068]_ ) & (~\new_[6930]_  | ~\new_[19005]_ );
  assign \new_[21093]_  = ~\new_[11717]_  | ~\new_[18091]_  | ~\new_[17845]_ ;
  assign \new_[21094]_  = ~\new_[21095]_ ;
  assign \new_[21095]_  = \new_[19624]_  | \new_[21096]_ ;
  assign \new_[21096]_  = ~\new_[19329]_  | ~\new_[19644]_  | ~\new_[21097]_ ;
  assign \new_[21097]_  = \new_[997]_ ;
  assign \new_[21098]_  = ~\new_[21099]_ ;
  assign \new_[21099]_  = ~\new_[19329]_  | ~\new_[19644]_ ;
  assign \new_[21100]_  = ~\new_[21097]_ ;
  assign \new_[21101]_  = ~\new_[21102]_  & ~\new_[21105]_ ;
  assign \new_[21102]_  = ~\new_[21103]_  | ~\new_[21104]_ ;
  assign \new_[21103]_  = ~\new_[4078]_  | ~\new_[21180]_ ;
  assign \new_[21104]_  = ~\new_[19623]_  | (~\new_[4916]_  & ~\new_[6611]_ );
  assign \new_[21105]_  = ~\new_[21106]_  | ~\new_[21107]_ ;
  assign \new_[21106]_  = ~\new_[986]_  | ~\new_[3814]_ ;
  assign \new_[21107]_  = ~\new_[21108]_  | ~\new_[18983]_ ;
  assign \new_[21108]_  = ~\new_[5318]_  | ~\new_[20084]_ ;
  assign \new_[21109]_  = ~\new_[21117]_  | ~\new_[21110]_  | ~\new_[21116]_ ;
  assign \new_[21110]_  = ~\new_[21111]_  | ~\new_[21114]_ ;
  assign \new_[21111]_  = ~\new_[6887]_  | ~\new_[21113]_ ;
  assign \new_[21112]_  = ~\new_[10627]_  | ~\new_[12526]_ ;
  assign \new_[21113]_  = ~\new_[17941]_  | ~\new_[19042]_ ;
  assign \new_[21114]_  = \new_[21115]_ ;
  assign \new_[21115]_  = ~\new_[1084]_ ;
  assign \new_[21116]_  = \new_[21114]_  | \new_[12367]_ ;
  assign \new_[21117]_  = \new_[21118]_  & \new_[21119]_ ;
  assign \new_[21118]_  = ~\new_[15209]_  | ~\new_[17922]_ ;
  assign \new_[21119]_  = ~\new_[21120]_ ;
  assign \new_[21120]_  = \new_[13247]_  & \new_[21115]_ ;
  assign \new_[21121]_  = ~\new_[21122]_  | ~\new_[21125]_ ;
  assign \new_[21122]_  = ~\new_[21123]_  & ~\new_[21124]_ ;
  assign \new_[21123]_  = ~\new_[3948]_ ;
  assign \new_[21124]_  = ~\new_[20950]_  & ~\new_[3809]_ ;
  assign \new_[21125]_  = ~\new_[21126]_  & (~\new_[4336]_  | ~\new_[19659]_ );
  assign \new_[21126]_  = ~\new_[21128]_  | (~\new_[21127]_  & ~\new_[19659]_ );
  assign \new_[21127]_  = \new_[5697]_  & \new_[10590]_ ;
  assign \new_[21128]_  = \new_[13604]_  ? \new_[18650]_  : \new_[12499]_ ;
  assign \new_[21129]_  = \new_[21130]_  | \new_[21131]_ ;
  assign \new_[21130]_  = ~\new_[19128]_  & ~\new_[14815]_ ;
  assign \new_[21131]_  = ~\new_[21132]_  | ~\new_[21133]_ ;
  assign \new_[21132]_  = ~\new_[17094]_  | ~\new_[19268]_ ;
  assign \new_[21133]_  = ~\new_[21134]_  & ~\new_[21137]_ ;
  assign \new_[21134]_  = ~\new_[21135]_  | ~\new_[21136]_ ;
  assign \new_[21135]_  = \new_[20764]_  | \new_[20768]_ ;
  assign \new_[21136]_  = \new_[19568]_  | \new_[17706]_ ;
  assign \new_[21137]_  = ~\new_[18709]_  & ~\new_[16896]_ ;
  assign \new_[21138]_  = ~\new_[21135]_ ;
  assign \new_[21139]_  = ~\new_[21140]_  | ~\new_[21143]_ ;
  assign \new_[21140]_  = ~\new_[19022]_  | ~\new_[19912]_  | ~\new_[21141]_  | ~\new_[19910]_ ;
  assign \new_[21141]_  = \new_[10997]_  & \new_[13644]_ ;
  assign \new_[21142]_  = ~\new_[946]_ ;
  assign \new_[21143]_  = ~\new_[21142]_  | ~\new_[13097]_  | ~\new_[21144]_  | ~\new_[21146]_ ;
  assign \new_[21144]_  = ~\new_[14318]_  & ~\new_[21145]_ ;
  assign \new_[21145]_  = ~\new_[13744]_  | ~\new_[14417]_ ;
  assign \new_[21146]_  = ~\new_[12724]_  | ~\new_[16785]_ ;
  assign \new_[21147]_  = ~\new_[3942]_  | ~\new_[21152]_  | ~\new_[21148]_  | ~\new_[21151]_ ;
  assign \new_[21148]_  = ~\new_[937]_  | (~\new_[21149]_  & ~\new_[21150]_ );
  assign \new_[21149]_  = ~\new_[4458]_  | ~\new_[20470]_ ;
  assign \new_[21150]_  = ~\new_[5006]_  | ~\new_[20471]_ ;
  assign \new_[21151]_  = ~\new_[19054]_  | (~\new_[4317]_  & ~\new_[12707]_ );
  assign \new_[21152]_  = ~\new_[21153]_ ;
  assign \new_[21153]_  = ~\new_[6787]_  | ~\new_[20473]_  | ~\new_[5177]_ ;
  assign \new_[21154]_  = ~\new_[21155]_  | ~\new_[21157]_ ;
  assign \new_[21155]_  = ~\new_[21156]_  | (~\new_[3954]_  & ~\new_[1517]_ );
  assign \new_[21156]_  = \new_[19661]_  | \new_[3864]_ ;
  assign \new_[21157]_  = ~\new_[4025]_  & ~\new_[21158]_ ;
  assign \new_[21158]_  = ~\new_[21159]_ ;
  assign \new_[21159]_  = ~\new_[7311]_  & (~\new_[21160]_  | ~\new_[2500]_ );
  assign \new_[21160]_  = ~\new_[4846]_  | ~\new_[4670]_ ;
  assign \new_[21161]_  = ~\new_[21162]_  | ~\new_[21167]_ ;
  assign \new_[21162]_  = (~\new_[14951]_  | ~\new_[16267]_ ) & (~\new_[21163]_  | ~\new_[18973]_ );
  assign \new_[21163]_  = ~\new_[21164]_ ;
  assign \new_[21164]_  = ~\new_[19097]_  | ~\new_[16140]_ ;
  assign \new_[21165]_  = ~\new_[21166]_ ;
  assign \new_[21166]_  = ~\new_[1000]_ ;
  assign \new_[21167]_  = ~\new_[18385]_  | ~\new_[18927]_ ;
  assign \new_[21168]_  = ~\new_[21165]_ ;
  assign \new_[21169]_  = ~\new_[21170]_ ;
  assign \new_[21170]_  = ~\new_[9949]_  | ~\new_[21174]_  | ~\new_[21171]_  | ~\new_[21172]_ ;
  assign \new_[21171]_  = ~\new_[10738]_  | ~\new_[19145]_ ;
  assign \new_[21172]_  = \new_[14150]_  & \new_[21173]_ ;
  assign \new_[21173]_  = ~\new_[14439]_  | ~\new_[18807]_ ;
  assign \new_[21174]_  = ~\new_[21175]_ ;
  assign \new_[21175]_  = ~\new_[19249]_  & (~\new_[12928]_  | ~\new_[16185]_ );
  assign \new_[21176]_  = \new_[21177]_ ;
  assign \new_[21177]_  = ~\new_[21178]_  | ~\new_[21182]_ ;
  assign \new_[21178]_  = ~\new_[21181]_  & (~\new_[21179]_  | ~\new_[21180]_ );
  assign \new_[21179]_  = ~\new_[5927]_  | ~\new_[5651]_  | ~\new_[4485]_  | ~\new_[5956]_ ;
  assign \new_[21180]_  = ~\new_[986]_ ;
  assign \new_[21181]_  = ~\new_[21180]_  & (~\new_[4109]_  | ~\new_[4299]_ );
  assign \new_[21182]_  = ~\new_[21183]_  & ~\new_[21184]_ ;
  assign \new_[21183]_  = ~\new_[5037]_  | ~\new_[8512]_ ;
  assign \new_[21184]_  = ~\new_[6261]_  | ~\new_[21185]_  | ~\new_[4372]_  | ~\new_[6025]_ ;
  assign \new_[21185]_  = ~\new_[21186]_  & (~\new_[10546]_  | ~\new_[19102]_ );
  assign \new_[21186]_  = ~\new_[8572]_ ;
  assign \new_[21187]_  = ~\new_[21192]_  | ~\new_[21188]_  | ~\new_[21190]_ ;
  assign \new_[21188]_  = ~\new_[21189]_  & ~\new_[3830]_ ;
  assign \new_[21189]_  = ~\new_[20725]_  & (~\new_[6077]_  | ~\new_[14016]_ );
  assign \new_[21190]_  = ~\new_[21191]_ ;
  assign \new_[21191]_  = ~\new_[1004]_  & (~\new_[4398]_  | ~\new_[4532]_ );
  assign \new_[21192]_  = ~\new_[21193]_  & ~\new_[3999]_ ;
  assign \new_[21193]_  = ~\new_[21194]_  | (~\new_[9489]_  & ~\new_[19032]_ );
  assign \new_[21194]_  = \new_[21195]_  & \new_[21196]_ ;
  assign \new_[21195]_  = ~\new_[15461]_  | ~\new_[16998]_ ;
  assign \new_[21196]_  = ~\new_[17373]_  | ~\new_[11705]_ ;
  assign \new_[21197]_  = ~\new_[21195]_ ;
  assign \new_[21198]_  = ~\new_[4462]_  | ~\new_[21202]_  | ~\new_[3791]_  | ~\new_[21199]_ ;
  assign \new_[21199]_  = ~\new_[21200]_ ;
  assign \new_[21200]_  = ~\new_[21201]_  | ~\new_[4495]_  | ~\new_[12741]_ ;
  assign \new_[21201]_  = \new_[18609]_  | \new_[17155]_  | \new_[18683]_  | \new_[18542]_ ;
  assign \new_[21202]_  = ~\new_[21203]_  | ~\new_[19564]_ ;
  assign \new_[21203]_  = ~\new_[10415]_  | ~\new_[5668]_  | ~\new_[4995]_  | ~\new_[5546]_ ;
  assign \new_[21204]_  = ~\new_[8298]_  | ~\new_[5752]_  | ~\new_[5682]_ ;
  assign \new_[21205]_  = ~\new_[994]_ ;
  assign \new_[21206]_  = ~\new_[21208]_  | ~\new_[21294]_  | ~\new_[21207]_ ;
  assign \new_[21207]_  = ~\new_[19236]_  | (~\new_[6428]_  & ~\new_[15270]_ );
  assign \new_[21208]_  = \new_[18416]_  | \new_[21209]_ ;
  assign \new_[21209]_  = ~\new_[14312]_  & ~\new_[8559]_ ;
  assign \new_[21210]_  = ~\new_[21216]_  | ~\new_[21215]_  | ~\new_[21211]_  | ~\new_[21212]_ ;
  assign \new_[21211]_  = ~\new_[21071]_  | (~\new_[21069]_  & ~\new_[21070]_ );
  assign \new_[21212]_  = \new_[21072]_  & \new_[21213]_ ;
  assign \new_[21213]_  = ~\new_[21214]_  | ~\new_[19599]_ ;
  assign \new_[21214]_  = ~\new_[4999]_ ;
  assign \new_[21215]_  = ~\new_[950]_  | (~\new_[4366]_  & ~\new_[4949]_ );
  assign \new_[21216]_  = ~\new_[21217]_  & ~\new_[19864]_ ;
  assign \new_[21217]_  = ~\new_[6562]_ ;
  assign \new_[21218]_  = ~\new_[21219]_  | ~\new_[21225]_ ;
  assign \new_[21219]_  = ~\new_[21220]_  & ~\new_[21222]_ ;
  assign \new_[21220]_  = ~\new_[7235]_  | ~\new_[21221]_ ;
  assign \new_[21221]_  = \new_[14344]_  & \new_[16663]_ ;
  assign \new_[21222]_  = ~\new_[1033]_  & (~\new_[21224]_  | ~\new_[21223]_ );
  assign \new_[21223]_  = ~\new_[9097]_ ;
  assign \new_[21224]_  = ~\new_[6145]_ ;
  assign \new_[21225]_  = ~\new_[21226]_  & ~\new_[21227]_ ;
  assign \new_[21226]_  = ~\new_[19600]_  & (~\new_[11673]_  | ~\new_[9923]_ );
  assign \new_[21227]_  = ~\new_[21229]_  | (~\new_[21228]_  & ~\new_[18393]_ );
  assign \new_[21228]_  = \new_[12002]_  & \new_[12070]_ ;
  assign \new_[21229]_  = ~\new_[10669]_  | ~\new_[20099]_ ;
  assign \new_[21230]_  = ~\new_[21231]_  & ~\new_[21233]_ ;
  assign \new_[21231]_  = ~\new_[21232]_  | ~\new_[4208]_  | ~\new_[4727]_ ;
  assign \new_[21232]_  = \new_[10476]_  & \new_[9547]_ ;
  assign \new_[21233]_  = ~\new_[21236]_  & (~\new_[21234]_  | ~\new_[21235]_ );
  assign \new_[21234]_  = ~\new_[4467]_ ;
  assign \new_[21235]_  = ~\new_[932]_  & ~\new_[8105]_ ;
  assign \new_[21236]_  = ~\new_[21237]_  & ~\new_[3951]_ ;
  assign \new_[21237]_  = \new_[19786]_  | \new_[6869]_ ;
  assign \new_[21238]_  = \new_[21239]_  ^ \new_[21241]_ ;
  assign \new_[21239]_  = ~\new_[21240]_ ;
  assign \new_[21240]_  = \new_[20112]_  ? \new_[20114]_  : \new_[20113]_ ;
  assign \new_[21241]_  = \new_[21242]_  ? \new_[2543]_  : \new_[3168]_ ;
  assign \new_[21242]_  = ~\new_[3168]_ ;
  assign n1103 = ~\new_[21250]_  | ~\new_[21244]_  | ~\new_[21249]_ ;
  assign \new_[21244]_  = ~\new_[19874]_  | ~\new_[21245]_  | ~\new_[21247]_ ;
  assign \new_[21245]_  = ~\new_[21246]_ ;
  assign \new_[21246]_  = \new_[2989]_  ? \new_[2232]_  : \new_[2988]_ ;
  assign \new_[21247]_  = ~\new_[21248]_ ;
  assign \new_[21248]_  = ~\new_[1966]_  | ~\new_[2159]_ ;
  assign \new_[21249]_  = ~\new_[19874]_  | ~\new_[21246]_  | ~\new_[21248]_ ;
  assign \new_[21250]_  = \new_[15530]_  | \new_[17819]_ ;
  assign \new_[21251]_  = ~\new_[21252]_  & ~\new_[21253]_ ;
  assign \new_[21252]_  = ~\new_[947]_ ;
  assign \new_[21253]_  = ~\new_[21259]_  | ~\new_[21255]_ ;
  assign \new_[21254]_  = \new_[943]_ ;
  assign \new_[21255]_  = ~\new_[21256]_ ;
  assign \new_[21256]_  = ~\new_[19303]_  | ~\new_[18281]_ ;
  assign \new_[21257]_  = ~\new_[21259]_  | ~\new_[21255]_ ;
  assign \new_[21258]_  = ~\new_[21252]_ ;
  assign \new_[21259]_  = ~\new_[21254]_ ;
  assign \new_[21260]_  = ~\new_[21268]_  | ~\new_[21263]_  | ~\new_[21261]_  | ~\new_[21262]_ ;
  assign \new_[21261]_  = ~\new_[994]_  | (~\new_[4005]_  & ~\new_[4898]_ );
  assign \new_[21262]_  = ~\new_[4247]_  | ~\new_[21205]_ ;
  assign \new_[21263]_  = ~\new_[21264]_  | ~\new_[21267]_ ;
  assign \new_[21264]_  = ~\new_[21265]_  | ~\new_[21266]_ ;
  assign \new_[21265]_  = ~\new_[5801]_ ;
  assign \new_[21266]_  = ~\new_[7276]_  & ~\new_[12534]_  & ~\new_[12044]_ ;
  assign \new_[21267]_  = ~\new_[991]_ ;
  assign \new_[21268]_  = ~\new_[21269]_  & ~\new_[4856]_ ;
  assign \new_[21269]_  = ~\new_[21270]_  | ~\new_[21271]_ ;
  assign \new_[21270]_  = ~\new_[6569]_ ;
  assign \new_[21271]_  = ~\new_[8505]_  & (~\new_[21272]_  | ~\new_[21273]_ );
  assign \new_[21272]_  = ~\new_[17358]_  & ~\new_[21661]_ ;
  assign \new_[21273]_  = ~\new_[19236]_  & ~\new_[21628]_ ;
  assign \new_[21274]_  = ~\new_[21273]_ ;
  assign \new_[21275]_  = ~\new_[21276]_  | ~\new_[21284]_ ;
  assign \new_[21276]_  = ~\new_[21277]_ ;
  assign \new_[21277]_  = \new_[21278]_ ;
  assign \new_[21278]_  = ~\new_[21283]_  | ~\new_[21281]_  | ~\new_[21279]_  | ~\new_[21280]_ ;
  assign \new_[21279]_  = ~\new_[21206]_  & (~\new_[21204]_  | ~\new_[21205]_ );
  assign \new_[21280]_  = ~\new_[19304]_  | ~\new_[21309]_ ;
  assign \new_[21281]_  = ~\new_[20330]_  | ~\new_[21282]_ ;
  assign \new_[21282]_  = \new_[991]_  & \new_[21205]_ ;
  assign \new_[21283]_  = ~\new_[991]_  | (~\new_[5532]_  & ~\new_[5588]_ );
  assign \new_[21284]_  = ~\new_[21285]_ ;
  assign \new_[21285]_  = ~\new_[21286]_ ;
  assign \new_[21286]_  = ~\new_[20016]_  | ~\new_[20500]_  | ~\new_[20015]_ ;
  assign \new_[21287]_  = ~\new_[21288]_  | ~\new_[20616]_  | ~\new_[20615]_  | ~\new_[20617]_ ;
  assign \new_[21288]_  = ~\new_[21289]_  & ~\new_[21290]_ ;
  assign \new_[21289]_  = ~\new_[18875]_  & ~\new_[13715]_ ;
  assign \new_[21290]_  = ~\new_[18798]_  & ~\new_[9227]_ ;
  assign \new_[21291]_  = ~\new_[21292]_  | ~\new_[21293]_ ;
  assign \new_[21292]_  = ~\new_[4245]_  | ~\new_[19816]_ ;
  assign \new_[21293]_  = ~\new_[3968]_  | ~\new_[979]_ ;
  assign \new_[21294]_  = \new_[21630]_  | \new_[21295]_ ;
  assign \new_[21295]_  = \new_[21296]_  & \new_[21297]_ ;
  assign \new_[21296]_  = ~\new_[18126]_  | ~\new_[13271]_ ;
  assign \new_[21297]_  = \new_[14926]_  | \new_[18126]_ ;
  assign \new_[21298]_  = ~\new_[18126]_  | ~\new_[13271]_ ;
  assign \new_[21299]_  = ~\new_[21298]_ ;
  assign \new_[21300]_  = ~\new_[21301]_  | ~\new_[21306]_ ;
  assign \new_[21301]_  = ~\new_[21302]_ ;
  assign \new_[21302]_  = ~\new_[21655]_  | ~\new_[18327]_ ;
  assign \new_[21303]_  = ~\new_[21304]_ ;
  assign \new_[21304]_  = ~\new_[21305]_ ;
  assign \new_[21305]_  = ~\new_[941]_ ;
  assign \new_[21306]_  = ~\new_[21307]_ ;
  assign \new_[21307]_  = \new_[927]_ ;
  assign \new_[21308]_  = ~\new_[21536]_  & ~\new_[19678]_ ;
  assign \new_[21309]_  = ~\new_[21314]_  | ~\new_[21310]_  | ~\new_[21313]_ ;
  assign \new_[21310]_  = \new_[21311]_  & \new_[21312]_ ;
  assign \new_[21311]_  = ~\new_[8703]_  | ~\new_[991]_ ;
  assign \new_[21312]_  = ~\new_[21638]_  | ~\new_[10703]_ ;
  assign \new_[21313]_  = ~\new_[19236]_  | (~\new_[20517]_  & ~\new_[9102]_ );
  assign \new_[21314]_  = ~\new_[21315]_  & ~\new_[21317]_ ;
  assign \new_[21315]_  = ~\new_[7236]_  | ~\new_[21316]_ ;
  assign \new_[21316]_  = ~\new_[17909]_  | ~\new_[21653]_ ;
  assign \new_[21317]_  = ~\new_[13219]_  | ~\new_[21318]_ ;
  assign \new_[21318]_  = ~\new_[20922]_  | ~\new_[21273]_ ;
  assign \new_[21319]_  = ~\new_[21320]_  | ~\new_[21323]_ ;
  assign \new_[21320]_  = \new_[21321]_  & \new_[21322]_ ;
  assign \new_[21321]_  = ~\new_[17093]_  | ~\new_[18542]_ ;
  assign \new_[21322]_  = ~\new_[14483]_  | ~\new_[19233]_ ;
  assign \new_[21323]_  = ~\new_[21324]_  & ~\new_[21327]_ ;
  assign \new_[21324]_  = ~\new_[21325]_  & ~\new_[21326]_ ;
  assign \new_[21325]_  = \new_[1005]_ ;
  assign \new_[21326]_  = ~\new_[18375]_  | ~\new_[19136]_ ;
  assign \new_[21327]_  = ~\new_[21328]_  & ~\new_[16639]_ ;
  assign \new_[21328]_  = ~\new_[21325]_ ;
  assign \new_[21329]_  = ~\new_[21324]_ ;
  assign \new_[21330]_  = ~\new_[19233]_  | ~\new_[14483]_ ;
  assign \new_[21331]_  = ~\new_[21326]_ ;
  assign \new_[21332]_  = ~\new_[4086]_  | ~\new_[21335]_  | ~\new_[21333]_  | ~\new_[3796]_ ;
  assign \new_[21333]_  = ~\new_[21334]_  & (~\new_[4296]_  | ~\new_[19257]_ );
  assign \new_[21334]_  = ~\new_[6646]_  | ~\new_[10618]_ ;
  assign \new_[21335]_  = ~\new_[986]_  | ~\new_[21336]_ ;
  assign \new_[21336]_  = ~\new_[6283]_  | ~\new_[21338]_  | ~\new_[5939]_  | ~\new_[21337]_ ;
  assign \new_[21337]_  = ~\new_[5779]_  | ~\new_[18983]_ ;
  assign \new_[21338]_  = ~\new_[19623]_  | ~\new_[7134]_ ;
  assign \new_[21339]_  = ~\new_[21340]_  & ~\new_[21343]_ ;
  assign \new_[21340]_  = \new_[21341]_  & \new_[21342]_ ;
  assign \new_[21341]_  = ~\new_[21498]_  & ~\new_[17311]_ ;
  assign \new_[21342]_  = \new_[16879]_  & \new_[21142]_ ;
  assign \new_[21343]_  = ~\new_[19599]_  & (~\new_[21345]_  | ~\new_[21344]_ );
  assign \new_[21344]_  = ~\new_[7676]_  | ~\new_[18037]_ ;
  assign \new_[21345]_  = ~\new_[21346]_  & (~\new_[11378]_  | ~\new_[16879]_ );
  assign \new_[21346]_  = ~\new_[13530]_  & ~\new_[20704]_ ;
  assign \new_[21347]_  = ~\new_[21341]_ ;
  assign \new_[21348]_  = ~\new_[11378]_  | ~\new_[16879]_ ;
  assign \new_[21349]_  = ~\new_[21346]_ ;
  assign \new_[21350]_  = ~\new_[21356]_  | ~\new_[21351]_  | ~\new_[21352]_ ;
  assign \new_[21351]_  = ~\new_[19564]_  | (~\new_[4535]_  & ~\new_[4661]_ );
  assign \new_[21352]_  = ~\new_[21353]_  & ~\new_[21354]_ ;
  assign \new_[21353]_  = ~\new_[4926]_  | ~\new_[5190]_ ;
  assign \new_[21354]_  = ~\new_[21355]_  | ~\new_[4925]_ ;
  assign \new_[21355]_  = \new_[6750]_  & \new_[7298]_ ;
  assign \new_[21356]_  = ~\new_[20727]_  | ~\new_[935]_ ;
  assign \new_[21357]_  = ~\new_[21365]_  | ~\new_[21364]_  | ~\new_[21358]_  | ~\new_[21362]_ ;
  assign \new_[21358]_  = ~\new_[21359]_  & (~\new_[9242]_  | ~\new_[19170]_ );
  assign \new_[21359]_  = ~\new_[21360]_  | ~\new_[21361]_ ;
  assign \new_[21360]_  = ~\new_[10187]_  | ~\new_[19170]_ ;
  assign \new_[21361]_  = ~\new_[938]_  & (~\new_[8952]_  | ~\new_[18818]_ );
  assign \new_[21362]_  = ~\new_[21363]_ ;
  assign \new_[21363]_  = ~\new_[19619]_  & (~\new_[8451]_  | ~\new_[6575]_ );
  assign \new_[21364]_  = ~\new_[8453]_  & ~\new_[6499]_ ;
  assign \new_[21365]_  = ~\new_[18818]_  | ~\new_[12562]_ ;
  assign \new_[21366]_  = \new_[21367]_  ? \new_[21369]_  : \new_[21368]_ ;
  assign \new_[21367]_  = ~\new_[21368]_ ;
  assign \new_[21368]_  = ~\new_[3185]_  | ~\new_[2966]_ ;
  assign \new_[21369]_  = \new_[20053]_  ? \new_[2845]_  : \new_[3624]_ ;
  assign \new_[21370]_  = \new_[21371]_  ^ \new_[21374]_ ;
  assign \new_[21371]_  = ~\new_[21372]_  | ~\new_[21373]_ ;
  assign \new_[21372]_  = ~\new_[3911]_  & (~\new_[4229]_  | ~\new_[938]_ );
  assign \new_[21373]_  = ~\new_[5444]_  & ~\new_[3913]_ ;
  assign \new_[21374]_  = ~\new_[3834]_  | ~\new_[3749]_ ;
  assign \new_[21375]_  = ~\new_[21372]_  | ~\new_[21373]_ ;
  assign \new_[21376]_  = ~\new_[3749]_  | ~\new_[3834]_ ;
  assign \new_[21377]_  = ~\new_[21385]_  & (~\new_[21378]_  | ~\new_[21380]_ );
  assign \new_[21378]_  = ~\new_[21379]_  & (~\new_[21050]_  | ~\new_[18649]_ );
  assign \new_[21379]_  = \new_[20763]_  & \new_[6579]_ ;
  assign \new_[21380]_  = ~\new_[21381]_  & ~\new_[21384]_ ;
  assign \new_[21381]_  = \new_[21382]_  | \new_[21383]_ ;
  assign \new_[21382]_  = ~\new_[19073]_  & ~\new_[21055]_ ;
  assign \new_[21383]_  = ~\new_[21056]_  & ~\new_[14358]_ ;
  assign \new_[21384]_  = ~\new_[6861]_  | ~\new_[6485]_ ;
  assign \new_[21385]_  = ~\new_[21386]_ ;
  assign \new_[21386]_  = ~\new_[940]_ ;
  assign \new_[21387]_  = ~\new_[21388]_  & ~\new_[21389]_ ;
  assign \new_[21388]_  = ~\new_[19664]_  | ~\new_[21559]_ ;
  assign \new_[21389]_  = ~\new_[21390]_ ;
  assign \new_[21390]_  = ~\new_[21391]_ ;
  assign \new_[21391]_  = ~\new_[21392]_  | ~\new_[21394]_ ;
  assign \new_[21392]_  = ~\new_[21393]_ ;
  assign \new_[21393]_  = ~\new_[21493]_  | ~\new_[18457]_ ;
  assign \new_[21394]_  = ~\new_[21395]_ ;
  assign \new_[21395]_  = \new_[924]_ ;
  assign \new_[21396]_  = ~\new_[21395]_ ;
  assign \new_[21397]_  = ~\new_[924]_ ;
  assign \new_[21398]_  = ~\new_[21399]_  & ~\new_[19000]_ ;
  assign \new_[21399]_  = ~\new_[21400]_ ;
  assign \new_[21400]_  = ~\new_[1036]_  & ~\new_[21401]_ ;
  assign \new_[21401]_  = ~\new_[982]_ ;
  assign \new_[21402]_  = \new_[985]_ ;
  assign \new_[21403]_  = ~\new_[1036]_ ;
  assign \new_[21404]_  = ~\new_[21401]_ ;
  assign \new_[21405]_  = ~\new_[21409]_  | ~\new_[21406]_  | ~\new_[21408]_ ;
  assign \new_[21406]_  = ~\new_[21407]_ ;
  assign \new_[21407]_  = ~\new_[18007]_  & ~\new_[18564]_ ;
  assign \new_[21408]_  = ~\new_[17112]_  | ~\new_[18974]_ ;
  assign \new_[21409]_  = ~\new_[21410]_  | ~\new_[1089]_ ;
  assign \new_[21410]_  = ~\new_[21411]_ ;
  assign \new_[21411]_  = ~\new_[18218]_  | ~\new_[19359]_ ;
  assign \new_[21412]_  = ~\new_[21408]_ ;
  assign \new_[21413]_  = ~\new_[1089]_ ;
  assign \new_[21414]_  = ~\new_[937]_  & ~\new_[21415]_ ;
  assign \new_[21415]_  = ~\new_[21419]_  & (~\new_[21416]_  | ~\new_[21417]_ );
  assign \new_[21416]_  = ~\new_[20154]_  | ~\new_[20155]_  | ~\new_[20153]_ ;
  assign \new_[21417]_  = ~\new_[21418]_ ;
  assign \new_[21418]_  = ~\new_[959]_ ;
  assign \new_[21419]_  = ~\new_[7277]_  | ~\new_[21420]_  | ~\new_[21423]_ ;
  assign \new_[21420]_  = ~\new_[21421]_  | ~\new_[21422]_ ;
  assign \new_[21421]_  = ~\new_[10258]_  | ~\new_[8737]_  | ~\new_[7933]_ ;
  assign \new_[21422]_  = ~\new_[959]_ ;
  assign \new_[21423]_  = ~\new_[21424]_ ;
  assign \new_[21424]_  = ~\new_[13232]_  | ~\new_[9937]_  | ~\new_[11285]_ ;
  assign \new_[21425]_  = ~\new_[937]_ ;
  assign \new_[21426]_  = ~\new_[21427]_  & ~\new_[21433]_ ;
  assign \new_[21427]_  = ~\new_[3940]_  | ~\new_[21428]_ ;
  assign \new_[21428]_  = \new_[21429]_  & \new_[21432]_ ;
  assign \new_[21429]_  = ~\new_[21430]_  & ~\new_[20724]_ ;
  assign \new_[21430]_  = ~\new_[21431]_  | (~\new_[10485]_  & ~\new_[18941]_ );
  assign \new_[21431]_  = \new_[17615]_  | \new_[13468]_ ;
  assign \new_[21432]_  = ~\new_[8857]_  | ~\new_[16939]_ ;
  assign \new_[21433]_  = ~\new_[21434]_  | ~\new_[3807]_ ;
  assign \new_[21434]_  = \new_[21435]_  & \new_[21436]_ ;
  assign \new_[21435]_  = ~\new_[19442]_  | (~\new_[5057]_  & ~\new_[11645]_ );
  assign \new_[21436]_  = ~\new_[19271]_  | (~\new_[4309]_  & ~\new_[11706]_ );
  assign \new_[21437]_  = ~\new_[21443]_  | ~\new_[21438]_  | ~\new_[21442]_ ;
  assign \new_[21438]_  = ~\new_[21439]_  | ~\new_[21441]_ ;
  assign \new_[21439]_  = ~\new_[5069]_  | ~\new_[21440]_  | ~\new_[5010]_ ;
  assign \new_[21440]_  = \new_[6049]_  & \new_[6425]_ ;
  assign \new_[21441]_  = ~\new_[938]_ ;
  assign \new_[21442]_  = ~\new_[18409]_  | (~\new_[4188]_  & ~\new_[6313]_ );
  assign \new_[21443]_  = ~\new_[21444]_  | ~\new_[18599]_ ;
  assign \new_[21444]_  = ~\new_[6103]_  | ~\new_[10319]_ ;
  assign \new_[21445]_  = ~\new_[21455]_  | ~\new_[21454]_  | ~\new_[21447]_  | ~\new_[21446]_ ;
  assign \new_[21446]_  = ~\new_[20182]_  | ~\new_[20181]_ ;
  assign \new_[21447]_  = ~\new_[21448]_  | ~\new_[21452]_ ;
  assign \new_[21448]_  = ~\new_[21449]_  | ~\new_[4265]_ ;
  assign \new_[21449]_  = ~\new_[21450]_  & ~\new_[21451]_ ;
  assign \new_[21450]_  = ~\new_[10623]_  | ~\new_[6889]_  | ~\new_[6395]_ ;
  assign \new_[21451]_  = ~\new_[4958]_ ;
  assign \new_[21452]_  = ~\new_[21453]_ ;
  assign \new_[21453]_  = ~\new_[956]_ ;
  assign \new_[21454]_  = ~\new_[19748]_  | (~\new_[4316]_  & ~\new_[12635]_ );
  assign \new_[21455]_  = ~\new_[20183]_  & ~\new_[20184]_ ;
  assign \new_[21456]_  = ~\new_[21460]_  | ~\new_[21457]_  | ~\new_[21458]_ ;
  assign \new_[21457]_  = ~\new_[19490]_  | (~\new_[4613]_  & ~\new_[4936]_ );
  assign \new_[21458]_  = ~\new_[21459]_ ;
  assign \new_[21459]_  = ~\new_[932]_  & (~\new_[4625]_  | ~\new_[5078]_ );
  assign \new_[21460]_  = ~\new_[21461]_  & (~\new_[4618]_  | ~\new_[18406]_ );
  assign \new_[21461]_  = ~\new_[21467]_  | ~\new_[21464]_  | ~\new_[21463]_  | ~\new_[21462]_ ;
  assign \new_[21462]_  = ~\new_[20673]_ ;
  assign \new_[21463]_  = ~\new_[20674]_ ;
  assign \new_[21464]_  = ~\new_[21465]_  & (~\new_[10892]_  | ~\new_[20679]_ );
  assign \new_[21465]_  = ~\new_[21466]_ ;
  assign \new_[21466]_  = ~\new_[17954]_  | ~\new_[15412]_ ;
  assign \new_[21467]_  = ~\new_[21468]_  & ~\new_[21469]_ ;
  assign \new_[21468]_  = ~\new_[17523]_  & ~\new_[16183]_ ;
  assign \new_[21469]_  = ~\new_[21470]_ ;
  assign \new_[21470]_  = ~\new_[17357]_  | ~\new_[12812]_ ;
  assign \new_[21471]_  = ~\new_[21068]_  | ~\new_[21062]_  | ~\new_[21067]_ ;
  assign \new_[21472]_  = ~\new_[21068]_  | ~\new_[21062]_  | ~\new_[21067]_ ;
  assign \new_[21473]_  = ~\new_[4922]_  | ~\new_[3761]_  | ~\new_[3778]_  | ~\new_[4158]_ ;
  assign \new_[21474]_  = ~\new_[4922]_  | ~\new_[3761]_  | ~\new_[3778]_  | ~\new_[4158]_ ;
  assign \new_[21475]_  = ~\new_[21695]_  & ~\new_[12028]_ ;
  assign \new_[21476]_  = ~\new_[21697]_  & ~\new_[12028]_ ;
  assign \new_[21477]_  = ~\new_[19370]_  | ~\new_[19573]_ ;
  assign \new_[21478]_  = ~\new_[19370]_  | ~\new_[19573]_ ;
  assign \new_[21479]_  = \new_[21480]_ ;
  assign \new_[21480]_  = ~\new_[2399]_ ;
  assign \new_[21481]_  = ~\new_[2872]_ ;
  assign \new_[21482]_  = ~\new_[2872]_ ;
  assign \new_[21483]_  = \new_[20299]_ ;
  assign \new_[21484]_  = ~\new_[21488]_ ;
  assign \new_[21485]_  = ~\new_[21488]_ ;
  assign \new_[21486]_  = ~\new_[21487]_ ;
  assign \new_[21487]_  = ~\new_[21488]_ ;
  assign \new_[21488]_  = ~\new_[20101]_ ;
  assign \new_[21489]_  = ~\new_[21494]_ ;
  assign \new_[21490]_  = \new_[21494]_ ;
  assign \new_[21491]_  = ~\new_[21492]_ ;
  assign \new_[21492]_  = \new_[21493]_ ;
  assign \new_[21493]_  = ~\new_[21489]_ ;
  assign \new_[21494]_  = ~\new_[1021]_ ;
  assign \new_[21495]_  = \new_[21513]_ ;
  assign \new_[21496]_  = ~\new_[21497]_ ;
  assign \new_[21497]_  = ~\new_[21513]_ ;
  assign \new_[21498]_  = \new_[21501]_ ;
  assign \new_[21499]_  = \new_[21500]_ ;
  assign \new_[21500]_  = ~\new_[21503]_ ;
  assign \new_[21501]_  = ~\new_[21503]_ ;
  assign \new_[21502]_  = ~\new_[21503]_ ;
  assign \new_[21503]_  = ~\new_[21513]_ ;
  assign \new_[21504]_  = ~\new_[21505]_ ;
  assign \new_[21505]_  = \new_[21513]_ ;
  assign \new_[21506]_  = ~\new_[21512]_ ;
  assign \new_[21507]_  = ~\new_[21512]_ ;
  assign \new_[21508]_  = ~\new_[21509]_ ;
  assign \new_[21509]_  = ~\new_[21511]_ ;
  assign \new_[21510]_  = \new_[21511]_ ;
  assign \new_[21511]_  = ~\new_[21512]_ ;
  assign \new_[21512]_  = ~\new_[21513]_ ;
  assign \new_[21513]_  = ~\new_[928]_ ;
  assign \new_[21514]_  = ~\new_[21515]_ ;
  assign \new_[21515]_  = \new_[21517]_ ;
  assign \new_[21516]_  = ~\new_[21517]_ ;
  assign \new_[21517]_  = ~\new_[990]_ ;
  assign \new_[21518]_  = ~\new_[21523]_ ;
  assign \new_[21519]_  = ~\new_[21520]_ ;
  assign \new_[21520]_  = \new_[21521]_ ;
  assign \new_[21521]_  = ~\new_[21523]_ ;
  assign \new_[21522]_  = ~\new_[21523]_ ;
  assign \new_[21523]_  = ~\new_[21526]_ ;
  assign \new_[21524]_  = ~\new_[21525]_ ;
  assign \new_[21525]_  = \new_[21526]_ ;
  assign \new_[21526]_  = ~\new_[953]_ ;
  assign \new_[21527]_  = \new_[3694]_ ;
  assign \new_[21528]_  = ~\new_[21529]_ ;
  assign \new_[21529]_  = ~\new_[18282]_ ;
  assign \new_[21530]_  = ~\new_[5120]_  | ~\new_[4081]_  | ~\new_[3760]_  | ~\new_[3874]_ ;
  assign \new_[21531]_  = ~\new_[5120]_  | ~\new_[4081]_  | ~\new_[3760]_  | ~\new_[3874]_ ;
  assign \new_[21532]_  = ~\new_[21534]_ ;
  assign \new_[21533]_  = ~\new_[21534]_ ;
  assign \new_[21534]_  = \new_[21536]_ ;
  assign \new_[21535]_  = ~\new_[21536]_ ;
  assign \new_[21536]_  = ~\new_[987]_ ;
  assign \new_[21537]_  = ~\new_[21275]_  | ~\new_[3274]_ ;
  assign \new_[21538]_  = ~\new_[21275]_  | ~\new_[3274]_ ;
  assign \new_[21539]_  = ~\new_[21540]_ ;
  assign \new_[21540]_  = \new_[21545]_ ;
  assign \new_[21541]_  = ~\new_[21542]_ ;
  assign \new_[21542]_  = \new_[21543]_ ;
  assign \new_[21543]_  = ~\new_[21544]_ ;
  assign \new_[21544]_  = ~\new_[21545]_ ;
  assign \new_[21545]_  = ~\new_[1137]_ ;
  assign \new_[21546]_  = ~\new_[21547]_ ;
  assign \new_[21547]_  = ~\new_[12875]_ ;
  assign \new_[21548]_  = ~\new_[21549]_ ;
  assign \new_[21549]_  = ~\new_[16066]_ ;
  assign \new_[21550]_  = ~\new_[16791]_ ;
  assign \new_[21551]_  = ~\new_[21552]_ ;
  assign \new_[21552]_  = \new_[16791]_ ;
  assign \new_[21553]_  = ~\new_[21554]_ ;
  assign \new_[21554]_  = \new_[21555]_ ;
  assign \new_[21555]_  = ~\new_[12847]_ ;
  assign \new_[21556]_  = ~\new_[21559]_ ;
  assign \new_[21557]_  = ~\new_[21559]_ ;
  assign \new_[21558]_  = ~\new_[21559]_ ;
  assign \new_[21559]_  = ~\new_[21563]_ ;
  assign \new_[21560]_  = ~\new_[21559]_ ;
  assign \new_[21561]_  = ~\new_[21562]_ ;
  assign \new_[21562]_  = ~\new_[21559]_ ;
  assign \new_[21563]_  = ~\new_[1028]_ ;
  assign \new_[21564]_  = ~\new_[21565]_ ;
  assign \new_[21565]_  = ~\new_[21566]_ ;
  assign \new_[21566]_  = ~\new_[17627]_ ;
  assign \new_[21567]_  = ~\new_[21569]_ ;
  assign \new_[21568]_  = \new_[21569]_ ;
  assign \new_[21569]_  = \new_[21575]_ ;
  assign \new_[21570]_  = \new_[21575]_ ;
  assign \new_[21571]_  = \new_[21572]_ ;
  assign \new_[21572]_  = ~\new_[1040]_ ;
  assign \new_[21573]_  = ~\new_[21575]_ ;
  assign \new_[21574]_  = ~\new_[21573]_ ;
  assign \new_[21575]_  = ~\new_[1040]_ ;
  assign \new_[21576]_  = \new_[21577]_ ;
  assign \new_[21577]_  = ~\new_[20993]_ ;
  assign \new_[21578]_  = ~\new_[21583]_ ;
  assign \new_[21579]_  = ~\new_[21580]_ ;
  assign \new_[21580]_  = \new_[21581]_ ;
  assign \new_[21581]_  = \new_[21583]_ ;
  assign \new_[21582]_  = \new_[21583]_ ;
  assign \new_[21583]_  = ~\new_[1032]_ ;
  assign \new_[21584]_  = \new_[21585]_ ;
  assign \new_[21585]_  = ~\new_[1032]_ ;
  assign \new_[21586]_  = \new_[21147]_ ;
  assign \new_[21587]_  = ~\new_[21590]_ ;
  assign \new_[21588]_  = ~\new_[21589]_ ;
  assign \new_[21589]_  = \new_[21590]_ ;
  assign \new_[21590]_  = ~\new_[21147]_ ;
  assign \new_[21591]_  = ~\new_[10595]_ ;
  assign \new_[21592]_  = ~\new_[12406]_ ;
  assign \new_[21593]_  = ~\new_[15915]_ ;
  assign \new_[21594]_  = ~\new_[13224]_ ;
  assign \new_[21595]_  = ~\new_[21596]_ ;
  assign \new_[21596]_  = ~\new_[21597]_ ;
  assign \new_[21597]_  = \new_[21426]_ ;
  assign \new_[21598]_  = ~\new_[21599]_ ;
  assign \new_[21599]_  = ~\new_[21426]_ ;
  assign \new_[21600]_  = ~\new_[12970]_ ;
  assign \new_[21601]_  = ~\new_[14268]_ ;
  assign \new_[21602]_  = \new_[20749]_  | \new_[16604]_ ;
  assign \new_[21603]_  = \new_[20749]_  | \new_[16604]_ ;
  assign \new_[21604]_  = ~\new_[18417]_  | ~\new_[21518]_ ;
  assign \new_[21605]_  = ~\new_[18417]_  | ~\new_[21518]_ ;
  assign \new_[21606]_  = ~\new_[21607]_ ;
  assign \new_[21607]_  = \new_[17071]_ ;
  assign \new_[21608]_  = ~\new_[21609]_ ;
  assign \new_[21609]_  = \new_[21610]_ ;
  assign \new_[21610]_  = ~\new_[21611]_ ;
  assign \new_[21611]_  = ~\new_[18625]_ ;
  assign \new_[21612]_  = ~\new_[12295]_ ;
  assign \new_[21613]_  = ~\new_[3418]_  | ~\new_[5340]_ ;
  assign \new_[21614]_  = ~\new_[3418]_  | ~\new_[5340]_ ;
  assign \new_[21615]_  = ~\new_[17114]_  | ~\new_[21505]_ ;
  assign \new_[21616]_  = ~\new_[17114]_  | ~\new_[21505]_ ;
  assign \new_[21617]_  = \new_[3740]_  | \new_[4216]_  | \new_[5475]_  | \new_[4001]_ ;
  assign \new_[21618]_  = \new_[3740]_  | \new_[4216]_  | \new_[5475]_  | \new_[4001]_ ;
  assign \new_[21619]_  = \new_[3255]_ ;
  assign \new_[21620]_  = ~\new_[13546]_ ;
  assign \new_[21621]_  = ~\new_[21622]_ ;
  assign \new_[21622]_  = ~\new_[17149]_ ;
  assign \new_[21623]_  = ~\new_[12646]_ ;
  assign \new_[21624]_  = ~\new_[21625]_ ;
  assign \new_[21625]_  = ~\new_[21626]_ ;
  assign \new_[21626]_  = ~\new_[21627]_ ;
  assign \new_[21627]_  = \new_[20810]_ ;
  assign \new_[21628]_  = ~\new_[21632]_ ;
  assign \new_[21629]_  = ~\new_[21630]_ ;
  assign \new_[21630]_  = ~\new_[21631]_ ;
  assign \new_[21631]_  = ~\new_[21632]_ ;
  assign \new_[21632]_  = ~\new_[21635]_ ;
  assign \new_[21633]_  = ~\new_[21634]_ ;
  assign \new_[21634]_  = \new_[21635]_ ;
  assign \new_[21635]_  = ~\new_[1043]_ ;
  assign \new_[21636]_  = ~\new_[21637]_ ;
  assign \new_[21637]_  = ~\new_[21638]_ ;
  assign \new_[21638]_  = ~\new_[1043]_ ;
  assign \new_[21639]_  = ~\new_[20459]_ ;
  assign \new_[21640]_  = ~\new_[19129]_ ;
  assign \new_[21641]_  = ~\new_[21642]_ ;
  assign \new_[21642]_  = \new_[21643]_ ;
  assign \new_[21643]_  = \new_[19129]_ ;
  assign \new_[21644]_  = ~\new_[20171]_  | ~\new_[19516]_ ;
  assign \new_[21645]_  = ~\new_[20171]_  | ~\new_[19516]_ ;
  assign \new_[21646]_  = ~\new_[4122]_  | ~\new_[3767]_  | ~\new_[3800]_  | ~\new_[4469]_ ;
  assign \new_[21647]_  = ~\new_[4122]_  | ~\new_[3767]_  | ~\new_[3800]_  | ~\new_[4469]_ ;
  assign \new_[21648]_  = ~\new_[20282]_  | ~\new_[20288]_ ;
  assign \new_[21649]_  = ~\new_[20282]_  | ~\new_[20288]_ ;
  assign \new_[21650]_  = ~\new_[21651]_ ;
  assign \new_[21651]_  = \new_[17162]_ ;
  assign \new_[21652]_  = ~\new_[17162]_ ;
  assign \new_[21653]_  = \new_[21654]_ ;
  assign \new_[21654]_  = ~\new_[18095]_ ;
  assign \new_[21655]_  = ~\new_[21656]_ ;
  assign \new_[21656]_  = ~\new_[21657]_ ;
  assign \new_[21657]_  = ~\new_[980]_ ;
  assign \new_[21658]_  = ~\new_[21659]_ ;
  assign \new_[21659]_  = \new_[21660]_ ;
  assign \new_[21660]_  = ~\new_[980]_ ;
  assign \new_[21661]_  = ~\new_[21662]_ ;
  assign \new_[21662]_  = ~\new_[13855]_ ;
  assign \new_[21663]_  = ~\new_[21610]_  & ~\new_[18968]_ ;
  assign \new_[21664]_  = ~\new_[21610]_  & ~\new_[18968]_ ;
  assign \new_[21665]_  = ~\new_[15038]_  & ~\new_[19697]_ ;
  assign \new_[21666]_  = ~\new_[15038]_  & ~\new_[19697]_ ;
  assign \new_[21667]_  = \new_[10730]_  ^ \new_[3484]_ ;
  assign \new_[21668]_  = \new_[10730]_  ^ \new_[3484]_ ;
  assign \new_[21669]_  = ~\new_[16609]_ ;
  assign \new_[21670]_  = ~\new_[21671]_ ;
  assign \new_[21671]_  = \new_[21673]_ ;
  assign \new_[21672]_  = ~\new_[21673]_ ;
  assign \new_[21673]_  = \new_[16609]_ ;
  assign \new_[21674]_  = ~\new_[15514]_  | ~\new_[19084]_ ;
  assign \new_[21675]_  = ~\new_[15514]_  | ~\new_[19084]_ ;
  assign \new_[21676]_  = ~\new_[21287]_  & ~\new_[21291]_ ;
  assign \new_[21677]_  = ~\new_[21287]_  & ~\new_[21291]_ ;
  assign \new_[21678]_  = ~\new_[21679]_ ;
  assign \new_[21679]_  = ~\new_[21680]_ ;
  assign \new_[21680]_  = ~\new_[21681]_ ;
  assign \new_[21681]_  = ~\new_[19913]_ ;
  assign \new_[21682]_  = ~\new_[18432]_ ;
  assign \new_[21683]_  = \new_[3683]_ ;
  assign \new_[21684]_  = \new_[21686]_ ;
  assign \new_[21685]_  = ~\new_[21687]_ ;
  assign \new_[21686]_  = ~\new_[21687]_ ;
  assign \new_[21687]_  = \new_[933]_ ;
  assign \new_[21688]_  = ~\new_[21691]_ ;
  assign \new_[21689]_  = ~\new_[21690]_ ;
  assign \new_[21690]_  = \new_[21691]_ ;
  assign \new_[21691]_  = ~\new_[21698]_ ;
  assign \new_[21692]_  = \new_[21693]_ ;
  assign \new_[21693]_  = \new_[21698]_ ;
  assign \new_[21694]_  = ~\new_[21696]_ ;
  assign \new_[21695]_  = ~\new_[21696]_ ;
  assign \new_[21696]_  = ~\new_[21697]_ ;
  assign \new_[21697]_  = \new_[21698]_ ;
  assign \new_[21698]_  = ~\new_[933]_ ;
  assign \new_[21699]_  = ~\new_[20042]_  | ~\new_[20041]_  | ~\new_[20038]_  | ~\new_[20039]_ ;
  assign \new_[21700]_  = ~\new_[20042]_  | ~\new_[20041]_  | ~\new_[20038]_  | ~\new_[20039]_ ;
  assign \new_[21701]_  = ~\new_[21704]_ ;
  assign \new_[21702]_  = ~\new_[21703]_ ;
  assign \new_[21703]_  = \new_[21704]_ ;
  assign \new_[21704]_  = ~\new_[17018]_ ;
  assign \new_[21705]_  = ~\new_[14102]_ ;
  assign \new_[21706]_  = ~\new_[14935]_ ;
  assign \new_[21707]_  = ~\new_[21710]_ ;
  assign \new_[21708]_  = ~\new_[21710]_ ;
  assign \new_[21709]_  = ~\new_[21710]_ ;
  assign \new_[21710]_  = ~\new_[3214]_ ;
  assign \new_[21711]_  = ~\new_[21712]_ ;
  assign \new_[21712]_  = \new_[18211]_ ;
  assign \new_[21713]_  = ~\new_[18211]_ ;
  assign \new_[21714]_  = ~\new_[16174]_ ;
  always @ (posedge clock) begin
    \\sa22_reg[4]  <= n778;
    \\sa02_reg[1]  <= n783;
    \\sa01_reg[1]  <= n788;
    \\sa00_reg[1]  <= n793;
    \\sa03_reg[4]  <= n798;
    \\sa03_reg[3]  <= n803;
    \\sa33_reg[0]  <= n808;
    \\sa02_reg[4]  <= n813;
    \\sa12_reg[3]  <= n818;
    \\sa32_reg[3]  <= n823;
    \\sa32_reg[0]  <= n828;
    \\sa22_reg[3]  <= n833;
    \\sa31_reg[0]  <= n838;
    \\sa02_reg[3]  <= n843;
    \\sa20_reg[3]  <= n848;
    \\sa30_reg[0]  <= n853;
    \\sa00_reg[4]  <= n858;
    \\sa10_reg[0]  <= n863;
    \\sa03_reg[0]  <= n868;
    \\sa33_reg[3]  <= n873;
    \\sa13_reg[0]  <= n878;
    \\sa02_reg[6]  <= n883;
    \\sa22_reg[5]  <= n888;
    \\sa13_reg[4]  <= n893;
    \\sa03_reg[1]  <= n898;
    \\sa32_reg[5]  <= n903;
    \\sa12_reg[1]  <= n908;
    \\sa13_reg[3]  <= n913;
    \\sa23_reg[3]  <= n918;
    \\sa02_reg[0]  <= n923;
    \\sa12_reg[0]  <= n928;
    \\sa21_reg[4]  <= n933;
    \\sa01_reg[4]  <= n938;
    \\sa31_reg[5]  <= n943;
    \\sa11_reg[1]  <= n948;
    \\sa21_reg[3]  <= n953;
    \\sa01_reg[0]  <= n958;
    \\sa21_reg[5]  <= n963;
    \\sa11_reg[0]  <= n968;
    \\sa10_reg[1]  <= n973;
    \\sa20_reg[1]  <= n978;
    \\sa00_reg[5]  <= n983;
    \\sa30_reg[6]  <= n988;
    \\sa10_reg[3]  <= n993;
    \\sa00_reg[0]  <= n998;
    \\sa00_reg[7]  <= n1003;
    \\sa23_reg[6]  <= n1008;
    \\sa13_reg[6]  <= n1013;
    \\sa13_reg[1]  <= n1018;
    \\sa33_reg[4]  <= n1023;
    \\sa23_reg[7]  <= n1028;
    \\sa33_reg[7]  <= n1033;
    \\sa03_reg[6]  <= n1038;
    \\sa23_reg[0]  <= n1043;
    \\sa02_reg[5]  <= n1048;
    \\sa32_reg[6]  <= n1053;
    \\sa12_reg[6]  <= n1058;
    \\sa22_reg[6]  <= n1063;
    \\sa22_reg[1]  <= n1068;
    \\sa12_reg[4]  <= n1073;
    \\sa22_reg[0]  <= n1078;
    \\sa01_reg[6]  <= n1083;
    \\sa11_reg[6]  <= n1088;
    \\sa31_reg[6]  <= n1093;
    \\sa01_reg[5]  <= n1098;
    \\sa21_reg[1]  <= n1103;
    \\sa11_reg[3]  <= n1108;
    \\sa01_reg[3]  <= n1113;
    \\sa21_reg[0]  <= n1118;
    \\sa31_reg[3]  <= n1123;
    \\sa10_reg[5]  <= n1128;
    \\sa30_reg[5]  <= n1133;
    \\sa20_reg[5]  <= n1138;
    \\sa30_reg[1]  <= n1143;
    \\sa00_reg[3]  <= n1148;
    \\sa30_reg[4]  <= n1153;
    \\sa10_reg[4]  <= n1158;
    \\sa10_reg[6]  <= n1163;
    \\sa20_reg[0]  <= n1168;
    \\sa30_reg[3]  <= n1173;
    \\sa30_reg[2]  <= n1178;
    \\sa00_reg[6]  <= n1183;
    \\sa20_reg[6]  <= n1188;
    \\sa20_reg[2]  <= n1193;
    \\sa03_reg[5]  <= n1198;
    \\sa23_reg[4]  <= n1203;
    \\sa33_reg[5]  <= n1208;
    \\sa23_reg[5]  <= n1213;
    \\sa33_reg[1]  <= n1218;
    \\sa23_reg[1]  <= n1223;
    \\sa33_reg[2]  <= n1228;
    \\sa03_reg[2]  <= n1233;
    \\sa23_reg[2]  <= n1238;
    \\sa13_reg[7]  <= n1243;
    \\sa03_reg[7]  <= n1248;
    \\sa12_reg[5]  <= n1253;
    \\sa32_reg[1]  <= n1258;
    \\sa22_reg[7]  <= n1263;
    \\sa02_reg[7]  <= n1268;
    \\sa12_reg[7]  <= n1273;
    \\sa21_reg[6]  <= n1278;
    \\sa11_reg[5]  <= n1283;
    \\sa31_reg[1]  <= n1288;
    \\sa11_reg[4]  <= n1293;
    \\sa31_reg[2]  <= n1298;
    \\sa01_reg[7]  <= n1303;
    \\sa21_reg[2]  <= n1308;
    \\sa20_reg[4]  <= n1313;
    \\sa20_reg[7]  <= n1318;
    \\sa10_reg[7]  <= n1323;
    \\sa30_reg[7]  <= n1328;
    \\sa13_reg[5]  <= n1333;
    \\sa33_reg[6]  <= n1338;
    \\sa32_reg[2]  <= n1343;
    \\sa02_reg[2]  <= n1348;
    \\sa12_reg[2]  <= n1353;
    \\sa22_reg[2]  <= n1358;
    \\sa01_reg[2]  <= n1363;
    \\sa11_reg[2]  <= n1368;
    \\sa11_reg[7]  <= n1373;
    \\sa00_reg[2]  <= n1378;
    \\u0_w_reg[2][19]  <= n1383;
    \\sa10_reg[2]  <= n1388;
    \\sa13_reg[2]  <= n1393;
    \\sa32_reg[7]  <= n1398;
    \\sa32_reg[4]  <= n1403;
    \\sa31_reg[7]  <= n1408;
    \\sa31_reg[4]  <= n1413;
    \\sa21_reg[7]  <= n1418;
    \\u0_w_reg[3][29]  <= n1423;
    \\u0_w_reg[0][19]  <= n1428;
    \\u0_w_reg[1][19]  <= n1433;
    \\u0_w_reg[3][19]  <= n1438;
    \\u0_w_reg[2][21]  <= n1443;
    \\u0_w_reg[0][27]  <= n1448;
    \\u0_w_reg[1][27]  <= n1453;
    \\u0_w_reg[2][27]  <= n1458;
    \\u0_w_reg[2][11]  <= n1463;
    \\u0_w_reg[3][27]  <= n1468;
    \\u0_w_reg[3][24]  <= n1473;
    \\u0_w_reg[2][29]  <= n1478;
    \\u0_w_reg[0][29]  <= n1483;
    \\u0_w_reg[2][5]  <= n1488;
    \\u0_w_reg[2][3]  <= n1493;
    \\u0_w_reg[1][29]  <= n1498;
    \\u0_w_reg[0][30]  <= n1503;
    \\u0_w_reg[1][30]  <= n1508;
    \\u0_w_reg[3][30]  <= n1513;
    \\u0_w_reg[0][21]  <= n1518;
    \\u0_w_reg[1][21]  <= n1523;
    \\u0_w_reg[2][0]  <= n1528;
    \\u0_w_reg[2][10]  <= n1533;
    \\u0_w_reg[2][14]  <= n1538;
    \\u0_w_reg[2][30]  <= n1543;
    \\u0_w_reg[2][16]  <= n1548;
    \\u0_w_reg[2][8]  <= n1553;
    \\u0_w_reg[2][15]  <= n1558;
    \\u0_w_reg[3][21]  <= n1563;
    \\text_out_reg[12]  <= n1568;
    \\u0_w_reg[2][12]  <= n1573;
    \\u0_w_reg[0][24]  <= n1578;
    \\u0_w_reg[0][31]  <= n1583;
    \\u0_w_reg[1][24]  <= n1588;
    \\u0_w_reg[1][31]  <= n1593;
    \\u0_w_reg[2][24]  <= n1598;
    \\u0_w_reg[2][31]  <= n1603;
    \\u0_w_reg[3][31]  <= n1608;
    \\u0_w_reg[0][5]  <= n1613;
    \\u0_w_reg[2][22]  <= n1618;
    \\u0_w_reg[2][6]  <= n1623;
    \\u0_w_reg[3][5]  <= n1628;
    \\u0_w_reg[0][11]  <= n1633;
    \\u0_w_reg[1][11]  <= n1638;
    \\u0_w_reg[2][17]  <= n1643;
    \\u0_w_reg[2][9]  <= n1648;
    \\u0_w_reg[3][11]  <= n1653;
    \\text_out_reg[125]  <= n1658;
    \\text_out_reg[44]  <= n1663;
    \\u0_w_reg[1][5]  <= n1668;
    \\u0_w_reg[2][13]  <= n1673;
    \\u0_w_reg[1][3]  <= n1678;
    \\u0_w_reg[0][3]  <= n1683;
    \\u0_w_reg[3][3]  <= n1688;
    \\u0_w_reg[2][4]  <= n1693;
    \\u0_w_reg[1][28]  <= n1698;
    \\u0_w_reg[3][28]  <= n1703;
    \\text_out_reg[93]  <= n1708;
    \\u0_w_reg[0][0]  <= n1713;
    \\text_out_reg[61]  <= n1718;
    \\u0_w_reg[0][16]  <= n1723;
    \\u0_w_reg[1][0]  <= n1728;
    \\u0_w_reg[3][0]  <= n1733;
    \\u0_w_reg[1][16]  <= n1738;
    \\u0_w_reg[3][16]  <= n1743;
    \\text_out_reg[101]  <= n1748;
    \\text_out_reg[108]  <= n1753;
    \\text_out_reg[43]  <= n1758;
    \\text_out_reg[109]  <= n1763;
    \\text_out_reg[117]  <= n1768;
    \\text_out_reg[76]  <= n1773;
    \\text_out_reg[111]  <= n1778;
    \\text_out_reg[48]  <= n1783;
    \\text_out_reg[80]  <= n1788;
    \\text_out_reg[112]  <= n1793;
    \\text_out_reg[46]  <= n1798;
    \\text_out_reg[126]  <= n1803;
    \\text_out_reg[10]  <= n1808;
    \\u0_w_reg[3][26]  <= n1813;
    \\u0_w_reg[1][26]  <= n1818;
    \\u0_w_reg[2][26]  <= n1823;
    \\u0_w_reg[0][26]  <= n1828;
    \\text_out_reg[0]  <= n1833;
    \\text_out_reg[4]  <= n1838;
    \\text_out_reg[6]  <= n1843;
    \\text_out_reg[32]  <= n1848;
    \\u0_w_reg[3][14]  <= n1853;
    \\text_out_reg[64]  <= n1858;
    \\u0_w_reg[2][18]  <= n1863;
    \\u0_w_reg[2][2]  <= n1868;
    \\u0_w_reg[2][23]  <= n1873;
    \\u0_w_reg[2][20]  <= n1878;
    \\u0_w_reg[2][28]  <= n1883;
    \\u0_w_reg[0][10]  <= n1888;
    \\u0_w_reg[0][13]  <= n1893;
    \\u0_w_reg[0][15]  <= n1898;
    \\u0_w_reg[0][8]  <= n1903;
    \\u0_w_reg[1][13]  <= n1908;
    \\u0_w_reg[1][14]  <= n1913;
    \\u0_w_reg[1][15]  <= n1918;
    \\u0_w_reg[1][10]  <= n1923;
    \\u0_w_reg[1][8]  <= n1928;
    \\u0_w_reg[3][10]  <= n1933;
    \\u0_w_reg[3][13]  <= n1938;
    \\u0_w_reg[3][15]  <= n1943;
    \\u0_w_reg[3][8]  <= n1948;
    \\text_out_reg[29]  <= n1953;
    \\text_out_reg[51]  <= n1958;
    \\text_out_reg[45]  <= n1963;
    \\text_out_reg[105]  <= n1968;
    \\text_out_reg[104]  <= n1973;
    \\text_out_reg[77]  <= n1978;
    \\text_out_reg[13]  <= n1983;
    \\text_out_reg[115]  <= n1988;
    \\text_out_reg[19]  <= n1993;
    \\text_out_reg[47]  <= n1998;
    \\text_out_reg[42]  <= n2003;
    \\text_out_reg[79]  <= n2008;
    \\text_out_reg[74]  <= n2013;
    \\text_out_reg[100]  <= n2018;
    \\text_out_reg[62]  <= n2023;
    \\text_out_reg[94]  <= n2028;
    \\text_out_reg[110]  <= n2033;
    \\text_out_reg[78]  <= n2038;
    \\text_out_reg[121]  <= n2043;
    \\text_out_reg[124]  <= n2048;
    \\u0_w_reg[0][28]  <= n2053;
    \\u0_w_reg[0][14]  <= n2058;
    \\u0_w_reg[2][1]  <= n2063;
    \\u0_w_reg[2][7]  <= n2068;
    \\text_out_reg[21]  <= n2073;
    \\text_out_reg[120]  <= n2078;
    \\text_out_reg[16]  <= n2083;
    \\text_out_reg[5]  <= n2088;
    \\text_out_reg[37]  <= n2093;
    \\text_out_reg[35]  <= n2098;
    \\text_out_reg[69]  <= n2103;
    \\text_out_reg[67]  <= n2108;
    \\u0_w_reg[2][25]  <= n2113;
    \\u0_w_reg[1][25]  <= n2118;
    \\u0_w_reg[0][12]  <= n2123;
    \\u0_w_reg[3][12]  <= n2128;
    \\u0_w_reg[0][22]  <= n2133;
    \\u0_w_reg[0][6]  <= n2138;
    \\u0_w_reg[1][22]  <= n2143;
    \\u0_w_reg[1][6]  <= n2148;
    \\u0_w_reg[3][22]  <= n2153;
    \\u0_w_reg[3][6]  <= n2158;
    \\text_out_reg[56]  <= n2163;
    \\u0_w_reg[0][17]  <= n2168;
    \\text_out_reg[88]  <= n2173;
    \\u0_w_reg[0][9]  <= n2178;
    \\u0_w_reg[1][17]  <= n2183;
    \\text_out_reg[53]  <= n2188;
    \\u0_w_reg[1][9]  <= n2193;
    \\u0_w_reg[3][17]  <= n2198;
    \\u0_w_reg[3][9]  <= n2203;
    \\text_out_reg[85]  <= n2208;
    \\text_out_reg[83]  <= n2213;
    \\text_out_reg[24]  <= n2218;
    \\text_out_reg[75]  <= n2223;
    \\text_out_reg[123]  <= n2228;
    \\text_out_reg[73]  <= n2233;
    \\text_out_reg[106]  <= n2238;
    \\text_out_reg[82]  <= n2243;
    \\text_out_reg[30]  <= n2248;
    \\text_out_reg[23]  <= n2253;
    \\text_out_reg[18]  <= n2258;
    \\text_out_reg[114]  <= n2263;
    \\text_out_reg[57]  <= n2268;
    \\text_out_reg[89]  <= n2273;
    \\text_out_reg[60]  <= n2278;
    \\u0_w_reg[1][12]  <= n2283;
    \\u0_w_reg[3][25]  <= n2288;
    \\u0_w_reg[0][25]  <= n2293;
    \\text_out_reg[41]  <= n2298;
    \\text_out_reg[1]  <= n2303;
    \\text_out_reg[7]  <= n2308;
    \\text_out_reg[38]  <= n2313;
    \\text_out_reg[36]  <= n2318;
    \\text_out_reg[33]  <= n2323;
    \\text_out_reg[39]  <= n2328;
    \\text_out_reg[68]  <= n2333;
    \\text_out_reg[70]  <= n2338;
    \\text_out_reg[71]  <= n2343;
    \\text_out_reg[50]  <= n2348;
    \\text_out_reg[59]  <= n2353;
    \\text_out_reg[91]  <= n2358;
    \\text_out_reg[40]  <= n2363;
    \\text_out_reg[72]  <= n2368;
    \\u0_w_reg[0][4]  <= n2373;
    \\u0_w_reg[1][4]  <= n2378;
    \\u0_w_reg[3][4]  <= n2383;
    \\text_out_reg[9]  <= n2388;
    \\text_out_reg[31]  <= n2393;
    \\text_out_reg[102]  <= n2398;
    \\text_out_reg[55]  <= n2403;
    \\text_out_reg[54]  <= n2408;
    \\text_out_reg[90]  <= n2413;
    \\text_out_reg[119]  <= n2418;
    \\text_out_reg[22]  <= n2423;
    \\text_out_reg[103]  <= n2428;
    \\text_out_reg[15]  <= n2433;
    \\text_out_reg[14]  <= n2438;
    \\text_out_reg[92]  <= n2443;
    \\text_out_reg[116]  <= n2448;
    \\text_out_reg[66]  <= n2453;
    \\text_out_reg[11]  <= n2458;
    \\text_out_reg[34]  <= n2463;
    \\text_out_reg[27]  <= n2468;
    \\text_out_reg[2]  <= n2473;
    \\text_out_reg[28]  <= n2478;
    \\text_out_reg[25]  <= n2483;
    \\u0_w_reg[3][7]  <= n2488;
    \\text_out_reg[58]  <= n2493;
    \\text_out_reg[122]  <= n2498;
    \\text_out_reg[3]  <= n2503;
    \\u0_w_reg[1][18]  <= n2508;
    \\text_out_reg[65]  <= n2513;
    \\u0_w_reg[1][7]  <= n2518;
    \\u0_w_reg[0][2]  <= n2523;
    \\u0_w_reg[1][2]  <= n2528;
    \\u0_w_reg[3][18]  <= n2533;
    \\u0_w_reg[3][2]  <= n2538;
    \\u0_w_reg[0][23]  <= n2543;
    \\u0_w_reg[3][23]  <= n2548;
    \\text_out_reg[107]  <= n2553;
    \\u0_w_reg[0][20]  <= n2558;
    \\u0_w_reg[1][20]  <= n2563;
    \\u0_w_reg[3][20]  <= n2568;
    \\text_out_reg[97]  <= n2573;
    \\text_out_reg[63]  <= n2578;
    \\text_out_reg[96]  <= n2583;
    \\text_out_reg[113]  <= n2588;
    \\text_out_reg[127]  <= n2593;
    \\text_out_reg[118]  <= n2598;
    \\text_out_reg[26]  <= n2603;
    \\text_out_reg[98]  <= n2608;
    \\text_out_reg[52]  <= n2613;
    \\text_out_reg[84]  <= n2618;
    \\text_out_reg[95]  <= n2623;
    \\u0_w_reg[0][7]  <= n2628;
    \\u0_w_reg[0][18]  <= n2633;
    \\u0_w_reg[3][1]  <= n2638;
    \\u0_w_reg[1][1]  <= n2643;
    \\text_out_reg[20]  <= n2648;
    \\u0_w_reg[1][23]  <= n2653;
    \\u0_w_reg[0][1]  <= n2658;
    \\text_out_reg[86]  <= n2663;
    \\text_out_reg[81]  <= n2668;
    \\text_out_reg[99]  <= n2673;
    \\text_out_reg[87]  <= n2678;
    \\text_out_reg[17]  <= n2683;
    \\text_out_reg[49]  <= n2688;
    \\text_out_reg[8]  <= n2693;
    \\u0_r0_out_reg[28]  <= n2698;
    \\u0_r0_out_reg[26]  <= n2703;
    \\u0_r0_out_reg[27]  <= n2708;
    \\dcnt_reg[3]  <= n2713;
    \\u0_r0_out_reg[29]  <= n2718;
    \\u0_r0_out_reg[25]  <= n2723;
    \\dcnt_reg[2]  <= n2728;
    \\u0_r0_out_reg[30]  <= n2733;
    \\u0_r0_out_reg[31]  <= n2738;
    \\dcnt_reg[1]  <= n2743;
    \\u0_r0_out_reg[24]  <= n2748;
    \\dcnt_reg[0]  <= n2753;
    \\u0_r0_rcnt_reg[3]  <= n2758;
    done_reg <= n2763;
    \\text_in_r_reg[116]  <= n2768;
    \\text_in_r_reg[111]  <= n2773;
    \\text_in_r_reg[37]  <= n2778;
    \\text_in_r_reg[14]  <= n2783;
    \\text_in_r_reg[67]  <= n2788;
    \\text_in_r_reg[47]  <= n2793;
    \\text_in_r_reg[18]  <= n2798;
    \\text_in_r_reg[0]  <= n2803;
    \\text_in_r_reg[68]  <= n2808;
    \\text_in_r_reg[49]  <= n2813;
    \\text_in_r_reg[42]  <= n2818;
    \\text_in_r_reg[127]  <= n2823;
    \\text_in_r_reg[64]  <= n2828;
    \\text_in_r_reg[54]  <= n2833;
    \\text_in_r_reg[35]  <= n2838;
    \\text_in_r_reg[6]  <= n2843;
    \\text_in_r_reg[17]  <= n2848;
    \\text_in_r_reg[108]  <= n2853;
    \\text_in_r_reg[11]  <= n2858;
    \\text_in_r_reg[123]  <= n2863;
    \\text_in_r_reg[24]  <= n2868;
    \\text_in_r_reg[26]  <= n2873;
    \\text_in_r_reg[29]  <= n2878;
    \\text_in_r_reg[46]  <= n2883;
    \\text_in_r_reg[55]  <= n2888;
    \\text_in_r_reg[61]  <= n2893;
    \\text_in_r_reg[63]  <= n2898;
    \\text_in_r_reg[78]  <= n2903;
    \\text_in_r_reg[81]  <= n2908;
    \\text_in_r_reg[86]  <= n2913;
    \\text_in_r_reg[8]  <= n2918;
    \\text_in_r_reg[99]  <= n2923;
    \\text_in_r_reg[91]  <= n2928;
    \\text_in_r_reg[39]  <= n2933;
    \\text_in_r_reg[60]  <= n2938;
    \\text_in_r_reg[103]  <= n2943;
    \\text_in_r_reg[23]  <= n2948;
    \\text_in_r_reg[58]  <= n2953;
    \\text_in_r_reg[3]  <= n2958;
    \\text_in_r_reg[118]  <= n2963;
    \\text_in_r_reg[59]  <= n2968;
    \\text_in_r_reg[96]  <= n2973;
    \\text_in_r_reg[70]  <= n2978;
    \\text_in_r_reg[51]  <= n2983;
    \\text_in_r_reg[92]  <= n2988;
    \\text_in_r_reg[107]  <= n2993;
    \\text_in_r_reg[28]  <= n2998;
    \\text_in_r_reg[77]  <= n3003;
    \\text_in_r_reg[1]  <= n3008;
    \\text_in_r_reg[19]  <= n3013;
    \\text_in_r_reg[56]  <= n3018;
    \\text_in_r_reg[90]  <= n3023;
    \\text_in_r_reg[69]  <= n3028;
    \\text_in_r_reg[12]  <= n3033;
    \\text_in_r_reg[85]  <= n3038;
    \\text_in_r_reg[80]  <= n3043;
    \\text_in_r_reg[66]  <= n3048;
    \\text_in_r_reg[9]  <= n3053;
    \\text_in_r_reg[53]  <= n3058;
    \\text_in_r_reg[45]  <= n3063;
    \\text_in_r_reg[52]  <= n3068;
    \\text_in_r_reg[97]  <= n3073;
    \\text_in_r_reg[10]  <= n3078;
    \\text_in_r_reg[34]  <= n3083;
    \\text_in_r_reg[110]  <= n3088;
    \\text_in_r_reg[30]  <= n3093;
    \\text_in_r_reg[104]  <= n3098;
    \\text_in_r_reg[65]  <= n3103;
    \\text_in_r_reg[79]  <= n3108;
    \\text_in_r_reg[7]  <= n3113;
    \\text_in_r_reg[82]  <= n3118;
    \\text_in_r_reg[126]  <= n3123;
    \\text_in_r_reg[105]  <= n3128;
    \\text_in_r_reg[13]  <= n3133;
    \\text_in_r_reg[120]  <= n3138;
    \\text_in_r_reg[84]  <= n3143;
    \\text_in_r_reg[74]  <= n3148;
    \\text_in_r_reg[16]  <= n3153;
    \\text_in_r_reg[40]  <= n3158;
    \\text_in_r_reg[15]  <= n3163;
    \\text_in_r_reg[121]  <= n3168;
    \\text_in_r_reg[41]  <= n3173;
    \\text_in_r_reg[36]  <= n3178;
    \\text_in_r_reg[20]  <= n3183;
    \\u0_r0_rcnt_reg[2]  <= n3188;
    \\text_in_r_reg[32]  <= n3193;
    \\text_in_r_reg[75]  <= n3198;
    \\text_in_r_reg[88]  <= n3203;
    \\text_in_r_reg[33]  <= n3208;
    \\u0_r0_rcnt_reg[1]  <= n3213;
    \\text_in_r_reg[125]  <= n3218;
    \\text_in_r_reg[2]  <= n3223;
    \\text_in_r_reg[44]  <= n3228;
    \\text_in_r_reg[72]  <= n3233;
    \\text_in_r_reg[101]  <= n3238;
    \\text_in_r_reg[106]  <= n3243;
    \\text_in_r_reg[4]  <= n3248;
    \\text_in_r_reg[43]  <= n3253;
    \\text_in_r_reg[112]  <= n3258;
    \\text_in_r_reg[93]  <= n3263;
    \\text_in_r_reg[73]  <= n3268;
    \\text_in_r_reg[50]  <= n3273;
    \\text_in_r_reg[100]  <= n3278;
    \\text_in_r_reg[114]  <= n3283;
    \\text_in_r_reg[25]  <= n3288;
    \\text_in_r_reg[57]  <= n3293;
    \\text_in_r_reg[95]  <= n3298;
    \\text_in_r_reg[124]  <= n3303;
    \\text_in_r_reg[115]  <= n3308;
    \\text_in_r_reg[98]  <= n3313;
    \\text_in_r_reg[31]  <= n3318;
    \\text_in_r_reg[122]  <= n3323;
    \\text_in_r_reg[119]  <= n3328;
    \\text_in_r_reg[102]  <= n3333;
    \\text_in_r_reg[76]  <= n3338;
    \\text_in_r_reg[113]  <= n3343;
    \\text_in_r_reg[94]  <= n3348;
    \\text_in_r_reg[62]  <= n3353;
    \\text_in_r_reg[48]  <= n3358;
    \\text_in_r_reg[27]  <= n3363;
    \\text_in_r_reg[109]  <= n3368;
    \\text_in_r_reg[117]  <= n3373;
    \\u0_r0_rcnt_reg[0]  <= n3378;
    \\text_in_r_reg[21]  <= n3383;
    \\text_in_r_reg[5]  <= n3388;
    \\text_in_r_reg[22]  <= n3393;
    \\text_in_r_reg[83]  <= n3398;
    \\text_in_r_reg[38]  <= n3403;
    \\text_in_r_reg[71]  <= n3408;
    \\text_in_r_reg[89]  <= n3413;
    \\text_in_r_reg[87]  <= n3418;
    ld_r_reg <= n3423;
  end
endmodule


