// Benchmark "testing" written by ABC on Thu Oct  8 22:16:38 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A9  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A9;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ , \new_[350]_ ,
    \new_[351]_ , \new_[352]_ , \new_[353]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[405]_ ,
    \new_[406]_ , \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ ,
    \new_[411]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[436]_ , \new_[437]_ , \new_[438]_ , \new_[439]_ , \new_[440]_ ,
    \new_[441]_ , \new_[442]_ , \new_[443]_ , \new_[444]_ , \new_[445]_ ,
    \new_[446]_ , \new_[447]_ , \new_[448]_ , \new_[449]_ , \new_[450]_ ,
    \new_[451]_ , \new_[452]_ , \new_[453]_ , \new_[454]_ , \new_[455]_ ,
    \new_[456]_ , \new_[457]_ , \new_[458]_ , \new_[459]_ , \new_[460]_ ,
    \new_[461]_ , \new_[462]_ , \new_[463]_ , \new_[464]_ , \new_[465]_ ,
    \new_[466]_ , \new_[467]_ , \new_[468]_ , \new_[469]_ , \new_[470]_ ,
    \new_[471]_ , \new_[472]_ , \new_[473]_ , \new_[474]_ , \new_[475]_ ,
    \new_[476]_ , \new_[477]_ , \new_[478]_ , \new_[479]_ , \new_[480]_ ,
    \new_[481]_ , \new_[482]_ , \new_[483]_ , \new_[484]_ , \new_[485]_ ,
    \new_[486]_ , \new_[487]_ , \new_[488]_ , \new_[489]_ , \new_[490]_ ,
    \new_[491]_ , \new_[492]_ , \new_[493]_ , \new_[494]_ , \new_[495]_ ,
    \new_[496]_ , \new_[497]_ , \new_[498]_ , \new_[499]_ , \new_[500]_ ,
    \new_[501]_ , \new_[502]_ , \new_[503]_ , \new_[504]_ , \new_[505]_ ,
    \new_[506]_ , \new_[507]_ , \new_[508]_ , \new_[509]_ , \new_[510]_ ,
    \new_[511]_ , \new_[512]_ , \new_[513]_ , \new_[514]_ , \new_[515]_ ,
    \new_[516]_ , \new_[517]_ , \new_[518]_ , \new_[519]_ , \new_[520]_ ,
    \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[525]_ ,
    \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ , \new_[530]_ ,
    \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ , \new_[535]_ ,
    \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ , \new_[540]_ ,
    \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ , \new_[545]_ ,
    \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ , \new_[550]_ ,
    \new_[551]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[566]_ , \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ ,
    \new_[571]_ , \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ ,
    \new_[576]_ , \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ ,
    \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[584]_ , \new_[585]_ ,
    \new_[586]_ , \new_[587]_ , \new_[588]_ , \new_[589]_ , \new_[590]_ ,
    \new_[591]_ , \new_[592]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[598]_ , \new_[599]_ , \new_[600]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ ,
    \new_[611]_ , \new_[612]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[616]_ , \new_[617]_ , \new_[618]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[626]_ , \new_[627]_ , \new_[628]_ , \new_[629]_ , \new_[630]_ ,
    \new_[631]_ , \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ ,
    \new_[636]_ , \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ ,
    \new_[641]_ , \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ ,
    \new_[646]_ , \new_[647]_ , \new_[648]_ , \new_[649]_ , \new_[650]_ ,
    \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[655]_ ,
    \new_[656]_ , \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ ,
    \new_[661]_ , \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ ,
    \new_[666]_ , \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ ,
    \new_[671]_ , \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ ,
    \new_[676]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ ,
    \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ ,
    \new_[686]_ , \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ ,
    \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ ,
    \new_[696]_ , \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ ,
    \new_[701]_ , \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ ,
    \new_[706]_ , \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ ,
    \new_[711]_ , \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ ,
    \new_[716]_ , \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ ,
    \new_[726]_ , \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ ,
    \new_[731]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[736]_ , \new_[737]_ , \new_[738]_ , \new_[739]_ , \new_[740]_ ,
    \new_[741]_ , \new_[742]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ ,
    \new_[746]_ , \new_[747]_ , \new_[748]_ , \new_[749]_ , \new_[750]_ ,
    \new_[751]_ , \new_[752]_ , \new_[753]_ , \new_[754]_ , \new_[755]_ ,
    \new_[756]_ , \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ ,
    \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ ,
    \new_[766]_ , \new_[767]_ , \new_[768]_ , \new_[769]_ , \new_[770]_ ,
    \new_[771]_ , \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ ,
    \new_[776]_ , \new_[777]_ , \new_[778]_ , \new_[779]_ , \new_[780]_ ,
    \new_[781]_ , \new_[782]_ , \new_[783]_ , \new_[784]_ , \new_[785]_ ,
    \new_[786]_ , \new_[787]_ , \new_[788]_ , \new_[789]_ , \new_[790]_ ,
    \new_[791]_ , \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ ,
    \new_[796]_ , \new_[797]_ , \new_[798]_ , \new_[799]_ , \new_[800]_ ,
    \new_[801]_ , \new_[802]_ , \new_[803]_ , \new_[804]_ , \new_[805]_ ,
    \new_[806]_ , \new_[807]_ , \new_[808]_ , \new_[809]_ , \new_[810]_ ,
    \new_[811]_ , \new_[812]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ ,
    \new_[816]_ , \new_[817]_ , \new_[818]_ , \new_[819]_ , \new_[820]_ ,
    \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[824]_ , \new_[825]_ ,
    \new_[826]_ , \new_[827]_ , \new_[828]_ , \new_[829]_ , \new_[830]_ ,
    \new_[831]_ , \new_[832]_ , \new_[833]_ , \new_[834]_ , \new_[835]_ ,
    \new_[836]_ , \new_[837]_ , \new_[838]_ , \new_[839]_ , \new_[840]_ ,
    \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[845]_ ,
    \new_[846]_ , \new_[847]_ , \new_[848]_ , \new_[849]_ , \new_[850]_ ,
    \new_[851]_ , \new_[852]_ , \new_[853]_ , \new_[854]_ , \new_[855]_ ,
    \new_[856]_ , \new_[857]_ , \new_[858]_ , \new_[859]_ , \new_[860]_ ,
    \new_[861]_ , \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[865]_ ,
    \new_[866]_ , \new_[867]_ , \new_[868]_ , \new_[869]_ , \new_[870]_ ,
    \new_[871]_ , \new_[872]_ , \new_[873]_ , \new_[874]_ , \new_[875]_ ,
    \new_[876]_ , \new_[877]_ , \new_[878]_ , \new_[879]_ , \new_[880]_ ,
    \new_[881]_ , \new_[882]_ , \new_[883]_ , \new_[884]_ , \new_[885]_ ,
    \new_[886]_ , \new_[887]_ , \new_[888]_ , \new_[889]_ , \new_[890]_ ,
    \new_[891]_ , \new_[892]_ , \new_[893]_ , \new_[894]_ , \new_[895]_ ,
    \new_[896]_ , \new_[897]_ , \new_[898]_ , \new_[899]_ , \new_[900]_ ,
    \new_[901]_ , \new_[902]_ , \new_[903]_ , \new_[904]_ , \new_[905]_ ,
    \new_[906]_ , \new_[907]_ , \new_[908]_ , \new_[909]_ , \new_[910]_ ,
    \new_[911]_ , \new_[912]_ , \new_[913]_ , \new_[914]_ , \new_[915]_ ,
    \new_[916]_ , \new_[917]_ , \new_[918]_ , \new_[919]_ , \new_[920]_ ,
    \new_[921]_ , \new_[922]_ , \new_[923]_ , \new_[924]_ , \new_[925]_ ,
    \new_[926]_ , \new_[927]_ , \new_[928]_ , \new_[929]_ , \new_[930]_ ,
    \new_[931]_ , \new_[932]_ , \new_[933]_ , \new_[934]_ , \new_[935]_ ,
    \new_[936]_ , \new_[937]_ , \new_[938]_ , \new_[939]_ , \new_[940]_ ,
    \new_[941]_ , \new_[942]_ , \new_[943]_ , \new_[944]_ , \new_[945]_ ,
    \new_[946]_ , \new_[947]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ ,
    \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[955]_ ,
    \new_[956]_ , \new_[957]_ , \new_[958]_ , \new_[959]_ , \new_[960]_ ,
    \new_[961]_ , \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ ,
    \new_[966]_ , \new_[967]_ , \new_[968]_ , \new_[969]_ , \new_[970]_ ,
    \new_[971]_ , \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[975]_ ,
    \new_[976]_ , \new_[977]_ , \new_[978]_ , \new_[979]_ , \new_[980]_ ,
    \new_[981]_ , \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ ,
    \new_[986]_ , \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ ,
    \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ ,
    \new_[996]_ , \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ ,
    \new_[1001]_ , \new_[1002]_ , \new_[1003]_ , \new_[1004]_ ,
    \new_[1005]_ , \new_[1006]_ , \new_[1007]_ , \new_[1008]_ ,
    \new_[1009]_ , \new_[1010]_ , \new_[1011]_ , \new_[1012]_ ,
    \new_[1013]_ , \new_[1014]_ , \new_[1015]_ , \new_[1016]_ ,
    \new_[1017]_ , \new_[1018]_ , \new_[1019]_ , \new_[1020]_ ,
    \new_[1021]_ , \new_[1022]_ , \new_[1023]_ , \new_[1024]_ ,
    \new_[1025]_ , \new_[1026]_ , \new_[1027]_ , \new_[1028]_ ,
    \new_[1029]_ , \new_[1030]_ , \new_[1031]_ , \new_[1032]_ ,
    \new_[1033]_ , \new_[1034]_ , \new_[1035]_ , \new_[1036]_ ,
    \new_[1037]_ , \new_[1038]_ , \new_[1039]_ , \new_[1040]_ ,
    \new_[1041]_ , \new_[1042]_ , \new_[1043]_ , \new_[1044]_ ,
    \new_[1045]_ , \new_[1046]_ , \new_[1047]_ , \new_[1048]_ ,
    \new_[1049]_ , \new_[1050]_ , \new_[1051]_ , \new_[1052]_ ,
    \new_[1053]_ , \new_[1054]_ , \new_[1055]_ , \new_[1056]_ ,
    \new_[1057]_ , \new_[1058]_ , \new_[1059]_ , \new_[1060]_ ,
    \new_[1061]_ , \new_[1062]_ , \new_[1063]_ , \new_[1064]_ ,
    \new_[1065]_ , \new_[1066]_ , \new_[1067]_ , \new_[1068]_ ,
    \new_[1069]_ , \new_[1070]_ , \new_[1071]_ , \new_[1072]_ ,
    \new_[1073]_ , \new_[1074]_ , \new_[1075]_ , \new_[1076]_ ,
    \new_[1077]_ , \new_[1078]_ , \new_[1079]_ , \new_[1080]_ ,
    \new_[1081]_ , \new_[1082]_ , \new_[1083]_ , \new_[1084]_ ,
    \new_[1085]_ , \new_[1086]_ , \new_[1087]_ , \new_[1088]_ ,
    \new_[1089]_ , \new_[1090]_ , \new_[1091]_ , \new_[1092]_ ,
    \new_[1093]_ , \new_[1094]_ , \new_[1095]_ , \new_[1096]_ ,
    \new_[1097]_ , \new_[1098]_ , \new_[1099]_ , \new_[1100]_ ,
    \new_[1101]_ , \new_[1102]_ , \new_[1103]_ , \new_[1104]_ ,
    \new_[1105]_ , \new_[1106]_ , \new_[1107]_ , \new_[1108]_ ,
    \new_[1109]_ , \new_[1110]_ , \new_[1111]_ , \new_[1112]_ ,
    \new_[1113]_ , \new_[1114]_ , \new_[1115]_ , \new_[1116]_ ,
    \new_[1117]_ , \new_[1118]_ , \new_[1119]_ , \new_[1120]_ ,
    \new_[1121]_ , \new_[1122]_ , \new_[1123]_ , \new_[1124]_ ,
    \new_[1125]_ , \new_[1126]_ , \new_[1127]_ , \new_[1128]_ ,
    \new_[1129]_ , \new_[1130]_ , \new_[1131]_ , \new_[1132]_ ,
    \new_[1133]_ , \new_[1134]_ , \new_[1135]_ , \new_[1136]_ ,
    \new_[1137]_ , \new_[1138]_ , \new_[1139]_ , \new_[1140]_ ,
    \new_[1141]_ , \new_[1142]_ , \new_[1143]_ , \new_[1144]_ ,
    \new_[1145]_ , \new_[1146]_ , \new_[1147]_ , \new_[1148]_ ,
    \new_[1149]_ , \new_[1150]_ , \new_[1151]_ , \new_[1152]_ ,
    \new_[1153]_ , \new_[1154]_ , \new_[1155]_ , \new_[1156]_ ,
    \new_[1157]_ , \new_[1158]_ , \new_[1159]_ , \new_[1160]_ ,
    \new_[1161]_ , \new_[1162]_ , \new_[1163]_ , \new_[1164]_ ,
    \new_[1165]_ , \new_[1166]_ , \new_[1167]_ , \new_[1168]_ ,
    \new_[1169]_ , \new_[1170]_ , \new_[1171]_ , \new_[1172]_ ,
    \new_[1173]_ , \new_[1174]_ , \new_[1175]_ , \new_[1176]_ ,
    \new_[1177]_ , \new_[1178]_ , \new_[1179]_ , \new_[1180]_ ,
    \new_[1181]_ , \new_[1182]_ , \new_[1183]_ , \new_[1184]_ ,
    \new_[1185]_ , \new_[1186]_ , \new_[1187]_ , \new_[1188]_ ,
    \new_[1189]_ , \new_[1190]_ , \new_[1191]_ , \new_[1192]_ ,
    \new_[1193]_ , \new_[1194]_ , \new_[1195]_ , \new_[1196]_ ,
    \new_[1197]_ , \new_[1198]_ , \new_[1199]_ , \new_[1200]_ ,
    \new_[1201]_ , \new_[1202]_ , \new_[1203]_ , \new_[1204]_ ,
    \new_[1205]_ , \new_[1206]_ , \new_[1207]_ , \new_[1208]_ ,
    \new_[1209]_ , \new_[1210]_ , \new_[1211]_ , \new_[1212]_ ,
    \new_[1213]_ , \new_[1214]_ , \new_[1215]_ , \new_[1216]_ ,
    \new_[1217]_ , \new_[1218]_ , \new_[1219]_ , \new_[1220]_ ,
    \new_[1221]_ , \new_[1222]_ , \new_[1223]_ , \new_[1224]_ ,
    \new_[1225]_ , \new_[1226]_ , \new_[1227]_ , \new_[1228]_ ,
    \new_[1229]_ , \new_[1230]_ , \new_[1231]_ , \new_[1232]_ ,
    \new_[1233]_ , \new_[1234]_ , \new_[1235]_ , \new_[1236]_ ,
    \new_[1237]_ , \new_[1238]_ , \new_[1239]_ , \new_[1240]_ ,
    \new_[1241]_ , \new_[1242]_ , \new_[1243]_ , \new_[1244]_ ,
    \new_[1245]_ , \new_[1246]_ , \new_[1247]_ , \new_[1248]_ ,
    \new_[1249]_ , \new_[1250]_ , \new_[1251]_ , \new_[1252]_ ,
    \new_[1253]_ , \new_[1254]_ , \new_[1255]_ , \new_[1256]_ ,
    \new_[1257]_ , \new_[1258]_ , \new_[1259]_ , \new_[1260]_ ,
    \new_[1261]_ , \new_[1262]_ , \new_[1263]_ , \new_[1264]_ ,
    \new_[1265]_ , \new_[1266]_ , \new_[1267]_ , \new_[1268]_ ,
    \new_[1269]_ , \new_[1270]_ , \new_[1271]_ , \new_[1272]_ ,
    \new_[1273]_ , \new_[1274]_ , \new_[1275]_ , \new_[1276]_ ,
    \new_[1277]_ , \new_[1278]_ , \new_[1279]_ , \new_[1280]_ ,
    \new_[1281]_ , \new_[1282]_ , \new_[1283]_ , \new_[1284]_ ,
    \new_[1285]_ , \new_[1286]_ , \new_[1287]_ , \new_[1288]_ ,
    \new_[1289]_ , \new_[1290]_ , \new_[1291]_ , \new_[1292]_ ,
    \new_[1293]_ , \new_[1294]_ , \new_[1295]_ , \new_[1296]_ ,
    \new_[1297]_ , \new_[1298]_ , \new_[1299]_ , \new_[1300]_ ,
    \new_[1301]_ , \new_[1302]_ , \new_[1303]_ , \new_[1304]_ ,
    \new_[1305]_ , \new_[1306]_ , \new_[1307]_ , \new_[1308]_ ,
    \new_[1309]_ , \new_[1310]_ , \new_[1311]_ , \new_[1312]_ ,
    \new_[1313]_ , \new_[1314]_ , \new_[1315]_ , \new_[1316]_ ,
    \new_[1317]_ , \new_[1318]_ , \new_[1319]_ , \new_[1320]_ ,
    \new_[1321]_ , \new_[1322]_ , \new_[1323]_ , \new_[1324]_ ,
    \new_[1325]_ , \new_[1326]_ , \new_[1327]_ , \new_[1328]_ ,
    \new_[1329]_ , \new_[1330]_ , \new_[1331]_ , \new_[1332]_ ,
    \new_[1333]_ , \new_[1334]_ , \new_[1335]_ , \new_[1336]_ ,
    \new_[1337]_ , \new_[1338]_ , \new_[1339]_ , \new_[1340]_ ,
    \new_[1341]_ , \new_[1342]_ , \new_[1343]_ , \new_[1344]_ ,
    \new_[1345]_ , \new_[1346]_ , \new_[1347]_ , \new_[1348]_ ,
    \new_[1349]_ , \new_[1350]_ , \new_[1351]_ , \new_[1352]_ ,
    \new_[1353]_ , \new_[1354]_ , \new_[1355]_ , \new_[1356]_ ,
    \new_[1357]_ , \new_[1358]_ , \new_[1359]_ , \new_[1360]_ ,
    \new_[1361]_ , \new_[1362]_ , \new_[1363]_ , \new_[1364]_ ,
    \new_[1365]_ , \new_[1366]_ , \new_[1367]_ , \new_[1368]_ ,
    \new_[1369]_ , \new_[1370]_ , \new_[1371]_ , \new_[1372]_ ,
    \new_[1373]_ , \new_[1374]_ , \new_[1375]_ , \new_[1376]_ ,
    \new_[1377]_ , \new_[1378]_ , \new_[1379]_ , \new_[1380]_ ,
    \new_[1381]_ , \new_[1382]_ , \new_[1383]_ , \new_[1384]_ ,
    \new_[1385]_ , \new_[1386]_ , \new_[1387]_ , \new_[1388]_ ,
    \new_[1389]_ , \new_[1390]_ , \new_[1391]_ , \new_[1392]_ ,
    \new_[1393]_ , \new_[1394]_ , \new_[1395]_ , \new_[1396]_ ,
    \new_[1397]_ , \new_[1398]_ , \new_[1399]_ , \new_[1400]_ ,
    \new_[1401]_ , \new_[1402]_ , \new_[1403]_ , \new_[1404]_ ,
    \new_[1405]_ , \new_[1406]_ , \new_[1407]_ , \new_[1408]_ ,
    \new_[1409]_ , \new_[1410]_ , \new_[1411]_ , \new_[1412]_ ,
    \new_[1413]_ , \new_[1414]_ , \new_[1415]_ , \new_[1416]_ ,
    \new_[1417]_ , \new_[1418]_ , \new_[1419]_ , \new_[1420]_ ,
    \new_[1421]_ , \new_[1422]_ , \new_[1423]_ , \new_[1424]_ ,
    \new_[1425]_ , \new_[1426]_ , \new_[1427]_ , \new_[1428]_ ,
    \new_[1429]_ , \new_[1430]_ , \new_[1431]_ , \new_[1432]_ ,
    \new_[1433]_ , \new_[1434]_ , \new_[1435]_ , \new_[1436]_ ,
    \new_[1437]_ , \new_[1438]_ , \new_[1439]_ , \new_[1440]_ ,
    \new_[1441]_ , \new_[1442]_ , \new_[1443]_ , \new_[1444]_ ,
    \new_[1445]_ , \new_[1446]_ , \new_[1447]_ , \new_[1448]_ ,
    \new_[1449]_ , \new_[1450]_ , \new_[1451]_ , \new_[1452]_ ,
    \new_[1453]_ , \new_[1454]_ , \new_[1455]_ , \new_[1456]_ ,
    \new_[1457]_ , \new_[1458]_ , \new_[1459]_ , \new_[1460]_ ,
    \new_[1461]_ , \new_[1462]_ , \new_[1463]_ , \new_[1464]_ ,
    \new_[1465]_ , \new_[1466]_ , \new_[1467]_ , \new_[1468]_ ,
    \new_[1469]_ , \new_[1470]_ , \new_[1471]_ , \new_[1472]_ ,
    \new_[1473]_ , \new_[1474]_ , \new_[1475]_ , \new_[1476]_ ,
    \new_[1477]_ , \new_[1478]_ , \new_[1479]_ , \new_[1480]_ ,
    \new_[1481]_ , \new_[1482]_ , \new_[1483]_ , \new_[1484]_ ,
    \new_[1485]_ , \new_[1486]_ , \new_[1487]_ , \new_[1488]_ ,
    \new_[1489]_ , \new_[1490]_ , \new_[1491]_ , \new_[1492]_ ,
    \new_[1493]_ , \new_[1494]_ , \new_[1495]_ , \new_[1496]_ ,
    \new_[1497]_ , \new_[1498]_ , \new_[1499]_ , \new_[1500]_ ,
    \new_[1501]_ , \new_[1502]_ , \new_[1503]_ , \new_[1504]_ ,
    \new_[1505]_ , \new_[1506]_ , \new_[1507]_ , \new_[1508]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1512]_ ,
    \new_[1513]_ , \new_[1514]_ , \new_[1515]_ , \new_[1516]_ ,
    \new_[1517]_ , \new_[1518]_ , \new_[1519]_ , \new_[1520]_ ,
    \new_[1521]_ , \new_[1522]_ , \new_[1523]_ , \new_[1524]_ ,
    \new_[1525]_ , \new_[1526]_ , \new_[1527]_ , \new_[1528]_ ,
    \new_[1529]_ , \new_[1530]_ , \new_[1531]_ , \new_[1532]_ ,
    \new_[1533]_ , \new_[1534]_ , \new_[1535]_ , \new_[1536]_ ,
    \new_[1537]_ , \new_[1538]_ , \new_[1539]_ , \new_[1540]_ ,
    \new_[1541]_ , \new_[1542]_ , \new_[1543]_ , \new_[1544]_ ,
    \new_[1545]_ , \new_[1546]_ , \new_[1547]_ , \new_[1548]_ ,
    \new_[1549]_ , \new_[1550]_ , \new_[1551]_ , \new_[1552]_ ,
    \new_[1553]_ , \new_[1554]_ , \new_[1555]_ , \new_[1556]_ ,
    \new_[1557]_ , \new_[1558]_ , \new_[1559]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1562]_ , \new_[1563]_ , \new_[1564]_ ,
    \new_[1565]_ , \new_[1566]_ , \new_[1567]_ , \new_[1568]_ ,
    \new_[1569]_ , \new_[1570]_ , \new_[1571]_ , \new_[1572]_ ,
    \new_[1573]_ , \new_[1574]_ , \new_[1575]_ , \new_[1576]_ ,
    \new_[1577]_ , \new_[1578]_ , \new_[1579]_ , \new_[1580]_ ,
    \new_[1581]_ , \new_[1582]_ , \new_[1583]_ , \new_[1584]_ ,
    \new_[1585]_ , \new_[1586]_ , \new_[1587]_ , \new_[1588]_ ,
    \new_[1589]_ , \new_[1590]_ , \new_[1591]_ , \new_[1592]_ ,
    \new_[1593]_ , \new_[1594]_ , \new_[1595]_ , \new_[1596]_ ,
    \new_[1597]_ , \new_[1598]_ , \new_[1599]_ , \new_[1600]_ ,
    \new_[1601]_ , \new_[1602]_ , \new_[1603]_ , \new_[1604]_ ,
    \new_[1605]_ , \new_[1606]_ , \new_[1607]_ , \new_[1608]_ ,
    \new_[1609]_ , \new_[1610]_ , \new_[1611]_ , \new_[1612]_ ,
    \new_[1613]_ , \new_[1614]_ , \new_[1615]_ , \new_[1616]_ ,
    \new_[1617]_ , \new_[1618]_ , \new_[1619]_ , \new_[1620]_ ,
    \new_[1621]_ , \new_[1622]_ , \new_[1623]_ , \new_[1624]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1627]_ , \new_[1628]_ ,
    \new_[1629]_ , \new_[1630]_ , \new_[1631]_ , \new_[1632]_ ,
    \new_[1633]_ , \new_[1634]_ , \new_[1635]_ , \new_[1636]_ ,
    \new_[1637]_ , \new_[1638]_ , \new_[1639]_ , \new_[1640]_ ,
    \new_[1641]_ , \new_[1642]_ , \new_[1643]_ , \new_[1644]_ ,
    \new_[1645]_ , \new_[1646]_ , \new_[1647]_ , \new_[1648]_ ,
    \new_[1649]_ , \new_[1650]_ , \new_[1651]_ , \new_[1652]_ ,
    \new_[1653]_ , \new_[1654]_ , \new_[1655]_ , \new_[1656]_ ,
    \new_[1657]_ , \new_[1658]_ , \new_[1659]_ , \new_[1660]_ ,
    \new_[1661]_ , \new_[1662]_ , \new_[1663]_ , \new_[1664]_ ,
    \new_[1665]_ , \new_[1666]_ , \new_[1667]_ , \new_[1668]_ ,
    \new_[1669]_ , \new_[1670]_ , \new_[1671]_ , \new_[1672]_ ,
    \new_[1673]_ , \new_[1674]_ , \new_[1675]_ , \new_[1676]_ ,
    \new_[1677]_ , \new_[1678]_ , \new_[1679]_ , \new_[1680]_ ,
    \new_[1681]_ , \new_[1682]_ , \new_[1683]_ , \new_[1684]_ ,
    \new_[1685]_ , \new_[1686]_ , \new_[1687]_ , \new_[1688]_ ,
    \new_[1689]_ , \new_[1690]_ , \new_[1691]_ , \new_[1692]_ ,
    \new_[1693]_ , \new_[1694]_ , \new_[1695]_ , \new_[1696]_ ,
    \new_[1697]_ , \new_[1698]_ , \new_[1699]_ , \new_[1700]_ ,
    \new_[1701]_ , \new_[1702]_ , \new_[1703]_ , \new_[1704]_ ,
    \new_[1705]_ , \new_[1706]_ , \new_[1707]_ , \new_[1708]_ ,
    \new_[1709]_ , \new_[1710]_ , \new_[1711]_ , \new_[1712]_ ,
    \new_[1713]_ , \new_[1714]_ , \new_[1715]_ , \new_[1716]_ ,
    \new_[1717]_ , \new_[1718]_ , \new_[1719]_ , \new_[1720]_ ,
    \new_[1721]_ , \new_[1722]_ , \new_[1723]_ , \new_[1724]_ ,
    \new_[1725]_ , \new_[1726]_ , \new_[1727]_ , \new_[1728]_ ,
    \new_[1729]_ , \new_[1730]_ , \new_[1731]_ , \new_[1732]_ ,
    \new_[1733]_ , \new_[1734]_ , \new_[1735]_ , \new_[1736]_ ,
    \new_[1737]_ , \new_[1738]_ , \new_[1739]_ , \new_[1740]_ ,
    \new_[1741]_ , \new_[1742]_ , \new_[1743]_ , \new_[1744]_ ,
    \new_[1745]_ , \new_[1746]_ , \new_[1747]_ , \new_[1748]_ ,
    \new_[1749]_ , \new_[1750]_ , \new_[1751]_ , \new_[1752]_ ,
    \new_[1753]_ , \new_[1754]_ , \new_[1755]_ , \new_[1756]_ ,
    \new_[1757]_ , \new_[1758]_ , \new_[1759]_ , \new_[1760]_ ,
    \new_[1761]_ , \new_[1762]_ , \new_[1763]_ , \new_[1764]_ ,
    \new_[1765]_ , \new_[1766]_ , \new_[1767]_ , \new_[1768]_ ,
    \new_[1769]_ , \new_[1770]_ , \new_[1771]_ , \new_[1772]_ ,
    \new_[1773]_ , \new_[1774]_ , \new_[1775]_ , \new_[1776]_ ,
    \new_[1777]_ , \new_[1778]_ , \new_[1779]_ , \new_[1780]_ ,
    \new_[1781]_ , \new_[1782]_ , \new_[1783]_ , \new_[1784]_ ,
    \new_[1785]_ , \new_[1786]_ , \new_[1787]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1791]_ , \new_[1792]_ ,
    \new_[1793]_ , \new_[1794]_ , \new_[1795]_ , \new_[1796]_ ,
    \new_[1797]_ , \new_[1798]_ , \new_[1799]_ , \new_[1800]_ ,
    \new_[1801]_ , \new_[1802]_ , \new_[1803]_ , \new_[1804]_ ,
    \new_[1805]_ , \new_[1806]_ , \new_[1807]_ , \new_[1808]_ ,
    \new_[1809]_ , \new_[1810]_ , \new_[1811]_ , \new_[1812]_ ,
    \new_[1813]_ , \new_[1814]_ , \new_[1815]_ , \new_[1816]_ ,
    \new_[1817]_ , \new_[1818]_ , \new_[1819]_ , \new_[1820]_ ,
    \new_[1821]_ , \new_[1822]_ , \new_[1823]_ , \new_[1824]_ ,
    \new_[1825]_ , \new_[1826]_ , \new_[1827]_ , \new_[1828]_ ,
    \new_[1829]_ , \new_[1830]_ , \new_[1831]_ , \new_[1832]_ ,
    \new_[1833]_ , \new_[1834]_ , \new_[1835]_ , \new_[1836]_ ,
    \new_[1837]_ , \new_[1838]_ , \new_[1839]_ , \new_[1840]_ ,
    \new_[1841]_ , \new_[1842]_ , \new_[1843]_ , \new_[1844]_ ,
    \new_[1845]_ , \new_[1846]_ , \new_[1847]_ , \new_[1848]_ ,
    \new_[1849]_ , \new_[1850]_ , \new_[1851]_ , \new_[1852]_ ,
    \new_[1853]_ , \new_[1854]_ , \new_[1855]_ , \new_[1856]_ ,
    \new_[1857]_ , \new_[1858]_ , \new_[1859]_ , \new_[1860]_ ,
    \new_[1861]_ , \new_[1862]_ , \new_[1863]_ , \new_[1864]_ ,
    \new_[1865]_ , \new_[1866]_ , \new_[1867]_ , \new_[1868]_ ,
    \new_[1869]_ , \new_[1870]_ , \new_[1871]_ , \new_[1872]_ ,
    \new_[1873]_ , \new_[1874]_ , \new_[1875]_ , \new_[1876]_ ,
    \new_[1877]_ , \new_[1878]_ , \new_[1879]_ , \new_[1880]_ ,
    \new_[1881]_ , \new_[1882]_ , \new_[1883]_ , \new_[1884]_ ,
    \new_[1885]_ , \new_[1886]_ , \new_[1887]_ , \new_[1888]_ ,
    \new_[1889]_ , \new_[1890]_ , \new_[1891]_ , \new_[1892]_ ,
    \new_[1893]_ , \new_[1894]_ , \new_[1895]_ , \new_[1896]_ ,
    \new_[1897]_ , \new_[1898]_ , \new_[1899]_ , \new_[1900]_ ,
    \new_[1901]_ , \new_[1902]_ , \new_[1903]_ , \new_[1904]_ ,
    \new_[1905]_ , \new_[1906]_ , \new_[1907]_ , \new_[1908]_ ,
    \new_[1909]_ , \new_[1910]_ , \new_[1911]_ , \new_[1912]_ ,
    \new_[1913]_ , \new_[1914]_ , \new_[1915]_ , \new_[1916]_ ,
    \new_[1917]_ , \new_[1918]_ , \new_[1919]_ , \new_[1920]_ ,
    \new_[1921]_ , \new_[1922]_ , \new_[1923]_ , \new_[1924]_ ,
    \new_[1925]_ , \new_[1926]_ , \new_[1927]_ , \new_[1928]_ ,
    \new_[1929]_ , \new_[1930]_ , \new_[1931]_ , \new_[1932]_ ,
    \new_[1933]_ , \new_[1934]_ , \new_[1935]_ , \new_[1936]_ ,
    \new_[1937]_ , \new_[1938]_ , \new_[1939]_ , \new_[1940]_ ,
    \new_[1941]_ , \new_[1942]_ , \new_[1943]_ , \new_[1944]_ ,
    \new_[1945]_ , \new_[1946]_ , \new_[1947]_ , \new_[1948]_ ,
    \new_[1949]_ , \new_[1950]_ , \new_[1951]_ , \new_[1952]_ ,
    \new_[1953]_ , \new_[1954]_ , \new_[1955]_ , \new_[1956]_ ,
    \new_[1957]_ , \new_[1958]_ , \new_[1959]_ , \new_[1960]_ ,
    \new_[1961]_ , \new_[1962]_ , \new_[1963]_ , \new_[1964]_ ,
    \new_[1965]_ , \new_[1966]_ , \new_[1967]_ , \new_[1968]_ ,
    \new_[1969]_ , \new_[1970]_ , \new_[1971]_ , \new_[1972]_ ,
    \new_[1973]_ , \new_[1974]_ , \new_[1975]_ , \new_[1976]_ ,
    \new_[1977]_ , \new_[1978]_ , \new_[1979]_ , \new_[1980]_ ,
    \new_[1981]_ , \new_[1982]_ , \new_[1983]_ , \new_[1984]_ ,
    \new_[1985]_ , \new_[1986]_ , \new_[1987]_ , \new_[1988]_ ,
    \new_[1989]_ , \new_[1990]_ , \new_[1991]_ , \new_[1992]_ ,
    \new_[1993]_ , \new_[1994]_ , \new_[1995]_ , \new_[1996]_ ,
    \new_[1997]_ , \new_[1998]_ , \new_[1999]_ , \new_[2000]_ ,
    \new_[2001]_ , \new_[2002]_ , \new_[2003]_ , \new_[2004]_ ,
    \new_[2005]_ , \new_[2006]_ , \new_[2007]_ , \new_[2008]_ ,
    \new_[2009]_ , \new_[2010]_ , \new_[2011]_ , \new_[2012]_ ,
    \new_[2013]_ , \new_[2014]_ , \new_[2015]_ , \new_[2016]_ ,
    \new_[2017]_ , \new_[2018]_ , \new_[2019]_ , \new_[2020]_ ,
    \new_[2021]_ , \new_[2022]_ , \new_[2023]_ , \new_[2024]_ ,
    \new_[2025]_ , \new_[2026]_ , \new_[2027]_ , \new_[2028]_ ,
    \new_[2029]_ , \new_[2030]_ , \new_[2031]_ , \new_[2032]_ ,
    \new_[2033]_ , \new_[2034]_ , \new_[2035]_ , \new_[2036]_ ,
    \new_[2037]_ , \new_[2038]_ , \new_[2039]_ , \new_[2040]_ ,
    \new_[2041]_ , \new_[2042]_ , \new_[2043]_ , \new_[2044]_ ,
    \new_[2045]_ , \new_[2046]_ , \new_[2047]_ , \new_[2048]_ ,
    \new_[2049]_ , \new_[2050]_ , \new_[2051]_ , \new_[2052]_ ,
    \new_[2053]_ , \new_[2054]_ , \new_[2055]_ , \new_[2056]_ ,
    \new_[2057]_ , \new_[2058]_ , \new_[2059]_ , \new_[2060]_ ,
    \new_[2061]_ , \new_[2062]_ , \new_[2063]_ , \new_[2064]_ ,
    \new_[2065]_ , \new_[2066]_ , \new_[2067]_ , \new_[2068]_ ,
    \new_[2069]_ , \new_[2070]_ , \new_[2071]_ , \new_[2072]_ ,
    \new_[2073]_ , \new_[2074]_ , \new_[2075]_ , \new_[2076]_ ,
    \new_[2077]_ , \new_[2078]_ , \new_[2079]_ , \new_[2080]_ ,
    \new_[2081]_ , \new_[2082]_ , \new_[2083]_ , \new_[2084]_ ,
    \new_[2085]_ , \new_[2086]_ , \new_[2087]_ , \new_[2088]_ ,
    \new_[2089]_ , \new_[2090]_ , \new_[2091]_ , \new_[2092]_ ,
    \new_[2093]_ , \new_[2094]_ , \new_[2095]_ , \new_[2096]_ ,
    \new_[2097]_ , \new_[2098]_ , \new_[2099]_ , \new_[2100]_ ,
    \new_[2101]_ , \new_[2102]_ , \new_[2103]_ , \new_[2104]_ ,
    \new_[2105]_ , \new_[2106]_ , \new_[2107]_ , \new_[2108]_ ,
    \new_[2109]_ , \new_[2110]_ , \new_[2111]_ , \new_[2112]_ ,
    \new_[2113]_ , \new_[2114]_ , \new_[2115]_ , \new_[2116]_ ,
    \new_[2117]_ , \new_[2118]_ , \new_[2119]_ , \new_[2120]_ ,
    \new_[2121]_ , \new_[2122]_ , \new_[2123]_ , \new_[2124]_ ,
    \new_[2125]_ , \new_[2126]_ , \new_[2127]_ , \new_[2128]_ ,
    \new_[2129]_ , \new_[2130]_ , \new_[2131]_ , \new_[2132]_ ,
    \new_[2133]_ , \new_[2134]_ , \new_[2135]_ , \new_[2136]_ ,
    \new_[2137]_ , \new_[2138]_ , \new_[2139]_ , \new_[2140]_ ,
    \new_[2141]_ , \new_[2142]_ , \new_[2143]_ , \new_[2144]_ ,
    \new_[2145]_ , \new_[2146]_ , \new_[2147]_ , \new_[2148]_ ,
    \new_[2149]_ , \new_[2150]_ , \new_[2151]_ , \new_[2152]_ ,
    \new_[2153]_ , \new_[2154]_ , \new_[2155]_ , \new_[2156]_ ,
    \new_[2157]_ , \new_[2158]_ , \new_[2159]_ , \new_[2160]_ ,
    \new_[2161]_ , \new_[2162]_ , \new_[2163]_ , \new_[2164]_ ,
    \new_[2165]_ , \new_[2166]_ , \new_[2167]_ , \new_[2168]_ ,
    \new_[2169]_ , \new_[2170]_ , \new_[2171]_ , \new_[2172]_ ,
    \new_[2173]_ , \new_[2174]_ , \new_[2175]_ , \new_[2176]_ ,
    \new_[2177]_ , \new_[2178]_ , \new_[2179]_ , \new_[2180]_ ,
    \new_[2181]_ , \new_[2182]_ , \new_[2183]_ , \new_[2184]_ ,
    \new_[2185]_ , \new_[2186]_ , \new_[2187]_ , \new_[2188]_ ,
    \new_[2189]_ , \new_[2190]_ , \new_[2193]_ , \new_[2196]_ ,
    \new_[2197]_ , \new_[2200]_ , \new_[2203]_ , \new_[2204]_ ,
    \new_[2205]_ , \new_[2208]_ , \new_[2211]_ , \new_[2212]_ ,
    \new_[2215]_ , \new_[2219]_ , \new_[2220]_ , \new_[2221]_ ,
    \new_[2222]_ , \new_[2223]_ , \new_[2226]_ , \new_[2229]_ ,
    \new_[2230]_ , \new_[2233]_ , \new_[2236]_ , \new_[2237]_ ,
    \new_[2238]_ , \new_[2241]_ , \new_[2244]_ , \new_[2245]_ ,
    \new_[2248]_ , \new_[2252]_ , \new_[2253]_ , \new_[2254]_ ,
    \new_[2255]_ , \new_[2256]_ , \new_[2257]_ , \new_[2260]_ ,
    \new_[2263]_ , \new_[2264]_ , \new_[2267]_ , \new_[2270]_ ,
    \new_[2271]_ , \new_[2272]_ , \new_[2275]_ , \new_[2278]_ ,
    \new_[2279]_ , \new_[2282]_ , \new_[2286]_ , \new_[2287]_ ,
    \new_[2288]_ , \new_[2289]_ , \new_[2290]_ , \new_[2293]_ ,
    \new_[2296]_ , \new_[2297]_ , \new_[2300]_ , \new_[2303]_ ,
    \new_[2304]_ , \new_[2305]_ , \new_[2308]_ , \new_[2311]_ ,
    \new_[2312]_ , \new_[2315]_ , \new_[2319]_ , \new_[2320]_ ,
    \new_[2321]_ , \new_[2322]_ , \new_[2323]_ , \new_[2324]_ ,
    \new_[2325]_ , \new_[2328]_ , \new_[2331]_ , \new_[2332]_ ,
    \new_[2335]_ , \new_[2338]_ , \new_[2339]_ , \new_[2340]_ ,
    \new_[2343]_ , \new_[2346]_ , \new_[2347]_ , \new_[2350]_ ,
    \new_[2354]_ , \new_[2355]_ , \new_[2356]_ , \new_[2357]_ ,
    \new_[2358]_ , \new_[2361]_ , \new_[2364]_ , \new_[2365]_ ,
    \new_[2368]_ , \new_[2371]_ , \new_[2372]_ , \new_[2373]_ ,
    \new_[2376]_ , \new_[2379]_ , \new_[2380]_ , \new_[2383]_ ,
    \new_[2387]_ , \new_[2388]_ , \new_[2389]_ , \new_[2390]_ ,
    \new_[2391]_ , \new_[2392]_ , \new_[2395]_ , \new_[2398]_ ,
    \new_[2399]_ , \new_[2402]_ , \new_[2405]_ , \new_[2406]_ ,
    \new_[2407]_ , \new_[2410]_ , \new_[2413]_ , \new_[2414]_ ,
    \new_[2417]_ , \new_[2421]_ , \new_[2422]_ , \new_[2423]_ ,
    \new_[2424]_ , \new_[2425]_ , \new_[2428]_ , \new_[2431]_ ,
    \new_[2432]_ , \new_[2435]_ , \new_[2438]_ , \new_[2439]_ ,
    \new_[2440]_ , \new_[2443]_ , \new_[2446]_ , \new_[2447]_ ,
    \new_[2450]_ , \new_[2454]_ , \new_[2455]_ , \new_[2456]_ ,
    \new_[2457]_ , \new_[2458]_ , \new_[2459]_ , \new_[2460]_ ,
    \new_[2461]_ , \new_[2464]_ , \new_[2467]_ , \new_[2468]_ ,
    \new_[2471]_ , \new_[2474]_ , \new_[2475]_ , \new_[2476]_ ,
    \new_[2479]_ , \new_[2482]_ , \new_[2483]_ , \new_[2486]_ ,
    \new_[2490]_ , \new_[2491]_ , \new_[2492]_ , \new_[2493]_ ,
    \new_[2494]_ , \new_[2497]_ , \new_[2500]_ , \new_[2501]_ ,
    \new_[2504]_ , \new_[2507]_ , \new_[2508]_ , \new_[2509]_ ,
    \new_[2512]_ , \new_[2515]_ , \new_[2516]_ , \new_[2519]_ ,
    \new_[2523]_ , \new_[2524]_ , \new_[2525]_ , \new_[2526]_ ,
    \new_[2527]_ , \new_[2528]_ , \new_[2531]_ , \new_[2534]_ ,
    \new_[2535]_ , \new_[2538]_ , \new_[2541]_ , \new_[2542]_ ,
    \new_[2543]_ , \new_[2546]_ , \new_[2549]_ , \new_[2550]_ ,
    \new_[2553]_ , \new_[2557]_ , \new_[2558]_ , \new_[2559]_ ,
    \new_[2560]_ , \new_[2561]_ , \new_[2564]_ , \new_[2567]_ ,
    \new_[2568]_ , \new_[2571]_ , \new_[2574]_ , \new_[2575]_ ,
    \new_[2576]_ , \new_[2579]_ , \new_[2582]_ , \new_[2583]_ ,
    \new_[2586]_ , \new_[2590]_ , \new_[2591]_ , \new_[2592]_ ,
    \new_[2593]_ , \new_[2594]_ , \new_[2595]_ , \new_[2596]_ ,
    \new_[2599]_ , \new_[2602]_ , \new_[2603]_ , \new_[2606]_ ,
    \new_[2609]_ , \new_[2610]_ , \new_[2611]_ , \new_[2614]_ ,
    \new_[2617]_ , \new_[2618]_ , \new_[2621]_ , \new_[2625]_ ,
    \new_[2626]_ , \new_[2627]_ , \new_[2628]_ , \new_[2629]_ ,
    \new_[2632]_ , \new_[2635]_ , \new_[2636]_ , \new_[2639]_ ,
    \new_[2642]_ , \new_[2643]_ , \new_[2644]_ , \new_[2647]_ ,
    \new_[2650]_ , \new_[2651]_ , \new_[2654]_ , \new_[2658]_ ,
    \new_[2659]_ , \new_[2660]_ , \new_[2661]_ , \new_[2662]_ ,
    \new_[2663]_ , \new_[2666]_ , \new_[2669]_ , \new_[2670]_ ,
    \new_[2673]_ , \new_[2676]_ , \new_[2677]_ , \new_[2678]_ ,
    \new_[2681]_ , \new_[2684]_ , \new_[2685]_ , \new_[2688]_ ,
    \new_[2692]_ , \new_[2693]_ , \new_[2694]_ , \new_[2695]_ ,
    \new_[2696]_ , \new_[2699]_ , \new_[2702]_ , \new_[2703]_ ,
    \new_[2706]_ , \new_[2710]_ , \new_[2711]_ , \new_[2712]_ ,
    \new_[2713]_ , \new_[2716]_ , \new_[2719]_ , \new_[2720]_ ,
    \new_[2723]_ , \new_[2727]_ , \new_[2728]_ , \new_[2729]_ ,
    \new_[2730]_ , \new_[2731]_ , \new_[2732]_ , \new_[2733]_ ,
    \new_[2734]_ , \new_[2735]_ , \new_[2738]_ , \new_[2741]_ ,
    \new_[2742]_ , \new_[2745]_ , \new_[2748]_ , \new_[2749]_ ,
    \new_[2750]_ , \new_[2753]_ , \new_[2756]_ , \new_[2757]_ ,
    \new_[2760]_ , \new_[2764]_ , \new_[2765]_ , \new_[2766]_ ,
    \new_[2767]_ , \new_[2768]_ , \new_[2771]_ , \new_[2774]_ ,
    \new_[2775]_ , \new_[2778]_ , \new_[2781]_ , \new_[2782]_ ,
    \new_[2783]_ , \new_[2786]_ , \new_[2789]_ , \new_[2790]_ ,
    \new_[2793]_ , \new_[2797]_ , \new_[2798]_ , \new_[2799]_ ,
    \new_[2800]_ , \new_[2801]_ , \new_[2802]_ , \new_[2805]_ ,
    \new_[2808]_ , \new_[2809]_ , \new_[2812]_ , \new_[2815]_ ,
    \new_[2816]_ , \new_[2817]_ , \new_[2820]_ , \new_[2823]_ ,
    \new_[2824]_ , \new_[2827]_ , \new_[2831]_ , \new_[2832]_ ,
    \new_[2833]_ , \new_[2834]_ , \new_[2835]_ , \new_[2838]_ ,
    \new_[2841]_ , \new_[2842]_ , \new_[2845]_ , \new_[2848]_ ,
    \new_[2849]_ , \new_[2850]_ , \new_[2853]_ , \new_[2856]_ ,
    \new_[2857]_ , \new_[2860]_ , \new_[2864]_ , \new_[2865]_ ,
    \new_[2866]_ , \new_[2867]_ , \new_[2868]_ , \new_[2869]_ ,
    \new_[2870]_ , \new_[2873]_ , \new_[2876]_ , \new_[2877]_ ,
    \new_[2880]_ , \new_[2883]_ , \new_[2884]_ , \new_[2885]_ ,
    \new_[2888]_ , \new_[2891]_ , \new_[2892]_ , \new_[2895]_ ,
    \new_[2899]_ , \new_[2900]_ , \new_[2901]_ , \new_[2902]_ ,
    \new_[2903]_ , \new_[2906]_ , \new_[2909]_ , \new_[2910]_ ,
    \new_[2913]_ , \new_[2916]_ , \new_[2917]_ , \new_[2918]_ ,
    \new_[2921]_ , \new_[2924]_ , \new_[2925]_ , \new_[2928]_ ,
    \new_[2932]_ , \new_[2933]_ , \new_[2934]_ , \new_[2935]_ ,
    \new_[2936]_ , \new_[2937]_ , \new_[2940]_ , \new_[2943]_ ,
    \new_[2944]_ , \new_[2947]_ , \new_[2950]_ , \new_[2951]_ ,
    \new_[2952]_ , \new_[2955]_ , \new_[2958]_ , \new_[2959]_ ,
    \new_[2962]_ , \new_[2966]_ , \new_[2967]_ , \new_[2968]_ ,
    \new_[2969]_ , \new_[2970]_ , \new_[2973]_ , \new_[2976]_ ,
    \new_[2977]_ , \new_[2980]_ , \new_[2984]_ , \new_[2985]_ ,
    \new_[2986]_ , \new_[2987]_ , \new_[2990]_ , \new_[2993]_ ,
    \new_[2994]_ , \new_[2997]_ , \new_[3001]_ , \new_[3002]_ ,
    \new_[3003]_ , \new_[3004]_ , \new_[3005]_ , \new_[3006]_ ,
    \new_[3007]_ , \new_[3008]_ , \new_[3011]_ , \new_[3014]_ ,
    \new_[3015]_ , \new_[3018]_ , \new_[3021]_ , \new_[3022]_ ,
    \new_[3023]_ , \new_[3026]_ , \new_[3029]_ , \new_[3030]_ ,
    \new_[3033]_ , \new_[3037]_ , \new_[3038]_ , \new_[3039]_ ,
    \new_[3040]_ , \new_[3041]_ , \new_[3044]_ , \new_[3047]_ ,
    \new_[3048]_ , \new_[3051]_ , \new_[3054]_ , \new_[3055]_ ,
    \new_[3056]_ , \new_[3059]_ , \new_[3062]_ , \new_[3063]_ ,
    \new_[3066]_ , \new_[3070]_ , \new_[3071]_ , \new_[3072]_ ,
    \new_[3073]_ , \new_[3074]_ , \new_[3075]_ , \new_[3078]_ ,
    \new_[3081]_ , \new_[3082]_ , \new_[3085]_ , \new_[3088]_ ,
    \new_[3089]_ , \new_[3090]_ , \new_[3093]_ , \new_[3096]_ ,
    \new_[3097]_ , \new_[3100]_ , \new_[3104]_ , \new_[3105]_ ,
    \new_[3106]_ , \new_[3107]_ , \new_[3108]_ , \new_[3111]_ ,
    \new_[3114]_ , \new_[3115]_ , \new_[3118]_ , \new_[3121]_ ,
    \new_[3122]_ , \new_[3123]_ , \new_[3126]_ , \new_[3129]_ ,
    \new_[3130]_ , \new_[3133]_ , \new_[3137]_ , \new_[3138]_ ,
    \new_[3139]_ , \new_[3140]_ , \new_[3141]_ , \new_[3142]_ ,
    \new_[3143]_ , \new_[3146]_ , \new_[3149]_ , \new_[3150]_ ,
    \new_[3153]_ , \new_[3156]_ , \new_[3157]_ , \new_[3158]_ ,
    \new_[3161]_ , \new_[3164]_ , \new_[3165]_ , \new_[3168]_ ,
    \new_[3172]_ , \new_[3173]_ , \new_[3174]_ , \new_[3175]_ ,
    \new_[3176]_ , \new_[3179]_ , \new_[3182]_ , \new_[3183]_ ,
    \new_[3186]_ , \new_[3189]_ , \new_[3190]_ , \new_[3191]_ ,
    \new_[3194]_ , \new_[3197]_ , \new_[3198]_ , \new_[3201]_ ,
    \new_[3205]_ , \new_[3206]_ , \new_[3207]_ , \new_[3208]_ ,
    \new_[3209]_ , \new_[3210]_ , \new_[3213]_ , \new_[3216]_ ,
    \new_[3217]_ , \new_[3220]_ , \new_[3223]_ , \new_[3224]_ ,
    \new_[3225]_ , \new_[3228]_ , \new_[3231]_ , \new_[3232]_ ,
    \new_[3235]_ , \new_[3239]_ , \new_[3240]_ , \new_[3241]_ ,
    \new_[3242]_ , \new_[3243]_ , \new_[3246]_ , \new_[3249]_ ,
    \new_[3250]_ , \new_[3253]_ , \new_[3257]_ , \new_[3258]_ ,
    \new_[3259]_ , \new_[3260]_ , \new_[3263]_ , \new_[3266]_ ,
    \new_[3267]_ , \new_[3270]_ , \new_[3274]_ , \new_[3275]_ ,
    \new_[3276]_ , \new_[3277]_ , \new_[3278]_ , \new_[3279]_ ,
    \new_[3280]_ , \new_[3281]_ , \new_[3282]_ , \new_[3283]_ ,
    \new_[3286]_ , \new_[3289]_ , \new_[3290]_ , \new_[3293]_ ,
    \new_[3296]_ , \new_[3297]_ , \new_[3298]_ , \new_[3301]_ ,
    \new_[3304]_ , \new_[3305]_ , \new_[3308]_ , \new_[3312]_ ,
    \new_[3313]_ , \new_[3314]_ , \new_[3315]_ , \new_[3316]_ ,
    \new_[3319]_ , \new_[3322]_ , \new_[3323]_ , \new_[3326]_ ,
    \new_[3329]_ , \new_[3330]_ , \new_[3331]_ , \new_[3334]_ ,
    \new_[3337]_ , \new_[3338]_ , \new_[3341]_ , \new_[3345]_ ,
    \new_[3346]_ , \new_[3347]_ , \new_[3348]_ , \new_[3349]_ ,
    \new_[3350]_ , \new_[3353]_ , \new_[3356]_ , \new_[3357]_ ,
    \new_[3360]_ , \new_[3363]_ , \new_[3364]_ , \new_[3365]_ ,
    \new_[3368]_ , \new_[3371]_ , \new_[3372]_ , \new_[3375]_ ,
    \new_[3379]_ , \new_[3380]_ , \new_[3381]_ , \new_[3382]_ ,
    \new_[3383]_ , \new_[3386]_ , \new_[3389]_ , \new_[3390]_ ,
    \new_[3393]_ , \new_[3396]_ , \new_[3397]_ , \new_[3398]_ ,
    \new_[3401]_ , \new_[3404]_ , \new_[3405]_ , \new_[3408]_ ,
    \new_[3412]_ , \new_[3413]_ , \new_[3414]_ , \new_[3415]_ ,
    \new_[3416]_ , \new_[3417]_ , \new_[3418]_ , \new_[3421]_ ,
    \new_[3424]_ , \new_[3425]_ , \new_[3428]_ , \new_[3431]_ ,
    \new_[3432]_ , \new_[3433]_ , \new_[3436]_ , \new_[3439]_ ,
    \new_[3440]_ , \new_[3443]_ , \new_[3447]_ , \new_[3448]_ ,
    \new_[3449]_ , \new_[3450]_ , \new_[3451]_ , \new_[3454]_ ,
    \new_[3457]_ , \new_[3458]_ , \new_[3461]_ , \new_[3464]_ ,
    \new_[3465]_ , \new_[3466]_ , \new_[3469]_ , \new_[3472]_ ,
    \new_[3473]_ , \new_[3476]_ , \new_[3480]_ , \new_[3481]_ ,
    \new_[3482]_ , \new_[3483]_ , \new_[3484]_ , \new_[3485]_ ,
    \new_[3488]_ , \new_[3491]_ , \new_[3492]_ , \new_[3495]_ ,
    \new_[3498]_ , \new_[3499]_ , \new_[3500]_ , \new_[3503]_ ,
    \new_[3506]_ , \new_[3507]_ , \new_[3510]_ , \new_[3514]_ ,
    \new_[3515]_ , \new_[3516]_ , \new_[3517]_ , \new_[3518]_ ,
    \new_[3521]_ , \new_[3524]_ , \new_[3525]_ , \new_[3528]_ ,
    \new_[3532]_ , \new_[3533]_ , \new_[3534]_ , \new_[3535]_ ,
    \new_[3538]_ , \new_[3541]_ , \new_[3542]_ , \new_[3545]_ ,
    \new_[3549]_ , \new_[3550]_ , \new_[3551]_ , \new_[3552]_ ,
    \new_[3553]_ , \new_[3554]_ , \new_[3555]_ , \new_[3556]_ ,
    \new_[3559]_ , \new_[3562]_ , \new_[3563]_ , \new_[3566]_ ,
    \new_[3569]_ , \new_[3570]_ , \new_[3571]_ , \new_[3574]_ ,
    \new_[3577]_ , \new_[3578]_ , \new_[3581]_ , \new_[3585]_ ,
    \new_[3586]_ , \new_[3587]_ , \new_[3588]_ , \new_[3589]_ ,
    \new_[3592]_ , \new_[3595]_ , \new_[3596]_ , \new_[3599]_ ,
    \new_[3602]_ , \new_[3603]_ , \new_[3604]_ , \new_[3607]_ ,
    \new_[3610]_ , \new_[3611]_ , \new_[3614]_ , \new_[3618]_ ,
    \new_[3619]_ , \new_[3620]_ , \new_[3621]_ , \new_[3622]_ ,
    \new_[3623]_ , \new_[3626]_ , \new_[3629]_ , \new_[3630]_ ,
    \new_[3633]_ , \new_[3636]_ , \new_[3637]_ , \new_[3638]_ ,
    \new_[3641]_ , \new_[3644]_ , \new_[3645]_ , \new_[3648]_ ,
    \new_[3652]_ , \new_[3653]_ , \new_[3654]_ , \new_[3655]_ ,
    \new_[3656]_ , \new_[3659]_ , \new_[3662]_ , \new_[3663]_ ,
    \new_[3666]_ , \new_[3669]_ , \new_[3670]_ , \new_[3671]_ ,
    \new_[3674]_ , \new_[3677]_ , \new_[3678]_ , \new_[3681]_ ,
    \new_[3685]_ , \new_[3686]_ , \new_[3687]_ , \new_[3688]_ ,
    \new_[3689]_ , \new_[3690]_ , \new_[3691]_ , \new_[3694]_ ,
    \new_[3697]_ , \new_[3698]_ , \new_[3701]_ , \new_[3704]_ ,
    \new_[3705]_ , \new_[3706]_ , \new_[3709]_ , \new_[3712]_ ,
    \new_[3713]_ , \new_[3716]_ , \new_[3720]_ , \new_[3721]_ ,
    \new_[3722]_ , \new_[3723]_ , \new_[3724]_ , \new_[3727]_ ,
    \new_[3730]_ , \new_[3731]_ , \new_[3734]_ , \new_[3737]_ ,
    \new_[3738]_ , \new_[3739]_ , \new_[3742]_ , \new_[3745]_ ,
    \new_[3746]_ , \new_[3749]_ , \new_[3753]_ , \new_[3754]_ ,
    \new_[3755]_ , \new_[3756]_ , \new_[3757]_ , \new_[3758]_ ,
    \new_[3761]_ , \new_[3764]_ , \new_[3765]_ , \new_[3768]_ ,
    \new_[3771]_ , \new_[3772]_ , \new_[3773]_ , \new_[3776]_ ,
    \new_[3779]_ , \new_[3780]_ , \new_[3783]_ , \new_[3787]_ ,
    \new_[3788]_ , \new_[3789]_ , \new_[3790]_ , \new_[3791]_ ,
    \new_[3794]_ , \new_[3797]_ , \new_[3798]_ , \new_[3801]_ ,
    \new_[3805]_ , \new_[3806]_ , \new_[3807]_ , \new_[3808]_ ,
    \new_[3811]_ , \new_[3814]_ , \new_[3815]_ , \new_[3818]_ ,
    \new_[3822]_ , \new_[3823]_ , \new_[3824]_ , \new_[3825]_ ,
    \new_[3826]_ , \new_[3827]_ , \new_[3828]_ , \new_[3829]_ ,
    \new_[3830]_ , \new_[3833]_ , \new_[3836]_ , \new_[3837]_ ,
    \new_[3840]_ , \new_[3843]_ , \new_[3844]_ , \new_[3845]_ ,
    \new_[3848]_ , \new_[3851]_ , \new_[3852]_ , \new_[3855]_ ,
    \new_[3859]_ , \new_[3860]_ , \new_[3861]_ , \new_[3862]_ ,
    \new_[3863]_ , \new_[3866]_ , \new_[3869]_ , \new_[3870]_ ,
    \new_[3873]_ , \new_[3876]_ , \new_[3877]_ , \new_[3878]_ ,
    \new_[3881]_ , \new_[3884]_ , \new_[3885]_ , \new_[3888]_ ,
    \new_[3892]_ , \new_[3893]_ , \new_[3894]_ , \new_[3895]_ ,
    \new_[3896]_ , \new_[3897]_ , \new_[3900]_ , \new_[3903]_ ,
    \new_[3904]_ , \new_[3907]_ , \new_[3910]_ , \new_[3911]_ ,
    \new_[3912]_ , \new_[3915]_ , \new_[3918]_ , \new_[3919]_ ,
    \new_[3922]_ , \new_[3926]_ , \new_[3927]_ , \new_[3928]_ ,
    \new_[3929]_ , \new_[3930]_ , \new_[3933]_ , \new_[3936]_ ,
    \new_[3937]_ , \new_[3940]_ , \new_[3943]_ , \new_[3944]_ ,
    \new_[3945]_ , \new_[3948]_ , \new_[3951]_ , \new_[3952]_ ,
    \new_[3955]_ , \new_[3959]_ , \new_[3960]_ , \new_[3961]_ ,
    \new_[3962]_ , \new_[3963]_ , \new_[3964]_ , \new_[3965]_ ,
    \new_[3968]_ , \new_[3971]_ , \new_[3972]_ , \new_[3975]_ ,
    \new_[3978]_ , \new_[3979]_ , \new_[3980]_ , \new_[3983]_ ,
    \new_[3986]_ , \new_[3987]_ , \new_[3990]_ , \new_[3994]_ ,
    \new_[3995]_ , \new_[3996]_ , \new_[3997]_ , \new_[3998]_ ,
    \new_[4001]_ , \new_[4004]_ , \new_[4005]_ , \new_[4008]_ ,
    \new_[4011]_ , \new_[4012]_ , \new_[4013]_ , \new_[4016]_ ,
    \new_[4019]_ , \new_[4020]_ , \new_[4023]_ , \new_[4027]_ ,
    \new_[4028]_ , \new_[4029]_ , \new_[4030]_ , \new_[4031]_ ,
    \new_[4032]_ , \new_[4035]_ , \new_[4038]_ , \new_[4039]_ ,
    \new_[4042]_ , \new_[4045]_ , \new_[4046]_ , \new_[4047]_ ,
    \new_[4050]_ , \new_[4053]_ , \new_[4054]_ , \new_[4057]_ ,
    \new_[4061]_ , \new_[4062]_ , \new_[4063]_ , \new_[4064]_ ,
    \new_[4065]_ , \new_[4068]_ , \new_[4071]_ , \new_[4072]_ ,
    \new_[4075]_ , \new_[4079]_ , \new_[4080]_ , \new_[4081]_ ,
    \new_[4082]_ , \new_[4085]_ , \new_[4088]_ , \new_[4089]_ ,
    \new_[4092]_ , \new_[4096]_ , \new_[4097]_ , \new_[4098]_ ,
    \new_[4099]_ , \new_[4100]_ , \new_[4101]_ , \new_[4102]_ ,
    \new_[4103]_ , \new_[4106]_ , \new_[4109]_ , \new_[4110]_ ,
    \new_[4113]_ , \new_[4116]_ , \new_[4117]_ , \new_[4118]_ ,
    \new_[4121]_ , \new_[4124]_ , \new_[4125]_ , \new_[4128]_ ,
    \new_[4132]_ , \new_[4133]_ , \new_[4134]_ , \new_[4135]_ ,
    \new_[4136]_ , \new_[4139]_ , \new_[4142]_ , \new_[4143]_ ,
    \new_[4146]_ , \new_[4149]_ , \new_[4150]_ , \new_[4151]_ ,
    \new_[4154]_ , \new_[4157]_ , \new_[4158]_ , \new_[4161]_ ,
    \new_[4165]_ , \new_[4166]_ , \new_[4167]_ , \new_[4168]_ ,
    \new_[4169]_ , \new_[4170]_ , \new_[4173]_ , \new_[4176]_ ,
    \new_[4177]_ , \new_[4180]_ , \new_[4183]_ , \new_[4184]_ ,
    \new_[4185]_ , \new_[4188]_ , \new_[4191]_ , \new_[4192]_ ,
    \new_[4195]_ , \new_[4199]_ , \new_[4200]_ , \new_[4201]_ ,
    \new_[4202]_ , \new_[4203]_ , \new_[4206]_ , \new_[4209]_ ,
    \new_[4210]_ , \new_[4213]_ , \new_[4216]_ , \new_[4217]_ ,
    \new_[4218]_ , \new_[4221]_ , \new_[4224]_ , \new_[4225]_ ,
    \new_[4228]_ , \new_[4232]_ , \new_[4233]_ , \new_[4234]_ ,
    \new_[4235]_ , \new_[4236]_ , \new_[4237]_ , \new_[4238]_ ,
    \new_[4241]_ , \new_[4244]_ , \new_[4245]_ , \new_[4248]_ ,
    \new_[4251]_ , \new_[4252]_ , \new_[4253]_ , \new_[4256]_ ,
    \new_[4259]_ , \new_[4260]_ , \new_[4263]_ , \new_[4267]_ ,
    \new_[4268]_ , \new_[4269]_ , \new_[4270]_ , \new_[4271]_ ,
    \new_[4274]_ , \new_[4277]_ , \new_[4278]_ , \new_[4281]_ ,
    \new_[4284]_ , \new_[4285]_ , \new_[4286]_ , \new_[4289]_ ,
    \new_[4292]_ , \new_[4293]_ , \new_[4296]_ , \new_[4300]_ ,
    \new_[4301]_ , \new_[4302]_ , \new_[4303]_ , \new_[4304]_ ,
    \new_[4305]_ , \new_[4308]_ , \new_[4311]_ , \new_[4312]_ ,
    \new_[4315]_ , \new_[4318]_ , \new_[4319]_ , \new_[4320]_ ,
    \new_[4323]_ , \new_[4326]_ , \new_[4327]_ , \new_[4330]_ ,
    \new_[4334]_ , \new_[4335]_ , \new_[4336]_ , \new_[4337]_ ,
    \new_[4338]_ , \new_[4341]_ , \new_[4344]_ , \new_[4345]_ ,
    \new_[4348]_ , \new_[4352]_ , \new_[4353]_ , \new_[4354]_ ,
    \new_[4355]_ , \new_[4358]_ , \new_[4361]_ , \new_[4362]_ ,
    \new_[4365]_ , \new_[4369]_ , \new_[4370]_ , \new_[4371]_ ,
    \new_[4372]_ , \new_[4373]_ , \new_[4374]_ , \new_[4375]_ ,
    \new_[4376]_ , \new_[4377]_ , \new_[4378]_ , \new_[4379]_ ,
    \new_[4382]_ , \new_[4385]_ , \new_[4386]_ , \new_[4389]_ ,
    \new_[4392]_ , \new_[4393]_ , \new_[4394]_ , \new_[4397]_ ,
    \new_[4400]_ , \new_[4401]_ , \new_[4404]_ , \new_[4408]_ ,
    \new_[4409]_ , \new_[4410]_ , \new_[4411]_ , \new_[4412]_ ,
    \new_[4415]_ , \new_[4418]_ , \new_[4419]_ , \new_[4422]_ ,
    \new_[4425]_ , \new_[4426]_ , \new_[4427]_ , \new_[4430]_ ,
    \new_[4433]_ , \new_[4434]_ , \new_[4437]_ , \new_[4441]_ ,
    \new_[4442]_ , \new_[4443]_ , \new_[4444]_ , \new_[4445]_ ,
    \new_[4446]_ , \new_[4449]_ , \new_[4452]_ , \new_[4453]_ ,
    \new_[4456]_ , \new_[4459]_ , \new_[4460]_ , \new_[4461]_ ,
    \new_[4464]_ , \new_[4467]_ , \new_[4468]_ , \new_[4471]_ ,
    \new_[4475]_ , \new_[4476]_ , \new_[4477]_ , \new_[4478]_ ,
    \new_[4479]_ , \new_[4482]_ , \new_[4485]_ , \new_[4486]_ ,
    \new_[4489]_ , \new_[4492]_ , \new_[4493]_ , \new_[4494]_ ,
    \new_[4497]_ , \new_[4500]_ , \new_[4501]_ , \new_[4504]_ ,
    \new_[4508]_ , \new_[4509]_ , \new_[4510]_ , \new_[4511]_ ,
    \new_[4512]_ , \new_[4513]_ , \new_[4514]_ , \new_[4517]_ ,
    \new_[4520]_ , \new_[4521]_ , \new_[4524]_ , \new_[4527]_ ,
    \new_[4528]_ , \new_[4529]_ , \new_[4532]_ , \new_[4535]_ ,
    \new_[4536]_ , \new_[4539]_ , \new_[4543]_ , \new_[4544]_ ,
    \new_[4545]_ , \new_[4546]_ , \new_[4547]_ , \new_[4550]_ ,
    \new_[4553]_ , \new_[4554]_ , \new_[4557]_ , \new_[4560]_ ,
    \new_[4561]_ , \new_[4562]_ , \new_[4565]_ , \new_[4568]_ ,
    \new_[4569]_ , \new_[4572]_ , \new_[4576]_ , \new_[4577]_ ,
    \new_[4578]_ , \new_[4579]_ , \new_[4580]_ , \new_[4581]_ ,
    \new_[4584]_ , \new_[4587]_ , \new_[4588]_ , \new_[4591]_ ,
    \new_[4594]_ , \new_[4595]_ , \new_[4596]_ , \new_[4599]_ ,
    \new_[4602]_ , \new_[4603]_ , \new_[4606]_ , \new_[4610]_ ,
    \new_[4611]_ , \new_[4612]_ , \new_[4613]_ , \new_[4614]_ ,
    \new_[4617]_ , \new_[4620]_ , \new_[4621]_ , \new_[4624]_ ,
    \new_[4627]_ , \new_[4628]_ , \new_[4629]_ , \new_[4632]_ ,
    \new_[4635]_ , \new_[4636]_ , \new_[4639]_ , \new_[4643]_ ,
    \new_[4644]_ , \new_[4645]_ , \new_[4646]_ , \new_[4647]_ ,
    \new_[4648]_ , \new_[4649]_ , \new_[4650]_ , \new_[4653]_ ,
    \new_[4656]_ , \new_[4657]_ , \new_[4660]_ , \new_[4663]_ ,
    \new_[4664]_ , \new_[4665]_ , \new_[4668]_ , \new_[4671]_ ,
    \new_[4672]_ , \new_[4675]_ , \new_[4679]_ , \new_[4680]_ ,
    \new_[4681]_ , \new_[4682]_ , \new_[4683]_ , \new_[4686]_ ,
    \new_[4689]_ , \new_[4690]_ , \new_[4693]_ , \new_[4696]_ ,
    \new_[4697]_ , \new_[4698]_ , \new_[4701]_ , \new_[4704]_ ,
    \new_[4705]_ , \new_[4708]_ , \new_[4712]_ , \new_[4713]_ ,
    \new_[4714]_ , \new_[4715]_ , \new_[4716]_ , \new_[4717]_ ,
    \new_[4720]_ , \new_[4723]_ , \new_[4724]_ , \new_[4727]_ ,
    \new_[4730]_ , \new_[4731]_ , \new_[4732]_ , \new_[4735]_ ,
    \new_[4738]_ , \new_[4739]_ , \new_[4742]_ , \new_[4746]_ ,
    \new_[4747]_ , \new_[4748]_ , \new_[4749]_ , \new_[4750]_ ,
    \new_[4753]_ , \new_[4756]_ , \new_[4757]_ , \new_[4760]_ ,
    \new_[4763]_ , \new_[4764]_ , \new_[4765]_ , \new_[4768]_ ,
    \new_[4771]_ , \new_[4772]_ , \new_[4775]_ , \new_[4779]_ ,
    \new_[4780]_ , \new_[4781]_ , \new_[4782]_ , \new_[4783]_ ,
    \new_[4784]_ , \new_[4785]_ , \new_[4788]_ , \new_[4791]_ ,
    \new_[4792]_ , \new_[4795]_ , \new_[4798]_ , \new_[4799]_ ,
    \new_[4800]_ , \new_[4803]_ , \new_[4806]_ , \new_[4807]_ ,
    \new_[4810]_ , \new_[4814]_ , \new_[4815]_ , \new_[4816]_ ,
    \new_[4817]_ , \new_[4818]_ , \new_[4821]_ , \new_[4824]_ ,
    \new_[4825]_ , \new_[4828]_ , \new_[4831]_ , \new_[4832]_ ,
    \new_[4833]_ , \new_[4836]_ , \new_[4839]_ , \new_[4840]_ ,
    \new_[4843]_ , \new_[4847]_ , \new_[4848]_ , \new_[4849]_ ,
    \new_[4850]_ , \new_[4851]_ , \new_[4852]_ , \new_[4855]_ ,
    \new_[4858]_ , \new_[4859]_ , \new_[4862]_ , \new_[4865]_ ,
    \new_[4866]_ , \new_[4867]_ , \new_[4870]_ , \new_[4873]_ ,
    \new_[4874]_ , \new_[4877]_ , \new_[4881]_ , \new_[4882]_ ,
    \new_[4883]_ , \new_[4884]_ , \new_[4885]_ , \new_[4888]_ ,
    \new_[4891]_ , \new_[4892]_ , \new_[4895]_ , \new_[4899]_ ,
    \new_[4900]_ , \new_[4901]_ , \new_[4902]_ , \new_[4905]_ ,
    \new_[4908]_ , \new_[4909]_ , \new_[4912]_ , \new_[4916]_ ,
    \new_[4917]_ , \new_[4918]_ , \new_[4919]_ , \new_[4920]_ ,
    \new_[4921]_ , \new_[4922]_ , \new_[4923]_ , \new_[4924]_ ,
    \new_[4927]_ , \new_[4930]_ , \new_[4931]_ , \new_[4934]_ ,
    \new_[4937]_ , \new_[4938]_ , \new_[4939]_ , \new_[4942]_ ,
    \new_[4945]_ , \new_[4946]_ , \new_[4949]_ , \new_[4953]_ ,
    \new_[4954]_ , \new_[4955]_ , \new_[4956]_ , \new_[4957]_ ,
    \new_[4960]_ , \new_[4963]_ , \new_[4964]_ , \new_[4967]_ ,
    \new_[4970]_ , \new_[4971]_ , \new_[4972]_ , \new_[4975]_ ,
    \new_[4978]_ , \new_[4979]_ , \new_[4982]_ , \new_[4986]_ ,
    \new_[4987]_ , \new_[4988]_ , \new_[4989]_ , \new_[4990]_ ,
    \new_[4991]_ , \new_[4994]_ , \new_[4997]_ , \new_[4998]_ ,
    \new_[5001]_ , \new_[5004]_ , \new_[5005]_ , \new_[5006]_ ,
    \new_[5009]_ , \new_[5012]_ , \new_[5013]_ , \new_[5016]_ ,
    \new_[5020]_ , \new_[5021]_ , \new_[5022]_ , \new_[5023]_ ,
    \new_[5024]_ , \new_[5027]_ , \new_[5030]_ , \new_[5031]_ ,
    \new_[5034]_ , \new_[5037]_ , \new_[5038]_ , \new_[5039]_ ,
    \new_[5042]_ , \new_[5045]_ , \new_[5046]_ , \new_[5049]_ ,
    \new_[5053]_ , \new_[5054]_ , \new_[5055]_ , \new_[5056]_ ,
    \new_[5057]_ , \new_[5058]_ , \new_[5059]_ , \new_[5062]_ ,
    \new_[5065]_ , \new_[5066]_ , \new_[5069]_ , \new_[5072]_ ,
    \new_[5073]_ , \new_[5074]_ , \new_[5077]_ , \new_[5080]_ ,
    \new_[5081]_ , \new_[5084]_ , \new_[5088]_ , \new_[5089]_ ,
    \new_[5090]_ , \new_[5091]_ , \new_[5092]_ , \new_[5095]_ ,
    \new_[5098]_ , \new_[5099]_ , \new_[5102]_ , \new_[5105]_ ,
    \new_[5106]_ , \new_[5107]_ , \new_[5110]_ , \new_[5113]_ ,
    \new_[5114]_ , \new_[5117]_ , \new_[5121]_ , \new_[5122]_ ,
    \new_[5123]_ , \new_[5124]_ , \new_[5125]_ , \new_[5126]_ ,
    \new_[5129]_ , \new_[5132]_ , \new_[5133]_ , \new_[5136]_ ,
    \new_[5139]_ , \new_[5140]_ , \new_[5141]_ , \new_[5144]_ ,
    \new_[5147]_ , \new_[5148]_ , \new_[5151]_ , \new_[5155]_ ,
    \new_[5156]_ , \new_[5157]_ , \new_[5158]_ , \new_[5159]_ ,
    \new_[5162]_ , \new_[5165]_ , \new_[5166]_ , \new_[5169]_ ,
    \new_[5173]_ , \new_[5174]_ , \new_[5175]_ , \new_[5176]_ ,
    \new_[5179]_ , \new_[5182]_ , \new_[5183]_ , \new_[5186]_ ,
    \new_[5190]_ , \new_[5191]_ , \new_[5192]_ , \new_[5193]_ ,
    \new_[5194]_ , \new_[5195]_ , \new_[5196]_ , \new_[5197]_ ,
    \new_[5200]_ , \new_[5203]_ , \new_[5204]_ , \new_[5207]_ ,
    \new_[5210]_ , \new_[5211]_ , \new_[5212]_ , \new_[5215]_ ,
    \new_[5218]_ , \new_[5219]_ , \new_[5222]_ , \new_[5226]_ ,
    \new_[5227]_ , \new_[5228]_ , \new_[5229]_ , \new_[5230]_ ,
    \new_[5233]_ , \new_[5236]_ , \new_[5237]_ , \new_[5240]_ ,
    \new_[5243]_ , \new_[5244]_ , \new_[5245]_ , \new_[5248]_ ,
    \new_[5251]_ , \new_[5252]_ , \new_[5255]_ , \new_[5259]_ ,
    \new_[5260]_ , \new_[5261]_ , \new_[5262]_ , \new_[5263]_ ,
    \new_[5264]_ , \new_[5267]_ , \new_[5270]_ , \new_[5271]_ ,
    \new_[5274]_ , \new_[5277]_ , \new_[5278]_ , \new_[5279]_ ,
    \new_[5282]_ , \new_[5285]_ , \new_[5286]_ , \new_[5289]_ ,
    \new_[5293]_ , \new_[5294]_ , \new_[5295]_ , \new_[5296]_ ,
    \new_[5297]_ , \new_[5300]_ , \new_[5303]_ , \new_[5304]_ ,
    \new_[5307]_ , \new_[5310]_ , \new_[5311]_ , \new_[5312]_ ,
    \new_[5315]_ , \new_[5318]_ , \new_[5319]_ , \new_[5322]_ ,
    \new_[5326]_ , \new_[5327]_ , \new_[5328]_ , \new_[5329]_ ,
    \new_[5330]_ , \new_[5331]_ , \new_[5332]_ , \new_[5335]_ ,
    \new_[5338]_ , \new_[5339]_ , \new_[5342]_ , \new_[5345]_ ,
    \new_[5346]_ , \new_[5347]_ , \new_[5350]_ , \new_[5353]_ ,
    \new_[5354]_ , \new_[5357]_ , \new_[5361]_ , \new_[5362]_ ,
    \new_[5363]_ , \new_[5364]_ , \new_[5365]_ , \new_[5368]_ ,
    \new_[5371]_ , \new_[5372]_ , \new_[5375]_ , \new_[5378]_ ,
    \new_[5379]_ , \new_[5380]_ , \new_[5383]_ , \new_[5386]_ ,
    \new_[5387]_ , \new_[5390]_ , \new_[5394]_ , \new_[5395]_ ,
    \new_[5396]_ , \new_[5397]_ , \new_[5398]_ , \new_[5399]_ ,
    \new_[5402]_ , \new_[5405]_ , \new_[5406]_ , \new_[5409]_ ,
    \new_[5412]_ , \new_[5413]_ , \new_[5414]_ , \new_[5417]_ ,
    \new_[5420]_ , \new_[5421]_ , \new_[5424]_ , \new_[5428]_ ,
    \new_[5429]_ , \new_[5430]_ , \new_[5431]_ , \new_[5432]_ ,
    \new_[5435]_ , \new_[5438]_ , \new_[5439]_ , \new_[5442]_ ,
    \new_[5446]_ , \new_[5447]_ , \new_[5448]_ , \new_[5449]_ ,
    \new_[5452]_ , \new_[5455]_ , \new_[5456]_ , \new_[5459]_ ,
    \new_[5463]_ , \new_[5464]_ , \new_[5465]_ , \new_[5466]_ ,
    \new_[5467]_ , \new_[5468]_ , \new_[5469]_ , \new_[5470]_ ,
    \new_[5471]_ , \new_[5472]_ , \new_[5475]_ , \new_[5478]_ ,
    \new_[5479]_ , \new_[5482]_ , \new_[5485]_ , \new_[5486]_ ,
    \new_[5487]_ , \new_[5490]_ , \new_[5493]_ , \new_[5494]_ ,
    \new_[5497]_ , \new_[5501]_ , \new_[5502]_ , \new_[5503]_ ,
    \new_[5504]_ , \new_[5505]_ , \new_[5508]_ , \new_[5511]_ ,
    \new_[5512]_ , \new_[5515]_ , \new_[5518]_ , \new_[5519]_ ,
    \new_[5520]_ , \new_[5523]_ , \new_[5526]_ , \new_[5527]_ ,
    \new_[5530]_ , \new_[5534]_ , \new_[5535]_ , \new_[5536]_ ,
    \new_[5537]_ , \new_[5538]_ , \new_[5539]_ , \new_[5542]_ ,
    \new_[5545]_ , \new_[5546]_ , \new_[5549]_ , \new_[5552]_ ,
    \new_[5553]_ , \new_[5554]_ , \new_[5557]_ , \new_[5560]_ ,
    \new_[5561]_ , \new_[5564]_ , \new_[5568]_ , \new_[5569]_ ,
    \new_[5570]_ , \new_[5571]_ , \new_[5572]_ , \new_[5575]_ ,
    \new_[5578]_ , \new_[5579]_ , \new_[5582]_ , \new_[5585]_ ,
    \new_[5586]_ , \new_[5587]_ , \new_[5590]_ , \new_[5593]_ ,
    \new_[5594]_ , \new_[5597]_ , \new_[5601]_ , \new_[5602]_ ,
    \new_[5603]_ , \new_[5604]_ , \new_[5605]_ , \new_[5606]_ ,
    \new_[5607]_ , \new_[5610]_ , \new_[5613]_ , \new_[5614]_ ,
    \new_[5617]_ , \new_[5620]_ , \new_[5621]_ , \new_[5622]_ ,
    \new_[5625]_ , \new_[5628]_ , \new_[5629]_ , \new_[5632]_ ,
    \new_[5636]_ , \new_[5637]_ , \new_[5638]_ , \new_[5639]_ ,
    \new_[5640]_ , \new_[5643]_ , \new_[5646]_ , \new_[5647]_ ,
    \new_[5650]_ , \new_[5653]_ , \new_[5654]_ , \new_[5655]_ ,
    \new_[5658]_ , \new_[5661]_ , \new_[5662]_ , \new_[5665]_ ,
    \new_[5669]_ , \new_[5670]_ , \new_[5671]_ , \new_[5672]_ ,
    \new_[5673]_ , \new_[5674]_ , \new_[5677]_ , \new_[5680]_ ,
    \new_[5681]_ , \new_[5684]_ , \new_[5687]_ , \new_[5688]_ ,
    \new_[5689]_ , \new_[5692]_ , \new_[5695]_ , \new_[5696]_ ,
    \new_[5699]_ , \new_[5703]_ , \new_[5704]_ , \new_[5705]_ ,
    \new_[5706]_ , \new_[5707]_ , \new_[5710]_ , \new_[5713]_ ,
    \new_[5714]_ , \new_[5717]_ , \new_[5721]_ , \new_[5722]_ ,
    \new_[5723]_ , \new_[5724]_ , \new_[5727]_ , \new_[5730]_ ,
    \new_[5731]_ , \new_[5734]_ , \new_[5738]_ , \new_[5739]_ ,
    \new_[5740]_ , \new_[5741]_ , \new_[5742]_ , \new_[5743]_ ,
    \new_[5744]_ , \new_[5745]_ , \new_[5748]_ , \new_[5751]_ ,
    \new_[5752]_ , \new_[5755]_ , \new_[5758]_ , \new_[5759]_ ,
    \new_[5760]_ , \new_[5763]_ , \new_[5766]_ , \new_[5767]_ ,
    \new_[5770]_ , \new_[5774]_ , \new_[5775]_ , \new_[5776]_ ,
    \new_[5777]_ , \new_[5778]_ , \new_[5781]_ , \new_[5784]_ ,
    \new_[5785]_ , \new_[5788]_ , \new_[5791]_ , \new_[5792]_ ,
    \new_[5793]_ , \new_[5796]_ , \new_[5799]_ , \new_[5800]_ ,
    \new_[5803]_ , \new_[5807]_ , \new_[5808]_ , \new_[5809]_ ,
    \new_[5810]_ , \new_[5811]_ , \new_[5812]_ , \new_[5815]_ ,
    \new_[5818]_ , \new_[5819]_ , \new_[5822]_ , \new_[5825]_ ,
    \new_[5826]_ , \new_[5827]_ , \new_[5830]_ , \new_[5833]_ ,
    \new_[5834]_ , \new_[5837]_ , \new_[5841]_ , \new_[5842]_ ,
    \new_[5843]_ , \new_[5844]_ , \new_[5845]_ , \new_[5848]_ ,
    \new_[5851]_ , \new_[5852]_ , \new_[5855]_ , \new_[5858]_ ,
    \new_[5859]_ , \new_[5860]_ , \new_[5863]_ , \new_[5866]_ ,
    \new_[5867]_ , \new_[5870]_ , \new_[5874]_ , \new_[5875]_ ,
    \new_[5876]_ , \new_[5877]_ , \new_[5878]_ , \new_[5879]_ ,
    \new_[5880]_ , \new_[5883]_ , \new_[5886]_ , \new_[5887]_ ,
    \new_[5890]_ , \new_[5893]_ , \new_[5894]_ , \new_[5895]_ ,
    \new_[5898]_ , \new_[5901]_ , \new_[5902]_ , \new_[5905]_ ,
    \new_[5909]_ , \new_[5910]_ , \new_[5911]_ , \new_[5912]_ ,
    \new_[5913]_ , \new_[5916]_ , \new_[5919]_ , \new_[5920]_ ,
    \new_[5923]_ , \new_[5926]_ , \new_[5927]_ , \new_[5928]_ ,
    \new_[5931]_ , \new_[5934]_ , \new_[5935]_ , \new_[5938]_ ,
    \new_[5942]_ , \new_[5943]_ , \new_[5944]_ , \new_[5945]_ ,
    \new_[5946]_ , \new_[5947]_ , \new_[5950]_ , \new_[5953]_ ,
    \new_[5954]_ , \new_[5957]_ , \new_[5960]_ , \new_[5961]_ ,
    \new_[5962]_ , \new_[5965]_ , \new_[5968]_ , \new_[5969]_ ,
    \new_[5972]_ , \new_[5976]_ , \new_[5977]_ , \new_[5978]_ ,
    \new_[5979]_ , \new_[5980]_ , \new_[5983]_ , \new_[5986]_ ,
    \new_[5987]_ , \new_[5990]_ , \new_[5994]_ , \new_[5995]_ ,
    \new_[5996]_ , \new_[5997]_ , \new_[6000]_ , \new_[6003]_ ,
    \new_[6004]_ , \new_[6007]_ , \new_[6011]_ , \new_[6012]_ ,
    \new_[6013]_ , \new_[6014]_ , \new_[6015]_ , \new_[6016]_ ,
    \new_[6017]_ , \new_[6018]_ , \new_[6019]_ , \new_[6022]_ ,
    \new_[6025]_ , \new_[6026]_ , \new_[6029]_ , \new_[6032]_ ,
    \new_[6033]_ , \new_[6034]_ , \new_[6037]_ , \new_[6040]_ ,
    \new_[6041]_ , \new_[6044]_ , \new_[6048]_ , \new_[6049]_ ,
    \new_[6050]_ , \new_[6051]_ , \new_[6052]_ , \new_[6055]_ ,
    \new_[6058]_ , \new_[6059]_ , \new_[6062]_ , \new_[6065]_ ,
    \new_[6066]_ , \new_[6067]_ , \new_[6070]_ , \new_[6073]_ ,
    \new_[6074]_ , \new_[6077]_ , \new_[6081]_ , \new_[6082]_ ,
    \new_[6083]_ , \new_[6084]_ , \new_[6085]_ , \new_[6086]_ ,
    \new_[6089]_ , \new_[6092]_ , \new_[6093]_ , \new_[6096]_ ,
    \new_[6099]_ , \new_[6100]_ , \new_[6101]_ , \new_[6104]_ ,
    \new_[6107]_ , \new_[6108]_ , \new_[6111]_ , \new_[6115]_ ,
    \new_[6116]_ , \new_[6117]_ , \new_[6118]_ , \new_[6119]_ ,
    \new_[6122]_ , \new_[6125]_ , \new_[6126]_ , \new_[6129]_ ,
    \new_[6132]_ , \new_[6133]_ , \new_[6134]_ , \new_[6137]_ ,
    \new_[6140]_ , \new_[6141]_ , \new_[6144]_ , \new_[6148]_ ,
    \new_[6149]_ , \new_[6150]_ , \new_[6151]_ , \new_[6152]_ ,
    \new_[6153]_ , \new_[6154]_ , \new_[6157]_ , \new_[6160]_ ,
    \new_[6161]_ , \new_[6164]_ , \new_[6167]_ , \new_[6168]_ ,
    \new_[6169]_ , \new_[6172]_ , \new_[6175]_ , \new_[6176]_ ,
    \new_[6179]_ , \new_[6183]_ , \new_[6184]_ , \new_[6185]_ ,
    \new_[6186]_ , \new_[6187]_ , \new_[6190]_ , \new_[6193]_ ,
    \new_[6194]_ , \new_[6197]_ , \new_[6200]_ , \new_[6201]_ ,
    \new_[6202]_ , \new_[6205]_ , \new_[6208]_ , \new_[6209]_ ,
    \new_[6212]_ , \new_[6216]_ , \new_[6217]_ , \new_[6218]_ ,
    \new_[6219]_ , \new_[6220]_ , \new_[6221]_ , \new_[6224]_ ,
    \new_[6227]_ , \new_[6228]_ , \new_[6231]_ , \new_[6234]_ ,
    \new_[6235]_ , \new_[6236]_ , \new_[6239]_ , \new_[6242]_ ,
    \new_[6243]_ , \new_[6246]_ , \new_[6250]_ , \new_[6251]_ ,
    \new_[6252]_ , \new_[6253]_ , \new_[6254]_ , \new_[6257]_ ,
    \new_[6260]_ , \new_[6261]_ , \new_[6264]_ , \new_[6268]_ ,
    \new_[6269]_ , \new_[6270]_ , \new_[6271]_ , \new_[6274]_ ,
    \new_[6277]_ , \new_[6278]_ , \new_[6281]_ , \new_[6285]_ ,
    \new_[6286]_ , \new_[6287]_ , \new_[6288]_ , \new_[6289]_ ,
    \new_[6290]_ , \new_[6291]_ , \new_[6292]_ , \new_[6295]_ ,
    \new_[6298]_ , \new_[6299]_ , \new_[6302]_ , \new_[6305]_ ,
    \new_[6306]_ , \new_[6307]_ , \new_[6310]_ , \new_[6313]_ ,
    \new_[6314]_ , \new_[6317]_ , \new_[6321]_ , \new_[6322]_ ,
    \new_[6323]_ , \new_[6324]_ , \new_[6325]_ , \new_[6328]_ ,
    \new_[6331]_ , \new_[6332]_ , \new_[6335]_ , \new_[6338]_ ,
    \new_[6339]_ , \new_[6340]_ , \new_[6343]_ , \new_[6346]_ ,
    \new_[6347]_ , \new_[6350]_ , \new_[6354]_ , \new_[6355]_ ,
    \new_[6356]_ , \new_[6357]_ , \new_[6358]_ , \new_[6359]_ ,
    \new_[6362]_ , \new_[6365]_ , \new_[6366]_ , \new_[6369]_ ,
    \new_[6372]_ , \new_[6373]_ , \new_[6374]_ , \new_[6377]_ ,
    \new_[6380]_ , \new_[6381]_ , \new_[6384]_ , \new_[6388]_ ,
    \new_[6389]_ , \new_[6390]_ , \new_[6391]_ , \new_[6392]_ ,
    \new_[6395]_ , \new_[6398]_ , \new_[6399]_ , \new_[6402]_ ,
    \new_[6405]_ , \new_[6406]_ , \new_[6407]_ , \new_[6410]_ ,
    \new_[6413]_ , \new_[6414]_ , \new_[6417]_ , \new_[6421]_ ,
    \new_[6422]_ , \new_[6423]_ , \new_[6424]_ , \new_[6425]_ ,
    \new_[6426]_ , \new_[6427]_ , \new_[6430]_ , \new_[6433]_ ,
    \new_[6434]_ , \new_[6437]_ , \new_[6440]_ , \new_[6441]_ ,
    \new_[6442]_ , \new_[6445]_ , \new_[6448]_ , \new_[6449]_ ,
    \new_[6452]_ , \new_[6456]_ , \new_[6457]_ , \new_[6458]_ ,
    \new_[6459]_ , \new_[6460]_ , \new_[6463]_ , \new_[6466]_ ,
    \new_[6467]_ , \new_[6470]_ , \new_[6473]_ , \new_[6474]_ ,
    \new_[6475]_ , \new_[6478]_ , \new_[6481]_ , \new_[6482]_ ,
    \new_[6485]_ , \new_[6489]_ , \new_[6490]_ , \new_[6491]_ ,
    \new_[6492]_ , \new_[6493]_ , \new_[6494]_ , \new_[6497]_ ,
    \new_[6500]_ , \new_[6501]_ , \new_[6504]_ , \new_[6507]_ ,
    \new_[6508]_ , \new_[6509]_ , \new_[6512]_ , \new_[6515]_ ,
    \new_[6516]_ , \new_[6519]_ , \new_[6523]_ , \new_[6524]_ ,
    \new_[6525]_ , \new_[6526]_ , \new_[6527]_ , \new_[6530]_ ,
    \new_[6533]_ , \new_[6534]_ , \new_[6537]_ , \new_[6541]_ ,
    \new_[6542]_ , \new_[6543]_ , \new_[6544]_ , \new_[6547]_ ,
    \new_[6550]_ , \new_[6551]_ , \new_[6554]_ , \new_[6558]_ ,
    \new_[6559]_ , \new_[6560]_ , \new_[6561]_ , \new_[6562]_ ,
    \new_[6563]_ , \new_[6564]_ , \new_[6565]_ , \new_[6566]_ ,
    \new_[6567]_ , \new_[6568]_ , \new_[6572]_ , \new_[6573]_ ,
    \new_[6577]_ , \new_[6578]_ , \new_[6582]_ , \new_[6583]_ ,
    \new_[6587]_ , \new_[6588]_ , \new_[6592]_ , \new_[6593]_ ,
    \new_[6597]_ , \new_[6598]_ , \new_[6602]_ , \new_[6603]_ ,
    \new_[6607]_ , \new_[6608]_ , \new_[6612]_ , \new_[6613]_ ,
    \new_[6617]_ , \new_[6618]_ , \new_[6622]_ , \new_[6623]_ ,
    \new_[6627]_ , \new_[6628]_ , \new_[6632]_ , \new_[6633]_ ,
    \new_[6637]_ , \new_[6638]_ , \new_[6642]_ , \new_[6643]_ ,
    \new_[6647]_ , \new_[6648]_ , \new_[6652]_ , \new_[6653]_ ,
    \new_[6657]_ , \new_[6658]_ , \new_[6662]_ , \new_[6663]_ ,
    \new_[6667]_ , \new_[6668]_ , \new_[6672]_ , \new_[6673]_ ,
    \new_[6677]_ , \new_[6678]_ , \new_[6682]_ , \new_[6683]_ ,
    \new_[6687]_ , \new_[6688]_ , \new_[6692]_ , \new_[6693]_ ,
    \new_[6697]_ , \new_[6698]_ , \new_[6702]_ , \new_[6703]_ ,
    \new_[6707]_ , \new_[6708]_ , \new_[6712]_ , \new_[6713]_ ,
    \new_[6717]_ , \new_[6718]_ , \new_[6722]_ , \new_[6723]_ ,
    \new_[6727]_ , \new_[6728]_ , \new_[6732]_ , \new_[6733]_ ,
    \new_[6736]_ , \new_[6739]_ , \new_[6740]_ , \new_[6744]_ ,
    \new_[6745]_ , \new_[6748]_ , \new_[6751]_ , \new_[6752]_ ,
    \new_[6756]_ , \new_[6757]_ , \new_[6760]_ , \new_[6763]_ ,
    \new_[6764]_ , \new_[6768]_ , \new_[6769]_ , \new_[6772]_ ,
    \new_[6775]_ , \new_[6776]_ , \new_[6780]_ , \new_[6781]_ ,
    \new_[6784]_ , \new_[6787]_ , \new_[6788]_ , \new_[6792]_ ,
    \new_[6793]_ , \new_[6796]_ , \new_[6799]_ , \new_[6800]_ ,
    \new_[6804]_ , \new_[6805]_ , \new_[6808]_ , \new_[6811]_ ,
    \new_[6812]_ , \new_[6816]_ , \new_[6817]_ , \new_[6820]_ ,
    \new_[6823]_ , \new_[6824]_ , \new_[6828]_ , \new_[6829]_ ,
    \new_[6832]_ , \new_[6835]_ , \new_[6836]_ , \new_[6840]_ ,
    \new_[6841]_ , \new_[6844]_ , \new_[6847]_ , \new_[6848]_ ,
    \new_[6852]_ , \new_[6853]_ , \new_[6856]_ , \new_[6859]_ ,
    \new_[6860]_ , \new_[6864]_ , \new_[6865]_ , \new_[6868]_ ,
    \new_[6871]_ , \new_[6872]_ , \new_[6875]_ , \new_[6878]_ ,
    \new_[6879]_ , \new_[6882]_ , \new_[6885]_ , \new_[6886]_ ,
    \new_[6889]_ , \new_[6892]_ , \new_[6893]_ , \new_[6896]_ ,
    \new_[6899]_ , \new_[6900]_ , \new_[6904]_ , \new_[6905]_ ,
    \new_[6908]_ , \new_[6911]_ , \new_[6912]_ , \new_[6913]_ ,
    \new_[6917]_ , \new_[6918]_ , \new_[6921]_ , \new_[6924]_ ,
    \new_[6925]_ , \new_[6926]_ , \new_[6930]_ , \new_[6931]_ ,
    \new_[6934]_ , \new_[6937]_ , \new_[6938]_ , \new_[6939]_ ,
    \new_[6943]_ , \new_[6944]_ , \new_[6947]_ , \new_[6950]_ ,
    \new_[6951]_ , \new_[6952]_ , \new_[6956]_ , \new_[6957]_ ,
    \new_[6960]_ , \new_[6963]_ , \new_[6964]_ , \new_[6965]_ ,
    \new_[6969]_ , \new_[6970]_ , \new_[6973]_ , \new_[6976]_ ,
    \new_[6977]_ , \new_[6978]_ , \new_[6982]_ , \new_[6983]_ ,
    \new_[6986]_ , \new_[6989]_ , \new_[6990]_ , \new_[6991]_ ,
    \new_[6995]_ , \new_[6996]_ , \new_[6999]_ , \new_[7002]_ ,
    \new_[7003]_ , \new_[7004]_ , \new_[7008]_ , \new_[7009]_ ,
    \new_[7012]_ , \new_[7015]_ , \new_[7016]_ , \new_[7017]_ ,
    \new_[7021]_ , \new_[7022]_ , \new_[7025]_ , \new_[7028]_ ,
    \new_[7029]_ , \new_[7030]_ , \new_[7034]_ , \new_[7035]_ ,
    \new_[7038]_ , \new_[7041]_ , \new_[7042]_ , \new_[7043]_ ,
    \new_[7047]_ , \new_[7048]_ , \new_[7051]_ , \new_[7054]_ ,
    \new_[7055]_ , \new_[7056]_ , \new_[7060]_ , \new_[7061]_ ,
    \new_[7064]_ , \new_[7067]_ , \new_[7068]_ , \new_[7069]_ ,
    \new_[7073]_ , \new_[7074]_ , \new_[7077]_ , \new_[7080]_ ,
    \new_[7081]_ , \new_[7082]_ , \new_[7086]_ , \new_[7087]_ ,
    \new_[7090]_ , \new_[7093]_ , \new_[7094]_ , \new_[7095]_ ,
    \new_[7099]_ , \new_[7100]_ , \new_[7103]_ , \new_[7106]_ ,
    \new_[7107]_ , \new_[7108]_ , \new_[7112]_ , \new_[7113]_ ,
    \new_[7116]_ , \new_[7119]_ , \new_[7120]_ , \new_[7121]_ ,
    \new_[7125]_ , \new_[7126]_ , \new_[7129]_ , \new_[7132]_ ,
    \new_[7133]_ , \new_[7134]_ , \new_[7138]_ , \new_[7139]_ ,
    \new_[7142]_ , \new_[7145]_ , \new_[7146]_ , \new_[7147]_ ,
    \new_[7151]_ , \new_[7152]_ , \new_[7155]_ , \new_[7158]_ ,
    \new_[7159]_ , \new_[7160]_ , \new_[7164]_ , \new_[7165]_ ,
    \new_[7168]_ , \new_[7171]_ , \new_[7172]_ , \new_[7173]_ ,
    \new_[7177]_ , \new_[7178]_ , \new_[7181]_ , \new_[7184]_ ,
    \new_[7185]_ , \new_[7186]_ , \new_[7190]_ , \new_[7191]_ ,
    \new_[7194]_ , \new_[7197]_ , \new_[7198]_ , \new_[7199]_ ,
    \new_[7203]_ , \new_[7204]_ , \new_[7207]_ , \new_[7210]_ ,
    \new_[7211]_ , \new_[7212]_ , \new_[7216]_ , \new_[7217]_ ,
    \new_[7220]_ , \new_[7223]_ , \new_[7224]_ , \new_[7225]_ ,
    \new_[7229]_ , \new_[7230]_ , \new_[7233]_ , \new_[7236]_ ,
    \new_[7237]_ , \new_[7238]_ , \new_[7242]_ , \new_[7243]_ ,
    \new_[7246]_ , \new_[7249]_ , \new_[7250]_ , \new_[7251]_ ,
    \new_[7255]_ , \new_[7256]_ , \new_[7259]_ , \new_[7262]_ ,
    \new_[7263]_ , \new_[7264]_ , \new_[7268]_ , \new_[7269]_ ,
    \new_[7272]_ , \new_[7275]_ , \new_[7276]_ , \new_[7277]_ ,
    \new_[7281]_ , \new_[7282]_ , \new_[7285]_ , \new_[7288]_ ,
    \new_[7289]_ , \new_[7290]_ , \new_[7294]_ , \new_[7295]_ ,
    \new_[7298]_ , \new_[7301]_ , \new_[7302]_ , \new_[7303]_ ,
    \new_[7307]_ , \new_[7308]_ , \new_[7311]_ , \new_[7314]_ ,
    \new_[7315]_ , \new_[7316]_ , \new_[7320]_ , \new_[7321]_ ,
    \new_[7324]_ , \new_[7327]_ , \new_[7328]_ , \new_[7329]_ ,
    \new_[7333]_ , \new_[7334]_ , \new_[7337]_ , \new_[7340]_ ,
    \new_[7341]_ , \new_[7342]_ , \new_[7346]_ , \new_[7347]_ ,
    \new_[7350]_ , \new_[7353]_ , \new_[7354]_ , \new_[7355]_ ,
    \new_[7359]_ , \new_[7360]_ , \new_[7363]_ , \new_[7366]_ ,
    \new_[7367]_ , \new_[7368]_ , \new_[7372]_ , \new_[7373]_ ,
    \new_[7376]_ , \new_[7379]_ , \new_[7380]_ , \new_[7381]_ ,
    \new_[7385]_ , \new_[7386]_ , \new_[7389]_ , \new_[7392]_ ,
    \new_[7393]_ , \new_[7394]_ , \new_[7398]_ , \new_[7399]_ ,
    \new_[7402]_ , \new_[7405]_ , \new_[7406]_ , \new_[7407]_ ,
    \new_[7411]_ , \new_[7412]_ , \new_[7415]_ , \new_[7418]_ ,
    \new_[7419]_ , \new_[7420]_ , \new_[7424]_ , \new_[7425]_ ,
    \new_[7428]_ , \new_[7431]_ , \new_[7432]_ , \new_[7433]_ ,
    \new_[7437]_ , \new_[7438]_ , \new_[7441]_ , \new_[7444]_ ,
    \new_[7445]_ , \new_[7446]_ , \new_[7450]_ , \new_[7451]_ ,
    \new_[7454]_ , \new_[7457]_ , \new_[7458]_ , \new_[7459]_ ,
    \new_[7463]_ , \new_[7464]_ , \new_[7467]_ , \new_[7470]_ ,
    \new_[7471]_ , \new_[7472]_ , \new_[7476]_ , \new_[7477]_ ,
    \new_[7480]_ , \new_[7483]_ , \new_[7484]_ , \new_[7485]_ ,
    \new_[7489]_ , \new_[7490]_ , \new_[7493]_ , \new_[7496]_ ,
    \new_[7497]_ , \new_[7498]_ , \new_[7502]_ , \new_[7503]_ ,
    \new_[7506]_ , \new_[7509]_ , \new_[7510]_ , \new_[7511]_ ,
    \new_[7515]_ , \new_[7516]_ , \new_[7519]_ , \new_[7522]_ ,
    \new_[7523]_ , \new_[7524]_ , \new_[7528]_ , \new_[7529]_ ,
    \new_[7532]_ , \new_[7535]_ , \new_[7536]_ , \new_[7537]_ ,
    \new_[7541]_ , \new_[7542]_ , \new_[7545]_ , \new_[7548]_ ,
    \new_[7549]_ , \new_[7550]_ , \new_[7554]_ , \new_[7555]_ ,
    \new_[7558]_ , \new_[7561]_ , \new_[7562]_ , \new_[7563]_ ,
    \new_[7567]_ , \new_[7568]_ , \new_[7571]_ , \new_[7574]_ ,
    \new_[7575]_ , \new_[7576]_ , \new_[7580]_ , \new_[7581]_ ,
    \new_[7584]_ , \new_[7587]_ , \new_[7588]_ , \new_[7589]_ ,
    \new_[7593]_ , \new_[7594]_ , \new_[7597]_ , \new_[7600]_ ,
    \new_[7601]_ , \new_[7602]_ , \new_[7606]_ , \new_[7607]_ ,
    \new_[7610]_ , \new_[7613]_ , \new_[7614]_ , \new_[7615]_ ,
    \new_[7619]_ , \new_[7620]_ , \new_[7623]_ , \new_[7626]_ ,
    \new_[7627]_ , \new_[7628]_ , \new_[7632]_ , \new_[7633]_ ,
    \new_[7636]_ , \new_[7639]_ , \new_[7640]_ , \new_[7641]_ ,
    \new_[7645]_ , \new_[7646]_ , \new_[7649]_ , \new_[7652]_ ,
    \new_[7653]_ , \new_[7654]_ , \new_[7658]_ , \new_[7659]_ ,
    \new_[7662]_ , \new_[7665]_ , \new_[7666]_ , \new_[7667]_ ,
    \new_[7671]_ , \new_[7672]_ , \new_[7675]_ , \new_[7678]_ ,
    \new_[7679]_ , \new_[7680]_ , \new_[7684]_ , \new_[7685]_ ,
    \new_[7688]_ , \new_[7691]_ , \new_[7692]_ , \new_[7693]_ ,
    \new_[7697]_ , \new_[7698]_ , \new_[7701]_ , \new_[7704]_ ,
    \new_[7705]_ , \new_[7706]_ , \new_[7710]_ , \new_[7711]_ ,
    \new_[7714]_ , \new_[7717]_ , \new_[7718]_ , \new_[7719]_ ,
    \new_[7723]_ , \new_[7724]_ , \new_[7727]_ , \new_[7730]_ ,
    \new_[7731]_ , \new_[7732]_ , \new_[7736]_ , \new_[7737]_ ,
    \new_[7740]_ , \new_[7743]_ , \new_[7744]_ , \new_[7745]_ ,
    \new_[7749]_ , \new_[7750]_ , \new_[7753]_ , \new_[7756]_ ,
    \new_[7757]_ , \new_[7758]_ , \new_[7762]_ , \new_[7763]_ ,
    \new_[7766]_ , \new_[7769]_ , \new_[7770]_ , \new_[7771]_ ,
    \new_[7775]_ , \new_[7776]_ , \new_[7779]_ , \new_[7782]_ ,
    \new_[7783]_ , \new_[7784]_ , \new_[7788]_ , \new_[7789]_ ,
    \new_[7792]_ , \new_[7795]_ , \new_[7796]_ , \new_[7797]_ ,
    \new_[7801]_ , \new_[7802]_ , \new_[7805]_ , \new_[7808]_ ,
    \new_[7809]_ , \new_[7810]_ , \new_[7814]_ , \new_[7815]_ ,
    \new_[7818]_ , \new_[7821]_ , \new_[7822]_ , \new_[7823]_ ,
    \new_[7827]_ , \new_[7828]_ , \new_[7831]_ , \new_[7834]_ ,
    \new_[7835]_ , \new_[7836]_ , \new_[7840]_ , \new_[7841]_ ,
    \new_[7844]_ , \new_[7847]_ , \new_[7848]_ , \new_[7849]_ ,
    \new_[7853]_ , \new_[7854]_ , \new_[7857]_ , \new_[7860]_ ,
    \new_[7861]_ , \new_[7862]_ , \new_[7866]_ , \new_[7867]_ ,
    \new_[7870]_ , \new_[7873]_ , \new_[7874]_ , \new_[7875]_ ,
    \new_[7879]_ , \new_[7880]_ , \new_[7883]_ , \new_[7886]_ ,
    \new_[7887]_ , \new_[7888]_ , \new_[7892]_ , \new_[7893]_ ,
    \new_[7896]_ , \new_[7899]_ , \new_[7900]_ , \new_[7901]_ ,
    \new_[7905]_ , \new_[7906]_ , \new_[7909]_ , \new_[7912]_ ,
    \new_[7913]_ , \new_[7914]_ , \new_[7918]_ , \new_[7919]_ ,
    \new_[7922]_ , \new_[7925]_ , \new_[7926]_ , \new_[7927]_ ,
    \new_[7931]_ , \new_[7932]_ , \new_[7935]_ , \new_[7938]_ ,
    \new_[7939]_ , \new_[7940]_ , \new_[7944]_ , \new_[7945]_ ,
    \new_[7948]_ , \new_[7951]_ , \new_[7952]_ , \new_[7953]_ ,
    \new_[7957]_ , \new_[7958]_ , \new_[7961]_ , \new_[7964]_ ,
    \new_[7965]_ , \new_[7966]_ , \new_[7970]_ , \new_[7971]_ ,
    \new_[7974]_ , \new_[7977]_ , \new_[7978]_ , \new_[7979]_ ,
    \new_[7983]_ , \new_[7984]_ , \new_[7987]_ , \new_[7990]_ ,
    \new_[7991]_ , \new_[7992]_ , \new_[7996]_ , \new_[7997]_ ,
    \new_[8000]_ , \new_[8003]_ , \new_[8004]_ , \new_[8005]_ ,
    \new_[8009]_ , \new_[8010]_ , \new_[8013]_ , \new_[8016]_ ,
    \new_[8017]_ , \new_[8018]_ , \new_[8022]_ , \new_[8023]_ ,
    \new_[8026]_ , \new_[8029]_ , \new_[8030]_ , \new_[8031]_ ,
    \new_[8035]_ , \new_[8036]_ , \new_[8039]_ , \new_[8042]_ ,
    \new_[8043]_ , \new_[8044]_ , \new_[8048]_ , \new_[8049]_ ,
    \new_[8052]_ , \new_[8055]_ , \new_[8056]_ , \new_[8057]_ ,
    \new_[8061]_ , \new_[8062]_ , \new_[8065]_ , \new_[8068]_ ,
    \new_[8069]_ , \new_[8070]_ , \new_[8074]_ , \new_[8075]_ ,
    \new_[8078]_ , \new_[8081]_ , \new_[8082]_ , \new_[8083]_ ,
    \new_[8087]_ , \new_[8088]_ , \new_[8091]_ , \new_[8094]_ ,
    \new_[8095]_ , \new_[8096]_ , \new_[8100]_ , \new_[8101]_ ,
    \new_[8104]_ , \new_[8107]_ , \new_[8108]_ , \new_[8109]_ ,
    \new_[8113]_ , \new_[8114]_ , \new_[8117]_ , \new_[8120]_ ,
    \new_[8121]_ , \new_[8122]_ , \new_[8126]_ , \new_[8127]_ ,
    \new_[8130]_ , \new_[8133]_ , \new_[8134]_ , \new_[8135]_ ,
    \new_[8139]_ , \new_[8140]_ , \new_[8143]_ , \new_[8146]_ ,
    \new_[8147]_ , \new_[8148]_ , \new_[8152]_ , \new_[8153]_ ,
    \new_[8156]_ , \new_[8159]_ , \new_[8160]_ , \new_[8161]_ ,
    \new_[8165]_ , \new_[8166]_ , \new_[8169]_ , \new_[8172]_ ,
    \new_[8173]_ , \new_[8174]_ , \new_[8178]_ , \new_[8179]_ ,
    \new_[8182]_ , \new_[8185]_ , \new_[8186]_ , \new_[8187]_ ,
    \new_[8191]_ , \new_[8192]_ , \new_[8195]_ , \new_[8198]_ ,
    \new_[8199]_ , \new_[8200]_ , \new_[8204]_ , \new_[8205]_ ,
    \new_[8208]_ , \new_[8211]_ , \new_[8212]_ , \new_[8213]_ ,
    \new_[8217]_ , \new_[8218]_ , \new_[8221]_ , \new_[8224]_ ,
    \new_[8225]_ , \new_[8226]_ , \new_[8230]_ , \new_[8231]_ ,
    \new_[8234]_ , \new_[8237]_ , \new_[8238]_ , \new_[8239]_ ,
    \new_[8243]_ , \new_[8244]_ , \new_[8247]_ , \new_[8250]_ ,
    \new_[8251]_ , \new_[8252]_ , \new_[8256]_ , \new_[8257]_ ,
    \new_[8260]_ , \new_[8263]_ , \new_[8264]_ , \new_[8265]_ ,
    \new_[8269]_ , \new_[8270]_ , \new_[8273]_ , \new_[8276]_ ,
    \new_[8277]_ , \new_[8278]_ , \new_[8282]_ , \new_[8283]_ ,
    \new_[8286]_ , \new_[8289]_ , \new_[8290]_ , \new_[8291]_ ,
    \new_[8295]_ , \new_[8296]_ , \new_[8299]_ , \new_[8302]_ ,
    \new_[8303]_ , \new_[8304]_ , \new_[8308]_ , \new_[8309]_ ,
    \new_[8312]_ , \new_[8315]_ , \new_[8316]_ , \new_[8317]_ ,
    \new_[8321]_ , \new_[8322]_ , \new_[8325]_ , \new_[8328]_ ,
    \new_[8329]_ , \new_[8330]_ , \new_[8334]_ , \new_[8335]_ ,
    \new_[8338]_ , \new_[8341]_ , \new_[8342]_ , \new_[8343]_ ,
    \new_[8347]_ , \new_[8348]_ , \new_[8351]_ , \new_[8354]_ ,
    \new_[8355]_ , \new_[8356]_ , \new_[8360]_ , \new_[8361]_ ,
    \new_[8364]_ , \new_[8367]_ , \new_[8368]_ , \new_[8369]_ ,
    \new_[8373]_ , \new_[8374]_ , \new_[8377]_ , \new_[8380]_ ,
    \new_[8381]_ , \new_[8382]_ , \new_[8386]_ , \new_[8387]_ ,
    \new_[8390]_ , \new_[8393]_ , \new_[8394]_ , \new_[8395]_ ,
    \new_[8399]_ , \new_[8400]_ , \new_[8403]_ , \new_[8406]_ ,
    \new_[8407]_ , \new_[8408]_ , \new_[8412]_ , \new_[8413]_ ,
    \new_[8416]_ , \new_[8419]_ , \new_[8420]_ , \new_[8421]_ ,
    \new_[8425]_ , \new_[8426]_ , \new_[8429]_ , \new_[8432]_ ,
    \new_[8433]_ , \new_[8434]_ , \new_[8438]_ , \new_[8439]_ ,
    \new_[8442]_ , \new_[8445]_ , \new_[8446]_ , \new_[8447]_ ,
    \new_[8451]_ , \new_[8452]_ , \new_[8455]_ , \new_[8458]_ ,
    \new_[8459]_ , \new_[8460]_ , \new_[8464]_ , \new_[8465]_ ,
    \new_[8468]_ , \new_[8471]_ , \new_[8472]_ , \new_[8473]_ ,
    \new_[8477]_ , \new_[8478]_ , \new_[8481]_ , \new_[8484]_ ,
    \new_[8485]_ , \new_[8486]_ , \new_[8490]_ , \new_[8491]_ ,
    \new_[8494]_ , \new_[8497]_ , \new_[8498]_ , \new_[8499]_ ,
    \new_[8503]_ , \new_[8504]_ , \new_[8507]_ , \new_[8510]_ ,
    \new_[8511]_ , \new_[8512]_ , \new_[8516]_ , \new_[8517]_ ,
    \new_[8520]_ , \new_[8523]_ , \new_[8524]_ , \new_[8525]_ ,
    \new_[8529]_ , \new_[8530]_ , \new_[8533]_ , \new_[8536]_ ,
    \new_[8537]_ , \new_[8538]_ , \new_[8542]_ , \new_[8543]_ ,
    \new_[8546]_ , \new_[8549]_ , \new_[8550]_ , \new_[8551]_ ,
    \new_[8555]_ , \new_[8556]_ , \new_[8559]_ , \new_[8562]_ ,
    \new_[8563]_ , \new_[8564]_ , \new_[8568]_ , \new_[8569]_ ,
    \new_[8572]_ , \new_[8575]_ , \new_[8576]_ , \new_[8577]_ ,
    \new_[8581]_ , \new_[8582]_ , \new_[8585]_ , \new_[8588]_ ,
    \new_[8589]_ , \new_[8590]_ , \new_[8594]_ , \new_[8595]_ ,
    \new_[8598]_ , \new_[8601]_ , \new_[8602]_ , \new_[8603]_ ,
    \new_[8607]_ , \new_[8608]_ , \new_[8611]_ , \new_[8614]_ ,
    \new_[8615]_ , \new_[8616]_ , \new_[8620]_ , \new_[8621]_ ,
    \new_[8624]_ , \new_[8627]_ , \new_[8628]_ , \new_[8629]_ ,
    \new_[8633]_ , \new_[8634]_ , \new_[8637]_ , \new_[8640]_ ,
    \new_[8641]_ , \new_[8642]_ , \new_[8646]_ , \new_[8647]_ ,
    \new_[8650]_ , \new_[8653]_ , \new_[8654]_ , \new_[8655]_ ,
    \new_[8659]_ , \new_[8660]_ , \new_[8663]_ , \new_[8666]_ ,
    \new_[8667]_ , \new_[8668]_ , \new_[8672]_ , \new_[8673]_ ,
    \new_[8676]_ , \new_[8679]_ , \new_[8680]_ , \new_[8681]_ ,
    \new_[8685]_ , \new_[8686]_ , \new_[8689]_ , \new_[8692]_ ,
    \new_[8693]_ , \new_[8694]_ , \new_[8698]_ , \new_[8699]_ ,
    \new_[8702]_ , \new_[8705]_ , \new_[8706]_ , \new_[8707]_ ,
    \new_[8711]_ , \new_[8712]_ , \new_[8715]_ , \new_[8718]_ ,
    \new_[8719]_ , \new_[8720]_ , \new_[8724]_ , \new_[8725]_ ,
    \new_[8728]_ , \new_[8731]_ , \new_[8732]_ , \new_[8733]_ ,
    \new_[8737]_ , \new_[8738]_ , \new_[8741]_ , \new_[8744]_ ,
    \new_[8745]_ , \new_[8746]_ , \new_[8750]_ , \new_[8751]_ ,
    \new_[8754]_ , \new_[8757]_ , \new_[8758]_ , \new_[8759]_ ,
    \new_[8763]_ , \new_[8764]_ , \new_[8767]_ , \new_[8770]_ ,
    \new_[8771]_ , \new_[8772]_ , \new_[8776]_ , \new_[8777]_ ,
    \new_[8780]_ , \new_[8783]_ , \new_[8784]_ , \new_[8785]_ ,
    \new_[8789]_ , \new_[8790]_ , \new_[8793]_ , \new_[8796]_ ,
    \new_[8797]_ , \new_[8798]_ , \new_[8802]_ , \new_[8803]_ ,
    \new_[8806]_ , \new_[8809]_ , \new_[8810]_ , \new_[8811]_ ,
    \new_[8815]_ , \new_[8816]_ , \new_[8819]_ , \new_[8822]_ ,
    \new_[8823]_ , \new_[8824]_ , \new_[8828]_ , \new_[8829]_ ,
    \new_[8832]_ , \new_[8835]_ , \new_[8836]_ , \new_[8837]_ ,
    \new_[8841]_ , \new_[8842]_ , \new_[8845]_ , \new_[8848]_ ,
    \new_[8849]_ , \new_[8850]_ , \new_[8854]_ , \new_[8855]_ ,
    \new_[8858]_ , \new_[8861]_ , \new_[8862]_ , \new_[8863]_ ,
    \new_[8867]_ , \new_[8868]_ , \new_[8871]_ , \new_[8874]_ ,
    \new_[8875]_ , \new_[8876]_ , \new_[8880]_ , \new_[8881]_ ,
    \new_[8884]_ , \new_[8887]_ , \new_[8888]_ , \new_[8889]_ ,
    \new_[8893]_ , \new_[8894]_ , \new_[8897]_ , \new_[8900]_ ,
    \new_[8901]_ , \new_[8902]_ , \new_[8906]_ , \new_[8907]_ ,
    \new_[8910]_ , \new_[8913]_ , \new_[8914]_ , \new_[8915]_ ,
    \new_[8919]_ , \new_[8920]_ , \new_[8923]_ , \new_[8926]_ ,
    \new_[8927]_ , \new_[8928]_ , \new_[8932]_ , \new_[8933]_ ,
    \new_[8936]_ , \new_[8939]_ , \new_[8940]_ , \new_[8941]_ ,
    \new_[8945]_ , \new_[8946]_ , \new_[8949]_ , \new_[8952]_ ,
    \new_[8953]_ , \new_[8954]_ , \new_[8958]_ , \new_[8959]_ ,
    \new_[8962]_ , \new_[8965]_ , \new_[8966]_ , \new_[8967]_ ,
    \new_[8971]_ , \new_[8972]_ , \new_[8975]_ , \new_[8978]_ ,
    \new_[8979]_ , \new_[8980]_ , \new_[8984]_ , \new_[8985]_ ,
    \new_[8988]_ , \new_[8991]_ , \new_[8992]_ , \new_[8993]_ ,
    \new_[8997]_ , \new_[8998]_ , \new_[9001]_ , \new_[9004]_ ,
    \new_[9005]_ , \new_[9006]_ , \new_[9010]_ , \new_[9011]_ ,
    \new_[9014]_ , \new_[9017]_ , \new_[9018]_ , \new_[9019]_ ,
    \new_[9023]_ , \new_[9024]_ , \new_[9027]_ , \new_[9030]_ ,
    \new_[9031]_ , \new_[9032]_ , \new_[9036]_ , \new_[9037]_ ,
    \new_[9040]_ , \new_[9043]_ , \new_[9044]_ , \new_[9045]_ ,
    \new_[9049]_ , \new_[9050]_ , \new_[9053]_ , \new_[9056]_ ,
    \new_[9057]_ , \new_[9058]_ , \new_[9062]_ , \new_[9063]_ ,
    \new_[9066]_ , \new_[9069]_ , \new_[9070]_ , \new_[9071]_ ,
    \new_[9075]_ , \new_[9076]_ , \new_[9079]_ , \new_[9082]_ ,
    \new_[9083]_ , \new_[9084]_ , \new_[9088]_ , \new_[9089]_ ,
    \new_[9092]_ , \new_[9095]_ , \new_[9096]_ , \new_[9097]_ ,
    \new_[9101]_ , \new_[9102]_ , \new_[9105]_ , \new_[9108]_ ,
    \new_[9109]_ , \new_[9110]_ , \new_[9114]_ , \new_[9115]_ ,
    \new_[9118]_ , \new_[9121]_ , \new_[9122]_ , \new_[9123]_ ,
    \new_[9127]_ , \new_[9128]_ , \new_[9131]_ , \new_[9134]_ ,
    \new_[9135]_ , \new_[9136]_ , \new_[9140]_ , \new_[9141]_ ,
    \new_[9144]_ , \new_[9147]_ , \new_[9148]_ , \new_[9149]_ ,
    \new_[9153]_ , \new_[9154]_ , \new_[9157]_ , \new_[9160]_ ,
    \new_[9161]_ , \new_[9162]_ , \new_[9166]_ , \new_[9167]_ ,
    \new_[9170]_ , \new_[9173]_ , \new_[9174]_ , \new_[9175]_ ,
    \new_[9179]_ , \new_[9180]_ , \new_[9183]_ , \new_[9186]_ ,
    \new_[9187]_ , \new_[9188]_ , \new_[9192]_ , \new_[9193]_ ,
    \new_[9196]_ , \new_[9199]_ , \new_[9200]_ , \new_[9201]_ ,
    \new_[9205]_ , \new_[9206]_ , \new_[9209]_ , \new_[9212]_ ,
    \new_[9213]_ , \new_[9214]_ , \new_[9218]_ , \new_[9219]_ ,
    \new_[9222]_ , \new_[9225]_ , \new_[9226]_ , \new_[9227]_ ,
    \new_[9231]_ , \new_[9232]_ , \new_[9235]_ , \new_[9238]_ ,
    \new_[9239]_ , \new_[9240]_ , \new_[9244]_ , \new_[9245]_ ,
    \new_[9248]_ , \new_[9251]_ , \new_[9252]_ , \new_[9253]_ ,
    \new_[9257]_ , \new_[9258]_ , \new_[9261]_ , \new_[9264]_ ,
    \new_[9265]_ , \new_[9266]_ , \new_[9270]_ , \new_[9271]_ ,
    \new_[9274]_ , \new_[9277]_ , \new_[9278]_ , \new_[9279]_ ,
    \new_[9283]_ , \new_[9284]_ , \new_[9287]_ , \new_[9290]_ ,
    \new_[9291]_ , \new_[9292]_ , \new_[9296]_ , \new_[9297]_ ,
    \new_[9300]_ , \new_[9303]_ , \new_[9304]_ , \new_[9305]_ ,
    \new_[9309]_ , \new_[9310]_ , \new_[9313]_ , \new_[9316]_ ,
    \new_[9317]_ , \new_[9318]_ , \new_[9322]_ , \new_[9323]_ ,
    \new_[9326]_ , \new_[9329]_ , \new_[9330]_ , \new_[9331]_ ,
    \new_[9335]_ , \new_[9336]_ , \new_[9339]_ , \new_[9342]_ ,
    \new_[9343]_ , \new_[9344]_ , \new_[9348]_ , \new_[9349]_ ,
    \new_[9352]_ , \new_[9355]_ , \new_[9356]_ , \new_[9357]_ ,
    \new_[9361]_ , \new_[9362]_ , \new_[9365]_ , \new_[9368]_ ,
    \new_[9369]_ , \new_[9370]_ , \new_[9374]_ , \new_[9375]_ ,
    \new_[9378]_ , \new_[9381]_ , \new_[9382]_ , \new_[9383]_ ,
    \new_[9387]_ , \new_[9388]_ , \new_[9391]_ , \new_[9394]_ ,
    \new_[9395]_ , \new_[9396]_ , \new_[9400]_ , \new_[9401]_ ,
    \new_[9404]_ , \new_[9407]_ , \new_[9408]_ , \new_[9409]_ ,
    \new_[9413]_ , \new_[9414]_ , \new_[9417]_ , \new_[9420]_ ,
    \new_[9421]_ , \new_[9422]_ , \new_[9426]_ , \new_[9427]_ ,
    \new_[9430]_ , \new_[9433]_ , \new_[9434]_ , \new_[9435]_ ,
    \new_[9439]_ , \new_[9440]_ , \new_[9443]_ , \new_[9446]_ ,
    \new_[9447]_ , \new_[9448]_ , \new_[9452]_ , \new_[9453]_ ,
    \new_[9456]_ , \new_[9459]_ , \new_[9460]_ , \new_[9461]_ ,
    \new_[9465]_ , \new_[9466]_ , \new_[9469]_ , \new_[9472]_ ,
    \new_[9473]_ , \new_[9474]_ , \new_[9478]_ , \new_[9479]_ ,
    \new_[9482]_ , \new_[9485]_ , \new_[9486]_ , \new_[9487]_ ,
    \new_[9491]_ , \new_[9492]_ , \new_[9495]_ , \new_[9498]_ ,
    \new_[9499]_ , \new_[9500]_ , \new_[9504]_ , \new_[9505]_ ,
    \new_[9508]_ , \new_[9511]_ , \new_[9512]_ , \new_[9513]_ ,
    \new_[9517]_ , \new_[9518]_ , \new_[9521]_ , \new_[9524]_ ,
    \new_[9525]_ , \new_[9526]_ , \new_[9530]_ , \new_[9531]_ ,
    \new_[9534]_ , \new_[9537]_ , \new_[9538]_ , \new_[9539]_ ,
    \new_[9543]_ , \new_[9544]_ , \new_[9547]_ , \new_[9550]_ ,
    \new_[9551]_ , \new_[9552]_ , \new_[9556]_ , \new_[9557]_ ,
    \new_[9560]_ , \new_[9563]_ , \new_[9564]_ , \new_[9565]_ ,
    \new_[9569]_ , \new_[9570]_ , \new_[9573]_ , \new_[9576]_ ,
    \new_[9577]_ , \new_[9578]_ , \new_[9582]_ , \new_[9583]_ ,
    \new_[9586]_ , \new_[9589]_ , \new_[9590]_ , \new_[9591]_ ,
    \new_[9595]_ , \new_[9596]_ , \new_[9599]_ , \new_[9602]_ ,
    \new_[9603]_ , \new_[9604]_ , \new_[9608]_ , \new_[9609]_ ,
    \new_[9612]_ , \new_[9615]_ , \new_[9616]_ , \new_[9617]_ ,
    \new_[9621]_ , \new_[9622]_ , \new_[9625]_ , \new_[9628]_ ,
    \new_[9629]_ , \new_[9630]_ , \new_[9634]_ , \new_[9635]_ ,
    \new_[9638]_ , \new_[9641]_ , \new_[9642]_ , \new_[9643]_ ,
    \new_[9647]_ , \new_[9648]_ , \new_[9651]_ , \new_[9654]_ ,
    \new_[9655]_ , \new_[9656]_ , \new_[9660]_ , \new_[9661]_ ,
    \new_[9664]_ , \new_[9667]_ , \new_[9668]_ , \new_[9669]_ ,
    \new_[9673]_ , \new_[9674]_ , \new_[9677]_ , \new_[9680]_ ,
    \new_[9681]_ , \new_[9682]_ , \new_[9686]_ , \new_[9687]_ ,
    \new_[9690]_ , \new_[9693]_ , \new_[9694]_ , \new_[9695]_ ,
    \new_[9699]_ , \new_[9700]_ , \new_[9703]_ , \new_[9706]_ ,
    \new_[9707]_ , \new_[9708]_ , \new_[9712]_ , \new_[9713]_ ,
    \new_[9716]_ , \new_[9719]_ , \new_[9720]_ , \new_[9721]_ ,
    \new_[9725]_ , \new_[9726]_ , \new_[9729]_ , \new_[9732]_ ,
    \new_[9733]_ , \new_[9734]_ , \new_[9738]_ , \new_[9739]_ ,
    \new_[9742]_ , \new_[9745]_ , \new_[9746]_ , \new_[9747]_ ,
    \new_[9751]_ , \new_[9752]_ , \new_[9755]_ , \new_[9758]_ ,
    \new_[9759]_ , \new_[9760]_ , \new_[9764]_ , \new_[9765]_ ,
    \new_[9768]_ , \new_[9771]_ , \new_[9772]_ , \new_[9773]_ ,
    \new_[9777]_ , \new_[9778]_ , \new_[9781]_ , \new_[9784]_ ,
    \new_[9785]_ , \new_[9786]_ , \new_[9790]_ , \new_[9791]_ ,
    \new_[9794]_ , \new_[9797]_ , \new_[9798]_ , \new_[9799]_ ,
    \new_[9803]_ , \new_[9804]_ , \new_[9807]_ , \new_[9810]_ ,
    \new_[9811]_ , \new_[9812]_ , \new_[9816]_ , \new_[9817]_ ,
    \new_[9820]_ , \new_[9823]_ , \new_[9824]_ , \new_[9825]_ ,
    \new_[9829]_ , \new_[9830]_ , \new_[9833]_ , \new_[9836]_ ,
    \new_[9837]_ , \new_[9838]_ , \new_[9842]_ , \new_[9843]_ ,
    \new_[9846]_ , \new_[9849]_ , \new_[9850]_ , \new_[9851]_ ,
    \new_[9855]_ , \new_[9856]_ , \new_[9859]_ , \new_[9862]_ ,
    \new_[9863]_ , \new_[9864]_ , \new_[9868]_ , \new_[9869]_ ,
    \new_[9872]_ , \new_[9875]_ , \new_[9876]_ , \new_[9877]_ ,
    \new_[9881]_ , \new_[9882]_ , \new_[9885]_ , \new_[9888]_ ,
    \new_[9889]_ , \new_[9890]_ , \new_[9894]_ , \new_[9895]_ ,
    \new_[9898]_ , \new_[9901]_ , \new_[9902]_ , \new_[9903]_ ,
    \new_[9907]_ , \new_[9908]_ , \new_[9911]_ , \new_[9914]_ ,
    \new_[9915]_ , \new_[9916]_ , \new_[9920]_ , \new_[9921]_ ,
    \new_[9924]_ , \new_[9927]_ , \new_[9928]_ , \new_[9929]_ ,
    \new_[9933]_ , \new_[9934]_ , \new_[9937]_ , \new_[9940]_ ,
    \new_[9941]_ , \new_[9942]_ , \new_[9946]_ , \new_[9947]_ ,
    \new_[9950]_ , \new_[9953]_ , \new_[9954]_ , \new_[9955]_ ,
    \new_[9959]_ , \new_[9960]_ , \new_[9963]_ , \new_[9966]_ ,
    \new_[9967]_ , \new_[9968]_ , \new_[9972]_ , \new_[9973]_ ,
    \new_[9976]_ , \new_[9979]_ , \new_[9980]_ , \new_[9981]_ ,
    \new_[9985]_ , \new_[9986]_ , \new_[9989]_ , \new_[9992]_ ,
    \new_[9993]_ , \new_[9994]_ , \new_[9998]_ , \new_[9999]_ ,
    \new_[10002]_ , \new_[10005]_ , \new_[10006]_ , \new_[10007]_ ,
    \new_[10011]_ , \new_[10012]_ , \new_[10015]_ , \new_[10018]_ ,
    \new_[10019]_ , \new_[10020]_ , \new_[10024]_ , \new_[10025]_ ,
    \new_[10028]_ , \new_[10031]_ , \new_[10032]_ , \new_[10033]_ ,
    \new_[10037]_ , \new_[10038]_ , \new_[10041]_ , \new_[10044]_ ,
    \new_[10045]_ , \new_[10046]_ , \new_[10050]_ , \new_[10051]_ ,
    \new_[10054]_ , \new_[10057]_ , \new_[10058]_ , \new_[10059]_ ,
    \new_[10063]_ , \new_[10064]_ , \new_[10067]_ , \new_[10070]_ ,
    \new_[10071]_ , \new_[10072]_ , \new_[10076]_ , \new_[10077]_ ,
    \new_[10080]_ , \new_[10083]_ , \new_[10084]_ , \new_[10085]_ ,
    \new_[10089]_ , \new_[10090]_ , \new_[10093]_ , \new_[10096]_ ,
    \new_[10097]_ , \new_[10098]_ , \new_[10102]_ , \new_[10103]_ ,
    \new_[10106]_ , \new_[10109]_ , \new_[10110]_ , \new_[10111]_ ,
    \new_[10115]_ , \new_[10116]_ , \new_[10119]_ , \new_[10122]_ ,
    \new_[10123]_ , \new_[10124]_ , \new_[10128]_ , \new_[10129]_ ,
    \new_[10132]_ , \new_[10135]_ , \new_[10136]_ , \new_[10137]_ ,
    \new_[10141]_ , \new_[10142]_ , \new_[10145]_ , \new_[10148]_ ,
    \new_[10149]_ , \new_[10150]_ , \new_[10154]_ , \new_[10155]_ ,
    \new_[10158]_ , \new_[10161]_ , \new_[10162]_ , \new_[10163]_ ,
    \new_[10167]_ , \new_[10168]_ , \new_[10171]_ , \new_[10174]_ ,
    \new_[10175]_ , \new_[10176]_ , \new_[10180]_ , \new_[10181]_ ,
    \new_[10184]_ , \new_[10187]_ , \new_[10188]_ , \new_[10189]_ ,
    \new_[10193]_ , \new_[10194]_ , \new_[10197]_ , \new_[10200]_ ,
    \new_[10201]_ , \new_[10202]_ , \new_[10206]_ , \new_[10207]_ ,
    \new_[10210]_ , \new_[10213]_ , \new_[10214]_ , \new_[10215]_ ,
    \new_[10219]_ , \new_[10220]_ , \new_[10223]_ , \new_[10226]_ ,
    \new_[10227]_ , \new_[10228]_ , \new_[10232]_ , \new_[10233]_ ,
    \new_[10236]_ , \new_[10239]_ , \new_[10240]_ , \new_[10241]_ ,
    \new_[10245]_ , \new_[10246]_ , \new_[10249]_ , \new_[10252]_ ,
    \new_[10253]_ , \new_[10254]_ , \new_[10258]_ , \new_[10259]_ ,
    \new_[10262]_ , \new_[10265]_ , \new_[10266]_ , \new_[10267]_ ,
    \new_[10271]_ , \new_[10272]_ , \new_[10275]_ , \new_[10278]_ ,
    \new_[10279]_ , \new_[10280]_ , \new_[10284]_ , \new_[10285]_ ,
    \new_[10288]_ , \new_[10291]_ , \new_[10292]_ , \new_[10293]_ ,
    \new_[10297]_ , \new_[10298]_ , \new_[10301]_ , \new_[10304]_ ,
    \new_[10305]_ , \new_[10306]_ , \new_[10310]_ , \new_[10311]_ ,
    \new_[10314]_ , \new_[10317]_ , \new_[10318]_ , \new_[10319]_ ,
    \new_[10323]_ , \new_[10324]_ , \new_[10327]_ , \new_[10330]_ ,
    \new_[10331]_ , \new_[10332]_ , \new_[10336]_ , \new_[10337]_ ,
    \new_[10340]_ , \new_[10343]_ , \new_[10344]_ , \new_[10345]_ ,
    \new_[10349]_ , \new_[10350]_ , \new_[10353]_ , \new_[10356]_ ,
    \new_[10357]_ , \new_[10358]_ , \new_[10362]_ , \new_[10363]_ ,
    \new_[10366]_ , \new_[10369]_ , \new_[10370]_ , \new_[10371]_ ,
    \new_[10375]_ , \new_[10376]_ , \new_[10379]_ , \new_[10382]_ ,
    \new_[10383]_ , \new_[10384]_ , \new_[10388]_ , \new_[10389]_ ,
    \new_[10392]_ , \new_[10395]_ , \new_[10396]_ , \new_[10397]_ ,
    \new_[10401]_ , \new_[10402]_ , \new_[10405]_ , \new_[10408]_ ,
    \new_[10409]_ , \new_[10410]_ , \new_[10414]_ , \new_[10415]_ ,
    \new_[10418]_ , \new_[10421]_ , \new_[10422]_ , \new_[10423]_ ,
    \new_[10427]_ , \new_[10428]_ , \new_[10431]_ , \new_[10434]_ ,
    \new_[10435]_ , \new_[10436]_ , \new_[10440]_ , \new_[10441]_ ,
    \new_[10444]_ , \new_[10447]_ , \new_[10448]_ , \new_[10449]_ ,
    \new_[10453]_ , \new_[10454]_ , \new_[10457]_ , \new_[10460]_ ,
    \new_[10461]_ , \new_[10462]_ , \new_[10466]_ , \new_[10467]_ ,
    \new_[10470]_ , \new_[10473]_ , \new_[10474]_ , \new_[10475]_ ,
    \new_[10479]_ , \new_[10480]_ , \new_[10483]_ , \new_[10486]_ ,
    \new_[10487]_ , \new_[10488]_ , \new_[10492]_ , \new_[10493]_ ,
    \new_[10496]_ , \new_[10499]_ , \new_[10500]_ , \new_[10501]_ ,
    \new_[10505]_ , \new_[10506]_ , \new_[10509]_ , \new_[10512]_ ,
    \new_[10513]_ , \new_[10514]_ , \new_[10518]_ , \new_[10519]_ ,
    \new_[10522]_ , \new_[10525]_ , \new_[10526]_ , \new_[10527]_ ,
    \new_[10531]_ , \new_[10532]_ , \new_[10535]_ , \new_[10538]_ ,
    \new_[10539]_ , \new_[10540]_ , \new_[10544]_ , \new_[10545]_ ,
    \new_[10548]_ , \new_[10551]_ , \new_[10552]_ , \new_[10553]_ ,
    \new_[10557]_ , \new_[10558]_ , \new_[10561]_ , \new_[10564]_ ,
    \new_[10565]_ , \new_[10566]_ , \new_[10570]_ , \new_[10571]_ ,
    \new_[10574]_ , \new_[10577]_ , \new_[10578]_ , \new_[10579]_ ,
    \new_[10583]_ , \new_[10584]_ , \new_[10587]_ , \new_[10590]_ ,
    \new_[10591]_ , \new_[10592]_ , \new_[10596]_ , \new_[10597]_ ,
    \new_[10600]_ , \new_[10603]_ , \new_[10604]_ , \new_[10605]_ ,
    \new_[10609]_ , \new_[10610]_ , \new_[10613]_ , \new_[10616]_ ,
    \new_[10617]_ , \new_[10618]_ , \new_[10622]_ , \new_[10623]_ ,
    \new_[10626]_ , \new_[10629]_ , \new_[10630]_ , \new_[10631]_ ,
    \new_[10635]_ , \new_[10636]_ , \new_[10639]_ , \new_[10642]_ ,
    \new_[10643]_ , \new_[10644]_ , \new_[10648]_ , \new_[10649]_ ,
    \new_[10652]_ , \new_[10655]_ , \new_[10656]_ , \new_[10657]_ ,
    \new_[10661]_ , \new_[10662]_ , \new_[10665]_ , \new_[10668]_ ,
    \new_[10669]_ , \new_[10670]_ , \new_[10674]_ , \new_[10675]_ ,
    \new_[10678]_ , \new_[10681]_ , \new_[10682]_ , \new_[10683]_ ,
    \new_[10687]_ , \new_[10688]_ , \new_[10691]_ , \new_[10694]_ ,
    \new_[10695]_ , \new_[10696]_ , \new_[10700]_ , \new_[10701]_ ,
    \new_[10704]_ , \new_[10707]_ , \new_[10708]_ , \new_[10709]_ ,
    \new_[10713]_ , \new_[10714]_ , \new_[10717]_ , \new_[10720]_ ,
    \new_[10721]_ , \new_[10722]_ , \new_[10726]_ , \new_[10727]_ ,
    \new_[10730]_ , \new_[10733]_ , \new_[10734]_ , \new_[10735]_ ,
    \new_[10739]_ , \new_[10740]_ , \new_[10743]_ , \new_[10746]_ ,
    \new_[10747]_ , \new_[10748]_ , \new_[10752]_ , \new_[10753]_ ,
    \new_[10756]_ , \new_[10759]_ , \new_[10760]_ , \new_[10761]_ ,
    \new_[10765]_ , \new_[10766]_ , \new_[10769]_ , \new_[10772]_ ,
    \new_[10773]_ , \new_[10774]_ , \new_[10778]_ , \new_[10779]_ ,
    \new_[10782]_ , \new_[10785]_ , \new_[10786]_ , \new_[10787]_ ,
    \new_[10791]_ , \new_[10792]_ , \new_[10795]_ , \new_[10798]_ ,
    \new_[10799]_ , \new_[10800]_ , \new_[10804]_ , \new_[10805]_ ,
    \new_[10808]_ , \new_[10811]_ , \new_[10812]_ , \new_[10813]_ ,
    \new_[10817]_ , \new_[10818]_ , \new_[10821]_ , \new_[10824]_ ,
    \new_[10825]_ , \new_[10826]_ , \new_[10830]_ , \new_[10831]_ ,
    \new_[10834]_ , \new_[10837]_ , \new_[10838]_ , \new_[10839]_ ,
    \new_[10843]_ , \new_[10844]_ , \new_[10847]_ , \new_[10850]_ ,
    \new_[10851]_ , \new_[10852]_ , \new_[10856]_ , \new_[10857]_ ,
    \new_[10860]_ , \new_[10863]_ , \new_[10864]_ , \new_[10865]_ ,
    \new_[10869]_ , \new_[10870]_ , \new_[10873]_ , \new_[10876]_ ,
    \new_[10877]_ , \new_[10878]_ , \new_[10882]_ , \new_[10883]_ ,
    \new_[10886]_ , \new_[10889]_ , \new_[10890]_ , \new_[10891]_ ,
    \new_[10895]_ , \new_[10896]_ , \new_[10899]_ , \new_[10902]_ ,
    \new_[10903]_ , \new_[10904]_ , \new_[10908]_ , \new_[10909]_ ,
    \new_[10912]_ , \new_[10915]_ , \new_[10916]_ , \new_[10917]_ ,
    \new_[10921]_ , \new_[10922]_ , \new_[10925]_ , \new_[10928]_ ,
    \new_[10929]_ , \new_[10930]_ , \new_[10934]_ , \new_[10935]_ ,
    \new_[10938]_ , \new_[10941]_ , \new_[10942]_ , \new_[10943]_ ,
    \new_[10947]_ , \new_[10948]_ , \new_[10951]_ , \new_[10954]_ ,
    \new_[10955]_ , \new_[10956]_ , \new_[10960]_ , \new_[10961]_ ,
    \new_[10964]_ , \new_[10967]_ , \new_[10968]_ , \new_[10969]_ ,
    \new_[10973]_ , \new_[10974]_ , \new_[10977]_ , \new_[10980]_ ,
    \new_[10981]_ , \new_[10982]_ , \new_[10986]_ , \new_[10987]_ ,
    \new_[10990]_ , \new_[10993]_ , \new_[10994]_ , \new_[10995]_ ,
    \new_[10999]_ , \new_[11000]_ , \new_[11003]_ , \new_[11006]_ ,
    \new_[11007]_ , \new_[11008]_ , \new_[11012]_ , \new_[11013]_ ,
    \new_[11016]_ , \new_[11019]_ , \new_[11020]_ , \new_[11021]_ ,
    \new_[11025]_ , \new_[11026]_ , \new_[11029]_ , \new_[11032]_ ,
    \new_[11033]_ , \new_[11034]_ , \new_[11038]_ , \new_[11039]_ ,
    \new_[11042]_ , \new_[11045]_ , \new_[11046]_ , \new_[11047]_ ,
    \new_[11051]_ , \new_[11052]_ , \new_[11055]_ , \new_[11058]_ ,
    \new_[11059]_ , \new_[11060]_ , \new_[11064]_ , \new_[11065]_ ,
    \new_[11068]_ , \new_[11071]_ , \new_[11072]_ , \new_[11073]_ ,
    \new_[11077]_ , \new_[11078]_ , \new_[11081]_ , \new_[11084]_ ,
    \new_[11085]_ , \new_[11086]_ , \new_[11090]_ , \new_[11091]_ ,
    \new_[11094]_ , \new_[11097]_ , \new_[11098]_ , \new_[11099]_ ,
    \new_[11103]_ , \new_[11104]_ , \new_[11107]_ , \new_[11110]_ ,
    \new_[11111]_ , \new_[11112]_ , \new_[11116]_ , \new_[11117]_ ,
    \new_[11120]_ , \new_[11123]_ , \new_[11124]_ , \new_[11125]_ ,
    \new_[11129]_ , \new_[11130]_ , \new_[11133]_ , \new_[11136]_ ,
    \new_[11137]_ , \new_[11138]_ , \new_[11142]_ , \new_[11143]_ ,
    \new_[11146]_ , \new_[11149]_ , \new_[11150]_ , \new_[11151]_ ,
    \new_[11155]_ , \new_[11156]_ , \new_[11159]_ , \new_[11162]_ ,
    \new_[11163]_ , \new_[11164]_ , \new_[11168]_ , \new_[11169]_ ,
    \new_[11172]_ , \new_[11175]_ , \new_[11176]_ , \new_[11177]_ ,
    \new_[11181]_ , \new_[11182]_ , \new_[11185]_ , \new_[11188]_ ,
    \new_[11189]_ , \new_[11190]_ , \new_[11194]_ , \new_[11195]_ ,
    \new_[11198]_ , \new_[11201]_ , \new_[11202]_ , \new_[11203]_ ,
    \new_[11207]_ , \new_[11208]_ , \new_[11211]_ , \new_[11214]_ ,
    \new_[11215]_ , \new_[11216]_ , \new_[11220]_ , \new_[11221]_ ,
    \new_[11224]_ , \new_[11227]_ , \new_[11228]_ , \new_[11229]_ ,
    \new_[11233]_ , \new_[11234]_ , \new_[11237]_ , \new_[11240]_ ,
    \new_[11241]_ , \new_[11242]_ , \new_[11246]_ , \new_[11247]_ ,
    \new_[11250]_ , \new_[11253]_ , \new_[11254]_ , \new_[11255]_ ,
    \new_[11259]_ , \new_[11260]_ , \new_[11263]_ , \new_[11266]_ ,
    \new_[11267]_ , \new_[11268]_ , \new_[11272]_ , \new_[11273]_ ,
    \new_[11276]_ , \new_[11279]_ , \new_[11280]_ , \new_[11281]_ ,
    \new_[11285]_ , \new_[11286]_ , \new_[11289]_ , \new_[11292]_ ,
    \new_[11293]_ , \new_[11294]_ , \new_[11298]_ , \new_[11299]_ ,
    \new_[11302]_ , \new_[11305]_ , \new_[11306]_ , \new_[11307]_ ,
    \new_[11311]_ , \new_[11312]_ , \new_[11315]_ , \new_[11318]_ ,
    \new_[11319]_ , \new_[11320]_ , \new_[11324]_ , \new_[11325]_ ,
    \new_[11328]_ , \new_[11331]_ , \new_[11332]_ , \new_[11333]_ ,
    \new_[11337]_ , \new_[11338]_ , \new_[11341]_ , \new_[11344]_ ,
    \new_[11345]_ , \new_[11346]_ , \new_[11350]_ , \new_[11351]_ ,
    \new_[11354]_ , \new_[11357]_ , \new_[11358]_ , \new_[11359]_ ,
    \new_[11363]_ , \new_[11364]_ , \new_[11367]_ , \new_[11370]_ ,
    \new_[11371]_ , \new_[11372]_ , \new_[11376]_ , \new_[11377]_ ,
    \new_[11380]_ , \new_[11383]_ , \new_[11384]_ , \new_[11385]_ ,
    \new_[11389]_ , \new_[11390]_ , \new_[11393]_ , \new_[11396]_ ,
    \new_[11397]_ , \new_[11398]_ , \new_[11402]_ , \new_[11403]_ ,
    \new_[11406]_ , \new_[11409]_ , \new_[11410]_ , \new_[11411]_ ,
    \new_[11415]_ , \new_[11416]_ , \new_[11419]_ , \new_[11422]_ ,
    \new_[11423]_ , \new_[11424]_ , \new_[11428]_ , \new_[11429]_ ,
    \new_[11432]_ , \new_[11435]_ , \new_[11436]_ , \new_[11437]_ ,
    \new_[11441]_ , \new_[11442]_ , \new_[11445]_ , \new_[11448]_ ,
    \new_[11449]_ , \new_[11450]_ , \new_[11454]_ , \new_[11455]_ ,
    \new_[11458]_ , \new_[11461]_ , \new_[11462]_ , \new_[11463]_ ,
    \new_[11467]_ , \new_[11468]_ , \new_[11471]_ , \new_[11474]_ ,
    \new_[11475]_ , \new_[11476]_ , \new_[11480]_ , \new_[11481]_ ,
    \new_[11484]_ , \new_[11487]_ , \new_[11488]_ , \new_[11489]_ ,
    \new_[11493]_ , \new_[11494]_ , \new_[11497]_ , \new_[11500]_ ,
    \new_[11501]_ , \new_[11502]_ , \new_[11506]_ , \new_[11507]_ ,
    \new_[11510]_ , \new_[11513]_ , \new_[11514]_ , \new_[11515]_ ,
    \new_[11519]_ , \new_[11520]_ , \new_[11523]_ , \new_[11526]_ ,
    \new_[11527]_ , \new_[11528]_ , \new_[11532]_ , \new_[11533]_ ,
    \new_[11536]_ , \new_[11539]_ , \new_[11540]_ , \new_[11541]_ ,
    \new_[11545]_ , \new_[11546]_ , \new_[11549]_ , \new_[11552]_ ,
    \new_[11553]_ , \new_[11554]_ , \new_[11558]_ , \new_[11559]_ ,
    \new_[11562]_ , \new_[11565]_ , \new_[11566]_ , \new_[11567]_ ,
    \new_[11571]_ , \new_[11572]_ , \new_[11575]_ , \new_[11578]_ ,
    \new_[11579]_ , \new_[11580]_ , \new_[11584]_ , \new_[11585]_ ,
    \new_[11588]_ , \new_[11591]_ , \new_[11592]_ , \new_[11593]_ ,
    \new_[11597]_ , \new_[11598]_ , \new_[11601]_ , \new_[11604]_ ,
    \new_[11605]_ , \new_[11606]_ , \new_[11610]_ , \new_[11611]_ ,
    \new_[11614]_ , \new_[11617]_ , \new_[11618]_ , \new_[11619]_ ,
    \new_[11623]_ , \new_[11624]_ , \new_[11627]_ , \new_[11630]_ ,
    \new_[11631]_ , \new_[11632]_ , \new_[11636]_ , \new_[11637]_ ,
    \new_[11640]_ , \new_[11643]_ , \new_[11644]_ , \new_[11645]_ ,
    \new_[11649]_ , \new_[11650]_ , \new_[11653]_ , \new_[11656]_ ,
    \new_[11657]_ , \new_[11658]_ , \new_[11662]_ , \new_[11663]_ ,
    \new_[11666]_ , \new_[11669]_ , \new_[11670]_ , \new_[11671]_ ,
    \new_[11675]_ , \new_[11676]_ , \new_[11679]_ , \new_[11682]_ ,
    \new_[11683]_ , \new_[11684]_ , \new_[11688]_ , \new_[11689]_ ,
    \new_[11692]_ , \new_[11695]_ , \new_[11696]_ , \new_[11697]_ ,
    \new_[11701]_ , \new_[11702]_ , \new_[11705]_ , \new_[11708]_ ,
    \new_[11709]_ , \new_[11710]_ , \new_[11714]_ , \new_[11715]_ ,
    \new_[11718]_ , \new_[11721]_ , \new_[11722]_ , \new_[11723]_ ,
    \new_[11727]_ , \new_[11728]_ , \new_[11731]_ , \new_[11734]_ ,
    \new_[11735]_ , \new_[11736]_ , \new_[11740]_ , \new_[11741]_ ,
    \new_[11744]_ , \new_[11747]_ , \new_[11748]_ , \new_[11749]_ ,
    \new_[11753]_ , \new_[11754]_ , \new_[11757]_ , \new_[11760]_ ,
    \new_[11761]_ , \new_[11762]_ , \new_[11766]_ , \new_[11767]_ ,
    \new_[11770]_ , \new_[11773]_ , \new_[11774]_ , \new_[11775]_ ,
    \new_[11779]_ , \new_[11780]_ , \new_[11783]_ , \new_[11786]_ ,
    \new_[11787]_ , \new_[11788]_ , \new_[11792]_ , \new_[11793]_ ,
    \new_[11796]_ , \new_[11799]_ , \new_[11800]_ , \new_[11801]_ ,
    \new_[11805]_ , \new_[11806]_ , \new_[11809]_ , \new_[11812]_ ,
    \new_[11813]_ , \new_[11814]_ , \new_[11818]_ , \new_[11819]_ ,
    \new_[11822]_ , \new_[11825]_ , \new_[11826]_ , \new_[11827]_ ,
    \new_[11831]_ , \new_[11832]_ , \new_[11835]_ , \new_[11838]_ ,
    \new_[11839]_ , \new_[11840]_ , \new_[11844]_ , \new_[11845]_ ,
    \new_[11848]_ , \new_[11851]_ , \new_[11852]_ , \new_[11853]_ ,
    \new_[11857]_ , \new_[11858]_ , \new_[11861]_ , \new_[11864]_ ,
    \new_[11865]_ , \new_[11866]_ , \new_[11870]_ , \new_[11871]_ ,
    \new_[11874]_ , \new_[11877]_ , \new_[11878]_ , \new_[11879]_ ,
    \new_[11883]_ , \new_[11884]_ , \new_[11887]_ , \new_[11890]_ ,
    \new_[11891]_ , \new_[11892]_ , \new_[11896]_ , \new_[11897]_ ,
    \new_[11900]_ , \new_[11903]_ , \new_[11904]_ , \new_[11905]_ ,
    \new_[11909]_ , \new_[11910]_ , \new_[11913]_ , \new_[11916]_ ,
    \new_[11917]_ , \new_[11918]_ , \new_[11922]_ , \new_[11923]_ ,
    \new_[11926]_ , \new_[11929]_ , \new_[11930]_ , \new_[11931]_ ,
    \new_[11935]_ , \new_[11936]_ , \new_[11939]_ , \new_[11942]_ ,
    \new_[11943]_ , \new_[11944]_ , \new_[11948]_ , \new_[11949]_ ,
    \new_[11952]_ , \new_[11955]_ , \new_[11956]_ , \new_[11957]_ ,
    \new_[11961]_ , \new_[11962]_ , \new_[11965]_ , \new_[11968]_ ,
    \new_[11969]_ , \new_[11970]_ , \new_[11974]_ , \new_[11975]_ ,
    \new_[11978]_ , \new_[11981]_ , \new_[11982]_ , \new_[11983]_ ,
    \new_[11987]_ , \new_[11988]_ , \new_[11991]_ , \new_[11994]_ ,
    \new_[11995]_ , \new_[11996]_ , \new_[12000]_ , \new_[12001]_ ,
    \new_[12004]_ , \new_[12007]_ , \new_[12008]_ , \new_[12009]_ ,
    \new_[12013]_ , \new_[12014]_ , \new_[12017]_ , \new_[12020]_ ,
    \new_[12021]_ , \new_[12022]_ , \new_[12026]_ , \new_[12027]_ ,
    \new_[12030]_ , \new_[12033]_ , \new_[12034]_ , \new_[12035]_ ,
    \new_[12039]_ , \new_[12040]_ , \new_[12043]_ , \new_[12046]_ ,
    \new_[12047]_ , \new_[12048]_ , \new_[12052]_ , \new_[12053]_ ,
    \new_[12056]_ , \new_[12059]_ , \new_[12060]_ , \new_[12061]_ ,
    \new_[12065]_ , \new_[12066]_ , \new_[12069]_ , \new_[12072]_ ,
    \new_[12073]_ , \new_[12074]_ , \new_[12078]_ , \new_[12079]_ ,
    \new_[12082]_ , \new_[12085]_ , \new_[12086]_ , \new_[12087]_ ,
    \new_[12091]_ , \new_[12092]_ , \new_[12095]_ , \new_[12098]_ ,
    \new_[12099]_ , \new_[12100]_ , \new_[12104]_ , \new_[12105]_ ,
    \new_[12108]_ , \new_[12111]_ , \new_[12112]_ , \new_[12113]_ ,
    \new_[12117]_ , \new_[12118]_ , \new_[12121]_ , \new_[12124]_ ,
    \new_[12125]_ , \new_[12126]_ , \new_[12130]_ , \new_[12131]_ ,
    \new_[12134]_ , \new_[12137]_ , \new_[12138]_ , \new_[12139]_ ,
    \new_[12143]_ , \new_[12144]_ , \new_[12147]_ , \new_[12150]_ ,
    \new_[12151]_ , \new_[12152]_ , \new_[12156]_ , \new_[12157]_ ,
    \new_[12160]_ , \new_[12163]_ , \new_[12164]_ , \new_[12165]_ ,
    \new_[12169]_ , \new_[12170]_ , \new_[12173]_ , \new_[12176]_ ,
    \new_[12177]_ , \new_[12178]_ , \new_[12182]_ , \new_[12183]_ ,
    \new_[12186]_ , \new_[12189]_ , \new_[12190]_ , \new_[12191]_ ,
    \new_[12195]_ , \new_[12196]_ , \new_[12199]_ , \new_[12202]_ ,
    \new_[12203]_ , \new_[12204]_ , \new_[12208]_ , \new_[12209]_ ,
    \new_[12212]_ , \new_[12215]_ , \new_[12216]_ , \new_[12217]_ ,
    \new_[12221]_ , \new_[12222]_ , \new_[12225]_ , \new_[12228]_ ,
    \new_[12229]_ , \new_[12230]_ , \new_[12234]_ , \new_[12235]_ ,
    \new_[12238]_ , \new_[12241]_ , \new_[12242]_ , \new_[12243]_ ,
    \new_[12247]_ , \new_[12248]_ , \new_[12251]_ , \new_[12254]_ ,
    \new_[12255]_ , \new_[12256]_ , \new_[12260]_ , \new_[12261]_ ,
    \new_[12264]_ , \new_[12267]_ , \new_[12268]_ , \new_[12269]_ ,
    \new_[12273]_ , \new_[12274]_ , \new_[12277]_ , \new_[12280]_ ,
    \new_[12281]_ , \new_[12282]_ , \new_[12286]_ , \new_[12287]_ ,
    \new_[12290]_ , \new_[12293]_ , \new_[12294]_ , \new_[12295]_ ,
    \new_[12299]_ , \new_[12300]_ , \new_[12303]_ , \new_[12306]_ ,
    \new_[12307]_ , \new_[12308]_ , \new_[12312]_ , \new_[12313]_ ,
    \new_[12316]_ , \new_[12319]_ , \new_[12320]_ , \new_[12321]_ ,
    \new_[12325]_ , \new_[12326]_ , \new_[12329]_ , \new_[12332]_ ,
    \new_[12333]_ , \new_[12334]_ , \new_[12338]_ , \new_[12339]_ ,
    \new_[12342]_ , \new_[12345]_ , \new_[12346]_ , \new_[12347]_ ,
    \new_[12351]_ , \new_[12352]_ , \new_[12355]_ , \new_[12358]_ ,
    \new_[12359]_ , \new_[12360]_ , \new_[12364]_ , \new_[12365]_ ,
    \new_[12368]_ , \new_[12371]_ , \new_[12372]_ , \new_[12373]_ ,
    \new_[12377]_ , \new_[12378]_ , \new_[12381]_ , \new_[12384]_ ,
    \new_[12385]_ , \new_[12386]_ , \new_[12390]_ , \new_[12391]_ ,
    \new_[12394]_ , \new_[12397]_ , \new_[12398]_ , \new_[12399]_ ,
    \new_[12403]_ , \new_[12404]_ , \new_[12407]_ , \new_[12410]_ ,
    \new_[12411]_ , \new_[12412]_ , \new_[12416]_ , \new_[12417]_ ,
    \new_[12420]_ , \new_[12423]_ , \new_[12424]_ , \new_[12425]_ ,
    \new_[12429]_ , \new_[12430]_ , \new_[12433]_ , \new_[12436]_ ,
    \new_[12437]_ , \new_[12438]_ , \new_[12442]_ , \new_[12443]_ ,
    \new_[12446]_ , \new_[12449]_ , \new_[12450]_ , \new_[12451]_ ,
    \new_[12455]_ , \new_[12456]_ , \new_[12459]_ , \new_[12462]_ ,
    \new_[12463]_ , \new_[12464]_ , \new_[12468]_ , \new_[12469]_ ,
    \new_[12472]_ , \new_[12475]_ , \new_[12476]_ , \new_[12477]_ ,
    \new_[12481]_ , \new_[12482]_ , \new_[12485]_ , \new_[12488]_ ,
    \new_[12489]_ , \new_[12490]_ , \new_[12494]_ , \new_[12495]_ ,
    \new_[12498]_ , \new_[12501]_ , \new_[12502]_ , \new_[12503]_ ,
    \new_[12507]_ , \new_[12508]_ , \new_[12511]_ , \new_[12514]_ ,
    \new_[12515]_ , \new_[12516]_ , \new_[12520]_ , \new_[12521]_ ,
    \new_[12524]_ , \new_[12527]_ , \new_[12528]_ , \new_[12529]_ ,
    \new_[12533]_ , \new_[12534]_ , \new_[12537]_ , \new_[12540]_ ,
    \new_[12541]_ , \new_[12542]_ , \new_[12546]_ , \new_[12547]_ ,
    \new_[12550]_ , \new_[12553]_ , \new_[12554]_ , \new_[12555]_ ,
    \new_[12559]_ , \new_[12560]_ , \new_[12563]_ , \new_[12566]_ ,
    \new_[12567]_ , \new_[12568]_ , \new_[12572]_ , \new_[12573]_ ,
    \new_[12576]_ , \new_[12579]_ , \new_[12580]_ , \new_[12581]_ ,
    \new_[12585]_ , \new_[12586]_ , \new_[12589]_ , \new_[12592]_ ,
    \new_[12593]_ , \new_[12594]_ , \new_[12598]_ , \new_[12599]_ ,
    \new_[12602]_ , \new_[12605]_ , \new_[12606]_ , \new_[12607]_ ,
    \new_[12611]_ , \new_[12612]_ , \new_[12615]_ , \new_[12618]_ ,
    \new_[12619]_ , \new_[12620]_ , \new_[12624]_ , \new_[12625]_ ,
    \new_[12628]_ , \new_[12631]_ , \new_[12632]_ , \new_[12633]_ ,
    \new_[12637]_ , \new_[12638]_ , \new_[12641]_ , \new_[12644]_ ,
    \new_[12645]_ , \new_[12646]_ , \new_[12650]_ , \new_[12651]_ ,
    \new_[12654]_ , \new_[12657]_ , \new_[12658]_ , \new_[12659]_ ,
    \new_[12663]_ , \new_[12664]_ , \new_[12667]_ , \new_[12670]_ ,
    \new_[12671]_ , \new_[12672]_ , \new_[12676]_ , \new_[12677]_ ,
    \new_[12680]_ , \new_[12683]_ , \new_[12684]_ , \new_[12685]_ ,
    \new_[12689]_ , \new_[12690]_ , \new_[12693]_ , \new_[12696]_ ,
    \new_[12697]_ , \new_[12698]_ , \new_[12702]_ , \new_[12703]_ ,
    \new_[12706]_ , \new_[12709]_ , \new_[12710]_ , \new_[12711]_ ,
    \new_[12715]_ , \new_[12716]_ , \new_[12719]_ , \new_[12722]_ ,
    \new_[12723]_ , \new_[12724]_ , \new_[12728]_ , \new_[12729]_ ,
    \new_[12732]_ , \new_[12735]_ , \new_[12736]_ , \new_[12737]_ ,
    \new_[12741]_ , \new_[12742]_ , \new_[12745]_ , \new_[12748]_ ,
    \new_[12749]_ , \new_[12750]_ , \new_[12754]_ , \new_[12755]_ ,
    \new_[12758]_ , \new_[12761]_ , \new_[12762]_ , \new_[12763]_ ,
    \new_[12767]_ , \new_[12768]_ , \new_[12771]_ , \new_[12774]_ ,
    \new_[12775]_ , \new_[12776]_ , \new_[12780]_ , \new_[12781]_ ,
    \new_[12784]_ , \new_[12787]_ , \new_[12788]_ , \new_[12789]_ ,
    \new_[12793]_ , \new_[12794]_ , \new_[12797]_ , \new_[12800]_ ,
    \new_[12801]_ , \new_[12802]_ , \new_[12806]_ , \new_[12807]_ ,
    \new_[12810]_ , \new_[12813]_ , \new_[12814]_ , \new_[12815]_ ,
    \new_[12819]_ , \new_[12820]_ , \new_[12823]_ , \new_[12826]_ ,
    \new_[12827]_ , \new_[12828]_ , \new_[12832]_ , \new_[12833]_ ,
    \new_[12836]_ , \new_[12839]_ , \new_[12840]_ , \new_[12841]_ ,
    \new_[12845]_ , \new_[12846]_ , \new_[12849]_ , \new_[12852]_ ,
    \new_[12853]_ , \new_[12854]_ , \new_[12858]_ , \new_[12859]_ ,
    \new_[12862]_ , \new_[12865]_ , \new_[12866]_ , \new_[12867]_ ,
    \new_[12871]_ , \new_[12872]_ , \new_[12875]_ , \new_[12878]_ ,
    \new_[12879]_ , \new_[12880]_ , \new_[12884]_ , \new_[12885]_ ,
    \new_[12888]_ , \new_[12891]_ , \new_[12892]_ , \new_[12893]_ ,
    \new_[12897]_ , \new_[12898]_ , \new_[12901]_ , \new_[12904]_ ,
    \new_[12905]_ , \new_[12906]_ , \new_[12910]_ , \new_[12911]_ ,
    \new_[12914]_ , \new_[12917]_ , \new_[12918]_ , \new_[12919]_ ,
    \new_[12923]_ , \new_[12924]_ , \new_[12927]_ , \new_[12930]_ ,
    \new_[12931]_ , \new_[12932]_ , \new_[12936]_ , \new_[12937]_ ,
    \new_[12940]_ , \new_[12943]_ , \new_[12944]_ , \new_[12945]_ ,
    \new_[12949]_ , \new_[12950]_ , \new_[12953]_ , \new_[12956]_ ,
    \new_[12957]_ , \new_[12958]_ , \new_[12962]_ , \new_[12963]_ ,
    \new_[12966]_ , \new_[12969]_ , \new_[12970]_ , \new_[12971]_ ,
    \new_[12975]_ , \new_[12976]_ , \new_[12979]_ , \new_[12982]_ ,
    \new_[12983]_ , \new_[12984]_ , \new_[12988]_ , \new_[12989]_ ,
    \new_[12992]_ , \new_[12995]_ , \new_[12996]_ , \new_[12997]_ ,
    \new_[13001]_ , \new_[13002]_ , \new_[13005]_ , \new_[13008]_ ,
    \new_[13009]_ , \new_[13010]_ , \new_[13014]_ , \new_[13015]_ ,
    \new_[13018]_ , \new_[13021]_ , \new_[13022]_ , \new_[13023]_ ,
    \new_[13027]_ , \new_[13028]_ , \new_[13031]_ , \new_[13034]_ ,
    \new_[13035]_ , \new_[13036]_ , \new_[13040]_ , \new_[13041]_ ,
    \new_[13044]_ , \new_[13047]_ , \new_[13048]_ , \new_[13049]_ ,
    \new_[13053]_ , \new_[13054]_ , \new_[13057]_ , \new_[13060]_ ,
    \new_[13061]_ , \new_[13062]_ , \new_[13066]_ , \new_[13067]_ ,
    \new_[13070]_ , \new_[13073]_ , \new_[13074]_ , \new_[13075]_ ,
    \new_[13079]_ , \new_[13080]_ , \new_[13083]_ , \new_[13086]_ ,
    \new_[13087]_ , \new_[13088]_ , \new_[13092]_ , \new_[13093]_ ,
    \new_[13096]_ , \new_[13099]_ , \new_[13100]_ , \new_[13101]_ ,
    \new_[13105]_ , \new_[13106]_ , \new_[13109]_ , \new_[13112]_ ,
    \new_[13113]_ , \new_[13114]_ , \new_[13118]_ , \new_[13119]_ ,
    \new_[13122]_ , \new_[13125]_ , \new_[13126]_ , \new_[13127]_ ,
    \new_[13131]_ , \new_[13132]_ , \new_[13135]_ , \new_[13138]_ ,
    \new_[13139]_ , \new_[13140]_ , \new_[13144]_ , \new_[13145]_ ,
    \new_[13148]_ , \new_[13151]_ , \new_[13152]_ , \new_[13153]_ ,
    \new_[13157]_ , \new_[13158]_ , \new_[13161]_ , \new_[13164]_ ,
    \new_[13165]_ , \new_[13166]_ , \new_[13170]_ , \new_[13171]_ ,
    \new_[13174]_ , \new_[13177]_ , \new_[13178]_ , \new_[13179]_ ,
    \new_[13183]_ , \new_[13184]_ , \new_[13187]_ , \new_[13190]_ ,
    \new_[13191]_ , \new_[13192]_ , \new_[13196]_ , \new_[13197]_ ,
    \new_[13200]_ , \new_[13203]_ , \new_[13204]_ , \new_[13205]_ ,
    \new_[13209]_ , \new_[13210]_ , \new_[13213]_ , \new_[13216]_ ,
    \new_[13217]_ , \new_[13218]_ , \new_[13222]_ , \new_[13223]_ ,
    \new_[13226]_ , \new_[13229]_ , \new_[13230]_ , \new_[13231]_ ,
    \new_[13235]_ , \new_[13236]_ , \new_[13239]_ , \new_[13242]_ ,
    \new_[13243]_ , \new_[13244]_ , \new_[13248]_ , \new_[13249]_ ,
    \new_[13252]_ , \new_[13255]_ , \new_[13256]_ , \new_[13257]_ ,
    \new_[13261]_ , \new_[13262]_ , \new_[13265]_ , \new_[13268]_ ,
    \new_[13269]_ , \new_[13270]_ , \new_[13274]_ , \new_[13275]_ ,
    \new_[13278]_ , \new_[13281]_ , \new_[13282]_ , \new_[13283]_ ,
    \new_[13287]_ , \new_[13288]_ , \new_[13291]_ , \new_[13294]_ ,
    \new_[13295]_ , \new_[13296]_ , \new_[13300]_ , \new_[13301]_ ,
    \new_[13304]_ , \new_[13307]_ , \new_[13308]_ , \new_[13309]_ ,
    \new_[13313]_ , \new_[13314]_ , \new_[13317]_ , \new_[13320]_ ,
    \new_[13321]_ , \new_[13322]_ , \new_[13326]_ , \new_[13327]_ ,
    \new_[13330]_ , \new_[13333]_ , \new_[13334]_ , \new_[13335]_ ,
    \new_[13339]_ , \new_[13340]_ , \new_[13343]_ , \new_[13346]_ ,
    \new_[13347]_ , \new_[13348]_ , \new_[13352]_ , \new_[13353]_ ,
    \new_[13356]_ , \new_[13359]_ , \new_[13360]_ , \new_[13361]_ ,
    \new_[13365]_ , \new_[13366]_ , \new_[13369]_ , \new_[13372]_ ,
    \new_[13373]_ , \new_[13374]_ , \new_[13378]_ , \new_[13379]_ ,
    \new_[13382]_ , \new_[13385]_ , \new_[13386]_ , \new_[13387]_ ,
    \new_[13391]_ , \new_[13392]_ , \new_[13395]_ , \new_[13398]_ ,
    \new_[13399]_ , \new_[13400]_ , \new_[13404]_ , \new_[13405]_ ,
    \new_[13408]_ , \new_[13411]_ , \new_[13412]_ , \new_[13413]_ ,
    \new_[13417]_ , \new_[13418]_ , \new_[13421]_ , \new_[13424]_ ,
    \new_[13425]_ , \new_[13426]_ , \new_[13430]_ , \new_[13431]_ ,
    \new_[13434]_ , \new_[13437]_ , \new_[13438]_ , \new_[13439]_ ,
    \new_[13443]_ , \new_[13444]_ , \new_[13447]_ , \new_[13450]_ ,
    \new_[13451]_ , \new_[13452]_ , \new_[13456]_ , \new_[13457]_ ,
    \new_[13460]_ , \new_[13463]_ , \new_[13464]_ , \new_[13465]_ ,
    \new_[13469]_ , \new_[13470]_ , \new_[13473]_ , \new_[13476]_ ,
    \new_[13477]_ , \new_[13478]_ , \new_[13482]_ , \new_[13483]_ ,
    \new_[13486]_ , \new_[13489]_ , \new_[13490]_ , \new_[13491]_ ,
    \new_[13495]_ , \new_[13496]_ , \new_[13499]_ , \new_[13502]_ ,
    \new_[13503]_ , \new_[13504]_ , \new_[13508]_ , \new_[13509]_ ,
    \new_[13512]_ , \new_[13515]_ , \new_[13516]_ , \new_[13517]_ ,
    \new_[13521]_ , \new_[13522]_ , \new_[13525]_ , \new_[13528]_ ,
    \new_[13529]_ , \new_[13530]_ , \new_[13534]_ , \new_[13535]_ ,
    \new_[13538]_ , \new_[13541]_ , \new_[13542]_ , \new_[13543]_ ,
    \new_[13547]_ , \new_[13548]_ , \new_[13551]_ , \new_[13554]_ ,
    \new_[13555]_ , \new_[13556]_ , \new_[13560]_ , \new_[13561]_ ,
    \new_[13564]_ , \new_[13567]_ , \new_[13568]_ , \new_[13569]_ ,
    \new_[13573]_ , \new_[13574]_ , \new_[13577]_ , \new_[13580]_ ,
    \new_[13581]_ , \new_[13582]_ , \new_[13586]_ , \new_[13587]_ ,
    \new_[13590]_ , \new_[13593]_ , \new_[13594]_ , \new_[13595]_ ,
    \new_[13599]_ , \new_[13600]_ , \new_[13603]_ , \new_[13606]_ ,
    \new_[13607]_ , \new_[13608]_ , \new_[13612]_ , \new_[13613]_ ,
    \new_[13616]_ , \new_[13619]_ , \new_[13620]_ , \new_[13621]_ ,
    \new_[13625]_ , \new_[13626]_ , \new_[13629]_ , \new_[13632]_ ,
    \new_[13633]_ , \new_[13634]_ , \new_[13638]_ , \new_[13639]_ ,
    \new_[13642]_ , \new_[13645]_ , \new_[13646]_ , \new_[13647]_ ,
    \new_[13651]_ , \new_[13652]_ , \new_[13655]_ , \new_[13658]_ ,
    \new_[13659]_ , \new_[13660]_ , \new_[13664]_ , \new_[13665]_ ,
    \new_[13668]_ , \new_[13671]_ , \new_[13672]_ , \new_[13673]_ ,
    \new_[13677]_ , \new_[13678]_ , \new_[13681]_ , \new_[13684]_ ,
    \new_[13685]_ , \new_[13686]_ , \new_[13690]_ , \new_[13691]_ ,
    \new_[13694]_ , \new_[13697]_ , \new_[13698]_ , \new_[13699]_ ,
    \new_[13703]_ , \new_[13704]_ , \new_[13707]_ , \new_[13710]_ ,
    \new_[13711]_ , \new_[13712]_ , \new_[13716]_ , \new_[13717]_ ,
    \new_[13720]_ , \new_[13723]_ , \new_[13724]_ , \new_[13725]_ ,
    \new_[13729]_ , \new_[13730]_ , \new_[13733]_ , \new_[13736]_ ,
    \new_[13737]_ , \new_[13738]_ , \new_[13742]_ , \new_[13743]_ ,
    \new_[13746]_ , \new_[13749]_ , \new_[13750]_ , \new_[13751]_ ,
    \new_[13755]_ , \new_[13756]_ , \new_[13759]_ , \new_[13762]_ ,
    \new_[13763]_ , \new_[13764]_ , \new_[13768]_ , \new_[13769]_ ,
    \new_[13772]_ , \new_[13775]_ , \new_[13776]_ , \new_[13777]_ ,
    \new_[13781]_ , \new_[13782]_ , \new_[13785]_ , \new_[13788]_ ,
    \new_[13789]_ , \new_[13790]_ , \new_[13794]_ , \new_[13795]_ ,
    \new_[13798]_ , \new_[13801]_ , \new_[13802]_ , \new_[13803]_ ,
    \new_[13807]_ , \new_[13808]_ , \new_[13811]_ , \new_[13814]_ ,
    \new_[13815]_ , \new_[13816]_ , \new_[13820]_ , \new_[13821]_ ,
    \new_[13824]_ , \new_[13827]_ , \new_[13828]_ , \new_[13829]_ ,
    \new_[13833]_ , \new_[13834]_ , \new_[13837]_ , \new_[13840]_ ,
    \new_[13841]_ , \new_[13842]_ , \new_[13846]_ , \new_[13847]_ ,
    \new_[13850]_ , \new_[13853]_ , \new_[13854]_ , \new_[13855]_ ,
    \new_[13859]_ , \new_[13860]_ , \new_[13863]_ , \new_[13866]_ ,
    \new_[13867]_ , \new_[13868]_ , \new_[13872]_ , \new_[13873]_ ,
    \new_[13876]_ , \new_[13879]_ , \new_[13880]_ , \new_[13881]_ ,
    \new_[13885]_ , \new_[13886]_ , \new_[13889]_ , \new_[13892]_ ,
    \new_[13893]_ , \new_[13894]_ , \new_[13898]_ , \new_[13899]_ ,
    \new_[13902]_ , \new_[13905]_ , \new_[13906]_ , \new_[13907]_ ,
    \new_[13911]_ , \new_[13912]_ , \new_[13915]_ , \new_[13918]_ ,
    \new_[13919]_ , \new_[13920]_ , \new_[13924]_ , \new_[13925]_ ,
    \new_[13928]_ , \new_[13931]_ , \new_[13932]_ , \new_[13933]_ ,
    \new_[13937]_ , \new_[13938]_ , \new_[13941]_ , \new_[13944]_ ,
    \new_[13945]_ , \new_[13946]_ , \new_[13950]_ , \new_[13951]_ ,
    \new_[13954]_ , \new_[13957]_ , \new_[13958]_ , \new_[13959]_ ,
    \new_[13963]_ , \new_[13964]_ , \new_[13967]_ , \new_[13970]_ ,
    \new_[13971]_ , \new_[13972]_ , \new_[13976]_ , \new_[13977]_ ,
    \new_[13980]_ , \new_[13983]_ , \new_[13984]_ , \new_[13985]_ ,
    \new_[13989]_ , \new_[13990]_ , \new_[13993]_ , \new_[13996]_ ,
    \new_[13997]_ , \new_[13998]_ , \new_[14002]_ , \new_[14003]_ ,
    \new_[14006]_ , \new_[14009]_ , \new_[14010]_ , \new_[14011]_ ,
    \new_[14015]_ , \new_[14016]_ , \new_[14019]_ , \new_[14022]_ ,
    \new_[14023]_ , \new_[14024]_ , \new_[14028]_ , \new_[14029]_ ,
    \new_[14032]_ , \new_[14035]_ , \new_[14036]_ , \new_[14037]_ ,
    \new_[14041]_ , \new_[14042]_ , \new_[14045]_ , \new_[14048]_ ,
    \new_[14049]_ , \new_[14050]_ , \new_[14054]_ , \new_[14055]_ ,
    \new_[14058]_ , \new_[14061]_ , \new_[14062]_ , \new_[14063]_ ,
    \new_[14067]_ , \new_[14068]_ , \new_[14071]_ , \new_[14074]_ ,
    \new_[14075]_ , \new_[14076]_ , \new_[14080]_ , \new_[14081]_ ,
    \new_[14084]_ , \new_[14087]_ , \new_[14088]_ , \new_[14089]_ ,
    \new_[14093]_ , \new_[14094]_ , \new_[14097]_ , \new_[14100]_ ,
    \new_[14101]_ , \new_[14102]_ , \new_[14106]_ , \new_[14107]_ ,
    \new_[14110]_ , \new_[14113]_ , \new_[14114]_ , \new_[14115]_ ,
    \new_[14119]_ , \new_[14120]_ , \new_[14123]_ , \new_[14126]_ ,
    \new_[14127]_ , \new_[14128]_ , \new_[14132]_ , \new_[14133]_ ,
    \new_[14136]_ , \new_[14139]_ , \new_[14140]_ , \new_[14141]_ ,
    \new_[14145]_ , \new_[14146]_ , \new_[14149]_ , \new_[14152]_ ,
    \new_[14153]_ , \new_[14154]_ , \new_[14158]_ , \new_[14159]_ ,
    \new_[14162]_ , \new_[14165]_ , \new_[14166]_ , \new_[14167]_ ,
    \new_[14171]_ , \new_[14172]_ , \new_[14175]_ , \new_[14178]_ ,
    \new_[14179]_ , \new_[14180]_ , \new_[14184]_ , \new_[14185]_ ,
    \new_[14188]_ , \new_[14191]_ , \new_[14192]_ , \new_[14193]_ ,
    \new_[14197]_ , \new_[14198]_ , \new_[14201]_ , \new_[14204]_ ,
    \new_[14205]_ , \new_[14206]_ , \new_[14210]_ , \new_[14211]_ ,
    \new_[14214]_ , \new_[14217]_ , \new_[14218]_ , \new_[14219]_ ,
    \new_[14223]_ , \new_[14224]_ , \new_[14227]_ , \new_[14230]_ ,
    \new_[14231]_ , \new_[14232]_ , \new_[14236]_ , \new_[14237]_ ,
    \new_[14240]_ , \new_[14243]_ , \new_[14244]_ , \new_[14245]_ ,
    \new_[14249]_ , \new_[14250]_ , \new_[14253]_ , \new_[14256]_ ,
    \new_[14257]_ , \new_[14258]_ , \new_[14262]_ , \new_[14263]_ ,
    \new_[14266]_ , \new_[14269]_ , \new_[14270]_ , \new_[14271]_ ,
    \new_[14275]_ , \new_[14276]_ , \new_[14279]_ , \new_[14282]_ ,
    \new_[14283]_ , \new_[14284]_ , \new_[14288]_ , \new_[14289]_ ,
    \new_[14292]_ , \new_[14295]_ , \new_[14296]_ , \new_[14297]_ ,
    \new_[14301]_ , \new_[14302]_ , \new_[14305]_ , \new_[14308]_ ,
    \new_[14309]_ , \new_[14310]_ , \new_[14314]_ , \new_[14315]_ ,
    \new_[14318]_ , \new_[14321]_ , \new_[14322]_ , \new_[14323]_ ,
    \new_[14327]_ , \new_[14328]_ , \new_[14331]_ , \new_[14334]_ ,
    \new_[14335]_ , \new_[14336]_ , \new_[14340]_ , \new_[14341]_ ,
    \new_[14344]_ , \new_[14347]_ , \new_[14348]_ , \new_[14349]_ ,
    \new_[14353]_ , \new_[14354]_ , \new_[14357]_ , \new_[14360]_ ,
    \new_[14361]_ , \new_[14362]_ , \new_[14366]_ , \new_[14367]_ ,
    \new_[14370]_ , \new_[14373]_ , \new_[14374]_ , \new_[14375]_ ,
    \new_[14379]_ , \new_[14380]_ , \new_[14383]_ , \new_[14386]_ ,
    \new_[14387]_ , \new_[14388]_ , \new_[14392]_ , \new_[14393]_ ,
    \new_[14396]_ , \new_[14399]_ , \new_[14400]_ , \new_[14401]_ ,
    \new_[14405]_ , \new_[14406]_ , \new_[14409]_ , \new_[14412]_ ,
    \new_[14413]_ , \new_[14414]_ , \new_[14418]_ , \new_[14419]_ ,
    \new_[14422]_ , \new_[14425]_ , \new_[14426]_ , \new_[14427]_ ,
    \new_[14431]_ , \new_[14432]_ , \new_[14435]_ , \new_[14438]_ ,
    \new_[14439]_ , \new_[14440]_ , \new_[14444]_ , \new_[14445]_ ,
    \new_[14448]_ , \new_[14451]_ , \new_[14452]_ , \new_[14453]_ ,
    \new_[14457]_ , \new_[14458]_ , \new_[14461]_ , \new_[14464]_ ,
    \new_[14465]_ , \new_[14466]_ , \new_[14470]_ , \new_[14471]_ ,
    \new_[14474]_ , \new_[14477]_ , \new_[14478]_ , \new_[14479]_ ,
    \new_[14483]_ , \new_[14484]_ , \new_[14487]_ , \new_[14490]_ ,
    \new_[14491]_ , \new_[14492]_ , \new_[14496]_ , \new_[14497]_ ,
    \new_[14500]_ , \new_[14503]_ , \new_[14504]_ , \new_[14505]_ ,
    \new_[14509]_ , \new_[14510]_ , \new_[14513]_ , \new_[14516]_ ,
    \new_[14517]_ , \new_[14518]_ , \new_[14522]_ , \new_[14523]_ ,
    \new_[14526]_ , \new_[14529]_ , \new_[14530]_ , \new_[14531]_ ,
    \new_[14535]_ , \new_[14536]_ , \new_[14539]_ , \new_[14542]_ ,
    \new_[14543]_ , \new_[14544]_ , \new_[14548]_ , \new_[14549]_ ,
    \new_[14552]_ , \new_[14555]_ , \new_[14556]_ , \new_[14557]_ ,
    \new_[14561]_ , \new_[14562]_ , \new_[14565]_ , \new_[14568]_ ,
    \new_[14569]_ , \new_[14570]_ , \new_[14574]_ , \new_[14575]_ ,
    \new_[14578]_ , \new_[14581]_ , \new_[14582]_ , \new_[14583]_ ,
    \new_[14587]_ , \new_[14588]_ , \new_[14591]_ , \new_[14594]_ ,
    \new_[14595]_ , \new_[14596]_ , \new_[14600]_ , \new_[14601]_ ,
    \new_[14604]_ , \new_[14607]_ , \new_[14608]_ , \new_[14609]_ ,
    \new_[14613]_ , \new_[14614]_ , \new_[14617]_ , \new_[14620]_ ,
    \new_[14621]_ , \new_[14622]_ , \new_[14626]_ , \new_[14627]_ ,
    \new_[14630]_ , \new_[14633]_ , \new_[14634]_ , \new_[14635]_ ,
    \new_[14639]_ , \new_[14640]_ , \new_[14643]_ , \new_[14646]_ ,
    \new_[14647]_ , \new_[14648]_ , \new_[14652]_ , \new_[14653]_ ,
    \new_[14656]_ , \new_[14659]_ , \new_[14660]_ , \new_[14661]_ ,
    \new_[14665]_ , \new_[14666]_ , \new_[14669]_ , \new_[14672]_ ,
    \new_[14673]_ , \new_[14674]_ , \new_[14678]_ , \new_[14679]_ ,
    \new_[14682]_ , \new_[14685]_ , \new_[14686]_ , \new_[14687]_ ,
    \new_[14691]_ , \new_[14692]_ , \new_[14695]_ , \new_[14698]_ ,
    \new_[14699]_ , \new_[14700]_ , \new_[14704]_ , \new_[14705]_ ,
    \new_[14708]_ , \new_[14711]_ , \new_[14712]_ , \new_[14713]_ ,
    \new_[14717]_ , \new_[14718]_ , \new_[14721]_ , \new_[14724]_ ,
    \new_[14725]_ , \new_[14726]_ , \new_[14730]_ , \new_[14731]_ ,
    \new_[14734]_ , \new_[14737]_ , \new_[14738]_ , \new_[14739]_ ,
    \new_[14743]_ , \new_[14744]_ , \new_[14747]_ , \new_[14750]_ ,
    \new_[14751]_ , \new_[14752]_ , \new_[14756]_ , \new_[14757]_ ,
    \new_[14760]_ , \new_[14763]_ , \new_[14764]_ , \new_[14765]_ ,
    \new_[14769]_ , \new_[14770]_ , \new_[14773]_ , \new_[14776]_ ,
    \new_[14777]_ , \new_[14778]_ , \new_[14782]_ , \new_[14783]_ ,
    \new_[14786]_ , \new_[14789]_ , \new_[14790]_ , \new_[14791]_ ,
    \new_[14795]_ , \new_[14796]_ , \new_[14799]_ , \new_[14802]_ ,
    \new_[14803]_ , \new_[14804]_ , \new_[14808]_ , \new_[14809]_ ,
    \new_[14812]_ , \new_[14815]_ , \new_[14816]_ , \new_[14817]_ ,
    \new_[14821]_ , \new_[14822]_ , \new_[14825]_ , \new_[14828]_ ,
    \new_[14829]_ , \new_[14830]_ , \new_[14834]_ , \new_[14835]_ ,
    \new_[14838]_ , \new_[14841]_ , \new_[14842]_ , \new_[14843]_ ,
    \new_[14847]_ , \new_[14848]_ , \new_[14851]_ , \new_[14854]_ ,
    \new_[14855]_ , \new_[14856]_ , \new_[14860]_ , \new_[14861]_ ,
    \new_[14864]_ , \new_[14867]_ , \new_[14868]_ , \new_[14869]_ ,
    \new_[14873]_ , \new_[14874]_ , \new_[14877]_ , \new_[14880]_ ,
    \new_[14881]_ , \new_[14882]_ , \new_[14886]_ , \new_[14887]_ ,
    \new_[14890]_ , \new_[14893]_ , \new_[14894]_ , \new_[14895]_ ,
    \new_[14899]_ , \new_[14900]_ , \new_[14903]_ , \new_[14906]_ ,
    \new_[14907]_ , \new_[14908]_ , \new_[14912]_ , \new_[14913]_ ,
    \new_[14916]_ , \new_[14919]_ , \new_[14920]_ , \new_[14921]_ ,
    \new_[14925]_ , \new_[14926]_ , \new_[14929]_ , \new_[14932]_ ,
    \new_[14933]_ , \new_[14934]_ , \new_[14938]_ , \new_[14939]_ ,
    \new_[14942]_ , \new_[14945]_ , \new_[14946]_ , \new_[14947]_ ,
    \new_[14951]_ , \new_[14952]_ , \new_[14955]_ , \new_[14958]_ ,
    \new_[14959]_ , \new_[14960]_ , \new_[14964]_ , \new_[14965]_ ,
    \new_[14968]_ , \new_[14971]_ , \new_[14972]_ , \new_[14973]_ ,
    \new_[14977]_ , \new_[14978]_ , \new_[14981]_ , \new_[14984]_ ,
    \new_[14985]_ , \new_[14986]_ , \new_[14990]_ , \new_[14991]_ ,
    \new_[14994]_ , \new_[14997]_ , \new_[14998]_ , \new_[14999]_ ,
    \new_[15003]_ , \new_[15004]_ , \new_[15007]_ , \new_[15010]_ ,
    \new_[15011]_ , \new_[15012]_ , \new_[15016]_ , \new_[15017]_ ,
    \new_[15020]_ , \new_[15023]_ , \new_[15024]_ , \new_[15025]_ ,
    \new_[15029]_ , \new_[15030]_ , \new_[15033]_ , \new_[15036]_ ,
    \new_[15037]_ , \new_[15038]_ , \new_[15042]_ , \new_[15043]_ ,
    \new_[15046]_ , \new_[15049]_ , \new_[15050]_ , \new_[15051]_ ,
    \new_[15055]_ , \new_[15056]_ , \new_[15059]_ , \new_[15062]_ ,
    \new_[15063]_ , \new_[15064]_ , \new_[15068]_ , \new_[15069]_ ,
    \new_[15072]_ , \new_[15075]_ , \new_[15076]_ , \new_[15077]_ ,
    \new_[15081]_ , \new_[15082]_ , \new_[15085]_ , \new_[15088]_ ,
    \new_[15089]_ , \new_[15090]_ , \new_[15094]_ , \new_[15095]_ ,
    \new_[15098]_ , \new_[15101]_ , \new_[15102]_ , \new_[15103]_ ,
    \new_[15107]_ , \new_[15108]_ , \new_[15111]_ , \new_[15114]_ ,
    \new_[15115]_ , \new_[15116]_ , \new_[15120]_ , \new_[15121]_ ,
    \new_[15124]_ , \new_[15127]_ , \new_[15128]_ , \new_[15129]_ ,
    \new_[15133]_ , \new_[15134]_ , \new_[15137]_ , \new_[15140]_ ,
    \new_[15141]_ , \new_[15142]_ , \new_[15146]_ , \new_[15147]_ ,
    \new_[15150]_ , \new_[15153]_ , \new_[15154]_ , \new_[15155]_ ,
    \new_[15159]_ , \new_[15160]_ , \new_[15163]_ , \new_[15166]_ ,
    \new_[15167]_ , \new_[15168]_ , \new_[15172]_ , \new_[15173]_ ,
    \new_[15176]_ , \new_[15179]_ , \new_[15180]_ , \new_[15181]_ ,
    \new_[15185]_ , \new_[15186]_ , \new_[15189]_ , \new_[15192]_ ,
    \new_[15193]_ , \new_[15194]_ , \new_[15198]_ , \new_[15199]_ ,
    \new_[15202]_ , \new_[15205]_ , \new_[15206]_ , \new_[15207]_ ,
    \new_[15211]_ , \new_[15212]_ , \new_[15215]_ , \new_[15218]_ ,
    \new_[15219]_ , \new_[15220]_ , \new_[15224]_ , \new_[15225]_ ,
    \new_[15228]_ , \new_[15231]_ , \new_[15232]_ , \new_[15233]_ ,
    \new_[15237]_ , \new_[15238]_ , \new_[15241]_ , \new_[15244]_ ,
    \new_[15245]_ , \new_[15246]_ , \new_[15250]_ , \new_[15251]_ ,
    \new_[15254]_ , \new_[15257]_ , \new_[15258]_ , \new_[15259]_ ,
    \new_[15263]_ , \new_[15264]_ , \new_[15267]_ , \new_[15270]_ ,
    \new_[15271]_ , \new_[15272]_ , \new_[15276]_ , \new_[15277]_ ,
    \new_[15280]_ , \new_[15283]_ , \new_[15284]_ , \new_[15285]_ ,
    \new_[15289]_ , \new_[15290]_ , \new_[15293]_ , \new_[15296]_ ,
    \new_[15297]_ , \new_[15298]_ , \new_[15302]_ , \new_[15303]_ ,
    \new_[15306]_ , \new_[15309]_ , \new_[15310]_ , \new_[15311]_ ,
    \new_[15315]_ , \new_[15316]_ , \new_[15319]_ , \new_[15322]_ ,
    \new_[15323]_ , \new_[15324]_ , \new_[15328]_ , \new_[15329]_ ,
    \new_[15332]_ , \new_[15335]_ , \new_[15336]_ , \new_[15337]_ ,
    \new_[15341]_ , \new_[15342]_ , \new_[15345]_ , \new_[15348]_ ,
    \new_[15349]_ , \new_[15350]_ , \new_[15354]_ , \new_[15355]_ ,
    \new_[15358]_ , \new_[15361]_ , \new_[15362]_ , \new_[15363]_ ,
    \new_[15367]_ , \new_[15368]_ , \new_[15371]_ , \new_[15374]_ ,
    \new_[15375]_ , \new_[15376]_ , \new_[15380]_ , \new_[15381]_ ,
    \new_[15384]_ , \new_[15387]_ , \new_[15388]_ , \new_[15389]_ ,
    \new_[15393]_ , \new_[15394]_ , \new_[15397]_ , \new_[15400]_ ,
    \new_[15401]_ , \new_[15402]_ , \new_[15406]_ , \new_[15407]_ ,
    \new_[15410]_ , \new_[15413]_ , \new_[15414]_ , \new_[15415]_ ,
    \new_[15419]_ , \new_[15420]_ , \new_[15423]_ , \new_[15426]_ ,
    \new_[15427]_ , \new_[15428]_ , \new_[15432]_ , \new_[15433]_ ,
    \new_[15436]_ , \new_[15439]_ , \new_[15440]_ , \new_[15441]_ ,
    \new_[15445]_ , \new_[15446]_ , \new_[15449]_ , \new_[15452]_ ,
    \new_[15453]_ , \new_[15454]_ , \new_[15458]_ , \new_[15459]_ ,
    \new_[15462]_ , \new_[15465]_ , \new_[15466]_ , \new_[15467]_ ,
    \new_[15471]_ , \new_[15472]_ , \new_[15475]_ , \new_[15478]_ ,
    \new_[15479]_ , \new_[15480]_ , \new_[15484]_ , \new_[15485]_ ,
    \new_[15488]_ , \new_[15491]_ , \new_[15492]_ , \new_[15493]_ ,
    \new_[15497]_ , \new_[15498]_ , \new_[15501]_ , \new_[15504]_ ,
    \new_[15505]_ , \new_[15506]_ , \new_[15510]_ , \new_[15511]_ ,
    \new_[15514]_ , \new_[15517]_ , \new_[15518]_ , \new_[15519]_ ,
    \new_[15523]_ , \new_[15524]_ , \new_[15527]_ , \new_[15530]_ ,
    \new_[15531]_ , \new_[15532]_ , \new_[15536]_ , \new_[15537]_ ,
    \new_[15540]_ , \new_[15543]_ , \new_[15544]_ , \new_[15545]_ ,
    \new_[15549]_ , \new_[15550]_ , \new_[15553]_ , \new_[15556]_ ,
    \new_[15557]_ , \new_[15558]_ , \new_[15562]_ , \new_[15563]_ ,
    \new_[15566]_ , \new_[15569]_ , \new_[15570]_ , \new_[15571]_ ,
    \new_[15575]_ , \new_[15576]_ , \new_[15579]_ , \new_[15582]_ ,
    \new_[15583]_ , \new_[15584]_ , \new_[15588]_ , \new_[15589]_ ,
    \new_[15592]_ , \new_[15595]_ , \new_[15596]_ , \new_[15597]_ ,
    \new_[15601]_ , \new_[15602]_ , \new_[15605]_ , \new_[15608]_ ,
    \new_[15609]_ , \new_[15610]_ , \new_[15614]_ , \new_[15615]_ ,
    \new_[15618]_ , \new_[15621]_ , \new_[15622]_ , \new_[15623]_ ,
    \new_[15627]_ , \new_[15628]_ , \new_[15631]_ , \new_[15634]_ ,
    \new_[15635]_ , \new_[15636]_ , \new_[15640]_ , \new_[15641]_ ,
    \new_[15644]_ , \new_[15647]_ , \new_[15648]_ , \new_[15649]_ ,
    \new_[15653]_ , \new_[15654]_ , \new_[15657]_ , \new_[15660]_ ,
    \new_[15661]_ , \new_[15662]_ , \new_[15666]_ , \new_[15667]_ ,
    \new_[15670]_ , \new_[15673]_ , \new_[15674]_ , \new_[15675]_ ,
    \new_[15679]_ , \new_[15680]_ , \new_[15683]_ , \new_[15686]_ ,
    \new_[15687]_ , \new_[15688]_ , \new_[15692]_ , \new_[15693]_ ,
    \new_[15696]_ , \new_[15699]_ , \new_[15700]_ , \new_[15701]_ ,
    \new_[15705]_ , \new_[15706]_ , \new_[15709]_ , \new_[15712]_ ,
    \new_[15713]_ , \new_[15714]_ , \new_[15718]_ , \new_[15719]_ ,
    \new_[15722]_ , \new_[15725]_ , \new_[15726]_ , \new_[15727]_ ,
    \new_[15731]_ , \new_[15732]_ , \new_[15735]_ , \new_[15738]_ ,
    \new_[15739]_ , \new_[15740]_ , \new_[15744]_ , \new_[15745]_ ,
    \new_[15748]_ , \new_[15751]_ , \new_[15752]_ , \new_[15753]_ ,
    \new_[15757]_ , \new_[15758]_ , \new_[15761]_ , \new_[15764]_ ,
    \new_[15765]_ , \new_[15766]_ , \new_[15770]_ , \new_[15771]_ ,
    \new_[15774]_ , \new_[15777]_ , \new_[15778]_ , \new_[15779]_ ,
    \new_[15783]_ , \new_[15784]_ , \new_[15787]_ , \new_[15790]_ ,
    \new_[15791]_ , \new_[15792]_ , \new_[15796]_ , \new_[15797]_ ,
    \new_[15800]_ , \new_[15803]_ , \new_[15804]_ , \new_[15805]_ ,
    \new_[15809]_ , \new_[15810]_ , \new_[15813]_ , \new_[15816]_ ,
    \new_[15817]_ , \new_[15818]_ , \new_[15822]_ , \new_[15823]_ ,
    \new_[15826]_ , \new_[15829]_ , \new_[15830]_ , \new_[15831]_ ,
    \new_[15835]_ , \new_[15836]_ , \new_[15839]_ , \new_[15842]_ ,
    \new_[15843]_ , \new_[15844]_ , \new_[15848]_ , \new_[15849]_ ,
    \new_[15852]_ , \new_[15855]_ , \new_[15856]_ , \new_[15857]_ ,
    \new_[15861]_ , \new_[15862]_ , \new_[15865]_ , \new_[15868]_ ,
    \new_[15869]_ , \new_[15870]_ , \new_[15874]_ , \new_[15875]_ ,
    \new_[15878]_ , \new_[15881]_ , \new_[15882]_ , \new_[15883]_ ,
    \new_[15887]_ , \new_[15888]_ , \new_[15891]_ , \new_[15894]_ ,
    \new_[15895]_ , \new_[15896]_ , \new_[15900]_ , \new_[15901]_ ,
    \new_[15904]_ , \new_[15907]_ , \new_[15908]_ , \new_[15909]_ ,
    \new_[15913]_ , \new_[15914]_ , \new_[15917]_ , \new_[15920]_ ,
    \new_[15921]_ , \new_[15922]_ , \new_[15926]_ , \new_[15927]_ ,
    \new_[15930]_ , \new_[15933]_ , \new_[15934]_ , \new_[15935]_ ,
    \new_[15939]_ , \new_[15940]_ , \new_[15943]_ , \new_[15946]_ ,
    \new_[15947]_ , \new_[15948]_ , \new_[15952]_ , \new_[15953]_ ,
    \new_[15956]_ , \new_[15959]_ , \new_[15960]_ , \new_[15961]_ ,
    \new_[15965]_ , \new_[15966]_ , \new_[15969]_ , \new_[15972]_ ,
    \new_[15973]_ , \new_[15974]_ , \new_[15978]_ , \new_[15979]_ ,
    \new_[15982]_ , \new_[15985]_ , \new_[15986]_ , \new_[15987]_ ,
    \new_[15991]_ , \new_[15992]_ , \new_[15995]_ , \new_[15998]_ ,
    \new_[15999]_ , \new_[16000]_ , \new_[16004]_ , \new_[16005]_ ,
    \new_[16008]_ , \new_[16011]_ , \new_[16012]_ , \new_[16013]_ ,
    \new_[16017]_ , \new_[16018]_ , \new_[16021]_ , \new_[16024]_ ,
    \new_[16025]_ , \new_[16026]_ , \new_[16030]_ , \new_[16031]_ ,
    \new_[16034]_ , \new_[16037]_ , \new_[16038]_ , \new_[16039]_ ,
    \new_[16043]_ , \new_[16044]_ , \new_[16047]_ , \new_[16050]_ ,
    \new_[16051]_ , \new_[16052]_ , \new_[16056]_ , \new_[16057]_ ,
    \new_[16060]_ , \new_[16063]_ , \new_[16064]_ , \new_[16065]_ ,
    \new_[16069]_ , \new_[16070]_ , \new_[16073]_ , \new_[16076]_ ,
    \new_[16077]_ , \new_[16078]_ , \new_[16082]_ , \new_[16083]_ ,
    \new_[16086]_ , \new_[16089]_ , \new_[16090]_ , \new_[16091]_ ,
    \new_[16095]_ , \new_[16096]_ , \new_[16099]_ , \new_[16102]_ ,
    \new_[16103]_ , \new_[16104]_ , \new_[16108]_ , \new_[16109]_ ,
    \new_[16112]_ , \new_[16115]_ , \new_[16116]_ , \new_[16117]_ ,
    \new_[16121]_ , \new_[16122]_ , \new_[16125]_ , \new_[16128]_ ,
    \new_[16129]_ , \new_[16130]_ , \new_[16134]_ , \new_[16135]_ ,
    \new_[16138]_ , \new_[16141]_ , \new_[16142]_ , \new_[16143]_ ,
    \new_[16147]_ , \new_[16148]_ , \new_[16151]_ , \new_[16154]_ ,
    \new_[16155]_ , \new_[16156]_ , \new_[16160]_ , \new_[16161]_ ,
    \new_[16164]_ , \new_[16167]_ , \new_[16168]_ , \new_[16169]_ ,
    \new_[16173]_ , \new_[16174]_ , \new_[16177]_ , \new_[16180]_ ,
    \new_[16181]_ , \new_[16182]_ , \new_[16186]_ , \new_[16187]_ ,
    \new_[16190]_ , \new_[16193]_ , \new_[16194]_ , \new_[16195]_ ,
    \new_[16199]_ , \new_[16200]_ , \new_[16203]_ , \new_[16206]_ ,
    \new_[16207]_ , \new_[16208]_ , \new_[16212]_ , \new_[16213]_ ,
    \new_[16216]_ , \new_[16219]_ , \new_[16220]_ , \new_[16221]_ ,
    \new_[16225]_ , \new_[16226]_ , \new_[16229]_ , \new_[16232]_ ,
    \new_[16233]_ , \new_[16234]_ , \new_[16238]_ , \new_[16239]_ ,
    \new_[16242]_ , \new_[16245]_ , \new_[16246]_ , \new_[16247]_ ,
    \new_[16251]_ , \new_[16252]_ , \new_[16255]_ , \new_[16258]_ ,
    \new_[16259]_ , \new_[16260]_ , \new_[16264]_ , \new_[16265]_ ,
    \new_[16268]_ , \new_[16271]_ , \new_[16272]_ , \new_[16273]_ ,
    \new_[16277]_ , \new_[16278]_ , \new_[16281]_ , \new_[16284]_ ,
    \new_[16285]_ , \new_[16286]_ , \new_[16290]_ , \new_[16291]_ ,
    \new_[16294]_ , \new_[16297]_ , \new_[16298]_ , \new_[16299]_ ,
    \new_[16303]_ , \new_[16304]_ , \new_[16307]_ , \new_[16310]_ ,
    \new_[16311]_ , \new_[16312]_ , \new_[16316]_ , \new_[16317]_ ,
    \new_[16320]_ , \new_[16323]_ , \new_[16324]_ , \new_[16325]_ ,
    \new_[16329]_ , \new_[16330]_ , \new_[16333]_ , \new_[16336]_ ,
    \new_[16337]_ , \new_[16338]_ , \new_[16342]_ , \new_[16343]_ ,
    \new_[16346]_ , \new_[16349]_ , \new_[16350]_ , \new_[16351]_ ,
    \new_[16355]_ , \new_[16356]_ , \new_[16359]_ , \new_[16362]_ ,
    \new_[16363]_ , \new_[16364]_ , \new_[16368]_ , \new_[16369]_ ,
    \new_[16372]_ , \new_[16375]_ , \new_[16376]_ , \new_[16377]_ ,
    \new_[16381]_ , \new_[16382]_ , \new_[16385]_ , \new_[16388]_ ,
    \new_[16389]_ , \new_[16390]_ , \new_[16394]_ , \new_[16395]_ ,
    \new_[16398]_ , \new_[16401]_ , \new_[16402]_ , \new_[16403]_ ,
    \new_[16407]_ , \new_[16408]_ , \new_[16411]_ , \new_[16414]_ ,
    \new_[16415]_ , \new_[16416]_ , \new_[16420]_ , \new_[16421]_ ,
    \new_[16424]_ , \new_[16427]_ , \new_[16428]_ , \new_[16429]_ ,
    \new_[16433]_ , \new_[16434]_ , \new_[16437]_ , \new_[16440]_ ,
    \new_[16441]_ , \new_[16442]_ , \new_[16446]_ , \new_[16447]_ ,
    \new_[16450]_ , \new_[16453]_ , \new_[16454]_ , \new_[16455]_ ,
    \new_[16459]_ , \new_[16460]_ , \new_[16463]_ , \new_[16466]_ ,
    \new_[16467]_ , \new_[16468]_ , \new_[16472]_ , \new_[16473]_ ,
    \new_[16476]_ , \new_[16479]_ , \new_[16480]_ , \new_[16481]_ ,
    \new_[16485]_ , \new_[16486]_ , \new_[16489]_ , \new_[16492]_ ,
    \new_[16493]_ , \new_[16494]_ , \new_[16498]_ , \new_[16499]_ ,
    \new_[16502]_ , \new_[16505]_ , \new_[16506]_ , \new_[16507]_ ,
    \new_[16511]_ , \new_[16512]_ , \new_[16515]_ , \new_[16518]_ ,
    \new_[16519]_ , \new_[16520]_ , \new_[16524]_ , \new_[16525]_ ,
    \new_[16528]_ , \new_[16531]_ , \new_[16532]_ , \new_[16533]_ ,
    \new_[16537]_ , \new_[16538]_ , \new_[16541]_ , \new_[16544]_ ,
    \new_[16545]_ , \new_[16546]_ , \new_[16550]_ , \new_[16551]_ ,
    \new_[16554]_ , \new_[16557]_ , \new_[16558]_ , \new_[16559]_ ,
    \new_[16563]_ , \new_[16564]_ , \new_[16567]_ , \new_[16570]_ ,
    \new_[16571]_ , \new_[16572]_ , \new_[16576]_ , \new_[16577]_ ,
    \new_[16580]_ , \new_[16583]_ , \new_[16584]_ , \new_[16585]_ ,
    \new_[16589]_ , \new_[16590]_ , \new_[16593]_ , \new_[16596]_ ,
    \new_[16597]_ , \new_[16598]_ , \new_[16602]_ , \new_[16603]_ ,
    \new_[16606]_ , \new_[16609]_ , \new_[16610]_ , \new_[16611]_ ,
    \new_[16615]_ , \new_[16616]_ , \new_[16619]_ , \new_[16622]_ ,
    \new_[16623]_ , \new_[16624]_ , \new_[16628]_ , \new_[16629]_ ,
    \new_[16632]_ , \new_[16635]_ , \new_[16636]_ , \new_[16637]_ ,
    \new_[16641]_ , \new_[16642]_ , \new_[16645]_ , \new_[16648]_ ,
    \new_[16649]_ , \new_[16650]_ , \new_[16654]_ , \new_[16655]_ ,
    \new_[16658]_ , \new_[16661]_ , \new_[16662]_ , \new_[16663]_ ,
    \new_[16667]_ , \new_[16668]_ , \new_[16671]_ , \new_[16674]_ ,
    \new_[16675]_ , \new_[16676]_ , \new_[16680]_ , \new_[16681]_ ,
    \new_[16684]_ , \new_[16687]_ , \new_[16688]_ , \new_[16689]_ ,
    \new_[16693]_ , \new_[16694]_ , \new_[16697]_ , \new_[16700]_ ,
    \new_[16701]_ , \new_[16702]_ , \new_[16706]_ , \new_[16707]_ ,
    \new_[16710]_ , \new_[16713]_ , \new_[16714]_ , \new_[16715]_ ,
    \new_[16719]_ , \new_[16720]_ , \new_[16723]_ , \new_[16726]_ ,
    \new_[16727]_ , \new_[16728]_ , \new_[16732]_ , \new_[16733]_ ,
    \new_[16736]_ , \new_[16739]_ , \new_[16740]_ , \new_[16741]_ ,
    \new_[16745]_ , \new_[16746]_ , \new_[16749]_ , \new_[16752]_ ,
    \new_[16753]_ , \new_[16754]_ , \new_[16758]_ , \new_[16759]_ ,
    \new_[16762]_ , \new_[16765]_ , \new_[16766]_ , \new_[16767]_ ,
    \new_[16771]_ , \new_[16772]_ , \new_[16775]_ , \new_[16778]_ ,
    \new_[16779]_ , \new_[16780]_ , \new_[16784]_ , \new_[16785]_ ,
    \new_[16788]_ , \new_[16791]_ , \new_[16792]_ , \new_[16793]_ ,
    \new_[16797]_ , \new_[16798]_ , \new_[16801]_ , \new_[16804]_ ,
    \new_[16805]_ , \new_[16806]_ , \new_[16810]_ , \new_[16811]_ ,
    \new_[16814]_ , \new_[16817]_ , \new_[16818]_ , \new_[16819]_ ,
    \new_[16823]_ , \new_[16824]_ , \new_[16827]_ , \new_[16830]_ ,
    \new_[16831]_ , \new_[16832]_ , \new_[16836]_ , \new_[16837]_ ,
    \new_[16840]_ , \new_[16843]_ , \new_[16844]_ , \new_[16845]_ ,
    \new_[16849]_ , \new_[16850]_ , \new_[16853]_ , \new_[16856]_ ,
    \new_[16857]_ , \new_[16858]_ , \new_[16862]_ , \new_[16863]_ ,
    \new_[16866]_ , \new_[16869]_ , \new_[16870]_ , \new_[16871]_ ,
    \new_[16875]_ , \new_[16876]_ , \new_[16879]_ , \new_[16882]_ ,
    \new_[16883]_ , \new_[16884]_ , \new_[16888]_ , \new_[16889]_ ,
    \new_[16892]_ , \new_[16895]_ , \new_[16896]_ , \new_[16897]_ ,
    \new_[16901]_ , \new_[16902]_ , \new_[16905]_ , \new_[16908]_ ,
    \new_[16909]_ , \new_[16910]_ , \new_[16914]_ , \new_[16915]_ ,
    \new_[16918]_ , \new_[16921]_ , \new_[16922]_ , \new_[16923]_ ,
    \new_[16927]_ , \new_[16928]_ , \new_[16931]_ , \new_[16934]_ ,
    \new_[16935]_ , \new_[16936]_ , \new_[16940]_ , \new_[16941]_ ,
    \new_[16944]_ , \new_[16947]_ , \new_[16948]_ , \new_[16949]_ ,
    \new_[16953]_ , \new_[16954]_ , \new_[16957]_ , \new_[16960]_ ,
    \new_[16961]_ , \new_[16962]_ , \new_[16966]_ , \new_[16967]_ ,
    \new_[16970]_ , \new_[16973]_ , \new_[16974]_ , \new_[16975]_ ,
    \new_[16979]_ , \new_[16980]_ , \new_[16983]_ , \new_[16986]_ ,
    \new_[16987]_ , \new_[16988]_ , \new_[16992]_ , \new_[16993]_ ,
    \new_[16996]_ , \new_[16999]_ , \new_[17000]_ , \new_[17001]_ ,
    \new_[17005]_ , \new_[17006]_ , \new_[17009]_ , \new_[17012]_ ,
    \new_[17013]_ , \new_[17014]_ , \new_[17018]_ , \new_[17019]_ ,
    \new_[17022]_ , \new_[17025]_ , \new_[17026]_ , \new_[17027]_ ,
    \new_[17031]_ , \new_[17032]_ , \new_[17035]_ , \new_[17038]_ ,
    \new_[17039]_ , \new_[17040]_ , \new_[17044]_ , \new_[17045]_ ,
    \new_[17048]_ , \new_[17051]_ , \new_[17052]_ , \new_[17053]_ ,
    \new_[17057]_ , \new_[17058]_ , \new_[17061]_ , \new_[17064]_ ,
    \new_[17065]_ , \new_[17066]_ , \new_[17070]_ , \new_[17071]_ ,
    \new_[17074]_ , \new_[17077]_ , \new_[17078]_ , \new_[17079]_ ,
    \new_[17083]_ , \new_[17084]_ , \new_[17087]_ , \new_[17090]_ ,
    \new_[17091]_ , \new_[17092]_ , \new_[17096]_ , \new_[17097]_ ,
    \new_[17100]_ , \new_[17103]_ , \new_[17104]_ , \new_[17105]_ ,
    \new_[17109]_ , \new_[17110]_ , \new_[17113]_ , \new_[17116]_ ,
    \new_[17117]_ , \new_[17118]_ , \new_[17122]_ , \new_[17123]_ ,
    \new_[17126]_ , \new_[17129]_ , \new_[17130]_ , \new_[17131]_ ,
    \new_[17135]_ , \new_[17136]_ , \new_[17139]_ , \new_[17142]_ ,
    \new_[17143]_ , \new_[17144]_ , \new_[17148]_ , \new_[17149]_ ,
    \new_[17152]_ , \new_[17155]_ , \new_[17156]_ , \new_[17157]_ ,
    \new_[17161]_ , \new_[17162]_ , \new_[17165]_ , \new_[17168]_ ,
    \new_[17169]_ , \new_[17170]_ , \new_[17174]_ , \new_[17175]_ ,
    \new_[17178]_ , \new_[17181]_ , \new_[17182]_ , \new_[17183]_ ,
    \new_[17187]_ , \new_[17188]_ , \new_[17191]_ , \new_[17194]_ ,
    \new_[17195]_ , \new_[17196]_ , \new_[17200]_ , \new_[17201]_ ,
    \new_[17204]_ , \new_[17207]_ , \new_[17208]_ , \new_[17209]_ ,
    \new_[17213]_ , \new_[17214]_ , \new_[17217]_ , \new_[17220]_ ,
    \new_[17221]_ , \new_[17222]_ , \new_[17226]_ , \new_[17227]_ ,
    \new_[17230]_ , \new_[17233]_ , \new_[17234]_ , \new_[17235]_ ,
    \new_[17239]_ , \new_[17240]_ , \new_[17243]_ , \new_[17246]_ ,
    \new_[17247]_ , \new_[17248]_ , \new_[17252]_ , \new_[17253]_ ,
    \new_[17256]_ , \new_[17259]_ , \new_[17260]_ , \new_[17261]_ ,
    \new_[17265]_ , \new_[17266]_ , \new_[17269]_ , \new_[17272]_ ,
    \new_[17273]_ , \new_[17274]_ , \new_[17278]_ , \new_[17279]_ ,
    \new_[17282]_ , \new_[17285]_ , \new_[17286]_ , \new_[17287]_ ,
    \new_[17291]_ , \new_[17292]_ , \new_[17295]_ , \new_[17298]_ ,
    \new_[17299]_ , \new_[17300]_ , \new_[17304]_ , \new_[17305]_ ,
    \new_[17308]_ , \new_[17311]_ , \new_[17312]_ , \new_[17313]_ ,
    \new_[17317]_ , \new_[17318]_ , \new_[17321]_ , \new_[17324]_ ,
    \new_[17325]_ , \new_[17326]_ , \new_[17330]_ , \new_[17331]_ ,
    \new_[17334]_ , \new_[17337]_ , \new_[17338]_ , \new_[17339]_ ,
    \new_[17343]_ , \new_[17344]_ , \new_[17347]_ , \new_[17350]_ ,
    \new_[17351]_ , \new_[17352]_ , \new_[17356]_ , \new_[17357]_ ,
    \new_[17360]_ , \new_[17363]_ , \new_[17364]_ , \new_[17365]_ ,
    \new_[17369]_ , \new_[17370]_ , \new_[17373]_ , \new_[17376]_ ,
    \new_[17377]_ , \new_[17378]_ , \new_[17382]_ , \new_[17383]_ ,
    \new_[17386]_ , \new_[17389]_ , \new_[17390]_ , \new_[17391]_ ,
    \new_[17395]_ , \new_[17396]_ , \new_[17399]_ , \new_[17402]_ ,
    \new_[17403]_ , \new_[17404]_ , \new_[17408]_ , \new_[17409]_ ,
    \new_[17412]_ , \new_[17415]_ , \new_[17416]_ , \new_[17417]_ ,
    \new_[17421]_ , \new_[17422]_ , \new_[17425]_ , \new_[17428]_ ,
    \new_[17429]_ , \new_[17430]_ , \new_[17434]_ , \new_[17435]_ ,
    \new_[17438]_ , \new_[17441]_ , \new_[17442]_ , \new_[17443]_ ,
    \new_[17447]_ , \new_[17448]_ , \new_[17451]_ , \new_[17454]_ ,
    \new_[17455]_ , \new_[17456]_ , \new_[17460]_ , \new_[17461]_ ,
    \new_[17464]_ , \new_[17467]_ , \new_[17468]_ , \new_[17469]_ ,
    \new_[17473]_ , \new_[17474]_ , \new_[17477]_ , \new_[17480]_ ,
    \new_[17481]_ , \new_[17482]_ , \new_[17486]_ , \new_[17487]_ ,
    \new_[17490]_ , \new_[17493]_ , \new_[17494]_ , \new_[17495]_ ,
    \new_[17499]_ , \new_[17500]_ , \new_[17503]_ , \new_[17506]_ ,
    \new_[17507]_ , \new_[17508]_ , \new_[17512]_ , \new_[17513]_ ,
    \new_[17516]_ , \new_[17519]_ , \new_[17520]_ , \new_[17521]_ ,
    \new_[17525]_ , \new_[17526]_ , \new_[17529]_ , \new_[17532]_ ,
    \new_[17533]_ , \new_[17534]_ , \new_[17538]_ , \new_[17539]_ ,
    \new_[17542]_ , \new_[17545]_ , \new_[17546]_ , \new_[17547]_ ,
    \new_[17551]_ , \new_[17552]_ , \new_[17555]_ , \new_[17558]_ ,
    \new_[17559]_ , \new_[17560]_ , \new_[17564]_ , \new_[17565]_ ,
    \new_[17568]_ , \new_[17571]_ , \new_[17572]_ , \new_[17573]_ ,
    \new_[17577]_ , \new_[17578]_ , \new_[17581]_ , \new_[17584]_ ,
    \new_[17585]_ , \new_[17586]_ , \new_[17590]_ , \new_[17591]_ ,
    \new_[17594]_ , \new_[17597]_ , \new_[17598]_ , \new_[17599]_ ,
    \new_[17603]_ , \new_[17604]_ , \new_[17607]_ , \new_[17610]_ ,
    \new_[17611]_ , \new_[17612]_ , \new_[17616]_ , \new_[17617]_ ,
    \new_[17620]_ , \new_[17623]_ , \new_[17624]_ , \new_[17625]_ ,
    \new_[17629]_ , \new_[17630]_ , \new_[17633]_ , \new_[17636]_ ,
    \new_[17637]_ , \new_[17638]_ , \new_[17642]_ , \new_[17643]_ ,
    \new_[17646]_ , \new_[17649]_ , \new_[17650]_ , \new_[17651]_ ,
    \new_[17655]_ , \new_[17656]_ , \new_[17659]_ , \new_[17662]_ ,
    \new_[17663]_ , \new_[17664]_ , \new_[17668]_ , \new_[17669]_ ,
    \new_[17672]_ , \new_[17675]_ , \new_[17676]_ , \new_[17677]_ ,
    \new_[17681]_ , \new_[17682]_ , \new_[17685]_ , \new_[17688]_ ,
    \new_[17689]_ , \new_[17690]_ , \new_[17694]_ , \new_[17695]_ ,
    \new_[17698]_ , \new_[17701]_ , \new_[17702]_ , \new_[17703]_ ,
    \new_[17707]_ , \new_[17708]_ , \new_[17711]_ , \new_[17714]_ ,
    \new_[17715]_ , \new_[17716]_ , \new_[17720]_ , \new_[17721]_ ,
    \new_[17724]_ , \new_[17727]_ , \new_[17728]_ , \new_[17729]_ ,
    \new_[17733]_ , \new_[17734]_ , \new_[17737]_ , \new_[17740]_ ,
    \new_[17741]_ , \new_[17742]_ , \new_[17746]_ , \new_[17747]_ ,
    \new_[17750]_ , \new_[17753]_ , \new_[17754]_ , \new_[17755]_ ,
    \new_[17759]_ , \new_[17760]_ , \new_[17763]_ , \new_[17766]_ ,
    \new_[17767]_ , \new_[17768]_ , \new_[17772]_ , \new_[17773]_ ,
    \new_[17776]_ , \new_[17779]_ , \new_[17780]_ , \new_[17781]_ ,
    \new_[17785]_ , \new_[17786]_ , \new_[17789]_ , \new_[17792]_ ,
    \new_[17793]_ , \new_[17794]_ , \new_[17798]_ , \new_[17799]_ ,
    \new_[17802]_ , \new_[17805]_ , \new_[17806]_ , \new_[17807]_ ,
    \new_[17811]_ , \new_[17812]_ , \new_[17815]_ , \new_[17818]_ ,
    \new_[17819]_ , \new_[17820]_ , \new_[17824]_ , \new_[17825]_ ,
    \new_[17828]_ , \new_[17831]_ , \new_[17832]_ , \new_[17833]_ ,
    \new_[17837]_ , \new_[17838]_ , \new_[17841]_ , \new_[17844]_ ,
    \new_[17845]_ , \new_[17846]_ , \new_[17850]_ , \new_[17851]_ ,
    \new_[17854]_ , \new_[17857]_ , \new_[17858]_ , \new_[17859]_ ,
    \new_[17863]_ , \new_[17864]_ , \new_[17867]_ , \new_[17870]_ ,
    \new_[17871]_ , \new_[17872]_ , \new_[17876]_ , \new_[17877]_ ,
    \new_[17880]_ , \new_[17883]_ , \new_[17884]_ , \new_[17885]_ ,
    \new_[17889]_ , \new_[17890]_ , \new_[17893]_ , \new_[17896]_ ,
    \new_[17897]_ , \new_[17898]_ , \new_[17902]_ , \new_[17903]_ ,
    \new_[17906]_ , \new_[17909]_ , \new_[17910]_ , \new_[17911]_ ,
    \new_[17915]_ , \new_[17916]_ , \new_[17919]_ , \new_[17922]_ ,
    \new_[17923]_ , \new_[17924]_ , \new_[17928]_ , \new_[17929]_ ,
    \new_[17932]_ , \new_[17935]_ , \new_[17936]_ , \new_[17937]_ ,
    \new_[17941]_ , \new_[17942]_ , \new_[17945]_ , \new_[17948]_ ,
    \new_[17949]_ , \new_[17950]_ , \new_[17954]_ , \new_[17955]_ ,
    \new_[17958]_ , \new_[17961]_ , \new_[17962]_ , \new_[17963]_ ,
    \new_[17967]_ , \new_[17968]_ , \new_[17971]_ , \new_[17974]_ ,
    \new_[17975]_ , \new_[17976]_ , \new_[17980]_ , \new_[17981]_ ,
    \new_[17984]_ , \new_[17987]_ , \new_[17988]_ , \new_[17989]_ ,
    \new_[17993]_ , \new_[17994]_ , \new_[17997]_ , \new_[18000]_ ,
    \new_[18001]_ , \new_[18002]_ , \new_[18006]_ , \new_[18007]_ ,
    \new_[18010]_ , \new_[18013]_ , \new_[18014]_ , \new_[18015]_ ,
    \new_[18019]_ , \new_[18020]_ , \new_[18023]_ , \new_[18026]_ ,
    \new_[18027]_ , \new_[18028]_ , \new_[18032]_ , \new_[18033]_ ,
    \new_[18036]_ , \new_[18039]_ , \new_[18040]_ , \new_[18041]_ ,
    \new_[18045]_ , \new_[18046]_ , \new_[18049]_ , \new_[18052]_ ,
    \new_[18053]_ , \new_[18054]_ , \new_[18058]_ , \new_[18059]_ ,
    \new_[18062]_ , \new_[18065]_ , \new_[18066]_ , \new_[18067]_ ,
    \new_[18071]_ , \new_[18072]_ , \new_[18075]_ , \new_[18078]_ ,
    \new_[18079]_ , \new_[18080]_ , \new_[18084]_ , \new_[18085]_ ,
    \new_[18088]_ , \new_[18091]_ , \new_[18092]_ , \new_[18093]_ ,
    \new_[18097]_ , \new_[18098]_ , \new_[18101]_ , \new_[18104]_ ,
    \new_[18105]_ , \new_[18106]_ , \new_[18110]_ , \new_[18111]_ ,
    \new_[18114]_ , \new_[18117]_ , \new_[18118]_ , \new_[18119]_ ,
    \new_[18123]_ , \new_[18124]_ , \new_[18127]_ , \new_[18130]_ ,
    \new_[18131]_ , \new_[18132]_ , \new_[18136]_ , \new_[18137]_ ,
    \new_[18140]_ , \new_[18143]_ , \new_[18144]_ , \new_[18145]_ ,
    \new_[18149]_ , \new_[18150]_ , \new_[18153]_ , \new_[18156]_ ,
    \new_[18157]_ , \new_[18158]_ , \new_[18162]_ , \new_[18163]_ ,
    \new_[18166]_ , \new_[18169]_ , \new_[18170]_ , \new_[18171]_ ,
    \new_[18175]_ , \new_[18176]_ , \new_[18179]_ , \new_[18182]_ ,
    \new_[18183]_ , \new_[18184]_ , \new_[18188]_ , \new_[18189]_ ,
    \new_[18192]_ , \new_[18195]_ , \new_[18196]_ , \new_[18197]_ ,
    \new_[18201]_ , \new_[18202]_ , \new_[18205]_ , \new_[18208]_ ,
    \new_[18209]_ , \new_[18210]_ , \new_[18214]_ , \new_[18215]_ ,
    \new_[18218]_ , \new_[18221]_ , \new_[18222]_ , \new_[18223]_ ,
    \new_[18227]_ , \new_[18228]_ , \new_[18231]_ , \new_[18234]_ ,
    \new_[18235]_ , \new_[18236]_ , \new_[18240]_ , \new_[18241]_ ,
    \new_[18244]_ , \new_[18247]_ , \new_[18248]_ , \new_[18249]_ ,
    \new_[18253]_ , \new_[18254]_ , \new_[18257]_ , \new_[18260]_ ,
    \new_[18261]_ , \new_[18262]_ , \new_[18266]_ , \new_[18267]_ ,
    \new_[18270]_ , \new_[18273]_ , \new_[18274]_ , \new_[18275]_ ,
    \new_[18279]_ , \new_[18280]_ , \new_[18283]_ , \new_[18286]_ ,
    \new_[18287]_ , \new_[18288]_ , \new_[18292]_ , \new_[18293]_ ,
    \new_[18296]_ , \new_[18299]_ , \new_[18300]_ , \new_[18301]_ ,
    \new_[18305]_ , \new_[18306]_ , \new_[18309]_ , \new_[18312]_ ,
    \new_[18313]_ , \new_[18314]_ , \new_[18318]_ , \new_[18319]_ ,
    \new_[18322]_ , \new_[18325]_ , \new_[18326]_ , \new_[18327]_ ,
    \new_[18331]_ , \new_[18332]_ , \new_[18335]_ , \new_[18338]_ ,
    \new_[18339]_ , \new_[18340]_ , \new_[18344]_ , \new_[18345]_ ,
    \new_[18348]_ , \new_[18351]_ , \new_[18352]_ , \new_[18353]_ ,
    \new_[18357]_ , \new_[18358]_ , \new_[18361]_ , \new_[18364]_ ,
    \new_[18365]_ , \new_[18366]_ , \new_[18370]_ , \new_[18371]_ ,
    \new_[18374]_ , \new_[18377]_ , \new_[18378]_ , \new_[18379]_ ,
    \new_[18383]_ , \new_[18384]_ , \new_[18387]_ , \new_[18390]_ ,
    \new_[18391]_ , \new_[18392]_ , \new_[18396]_ , \new_[18397]_ ,
    \new_[18400]_ , \new_[18403]_ , \new_[18404]_ , \new_[18405]_ ,
    \new_[18409]_ , \new_[18410]_ , \new_[18413]_ , \new_[18416]_ ,
    \new_[18417]_ , \new_[18418]_ , \new_[18422]_ , \new_[18423]_ ,
    \new_[18426]_ , \new_[18429]_ , \new_[18430]_ , \new_[18431]_ ,
    \new_[18435]_ , \new_[18436]_ , \new_[18439]_ , \new_[18442]_ ,
    \new_[18443]_ , \new_[18444]_ , \new_[18448]_ , \new_[18449]_ ,
    \new_[18452]_ , \new_[18455]_ , \new_[18456]_ , \new_[18457]_ ,
    \new_[18461]_ , \new_[18462]_ , \new_[18465]_ , \new_[18468]_ ,
    \new_[18469]_ , \new_[18470]_ , \new_[18474]_ , \new_[18475]_ ,
    \new_[18478]_ , \new_[18481]_ , \new_[18482]_ , \new_[18483]_ ,
    \new_[18487]_ , \new_[18488]_ , \new_[18491]_ , \new_[18494]_ ,
    \new_[18495]_ , \new_[18496]_ , \new_[18500]_ , \new_[18501]_ ,
    \new_[18504]_ , \new_[18507]_ , \new_[18508]_ , \new_[18509]_ ,
    \new_[18513]_ , \new_[18514]_ , \new_[18517]_ , \new_[18520]_ ,
    \new_[18521]_ , \new_[18522]_ , \new_[18526]_ , \new_[18527]_ ,
    \new_[18530]_ , \new_[18533]_ , \new_[18534]_ , \new_[18535]_ ,
    \new_[18539]_ , \new_[18540]_ , \new_[18543]_ , \new_[18546]_ ,
    \new_[18547]_ , \new_[18548]_ , \new_[18552]_ , \new_[18553]_ ,
    \new_[18556]_ , \new_[18559]_ , \new_[18560]_ , \new_[18561]_ ,
    \new_[18565]_ , \new_[18566]_ , \new_[18569]_ , \new_[18572]_ ,
    \new_[18573]_ , \new_[18574]_ , \new_[18578]_ , \new_[18579]_ ,
    \new_[18582]_ , \new_[18585]_ , \new_[18586]_ , \new_[18587]_ ,
    \new_[18591]_ , \new_[18592]_ , \new_[18595]_ , \new_[18598]_ ,
    \new_[18599]_ , \new_[18600]_ , \new_[18604]_ , \new_[18605]_ ,
    \new_[18608]_ , \new_[18611]_ , \new_[18612]_ , \new_[18613]_ ,
    \new_[18617]_ , \new_[18618]_ , \new_[18621]_ , \new_[18624]_ ,
    \new_[18625]_ , \new_[18626]_ , \new_[18630]_ , \new_[18631]_ ,
    \new_[18634]_ , \new_[18637]_ , \new_[18638]_ , \new_[18639]_ ,
    \new_[18643]_ , \new_[18644]_ , \new_[18647]_ , \new_[18650]_ ,
    \new_[18651]_ , \new_[18652]_ , \new_[18656]_ , \new_[18657]_ ,
    \new_[18660]_ , \new_[18663]_ , \new_[18664]_ , \new_[18665]_ ,
    \new_[18669]_ , \new_[18670]_ , \new_[18673]_ , \new_[18676]_ ,
    \new_[18677]_ , \new_[18678]_ , \new_[18682]_ , \new_[18683]_ ,
    \new_[18686]_ , \new_[18689]_ , \new_[18690]_ , \new_[18691]_ ,
    \new_[18695]_ , \new_[18696]_ , \new_[18699]_ , \new_[18702]_ ,
    \new_[18703]_ , \new_[18704]_ , \new_[18708]_ , \new_[18709]_ ,
    \new_[18712]_ , \new_[18715]_ , \new_[18716]_ , \new_[18717]_ ,
    \new_[18721]_ , \new_[18722]_ , \new_[18725]_ , \new_[18728]_ ,
    \new_[18729]_ , \new_[18730]_ , \new_[18734]_ , \new_[18735]_ ,
    \new_[18738]_ , \new_[18741]_ , \new_[18742]_ , \new_[18743]_ ,
    \new_[18747]_ , \new_[18748]_ , \new_[18751]_ , \new_[18754]_ ,
    \new_[18755]_ , \new_[18756]_ , \new_[18760]_ , \new_[18761]_ ,
    \new_[18764]_ , \new_[18767]_ , \new_[18768]_ , \new_[18769]_ ,
    \new_[18773]_ , \new_[18774]_ , \new_[18777]_ , \new_[18780]_ ,
    \new_[18781]_ , \new_[18782]_ , \new_[18786]_ , \new_[18787]_ ,
    \new_[18790]_ , \new_[18793]_ , \new_[18794]_ , \new_[18795]_ ,
    \new_[18799]_ , \new_[18800]_ , \new_[18803]_ , \new_[18806]_ ,
    \new_[18807]_ , \new_[18808]_ , \new_[18812]_ , \new_[18813]_ ,
    \new_[18816]_ , \new_[18819]_ , \new_[18820]_ , \new_[18821]_ ,
    \new_[18825]_ , \new_[18826]_ , \new_[18829]_ , \new_[18832]_ ,
    \new_[18833]_ , \new_[18834]_ , \new_[18838]_ , \new_[18839]_ ,
    \new_[18842]_ , \new_[18845]_ , \new_[18846]_ , \new_[18847]_ ,
    \new_[18851]_ , \new_[18852]_ , \new_[18855]_ , \new_[18858]_ ,
    \new_[18859]_ , \new_[18860]_ , \new_[18864]_ , \new_[18865]_ ,
    \new_[18868]_ , \new_[18871]_ , \new_[18872]_ , \new_[18873]_ ,
    \new_[18877]_ , \new_[18878]_ , \new_[18881]_ , \new_[18884]_ ,
    \new_[18885]_ , \new_[18886]_ , \new_[18890]_ , \new_[18891]_ ,
    \new_[18894]_ , \new_[18897]_ , \new_[18898]_ , \new_[18899]_ ,
    \new_[18903]_ , \new_[18904]_ , \new_[18907]_ , \new_[18910]_ ,
    \new_[18911]_ , \new_[18912]_ , \new_[18916]_ , \new_[18917]_ ,
    \new_[18920]_ , \new_[18923]_ , \new_[18924]_ , \new_[18925]_ ,
    \new_[18929]_ , \new_[18930]_ , \new_[18933]_ , \new_[18936]_ ,
    \new_[18937]_ , \new_[18938]_ , \new_[18942]_ , \new_[18943]_ ,
    \new_[18946]_ , \new_[18949]_ , \new_[18950]_ , \new_[18951]_ ,
    \new_[18955]_ , \new_[18956]_ , \new_[18959]_ , \new_[18962]_ ,
    \new_[18963]_ , \new_[18964]_ , \new_[18968]_ , \new_[18969]_ ,
    \new_[18972]_ , \new_[18975]_ , \new_[18976]_ , \new_[18977]_ ,
    \new_[18981]_ , \new_[18982]_ , \new_[18985]_ , \new_[18988]_ ,
    \new_[18989]_ , \new_[18990]_ , \new_[18994]_ , \new_[18995]_ ,
    \new_[18998]_ , \new_[19001]_ , \new_[19002]_ , \new_[19003]_ ,
    \new_[19007]_ , \new_[19008]_ , \new_[19011]_ , \new_[19014]_ ,
    \new_[19015]_ , \new_[19016]_ , \new_[19020]_ , \new_[19021]_ ,
    \new_[19024]_ , \new_[19027]_ , \new_[19028]_ , \new_[19029]_ ,
    \new_[19033]_ , \new_[19034]_ , \new_[19037]_ , \new_[19040]_ ,
    \new_[19041]_ , \new_[19042]_ , \new_[19046]_ , \new_[19047]_ ,
    \new_[19050]_ , \new_[19053]_ , \new_[19054]_ , \new_[19055]_ ,
    \new_[19059]_ , \new_[19060]_ , \new_[19063]_ , \new_[19066]_ ,
    \new_[19067]_ , \new_[19068]_ , \new_[19072]_ , \new_[19073]_ ,
    \new_[19076]_ , \new_[19079]_ , \new_[19080]_ , \new_[19081]_ ,
    \new_[19085]_ , \new_[19086]_ , \new_[19089]_ , \new_[19092]_ ,
    \new_[19093]_ , \new_[19094]_ , \new_[19098]_ , \new_[19099]_ ,
    \new_[19102]_ , \new_[19105]_ , \new_[19106]_ , \new_[19107]_ ,
    \new_[19111]_ , \new_[19112]_ , \new_[19115]_ , \new_[19118]_ ,
    \new_[19119]_ , \new_[19120]_ , \new_[19124]_ , \new_[19125]_ ,
    \new_[19128]_ , \new_[19131]_ , \new_[19132]_ , \new_[19133]_ ,
    \new_[19137]_ , \new_[19138]_ , \new_[19141]_ , \new_[19144]_ ,
    \new_[19145]_ , \new_[19146]_ , \new_[19150]_ , \new_[19151]_ ,
    \new_[19154]_ , \new_[19157]_ , \new_[19158]_ , \new_[19159]_ ,
    \new_[19163]_ , \new_[19164]_ , \new_[19167]_ , \new_[19170]_ ,
    \new_[19171]_ , \new_[19172]_ , \new_[19176]_ , \new_[19177]_ ,
    \new_[19180]_ , \new_[19183]_ , \new_[19184]_ , \new_[19185]_ ,
    \new_[19189]_ , \new_[19190]_ , \new_[19193]_ , \new_[19196]_ ,
    \new_[19197]_ , \new_[19198]_ , \new_[19202]_ , \new_[19203]_ ,
    \new_[19206]_ , \new_[19209]_ , \new_[19210]_ , \new_[19211]_ ,
    \new_[19215]_ , \new_[19216]_ , \new_[19219]_ , \new_[19222]_ ,
    \new_[19223]_ , \new_[19224]_ , \new_[19228]_ , \new_[19229]_ ,
    \new_[19232]_ , \new_[19235]_ , \new_[19236]_ , \new_[19237]_ ,
    \new_[19241]_ , \new_[19242]_ , \new_[19245]_ , \new_[19248]_ ,
    \new_[19249]_ , \new_[19250]_ , \new_[19254]_ , \new_[19255]_ ,
    \new_[19258]_ , \new_[19261]_ , \new_[19262]_ , \new_[19263]_ ,
    \new_[19267]_ , \new_[19268]_ , \new_[19271]_ , \new_[19274]_ ,
    \new_[19275]_ , \new_[19276]_ , \new_[19280]_ , \new_[19281]_ ,
    \new_[19284]_ , \new_[19287]_ , \new_[19288]_ , \new_[19289]_ ,
    \new_[19293]_ , \new_[19294]_ , \new_[19297]_ , \new_[19300]_ ,
    \new_[19301]_ , \new_[19302]_ , \new_[19306]_ , \new_[19307]_ ,
    \new_[19310]_ , \new_[19313]_ , \new_[19314]_ , \new_[19315]_ ,
    \new_[19319]_ , \new_[19320]_ , \new_[19323]_ , \new_[19326]_ ,
    \new_[19327]_ , \new_[19328]_ , \new_[19332]_ , \new_[19333]_ ,
    \new_[19336]_ , \new_[19339]_ , \new_[19340]_ , \new_[19341]_ ,
    \new_[19345]_ , \new_[19346]_ , \new_[19349]_ , \new_[19352]_ ,
    \new_[19353]_ , \new_[19354]_ , \new_[19358]_ , \new_[19359]_ ,
    \new_[19362]_ , \new_[19365]_ , \new_[19366]_ , \new_[19367]_ ,
    \new_[19371]_ , \new_[19372]_ , \new_[19375]_ , \new_[19378]_ ,
    \new_[19379]_ , \new_[19380]_ , \new_[19384]_ , \new_[19385]_ ,
    \new_[19388]_ , \new_[19391]_ , \new_[19392]_ , \new_[19393]_ ,
    \new_[19397]_ , \new_[19398]_ , \new_[19401]_ , \new_[19404]_ ,
    \new_[19405]_ , \new_[19406]_ , \new_[19410]_ , \new_[19411]_ ,
    \new_[19414]_ , \new_[19417]_ , \new_[19418]_ , \new_[19419]_ ,
    \new_[19423]_ , \new_[19424]_ , \new_[19427]_ , \new_[19430]_ ,
    \new_[19431]_ , \new_[19432]_ , \new_[19436]_ , \new_[19437]_ ,
    \new_[19440]_ , \new_[19443]_ , \new_[19444]_ , \new_[19445]_ ,
    \new_[19449]_ , \new_[19450]_ , \new_[19453]_ , \new_[19456]_ ,
    \new_[19457]_ , \new_[19458]_ , \new_[19462]_ , \new_[19463]_ ,
    \new_[19466]_ , \new_[19469]_ , \new_[19470]_ , \new_[19471]_ ,
    \new_[19475]_ , \new_[19476]_ , \new_[19479]_ , \new_[19482]_ ,
    \new_[19483]_ , \new_[19484]_ , \new_[19488]_ , \new_[19489]_ ,
    \new_[19492]_ , \new_[19495]_ , \new_[19496]_ , \new_[19497]_ ,
    \new_[19501]_ , \new_[19502]_ , \new_[19505]_ , \new_[19508]_ ,
    \new_[19509]_ , \new_[19510]_ , \new_[19514]_ , \new_[19515]_ ,
    \new_[19518]_ , \new_[19521]_ , \new_[19522]_ , \new_[19523]_ ,
    \new_[19527]_ , \new_[19528]_ , \new_[19531]_ , \new_[19534]_ ,
    \new_[19535]_ , \new_[19536]_ , \new_[19540]_ , \new_[19541]_ ,
    \new_[19544]_ , \new_[19547]_ , \new_[19548]_ , \new_[19549]_ ,
    \new_[19553]_ , \new_[19554]_ , \new_[19557]_ , \new_[19560]_ ,
    \new_[19561]_ , \new_[19562]_ , \new_[19566]_ , \new_[19567]_ ,
    \new_[19570]_ , \new_[19573]_ , \new_[19574]_ , \new_[19575]_ ,
    \new_[19579]_ , \new_[19580]_ , \new_[19583]_ , \new_[19586]_ ,
    \new_[19587]_ , \new_[19588]_ , \new_[19592]_ , \new_[19593]_ ,
    \new_[19596]_ , \new_[19599]_ , \new_[19600]_ , \new_[19601]_ ,
    \new_[19605]_ , \new_[19606]_ , \new_[19609]_ , \new_[19612]_ ,
    \new_[19613]_ , \new_[19614]_ , \new_[19618]_ , \new_[19619]_ ,
    \new_[19622]_ , \new_[19625]_ , \new_[19626]_ , \new_[19627]_ ,
    \new_[19631]_ , \new_[19632]_ , \new_[19635]_ , \new_[19638]_ ,
    \new_[19639]_ , \new_[19640]_ , \new_[19644]_ , \new_[19645]_ ,
    \new_[19648]_ , \new_[19651]_ , \new_[19652]_ , \new_[19653]_ ,
    \new_[19657]_ , \new_[19658]_ , \new_[19661]_ , \new_[19664]_ ,
    \new_[19665]_ , \new_[19666]_ , \new_[19670]_ , \new_[19671]_ ,
    \new_[19674]_ , \new_[19677]_ , \new_[19678]_ , \new_[19679]_ ,
    \new_[19683]_ , \new_[19684]_ , \new_[19687]_ , \new_[19690]_ ,
    \new_[19691]_ , \new_[19692]_ , \new_[19696]_ , \new_[19697]_ ,
    \new_[19700]_ , \new_[19703]_ , \new_[19704]_ , \new_[19705]_ ,
    \new_[19709]_ , \new_[19710]_ , \new_[19713]_ , \new_[19716]_ ,
    \new_[19717]_ , \new_[19718]_ , \new_[19722]_ , \new_[19723]_ ,
    \new_[19726]_ , \new_[19729]_ , \new_[19730]_ , \new_[19731]_ ,
    \new_[19735]_ , \new_[19736]_ , \new_[19739]_ , \new_[19742]_ ,
    \new_[19743]_ , \new_[19744]_ , \new_[19748]_ , \new_[19749]_ ,
    \new_[19752]_ , \new_[19755]_ , \new_[19756]_ , \new_[19757]_ ,
    \new_[19761]_ , \new_[19762]_ , \new_[19765]_ , \new_[19768]_ ,
    \new_[19769]_ , \new_[19770]_ , \new_[19774]_ , \new_[19775]_ ,
    \new_[19778]_ , \new_[19781]_ , \new_[19782]_ , \new_[19783]_ ,
    \new_[19787]_ , \new_[19788]_ , \new_[19791]_ , \new_[19794]_ ,
    \new_[19795]_ , \new_[19796]_ , \new_[19800]_ , \new_[19801]_ ,
    \new_[19804]_ , \new_[19807]_ , \new_[19808]_ , \new_[19809]_ ,
    \new_[19813]_ , \new_[19814]_ , \new_[19817]_ , \new_[19820]_ ,
    \new_[19821]_ , \new_[19822]_ , \new_[19826]_ , \new_[19827]_ ,
    \new_[19830]_ , \new_[19833]_ , \new_[19834]_ , \new_[19835]_ ,
    \new_[19839]_ , \new_[19840]_ , \new_[19843]_ , \new_[19846]_ ,
    \new_[19847]_ , \new_[19848]_ , \new_[19852]_ , \new_[19853]_ ,
    \new_[19856]_ , \new_[19859]_ , \new_[19860]_ , \new_[19861]_ ,
    \new_[19865]_ , \new_[19866]_ , \new_[19869]_ , \new_[19872]_ ,
    \new_[19873]_ , \new_[19874]_ , \new_[19878]_ , \new_[19879]_ ,
    \new_[19882]_ , \new_[19885]_ , \new_[19886]_ , \new_[19887]_ ,
    \new_[19891]_ , \new_[19892]_ , \new_[19895]_ , \new_[19898]_ ,
    \new_[19899]_ , \new_[19900]_ , \new_[19904]_ , \new_[19905]_ ,
    \new_[19908]_ , \new_[19911]_ , \new_[19912]_ , \new_[19913]_ ,
    \new_[19917]_ , \new_[19918]_ , \new_[19921]_ , \new_[19924]_ ,
    \new_[19925]_ , \new_[19926]_ , \new_[19930]_ , \new_[19931]_ ,
    \new_[19934]_ , \new_[19937]_ , \new_[19938]_ , \new_[19939]_ ,
    \new_[19943]_ , \new_[19944]_ , \new_[19947]_ , \new_[19950]_ ,
    \new_[19951]_ , \new_[19952]_ , \new_[19956]_ , \new_[19957]_ ,
    \new_[19960]_ , \new_[19963]_ , \new_[19964]_ , \new_[19965]_ ,
    \new_[19969]_ , \new_[19970]_ , \new_[19973]_ , \new_[19976]_ ,
    \new_[19977]_ , \new_[19978]_ , \new_[19982]_ , \new_[19983]_ ,
    \new_[19986]_ , \new_[19989]_ , \new_[19990]_ , \new_[19991]_ ,
    \new_[19995]_ , \new_[19996]_ , \new_[19999]_ , \new_[20002]_ ,
    \new_[20003]_ , \new_[20004]_ , \new_[20008]_ , \new_[20009]_ ,
    \new_[20012]_ , \new_[20015]_ , \new_[20016]_ , \new_[20017]_ ,
    \new_[20021]_ , \new_[20022]_ , \new_[20025]_ , \new_[20028]_ ,
    \new_[20029]_ , \new_[20030]_ , \new_[20034]_ , \new_[20035]_ ,
    \new_[20038]_ , \new_[20041]_ , \new_[20042]_ , \new_[20043]_ ,
    \new_[20047]_ , \new_[20048]_ , \new_[20051]_ , \new_[20054]_ ,
    \new_[20055]_ , \new_[20056]_ , \new_[20060]_ , \new_[20061]_ ,
    \new_[20064]_ , \new_[20067]_ , \new_[20068]_ , \new_[20069]_ ,
    \new_[20073]_ , \new_[20074]_ , \new_[20077]_ , \new_[20080]_ ,
    \new_[20081]_ , \new_[20082]_ , \new_[20086]_ , \new_[20087]_ ,
    \new_[20090]_ , \new_[20093]_ , \new_[20094]_ , \new_[20095]_ ,
    \new_[20099]_ , \new_[20100]_ , \new_[20103]_ , \new_[20106]_ ,
    \new_[20107]_ , \new_[20108]_ , \new_[20112]_ , \new_[20113]_ ,
    \new_[20116]_ , \new_[20119]_ , \new_[20120]_ , \new_[20121]_ ,
    \new_[20125]_ , \new_[20126]_ , \new_[20129]_ , \new_[20132]_ ,
    \new_[20133]_ , \new_[20134]_ , \new_[20138]_ , \new_[20139]_ ,
    \new_[20142]_ , \new_[20145]_ , \new_[20146]_ , \new_[20147]_ ,
    \new_[20151]_ , \new_[20152]_ , \new_[20155]_ , \new_[20158]_ ,
    \new_[20159]_ , \new_[20160]_ , \new_[20164]_ , \new_[20165]_ ,
    \new_[20168]_ , \new_[20171]_ , \new_[20172]_ , \new_[20173]_ ,
    \new_[20177]_ , \new_[20178]_ , \new_[20181]_ , \new_[20184]_ ,
    \new_[20185]_ , \new_[20186]_ , \new_[20190]_ , \new_[20191]_ ,
    \new_[20194]_ , \new_[20197]_ , \new_[20198]_ , \new_[20199]_ ,
    \new_[20203]_ , \new_[20204]_ , \new_[20207]_ , \new_[20210]_ ,
    \new_[20211]_ , \new_[20212]_ , \new_[20216]_ , \new_[20217]_ ,
    \new_[20220]_ , \new_[20223]_ , \new_[20224]_ , \new_[20225]_ ,
    \new_[20228]_ , \new_[20231]_ , \new_[20232]_ , \new_[20235]_ ,
    \new_[20238]_ , \new_[20239]_ , \new_[20240]_ , \new_[20244]_ ,
    \new_[20245]_ , \new_[20248]_ , \new_[20251]_ , \new_[20252]_ ,
    \new_[20253]_ , \new_[20256]_ , \new_[20259]_ , \new_[20260]_ ,
    \new_[20263]_ , \new_[20266]_ , \new_[20267]_ , \new_[20268]_ ,
    \new_[20272]_ , \new_[20273]_ , \new_[20276]_ , \new_[20279]_ ,
    \new_[20280]_ , \new_[20281]_ , \new_[20284]_ , \new_[20287]_ ,
    \new_[20288]_ , \new_[20291]_ , \new_[20294]_ , \new_[20295]_ ,
    \new_[20296]_ , \new_[20300]_ , \new_[20301]_ , \new_[20304]_ ,
    \new_[20307]_ , \new_[20308]_ , \new_[20309]_ , \new_[20312]_ ,
    \new_[20315]_ , \new_[20316]_ , \new_[20319]_ , \new_[20322]_ ,
    \new_[20323]_ , \new_[20324]_ , \new_[20328]_ , \new_[20329]_ ,
    \new_[20332]_ , \new_[20335]_ , \new_[20336]_ , \new_[20337]_ ,
    \new_[20340]_ , \new_[20343]_ , \new_[20344]_ , \new_[20347]_ ,
    \new_[20350]_ , \new_[20351]_ , \new_[20352]_ , \new_[20356]_ ,
    \new_[20357]_ , \new_[20360]_ , \new_[20363]_ , \new_[20364]_ ,
    \new_[20365]_ , \new_[20368]_ , \new_[20371]_ , \new_[20372]_ ,
    \new_[20375]_ , \new_[20378]_ , \new_[20379]_ , \new_[20380]_ ,
    \new_[20384]_ , \new_[20385]_ , \new_[20388]_ , \new_[20391]_ ,
    \new_[20392]_ , \new_[20393]_ , \new_[20396]_ , \new_[20399]_ ,
    \new_[20400]_ , \new_[20403]_ , \new_[20406]_ , \new_[20407]_ ,
    \new_[20408]_ , \new_[20412]_ , \new_[20413]_ , \new_[20416]_ ,
    \new_[20419]_ , \new_[20420]_ , \new_[20421]_ , \new_[20424]_ ,
    \new_[20427]_ , \new_[20428]_ , \new_[20431]_ , \new_[20434]_ ,
    \new_[20435]_ , \new_[20436]_ , \new_[20440]_ , \new_[20441]_ ,
    \new_[20444]_ , \new_[20447]_ , \new_[20448]_ , \new_[20449]_ ,
    \new_[20452]_ , \new_[20455]_ , \new_[20456]_ , \new_[20459]_ ,
    \new_[20462]_ , \new_[20463]_ , \new_[20464]_ , \new_[20468]_ ,
    \new_[20469]_ , \new_[20472]_ , \new_[20475]_ , \new_[20476]_ ,
    \new_[20477]_ , \new_[20480]_ , \new_[20483]_ , \new_[20484]_ ,
    \new_[20487]_ , \new_[20490]_ , \new_[20491]_ , \new_[20492]_ ,
    \new_[20496]_ , \new_[20497]_ , \new_[20500]_ , \new_[20503]_ ,
    \new_[20504]_ , \new_[20505]_ , \new_[20508]_ , \new_[20511]_ ,
    \new_[20512]_ , \new_[20515]_ , \new_[20518]_ , \new_[20519]_ ,
    \new_[20520]_ , \new_[20524]_ , \new_[20525]_ , \new_[20528]_ ,
    \new_[20531]_ , \new_[20532]_ , \new_[20533]_ , \new_[20536]_ ,
    \new_[20539]_ , \new_[20540]_ , \new_[20543]_ , \new_[20546]_ ,
    \new_[20547]_ , \new_[20548]_ , \new_[20552]_ , \new_[20553]_ ,
    \new_[20556]_ , \new_[20559]_ , \new_[20560]_ , \new_[20561]_ ,
    \new_[20564]_ , \new_[20567]_ , \new_[20568]_ , \new_[20571]_ ,
    \new_[20574]_ , \new_[20575]_ , \new_[20576]_ , \new_[20580]_ ,
    \new_[20581]_ , \new_[20584]_ , \new_[20587]_ , \new_[20588]_ ,
    \new_[20589]_ , \new_[20592]_ , \new_[20595]_ , \new_[20596]_ ,
    \new_[20599]_ , \new_[20602]_ , \new_[20603]_ , \new_[20604]_ ,
    \new_[20608]_ , \new_[20609]_ , \new_[20612]_ , \new_[20615]_ ,
    \new_[20616]_ , \new_[20617]_ , \new_[20620]_ , \new_[20623]_ ,
    \new_[20624]_ , \new_[20627]_ , \new_[20630]_ , \new_[20631]_ ,
    \new_[20632]_ , \new_[20636]_ , \new_[20637]_ , \new_[20640]_ ,
    \new_[20643]_ , \new_[20644]_ , \new_[20645]_ , \new_[20648]_ ,
    \new_[20651]_ , \new_[20652]_ , \new_[20655]_ , \new_[20658]_ ,
    \new_[20659]_ , \new_[20660]_ , \new_[20664]_ , \new_[20665]_ ,
    \new_[20668]_ , \new_[20671]_ , \new_[20672]_ , \new_[20673]_ ,
    \new_[20676]_ , \new_[20679]_ , \new_[20680]_ , \new_[20683]_ ,
    \new_[20686]_ , \new_[20687]_ , \new_[20688]_ , \new_[20692]_ ,
    \new_[20693]_ , \new_[20696]_ , \new_[20699]_ , \new_[20700]_ ,
    \new_[20701]_ , \new_[20704]_ , \new_[20707]_ , \new_[20708]_ ,
    \new_[20711]_ , \new_[20714]_ , \new_[20715]_ , \new_[20716]_ ,
    \new_[20720]_ , \new_[20721]_ , \new_[20724]_ , \new_[20727]_ ,
    \new_[20728]_ , \new_[20729]_ , \new_[20732]_ , \new_[20735]_ ,
    \new_[20736]_ , \new_[20739]_ , \new_[20742]_ , \new_[20743]_ ,
    \new_[20744]_ , \new_[20748]_ , \new_[20749]_ , \new_[20752]_ ,
    \new_[20755]_ , \new_[20756]_ , \new_[20757]_ , \new_[20760]_ ,
    \new_[20763]_ , \new_[20764]_ , \new_[20767]_ , \new_[20770]_ ,
    \new_[20771]_ , \new_[20772]_ , \new_[20776]_ , \new_[20777]_ ,
    \new_[20780]_ , \new_[20783]_ , \new_[20784]_ , \new_[20785]_ ,
    \new_[20788]_ , \new_[20791]_ , \new_[20792]_ , \new_[20795]_ ,
    \new_[20798]_ , \new_[20799]_ , \new_[20800]_ , \new_[20804]_ ,
    \new_[20805]_ , \new_[20808]_ , \new_[20811]_ , \new_[20812]_ ,
    \new_[20813]_ , \new_[20816]_ , \new_[20819]_ , \new_[20820]_ ,
    \new_[20823]_ , \new_[20826]_ , \new_[20827]_ , \new_[20828]_ ,
    \new_[20832]_ , \new_[20833]_ , \new_[20836]_ , \new_[20839]_ ,
    \new_[20840]_ , \new_[20841]_ , \new_[20844]_ , \new_[20847]_ ,
    \new_[20848]_ , \new_[20851]_ , \new_[20854]_ , \new_[20855]_ ,
    \new_[20856]_ , \new_[20860]_ , \new_[20861]_ , \new_[20864]_ ,
    \new_[20867]_ , \new_[20868]_ , \new_[20869]_ , \new_[20872]_ ,
    \new_[20875]_ , \new_[20876]_ , \new_[20879]_ , \new_[20882]_ ,
    \new_[20883]_ , \new_[20884]_ , \new_[20888]_ , \new_[20889]_ ,
    \new_[20892]_ , \new_[20895]_ , \new_[20896]_ , \new_[20897]_ ,
    \new_[20900]_ , \new_[20903]_ , \new_[20904]_ , \new_[20907]_ ,
    \new_[20910]_ , \new_[20911]_ , \new_[20912]_ , \new_[20916]_ ,
    \new_[20917]_ , \new_[20920]_ , \new_[20923]_ , \new_[20924]_ ,
    \new_[20925]_ , \new_[20928]_ , \new_[20931]_ , \new_[20932]_ ,
    \new_[20935]_ , \new_[20938]_ , \new_[20939]_ , \new_[20940]_ ,
    \new_[20944]_ , \new_[20945]_ , \new_[20948]_ , \new_[20951]_ ,
    \new_[20952]_ , \new_[20953]_ , \new_[20956]_ , \new_[20959]_ ,
    \new_[20960]_ , \new_[20963]_ , \new_[20966]_ , \new_[20967]_ ,
    \new_[20968]_ , \new_[20972]_ , \new_[20973]_ , \new_[20976]_ ,
    \new_[20979]_ , \new_[20980]_ , \new_[20981]_ , \new_[20984]_ ,
    \new_[20987]_ , \new_[20988]_ , \new_[20991]_ , \new_[20994]_ ,
    \new_[20995]_ , \new_[20996]_ , \new_[21000]_ , \new_[21001]_ ,
    \new_[21004]_ , \new_[21007]_ , \new_[21008]_ , \new_[21009]_ ,
    \new_[21012]_ , \new_[21015]_ , \new_[21016]_ , \new_[21019]_ ,
    \new_[21022]_ , \new_[21023]_ , \new_[21024]_ , \new_[21028]_ ,
    \new_[21029]_ , \new_[21032]_ , \new_[21035]_ , \new_[21036]_ ,
    \new_[21037]_ , \new_[21040]_ , \new_[21043]_ , \new_[21044]_ ,
    \new_[21047]_ , \new_[21050]_ , \new_[21051]_ , \new_[21052]_ ,
    \new_[21056]_ , \new_[21057]_ , \new_[21060]_ , \new_[21063]_ ,
    \new_[21064]_ , \new_[21065]_ , \new_[21068]_ , \new_[21071]_ ,
    \new_[21072]_ , \new_[21075]_ , \new_[21078]_ , \new_[21079]_ ,
    \new_[21080]_ , \new_[21084]_ , \new_[21085]_ , \new_[21088]_ ,
    \new_[21091]_ , \new_[21092]_ , \new_[21093]_ , \new_[21096]_ ,
    \new_[21099]_ , \new_[21100]_ , \new_[21103]_ , \new_[21106]_ ,
    \new_[21107]_ , \new_[21108]_ , \new_[21112]_ , \new_[21113]_ ,
    \new_[21116]_ , \new_[21119]_ , \new_[21120]_ , \new_[21121]_ ,
    \new_[21124]_ , \new_[21127]_ , \new_[21128]_ , \new_[21131]_ ,
    \new_[21134]_ , \new_[21135]_ , \new_[21136]_ , \new_[21140]_ ,
    \new_[21141]_ , \new_[21144]_ , \new_[21147]_ , \new_[21148]_ ,
    \new_[21149]_ , \new_[21152]_ , \new_[21155]_ , \new_[21156]_ ,
    \new_[21159]_ , \new_[21162]_ , \new_[21163]_ , \new_[21164]_ ,
    \new_[21168]_ , \new_[21169]_ , \new_[21172]_ , \new_[21175]_ ,
    \new_[21176]_ , \new_[21177]_ , \new_[21180]_ , \new_[21183]_ ,
    \new_[21184]_ , \new_[21187]_ , \new_[21190]_ , \new_[21191]_ ,
    \new_[21192]_ , \new_[21196]_ , \new_[21197]_ , \new_[21200]_ ,
    \new_[21203]_ , \new_[21204]_ , \new_[21205]_ , \new_[21208]_ ,
    \new_[21211]_ , \new_[21212]_ , \new_[21215]_ , \new_[21218]_ ,
    \new_[21219]_ , \new_[21220]_ , \new_[21224]_ , \new_[21225]_ ,
    \new_[21228]_ , \new_[21231]_ , \new_[21232]_ , \new_[21233]_ ,
    \new_[21236]_ , \new_[21239]_ , \new_[21240]_ , \new_[21243]_ ,
    \new_[21246]_ , \new_[21247]_ , \new_[21248]_ , \new_[21252]_ ,
    \new_[21253]_ , \new_[21256]_ , \new_[21259]_ , \new_[21260]_ ,
    \new_[21261]_ , \new_[21264]_ , \new_[21267]_ , \new_[21268]_ ,
    \new_[21271]_ , \new_[21274]_ , \new_[21275]_ , \new_[21276]_ ,
    \new_[21280]_ , \new_[21281]_ , \new_[21284]_ , \new_[21287]_ ,
    \new_[21288]_ , \new_[21289]_ , \new_[21292]_ , \new_[21295]_ ,
    \new_[21296]_ , \new_[21299]_ , \new_[21302]_ , \new_[21303]_ ,
    \new_[21304]_ , \new_[21308]_ , \new_[21309]_ , \new_[21312]_ ,
    \new_[21315]_ , \new_[21316]_ , \new_[21317]_ , \new_[21320]_ ,
    \new_[21323]_ , \new_[21324]_ , \new_[21327]_ , \new_[21330]_ ,
    \new_[21331]_ , \new_[21332]_ , \new_[21336]_ , \new_[21337]_ ,
    \new_[21340]_ , \new_[21343]_ , \new_[21344]_ , \new_[21345]_ ,
    \new_[21348]_ , \new_[21351]_ , \new_[21352]_ , \new_[21355]_ ,
    \new_[21358]_ , \new_[21359]_ , \new_[21360]_ , \new_[21364]_ ,
    \new_[21365]_ , \new_[21368]_ , \new_[21371]_ , \new_[21372]_ ,
    \new_[21373]_ , \new_[21376]_ , \new_[21379]_ , \new_[21380]_ ,
    \new_[21383]_ , \new_[21386]_ , \new_[21387]_ , \new_[21388]_ ,
    \new_[21392]_ , \new_[21393]_ , \new_[21396]_ , \new_[21399]_ ,
    \new_[21400]_ , \new_[21401]_ , \new_[21404]_ , \new_[21407]_ ,
    \new_[21408]_ , \new_[21411]_ , \new_[21414]_ , \new_[21415]_ ,
    \new_[21416]_ , \new_[21420]_ , \new_[21421]_ , \new_[21424]_ ,
    \new_[21427]_ , \new_[21428]_ , \new_[21429]_ , \new_[21432]_ ,
    \new_[21435]_ , \new_[21436]_ , \new_[21439]_ , \new_[21442]_ ,
    \new_[21443]_ , \new_[21444]_ , \new_[21448]_ , \new_[21449]_ ,
    \new_[21452]_ , \new_[21455]_ , \new_[21456]_ , \new_[21457]_ ,
    \new_[21460]_ , \new_[21463]_ , \new_[21464]_ , \new_[21467]_ ,
    \new_[21470]_ , \new_[21471]_ , \new_[21472]_ , \new_[21476]_ ,
    \new_[21477]_ , \new_[21480]_ , \new_[21483]_ , \new_[21484]_ ,
    \new_[21485]_ , \new_[21488]_ , \new_[21491]_ , \new_[21492]_ ,
    \new_[21495]_ , \new_[21498]_ , \new_[21499]_ , \new_[21500]_ ,
    \new_[21504]_ , \new_[21505]_ , \new_[21508]_ , \new_[21511]_ ,
    \new_[21512]_ , \new_[21513]_ , \new_[21516]_ , \new_[21519]_ ,
    \new_[21520]_ , \new_[21523]_ , \new_[21526]_ , \new_[21527]_ ,
    \new_[21528]_ , \new_[21532]_ , \new_[21533]_ , \new_[21536]_ ,
    \new_[21539]_ , \new_[21540]_ , \new_[21541]_ , \new_[21544]_ ,
    \new_[21547]_ , \new_[21548]_ , \new_[21551]_ , \new_[21554]_ ,
    \new_[21555]_ , \new_[21556]_ , \new_[21560]_ , \new_[21561]_ ,
    \new_[21564]_ , \new_[21567]_ , \new_[21568]_ , \new_[21569]_ ,
    \new_[21572]_ , \new_[21575]_ , \new_[21576]_ , \new_[21579]_ ,
    \new_[21582]_ , \new_[21583]_ , \new_[21584]_ , \new_[21588]_ ,
    \new_[21589]_ , \new_[21592]_ , \new_[21595]_ , \new_[21596]_ ,
    \new_[21597]_ , \new_[21600]_ , \new_[21603]_ , \new_[21604]_ ,
    \new_[21607]_ , \new_[21610]_ , \new_[21611]_ , \new_[21612]_ ,
    \new_[21616]_ , \new_[21617]_ , \new_[21620]_ , \new_[21623]_ ,
    \new_[21624]_ , \new_[21625]_ , \new_[21628]_ , \new_[21631]_ ,
    \new_[21632]_ , \new_[21635]_ , \new_[21638]_ , \new_[21639]_ ,
    \new_[21640]_ , \new_[21644]_ , \new_[21645]_ , \new_[21648]_ ,
    \new_[21651]_ , \new_[21652]_ , \new_[21653]_ , \new_[21656]_ ,
    \new_[21659]_ , \new_[21660]_ , \new_[21663]_ , \new_[21666]_ ,
    \new_[21667]_ , \new_[21668]_ , \new_[21672]_ , \new_[21673]_ ,
    \new_[21676]_ , \new_[21679]_ , \new_[21680]_ , \new_[21681]_ ,
    \new_[21684]_ , \new_[21687]_ , \new_[21688]_ , \new_[21691]_ ,
    \new_[21694]_ , \new_[21695]_ , \new_[21696]_ , \new_[21700]_ ,
    \new_[21701]_ , \new_[21704]_ , \new_[21707]_ , \new_[21708]_ ,
    \new_[21709]_ , \new_[21712]_ , \new_[21715]_ , \new_[21716]_ ,
    \new_[21719]_ , \new_[21722]_ , \new_[21723]_ , \new_[21724]_ ,
    \new_[21728]_ , \new_[21729]_ , \new_[21732]_ , \new_[21735]_ ,
    \new_[21736]_ , \new_[21737]_ , \new_[21740]_ , \new_[21743]_ ,
    \new_[21744]_ , \new_[21747]_ , \new_[21750]_ , \new_[21751]_ ,
    \new_[21752]_ , \new_[21756]_ , \new_[21757]_ , \new_[21760]_ ,
    \new_[21763]_ , \new_[21764]_ , \new_[21765]_ , \new_[21768]_ ,
    \new_[21771]_ , \new_[21772]_ , \new_[21775]_ , \new_[21778]_ ,
    \new_[21779]_ , \new_[21780]_ , \new_[21784]_ , \new_[21785]_ ,
    \new_[21788]_ , \new_[21791]_ , \new_[21792]_ , \new_[21793]_ ,
    \new_[21796]_ , \new_[21799]_ , \new_[21800]_ , \new_[21803]_ ,
    \new_[21806]_ , \new_[21807]_ , \new_[21808]_ , \new_[21812]_ ,
    \new_[21813]_ , \new_[21816]_ , \new_[21819]_ , \new_[21820]_ ,
    \new_[21821]_ , \new_[21824]_ , \new_[21827]_ , \new_[21828]_ ,
    \new_[21831]_ , \new_[21834]_ , \new_[21835]_ , \new_[21836]_ ,
    \new_[21840]_ , \new_[21841]_ , \new_[21844]_ , \new_[21847]_ ,
    \new_[21848]_ , \new_[21849]_ , \new_[21852]_ , \new_[21855]_ ,
    \new_[21856]_ , \new_[21859]_ , \new_[21862]_ , \new_[21863]_ ,
    \new_[21864]_ , \new_[21868]_ , \new_[21869]_ , \new_[21872]_ ,
    \new_[21875]_ , \new_[21876]_ , \new_[21877]_ , \new_[21880]_ ,
    \new_[21883]_ , \new_[21884]_ , \new_[21887]_ , \new_[21890]_ ,
    \new_[21891]_ , \new_[21892]_ , \new_[21896]_ , \new_[21897]_ ,
    \new_[21900]_ , \new_[21903]_ , \new_[21904]_ , \new_[21905]_ ,
    \new_[21908]_ , \new_[21911]_ , \new_[21912]_ , \new_[21915]_ ,
    \new_[21918]_ , \new_[21919]_ , \new_[21920]_ , \new_[21924]_ ,
    \new_[21925]_ , \new_[21928]_ , \new_[21931]_ , \new_[21932]_ ,
    \new_[21933]_ , \new_[21936]_ , \new_[21939]_ , \new_[21940]_ ,
    \new_[21943]_ , \new_[21946]_ , \new_[21947]_ , \new_[21948]_ ,
    \new_[21952]_ , \new_[21953]_ , \new_[21956]_ , \new_[21959]_ ,
    \new_[21960]_ , \new_[21961]_ , \new_[21964]_ , \new_[21967]_ ,
    \new_[21968]_ , \new_[21971]_ , \new_[21974]_ , \new_[21975]_ ,
    \new_[21976]_ , \new_[21980]_ , \new_[21981]_ , \new_[21984]_ ,
    \new_[21987]_ , \new_[21988]_ , \new_[21989]_ , \new_[21992]_ ,
    \new_[21995]_ , \new_[21996]_ , \new_[21999]_ , \new_[22002]_ ,
    \new_[22003]_ , \new_[22004]_ , \new_[22008]_ , \new_[22009]_ ,
    \new_[22012]_ , \new_[22015]_ , \new_[22016]_ , \new_[22017]_ ,
    \new_[22020]_ , \new_[22023]_ , \new_[22024]_ , \new_[22027]_ ,
    \new_[22030]_ , \new_[22031]_ , \new_[22032]_ , \new_[22036]_ ,
    \new_[22037]_ , \new_[22040]_ , \new_[22043]_ , \new_[22044]_ ,
    \new_[22045]_ , \new_[22048]_ , \new_[22051]_ , \new_[22052]_ ,
    \new_[22055]_ , \new_[22058]_ , \new_[22059]_ , \new_[22060]_ ,
    \new_[22064]_ , \new_[22065]_ , \new_[22068]_ , \new_[22071]_ ,
    \new_[22072]_ , \new_[22073]_ , \new_[22076]_ , \new_[22079]_ ,
    \new_[22080]_ , \new_[22083]_ , \new_[22086]_ , \new_[22087]_ ,
    \new_[22088]_ , \new_[22092]_ , \new_[22093]_ , \new_[22096]_ ,
    \new_[22099]_ , \new_[22100]_ , \new_[22101]_ , \new_[22104]_ ,
    \new_[22107]_ , \new_[22108]_ , \new_[22111]_ , \new_[22114]_ ,
    \new_[22115]_ , \new_[22116]_ , \new_[22120]_ , \new_[22121]_ ,
    \new_[22124]_ , \new_[22127]_ , \new_[22128]_ , \new_[22129]_ ,
    \new_[22132]_ , \new_[22135]_ , \new_[22136]_ , \new_[22139]_ ,
    \new_[22142]_ , \new_[22143]_ , \new_[22144]_ , \new_[22148]_ ,
    \new_[22149]_ , \new_[22152]_ , \new_[22155]_ , \new_[22156]_ ,
    \new_[22157]_ , \new_[22160]_ , \new_[22163]_ , \new_[22164]_ ,
    \new_[22167]_ , \new_[22170]_ , \new_[22171]_ , \new_[22172]_ ,
    \new_[22176]_ , \new_[22177]_ , \new_[22180]_ , \new_[22183]_ ,
    \new_[22184]_ , \new_[22185]_ , \new_[22188]_ , \new_[22191]_ ,
    \new_[22192]_ , \new_[22195]_ , \new_[22198]_ , \new_[22199]_ ,
    \new_[22200]_ , \new_[22204]_ , \new_[22205]_ , \new_[22208]_ ,
    \new_[22211]_ , \new_[22212]_ , \new_[22213]_ , \new_[22216]_ ,
    \new_[22219]_ , \new_[22220]_ , \new_[22223]_ , \new_[22226]_ ,
    \new_[22227]_ , \new_[22228]_ , \new_[22232]_ , \new_[22233]_ ,
    \new_[22236]_ , \new_[22239]_ , \new_[22240]_ , \new_[22241]_ ,
    \new_[22244]_ , \new_[22247]_ , \new_[22248]_ , \new_[22251]_ ,
    \new_[22254]_ , \new_[22255]_ , \new_[22256]_ , \new_[22260]_ ,
    \new_[22261]_ , \new_[22264]_ , \new_[22267]_ , \new_[22268]_ ,
    \new_[22269]_ , \new_[22272]_ , \new_[22275]_ , \new_[22276]_ ,
    \new_[22279]_ , \new_[22282]_ , \new_[22283]_ , \new_[22284]_ ,
    \new_[22288]_ , \new_[22289]_ , \new_[22292]_ , \new_[22295]_ ,
    \new_[22296]_ , \new_[22297]_ , \new_[22300]_ , \new_[22303]_ ,
    \new_[22304]_ , \new_[22307]_ , \new_[22310]_ , \new_[22311]_ ,
    \new_[22312]_ , \new_[22316]_ , \new_[22317]_ , \new_[22320]_ ,
    \new_[22323]_ , \new_[22324]_ , \new_[22325]_ , \new_[22328]_ ,
    \new_[22331]_ , \new_[22332]_ , \new_[22335]_ , \new_[22338]_ ,
    \new_[22339]_ , \new_[22340]_ , \new_[22344]_ , \new_[22345]_ ,
    \new_[22348]_ , \new_[22351]_ , \new_[22352]_ , \new_[22353]_ ,
    \new_[22356]_ , \new_[22359]_ , \new_[22360]_ , \new_[22363]_ ,
    \new_[22366]_ , \new_[22367]_ , \new_[22368]_ , \new_[22372]_ ,
    \new_[22373]_ , \new_[22376]_ , \new_[22379]_ , \new_[22380]_ ,
    \new_[22381]_ , \new_[22384]_ , \new_[22387]_ , \new_[22388]_ ,
    \new_[22391]_ , \new_[22394]_ , \new_[22395]_ , \new_[22396]_ ,
    \new_[22400]_ , \new_[22401]_ , \new_[22404]_ , \new_[22407]_ ,
    \new_[22408]_ , \new_[22409]_ , \new_[22412]_ , \new_[22415]_ ,
    \new_[22416]_ , \new_[22419]_ , \new_[22422]_ , \new_[22423]_ ,
    \new_[22424]_ , \new_[22428]_ , \new_[22429]_ , \new_[22432]_ ,
    \new_[22435]_ , \new_[22436]_ , \new_[22437]_ , \new_[22440]_ ,
    \new_[22443]_ , \new_[22444]_ , \new_[22447]_ , \new_[22450]_ ,
    \new_[22451]_ , \new_[22452]_ , \new_[22456]_ , \new_[22457]_ ,
    \new_[22460]_ , \new_[22463]_ , \new_[22464]_ , \new_[22465]_ ,
    \new_[22468]_ , \new_[22471]_ , \new_[22472]_ , \new_[22475]_ ,
    \new_[22478]_ , \new_[22479]_ , \new_[22480]_ , \new_[22484]_ ,
    \new_[22485]_ , \new_[22488]_ , \new_[22491]_ , \new_[22492]_ ,
    \new_[22493]_ , \new_[22496]_ , \new_[22499]_ , \new_[22500]_ ,
    \new_[22503]_ , \new_[22506]_ , \new_[22507]_ , \new_[22508]_ ,
    \new_[22512]_ , \new_[22513]_ , \new_[22516]_ , \new_[22519]_ ,
    \new_[22520]_ , \new_[22521]_ , \new_[22524]_ , \new_[22527]_ ,
    \new_[22528]_ , \new_[22531]_ , \new_[22534]_ , \new_[22535]_ ,
    \new_[22536]_ , \new_[22540]_ , \new_[22541]_ , \new_[22544]_ ,
    \new_[22547]_ , \new_[22548]_ , \new_[22549]_ , \new_[22552]_ ,
    \new_[22555]_ , \new_[22556]_ , \new_[22559]_ , \new_[22562]_ ,
    \new_[22563]_ , \new_[22564]_ , \new_[22568]_ , \new_[22569]_ ,
    \new_[22572]_ , \new_[22575]_ , \new_[22576]_ , \new_[22577]_ ,
    \new_[22580]_ , \new_[22583]_ , \new_[22584]_ , \new_[22587]_ ,
    \new_[22590]_ , \new_[22591]_ , \new_[22592]_ , \new_[22596]_ ,
    \new_[22597]_ , \new_[22600]_ , \new_[22603]_ , \new_[22604]_ ,
    \new_[22605]_ , \new_[22608]_ , \new_[22611]_ , \new_[22612]_ ,
    \new_[22615]_ , \new_[22618]_ , \new_[22619]_ , \new_[22620]_ ,
    \new_[22624]_ , \new_[22625]_ , \new_[22628]_ , \new_[22631]_ ,
    \new_[22632]_ , \new_[22633]_ , \new_[22636]_ , \new_[22639]_ ,
    \new_[22640]_ , \new_[22643]_ , \new_[22646]_ , \new_[22647]_ ,
    \new_[22648]_ , \new_[22652]_ , \new_[22653]_ , \new_[22656]_ ,
    \new_[22659]_ , \new_[22660]_ , \new_[22661]_ , \new_[22664]_ ,
    \new_[22667]_ , \new_[22668]_ , \new_[22671]_ , \new_[22674]_ ,
    \new_[22675]_ , \new_[22676]_ , \new_[22680]_ , \new_[22681]_ ,
    \new_[22684]_ , \new_[22687]_ , \new_[22688]_ , \new_[22689]_ ,
    \new_[22692]_ , \new_[22695]_ , \new_[22696]_ , \new_[22699]_ ,
    \new_[22702]_ , \new_[22703]_ , \new_[22704]_ , \new_[22708]_ ,
    \new_[22709]_ , \new_[22712]_ , \new_[22715]_ , \new_[22716]_ ,
    \new_[22717]_ , \new_[22720]_ , \new_[22723]_ , \new_[22724]_ ,
    \new_[22727]_ , \new_[22730]_ , \new_[22731]_ , \new_[22732]_ ,
    \new_[22736]_ , \new_[22737]_ , \new_[22740]_ , \new_[22743]_ ,
    \new_[22744]_ , \new_[22745]_ , \new_[22748]_ , \new_[22751]_ ,
    \new_[22752]_ , \new_[22755]_ , \new_[22758]_ , \new_[22759]_ ,
    \new_[22760]_ , \new_[22764]_ , \new_[22765]_ , \new_[22768]_ ,
    \new_[22771]_ , \new_[22772]_ , \new_[22773]_ , \new_[22776]_ ,
    \new_[22779]_ , \new_[22780]_ , \new_[22783]_ , \new_[22786]_ ,
    \new_[22787]_ , \new_[22788]_ , \new_[22792]_ , \new_[22793]_ ,
    \new_[22796]_ , \new_[22799]_ , \new_[22800]_ , \new_[22801]_ ,
    \new_[22804]_ , \new_[22807]_ , \new_[22808]_ , \new_[22811]_ ,
    \new_[22814]_ , \new_[22815]_ , \new_[22816]_ , \new_[22820]_ ,
    \new_[22821]_ , \new_[22824]_ , \new_[22827]_ , \new_[22828]_ ,
    \new_[22829]_ , \new_[22832]_ , \new_[22835]_ , \new_[22836]_ ,
    \new_[22839]_ , \new_[22842]_ , \new_[22843]_ , \new_[22844]_ ,
    \new_[22848]_ , \new_[22849]_ , \new_[22852]_ , \new_[22855]_ ,
    \new_[22856]_ , \new_[22857]_ , \new_[22860]_ , \new_[22863]_ ,
    \new_[22864]_ , \new_[22867]_ , \new_[22870]_ , \new_[22871]_ ,
    \new_[22872]_ , \new_[22876]_ , \new_[22877]_ , \new_[22880]_ ,
    \new_[22883]_ , \new_[22884]_ , \new_[22885]_ , \new_[22888]_ ,
    \new_[22891]_ , \new_[22892]_ , \new_[22895]_ , \new_[22898]_ ,
    \new_[22899]_ , \new_[22900]_ , \new_[22904]_ , \new_[22905]_ ,
    \new_[22908]_ , \new_[22911]_ , \new_[22912]_ , \new_[22913]_ ,
    \new_[22916]_ , \new_[22919]_ , \new_[22920]_ , \new_[22923]_ ,
    \new_[22926]_ , \new_[22927]_ , \new_[22928]_ , \new_[22932]_ ,
    \new_[22933]_ , \new_[22936]_ , \new_[22939]_ , \new_[22940]_ ,
    \new_[22941]_ , \new_[22944]_ , \new_[22947]_ , \new_[22948]_ ,
    \new_[22951]_ , \new_[22954]_ , \new_[22955]_ , \new_[22956]_ ,
    \new_[22960]_ , \new_[22961]_ , \new_[22964]_ , \new_[22967]_ ,
    \new_[22968]_ , \new_[22969]_ , \new_[22972]_ , \new_[22975]_ ,
    \new_[22976]_ , \new_[22979]_ , \new_[22982]_ , \new_[22983]_ ,
    \new_[22984]_ , \new_[22988]_ , \new_[22989]_ , \new_[22992]_ ,
    \new_[22995]_ , \new_[22996]_ , \new_[22997]_ , \new_[23000]_ ,
    \new_[23003]_ , \new_[23004]_ , \new_[23007]_ , \new_[23010]_ ,
    \new_[23011]_ , \new_[23012]_ , \new_[23016]_ , \new_[23017]_ ,
    \new_[23020]_ , \new_[23023]_ , \new_[23024]_ , \new_[23025]_ ,
    \new_[23028]_ , \new_[23031]_ , \new_[23032]_ , \new_[23035]_ ,
    \new_[23038]_ , \new_[23039]_ , \new_[23040]_ , \new_[23044]_ ,
    \new_[23045]_ , \new_[23048]_ , \new_[23051]_ , \new_[23052]_ ,
    \new_[23053]_ , \new_[23056]_ , \new_[23059]_ , \new_[23060]_ ,
    \new_[23063]_ , \new_[23066]_ , \new_[23067]_ , \new_[23068]_ ,
    \new_[23072]_ , \new_[23073]_ , \new_[23076]_ , \new_[23079]_ ,
    \new_[23080]_ , \new_[23081]_ , \new_[23084]_ , \new_[23087]_ ,
    \new_[23088]_ , \new_[23091]_ , \new_[23094]_ , \new_[23095]_ ,
    \new_[23096]_ , \new_[23100]_ , \new_[23101]_ , \new_[23104]_ ,
    \new_[23107]_ , \new_[23108]_ , \new_[23109]_ , \new_[23112]_ ,
    \new_[23115]_ , \new_[23116]_ , \new_[23119]_ , \new_[23122]_ ,
    \new_[23123]_ , \new_[23124]_ , \new_[23128]_ , \new_[23129]_ ,
    \new_[23132]_ , \new_[23135]_ , \new_[23136]_ , \new_[23137]_ ,
    \new_[23140]_ , \new_[23143]_ , \new_[23144]_ , \new_[23147]_ ,
    \new_[23150]_ , \new_[23151]_ , \new_[23152]_ , \new_[23156]_ ,
    \new_[23157]_ , \new_[23160]_ , \new_[23163]_ , \new_[23164]_ ,
    \new_[23165]_ , \new_[23168]_ , \new_[23171]_ , \new_[23172]_ ,
    \new_[23175]_ , \new_[23178]_ , \new_[23179]_ , \new_[23180]_ ,
    \new_[23184]_ , \new_[23185]_ , \new_[23188]_ , \new_[23191]_ ,
    \new_[23192]_ , \new_[23193]_ , \new_[23196]_ , \new_[23199]_ ,
    \new_[23200]_ , \new_[23203]_ , \new_[23206]_ , \new_[23207]_ ,
    \new_[23208]_ , \new_[23212]_ , \new_[23213]_ , \new_[23216]_ ,
    \new_[23219]_ , \new_[23220]_ , \new_[23221]_ , \new_[23224]_ ,
    \new_[23227]_ , \new_[23228]_ , \new_[23231]_ , \new_[23234]_ ,
    \new_[23235]_ , \new_[23236]_ , \new_[23240]_ , \new_[23241]_ ,
    \new_[23244]_ , \new_[23247]_ , \new_[23248]_ , \new_[23249]_ ,
    \new_[23252]_ , \new_[23255]_ , \new_[23256]_ , \new_[23259]_ ,
    \new_[23262]_ , \new_[23263]_ , \new_[23264]_ , \new_[23268]_ ,
    \new_[23269]_ , \new_[23272]_ , \new_[23275]_ , \new_[23276]_ ,
    \new_[23277]_ , \new_[23280]_ , \new_[23283]_ , \new_[23284]_ ,
    \new_[23287]_ , \new_[23290]_ , \new_[23291]_ , \new_[23292]_ ,
    \new_[23296]_ , \new_[23297]_ , \new_[23300]_ , \new_[23303]_ ,
    \new_[23304]_ , \new_[23305]_ , \new_[23308]_ , \new_[23311]_ ,
    \new_[23312]_ , \new_[23315]_ , \new_[23318]_ , \new_[23319]_ ,
    \new_[23320]_ , \new_[23324]_ , \new_[23325]_ , \new_[23328]_ ,
    \new_[23331]_ , \new_[23332]_ , \new_[23333]_ , \new_[23336]_ ,
    \new_[23339]_ , \new_[23340]_ , \new_[23343]_ , \new_[23346]_ ,
    \new_[23347]_ , \new_[23348]_ , \new_[23352]_ , \new_[23353]_ ,
    \new_[23356]_ , \new_[23359]_ , \new_[23360]_ , \new_[23361]_ ,
    \new_[23364]_ , \new_[23367]_ , \new_[23368]_ , \new_[23371]_ ,
    \new_[23374]_ , \new_[23375]_ , \new_[23376]_ , \new_[23380]_ ,
    \new_[23381]_ , \new_[23384]_ , \new_[23387]_ , \new_[23388]_ ,
    \new_[23389]_ , \new_[23392]_ , \new_[23395]_ , \new_[23396]_ ,
    \new_[23399]_ , \new_[23402]_ , \new_[23403]_ , \new_[23404]_ ,
    \new_[23408]_ , \new_[23409]_ , \new_[23412]_ , \new_[23415]_ ,
    \new_[23416]_ , \new_[23417]_ , \new_[23420]_ , \new_[23423]_ ,
    \new_[23424]_ , \new_[23427]_ , \new_[23430]_ , \new_[23431]_ ,
    \new_[23432]_ , \new_[23436]_ , \new_[23437]_ , \new_[23440]_ ,
    \new_[23443]_ , \new_[23444]_ , \new_[23445]_ , \new_[23448]_ ,
    \new_[23451]_ , \new_[23452]_ , \new_[23455]_ , \new_[23458]_ ,
    \new_[23459]_ , \new_[23460]_ , \new_[23464]_ , \new_[23465]_ ,
    \new_[23468]_ , \new_[23471]_ , \new_[23472]_ , \new_[23473]_ ,
    \new_[23476]_ , \new_[23479]_ , \new_[23480]_ , \new_[23483]_ ,
    \new_[23486]_ , \new_[23487]_ , \new_[23488]_ , \new_[23492]_ ,
    \new_[23493]_ , \new_[23496]_ , \new_[23499]_ , \new_[23500]_ ,
    \new_[23501]_ , \new_[23504]_ , \new_[23507]_ , \new_[23508]_ ,
    \new_[23511]_ , \new_[23514]_ , \new_[23515]_ , \new_[23516]_ ,
    \new_[23520]_ , \new_[23521]_ , \new_[23524]_ , \new_[23527]_ ,
    \new_[23528]_ , \new_[23529]_ , \new_[23532]_ , \new_[23535]_ ,
    \new_[23536]_ , \new_[23539]_ , \new_[23542]_ , \new_[23543]_ ,
    \new_[23544]_ , \new_[23548]_ , \new_[23549]_ , \new_[23552]_ ,
    \new_[23555]_ , \new_[23556]_ , \new_[23557]_ , \new_[23560]_ ,
    \new_[23563]_ , \new_[23564]_ , \new_[23567]_ , \new_[23570]_ ,
    \new_[23571]_ , \new_[23572]_ , \new_[23576]_ , \new_[23577]_ ,
    \new_[23580]_ , \new_[23583]_ , \new_[23584]_ , \new_[23585]_ ,
    \new_[23588]_ , \new_[23591]_ , \new_[23592]_ , \new_[23595]_ ,
    \new_[23598]_ , \new_[23599]_ , \new_[23600]_ , \new_[23604]_ ,
    \new_[23605]_ , \new_[23608]_ , \new_[23611]_ , \new_[23612]_ ,
    \new_[23613]_ , \new_[23616]_ , \new_[23619]_ , \new_[23620]_ ,
    \new_[23623]_ , \new_[23626]_ , \new_[23627]_ , \new_[23628]_ ,
    \new_[23632]_ , \new_[23633]_ , \new_[23636]_ , \new_[23639]_ ,
    \new_[23640]_ , \new_[23641]_ , \new_[23644]_ , \new_[23647]_ ,
    \new_[23648]_ , \new_[23651]_ , \new_[23654]_ , \new_[23655]_ ,
    \new_[23656]_ , \new_[23660]_ , \new_[23661]_ , \new_[23664]_ ,
    \new_[23667]_ , \new_[23668]_ , \new_[23669]_ , \new_[23672]_ ,
    \new_[23675]_ , \new_[23676]_ , \new_[23679]_ , \new_[23682]_ ,
    \new_[23683]_ , \new_[23684]_ , \new_[23688]_ , \new_[23689]_ ,
    \new_[23692]_ , \new_[23695]_ , \new_[23696]_ , \new_[23697]_ ,
    \new_[23700]_ , \new_[23703]_ , \new_[23704]_ , \new_[23707]_ ,
    \new_[23710]_ , \new_[23711]_ , \new_[23712]_ , \new_[23716]_ ,
    \new_[23717]_ , \new_[23720]_ , \new_[23723]_ , \new_[23724]_ ,
    \new_[23725]_ , \new_[23728]_ , \new_[23731]_ , \new_[23732]_ ,
    \new_[23735]_ , \new_[23738]_ , \new_[23739]_ , \new_[23740]_ ,
    \new_[23744]_ , \new_[23745]_ , \new_[23748]_ , \new_[23751]_ ,
    \new_[23752]_ , \new_[23753]_ , \new_[23756]_ , \new_[23759]_ ,
    \new_[23760]_ , \new_[23763]_ , \new_[23766]_ , \new_[23767]_ ,
    \new_[23768]_ , \new_[23772]_ , \new_[23773]_ , \new_[23776]_ ,
    \new_[23779]_ , \new_[23780]_ , \new_[23781]_ , \new_[23784]_ ,
    \new_[23787]_ , \new_[23788]_ , \new_[23791]_ , \new_[23794]_ ,
    \new_[23795]_ , \new_[23796]_ , \new_[23800]_ , \new_[23801]_ ,
    \new_[23804]_ , \new_[23807]_ , \new_[23808]_ , \new_[23809]_ ,
    \new_[23812]_ , \new_[23815]_ , \new_[23816]_ , \new_[23819]_ ,
    \new_[23822]_ , \new_[23823]_ , \new_[23824]_ , \new_[23828]_ ,
    \new_[23829]_ , \new_[23832]_ , \new_[23835]_ , \new_[23836]_ ,
    \new_[23837]_ , \new_[23840]_ , \new_[23843]_ , \new_[23844]_ ,
    \new_[23847]_ , \new_[23850]_ , \new_[23851]_ , \new_[23852]_ ,
    \new_[23856]_ , \new_[23857]_ , \new_[23860]_ , \new_[23863]_ ,
    \new_[23864]_ , \new_[23865]_ , \new_[23868]_ , \new_[23871]_ ,
    \new_[23872]_ , \new_[23875]_ , \new_[23878]_ , \new_[23879]_ ,
    \new_[23880]_ , \new_[23884]_ , \new_[23885]_ , \new_[23888]_ ,
    \new_[23891]_ , \new_[23892]_ , \new_[23893]_ , \new_[23896]_ ,
    \new_[23899]_ , \new_[23900]_ , \new_[23903]_ , \new_[23906]_ ,
    \new_[23907]_ , \new_[23908]_ , \new_[23912]_ , \new_[23913]_ ,
    \new_[23916]_ , \new_[23919]_ , \new_[23920]_ , \new_[23921]_ ,
    \new_[23924]_ , \new_[23927]_ , \new_[23928]_ , \new_[23931]_ ,
    \new_[23934]_ , \new_[23935]_ , \new_[23936]_ , \new_[23940]_ ,
    \new_[23941]_ , \new_[23944]_ , \new_[23947]_ , \new_[23948]_ ,
    \new_[23949]_ , \new_[23952]_ , \new_[23955]_ , \new_[23956]_ ,
    \new_[23959]_ , \new_[23962]_ , \new_[23963]_ , \new_[23964]_ ,
    \new_[23968]_ , \new_[23969]_ , \new_[23972]_ , \new_[23975]_ ,
    \new_[23976]_ , \new_[23977]_ , \new_[23980]_ , \new_[23983]_ ,
    \new_[23984]_ , \new_[23987]_ , \new_[23990]_ , \new_[23991]_ ,
    \new_[23992]_ , \new_[23996]_ , \new_[23997]_ , \new_[24000]_ ,
    \new_[24003]_ , \new_[24004]_ , \new_[24005]_ , \new_[24008]_ ,
    \new_[24011]_ , \new_[24012]_ , \new_[24015]_ , \new_[24018]_ ,
    \new_[24019]_ , \new_[24020]_ , \new_[24024]_ , \new_[24025]_ ,
    \new_[24028]_ , \new_[24031]_ , \new_[24032]_ , \new_[24033]_ ,
    \new_[24036]_ , \new_[24039]_ , \new_[24040]_ , \new_[24043]_ ,
    \new_[24046]_ , \new_[24047]_ , \new_[24048]_ , \new_[24052]_ ,
    \new_[24053]_ , \new_[24056]_ , \new_[24059]_ , \new_[24060]_ ,
    \new_[24061]_ , \new_[24064]_ , \new_[24067]_ , \new_[24068]_ ,
    \new_[24071]_ , \new_[24074]_ , \new_[24075]_ , \new_[24076]_ ,
    \new_[24080]_ , \new_[24081]_ , \new_[24084]_ , \new_[24087]_ ,
    \new_[24088]_ , \new_[24089]_ , \new_[24092]_ , \new_[24095]_ ,
    \new_[24096]_ , \new_[24099]_ , \new_[24102]_ , \new_[24103]_ ,
    \new_[24104]_ , \new_[24108]_ , \new_[24109]_ , \new_[24112]_ ,
    \new_[24115]_ , \new_[24116]_ , \new_[24117]_ , \new_[24120]_ ,
    \new_[24123]_ , \new_[24124]_ , \new_[24127]_ , \new_[24130]_ ,
    \new_[24131]_ , \new_[24132]_ , \new_[24136]_ , \new_[24137]_ ,
    \new_[24140]_ , \new_[24143]_ , \new_[24144]_ , \new_[24145]_ ,
    \new_[24148]_ , \new_[24151]_ , \new_[24152]_ , \new_[24155]_ ,
    \new_[24158]_ , \new_[24159]_ , \new_[24160]_ , \new_[24164]_ ,
    \new_[24165]_ , \new_[24168]_ , \new_[24171]_ , \new_[24172]_ ,
    \new_[24173]_ , \new_[24176]_ , \new_[24179]_ , \new_[24180]_ ,
    \new_[24183]_ , \new_[24186]_ , \new_[24187]_ , \new_[24188]_ ,
    \new_[24192]_ , \new_[24193]_ , \new_[24196]_ , \new_[24199]_ ,
    \new_[24200]_ , \new_[24201]_ , \new_[24204]_ , \new_[24207]_ ,
    \new_[24208]_ , \new_[24211]_ , \new_[24214]_ , \new_[24215]_ ,
    \new_[24216]_ , \new_[24220]_ , \new_[24221]_ , \new_[24224]_ ,
    \new_[24227]_ , \new_[24228]_ , \new_[24229]_ , \new_[24232]_ ,
    \new_[24235]_ , \new_[24236]_ , \new_[24239]_ , \new_[24242]_ ,
    \new_[24243]_ , \new_[24244]_ , \new_[24248]_ , \new_[24249]_ ,
    \new_[24252]_ , \new_[24255]_ , \new_[24256]_ , \new_[24257]_ ,
    \new_[24260]_ , \new_[24263]_ , \new_[24264]_ , \new_[24267]_ ,
    \new_[24270]_ , \new_[24271]_ , \new_[24272]_ , \new_[24276]_ ,
    \new_[24277]_ , \new_[24280]_ , \new_[24283]_ , \new_[24284]_ ,
    \new_[24285]_ , \new_[24288]_ , \new_[24291]_ , \new_[24292]_ ,
    \new_[24295]_ , \new_[24298]_ , \new_[24299]_ , \new_[24300]_ ,
    \new_[24304]_ , \new_[24305]_ , \new_[24308]_ , \new_[24311]_ ,
    \new_[24312]_ , \new_[24313]_ , \new_[24316]_ , \new_[24319]_ ,
    \new_[24320]_ , \new_[24323]_ , \new_[24326]_ , \new_[24327]_ ,
    \new_[24328]_ , \new_[24332]_ , \new_[24333]_ , \new_[24336]_ ,
    \new_[24339]_ , \new_[24340]_ , \new_[24341]_ , \new_[24344]_ ,
    \new_[24347]_ , \new_[24348]_ , \new_[24351]_ , \new_[24354]_ ,
    \new_[24355]_ , \new_[24356]_ , \new_[24360]_ , \new_[24361]_ ,
    \new_[24364]_ , \new_[24367]_ , \new_[24368]_ , \new_[24369]_ ,
    \new_[24372]_ , \new_[24375]_ , \new_[24376]_ , \new_[24379]_ ,
    \new_[24382]_ , \new_[24383]_ , \new_[24384]_ , \new_[24388]_ ,
    \new_[24389]_ , \new_[24392]_ , \new_[24395]_ , \new_[24396]_ ,
    \new_[24397]_ , \new_[24400]_ , \new_[24403]_ , \new_[24404]_ ,
    \new_[24407]_ , \new_[24410]_ , \new_[24411]_ , \new_[24412]_ ,
    \new_[24416]_ , \new_[24417]_ , \new_[24420]_ , \new_[24423]_ ,
    \new_[24424]_ , \new_[24425]_ , \new_[24428]_ , \new_[24431]_ ,
    \new_[24432]_ , \new_[24435]_ , \new_[24438]_ , \new_[24439]_ ,
    \new_[24440]_ , \new_[24444]_ , \new_[24445]_ , \new_[24448]_ ,
    \new_[24451]_ , \new_[24452]_ , \new_[24453]_ , \new_[24456]_ ,
    \new_[24459]_ , \new_[24460]_ , \new_[24463]_ , \new_[24466]_ ,
    \new_[24467]_ , \new_[24468]_ , \new_[24472]_ , \new_[24473]_ ,
    \new_[24476]_ , \new_[24479]_ , \new_[24480]_ , \new_[24481]_ ,
    \new_[24484]_ , \new_[24487]_ , \new_[24488]_ , \new_[24491]_ ,
    \new_[24494]_ , \new_[24495]_ , \new_[24496]_ , \new_[24500]_ ,
    \new_[24501]_ , \new_[24504]_ , \new_[24507]_ , \new_[24508]_ ,
    \new_[24509]_ , \new_[24512]_ , \new_[24515]_ , \new_[24516]_ ,
    \new_[24519]_ , \new_[24522]_ , \new_[24523]_ , \new_[24524]_ ,
    \new_[24528]_ , \new_[24529]_ , \new_[24532]_ , \new_[24535]_ ,
    \new_[24536]_ , \new_[24537]_ , \new_[24540]_ , \new_[24543]_ ,
    \new_[24544]_ , \new_[24547]_ , \new_[24550]_ , \new_[24551]_ ,
    \new_[24552]_ , \new_[24556]_ , \new_[24557]_ , \new_[24560]_ ,
    \new_[24563]_ , \new_[24564]_ , \new_[24565]_ , \new_[24568]_ ,
    \new_[24571]_ , \new_[24572]_ , \new_[24575]_ , \new_[24578]_ ,
    \new_[24579]_ , \new_[24580]_ , \new_[24584]_ , \new_[24585]_ ,
    \new_[24588]_ , \new_[24591]_ , \new_[24592]_ , \new_[24593]_ ,
    \new_[24596]_ , \new_[24599]_ , \new_[24600]_ , \new_[24603]_ ,
    \new_[24606]_ , \new_[24607]_ , \new_[24608]_ , \new_[24612]_ ,
    \new_[24613]_ , \new_[24616]_ , \new_[24619]_ , \new_[24620]_ ,
    \new_[24621]_ , \new_[24624]_ , \new_[24627]_ , \new_[24628]_ ,
    \new_[24631]_ , \new_[24634]_ , \new_[24635]_ , \new_[24636]_ ,
    \new_[24640]_ , \new_[24641]_ , \new_[24644]_ , \new_[24647]_ ,
    \new_[24648]_ , \new_[24649]_ , \new_[24652]_ , \new_[24655]_ ,
    \new_[24656]_ , \new_[24659]_ , \new_[24662]_ , \new_[24663]_ ,
    \new_[24664]_ , \new_[24668]_ , \new_[24669]_ , \new_[24672]_ ,
    \new_[24675]_ , \new_[24676]_ , \new_[24677]_ , \new_[24680]_ ,
    \new_[24683]_ , \new_[24684]_ , \new_[24687]_ , \new_[24690]_ ,
    \new_[24691]_ , \new_[24692]_ , \new_[24696]_ , \new_[24697]_ ,
    \new_[24700]_ , \new_[24703]_ , \new_[24704]_ , \new_[24705]_ ,
    \new_[24708]_ , \new_[24711]_ , \new_[24712]_ , \new_[24715]_ ,
    \new_[24718]_ , \new_[24719]_ , \new_[24720]_ , \new_[24724]_ ,
    \new_[24725]_ , \new_[24728]_ , \new_[24731]_ , \new_[24732]_ ,
    \new_[24733]_ , \new_[24736]_ , \new_[24739]_ , \new_[24740]_ ,
    \new_[24743]_ , \new_[24746]_ , \new_[24747]_ , \new_[24748]_ ,
    \new_[24752]_ , \new_[24753]_ , \new_[24756]_ , \new_[24759]_ ,
    \new_[24760]_ , \new_[24761]_ , \new_[24764]_ , \new_[24767]_ ,
    \new_[24768]_ , \new_[24771]_ , \new_[24774]_ , \new_[24775]_ ,
    \new_[24776]_ , \new_[24780]_ , \new_[24781]_ , \new_[24784]_ ,
    \new_[24787]_ , \new_[24788]_ , \new_[24789]_ , \new_[24792]_ ,
    \new_[24795]_ , \new_[24796]_ , \new_[24799]_ , \new_[24802]_ ,
    \new_[24803]_ , \new_[24804]_ , \new_[24808]_ , \new_[24809]_ ,
    \new_[24812]_ , \new_[24815]_ , \new_[24816]_ , \new_[24817]_ ,
    \new_[24820]_ , \new_[24823]_ , \new_[24824]_ , \new_[24827]_ ,
    \new_[24830]_ , \new_[24831]_ , \new_[24832]_ , \new_[24836]_ ,
    \new_[24837]_ , \new_[24840]_ , \new_[24843]_ , \new_[24844]_ ,
    \new_[24845]_ , \new_[24848]_ , \new_[24851]_ , \new_[24852]_ ,
    \new_[24855]_ , \new_[24858]_ , \new_[24859]_ , \new_[24860]_ ,
    \new_[24864]_ , \new_[24865]_ , \new_[24868]_ , \new_[24871]_ ,
    \new_[24872]_ , \new_[24873]_ , \new_[24876]_ , \new_[24879]_ ,
    \new_[24880]_ , \new_[24883]_ , \new_[24886]_ , \new_[24887]_ ,
    \new_[24888]_ , \new_[24892]_ , \new_[24893]_ , \new_[24896]_ ,
    \new_[24899]_ , \new_[24900]_ , \new_[24901]_ , \new_[24904]_ ,
    \new_[24907]_ , \new_[24908]_ , \new_[24911]_ , \new_[24914]_ ,
    \new_[24915]_ , \new_[24916]_ , \new_[24920]_ , \new_[24921]_ ,
    \new_[24924]_ , \new_[24927]_ , \new_[24928]_ , \new_[24929]_ ,
    \new_[24932]_ , \new_[24935]_ , \new_[24936]_ , \new_[24939]_ ,
    \new_[24942]_ , \new_[24943]_ , \new_[24944]_ , \new_[24948]_ ,
    \new_[24949]_ , \new_[24952]_ , \new_[24955]_ , \new_[24956]_ ,
    \new_[24957]_ , \new_[24960]_ , \new_[24963]_ , \new_[24964]_ ,
    \new_[24967]_ , \new_[24970]_ , \new_[24971]_ , \new_[24972]_ ,
    \new_[24976]_ , \new_[24977]_ , \new_[24980]_ , \new_[24983]_ ,
    \new_[24984]_ , \new_[24985]_ , \new_[24988]_ , \new_[24991]_ ,
    \new_[24992]_ , \new_[24995]_ , \new_[24998]_ , \new_[24999]_ ,
    \new_[25000]_ , \new_[25004]_ , \new_[25005]_ , \new_[25008]_ ,
    \new_[25011]_ , \new_[25012]_ , \new_[25013]_ , \new_[25016]_ ,
    \new_[25019]_ , \new_[25020]_ , \new_[25023]_ , \new_[25026]_ ,
    \new_[25027]_ , \new_[25028]_ , \new_[25032]_ , \new_[25033]_ ,
    \new_[25036]_ , \new_[25039]_ , \new_[25040]_ , \new_[25041]_ ,
    \new_[25044]_ , \new_[25047]_ , \new_[25048]_ , \new_[25051]_ ,
    \new_[25054]_ , \new_[25055]_ , \new_[25056]_ , \new_[25060]_ ,
    \new_[25061]_ , \new_[25064]_ , \new_[25067]_ , \new_[25068]_ ,
    \new_[25069]_ , \new_[25072]_ , \new_[25075]_ , \new_[25076]_ ,
    \new_[25079]_ , \new_[25082]_ , \new_[25083]_ , \new_[25084]_ ,
    \new_[25088]_ , \new_[25089]_ , \new_[25092]_ , \new_[25095]_ ,
    \new_[25096]_ , \new_[25097]_ , \new_[25100]_ , \new_[25103]_ ,
    \new_[25104]_ , \new_[25107]_ , \new_[25110]_ , \new_[25111]_ ,
    \new_[25112]_ , \new_[25116]_ , \new_[25117]_ , \new_[25120]_ ,
    \new_[25123]_ , \new_[25124]_ , \new_[25125]_ , \new_[25128]_ ,
    \new_[25131]_ , \new_[25132]_ , \new_[25135]_ , \new_[25138]_ ,
    \new_[25139]_ , \new_[25140]_ , \new_[25144]_ , \new_[25145]_ ,
    \new_[25148]_ , \new_[25151]_ , \new_[25152]_ , \new_[25153]_ ,
    \new_[25156]_ , \new_[25159]_ , \new_[25160]_ , \new_[25163]_ ,
    \new_[25166]_ , \new_[25167]_ , \new_[25168]_ , \new_[25172]_ ,
    \new_[25173]_ , \new_[25176]_ , \new_[25179]_ , \new_[25180]_ ,
    \new_[25181]_ , \new_[25184]_ , \new_[25187]_ , \new_[25188]_ ,
    \new_[25191]_ , \new_[25194]_ , \new_[25195]_ , \new_[25196]_ ,
    \new_[25200]_ , \new_[25201]_ , \new_[25204]_ , \new_[25207]_ ,
    \new_[25208]_ , \new_[25209]_ , \new_[25212]_ , \new_[25215]_ ,
    \new_[25216]_ , \new_[25219]_ , \new_[25222]_ , \new_[25223]_ ,
    \new_[25224]_ , \new_[25228]_ , \new_[25229]_ , \new_[25232]_ ,
    \new_[25235]_ , \new_[25236]_ , \new_[25237]_ , \new_[25240]_ ,
    \new_[25243]_ , \new_[25244]_ , \new_[25247]_ , \new_[25250]_ ,
    \new_[25251]_ , \new_[25252]_ , \new_[25256]_ , \new_[25257]_ ,
    \new_[25260]_ , \new_[25263]_ , \new_[25264]_ , \new_[25265]_ ,
    \new_[25268]_ , \new_[25271]_ , \new_[25272]_ , \new_[25275]_ ,
    \new_[25278]_ , \new_[25279]_ , \new_[25280]_ , \new_[25284]_ ,
    \new_[25285]_ , \new_[25288]_ , \new_[25291]_ , \new_[25292]_ ,
    \new_[25293]_ , \new_[25296]_ , \new_[25299]_ , \new_[25300]_ ,
    \new_[25303]_ , \new_[25306]_ , \new_[25307]_ , \new_[25308]_ ,
    \new_[25312]_ , \new_[25313]_ , \new_[25316]_ , \new_[25319]_ ,
    \new_[25320]_ , \new_[25321]_ , \new_[25324]_ , \new_[25327]_ ,
    \new_[25328]_ , \new_[25331]_ , \new_[25334]_ , \new_[25335]_ ,
    \new_[25336]_ , \new_[25340]_ , \new_[25341]_ , \new_[25344]_ ,
    \new_[25347]_ , \new_[25348]_ , \new_[25349]_ , \new_[25352]_ ,
    \new_[25355]_ , \new_[25356]_ , \new_[25359]_ , \new_[25362]_ ,
    \new_[25363]_ , \new_[25364]_ , \new_[25368]_ , \new_[25369]_ ,
    \new_[25372]_ , \new_[25375]_ , \new_[25376]_ , \new_[25377]_ ,
    \new_[25380]_ , \new_[25383]_ , \new_[25384]_ , \new_[25387]_ ,
    \new_[25390]_ , \new_[25391]_ , \new_[25392]_ , \new_[25396]_ ,
    \new_[25397]_ , \new_[25400]_ , \new_[25403]_ , \new_[25404]_ ,
    \new_[25405]_ , \new_[25408]_ , \new_[25411]_ , \new_[25412]_ ,
    \new_[25415]_ , \new_[25418]_ , \new_[25419]_ , \new_[25420]_ ,
    \new_[25424]_ , \new_[25425]_ , \new_[25428]_ , \new_[25431]_ ,
    \new_[25432]_ , \new_[25433]_ , \new_[25436]_ , \new_[25439]_ ,
    \new_[25440]_ , \new_[25443]_ , \new_[25446]_ , \new_[25447]_ ,
    \new_[25448]_ , \new_[25452]_ , \new_[25453]_ , \new_[25456]_ ,
    \new_[25459]_ , \new_[25460]_ , \new_[25461]_ , \new_[25464]_ ,
    \new_[25467]_ , \new_[25468]_ , \new_[25471]_ , \new_[25474]_ ,
    \new_[25475]_ , \new_[25476]_ , \new_[25480]_ , \new_[25481]_ ,
    \new_[25484]_ , \new_[25487]_ , \new_[25488]_ , \new_[25489]_ ,
    \new_[25492]_ , \new_[25495]_ , \new_[25496]_ , \new_[25499]_ ,
    \new_[25502]_ , \new_[25503]_ , \new_[25504]_ , \new_[25508]_ ,
    \new_[25509]_ , \new_[25512]_ , \new_[25515]_ , \new_[25516]_ ,
    \new_[25517]_ , \new_[25520]_ , \new_[25523]_ , \new_[25524]_ ,
    \new_[25527]_ , \new_[25530]_ , \new_[25531]_ , \new_[25532]_ ,
    \new_[25536]_ , \new_[25537]_ , \new_[25540]_ , \new_[25543]_ ,
    \new_[25544]_ , \new_[25545]_ , \new_[25548]_ , \new_[25551]_ ,
    \new_[25552]_ , \new_[25555]_ , \new_[25558]_ , \new_[25559]_ ,
    \new_[25560]_ , \new_[25564]_ , \new_[25565]_ , \new_[25568]_ ,
    \new_[25571]_ , \new_[25572]_ , \new_[25573]_ , \new_[25576]_ ,
    \new_[25579]_ , \new_[25580]_ , \new_[25583]_ , \new_[25586]_ ,
    \new_[25587]_ , \new_[25588]_ , \new_[25592]_ , \new_[25593]_ ,
    \new_[25596]_ , \new_[25599]_ , \new_[25600]_ , \new_[25601]_ ,
    \new_[25604]_ , \new_[25607]_ , \new_[25608]_ , \new_[25611]_ ,
    \new_[25614]_ , \new_[25615]_ , \new_[25616]_ , \new_[25620]_ ,
    \new_[25621]_ , \new_[25624]_ , \new_[25627]_ , \new_[25628]_ ,
    \new_[25629]_ , \new_[25632]_ , \new_[25635]_ , \new_[25636]_ ,
    \new_[25639]_ , \new_[25642]_ , \new_[25643]_ , \new_[25644]_ ,
    \new_[25648]_ , \new_[25649]_ , \new_[25652]_ , \new_[25655]_ ,
    \new_[25656]_ , \new_[25657]_ , \new_[25660]_ , \new_[25663]_ ,
    \new_[25664]_ , \new_[25667]_ , \new_[25670]_ , \new_[25671]_ ,
    \new_[25672]_ , \new_[25676]_ , \new_[25677]_ , \new_[25680]_ ,
    \new_[25683]_ , \new_[25684]_ , \new_[25685]_ , \new_[25688]_ ,
    \new_[25691]_ , \new_[25692]_ , \new_[25695]_ , \new_[25698]_ ,
    \new_[25699]_ , \new_[25700]_ , \new_[25704]_ , \new_[25705]_ ,
    \new_[25708]_ , \new_[25711]_ , \new_[25712]_ , \new_[25713]_ ,
    \new_[25716]_ , \new_[25719]_ , \new_[25720]_ , \new_[25723]_ ,
    \new_[25726]_ , \new_[25727]_ , \new_[25728]_ , \new_[25732]_ ,
    \new_[25733]_ , \new_[25736]_ , \new_[25739]_ , \new_[25740]_ ,
    \new_[25741]_ , \new_[25744]_ , \new_[25747]_ , \new_[25748]_ ,
    \new_[25751]_ , \new_[25754]_ , \new_[25755]_ , \new_[25756]_ ,
    \new_[25760]_ , \new_[25761]_ , \new_[25764]_ , \new_[25767]_ ,
    \new_[25768]_ , \new_[25769]_ , \new_[25772]_ , \new_[25775]_ ,
    \new_[25776]_ , \new_[25779]_ , \new_[25782]_ , \new_[25783]_ ,
    \new_[25784]_ , \new_[25788]_ , \new_[25789]_ , \new_[25792]_ ,
    \new_[25795]_ , \new_[25796]_ , \new_[25797]_ , \new_[25800]_ ,
    \new_[25803]_ , \new_[25804]_ , \new_[25807]_ , \new_[25810]_ ,
    \new_[25811]_ , \new_[25812]_ , \new_[25816]_ , \new_[25817]_ ,
    \new_[25820]_ , \new_[25823]_ , \new_[25824]_ , \new_[25825]_ ,
    \new_[25828]_ , \new_[25831]_ , \new_[25832]_ , \new_[25835]_ ,
    \new_[25838]_ , \new_[25839]_ , \new_[25840]_ , \new_[25844]_ ,
    \new_[25845]_ , \new_[25848]_ , \new_[25851]_ , \new_[25852]_ ,
    \new_[25853]_ , \new_[25856]_ , \new_[25859]_ , \new_[25860]_ ,
    \new_[25863]_ , \new_[25866]_ , \new_[25867]_ , \new_[25868]_ ,
    \new_[25872]_ , \new_[25873]_ , \new_[25876]_ , \new_[25879]_ ,
    \new_[25880]_ , \new_[25881]_ , \new_[25884]_ , \new_[25887]_ ,
    \new_[25888]_ , \new_[25891]_ , \new_[25894]_ , \new_[25895]_ ,
    \new_[25896]_ , \new_[25900]_ , \new_[25901]_ , \new_[25904]_ ,
    \new_[25907]_ , \new_[25908]_ , \new_[25909]_ , \new_[25912]_ ,
    \new_[25915]_ , \new_[25916]_ , \new_[25919]_ , \new_[25922]_ ,
    \new_[25923]_ , \new_[25924]_ , \new_[25928]_ , \new_[25929]_ ,
    \new_[25932]_ , \new_[25935]_ , \new_[25936]_ , \new_[25937]_ ,
    \new_[25940]_ , \new_[25943]_ , \new_[25944]_ , \new_[25947]_ ,
    \new_[25950]_ , \new_[25951]_ , \new_[25952]_ , \new_[25956]_ ,
    \new_[25957]_ , \new_[25960]_ , \new_[25963]_ , \new_[25964]_ ,
    \new_[25965]_ , \new_[25968]_ , \new_[25971]_ , \new_[25972]_ ,
    \new_[25975]_ , \new_[25978]_ , \new_[25979]_ , \new_[25980]_ ,
    \new_[25984]_ , \new_[25985]_ , \new_[25988]_ , \new_[25991]_ ,
    \new_[25992]_ , \new_[25993]_ , \new_[25996]_ , \new_[25999]_ ,
    \new_[26000]_ , \new_[26003]_ , \new_[26006]_ , \new_[26007]_ ,
    \new_[26008]_ , \new_[26012]_ , \new_[26013]_ , \new_[26016]_ ,
    \new_[26019]_ , \new_[26020]_ , \new_[26021]_ , \new_[26024]_ ,
    \new_[26027]_ , \new_[26028]_ , \new_[26031]_ , \new_[26034]_ ,
    \new_[26035]_ , \new_[26036]_ , \new_[26040]_ , \new_[26041]_ ,
    \new_[26044]_ , \new_[26047]_ , \new_[26048]_ , \new_[26049]_ ,
    \new_[26052]_ , \new_[26055]_ , \new_[26056]_ , \new_[26059]_ ,
    \new_[26062]_ , \new_[26063]_ , \new_[26064]_ , \new_[26068]_ ,
    \new_[26069]_ , \new_[26072]_ , \new_[26075]_ , \new_[26076]_ ,
    \new_[26077]_ , \new_[26080]_ , \new_[26083]_ , \new_[26084]_ ,
    \new_[26087]_ , \new_[26090]_ , \new_[26091]_ , \new_[26092]_ ,
    \new_[26096]_ , \new_[26097]_ , \new_[26100]_ , \new_[26103]_ ,
    \new_[26104]_ , \new_[26105]_ , \new_[26108]_ , \new_[26111]_ ,
    \new_[26112]_ , \new_[26115]_ , \new_[26118]_ , \new_[26119]_ ,
    \new_[26120]_ , \new_[26124]_ , \new_[26125]_ , \new_[26128]_ ,
    \new_[26131]_ , \new_[26132]_ , \new_[26133]_ , \new_[26136]_ ,
    \new_[26139]_ , \new_[26140]_ , \new_[26143]_ , \new_[26146]_ ,
    \new_[26147]_ , \new_[26148]_ , \new_[26152]_ , \new_[26153]_ ,
    \new_[26156]_ , \new_[26159]_ , \new_[26160]_ , \new_[26161]_ ,
    \new_[26164]_ , \new_[26167]_ , \new_[26168]_ , \new_[26171]_ ,
    \new_[26174]_ , \new_[26175]_ , \new_[26176]_ , \new_[26180]_ ,
    \new_[26181]_ , \new_[26184]_ , \new_[26187]_ , \new_[26188]_ ,
    \new_[26189]_ , \new_[26192]_ , \new_[26195]_ , \new_[26196]_ ,
    \new_[26199]_ , \new_[26202]_ , \new_[26203]_ , \new_[26204]_ ,
    \new_[26208]_ , \new_[26209]_ , \new_[26212]_ , \new_[26215]_ ,
    \new_[26216]_ , \new_[26217]_ , \new_[26220]_ , \new_[26223]_ ,
    \new_[26224]_ , \new_[26227]_ , \new_[26230]_ , \new_[26231]_ ,
    \new_[26232]_ , \new_[26236]_ , \new_[26237]_ , \new_[26240]_ ,
    \new_[26243]_ , \new_[26244]_ , \new_[26245]_ , \new_[26248]_ ,
    \new_[26251]_ , \new_[26252]_ , \new_[26255]_ , \new_[26258]_ ,
    \new_[26259]_ , \new_[26260]_ , \new_[26264]_ , \new_[26265]_ ,
    \new_[26268]_ , \new_[26271]_ , \new_[26272]_ , \new_[26273]_ ,
    \new_[26276]_ , \new_[26279]_ , \new_[26280]_ , \new_[26283]_ ,
    \new_[26286]_ , \new_[26287]_ , \new_[26288]_ , \new_[26292]_ ,
    \new_[26293]_ , \new_[26296]_ , \new_[26299]_ , \new_[26300]_ ,
    \new_[26301]_ , \new_[26304]_ , \new_[26307]_ , \new_[26308]_ ,
    \new_[26311]_ , \new_[26314]_ , \new_[26315]_ , \new_[26316]_ ,
    \new_[26320]_ , \new_[26321]_ , \new_[26324]_ , \new_[26327]_ ,
    \new_[26328]_ , \new_[26329]_ , \new_[26332]_ , \new_[26335]_ ,
    \new_[26336]_ , \new_[26339]_ , \new_[26342]_ , \new_[26343]_ ,
    \new_[26344]_ , \new_[26348]_ , \new_[26349]_ , \new_[26352]_ ,
    \new_[26355]_ , \new_[26356]_ , \new_[26357]_ , \new_[26360]_ ,
    \new_[26363]_ , \new_[26364]_ , \new_[26367]_ , \new_[26370]_ ,
    \new_[26371]_ , \new_[26372]_ , \new_[26376]_ , \new_[26377]_ ,
    \new_[26380]_ , \new_[26383]_ , \new_[26384]_ , \new_[26385]_ ,
    \new_[26388]_ , \new_[26391]_ , \new_[26392]_ , \new_[26395]_ ,
    \new_[26398]_ , \new_[26399]_ , \new_[26400]_ , \new_[26404]_ ,
    \new_[26405]_ , \new_[26408]_ , \new_[26411]_ , \new_[26412]_ ,
    \new_[26413]_ , \new_[26416]_ , \new_[26419]_ , \new_[26420]_ ,
    \new_[26423]_ , \new_[26426]_ , \new_[26427]_ , \new_[26428]_ ,
    \new_[26432]_ , \new_[26433]_ , \new_[26436]_ , \new_[26439]_ ,
    \new_[26440]_ , \new_[26441]_ , \new_[26444]_ , \new_[26447]_ ,
    \new_[26448]_ , \new_[26451]_ , \new_[26454]_ , \new_[26455]_ ,
    \new_[26456]_ , \new_[26460]_ , \new_[26461]_ , \new_[26464]_ ,
    \new_[26467]_ , \new_[26468]_ , \new_[26469]_ , \new_[26472]_ ,
    \new_[26475]_ , \new_[26476]_ , \new_[26479]_ , \new_[26482]_ ,
    \new_[26483]_ , \new_[26484]_ , \new_[26488]_ , \new_[26489]_ ,
    \new_[26492]_ , \new_[26495]_ , \new_[26496]_ , \new_[26497]_ ,
    \new_[26500]_ , \new_[26503]_ , \new_[26504]_ , \new_[26507]_ ,
    \new_[26510]_ , \new_[26511]_ , \new_[26512]_ , \new_[26516]_ ,
    \new_[26517]_ , \new_[26520]_ , \new_[26523]_ , \new_[26524]_ ,
    \new_[26525]_ , \new_[26528]_ , \new_[26531]_ , \new_[26532]_ ,
    \new_[26535]_ , \new_[26538]_ , \new_[26539]_ , \new_[26540]_ ,
    \new_[26544]_ , \new_[26545]_ , \new_[26548]_ , \new_[26551]_ ,
    \new_[26552]_ , \new_[26553]_ , \new_[26556]_ , \new_[26559]_ ,
    \new_[26560]_ , \new_[26563]_ , \new_[26566]_ , \new_[26567]_ ,
    \new_[26568]_ , \new_[26572]_ , \new_[26573]_ , \new_[26576]_ ,
    \new_[26579]_ , \new_[26580]_ , \new_[26581]_ , \new_[26584]_ ,
    \new_[26587]_ , \new_[26588]_ , \new_[26591]_ , \new_[26594]_ ,
    \new_[26595]_ , \new_[26596]_ , \new_[26600]_ , \new_[26601]_ ,
    \new_[26604]_ , \new_[26607]_ , \new_[26608]_ , \new_[26609]_ ,
    \new_[26612]_ , \new_[26615]_ , \new_[26616]_ , \new_[26619]_ ,
    \new_[26622]_ , \new_[26623]_ , \new_[26624]_ , \new_[26628]_ ,
    \new_[26629]_ , \new_[26632]_ , \new_[26635]_ , \new_[26636]_ ,
    \new_[26637]_ , \new_[26640]_ , \new_[26643]_ , \new_[26644]_ ,
    \new_[26647]_ , \new_[26650]_ , \new_[26651]_ , \new_[26652]_ ,
    \new_[26656]_ , \new_[26657]_ , \new_[26660]_ , \new_[26663]_ ,
    \new_[26664]_ , \new_[26665]_ , \new_[26668]_ , \new_[26671]_ ,
    \new_[26672]_ , \new_[26675]_ , \new_[26678]_ , \new_[26679]_ ,
    \new_[26680]_ , \new_[26684]_ , \new_[26685]_ , \new_[26688]_ ,
    \new_[26691]_ , \new_[26692]_ , \new_[26693]_ , \new_[26696]_ ,
    \new_[26699]_ , \new_[26700]_ , \new_[26703]_ , \new_[26706]_ ,
    \new_[26707]_ , \new_[26708]_ , \new_[26712]_ , \new_[26713]_ ,
    \new_[26716]_ , \new_[26719]_ , \new_[26720]_ , \new_[26721]_ ,
    \new_[26724]_ , \new_[26727]_ , \new_[26728]_ , \new_[26731]_ ,
    \new_[26734]_ , \new_[26735]_ , \new_[26736]_ , \new_[26740]_ ,
    \new_[26741]_ , \new_[26744]_ , \new_[26747]_ , \new_[26748]_ ,
    \new_[26749]_ , \new_[26752]_ , \new_[26755]_ , \new_[26756]_ ,
    \new_[26759]_ , \new_[26762]_ , \new_[26763]_ , \new_[26764]_ ,
    \new_[26768]_ , \new_[26769]_ , \new_[26772]_ , \new_[26775]_ ,
    \new_[26776]_ , \new_[26777]_ , \new_[26780]_ , \new_[26783]_ ,
    \new_[26784]_ , \new_[26787]_ , \new_[26790]_ , \new_[26791]_ ,
    \new_[26792]_ , \new_[26796]_ , \new_[26797]_ , \new_[26800]_ ,
    \new_[26803]_ , \new_[26804]_ , \new_[26805]_ , \new_[26808]_ ,
    \new_[26811]_ , \new_[26812]_ , \new_[26815]_ , \new_[26818]_ ,
    \new_[26819]_ , \new_[26820]_ , \new_[26824]_ , \new_[26825]_ ,
    \new_[26828]_ , \new_[26831]_ , \new_[26832]_ , \new_[26833]_ ,
    \new_[26836]_ , \new_[26839]_ , \new_[26840]_ , \new_[26843]_ ,
    \new_[26846]_ , \new_[26847]_ , \new_[26848]_ , \new_[26852]_ ,
    \new_[26853]_ , \new_[26856]_ , \new_[26859]_ , \new_[26860]_ ,
    \new_[26861]_ , \new_[26864]_ , \new_[26867]_ , \new_[26868]_ ,
    \new_[26871]_ , \new_[26874]_ , \new_[26875]_ , \new_[26876]_ ,
    \new_[26880]_ , \new_[26881]_ , \new_[26884]_ , \new_[26887]_ ,
    \new_[26888]_ , \new_[26889]_ , \new_[26892]_ , \new_[26895]_ ,
    \new_[26896]_ , \new_[26899]_ , \new_[26902]_ , \new_[26903]_ ,
    \new_[26904]_ , \new_[26908]_ , \new_[26909]_ , \new_[26912]_ ,
    \new_[26915]_ , \new_[26916]_ , \new_[26917]_ , \new_[26920]_ ,
    \new_[26923]_ , \new_[26924]_ , \new_[26927]_ , \new_[26930]_ ,
    \new_[26931]_ , \new_[26932]_ , \new_[26936]_ , \new_[26937]_ ,
    \new_[26940]_ , \new_[26943]_ , \new_[26944]_ , \new_[26945]_ ,
    \new_[26948]_ , \new_[26951]_ , \new_[26952]_ , \new_[26955]_ ,
    \new_[26958]_ , \new_[26959]_ , \new_[26960]_ , \new_[26964]_ ,
    \new_[26965]_ , \new_[26968]_ , \new_[26971]_ , \new_[26972]_ ,
    \new_[26973]_ , \new_[26976]_ , \new_[26979]_ , \new_[26980]_ ,
    \new_[26983]_ , \new_[26986]_ , \new_[26987]_ , \new_[26988]_ ,
    \new_[26992]_ , \new_[26993]_ , \new_[26996]_ , \new_[26999]_ ,
    \new_[27000]_ , \new_[27001]_ , \new_[27004]_ , \new_[27007]_ ,
    \new_[27008]_ , \new_[27011]_ , \new_[27014]_ , \new_[27015]_ ,
    \new_[27016]_ , \new_[27020]_ , \new_[27021]_ , \new_[27024]_ ,
    \new_[27027]_ , \new_[27028]_ , \new_[27029]_ , \new_[27032]_ ,
    \new_[27035]_ , \new_[27036]_ , \new_[27039]_ , \new_[27042]_ ,
    \new_[27043]_ , \new_[27044]_ , \new_[27048]_ , \new_[27049]_ ,
    \new_[27052]_ , \new_[27055]_ , \new_[27056]_ , \new_[27057]_ ,
    \new_[27060]_ , \new_[27063]_ , \new_[27064]_ , \new_[27067]_ ,
    \new_[27070]_ , \new_[27071]_ , \new_[27072]_ , \new_[27076]_ ,
    \new_[27077]_ , \new_[27080]_ , \new_[27083]_ , \new_[27084]_ ,
    \new_[27085]_ , \new_[27088]_ , \new_[27091]_ , \new_[27092]_ ,
    \new_[27095]_ , \new_[27098]_ , \new_[27099]_ , \new_[27100]_ ,
    \new_[27104]_ , \new_[27105]_ , \new_[27108]_ , \new_[27111]_ ,
    \new_[27112]_ , \new_[27113]_ , \new_[27116]_ , \new_[27119]_ ,
    \new_[27120]_ , \new_[27123]_ , \new_[27126]_ , \new_[27127]_ ,
    \new_[27128]_ , \new_[27132]_ , \new_[27133]_ , \new_[27136]_ ,
    \new_[27139]_ , \new_[27140]_ , \new_[27141]_ , \new_[27144]_ ,
    \new_[27147]_ , \new_[27148]_ , \new_[27151]_ , \new_[27154]_ ,
    \new_[27155]_ , \new_[27156]_ , \new_[27160]_ , \new_[27161]_ ,
    \new_[27164]_ , \new_[27167]_ , \new_[27168]_ , \new_[27169]_ ,
    \new_[27172]_ , \new_[27175]_ , \new_[27176]_ , \new_[27179]_ ,
    \new_[27182]_ , \new_[27183]_ , \new_[27184]_ , \new_[27188]_ ,
    \new_[27189]_ , \new_[27192]_ , \new_[27195]_ , \new_[27196]_ ,
    \new_[27197]_ , \new_[27200]_ , \new_[27203]_ , \new_[27204]_ ,
    \new_[27207]_ , \new_[27210]_ , \new_[27211]_ , \new_[27212]_ ,
    \new_[27216]_ , \new_[27217]_ , \new_[27220]_ , \new_[27223]_ ,
    \new_[27224]_ , \new_[27225]_ , \new_[27228]_ , \new_[27231]_ ,
    \new_[27232]_ , \new_[27235]_ , \new_[27238]_ , \new_[27239]_ ,
    \new_[27240]_ , \new_[27244]_ , \new_[27245]_ , \new_[27248]_ ,
    \new_[27251]_ , \new_[27252]_ , \new_[27253]_ , \new_[27256]_ ,
    \new_[27259]_ , \new_[27260]_ , \new_[27263]_ , \new_[27266]_ ,
    \new_[27267]_ , \new_[27268]_ , \new_[27272]_ , \new_[27273]_ ,
    \new_[27276]_ , \new_[27279]_ , \new_[27280]_ , \new_[27281]_ ,
    \new_[27284]_ , \new_[27287]_ , \new_[27288]_ , \new_[27291]_ ,
    \new_[27294]_ , \new_[27295]_ , \new_[27296]_ , \new_[27300]_ ,
    \new_[27301]_ , \new_[27304]_ , \new_[27307]_ , \new_[27308]_ ,
    \new_[27309]_ , \new_[27312]_ , \new_[27315]_ , \new_[27316]_ ,
    \new_[27319]_ , \new_[27322]_ , \new_[27323]_ , \new_[27324]_ ,
    \new_[27328]_ , \new_[27329]_ , \new_[27332]_ , \new_[27335]_ ,
    \new_[27336]_ , \new_[27337]_ , \new_[27340]_ , \new_[27343]_ ,
    \new_[27344]_ , \new_[27347]_ , \new_[27350]_ , \new_[27351]_ ,
    \new_[27352]_ , \new_[27356]_ , \new_[27357]_ , \new_[27360]_ ,
    \new_[27363]_ , \new_[27364]_ , \new_[27365]_ , \new_[27368]_ ,
    \new_[27371]_ , \new_[27372]_ , \new_[27375]_ , \new_[27378]_ ,
    \new_[27379]_ , \new_[27380]_ , \new_[27384]_ , \new_[27385]_ ,
    \new_[27388]_ , \new_[27391]_ , \new_[27392]_ , \new_[27393]_ ,
    \new_[27396]_ , \new_[27399]_ , \new_[27400]_ , \new_[27403]_ ,
    \new_[27406]_ , \new_[27407]_ , \new_[27408]_ , \new_[27412]_ ,
    \new_[27413]_ , \new_[27416]_ , \new_[27419]_ , \new_[27420]_ ,
    \new_[27421]_ , \new_[27424]_ , \new_[27427]_ , \new_[27428]_ ,
    \new_[27431]_ , \new_[27434]_ , \new_[27435]_ , \new_[27436]_ ,
    \new_[27440]_ , \new_[27441]_ , \new_[27444]_ , \new_[27447]_ ,
    \new_[27448]_ , \new_[27449]_ , \new_[27452]_ , \new_[27455]_ ,
    \new_[27456]_ , \new_[27459]_ , \new_[27462]_ , \new_[27463]_ ,
    \new_[27464]_ , \new_[27468]_ , \new_[27469]_ , \new_[27472]_ ,
    \new_[27475]_ , \new_[27476]_ , \new_[27477]_ , \new_[27480]_ ,
    \new_[27483]_ , \new_[27484]_ , \new_[27487]_ , \new_[27490]_ ,
    \new_[27491]_ , \new_[27492]_ , \new_[27496]_ , \new_[27497]_ ,
    \new_[27500]_ , \new_[27503]_ , \new_[27504]_ , \new_[27505]_ ,
    \new_[27508]_ , \new_[27511]_ , \new_[27512]_ , \new_[27515]_ ,
    \new_[27518]_ , \new_[27519]_ , \new_[27520]_ , \new_[27524]_ ,
    \new_[27525]_ , \new_[27528]_ , \new_[27531]_ , \new_[27532]_ ,
    \new_[27533]_ , \new_[27536]_ , \new_[27539]_ , \new_[27540]_ ,
    \new_[27543]_ , \new_[27546]_ , \new_[27547]_ , \new_[27548]_ ,
    \new_[27552]_ , \new_[27553]_ , \new_[27556]_ , \new_[27559]_ ,
    \new_[27560]_ , \new_[27561]_ , \new_[27564]_ , \new_[27567]_ ,
    \new_[27568]_ , \new_[27571]_ , \new_[27574]_ , \new_[27575]_ ,
    \new_[27576]_ , \new_[27580]_ , \new_[27581]_ , \new_[27584]_ ,
    \new_[27587]_ , \new_[27588]_ , \new_[27589]_ , \new_[27592]_ ,
    \new_[27595]_ , \new_[27596]_ , \new_[27599]_ , \new_[27602]_ ,
    \new_[27603]_ , \new_[27604]_ , \new_[27608]_ , \new_[27609]_ ,
    \new_[27612]_ , \new_[27615]_ , \new_[27616]_ , \new_[27617]_ ,
    \new_[27620]_ , \new_[27623]_ , \new_[27624]_ , \new_[27627]_ ,
    \new_[27630]_ , \new_[27631]_ , \new_[27632]_ , \new_[27636]_ ,
    \new_[27637]_ , \new_[27640]_ , \new_[27643]_ , \new_[27644]_ ,
    \new_[27645]_ , \new_[27648]_ , \new_[27651]_ , \new_[27652]_ ,
    \new_[27655]_ , \new_[27658]_ , \new_[27659]_ , \new_[27660]_ ,
    \new_[27664]_ , \new_[27665]_ , \new_[27668]_ , \new_[27671]_ ,
    \new_[27672]_ , \new_[27673]_ , \new_[27676]_ , \new_[27679]_ ,
    \new_[27680]_ , \new_[27683]_ , \new_[27686]_ , \new_[27687]_ ,
    \new_[27688]_ , \new_[27692]_ , \new_[27693]_ , \new_[27696]_ ,
    \new_[27699]_ , \new_[27700]_ , \new_[27701]_ , \new_[27704]_ ,
    \new_[27707]_ , \new_[27708]_ , \new_[27711]_ , \new_[27714]_ ,
    \new_[27715]_ , \new_[27716]_ , \new_[27720]_ , \new_[27721]_ ,
    \new_[27724]_ , \new_[27727]_ , \new_[27728]_ , \new_[27729]_ ,
    \new_[27732]_ , \new_[27735]_ , \new_[27736]_ , \new_[27739]_ ,
    \new_[27742]_ , \new_[27743]_ , \new_[27744]_ , \new_[27748]_ ,
    \new_[27749]_ , \new_[27752]_ , \new_[27755]_ , \new_[27756]_ ,
    \new_[27757]_ , \new_[27760]_ , \new_[27763]_ , \new_[27764]_ ,
    \new_[27767]_ , \new_[27770]_ , \new_[27771]_ , \new_[27772]_ ,
    \new_[27776]_ , \new_[27777]_ , \new_[27780]_ , \new_[27783]_ ,
    \new_[27784]_ , \new_[27785]_ , \new_[27788]_ , \new_[27791]_ ,
    \new_[27792]_ , \new_[27795]_ , \new_[27798]_ , \new_[27799]_ ,
    \new_[27800]_ , \new_[27804]_ , \new_[27805]_ , \new_[27808]_ ,
    \new_[27811]_ , \new_[27812]_ , \new_[27813]_ , \new_[27816]_ ,
    \new_[27819]_ , \new_[27820]_ , \new_[27823]_ , \new_[27826]_ ,
    \new_[27827]_ , \new_[27828]_ , \new_[27832]_ , \new_[27833]_ ,
    \new_[27836]_ , \new_[27839]_ , \new_[27840]_ , \new_[27841]_ ,
    \new_[27844]_ , \new_[27847]_ , \new_[27848]_ , \new_[27851]_ ,
    \new_[27854]_ , \new_[27855]_ , \new_[27856]_ , \new_[27860]_ ,
    \new_[27861]_ , \new_[27864]_ , \new_[27867]_ , \new_[27868]_ ,
    \new_[27869]_ , \new_[27872]_ , \new_[27875]_ , \new_[27876]_ ,
    \new_[27879]_ , \new_[27882]_ , \new_[27883]_ , \new_[27884]_ ,
    \new_[27888]_ , \new_[27889]_ , \new_[27892]_ , \new_[27895]_ ,
    \new_[27896]_ , \new_[27897]_ , \new_[27900]_ , \new_[27903]_ ,
    \new_[27904]_ , \new_[27907]_ , \new_[27910]_ , \new_[27911]_ ,
    \new_[27912]_ , \new_[27916]_ , \new_[27917]_ , \new_[27920]_ ,
    \new_[27923]_ , \new_[27924]_ , \new_[27925]_ , \new_[27928]_ ,
    \new_[27931]_ , \new_[27932]_ , \new_[27935]_ , \new_[27938]_ ,
    \new_[27939]_ , \new_[27940]_ , \new_[27944]_ , \new_[27945]_ ,
    \new_[27948]_ , \new_[27951]_ , \new_[27952]_ , \new_[27953]_ ,
    \new_[27956]_ , \new_[27959]_ , \new_[27960]_ , \new_[27963]_ ,
    \new_[27966]_ , \new_[27967]_ , \new_[27968]_ , \new_[27972]_ ,
    \new_[27973]_ , \new_[27976]_ , \new_[27979]_ , \new_[27980]_ ,
    \new_[27981]_ , \new_[27984]_ , \new_[27987]_ , \new_[27988]_ ,
    \new_[27991]_ , \new_[27994]_ , \new_[27995]_ , \new_[27996]_ ,
    \new_[28000]_ , \new_[28001]_ , \new_[28004]_ , \new_[28007]_ ,
    \new_[28008]_ , \new_[28009]_ , \new_[28012]_ , \new_[28015]_ ,
    \new_[28016]_ , \new_[28019]_ , \new_[28022]_ , \new_[28023]_ ,
    \new_[28024]_ , \new_[28028]_ , \new_[28029]_ , \new_[28032]_ ,
    \new_[28035]_ , \new_[28036]_ , \new_[28037]_ , \new_[28040]_ ,
    \new_[28043]_ , \new_[28044]_ , \new_[28047]_ , \new_[28050]_ ,
    \new_[28051]_ , \new_[28052]_ , \new_[28056]_ , \new_[28057]_ ,
    \new_[28060]_ , \new_[28063]_ , \new_[28064]_ , \new_[28065]_ ,
    \new_[28068]_ , \new_[28071]_ , \new_[28072]_ , \new_[28075]_ ,
    \new_[28078]_ , \new_[28079]_ , \new_[28080]_ , \new_[28084]_ ,
    \new_[28085]_ , \new_[28088]_ , \new_[28091]_ , \new_[28092]_ ,
    \new_[28093]_ , \new_[28096]_ , \new_[28099]_ , \new_[28100]_ ,
    \new_[28103]_ , \new_[28106]_ , \new_[28107]_ , \new_[28108]_ ,
    \new_[28112]_ , \new_[28113]_ , \new_[28116]_ , \new_[28119]_ ,
    \new_[28120]_ , \new_[28121]_ , \new_[28124]_ , \new_[28127]_ ,
    \new_[28128]_ , \new_[28131]_ , \new_[28134]_ , \new_[28135]_ ,
    \new_[28136]_ , \new_[28140]_ , \new_[28141]_ , \new_[28144]_ ,
    \new_[28147]_ , \new_[28148]_ , \new_[28149]_ , \new_[28152]_ ,
    \new_[28155]_ , \new_[28156]_ , \new_[28159]_ , \new_[28162]_ ,
    \new_[28163]_ , \new_[28164]_ , \new_[28168]_ , \new_[28169]_ ,
    \new_[28172]_ , \new_[28175]_ , \new_[28176]_ , \new_[28177]_ ,
    \new_[28180]_ , \new_[28183]_ , \new_[28184]_ , \new_[28187]_ ,
    \new_[28190]_ , \new_[28191]_ , \new_[28192]_ , \new_[28196]_ ,
    \new_[28197]_ , \new_[28200]_ , \new_[28203]_ , \new_[28204]_ ,
    \new_[28205]_ , \new_[28208]_ , \new_[28211]_ , \new_[28212]_ ,
    \new_[28215]_ , \new_[28218]_ , \new_[28219]_ , \new_[28220]_ ,
    \new_[28224]_ , \new_[28225]_ , \new_[28228]_ , \new_[28231]_ ,
    \new_[28232]_ , \new_[28233]_ , \new_[28236]_ , \new_[28239]_ ,
    \new_[28240]_ , \new_[28243]_ , \new_[28246]_ , \new_[28247]_ ,
    \new_[28248]_ , \new_[28252]_ , \new_[28253]_ , \new_[28256]_ ,
    \new_[28259]_ , \new_[28260]_ , \new_[28261]_ , \new_[28264]_ ,
    \new_[28267]_ , \new_[28268]_ , \new_[28271]_ , \new_[28274]_ ,
    \new_[28275]_ , \new_[28276]_ , \new_[28280]_ , \new_[28281]_ ,
    \new_[28284]_ , \new_[28287]_ , \new_[28288]_ , \new_[28289]_ ,
    \new_[28292]_ , \new_[28295]_ , \new_[28296]_ , \new_[28299]_ ,
    \new_[28302]_ , \new_[28303]_ , \new_[28304]_ , \new_[28308]_ ,
    \new_[28309]_ , \new_[28312]_ , \new_[28315]_ , \new_[28316]_ ,
    \new_[28317]_ , \new_[28320]_ , \new_[28323]_ , \new_[28324]_ ,
    \new_[28327]_ , \new_[28330]_ , \new_[28331]_ , \new_[28332]_ ,
    \new_[28336]_ , \new_[28337]_ , \new_[28340]_ , \new_[28343]_ ,
    \new_[28344]_ , \new_[28345]_ , \new_[28348]_ , \new_[28351]_ ,
    \new_[28352]_ , \new_[28355]_ , \new_[28358]_ , \new_[28359]_ ,
    \new_[28360]_ , \new_[28364]_ , \new_[28365]_ , \new_[28368]_ ,
    \new_[28371]_ , \new_[28372]_ , \new_[28373]_ , \new_[28376]_ ,
    \new_[28379]_ , \new_[28380]_ , \new_[28383]_ , \new_[28386]_ ,
    \new_[28387]_ , \new_[28388]_ , \new_[28392]_ , \new_[28393]_ ,
    \new_[28396]_ , \new_[28399]_ , \new_[28400]_ , \new_[28401]_ ,
    \new_[28404]_ , \new_[28407]_ , \new_[28408]_ , \new_[28411]_ ,
    \new_[28414]_ , \new_[28415]_ , \new_[28416]_ , \new_[28420]_ ,
    \new_[28421]_ , \new_[28424]_ , \new_[28427]_ , \new_[28428]_ ,
    \new_[28429]_ , \new_[28432]_ , \new_[28435]_ , \new_[28436]_ ,
    \new_[28439]_ , \new_[28442]_ , \new_[28443]_ , \new_[28444]_ ,
    \new_[28448]_ , \new_[28449]_ , \new_[28452]_ , \new_[28455]_ ,
    \new_[28456]_ , \new_[28457]_ , \new_[28460]_ , \new_[28463]_ ,
    \new_[28464]_ , \new_[28467]_ , \new_[28470]_ , \new_[28471]_ ,
    \new_[28472]_ , \new_[28476]_ , \new_[28477]_ , \new_[28480]_ ,
    \new_[28483]_ , \new_[28484]_ , \new_[28485]_ , \new_[28488]_ ,
    \new_[28491]_ , \new_[28492]_ , \new_[28495]_ , \new_[28498]_ ,
    \new_[28499]_ , \new_[28500]_ , \new_[28504]_ , \new_[28505]_ ,
    \new_[28508]_ , \new_[28511]_ , \new_[28512]_ , \new_[28513]_ ,
    \new_[28516]_ , \new_[28519]_ , \new_[28520]_ , \new_[28523]_ ,
    \new_[28526]_ , \new_[28527]_ , \new_[28528]_ , \new_[28532]_ ,
    \new_[28533]_ , \new_[28536]_ , \new_[28539]_ , \new_[28540]_ ,
    \new_[28541]_ , \new_[28544]_ , \new_[28547]_ , \new_[28548]_ ,
    \new_[28551]_ , \new_[28554]_ , \new_[28555]_ , \new_[28556]_ ,
    \new_[28560]_ , \new_[28561]_ , \new_[28564]_ , \new_[28567]_ ,
    \new_[28568]_ , \new_[28569]_ , \new_[28572]_ , \new_[28575]_ ,
    \new_[28576]_ , \new_[28579]_ , \new_[28582]_ , \new_[28583]_ ,
    \new_[28584]_ , \new_[28588]_ , \new_[28589]_ , \new_[28592]_ ,
    \new_[28595]_ , \new_[28596]_ , \new_[28597]_ , \new_[28600]_ ,
    \new_[28603]_ , \new_[28604]_ , \new_[28607]_ , \new_[28610]_ ,
    \new_[28611]_ , \new_[28612]_ , \new_[28616]_ , \new_[28617]_ ,
    \new_[28620]_ , \new_[28623]_ , \new_[28624]_ , \new_[28625]_ ,
    \new_[28628]_ , \new_[28631]_ , \new_[28632]_ , \new_[28635]_ ,
    \new_[28638]_ , \new_[28639]_ , \new_[28640]_ , \new_[28644]_ ,
    \new_[28645]_ , \new_[28648]_ , \new_[28651]_ , \new_[28652]_ ,
    \new_[28653]_ , \new_[28656]_ , \new_[28659]_ , \new_[28660]_ ,
    \new_[28663]_ , \new_[28666]_ , \new_[28667]_ , \new_[28668]_ ,
    \new_[28672]_ , \new_[28673]_ , \new_[28676]_ , \new_[28679]_ ,
    \new_[28680]_ , \new_[28681]_ , \new_[28684]_ , \new_[28687]_ ,
    \new_[28688]_ , \new_[28691]_ , \new_[28694]_ , \new_[28695]_ ,
    \new_[28696]_ , \new_[28700]_ , \new_[28701]_ , \new_[28704]_ ,
    \new_[28707]_ , \new_[28708]_ , \new_[28709]_ , \new_[28712]_ ,
    \new_[28715]_ , \new_[28716]_ , \new_[28719]_ , \new_[28722]_ ,
    \new_[28723]_ , \new_[28724]_ , \new_[28728]_ , \new_[28729]_ ,
    \new_[28732]_ , \new_[28735]_ , \new_[28736]_ , \new_[28737]_ ,
    \new_[28740]_ , \new_[28743]_ , \new_[28744]_ , \new_[28747]_ ,
    \new_[28750]_ , \new_[28751]_ , \new_[28752]_ , \new_[28756]_ ,
    \new_[28757]_ , \new_[28760]_ , \new_[28763]_ , \new_[28764]_ ,
    \new_[28765]_ , \new_[28768]_ , \new_[28771]_ , \new_[28772]_ ,
    \new_[28775]_ , \new_[28778]_ , \new_[28779]_ , \new_[28780]_ ,
    \new_[28784]_ , \new_[28785]_ , \new_[28788]_ , \new_[28791]_ ,
    \new_[28792]_ , \new_[28793]_ , \new_[28796]_ , \new_[28799]_ ,
    \new_[28800]_ , \new_[28803]_ , \new_[28806]_ , \new_[28807]_ ,
    \new_[28808]_ , \new_[28812]_ , \new_[28813]_ , \new_[28816]_ ,
    \new_[28819]_ , \new_[28820]_ , \new_[28821]_ , \new_[28824]_ ,
    \new_[28827]_ , \new_[28828]_ , \new_[28831]_ , \new_[28834]_ ,
    \new_[28835]_ , \new_[28836]_ , \new_[28840]_ , \new_[28841]_ ,
    \new_[28844]_ , \new_[28847]_ , \new_[28848]_ , \new_[28849]_ ,
    \new_[28852]_ , \new_[28855]_ , \new_[28856]_ , \new_[28859]_ ,
    \new_[28862]_ , \new_[28863]_ , \new_[28864]_ , \new_[28868]_ ,
    \new_[28869]_ , \new_[28872]_ , \new_[28875]_ , \new_[28876]_ ,
    \new_[28877]_ , \new_[28880]_ , \new_[28883]_ , \new_[28884]_ ,
    \new_[28887]_ , \new_[28890]_ , \new_[28891]_ , \new_[28892]_ ,
    \new_[28896]_ , \new_[28897]_ , \new_[28900]_ , \new_[28903]_ ,
    \new_[28904]_ , \new_[28905]_ , \new_[28908]_ , \new_[28911]_ ,
    \new_[28912]_ , \new_[28915]_ , \new_[28918]_ , \new_[28919]_ ,
    \new_[28920]_ , \new_[28924]_ , \new_[28925]_ , \new_[28928]_ ,
    \new_[28931]_ , \new_[28932]_ , \new_[28933]_ , \new_[28936]_ ,
    \new_[28939]_ , \new_[28940]_ , \new_[28943]_ , \new_[28946]_ ,
    \new_[28947]_ , \new_[28948]_ , \new_[28952]_ , \new_[28953]_ ,
    \new_[28956]_ , \new_[28959]_ , \new_[28960]_ , \new_[28961]_ ,
    \new_[28964]_ , \new_[28967]_ , \new_[28968]_ , \new_[28971]_ ,
    \new_[28974]_ , \new_[28975]_ , \new_[28976]_ , \new_[28980]_ ,
    \new_[28981]_ , \new_[28984]_ , \new_[28987]_ , \new_[28988]_ ,
    \new_[28989]_ , \new_[28992]_ , \new_[28995]_ , \new_[28996]_ ,
    \new_[28999]_ , \new_[29002]_ , \new_[29003]_ , \new_[29004]_ ,
    \new_[29008]_ , \new_[29009]_ , \new_[29012]_ , \new_[29015]_ ,
    \new_[29016]_ , \new_[29017]_ , \new_[29020]_ , \new_[29023]_ ,
    \new_[29024]_ , \new_[29027]_ , \new_[29030]_ , \new_[29031]_ ,
    \new_[29032]_ , \new_[29036]_ , \new_[29037]_ , \new_[29040]_ ,
    \new_[29043]_ , \new_[29044]_ , \new_[29045]_ , \new_[29048]_ ,
    \new_[29051]_ , \new_[29052]_ , \new_[29055]_ , \new_[29058]_ ,
    \new_[29059]_ , \new_[29060]_ , \new_[29064]_ , \new_[29065]_ ,
    \new_[29068]_ , \new_[29071]_ , \new_[29072]_ , \new_[29073]_ ,
    \new_[29076]_ , \new_[29079]_ , \new_[29080]_ , \new_[29083]_ ,
    \new_[29086]_ , \new_[29087]_ , \new_[29088]_ , \new_[29092]_ ,
    \new_[29093]_ , \new_[29096]_ , \new_[29099]_ , \new_[29100]_ ,
    \new_[29101]_ , \new_[29104]_ , \new_[29107]_ , \new_[29108]_ ,
    \new_[29111]_ , \new_[29114]_ , \new_[29115]_ , \new_[29116]_ ,
    \new_[29120]_ , \new_[29121]_ , \new_[29124]_ , \new_[29127]_ ,
    \new_[29128]_ , \new_[29129]_ , \new_[29132]_ , \new_[29135]_ ,
    \new_[29136]_ , \new_[29139]_ , \new_[29142]_ , \new_[29143]_ ,
    \new_[29144]_ , \new_[29148]_ , \new_[29149]_ , \new_[29152]_ ,
    \new_[29155]_ , \new_[29156]_ , \new_[29157]_ , \new_[29160]_ ,
    \new_[29163]_ , \new_[29164]_ , \new_[29167]_ , \new_[29170]_ ,
    \new_[29171]_ , \new_[29172]_ , \new_[29176]_ , \new_[29177]_ ,
    \new_[29180]_ , \new_[29183]_ , \new_[29184]_ , \new_[29185]_ ,
    \new_[29188]_ , \new_[29191]_ , \new_[29192]_ , \new_[29195]_ ,
    \new_[29198]_ , \new_[29199]_ , \new_[29200]_ , \new_[29204]_ ,
    \new_[29205]_ , \new_[29208]_ , \new_[29211]_ , \new_[29212]_ ,
    \new_[29213]_ , \new_[29216]_ , \new_[29219]_ , \new_[29220]_ ,
    \new_[29223]_ , \new_[29226]_ , \new_[29227]_ , \new_[29228]_ ,
    \new_[29232]_ , \new_[29233]_ , \new_[29236]_ , \new_[29239]_ ,
    \new_[29240]_ , \new_[29241]_ , \new_[29244]_ , \new_[29247]_ ,
    \new_[29248]_ , \new_[29251]_ , \new_[29254]_ , \new_[29255]_ ,
    \new_[29256]_ , \new_[29260]_ , \new_[29261]_ , \new_[29264]_ ,
    \new_[29267]_ , \new_[29268]_ , \new_[29269]_ , \new_[29272]_ ,
    \new_[29275]_ , \new_[29276]_ , \new_[29279]_ , \new_[29282]_ ,
    \new_[29283]_ , \new_[29284]_ , \new_[29288]_ , \new_[29289]_ ,
    \new_[29292]_ , \new_[29295]_ , \new_[29296]_ , \new_[29297]_ ,
    \new_[29300]_ , \new_[29303]_ , \new_[29304]_ , \new_[29307]_ ,
    \new_[29310]_ , \new_[29311]_ , \new_[29312]_ , \new_[29316]_ ,
    \new_[29317]_ , \new_[29320]_ , \new_[29323]_ , \new_[29324]_ ,
    \new_[29325]_ , \new_[29328]_ , \new_[29331]_ , \new_[29332]_ ,
    \new_[29335]_ , \new_[29338]_ , \new_[29339]_ , \new_[29340]_ ,
    \new_[29344]_ , \new_[29345]_ , \new_[29348]_ , \new_[29351]_ ,
    \new_[29352]_ , \new_[29353]_ , \new_[29356]_ , \new_[29359]_ ,
    \new_[29360]_ , \new_[29363]_ , \new_[29366]_ , \new_[29367]_ ,
    \new_[29368]_ , \new_[29372]_ , \new_[29373]_ , \new_[29376]_ ,
    \new_[29379]_ , \new_[29380]_ , \new_[29381]_ , \new_[29384]_ ,
    \new_[29387]_ , \new_[29388]_ , \new_[29391]_ , \new_[29394]_ ,
    \new_[29395]_ , \new_[29396]_ , \new_[29400]_ , \new_[29401]_ ,
    \new_[29404]_ , \new_[29407]_ , \new_[29408]_ , \new_[29409]_ ,
    \new_[29412]_ , \new_[29415]_ , \new_[29416]_ , \new_[29419]_ ,
    \new_[29422]_ , \new_[29423]_ , \new_[29424]_ , \new_[29428]_ ,
    \new_[29429]_ , \new_[29432]_ , \new_[29435]_ , \new_[29436]_ ,
    \new_[29437]_ , \new_[29440]_ , \new_[29443]_ , \new_[29444]_ ,
    \new_[29447]_ , \new_[29450]_ , \new_[29451]_ , \new_[29452]_ ,
    \new_[29456]_ , \new_[29457]_ , \new_[29460]_ , \new_[29463]_ ,
    \new_[29464]_ , \new_[29465]_ , \new_[29468]_ , \new_[29471]_ ,
    \new_[29472]_ , \new_[29475]_ , \new_[29478]_ , \new_[29479]_ ,
    \new_[29480]_ , \new_[29484]_ , \new_[29485]_ , \new_[29488]_ ,
    \new_[29491]_ , \new_[29492]_ , \new_[29493]_ , \new_[29496]_ ,
    \new_[29499]_ , \new_[29500]_ , \new_[29503]_ , \new_[29506]_ ,
    \new_[29507]_ , \new_[29508]_ , \new_[29512]_ , \new_[29513]_ ,
    \new_[29516]_ , \new_[29519]_ , \new_[29520]_ , \new_[29521]_ ,
    \new_[29524]_ , \new_[29527]_ , \new_[29528]_ , \new_[29531]_ ,
    \new_[29534]_ , \new_[29535]_ , \new_[29536]_ , \new_[29540]_ ,
    \new_[29541]_ , \new_[29544]_ , \new_[29547]_ , \new_[29548]_ ,
    \new_[29549]_ , \new_[29552]_ , \new_[29555]_ , \new_[29556]_ ,
    \new_[29559]_ , \new_[29562]_ , \new_[29563]_ , \new_[29564]_ ,
    \new_[29568]_ , \new_[29569]_ , \new_[29572]_ , \new_[29575]_ ,
    \new_[29576]_ , \new_[29577]_ , \new_[29580]_ , \new_[29583]_ ,
    \new_[29584]_ , \new_[29587]_ , \new_[29590]_ , \new_[29591]_ ,
    \new_[29592]_ , \new_[29596]_ , \new_[29597]_ , \new_[29600]_ ,
    \new_[29603]_ , \new_[29604]_ , \new_[29605]_ , \new_[29608]_ ,
    \new_[29611]_ , \new_[29612]_ , \new_[29615]_ , \new_[29618]_ ,
    \new_[29619]_ , \new_[29620]_ , \new_[29624]_ , \new_[29625]_ ,
    \new_[29628]_ , \new_[29631]_ , \new_[29632]_ , \new_[29633]_ ,
    \new_[29636]_ , \new_[29639]_ , \new_[29640]_ , \new_[29643]_ ,
    \new_[29646]_ , \new_[29647]_ , \new_[29648]_ , \new_[29652]_ ,
    \new_[29653]_ , \new_[29656]_ , \new_[29659]_ , \new_[29660]_ ,
    \new_[29661]_ , \new_[29664]_ , \new_[29667]_ , \new_[29668]_ ,
    \new_[29671]_ , \new_[29674]_ , \new_[29675]_ , \new_[29676]_ ,
    \new_[29680]_ , \new_[29681]_ , \new_[29684]_ , \new_[29687]_ ,
    \new_[29688]_ , \new_[29689]_ , \new_[29692]_ , \new_[29695]_ ,
    \new_[29696]_ , \new_[29699]_ , \new_[29702]_ , \new_[29703]_ ,
    \new_[29704]_ , \new_[29708]_ , \new_[29709]_ , \new_[29712]_ ,
    \new_[29715]_ , \new_[29716]_ , \new_[29717]_ , \new_[29720]_ ,
    \new_[29723]_ , \new_[29724]_ , \new_[29727]_ , \new_[29730]_ ,
    \new_[29731]_ , \new_[29732]_ , \new_[29736]_ , \new_[29737]_ ,
    \new_[29740]_ , \new_[29743]_ , \new_[29744]_ , \new_[29745]_ ,
    \new_[29748]_ , \new_[29751]_ , \new_[29752]_ , \new_[29755]_ ,
    \new_[29758]_ , \new_[29759]_ , \new_[29760]_ , \new_[29764]_ ,
    \new_[29765]_ , \new_[29768]_ , \new_[29771]_ , \new_[29772]_ ,
    \new_[29773]_ , \new_[29776]_ , \new_[29779]_ , \new_[29780]_ ,
    \new_[29783]_ , \new_[29786]_ , \new_[29787]_ , \new_[29788]_ ,
    \new_[29792]_ , \new_[29793]_ , \new_[29796]_ , \new_[29799]_ ,
    \new_[29800]_ , \new_[29801]_ , \new_[29804]_ , \new_[29807]_ ,
    \new_[29808]_ , \new_[29811]_ , \new_[29814]_ , \new_[29815]_ ,
    \new_[29816]_ , \new_[29820]_ , \new_[29821]_ , \new_[29824]_ ,
    \new_[29827]_ , \new_[29828]_ , \new_[29829]_ , \new_[29832]_ ,
    \new_[29835]_ , \new_[29836]_ , \new_[29839]_ , \new_[29842]_ ,
    \new_[29843]_ , \new_[29844]_ , \new_[29848]_ , \new_[29849]_ ,
    \new_[29852]_ , \new_[29855]_ , \new_[29856]_ , \new_[29857]_ ,
    \new_[29860]_ , \new_[29863]_ , \new_[29864]_ , \new_[29867]_ ,
    \new_[29870]_ , \new_[29871]_ , \new_[29872]_ , \new_[29876]_ ,
    \new_[29877]_ , \new_[29880]_ , \new_[29883]_ , \new_[29884]_ ,
    \new_[29885]_ , \new_[29888]_ , \new_[29891]_ , \new_[29892]_ ,
    \new_[29895]_ , \new_[29898]_ , \new_[29899]_ , \new_[29900]_ ,
    \new_[29904]_ , \new_[29905]_ , \new_[29908]_ , \new_[29911]_ ,
    \new_[29912]_ , \new_[29913]_ , \new_[29916]_ , \new_[29919]_ ,
    \new_[29920]_ , \new_[29923]_ , \new_[29926]_ , \new_[29927]_ ,
    \new_[29928]_ , \new_[29932]_ , \new_[29933]_ , \new_[29936]_ ,
    \new_[29939]_ , \new_[29940]_ , \new_[29941]_ , \new_[29944]_ ,
    \new_[29947]_ , \new_[29948]_ , \new_[29951]_ , \new_[29954]_ ,
    \new_[29955]_ , \new_[29956]_ , \new_[29960]_ , \new_[29961]_ ,
    \new_[29964]_ , \new_[29967]_ , \new_[29968]_ , \new_[29969]_ ,
    \new_[29972]_ , \new_[29975]_ , \new_[29976]_ , \new_[29979]_ ,
    \new_[29982]_ , \new_[29983]_ , \new_[29984]_ , \new_[29988]_ ,
    \new_[29989]_ , \new_[29992]_ , \new_[29995]_ , \new_[29996]_ ,
    \new_[29997]_ , \new_[30000]_ , \new_[30003]_ , \new_[30004]_ ,
    \new_[30007]_ , \new_[30010]_ , \new_[30011]_ , \new_[30012]_ ,
    \new_[30016]_ , \new_[30017]_ , \new_[30020]_ , \new_[30023]_ ,
    \new_[30024]_ , \new_[30025]_ , \new_[30028]_ , \new_[30031]_ ,
    \new_[30032]_ , \new_[30035]_ , \new_[30038]_ , \new_[30039]_ ,
    \new_[30040]_ , \new_[30044]_ , \new_[30045]_ , \new_[30048]_ ,
    \new_[30051]_ , \new_[30052]_ , \new_[30053]_ , \new_[30056]_ ,
    \new_[30059]_ , \new_[30060]_ , \new_[30063]_ , \new_[30066]_ ,
    \new_[30067]_ , \new_[30068]_ , \new_[30072]_ , \new_[30073]_ ,
    \new_[30076]_ , \new_[30079]_ , \new_[30080]_ , \new_[30081]_ ,
    \new_[30084]_ , \new_[30087]_ , \new_[30088]_ , \new_[30091]_ ,
    \new_[30094]_ , \new_[30095]_ , \new_[30096]_ , \new_[30100]_ ,
    \new_[30101]_ , \new_[30104]_ , \new_[30107]_ , \new_[30108]_ ,
    \new_[30109]_ , \new_[30112]_ , \new_[30115]_ , \new_[30116]_ ,
    \new_[30119]_ , \new_[30122]_ , \new_[30123]_ , \new_[30124]_ ,
    \new_[30128]_ , \new_[30129]_ , \new_[30132]_ , \new_[30135]_ ,
    \new_[30136]_ , \new_[30137]_ , \new_[30140]_ , \new_[30143]_ ,
    \new_[30144]_ , \new_[30147]_ , \new_[30150]_ , \new_[30151]_ ,
    \new_[30152]_ , \new_[30156]_ , \new_[30157]_ , \new_[30160]_ ,
    \new_[30163]_ , \new_[30164]_ , \new_[30165]_ , \new_[30168]_ ,
    \new_[30171]_ , \new_[30172]_ , \new_[30175]_ , \new_[30178]_ ,
    \new_[30179]_ , \new_[30180]_ , \new_[30184]_ , \new_[30185]_ ,
    \new_[30188]_ , \new_[30191]_ , \new_[30192]_ , \new_[30193]_ ,
    \new_[30196]_ , \new_[30199]_ , \new_[30200]_ , \new_[30203]_ ,
    \new_[30206]_ , \new_[30207]_ , \new_[30208]_ , \new_[30212]_ ,
    \new_[30213]_ , \new_[30216]_ , \new_[30219]_ , \new_[30220]_ ,
    \new_[30221]_ , \new_[30224]_ , \new_[30227]_ , \new_[30228]_ ,
    \new_[30231]_ , \new_[30234]_ , \new_[30235]_ , \new_[30236]_ ,
    \new_[30240]_ , \new_[30241]_ , \new_[30244]_ , \new_[30247]_ ,
    \new_[30248]_ , \new_[30249]_ , \new_[30252]_ , \new_[30255]_ ,
    \new_[30256]_ , \new_[30259]_ , \new_[30262]_ , \new_[30263]_ ,
    \new_[30264]_ , \new_[30268]_ , \new_[30269]_ , \new_[30272]_ ,
    \new_[30275]_ , \new_[30276]_ , \new_[30277]_ , \new_[30280]_ ,
    \new_[30283]_ , \new_[30284]_ , \new_[30287]_ , \new_[30290]_ ,
    \new_[30291]_ , \new_[30292]_ , \new_[30296]_ , \new_[30297]_ ,
    \new_[30300]_ , \new_[30303]_ , \new_[30304]_ , \new_[30305]_ ,
    \new_[30308]_ , \new_[30311]_ , \new_[30312]_ , \new_[30315]_ ,
    \new_[30318]_ , \new_[30319]_ , \new_[30320]_ , \new_[30324]_ ,
    \new_[30325]_ , \new_[30328]_ , \new_[30331]_ , \new_[30332]_ ,
    \new_[30333]_ , \new_[30336]_ , \new_[30339]_ , \new_[30340]_ ,
    \new_[30343]_ , \new_[30346]_ , \new_[30347]_ , \new_[30348]_ ,
    \new_[30352]_ , \new_[30353]_ , \new_[30356]_ , \new_[30359]_ ,
    \new_[30360]_ , \new_[30361]_ , \new_[30364]_ , \new_[30367]_ ,
    \new_[30368]_ , \new_[30371]_ , \new_[30374]_ , \new_[30375]_ ,
    \new_[30376]_ , \new_[30380]_ , \new_[30381]_ , \new_[30384]_ ,
    \new_[30387]_ , \new_[30388]_ , \new_[30389]_ , \new_[30392]_ ,
    \new_[30395]_ , \new_[30396]_ , \new_[30399]_ , \new_[30402]_ ,
    \new_[30403]_ , \new_[30404]_ , \new_[30408]_ , \new_[30409]_ ,
    \new_[30412]_ , \new_[30415]_ , \new_[30416]_ , \new_[30417]_ ,
    \new_[30420]_ , \new_[30423]_ , \new_[30424]_ , \new_[30427]_ ,
    \new_[30430]_ , \new_[30431]_ , \new_[30432]_ , \new_[30436]_ ,
    \new_[30437]_ , \new_[30440]_ , \new_[30443]_ , \new_[30444]_ ,
    \new_[30445]_ , \new_[30448]_ , \new_[30451]_ , \new_[30452]_ ,
    \new_[30455]_ , \new_[30458]_ , \new_[30459]_ , \new_[30460]_ ,
    \new_[30464]_ , \new_[30465]_ , \new_[30468]_ , \new_[30471]_ ,
    \new_[30472]_ , \new_[30473]_ , \new_[30476]_ , \new_[30479]_ ,
    \new_[30480]_ , \new_[30483]_ , \new_[30486]_ , \new_[30487]_ ,
    \new_[30488]_ , \new_[30492]_ , \new_[30493]_ , \new_[30496]_ ,
    \new_[30499]_ , \new_[30500]_ , \new_[30501]_ , \new_[30504]_ ,
    \new_[30507]_ , \new_[30508]_ , \new_[30511]_ , \new_[30514]_ ,
    \new_[30515]_ , \new_[30516]_ , \new_[30520]_ , \new_[30521]_ ,
    \new_[30524]_ , \new_[30527]_ , \new_[30528]_ , \new_[30529]_ ,
    \new_[30532]_ , \new_[30535]_ , \new_[30536]_ , \new_[30539]_ ,
    \new_[30542]_ , \new_[30543]_ , \new_[30544]_ , \new_[30548]_ ,
    \new_[30549]_ , \new_[30552]_ , \new_[30555]_ , \new_[30556]_ ,
    \new_[30557]_ , \new_[30560]_ , \new_[30563]_ , \new_[30564]_ ,
    \new_[30567]_ , \new_[30570]_ , \new_[30571]_ , \new_[30572]_ ,
    \new_[30576]_ , \new_[30577]_ , \new_[30580]_ , \new_[30583]_ ,
    \new_[30584]_ , \new_[30585]_ , \new_[30588]_ , \new_[30591]_ ,
    \new_[30592]_ , \new_[30595]_ , \new_[30598]_ , \new_[30599]_ ,
    \new_[30600]_ , \new_[30604]_ , \new_[30605]_ , \new_[30608]_ ,
    \new_[30611]_ , \new_[30612]_ , \new_[30613]_ , \new_[30616]_ ,
    \new_[30619]_ , \new_[30620]_ , \new_[30623]_ , \new_[30626]_ ,
    \new_[30627]_ , \new_[30628]_ , \new_[30632]_ , \new_[30633]_ ,
    \new_[30636]_ , \new_[30639]_ , \new_[30640]_ , \new_[30641]_ ,
    \new_[30644]_ , \new_[30647]_ , \new_[30648]_ , \new_[30651]_ ,
    \new_[30654]_ , \new_[30655]_ , \new_[30656]_ , \new_[30660]_ ,
    \new_[30661]_ , \new_[30664]_ , \new_[30667]_ , \new_[30668]_ ,
    \new_[30669]_ , \new_[30672]_ , \new_[30675]_ , \new_[30676]_ ,
    \new_[30679]_ , \new_[30682]_ , \new_[30683]_ , \new_[30684]_ ,
    \new_[30688]_ , \new_[30689]_ , \new_[30692]_ , \new_[30695]_ ,
    \new_[30696]_ , \new_[30697]_ , \new_[30700]_ , \new_[30703]_ ,
    \new_[30704]_ , \new_[30707]_ , \new_[30710]_ , \new_[30711]_ ,
    \new_[30712]_ , \new_[30716]_ , \new_[30717]_ , \new_[30720]_ ,
    \new_[30723]_ , \new_[30724]_ , \new_[30725]_ , \new_[30728]_ ,
    \new_[30731]_ , \new_[30732]_ , \new_[30735]_ , \new_[30738]_ ,
    \new_[30739]_ , \new_[30740]_ , \new_[30744]_ , \new_[30745]_ ,
    \new_[30748]_ , \new_[30751]_ , \new_[30752]_ , \new_[30753]_ ,
    \new_[30756]_ , \new_[30759]_ , \new_[30760]_ , \new_[30763]_ ,
    \new_[30766]_ , \new_[30767]_ , \new_[30768]_ , \new_[30772]_ ,
    \new_[30773]_ , \new_[30776]_ , \new_[30779]_ , \new_[30780]_ ,
    \new_[30781]_ , \new_[30784]_ , \new_[30787]_ , \new_[30788]_ ,
    \new_[30791]_ , \new_[30794]_ , \new_[30795]_ , \new_[30796]_ ,
    \new_[30800]_ , \new_[30801]_ , \new_[30804]_ , \new_[30807]_ ,
    \new_[30808]_ , \new_[30809]_ , \new_[30812]_ , \new_[30815]_ ,
    \new_[30816]_ , \new_[30819]_ , \new_[30822]_ , \new_[30823]_ ,
    \new_[30824]_ , \new_[30828]_ , \new_[30829]_ , \new_[30832]_ ,
    \new_[30835]_ , \new_[30836]_ , \new_[30837]_ , \new_[30840]_ ,
    \new_[30843]_ , \new_[30844]_ , \new_[30847]_ , \new_[30850]_ ,
    \new_[30851]_ , \new_[30852]_ , \new_[30856]_ , \new_[30857]_ ,
    \new_[30860]_ , \new_[30863]_ , \new_[30864]_ , \new_[30865]_ ,
    \new_[30868]_ , \new_[30871]_ , \new_[30872]_ , \new_[30875]_ ,
    \new_[30878]_ , \new_[30879]_ , \new_[30880]_ , \new_[30884]_ ,
    \new_[30885]_ , \new_[30888]_ , \new_[30891]_ , \new_[30892]_ ,
    \new_[30893]_ , \new_[30896]_ , \new_[30899]_ , \new_[30900]_ ,
    \new_[30903]_ , \new_[30906]_ , \new_[30907]_ , \new_[30908]_ ,
    \new_[30912]_ , \new_[30913]_ , \new_[30916]_ , \new_[30919]_ ,
    \new_[30920]_ , \new_[30921]_ , \new_[30924]_ , \new_[30927]_ ,
    \new_[30928]_ , \new_[30931]_ , \new_[30934]_ , \new_[30935]_ ,
    \new_[30936]_ , \new_[30940]_ , \new_[30941]_ , \new_[30944]_ ,
    \new_[30947]_ , \new_[30948]_ , \new_[30949]_ , \new_[30952]_ ,
    \new_[30955]_ , \new_[30956]_ , \new_[30959]_ , \new_[30962]_ ,
    \new_[30963]_ , \new_[30964]_ , \new_[30968]_ , \new_[30969]_ ,
    \new_[30972]_ , \new_[30975]_ , \new_[30976]_ , \new_[30977]_ ,
    \new_[30980]_ , \new_[30983]_ , \new_[30984]_ , \new_[30987]_ ,
    \new_[30990]_ , \new_[30991]_ , \new_[30992]_ , \new_[30996]_ ,
    \new_[30997]_ , \new_[31000]_ , \new_[31003]_ , \new_[31004]_ ,
    \new_[31005]_ , \new_[31008]_ , \new_[31011]_ , \new_[31012]_ ,
    \new_[31015]_ , \new_[31018]_ , \new_[31019]_ , \new_[31020]_ ,
    \new_[31024]_ , \new_[31025]_ , \new_[31028]_ , \new_[31031]_ ,
    \new_[31032]_ , \new_[31033]_ , \new_[31036]_ , \new_[31039]_ ,
    \new_[31040]_ , \new_[31043]_ , \new_[31046]_ , \new_[31047]_ ,
    \new_[31048]_ , \new_[31052]_ , \new_[31053]_ , \new_[31056]_ ,
    \new_[31059]_ , \new_[31060]_ , \new_[31061]_ , \new_[31064]_ ,
    \new_[31067]_ , \new_[31068]_ , \new_[31071]_ , \new_[31074]_ ,
    \new_[31075]_ , \new_[31076]_ , \new_[31080]_ , \new_[31081]_ ,
    \new_[31084]_ , \new_[31087]_ , \new_[31088]_ , \new_[31089]_ ,
    \new_[31092]_ , \new_[31095]_ , \new_[31096]_ , \new_[31099]_ ,
    \new_[31102]_ , \new_[31103]_ , \new_[31104]_ , \new_[31108]_ ,
    \new_[31109]_ , \new_[31112]_ , \new_[31115]_ , \new_[31116]_ ,
    \new_[31117]_ , \new_[31120]_ , \new_[31123]_ , \new_[31124]_ ,
    \new_[31127]_ , \new_[31130]_ , \new_[31131]_ , \new_[31132]_ ,
    \new_[31136]_ , \new_[31137]_ , \new_[31140]_ , \new_[31143]_ ,
    \new_[31144]_ , \new_[31145]_ , \new_[31148]_ , \new_[31151]_ ,
    \new_[31152]_ , \new_[31155]_ , \new_[31158]_ , \new_[31159]_ ,
    \new_[31160]_ , \new_[31164]_ , \new_[31165]_ , \new_[31168]_ ,
    \new_[31171]_ , \new_[31172]_ , \new_[31173]_ , \new_[31176]_ ,
    \new_[31179]_ , \new_[31180]_ , \new_[31183]_ , \new_[31186]_ ,
    \new_[31187]_ , \new_[31188]_ , \new_[31192]_ , \new_[31193]_ ,
    \new_[31196]_ , \new_[31199]_ , \new_[31200]_ , \new_[31201]_ ,
    \new_[31204]_ , \new_[31207]_ , \new_[31208]_ , \new_[31211]_ ,
    \new_[31214]_ , \new_[31215]_ , \new_[31216]_ , \new_[31220]_ ,
    \new_[31221]_ , \new_[31224]_ , \new_[31227]_ , \new_[31228]_ ,
    \new_[31229]_ , \new_[31232]_ , \new_[31235]_ , \new_[31236]_ ,
    \new_[31239]_ , \new_[31242]_ , \new_[31243]_ , \new_[31244]_ ,
    \new_[31248]_ , \new_[31249]_ , \new_[31252]_ , \new_[31255]_ ,
    \new_[31256]_ , \new_[31257]_ , \new_[31260]_ , \new_[31263]_ ,
    \new_[31264]_ , \new_[31267]_ , \new_[31270]_ , \new_[31271]_ ,
    \new_[31272]_ , \new_[31276]_ , \new_[31277]_ , \new_[31280]_ ,
    \new_[31283]_ , \new_[31284]_ , \new_[31285]_ , \new_[31288]_ ,
    \new_[31291]_ , \new_[31292]_ , \new_[31295]_ , \new_[31298]_ ,
    \new_[31299]_ , \new_[31300]_ , \new_[31304]_ , \new_[31305]_ ,
    \new_[31308]_ , \new_[31311]_ , \new_[31312]_ , \new_[31313]_ ,
    \new_[31316]_ , \new_[31319]_ , \new_[31320]_ , \new_[31323]_ ,
    \new_[31326]_ , \new_[31327]_ , \new_[31328]_ , \new_[31332]_ ,
    \new_[31333]_ , \new_[31336]_ , \new_[31339]_ , \new_[31340]_ ,
    \new_[31341]_ , \new_[31344]_ , \new_[31347]_ , \new_[31348]_ ,
    \new_[31351]_ , \new_[31354]_ , \new_[31355]_ , \new_[31356]_ ,
    \new_[31360]_ , \new_[31361]_ , \new_[31364]_ , \new_[31367]_ ,
    \new_[31368]_ , \new_[31369]_ , \new_[31372]_ , \new_[31375]_ ,
    \new_[31376]_ , \new_[31379]_ , \new_[31382]_ , \new_[31383]_ ,
    \new_[31384]_ , \new_[31388]_ , \new_[31389]_ , \new_[31392]_ ,
    \new_[31395]_ , \new_[31396]_ , \new_[31397]_ , \new_[31400]_ ,
    \new_[31403]_ , \new_[31404]_ , \new_[31407]_ , \new_[31410]_ ,
    \new_[31411]_ , \new_[31412]_ , \new_[31416]_ , \new_[31417]_ ,
    \new_[31420]_ , \new_[31423]_ , \new_[31424]_ , \new_[31425]_ ,
    \new_[31428]_ , \new_[31431]_ , \new_[31432]_ , \new_[31435]_ ,
    \new_[31438]_ , \new_[31439]_ , \new_[31440]_ , \new_[31444]_ ,
    \new_[31445]_ , \new_[31448]_ , \new_[31451]_ , \new_[31452]_ ,
    \new_[31453]_ , \new_[31456]_ , \new_[31459]_ , \new_[31460]_ ,
    \new_[31463]_ , \new_[31466]_ , \new_[31467]_ , \new_[31468]_ ,
    \new_[31472]_ , \new_[31473]_ , \new_[31476]_ , \new_[31479]_ ,
    \new_[31480]_ , \new_[31481]_ , \new_[31484]_ , \new_[31487]_ ,
    \new_[31488]_ , \new_[31491]_ , \new_[31494]_ , \new_[31495]_ ,
    \new_[31496]_ , \new_[31500]_ , \new_[31501]_ , \new_[31504]_ ,
    \new_[31507]_ , \new_[31508]_ , \new_[31509]_ , \new_[31512]_ ,
    \new_[31515]_ , \new_[31516]_ , \new_[31519]_ , \new_[31522]_ ,
    \new_[31523]_ , \new_[31524]_ , \new_[31528]_ , \new_[31529]_ ,
    \new_[31532]_ , \new_[31535]_ , \new_[31536]_ , \new_[31537]_ ,
    \new_[31540]_ , \new_[31543]_ , \new_[31544]_ , \new_[31547]_ ,
    \new_[31550]_ , \new_[31551]_ , \new_[31552]_ , \new_[31556]_ ,
    \new_[31557]_ , \new_[31560]_ , \new_[31563]_ , \new_[31564]_ ,
    \new_[31565]_ , \new_[31568]_ , \new_[31571]_ , \new_[31572]_ ,
    \new_[31575]_ , \new_[31578]_ , \new_[31579]_ , \new_[31580]_ ,
    \new_[31584]_ , \new_[31585]_ , \new_[31588]_ , \new_[31591]_ ,
    \new_[31592]_ , \new_[31593]_ , \new_[31596]_ , \new_[31599]_ ,
    \new_[31600]_ , \new_[31603]_ , \new_[31606]_ , \new_[31607]_ ,
    \new_[31608]_ , \new_[31612]_ , \new_[31613]_ , \new_[31616]_ ,
    \new_[31619]_ , \new_[31620]_ , \new_[31621]_ , \new_[31624]_ ,
    \new_[31627]_ , \new_[31628]_ , \new_[31631]_ , \new_[31634]_ ,
    \new_[31635]_ , \new_[31636]_ , \new_[31640]_ , \new_[31641]_ ,
    \new_[31644]_ , \new_[31647]_ , \new_[31648]_ , \new_[31649]_ ,
    \new_[31652]_ , \new_[31655]_ , \new_[31656]_ , \new_[31659]_ ,
    \new_[31662]_ , \new_[31663]_ , \new_[31664]_ , \new_[31668]_ ,
    \new_[31669]_ , \new_[31672]_ , \new_[31675]_ , \new_[31676]_ ,
    \new_[31677]_ , \new_[31680]_ , \new_[31683]_ , \new_[31684]_ ,
    \new_[31687]_ , \new_[31690]_ , \new_[31691]_ , \new_[31692]_ ,
    \new_[31696]_ , \new_[31697]_ , \new_[31700]_ , \new_[31703]_ ,
    \new_[31704]_ , \new_[31705]_ , \new_[31708]_ , \new_[31711]_ ,
    \new_[31712]_ , \new_[31715]_ , \new_[31718]_ , \new_[31719]_ ,
    \new_[31720]_ , \new_[31724]_ , \new_[31725]_ , \new_[31728]_ ,
    \new_[31731]_ , \new_[31732]_ , \new_[31733]_ , \new_[31736]_ ,
    \new_[31739]_ , \new_[31740]_ , \new_[31743]_ , \new_[31746]_ ,
    \new_[31747]_ , \new_[31748]_ , \new_[31752]_ , \new_[31753]_ ,
    \new_[31756]_ , \new_[31759]_ , \new_[31760]_ , \new_[31761]_ ,
    \new_[31764]_ , \new_[31767]_ , \new_[31768]_ , \new_[31771]_ ,
    \new_[31774]_ , \new_[31775]_ , \new_[31776]_ , \new_[31780]_ ,
    \new_[31781]_ , \new_[31784]_ , \new_[31787]_ , \new_[31788]_ ,
    \new_[31789]_ , \new_[31792]_ , \new_[31795]_ , \new_[31796]_ ,
    \new_[31799]_ , \new_[31802]_ , \new_[31803]_ , \new_[31804]_ ,
    \new_[31808]_ , \new_[31809]_ , \new_[31812]_ , \new_[31815]_ ,
    \new_[31816]_ , \new_[31817]_ , \new_[31820]_ , \new_[31823]_ ,
    \new_[31824]_ , \new_[31827]_ , \new_[31830]_ , \new_[31831]_ ,
    \new_[31832]_ , \new_[31836]_ , \new_[31837]_ , \new_[31840]_ ,
    \new_[31843]_ , \new_[31844]_ , \new_[31845]_ , \new_[31848]_ ,
    \new_[31851]_ , \new_[31852]_ , \new_[31855]_ , \new_[31858]_ ,
    \new_[31859]_ , \new_[31860]_ , \new_[31864]_ , \new_[31865]_ ,
    \new_[31868]_ , \new_[31871]_ , \new_[31872]_ , \new_[31873]_ ,
    \new_[31876]_ , \new_[31879]_ , \new_[31880]_ , \new_[31883]_ ,
    \new_[31886]_ , \new_[31887]_ , \new_[31888]_ , \new_[31892]_ ,
    \new_[31893]_ , \new_[31896]_ , \new_[31899]_ , \new_[31900]_ ,
    \new_[31901]_ , \new_[31904]_ , \new_[31907]_ , \new_[31908]_ ,
    \new_[31911]_ , \new_[31914]_ , \new_[31915]_ , \new_[31916]_ ,
    \new_[31920]_ , \new_[31921]_ , \new_[31924]_ , \new_[31927]_ ,
    \new_[31928]_ , \new_[31929]_ , \new_[31932]_ , \new_[31935]_ ,
    \new_[31936]_ , \new_[31939]_ , \new_[31942]_ , \new_[31943]_ ,
    \new_[31944]_ , \new_[31948]_ , \new_[31949]_ , \new_[31952]_ ,
    \new_[31955]_ , \new_[31956]_ , \new_[31957]_ , \new_[31960]_ ,
    \new_[31963]_ , \new_[31964]_ , \new_[31967]_ , \new_[31970]_ ,
    \new_[31971]_ , \new_[31972]_ , \new_[31976]_ , \new_[31977]_ ,
    \new_[31980]_ , \new_[31983]_ , \new_[31984]_ , \new_[31985]_ ,
    \new_[31988]_ , \new_[31991]_ , \new_[31992]_ , \new_[31995]_ ,
    \new_[31998]_ , \new_[31999]_ , \new_[32000]_ , \new_[32004]_ ,
    \new_[32005]_ , \new_[32008]_ , \new_[32011]_ , \new_[32012]_ ,
    \new_[32013]_ , \new_[32016]_ , \new_[32019]_ , \new_[32020]_ ,
    \new_[32023]_ , \new_[32026]_ , \new_[32027]_ , \new_[32028]_ ,
    \new_[32032]_ , \new_[32033]_ , \new_[32036]_ , \new_[32039]_ ,
    \new_[32040]_ , \new_[32041]_ , \new_[32044]_ , \new_[32047]_ ,
    \new_[32048]_ , \new_[32051]_ , \new_[32054]_ , \new_[32055]_ ,
    \new_[32056]_ , \new_[32060]_ , \new_[32061]_ , \new_[32064]_ ,
    \new_[32067]_ , \new_[32068]_ , \new_[32069]_ , \new_[32072]_ ,
    \new_[32075]_ , \new_[32076]_ , \new_[32079]_ , \new_[32082]_ ,
    \new_[32083]_ , \new_[32084]_ , \new_[32088]_ , \new_[32089]_ ,
    \new_[32092]_ , \new_[32095]_ , \new_[32096]_ , \new_[32097]_ ,
    \new_[32100]_ , \new_[32103]_ , \new_[32104]_ , \new_[32107]_ ,
    \new_[32110]_ , \new_[32111]_ , \new_[32112]_ , \new_[32116]_ ,
    \new_[32117]_ , \new_[32120]_ , \new_[32123]_ , \new_[32124]_ ,
    \new_[32125]_ , \new_[32128]_ , \new_[32131]_ , \new_[32132]_ ,
    \new_[32135]_ , \new_[32138]_ , \new_[32139]_ , \new_[32140]_ ,
    \new_[32144]_ , \new_[32145]_ , \new_[32148]_ , \new_[32151]_ ,
    \new_[32152]_ , \new_[32153]_ , \new_[32156]_ , \new_[32159]_ ,
    \new_[32160]_ , \new_[32163]_ , \new_[32166]_ , \new_[32167]_ ,
    \new_[32168]_ , \new_[32172]_ , \new_[32173]_ , \new_[32176]_ ,
    \new_[32179]_ , \new_[32180]_ , \new_[32181]_ , \new_[32184]_ ,
    \new_[32187]_ , \new_[32188]_ , \new_[32191]_ , \new_[32194]_ ,
    \new_[32195]_ , \new_[32196]_ , \new_[32200]_ , \new_[32201]_ ,
    \new_[32204]_ , \new_[32207]_ , \new_[32208]_ , \new_[32209]_ ,
    \new_[32212]_ , \new_[32215]_ , \new_[32216]_ , \new_[32219]_ ,
    \new_[32222]_ , \new_[32223]_ , \new_[32224]_ , \new_[32228]_ ,
    \new_[32229]_ , \new_[32232]_ , \new_[32235]_ , \new_[32236]_ ,
    \new_[32237]_ , \new_[32240]_ , \new_[32243]_ , \new_[32244]_ ,
    \new_[32247]_ , \new_[32250]_ , \new_[32251]_ , \new_[32252]_ ,
    \new_[32256]_ , \new_[32257]_ , \new_[32260]_ , \new_[32263]_ ,
    \new_[32264]_ , \new_[32265]_ , \new_[32268]_ , \new_[32271]_ ,
    \new_[32272]_ , \new_[32275]_ , \new_[32278]_ , \new_[32279]_ ,
    \new_[32280]_ , \new_[32284]_ , \new_[32285]_ , \new_[32288]_ ,
    \new_[32291]_ , \new_[32292]_ , \new_[32293]_ , \new_[32296]_ ,
    \new_[32299]_ , \new_[32300]_ , \new_[32303]_ , \new_[32306]_ ,
    \new_[32307]_ , \new_[32308]_ , \new_[32312]_ , \new_[32313]_ ,
    \new_[32316]_ , \new_[32319]_ , \new_[32320]_ , \new_[32321]_ ,
    \new_[32324]_ , \new_[32327]_ , \new_[32328]_ , \new_[32331]_ ,
    \new_[32334]_ , \new_[32335]_ , \new_[32336]_ , \new_[32340]_ ,
    \new_[32341]_ , \new_[32344]_ , \new_[32347]_ , \new_[32348]_ ,
    \new_[32349]_ , \new_[32352]_ , \new_[32355]_ , \new_[32356]_ ,
    \new_[32359]_ , \new_[32362]_ , \new_[32363]_ , \new_[32364]_ ,
    \new_[32368]_ , \new_[32369]_ , \new_[32372]_ , \new_[32375]_ ,
    \new_[32376]_ , \new_[32377]_ , \new_[32380]_ , \new_[32383]_ ,
    \new_[32384]_ , \new_[32387]_ , \new_[32390]_ , \new_[32391]_ ,
    \new_[32392]_ , \new_[32396]_ , \new_[32397]_ , \new_[32400]_ ,
    \new_[32403]_ , \new_[32404]_ , \new_[32405]_ , \new_[32408]_ ,
    \new_[32411]_ , \new_[32412]_ , \new_[32415]_ , \new_[32418]_ ,
    \new_[32419]_ , \new_[32420]_ , \new_[32424]_ , \new_[32425]_ ,
    \new_[32428]_ , \new_[32431]_ , \new_[32432]_ , \new_[32433]_ ,
    \new_[32436]_ , \new_[32439]_ , \new_[32440]_ , \new_[32443]_ ,
    \new_[32446]_ , \new_[32447]_ , \new_[32448]_ , \new_[32452]_ ,
    \new_[32453]_ , \new_[32456]_ , \new_[32459]_ , \new_[32460]_ ,
    \new_[32461]_ , \new_[32464]_ , \new_[32467]_ , \new_[32468]_ ,
    \new_[32471]_ , \new_[32474]_ , \new_[32475]_ , \new_[32476]_ ,
    \new_[32480]_ , \new_[32481]_ , \new_[32484]_ , \new_[32487]_ ,
    \new_[32488]_ , \new_[32489]_ , \new_[32492]_ , \new_[32495]_ ,
    \new_[32496]_ , \new_[32499]_ , \new_[32502]_ , \new_[32503]_ ,
    \new_[32504]_ , \new_[32508]_ , \new_[32509]_ , \new_[32512]_ ,
    \new_[32515]_ , \new_[32516]_ , \new_[32517]_ , \new_[32520]_ ,
    \new_[32523]_ , \new_[32524]_ , \new_[32527]_ , \new_[32530]_ ,
    \new_[32531]_ , \new_[32532]_ , \new_[32536]_ , \new_[32537]_ ,
    \new_[32540]_ , \new_[32543]_ , \new_[32544]_ , \new_[32545]_ ,
    \new_[32548]_ , \new_[32551]_ , \new_[32552]_ , \new_[32555]_ ,
    \new_[32558]_ , \new_[32559]_ , \new_[32560]_ , \new_[32564]_ ,
    \new_[32565]_ , \new_[32568]_ , \new_[32571]_ , \new_[32572]_ ,
    \new_[32573]_ , \new_[32576]_ , \new_[32579]_ , \new_[32580]_ ,
    \new_[32583]_ , \new_[32586]_ , \new_[32587]_ , \new_[32588]_ ,
    \new_[32592]_ , \new_[32593]_ , \new_[32596]_ , \new_[32599]_ ,
    \new_[32600]_ , \new_[32601]_ , \new_[32604]_ , \new_[32607]_ ,
    \new_[32608]_ , \new_[32611]_ , \new_[32614]_ , \new_[32615]_ ,
    \new_[32616]_ , \new_[32620]_ , \new_[32621]_ , \new_[32624]_ ,
    \new_[32627]_ , \new_[32628]_ , \new_[32629]_ , \new_[32632]_ ,
    \new_[32635]_ , \new_[32636]_ , \new_[32639]_ , \new_[32642]_ ,
    \new_[32643]_ , \new_[32644]_ , \new_[32648]_ , \new_[32649]_ ,
    \new_[32652]_ , \new_[32655]_ , \new_[32656]_ , \new_[32657]_ ,
    \new_[32660]_ , \new_[32663]_ , \new_[32664]_ , \new_[32667]_ ,
    \new_[32670]_ , \new_[32671]_ , \new_[32672]_ , \new_[32676]_ ,
    \new_[32677]_ , \new_[32680]_ , \new_[32683]_ , \new_[32684]_ ,
    \new_[32685]_ , \new_[32688]_ , \new_[32691]_ , \new_[32692]_ ,
    \new_[32695]_ , \new_[32698]_ , \new_[32699]_ , \new_[32700]_ ,
    \new_[32704]_ , \new_[32705]_ , \new_[32708]_ , \new_[32711]_ ,
    \new_[32712]_ , \new_[32713]_ , \new_[32716]_ , \new_[32719]_ ,
    \new_[32720]_ , \new_[32723]_ , \new_[32726]_ , \new_[32727]_ ,
    \new_[32728]_ , \new_[32732]_ , \new_[32733]_ , \new_[32736]_ ,
    \new_[32739]_ , \new_[32740]_ , \new_[32741]_ , \new_[32744]_ ,
    \new_[32747]_ , \new_[32748]_ , \new_[32751]_ , \new_[32754]_ ,
    \new_[32755]_ , \new_[32756]_ , \new_[32760]_ , \new_[32761]_ ,
    \new_[32764]_ , \new_[32767]_ , \new_[32768]_ , \new_[32769]_ ,
    \new_[32772]_ , \new_[32775]_ , \new_[32776]_ , \new_[32779]_ ,
    \new_[32782]_ , \new_[32783]_ , \new_[32784]_ , \new_[32788]_ ,
    \new_[32789]_ , \new_[32792]_ , \new_[32795]_ , \new_[32796]_ ,
    \new_[32797]_ , \new_[32800]_ , \new_[32803]_ , \new_[32804]_ ,
    \new_[32807]_ , \new_[32810]_ , \new_[32811]_ , \new_[32812]_ ,
    \new_[32816]_ , \new_[32817]_ , \new_[32820]_ , \new_[32823]_ ,
    \new_[32824]_ , \new_[32825]_ , \new_[32828]_ , \new_[32831]_ ,
    \new_[32832]_ , \new_[32835]_ , \new_[32838]_ , \new_[32839]_ ,
    \new_[32840]_ , \new_[32844]_ , \new_[32845]_ , \new_[32848]_ ,
    \new_[32851]_ , \new_[32852]_ , \new_[32853]_ , \new_[32856]_ ,
    \new_[32859]_ , \new_[32860]_ , \new_[32863]_ , \new_[32866]_ ,
    \new_[32867]_ , \new_[32868]_ , \new_[32872]_ , \new_[32873]_ ,
    \new_[32876]_ , \new_[32879]_ , \new_[32880]_ , \new_[32881]_ ,
    \new_[32884]_ , \new_[32887]_ , \new_[32888]_ , \new_[32891]_ ,
    \new_[32894]_ , \new_[32895]_ , \new_[32896]_ , \new_[32900]_ ,
    \new_[32901]_ , \new_[32904]_ , \new_[32907]_ , \new_[32908]_ ,
    \new_[32909]_ , \new_[32912]_ , \new_[32915]_ , \new_[32916]_ ,
    \new_[32919]_ , \new_[32922]_ , \new_[32923]_ , \new_[32924]_ ,
    \new_[32928]_ , \new_[32929]_ , \new_[32932]_ , \new_[32935]_ ,
    \new_[32936]_ , \new_[32937]_ , \new_[32940]_ , \new_[32943]_ ,
    \new_[32944]_ , \new_[32947]_ , \new_[32950]_ , \new_[32951]_ ,
    \new_[32952]_ , \new_[32956]_ , \new_[32957]_ , \new_[32960]_ ,
    \new_[32963]_ , \new_[32964]_ , \new_[32965]_ , \new_[32968]_ ,
    \new_[32971]_ , \new_[32972]_ , \new_[32975]_ , \new_[32978]_ ,
    \new_[32979]_ , \new_[32980]_ , \new_[32984]_ , \new_[32985]_ ,
    \new_[32988]_ , \new_[32991]_ , \new_[32992]_ , \new_[32993]_ ,
    \new_[32996]_ , \new_[32999]_ , \new_[33000]_ , \new_[33003]_ ,
    \new_[33006]_ , \new_[33007]_ , \new_[33008]_ , \new_[33012]_ ,
    \new_[33013]_ , \new_[33016]_ , \new_[33019]_ , \new_[33020]_ ,
    \new_[33021]_ , \new_[33024]_ , \new_[33027]_ , \new_[33028]_ ,
    \new_[33031]_ , \new_[33034]_ , \new_[33035]_ , \new_[33036]_ ,
    \new_[33040]_ , \new_[33041]_ , \new_[33044]_ , \new_[33047]_ ,
    \new_[33048]_ , \new_[33049]_ , \new_[33052]_ , \new_[33055]_ ,
    \new_[33056]_ , \new_[33059]_ , \new_[33062]_ , \new_[33063]_ ,
    \new_[33064]_ , \new_[33068]_ , \new_[33069]_ , \new_[33072]_ ,
    \new_[33075]_ , \new_[33076]_ , \new_[33077]_ , \new_[33080]_ ,
    \new_[33083]_ , \new_[33084]_ , \new_[33087]_ , \new_[33090]_ ,
    \new_[33091]_ , \new_[33092]_ , \new_[33096]_ , \new_[33097]_ ,
    \new_[33100]_ , \new_[33103]_ , \new_[33104]_ , \new_[33105]_ ,
    \new_[33108]_ , \new_[33111]_ , \new_[33112]_ , \new_[33115]_ ,
    \new_[33118]_ , \new_[33119]_ , \new_[33120]_ , \new_[33124]_ ,
    \new_[33125]_ , \new_[33128]_ , \new_[33131]_ , \new_[33132]_ ,
    \new_[33133]_ , \new_[33136]_ , \new_[33139]_ , \new_[33140]_ ,
    \new_[33143]_ , \new_[33146]_ , \new_[33147]_ , \new_[33148]_ ,
    \new_[33152]_ , \new_[33153]_ , \new_[33156]_ , \new_[33159]_ ,
    \new_[33160]_ , \new_[33161]_ , \new_[33164]_ , \new_[33167]_ ,
    \new_[33168]_ , \new_[33171]_ , \new_[33174]_ , \new_[33175]_ ,
    \new_[33176]_ , \new_[33180]_ , \new_[33181]_ , \new_[33184]_ ,
    \new_[33187]_ , \new_[33188]_ , \new_[33189]_ , \new_[33192]_ ,
    \new_[33195]_ , \new_[33196]_ , \new_[33199]_ , \new_[33202]_ ,
    \new_[33203]_ , \new_[33204]_ , \new_[33208]_ , \new_[33209]_ ,
    \new_[33212]_ , \new_[33215]_ , \new_[33216]_ , \new_[33217]_ ,
    \new_[33220]_ , \new_[33223]_ , \new_[33224]_ , \new_[33227]_ ,
    \new_[33230]_ , \new_[33231]_ , \new_[33232]_ , \new_[33236]_ ,
    \new_[33237]_ , \new_[33240]_ , \new_[33243]_ , \new_[33244]_ ,
    \new_[33245]_ , \new_[33248]_ , \new_[33251]_ , \new_[33252]_ ,
    \new_[33255]_ , \new_[33258]_ , \new_[33259]_ , \new_[33260]_ ,
    \new_[33264]_ , \new_[33265]_ , \new_[33268]_ , \new_[33271]_ ,
    \new_[33272]_ , \new_[33273]_ , \new_[33276]_ , \new_[33279]_ ,
    \new_[33280]_ , \new_[33283]_ , \new_[33286]_ , \new_[33287]_ ,
    \new_[33288]_ , \new_[33292]_ , \new_[33293]_ , \new_[33296]_ ,
    \new_[33299]_ , \new_[33300]_ , \new_[33301]_ , \new_[33304]_ ,
    \new_[33307]_ , \new_[33308]_ , \new_[33311]_ , \new_[33314]_ ,
    \new_[33315]_ , \new_[33316]_ , \new_[33320]_ , \new_[33321]_ ,
    \new_[33324]_ , \new_[33327]_ , \new_[33328]_ , \new_[33329]_ ,
    \new_[33332]_ , \new_[33335]_ , \new_[33336]_ , \new_[33339]_ ,
    \new_[33342]_ , \new_[33343]_ , \new_[33344]_ , \new_[33348]_ ,
    \new_[33349]_ , \new_[33352]_ , \new_[33355]_ , \new_[33356]_ ,
    \new_[33357]_ , \new_[33360]_ , \new_[33363]_ , \new_[33364]_ ,
    \new_[33367]_ , \new_[33370]_ , \new_[33371]_ , \new_[33372]_ ,
    \new_[33376]_ , \new_[33377]_ , \new_[33380]_ , \new_[33383]_ ,
    \new_[33384]_ , \new_[33385]_ , \new_[33388]_ , \new_[33391]_ ,
    \new_[33392]_ , \new_[33395]_ , \new_[33398]_ , \new_[33399]_ ,
    \new_[33400]_ , \new_[33404]_ , \new_[33405]_ , \new_[33408]_ ,
    \new_[33411]_ , \new_[33412]_ , \new_[33413]_ , \new_[33416]_ ,
    \new_[33419]_ , \new_[33420]_ , \new_[33423]_ , \new_[33426]_ ,
    \new_[33427]_ , \new_[33428]_ , \new_[33432]_ , \new_[33433]_ ,
    \new_[33436]_ , \new_[33439]_ , \new_[33440]_ , \new_[33441]_ ,
    \new_[33444]_ , \new_[33447]_ , \new_[33448]_ , \new_[33451]_ ,
    \new_[33454]_ , \new_[33455]_ , \new_[33456]_ , \new_[33460]_ ,
    \new_[33461]_ , \new_[33464]_ , \new_[33467]_ , \new_[33468]_ ,
    \new_[33469]_ , \new_[33472]_ , \new_[33475]_ , \new_[33476]_ ,
    \new_[33479]_ , \new_[33482]_ , \new_[33483]_ , \new_[33484]_ ,
    \new_[33488]_ , \new_[33489]_ , \new_[33492]_ , \new_[33495]_ ,
    \new_[33496]_ , \new_[33497]_ , \new_[33500]_ , \new_[33503]_ ,
    \new_[33504]_ , \new_[33507]_ , \new_[33510]_ , \new_[33511]_ ,
    \new_[33512]_ , \new_[33516]_ , \new_[33517]_ , \new_[33520]_ ,
    \new_[33523]_ , \new_[33524]_ , \new_[33525]_ , \new_[33528]_ ,
    \new_[33531]_ , \new_[33532]_ , \new_[33535]_ , \new_[33538]_ ,
    \new_[33539]_ , \new_[33540]_ , \new_[33544]_ , \new_[33545]_ ,
    \new_[33548]_ , \new_[33551]_ , \new_[33552]_ , \new_[33553]_ ,
    \new_[33556]_ , \new_[33559]_ , \new_[33560]_ , \new_[33563]_ ,
    \new_[33566]_ , \new_[33567]_ , \new_[33568]_ , \new_[33572]_ ,
    \new_[33573]_ , \new_[33576]_ , \new_[33579]_ , \new_[33580]_ ,
    \new_[33581]_ , \new_[33584]_ , \new_[33587]_ , \new_[33588]_ ,
    \new_[33591]_ , \new_[33594]_ , \new_[33595]_ , \new_[33596]_ ,
    \new_[33600]_ , \new_[33601]_ , \new_[33604]_ , \new_[33607]_ ,
    \new_[33608]_ , \new_[33609]_ , \new_[33612]_ , \new_[33615]_ ,
    \new_[33616]_ , \new_[33619]_ , \new_[33622]_ , \new_[33623]_ ,
    \new_[33624]_ , \new_[33628]_ , \new_[33629]_ , \new_[33632]_ ,
    \new_[33635]_ , \new_[33636]_ , \new_[33637]_ , \new_[33640]_ ,
    \new_[33643]_ , \new_[33644]_ , \new_[33647]_ , \new_[33650]_ ,
    \new_[33651]_ , \new_[33652]_ , \new_[33656]_ , \new_[33657]_ ,
    \new_[33660]_ , \new_[33663]_ , \new_[33664]_ , \new_[33665]_ ,
    \new_[33668]_ , \new_[33671]_ , \new_[33672]_ , \new_[33675]_ ,
    \new_[33678]_ , \new_[33679]_ , \new_[33680]_ , \new_[33684]_ ,
    \new_[33685]_ , \new_[33688]_ , \new_[33691]_ , \new_[33692]_ ,
    \new_[33693]_ , \new_[33696]_ , \new_[33699]_ , \new_[33700]_ ,
    \new_[33703]_ , \new_[33706]_ , \new_[33707]_ , \new_[33708]_ ,
    \new_[33712]_ , \new_[33713]_ , \new_[33716]_ , \new_[33719]_ ,
    \new_[33720]_ , \new_[33721]_ , \new_[33724]_ , \new_[33727]_ ,
    \new_[33728]_ , \new_[33731]_ , \new_[33734]_ , \new_[33735]_ ,
    \new_[33736]_ , \new_[33740]_ , \new_[33741]_ , \new_[33744]_ ,
    \new_[33747]_ , \new_[33748]_ , \new_[33749]_ , \new_[33752]_ ,
    \new_[33755]_ , \new_[33756]_ , \new_[33759]_ , \new_[33762]_ ,
    \new_[33763]_ , \new_[33764]_ , \new_[33768]_ , \new_[33769]_ ,
    \new_[33772]_ , \new_[33775]_ , \new_[33776]_ , \new_[33777]_ ,
    \new_[33780]_ , \new_[33783]_ , \new_[33784]_ , \new_[33787]_ ,
    \new_[33790]_ , \new_[33791]_ , \new_[33792]_ , \new_[33796]_ ,
    \new_[33797]_ , \new_[33800]_ , \new_[33803]_ , \new_[33804]_ ,
    \new_[33805]_ , \new_[33808]_ , \new_[33811]_ , \new_[33812]_ ,
    \new_[33815]_ , \new_[33818]_ , \new_[33819]_ , \new_[33820]_ ,
    \new_[33824]_ , \new_[33825]_ , \new_[33828]_ , \new_[33831]_ ,
    \new_[33832]_ , \new_[33833]_ , \new_[33836]_ , \new_[33839]_ ,
    \new_[33840]_ , \new_[33843]_ , \new_[33846]_ , \new_[33847]_ ,
    \new_[33848]_ , \new_[33852]_ , \new_[33853]_ , \new_[33856]_ ,
    \new_[33859]_ , \new_[33860]_ , \new_[33861]_ , \new_[33864]_ ,
    \new_[33867]_ , \new_[33868]_ , \new_[33871]_ , \new_[33874]_ ,
    \new_[33875]_ , \new_[33876]_ , \new_[33880]_ , \new_[33881]_ ,
    \new_[33884]_ , \new_[33887]_ , \new_[33888]_ , \new_[33889]_ ,
    \new_[33892]_ , \new_[33895]_ , \new_[33896]_ , \new_[33899]_ ,
    \new_[33902]_ , \new_[33903]_ , \new_[33904]_ , \new_[33908]_ ,
    \new_[33909]_ , \new_[33912]_ , \new_[33915]_ , \new_[33916]_ ,
    \new_[33917]_ , \new_[33920]_ , \new_[33923]_ , \new_[33924]_ ,
    \new_[33927]_ , \new_[33930]_ , \new_[33931]_ , \new_[33932]_ ,
    \new_[33936]_ , \new_[33937]_ , \new_[33940]_ , \new_[33943]_ ,
    \new_[33944]_ , \new_[33945]_ , \new_[33948]_ , \new_[33951]_ ,
    \new_[33952]_ , \new_[33955]_ , \new_[33958]_ , \new_[33959]_ ,
    \new_[33960]_ , \new_[33964]_ , \new_[33965]_ , \new_[33968]_ ,
    \new_[33971]_ , \new_[33972]_ , \new_[33973]_ , \new_[33976]_ ,
    \new_[33979]_ , \new_[33980]_ , \new_[33983]_ , \new_[33986]_ ,
    \new_[33987]_ , \new_[33988]_ , \new_[33992]_ , \new_[33993]_ ,
    \new_[33996]_ , \new_[33999]_ , \new_[34000]_ , \new_[34001]_ ,
    \new_[34004]_ , \new_[34007]_ , \new_[34008]_ , \new_[34011]_ ,
    \new_[34014]_ , \new_[34015]_ , \new_[34016]_ , \new_[34020]_ ,
    \new_[34021]_ , \new_[34024]_ , \new_[34027]_ , \new_[34028]_ ,
    \new_[34029]_ , \new_[34032]_ , \new_[34035]_ , \new_[34036]_ ,
    \new_[34039]_ , \new_[34042]_ , \new_[34043]_ , \new_[34044]_ ,
    \new_[34048]_ , \new_[34049]_ , \new_[34052]_ , \new_[34055]_ ,
    \new_[34056]_ , \new_[34057]_ , \new_[34060]_ , \new_[34063]_ ,
    \new_[34064]_ , \new_[34067]_ , \new_[34070]_ , \new_[34071]_ ,
    \new_[34072]_ , \new_[34076]_ , \new_[34077]_ , \new_[34080]_ ,
    \new_[34083]_ , \new_[34084]_ , \new_[34085]_ , \new_[34088]_ ,
    \new_[34091]_ , \new_[34092]_ , \new_[34095]_ , \new_[34098]_ ,
    \new_[34099]_ , \new_[34100]_ , \new_[34104]_ , \new_[34105]_ ,
    \new_[34108]_ , \new_[34111]_ , \new_[34112]_ , \new_[34113]_ ,
    \new_[34116]_ , \new_[34119]_ , \new_[34120]_ , \new_[34123]_ ,
    \new_[34126]_ , \new_[34127]_ , \new_[34128]_ , \new_[34132]_ ,
    \new_[34133]_ , \new_[34136]_ , \new_[34139]_ , \new_[34140]_ ,
    \new_[34141]_ , \new_[34144]_ , \new_[34147]_ , \new_[34148]_ ,
    \new_[34151]_ , \new_[34154]_ , \new_[34155]_ , \new_[34156]_ ,
    \new_[34160]_ , \new_[34161]_ , \new_[34164]_ , \new_[34167]_ ,
    \new_[34168]_ , \new_[34169]_ , \new_[34172]_ , \new_[34175]_ ,
    \new_[34176]_ , \new_[34179]_ , \new_[34182]_ , \new_[34183]_ ,
    \new_[34184]_ , \new_[34188]_ , \new_[34189]_ , \new_[34192]_ ,
    \new_[34195]_ , \new_[34196]_ , \new_[34197]_ , \new_[34200]_ ,
    \new_[34203]_ , \new_[34204]_ , \new_[34207]_ , \new_[34210]_ ,
    \new_[34211]_ , \new_[34212]_ , \new_[34216]_ , \new_[34217]_ ,
    \new_[34220]_ , \new_[34223]_ , \new_[34224]_ , \new_[34225]_ ,
    \new_[34228]_ , \new_[34231]_ , \new_[34232]_ , \new_[34235]_ ,
    \new_[34238]_ , \new_[34239]_ , \new_[34240]_ , \new_[34244]_ ,
    \new_[34245]_ , \new_[34248]_ , \new_[34251]_ , \new_[34252]_ ,
    \new_[34253]_ , \new_[34256]_ , \new_[34259]_ , \new_[34260]_ ,
    \new_[34263]_ , \new_[34266]_ , \new_[34267]_ , \new_[34268]_ ,
    \new_[34272]_ , \new_[34273]_ , \new_[34276]_ , \new_[34279]_ ,
    \new_[34280]_ , \new_[34281]_ , \new_[34284]_ , \new_[34287]_ ,
    \new_[34288]_ , \new_[34291]_ , \new_[34294]_ , \new_[34295]_ ,
    \new_[34296]_ , \new_[34300]_ , \new_[34301]_ , \new_[34304]_ ,
    \new_[34307]_ , \new_[34308]_ , \new_[34309]_ , \new_[34312]_ ,
    \new_[34315]_ , \new_[34316]_ , \new_[34319]_ , \new_[34322]_ ,
    \new_[34323]_ , \new_[34324]_ , \new_[34328]_ , \new_[34329]_ ,
    \new_[34332]_ , \new_[34335]_ , \new_[34336]_ , \new_[34337]_ ,
    \new_[34340]_ , \new_[34343]_ , \new_[34344]_ , \new_[34347]_ ,
    \new_[34350]_ , \new_[34351]_ , \new_[34352]_ , \new_[34356]_ ,
    \new_[34357]_ , \new_[34360]_ , \new_[34363]_ , \new_[34364]_ ,
    \new_[34365]_ , \new_[34368]_ , \new_[34371]_ , \new_[34372]_ ,
    \new_[34375]_ , \new_[34378]_ , \new_[34379]_ , \new_[34380]_ ,
    \new_[34384]_ , \new_[34385]_ , \new_[34388]_ , \new_[34391]_ ,
    \new_[34392]_ , \new_[34393]_ , \new_[34396]_ , \new_[34399]_ ,
    \new_[34400]_ , \new_[34403]_ , \new_[34406]_ , \new_[34407]_ ,
    \new_[34408]_ , \new_[34412]_ , \new_[34413]_ , \new_[34416]_ ,
    \new_[34419]_ , \new_[34420]_ , \new_[34421]_ , \new_[34424]_ ,
    \new_[34427]_ , \new_[34428]_ , \new_[34431]_ , \new_[34434]_ ,
    \new_[34435]_ , \new_[34436]_ , \new_[34440]_ , \new_[34441]_ ,
    \new_[34444]_ , \new_[34447]_ , \new_[34448]_ , \new_[34449]_ ,
    \new_[34452]_ , \new_[34455]_ , \new_[34456]_ , \new_[34459]_ ,
    \new_[34462]_ , \new_[34463]_ , \new_[34464]_ , \new_[34468]_ ,
    \new_[34469]_ , \new_[34472]_ , \new_[34475]_ , \new_[34476]_ ,
    \new_[34477]_ , \new_[34480]_ , \new_[34483]_ , \new_[34484]_ ,
    \new_[34487]_ , \new_[34490]_ , \new_[34491]_ , \new_[34492]_ ,
    \new_[34496]_ , \new_[34497]_ , \new_[34500]_ , \new_[34503]_ ,
    \new_[34504]_ , \new_[34505]_ , \new_[34508]_ , \new_[34511]_ ,
    \new_[34512]_ , \new_[34515]_ , \new_[34518]_ , \new_[34519]_ ,
    \new_[34520]_ , \new_[34524]_ , \new_[34525]_ , \new_[34528]_ ,
    \new_[34531]_ , \new_[34532]_ , \new_[34533]_ , \new_[34536]_ ,
    \new_[34539]_ , \new_[34540]_ , \new_[34543]_ , \new_[34546]_ ,
    \new_[34547]_ , \new_[34548]_ , \new_[34552]_ , \new_[34553]_ ,
    \new_[34556]_ , \new_[34559]_ , \new_[34560]_ , \new_[34561]_ ,
    \new_[34564]_ , \new_[34567]_ , \new_[34568]_ , \new_[34571]_ ,
    \new_[34574]_ , \new_[34575]_ , \new_[34576]_ , \new_[34580]_ ,
    \new_[34581]_ , \new_[34584]_ , \new_[34587]_ , \new_[34588]_ ,
    \new_[34589]_ , \new_[34592]_ , \new_[34595]_ , \new_[34596]_ ,
    \new_[34599]_ , \new_[34602]_ , \new_[34603]_ , \new_[34604]_ ,
    \new_[34608]_ , \new_[34609]_ , \new_[34612]_ , \new_[34615]_ ,
    \new_[34616]_ , \new_[34617]_ , \new_[34620]_ , \new_[34623]_ ,
    \new_[34624]_ , \new_[34627]_ , \new_[34630]_ , \new_[34631]_ ,
    \new_[34632]_ , \new_[34636]_ , \new_[34637]_ , \new_[34640]_ ,
    \new_[34643]_ , \new_[34644]_ , \new_[34645]_ , \new_[34648]_ ,
    \new_[34651]_ , \new_[34652]_ , \new_[34655]_ , \new_[34658]_ ,
    \new_[34659]_ , \new_[34660]_ , \new_[34664]_ , \new_[34665]_ ,
    \new_[34668]_ , \new_[34671]_ , \new_[34672]_ , \new_[34673]_ ,
    \new_[34676]_ , \new_[34679]_ , \new_[34680]_ , \new_[34683]_ ,
    \new_[34686]_ , \new_[34687]_ , \new_[34688]_ , \new_[34692]_ ,
    \new_[34693]_ , \new_[34696]_ , \new_[34699]_ , \new_[34700]_ ,
    \new_[34701]_ , \new_[34704]_ , \new_[34707]_ , \new_[34708]_ ,
    \new_[34711]_ , \new_[34714]_ , \new_[34715]_ , \new_[34716]_ ,
    \new_[34720]_ , \new_[34721]_ , \new_[34724]_ , \new_[34727]_ ,
    \new_[34728]_ , \new_[34729]_ , \new_[34732]_ , \new_[34735]_ ,
    \new_[34736]_ , \new_[34739]_ , \new_[34742]_ , \new_[34743]_ ,
    \new_[34744]_ , \new_[34748]_ , \new_[34749]_ , \new_[34752]_ ,
    \new_[34755]_ , \new_[34756]_ , \new_[34757]_ , \new_[34760]_ ,
    \new_[34763]_ , \new_[34764]_ , \new_[34767]_ , \new_[34770]_ ,
    \new_[34771]_ , \new_[34772]_ , \new_[34776]_ , \new_[34777]_ ,
    \new_[34780]_ , \new_[34783]_ , \new_[34784]_ , \new_[34785]_ ,
    \new_[34788]_ , \new_[34791]_ , \new_[34792]_ , \new_[34795]_ ,
    \new_[34798]_ , \new_[34799]_ , \new_[34800]_ , \new_[34804]_ ,
    \new_[34805]_ , \new_[34808]_ , \new_[34811]_ , \new_[34812]_ ,
    \new_[34813]_ , \new_[34816]_ , \new_[34819]_ , \new_[34820]_ ,
    \new_[34823]_ , \new_[34826]_ , \new_[34827]_ , \new_[34828]_ ,
    \new_[34832]_ , \new_[34833]_ , \new_[34836]_ , \new_[34839]_ ,
    \new_[34840]_ , \new_[34841]_ , \new_[34844]_ , \new_[34847]_ ,
    \new_[34848]_ , \new_[34851]_ , \new_[34854]_ , \new_[34855]_ ,
    \new_[34856]_ , \new_[34860]_ , \new_[34861]_ , \new_[34864]_ ,
    \new_[34867]_ , \new_[34868]_ , \new_[34869]_ , \new_[34872]_ ,
    \new_[34875]_ , \new_[34876]_ , \new_[34879]_ , \new_[34882]_ ,
    \new_[34883]_ , \new_[34884]_ , \new_[34888]_ , \new_[34889]_ ,
    \new_[34892]_ , \new_[34895]_ , \new_[34896]_ , \new_[34897]_ ,
    \new_[34900]_ , \new_[34903]_ , \new_[34904]_ , \new_[34907]_ ,
    \new_[34910]_ , \new_[34911]_ , \new_[34912]_ , \new_[34916]_ ,
    \new_[34917]_ , \new_[34920]_ , \new_[34923]_ , \new_[34924]_ ,
    \new_[34925]_ , \new_[34928]_ , \new_[34931]_ , \new_[34932]_ ,
    \new_[34935]_ , \new_[34938]_ , \new_[34939]_ , \new_[34940]_ ,
    \new_[34944]_ , \new_[34945]_ , \new_[34948]_ , \new_[34951]_ ,
    \new_[34952]_ , \new_[34953]_ , \new_[34956]_ , \new_[34959]_ ,
    \new_[34960]_ , \new_[34963]_ , \new_[34966]_ , \new_[34967]_ ,
    \new_[34968]_ , \new_[34972]_ , \new_[34973]_ , \new_[34976]_ ,
    \new_[34979]_ , \new_[34980]_ , \new_[34981]_ , \new_[34984]_ ,
    \new_[34987]_ , \new_[34988]_ , \new_[34991]_ , \new_[34994]_ ,
    \new_[34995]_ , \new_[34996]_ , \new_[35000]_ , \new_[35001]_ ,
    \new_[35004]_ , \new_[35007]_ , \new_[35008]_ , \new_[35009]_ ,
    \new_[35012]_ , \new_[35015]_ , \new_[35016]_ , \new_[35019]_ ,
    \new_[35022]_ , \new_[35023]_ , \new_[35024]_ , \new_[35028]_ ,
    \new_[35029]_ , \new_[35032]_ , \new_[35035]_ , \new_[35036]_ ,
    \new_[35037]_ , \new_[35040]_ , \new_[35043]_ , \new_[35044]_ ,
    \new_[35047]_ , \new_[35050]_ , \new_[35051]_ , \new_[35052]_ ,
    \new_[35056]_ , \new_[35057]_ , \new_[35060]_ , \new_[35063]_ ,
    \new_[35064]_ , \new_[35065]_ , \new_[35068]_ , \new_[35071]_ ,
    \new_[35072]_ , \new_[35075]_ , \new_[35078]_ , \new_[35079]_ ,
    \new_[35080]_ , \new_[35084]_ , \new_[35085]_ , \new_[35088]_ ,
    \new_[35091]_ , \new_[35092]_ , \new_[35093]_ , \new_[35096]_ ,
    \new_[35099]_ , \new_[35100]_ , \new_[35103]_ , \new_[35106]_ ,
    \new_[35107]_ , \new_[35108]_ , \new_[35112]_ , \new_[35113]_ ,
    \new_[35116]_ , \new_[35119]_ , \new_[35120]_ , \new_[35121]_ ,
    \new_[35124]_ , \new_[35127]_ , \new_[35128]_ , \new_[35131]_ ,
    \new_[35134]_ , \new_[35135]_ , \new_[35136]_ , \new_[35140]_ ,
    \new_[35141]_ , \new_[35144]_ , \new_[35147]_ , \new_[35148]_ ,
    \new_[35149]_ , \new_[35152]_ , \new_[35155]_ , \new_[35156]_ ,
    \new_[35159]_ , \new_[35162]_ , \new_[35163]_ , \new_[35164]_ ,
    \new_[35168]_ , \new_[35169]_ , \new_[35172]_ , \new_[35175]_ ,
    \new_[35176]_ , \new_[35177]_ , \new_[35180]_ , \new_[35183]_ ,
    \new_[35184]_ , \new_[35187]_ , \new_[35190]_ , \new_[35191]_ ,
    \new_[35192]_ , \new_[35196]_ , \new_[35197]_ , \new_[35200]_ ,
    \new_[35203]_ , \new_[35204]_ , \new_[35205]_ , \new_[35208]_ ,
    \new_[35211]_ , \new_[35212]_ , \new_[35215]_ , \new_[35218]_ ,
    \new_[35219]_ , \new_[35220]_ , \new_[35224]_ , \new_[35225]_ ,
    \new_[35228]_ , \new_[35231]_ , \new_[35232]_ , \new_[35233]_ ,
    \new_[35236]_ , \new_[35239]_ , \new_[35240]_ , \new_[35243]_ ,
    \new_[35246]_ , \new_[35247]_ , \new_[35248]_ , \new_[35252]_ ,
    \new_[35253]_ , \new_[35256]_ , \new_[35259]_ , \new_[35260]_ ,
    \new_[35261]_ , \new_[35264]_ , \new_[35267]_ , \new_[35268]_ ,
    \new_[35271]_ , \new_[35274]_ , \new_[35275]_ , \new_[35276]_ ,
    \new_[35280]_ , \new_[35281]_ , \new_[35284]_ , \new_[35287]_ ,
    \new_[35288]_ , \new_[35289]_ , \new_[35292]_ , \new_[35295]_ ,
    \new_[35296]_ , \new_[35299]_ , \new_[35302]_ , \new_[35303]_ ,
    \new_[35304]_ , \new_[35308]_ , \new_[35309]_ , \new_[35312]_ ,
    \new_[35315]_ , \new_[35316]_ , \new_[35317]_ , \new_[35320]_ ,
    \new_[35323]_ , \new_[35324]_ , \new_[35327]_ , \new_[35330]_ ,
    \new_[35331]_ , \new_[35332]_ , \new_[35336]_ , \new_[35337]_ ,
    \new_[35340]_ , \new_[35343]_ , \new_[35344]_ , \new_[35345]_ ,
    \new_[35348]_ , \new_[35351]_ , \new_[35352]_ , \new_[35355]_ ,
    \new_[35358]_ , \new_[35359]_ , \new_[35360]_ , \new_[35364]_ ,
    \new_[35365]_ , \new_[35368]_ , \new_[35371]_ , \new_[35372]_ ,
    \new_[35373]_ , \new_[35376]_ , \new_[35379]_ , \new_[35380]_ ,
    \new_[35383]_ , \new_[35386]_ , \new_[35387]_ , \new_[35388]_ ,
    \new_[35392]_ , \new_[35393]_ , \new_[35396]_ , \new_[35399]_ ,
    \new_[35400]_ , \new_[35401]_ , \new_[35404]_ , \new_[35407]_ ,
    \new_[35408]_ , \new_[35411]_ , \new_[35414]_ , \new_[35415]_ ,
    \new_[35416]_ , \new_[35420]_ , \new_[35421]_ , \new_[35424]_ ,
    \new_[35427]_ , \new_[35428]_ , \new_[35429]_ , \new_[35432]_ ,
    \new_[35435]_ , \new_[35436]_ , \new_[35439]_ , \new_[35442]_ ,
    \new_[35443]_ , \new_[35444]_ , \new_[35448]_ , \new_[35449]_ ,
    \new_[35452]_ , \new_[35455]_ , \new_[35456]_ , \new_[35457]_ ,
    \new_[35460]_ , \new_[35463]_ , \new_[35464]_ , \new_[35467]_ ,
    \new_[35470]_ , \new_[35471]_ , \new_[35472]_ , \new_[35476]_ ,
    \new_[35477]_ , \new_[35480]_ , \new_[35483]_ , \new_[35484]_ ,
    \new_[35485]_ , \new_[35488]_ , \new_[35491]_ , \new_[35492]_ ,
    \new_[35495]_ , \new_[35498]_ , \new_[35499]_ , \new_[35500]_ ,
    \new_[35504]_ , \new_[35505]_ , \new_[35508]_ , \new_[35511]_ ,
    \new_[35512]_ , \new_[35513]_ , \new_[35516]_ , \new_[35519]_ ,
    \new_[35520]_ , \new_[35523]_ , \new_[35526]_ , \new_[35527]_ ,
    \new_[35528]_ , \new_[35532]_ , \new_[35533]_ , \new_[35536]_ ,
    \new_[35539]_ , \new_[35540]_ , \new_[35541]_ , \new_[35544]_ ,
    \new_[35547]_ , \new_[35548]_ , \new_[35551]_ , \new_[35554]_ ,
    \new_[35555]_ , \new_[35556]_ , \new_[35560]_ , \new_[35561]_ ,
    \new_[35564]_ , \new_[35567]_ , \new_[35568]_ , \new_[35569]_ ,
    \new_[35572]_ , \new_[35575]_ , \new_[35576]_ , \new_[35579]_ ,
    \new_[35582]_ , \new_[35583]_ , \new_[35584]_ , \new_[35588]_ ,
    \new_[35589]_ , \new_[35592]_ , \new_[35595]_ , \new_[35596]_ ,
    \new_[35597]_ , \new_[35600]_ , \new_[35603]_ , \new_[35604]_ ,
    \new_[35607]_ , \new_[35610]_ , \new_[35611]_ , \new_[35612]_ ,
    \new_[35616]_ , \new_[35617]_ , \new_[35620]_ , \new_[35623]_ ,
    \new_[35624]_ , \new_[35625]_ , \new_[35628]_ , \new_[35631]_ ,
    \new_[35632]_ , \new_[35635]_ , \new_[35638]_ , \new_[35639]_ ,
    \new_[35640]_ , \new_[35644]_ , \new_[35645]_ , \new_[35648]_ ,
    \new_[35651]_ , \new_[35652]_ , \new_[35653]_ , \new_[35656]_ ,
    \new_[35659]_ , \new_[35660]_ , \new_[35663]_ , \new_[35666]_ ,
    \new_[35667]_ , \new_[35668]_ , \new_[35672]_ , \new_[35673]_ ,
    \new_[35676]_ , \new_[35679]_ , \new_[35680]_ , \new_[35681]_ ,
    \new_[35684]_ , \new_[35687]_ , \new_[35688]_ , \new_[35691]_ ,
    \new_[35694]_ , \new_[35695]_ , \new_[35696]_ , \new_[35700]_ ,
    \new_[35701]_ , \new_[35704]_ , \new_[35707]_ , \new_[35708]_ ,
    \new_[35709]_ , \new_[35712]_ , \new_[35715]_ , \new_[35716]_ ,
    \new_[35719]_ , \new_[35722]_ , \new_[35723]_ , \new_[35724]_ ,
    \new_[35728]_ , \new_[35729]_ , \new_[35732]_ , \new_[35735]_ ,
    \new_[35736]_ , \new_[35737]_ , \new_[35740]_ , \new_[35743]_ ,
    \new_[35744]_ , \new_[35747]_ , \new_[35750]_ , \new_[35751]_ ,
    \new_[35752]_ , \new_[35756]_ , \new_[35757]_ , \new_[35760]_ ,
    \new_[35763]_ , \new_[35764]_ , \new_[35765]_ , \new_[35768]_ ,
    \new_[35771]_ , \new_[35772]_ , \new_[35775]_ , \new_[35778]_ ,
    \new_[35779]_ , \new_[35780]_ , \new_[35784]_ , \new_[35785]_ ,
    \new_[35788]_ , \new_[35791]_ , \new_[35792]_ , \new_[35793]_ ,
    \new_[35796]_ , \new_[35799]_ , \new_[35800]_ , \new_[35803]_ ,
    \new_[35806]_ , \new_[35807]_ , \new_[35808]_ , \new_[35812]_ ,
    \new_[35813]_ , \new_[35816]_ , \new_[35819]_ , \new_[35820]_ ,
    \new_[35821]_ , \new_[35824]_ , \new_[35827]_ , \new_[35828]_ ,
    \new_[35831]_ , \new_[35834]_ , \new_[35835]_ , \new_[35836]_ ,
    \new_[35840]_ , \new_[35841]_ , \new_[35844]_ , \new_[35847]_ ,
    \new_[35848]_ , \new_[35849]_ , \new_[35852]_ , \new_[35855]_ ,
    \new_[35856]_ , \new_[35859]_ , \new_[35862]_ , \new_[35863]_ ,
    \new_[35864]_ , \new_[35868]_ , \new_[35869]_ , \new_[35872]_ ,
    \new_[35875]_ , \new_[35876]_ , \new_[35877]_ , \new_[35880]_ ,
    \new_[35883]_ , \new_[35884]_ , \new_[35887]_ , \new_[35890]_ ,
    \new_[35891]_ , \new_[35892]_ , \new_[35896]_ , \new_[35897]_ ,
    \new_[35900]_ , \new_[35903]_ , \new_[35904]_ , \new_[35905]_ ,
    \new_[35908]_ , \new_[35911]_ , \new_[35912]_ , \new_[35915]_ ,
    \new_[35918]_ , \new_[35919]_ , \new_[35920]_ , \new_[35924]_ ,
    \new_[35925]_ , \new_[35928]_ , \new_[35931]_ , \new_[35932]_ ,
    \new_[35933]_ , \new_[35936]_ , \new_[35939]_ , \new_[35940]_ ,
    \new_[35943]_ , \new_[35946]_ , \new_[35947]_ , \new_[35948]_ ,
    \new_[35952]_ , \new_[35953]_ , \new_[35956]_ , \new_[35959]_ ,
    \new_[35960]_ , \new_[35961]_ , \new_[35964]_ , \new_[35967]_ ,
    \new_[35968]_ , \new_[35971]_ , \new_[35974]_ , \new_[35975]_ ,
    \new_[35976]_ , \new_[35980]_ , \new_[35981]_ , \new_[35984]_ ,
    \new_[35987]_ , \new_[35988]_ , \new_[35989]_ , \new_[35992]_ ,
    \new_[35995]_ , \new_[35996]_ , \new_[35999]_ , \new_[36002]_ ,
    \new_[36003]_ , \new_[36004]_ , \new_[36008]_ , \new_[36009]_ ,
    \new_[36012]_ , \new_[36015]_ , \new_[36016]_ , \new_[36017]_ ,
    \new_[36020]_ , \new_[36023]_ , \new_[36024]_ , \new_[36027]_ ,
    \new_[36030]_ , \new_[36031]_ , \new_[36032]_ , \new_[36036]_ ,
    \new_[36037]_ , \new_[36040]_ , \new_[36043]_ , \new_[36044]_ ,
    \new_[36045]_ , \new_[36048]_ , \new_[36051]_ , \new_[36052]_ ,
    \new_[36055]_ , \new_[36058]_ , \new_[36059]_ , \new_[36060]_ ,
    \new_[36064]_ , \new_[36065]_ , \new_[36068]_ , \new_[36071]_ ,
    \new_[36072]_ , \new_[36073]_ , \new_[36076]_ , \new_[36079]_ ,
    \new_[36080]_ , \new_[36083]_ , \new_[36086]_ , \new_[36087]_ ,
    \new_[36088]_ , \new_[36092]_ , \new_[36093]_ , \new_[36096]_ ,
    \new_[36099]_ , \new_[36100]_ , \new_[36101]_ , \new_[36104]_ ,
    \new_[36107]_ , \new_[36108]_ , \new_[36111]_ , \new_[36114]_ ,
    \new_[36115]_ , \new_[36116]_ , \new_[36120]_ , \new_[36121]_ ,
    \new_[36124]_ , \new_[36127]_ , \new_[36128]_ , \new_[36129]_ ,
    \new_[36132]_ , \new_[36135]_ , \new_[36136]_ , \new_[36139]_ ,
    \new_[36142]_ , \new_[36143]_ , \new_[36144]_ , \new_[36148]_ ,
    \new_[36149]_ , \new_[36152]_ , \new_[36155]_ , \new_[36156]_ ,
    \new_[36157]_ , \new_[36160]_ , \new_[36163]_ , \new_[36164]_ ,
    \new_[36167]_ , \new_[36170]_ , \new_[36171]_ , \new_[36172]_ ,
    \new_[36176]_ , \new_[36177]_ , \new_[36180]_ , \new_[36183]_ ,
    \new_[36184]_ , \new_[36185]_ , \new_[36188]_ , \new_[36191]_ ,
    \new_[36192]_ , \new_[36195]_ , \new_[36198]_ , \new_[36199]_ ,
    \new_[36200]_ , \new_[36204]_ , \new_[36205]_ , \new_[36208]_ ,
    \new_[36211]_ , \new_[36212]_ , \new_[36213]_ , \new_[36216]_ ,
    \new_[36219]_ , \new_[36220]_ , \new_[36223]_ , \new_[36226]_ ,
    \new_[36227]_ , \new_[36228]_ , \new_[36232]_ , \new_[36233]_ ,
    \new_[36236]_ , \new_[36239]_ , \new_[36240]_ , \new_[36241]_ ,
    \new_[36244]_ , \new_[36247]_ , \new_[36248]_ , \new_[36251]_ ,
    \new_[36254]_ , \new_[36255]_ , \new_[36256]_ , \new_[36260]_ ,
    \new_[36261]_ , \new_[36264]_ , \new_[36267]_ , \new_[36268]_ ,
    \new_[36269]_ , \new_[36272]_ , \new_[36275]_ , \new_[36276]_ ,
    \new_[36279]_ , \new_[36282]_ , \new_[36283]_ , \new_[36284]_ ,
    \new_[36288]_ , \new_[36289]_ , \new_[36292]_ , \new_[36295]_ ,
    \new_[36296]_ , \new_[36297]_ , \new_[36300]_ , \new_[36303]_ ,
    \new_[36304]_ , \new_[36307]_ , \new_[36310]_ , \new_[36311]_ ,
    \new_[36312]_ , \new_[36316]_ , \new_[36317]_ , \new_[36320]_ ,
    \new_[36323]_ , \new_[36324]_ , \new_[36325]_ , \new_[36328]_ ,
    \new_[36331]_ , \new_[36332]_ , \new_[36335]_ , \new_[36338]_ ,
    \new_[36339]_ , \new_[36340]_ , \new_[36344]_ , \new_[36345]_ ,
    \new_[36348]_ , \new_[36351]_ , \new_[36352]_ , \new_[36353]_ ,
    \new_[36356]_ , \new_[36359]_ , \new_[36360]_ , \new_[36363]_ ,
    \new_[36366]_ , \new_[36367]_ , \new_[36368]_ , \new_[36372]_ ,
    \new_[36373]_ , \new_[36376]_ , \new_[36379]_ , \new_[36380]_ ,
    \new_[36381]_ , \new_[36384]_ , \new_[36387]_ , \new_[36388]_ ,
    \new_[36391]_ , \new_[36394]_ , \new_[36395]_ , \new_[36396]_ ,
    \new_[36400]_ , \new_[36401]_ , \new_[36404]_ , \new_[36407]_ ,
    \new_[36408]_ , \new_[36409]_ , \new_[36412]_ , \new_[36415]_ ,
    \new_[36416]_ , \new_[36419]_ , \new_[36422]_ , \new_[36423]_ ,
    \new_[36424]_ , \new_[36428]_ , \new_[36429]_ , \new_[36432]_ ,
    \new_[36435]_ , \new_[36436]_ , \new_[36437]_ , \new_[36440]_ ,
    \new_[36443]_ , \new_[36444]_ , \new_[36447]_ , \new_[36450]_ ,
    \new_[36451]_ , \new_[36452]_ , \new_[36456]_ , \new_[36457]_ ,
    \new_[36460]_ , \new_[36463]_ , \new_[36464]_ , \new_[36465]_ ,
    \new_[36468]_ , \new_[36471]_ , \new_[36472]_ , \new_[36475]_ ,
    \new_[36478]_ , \new_[36479]_ , \new_[36480]_ , \new_[36484]_ ,
    \new_[36485]_ , \new_[36488]_ , \new_[36491]_ , \new_[36492]_ ,
    \new_[36493]_ , \new_[36496]_ , \new_[36499]_ , \new_[36500]_ ,
    \new_[36503]_ , \new_[36506]_ , \new_[36507]_ , \new_[36508]_ ,
    \new_[36512]_ , \new_[36513]_ , \new_[36516]_ , \new_[36519]_ ,
    \new_[36520]_ , \new_[36521]_ , \new_[36524]_ , \new_[36527]_ ,
    \new_[36528]_ , \new_[36531]_ , \new_[36534]_ , \new_[36535]_ ,
    \new_[36536]_ , \new_[36540]_ , \new_[36541]_ , \new_[36544]_ ,
    \new_[36547]_ , \new_[36548]_ , \new_[36549]_ , \new_[36552]_ ,
    \new_[36555]_ , \new_[36556]_ , \new_[36559]_ , \new_[36562]_ ,
    \new_[36563]_ , \new_[36564]_ , \new_[36568]_ , \new_[36569]_ ,
    \new_[36572]_ , \new_[36575]_ , \new_[36576]_ , \new_[36577]_ ,
    \new_[36580]_ , \new_[36583]_ , \new_[36584]_ , \new_[36587]_ ,
    \new_[36590]_ , \new_[36591]_ , \new_[36592]_ , \new_[36596]_ ,
    \new_[36597]_ , \new_[36600]_ , \new_[36603]_ , \new_[36604]_ ,
    \new_[36605]_ , \new_[36608]_ , \new_[36611]_ , \new_[36612]_ ,
    \new_[36615]_ , \new_[36618]_ , \new_[36619]_ , \new_[36620]_ ,
    \new_[36624]_ , \new_[36625]_ , \new_[36628]_ , \new_[36631]_ ,
    \new_[36632]_ , \new_[36633]_ , \new_[36636]_ , \new_[36639]_ ,
    \new_[36640]_ , \new_[36643]_ , \new_[36646]_ , \new_[36647]_ ,
    \new_[36648]_ , \new_[36652]_ , \new_[36653]_ , \new_[36656]_ ,
    \new_[36659]_ , \new_[36660]_ , \new_[36661]_ , \new_[36664]_ ,
    \new_[36667]_ , \new_[36668]_ , \new_[36671]_ , \new_[36674]_ ,
    \new_[36675]_ , \new_[36676]_ , \new_[36680]_ , \new_[36681]_ ,
    \new_[36684]_ , \new_[36687]_ , \new_[36688]_ , \new_[36689]_ ,
    \new_[36692]_ , \new_[36695]_ , \new_[36696]_ , \new_[36699]_ ,
    \new_[36702]_ , \new_[36703]_ , \new_[36704]_ , \new_[36708]_ ,
    \new_[36709]_ , \new_[36712]_ , \new_[36715]_ , \new_[36716]_ ,
    \new_[36717]_ , \new_[36720]_ , \new_[36723]_ , \new_[36724]_ ,
    \new_[36727]_ , \new_[36730]_ , \new_[36731]_ , \new_[36732]_ ,
    \new_[36736]_ , \new_[36737]_ , \new_[36740]_ , \new_[36743]_ ,
    \new_[36744]_ , \new_[36745]_ , \new_[36748]_ , \new_[36751]_ ,
    \new_[36752]_ , \new_[36755]_ , \new_[36758]_ , \new_[36759]_ ,
    \new_[36760]_ , \new_[36764]_ , \new_[36765]_ , \new_[36768]_ ,
    \new_[36771]_ , \new_[36772]_ , \new_[36773]_ , \new_[36776]_ ,
    \new_[36779]_ , \new_[36780]_ , \new_[36783]_ , \new_[36786]_ ,
    \new_[36787]_ , \new_[36788]_ , \new_[36792]_ , \new_[36793]_ ,
    \new_[36796]_ , \new_[36799]_ , \new_[36800]_ , \new_[36801]_ ,
    \new_[36804]_ , \new_[36807]_ , \new_[36808]_ , \new_[36811]_ ,
    \new_[36814]_ , \new_[36815]_ , \new_[36816]_ , \new_[36820]_ ,
    \new_[36821]_ , \new_[36824]_ , \new_[36827]_ , \new_[36828]_ ,
    \new_[36829]_ , \new_[36832]_ , \new_[36835]_ , \new_[36836]_ ,
    \new_[36839]_ , \new_[36842]_ , \new_[36843]_ , \new_[36844]_ ,
    \new_[36848]_ , \new_[36849]_ , \new_[36852]_ , \new_[36855]_ ,
    \new_[36856]_ , \new_[36857]_ , \new_[36860]_ , \new_[36863]_ ,
    \new_[36864]_ , \new_[36867]_ , \new_[36870]_ , \new_[36871]_ ,
    \new_[36872]_ , \new_[36876]_ , \new_[36877]_ , \new_[36880]_ ,
    \new_[36883]_ , \new_[36884]_ , \new_[36885]_ , \new_[36888]_ ,
    \new_[36891]_ , \new_[36892]_ , \new_[36895]_ , \new_[36898]_ ,
    \new_[36899]_ , \new_[36900]_ , \new_[36904]_ , \new_[36905]_ ,
    \new_[36908]_ , \new_[36911]_ , \new_[36912]_ , \new_[36913]_ ,
    \new_[36916]_ , \new_[36919]_ , \new_[36920]_ , \new_[36923]_ ,
    \new_[36926]_ , \new_[36927]_ , \new_[36928]_ , \new_[36932]_ ,
    \new_[36933]_ , \new_[36936]_ , \new_[36939]_ , \new_[36940]_ ,
    \new_[36941]_ , \new_[36944]_ , \new_[36947]_ , \new_[36948]_ ,
    \new_[36951]_ , \new_[36954]_ , \new_[36955]_ , \new_[36956]_ ,
    \new_[36960]_ , \new_[36961]_ , \new_[36964]_ , \new_[36967]_ ,
    \new_[36968]_ , \new_[36969]_ , \new_[36972]_ , \new_[36975]_ ,
    \new_[36976]_ , \new_[36979]_ , \new_[36982]_ , \new_[36983]_ ,
    \new_[36984]_ , \new_[36988]_ , \new_[36989]_ , \new_[36992]_ ,
    \new_[36995]_ , \new_[36996]_ , \new_[36997]_ , \new_[37000]_ ,
    \new_[37003]_ , \new_[37004]_ , \new_[37007]_ , \new_[37010]_ ,
    \new_[37011]_ , \new_[37012]_ , \new_[37016]_ , \new_[37017]_ ,
    \new_[37020]_ , \new_[37023]_ , \new_[37024]_ , \new_[37025]_ ,
    \new_[37028]_ , \new_[37031]_ , \new_[37032]_ , \new_[37035]_ ,
    \new_[37038]_ , \new_[37039]_ , \new_[37040]_ , \new_[37044]_ ,
    \new_[37045]_ , \new_[37048]_ , \new_[37051]_ , \new_[37052]_ ,
    \new_[37053]_ , \new_[37056]_ , \new_[37059]_ , \new_[37060]_ ,
    \new_[37063]_ , \new_[37066]_ , \new_[37067]_ , \new_[37068]_ ,
    \new_[37072]_ , \new_[37073]_ , \new_[37076]_ , \new_[37079]_ ,
    \new_[37080]_ , \new_[37081]_ , \new_[37084]_ , \new_[37087]_ ,
    \new_[37088]_ , \new_[37091]_ , \new_[37094]_ , \new_[37095]_ ,
    \new_[37096]_ , \new_[37100]_ , \new_[37101]_ , \new_[37104]_ ,
    \new_[37107]_ , \new_[37108]_ , \new_[37109]_ , \new_[37112]_ ,
    \new_[37115]_ , \new_[37116]_ , \new_[37119]_ , \new_[37122]_ ,
    \new_[37123]_ , \new_[37124]_ , \new_[37128]_ , \new_[37129]_ ,
    \new_[37132]_ , \new_[37135]_ , \new_[37136]_ , \new_[37137]_ ,
    \new_[37140]_ , \new_[37143]_ , \new_[37144]_ , \new_[37147]_ ,
    \new_[37150]_ , \new_[37151]_ , \new_[37152]_ , \new_[37156]_ ,
    \new_[37157]_ , \new_[37160]_ , \new_[37163]_ , \new_[37164]_ ,
    \new_[37165]_ , \new_[37168]_ , \new_[37171]_ , \new_[37172]_ ,
    \new_[37175]_ , \new_[37178]_ , \new_[37179]_ , \new_[37180]_ ,
    \new_[37184]_ , \new_[37185]_ , \new_[37188]_ , \new_[37191]_ ,
    \new_[37192]_ , \new_[37193]_ , \new_[37196]_ , \new_[37199]_ ,
    \new_[37200]_ , \new_[37203]_ , \new_[37206]_ , \new_[37207]_ ,
    \new_[37208]_ , \new_[37212]_ , \new_[37213]_ , \new_[37216]_ ,
    \new_[37219]_ , \new_[37220]_ , \new_[37221]_ , \new_[37224]_ ,
    \new_[37227]_ , \new_[37228]_ , \new_[37231]_ , \new_[37234]_ ,
    \new_[37235]_ , \new_[37236]_ , \new_[37240]_ , \new_[37241]_ ,
    \new_[37244]_ , \new_[37247]_ , \new_[37248]_ , \new_[37249]_ ,
    \new_[37252]_ , \new_[37255]_ , \new_[37256]_ , \new_[37259]_ ,
    \new_[37262]_ , \new_[37263]_ , \new_[37264]_ , \new_[37268]_ ,
    \new_[37269]_ , \new_[37272]_ , \new_[37275]_ , \new_[37276]_ ,
    \new_[37277]_ , \new_[37280]_ , \new_[37283]_ , \new_[37284]_ ,
    \new_[37287]_ , \new_[37290]_ , \new_[37291]_ , \new_[37292]_ ,
    \new_[37296]_ , \new_[37297]_ , \new_[37300]_ , \new_[37303]_ ,
    \new_[37304]_ , \new_[37305]_ , \new_[37308]_ , \new_[37311]_ ,
    \new_[37312]_ , \new_[37315]_ , \new_[37318]_ , \new_[37319]_ ,
    \new_[37320]_ , \new_[37324]_ , \new_[37325]_ , \new_[37328]_ ,
    \new_[37331]_ , \new_[37332]_ , \new_[37333]_ , \new_[37336]_ ,
    \new_[37339]_ , \new_[37340]_ , \new_[37343]_ , \new_[37346]_ ,
    \new_[37347]_ , \new_[37348]_ , \new_[37352]_ , \new_[37353]_ ,
    \new_[37356]_ , \new_[37359]_ , \new_[37360]_ , \new_[37361]_ ,
    \new_[37364]_ , \new_[37367]_ , \new_[37368]_ , \new_[37371]_ ,
    \new_[37374]_ , \new_[37375]_ , \new_[37376]_ , \new_[37380]_ ,
    \new_[37381]_ , \new_[37384]_ , \new_[37387]_ , \new_[37388]_ ,
    \new_[37389]_ , \new_[37392]_ , \new_[37395]_ , \new_[37396]_ ,
    \new_[37399]_ , \new_[37402]_ , \new_[37403]_ , \new_[37404]_ ,
    \new_[37408]_ , \new_[37409]_ , \new_[37412]_ , \new_[37415]_ ,
    \new_[37416]_ , \new_[37417]_ , \new_[37420]_ , \new_[37423]_ ,
    \new_[37424]_ , \new_[37427]_ , \new_[37430]_ , \new_[37431]_ ,
    \new_[37432]_ , \new_[37436]_ , \new_[37437]_ , \new_[37440]_ ,
    \new_[37443]_ , \new_[37444]_ , \new_[37445]_ , \new_[37448]_ ,
    \new_[37451]_ , \new_[37452]_ , \new_[37455]_ , \new_[37458]_ ,
    \new_[37459]_ , \new_[37460]_ , \new_[37464]_ , \new_[37465]_ ,
    \new_[37468]_ , \new_[37471]_ , \new_[37472]_ , \new_[37473]_ ,
    \new_[37476]_ , \new_[37479]_ , \new_[37480]_ , \new_[37483]_ ,
    \new_[37486]_ , \new_[37487]_ , \new_[37488]_ , \new_[37492]_ ,
    \new_[37493]_ , \new_[37496]_ , \new_[37499]_ , \new_[37500]_ ,
    \new_[37501]_ , \new_[37504]_ , \new_[37507]_ , \new_[37508]_ ,
    \new_[37511]_ , \new_[37514]_ , \new_[37515]_ , \new_[37516]_ ,
    \new_[37520]_ , \new_[37521]_ , \new_[37524]_ , \new_[37527]_ ,
    \new_[37528]_ , \new_[37529]_ , \new_[37532]_ , \new_[37535]_ ,
    \new_[37536]_ , \new_[37539]_ , \new_[37542]_ , \new_[37543]_ ,
    \new_[37544]_ , \new_[37548]_ , \new_[37549]_ , \new_[37552]_ ,
    \new_[37555]_ , \new_[37556]_ , \new_[37557]_ , \new_[37560]_ ,
    \new_[37563]_ , \new_[37564]_ , \new_[37567]_ , \new_[37570]_ ,
    \new_[37571]_ , \new_[37572]_ , \new_[37576]_ , \new_[37577]_ ,
    \new_[37580]_ , \new_[37583]_ , \new_[37584]_ , \new_[37585]_ ,
    \new_[37588]_ , \new_[37591]_ , \new_[37592]_ , \new_[37595]_ ,
    \new_[37598]_ , \new_[37599]_ , \new_[37600]_ , \new_[37604]_ ,
    \new_[37605]_ , \new_[37608]_ , \new_[37611]_ , \new_[37612]_ ,
    \new_[37613]_ , \new_[37616]_ , \new_[37619]_ , \new_[37620]_ ,
    \new_[37623]_ , \new_[37626]_ , \new_[37627]_ , \new_[37628]_ ,
    \new_[37632]_ , \new_[37633]_ , \new_[37636]_ , \new_[37639]_ ,
    \new_[37640]_ , \new_[37641]_ , \new_[37644]_ , \new_[37647]_ ,
    \new_[37648]_ , \new_[37651]_ , \new_[37654]_ , \new_[37655]_ ,
    \new_[37656]_ , \new_[37660]_ , \new_[37661]_ , \new_[37664]_ ,
    \new_[37667]_ , \new_[37668]_ , \new_[37669]_ , \new_[37672]_ ,
    \new_[37675]_ , \new_[37676]_ , \new_[37679]_ , \new_[37682]_ ,
    \new_[37683]_ , \new_[37684]_ , \new_[37688]_ , \new_[37689]_ ,
    \new_[37692]_ , \new_[37695]_ , \new_[37696]_ , \new_[37697]_ ,
    \new_[37700]_ , \new_[37703]_ , \new_[37704]_ , \new_[37707]_ ,
    \new_[37710]_ , \new_[37711]_ , \new_[37712]_ , \new_[37716]_ ,
    \new_[37717]_ , \new_[37720]_ , \new_[37723]_ , \new_[37724]_ ,
    \new_[37725]_ , \new_[37728]_ , \new_[37731]_ , \new_[37732]_ ,
    \new_[37735]_ , \new_[37738]_ , \new_[37739]_ , \new_[37740]_ ,
    \new_[37744]_ , \new_[37745]_ , \new_[37748]_ , \new_[37751]_ ,
    \new_[37752]_ , \new_[37753]_ , \new_[37756]_ , \new_[37759]_ ,
    \new_[37760]_ , \new_[37763]_ , \new_[37766]_ , \new_[37767]_ ,
    \new_[37768]_ , \new_[37772]_ , \new_[37773]_ , \new_[37776]_ ,
    \new_[37779]_ , \new_[37780]_ , \new_[37781]_ , \new_[37784]_ ,
    \new_[37787]_ , \new_[37788]_ , \new_[37791]_ , \new_[37794]_ ,
    \new_[37795]_ , \new_[37796]_ , \new_[37800]_ , \new_[37801]_ ,
    \new_[37804]_ , \new_[37807]_ , \new_[37808]_ , \new_[37809]_ ,
    \new_[37812]_ , \new_[37815]_ , \new_[37816]_ , \new_[37819]_ ,
    \new_[37822]_ , \new_[37823]_ , \new_[37824]_ , \new_[37828]_ ,
    \new_[37829]_ , \new_[37832]_ , \new_[37835]_ , \new_[37836]_ ,
    \new_[37837]_ , \new_[37840]_ , \new_[37843]_ , \new_[37844]_ ,
    \new_[37847]_ , \new_[37850]_ , \new_[37851]_ , \new_[37852]_ ,
    \new_[37856]_ , \new_[37857]_ , \new_[37860]_ , \new_[37863]_ ,
    \new_[37864]_ , \new_[37865]_ , \new_[37868]_ , \new_[37871]_ ,
    \new_[37872]_ , \new_[37875]_ , \new_[37878]_ , \new_[37879]_ ,
    \new_[37880]_ , \new_[37884]_ , \new_[37885]_ , \new_[37888]_ ,
    \new_[37891]_ , \new_[37892]_ , \new_[37893]_ , \new_[37896]_ ,
    \new_[37899]_ , \new_[37900]_ , \new_[37903]_ , \new_[37906]_ ,
    \new_[37907]_ , \new_[37908]_ , \new_[37912]_ , \new_[37913]_ ,
    \new_[37916]_ , \new_[37919]_ , \new_[37920]_ , \new_[37921]_ ,
    \new_[37924]_ , \new_[37927]_ , \new_[37928]_ , \new_[37931]_ ,
    \new_[37934]_ , \new_[37935]_ , \new_[37936]_ , \new_[37940]_ ,
    \new_[37941]_ , \new_[37944]_ , \new_[37947]_ , \new_[37948]_ ,
    \new_[37949]_ , \new_[37952]_ , \new_[37955]_ , \new_[37956]_ ,
    \new_[37959]_ , \new_[37962]_ , \new_[37963]_ , \new_[37964]_ ,
    \new_[37968]_ , \new_[37969]_ , \new_[37972]_ , \new_[37975]_ ,
    \new_[37976]_ , \new_[37977]_ , \new_[37980]_ , \new_[37983]_ ,
    \new_[37984]_ , \new_[37987]_ , \new_[37990]_ , \new_[37991]_ ,
    \new_[37992]_ , \new_[37996]_ , \new_[37997]_ , \new_[38000]_ ,
    \new_[38003]_ , \new_[38004]_ , \new_[38005]_ , \new_[38008]_ ,
    \new_[38011]_ , \new_[38012]_ , \new_[38015]_ , \new_[38018]_ ,
    \new_[38019]_ , \new_[38020]_ , \new_[38024]_ , \new_[38025]_ ,
    \new_[38028]_ , \new_[38031]_ , \new_[38032]_ , \new_[38033]_ ,
    \new_[38036]_ , \new_[38039]_ , \new_[38040]_ , \new_[38043]_ ,
    \new_[38046]_ , \new_[38047]_ , \new_[38048]_ , \new_[38052]_ ,
    \new_[38053]_ , \new_[38056]_ , \new_[38059]_ , \new_[38060]_ ,
    \new_[38061]_ , \new_[38064]_ , \new_[38067]_ , \new_[38068]_ ,
    \new_[38071]_ , \new_[38074]_ , \new_[38075]_ , \new_[38076]_ ,
    \new_[38080]_ , \new_[38081]_ , \new_[38084]_ , \new_[38087]_ ,
    \new_[38088]_ , \new_[38089]_ , \new_[38092]_ , \new_[38095]_ ,
    \new_[38096]_ , \new_[38099]_ , \new_[38102]_ , \new_[38103]_ ,
    \new_[38104]_ , \new_[38108]_ , \new_[38109]_ , \new_[38112]_ ,
    \new_[38115]_ , \new_[38116]_ , \new_[38117]_ , \new_[38120]_ ,
    \new_[38123]_ , \new_[38124]_ , \new_[38127]_ , \new_[38130]_ ,
    \new_[38131]_ , \new_[38132]_ , \new_[38136]_ , \new_[38137]_ ,
    \new_[38140]_ , \new_[38143]_ , \new_[38144]_ , \new_[38145]_ ,
    \new_[38148]_ , \new_[38151]_ , \new_[38152]_ , \new_[38155]_ ,
    \new_[38158]_ , \new_[38159]_ , \new_[38160]_ , \new_[38164]_ ,
    \new_[38165]_ , \new_[38168]_ , \new_[38171]_ , \new_[38172]_ ,
    \new_[38173]_ , \new_[38176]_ , \new_[38179]_ , \new_[38180]_ ,
    \new_[38183]_ , \new_[38186]_ , \new_[38187]_ , \new_[38188]_ ,
    \new_[38192]_ , \new_[38193]_ , \new_[38196]_ , \new_[38199]_ ,
    \new_[38200]_ , \new_[38201]_ , \new_[38204]_ , \new_[38207]_ ,
    \new_[38208]_ , \new_[38211]_ , \new_[38214]_ , \new_[38215]_ ,
    \new_[38216]_ , \new_[38220]_ , \new_[38221]_ , \new_[38224]_ ,
    \new_[38227]_ , \new_[38228]_ , \new_[38229]_ , \new_[38232]_ ,
    \new_[38235]_ , \new_[38236]_ , \new_[38239]_ , \new_[38242]_ ,
    \new_[38243]_ , \new_[38244]_ , \new_[38248]_ , \new_[38249]_ ,
    \new_[38252]_ , \new_[38255]_ , \new_[38256]_ , \new_[38257]_ ,
    \new_[38260]_ , \new_[38263]_ , \new_[38264]_ , \new_[38267]_ ,
    \new_[38270]_ , \new_[38271]_ , \new_[38272]_ , \new_[38276]_ ,
    \new_[38277]_ , \new_[38280]_ , \new_[38283]_ , \new_[38284]_ ,
    \new_[38285]_ , \new_[38288]_ , \new_[38291]_ , \new_[38292]_ ,
    \new_[38295]_ , \new_[38298]_ , \new_[38299]_ , \new_[38300]_ ,
    \new_[38304]_ , \new_[38305]_ , \new_[38308]_ , \new_[38311]_ ,
    \new_[38312]_ , \new_[38313]_ , \new_[38316]_ , \new_[38319]_ ,
    \new_[38320]_ , \new_[38323]_ , \new_[38326]_ , \new_[38327]_ ,
    \new_[38328]_ , \new_[38332]_ , \new_[38333]_ , \new_[38336]_ ,
    \new_[38339]_ , \new_[38340]_ , \new_[38341]_ , \new_[38344]_ ,
    \new_[38347]_ , \new_[38348]_ , \new_[38351]_ , \new_[38354]_ ,
    \new_[38355]_ , \new_[38356]_ , \new_[38360]_ , \new_[38361]_ ,
    \new_[38364]_ , \new_[38367]_ , \new_[38368]_ , \new_[38369]_ ,
    \new_[38372]_ , \new_[38375]_ , \new_[38376]_ , \new_[38379]_ ,
    \new_[38382]_ , \new_[38383]_ , \new_[38384]_ , \new_[38388]_ ,
    \new_[38389]_ , \new_[38392]_ , \new_[38395]_ , \new_[38396]_ ,
    \new_[38397]_ , \new_[38400]_ , \new_[38403]_ , \new_[38404]_ ,
    \new_[38407]_ , \new_[38410]_ , \new_[38411]_ , \new_[38412]_ ,
    \new_[38416]_ , \new_[38417]_ , \new_[38420]_ , \new_[38423]_ ,
    \new_[38424]_ , \new_[38425]_ , \new_[38428]_ , \new_[38431]_ ,
    \new_[38432]_ , \new_[38435]_ , \new_[38438]_ , \new_[38439]_ ,
    \new_[38440]_ , \new_[38444]_ , \new_[38445]_ , \new_[38448]_ ,
    \new_[38451]_ , \new_[38452]_ , \new_[38453]_ , \new_[38456]_ ,
    \new_[38459]_ , \new_[38460]_ , \new_[38463]_ , \new_[38466]_ ,
    \new_[38467]_ , \new_[38468]_ , \new_[38472]_ , \new_[38473]_ ,
    \new_[38476]_ , \new_[38479]_ , \new_[38480]_ , \new_[38481]_ ,
    \new_[38484]_ , \new_[38487]_ , \new_[38488]_ , \new_[38491]_ ,
    \new_[38494]_ , \new_[38495]_ , \new_[38496]_ , \new_[38500]_ ,
    \new_[38501]_ , \new_[38504]_ , \new_[38507]_ , \new_[38508]_ ,
    \new_[38509]_ , \new_[38512]_ , \new_[38515]_ , \new_[38516]_ ,
    \new_[38519]_ , \new_[38522]_ , \new_[38523]_ , \new_[38524]_ ,
    \new_[38528]_ , \new_[38529]_ , \new_[38532]_ , \new_[38535]_ ,
    \new_[38536]_ , \new_[38537]_ , \new_[38540]_ , \new_[38543]_ ,
    \new_[38544]_ , \new_[38547]_ , \new_[38550]_ , \new_[38551]_ ,
    \new_[38552]_ , \new_[38556]_ , \new_[38557]_ , \new_[38560]_ ,
    \new_[38563]_ , \new_[38564]_ , \new_[38565]_ , \new_[38568]_ ,
    \new_[38571]_ , \new_[38572]_ , \new_[38575]_ , \new_[38578]_ ,
    \new_[38579]_ , \new_[38580]_ , \new_[38584]_ , \new_[38585]_ ,
    \new_[38588]_ , \new_[38591]_ , \new_[38592]_ , \new_[38593]_ ,
    \new_[38596]_ , \new_[38599]_ , \new_[38600]_ , \new_[38603]_ ,
    \new_[38606]_ , \new_[38607]_ , \new_[38608]_ , \new_[38612]_ ,
    \new_[38613]_ , \new_[38616]_ , \new_[38619]_ , \new_[38620]_ ,
    \new_[38621]_ , \new_[38624]_ , \new_[38627]_ , \new_[38628]_ ,
    \new_[38631]_ , \new_[38634]_ , \new_[38635]_ , \new_[38636]_ ,
    \new_[38640]_ , \new_[38641]_ , \new_[38644]_ , \new_[38647]_ ,
    \new_[38648]_ , \new_[38649]_ , \new_[38652]_ , \new_[38655]_ ,
    \new_[38656]_ , \new_[38659]_ , \new_[38662]_ , \new_[38663]_ ,
    \new_[38664]_ , \new_[38668]_ , \new_[38669]_ , \new_[38672]_ ,
    \new_[38675]_ , \new_[38676]_ , \new_[38677]_ , \new_[38680]_ ,
    \new_[38683]_ , \new_[38684]_ , \new_[38687]_ , \new_[38690]_ ,
    \new_[38691]_ , \new_[38692]_ , \new_[38696]_ , \new_[38697]_ ,
    \new_[38700]_ , \new_[38703]_ , \new_[38704]_ , \new_[38705]_ ,
    \new_[38708]_ , \new_[38711]_ , \new_[38712]_ , \new_[38715]_ ,
    \new_[38718]_ , \new_[38719]_ , \new_[38720]_ , \new_[38724]_ ,
    \new_[38725]_ , \new_[38728]_ , \new_[38731]_ , \new_[38732]_ ,
    \new_[38733]_ , \new_[38736]_ , \new_[38739]_ , \new_[38740]_ ,
    \new_[38743]_ , \new_[38746]_ , \new_[38747]_ , \new_[38748]_ ,
    \new_[38752]_ , \new_[38753]_ , \new_[38756]_ , \new_[38759]_ ,
    \new_[38760]_ , \new_[38761]_ , \new_[38764]_ , \new_[38767]_ ,
    \new_[38768]_ , \new_[38771]_ , \new_[38774]_ , \new_[38775]_ ,
    \new_[38776]_ , \new_[38780]_ , \new_[38781]_ , \new_[38784]_ ,
    \new_[38787]_ , \new_[38788]_ , \new_[38789]_ , \new_[38792]_ ,
    \new_[38795]_ , \new_[38796]_ , \new_[38799]_ , \new_[38802]_ ,
    \new_[38803]_ , \new_[38804]_ , \new_[38808]_ , \new_[38809]_ ,
    \new_[38812]_ , \new_[38815]_ , \new_[38816]_ , \new_[38817]_ ,
    \new_[38820]_ , \new_[38823]_ , \new_[38824]_ , \new_[38827]_ ,
    \new_[38830]_ , \new_[38831]_ , \new_[38832]_ , \new_[38836]_ ,
    \new_[38837]_ , \new_[38840]_ , \new_[38843]_ , \new_[38844]_ ,
    \new_[38845]_ , \new_[38848]_ , \new_[38851]_ , \new_[38852]_ ,
    \new_[38855]_ , \new_[38858]_ , \new_[38859]_ , \new_[38860]_ ,
    \new_[38864]_ , \new_[38865]_ , \new_[38868]_ , \new_[38871]_ ,
    \new_[38872]_ , \new_[38873]_ , \new_[38876]_ , \new_[38879]_ ,
    \new_[38880]_ , \new_[38883]_ , \new_[38886]_ , \new_[38887]_ ,
    \new_[38888]_ , \new_[38892]_ , \new_[38893]_ , \new_[38896]_ ,
    \new_[38899]_ , \new_[38900]_ , \new_[38901]_ , \new_[38904]_ ,
    \new_[38907]_ , \new_[38908]_ , \new_[38911]_ , \new_[38914]_ ,
    \new_[38915]_ , \new_[38916]_ , \new_[38920]_ , \new_[38921]_ ,
    \new_[38924]_ , \new_[38927]_ , \new_[38928]_ , \new_[38929]_ ,
    \new_[38932]_ , \new_[38935]_ , \new_[38936]_ , \new_[38939]_ ,
    \new_[38942]_ , \new_[38943]_ , \new_[38944]_ , \new_[38948]_ ,
    \new_[38949]_ , \new_[38952]_ , \new_[38955]_ , \new_[38956]_ ,
    \new_[38957]_ , \new_[38960]_ , \new_[38963]_ , \new_[38964]_ ,
    \new_[38967]_ , \new_[38970]_ , \new_[38971]_ , \new_[38972]_ ,
    \new_[38976]_ , \new_[38977]_ , \new_[38980]_ , \new_[38983]_ ,
    \new_[38984]_ , \new_[38985]_ , \new_[38988]_ , \new_[38991]_ ,
    \new_[38992]_ , \new_[38995]_ , \new_[38998]_ , \new_[38999]_ ,
    \new_[39000]_ , \new_[39004]_ , \new_[39005]_ , \new_[39008]_ ,
    \new_[39011]_ , \new_[39012]_ , \new_[39013]_ , \new_[39016]_ ,
    \new_[39019]_ , \new_[39020]_ , \new_[39023]_ , \new_[39026]_ ,
    \new_[39027]_ , \new_[39028]_ , \new_[39032]_ , \new_[39033]_ ,
    \new_[39036]_ , \new_[39039]_ , \new_[39040]_ , \new_[39041]_ ,
    \new_[39044]_ , \new_[39047]_ , \new_[39048]_ , \new_[39051]_ ,
    \new_[39054]_ , \new_[39055]_ , \new_[39056]_ , \new_[39060]_ ,
    \new_[39061]_ , \new_[39064]_ , \new_[39067]_ , \new_[39068]_ ,
    \new_[39069]_ , \new_[39072]_ , \new_[39075]_ , \new_[39076]_ ,
    \new_[39079]_ , \new_[39082]_ , \new_[39083]_ , \new_[39084]_ ,
    \new_[39088]_ , \new_[39089]_ , \new_[39092]_ , \new_[39095]_ ,
    \new_[39096]_ , \new_[39097]_ , \new_[39100]_ , \new_[39103]_ ,
    \new_[39104]_ , \new_[39107]_ , \new_[39110]_ , \new_[39111]_ ,
    \new_[39112]_ , \new_[39116]_ , \new_[39117]_ , \new_[39120]_ ,
    \new_[39123]_ , \new_[39124]_ , \new_[39125]_ , \new_[39128]_ ,
    \new_[39131]_ , \new_[39132]_ , \new_[39135]_ , \new_[39138]_ ,
    \new_[39139]_ , \new_[39140]_ , \new_[39144]_ , \new_[39145]_ ,
    \new_[39148]_ , \new_[39151]_ , \new_[39152]_ , \new_[39153]_ ,
    \new_[39156]_ , \new_[39159]_ , \new_[39160]_ , \new_[39163]_ ,
    \new_[39166]_ , \new_[39167]_ , \new_[39168]_ , \new_[39172]_ ,
    \new_[39173]_ , \new_[39176]_ , \new_[39179]_ , \new_[39180]_ ,
    \new_[39181]_ , \new_[39184]_ , \new_[39187]_ , \new_[39188]_ ,
    \new_[39191]_ , \new_[39194]_ , \new_[39195]_ , \new_[39196]_ ,
    \new_[39200]_ , \new_[39201]_ , \new_[39204]_ , \new_[39207]_ ,
    \new_[39208]_ , \new_[39209]_ , \new_[39212]_ , \new_[39215]_ ,
    \new_[39216]_ , \new_[39219]_ , \new_[39222]_ , \new_[39223]_ ,
    \new_[39224]_ , \new_[39228]_ , \new_[39229]_ , \new_[39232]_ ,
    \new_[39235]_ , \new_[39236]_ , \new_[39237]_ , \new_[39240]_ ,
    \new_[39243]_ , \new_[39244]_ , \new_[39247]_ , \new_[39250]_ ,
    \new_[39251]_ , \new_[39252]_ , \new_[39256]_ , \new_[39257]_ ,
    \new_[39260]_ , \new_[39263]_ , \new_[39264]_ , \new_[39265]_ ,
    \new_[39268]_ , \new_[39271]_ , \new_[39272]_ , \new_[39275]_ ,
    \new_[39278]_ , \new_[39279]_ , \new_[39280]_ , \new_[39284]_ ,
    \new_[39285]_ , \new_[39288]_ , \new_[39291]_ , \new_[39292]_ ,
    \new_[39293]_ , \new_[39296]_ , \new_[39299]_ , \new_[39300]_ ,
    \new_[39303]_ , \new_[39306]_ , \new_[39307]_ , \new_[39308]_ ,
    \new_[39312]_ , \new_[39313]_ , \new_[39316]_ , \new_[39319]_ ,
    \new_[39320]_ , \new_[39321]_ , \new_[39324]_ , \new_[39327]_ ,
    \new_[39328]_ , \new_[39331]_ , \new_[39334]_ , \new_[39335]_ ,
    \new_[39336]_ , \new_[39340]_ , \new_[39341]_ , \new_[39344]_ ,
    \new_[39347]_ , \new_[39348]_ , \new_[39349]_ , \new_[39352]_ ,
    \new_[39355]_ , \new_[39356]_ , \new_[39359]_ , \new_[39362]_ ,
    \new_[39363]_ , \new_[39364]_ , \new_[39368]_ , \new_[39369]_ ,
    \new_[39372]_ , \new_[39375]_ , \new_[39376]_ , \new_[39377]_ ,
    \new_[39380]_ , \new_[39383]_ , \new_[39384]_ , \new_[39387]_ ,
    \new_[39390]_ , \new_[39391]_ , \new_[39392]_ , \new_[39396]_ ,
    \new_[39397]_ , \new_[39400]_ , \new_[39403]_ , \new_[39404]_ ,
    \new_[39405]_ , \new_[39408]_ , \new_[39411]_ , \new_[39412]_ ,
    \new_[39415]_ , \new_[39418]_ , \new_[39419]_ , \new_[39420]_ ,
    \new_[39424]_ , \new_[39425]_ , \new_[39428]_ , \new_[39431]_ ,
    \new_[39432]_ , \new_[39433]_ , \new_[39436]_ , \new_[39439]_ ,
    \new_[39440]_ , \new_[39443]_ , \new_[39446]_ , \new_[39447]_ ,
    \new_[39448]_ , \new_[39452]_ , \new_[39453]_ , \new_[39456]_ ,
    \new_[39459]_ , \new_[39460]_ , \new_[39461]_ , \new_[39464]_ ,
    \new_[39467]_ , \new_[39468]_ , \new_[39471]_ , \new_[39474]_ ,
    \new_[39475]_ , \new_[39476]_ , \new_[39480]_ , \new_[39481]_ ,
    \new_[39484]_ , \new_[39487]_ , \new_[39488]_ , \new_[39489]_ ,
    \new_[39492]_ , \new_[39495]_ , \new_[39496]_ , \new_[39499]_ ,
    \new_[39502]_ , \new_[39503]_ , \new_[39504]_ , \new_[39508]_ ,
    \new_[39509]_ , \new_[39512]_ , \new_[39515]_ , \new_[39516]_ ,
    \new_[39517]_ , \new_[39520]_ , \new_[39523]_ , \new_[39524]_ ,
    \new_[39527]_ , \new_[39530]_ , \new_[39531]_ , \new_[39532]_ ,
    \new_[39536]_ , \new_[39537]_ , \new_[39540]_ , \new_[39543]_ ,
    \new_[39544]_ , \new_[39545]_ , \new_[39548]_ , \new_[39551]_ ,
    \new_[39552]_ , \new_[39555]_ , \new_[39558]_ , \new_[39559]_ ,
    \new_[39560]_ , \new_[39564]_ , \new_[39565]_ , \new_[39568]_ ,
    \new_[39571]_ , \new_[39572]_ , \new_[39573]_ , \new_[39576]_ ,
    \new_[39579]_ , \new_[39580]_ , \new_[39583]_ , \new_[39586]_ ,
    \new_[39587]_ , \new_[39588]_ , \new_[39592]_ , \new_[39593]_ ,
    \new_[39596]_ , \new_[39599]_ , \new_[39600]_ , \new_[39601]_ ,
    \new_[39604]_ , \new_[39607]_ , \new_[39608]_ , \new_[39611]_ ,
    \new_[39614]_ , \new_[39615]_ , \new_[39616]_ , \new_[39620]_ ,
    \new_[39621]_ , \new_[39624]_ , \new_[39627]_ , \new_[39628]_ ,
    \new_[39629]_ , \new_[39632]_ , \new_[39635]_ , \new_[39636]_ ,
    \new_[39639]_ , \new_[39642]_ , \new_[39643]_ , \new_[39644]_ ,
    \new_[39648]_ , \new_[39649]_ , \new_[39652]_ , \new_[39655]_ ,
    \new_[39656]_ , \new_[39657]_ , \new_[39660]_ , \new_[39663]_ ,
    \new_[39664]_ , \new_[39667]_ , \new_[39670]_ , \new_[39671]_ ,
    \new_[39672]_ , \new_[39676]_ , \new_[39677]_ , \new_[39680]_ ,
    \new_[39683]_ , \new_[39684]_ , \new_[39685]_ , \new_[39688]_ ,
    \new_[39691]_ , \new_[39692]_ , \new_[39695]_ , \new_[39698]_ ,
    \new_[39699]_ , \new_[39700]_ , \new_[39704]_ , \new_[39705]_ ,
    \new_[39708]_ , \new_[39711]_ , \new_[39712]_ , \new_[39713]_ ,
    \new_[39716]_ , \new_[39719]_ , \new_[39720]_ , \new_[39723]_ ,
    \new_[39726]_ , \new_[39727]_ , \new_[39728]_ , \new_[39732]_ ,
    \new_[39733]_ , \new_[39736]_ , \new_[39739]_ , \new_[39740]_ ,
    \new_[39741]_ , \new_[39744]_ , \new_[39747]_ , \new_[39748]_ ,
    \new_[39751]_ , \new_[39754]_ , \new_[39755]_ , \new_[39756]_ ,
    \new_[39760]_ , \new_[39761]_ , \new_[39764]_ , \new_[39767]_ ,
    \new_[39768]_ , \new_[39769]_ , \new_[39772]_ , \new_[39775]_ ,
    \new_[39776]_ , \new_[39779]_ , \new_[39782]_ , \new_[39783]_ ,
    \new_[39784]_ , \new_[39788]_ , \new_[39789]_ , \new_[39792]_ ,
    \new_[39795]_ , \new_[39796]_ , \new_[39797]_ , \new_[39800]_ ,
    \new_[39803]_ , \new_[39804]_ , \new_[39807]_ , \new_[39810]_ ,
    \new_[39811]_ , \new_[39812]_ , \new_[39816]_ , \new_[39817]_ ,
    \new_[39820]_ , \new_[39823]_ , \new_[39824]_ , \new_[39825]_ ,
    \new_[39828]_ , \new_[39831]_ , \new_[39832]_ , \new_[39835]_ ,
    \new_[39838]_ , \new_[39839]_ , \new_[39840]_ , \new_[39844]_ ,
    \new_[39845]_ , \new_[39848]_ , \new_[39851]_ , \new_[39852]_ ,
    \new_[39853]_ , \new_[39856]_ , \new_[39859]_ , \new_[39860]_ ,
    \new_[39863]_ , \new_[39866]_ , \new_[39867]_ , \new_[39868]_ ,
    \new_[39872]_ , \new_[39873]_ , \new_[39876]_ , \new_[39879]_ ,
    \new_[39880]_ , \new_[39881]_ , \new_[39884]_ , \new_[39887]_ ,
    \new_[39888]_ , \new_[39891]_ , \new_[39894]_ , \new_[39895]_ ,
    \new_[39896]_ , \new_[39900]_ , \new_[39901]_ , \new_[39904]_ ,
    \new_[39907]_ , \new_[39908]_ , \new_[39909]_ , \new_[39912]_ ,
    \new_[39915]_ , \new_[39916]_ , \new_[39919]_ , \new_[39922]_ ,
    \new_[39923]_ , \new_[39924]_ , \new_[39928]_ , \new_[39929]_ ,
    \new_[39932]_ , \new_[39935]_ , \new_[39936]_ , \new_[39937]_ ,
    \new_[39940]_ , \new_[39943]_ , \new_[39944]_ , \new_[39947]_ ,
    \new_[39950]_ , \new_[39951]_ , \new_[39952]_ , \new_[39956]_ ,
    \new_[39957]_ , \new_[39960]_ , \new_[39963]_ , \new_[39964]_ ,
    \new_[39965]_ , \new_[39968]_ , \new_[39971]_ , \new_[39972]_ ,
    \new_[39975]_ , \new_[39978]_ , \new_[39979]_ , \new_[39980]_ ,
    \new_[39984]_ , \new_[39985]_ , \new_[39988]_ , \new_[39991]_ ,
    \new_[39992]_ , \new_[39993]_ , \new_[39996]_ , \new_[39999]_ ,
    \new_[40000]_ , \new_[40003]_ , \new_[40006]_ , \new_[40007]_ ,
    \new_[40008]_ , \new_[40012]_ , \new_[40013]_ , \new_[40016]_ ,
    \new_[40019]_ , \new_[40020]_ , \new_[40021]_ , \new_[40024]_ ,
    \new_[40027]_ , \new_[40028]_ , \new_[40031]_ , \new_[40034]_ ,
    \new_[40035]_ , \new_[40036]_ , \new_[40040]_ , \new_[40041]_ ,
    \new_[40044]_ , \new_[40047]_ , \new_[40048]_ , \new_[40049]_ ,
    \new_[40052]_ , \new_[40055]_ , \new_[40056]_ , \new_[40059]_ ,
    \new_[40062]_ , \new_[40063]_ , \new_[40064]_ , \new_[40068]_ ,
    \new_[40069]_ , \new_[40072]_ , \new_[40075]_ , \new_[40076]_ ,
    \new_[40077]_ , \new_[40080]_ , \new_[40083]_ , \new_[40084]_ ,
    \new_[40087]_ , \new_[40090]_ , \new_[40091]_ , \new_[40092]_ ,
    \new_[40096]_ , \new_[40097]_ , \new_[40100]_ , \new_[40103]_ ,
    \new_[40104]_ , \new_[40105]_ , \new_[40108]_ , \new_[40111]_ ,
    \new_[40112]_ , \new_[40115]_ , \new_[40118]_ , \new_[40119]_ ,
    \new_[40120]_ , \new_[40124]_ , \new_[40125]_ , \new_[40128]_ ,
    \new_[40131]_ , \new_[40132]_ , \new_[40133]_ , \new_[40136]_ ,
    \new_[40139]_ , \new_[40140]_ , \new_[40143]_ , \new_[40146]_ ,
    \new_[40147]_ , \new_[40148]_ , \new_[40152]_ , \new_[40153]_ ,
    \new_[40156]_ , \new_[40159]_ , \new_[40160]_ , \new_[40161]_ ,
    \new_[40164]_ , \new_[40167]_ , \new_[40168]_ , \new_[40171]_ ,
    \new_[40174]_ , \new_[40175]_ , \new_[40176]_ , \new_[40180]_ ,
    \new_[40181]_ , \new_[40184]_ , \new_[40187]_ , \new_[40188]_ ,
    \new_[40189]_ , \new_[40192]_ , \new_[40195]_ , \new_[40196]_ ,
    \new_[40199]_ , \new_[40202]_ , \new_[40203]_ , \new_[40204]_ ,
    \new_[40208]_ , \new_[40209]_ , \new_[40212]_ , \new_[40215]_ ,
    \new_[40216]_ , \new_[40217]_ , \new_[40220]_ , \new_[40223]_ ,
    \new_[40224]_ , \new_[40227]_ , \new_[40230]_ , \new_[40231]_ ,
    \new_[40232]_ , \new_[40236]_ , \new_[40237]_ , \new_[40240]_ ,
    \new_[40243]_ , \new_[40244]_ , \new_[40245]_ , \new_[40248]_ ,
    \new_[40251]_ , \new_[40252]_ , \new_[40255]_ , \new_[40258]_ ,
    \new_[40259]_ , \new_[40260]_ , \new_[40264]_ , \new_[40265]_ ,
    \new_[40268]_ , \new_[40271]_ , \new_[40272]_ , \new_[40273]_ ,
    \new_[40276]_ , \new_[40279]_ , \new_[40280]_ , \new_[40283]_ ,
    \new_[40286]_ , \new_[40287]_ , \new_[40288]_ , \new_[40292]_ ,
    \new_[40293]_ , \new_[40296]_ , \new_[40299]_ , \new_[40300]_ ,
    \new_[40301]_ , \new_[40304]_ , \new_[40307]_ , \new_[40308]_ ,
    \new_[40311]_ , \new_[40314]_ , \new_[40315]_ , \new_[40316]_ ,
    \new_[40320]_ , \new_[40321]_ , \new_[40324]_ , \new_[40327]_ ,
    \new_[40328]_ , \new_[40329]_ , \new_[40332]_ , \new_[40335]_ ,
    \new_[40336]_ , \new_[40339]_ , \new_[40342]_ , \new_[40343]_ ,
    \new_[40344]_ , \new_[40348]_ , \new_[40349]_ , \new_[40352]_ ,
    \new_[40355]_ , \new_[40356]_ , \new_[40357]_ , \new_[40360]_ ,
    \new_[40363]_ , \new_[40364]_ , \new_[40367]_ , \new_[40370]_ ,
    \new_[40371]_ , \new_[40372]_ , \new_[40376]_ , \new_[40377]_ ,
    \new_[40380]_ , \new_[40383]_ , \new_[40384]_ , \new_[40385]_ ,
    \new_[40388]_ , \new_[40391]_ , \new_[40392]_ , \new_[40395]_ ,
    \new_[40398]_ , \new_[40399]_ , \new_[40400]_ , \new_[40404]_ ,
    \new_[40405]_ , \new_[40408]_ , \new_[40411]_ , \new_[40412]_ ,
    \new_[40413]_ , \new_[40416]_ , \new_[40419]_ , \new_[40420]_ ,
    \new_[40423]_ , \new_[40426]_ , \new_[40427]_ , \new_[40428]_ ,
    \new_[40432]_ , \new_[40433]_ , \new_[40436]_ , \new_[40439]_ ,
    \new_[40440]_ , \new_[40441]_ , \new_[40444]_ , \new_[40447]_ ,
    \new_[40448]_ , \new_[40451]_ , \new_[40454]_ , \new_[40455]_ ,
    \new_[40456]_ , \new_[40460]_ , \new_[40461]_ , \new_[40464]_ ,
    \new_[40467]_ , \new_[40468]_ , \new_[40469]_ , \new_[40472]_ ,
    \new_[40475]_ , \new_[40476]_ , \new_[40479]_ , \new_[40482]_ ,
    \new_[40483]_ , \new_[40484]_ , \new_[40488]_ , \new_[40489]_ ,
    \new_[40492]_ , \new_[40495]_ , \new_[40496]_ , \new_[40497]_ ,
    \new_[40500]_ , \new_[40503]_ , \new_[40504]_ , \new_[40507]_ ,
    \new_[40510]_ , \new_[40511]_ , \new_[40512]_ , \new_[40516]_ ,
    \new_[40517]_ , \new_[40520]_ , \new_[40523]_ , \new_[40524]_ ,
    \new_[40525]_ , \new_[40528]_ , \new_[40531]_ , \new_[40532]_ ,
    \new_[40535]_ , \new_[40538]_ , \new_[40539]_ , \new_[40540]_ ,
    \new_[40544]_ , \new_[40545]_ , \new_[40548]_ , \new_[40551]_ ,
    \new_[40552]_ , \new_[40553]_ , \new_[40556]_ , \new_[40559]_ ,
    \new_[40560]_ , \new_[40563]_ , \new_[40566]_ , \new_[40567]_ ,
    \new_[40568]_ , \new_[40572]_ , \new_[40573]_ , \new_[40576]_ ,
    \new_[40579]_ , \new_[40580]_ , \new_[40581]_ , \new_[40584]_ ,
    \new_[40587]_ , \new_[40588]_ , \new_[40591]_ , \new_[40594]_ ,
    \new_[40595]_ , \new_[40596]_ , \new_[40600]_ , \new_[40601]_ ,
    \new_[40604]_ , \new_[40607]_ , \new_[40608]_ , \new_[40609]_ ,
    \new_[40612]_ , \new_[40615]_ , \new_[40616]_ , \new_[40619]_ ,
    \new_[40622]_ , \new_[40623]_ , \new_[40624]_ , \new_[40628]_ ,
    \new_[40629]_ , \new_[40632]_ , \new_[40635]_ , \new_[40636]_ ,
    \new_[40637]_ , \new_[40640]_ , \new_[40643]_ , \new_[40644]_ ,
    \new_[40647]_ , \new_[40650]_ , \new_[40651]_ , \new_[40652]_ ,
    \new_[40656]_ , \new_[40657]_ , \new_[40660]_ , \new_[40663]_ ,
    \new_[40664]_ , \new_[40665]_ , \new_[40668]_ , \new_[40671]_ ,
    \new_[40672]_ , \new_[40675]_ , \new_[40678]_ , \new_[40679]_ ,
    \new_[40680]_ , \new_[40684]_ , \new_[40685]_ , \new_[40688]_ ,
    \new_[40691]_ , \new_[40692]_ , \new_[40693]_ , \new_[40696]_ ,
    \new_[40699]_ , \new_[40700]_ , \new_[40703]_ , \new_[40706]_ ,
    \new_[40707]_ , \new_[40708]_ , \new_[40712]_ , \new_[40713]_ ,
    \new_[40716]_ , \new_[40719]_ , \new_[40720]_ , \new_[40721]_ ,
    \new_[40724]_ , \new_[40727]_ , \new_[40728]_ , \new_[40731]_ ,
    \new_[40734]_ , \new_[40735]_ , \new_[40736]_ , \new_[40740]_ ,
    \new_[40741]_ , \new_[40744]_ , \new_[40747]_ , \new_[40748]_ ,
    \new_[40749]_ , \new_[40752]_ , \new_[40755]_ , \new_[40756]_ ,
    \new_[40759]_ , \new_[40762]_ , \new_[40763]_ , \new_[40764]_ ,
    \new_[40768]_ , \new_[40769]_ , \new_[40772]_ , \new_[40775]_ ,
    \new_[40776]_ , \new_[40777]_ , \new_[40780]_ , \new_[40783]_ ,
    \new_[40784]_ , \new_[40787]_ , \new_[40790]_ , \new_[40791]_ ,
    \new_[40792]_ , \new_[40796]_ , \new_[40797]_ , \new_[40800]_ ,
    \new_[40803]_ , \new_[40804]_ , \new_[40805]_ , \new_[40808]_ ,
    \new_[40811]_ , \new_[40812]_ , \new_[40815]_ , \new_[40818]_ ,
    \new_[40819]_ , \new_[40820]_ , \new_[40824]_ , \new_[40825]_ ,
    \new_[40828]_ , \new_[40831]_ , \new_[40832]_ , \new_[40833]_ ,
    \new_[40836]_ , \new_[40839]_ , \new_[40840]_ , \new_[40843]_ ,
    \new_[40846]_ , \new_[40847]_ , \new_[40848]_ , \new_[40852]_ ,
    \new_[40853]_ , \new_[40856]_ , \new_[40859]_ , \new_[40860]_ ,
    \new_[40861]_ , \new_[40864]_ , \new_[40867]_ , \new_[40868]_ ,
    \new_[40871]_ , \new_[40874]_ , \new_[40875]_ , \new_[40876]_ ,
    \new_[40880]_ , \new_[40881]_ , \new_[40884]_ , \new_[40887]_ ,
    \new_[40888]_ , \new_[40889]_ , \new_[40892]_ , \new_[40895]_ ,
    \new_[40896]_ , \new_[40899]_ , \new_[40902]_ , \new_[40903]_ ,
    \new_[40904]_ , \new_[40908]_ , \new_[40909]_ , \new_[40912]_ ,
    \new_[40915]_ , \new_[40916]_ , \new_[40917]_ , \new_[40920]_ ,
    \new_[40923]_ , \new_[40924]_ , \new_[40927]_ , \new_[40930]_ ,
    \new_[40931]_ , \new_[40932]_ , \new_[40936]_ , \new_[40937]_ ,
    \new_[40940]_ , \new_[40943]_ , \new_[40944]_ , \new_[40945]_ ,
    \new_[40948]_ , \new_[40951]_ , \new_[40952]_ , \new_[40955]_ ,
    \new_[40958]_ , \new_[40959]_ , \new_[40960]_ , \new_[40964]_ ,
    \new_[40965]_ , \new_[40968]_ , \new_[40971]_ , \new_[40972]_ ,
    \new_[40973]_ , \new_[40976]_ , \new_[40979]_ , \new_[40980]_ ,
    \new_[40983]_ , \new_[40986]_ , \new_[40987]_ , \new_[40988]_ ,
    \new_[40992]_ , \new_[40993]_ , \new_[40996]_ , \new_[40999]_ ,
    \new_[41000]_ , \new_[41001]_ , \new_[41004]_ , \new_[41007]_ ,
    \new_[41008]_ , \new_[41011]_ , \new_[41014]_ , \new_[41015]_ ,
    \new_[41016]_ , \new_[41020]_ , \new_[41021]_ , \new_[41024]_ ,
    \new_[41027]_ , \new_[41028]_ , \new_[41029]_ , \new_[41032]_ ,
    \new_[41035]_ , \new_[41036]_ , \new_[41039]_ , \new_[41042]_ ,
    \new_[41043]_ , \new_[41044]_ , \new_[41048]_ , \new_[41049]_ ,
    \new_[41052]_ , \new_[41055]_ , \new_[41056]_ , \new_[41057]_ ,
    \new_[41060]_ , \new_[41063]_ , \new_[41064]_ , \new_[41067]_ ,
    \new_[41070]_ , \new_[41071]_ , \new_[41072]_ , \new_[41076]_ ,
    \new_[41077]_ , \new_[41080]_ , \new_[41083]_ , \new_[41084]_ ,
    \new_[41085]_ , \new_[41088]_ , \new_[41091]_ , \new_[41092]_ ,
    \new_[41095]_ , \new_[41098]_ , \new_[41099]_ , \new_[41100]_ ,
    \new_[41104]_ , \new_[41105]_ , \new_[41108]_ , \new_[41111]_ ,
    \new_[41112]_ , \new_[41113]_ , \new_[41116]_ , \new_[41119]_ ,
    \new_[41120]_ , \new_[41123]_ , \new_[41126]_ , \new_[41127]_ ,
    \new_[41128]_ , \new_[41132]_ , \new_[41133]_ , \new_[41136]_ ,
    \new_[41139]_ , \new_[41140]_ , \new_[41141]_ , \new_[41144]_ ,
    \new_[41147]_ , \new_[41148]_ , \new_[41151]_ , \new_[41154]_ ,
    \new_[41155]_ , \new_[41156]_ , \new_[41160]_ , \new_[41161]_ ,
    \new_[41164]_ , \new_[41167]_ , \new_[41168]_ , \new_[41169]_ ,
    \new_[41172]_ , \new_[41175]_ , \new_[41176]_ , \new_[41179]_ ,
    \new_[41182]_ , \new_[41183]_ , \new_[41184]_ , \new_[41188]_ ,
    \new_[41189]_ , \new_[41192]_ , \new_[41195]_ , \new_[41196]_ ,
    \new_[41197]_ , \new_[41200]_ , \new_[41203]_ , \new_[41204]_ ,
    \new_[41207]_ , \new_[41210]_ , \new_[41211]_ , \new_[41212]_ ,
    \new_[41216]_ , \new_[41217]_ , \new_[41220]_ , \new_[41223]_ ,
    \new_[41224]_ , \new_[41225]_ , \new_[41228]_ , \new_[41231]_ ,
    \new_[41232]_ , \new_[41235]_ , \new_[41238]_ , \new_[41239]_ ,
    \new_[41240]_ , \new_[41244]_ , \new_[41245]_ , \new_[41248]_ ,
    \new_[41251]_ , \new_[41252]_ , \new_[41253]_ , \new_[41256]_ ,
    \new_[41259]_ , \new_[41260]_ , \new_[41263]_ , \new_[41266]_ ,
    \new_[41267]_ , \new_[41268]_ , \new_[41272]_ , \new_[41273]_ ,
    \new_[41276]_ , \new_[41279]_ , \new_[41280]_ , \new_[41281]_ ,
    \new_[41284]_ , \new_[41287]_ , \new_[41288]_ , \new_[41291]_ ,
    \new_[41294]_ , \new_[41295]_ , \new_[41296]_ , \new_[41300]_ ,
    \new_[41301]_ , \new_[41304]_ , \new_[41307]_ , \new_[41308]_ ,
    \new_[41309]_ , \new_[41312]_ , \new_[41315]_ , \new_[41316]_ ,
    \new_[41319]_ , \new_[41322]_ , \new_[41323]_ , \new_[41324]_ ,
    \new_[41328]_ , \new_[41329]_ , \new_[41332]_ , \new_[41335]_ ,
    \new_[41336]_ , \new_[41337]_ , \new_[41340]_ , \new_[41343]_ ,
    \new_[41344]_ , \new_[41347]_ , \new_[41350]_ , \new_[41351]_ ,
    \new_[41352]_ , \new_[41356]_ , \new_[41357]_ , \new_[41360]_ ,
    \new_[41363]_ , \new_[41364]_ , \new_[41365]_ , \new_[41368]_ ,
    \new_[41371]_ , \new_[41372]_ , \new_[41375]_ , \new_[41378]_ ,
    \new_[41379]_ , \new_[41380]_ , \new_[41384]_ , \new_[41385]_ ,
    \new_[41388]_ , \new_[41391]_ , \new_[41392]_ , \new_[41393]_ ,
    \new_[41396]_ , \new_[41399]_ , \new_[41400]_ , \new_[41403]_ ,
    \new_[41406]_ , \new_[41407]_ , \new_[41408]_ , \new_[41412]_ ,
    \new_[41413]_ , \new_[41416]_ , \new_[41419]_ , \new_[41420]_ ,
    \new_[41421]_ , \new_[41424]_ , \new_[41427]_ , \new_[41428]_ ,
    \new_[41431]_ , \new_[41434]_ , \new_[41435]_ , \new_[41436]_ ,
    \new_[41440]_ , \new_[41441]_ , \new_[41444]_ , \new_[41447]_ ,
    \new_[41448]_ , \new_[41449]_ , \new_[41452]_ , \new_[41455]_ ,
    \new_[41456]_ , \new_[41459]_ , \new_[41462]_ , \new_[41463]_ ,
    \new_[41464]_ , \new_[41468]_ , \new_[41469]_ , \new_[41472]_ ,
    \new_[41475]_ , \new_[41476]_ , \new_[41477]_ , \new_[41480]_ ,
    \new_[41483]_ , \new_[41484]_ , \new_[41487]_ , \new_[41490]_ ,
    \new_[41491]_ , \new_[41492]_ , \new_[41496]_ , \new_[41497]_ ,
    \new_[41500]_ , \new_[41503]_ , \new_[41504]_ , \new_[41505]_ ,
    \new_[41508]_ , \new_[41511]_ , \new_[41512]_ , \new_[41515]_ ,
    \new_[41518]_ , \new_[41519]_ , \new_[41520]_ , \new_[41524]_ ,
    \new_[41525]_ , \new_[41528]_ , \new_[41531]_ , \new_[41532]_ ,
    \new_[41533]_ , \new_[41536]_ , \new_[41539]_ , \new_[41540]_ ,
    \new_[41543]_ , \new_[41546]_ , \new_[41547]_ , \new_[41548]_ ,
    \new_[41552]_ , \new_[41553]_ , \new_[41556]_ , \new_[41559]_ ,
    \new_[41560]_ , \new_[41561]_ , \new_[41564]_ , \new_[41567]_ ,
    \new_[41568]_ , \new_[41571]_ , \new_[41574]_ , \new_[41575]_ ,
    \new_[41576]_ , \new_[41580]_ , \new_[41581]_ , \new_[41584]_ ,
    \new_[41587]_ , \new_[41588]_ , \new_[41589]_ , \new_[41592]_ ,
    \new_[41595]_ , \new_[41596]_ , \new_[41599]_ , \new_[41602]_ ,
    \new_[41603]_ , \new_[41604]_ , \new_[41608]_ , \new_[41609]_ ,
    \new_[41612]_ , \new_[41615]_ , \new_[41616]_ , \new_[41617]_ ,
    \new_[41620]_ , \new_[41623]_ , \new_[41624]_ , \new_[41627]_ ,
    \new_[41630]_ , \new_[41631]_ , \new_[41632]_ , \new_[41636]_ ,
    \new_[41637]_ , \new_[41640]_ , \new_[41643]_ , \new_[41644]_ ,
    \new_[41645]_ , \new_[41648]_ , \new_[41651]_ , \new_[41652]_ ,
    \new_[41655]_ , \new_[41658]_ , \new_[41659]_ , \new_[41660]_ ,
    \new_[41664]_ , \new_[41665]_ , \new_[41668]_ , \new_[41671]_ ,
    \new_[41672]_ , \new_[41673]_ , \new_[41676]_ , \new_[41679]_ ,
    \new_[41680]_ , \new_[41683]_ , \new_[41686]_ , \new_[41687]_ ,
    \new_[41688]_ , \new_[41692]_ , \new_[41693]_ , \new_[41696]_ ,
    \new_[41699]_ , \new_[41700]_ , \new_[41701]_ , \new_[41704]_ ,
    \new_[41707]_ , \new_[41708]_ , \new_[41711]_ , \new_[41714]_ ,
    \new_[41715]_ , \new_[41716]_ , \new_[41720]_ , \new_[41721]_ ,
    \new_[41724]_ , \new_[41727]_ , \new_[41728]_ , \new_[41729]_ ,
    \new_[41732]_ , \new_[41735]_ , \new_[41736]_ , \new_[41739]_ ,
    \new_[41742]_ , \new_[41743]_ , \new_[41744]_ , \new_[41748]_ ,
    \new_[41749]_ , \new_[41752]_ , \new_[41755]_ , \new_[41756]_ ,
    \new_[41757]_ , \new_[41760]_ , \new_[41763]_ , \new_[41764]_ ,
    \new_[41767]_ , \new_[41770]_ , \new_[41771]_ , \new_[41772]_ ,
    \new_[41776]_ , \new_[41777]_ , \new_[41780]_ , \new_[41783]_ ,
    \new_[41784]_ , \new_[41785]_ , \new_[41788]_ , \new_[41791]_ ,
    \new_[41792]_ , \new_[41795]_ , \new_[41798]_ , \new_[41799]_ ,
    \new_[41800]_ , \new_[41804]_ , \new_[41805]_ , \new_[41808]_ ,
    \new_[41811]_ , \new_[41812]_ , \new_[41813]_ , \new_[41816]_ ,
    \new_[41819]_ , \new_[41820]_ , \new_[41823]_ , \new_[41826]_ ,
    \new_[41827]_ , \new_[41828]_ , \new_[41832]_ , \new_[41833]_ ,
    \new_[41836]_ , \new_[41839]_ , \new_[41840]_ , \new_[41841]_ ,
    \new_[41844]_ , \new_[41847]_ , \new_[41848]_ , \new_[41851]_ ,
    \new_[41854]_ , \new_[41855]_ , \new_[41856]_ , \new_[41860]_ ,
    \new_[41861]_ , \new_[41864]_ , \new_[41867]_ , \new_[41868]_ ,
    \new_[41869]_ , \new_[41872]_ , \new_[41875]_ , \new_[41876]_ ,
    \new_[41879]_ , \new_[41882]_ , \new_[41883]_ , \new_[41884]_ ,
    \new_[41888]_ , \new_[41889]_ , \new_[41892]_ , \new_[41895]_ ,
    \new_[41896]_ , \new_[41897]_ , \new_[41900]_ , \new_[41903]_ ,
    \new_[41904]_ , \new_[41907]_ , \new_[41910]_ , \new_[41911]_ ,
    \new_[41912]_ , \new_[41916]_ , \new_[41917]_ , \new_[41920]_ ,
    \new_[41923]_ , \new_[41924]_ , \new_[41925]_ , \new_[41928]_ ,
    \new_[41931]_ , \new_[41932]_ , \new_[41935]_ , \new_[41938]_ ,
    \new_[41939]_ , \new_[41940]_ , \new_[41944]_ , \new_[41945]_ ,
    \new_[41948]_ , \new_[41951]_ , \new_[41952]_ , \new_[41953]_ ,
    \new_[41956]_ , \new_[41959]_ , \new_[41960]_ , \new_[41963]_ ,
    \new_[41966]_ , \new_[41967]_ , \new_[41968]_ , \new_[41972]_ ,
    \new_[41973]_ , \new_[41976]_ , \new_[41979]_ , \new_[41980]_ ,
    \new_[41981]_ , \new_[41984]_ , \new_[41987]_ , \new_[41988]_ ,
    \new_[41991]_ , \new_[41994]_ , \new_[41995]_ , \new_[41996]_ ,
    \new_[42000]_ , \new_[42001]_ , \new_[42004]_ , \new_[42007]_ ,
    \new_[42008]_ , \new_[42009]_ , \new_[42012]_ , \new_[42015]_ ,
    \new_[42016]_ , \new_[42019]_ , \new_[42022]_ , \new_[42023]_ ,
    \new_[42024]_ , \new_[42028]_ , \new_[42029]_ , \new_[42032]_ ,
    \new_[42035]_ , \new_[42036]_ , \new_[42037]_ , \new_[42040]_ ,
    \new_[42043]_ , \new_[42044]_ , \new_[42047]_ , \new_[42050]_ ,
    \new_[42051]_ , \new_[42052]_ , \new_[42056]_ , \new_[42057]_ ,
    \new_[42060]_ , \new_[42063]_ , \new_[42064]_ , \new_[42065]_ ,
    \new_[42068]_ , \new_[42071]_ , \new_[42072]_ , \new_[42075]_ ,
    \new_[42078]_ , \new_[42079]_ , \new_[42080]_ , \new_[42084]_ ,
    \new_[42085]_ , \new_[42088]_ , \new_[42091]_ , \new_[42092]_ ,
    \new_[42093]_ , \new_[42096]_ , \new_[42099]_ , \new_[42100]_ ,
    \new_[42103]_ , \new_[42106]_ , \new_[42107]_ , \new_[42108]_ ,
    \new_[42112]_ , \new_[42113]_ , \new_[42116]_ , \new_[42119]_ ,
    \new_[42120]_ , \new_[42121]_ , \new_[42124]_ , \new_[42127]_ ,
    \new_[42128]_ , \new_[42131]_ , \new_[42134]_ , \new_[42135]_ ,
    \new_[42136]_ , \new_[42140]_ , \new_[42141]_ , \new_[42144]_ ,
    \new_[42147]_ , \new_[42148]_ , \new_[42149]_ , \new_[42152]_ ,
    \new_[42155]_ , \new_[42156]_ , \new_[42159]_ , \new_[42162]_ ,
    \new_[42163]_ , \new_[42164]_ , \new_[42168]_ , \new_[42169]_ ,
    \new_[42172]_ , \new_[42175]_ , \new_[42176]_ , \new_[42177]_ ,
    \new_[42180]_ , \new_[42183]_ , \new_[42184]_ , \new_[42187]_ ,
    \new_[42190]_ , \new_[42191]_ , \new_[42192]_ , \new_[42196]_ ,
    \new_[42197]_ , \new_[42200]_ , \new_[42203]_ , \new_[42204]_ ,
    \new_[42205]_ , \new_[42208]_ , \new_[42211]_ , \new_[42212]_ ,
    \new_[42215]_ , \new_[42218]_ , \new_[42219]_ , \new_[42220]_ ,
    \new_[42224]_ , \new_[42225]_ , \new_[42228]_ , \new_[42231]_ ,
    \new_[42232]_ , \new_[42233]_ , \new_[42236]_ , \new_[42239]_ ,
    \new_[42240]_ , \new_[42243]_ , \new_[42246]_ , \new_[42247]_ ,
    \new_[42248]_ , \new_[42252]_ , \new_[42253]_ , \new_[42256]_ ,
    \new_[42259]_ , \new_[42260]_ , \new_[42261]_ , \new_[42264]_ ,
    \new_[42267]_ , \new_[42268]_ , \new_[42271]_ , \new_[42274]_ ,
    \new_[42275]_ , \new_[42276]_ , \new_[42280]_ , \new_[42281]_ ,
    \new_[42284]_ , \new_[42287]_ , \new_[42288]_ , \new_[42289]_ ,
    \new_[42292]_ , \new_[42295]_ , \new_[42296]_ , \new_[42299]_ ,
    \new_[42302]_ , \new_[42303]_ , \new_[42304]_ , \new_[42308]_ ,
    \new_[42309]_ , \new_[42312]_ , \new_[42315]_ , \new_[42316]_ ,
    \new_[42317]_ , \new_[42320]_ , \new_[42323]_ , \new_[42324]_ ,
    \new_[42327]_ , \new_[42330]_ , \new_[42331]_ , \new_[42332]_ ,
    \new_[42336]_ , \new_[42337]_ , \new_[42340]_ , \new_[42343]_ ,
    \new_[42344]_ , \new_[42345]_ , \new_[42348]_ , \new_[42351]_ ,
    \new_[42352]_ , \new_[42355]_ , \new_[42358]_ , \new_[42359]_ ,
    \new_[42360]_ , \new_[42364]_ , \new_[42365]_ , \new_[42368]_ ,
    \new_[42371]_ , \new_[42372]_ , \new_[42373]_ , \new_[42376]_ ,
    \new_[42379]_ , \new_[42380]_ , \new_[42383]_ , \new_[42386]_ ,
    \new_[42387]_ , \new_[42388]_ , \new_[42392]_ , \new_[42393]_ ,
    \new_[42396]_ , \new_[42399]_ , \new_[42400]_ , \new_[42401]_ ,
    \new_[42404]_ , \new_[42407]_ , \new_[42408]_ , \new_[42411]_ ,
    \new_[42414]_ , \new_[42415]_ , \new_[42416]_ , \new_[42420]_ ,
    \new_[42421]_ , \new_[42424]_ , \new_[42427]_ , \new_[42428]_ ,
    \new_[42429]_ , \new_[42432]_ , \new_[42435]_ , \new_[42436]_ ,
    \new_[42439]_ , \new_[42442]_ , \new_[42443]_ , \new_[42444]_ ,
    \new_[42448]_ , \new_[42449]_ , \new_[42452]_ , \new_[42455]_ ,
    \new_[42456]_ , \new_[42457]_ , \new_[42460]_ , \new_[42463]_ ,
    \new_[42464]_ , \new_[42467]_ , \new_[42470]_ , \new_[42471]_ ,
    \new_[42472]_ , \new_[42476]_ , \new_[42477]_ , \new_[42480]_ ,
    \new_[42483]_ , \new_[42484]_ , \new_[42485]_ , \new_[42488]_ ,
    \new_[42491]_ , \new_[42492]_ , \new_[42495]_ , \new_[42498]_ ,
    \new_[42499]_ , \new_[42500]_ , \new_[42504]_ , \new_[42505]_ ,
    \new_[42508]_ , \new_[42511]_ , \new_[42512]_ , \new_[42513]_ ,
    \new_[42516]_ , \new_[42519]_ , \new_[42520]_ , \new_[42523]_ ,
    \new_[42526]_ , \new_[42527]_ , \new_[42528]_ , \new_[42532]_ ,
    \new_[42533]_ , \new_[42536]_ , \new_[42539]_ , \new_[42540]_ ,
    \new_[42541]_ , \new_[42544]_ , \new_[42547]_ , \new_[42548]_ ,
    \new_[42551]_ , \new_[42554]_ , \new_[42555]_ , \new_[42556]_ ,
    \new_[42560]_ , \new_[42561]_ , \new_[42564]_ , \new_[42567]_ ,
    \new_[42568]_ , \new_[42569]_ , \new_[42572]_ , \new_[42575]_ ,
    \new_[42576]_ , \new_[42579]_ , \new_[42582]_ , \new_[42583]_ ,
    \new_[42584]_ , \new_[42588]_ , \new_[42589]_ , \new_[42592]_ ,
    \new_[42595]_ , \new_[42596]_ , \new_[42597]_ , \new_[42600]_ ,
    \new_[42603]_ , \new_[42604]_ , \new_[42607]_ , \new_[42610]_ ,
    \new_[42611]_ , \new_[42612]_ , \new_[42616]_ , \new_[42617]_ ,
    \new_[42620]_ , \new_[42623]_ , \new_[42624]_ , \new_[42625]_ ,
    \new_[42628]_ , \new_[42631]_ , \new_[42632]_ , \new_[42635]_ ,
    \new_[42638]_ , \new_[42639]_ , \new_[42640]_ , \new_[42644]_ ,
    \new_[42645]_ , \new_[42648]_ , \new_[42651]_ , \new_[42652]_ ,
    \new_[42653]_ , \new_[42656]_ , \new_[42659]_ , \new_[42660]_ ,
    \new_[42663]_ , \new_[42666]_ , \new_[42667]_ , \new_[42668]_ ,
    \new_[42672]_ , \new_[42673]_ , \new_[42676]_ , \new_[42679]_ ,
    \new_[42680]_ , \new_[42681]_ , \new_[42684]_ , \new_[42687]_ ,
    \new_[42688]_ , \new_[42691]_ , \new_[42694]_ , \new_[42695]_ ,
    \new_[42696]_ , \new_[42700]_ , \new_[42701]_ , \new_[42704]_ ,
    \new_[42707]_ , \new_[42708]_ , \new_[42709]_ , \new_[42712]_ ,
    \new_[42715]_ , \new_[42716]_ , \new_[42719]_ , \new_[42722]_ ,
    \new_[42723]_ , \new_[42724]_ , \new_[42728]_ , \new_[42729]_ ,
    \new_[42732]_ , \new_[42735]_ , \new_[42736]_ , \new_[42737]_ ,
    \new_[42740]_ , \new_[42743]_ , \new_[42744]_ , \new_[42747]_ ,
    \new_[42750]_ , \new_[42751]_ , \new_[42752]_ , \new_[42756]_ ,
    \new_[42757]_ , \new_[42760]_ , \new_[42763]_ , \new_[42764]_ ,
    \new_[42765]_ , \new_[42768]_ , \new_[42771]_ , \new_[42772]_ ,
    \new_[42775]_ , \new_[42778]_ , \new_[42779]_ , \new_[42780]_ ,
    \new_[42784]_ , \new_[42785]_ , \new_[42788]_ , \new_[42791]_ ,
    \new_[42792]_ , \new_[42793]_ , \new_[42796]_ , \new_[42799]_ ,
    \new_[42800]_ , \new_[42803]_ , \new_[42806]_ , \new_[42807]_ ,
    \new_[42808]_ , \new_[42812]_ , \new_[42813]_ , \new_[42816]_ ,
    \new_[42819]_ , \new_[42820]_ , \new_[42821]_ , \new_[42824]_ ,
    \new_[42827]_ , \new_[42828]_ , \new_[42831]_ , \new_[42834]_ ,
    \new_[42835]_ , \new_[42836]_ , \new_[42840]_ , \new_[42841]_ ,
    \new_[42844]_ , \new_[42847]_ , \new_[42848]_ , \new_[42849]_ ,
    \new_[42852]_ , \new_[42855]_ , \new_[42856]_ , \new_[42859]_ ,
    \new_[42862]_ , \new_[42863]_ , \new_[42864]_ , \new_[42868]_ ,
    \new_[42869]_ , \new_[42872]_ , \new_[42875]_ , \new_[42876]_ ,
    \new_[42877]_ , \new_[42880]_ , \new_[42883]_ , \new_[42884]_ ,
    \new_[42887]_ , \new_[42890]_ , \new_[42891]_ , \new_[42892]_ ,
    \new_[42896]_ , \new_[42897]_ , \new_[42900]_ , \new_[42903]_ ,
    \new_[42904]_ , \new_[42905]_ , \new_[42908]_ , \new_[42911]_ ,
    \new_[42912]_ , \new_[42915]_ , \new_[42918]_ , \new_[42919]_ ,
    \new_[42920]_ , \new_[42924]_ , \new_[42925]_ , \new_[42928]_ ,
    \new_[42931]_ , \new_[42932]_ , \new_[42933]_ , \new_[42936]_ ,
    \new_[42939]_ , \new_[42940]_ , \new_[42943]_ , \new_[42946]_ ,
    \new_[42947]_ , \new_[42948]_ , \new_[42952]_ , \new_[42953]_ ,
    \new_[42956]_ , \new_[42959]_ , \new_[42960]_ , \new_[42961]_ ,
    \new_[42964]_ , \new_[42967]_ , \new_[42968]_ , \new_[42971]_ ,
    \new_[42974]_ , \new_[42975]_ , \new_[42976]_ , \new_[42980]_ ,
    \new_[42981]_ , \new_[42984]_ , \new_[42987]_ , \new_[42988]_ ,
    \new_[42989]_ , \new_[42992]_ , \new_[42995]_ , \new_[42996]_ ,
    \new_[42999]_ , \new_[43002]_ , \new_[43003]_ , \new_[43004]_ ,
    \new_[43008]_ , \new_[43009]_ , \new_[43012]_ , \new_[43015]_ ,
    \new_[43016]_ , \new_[43017]_ , \new_[43020]_ , \new_[43023]_ ,
    \new_[43024]_ , \new_[43027]_ , \new_[43030]_ , \new_[43031]_ ,
    \new_[43032]_ , \new_[43036]_ , \new_[43037]_ , \new_[43040]_ ,
    \new_[43043]_ , \new_[43044]_ , \new_[43045]_ , \new_[43048]_ ,
    \new_[43051]_ , \new_[43052]_ , \new_[43055]_ , \new_[43058]_ ,
    \new_[43059]_ , \new_[43060]_ , \new_[43064]_ , \new_[43065]_ ,
    \new_[43068]_ , \new_[43071]_ , \new_[43072]_ , \new_[43073]_ ,
    \new_[43076]_ , \new_[43079]_ , \new_[43080]_ , \new_[43083]_ ,
    \new_[43086]_ , \new_[43087]_ , \new_[43088]_ , \new_[43092]_ ,
    \new_[43093]_ , \new_[43096]_ , \new_[43099]_ , \new_[43100]_ ,
    \new_[43101]_ , \new_[43104]_ , \new_[43107]_ , \new_[43108]_ ,
    \new_[43111]_ , \new_[43114]_ , \new_[43115]_ , \new_[43116]_ ,
    \new_[43120]_ , \new_[43121]_ , \new_[43124]_ , \new_[43127]_ ,
    \new_[43128]_ , \new_[43129]_ , \new_[43132]_ , \new_[43135]_ ,
    \new_[43136]_ , \new_[43139]_ , \new_[43142]_ , \new_[43143]_ ,
    \new_[43144]_ , \new_[43148]_ , \new_[43149]_ , \new_[43152]_ ,
    \new_[43155]_ , \new_[43156]_ , \new_[43157]_ , \new_[43160]_ ,
    \new_[43163]_ , \new_[43164]_ , \new_[43167]_ , \new_[43170]_ ,
    \new_[43171]_ , \new_[43172]_ , \new_[43176]_ , \new_[43177]_ ,
    \new_[43180]_ , \new_[43183]_ , \new_[43184]_ , \new_[43185]_ ,
    \new_[43188]_ , \new_[43191]_ , \new_[43192]_ , \new_[43195]_ ,
    \new_[43198]_ , \new_[43199]_ , \new_[43200]_ , \new_[43204]_ ,
    \new_[43205]_ , \new_[43208]_ , \new_[43211]_ , \new_[43212]_ ,
    \new_[43213]_ , \new_[43216]_ , \new_[43219]_ , \new_[43220]_ ,
    \new_[43223]_ , \new_[43226]_ , \new_[43227]_ , \new_[43228]_ ,
    \new_[43232]_ , \new_[43233]_ , \new_[43236]_ , \new_[43239]_ ,
    \new_[43240]_ , \new_[43241]_ , \new_[43244]_ , \new_[43247]_ ,
    \new_[43248]_ , \new_[43251]_ , \new_[43254]_ , \new_[43255]_ ,
    \new_[43256]_ , \new_[43260]_ , \new_[43261]_ , \new_[43264]_ ,
    \new_[43267]_ , \new_[43268]_ , \new_[43269]_ , \new_[43272]_ ,
    \new_[43275]_ , \new_[43276]_ , \new_[43279]_ , \new_[43282]_ ,
    \new_[43283]_ , \new_[43284]_ , \new_[43288]_ , \new_[43289]_ ,
    \new_[43292]_ , \new_[43295]_ , \new_[43296]_ , \new_[43297]_ ,
    \new_[43300]_ , \new_[43303]_ , \new_[43304]_ , \new_[43307]_ ,
    \new_[43310]_ , \new_[43311]_ , \new_[43312]_ , \new_[43316]_ ,
    \new_[43317]_ , \new_[43320]_ , \new_[43323]_ , \new_[43324]_ ,
    \new_[43325]_ , \new_[43328]_ , \new_[43331]_ , \new_[43332]_ ,
    \new_[43335]_ , \new_[43338]_ , \new_[43339]_ , \new_[43340]_ ,
    \new_[43344]_ , \new_[43345]_ , \new_[43348]_ , \new_[43351]_ ,
    \new_[43352]_ , \new_[43353]_ , \new_[43356]_ , \new_[43359]_ ,
    \new_[43360]_ , \new_[43363]_ , \new_[43366]_ , \new_[43367]_ ,
    \new_[43368]_ , \new_[43372]_ , \new_[43373]_ , \new_[43376]_ ,
    \new_[43379]_ , \new_[43380]_ , \new_[43381]_ , \new_[43384]_ ,
    \new_[43387]_ , \new_[43388]_ , \new_[43391]_ , \new_[43394]_ ,
    \new_[43395]_ , \new_[43396]_ , \new_[43400]_ , \new_[43401]_ ,
    \new_[43404]_ , \new_[43407]_ , \new_[43408]_ , \new_[43409]_ ,
    \new_[43412]_ , \new_[43415]_ , \new_[43416]_ , \new_[43419]_ ,
    \new_[43422]_ , \new_[43423]_ , \new_[43424]_ , \new_[43428]_ ,
    \new_[43429]_ , \new_[43432]_ , \new_[43435]_ , \new_[43436]_ ,
    \new_[43437]_ , \new_[43440]_ , \new_[43443]_ , \new_[43444]_ ,
    \new_[43447]_ , \new_[43450]_ , \new_[43451]_ , \new_[43452]_ ,
    \new_[43456]_ , \new_[43457]_ , \new_[43460]_ , \new_[43463]_ ,
    \new_[43464]_ , \new_[43465]_ , \new_[43468]_ , \new_[43471]_ ,
    \new_[43472]_ , \new_[43475]_ , \new_[43478]_ , \new_[43479]_ ,
    \new_[43480]_ , \new_[43484]_ , \new_[43485]_ , \new_[43488]_ ,
    \new_[43491]_ , \new_[43492]_ , \new_[43493]_ , \new_[43496]_ ,
    \new_[43499]_ , \new_[43500]_ , \new_[43503]_ , \new_[43506]_ ,
    \new_[43507]_ , \new_[43508]_ , \new_[43512]_ , \new_[43513]_ ,
    \new_[43516]_ , \new_[43519]_ , \new_[43520]_ , \new_[43521]_ ,
    \new_[43524]_ , \new_[43527]_ , \new_[43528]_ , \new_[43531]_ ,
    \new_[43534]_ , \new_[43535]_ , \new_[43536]_ , \new_[43540]_ ,
    \new_[43541]_ , \new_[43544]_ , \new_[43547]_ , \new_[43548]_ ,
    \new_[43549]_ , \new_[43552]_ , \new_[43555]_ , \new_[43556]_ ,
    \new_[43559]_ , \new_[43562]_ , \new_[43563]_ , \new_[43564]_ ,
    \new_[43568]_ , \new_[43569]_ , \new_[43572]_ , \new_[43575]_ ,
    \new_[43576]_ , \new_[43577]_ , \new_[43580]_ , \new_[43583]_ ,
    \new_[43584]_ , \new_[43587]_ , \new_[43590]_ , \new_[43591]_ ,
    \new_[43592]_ , \new_[43596]_ , \new_[43597]_ , \new_[43600]_ ,
    \new_[43603]_ , \new_[43604]_ , \new_[43605]_ , \new_[43608]_ ,
    \new_[43611]_ , \new_[43612]_ , \new_[43615]_ , \new_[43618]_ ,
    \new_[43619]_ , \new_[43620]_ , \new_[43624]_ , \new_[43625]_ ,
    \new_[43628]_ , \new_[43631]_ , \new_[43632]_ , \new_[43633]_ ,
    \new_[43636]_ , \new_[43639]_ , \new_[43640]_ , \new_[43643]_ ,
    \new_[43646]_ , \new_[43647]_ , \new_[43648]_ , \new_[43652]_ ,
    \new_[43653]_ , \new_[43656]_ , \new_[43659]_ , \new_[43660]_ ,
    \new_[43661]_ , \new_[43664]_ , \new_[43667]_ , \new_[43668]_ ,
    \new_[43671]_ , \new_[43674]_ , \new_[43675]_ , \new_[43676]_ ,
    \new_[43680]_ , \new_[43681]_ , \new_[43684]_ , \new_[43687]_ ,
    \new_[43688]_ , \new_[43689]_ , \new_[43692]_ , \new_[43695]_ ,
    \new_[43696]_ , \new_[43699]_ , \new_[43702]_ , \new_[43703]_ ,
    \new_[43704]_ , \new_[43708]_ , \new_[43709]_ , \new_[43712]_ ,
    \new_[43715]_ , \new_[43716]_ , \new_[43717]_ , \new_[43720]_ ,
    \new_[43723]_ , \new_[43724]_ , \new_[43727]_ , \new_[43730]_ ,
    \new_[43731]_ , \new_[43732]_ , \new_[43736]_ , \new_[43737]_ ,
    \new_[43740]_ , \new_[43743]_ , \new_[43744]_ , \new_[43745]_ ,
    \new_[43748]_ , \new_[43751]_ , \new_[43752]_ , \new_[43755]_ ,
    \new_[43758]_ , \new_[43759]_ , \new_[43760]_ , \new_[43764]_ ,
    \new_[43765]_ , \new_[43768]_ , \new_[43771]_ , \new_[43772]_ ,
    \new_[43773]_ , \new_[43776]_ , \new_[43779]_ , \new_[43780]_ ,
    \new_[43783]_ , \new_[43786]_ , \new_[43787]_ , \new_[43788]_ ,
    \new_[43792]_ , \new_[43793]_ , \new_[43796]_ , \new_[43799]_ ,
    \new_[43800]_ , \new_[43801]_ , \new_[43804]_ , \new_[43807]_ ,
    \new_[43808]_ , \new_[43811]_ , \new_[43814]_ , \new_[43815]_ ,
    \new_[43816]_ , \new_[43820]_ , \new_[43821]_ , \new_[43824]_ ,
    \new_[43827]_ , \new_[43828]_ , \new_[43829]_ , \new_[43832]_ ,
    \new_[43835]_ , \new_[43836]_ , \new_[43839]_ , \new_[43842]_ ,
    \new_[43843]_ , \new_[43844]_ , \new_[43848]_ , \new_[43849]_ ,
    \new_[43852]_ , \new_[43855]_ , \new_[43856]_ , \new_[43857]_ ,
    \new_[43860]_ , \new_[43863]_ , \new_[43864]_ , \new_[43867]_ ,
    \new_[43870]_ , \new_[43871]_ , \new_[43872]_ , \new_[43876]_ ,
    \new_[43877]_ , \new_[43880]_ , \new_[43883]_ , \new_[43884]_ ,
    \new_[43885]_ , \new_[43888]_ , \new_[43891]_ , \new_[43892]_ ,
    \new_[43895]_ , \new_[43898]_ , \new_[43899]_ , \new_[43900]_ ,
    \new_[43904]_ , \new_[43905]_ , \new_[43908]_ , \new_[43911]_ ,
    \new_[43912]_ , \new_[43913]_ , \new_[43916]_ , \new_[43919]_ ,
    \new_[43920]_ , \new_[43923]_ , \new_[43926]_ , \new_[43927]_ ,
    \new_[43928]_ , \new_[43932]_ , \new_[43933]_ , \new_[43936]_ ,
    \new_[43939]_ , \new_[43940]_ , \new_[43941]_ , \new_[43944]_ ,
    \new_[43947]_ , \new_[43948]_ , \new_[43951]_ , \new_[43954]_ ,
    \new_[43955]_ , \new_[43956]_ , \new_[43960]_ , \new_[43961]_ ,
    \new_[43964]_ , \new_[43967]_ , \new_[43968]_ , \new_[43969]_ ,
    \new_[43972]_ , \new_[43975]_ , \new_[43976]_ , \new_[43979]_ ,
    \new_[43982]_ , \new_[43983]_ , \new_[43984]_ , \new_[43988]_ ,
    \new_[43989]_ , \new_[43992]_ , \new_[43995]_ , \new_[43996]_ ,
    \new_[43997]_ , \new_[44000]_ , \new_[44003]_ , \new_[44004]_ ,
    \new_[44007]_ , \new_[44010]_ , \new_[44011]_ , \new_[44012]_ ,
    \new_[44016]_ , \new_[44017]_ , \new_[44020]_ , \new_[44023]_ ,
    \new_[44024]_ , \new_[44025]_ , \new_[44028]_ , \new_[44031]_ ,
    \new_[44032]_ , \new_[44035]_ , \new_[44038]_ , \new_[44039]_ ,
    \new_[44040]_ , \new_[44044]_ , \new_[44045]_ , \new_[44048]_ ,
    \new_[44051]_ , \new_[44052]_ , \new_[44053]_ , \new_[44056]_ ,
    \new_[44059]_ , \new_[44060]_ , \new_[44063]_ , \new_[44066]_ ,
    \new_[44067]_ , \new_[44068]_ , \new_[44072]_ , \new_[44073]_ ,
    \new_[44076]_ , \new_[44079]_ , \new_[44080]_ , \new_[44081]_ ,
    \new_[44084]_ , \new_[44087]_ , \new_[44088]_ , \new_[44091]_ ,
    \new_[44094]_ , \new_[44095]_ , \new_[44096]_ , \new_[44100]_ ,
    \new_[44101]_ , \new_[44104]_ , \new_[44107]_ , \new_[44108]_ ,
    \new_[44109]_ , \new_[44112]_ , \new_[44115]_ , \new_[44116]_ ,
    \new_[44119]_ , \new_[44122]_ , \new_[44123]_ , \new_[44124]_ ,
    \new_[44128]_ , \new_[44129]_ , \new_[44132]_ , \new_[44135]_ ,
    \new_[44136]_ , \new_[44137]_ , \new_[44140]_ , \new_[44143]_ ,
    \new_[44144]_ , \new_[44147]_ , \new_[44150]_ , \new_[44151]_ ,
    \new_[44152]_ , \new_[44156]_ , \new_[44157]_ , \new_[44160]_ ,
    \new_[44163]_ , \new_[44164]_ , \new_[44165]_ , \new_[44168]_ ,
    \new_[44171]_ , \new_[44172]_ , \new_[44175]_ , \new_[44178]_ ,
    \new_[44179]_ , \new_[44180]_ , \new_[44184]_ , \new_[44185]_ ,
    \new_[44188]_ , \new_[44191]_ , \new_[44192]_ , \new_[44193]_ ,
    \new_[44196]_ , \new_[44199]_ , \new_[44200]_ , \new_[44203]_ ,
    \new_[44206]_ , \new_[44207]_ , \new_[44208]_ , \new_[44212]_ ,
    \new_[44213]_ , \new_[44216]_ , \new_[44219]_ , \new_[44220]_ ,
    \new_[44221]_ , \new_[44224]_ , \new_[44227]_ , \new_[44228]_ ,
    \new_[44231]_ , \new_[44234]_ , \new_[44235]_ , \new_[44236]_ ,
    \new_[44240]_ , \new_[44241]_ , \new_[44244]_ , \new_[44247]_ ,
    \new_[44248]_ , \new_[44249]_ , \new_[44252]_ , \new_[44255]_ ,
    \new_[44256]_ , \new_[44259]_ , \new_[44262]_ , \new_[44263]_ ,
    \new_[44264]_ , \new_[44268]_ , \new_[44269]_ , \new_[44272]_ ,
    \new_[44275]_ , \new_[44276]_ , \new_[44277]_ , \new_[44280]_ ,
    \new_[44283]_ , \new_[44284]_ , \new_[44287]_ , \new_[44290]_ ,
    \new_[44291]_ , \new_[44292]_ , \new_[44296]_ , \new_[44297]_ ,
    \new_[44300]_ , \new_[44303]_ , \new_[44304]_ , \new_[44305]_ ,
    \new_[44308]_ , \new_[44311]_ , \new_[44312]_ , \new_[44315]_ ,
    \new_[44318]_ , \new_[44319]_ , \new_[44320]_ , \new_[44324]_ ,
    \new_[44325]_ , \new_[44328]_ , \new_[44331]_ , \new_[44332]_ ,
    \new_[44333]_ , \new_[44336]_ , \new_[44339]_ , \new_[44340]_ ,
    \new_[44343]_ , \new_[44346]_ , \new_[44347]_ , \new_[44348]_ ,
    \new_[44352]_ , \new_[44353]_ , \new_[44356]_ , \new_[44359]_ ,
    \new_[44360]_ , \new_[44361]_ , \new_[44364]_ , \new_[44367]_ ,
    \new_[44368]_ , \new_[44371]_ , \new_[44374]_ , \new_[44375]_ ,
    \new_[44376]_ , \new_[44380]_ , \new_[44381]_ , \new_[44384]_ ,
    \new_[44387]_ , \new_[44388]_ , \new_[44389]_ , \new_[44392]_ ,
    \new_[44395]_ , \new_[44396]_ , \new_[44399]_ , \new_[44402]_ ,
    \new_[44403]_ , \new_[44404]_ , \new_[44408]_ , \new_[44409]_ ,
    \new_[44412]_ , \new_[44415]_ , \new_[44416]_ , \new_[44417]_ ,
    \new_[44420]_ , \new_[44423]_ , \new_[44424]_ , \new_[44427]_ ,
    \new_[44430]_ , \new_[44431]_ , \new_[44432]_ , \new_[44436]_ ,
    \new_[44437]_ , \new_[44440]_ , \new_[44443]_ , \new_[44444]_ ,
    \new_[44445]_ , \new_[44448]_ , \new_[44451]_ , \new_[44452]_ ,
    \new_[44455]_ , \new_[44458]_ , \new_[44459]_ , \new_[44460]_ ,
    \new_[44464]_ , \new_[44465]_ , \new_[44468]_ , \new_[44471]_ ,
    \new_[44472]_ , \new_[44473]_ , \new_[44476]_ , \new_[44479]_ ,
    \new_[44480]_ , \new_[44483]_ , \new_[44486]_ , \new_[44487]_ ,
    \new_[44488]_ , \new_[44492]_ , \new_[44493]_ , \new_[44496]_ ,
    \new_[44499]_ , \new_[44500]_ , \new_[44501]_ , \new_[44504]_ ,
    \new_[44507]_ , \new_[44508]_ , \new_[44511]_ , \new_[44514]_ ,
    \new_[44515]_ , \new_[44516]_ , \new_[44520]_ , \new_[44521]_ ,
    \new_[44524]_ , \new_[44527]_ , \new_[44528]_ , \new_[44529]_ ,
    \new_[44532]_ , \new_[44535]_ , \new_[44536]_ , \new_[44539]_ ,
    \new_[44542]_ , \new_[44543]_ , \new_[44544]_ , \new_[44548]_ ,
    \new_[44549]_ , \new_[44552]_ , \new_[44555]_ , \new_[44556]_ ,
    \new_[44557]_ , \new_[44560]_ , \new_[44563]_ , \new_[44564]_ ,
    \new_[44567]_ , \new_[44570]_ , \new_[44571]_ , \new_[44572]_ ,
    \new_[44576]_ , \new_[44577]_ , \new_[44580]_ , \new_[44583]_ ,
    \new_[44584]_ , \new_[44585]_ , \new_[44588]_ , \new_[44591]_ ,
    \new_[44592]_ , \new_[44595]_ , \new_[44598]_ , \new_[44599]_ ,
    \new_[44600]_ , \new_[44604]_ , \new_[44605]_ , \new_[44608]_ ,
    \new_[44611]_ , \new_[44612]_ , \new_[44613]_ , \new_[44616]_ ,
    \new_[44619]_ , \new_[44620]_ , \new_[44623]_ , \new_[44626]_ ,
    \new_[44627]_ , \new_[44628]_ , \new_[44632]_ , \new_[44633]_ ,
    \new_[44636]_ , \new_[44639]_ , \new_[44640]_ , \new_[44641]_ ,
    \new_[44644]_ , \new_[44647]_ , \new_[44648]_ , \new_[44651]_ ,
    \new_[44654]_ , \new_[44655]_ , \new_[44656]_ , \new_[44660]_ ,
    \new_[44661]_ , \new_[44664]_ , \new_[44667]_ , \new_[44668]_ ,
    \new_[44669]_ , \new_[44672]_ , \new_[44675]_ , \new_[44676]_ ,
    \new_[44679]_ , \new_[44682]_ , \new_[44683]_ , \new_[44684]_ ,
    \new_[44688]_ , \new_[44689]_ , \new_[44692]_ , \new_[44695]_ ,
    \new_[44696]_ , \new_[44697]_ , \new_[44700]_ , \new_[44703]_ ,
    \new_[44704]_ , \new_[44707]_ , \new_[44710]_ , \new_[44711]_ ,
    \new_[44712]_ , \new_[44716]_ , \new_[44717]_ , \new_[44720]_ ,
    \new_[44723]_ , \new_[44724]_ , \new_[44725]_ , \new_[44728]_ ,
    \new_[44731]_ , \new_[44732]_ , \new_[44735]_ , \new_[44738]_ ,
    \new_[44739]_ , \new_[44740]_ , \new_[44744]_ , \new_[44745]_ ,
    \new_[44748]_ , \new_[44751]_ , \new_[44752]_ , \new_[44753]_ ,
    \new_[44756]_ , \new_[44759]_ , \new_[44760]_ , \new_[44763]_ ,
    \new_[44766]_ , \new_[44767]_ , \new_[44768]_ , \new_[44772]_ ,
    \new_[44773]_ , \new_[44776]_ , \new_[44779]_ , \new_[44780]_ ,
    \new_[44781]_ , \new_[44784]_ , \new_[44787]_ , \new_[44788]_ ,
    \new_[44791]_ , \new_[44794]_ , \new_[44795]_ , \new_[44796]_ ,
    \new_[44800]_ , \new_[44801]_ , \new_[44804]_ , \new_[44807]_ ,
    \new_[44808]_ , \new_[44809]_ , \new_[44812]_ , \new_[44815]_ ,
    \new_[44816]_ , \new_[44819]_ , \new_[44822]_ , \new_[44823]_ ,
    \new_[44824]_ , \new_[44828]_ , \new_[44829]_ , \new_[44832]_ ,
    \new_[44835]_ , \new_[44836]_ , \new_[44837]_ , \new_[44840]_ ,
    \new_[44843]_ , \new_[44844]_ , \new_[44847]_ , \new_[44850]_ ,
    \new_[44851]_ , \new_[44852]_ , \new_[44856]_ , \new_[44857]_ ,
    \new_[44860]_ , \new_[44863]_ , \new_[44864]_ , \new_[44865]_ ,
    \new_[44868]_ , \new_[44871]_ , \new_[44872]_ , \new_[44875]_ ,
    \new_[44878]_ , \new_[44879]_ , \new_[44880]_ , \new_[44884]_ ,
    \new_[44885]_ , \new_[44888]_ , \new_[44891]_ , \new_[44892]_ ,
    \new_[44893]_ , \new_[44896]_ , \new_[44899]_ , \new_[44900]_ ,
    \new_[44903]_ , \new_[44906]_ , \new_[44907]_ , \new_[44908]_ ,
    \new_[44912]_ , \new_[44913]_ , \new_[44916]_ , \new_[44919]_ ,
    \new_[44920]_ , \new_[44921]_ , \new_[44924]_ , \new_[44927]_ ,
    \new_[44928]_ , \new_[44931]_ , \new_[44934]_ , \new_[44935]_ ,
    \new_[44936]_ , \new_[44940]_ , \new_[44941]_ , \new_[44944]_ ,
    \new_[44947]_ , \new_[44948]_ , \new_[44949]_ , \new_[44952]_ ,
    \new_[44955]_ , \new_[44956]_ , \new_[44959]_ , \new_[44962]_ ,
    \new_[44963]_ , \new_[44964]_ , \new_[44968]_ , \new_[44969]_ ,
    \new_[44972]_ , \new_[44975]_ , \new_[44976]_ , \new_[44977]_ ,
    \new_[44980]_ , \new_[44983]_ , \new_[44984]_ , \new_[44987]_ ,
    \new_[44990]_ , \new_[44991]_ , \new_[44992]_ , \new_[44996]_ ,
    \new_[44997]_ , \new_[45000]_ , \new_[45003]_ , \new_[45004]_ ,
    \new_[45005]_ , \new_[45008]_ , \new_[45011]_ , \new_[45012]_ ,
    \new_[45015]_ , \new_[45018]_ , \new_[45019]_ , \new_[45020]_ ,
    \new_[45024]_ , \new_[45025]_ , \new_[45028]_ , \new_[45031]_ ,
    \new_[45032]_ , \new_[45033]_ , \new_[45036]_ , \new_[45039]_ ,
    \new_[45040]_ , \new_[45043]_ , \new_[45046]_ , \new_[45047]_ ,
    \new_[45048]_ , \new_[45052]_ , \new_[45053]_ , \new_[45056]_ ,
    \new_[45059]_ , \new_[45060]_ , \new_[45061]_ , \new_[45064]_ ,
    \new_[45067]_ , \new_[45068]_ , \new_[45071]_ , \new_[45074]_ ,
    \new_[45075]_ , \new_[45076]_ , \new_[45080]_ , \new_[45081]_ ,
    \new_[45084]_ , \new_[45087]_ , \new_[45088]_ , \new_[45089]_ ,
    \new_[45092]_ , \new_[45095]_ , \new_[45096]_ , \new_[45099]_ ,
    \new_[45102]_ , \new_[45103]_ , \new_[45104]_ , \new_[45108]_ ,
    \new_[45109]_ , \new_[45112]_ , \new_[45115]_ , \new_[45116]_ ,
    \new_[45117]_ , \new_[45120]_ , \new_[45123]_ , \new_[45124]_ ,
    \new_[45127]_ , \new_[45130]_ , \new_[45131]_ , \new_[45132]_ ,
    \new_[45136]_ , \new_[45137]_ , \new_[45140]_ , \new_[45143]_ ,
    \new_[45144]_ , \new_[45145]_ , \new_[45148]_ , \new_[45151]_ ,
    \new_[45152]_ , \new_[45155]_ , \new_[45158]_ , \new_[45159]_ ,
    \new_[45160]_ , \new_[45164]_ , \new_[45165]_ , \new_[45168]_ ,
    \new_[45171]_ , \new_[45172]_ , \new_[45173]_ , \new_[45176]_ ,
    \new_[45179]_ , \new_[45180]_ , \new_[45183]_ , \new_[45186]_ ,
    \new_[45187]_ , \new_[45188]_ , \new_[45192]_ , \new_[45193]_ ,
    \new_[45196]_ , \new_[45199]_ , \new_[45200]_ , \new_[45201]_ ,
    \new_[45204]_ , \new_[45207]_ , \new_[45208]_ , \new_[45211]_ ,
    \new_[45214]_ , \new_[45215]_ , \new_[45216]_ , \new_[45220]_ ,
    \new_[45221]_ , \new_[45224]_ , \new_[45227]_ , \new_[45228]_ ,
    \new_[45229]_ , \new_[45232]_ , \new_[45235]_ , \new_[45236]_ ,
    \new_[45239]_ , \new_[45242]_ , \new_[45243]_ , \new_[45244]_ ,
    \new_[45248]_ , \new_[45249]_ , \new_[45252]_ , \new_[45255]_ ,
    \new_[45256]_ , \new_[45257]_ , \new_[45260]_ , \new_[45263]_ ,
    \new_[45264]_ , \new_[45267]_ , \new_[45270]_ , \new_[45271]_ ,
    \new_[45272]_ , \new_[45276]_ , \new_[45277]_ , \new_[45280]_ ,
    \new_[45283]_ , \new_[45284]_ , \new_[45285]_ , \new_[45288]_ ,
    \new_[45291]_ , \new_[45292]_ , \new_[45295]_ , \new_[45298]_ ,
    \new_[45299]_ , \new_[45300]_ , \new_[45303]_ , \new_[45306]_ ,
    \new_[45307]_ , \new_[45310]_ , \new_[45313]_ , \new_[45314]_ ,
    \new_[45315]_ , \new_[45318]_ , \new_[45321]_ , \new_[45322]_ ,
    \new_[45325]_ , \new_[45328]_ , \new_[45329]_ , \new_[45330]_ ,
    \new_[45333]_ , \new_[45336]_ , \new_[45337]_ , \new_[45340]_ ,
    \new_[45343]_ , \new_[45344]_ , \new_[45345]_ , \new_[45348]_ ,
    \new_[45351]_ , \new_[45352]_ , \new_[45355]_ , \new_[45358]_ ,
    \new_[45359]_ , \new_[45360]_ , \new_[45363]_ , \new_[45366]_ ,
    \new_[45367]_ , \new_[45370]_ , \new_[45373]_ , \new_[45374]_ ,
    \new_[45375]_ , \new_[45378]_ , \new_[45381]_ , \new_[45382]_ ,
    \new_[45385]_ , \new_[45388]_ , \new_[45389]_ , \new_[45390]_ ,
    \new_[45393]_ , \new_[45396]_ , \new_[45397]_ , \new_[45400]_ ,
    \new_[45403]_ , \new_[45404]_ , \new_[45405]_ , \new_[45408]_ ,
    \new_[45411]_ , \new_[45412]_ , \new_[45415]_ , \new_[45418]_ ,
    \new_[45419]_ , \new_[45420]_ , \new_[45423]_ , \new_[45426]_ ,
    \new_[45427]_ , \new_[45430]_ , \new_[45433]_ , \new_[45434]_ ,
    \new_[45435]_ , \new_[45438]_ , \new_[45441]_ , \new_[45442]_ ,
    \new_[45445]_ , \new_[45448]_ , \new_[45449]_ , \new_[45450]_ ,
    \new_[45453]_ , \new_[45456]_ , \new_[45457]_ , \new_[45460]_ ,
    \new_[45463]_ , \new_[45464]_ , \new_[45465]_ , \new_[45468]_ ,
    \new_[45471]_ , \new_[45472]_ , \new_[45475]_ , \new_[45478]_ ,
    \new_[45479]_ , \new_[45480]_ , \new_[45483]_ , \new_[45486]_ ,
    \new_[45487]_ , \new_[45490]_ , \new_[45493]_ , \new_[45494]_ ,
    \new_[45495]_ , \new_[45498]_ , \new_[45501]_ , \new_[45502]_ ,
    \new_[45505]_ , \new_[45508]_ , \new_[45509]_ , \new_[45510]_ ,
    \new_[45513]_ , \new_[45516]_ , \new_[45517]_ , \new_[45520]_ ,
    \new_[45523]_ , \new_[45524]_ , \new_[45525]_ , \new_[45528]_ ,
    \new_[45531]_ , \new_[45532]_ , \new_[45535]_ , \new_[45538]_ ,
    \new_[45539]_ , \new_[45540]_ , \new_[45543]_ , \new_[45546]_ ,
    \new_[45547]_ , \new_[45550]_ , \new_[45553]_ , \new_[45554]_ ,
    \new_[45555]_ , \new_[45558]_ , \new_[45561]_ , \new_[45562]_ ,
    \new_[45565]_ , \new_[45568]_ , \new_[45569]_ , \new_[45570]_ ,
    \new_[45573]_ , \new_[45576]_ , \new_[45577]_ , \new_[45580]_ ,
    \new_[45583]_ , \new_[45584]_ , \new_[45585]_ , \new_[45588]_ ,
    \new_[45591]_ , \new_[45592]_ , \new_[45595]_ , \new_[45598]_ ,
    \new_[45599]_ , \new_[45600]_ , \new_[45603]_ , \new_[45606]_ ,
    \new_[45607]_ , \new_[45610]_ , \new_[45613]_ , \new_[45614]_ ,
    \new_[45615]_ , \new_[45618]_ , \new_[45621]_ , \new_[45622]_ ,
    \new_[45625]_ , \new_[45628]_ , \new_[45629]_ , \new_[45630]_ ,
    \new_[45633]_ , \new_[45636]_ , \new_[45637]_ , \new_[45640]_ ,
    \new_[45643]_ , \new_[45644]_ , \new_[45645]_ , \new_[45648]_ ,
    \new_[45651]_ , \new_[45652]_ , \new_[45655]_ , \new_[45658]_ ,
    \new_[45659]_ , \new_[45660]_ , \new_[45663]_ , \new_[45666]_ ,
    \new_[45667]_ , \new_[45670]_ , \new_[45673]_ , \new_[45674]_ ,
    \new_[45675]_ , \new_[45678]_ , \new_[45681]_ , \new_[45682]_ ,
    \new_[45685]_ , \new_[45688]_ , \new_[45689]_ , \new_[45690]_ ,
    \new_[45693]_ , \new_[45696]_ , \new_[45697]_ , \new_[45700]_ ,
    \new_[45703]_ , \new_[45704]_ , \new_[45705]_ , \new_[45708]_ ,
    \new_[45711]_ , \new_[45712]_ , \new_[45715]_ , \new_[45718]_ ,
    \new_[45719]_ , \new_[45720]_ , \new_[45723]_ , \new_[45726]_ ,
    \new_[45727]_ , \new_[45730]_ , \new_[45733]_ , \new_[45734]_ ,
    \new_[45735]_ , \new_[45738]_ , \new_[45741]_ , \new_[45742]_ ,
    \new_[45745]_ , \new_[45748]_ , \new_[45749]_ , \new_[45750]_ ,
    \new_[45753]_ , \new_[45756]_ , \new_[45757]_ , \new_[45760]_ ,
    \new_[45763]_ , \new_[45764]_ , \new_[45765]_ , \new_[45768]_ ,
    \new_[45771]_ , \new_[45772]_ , \new_[45775]_ , \new_[45778]_ ,
    \new_[45779]_ , \new_[45780]_ , \new_[45783]_ , \new_[45786]_ ,
    \new_[45787]_ , \new_[45790]_ , \new_[45793]_ , \new_[45794]_ ,
    \new_[45795]_ , \new_[45798]_ , \new_[45801]_ , \new_[45802]_ ,
    \new_[45805]_ , \new_[45808]_ , \new_[45809]_ , \new_[45810]_ ,
    \new_[45813]_ , \new_[45816]_ , \new_[45817]_ , \new_[45820]_ ,
    \new_[45823]_ , \new_[45824]_ , \new_[45825]_ , \new_[45828]_ ,
    \new_[45831]_ , \new_[45832]_ , \new_[45835]_ , \new_[45838]_ ,
    \new_[45839]_ , \new_[45840]_ , \new_[45843]_ , \new_[45846]_ ,
    \new_[45847]_ , \new_[45850]_ , \new_[45853]_ , \new_[45854]_ ,
    \new_[45855]_ , \new_[45858]_ , \new_[45861]_ , \new_[45862]_ ,
    \new_[45865]_ , \new_[45868]_ , \new_[45869]_ , \new_[45870]_ ,
    \new_[45873]_ , \new_[45876]_ , \new_[45877]_ , \new_[45880]_ ,
    \new_[45883]_ , \new_[45884]_ , \new_[45885]_ , \new_[45888]_ ,
    \new_[45891]_ , \new_[45892]_ , \new_[45895]_ , \new_[45898]_ ,
    \new_[45899]_ , \new_[45900]_ , \new_[45903]_ , \new_[45906]_ ,
    \new_[45907]_ , \new_[45910]_ , \new_[45913]_ , \new_[45914]_ ,
    \new_[45915]_ , \new_[45918]_ , \new_[45921]_ , \new_[45922]_ ,
    \new_[45925]_ , \new_[45928]_ , \new_[45929]_ , \new_[45930]_ ,
    \new_[45933]_ , \new_[45936]_ , \new_[45937]_ , \new_[45940]_ ,
    \new_[45943]_ , \new_[45944]_ , \new_[45945]_ , \new_[45948]_ ,
    \new_[45951]_ , \new_[45952]_ , \new_[45955]_ , \new_[45958]_ ,
    \new_[45959]_ , \new_[45960]_ , \new_[45963]_ , \new_[45966]_ ,
    \new_[45967]_ , \new_[45970]_ , \new_[45973]_ , \new_[45974]_ ,
    \new_[45975]_ , \new_[45978]_ , \new_[45981]_ , \new_[45982]_ ,
    \new_[45985]_ , \new_[45988]_ , \new_[45989]_ , \new_[45990]_ ,
    \new_[45993]_ , \new_[45996]_ , \new_[45997]_ , \new_[46000]_ ,
    \new_[46003]_ , \new_[46004]_ , \new_[46005]_ , \new_[46008]_ ,
    \new_[46011]_ , \new_[46012]_ , \new_[46015]_ , \new_[46018]_ ,
    \new_[46019]_ , \new_[46020]_ , \new_[46023]_ , \new_[46026]_ ,
    \new_[46027]_ , \new_[46030]_ , \new_[46033]_ , \new_[46034]_ ,
    \new_[46035]_ , \new_[46038]_ , \new_[46041]_ , \new_[46042]_ ,
    \new_[46045]_ , \new_[46048]_ , \new_[46049]_ , \new_[46050]_ ,
    \new_[46053]_ , \new_[46056]_ , \new_[46057]_ , \new_[46060]_ ,
    \new_[46063]_ , \new_[46064]_ , \new_[46065]_ , \new_[46068]_ ,
    \new_[46071]_ , \new_[46072]_ , \new_[46075]_ , \new_[46078]_ ,
    \new_[46079]_ , \new_[46080]_ , \new_[46083]_ , \new_[46086]_ ,
    \new_[46087]_ , \new_[46090]_ , \new_[46093]_ , \new_[46094]_ ,
    \new_[46095]_ , \new_[46098]_ , \new_[46101]_ , \new_[46102]_ ,
    \new_[46105]_ , \new_[46108]_ , \new_[46109]_ , \new_[46110]_ ,
    \new_[46113]_ , \new_[46116]_ , \new_[46117]_ , \new_[46120]_ ,
    \new_[46123]_ , \new_[46124]_ , \new_[46125]_ , \new_[46128]_ ,
    \new_[46131]_ , \new_[46132]_ , \new_[46135]_ , \new_[46138]_ ,
    \new_[46139]_ , \new_[46140]_ , \new_[46143]_ , \new_[46146]_ ,
    \new_[46147]_ , \new_[46150]_ , \new_[46153]_ , \new_[46154]_ ,
    \new_[46155]_ , \new_[46158]_ , \new_[46161]_ , \new_[46162]_ ,
    \new_[46165]_ , \new_[46168]_ , \new_[46169]_ , \new_[46170]_ ,
    \new_[46173]_ , \new_[46176]_ , \new_[46177]_ , \new_[46180]_ ,
    \new_[46183]_ , \new_[46184]_ , \new_[46185]_ , \new_[46188]_ ,
    \new_[46191]_ , \new_[46192]_ , \new_[46195]_ , \new_[46198]_ ,
    \new_[46199]_ , \new_[46200]_ , \new_[46203]_ , \new_[46206]_ ,
    \new_[46207]_ , \new_[46210]_ , \new_[46213]_ , \new_[46214]_ ,
    \new_[46215]_ , \new_[46218]_ , \new_[46221]_ , \new_[46222]_ ,
    \new_[46225]_ , \new_[46228]_ , \new_[46229]_ , \new_[46230]_ ,
    \new_[46233]_ , \new_[46236]_ , \new_[46237]_ , \new_[46240]_ ,
    \new_[46243]_ , \new_[46244]_ , \new_[46245]_ , \new_[46248]_ ,
    \new_[46251]_ , \new_[46252]_ , \new_[46255]_ , \new_[46258]_ ,
    \new_[46259]_ , \new_[46260]_ , \new_[46263]_ , \new_[46266]_ ,
    \new_[46267]_ , \new_[46270]_ , \new_[46273]_ , \new_[46274]_ ,
    \new_[46275]_ , \new_[46278]_ , \new_[46281]_ , \new_[46282]_ ,
    \new_[46285]_ , \new_[46288]_ , \new_[46289]_ , \new_[46290]_ ,
    \new_[46293]_ , \new_[46296]_ , \new_[46297]_ , \new_[46300]_ ,
    \new_[46303]_ , \new_[46304]_ , \new_[46305]_ , \new_[46308]_ ,
    \new_[46311]_ , \new_[46312]_ , \new_[46315]_ , \new_[46318]_ ,
    \new_[46319]_ , \new_[46320]_ , \new_[46323]_ , \new_[46326]_ ,
    \new_[46327]_ , \new_[46330]_ , \new_[46333]_ , \new_[46334]_ ,
    \new_[46335]_ , \new_[46338]_ , \new_[46341]_ , \new_[46342]_ ,
    \new_[46345]_ , \new_[46348]_ , \new_[46349]_ , \new_[46350]_ ,
    \new_[46353]_ , \new_[46356]_ , \new_[46357]_ , \new_[46360]_ ,
    \new_[46363]_ , \new_[46364]_ , \new_[46365]_ , \new_[46368]_ ,
    \new_[46371]_ , \new_[46372]_ , \new_[46375]_ , \new_[46378]_ ,
    \new_[46379]_ , \new_[46380]_ , \new_[46383]_ , \new_[46386]_ ,
    \new_[46387]_ , \new_[46390]_ , \new_[46393]_ , \new_[46394]_ ,
    \new_[46395]_ , \new_[46398]_ , \new_[46401]_ , \new_[46402]_ ,
    \new_[46405]_ , \new_[46408]_ , \new_[46409]_ , \new_[46410]_ ,
    \new_[46413]_ , \new_[46416]_ , \new_[46417]_ , \new_[46420]_ ,
    \new_[46423]_ , \new_[46424]_ , \new_[46425]_ , \new_[46428]_ ,
    \new_[46431]_ , \new_[46432]_ , \new_[46435]_ , \new_[46438]_ ,
    \new_[46439]_ , \new_[46440]_ , \new_[46443]_ , \new_[46446]_ ,
    \new_[46447]_ , \new_[46450]_ , \new_[46453]_ , \new_[46454]_ ,
    \new_[46455]_ , \new_[46458]_ , \new_[46461]_ , \new_[46462]_ ,
    \new_[46465]_ , \new_[46468]_ , \new_[46469]_ , \new_[46470]_ ,
    \new_[46473]_ , \new_[46476]_ , \new_[46477]_ , \new_[46480]_ ,
    \new_[46483]_ , \new_[46484]_ , \new_[46485]_ , \new_[46488]_ ,
    \new_[46491]_ , \new_[46492]_ , \new_[46495]_ , \new_[46498]_ ,
    \new_[46499]_ , \new_[46500]_ , \new_[46503]_ , \new_[46506]_ ,
    \new_[46507]_ , \new_[46510]_ , \new_[46513]_ , \new_[46514]_ ,
    \new_[46515]_ , \new_[46518]_ , \new_[46521]_ , \new_[46522]_ ,
    \new_[46525]_ , \new_[46528]_ , \new_[46529]_ , \new_[46530]_ ,
    \new_[46533]_ , \new_[46536]_ , \new_[46537]_ , \new_[46540]_ ,
    \new_[46543]_ , \new_[46544]_ , \new_[46545]_ , \new_[46548]_ ,
    \new_[46551]_ , \new_[46552]_ , \new_[46555]_ , \new_[46558]_ ,
    \new_[46559]_ , \new_[46560]_ , \new_[46563]_ , \new_[46566]_ ,
    \new_[46567]_ , \new_[46570]_ , \new_[46573]_ , \new_[46574]_ ,
    \new_[46575]_ , \new_[46578]_ , \new_[46581]_ , \new_[46582]_ ,
    \new_[46585]_ , \new_[46588]_ , \new_[46589]_ , \new_[46590]_ ,
    \new_[46593]_ , \new_[46596]_ , \new_[46597]_ , \new_[46600]_ ,
    \new_[46603]_ , \new_[46604]_ , \new_[46605]_ , \new_[46608]_ ,
    \new_[46611]_ , \new_[46612]_ , \new_[46615]_ , \new_[46618]_ ,
    \new_[46619]_ , \new_[46620]_ , \new_[46623]_ , \new_[46626]_ ,
    \new_[46627]_ , \new_[46630]_ , \new_[46633]_ , \new_[46634]_ ,
    \new_[46635]_ , \new_[46638]_ , \new_[46641]_ , \new_[46642]_ ,
    \new_[46645]_ , \new_[46648]_ , \new_[46649]_ , \new_[46650]_ ,
    \new_[46653]_ , \new_[46656]_ , \new_[46657]_ , \new_[46660]_ ,
    \new_[46663]_ , \new_[46664]_ , \new_[46665]_ , \new_[46668]_ ,
    \new_[46671]_ , \new_[46672]_ , \new_[46675]_ , \new_[46678]_ ,
    \new_[46679]_ , \new_[46680]_ , \new_[46683]_ , \new_[46686]_ ,
    \new_[46687]_ , \new_[46690]_ , \new_[46693]_ , \new_[46694]_ ,
    \new_[46695]_ , \new_[46698]_ , \new_[46701]_ , \new_[46702]_ ,
    \new_[46705]_ , \new_[46708]_ , \new_[46709]_ , \new_[46710]_ ,
    \new_[46713]_ , \new_[46716]_ , \new_[46717]_ , \new_[46720]_ ,
    \new_[46723]_ , \new_[46724]_ , \new_[46725]_ , \new_[46728]_ ,
    \new_[46731]_ , \new_[46732]_ , \new_[46735]_ , \new_[46738]_ ,
    \new_[46739]_ , \new_[46740]_ , \new_[46743]_ , \new_[46746]_ ,
    \new_[46747]_ , \new_[46750]_ , \new_[46753]_ , \new_[46754]_ ,
    \new_[46755]_ , \new_[46758]_ , \new_[46761]_ , \new_[46762]_ ,
    \new_[46765]_ , \new_[46768]_ , \new_[46769]_ , \new_[46770]_ ,
    \new_[46773]_ , \new_[46776]_ , \new_[46777]_ , \new_[46780]_ ,
    \new_[46783]_ , \new_[46784]_ , \new_[46785]_ , \new_[46788]_ ,
    \new_[46791]_ , \new_[46792]_ , \new_[46795]_ , \new_[46798]_ ,
    \new_[46799]_ , \new_[46800]_ , \new_[46803]_ , \new_[46806]_ ,
    \new_[46807]_ , \new_[46810]_ , \new_[46813]_ , \new_[46814]_ ,
    \new_[46815]_ , \new_[46818]_ , \new_[46821]_ , \new_[46822]_ ,
    \new_[46825]_ , \new_[46828]_ , \new_[46829]_ , \new_[46830]_ ,
    \new_[46833]_ , \new_[46836]_ , \new_[46837]_ , \new_[46840]_ ,
    \new_[46843]_ , \new_[46844]_ , \new_[46845]_ , \new_[46848]_ ,
    \new_[46851]_ , \new_[46852]_ , \new_[46855]_ , \new_[46858]_ ,
    \new_[46859]_ , \new_[46860]_ , \new_[46863]_ , \new_[46866]_ ,
    \new_[46867]_ , \new_[46870]_ , \new_[46873]_ , \new_[46874]_ ,
    \new_[46875]_ , \new_[46878]_ , \new_[46881]_ , \new_[46882]_ ,
    \new_[46885]_ , \new_[46888]_ , \new_[46889]_ , \new_[46890]_ ,
    \new_[46893]_ , \new_[46896]_ , \new_[46897]_ , \new_[46900]_ ,
    \new_[46903]_ , \new_[46904]_ , \new_[46905]_ , \new_[46908]_ ,
    \new_[46911]_ , \new_[46912]_ , \new_[46915]_ , \new_[46918]_ ,
    \new_[46919]_ , \new_[46920]_ , \new_[46923]_ , \new_[46926]_ ,
    \new_[46927]_ , \new_[46930]_ , \new_[46933]_ , \new_[46934]_ ,
    \new_[46935]_ , \new_[46938]_ , \new_[46941]_ , \new_[46942]_ ,
    \new_[46945]_ , \new_[46948]_ , \new_[46949]_ , \new_[46950]_ ,
    \new_[46953]_ , \new_[46956]_ , \new_[46957]_ , \new_[46960]_ ,
    \new_[46963]_ , \new_[46964]_ , \new_[46965]_ , \new_[46968]_ ,
    \new_[46971]_ , \new_[46972]_ , \new_[46975]_ , \new_[46978]_ ,
    \new_[46979]_ , \new_[46980]_ , \new_[46983]_ , \new_[46986]_ ,
    \new_[46987]_ , \new_[46990]_ , \new_[46993]_ , \new_[46994]_ ,
    \new_[46995]_ , \new_[46998]_ , \new_[47001]_ , \new_[47002]_ ,
    \new_[47005]_ , \new_[47008]_ , \new_[47009]_ , \new_[47010]_ ,
    \new_[47013]_ , \new_[47016]_ , \new_[47017]_ , \new_[47020]_ ,
    \new_[47023]_ , \new_[47024]_ , \new_[47025]_ , \new_[47028]_ ,
    \new_[47031]_ , \new_[47032]_ , \new_[47035]_ , \new_[47038]_ ,
    \new_[47039]_ , \new_[47040]_ , \new_[47043]_ , \new_[47046]_ ,
    \new_[47047]_ , \new_[47050]_ , \new_[47053]_ , \new_[47054]_ ,
    \new_[47055]_ , \new_[47058]_ , \new_[47061]_ , \new_[47062]_ ,
    \new_[47065]_ , \new_[47068]_ , \new_[47069]_ , \new_[47070]_ ,
    \new_[47073]_ , \new_[47076]_ , \new_[47077]_ , \new_[47080]_ ,
    \new_[47083]_ , \new_[47084]_ , \new_[47085]_ , \new_[47088]_ ,
    \new_[47091]_ , \new_[47092]_ , \new_[47095]_ , \new_[47098]_ ,
    \new_[47099]_ , \new_[47100]_ , \new_[47103]_ , \new_[47106]_ ,
    \new_[47107]_ , \new_[47110]_ , \new_[47113]_ , \new_[47114]_ ,
    \new_[47115]_ , \new_[47118]_ , \new_[47121]_ , \new_[47122]_ ,
    \new_[47125]_ , \new_[47128]_ , \new_[47129]_ , \new_[47130]_ ,
    \new_[47133]_ , \new_[47136]_ , \new_[47137]_ , \new_[47140]_ ,
    \new_[47143]_ , \new_[47144]_ , \new_[47145]_ , \new_[47148]_ ,
    \new_[47151]_ , \new_[47152]_ , \new_[47155]_ , \new_[47158]_ ,
    \new_[47159]_ , \new_[47160]_ , \new_[47163]_ , \new_[47166]_ ,
    \new_[47167]_ , \new_[47170]_ , \new_[47173]_ , \new_[47174]_ ,
    \new_[47175]_ , \new_[47178]_ , \new_[47181]_ , \new_[47182]_ ,
    \new_[47185]_ , \new_[47188]_ , \new_[47189]_ , \new_[47190]_ ,
    \new_[47193]_ , \new_[47196]_ , \new_[47197]_ , \new_[47200]_ ,
    \new_[47203]_ , \new_[47204]_ , \new_[47205]_ , \new_[47208]_ ,
    \new_[47211]_ , \new_[47212]_ , \new_[47215]_ , \new_[47218]_ ,
    \new_[47219]_ , \new_[47220]_ , \new_[47223]_ , \new_[47226]_ ,
    \new_[47227]_ , \new_[47230]_ , \new_[47233]_ , \new_[47234]_ ,
    \new_[47235]_ , \new_[47238]_ , \new_[47241]_ , \new_[47242]_ ,
    \new_[47245]_ , \new_[47248]_ , \new_[47249]_ , \new_[47250]_ ,
    \new_[47253]_ , \new_[47256]_ , \new_[47257]_ , \new_[47260]_ ,
    \new_[47263]_ , \new_[47264]_ , \new_[47265]_ , \new_[47268]_ ,
    \new_[47271]_ , \new_[47272]_ , \new_[47275]_ , \new_[47278]_ ,
    \new_[47279]_ , \new_[47280]_ , \new_[47283]_ , \new_[47286]_ ,
    \new_[47287]_ , \new_[47290]_ , \new_[47293]_ , \new_[47294]_ ,
    \new_[47295]_ , \new_[47298]_ , \new_[47301]_ , \new_[47302]_ ,
    \new_[47305]_ , \new_[47308]_ , \new_[47309]_ , \new_[47310]_ ,
    \new_[47313]_ , \new_[47316]_ , \new_[47317]_ , \new_[47320]_ ,
    \new_[47323]_ , \new_[47324]_ , \new_[47325]_ , \new_[47328]_ ,
    \new_[47331]_ , \new_[47332]_ , \new_[47335]_ , \new_[47338]_ ,
    \new_[47339]_ , \new_[47340]_ , \new_[47343]_ , \new_[47346]_ ,
    \new_[47347]_ , \new_[47350]_ , \new_[47353]_ , \new_[47354]_ ,
    \new_[47355]_ , \new_[47358]_ , \new_[47361]_ , \new_[47362]_ ,
    \new_[47365]_ , \new_[47368]_ , \new_[47369]_ , \new_[47370]_ ,
    \new_[47373]_ , \new_[47376]_ , \new_[47377]_ , \new_[47380]_ ,
    \new_[47383]_ , \new_[47384]_ , \new_[47385]_ , \new_[47388]_ ,
    \new_[47391]_ , \new_[47392]_ , \new_[47395]_ , \new_[47398]_ ,
    \new_[47399]_ , \new_[47400]_ , \new_[47403]_ , \new_[47406]_ ,
    \new_[47407]_ , \new_[47410]_ , \new_[47413]_ , \new_[47414]_ ,
    \new_[47415]_ , \new_[47418]_ , \new_[47421]_ , \new_[47422]_ ,
    \new_[47425]_ , \new_[47428]_ , \new_[47429]_ , \new_[47430]_ ,
    \new_[47433]_ , \new_[47436]_ , \new_[47437]_ , \new_[47440]_ ,
    \new_[47443]_ , \new_[47444]_ , \new_[47445]_ , \new_[47448]_ ,
    \new_[47451]_ , \new_[47452]_ , \new_[47455]_ , \new_[47458]_ ,
    \new_[47459]_ , \new_[47460]_ , \new_[47463]_ , \new_[47466]_ ,
    \new_[47467]_ , \new_[47470]_ , \new_[47473]_ , \new_[47474]_ ,
    \new_[47475]_ , \new_[47478]_ , \new_[47481]_ , \new_[47482]_ ,
    \new_[47485]_ , \new_[47488]_ , \new_[47489]_ , \new_[47490]_ ,
    \new_[47493]_ , \new_[47496]_ , \new_[47497]_ , \new_[47500]_ ,
    \new_[47503]_ , \new_[47504]_ , \new_[47505]_ , \new_[47508]_ ,
    \new_[47511]_ , \new_[47512]_ , \new_[47515]_ , \new_[47518]_ ,
    \new_[47519]_ , \new_[47520]_ , \new_[47523]_ , \new_[47526]_ ,
    \new_[47527]_ , \new_[47530]_ , \new_[47533]_ , \new_[47534]_ ,
    \new_[47535]_ , \new_[47538]_ , \new_[47541]_ , \new_[47542]_ ,
    \new_[47545]_ , \new_[47548]_ , \new_[47549]_ , \new_[47550]_ ,
    \new_[47553]_ , \new_[47556]_ , \new_[47557]_ , \new_[47560]_ ,
    \new_[47563]_ , \new_[47564]_ , \new_[47565]_ , \new_[47568]_ ,
    \new_[47571]_ , \new_[47572]_ , \new_[47575]_ , \new_[47578]_ ,
    \new_[47579]_ , \new_[47580]_ , \new_[47583]_ , \new_[47586]_ ,
    \new_[47587]_ , \new_[47590]_ , \new_[47593]_ , \new_[47594]_ ,
    \new_[47595]_ , \new_[47598]_ , \new_[47601]_ , \new_[47602]_ ,
    \new_[47605]_ , \new_[47608]_ , \new_[47609]_ , \new_[47610]_ ,
    \new_[47613]_ , \new_[47616]_ , \new_[47617]_ , \new_[47620]_ ,
    \new_[47623]_ , \new_[47624]_ , \new_[47625]_ , \new_[47628]_ ,
    \new_[47631]_ , \new_[47632]_ , \new_[47635]_ , \new_[47638]_ ,
    \new_[47639]_ , \new_[47640]_ , \new_[47643]_ , \new_[47646]_ ,
    \new_[47647]_ , \new_[47650]_ , \new_[47653]_ , \new_[47654]_ ,
    \new_[47655]_ , \new_[47658]_ , \new_[47661]_ , \new_[47662]_ ,
    \new_[47665]_ , \new_[47668]_ , \new_[47669]_ , \new_[47670]_ ,
    \new_[47673]_ , \new_[47676]_ , \new_[47677]_ , \new_[47680]_ ,
    \new_[47683]_ , \new_[47684]_ , \new_[47685]_ , \new_[47688]_ ,
    \new_[47691]_ , \new_[47692]_ , \new_[47695]_ , \new_[47698]_ ,
    \new_[47699]_ , \new_[47700]_ , \new_[47703]_ , \new_[47706]_ ,
    \new_[47707]_ , \new_[47710]_ , \new_[47713]_ , \new_[47714]_ ,
    \new_[47715]_ , \new_[47718]_ , \new_[47721]_ , \new_[47722]_ ,
    \new_[47725]_ , \new_[47728]_ , \new_[47729]_ , \new_[47730]_ ,
    \new_[47733]_ , \new_[47736]_ , \new_[47737]_ , \new_[47740]_ ,
    \new_[47743]_ , \new_[47744]_ , \new_[47745]_ , \new_[47748]_ ,
    \new_[47751]_ , \new_[47752]_ , \new_[47755]_ , \new_[47758]_ ,
    \new_[47759]_ , \new_[47760]_ , \new_[47763]_ , \new_[47766]_ ,
    \new_[47767]_ , \new_[47770]_ , \new_[47773]_ , \new_[47774]_ ,
    \new_[47775]_ , \new_[47778]_ , \new_[47781]_ , \new_[47782]_ ,
    \new_[47785]_ , \new_[47788]_ , \new_[47789]_ , \new_[47790]_ ,
    \new_[47793]_ , \new_[47796]_ , \new_[47797]_ , \new_[47800]_ ,
    \new_[47803]_ , \new_[47804]_ , \new_[47805]_ , \new_[47808]_ ,
    \new_[47811]_ , \new_[47812]_ , \new_[47815]_ , \new_[47818]_ ,
    \new_[47819]_ , \new_[47820]_ , \new_[47823]_ , \new_[47826]_ ,
    \new_[47827]_ , \new_[47830]_ , \new_[47833]_ , \new_[47834]_ ,
    \new_[47835]_ , \new_[47838]_ , \new_[47841]_ , \new_[47842]_ ,
    \new_[47845]_ , \new_[47848]_ , \new_[47849]_ , \new_[47850]_ ,
    \new_[47853]_ , \new_[47856]_ , \new_[47857]_ , \new_[47860]_ ,
    \new_[47863]_ , \new_[47864]_ , \new_[47865]_ , \new_[47868]_ ,
    \new_[47871]_ , \new_[47872]_ , \new_[47875]_ , \new_[47878]_ ,
    \new_[47879]_ , \new_[47880]_ , \new_[47883]_ , \new_[47886]_ ,
    \new_[47887]_ , \new_[47890]_ , \new_[47893]_ , \new_[47894]_ ,
    \new_[47895]_ , \new_[47898]_ , \new_[47901]_ , \new_[47902]_ ,
    \new_[47905]_ , \new_[47908]_ , \new_[47909]_ , \new_[47910]_ ,
    \new_[47913]_ , \new_[47916]_ , \new_[47917]_ , \new_[47920]_ ,
    \new_[47923]_ , \new_[47924]_ , \new_[47925]_ , \new_[47928]_ ,
    \new_[47931]_ , \new_[47932]_ , \new_[47935]_ , \new_[47938]_ ,
    \new_[47939]_ , \new_[47940]_ , \new_[47943]_ , \new_[47946]_ ,
    \new_[47947]_ , \new_[47950]_ , \new_[47953]_ , \new_[47954]_ ,
    \new_[47955]_ , \new_[47958]_ , \new_[47961]_ , \new_[47962]_ ,
    \new_[47965]_ , \new_[47968]_ , \new_[47969]_ , \new_[47970]_ ,
    \new_[47973]_ , \new_[47976]_ , \new_[47977]_ , \new_[47980]_ ,
    \new_[47983]_ , \new_[47984]_ , \new_[47985]_ , \new_[47988]_ ,
    \new_[47991]_ , \new_[47992]_ , \new_[47995]_ , \new_[47998]_ ,
    \new_[47999]_ , \new_[48000]_ , \new_[48003]_ , \new_[48006]_ ,
    \new_[48007]_ , \new_[48010]_ , \new_[48013]_ , \new_[48014]_ ,
    \new_[48015]_ , \new_[48018]_ , \new_[48021]_ , \new_[48022]_ ,
    \new_[48025]_ , \new_[48028]_ , \new_[48029]_ , \new_[48030]_ ,
    \new_[48033]_ , \new_[48036]_ , \new_[48037]_ , \new_[48040]_ ,
    \new_[48043]_ , \new_[48044]_ , \new_[48045]_ , \new_[48048]_ ,
    \new_[48051]_ , \new_[48052]_ , \new_[48055]_ , \new_[48058]_ ,
    \new_[48059]_ , \new_[48060]_ , \new_[48063]_ , \new_[48066]_ ,
    \new_[48067]_ , \new_[48070]_ , \new_[48073]_ , \new_[48074]_ ,
    \new_[48075]_ , \new_[48078]_ , \new_[48081]_ , \new_[48082]_ ,
    \new_[48085]_ , \new_[48088]_ , \new_[48089]_ , \new_[48090]_ ,
    \new_[48093]_ , \new_[48096]_ , \new_[48097]_ , \new_[48100]_ ,
    \new_[48103]_ , \new_[48104]_ , \new_[48105]_ , \new_[48108]_ ,
    \new_[48111]_ , \new_[48112]_ , \new_[48115]_ , \new_[48118]_ ,
    \new_[48119]_ , \new_[48120]_ , \new_[48123]_ , \new_[48126]_ ,
    \new_[48127]_ , \new_[48130]_ , \new_[48133]_ , \new_[48134]_ ,
    \new_[48135]_ , \new_[48138]_ , \new_[48141]_ , \new_[48142]_ ,
    \new_[48145]_ , \new_[48148]_ , \new_[48149]_ , \new_[48150]_ ,
    \new_[48153]_ , \new_[48156]_ , \new_[48157]_ , \new_[48160]_ ,
    \new_[48163]_ , \new_[48164]_ , \new_[48165]_ , \new_[48168]_ ,
    \new_[48171]_ , \new_[48172]_ , \new_[48175]_ , \new_[48178]_ ,
    \new_[48179]_ , \new_[48180]_ , \new_[48183]_ , \new_[48186]_ ,
    \new_[48187]_ , \new_[48190]_ , \new_[48193]_ , \new_[48194]_ ,
    \new_[48195]_ , \new_[48198]_ , \new_[48201]_ , \new_[48202]_ ,
    \new_[48205]_ , \new_[48208]_ , \new_[48209]_ , \new_[48210]_ ,
    \new_[48213]_ , \new_[48216]_ , \new_[48217]_ , \new_[48220]_ ,
    \new_[48223]_ , \new_[48224]_ , \new_[48225]_ , \new_[48228]_ ,
    \new_[48231]_ , \new_[48232]_ , \new_[48235]_ , \new_[48238]_ ,
    \new_[48239]_ , \new_[48240]_ , \new_[48243]_ , \new_[48246]_ ,
    \new_[48247]_ , \new_[48250]_ , \new_[48253]_ , \new_[48254]_ ,
    \new_[48255]_ , \new_[48258]_ , \new_[48261]_ , \new_[48262]_ ,
    \new_[48265]_ , \new_[48268]_ , \new_[48269]_ , \new_[48270]_ ,
    \new_[48273]_ , \new_[48276]_ , \new_[48277]_ , \new_[48280]_ ,
    \new_[48283]_ , \new_[48284]_ , \new_[48285]_ , \new_[48288]_ ,
    \new_[48291]_ , \new_[48292]_ , \new_[48295]_ , \new_[48298]_ ,
    \new_[48299]_ , \new_[48300]_ , \new_[48303]_ , \new_[48306]_ ,
    \new_[48307]_ , \new_[48310]_ , \new_[48313]_ , \new_[48314]_ ,
    \new_[48315]_ , \new_[48318]_ , \new_[48321]_ , \new_[48322]_ ,
    \new_[48325]_ , \new_[48328]_ , \new_[48329]_ , \new_[48330]_ ,
    \new_[48333]_ , \new_[48336]_ , \new_[48337]_ , \new_[48340]_ ,
    \new_[48343]_ , \new_[48344]_ , \new_[48345]_ , \new_[48348]_ ,
    \new_[48351]_ , \new_[48352]_ , \new_[48355]_ , \new_[48358]_ ,
    \new_[48359]_ , \new_[48360]_ , \new_[48363]_ , \new_[48366]_ ,
    \new_[48367]_ , \new_[48370]_ , \new_[48373]_ , \new_[48374]_ ,
    \new_[48375]_ , \new_[48378]_ , \new_[48381]_ , \new_[48382]_ ,
    \new_[48385]_ , \new_[48388]_ , \new_[48389]_ , \new_[48390]_ ,
    \new_[48393]_ , \new_[48396]_ , \new_[48397]_ , \new_[48400]_ ,
    \new_[48403]_ , \new_[48404]_ , \new_[48405]_ , \new_[48408]_ ,
    \new_[48411]_ , \new_[48412]_ , \new_[48415]_ , \new_[48418]_ ,
    \new_[48419]_ , \new_[48420]_ , \new_[48423]_ , \new_[48426]_ ,
    \new_[48427]_ , \new_[48430]_ , \new_[48433]_ , \new_[48434]_ ,
    \new_[48435]_ , \new_[48438]_ , \new_[48441]_ , \new_[48442]_ ,
    \new_[48445]_ , \new_[48448]_ , \new_[48449]_ , \new_[48450]_ ,
    \new_[48453]_ , \new_[48456]_ , \new_[48457]_ , \new_[48460]_ ,
    \new_[48463]_ , \new_[48464]_ , \new_[48465]_ , \new_[48468]_ ,
    \new_[48471]_ , \new_[48472]_ , \new_[48475]_ , \new_[48478]_ ,
    \new_[48479]_ , \new_[48480]_ , \new_[48483]_ , \new_[48486]_ ,
    \new_[48487]_ , \new_[48490]_ , \new_[48493]_ , \new_[48494]_ ,
    \new_[48495]_ , \new_[48498]_ , \new_[48501]_ , \new_[48502]_ ,
    \new_[48505]_ , \new_[48508]_ , \new_[48509]_ , \new_[48510]_ ,
    \new_[48513]_ , \new_[48516]_ , \new_[48517]_ , \new_[48520]_ ,
    \new_[48523]_ , \new_[48524]_ , \new_[48525]_ , \new_[48528]_ ,
    \new_[48531]_ , \new_[48532]_ , \new_[48535]_ , \new_[48538]_ ,
    \new_[48539]_ , \new_[48540]_ , \new_[48543]_ , \new_[48546]_ ,
    \new_[48547]_ , \new_[48550]_ , \new_[48553]_ , \new_[48554]_ ,
    \new_[48555]_ , \new_[48558]_ , \new_[48561]_ , \new_[48562]_ ,
    \new_[48565]_ , \new_[48568]_ , \new_[48569]_ , \new_[48570]_ ,
    \new_[48573]_ , \new_[48576]_ , \new_[48577]_ , \new_[48580]_ ,
    \new_[48583]_ , \new_[48584]_ , \new_[48585]_ , \new_[48588]_ ,
    \new_[48591]_ , \new_[48592]_ , \new_[48595]_ , \new_[48598]_ ,
    \new_[48599]_ , \new_[48600]_ , \new_[48603]_ , \new_[48606]_ ,
    \new_[48607]_ , \new_[48610]_ , \new_[48613]_ , \new_[48614]_ ,
    \new_[48615]_ , \new_[48618]_ , \new_[48621]_ , \new_[48622]_ ,
    \new_[48625]_ , \new_[48628]_ , \new_[48629]_ , \new_[48630]_ ,
    \new_[48633]_ , \new_[48636]_ , \new_[48637]_ , \new_[48640]_ ,
    \new_[48643]_ , \new_[48644]_ , \new_[48645]_ , \new_[48648]_ ,
    \new_[48651]_ , \new_[48652]_ , \new_[48655]_ , \new_[48658]_ ,
    \new_[48659]_ , \new_[48660]_ , \new_[48663]_ , \new_[48666]_ ,
    \new_[48667]_ , \new_[48670]_ , \new_[48673]_ , \new_[48674]_ ,
    \new_[48675]_ , \new_[48678]_ , \new_[48681]_ , \new_[48682]_ ,
    \new_[48685]_ , \new_[48688]_ , \new_[48689]_ , \new_[48690]_ ,
    \new_[48693]_ , \new_[48696]_ , \new_[48697]_ , \new_[48700]_ ,
    \new_[48703]_ , \new_[48704]_ , \new_[48705]_ , \new_[48708]_ ,
    \new_[48711]_ , \new_[48712]_ , \new_[48715]_ , \new_[48718]_ ,
    \new_[48719]_ , \new_[48720]_ , \new_[48723]_ , \new_[48726]_ ,
    \new_[48727]_ , \new_[48730]_ , \new_[48733]_ , \new_[48734]_ ,
    \new_[48735]_ , \new_[48738]_ , \new_[48741]_ , \new_[48742]_ ,
    \new_[48745]_ , \new_[48748]_ , \new_[48749]_ , \new_[48750]_ ,
    \new_[48753]_ , \new_[48756]_ , \new_[48757]_ , \new_[48760]_ ,
    \new_[48763]_ , \new_[48764]_ , \new_[48765]_ , \new_[48768]_ ,
    \new_[48771]_ , \new_[48772]_ , \new_[48775]_ , \new_[48778]_ ,
    \new_[48779]_ , \new_[48780]_ , \new_[48783]_ , \new_[48786]_ ,
    \new_[48787]_ , \new_[48790]_ , \new_[48793]_ , \new_[48794]_ ,
    \new_[48795]_ , \new_[48798]_ , \new_[48801]_ , \new_[48802]_ ,
    \new_[48805]_ , \new_[48808]_ , \new_[48809]_ , \new_[48810]_ ,
    \new_[48813]_ , \new_[48816]_ , \new_[48817]_ , \new_[48820]_ ,
    \new_[48823]_ , \new_[48824]_ , \new_[48825]_ , \new_[48828]_ ,
    \new_[48831]_ , \new_[48832]_ , \new_[48835]_ , \new_[48838]_ ,
    \new_[48839]_ , \new_[48840]_ , \new_[48843]_ , \new_[48846]_ ,
    \new_[48847]_ , \new_[48850]_ , \new_[48853]_ , \new_[48854]_ ,
    \new_[48855]_ , \new_[48858]_ , \new_[48861]_ , \new_[48862]_ ,
    \new_[48865]_ , \new_[48868]_ , \new_[48869]_ , \new_[48870]_ ,
    \new_[48873]_ , \new_[48876]_ , \new_[48877]_ , \new_[48880]_ ,
    \new_[48883]_ , \new_[48884]_ , \new_[48885]_ , \new_[48888]_ ,
    \new_[48891]_ , \new_[48892]_ , \new_[48895]_ , \new_[48898]_ ,
    \new_[48899]_ , \new_[48900]_ , \new_[48903]_ , \new_[48906]_ ,
    \new_[48907]_ , \new_[48910]_ , \new_[48913]_ , \new_[48914]_ ,
    \new_[48915]_ , \new_[48918]_ , \new_[48921]_ , \new_[48922]_ ,
    \new_[48925]_ , \new_[48928]_ , \new_[48929]_ , \new_[48930]_ ,
    \new_[48933]_ , \new_[48936]_ , \new_[48937]_ , \new_[48940]_ ,
    \new_[48943]_ , \new_[48944]_ , \new_[48945]_ , \new_[48948]_ ,
    \new_[48951]_ , \new_[48952]_ , \new_[48955]_ , \new_[48958]_ ,
    \new_[48959]_ , \new_[48960]_ , \new_[48963]_ , \new_[48966]_ ,
    \new_[48967]_ , \new_[48970]_ , \new_[48973]_ , \new_[48974]_ ,
    \new_[48975]_ , \new_[48978]_ , \new_[48981]_ , \new_[48982]_ ,
    \new_[48985]_ , \new_[48988]_ , \new_[48989]_ , \new_[48990]_ ,
    \new_[48993]_ , \new_[48996]_ , \new_[48997]_ , \new_[49000]_ ,
    \new_[49003]_ , \new_[49004]_ , \new_[49005]_ , \new_[49008]_ ,
    \new_[49011]_ , \new_[49012]_ , \new_[49015]_ , \new_[49018]_ ,
    \new_[49019]_ , \new_[49020]_ , \new_[49023]_ , \new_[49026]_ ,
    \new_[49027]_ , \new_[49030]_ , \new_[49033]_ , \new_[49034]_ ,
    \new_[49035]_ , \new_[49038]_ , \new_[49041]_ , \new_[49042]_ ,
    \new_[49045]_ , \new_[49048]_ , \new_[49049]_ , \new_[49050]_ ,
    \new_[49053]_ , \new_[49056]_ , \new_[49057]_ , \new_[49060]_ ,
    \new_[49063]_ , \new_[49064]_ , \new_[49065]_ , \new_[49068]_ ,
    \new_[49071]_ , \new_[49072]_ , \new_[49075]_ , \new_[49078]_ ,
    \new_[49079]_ , \new_[49080]_ , \new_[49083]_ , \new_[49086]_ ,
    \new_[49087]_ , \new_[49090]_ , \new_[49093]_ , \new_[49094]_ ,
    \new_[49095]_ , \new_[49098]_ , \new_[49101]_ , \new_[49102]_ ,
    \new_[49105]_ , \new_[49108]_ , \new_[49109]_ , \new_[49110]_ ,
    \new_[49113]_ , \new_[49116]_ , \new_[49117]_ , \new_[49120]_ ,
    \new_[49123]_ , \new_[49124]_ , \new_[49125]_ , \new_[49128]_ ,
    \new_[49131]_ , \new_[49132]_ , \new_[49135]_ , \new_[49138]_ ,
    \new_[49139]_ , \new_[49140]_ , \new_[49143]_ , \new_[49146]_ ,
    \new_[49147]_ , \new_[49150]_ , \new_[49153]_ , \new_[49154]_ ,
    \new_[49155]_ , \new_[49158]_ , \new_[49161]_ , \new_[49162]_ ,
    \new_[49165]_ , \new_[49168]_ , \new_[49169]_ , \new_[49170]_ ,
    \new_[49173]_ , \new_[49176]_ , \new_[49177]_ , \new_[49180]_ ,
    \new_[49183]_ , \new_[49184]_ , \new_[49185]_ , \new_[49188]_ ,
    \new_[49191]_ , \new_[49192]_ , \new_[49195]_ , \new_[49198]_ ,
    \new_[49199]_ , \new_[49200]_ , \new_[49203]_ , \new_[49206]_ ,
    \new_[49207]_ , \new_[49210]_ , \new_[49213]_ , \new_[49214]_ ,
    \new_[49215]_ , \new_[49218]_ , \new_[49221]_ , \new_[49222]_ ,
    \new_[49225]_ , \new_[49228]_ , \new_[49229]_ , \new_[49230]_ ,
    \new_[49233]_ , \new_[49236]_ , \new_[49237]_ , \new_[49240]_ ,
    \new_[49243]_ , \new_[49244]_ , \new_[49245]_ , \new_[49248]_ ,
    \new_[49251]_ , \new_[49252]_ , \new_[49255]_ , \new_[49258]_ ,
    \new_[49259]_ , \new_[49260]_ , \new_[49263]_ , \new_[49266]_ ,
    \new_[49267]_ , \new_[49270]_ , \new_[49273]_ , \new_[49274]_ ,
    \new_[49275]_ , \new_[49278]_ , \new_[49281]_ , \new_[49282]_ ,
    \new_[49285]_ , \new_[49288]_ , \new_[49289]_ , \new_[49290]_ ,
    \new_[49293]_ , \new_[49296]_ , \new_[49297]_ , \new_[49300]_ ,
    \new_[49303]_ , \new_[49304]_ , \new_[49305]_ , \new_[49308]_ ,
    \new_[49311]_ , \new_[49312]_ , \new_[49315]_ , \new_[49318]_ ,
    \new_[49319]_ , \new_[49320]_ , \new_[49323]_ , \new_[49326]_ ,
    \new_[49327]_ , \new_[49330]_ , \new_[49333]_ , \new_[49334]_ ,
    \new_[49335]_ , \new_[49338]_ , \new_[49341]_ , \new_[49342]_ ,
    \new_[49345]_ , \new_[49348]_ , \new_[49349]_ , \new_[49350]_ ,
    \new_[49353]_ , \new_[49356]_ , \new_[49357]_ , \new_[49360]_ ,
    \new_[49363]_ , \new_[49364]_ , \new_[49365]_ , \new_[49368]_ ,
    \new_[49371]_ , \new_[49372]_ , \new_[49375]_ , \new_[49378]_ ,
    \new_[49379]_ , \new_[49380]_ , \new_[49383]_ , \new_[49386]_ ,
    \new_[49387]_ , \new_[49390]_ , \new_[49393]_ , \new_[49394]_ ,
    \new_[49395]_ , \new_[49398]_ , \new_[49401]_ , \new_[49402]_ ,
    \new_[49405]_ , \new_[49408]_ , \new_[49409]_ , \new_[49410]_ ,
    \new_[49413]_ , \new_[49416]_ , \new_[49417]_ , \new_[49420]_ ,
    \new_[49423]_ , \new_[49424]_ , \new_[49425]_ , \new_[49428]_ ,
    \new_[49431]_ , \new_[49432]_ , \new_[49435]_ , \new_[49438]_ ,
    \new_[49439]_ , \new_[49440]_ , \new_[49443]_ , \new_[49446]_ ,
    \new_[49447]_ , \new_[49450]_ , \new_[49453]_ , \new_[49454]_ ,
    \new_[49455]_ , \new_[49458]_ , \new_[49461]_ , \new_[49462]_ ,
    \new_[49465]_ , \new_[49468]_ , \new_[49469]_ , \new_[49470]_ ,
    \new_[49473]_ , \new_[49476]_ , \new_[49477]_ , \new_[49480]_ ,
    \new_[49483]_ , \new_[49484]_ , \new_[49485]_ , \new_[49488]_ ,
    \new_[49491]_ , \new_[49492]_ , \new_[49495]_ , \new_[49498]_ ,
    \new_[49499]_ , \new_[49500]_ , \new_[49503]_ , \new_[49506]_ ,
    \new_[49507]_ , \new_[49510]_ , \new_[49513]_ , \new_[49514]_ ,
    \new_[49515]_ , \new_[49518]_ , \new_[49521]_ , \new_[49522]_ ,
    \new_[49525]_ , \new_[49528]_ , \new_[49529]_ , \new_[49530]_ ,
    \new_[49533]_ , \new_[49536]_ , \new_[49537]_ , \new_[49540]_ ,
    \new_[49543]_ , \new_[49544]_ , \new_[49545]_ , \new_[49548]_ ,
    \new_[49551]_ , \new_[49552]_ , \new_[49555]_ , \new_[49558]_ ,
    \new_[49559]_ , \new_[49560]_ , \new_[49563]_ , \new_[49566]_ ,
    \new_[49567]_ , \new_[49570]_ , \new_[49573]_ , \new_[49574]_ ,
    \new_[49575]_ , \new_[49578]_ , \new_[49581]_ , \new_[49582]_ ,
    \new_[49585]_ , \new_[49588]_ , \new_[49589]_ , \new_[49590]_ ,
    \new_[49593]_ , \new_[49596]_ , \new_[49597]_ , \new_[49600]_ ,
    \new_[49603]_ , \new_[49604]_ , \new_[49605]_ , \new_[49608]_ ,
    \new_[49611]_ , \new_[49612]_ , \new_[49615]_ , \new_[49618]_ ,
    \new_[49619]_ , \new_[49620]_ , \new_[49623]_ , \new_[49626]_ ,
    \new_[49627]_ , \new_[49630]_ , \new_[49633]_ , \new_[49634]_ ,
    \new_[49635]_ , \new_[49638]_ , \new_[49641]_ , \new_[49642]_ ,
    \new_[49645]_ , \new_[49648]_ , \new_[49649]_ , \new_[49650]_ ,
    \new_[49653]_ , \new_[49656]_ , \new_[49657]_ , \new_[49660]_ ,
    \new_[49663]_ , \new_[49664]_ , \new_[49665]_ , \new_[49668]_ ,
    \new_[49671]_ , \new_[49672]_ , \new_[49675]_ , \new_[49678]_ ,
    \new_[49679]_ , \new_[49680]_ , \new_[49683]_ , \new_[49686]_ ,
    \new_[49687]_ , \new_[49690]_ , \new_[49693]_ , \new_[49694]_ ,
    \new_[49695]_ , \new_[49698]_ , \new_[49701]_ , \new_[49702]_ ,
    \new_[49705]_ , \new_[49708]_ , \new_[49709]_ , \new_[49710]_ ,
    \new_[49713]_ , \new_[49716]_ , \new_[49717]_ , \new_[49720]_ ,
    \new_[49723]_ , \new_[49724]_ , \new_[49725]_ , \new_[49728]_ ,
    \new_[49731]_ , \new_[49732]_ , \new_[49735]_ , \new_[49738]_ ,
    \new_[49739]_ , \new_[49740]_ , \new_[49743]_ , \new_[49746]_ ,
    \new_[49747]_ , \new_[49750]_ , \new_[49753]_ , \new_[49754]_ ,
    \new_[49755]_ , \new_[49758]_ , \new_[49761]_ , \new_[49762]_ ,
    \new_[49765]_ , \new_[49768]_ , \new_[49769]_ , \new_[49770]_ ,
    \new_[49773]_ , \new_[49776]_ , \new_[49777]_ , \new_[49780]_ ,
    \new_[49783]_ , \new_[49784]_ , \new_[49785]_ , \new_[49788]_ ,
    \new_[49791]_ , \new_[49792]_ , \new_[49795]_ , \new_[49798]_ ,
    \new_[49799]_ , \new_[49800]_ , \new_[49803]_ , \new_[49806]_ ,
    \new_[49807]_ , \new_[49810]_ , \new_[49813]_ , \new_[49814]_ ,
    \new_[49815]_ , \new_[49818]_ , \new_[49821]_ , \new_[49822]_ ,
    \new_[49825]_ , \new_[49828]_ , \new_[49829]_ , \new_[49830]_ ,
    \new_[49833]_ , \new_[49836]_ , \new_[49837]_ , \new_[49840]_ ,
    \new_[49843]_ , \new_[49844]_ , \new_[49845]_ , \new_[49848]_ ,
    \new_[49851]_ , \new_[49852]_ , \new_[49855]_ , \new_[49858]_ ,
    \new_[49859]_ , \new_[49860]_ , \new_[49863]_ , \new_[49866]_ ,
    \new_[49867]_ , \new_[49870]_ , \new_[49873]_ , \new_[49874]_ ,
    \new_[49875]_ , \new_[49878]_ , \new_[49881]_ , \new_[49882]_ ,
    \new_[49885]_ , \new_[49888]_ , \new_[49889]_ , \new_[49890]_ ,
    \new_[49893]_ , \new_[49896]_ , \new_[49897]_ , \new_[49900]_ ,
    \new_[49903]_ , \new_[49904]_ , \new_[49905]_ , \new_[49908]_ ,
    \new_[49911]_ , \new_[49912]_ , \new_[49915]_ , \new_[49918]_ ,
    \new_[49919]_ , \new_[49920]_ , \new_[49923]_ , \new_[49926]_ ,
    \new_[49927]_ , \new_[49930]_ , \new_[49933]_ , \new_[49934]_ ,
    \new_[49935]_ , \new_[49938]_ , \new_[49941]_ , \new_[49942]_ ,
    \new_[49945]_ , \new_[49948]_ , \new_[49949]_ , \new_[49950]_ ,
    \new_[49953]_ , \new_[49956]_ , \new_[49957]_ , \new_[49960]_ ,
    \new_[49963]_ , \new_[49964]_ , \new_[49965]_ , \new_[49968]_ ,
    \new_[49971]_ , \new_[49972]_ , \new_[49975]_ , \new_[49978]_ ,
    \new_[49979]_ , \new_[49980]_ , \new_[49983]_ , \new_[49986]_ ,
    \new_[49987]_ , \new_[49990]_ , \new_[49993]_ , \new_[49994]_ ,
    \new_[49995]_ , \new_[49998]_ , \new_[50001]_ , \new_[50002]_ ,
    \new_[50005]_ , \new_[50008]_ , \new_[50009]_ , \new_[50010]_ ,
    \new_[50013]_ , \new_[50016]_ , \new_[50017]_ , \new_[50020]_ ,
    \new_[50023]_ , \new_[50024]_ , \new_[50025]_ , \new_[50028]_ ,
    \new_[50031]_ , \new_[50032]_ , \new_[50035]_ , \new_[50038]_ ,
    \new_[50039]_ , \new_[50040]_ , \new_[50043]_ , \new_[50046]_ ,
    \new_[50047]_ , \new_[50050]_ , \new_[50053]_ , \new_[50054]_ ,
    \new_[50055]_ , \new_[50058]_ , \new_[50061]_ , \new_[50062]_ ,
    \new_[50065]_ , \new_[50068]_ , \new_[50069]_ , \new_[50070]_ ,
    \new_[50073]_ , \new_[50076]_ , \new_[50077]_ , \new_[50080]_ ,
    \new_[50083]_ , \new_[50084]_ , \new_[50085]_ , \new_[50088]_ ,
    \new_[50091]_ , \new_[50092]_ , \new_[50095]_ , \new_[50098]_ ,
    \new_[50099]_ , \new_[50100]_ , \new_[50103]_ , \new_[50106]_ ,
    \new_[50107]_ , \new_[50110]_ , \new_[50113]_ , \new_[50114]_ ,
    \new_[50115]_ , \new_[50118]_ , \new_[50121]_ , \new_[50122]_ ,
    \new_[50125]_ , \new_[50128]_ , \new_[50129]_ , \new_[50130]_ ,
    \new_[50133]_ , \new_[50136]_ , \new_[50137]_ , \new_[50140]_ ,
    \new_[50143]_ , \new_[50144]_ , \new_[50145]_ , \new_[50148]_ ,
    \new_[50151]_ , \new_[50152]_ , \new_[50155]_ , \new_[50158]_ ,
    \new_[50159]_ , \new_[50160]_ , \new_[50163]_ , \new_[50166]_ ,
    \new_[50167]_ , \new_[50170]_ , \new_[50173]_ , \new_[50174]_ ,
    \new_[50175]_ , \new_[50178]_ , \new_[50181]_ , \new_[50182]_ ,
    \new_[50185]_ , \new_[50188]_ , \new_[50189]_ , \new_[50190]_ ,
    \new_[50193]_ , \new_[50196]_ , \new_[50197]_ , \new_[50200]_ ,
    \new_[50203]_ , \new_[50204]_ , \new_[50205]_ , \new_[50208]_ ,
    \new_[50211]_ , \new_[50212]_ , \new_[50215]_ , \new_[50218]_ ,
    \new_[50219]_ , \new_[50220]_ , \new_[50223]_ , \new_[50226]_ ,
    \new_[50227]_ , \new_[50230]_ , \new_[50233]_ , \new_[50234]_ ,
    \new_[50235]_ , \new_[50238]_ , \new_[50241]_ , \new_[50242]_ ,
    \new_[50245]_ , \new_[50248]_ , \new_[50249]_ , \new_[50250]_ ,
    \new_[50253]_ , \new_[50256]_ , \new_[50257]_ , \new_[50260]_ ,
    \new_[50263]_ , \new_[50264]_ , \new_[50265]_ , \new_[50268]_ ,
    \new_[50271]_ , \new_[50272]_ , \new_[50275]_ , \new_[50278]_ ,
    \new_[50279]_ , \new_[50280]_ , \new_[50283]_ , \new_[50286]_ ,
    \new_[50287]_ , \new_[50290]_ , \new_[50293]_ , \new_[50294]_ ,
    \new_[50295]_ , \new_[50298]_ , \new_[50301]_ , \new_[50302]_ ,
    \new_[50305]_ , \new_[50308]_ , \new_[50309]_ , \new_[50310]_ ,
    \new_[50313]_ , \new_[50316]_ , \new_[50317]_ , \new_[50320]_ ,
    \new_[50323]_ , \new_[50324]_ , \new_[50325]_ , \new_[50328]_ ,
    \new_[50331]_ , \new_[50332]_ , \new_[50335]_ , \new_[50338]_ ,
    \new_[50339]_ , \new_[50340]_ , \new_[50343]_ , \new_[50346]_ ,
    \new_[50347]_ , \new_[50350]_ , \new_[50353]_ , \new_[50354]_ ,
    \new_[50355]_ , \new_[50358]_ , \new_[50361]_ , \new_[50362]_ ,
    \new_[50365]_ , \new_[50368]_ , \new_[50369]_ , \new_[50370]_ ,
    \new_[50373]_ , \new_[50376]_ , \new_[50377]_ , \new_[50380]_ ,
    \new_[50383]_ , \new_[50384]_ , \new_[50385]_ , \new_[50388]_ ,
    \new_[50391]_ , \new_[50392]_ , \new_[50395]_ , \new_[50398]_ ,
    \new_[50399]_ , \new_[50400]_ , \new_[50403]_ , \new_[50406]_ ,
    \new_[50407]_ , \new_[50410]_ , \new_[50413]_ , \new_[50414]_ ,
    \new_[50415]_ , \new_[50418]_ , \new_[50421]_ , \new_[50422]_ ,
    \new_[50425]_ , \new_[50428]_ , \new_[50429]_ , \new_[50430]_ ,
    \new_[50433]_ , \new_[50436]_ , \new_[50437]_ , \new_[50440]_ ,
    \new_[50443]_ , \new_[50444]_ , \new_[50445]_ , \new_[50448]_ ,
    \new_[50451]_ , \new_[50452]_ , \new_[50455]_ , \new_[50458]_ ,
    \new_[50459]_ , \new_[50460]_ , \new_[50463]_ , \new_[50466]_ ,
    \new_[50467]_ , \new_[50470]_ , \new_[50473]_ , \new_[50474]_ ,
    \new_[50475]_ , \new_[50478]_ , \new_[50481]_ , \new_[50482]_ ,
    \new_[50485]_ , \new_[50488]_ , \new_[50489]_ , \new_[50490]_ ,
    \new_[50493]_ , \new_[50496]_ , \new_[50497]_ , \new_[50500]_ ,
    \new_[50503]_ , \new_[50504]_ , \new_[50505]_ , \new_[50508]_ ,
    \new_[50511]_ , \new_[50512]_ , \new_[50515]_ , \new_[50518]_ ,
    \new_[50519]_ , \new_[50520]_ , \new_[50523]_ , \new_[50526]_ ,
    \new_[50527]_ , \new_[50530]_ , \new_[50533]_ , \new_[50534]_ ,
    \new_[50535]_ , \new_[50538]_ , \new_[50541]_ , \new_[50542]_ ,
    \new_[50545]_ , \new_[50548]_ , \new_[50549]_ , \new_[50550]_ ,
    \new_[50553]_ , \new_[50556]_ , \new_[50557]_ , \new_[50560]_ ,
    \new_[50563]_ , \new_[50564]_ , \new_[50565]_ , \new_[50568]_ ,
    \new_[50571]_ , \new_[50572]_ , \new_[50575]_ , \new_[50578]_ ,
    \new_[50579]_ , \new_[50580]_ , \new_[50583]_ , \new_[50586]_ ,
    \new_[50587]_ , \new_[50590]_ , \new_[50593]_ , \new_[50594]_ ,
    \new_[50595]_ , \new_[50598]_ , \new_[50601]_ , \new_[50602]_ ,
    \new_[50605]_ , \new_[50608]_ , \new_[50609]_ , \new_[50610]_ ,
    \new_[50613]_ , \new_[50616]_ , \new_[50617]_ , \new_[50620]_ ,
    \new_[50623]_ , \new_[50624]_ , \new_[50625]_ , \new_[50628]_ ,
    \new_[50631]_ , \new_[50632]_ , \new_[50635]_ , \new_[50638]_ ,
    \new_[50639]_ , \new_[50640]_ , \new_[50643]_ , \new_[50646]_ ,
    \new_[50647]_ , \new_[50650]_ , \new_[50653]_ , \new_[50654]_ ,
    \new_[50655]_ , \new_[50658]_ , \new_[50661]_ , \new_[50662]_ ,
    \new_[50665]_ , \new_[50668]_ , \new_[50669]_ , \new_[50670]_ ,
    \new_[50673]_ , \new_[50676]_ , \new_[50677]_ , \new_[50680]_ ,
    \new_[50683]_ , \new_[50684]_ , \new_[50685]_ , \new_[50688]_ ,
    \new_[50691]_ , \new_[50692]_ , \new_[50695]_ , \new_[50698]_ ,
    \new_[50699]_ , \new_[50700]_ , \new_[50703]_ , \new_[50706]_ ,
    \new_[50707]_ , \new_[50710]_ , \new_[50713]_ , \new_[50714]_ ,
    \new_[50715]_ , \new_[50718]_ , \new_[50721]_ , \new_[50722]_ ,
    \new_[50725]_ , \new_[50728]_ , \new_[50729]_ , \new_[50730]_ ,
    \new_[50733]_ , \new_[50736]_ , \new_[50737]_ , \new_[50740]_ ,
    \new_[50743]_ , \new_[50744]_ , \new_[50745]_ , \new_[50748]_ ,
    \new_[50751]_ , \new_[50752]_ , \new_[50755]_ , \new_[50758]_ ,
    \new_[50759]_ , \new_[50760]_ , \new_[50763]_ , \new_[50766]_ ,
    \new_[50767]_ , \new_[50770]_ , \new_[50773]_ , \new_[50774]_ ,
    \new_[50775]_ , \new_[50778]_ , \new_[50781]_ , \new_[50782]_ ,
    \new_[50785]_ , \new_[50788]_ , \new_[50789]_ , \new_[50790]_ ,
    \new_[50793]_ , \new_[50796]_ , \new_[50797]_ , \new_[50800]_ ,
    \new_[50803]_ , \new_[50804]_ , \new_[50805]_ , \new_[50808]_ ,
    \new_[50811]_ , \new_[50812]_ , \new_[50815]_ , \new_[50818]_ ,
    \new_[50819]_ , \new_[50820]_ , \new_[50823]_ , \new_[50826]_ ,
    \new_[50827]_ , \new_[50830]_ , \new_[50833]_ , \new_[50834]_ ,
    \new_[50835]_ , \new_[50838]_ , \new_[50841]_ , \new_[50842]_ ,
    \new_[50845]_ , \new_[50848]_ , \new_[50849]_ , \new_[50850]_ ,
    \new_[50853]_ , \new_[50856]_ , \new_[50857]_ , \new_[50860]_ ,
    \new_[50863]_ , \new_[50864]_ , \new_[50865]_ , \new_[50868]_ ,
    \new_[50871]_ , \new_[50872]_ , \new_[50875]_ , \new_[50878]_ ,
    \new_[50879]_ , \new_[50880]_ , \new_[50883]_ , \new_[50886]_ ,
    \new_[50887]_ , \new_[50890]_ , \new_[50893]_ , \new_[50894]_ ,
    \new_[50895]_ , \new_[50898]_ , \new_[50901]_ , \new_[50902]_ ,
    \new_[50905]_ , \new_[50908]_ , \new_[50909]_ , \new_[50910]_ ,
    \new_[50913]_ , \new_[50916]_ , \new_[50917]_ , \new_[50920]_ ,
    \new_[50923]_ , \new_[50924]_ , \new_[50925]_ , \new_[50928]_ ,
    \new_[50931]_ , \new_[50932]_ , \new_[50935]_ , \new_[50938]_ ,
    \new_[50939]_ , \new_[50940]_ , \new_[50943]_ , \new_[50946]_ ,
    \new_[50947]_ , \new_[50950]_ , \new_[50953]_ , \new_[50954]_ ,
    \new_[50955]_ , \new_[50958]_ , \new_[50961]_ , \new_[50962]_ ,
    \new_[50965]_ , \new_[50968]_ , \new_[50969]_ , \new_[50970]_ ,
    \new_[50973]_ , \new_[50976]_ , \new_[50977]_ , \new_[50980]_ ,
    \new_[50983]_ , \new_[50984]_ , \new_[50985]_ , \new_[50988]_ ,
    \new_[50991]_ , \new_[50992]_ , \new_[50995]_ , \new_[50998]_ ,
    \new_[50999]_ , \new_[51000]_ , \new_[51003]_ , \new_[51006]_ ,
    \new_[51007]_ , \new_[51010]_ , \new_[51013]_ , \new_[51014]_ ,
    \new_[51015]_ , \new_[51018]_ , \new_[51021]_ , \new_[51022]_ ,
    \new_[51025]_ , \new_[51028]_ , \new_[51029]_ , \new_[51030]_ ,
    \new_[51033]_ , \new_[51036]_ , \new_[51037]_ , \new_[51040]_ ,
    \new_[51043]_ , \new_[51044]_ , \new_[51045]_ , \new_[51048]_ ,
    \new_[51051]_ , \new_[51052]_ , \new_[51055]_ , \new_[51058]_ ,
    \new_[51059]_ , \new_[51060]_ , \new_[51063]_ , \new_[51066]_ ,
    \new_[51067]_ , \new_[51070]_ , \new_[51073]_ , \new_[51074]_ ,
    \new_[51075]_ , \new_[51078]_ , \new_[51081]_ , \new_[51082]_ ,
    \new_[51085]_ , \new_[51088]_ , \new_[51089]_ , \new_[51090]_ ,
    \new_[51093]_ , \new_[51096]_ , \new_[51097]_ , \new_[51100]_ ,
    \new_[51103]_ , \new_[51104]_ , \new_[51105]_ , \new_[51108]_ ,
    \new_[51111]_ , \new_[51112]_ , \new_[51115]_ , \new_[51118]_ ,
    \new_[51119]_ , \new_[51120]_ , \new_[51123]_ , \new_[51126]_ ,
    \new_[51127]_ , \new_[51130]_ , \new_[51133]_ , \new_[51134]_ ,
    \new_[51135]_ , \new_[51138]_ , \new_[51141]_ , \new_[51142]_ ,
    \new_[51145]_ , \new_[51148]_ , \new_[51149]_ , \new_[51150]_ ,
    \new_[51153]_ , \new_[51156]_ , \new_[51157]_ , \new_[51160]_ ,
    \new_[51163]_ , \new_[51164]_ , \new_[51165]_ , \new_[51168]_ ,
    \new_[51171]_ , \new_[51172]_ , \new_[51175]_ , \new_[51178]_ ,
    \new_[51179]_ , \new_[51180]_ , \new_[51183]_ , \new_[51186]_ ,
    \new_[51187]_ , \new_[51190]_ , \new_[51193]_ , \new_[51194]_ ,
    \new_[51195]_ , \new_[51198]_ , \new_[51201]_ , \new_[51202]_ ,
    \new_[51205]_ , \new_[51208]_ , \new_[51209]_ , \new_[51210]_ ,
    \new_[51213]_ , \new_[51216]_ , \new_[51217]_ , \new_[51220]_ ,
    \new_[51223]_ , \new_[51224]_ , \new_[51225]_ , \new_[51228]_ ,
    \new_[51231]_ , \new_[51232]_ , \new_[51235]_ , \new_[51238]_ ,
    \new_[51239]_ , \new_[51240]_ , \new_[51243]_ , \new_[51246]_ ,
    \new_[51247]_ , \new_[51250]_ , \new_[51253]_ , \new_[51254]_ ,
    \new_[51255]_ , \new_[51258]_ , \new_[51261]_ , \new_[51262]_ ,
    \new_[51265]_ , \new_[51268]_ , \new_[51269]_ , \new_[51270]_ ,
    \new_[51273]_ , \new_[51276]_ , \new_[51277]_ , \new_[51280]_ ,
    \new_[51283]_ , \new_[51284]_ , \new_[51285]_ , \new_[51288]_ ,
    \new_[51291]_ , \new_[51292]_ , \new_[51295]_ , \new_[51298]_ ,
    \new_[51299]_ , \new_[51300]_ , \new_[51303]_ , \new_[51306]_ ,
    \new_[51307]_ , \new_[51310]_ , \new_[51313]_ , \new_[51314]_ ,
    \new_[51315]_ , \new_[51318]_ , \new_[51321]_ , \new_[51322]_ ,
    \new_[51325]_ , \new_[51328]_ , \new_[51329]_ , \new_[51330]_ ,
    \new_[51333]_ , \new_[51336]_ , \new_[51337]_ , \new_[51340]_ ,
    \new_[51343]_ , \new_[51344]_ , \new_[51345]_ , \new_[51348]_ ,
    \new_[51351]_ , \new_[51352]_ , \new_[51355]_ , \new_[51358]_ ,
    \new_[51359]_ , \new_[51360]_ , \new_[51363]_ , \new_[51366]_ ,
    \new_[51367]_ , \new_[51370]_ , \new_[51373]_ , \new_[51374]_ ,
    \new_[51375]_ , \new_[51378]_ , \new_[51381]_ , \new_[51382]_ ,
    \new_[51385]_ , \new_[51388]_ , \new_[51389]_ , \new_[51390]_ ,
    \new_[51393]_ , \new_[51396]_ , \new_[51397]_ , \new_[51400]_ ,
    \new_[51403]_ , \new_[51404]_ , \new_[51405]_ , \new_[51408]_ ,
    \new_[51411]_ , \new_[51412]_ , \new_[51415]_ , \new_[51418]_ ,
    \new_[51419]_ , \new_[51420]_ , \new_[51423]_ , \new_[51426]_ ,
    \new_[51427]_ , \new_[51430]_ , \new_[51433]_ , \new_[51434]_ ,
    \new_[51435]_ , \new_[51438]_ , \new_[51441]_ , \new_[51442]_ ,
    \new_[51445]_ , \new_[51448]_ , \new_[51449]_ , \new_[51450]_ ,
    \new_[51453]_ , \new_[51456]_ , \new_[51457]_ , \new_[51460]_ ,
    \new_[51463]_ , \new_[51464]_ , \new_[51465]_ , \new_[51468]_ ,
    \new_[51471]_ , \new_[51472]_ , \new_[51475]_ , \new_[51478]_ ,
    \new_[51479]_ , \new_[51480]_ , \new_[51483]_ , \new_[51486]_ ,
    \new_[51487]_ , \new_[51490]_ , \new_[51493]_ , \new_[51494]_ ,
    \new_[51495]_ , \new_[51498]_ , \new_[51501]_ , \new_[51502]_ ,
    \new_[51505]_ , \new_[51508]_ , \new_[51509]_ , \new_[51510]_ ,
    \new_[51513]_ , \new_[51516]_ , \new_[51517]_ , \new_[51520]_ ,
    \new_[51523]_ , \new_[51524]_ , \new_[51525]_ , \new_[51528]_ ,
    \new_[51531]_ , \new_[51532]_ , \new_[51535]_ , \new_[51538]_ ,
    \new_[51539]_ , \new_[51540]_ , \new_[51543]_ , \new_[51546]_ ,
    \new_[51547]_ , \new_[51550]_ , \new_[51553]_ , \new_[51554]_ ,
    \new_[51555]_ , \new_[51558]_ , \new_[51561]_ , \new_[51562]_ ,
    \new_[51565]_ , \new_[51568]_ , \new_[51569]_ , \new_[51570]_ ,
    \new_[51573]_ , \new_[51576]_ , \new_[51577]_ , \new_[51580]_ ,
    \new_[51583]_ , \new_[51584]_ , \new_[51585]_ , \new_[51588]_ ,
    \new_[51591]_ , \new_[51592]_ , \new_[51595]_ , \new_[51598]_ ,
    \new_[51599]_ , \new_[51600]_ , \new_[51603]_ , \new_[51606]_ ,
    \new_[51607]_ , \new_[51610]_ , \new_[51613]_ , \new_[51614]_ ,
    \new_[51615]_ , \new_[51618]_ , \new_[51621]_ , \new_[51622]_ ,
    \new_[51625]_ , \new_[51628]_ , \new_[51629]_ , \new_[51630]_ ,
    \new_[51633]_ , \new_[51636]_ , \new_[51637]_ , \new_[51640]_ ,
    \new_[51643]_ , \new_[51644]_ , \new_[51645]_ , \new_[51648]_ ,
    \new_[51651]_ , \new_[51652]_ , \new_[51655]_ , \new_[51658]_ ,
    \new_[51659]_ , \new_[51660]_ , \new_[51663]_ , \new_[51666]_ ,
    \new_[51667]_ , \new_[51670]_ , \new_[51673]_ , \new_[51674]_ ,
    \new_[51675]_ , \new_[51678]_ , \new_[51681]_ , \new_[51682]_ ,
    \new_[51685]_ , \new_[51688]_ , \new_[51689]_ , \new_[51690]_ ,
    \new_[51693]_ , \new_[51696]_ , \new_[51697]_ , \new_[51700]_ ,
    \new_[51703]_ , \new_[51704]_ , \new_[51705]_ , \new_[51708]_ ,
    \new_[51711]_ , \new_[51712]_ , \new_[51715]_ , \new_[51718]_ ,
    \new_[51719]_ , \new_[51720]_ , \new_[51723]_ , \new_[51726]_ ,
    \new_[51727]_ , \new_[51730]_ , \new_[51733]_ , \new_[51734]_ ,
    \new_[51735]_ , \new_[51738]_ , \new_[51741]_ , \new_[51742]_ ,
    \new_[51745]_ , \new_[51748]_ , \new_[51749]_ , \new_[51750]_ ,
    \new_[51753]_ , \new_[51756]_ , \new_[51757]_ , \new_[51760]_ ,
    \new_[51763]_ , \new_[51764]_ , \new_[51765]_ , \new_[51768]_ ,
    \new_[51771]_ , \new_[51772]_ , \new_[51775]_ , \new_[51778]_ ,
    \new_[51779]_ , \new_[51780]_ , \new_[51783]_ , \new_[51786]_ ,
    \new_[51787]_ , \new_[51790]_ , \new_[51793]_ , \new_[51794]_ ,
    \new_[51795]_ , \new_[51798]_ , \new_[51801]_ , \new_[51802]_ ,
    \new_[51805]_ , \new_[51808]_ , \new_[51809]_ , \new_[51810]_ ,
    \new_[51813]_ , \new_[51816]_ , \new_[51817]_ , \new_[51820]_ ,
    \new_[51823]_ , \new_[51824]_ , \new_[51825]_ , \new_[51828]_ ,
    \new_[51831]_ , \new_[51832]_ , \new_[51835]_ , \new_[51838]_ ,
    \new_[51839]_ , \new_[51840]_ , \new_[51843]_ , \new_[51846]_ ,
    \new_[51847]_ , \new_[51850]_ , \new_[51853]_ , \new_[51854]_ ,
    \new_[51855]_ , \new_[51858]_ , \new_[51861]_ , \new_[51862]_ ,
    \new_[51865]_ , \new_[51868]_ , \new_[51869]_ , \new_[51870]_ ,
    \new_[51873]_ , \new_[51876]_ , \new_[51877]_ , \new_[51880]_ ,
    \new_[51883]_ , \new_[51884]_ , \new_[51885]_ , \new_[51888]_ ,
    \new_[51891]_ , \new_[51892]_ , \new_[51895]_ , \new_[51898]_ ,
    \new_[51899]_ , \new_[51900]_ , \new_[51903]_ , \new_[51906]_ ,
    \new_[51907]_ , \new_[51910]_ , \new_[51913]_ , \new_[51914]_ ,
    \new_[51915]_ , \new_[51918]_ , \new_[51921]_ , \new_[51922]_ ,
    \new_[51925]_ , \new_[51928]_ , \new_[51929]_ , \new_[51930]_ ,
    \new_[51933]_ , \new_[51936]_ , \new_[51937]_ , \new_[51940]_ ,
    \new_[51943]_ , \new_[51944]_ , \new_[51945]_ , \new_[51948]_ ,
    \new_[51951]_ , \new_[51952]_ , \new_[51955]_ , \new_[51958]_ ,
    \new_[51959]_ , \new_[51960]_ , \new_[51963]_ , \new_[51966]_ ,
    \new_[51967]_ , \new_[51970]_ , \new_[51973]_ , \new_[51974]_ ,
    \new_[51975]_ , \new_[51978]_ , \new_[51981]_ , \new_[51982]_ ,
    \new_[51985]_ , \new_[51988]_ , \new_[51989]_ , \new_[51990]_ ,
    \new_[51993]_ , \new_[51996]_ , \new_[51997]_ , \new_[52000]_ ,
    \new_[52003]_ , \new_[52004]_ , \new_[52005]_ , \new_[52008]_ ,
    \new_[52011]_ , \new_[52012]_ , \new_[52015]_ , \new_[52018]_ ,
    \new_[52019]_ , \new_[52020]_ , \new_[52023]_ , \new_[52026]_ ,
    \new_[52027]_ , \new_[52030]_ , \new_[52033]_ , \new_[52034]_ ,
    \new_[52035]_ , \new_[52038]_ , \new_[52041]_ , \new_[52042]_ ,
    \new_[52045]_ , \new_[52048]_ , \new_[52049]_ , \new_[52050]_ ,
    \new_[52053]_ , \new_[52056]_ , \new_[52057]_ , \new_[52060]_ ,
    \new_[52063]_ , \new_[52064]_ , \new_[52065]_ , \new_[52068]_ ,
    \new_[52071]_ , \new_[52072]_ , \new_[52075]_ , \new_[52078]_ ,
    \new_[52079]_ , \new_[52080]_ , \new_[52083]_ , \new_[52086]_ ,
    \new_[52087]_ , \new_[52090]_ , \new_[52093]_ , \new_[52094]_ ,
    \new_[52095]_ , \new_[52098]_ , \new_[52101]_ , \new_[52102]_ ,
    \new_[52105]_ , \new_[52108]_ , \new_[52109]_ , \new_[52110]_ ,
    \new_[52113]_ , \new_[52116]_ , \new_[52117]_ , \new_[52120]_ ,
    \new_[52123]_ , \new_[52124]_ , \new_[52125]_ , \new_[52128]_ ,
    \new_[52131]_ , \new_[52132]_ , \new_[52135]_ , \new_[52138]_ ,
    \new_[52139]_ , \new_[52140]_ , \new_[52143]_ , \new_[52146]_ ,
    \new_[52147]_ , \new_[52150]_ , \new_[52153]_ , \new_[52154]_ ,
    \new_[52155]_ , \new_[52158]_ , \new_[52161]_ , \new_[52162]_ ,
    \new_[52165]_ , \new_[52168]_ , \new_[52169]_ , \new_[52170]_ ,
    \new_[52173]_ , \new_[52176]_ , \new_[52177]_ , \new_[52180]_ ,
    \new_[52183]_ , \new_[52184]_ , \new_[52185]_ , \new_[52188]_ ,
    \new_[52191]_ , \new_[52192]_ , \new_[52195]_ , \new_[52198]_ ,
    \new_[52199]_ , \new_[52200]_ , \new_[52203]_ , \new_[52206]_ ,
    \new_[52207]_ , \new_[52210]_ , \new_[52213]_ , \new_[52214]_ ,
    \new_[52215]_ , \new_[52218]_ , \new_[52221]_ , \new_[52222]_ ,
    \new_[52225]_ , \new_[52228]_ , \new_[52229]_ , \new_[52230]_ ,
    \new_[52233]_ , \new_[52236]_ , \new_[52237]_ , \new_[52240]_ ,
    \new_[52243]_ , \new_[52244]_ , \new_[52245]_ , \new_[52248]_ ,
    \new_[52251]_ , \new_[52252]_ , \new_[52255]_ , \new_[52258]_ ,
    \new_[52259]_ , \new_[52260]_ , \new_[52263]_ , \new_[52266]_ ,
    \new_[52267]_ , \new_[52270]_ , \new_[52273]_ , \new_[52274]_ ,
    \new_[52275]_ , \new_[52278]_ , \new_[52281]_ , \new_[52282]_ ,
    \new_[52285]_ , \new_[52288]_ , \new_[52289]_ , \new_[52290]_ ,
    \new_[52293]_ , \new_[52296]_ , \new_[52297]_ , \new_[52300]_ ,
    \new_[52303]_ , \new_[52304]_ , \new_[52305]_ , \new_[52308]_ ,
    \new_[52311]_ , \new_[52312]_ , \new_[52315]_ , \new_[52318]_ ,
    \new_[52319]_ , \new_[52320]_ , \new_[52323]_ , \new_[52326]_ ,
    \new_[52327]_ , \new_[52330]_ , \new_[52333]_ , \new_[52334]_ ,
    \new_[52335]_ , \new_[52338]_ , \new_[52341]_ , \new_[52342]_ ,
    \new_[52345]_ , \new_[52348]_ , \new_[52349]_ , \new_[52350]_ ,
    \new_[52353]_ , \new_[52356]_ , \new_[52357]_ , \new_[52360]_ ,
    \new_[52363]_ , \new_[52364]_ , \new_[52365]_ , \new_[52368]_ ,
    \new_[52371]_ , \new_[52372]_ , \new_[52375]_ , \new_[52378]_ ,
    \new_[52379]_ , \new_[52380]_ , \new_[52383]_ , \new_[52386]_ ,
    \new_[52387]_ , \new_[52390]_ , \new_[52393]_ , \new_[52394]_ ,
    \new_[52395]_ , \new_[52398]_ , \new_[52401]_ , \new_[52402]_ ,
    \new_[52405]_ , \new_[52408]_ , \new_[52409]_ , \new_[52410]_ ,
    \new_[52413]_ , \new_[52416]_ , \new_[52417]_ , \new_[52420]_ ,
    \new_[52423]_ , \new_[52424]_ , \new_[52425]_ , \new_[52428]_ ,
    \new_[52431]_ , \new_[52432]_ , \new_[52435]_ , \new_[52438]_ ,
    \new_[52439]_ , \new_[52440]_ , \new_[52443]_ , \new_[52446]_ ,
    \new_[52447]_ , \new_[52450]_ , \new_[52453]_ , \new_[52454]_ ,
    \new_[52455]_ , \new_[52458]_ , \new_[52461]_ , \new_[52462]_ ,
    \new_[52465]_ , \new_[52468]_ , \new_[52469]_ , \new_[52470]_ ,
    \new_[52473]_ , \new_[52476]_ , \new_[52477]_ , \new_[52480]_ ,
    \new_[52483]_ , \new_[52484]_ , \new_[52485]_ , \new_[52488]_ ,
    \new_[52491]_ , \new_[52492]_ , \new_[52495]_ , \new_[52498]_ ,
    \new_[52499]_ , \new_[52500]_ , \new_[52503]_ , \new_[52506]_ ,
    \new_[52507]_ , \new_[52510]_ , \new_[52513]_ , \new_[52514]_ ,
    \new_[52515]_ , \new_[52518]_ , \new_[52521]_ , \new_[52522]_ ,
    \new_[52525]_ , \new_[52528]_ , \new_[52529]_ , \new_[52530]_ ,
    \new_[52533]_ , \new_[52536]_ , \new_[52537]_ , \new_[52540]_ ,
    \new_[52543]_ , \new_[52544]_ , \new_[52545]_ , \new_[52548]_ ,
    \new_[52551]_ , \new_[52552]_ , \new_[52555]_ , \new_[52558]_ ,
    \new_[52559]_ , \new_[52560]_ , \new_[52563]_ , \new_[52566]_ ,
    \new_[52567]_ , \new_[52570]_ , \new_[52573]_ , \new_[52574]_ ,
    \new_[52575]_ , \new_[52578]_ , \new_[52581]_ , \new_[52582]_ ,
    \new_[52585]_ , \new_[52588]_ , \new_[52589]_ , \new_[52590]_ ,
    \new_[52593]_ , \new_[52596]_ , \new_[52597]_ , \new_[52600]_ ,
    \new_[52603]_ , \new_[52604]_ , \new_[52605]_ , \new_[52608]_ ,
    \new_[52611]_ , \new_[52612]_ , \new_[52615]_ , \new_[52618]_ ,
    \new_[52619]_ , \new_[52620]_ , \new_[52623]_ , \new_[52626]_ ,
    \new_[52627]_ , \new_[52630]_ , \new_[52633]_ , \new_[52634]_ ,
    \new_[52635]_ , \new_[52638]_ , \new_[52641]_ , \new_[52642]_ ,
    \new_[52645]_ , \new_[52648]_ , \new_[52649]_ , \new_[52650]_ ,
    \new_[52653]_ , \new_[52656]_ , \new_[52657]_ , \new_[52660]_ ,
    \new_[52663]_ , \new_[52664]_ , \new_[52665]_ , \new_[52668]_ ,
    \new_[52671]_ , \new_[52672]_ , \new_[52675]_ , \new_[52678]_ ,
    \new_[52679]_ , \new_[52680]_ , \new_[52683]_ , \new_[52686]_ ,
    \new_[52687]_ , \new_[52690]_ , \new_[52693]_ , \new_[52694]_ ,
    \new_[52695]_ , \new_[52698]_ , \new_[52701]_ , \new_[52702]_ ,
    \new_[52705]_ , \new_[52708]_ , \new_[52709]_ , \new_[52710]_ ,
    \new_[52713]_ , \new_[52716]_ , \new_[52717]_ , \new_[52720]_ ,
    \new_[52723]_ , \new_[52724]_ , \new_[52725]_ , \new_[52728]_ ,
    \new_[52731]_ , \new_[52732]_ , \new_[52735]_ , \new_[52738]_ ,
    \new_[52739]_ , \new_[52740]_ , \new_[52743]_ , \new_[52746]_ ,
    \new_[52747]_ , \new_[52750]_ , \new_[52753]_ , \new_[52754]_ ,
    \new_[52755]_ , \new_[52758]_ , \new_[52761]_ , \new_[52762]_ ,
    \new_[52765]_ , \new_[52768]_ , \new_[52769]_ , \new_[52770]_ ,
    \new_[52773]_ , \new_[52776]_ , \new_[52777]_ , \new_[52780]_ ,
    \new_[52783]_ , \new_[52784]_ , \new_[52785]_ , \new_[52788]_ ,
    \new_[52791]_ , \new_[52792]_ , \new_[52795]_ , \new_[52798]_ ,
    \new_[52799]_ , \new_[52800]_ , \new_[52803]_ , \new_[52806]_ ,
    \new_[52807]_ , \new_[52810]_ , \new_[52813]_ , \new_[52814]_ ,
    \new_[52815]_ , \new_[52818]_ , \new_[52821]_ , \new_[52822]_ ,
    \new_[52825]_ , \new_[52828]_ , \new_[52829]_ , \new_[52830]_ ,
    \new_[52833]_ , \new_[52836]_ , \new_[52837]_ , \new_[52840]_ ,
    \new_[52843]_ , \new_[52844]_ , \new_[52845]_ , \new_[52848]_ ,
    \new_[52851]_ , \new_[52852]_ , \new_[52855]_ , \new_[52858]_ ,
    \new_[52859]_ , \new_[52860]_ , \new_[52863]_ , \new_[52866]_ ,
    \new_[52867]_ , \new_[52870]_ , \new_[52873]_ , \new_[52874]_ ,
    \new_[52875]_ , \new_[52878]_ , \new_[52881]_ , \new_[52882]_ ,
    \new_[52885]_ , \new_[52888]_ , \new_[52889]_ , \new_[52890]_ ,
    \new_[52893]_ , \new_[52896]_ , \new_[52897]_ , \new_[52900]_ ,
    \new_[52903]_ , \new_[52904]_ , \new_[52905]_ , \new_[52908]_ ,
    \new_[52911]_ , \new_[52912]_ , \new_[52915]_ , \new_[52918]_ ,
    \new_[52919]_ , \new_[52920]_ , \new_[52923]_ , \new_[52926]_ ,
    \new_[52927]_ , \new_[52930]_ , \new_[52933]_ , \new_[52934]_ ,
    \new_[52935]_ , \new_[52938]_ , \new_[52941]_ , \new_[52942]_ ,
    \new_[52945]_ , \new_[52948]_ , \new_[52949]_ , \new_[52950]_ ,
    \new_[52953]_ , \new_[52956]_ , \new_[52957]_ , \new_[52960]_ ,
    \new_[52963]_ , \new_[52964]_ , \new_[52965]_ , \new_[52968]_ ,
    \new_[52971]_ , \new_[52972]_ , \new_[52975]_ , \new_[52978]_ ,
    \new_[52979]_ , \new_[52980]_ , \new_[52983]_ , \new_[52986]_ ,
    \new_[52987]_ , \new_[52990]_ , \new_[52993]_ , \new_[52994]_ ,
    \new_[52995]_ , \new_[52998]_ , \new_[53001]_ , \new_[53002]_ ,
    \new_[53005]_ , \new_[53008]_ , \new_[53009]_ , \new_[53010]_ ,
    \new_[53013]_ , \new_[53016]_ , \new_[53017]_ , \new_[53020]_ ,
    \new_[53023]_ , \new_[53024]_ , \new_[53025]_ , \new_[53028]_ ,
    \new_[53031]_ , \new_[53032]_ , \new_[53035]_ , \new_[53038]_ ,
    \new_[53039]_ , \new_[53040]_ , \new_[53043]_ , \new_[53046]_ ,
    \new_[53047]_ , \new_[53050]_ , \new_[53053]_ , \new_[53054]_ ,
    \new_[53055]_ , \new_[53058]_ , \new_[53061]_ , \new_[53062]_ ,
    \new_[53065]_ , \new_[53068]_ , \new_[53069]_ , \new_[53070]_ ,
    \new_[53073]_ , \new_[53076]_ , \new_[53077]_ , \new_[53080]_ ,
    \new_[53083]_ , \new_[53084]_ , \new_[53085]_ , \new_[53088]_ ,
    \new_[53091]_ , \new_[53092]_ , \new_[53095]_ , \new_[53098]_ ,
    \new_[53099]_ , \new_[53100]_ , \new_[53103]_ , \new_[53106]_ ,
    \new_[53107]_ , \new_[53110]_ , \new_[53113]_ , \new_[53114]_ ,
    \new_[53115]_ , \new_[53118]_ , \new_[53121]_ , \new_[53122]_ ,
    \new_[53125]_ , \new_[53128]_ , \new_[53129]_ , \new_[53130]_ ,
    \new_[53133]_ , \new_[53136]_ , \new_[53137]_ , \new_[53140]_ ,
    \new_[53143]_ , \new_[53144]_ , \new_[53145]_ , \new_[53148]_ ,
    \new_[53151]_ , \new_[53152]_ , \new_[53155]_ , \new_[53158]_ ,
    \new_[53159]_ , \new_[53160]_ , \new_[53163]_ , \new_[53166]_ ,
    \new_[53167]_ , \new_[53170]_ , \new_[53173]_ , \new_[53174]_ ,
    \new_[53175]_ , \new_[53178]_ , \new_[53181]_ , \new_[53182]_ ,
    \new_[53185]_ , \new_[53188]_ , \new_[53189]_ , \new_[53190]_ ,
    \new_[53193]_ , \new_[53196]_ , \new_[53197]_ , \new_[53200]_ ,
    \new_[53203]_ , \new_[53204]_ , \new_[53205]_ , \new_[53208]_ ,
    \new_[53211]_ , \new_[53212]_ , \new_[53215]_ , \new_[53218]_ ,
    \new_[53219]_ , \new_[53220]_ , \new_[53223]_ , \new_[53226]_ ,
    \new_[53227]_ , \new_[53230]_ , \new_[53233]_ , \new_[53234]_ ,
    \new_[53235]_ , \new_[53238]_ , \new_[53241]_ , \new_[53242]_ ,
    \new_[53245]_ , \new_[53248]_ , \new_[53249]_ , \new_[53250]_ ,
    \new_[53253]_ , \new_[53256]_ , \new_[53257]_ , \new_[53260]_ ,
    \new_[53263]_ , \new_[53264]_ , \new_[53265]_ , \new_[53268]_ ,
    \new_[53271]_ , \new_[53272]_ , \new_[53275]_ , \new_[53278]_ ,
    \new_[53279]_ , \new_[53280]_ , \new_[53283]_ , \new_[53286]_ ,
    \new_[53287]_ , \new_[53290]_ , \new_[53293]_ , \new_[53294]_ ,
    \new_[53295]_ , \new_[53298]_ , \new_[53301]_ , \new_[53302]_ ,
    \new_[53305]_ , \new_[53308]_ , \new_[53309]_ , \new_[53310]_ ,
    \new_[53313]_ , \new_[53316]_ , \new_[53317]_ , \new_[53320]_ ,
    \new_[53323]_ , \new_[53324]_ , \new_[53325]_ , \new_[53328]_ ,
    \new_[53331]_ , \new_[53332]_ , \new_[53335]_ , \new_[53338]_ ,
    \new_[53339]_ , \new_[53340]_ , \new_[53343]_ , \new_[53346]_ ,
    \new_[53347]_ , \new_[53350]_ , \new_[53353]_ , \new_[53354]_ ,
    \new_[53355]_ , \new_[53358]_ , \new_[53361]_ , \new_[53362]_ ,
    \new_[53365]_ , \new_[53368]_ , \new_[53369]_ , \new_[53370]_ ,
    \new_[53373]_ , \new_[53376]_ , \new_[53377]_ , \new_[53380]_ ,
    \new_[53383]_ , \new_[53384]_ , \new_[53385]_ , \new_[53388]_ ,
    \new_[53391]_ , \new_[53392]_ , \new_[53395]_ , \new_[53398]_ ,
    \new_[53399]_ , \new_[53400]_ , \new_[53403]_ , \new_[53406]_ ,
    \new_[53407]_ , \new_[53410]_ , \new_[53413]_ , \new_[53414]_ ,
    \new_[53415]_ , \new_[53418]_ , \new_[53421]_ , \new_[53422]_ ,
    \new_[53425]_ , \new_[53428]_ , \new_[53429]_ , \new_[53430]_ ,
    \new_[53433]_ , \new_[53436]_ , \new_[53437]_ , \new_[53440]_ ,
    \new_[53443]_ , \new_[53444]_ , \new_[53445]_ , \new_[53448]_ ,
    \new_[53451]_ , \new_[53452]_ , \new_[53455]_ , \new_[53458]_ ,
    \new_[53459]_ , \new_[53460]_ , \new_[53463]_ , \new_[53466]_ ,
    \new_[53467]_ , \new_[53470]_ , \new_[53473]_ , \new_[53474]_ ,
    \new_[53475]_ , \new_[53478]_ , \new_[53481]_ , \new_[53482]_ ,
    \new_[53485]_ , \new_[53488]_ , \new_[53489]_ , \new_[53490]_ ,
    \new_[53493]_ , \new_[53496]_ , \new_[53497]_ , \new_[53500]_ ,
    \new_[53503]_ , \new_[53504]_ , \new_[53505]_ , \new_[53508]_ ,
    \new_[53511]_ , \new_[53512]_ , \new_[53515]_ , \new_[53518]_ ,
    \new_[53519]_ , \new_[53520]_ , \new_[53523]_ , \new_[53526]_ ,
    \new_[53527]_ , \new_[53530]_ , \new_[53533]_ , \new_[53534]_ ,
    \new_[53535]_ , \new_[53538]_ , \new_[53541]_ , \new_[53542]_ ,
    \new_[53545]_ , \new_[53548]_ , \new_[53549]_ , \new_[53550]_ ,
    \new_[53553]_ , \new_[53556]_ , \new_[53557]_ , \new_[53560]_ ,
    \new_[53563]_ , \new_[53564]_ , \new_[53565]_ , \new_[53568]_ ,
    \new_[53571]_ , \new_[53572]_ , \new_[53575]_ , \new_[53578]_ ,
    \new_[53579]_ , \new_[53580]_ , \new_[53583]_ , \new_[53586]_ ,
    \new_[53587]_ , \new_[53590]_ , \new_[53593]_ , \new_[53594]_ ,
    \new_[53595]_ , \new_[53598]_ , \new_[53601]_ , \new_[53602]_ ,
    \new_[53605]_ , \new_[53608]_ , \new_[53609]_ , \new_[53610]_ ,
    \new_[53613]_ , \new_[53616]_ , \new_[53617]_ , \new_[53620]_ ,
    \new_[53623]_ , \new_[53624]_ , \new_[53625]_ , \new_[53628]_ ,
    \new_[53631]_ , \new_[53632]_ , \new_[53635]_ , \new_[53638]_ ,
    \new_[53639]_ , \new_[53640]_ , \new_[53643]_ , \new_[53646]_ ,
    \new_[53647]_ , \new_[53650]_ , \new_[53653]_ , \new_[53654]_ ,
    \new_[53655]_ , \new_[53658]_ , \new_[53661]_ , \new_[53662]_ ,
    \new_[53665]_ , \new_[53668]_ , \new_[53669]_ , \new_[53670]_ ,
    \new_[53673]_ , \new_[53676]_ , \new_[53677]_ , \new_[53680]_ ,
    \new_[53683]_ , \new_[53684]_ , \new_[53685]_ , \new_[53688]_ ,
    \new_[53691]_ , \new_[53692]_ , \new_[53695]_ , \new_[53698]_ ,
    \new_[53699]_ , \new_[53700]_ , \new_[53703]_ , \new_[53706]_ ,
    \new_[53707]_ , \new_[53710]_ , \new_[53713]_ , \new_[53714]_ ,
    \new_[53715]_ , \new_[53718]_ , \new_[53721]_ , \new_[53722]_ ,
    \new_[53725]_ , \new_[53728]_ , \new_[53729]_ , \new_[53730]_ ,
    \new_[53733]_ , \new_[53736]_ , \new_[53737]_ , \new_[53740]_ ,
    \new_[53743]_ , \new_[53744]_ , \new_[53745]_ , \new_[53748]_ ,
    \new_[53751]_ , \new_[53752]_ , \new_[53755]_ , \new_[53758]_ ,
    \new_[53759]_ , \new_[53760]_ , \new_[53763]_ , \new_[53766]_ ,
    \new_[53767]_ , \new_[53770]_ , \new_[53773]_ , \new_[53774]_ ,
    \new_[53775]_ , \new_[53778]_ , \new_[53781]_ , \new_[53782]_ ,
    \new_[53785]_ , \new_[53788]_ , \new_[53789]_ , \new_[53790]_ ,
    \new_[53793]_ , \new_[53796]_ , \new_[53797]_ , \new_[53800]_ ,
    \new_[53803]_ , \new_[53804]_ , \new_[53805]_ , \new_[53808]_ ,
    \new_[53811]_ , \new_[53812]_ , \new_[53815]_ , \new_[53818]_ ,
    \new_[53819]_ , \new_[53820]_ , \new_[53823]_ , \new_[53826]_ ,
    \new_[53827]_ , \new_[53830]_ , \new_[53833]_ , \new_[53834]_ ,
    \new_[53835]_ , \new_[53838]_ , \new_[53841]_ , \new_[53842]_ ,
    \new_[53845]_ , \new_[53848]_ , \new_[53849]_ , \new_[53850]_ ,
    \new_[53853]_ , \new_[53856]_ , \new_[53857]_ , \new_[53860]_ ,
    \new_[53863]_ , \new_[53864]_ , \new_[53865]_ , \new_[53868]_ ,
    \new_[53871]_ , \new_[53872]_ , \new_[53875]_ , \new_[53878]_ ,
    \new_[53879]_ , \new_[53880]_ , \new_[53883]_ , \new_[53886]_ ,
    \new_[53887]_ , \new_[53890]_ , \new_[53893]_ , \new_[53894]_ ,
    \new_[53895]_ , \new_[53898]_ , \new_[53901]_ , \new_[53902]_ ,
    \new_[53905]_ , \new_[53908]_ , \new_[53909]_ , \new_[53910]_ ,
    \new_[53913]_ , \new_[53916]_ , \new_[53917]_ , \new_[53920]_ ,
    \new_[53923]_ , \new_[53924]_ , \new_[53925]_ , \new_[53928]_ ,
    \new_[53931]_ , \new_[53932]_ , \new_[53935]_ , \new_[53938]_ ,
    \new_[53939]_ , \new_[53940]_ , \new_[53943]_ , \new_[53946]_ ,
    \new_[53947]_ , \new_[53950]_ , \new_[53953]_ , \new_[53954]_ ,
    \new_[53955]_ , \new_[53958]_ , \new_[53961]_ , \new_[53962]_ ,
    \new_[53965]_ , \new_[53968]_ , \new_[53969]_ , \new_[53970]_ ,
    \new_[53973]_ , \new_[53976]_ , \new_[53977]_ , \new_[53980]_ ,
    \new_[53983]_ , \new_[53984]_ , \new_[53985]_ , \new_[53988]_ ,
    \new_[53991]_ , \new_[53992]_ , \new_[53995]_ , \new_[53998]_ ,
    \new_[53999]_ , \new_[54000]_ , \new_[54003]_ , \new_[54006]_ ,
    \new_[54007]_ , \new_[54010]_ , \new_[54013]_ , \new_[54014]_ ,
    \new_[54015]_ , \new_[54018]_ , \new_[54021]_ , \new_[54022]_ ,
    \new_[54025]_ , \new_[54028]_ , \new_[54029]_ , \new_[54030]_ ,
    \new_[54033]_ , \new_[54036]_ , \new_[54037]_ , \new_[54040]_ ,
    \new_[54043]_ , \new_[54044]_ , \new_[54045]_ , \new_[54048]_ ,
    \new_[54051]_ , \new_[54052]_ , \new_[54055]_ , \new_[54058]_ ,
    \new_[54059]_ , \new_[54060]_ , \new_[54063]_ , \new_[54066]_ ,
    \new_[54067]_ , \new_[54070]_ , \new_[54073]_ , \new_[54074]_ ,
    \new_[54075]_ , \new_[54078]_ , \new_[54081]_ , \new_[54082]_ ,
    \new_[54085]_ , \new_[54088]_ , \new_[54089]_ , \new_[54090]_ ,
    \new_[54093]_ , \new_[54096]_ , \new_[54097]_ , \new_[54100]_ ,
    \new_[54103]_ , \new_[54104]_ , \new_[54105]_ , \new_[54108]_ ,
    \new_[54111]_ , \new_[54112]_ , \new_[54115]_ , \new_[54118]_ ,
    \new_[54119]_ , \new_[54120]_ , \new_[54123]_ , \new_[54126]_ ,
    \new_[54127]_ , \new_[54130]_ , \new_[54133]_ , \new_[54134]_ ,
    \new_[54135]_ , \new_[54138]_ , \new_[54141]_ , \new_[54142]_ ,
    \new_[54145]_ , \new_[54148]_ , \new_[54149]_ , \new_[54150]_ ,
    \new_[54153]_ , \new_[54156]_ , \new_[54157]_ , \new_[54160]_ ,
    \new_[54163]_ , \new_[54164]_ , \new_[54165]_ , \new_[54168]_ ,
    \new_[54171]_ , \new_[54172]_ , \new_[54175]_ , \new_[54178]_ ,
    \new_[54179]_ , \new_[54180]_ , \new_[54183]_ , \new_[54186]_ ,
    \new_[54187]_ , \new_[54190]_ , \new_[54193]_ , \new_[54194]_ ,
    \new_[54195]_ , \new_[54198]_ , \new_[54201]_ , \new_[54202]_ ,
    \new_[54205]_ , \new_[54208]_ , \new_[54209]_ , \new_[54210]_ ,
    \new_[54213]_ , \new_[54216]_ , \new_[54217]_ , \new_[54220]_ ,
    \new_[54223]_ , \new_[54224]_ , \new_[54225]_ , \new_[54228]_ ,
    \new_[54231]_ , \new_[54232]_ , \new_[54235]_ , \new_[54238]_ ,
    \new_[54239]_ , \new_[54240]_ , \new_[54243]_ , \new_[54246]_ ,
    \new_[54247]_ , \new_[54250]_ , \new_[54253]_ , \new_[54254]_ ,
    \new_[54255]_ , \new_[54258]_ , \new_[54261]_ , \new_[54262]_ ,
    \new_[54265]_ , \new_[54268]_ , \new_[54269]_ , \new_[54270]_ ,
    \new_[54273]_ , \new_[54276]_ , \new_[54277]_ , \new_[54280]_ ,
    \new_[54283]_ , \new_[54284]_ , \new_[54285]_ , \new_[54288]_ ,
    \new_[54291]_ , \new_[54292]_ , \new_[54295]_ , \new_[54298]_ ,
    \new_[54299]_ , \new_[54300]_ , \new_[54303]_ , \new_[54306]_ ,
    \new_[54307]_ , \new_[54310]_ , \new_[54313]_ , \new_[54314]_ ,
    \new_[54315]_ , \new_[54318]_ , \new_[54321]_ , \new_[54322]_ ,
    \new_[54325]_ , \new_[54328]_ , \new_[54329]_ , \new_[54330]_ ,
    \new_[54333]_ , \new_[54336]_ , \new_[54337]_ , \new_[54340]_ ,
    \new_[54343]_ , \new_[54344]_ , \new_[54345]_ , \new_[54348]_ ,
    \new_[54351]_ , \new_[54352]_ , \new_[54355]_ , \new_[54358]_ ,
    \new_[54359]_ , \new_[54360]_ , \new_[54363]_ , \new_[54366]_ ,
    \new_[54367]_ , \new_[54370]_ , \new_[54373]_ , \new_[54374]_ ,
    \new_[54375]_ , \new_[54378]_ , \new_[54381]_ , \new_[54382]_ ,
    \new_[54385]_ , \new_[54388]_ , \new_[54389]_ , \new_[54390]_ ,
    \new_[54393]_ , \new_[54396]_ , \new_[54397]_ , \new_[54400]_ ,
    \new_[54403]_ , \new_[54404]_ , \new_[54405]_ , \new_[54408]_ ,
    \new_[54411]_ , \new_[54412]_ , \new_[54415]_ , \new_[54418]_ ,
    \new_[54419]_ , \new_[54420]_ , \new_[54423]_ , \new_[54426]_ ,
    \new_[54427]_ , \new_[54430]_ , \new_[54433]_ , \new_[54434]_ ,
    \new_[54435]_ , \new_[54438]_ , \new_[54441]_ , \new_[54442]_ ,
    \new_[54445]_ , \new_[54448]_ , \new_[54449]_ , \new_[54450]_ ,
    \new_[54453]_ , \new_[54456]_ , \new_[54457]_ , \new_[54460]_ ,
    \new_[54463]_ , \new_[54464]_ , \new_[54465]_ , \new_[54468]_ ,
    \new_[54471]_ , \new_[54472]_ , \new_[54475]_ , \new_[54478]_ ,
    \new_[54479]_ , \new_[54480]_ , \new_[54483]_ , \new_[54486]_ ,
    \new_[54487]_ , \new_[54490]_ , \new_[54493]_ , \new_[54494]_ ,
    \new_[54495]_ , \new_[54498]_ , \new_[54501]_ , \new_[54502]_ ,
    \new_[54505]_ , \new_[54508]_ , \new_[54509]_ , \new_[54510]_ ,
    \new_[54513]_ , \new_[54516]_ , \new_[54517]_ , \new_[54520]_ ,
    \new_[54523]_ , \new_[54524]_ , \new_[54525]_ , \new_[54528]_ ,
    \new_[54531]_ , \new_[54532]_ , \new_[54535]_ , \new_[54538]_ ,
    \new_[54539]_ , \new_[54540]_ , \new_[54543]_ , \new_[54546]_ ,
    \new_[54547]_ , \new_[54550]_ , \new_[54553]_ , \new_[54554]_ ,
    \new_[54555]_ , \new_[54558]_ , \new_[54561]_ , \new_[54562]_ ,
    \new_[54565]_ , \new_[54568]_ , \new_[54569]_ , \new_[54570]_ ,
    \new_[54573]_ , \new_[54576]_ , \new_[54577]_ , \new_[54580]_ ,
    \new_[54583]_ , \new_[54584]_ , \new_[54585]_ , \new_[54588]_ ,
    \new_[54591]_ , \new_[54592]_ , \new_[54595]_ , \new_[54598]_ ,
    \new_[54599]_ , \new_[54600]_ , \new_[54603]_ , \new_[54606]_ ,
    \new_[54607]_ , \new_[54610]_ , \new_[54613]_ , \new_[54614]_ ,
    \new_[54615]_ , \new_[54618]_ , \new_[54621]_ , \new_[54622]_ ,
    \new_[54625]_ , \new_[54628]_ , \new_[54629]_ , \new_[54630]_ ,
    \new_[54633]_ , \new_[54636]_ , \new_[54637]_ , \new_[54640]_ ,
    \new_[54643]_ , \new_[54644]_ , \new_[54645]_ , \new_[54648]_ ,
    \new_[54651]_ , \new_[54652]_ , \new_[54655]_ , \new_[54658]_ ,
    \new_[54659]_ , \new_[54660]_ , \new_[54663]_ , \new_[54666]_ ,
    \new_[54667]_ , \new_[54670]_ , \new_[54673]_ , \new_[54674]_ ,
    \new_[54675]_ , \new_[54678]_ , \new_[54681]_ , \new_[54682]_ ,
    \new_[54685]_ , \new_[54688]_ , \new_[54689]_ , \new_[54690]_ ,
    \new_[54693]_ , \new_[54696]_ , \new_[54697]_ , \new_[54700]_ ,
    \new_[54703]_ , \new_[54704]_ , \new_[54705]_ , \new_[54708]_ ,
    \new_[54711]_ , \new_[54712]_ , \new_[54715]_ , \new_[54718]_ ,
    \new_[54719]_ , \new_[54720]_ , \new_[54723]_ , \new_[54726]_ ,
    \new_[54727]_ , \new_[54730]_ , \new_[54733]_ , \new_[54734]_ ,
    \new_[54735]_ , \new_[54738]_ , \new_[54741]_ , \new_[54742]_ ,
    \new_[54745]_ , \new_[54748]_ , \new_[54749]_ , \new_[54750]_ ,
    \new_[54753]_ , \new_[54756]_ , \new_[54757]_ , \new_[54760]_ ,
    \new_[54763]_ , \new_[54764]_ , \new_[54765]_ , \new_[54768]_ ,
    \new_[54771]_ , \new_[54772]_ , \new_[54775]_ , \new_[54778]_ ,
    \new_[54779]_ , \new_[54780]_ , \new_[54783]_ , \new_[54786]_ ,
    \new_[54787]_ , \new_[54790]_ , \new_[54793]_ , \new_[54794]_ ,
    \new_[54795]_ , \new_[54798]_ , \new_[54801]_ , \new_[54802]_ ,
    \new_[54805]_ , \new_[54808]_ , \new_[54809]_ , \new_[54810]_ ,
    \new_[54813]_ , \new_[54816]_ , \new_[54817]_ , \new_[54820]_ ,
    \new_[54823]_ , \new_[54824]_ , \new_[54825]_ , \new_[54828]_ ,
    \new_[54831]_ , \new_[54832]_ , \new_[54835]_ , \new_[54838]_ ,
    \new_[54839]_ , \new_[54840]_ , \new_[54843]_ , \new_[54846]_ ,
    \new_[54847]_ , \new_[54850]_ , \new_[54853]_ , \new_[54854]_ ,
    \new_[54855]_ , \new_[54858]_ , \new_[54861]_ , \new_[54862]_ ,
    \new_[54865]_ , \new_[54868]_ , \new_[54869]_ , \new_[54870]_ ,
    \new_[54873]_ , \new_[54876]_ , \new_[54877]_ , \new_[54880]_ ,
    \new_[54883]_ , \new_[54884]_ , \new_[54885]_ , \new_[54888]_ ,
    \new_[54891]_ , \new_[54892]_ , \new_[54895]_ , \new_[54898]_ ,
    \new_[54899]_ , \new_[54900]_ , \new_[54903]_ , \new_[54906]_ ,
    \new_[54907]_ , \new_[54910]_ , \new_[54913]_ , \new_[54914]_ ,
    \new_[54915]_ , \new_[54918]_ , \new_[54921]_ , \new_[54922]_ ,
    \new_[54925]_ , \new_[54928]_ , \new_[54929]_ , \new_[54930]_ ,
    \new_[54933]_ , \new_[54936]_ , \new_[54937]_ , \new_[54940]_ ,
    \new_[54943]_ , \new_[54944]_ , \new_[54945]_ , \new_[54948]_ ,
    \new_[54951]_ , \new_[54952]_ , \new_[54955]_ , \new_[54958]_ ,
    \new_[54959]_ , \new_[54960]_ , \new_[54963]_ , \new_[54966]_ ,
    \new_[54967]_ , \new_[54970]_ , \new_[54973]_ , \new_[54974]_ ,
    \new_[54975]_ , \new_[54978]_ , \new_[54981]_ , \new_[54982]_ ,
    \new_[54985]_ , \new_[54988]_ , \new_[54989]_ , \new_[54990]_ ,
    \new_[54993]_ , \new_[54996]_ , \new_[54997]_ , \new_[55000]_ ,
    \new_[55003]_ , \new_[55004]_ , \new_[55005]_ , \new_[55008]_ ,
    \new_[55011]_ , \new_[55012]_ , \new_[55015]_ , \new_[55018]_ ,
    \new_[55019]_ , \new_[55020]_ , \new_[55023]_ , \new_[55026]_ ,
    \new_[55027]_ , \new_[55030]_ , \new_[55033]_ , \new_[55034]_ ,
    \new_[55035]_ , \new_[55038]_ , \new_[55041]_ , \new_[55042]_ ,
    \new_[55045]_ , \new_[55048]_ , \new_[55049]_ , \new_[55050]_ ,
    \new_[55053]_ , \new_[55056]_ , \new_[55057]_ , \new_[55060]_ ,
    \new_[55063]_ , \new_[55064]_ , \new_[55065]_ , \new_[55068]_ ,
    \new_[55071]_ , \new_[55072]_ , \new_[55075]_ , \new_[55078]_ ,
    \new_[55079]_ , \new_[55080]_ , \new_[55083]_ , \new_[55086]_ ,
    \new_[55087]_ , \new_[55090]_ , \new_[55093]_ , \new_[55094]_ ,
    \new_[55095]_ , \new_[55098]_ , \new_[55101]_ , \new_[55102]_ ,
    \new_[55105]_ , \new_[55108]_ , \new_[55109]_ , \new_[55110]_ ,
    \new_[55113]_ , \new_[55116]_ , \new_[55117]_ , \new_[55120]_ ,
    \new_[55123]_ , \new_[55124]_ , \new_[55125]_ , \new_[55128]_ ,
    \new_[55131]_ , \new_[55132]_ , \new_[55135]_ , \new_[55138]_ ,
    \new_[55139]_ , \new_[55140]_ , \new_[55143]_ , \new_[55146]_ ,
    \new_[55147]_ , \new_[55150]_ , \new_[55153]_ , \new_[55154]_ ,
    \new_[55155]_ , \new_[55158]_ , \new_[55161]_ , \new_[55162]_ ,
    \new_[55165]_ , \new_[55168]_ , \new_[55169]_ , \new_[55170]_ ,
    \new_[55173]_ , \new_[55176]_ , \new_[55177]_ , \new_[55180]_ ,
    \new_[55183]_ , \new_[55184]_ , \new_[55185]_ , \new_[55188]_ ,
    \new_[55191]_ , \new_[55192]_ , \new_[55195]_ , \new_[55198]_ ,
    \new_[55199]_ , \new_[55200]_ , \new_[55203]_ , \new_[55206]_ ,
    \new_[55207]_ , \new_[55210]_ , \new_[55213]_ , \new_[55214]_ ,
    \new_[55215]_ , \new_[55218]_ , \new_[55221]_ , \new_[55222]_ ,
    \new_[55225]_ , \new_[55228]_ , \new_[55229]_ , \new_[55230]_ ,
    \new_[55233]_ , \new_[55236]_ , \new_[55237]_ , \new_[55240]_ ,
    \new_[55243]_ , \new_[55244]_ , \new_[55245]_ , \new_[55248]_ ,
    \new_[55251]_ , \new_[55252]_ , \new_[55255]_ , \new_[55258]_ ,
    \new_[55259]_ , \new_[55260]_ , \new_[55263]_ , \new_[55266]_ ,
    \new_[55267]_ , \new_[55270]_ , \new_[55273]_ , \new_[55274]_ ,
    \new_[55275]_ , \new_[55278]_ , \new_[55281]_ , \new_[55282]_ ,
    \new_[55285]_ , \new_[55288]_ , \new_[55289]_ , \new_[55290]_ ,
    \new_[55293]_ , \new_[55296]_ , \new_[55297]_ , \new_[55300]_ ,
    \new_[55303]_ , \new_[55304]_ , \new_[55305]_ , \new_[55308]_ ,
    \new_[55311]_ , \new_[55312]_ , \new_[55315]_ , \new_[55318]_ ,
    \new_[55319]_ , \new_[55320]_ , \new_[55323]_ , \new_[55326]_ ,
    \new_[55327]_ , \new_[55330]_ , \new_[55333]_ , \new_[55334]_ ,
    \new_[55335]_ , \new_[55338]_ , \new_[55341]_ , \new_[55342]_ ,
    \new_[55345]_ , \new_[55348]_ , \new_[55349]_ , \new_[55350]_ ,
    \new_[55353]_ , \new_[55356]_ , \new_[55357]_ , \new_[55360]_ ,
    \new_[55363]_ , \new_[55364]_ , \new_[55365]_ , \new_[55368]_ ,
    \new_[55371]_ , \new_[55372]_ , \new_[55375]_ , \new_[55378]_ ,
    \new_[55379]_ , \new_[55380]_ , \new_[55383]_ , \new_[55386]_ ,
    \new_[55387]_ , \new_[55390]_ , \new_[55393]_ , \new_[55394]_ ,
    \new_[55395]_ , \new_[55398]_ , \new_[55401]_ , \new_[55402]_ ,
    \new_[55405]_ , \new_[55408]_ , \new_[55409]_ , \new_[55410]_ ,
    \new_[55413]_ , \new_[55416]_ , \new_[55417]_ , \new_[55420]_ ,
    \new_[55423]_ , \new_[55424]_ , \new_[55425]_ , \new_[55428]_ ,
    \new_[55431]_ , \new_[55432]_ , \new_[55435]_ , \new_[55438]_ ,
    \new_[55439]_ , \new_[55440]_ , \new_[55443]_ , \new_[55446]_ ,
    \new_[55447]_ , \new_[55450]_ , \new_[55453]_ , \new_[55454]_ ,
    \new_[55455]_ , \new_[55458]_ , \new_[55461]_ , \new_[55462]_ ,
    \new_[55465]_ , \new_[55468]_ , \new_[55469]_ , \new_[55470]_ ,
    \new_[55473]_ , \new_[55476]_ , \new_[55477]_ , \new_[55480]_ ,
    \new_[55483]_ , \new_[55484]_ , \new_[55485]_ , \new_[55488]_ ,
    \new_[55491]_ , \new_[55492]_ , \new_[55495]_ , \new_[55498]_ ,
    \new_[55499]_ , \new_[55500]_ , \new_[55503]_ , \new_[55506]_ ,
    \new_[55507]_ , \new_[55510]_ , \new_[55513]_ , \new_[55514]_ ,
    \new_[55515]_ , \new_[55518]_ , \new_[55521]_ , \new_[55522]_ ,
    \new_[55525]_ , \new_[55528]_ , \new_[55529]_ , \new_[55530]_ ,
    \new_[55533]_ , \new_[55536]_ , \new_[55537]_ , \new_[55540]_ ,
    \new_[55543]_ , \new_[55544]_ , \new_[55545]_ , \new_[55548]_ ,
    \new_[55551]_ , \new_[55552]_ , \new_[55555]_ , \new_[55558]_ ,
    \new_[55559]_ , \new_[55560]_ , \new_[55563]_ , \new_[55566]_ ,
    \new_[55567]_ , \new_[55570]_ , \new_[55573]_ , \new_[55574]_ ,
    \new_[55575]_ , \new_[55578]_ , \new_[55581]_ , \new_[55582]_ ,
    \new_[55585]_ , \new_[55588]_ , \new_[55589]_ , \new_[55590]_ ,
    \new_[55593]_ , \new_[55596]_ , \new_[55597]_ , \new_[55600]_ ,
    \new_[55603]_ , \new_[55604]_ , \new_[55605]_ , \new_[55608]_ ,
    \new_[55611]_ , \new_[55612]_ , \new_[55615]_ , \new_[55618]_ ,
    \new_[55619]_ , \new_[55620]_ , \new_[55623]_ , \new_[55626]_ ,
    \new_[55627]_ , \new_[55630]_ , \new_[55633]_ , \new_[55634]_ ,
    \new_[55635]_ , \new_[55638]_ , \new_[55641]_ , \new_[55642]_ ,
    \new_[55645]_ , \new_[55648]_ , \new_[55649]_ , \new_[55650]_ ,
    \new_[55653]_ , \new_[55656]_ , \new_[55657]_ , \new_[55660]_ ,
    \new_[55663]_ , \new_[55664]_ , \new_[55665]_ , \new_[55668]_ ,
    \new_[55671]_ , \new_[55672]_ , \new_[55675]_ , \new_[55678]_ ,
    \new_[55679]_ , \new_[55680]_ , \new_[55683]_ , \new_[55686]_ ,
    \new_[55687]_ , \new_[55690]_ , \new_[55693]_ , \new_[55694]_ ,
    \new_[55695]_ , \new_[55698]_ , \new_[55701]_ , \new_[55702]_ ,
    \new_[55705]_ , \new_[55708]_ , \new_[55709]_ , \new_[55710]_ ,
    \new_[55713]_ , \new_[55716]_ , \new_[55717]_ , \new_[55720]_ ,
    \new_[55723]_ , \new_[55724]_ , \new_[55725]_ , \new_[55728]_ ,
    \new_[55731]_ , \new_[55732]_ , \new_[55735]_ , \new_[55738]_ ,
    \new_[55739]_ , \new_[55740]_ , \new_[55743]_ , \new_[55746]_ ,
    \new_[55747]_ , \new_[55750]_ , \new_[55753]_ , \new_[55754]_ ,
    \new_[55755]_ , \new_[55758]_ , \new_[55761]_ , \new_[55762]_ ,
    \new_[55765]_ , \new_[55768]_ , \new_[55769]_ , \new_[55770]_ ,
    \new_[55773]_ , \new_[55776]_ , \new_[55777]_ , \new_[55780]_ ,
    \new_[55783]_ , \new_[55784]_ , \new_[55785]_ , \new_[55788]_ ,
    \new_[55791]_ , \new_[55792]_ , \new_[55795]_ , \new_[55798]_ ,
    \new_[55799]_ , \new_[55800]_ , \new_[55803]_ , \new_[55806]_ ,
    \new_[55807]_ , \new_[55810]_ , \new_[55813]_ , \new_[55814]_ ,
    \new_[55815]_ , \new_[55818]_ , \new_[55821]_ , \new_[55822]_ ,
    \new_[55825]_ , \new_[55828]_ , \new_[55829]_ , \new_[55830]_ ,
    \new_[55833]_ , \new_[55836]_ , \new_[55837]_ , \new_[55840]_ ,
    \new_[55843]_ , \new_[55844]_ , \new_[55845]_ , \new_[55848]_ ,
    \new_[55851]_ , \new_[55852]_ , \new_[55855]_ , \new_[55858]_ ,
    \new_[55859]_ , \new_[55860]_ , \new_[55863]_ , \new_[55866]_ ,
    \new_[55867]_ , \new_[55870]_ , \new_[55873]_ , \new_[55874]_ ,
    \new_[55875]_ , \new_[55878]_ , \new_[55881]_ , \new_[55882]_ ,
    \new_[55885]_ , \new_[55888]_ , \new_[55889]_ , \new_[55890]_ ,
    \new_[55893]_ , \new_[55896]_ , \new_[55897]_ , \new_[55900]_ ,
    \new_[55903]_ , \new_[55904]_ , \new_[55905]_ , \new_[55908]_ ,
    \new_[55911]_ , \new_[55912]_ , \new_[55915]_ , \new_[55918]_ ,
    \new_[55919]_ , \new_[55920]_ , \new_[55923]_ , \new_[55926]_ ,
    \new_[55927]_ , \new_[55930]_ , \new_[55933]_ , \new_[55934]_ ,
    \new_[55935]_ , \new_[55938]_ , \new_[55941]_ , \new_[55942]_ ,
    \new_[55945]_ , \new_[55948]_ , \new_[55949]_ , \new_[55950]_ ,
    \new_[55953]_ , \new_[55956]_ , \new_[55957]_ , \new_[55960]_ ,
    \new_[55963]_ , \new_[55964]_ , \new_[55965]_ , \new_[55968]_ ,
    \new_[55971]_ , \new_[55972]_ , \new_[55975]_ , \new_[55978]_ ,
    \new_[55979]_ , \new_[55980]_ , \new_[55983]_ , \new_[55986]_ ,
    \new_[55987]_ , \new_[55990]_ , \new_[55993]_ , \new_[55994]_ ,
    \new_[55995]_ , \new_[55998]_ , \new_[56001]_ , \new_[56002]_ ,
    \new_[56005]_ , \new_[56008]_ , \new_[56009]_ , \new_[56010]_ ,
    \new_[56013]_ , \new_[56016]_ , \new_[56017]_ , \new_[56020]_ ,
    \new_[56023]_ , \new_[56024]_ , \new_[56025]_ , \new_[56028]_ ,
    \new_[56031]_ , \new_[56032]_ , \new_[56035]_ , \new_[56038]_ ,
    \new_[56039]_ , \new_[56040]_ , \new_[56043]_ , \new_[56046]_ ,
    \new_[56047]_ , \new_[56050]_ , \new_[56053]_ , \new_[56054]_ ,
    \new_[56055]_ , \new_[56058]_ , \new_[56061]_ , \new_[56062]_ ,
    \new_[56065]_ , \new_[56068]_ , \new_[56069]_ , \new_[56070]_ ,
    \new_[56073]_ , \new_[56076]_ , \new_[56077]_ , \new_[56080]_ ,
    \new_[56083]_ , \new_[56084]_ , \new_[56085]_ , \new_[56088]_ ,
    \new_[56091]_ , \new_[56092]_ , \new_[56095]_ , \new_[56098]_ ,
    \new_[56099]_ , \new_[56100]_ , \new_[56103]_ , \new_[56106]_ ,
    \new_[56107]_ , \new_[56110]_ , \new_[56113]_ , \new_[56114]_ ,
    \new_[56115]_ , \new_[56118]_ , \new_[56121]_ , \new_[56122]_ ,
    \new_[56125]_ , \new_[56128]_ , \new_[56129]_ , \new_[56130]_ ,
    \new_[56133]_ , \new_[56136]_ , \new_[56137]_ , \new_[56140]_ ,
    \new_[56143]_ , \new_[56144]_ , \new_[56145]_ , \new_[56148]_ ,
    \new_[56151]_ , \new_[56152]_ , \new_[56155]_ , \new_[56158]_ ,
    \new_[56159]_ , \new_[56160]_ , \new_[56163]_ , \new_[56166]_ ,
    \new_[56167]_ , \new_[56170]_ , \new_[56173]_ , \new_[56174]_ ,
    \new_[56175]_ , \new_[56178]_ , \new_[56181]_ , \new_[56182]_ ,
    \new_[56185]_ , \new_[56188]_ , \new_[56189]_ , \new_[56190]_ ,
    \new_[56193]_ , \new_[56196]_ , \new_[56197]_ , \new_[56200]_ ,
    \new_[56203]_ , \new_[56204]_ , \new_[56205]_ , \new_[56208]_ ,
    \new_[56211]_ , \new_[56212]_ , \new_[56215]_ , \new_[56218]_ ,
    \new_[56219]_ , \new_[56220]_ , \new_[56223]_ , \new_[56226]_ ,
    \new_[56227]_ , \new_[56230]_ , \new_[56233]_ , \new_[56234]_ ,
    \new_[56235]_ , \new_[56238]_ , \new_[56241]_ , \new_[56242]_ ,
    \new_[56245]_ , \new_[56248]_ , \new_[56249]_ , \new_[56250]_ ,
    \new_[56253]_ , \new_[56256]_ , \new_[56257]_ , \new_[56260]_ ,
    \new_[56263]_ , \new_[56264]_ , \new_[56265]_ , \new_[56268]_ ,
    \new_[56271]_ , \new_[56272]_ , \new_[56275]_ , \new_[56278]_ ,
    \new_[56279]_ , \new_[56280]_ , \new_[56283]_ , \new_[56286]_ ,
    \new_[56287]_ , \new_[56290]_ , \new_[56293]_ , \new_[56294]_ ,
    \new_[56295]_ , \new_[56298]_ , \new_[56301]_ , \new_[56302]_ ,
    \new_[56305]_ , \new_[56308]_ , \new_[56309]_ , \new_[56310]_ ,
    \new_[56313]_ , \new_[56316]_ , \new_[56317]_ , \new_[56320]_ ,
    \new_[56323]_ , \new_[56324]_ , \new_[56325]_ , \new_[56328]_ ,
    \new_[56331]_ , \new_[56332]_ , \new_[56335]_ , \new_[56338]_ ,
    \new_[56339]_ , \new_[56340]_ , \new_[56343]_ , \new_[56346]_ ,
    \new_[56347]_ , \new_[56350]_ , \new_[56353]_ , \new_[56354]_ ,
    \new_[56355]_ , \new_[56358]_ , \new_[56361]_ , \new_[56362]_ ,
    \new_[56365]_ , \new_[56368]_ , \new_[56369]_ , \new_[56370]_ ,
    \new_[56373]_ , \new_[56376]_ , \new_[56377]_ , \new_[56380]_ ,
    \new_[56383]_ , \new_[56384]_ , \new_[56385]_ , \new_[56388]_ ,
    \new_[56391]_ , \new_[56392]_ , \new_[56395]_ , \new_[56398]_ ,
    \new_[56399]_ , \new_[56400]_ , \new_[56403]_ , \new_[56406]_ ,
    \new_[56407]_ , \new_[56410]_ , \new_[56413]_ , \new_[56414]_ ,
    \new_[56415]_ , \new_[56418]_ , \new_[56421]_ , \new_[56422]_ ,
    \new_[56425]_ , \new_[56428]_ , \new_[56429]_ , \new_[56430]_ ,
    \new_[56433]_ , \new_[56436]_ , \new_[56437]_ , \new_[56440]_ ,
    \new_[56443]_ , \new_[56444]_ , \new_[56445]_ , \new_[56448]_ ,
    \new_[56451]_ , \new_[56452]_ , \new_[56455]_ , \new_[56458]_ ,
    \new_[56459]_ , \new_[56460]_ , \new_[56463]_ , \new_[56466]_ ,
    \new_[56467]_ , \new_[56470]_ , \new_[56473]_ , \new_[56474]_ ,
    \new_[56475]_ , \new_[56478]_ , \new_[56481]_ , \new_[56482]_ ,
    \new_[56485]_ , \new_[56488]_ , \new_[56489]_ , \new_[56490]_ ,
    \new_[56493]_ , \new_[56496]_ , \new_[56497]_ , \new_[56500]_ ,
    \new_[56503]_ , \new_[56504]_ , \new_[56505]_ , \new_[56508]_ ,
    \new_[56511]_ , \new_[56512]_ , \new_[56515]_ , \new_[56518]_ ,
    \new_[56519]_ , \new_[56520]_ , \new_[56523]_ , \new_[56526]_ ,
    \new_[56527]_ , \new_[56530]_ , \new_[56533]_ , \new_[56534]_ ,
    \new_[56535]_ , \new_[56538]_ , \new_[56541]_ , \new_[56542]_ ,
    \new_[56545]_ , \new_[56548]_ , \new_[56549]_ , \new_[56550]_ ,
    \new_[56553]_ , \new_[56556]_ , \new_[56557]_ , \new_[56560]_ ,
    \new_[56563]_ , \new_[56564]_ , \new_[56565]_ , \new_[56568]_ ,
    \new_[56571]_ , \new_[56572]_ , \new_[56575]_ , \new_[56578]_ ,
    \new_[56579]_ , \new_[56580]_ , \new_[56583]_ , \new_[56586]_ ,
    \new_[56587]_ , \new_[56590]_ , \new_[56593]_ , \new_[56594]_ ,
    \new_[56595]_ , \new_[56598]_ , \new_[56601]_ , \new_[56602]_ ,
    \new_[56605]_ , \new_[56608]_ , \new_[56609]_ , \new_[56610]_ ,
    \new_[56613]_ , \new_[56616]_ , \new_[56617]_ , \new_[56620]_ ,
    \new_[56623]_ , \new_[56624]_ , \new_[56625]_ , \new_[56628]_ ,
    \new_[56631]_ , \new_[56632]_ , \new_[56635]_ , \new_[56638]_ ,
    \new_[56639]_ , \new_[56640]_ , \new_[56643]_ , \new_[56646]_ ,
    \new_[56647]_ , \new_[56650]_ , \new_[56653]_ , \new_[56654]_ ,
    \new_[56655]_ , \new_[56658]_ , \new_[56661]_ , \new_[56662]_ ,
    \new_[56665]_ , \new_[56668]_ , \new_[56669]_ , \new_[56670]_ ,
    \new_[56673]_ , \new_[56676]_ , \new_[56677]_ , \new_[56680]_ ,
    \new_[56683]_ , \new_[56684]_ , \new_[56685]_ , \new_[56688]_ ,
    \new_[56691]_ , \new_[56692]_ , \new_[56695]_ , \new_[56698]_ ,
    \new_[56699]_ , \new_[56700]_ , \new_[56703]_ , \new_[56706]_ ,
    \new_[56707]_ , \new_[56710]_ , \new_[56713]_ , \new_[56714]_ ,
    \new_[56715]_ , \new_[56718]_ , \new_[56721]_ , \new_[56722]_ ,
    \new_[56725]_ , \new_[56728]_ , \new_[56729]_ , \new_[56730]_ ,
    \new_[56733]_ , \new_[56736]_ , \new_[56737]_ , \new_[56740]_ ,
    \new_[56743]_ , \new_[56744]_ , \new_[56745]_ , \new_[56748]_ ,
    \new_[56751]_ , \new_[56752]_ , \new_[56755]_ , \new_[56758]_ ,
    \new_[56759]_ , \new_[56760]_ , \new_[56763]_ , \new_[56766]_ ,
    \new_[56767]_ , \new_[56770]_ , \new_[56773]_ , \new_[56774]_ ,
    \new_[56775]_ , \new_[56778]_ , \new_[56781]_ , \new_[56782]_ ,
    \new_[56785]_ , \new_[56788]_ , \new_[56789]_ , \new_[56790]_ ,
    \new_[56793]_ , \new_[56796]_ , \new_[56797]_ , \new_[56800]_ ,
    \new_[56803]_ , \new_[56804]_ , \new_[56805]_ , \new_[56808]_ ,
    \new_[56811]_ , \new_[56812]_ , \new_[56815]_ , \new_[56818]_ ,
    \new_[56819]_ , \new_[56820]_ , \new_[56823]_ , \new_[56826]_ ,
    \new_[56827]_ , \new_[56830]_ , \new_[56833]_ , \new_[56834]_ ,
    \new_[56835]_ , \new_[56838]_ , \new_[56841]_ , \new_[56842]_ ,
    \new_[56845]_ , \new_[56848]_ , \new_[56849]_ , \new_[56850]_ ,
    \new_[56853]_ , \new_[56856]_ , \new_[56857]_ , \new_[56860]_ ,
    \new_[56863]_ , \new_[56864]_ , \new_[56865]_ , \new_[56868]_ ,
    \new_[56871]_ , \new_[56872]_ , \new_[56875]_ , \new_[56878]_ ,
    \new_[56879]_ , \new_[56880]_ , \new_[56883]_ , \new_[56886]_ ,
    \new_[56887]_ , \new_[56890]_ , \new_[56893]_ , \new_[56894]_ ,
    \new_[56895]_ , \new_[56898]_ , \new_[56901]_ , \new_[56902]_ ,
    \new_[56905]_ , \new_[56908]_ , \new_[56909]_ , \new_[56910]_ ,
    \new_[56913]_ , \new_[56916]_ , \new_[56917]_ , \new_[56920]_ ,
    \new_[56923]_ , \new_[56924]_ , \new_[56925]_ , \new_[56928]_ ,
    \new_[56931]_ , \new_[56932]_ , \new_[56935]_ , \new_[56938]_ ,
    \new_[56939]_ , \new_[56940]_ , \new_[56943]_ , \new_[56946]_ ,
    \new_[56947]_ , \new_[56950]_ , \new_[56953]_ , \new_[56954]_ ,
    \new_[56955]_ , \new_[56958]_ , \new_[56961]_ , \new_[56962]_ ,
    \new_[56965]_ , \new_[56968]_ , \new_[56969]_ , \new_[56970]_ ,
    \new_[56973]_ , \new_[56976]_ , \new_[56977]_ , \new_[56980]_ ,
    \new_[56983]_ , \new_[56984]_ , \new_[56985]_ , \new_[56988]_ ,
    \new_[56991]_ , \new_[56992]_ , \new_[56995]_ , \new_[56998]_ ,
    \new_[56999]_ , \new_[57000]_ , \new_[57003]_ , \new_[57006]_ ,
    \new_[57007]_ , \new_[57010]_ , \new_[57013]_ , \new_[57014]_ ,
    \new_[57015]_ , \new_[57018]_ , \new_[57021]_ , \new_[57022]_ ,
    \new_[57025]_ , \new_[57028]_ , \new_[57029]_ , \new_[57030]_ ,
    \new_[57033]_ , \new_[57036]_ , \new_[57037]_ , \new_[57040]_ ,
    \new_[57043]_ , \new_[57044]_ , \new_[57045]_ , \new_[57048]_ ,
    \new_[57051]_ , \new_[57052]_ , \new_[57055]_ , \new_[57058]_ ,
    \new_[57059]_ , \new_[57060]_ , \new_[57063]_ , \new_[57066]_ ,
    \new_[57067]_ , \new_[57070]_ , \new_[57073]_ , \new_[57074]_ ,
    \new_[57075]_ , \new_[57078]_ , \new_[57081]_ , \new_[57082]_ ,
    \new_[57085]_ , \new_[57088]_ , \new_[57089]_ , \new_[57090]_ ,
    \new_[57093]_ , \new_[57096]_ , \new_[57097]_ , \new_[57100]_ ,
    \new_[57103]_ , \new_[57104]_ , \new_[57105]_ , \new_[57108]_ ,
    \new_[57111]_ , \new_[57112]_ , \new_[57115]_ , \new_[57118]_ ,
    \new_[57119]_ , \new_[57120]_ , \new_[57123]_ , \new_[57126]_ ,
    \new_[57127]_ , \new_[57130]_ , \new_[57133]_ , \new_[57134]_ ,
    \new_[57135]_ , \new_[57138]_ , \new_[57141]_ , \new_[57142]_ ,
    \new_[57145]_ , \new_[57148]_ , \new_[57149]_ , \new_[57150]_ ,
    \new_[57153]_ , \new_[57156]_ , \new_[57157]_ , \new_[57160]_ ,
    \new_[57163]_ , \new_[57164]_ , \new_[57165]_ , \new_[57168]_ ,
    \new_[57171]_ , \new_[57172]_ , \new_[57175]_ , \new_[57178]_ ,
    \new_[57179]_ , \new_[57180]_ , \new_[57183]_ , \new_[57186]_ ,
    \new_[57187]_ , \new_[57190]_ , \new_[57193]_ , \new_[57194]_ ,
    \new_[57195]_ , \new_[57198]_ , \new_[57201]_ , \new_[57202]_ ,
    \new_[57205]_ , \new_[57208]_ , \new_[57209]_ , \new_[57210]_ ,
    \new_[57213]_ , \new_[57216]_ , \new_[57217]_ , \new_[57220]_ ,
    \new_[57223]_ , \new_[57224]_ , \new_[57225]_ , \new_[57228]_ ,
    \new_[57231]_ , \new_[57232]_ , \new_[57235]_ , \new_[57238]_ ,
    \new_[57239]_ , \new_[57240]_ , \new_[57243]_ , \new_[57246]_ ,
    \new_[57247]_ , \new_[57250]_ , \new_[57253]_ , \new_[57254]_ ,
    \new_[57255]_ , \new_[57258]_ , \new_[57261]_ , \new_[57262]_ ,
    \new_[57265]_ , \new_[57268]_ , \new_[57269]_ , \new_[57270]_ ,
    \new_[57273]_ , \new_[57276]_ , \new_[57277]_ , \new_[57280]_ ,
    \new_[57283]_ , \new_[57284]_ , \new_[57285]_ , \new_[57288]_ ,
    \new_[57291]_ , \new_[57292]_ , \new_[57295]_ , \new_[57298]_ ,
    \new_[57299]_ , \new_[57300]_ , \new_[57303]_ , \new_[57306]_ ,
    \new_[57307]_ , \new_[57310]_ , \new_[57313]_ , \new_[57314]_ ,
    \new_[57315]_ , \new_[57318]_ , \new_[57321]_ , \new_[57322]_ ,
    \new_[57325]_ , \new_[57328]_ , \new_[57329]_ , \new_[57330]_ ,
    \new_[57333]_ , \new_[57336]_ , \new_[57337]_ , \new_[57340]_ ,
    \new_[57343]_ , \new_[57344]_ , \new_[57345]_ , \new_[57348]_ ,
    \new_[57351]_ , \new_[57352]_ , \new_[57355]_ , \new_[57358]_ ,
    \new_[57359]_ , \new_[57360]_ , \new_[57363]_ , \new_[57366]_ ,
    \new_[57367]_ , \new_[57370]_ , \new_[57373]_ , \new_[57374]_ ,
    \new_[57375]_ , \new_[57378]_ , \new_[57381]_ , \new_[57382]_ ,
    \new_[57385]_ , \new_[57388]_ , \new_[57389]_ , \new_[57390]_ ,
    \new_[57393]_ , \new_[57396]_ , \new_[57397]_ , \new_[57400]_ ,
    \new_[57403]_ , \new_[57404]_ , \new_[57405]_ , \new_[57408]_ ,
    \new_[57411]_ , \new_[57412]_ , \new_[57415]_ , \new_[57418]_ ,
    \new_[57419]_ , \new_[57420]_ , \new_[57423]_ , \new_[57426]_ ,
    \new_[57427]_ , \new_[57430]_ , \new_[57433]_ , \new_[57434]_ ,
    \new_[57435]_ , \new_[57438]_ , \new_[57441]_ , \new_[57442]_ ,
    \new_[57445]_ , \new_[57448]_ , \new_[57449]_ , \new_[57450]_ ,
    \new_[57453]_ , \new_[57456]_ , \new_[57457]_ , \new_[57460]_ ,
    \new_[57463]_ , \new_[57464]_ , \new_[57465]_ , \new_[57468]_ ,
    \new_[57471]_ , \new_[57472]_ , \new_[57475]_ , \new_[57478]_ ,
    \new_[57479]_ , \new_[57480]_ , \new_[57483]_ , \new_[57486]_ ,
    \new_[57487]_ , \new_[57490]_ , \new_[57493]_ , \new_[57494]_ ,
    \new_[57495]_ , \new_[57498]_ , \new_[57501]_ , \new_[57502]_ ,
    \new_[57505]_ , \new_[57508]_ , \new_[57509]_ , \new_[57510]_ ,
    \new_[57513]_ , \new_[57516]_ , \new_[57517]_ , \new_[57520]_ ,
    \new_[57523]_ , \new_[57524]_ , \new_[57525]_ , \new_[57528]_ ,
    \new_[57531]_ , \new_[57532]_ , \new_[57535]_ , \new_[57538]_ ,
    \new_[57539]_ , \new_[57540]_ , \new_[57543]_ , \new_[57546]_ ,
    \new_[57547]_ , \new_[57550]_ , \new_[57553]_ , \new_[57554]_ ,
    \new_[57555]_ , \new_[57558]_ , \new_[57561]_ , \new_[57562]_ ,
    \new_[57565]_ , \new_[57568]_ , \new_[57569]_ , \new_[57570]_ ,
    \new_[57573]_ , \new_[57576]_ , \new_[57577]_ , \new_[57580]_ ,
    \new_[57583]_ , \new_[57584]_ , \new_[57585]_ , \new_[57588]_ ,
    \new_[57591]_ , \new_[57592]_ , \new_[57595]_ , \new_[57598]_ ,
    \new_[57599]_ , \new_[57600]_ , \new_[57603]_ , \new_[57606]_ ,
    \new_[57607]_ , \new_[57610]_ , \new_[57613]_ , \new_[57614]_ ,
    \new_[57615]_ , \new_[57618]_ , \new_[57621]_ , \new_[57622]_ ,
    \new_[57625]_ , \new_[57628]_ , \new_[57629]_ , \new_[57630]_ ,
    \new_[57633]_ , \new_[57636]_ , \new_[57637]_ , \new_[57640]_ ,
    \new_[57643]_ , \new_[57644]_ , \new_[57645]_ , \new_[57648]_ ,
    \new_[57651]_ , \new_[57652]_ , \new_[57655]_ , \new_[57658]_ ,
    \new_[57659]_ , \new_[57660]_ , \new_[57663]_ , \new_[57666]_ ,
    \new_[57667]_ , \new_[57670]_ , \new_[57673]_ , \new_[57674]_ ,
    \new_[57675]_ , \new_[57678]_ , \new_[57681]_ , \new_[57682]_ ,
    \new_[57685]_ , \new_[57688]_ , \new_[57689]_ , \new_[57690]_ ,
    \new_[57693]_ , \new_[57696]_ , \new_[57697]_ , \new_[57700]_ ,
    \new_[57703]_ , \new_[57704]_ , \new_[57705]_ , \new_[57708]_ ,
    \new_[57711]_ , \new_[57712]_ , \new_[57715]_ , \new_[57718]_ ,
    \new_[57719]_ , \new_[57720]_ , \new_[57723]_ , \new_[57726]_ ,
    \new_[57727]_ , \new_[57730]_ , \new_[57733]_ , \new_[57734]_ ,
    \new_[57735]_ , \new_[57738]_ , \new_[57741]_ , \new_[57742]_ ,
    \new_[57745]_ , \new_[57748]_ , \new_[57749]_ , \new_[57750]_ ,
    \new_[57753]_ , \new_[57756]_ , \new_[57757]_ , \new_[57760]_ ,
    \new_[57763]_ , \new_[57764]_ , \new_[57765]_ , \new_[57768]_ ,
    \new_[57771]_ , \new_[57772]_ , \new_[57775]_ , \new_[57778]_ ,
    \new_[57779]_ , \new_[57780]_ , \new_[57783]_ , \new_[57786]_ ,
    \new_[57787]_ , \new_[57790]_ , \new_[57793]_ , \new_[57794]_ ,
    \new_[57795]_ , \new_[57798]_ , \new_[57801]_ , \new_[57802]_ ,
    \new_[57805]_ , \new_[57808]_ , \new_[57809]_ , \new_[57810]_ ,
    \new_[57813]_ , \new_[57816]_ , \new_[57817]_ , \new_[57820]_ ,
    \new_[57823]_ , \new_[57824]_ , \new_[57825]_ , \new_[57828]_ ,
    \new_[57831]_ , \new_[57832]_ , \new_[57835]_ , \new_[57838]_ ,
    \new_[57839]_ , \new_[57840]_ , \new_[57843]_ , \new_[57846]_ ,
    \new_[57847]_ , \new_[57850]_ , \new_[57853]_ , \new_[57854]_ ,
    \new_[57855]_ , \new_[57858]_ , \new_[57861]_ , \new_[57862]_ ,
    \new_[57865]_ , \new_[57868]_ , \new_[57869]_ , \new_[57870]_ ,
    \new_[57873]_ , \new_[57876]_ , \new_[57877]_ , \new_[57880]_ ,
    \new_[57883]_ , \new_[57884]_ , \new_[57885]_ , \new_[57888]_ ,
    \new_[57891]_ , \new_[57892]_ , \new_[57895]_ , \new_[57898]_ ,
    \new_[57899]_ , \new_[57900]_ , \new_[57903]_ , \new_[57906]_ ,
    \new_[57907]_ , \new_[57910]_ , \new_[57913]_ , \new_[57914]_ ,
    \new_[57915]_ , \new_[57918]_ , \new_[57921]_ , \new_[57922]_ ,
    \new_[57925]_ , \new_[57928]_ , \new_[57929]_ , \new_[57930]_ ,
    \new_[57933]_ , \new_[57936]_ , \new_[57937]_ , \new_[57940]_ ,
    \new_[57943]_ , \new_[57944]_ , \new_[57945]_ , \new_[57948]_ ,
    \new_[57951]_ , \new_[57952]_ , \new_[57955]_ , \new_[57958]_ ,
    \new_[57959]_ , \new_[57960]_ , \new_[57963]_ , \new_[57966]_ ,
    \new_[57967]_ , \new_[57970]_ , \new_[57973]_ , \new_[57974]_ ,
    \new_[57975]_ , \new_[57978]_ , \new_[57981]_ , \new_[57982]_ ,
    \new_[57985]_ , \new_[57988]_ , \new_[57989]_ , \new_[57990]_ ,
    \new_[57993]_ , \new_[57996]_ , \new_[57997]_ , \new_[58000]_ ,
    \new_[58003]_ , \new_[58004]_ , \new_[58005]_ , \new_[58008]_ ,
    \new_[58011]_ , \new_[58012]_ , \new_[58015]_ , \new_[58018]_ ,
    \new_[58019]_ , \new_[58020]_ , \new_[58023]_ , \new_[58026]_ ,
    \new_[58027]_ , \new_[58030]_ , \new_[58033]_ , \new_[58034]_ ,
    \new_[58035]_ , \new_[58038]_ , \new_[58041]_ , \new_[58042]_ ,
    \new_[58045]_ , \new_[58048]_ , \new_[58049]_ , \new_[58050]_ ,
    \new_[58053]_ , \new_[58056]_ , \new_[58057]_ , \new_[58060]_ ,
    \new_[58063]_ , \new_[58064]_ , \new_[58065]_ , \new_[58068]_ ,
    \new_[58071]_ , \new_[58072]_ , \new_[58075]_ , \new_[58078]_ ,
    \new_[58079]_ , \new_[58080]_ , \new_[58083]_ , \new_[58086]_ ,
    \new_[58087]_ , \new_[58090]_ , \new_[58093]_ , \new_[58094]_ ,
    \new_[58095]_ , \new_[58098]_ , \new_[58101]_ , \new_[58102]_ ,
    \new_[58105]_ , \new_[58108]_ , \new_[58109]_ , \new_[58110]_ ,
    \new_[58113]_ , \new_[58116]_ , \new_[58117]_ , \new_[58120]_ ,
    \new_[58123]_ , \new_[58124]_ , \new_[58125]_ , \new_[58128]_ ,
    \new_[58131]_ , \new_[58132]_ , \new_[58135]_ , \new_[58138]_ ,
    \new_[58139]_ , \new_[58140]_ , \new_[58143]_ , \new_[58146]_ ,
    \new_[58147]_ , \new_[58150]_ , \new_[58153]_ , \new_[58154]_ ,
    \new_[58155]_ , \new_[58158]_ , \new_[58161]_ , \new_[58162]_ ,
    \new_[58165]_ , \new_[58168]_ , \new_[58169]_ , \new_[58170]_ ,
    \new_[58173]_ , \new_[58176]_ , \new_[58177]_ , \new_[58180]_ ,
    \new_[58183]_ , \new_[58184]_ , \new_[58185]_ , \new_[58188]_ ,
    \new_[58191]_ , \new_[58192]_ , \new_[58195]_ , \new_[58198]_ ,
    \new_[58199]_ , \new_[58200]_ , \new_[58203]_ , \new_[58206]_ ,
    \new_[58207]_ , \new_[58210]_ , \new_[58213]_ , \new_[58214]_ ,
    \new_[58215]_ , \new_[58218]_ , \new_[58221]_ , \new_[58222]_ ,
    \new_[58225]_ , \new_[58228]_ , \new_[58229]_ , \new_[58230]_ ,
    \new_[58233]_ , \new_[58236]_ , \new_[58237]_ , \new_[58240]_ ,
    \new_[58243]_ , \new_[58244]_ , \new_[58245]_ , \new_[58248]_ ,
    \new_[58251]_ , \new_[58252]_ , \new_[58255]_ , \new_[58258]_ ,
    \new_[58259]_ , \new_[58260]_ , \new_[58263]_ , \new_[58266]_ ,
    \new_[58267]_ , \new_[58270]_ , \new_[58273]_ , \new_[58274]_ ,
    \new_[58275]_ , \new_[58278]_ , \new_[58281]_ , \new_[58282]_ ,
    \new_[58285]_ , \new_[58288]_ , \new_[58289]_ , \new_[58290]_ ,
    \new_[58293]_ , \new_[58296]_ , \new_[58297]_ , \new_[58300]_ ,
    \new_[58303]_ , \new_[58304]_ , \new_[58305]_ , \new_[58308]_ ,
    \new_[58311]_ , \new_[58312]_ , \new_[58315]_ , \new_[58318]_ ,
    \new_[58319]_ , \new_[58320]_ , \new_[58323]_ , \new_[58326]_ ,
    \new_[58327]_ , \new_[58330]_ , \new_[58333]_ , \new_[58334]_ ,
    \new_[58335]_ , \new_[58338]_ , \new_[58341]_ , \new_[58342]_ ,
    \new_[58345]_ , \new_[58348]_ , \new_[58349]_ , \new_[58350]_ ,
    \new_[58353]_ , \new_[58356]_ , \new_[58357]_ , \new_[58360]_ ,
    \new_[58363]_ , \new_[58364]_ , \new_[58365]_ , \new_[58368]_ ,
    \new_[58371]_ , \new_[58372]_ , \new_[58375]_ , \new_[58378]_ ,
    \new_[58379]_ , \new_[58380]_ , \new_[58383]_ , \new_[58386]_ ,
    \new_[58387]_ , \new_[58390]_ , \new_[58393]_ , \new_[58394]_ ,
    \new_[58395]_ , \new_[58398]_ , \new_[58401]_ , \new_[58402]_ ,
    \new_[58405]_ , \new_[58408]_ , \new_[58409]_ , \new_[58410]_ ,
    \new_[58413]_ , \new_[58416]_ , \new_[58417]_ , \new_[58420]_ ,
    \new_[58423]_ , \new_[58424]_ , \new_[58425]_ , \new_[58428]_ ,
    \new_[58431]_ , \new_[58432]_ , \new_[58435]_ , \new_[58438]_ ,
    \new_[58439]_ , \new_[58440]_ , \new_[58443]_ , \new_[58446]_ ,
    \new_[58447]_ , \new_[58450]_ , \new_[58453]_ , \new_[58454]_ ,
    \new_[58455]_ , \new_[58458]_ , \new_[58461]_ , \new_[58462]_ ,
    \new_[58465]_ , \new_[58468]_ , \new_[58469]_ , \new_[58470]_ ,
    \new_[58473]_ , \new_[58476]_ , \new_[58477]_ , \new_[58480]_ ,
    \new_[58483]_ , \new_[58484]_ , \new_[58485]_ , \new_[58488]_ ,
    \new_[58491]_ , \new_[58492]_ , \new_[58495]_ , \new_[58498]_ ,
    \new_[58499]_ , \new_[58500]_ , \new_[58503]_ , \new_[58506]_ ,
    \new_[58507]_ , \new_[58510]_ , \new_[58513]_ , \new_[58514]_ ,
    \new_[58515]_ , \new_[58518]_ , \new_[58521]_ , \new_[58522]_ ,
    \new_[58525]_ , \new_[58528]_ , \new_[58529]_ , \new_[58530]_ ,
    \new_[58533]_ , \new_[58536]_ , \new_[58537]_ , \new_[58540]_ ,
    \new_[58543]_ , \new_[58544]_ , \new_[58545]_ , \new_[58548]_ ,
    \new_[58551]_ , \new_[58552]_ , \new_[58555]_ , \new_[58558]_ ,
    \new_[58559]_ , \new_[58560]_ , \new_[58563]_ , \new_[58566]_ ,
    \new_[58567]_ , \new_[58570]_ , \new_[58573]_ , \new_[58574]_ ,
    \new_[58575]_ , \new_[58578]_ , \new_[58581]_ , \new_[58582]_ ,
    \new_[58585]_ , \new_[58588]_ , \new_[58589]_ , \new_[58590]_ ,
    \new_[58593]_ , \new_[58596]_ , \new_[58597]_ , \new_[58600]_ ,
    \new_[58603]_ , \new_[58604]_ , \new_[58605]_ , \new_[58608]_ ,
    \new_[58611]_ , \new_[58612]_ , \new_[58615]_ , \new_[58618]_ ,
    \new_[58619]_ , \new_[58620]_ , \new_[58623]_ , \new_[58626]_ ,
    \new_[58627]_ , \new_[58630]_ , \new_[58633]_ , \new_[58634]_ ,
    \new_[58635]_ , \new_[58638]_ , \new_[58641]_ , \new_[58642]_ ,
    \new_[58645]_ , \new_[58648]_ , \new_[58649]_ , \new_[58650]_ ,
    \new_[58653]_ , \new_[58656]_ , \new_[58657]_ , \new_[58660]_ ,
    \new_[58663]_ , \new_[58664]_ , \new_[58665]_ , \new_[58668]_ ,
    \new_[58671]_ , \new_[58672]_ , \new_[58675]_ , \new_[58678]_ ,
    \new_[58679]_ , \new_[58680]_ , \new_[58683]_ , \new_[58686]_ ,
    \new_[58687]_ , \new_[58690]_ , \new_[58693]_ , \new_[58694]_ ,
    \new_[58695]_ , \new_[58698]_ , \new_[58701]_ , \new_[58702]_ ,
    \new_[58705]_ , \new_[58708]_ , \new_[58709]_ , \new_[58710]_ ,
    \new_[58713]_ , \new_[58716]_ , \new_[58717]_ , \new_[58720]_ ,
    \new_[58723]_ , \new_[58724]_ , \new_[58725]_ , \new_[58728]_ ,
    \new_[58731]_ , \new_[58732]_ , \new_[58735]_ , \new_[58738]_ ,
    \new_[58739]_ , \new_[58740]_ , \new_[58743]_ , \new_[58746]_ ,
    \new_[58747]_ , \new_[58750]_ , \new_[58753]_ , \new_[58754]_ ,
    \new_[58755]_ , \new_[58758]_ , \new_[58761]_ , \new_[58762]_ ,
    \new_[58765]_ , \new_[58768]_ , \new_[58769]_ , \new_[58770]_ ,
    \new_[58773]_ , \new_[58776]_ , \new_[58777]_ , \new_[58780]_ ,
    \new_[58783]_ , \new_[58784]_ , \new_[58785]_ , \new_[58788]_ ,
    \new_[58791]_ , \new_[58792]_ , \new_[58795]_ , \new_[58798]_ ,
    \new_[58799]_ , \new_[58800]_ , \new_[58803]_ , \new_[58806]_ ,
    \new_[58807]_ , \new_[58810]_ , \new_[58813]_ , \new_[58814]_ ,
    \new_[58815]_ , \new_[58818]_ , \new_[58821]_ , \new_[58822]_ ,
    \new_[58825]_ , \new_[58828]_ , \new_[58829]_ , \new_[58830]_ ,
    \new_[58833]_ , \new_[58836]_ , \new_[58837]_ , \new_[58840]_ ,
    \new_[58843]_ , \new_[58844]_ , \new_[58845]_ , \new_[58848]_ ,
    \new_[58851]_ , \new_[58852]_ , \new_[58855]_ , \new_[58858]_ ,
    \new_[58859]_ , \new_[58860]_ , \new_[58863]_ , \new_[58866]_ ,
    \new_[58867]_ , \new_[58870]_ , \new_[58873]_ , \new_[58874]_ ,
    \new_[58875]_ , \new_[58878]_ , \new_[58881]_ , \new_[58882]_ ,
    \new_[58885]_ , \new_[58888]_ , \new_[58889]_ , \new_[58890]_ ,
    \new_[58893]_ , \new_[58896]_ , \new_[58897]_ , \new_[58900]_ ,
    \new_[58903]_ , \new_[58904]_ , \new_[58905]_ , \new_[58908]_ ,
    \new_[58911]_ , \new_[58912]_ , \new_[58915]_ , \new_[58918]_ ,
    \new_[58919]_ , \new_[58920]_ , \new_[58923]_ , \new_[58926]_ ,
    \new_[58927]_ , \new_[58930]_ , \new_[58933]_ , \new_[58934]_ ,
    \new_[58935]_ , \new_[58938]_ , \new_[58941]_ , \new_[58942]_ ,
    \new_[58945]_ , \new_[58948]_ , \new_[58949]_ , \new_[58950]_ ,
    \new_[58953]_ , \new_[58956]_ , \new_[58957]_ , \new_[58960]_ ,
    \new_[58963]_ , \new_[58964]_ , \new_[58965]_ , \new_[58968]_ ,
    \new_[58971]_ , \new_[58972]_ , \new_[58975]_ , \new_[58978]_ ,
    \new_[58979]_ , \new_[58980]_ , \new_[58983]_ , \new_[58986]_ ,
    \new_[58987]_ , \new_[58990]_ , \new_[58993]_ , \new_[58994]_ ,
    \new_[58995]_ , \new_[58998]_ , \new_[59001]_ , \new_[59002]_ ,
    \new_[59005]_ , \new_[59008]_ , \new_[59009]_ , \new_[59010]_ ,
    \new_[59013]_ , \new_[59016]_ , \new_[59017]_ , \new_[59020]_ ,
    \new_[59023]_ , \new_[59024]_ , \new_[59025]_ , \new_[59028]_ ,
    \new_[59031]_ , \new_[59032]_ , \new_[59035]_ , \new_[59038]_ ,
    \new_[59039]_ , \new_[59040]_ , \new_[59043]_ , \new_[59046]_ ,
    \new_[59047]_ , \new_[59050]_ , \new_[59053]_ , \new_[59054]_ ,
    \new_[59055]_ , \new_[59058]_ , \new_[59061]_ , \new_[59062]_ ,
    \new_[59065]_ , \new_[59068]_ , \new_[59069]_ , \new_[59070]_ ,
    \new_[59073]_ , \new_[59076]_ , \new_[59077]_ , \new_[59080]_ ,
    \new_[59083]_ , \new_[59084]_ , \new_[59085]_ , \new_[59088]_ ,
    \new_[59091]_ , \new_[59092]_ , \new_[59095]_ , \new_[59098]_ ,
    \new_[59099]_ , \new_[59100]_ , \new_[59103]_ , \new_[59106]_ ,
    \new_[59107]_ , \new_[59110]_ , \new_[59113]_ , \new_[59114]_ ,
    \new_[59115]_ , \new_[59118]_ , \new_[59121]_ , \new_[59122]_ ,
    \new_[59125]_ , \new_[59128]_ , \new_[59129]_ , \new_[59130]_ ,
    \new_[59133]_ , \new_[59136]_ , \new_[59137]_ , \new_[59140]_ ,
    \new_[59143]_ , \new_[59144]_ , \new_[59145]_ , \new_[59148]_ ,
    \new_[59151]_ , \new_[59152]_ , \new_[59155]_ , \new_[59158]_ ,
    \new_[59159]_ , \new_[59160]_ , \new_[59163]_ , \new_[59166]_ ,
    \new_[59167]_ , \new_[59170]_ , \new_[59173]_ , \new_[59174]_ ,
    \new_[59175]_ , \new_[59178]_ , \new_[59181]_ , \new_[59182]_ ,
    \new_[59185]_ , \new_[59188]_ , \new_[59189]_ , \new_[59190]_ ,
    \new_[59193]_ , \new_[59196]_ , \new_[59197]_ , \new_[59200]_ ,
    \new_[59203]_ , \new_[59204]_ , \new_[59205]_ , \new_[59208]_ ,
    \new_[59211]_ , \new_[59212]_ , \new_[59215]_ , \new_[59218]_ ,
    \new_[59219]_ , \new_[59220]_ , \new_[59223]_ , \new_[59226]_ ,
    \new_[59227]_ , \new_[59230]_ , \new_[59233]_ , \new_[59234]_ ,
    \new_[59235]_ , \new_[59238]_ , \new_[59241]_ , \new_[59242]_ ,
    \new_[59245]_ , \new_[59248]_ , \new_[59249]_ , \new_[59250]_ ,
    \new_[59253]_ , \new_[59256]_ , \new_[59257]_ , \new_[59260]_ ,
    \new_[59263]_ , \new_[59264]_ , \new_[59265]_ , \new_[59268]_ ,
    \new_[59271]_ , \new_[59272]_ , \new_[59275]_ , \new_[59278]_ ,
    \new_[59279]_ , \new_[59280]_ , \new_[59283]_ , \new_[59286]_ ,
    \new_[59287]_ , \new_[59290]_ , \new_[59293]_ , \new_[59294]_ ,
    \new_[59295]_ , \new_[59298]_ , \new_[59301]_ , \new_[59302]_ ,
    \new_[59305]_ , \new_[59308]_ , \new_[59309]_ , \new_[59310]_ ,
    \new_[59313]_ , \new_[59316]_ , \new_[59317]_ , \new_[59320]_ ,
    \new_[59323]_ , \new_[59324]_ , \new_[59325]_ , \new_[59328]_ ,
    \new_[59331]_ , \new_[59332]_ , \new_[59335]_ , \new_[59338]_ ,
    \new_[59339]_ , \new_[59340]_ , \new_[59343]_ , \new_[59346]_ ,
    \new_[59347]_ , \new_[59350]_ , \new_[59353]_ , \new_[59354]_ ,
    \new_[59355]_ , \new_[59358]_ , \new_[59361]_ , \new_[59362]_ ,
    \new_[59365]_ , \new_[59368]_ , \new_[59369]_ , \new_[59370]_ ,
    \new_[59373]_ , \new_[59376]_ , \new_[59377]_ , \new_[59380]_ ,
    \new_[59383]_ , \new_[59384]_ , \new_[59385]_ , \new_[59388]_ ,
    \new_[59391]_ , \new_[59392]_ , \new_[59395]_ , \new_[59398]_ ,
    \new_[59399]_ , \new_[59400]_ , \new_[59403]_ , \new_[59406]_ ,
    \new_[59407]_ , \new_[59410]_ , \new_[59413]_ , \new_[59414]_ ,
    \new_[59415]_ , \new_[59418]_ , \new_[59421]_ , \new_[59422]_ ,
    \new_[59425]_ , \new_[59428]_ , \new_[59429]_ , \new_[59430]_ ,
    \new_[59433]_ , \new_[59436]_ , \new_[59437]_ , \new_[59440]_ ,
    \new_[59443]_ , \new_[59444]_ , \new_[59445]_ , \new_[59448]_ ,
    \new_[59451]_ , \new_[59452]_ , \new_[59455]_ , \new_[59458]_ ,
    \new_[59459]_ , \new_[59460]_ , \new_[59463]_ , \new_[59466]_ ,
    \new_[59467]_ , \new_[59470]_ , \new_[59473]_ , \new_[59474]_ ,
    \new_[59475]_ , \new_[59478]_ , \new_[59481]_ , \new_[59482]_ ,
    \new_[59485]_ , \new_[59488]_ , \new_[59489]_ , \new_[59490]_ ,
    \new_[59493]_ , \new_[59496]_ , \new_[59497]_ , \new_[59500]_ ,
    \new_[59503]_ , \new_[59504]_ , \new_[59505]_ , \new_[59508]_ ,
    \new_[59511]_ , \new_[59512]_ , \new_[59515]_ , \new_[59518]_ ,
    \new_[59519]_ , \new_[59520]_ , \new_[59523]_ , \new_[59526]_ ,
    \new_[59527]_ , \new_[59530]_ , \new_[59533]_ , \new_[59534]_ ,
    \new_[59535]_ , \new_[59538]_ , \new_[59541]_ , \new_[59542]_ ,
    \new_[59545]_ , \new_[59548]_ , \new_[59549]_ , \new_[59550]_ ,
    \new_[59553]_ , \new_[59556]_ , \new_[59557]_ , \new_[59560]_ ,
    \new_[59563]_ , \new_[59564]_ , \new_[59565]_ , \new_[59568]_ ,
    \new_[59571]_ , \new_[59572]_ , \new_[59575]_ , \new_[59578]_ ,
    \new_[59579]_ , \new_[59580]_ , \new_[59583]_ , \new_[59586]_ ,
    \new_[59587]_ , \new_[59590]_ , \new_[59593]_ , \new_[59594]_ ,
    \new_[59595]_ , \new_[59598]_ , \new_[59601]_ , \new_[59602]_ ,
    \new_[59605]_ , \new_[59608]_ , \new_[59609]_ , \new_[59610]_ ,
    \new_[59613]_ , \new_[59616]_ , \new_[59617]_ , \new_[59620]_ ,
    \new_[59623]_ , \new_[59624]_ , \new_[59625]_ , \new_[59628]_ ,
    \new_[59631]_ , \new_[59632]_ , \new_[59635]_ , \new_[59638]_ ,
    \new_[59639]_ , \new_[59640]_ , \new_[59643]_ , \new_[59646]_ ,
    \new_[59647]_ , \new_[59650]_ , \new_[59653]_ , \new_[59654]_ ,
    \new_[59655]_ , \new_[59658]_ , \new_[59661]_ , \new_[59662]_ ,
    \new_[59665]_ , \new_[59668]_ , \new_[59669]_ , \new_[59670]_ ,
    \new_[59673]_ , \new_[59676]_ , \new_[59677]_ , \new_[59680]_ ,
    \new_[59683]_ , \new_[59684]_ , \new_[59685]_ , \new_[59688]_ ,
    \new_[59691]_ , \new_[59692]_ , \new_[59695]_ , \new_[59698]_ ,
    \new_[59699]_ , \new_[59700]_ , \new_[59703]_ , \new_[59706]_ ,
    \new_[59707]_ , \new_[59710]_ , \new_[59713]_ , \new_[59714]_ ,
    \new_[59715]_ , \new_[59718]_ , \new_[59721]_ , \new_[59722]_ ,
    \new_[59725]_ , \new_[59728]_ , \new_[59729]_ , \new_[59730]_ ,
    \new_[59733]_ , \new_[59736]_ , \new_[59737]_ , \new_[59740]_ ,
    \new_[59743]_ , \new_[59744]_ , \new_[59745]_ , \new_[59748]_ ,
    \new_[59751]_ , \new_[59752]_ , \new_[59755]_ , \new_[59758]_ ,
    \new_[59759]_ , \new_[59760]_ , \new_[59763]_ , \new_[59766]_ ,
    \new_[59767]_ , \new_[59770]_ , \new_[59773]_ , \new_[59774]_ ,
    \new_[59775]_ , \new_[59778]_ , \new_[59781]_ , \new_[59782]_ ,
    \new_[59785]_ , \new_[59788]_ , \new_[59789]_ , \new_[59790]_ ,
    \new_[59793]_ , \new_[59796]_ , \new_[59797]_ , \new_[59800]_ ,
    \new_[59803]_ , \new_[59804]_ , \new_[59805]_ , \new_[59808]_ ,
    \new_[59811]_ , \new_[59812]_ , \new_[59815]_ , \new_[59818]_ ,
    \new_[59819]_ , \new_[59820]_ , \new_[59823]_ , \new_[59826]_ ,
    \new_[59827]_ , \new_[59830]_ , \new_[59833]_ , \new_[59834]_ ,
    \new_[59835]_ , \new_[59838]_ , \new_[59841]_ , \new_[59842]_ ,
    \new_[59845]_ , \new_[59848]_ , \new_[59849]_ , \new_[59850]_ ,
    \new_[59853]_ , \new_[59856]_ , \new_[59857]_ , \new_[59860]_ ,
    \new_[59863]_ , \new_[59864]_ , \new_[59865]_ , \new_[59868]_ ,
    \new_[59871]_ , \new_[59872]_ , \new_[59875]_ , \new_[59878]_ ,
    \new_[59879]_ , \new_[59880]_ , \new_[59883]_ , \new_[59886]_ ,
    \new_[59887]_ , \new_[59890]_ , \new_[59893]_ , \new_[59894]_ ,
    \new_[59895]_ , \new_[59898]_ , \new_[59901]_ , \new_[59902]_ ,
    \new_[59905]_ , \new_[59908]_ , \new_[59909]_ , \new_[59910]_ ,
    \new_[59913]_ , \new_[59916]_ , \new_[59917]_ , \new_[59920]_ ,
    \new_[59923]_ , \new_[59924]_ , \new_[59925]_ , \new_[59928]_ ,
    \new_[59931]_ , \new_[59932]_ , \new_[59935]_ , \new_[59938]_ ,
    \new_[59939]_ , \new_[59940]_ , \new_[59943]_ , \new_[59946]_ ,
    \new_[59947]_ , \new_[59950]_ , \new_[59953]_ , \new_[59954]_ ,
    \new_[59955]_ , \new_[59958]_ , \new_[59961]_ , \new_[59962]_ ,
    \new_[59965]_ , \new_[59968]_ , \new_[59969]_ , \new_[59970]_ ,
    \new_[59973]_ , \new_[59976]_ , \new_[59977]_ , \new_[59980]_ ,
    \new_[59983]_ , \new_[59984]_ , \new_[59985]_ , \new_[59988]_ ,
    \new_[59991]_ , \new_[59992]_ , \new_[59995]_ , \new_[59998]_ ,
    \new_[59999]_ , \new_[60000]_ , \new_[60003]_ , \new_[60006]_ ,
    \new_[60007]_ , \new_[60010]_ , \new_[60013]_ , \new_[60014]_ ,
    \new_[60015]_ , \new_[60018]_ , \new_[60021]_ , \new_[60022]_ ,
    \new_[60025]_ , \new_[60028]_ , \new_[60029]_ , \new_[60030]_ ,
    \new_[60033]_ , \new_[60036]_ , \new_[60037]_ , \new_[60040]_ ,
    \new_[60043]_ , \new_[60044]_ , \new_[60045]_ , \new_[60048]_ ,
    \new_[60051]_ , \new_[60052]_ , \new_[60055]_ , \new_[60058]_ ,
    \new_[60059]_ , \new_[60060]_ , \new_[60063]_ , \new_[60066]_ ,
    \new_[60067]_ , \new_[60070]_ , \new_[60073]_ , \new_[60074]_ ,
    \new_[60075]_ , \new_[60078]_ , \new_[60081]_ , \new_[60082]_ ,
    \new_[60085]_ , \new_[60088]_ , \new_[60089]_ , \new_[60090]_ ,
    \new_[60093]_ , \new_[60096]_ , \new_[60097]_ , \new_[60100]_ ,
    \new_[60103]_ , \new_[60104]_ , \new_[60105]_ , \new_[60108]_ ,
    \new_[60111]_ , \new_[60112]_ , \new_[60115]_ , \new_[60118]_ ,
    \new_[60119]_ , \new_[60120]_ , \new_[60123]_ , \new_[60126]_ ,
    \new_[60127]_ , \new_[60130]_ , \new_[60133]_ , \new_[60134]_ ,
    \new_[60135]_ , \new_[60138]_ , \new_[60141]_ , \new_[60142]_ ,
    \new_[60145]_ , \new_[60148]_ , \new_[60149]_ , \new_[60150]_ ,
    \new_[60153]_ , \new_[60156]_ , \new_[60157]_ , \new_[60160]_ ,
    \new_[60163]_ , \new_[60164]_ , \new_[60165]_ , \new_[60168]_ ,
    \new_[60171]_ , \new_[60172]_ , \new_[60175]_ , \new_[60178]_ ,
    \new_[60179]_ , \new_[60180]_ , \new_[60183]_ , \new_[60186]_ ,
    \new_[60187]_ , \new_[60190]_ , \new_[60193]_ , \new_[60194]_ ,
    \new_[60195]_ , \new_[60198]_ , \new_[60201]_ , \new_[60202]_ ,
    \new_[60205]_ , \new_[60208]_ , \new_[60209]_ , \new_[60210]_ ,
    \new_[60213]_ , \new_[60216]_ , \new_[60217]_ , \new_[60220]_ ,
    \new_[60223]_ , \new_[60224]_ , \new_[60225]_ , \new_[60228]_ ,
    \new_[60231]_ , \new_[60232]_ , \new_[60235]_ , \new_[60238]_ ,
    \new_[60239]_ , \new_[60240]_ , \new_[60243]_ , \new_[60246]_ ,
    \new_[60247]_ , \new_[60250]_ , \new_[60253]_ , \new_[60254]_ ,
    \new_[60255]_ , \new_[60258]_ , \new_[60261]_ , \new_[60262]_ ,
    \new_[60265]_ , \new_[60268]_ , \new_[60269]_ , \new_[60270]_ ,
    \new_[60273]_ , \new_[60276]_ , \new_[60277]_ , \new_[60280]_ ,
    \new_[60283]_ , \new_[60284]_ , \new_[60285]_ , \new_[60288]_ ,
    \new_[60291]_ , \new_[60292]_ , \new_[60295]_ , \new_[60298]_ ,
    \new_[60299]_ , \new_[60300]_ , \new_[60303]_ , \new_[60306]_ ,
    \new_[60307]_ , \new_[60310]_ , \new_[60313]_ , \new_[60314]_ ,
    \new_[60315]_ , \new_[60318]_ , \new_[60321]_ , \new_[60322]_ ,
    \new_[60325]_ , \new_[60328]_ , \new_[60329]_ , \new_[60330]_ ,
    \new_[60333]_ , \new_[60336]_ , \new_[60337]_ , \new_[60340]_ ,
    \new_[60343]_ , \new_[60344]_ , \new_[60345]_ , \new_[60348]_ ,
    \new_[60351]_ , \new_[60352]_ , \new_[60355]_ , \new_[60358]_ ,
    \new_[60359]_ , \new_[60360]_ , \new_[60363]_ , \new_[60366]_ ,
    \new_[60367]_ , \new_[60370]_ , \new_[60373]_ , \new_[60374]_ ,
    \new_[60375]_ , \new_[60378]_ , \new_[60381]_ , \new_[60382]_ ,
    \new_[60385]_ , \new_[60388]_ , \new_[60389]_ , \new_[60390]_ ,
    \new_[60393]_ , \new_[60396]_ , \new_[60397]_ , \new_[60400]_ ,
    \new_[60403]_ , \new_[60404]_ , \new_[60405]_ , \new_[60408]_ ,
    \new_[60411]_ , \new_[60412]_ , \new_[60415]_ , \new_[60418]_ ,
    \new_[60419]_ , \new_[60420]_ , \new_[60423]_ , \new_[60426]_ ,
    \new_[60427]_ , \new_[60430]_ , \new_[60433]_ , \new_[60434]_ ,
    \new_[60435]_ , \new_[60438]_ , \new_[60441]_ , \new_[60442]_ ,
    \new_[60445]_ , \new_[60448]_ , \new_[60449]_ , \new_[60450]_ ,
    \new_[60453]_ , \new_[60456]_ , \new_[60457]_ , \new_[60460]_ ,
    \new_[60463]_ , \new_[60464]_ , \new_[60465]_ , \new_[60468]_ ,
    \new_[60471]_ , \new_[60472]_ , \new_[60475]_ , \new_[60478]_ ,
    \new_[60479]_ , \new_[60480]_ , \new_[60483]_ , \new_[60486]_ ,
    \new_[60487]_ , \new_[60490]_ , \new_[60493]_ , \new_[60494]_ ,
    \new_[60495]_ , \new_[60498]_ , \new_[60501]_ , \new_[60502]_ ,
    \new_[60505]_ , \new_[60508]_ , \new_[60509]_ , \new_[60510]_ ,
    \new_[60513]_ , \new_[60516]_ , \new_[60517]_ , \new_[60520]_ ,
    \new_[60523]_ , \new_[60524]_ , \new_[60525]_ , \new_[60528]_ ,
    \new_[60531]_ , \new_[60532]_ , \new_[60535]_ , \new_[60538]_ ,
    \new_[60539]_ , \new_[60540]_ , \new_[60543]_ , \new_[60546]_ ,
    \new_[60547]_ , \new_[60550]_ , \new_[60553]_ , \new_[60554]_ ,
    \new_[60555]_ , \new_[60558]_ , \new_[60561]_ , \new_[60562]_ ,
    \new_[60565]_ , \new_[60568]_ , \new_[60569]_ , \new_[60570]_ ,
    \new_[60573]_ , \new_[60576]_ , \new_[60577]_ , \new_[60580]_ ,
    \new_[60583]_ , \new_[60584]_ , \new_[60585]_ , \new_[60588]_ ,
    \new_[60591]_ , \new_[60592]_ , \new_[60595]_ , \new_[60598]_ ,
    \new_[60599]_ , \new_[60600]_ , \new_[60603]_ , \new_[60606]_ ,
    \new_[60607]_ , \new_[60610]_ , \new_[60613]_ , \new_[60614]_ ,
    \new_[60615]_ , \new_[60618]_ , \new_[60621]_ , \new_[60622]_ ,
    \new_[60625]_ , \new_[60628]_ , \new_[60629]_ , \new_[60630]_ ,
    \new_[60633]_ , \new_[60636]_ , \new_[60637]_ , \new_[60640]_ ,
    \new_[60643]_ , \new_[60644]_ , \new_[60645]_ , \new_[60648]_ ,
    \new_[60651]_ , \new_[60652]_ , \new_[60655]_ , \new_[60658]_ ,
    \new_[60659]_ , \new_[60660]_ , \new_[60663]_ , \new_[60666]_ ,
    \new_[60667]_ , \new_[60670]_ , \new_[60673]_ , \new_[60674]_ ,
    \new_[60675]_ , \new_[60678]_ , \new_[60681]_ , \new_[60682]_ ,
    \new_[60685]_ , \new_[60688]_ , \new_[60689]_ , \new_[60690]_ ,
    \new_[60693]_ , \new_[60696]_ , \new_[60697]_ , \new_[60700]_ ,
    \new_[60703]_ , \new_[60704]_ , \new_[60705]_ , \new_[60708]_ ,
    \new_[60711]_ , \new_[60712]_ , \new_[60715]_ , \new_[60718]_ ,
    \new_[60719]_ , \new_[60720]_ , \new_[60723]_ , \new_[60726]_ ,
    \new_[60727]_ , \new_[60730]_ , \new_[60733]_ , \new_[60734]_ ,
    \new_[60735]_ , \new_[60738]_ , \new_[60741]_ , \new_[60742]_ ,
    \new_[60745]_ , \new_[60748]_ , \new_[60749]_ , \new_[60750]_ ,
    \new_[60753]_ , \new_[60756]_ , \new_[60757]_ , \new_[60760]_ ,
    \new_[60763]_ , \new_[60764]_ , \new_[60765]_ , \new_[60768]_ ,
    \new_[60771]_ , \new_[60772]_ , \new_[60775]_ , \new_[60778]_ ,
    \new_[60779]_ , \new_[60780]_ , \new_[60783]_ , \new_[60786]_ ,
    \new_[60787]_ , \new_[60790]_ , \new_[60793]_ , \new_[60794]_ ,
    \new_[60795]_ , \new_[60798]_ , \new_[60801]_ , \new_[60802]_ ,
    \new_[60805]_ , \new_[60808]_ , \new_[60809]_ , \new_[60810]_ ,
    \new_[60813]_ , \new_[60816]_ , \new_[60817]_ , \new_[60820]_ ,
    \new_[60823]_ , \new_[60824]_ , \new_[60825]_ , \new_[60828]_ ,
    \new_[60831]_ , \new_[60832]_ , \new_[60835]_ , \new_[60838]_ ,
    \new_[60839]_ , \new_[60840]_ , \new_[60843]_ , \new_[60846]_ ,
    \new_[60847]_ , \new_[60850]_ , \new_[60853]_ , \new_[60854]_ ,
    \new_[60855]_ , \new_[60858]_ , \new_[60861]_ , \new_[60862]_ ,
    \new_[60865]_ , \new_[60868]_ , \new_[60869]_ , \new_[60870]_ ,
    \new_[60873]_ , \new_[60876]_ , \new_[60877]_ , \new_[60880]_ ,
    \new_[60883]_ , \new_[60884]_ , \new_[60885]_ , \new_[60888]_ ,
    \new_[60891]_ , \new_[60892]_ , \new_[60895]_ , \new_[60898]_ ,
    \new_[60899]_ , \new_[60900]_ , \new_[60903]_ , \new_[60906]_ ,
    \new_[60907]_ , \new_[60910]_ , \new_[60913]_ , \new_[60914]_ ,
    \new_[60915]_ , \new_[60918]_ , \new_[60921]_ , \new_[60922]_ ,
    \new_[60925]_ , \new_[60928]_ , \new_[60929]_ , \new_[60930]_ ,
    \new_[60933]_ , \new_[60936]_ , \new_[60937]_ , \new_[60940]_ ,
    \new_[60943]_ , \new_[60944]_ , \new_[60945]_ , \new_[60948]_ ,
    \new_[60951]_ , \new_[60952]_ , \new_[60955]_ , \new_[60958]_ ,
    \new_[60959]_ , \new_[60960]_ , \new_[60963]_ , \new_[60966]_ ,
    \new_[60967]_ , \new_[60970]_ , \new_[60973]_ , \new_[60974]_ ,
    \new_[60975]_ , \new_[60978]_ , \new_[60981]_ , \new_[60982]_ ,
    \new_[60985]_ , \new_[60988]_ , \new_[60989]_ , \new_[60990]_ ,
    \new_[60993]_ , \new_[60996]_ , \new_[60997]_ , \new_[61000]_ ,
    \new_[61003]_ , \new_[61004]_ , \new_[61005]_ , \new_[61008]_ ,
    \new_[61011]_ , \new_[61012]_ , \new_[61015]_ , \new_[61018]_ ,
    \new_[61019]_ , \new_[61020]_ , \new_[61023]_ , \new_[61026]_ ,
    \new_[61027]_ , \new_[61030]_ , \new_[61033]_ , \new_[61034]_ ,
    \new_[61035]_ , \new_[61038]_ , \new_[61041]_ , \new_[61042]_ ,
    \new_[61045]_ , \new_[61048]_ , \new_[61049]_ , \new_[61050]_ ,
    \new_[61053]_ , \new_[61056]_ , \new_[61057]_ , \new_[61060]_ ,
    \new_[61063]_ , \new_[61064]_ , \new_[61065]_ , \new_[61068]_ ,
    \new_[61071]_ , \new_[61072]_ , \new_[61075]_ , \new_[61078]_ ,
    \new_[61079]_ , \new_[61080]_ , \new_[61083]_ , \new_[61086]_ ,
    \new_[61087]_ , \new_[61090]_ , \new_[61093]_ , \new_[61094]_ ,
    \new_[61095]_ , \new_[61098]_ , \new_[61101]_ , \new_[61102]_ ,
    \new_[61105]_ , \new_[61108]_ , \new_[61109]_ , \new_[61110]_ ,
    \new_[61113]_ , \new_[61116]_ , \new_[61117]_ , \new_[61120]_ ,
    \new_[61123]_ , \new_[61124]_ , \new_[61125]_ , \new_[61128]_ ,
    \new_[61131]_ , \new_[61132]_ , \new_[61135]_ , \new_[61138]_ ,
    \new_[61139]_ , \new_[61140]_ , \new_[61143]_ , \new_[61146]_ ,
    \new_[61147]_ , \new_[61150]_ , \new_[61153]_ , \new_[61154]_ ,
    \new_[61155]_ , \new_[61158]_ , \new_[61161]_ , \new_[61162]_ ,
    \new_[61165]_ , \new_[61168]_ , \new_[61169]_ , \new_[61170]_ ,
    \new_[61173]_ , \new_[61176]_ , \new_[61177]_ , \new_[61180]_ ,
    \new_[61183]_ , \new_[61184]_ , \new_[61185]_ , \new_[61188]_ ,
    \new_[61191]_ , \new_[61192]_ , \new_[61195]_ , \new_[61198]_ ,
    \new_[61199]_ , \new_[61200]_ , \new_[61203]_ , \new_[61206]_ ,
    \new_[61207]_ , \new_[61210]_ , \new_[61213]_ , \new_[61214]_ ,
    \new_[61215]_ , \new_[61218]_ , \new_[61221]_ , \new_[61222]_ ,
    \new_[61225]_ , \new_[61228]_ , \new_[61229]_ , \new_[61230]_ ,
    \new_[61233]_ , \new_[61236]_ , \new_[61237]_ , \new_[61240]_ ,
    \new_[61243]_ , \new_[61244]_ , \new_[61245]_ , \new_[61248]_ ,
    \new_[61251]_ , \new_[61252]_ , \new_[61255]_ , \new_[61258]_ ,
    \new_[61259]_ , \new_[61260]_ , \new_[61263]_ , \new_[61266]_ ,
    \new_[61267]_ , \new_[61270]_ , \new_[61273]_ , \new_[61274]_ ,
    \new_[61275]_ , \new_[61278]_ , \new_[61281]_ , \new_[61282]_ ,
    \new_[61285]_ , \new_[61288]_ , \new_[61289]_ , \new_[61290]_ ,
    \new_[61293]_ , \new_[61296]_ , \new_[61297]_ , \new_[61300]_ ,
    \new_[61303]_ , \new_[61304]_ , \new_[61305]_ , \new_[61308]_ ,
    \new_[61311]_ , \new_[61312]_ , \new_[61315]_ , \new_[61318]_ ,
    \new_[61319]_ , \new_[61320]_ , \new_[61323]_ , \new_[61326]_ ,
    \new_[61327]_ , \new_[61330]_ , \new_[61333]_ , \new_[61334]_ ,
    \new_[61335]_ , \new_[61338]_ , \new_[61341]_ , \new_[61342]_ ,
    \new_[61345]_ , \new_[61348]_ , \new_[61349]_ , \new_[61350]_ ,
    \new_[61353]_ , \new_[61356]_ , \new_[61357]_ , \new_[61360]_ ,
    \new_[61363]_ , \new_[61364]_ , \new_[61365]_ , \new_[61368]_ ,
    \new_[61371]_ , \new_[61372]_ , \new_[61375]_ , \new_[61378]_ ,
    \new_[61379]_ , \new_[61380]_ , \new_[61383]_ , \new_[61386]_ ,
    \new_[61387]_ , \new_[61390]_ , \new_[61393]_ , \new_[61394]_ ,
    \new_[61395]_ , \new_[61398]_ , \new_[61401]_ , \new_[61402]_ ,
    \new_[61405]_ , \new_[61408]_ , \new_[61409]_ , \new_[61410]_ ,
    \new_[61413]_ , \new_[61416]_ , \new_[61417]_ , \new_[61420]_ ,
    \new_[61423]_ , \new_[61424]_ , \new_[61425]_ , \new_[61428]_ ,
    \new_[61431]_ , \new_[61432]_ , \new_[61435]_ , \new_[61438]_ ,
    \new_[61439]_ , \new_[61440]_ , \new_[61443]_ , \new_[61446]_ ,
    \new_[61447]_ , \new_[61450]_ , \new_[61453]_ , \new_[61454]_ ,
    \new_[61455]_ , \new_[61458]_ , \new_[61461]_ , \new_[61462]_ ,
    \new_[61465]_ , \new_[61468]_ , \new_[61469]_ , \new_[61470]_ ,
    \new_[61473]_ , \new_[61476]_ , \new_[61477]_ , \new_[61480]_ ,
    \new_[61483]_ , \new_[61484]_ , \new_[61485]_ , \new_[61488]_ ,
    \new_[61491]_ , \new_[61492]_ , \new_[61495]_ , \new_[61498]_ ,
    \new_[61499]_ , \new_[61500]_ , \new_[61503]_ , \new_[61506]_ ,
    \new_[61507]_ , \new_[61510]_ , \new_[61513]_ , \new_[61514]_ ,
    \new_[61515]_ , \new_[61518]_ , \new_[61521]_ , \new_[61522]_ ,
    \new_[61525]_ , \new_[61528]_ , \new_[61529]_ , \new_[61530]_ ,
    \new_[61533]_ , \new_[61536]_ , \new_[61537]_ , \new_[61540]_ ,
    \new_[61543]_ , \new_[61544]_ , \new_[61545]_ , \new_[61548]_ ,
    \new_[61551]_ , \new_[61552]_ , \new_[61555]_ , \new_[61558]_ ,
    \new_[61559]_ , \new_[61560]_ , \new_[61563]_ , \new_[61566]_ ,
    \new_[61567]_ , \new_[61570]_ , \new_[61573]_ , \new_[61574]_ ,
    \new_[61575]_ , \new_[61578]_ , \new_[61581]_ , \new_[61582]_ ,
    \new_[61585]_ , \new_[61588]_ , \new_[61589]_ , \new_[61590]_ ,
    \new_[61593]_ , \new_[61596]_ , \new_[61597]_ , \new_[61600]_ ,
    \new_[61603]_ , \new_[61604]_ , \new_[61605]_ , \new_[61608]_ ,
    \new_[61611]_ , \new_[61612]_ , \new_[61615]_ , \new_[61618]_ ,
    \new_[61619]_ , \new_[61620]_ , \new_[61623]_ , \new_[61626]_ ,
    \new_[61627]_ , \new_[61630]_ , \new_[61633]_ , \new_[61634]_ ,
    \new_[61635]_ , \new_[61638]_ , \new_[61641]_ , \new_[61642]_ ,
    \new_[61645]_ , \new_[61648]_ , \new_[61649]_ , \new_[61650]_ ,
    \new_[61653]_ , \new_[61656]_ , \new_[61657]_ , \new_[61660]_ ,
    \new_[61663]_ , \new_[61664]_ , \new_[61665]_ , \new_[61668]_ ,
    \new_[61671]_ , \new_[61672]_ , \new_[61675]_ , \new_[61678]_ ,
    \new_[61679]_ , \new_[61680]_ , \new_[61683]_ , \new_[61686]_ ,
    \new_[61687]_ , \new_[61690]_ , \new_[61693]_ , \new_[61694]_ ,
    \new_[61695]_ , \new_[61698]_ , \new_[61701]_ , \new_[61702]_ ,
    \new_[61705]_ , \new_[61708]_ , \new_[61709]_ , \new_[61710]_ ,
    \new_[61713]_ , \new_[61716]_ , \new_[61717]_ , \new_[61720]_ ,
    \new_[61723]_ , \new_[61724]_ , \new_[61725]_ , \new_[61728]_ ,
    \new_[61731]_ , \new_[61732]_ , \new_[61735]_ , \new_[61738]_ ,
    \new_[61739]_ , \new_[61740]_ , \new_[61743]_ , \new_[61746]_ ,
    \new_[61747]_ , \new_[61750]_ , \new_[61753]_ , \new_[61754]_ ,
    \new_[61755]_ , \new_[61758]_ , \new_[61761]_ , \new_[61762]_ ,
    \new_[61765]_ , \new_[61768]_ , \new_[61769]_ , \new_[61770]_ ,
    \new_[61773]_ , \new_[61776]_ , \new_[61777]_ , \new_[61780]_ ,
    \new_[61783]_ , \new_[61784]_ , \new_[61785]_ , \new_[61788]_ ,
    \new_[61791]_ , \new_[61792]_ , \new_[61795]_ , \new_[61798]_ ,
    \new_[61799]_ , \new_[61800]_ , \new_[61803]_ , \new_[61806]_ ,
    \new_[61807]_ , \new_[61810]_ , \new_[61813]_ , \new_[61814]_ ,
    \new_[61815]_ , \new_[61818]_ , \new_[61821]_ , \new_[61822]_ ,
    \new_[61825]_ , \new_[61828]_ , \new_[61829]_ , \new_[61830]_ ,
    \new_[61833]_ , \new_[61836]_ , \new_[61837]_ , \new_[61840]_ ,
    \new_[61843]_ , \new_[61844]_ , \new_[61845]_ , \new_[61848]_ ,
    \new_[61851]_ , \new_[61852]_ , \new_[61855]_ , \new_[61858]_ ,
    \new_[61859]_ , \new_[61860]_ , \new_[61863]_ , \new_[61866]_ ,
    \new_[61867]_ , \new_[61870]_ , \new_[61873]_ , \new_[61874]_ ,
    \new_[61875]_ , \new_[61878]_ , \new_[61881]_ , \new_[61882]_ ,
    \new_[61885]_ , \new_[61888]_ , \new_[61889]_ , \new_[61890]_ ,
    \new_[61893]_ , \new_[61896]_ , \new_[61897]_ , \new_[61900]_ ,
    \new_[61903]_ , \new_[61904]_ , \new_[61905]_ , \new_[61908]_ ,
    \new_[61911]_ , \new_[61912]_ , \new_[61915]_ , \new_[61918]_ ,
    \new_[61919]_ , \new_[61920]_ , \new_[61923]_ , \new_[61926]_ ,
    \new_[61927]_ , \new_[61930]_ , \new_[61933]_ , \new_[61934]_ ,
    \new_[61935]_ , \new_[61938]_ , \new_[61941]_ , \new_[61942]_ ,
    \new_[61945]_ , \new_[61948]_ , \new_[61949]_ , \new_[61950]_ ,
    \new_[61953]_ , \new_[61956]_ , \new_[61957]_ , \new_[61960]_ ,
    \new_[61963]_ , \new_[61964]_ , \new_[61965]_ , \new_[61968]_ ,
    \new_[61971]_ , \new_[61972]_ , \new_[61975]_ , \new_[61978]_ ,
    \new_[61979]_ , \new_[61980]_ , \new_[61983]_ , \new_[61986]_ ,
    \new_[61987]_ , \new_[61990]_ , \new_[61993]_ , \new_[61994]_ ,
    \new_[61995]_ , \new_[61998]_ , \new_[62001]_ , \new_[62002]_ ,
    \new_[62005]_ , \new_[62008]_ , \new_[62009]_ , \new_[62010]_ ,
    \new_[62013]_ , \new_[62016]_ , \new_[62017]_ , \new_[62020]_ ,
    \new_[62023]_ , \new_[62024]_ , \new_[62025]_ , \new_[62028]_ ,
    \new_[62031]_ , \new_[62032]_ , \new_[62035]_ , \new_[62038]_ ,
    \new_[62039]_ , \new_[62040]_ , \new_[62043]_ , \new_[62046]_ ,
    \new_[62047]_ , \new_[62050]_ , \new_[62053]_ , \new_[62054]_ ,
    \new_[62055]_ , \new_[62058]_ , \new_[62061]_ , \new_[62062]_ ,
    \new_[62065]_ , \new_[62068]_ , \new_[62069]_ , \new_[62070]_ ,
    \new_[62073]_ , \new_[62076]_ , \new_[62077]_ , \new_[62080]_ ,
    \new_[62083]_ , \new_[62084]_ , \new_[62085]_ , \new_[62088]_ ,
    \new_[62091]_ , \new_[62092]_ , \new_[62095]_ , \new_[62098]_ ,
    \new_[62099]_ , \new_[62100]_ , \new_[62103]_ , \new_[62106]_ ,
    \new_[62107]_ , \new_[62110]_ , \new_[62113]_ , \new_[62114]_ ,
    \new_[62115]_ , \new_[62118]_ , \new_[62121]_ , \new_[62122]_ ,
    \new_[62125]_ , \new_[62128]_ , \new_[62129]_ , \new_[62130]_ ,
    \new_[62133]_ , \new_[62136]_ , \new_[62137]_ , \new_[62140]_ ,
    \new_[62143]_ , \new_[62144]_ , \new_[62145]_ , \new_[62148]_ ,
    \new_[62151]_ , \new_[62152]_ , \new_[62155]_ , \new_[62158]_ ,
    \new_[62159]_ , \new_[62160]_ , \new_[62163]_ , \new_[62166]_ ,
    \new_[62167]_ , \new_[62170]_ , \new_[62173]_ , \new_[62174]_ ,
    \new_[62175]_ , \new_[62178]_ , \new_[62181]_ , \new_[62182]_ ,
    \new_[62185]_ , \new_[62188]_ , \new_[62189]_ , \new_[62190]_ ,
    \new_[62193]_ , \new_[62196]_ , \new_[62197]_ , \new_[62200]_ ,
    \new_[62203]_ , \new_[62204]_ , \new_[62205]_ , \new_[62208]_ ,
    \new_[62211]_ , \new_[62212]_ , \new_[62215]_ , \new_[62218]_ ,
    \new_[62219]_ , \new_[62220]_ , \new_[62223]_ , \new_[62226]_ ,
    \new_[62227]_ , \new_[62230]_ , \new_[62233]_ , \new_[62234]_ ,
    \new_[62235]_ , \new_[62238]_ , \new_[62241]_ , \new_[62242]_ ,
    \new_[62245]_ , \new_[62248]_ , \new_[62249]_ , \new_[62250]_ ,
    \new_[62253]_ , \new_[62256]_ , \new_[62257]_ , \new_[62260]_ ,
    \new_[62263]_ , \new_[62264]_ , \new_[62265]_ , \new_[62268]_ ,
    \new_[62271]_ , \new_[62272]_ , \new_[62275]_ , \new_[62278]_ ,
    \new_[62279]_ , \new_[62280]_ , \new_[62283]_ , \new_[62286]_ ,
    \new_[62287]_ , \new_[62290]_ , \new_[62293]_ , \new_[62294]_ ,
    \new_[62295]_ , \new_[62298]_ , \new_[62301]_ , \new_[62302]_ ,
    \new_[62305]_ , \new_[62308]_ , \new_[62309]_ , \new_[62310]_ ,
    \new_[62313]_ , \new_[62316]_ , \new_[62317]_ , \new_[62320]_ ,
    \new_[62323]_ , \new_[62324]_ , \new_[62325]_ , \new_[62328]_ ,
    \new_[62331]_ , \new_[62332]_ , \new_[62335]_ , \new_[62338]_ ,
    \new_[62339]_ , \new_[62340]_ , \new_[62343]_ , \new_[62346]_ ,
    \new_[62347]_ , \new_[62350]_ , \new_[62353]_ , \new_[62354]_ ,
    \new_[62355]_ , \new_[62358]_ , \new_[62361]_ , \new_[62362]_ ,
    \new_[62365]_ , \new_[62368]_ , \new_[62369]_ , \new_[62370]_ ,
    \new_[62373]_ , \new_[62376]_ , \new_[62377]_ , \new_[62380]_ ,
    \new_[62383]_ , \new_[62384]_ , \new_[62385]_ , \new_[62388]_ ,
    \new_[62391]_ , \new_[62392]_ , \new_[62395]_ , \new_[62398]_ ,
    \new_[62399]_ , \new_[62400]_ , \new_[62403]_ , \new_[62406]_ ,
    \new_[62407]_ , \new_[62410]_ , \new_[62413]_ , \new_[62414]_ ,
    \new_[62415]_ , \new_[62418]_ , \new_[62421]_ , \new_[62422]_ ,
    \new_[62425]_ , \new_[62428]_ , \new_[62429]_ , \new_[62430]_ ,
    \new_[62433]_ , \new_[62436]_ , \new_[62437]_ , \new_[62440]_ ,
    \new_[62443]_ , \new_[62444]_ , \new_[62445]_ , \new_[62448]_ ,
    \new_[62451]_ , \new_[62452]_ , \new_[62455]_ , \new_[62458]_ ,
    \new_[62459]_ , \new_[62460]_ , \new_[62463]_ , \new_[62466]_ ,
    \new_[62467]_ , \new_[62470]_ , \new_[62473]_ , \new_[62474]_ ,
    \new_[62475]_ , \new_[62478]_ , \new_[62481]_ , \new_[62482]_ ,
    \new_[62485]_ , \new_[62488]_ , \new_[62489]_ , \new_[62490]_ ,
    \new_[62493]_ , \new_[62496]_ , \new_[62497]_ , \new_[62500]_ ,
    \new_[62503]_ , \new_[62504]_ , \new_[62505]_ , \new_[62508]_ ,
    \new_[62511]_ , \new_[62512]_ , \new_[62515]_ , \new_[62518]_ ,
    \new_[62519]_ , \new_[62520]_ , \new_[62523]_ , \new_[62526]_ ,
    \new_[62527]_ , \new_[62530]_ , \new_[62533]_ , \new_[62534]_ ,
    \new_[62535]_ , \new_[62538]_ , \new_[62541]_ , \new_[62542]_ ,
    \new_[62545]_ , \new_[62548]_ , \new_[62549]_ , \new_[62550]_ ,
    \new_[62553]_ , \new_[62556]_ , \new_[62557]_ , \new_[62560]_ ,
    \new_[62563]_ , \new_[62564]_ , \new_[62565]_ , \new_[62568]_ ,
    \new_[62571]_ , \new_[62572]_ , \new_[62575]_ , \new_[62578]_ ,
    \new_[62579]_ , \new_[62580]_ , \new_[62583]_ , \new_[62586]_ ,
    \new_[62587]_ , \new_[62590]_ , \new_[62593]_ , \new_[62594]_ ,
    \new_[62595]_ , \new_[62598]_ , \new_[62601]_ , \new_[62602]_ ,
    \new_[62605]_ , \new_[62609]_ , \new_[62610]_ , \new_[62611]_ ,
    \new_[62612]_ , \new_[62615]_ , \new_[62618]_ , \new_[62619]_ ,
    \new_[62622]_ , \new_[62625]_ , \new_[62626]_ , \new_[62627]_ ,
    \new_[62630]_ , \new_[62633]_ , \new_[62634]_ , \new_[62637]_ ,
    \new_[62641]_ , \new_[62642]_ , \new_[62643]_ , \new_[62644]_ ,
    \new_[62647]_ , \new_[62650]_ , \new_[62651]_ , \new_[62654]_ ,
    \new_[62657]_ , \new_[62658]_ , \new_[62659]_ , \new_[62662]_ ,
    \new_[62665]_ , \new_[62666]_ , \new_[62669]_ , \new_[62673]_ ,
    \new_[62674]_ , \new_[62675]_ , \new_[62676]_ , \new_[62679]_ ,
    \new_[62682]_ , \new_[62683]_ , \new_[62686]_ , \new_[62689]_ ,
    \new_[62690]_ , \new_[62691]_ , \new_[62694]_ , \new_[62697]_ ,
    \new_[62698]_ , \new_[62701]_ , \new_[62705]_ , \new_[62706]_ ,
    \new_[62707]_ , \new_[62708]_ , \new_[62711]_ , \new_[62714]_ ,
    \new_[62715]_ , \new_[62718]_ , \new_[62721]_ , \new_[62722]_ ,
    \new_[62723]_ , \new_[62726]_ , \new_[62729]_ , \new_[62730]_ ,
    \new_[62733]_ , \new_[62737]_ , \new_[62738]_ , \new_[62739]_ ,
    \new_[62740]_ , \new_[62743]_ , \new_[62746]_ , \new_[62747]_ ,
    \new_[62750]_ , \new_[62753]_ , \new_[62754]_ , \new_[62755]_ ,
    \new_[62758]_ , \new_[62761]_ , \new_[62762]_ , \new_[62765]_ ,
    \new_[62769]_ , \new_[62770]_ , \new_[62771]_ , \new_[62772]_ ,
    \new_[62775]_ , \new_[62778]_ , \new_[62779]_ , \new_[62782]_ ,
    \new_[62785]_ , \new_[62786]_ , \new_[62787]_ , \new_[62790]_ ,
    \new_[62793]_ , \new_[62794]_ , \new_[62797]_ , \new_[62801]_ ,
    \new_[62802]_ , \new_[62803]_ , \new_[62804]_ , \new_[62807]_ ,
    \new_[62810]_ , \new_[62811]_ , \new_[62814]_ , \new_[62817]_ ,
    \new_[62818]_ , \new_[62819]_ , \new_[62822]_ , \new_[62825]_ ,
    \new_[62826]_ , \new_[62829]_ , \new_[62833]_ , \new_[62834]_ ,
    \new_[62835]_ , \new_[62836]_ , \new_[62839]_ , \new_[62842]_ ,
    \new_[62843]_ , \new_[62846]_ , \new_[62849]_ , \new_[62850]_ ,
    \new_[62851]_ , \new_[62854]_ , \new_[62857]_ , \new_[62858]_ ,
    \new_[62861]_ , \new_[62865]_ , \new_[62866]_ , \new_[62867]_ ,
    \new_[62868]_ , \new_[62871]_ , \new_[62874]_ , \new_[62875]_ ,
    \new_[62878]_ , \new_[62881]_ , \new_[62882]_ , \new_[62883]_ ,
    \new_[62886]_ , \new_[62889]_ , \new_[62890]_ , \new_[62893]_ ,
    \new_[62897]_ , \new_[62898]_ , \new_[62899]_ , \new_[62900]_ ,
    \new_[62903]_ , \new_[62906]_ , \new_[62907]_ , \new_[62910]_ ,
    \new_[62913]_ , \new_[62914]_ , \new_[62915]_ , \new_[62918]_ ,
    \new_[62921]_ , \new_[62922]_ , \new_[62925]_ , \new_[62929]_ ,
    \new_[62930]_ , \new_[62931]_ , \new_[62932]_ , \new_[62935]_ ,
    \new_[62938]_ , \new_[62939]_ , \new_[62942]_ , \new_[62945]_ ,
    \new_[62946]_ , \new_[62947]_ , \new_[62950]_ , \new_[62953]_ ,
    \new_[62954]_ , \new_[62957]_ , \new_[62961]_ , \new_[62962]_ ,
    \new_[62963]_ , \new_[62964]_ , \new_[62967]_ , \new_[62970]_ ,
    \new_[62971]_ , \new_[62974]_ , \new_[62977]_ , \new_[62978]_ ,
    \new_[62979]_ , \new_[62982]_ , \new_[62985]_ , \new_[62986]_ ,
    \new_[62989]_ , \new_[62993]_ , \new_[62994]_ , \new_[62995]_ ,
    \new_[62996]_ , \new_[62999]_ , \new_[63002]_ , \new_[63003]_ ,
    \new_[63006]_ , \new_[63009]_ , \new_[63010]_ , \new_[63011]_ ,
    \new_[63014]_ , \new_[63017]_ , \new_[63018]_ , \new_[63021]_ ,
    \new_[63025]_ , \new_[63026]_ , \new_[63027]_ , \new_[63028]_ ,
    \new_[63031]_ , \new_[63034]_ , \new_[63035]_ , \new_[63038]_ ,
    \new_[63041]_ , \new_[63042]_ , \new_[63043]_ , \new_[63046]_ ,
    \new_[63049]_ , \new_[63050]_ , \new_[63053]_ , \new_[63057]_ ,
    \new_[63058]_ , \new_[63059]_ , \new_[63060]_ , \new_[63063]_ ,
    \new_[63066]_ , \new_[63067]_ , \new_[63070]_ , \new_[63073]_ ,
    \new_[63074]_ , \new_[63075]_ , \new_[63078]_ , \new_[63081]_ ,
    \new_[63082]_ , \new_[63085]_ , \new_[63089]_ , \new_[63090]_ ,
    \new_[63091]_ , \new_[63092]_ , \new_[63095]_ , \new_[63098]_ ,
    \new_[63099]_ , \new_[63102]_ , \new_[63105]_ , \new_[63106]_ ,
    \new_[63107]_ , \new_[63110]_ , \new_[63113]_ , \new_[63114]_ ,
    \new_[63117]_ , \new_[63121]_ , \new_[63122]_ , \new_[63123]_ ,
    \new_[63124]_ , \new_[63127]_ , \new_[63130]_ , \new_[63131]_ ,
    \new_[63134]_ , \new_[63137]_ , \new_[63138]_ , \new_[63139]_ ,
    \new_[63142]_ , \new_[63145]_ , \new_[63146]_ , \new_[63149]_ ,
    \new_[63153]_ , \new_[63154]_ , \new_[63155]_ , \new_[63156]_ ,
    \new_[63159]_ , \new_[63162]_ , \new_[63163]_ , \new_[63166]_ ,
    \new_[63169]_ , \new_[63170]_ , \new_[63171]_ , \new_[63174]_ ,
    \new_[63177]_ , \new_[63178]_ , \new_[63181]_ , \new_[63185]_ ,
    \new_[63186]_ , \new_[63187]_ , \new_[63188]_ , \new_[63191]_ ,
    \new_[63194]_ , \new_[63195]_ , \new_[63198]_ , \new_[63201]_ ,
    \new_[63202]_ , \new_[63203]_ , \new_[63206]_ , \new_[63209]_ ,
    \new_[63210]_ , \new_[63213]_ , \new_[63217]_ , \new_[63218]_ ,
    \new_[63219]_ , \new_[63220]_ , \new_[63223]_ , \new_[63226]_ ,
    \new_[63227]_ , \new_[63230]_ , \new_[63233]_ , \new_[63234]_ ,
    \new_[63235]_ , \new_[63238]_ , \new_[63241]_ , \new_[63242]_ ,
    \new_[63245]_ , \new_[63249]_ , \new_[63250]_ , \new_[63251]_ ,
    \new_[63252]_ , \new_[63255]_ , \new_[63258]_ , \new_[63259]_ ,
    \new_[63262]_ , \new_[63265]_ , \new_[63266]_ , \new_[63267]_ ,
    \new_[63270]_ , \new_[63273]_ , \new_[63274]_ , \new_[63277]_ ,
    \new_[63281]_ , \new_[63282]_ , \new_[63283]_ , \new_[63284]_ ,
    \new_[63287]_ , \new_[63290]_ , \new_[63291]_ , \new_[63294]_ ,
    \new_[63297]_ , \new_[63298]_ , \new_[63299]_ , \new_[63302]_ ,
    \new_[63305]_ , \new_[63306]_ , \new_[63309]_ , \new_[63313]_ ,
    \new_[63314]_ , \new_[63315]_ , \new_[63316]_ , \new_[63319]_ ,
    \new_[63322]_ , \new_[63323]_ , \new_[63326]_ , \new_[63329]_ ,
    \new_[63330]_ , \new_[63331]_ , \new_[63334]_ , \new_[63337]_ ,
    \new_[63338]_ , \new_[63341]_ , \new_[63345]_ , \new_[63346]_ ,
    \new_[63347]_ , \new_[63348]_ , \new_[63351]_ , \new_[63354]_ ,
    \new_[63355]_ , \new_[63358]_ , \new_[63361]_ , \new_[63362]_ ,
    \new_[63363]_ , \new_[63366]_ , \new_[63369]_ , \new_[63370]_ ,
    \new_[63373]_ , \new_[63377]_ , \new_[63378]_ , \new_[63379]_ ,
    \new_[63380]_ , \new_[63383]_ , \new_[63386]_ , \new_[63387]_ ,
    \new_[63390]_ , \new_[63393]_ , \new_[63394]_ , \new_[63395]_ ,
    \new_[63398]_ , \new_[63401]_ , \new_[63402]_ , \new_[63405]_ ,
    \new_[63409]_ , \new_[63410]_ , \new_[63411]_ , \new_[63412]_ ,
    \new_[63415]_ , \new_[63418]_ , \new_[63419]_ , \new_[63422]_ ,
    \new_[63425]_ , \new_[63426]_ , \new_[63427]_ , \new_[63430]_ ,
    \new_[63433]_ , \new_[63434]_ , \new_[63437]_ , \new_[63441]_ ,
    \new_[63442]_ , \new_[63443]_ , \new_[63444]_ , \new_[63447]_ ,
    \new_[63450]_ , \new_[63451]_ , \new_[63454]_ , \new_[63457]_ ,
    \new_[63458]_ , \new_[63459]_ , \new_[63462]_ , \new_[63465]_ ,
    \new_[63466]_ , \new_[63469]_ , \new_[63473]_ , \new_[63474]_ ,
    \new_[63475]_ , \new_[63476]_ , \new_[63479]_ , \new_[63482]_ ,
    \new_[63483]_ , \new_[63486]_ , \new_[63489]_ , \new_[63490]_ ,
    \new_[63491]_ , \new_[63494]_ , \new_[63497]_ , \new_[63498]_ ,
    \new_[63501]_ , \new_[63505]_ , \new_[63506]_ , \new_[63507]_ ,
    \new_[63508]_ , \new_[63511]_ , \new_[63514]_ , \new_[63515]_ ,
    \new_[63518]_ , \new_[63521]_ , \new_[63522]_ , \new_[63523]_ ,
    \new_[63526]_ , \new_[63529]_ , \new_[63530]_ , \new_[63533]_ ,
    \new_[63537]_ , \new_[63538]_ , \new_[63539]_ , \new_[63540]_ ,
    \new_[63543]_ , \new_[63546]_ , \new_[63547]_ , \new_[63550]_ ,
    \new_[63553]_ , \new_[63554]_ , \new_[63555]_ , \new_[63558]_ ,
    \new_[63561]_ , \new_[63562]_ , \new_[63565]_ , \new_[63569]_ ,
    \new_[63570]_ , \new_[63571]_ , \new_[63572]_ , \new_[63575]_ ,
    \new_[63578]_ , \new_[63579]_ , \new_[63582]_ , \new_[63585]_ ,
    \new_[63586]_ , \new_[63587]_ , \new_[63590]_ , \new_[63593]_ ,
    \new_[63594]_ , \new_[63597]_ , \new_[63601]_ , \new_[63602]_ ,
    \new_[63603]_ , \new_[63604]_ , \new_[63607]_ , \new_[63610]_ ,
    \new_[63611]_ , \new_[63614]_ , \new_[63617]_ , \new_[63618]_ ,
    \new_[63619]_ , \new_[63622]_ , \new_[63625]_ , \new_[63626]_ ,
    \new_[63629]_ , \new_[63633]_ , \new_[63634]_ , \new_[63635]_ ,
    \new_[63636]_ , \new_[63639]_ , \new_[63642]_ , \new_[63643]_ ,
    \new_[63646]_ , \new_[63649]_ , \new_[63650]_ , \new_[63651]_ ,
    \new_[63654]_ , \new_[63657]_ , \new_[63658]_ , \new_[63661]_ ,
    \new_[63665]_ , \new_[63666]_ , \new_[63667]_ , \new_[63668]_ ,
    \new_[63671]_ , \new_[63674]_ , \new_[63675]_ , \new_[63678]_ ,
    \new_[63681]_ , \new_[63682]_ , \new_[63683]_ , \new_[63686]_ ,
    \new_[63689]_ , \new_[63690]_ , \new_[63693]_ , \new_[63697]_ ,
    \new_[63698]_ , \new_[63699]_ , \new_[63700]_ , \new_[63703]_ ,
    \new_[63706]_ , \new_[63707]_ , \new_[63710]_ , \new_[63713]_ ,
    \new_[63714]_ , \new_[63715]_ , \new_[63718]_ , \new_[63721]_ ,
    \new_[63722]_ , \new_[63725]_ , \new_[63729]_ , \new_[63730]_ ,
    \new_[63731]_ , \new_[63732]_ , \new_[63735]_ , \new_[63738]_ ,
    \new_[63739]_ , \new_[63742]_ , \new_[63745]_ , \new_[63746]_ ,
    \new_[63747]_ , \new_[63750]_ , \new_[63753]_ , \new_[63754]_ ,
    \new_[63757]_ , \new_[63761]_ , \new_[63762]_ , \new_[63763]_ ,
    \new_[63764]_ , \new_[63767]_ , \new_[63770]_ , \new_[63771]_ ,
    \new_[63774]_ , \new_[63777]_ , \new_[63778]_ , \new_[63779]_ ,
    \new_[63782]_ , \new_[63785]_ , \new_[63786]_ , \new_[63789]_ ,
    \new_[63793]_ , \new_[63794]_ , \new_[63795]_ , \new_[63796]_ ,
    \new_[63799]_ , \new_[63802]_ , \new_[63803]_ , \new_[63806]_ ,
    \new_[63809]_ , \new_[63810]_ , \new_[63811]_ , \new_[63814]_ ,
    \new_[63817]_ , \new_[63818]_ , \new_[63821]_ , \new_[63825]_ ,
    \new_[63826]_ , \new_[63827]_ , \new_[63828]_ , \new_[63831]_ ,
    \new_[63834]_ , \new_[63835]_ , \new_[63838]_ , \new_[63841]_ ,
    \new_[63842]_ , \new_[63843]_ , \new_[63846]_ , \new_[63849]_ ,
    \new_[63850]_ , \new_[63853]_ , \new_[63857]_ , \new_[63858]_ ,
    \new_[63859]_ , \new_[63860]_ , \new_[63863]_ , \new_[63866]_ ,
    \new_[63867]_ , \new_[63870]_ , \new_[63873]_ , \new_[63874]_ ,
    \new_[63875]_ , \new_[63878]_ , \new_[63881]_ , \new_[63882]_ ,
    \new_[63885]_ , \new_[63889]_ , \new_[63890]_ , \new_[63891]_ ,
    \new_[63892]_ , \new_[63895]_ , \new_[63898]_ , \new_[63899]_ ,
    \new_[63902]_ , \new_[63905]_ , \new_[63906]_ , \new_[63907]_ ,
    \new_[63910]_ , \new_[63913]_ , \new_[63914]_ , \new_[63917]_ ,
    \new_[63921]_ , \new_[63922]_ , \new_[63923]_ , \new_[63924]_ ,
    \new_[63927]_ , \new_[63930]_ , \new_[63931]_ , \new_[63934]_ ,
    \new_[63937]_ , \new_[63938]_ , \new_[63939]_ , \new_[63942]_ ,
    \new_[63945]_ , \new_[63946]_ , \new_[63949]_ , \new_[63953]_ ,
    \new_[63954]_ , \new_[63955]_ , \new_[63956]_ , \new_[63959]_ ,
    \new_[63962]_ , \new_[63963]_ , \new_[63966]_ , \new_[63969]_ ,
    \new_[63970]_ , \new_[63971]_ , \new_[63974]_ , \new_[63977]_ ,
    \new_[63978]_ , \new_[63981]_ , \new_[63985]_ , \new_[63986]_ ,
    \new_[63987]_ , \new_[63988]_ , \new_[63991]_ , \new_[63994]_ ,
    \new_[63995]_ , \new_[63998]_ , \new_[64001]_ , \new_[64002]_ ,
    \new_[64003]_ , \new_[64006]_ , \new_[64009]_ , \new_[64010]_ ,
    \new_[64013]_ , \new_[64017]_ , \new_[64018]_ , \new_[64019]_ ,
    \new_[64020]_ , \new_[64023]_ , \new_[64026]_ , \new_[64027]_ ,
    \new_[64030]_ , \new_[64033]_ , \new_[64034]_ , \new_[64035]_ ,
    \new_[64038]_ , \new_[64041]_ , \new_[64042]_ , \new_[64045]_ ,
    \new_[64049]_ , \new_[64050]_ , \new_[64051]_ , \new_[64052]_ ,
    \new_[64055]_ , \new_[64058]_ , \new_[64059]_ , \new_[64062]_ ,
    \new_[64065]_ , \new_[64066]_ , \new_[64067]_ , \new_[64070]_ ,
    \new_[64073]_ , \new_[64074]_ , \new_[64077]_ , \new_[64081]_ ,
    \new_[64082]_ , \new_[64083]_ , \new_[64084]_ , \new_[64087]_ ,
    \new_[64090]_ , \new_[64091]_ , \new_[64094]_ , \new_[64097]_ ,
    \new_[64098]_ , \new_[64099]_ , \new_[64102]_ , \new_[64105]_ ,
    \new_[64106]_ , \new_[64109]_ , \new_[64113]_ , \new_[64114]_ ,
    \new_[64115]_ , \new_[64116]_ , \new_[64119]_ , \new_[64122]_ ,
    \new_[64123]_ , \new_[64126]_ , \new_[64129]_ , \new_[64130]_ ,
    \new_[64131]_ , \new_[64134]_ , \new_[64137]_ , \new_[64138]_ ,
    \new_[64141]_ , \new_[64145]_ , \new_[64146]_ , \new_[64147]_ ,
    \new_[64148]_ , \new_[64151]_ , \new_[64154]_ , \new_[64155]_ ,
    \new_[64158]_ , \new_[64161]_ , \new_[64162]_ , \new_[64163]_ ,
    \new_[64166]_ , \new_[64169]_ , \new_[64170]_ , \new_[64173]_ ,
    \new_[64177]_ , \new_[64178]_ , \new_[64179]_ , \new_[64180]_ ,
    \new_[64183]_ , \new_[64186]_ , \new_[64187]_ , \new_[64190]_ ,
    \new_[64193]_ , \new_[64194]_ , \new_[64195]_ , \new_[64198]_ ,
    \new_[64201]_ , \new_[64202]_ , \new_[64205]_ , \new_[64209]_ ,
    \new_[64210]_ , \new_[64211]_ , \new_[64212]_ , \new_[64215]_ ,
    \new_[64218]_ , \new_[64219]_ , \new_[64222]_ , \new_[64225]_ ,
    \new_[64226]_ , \new_[64227]_ , \new_[64230]_ , \new_[64233]_ ,
    \new_[64234]_ , \new_[64237]_ , \new_[64241]_ , \new_[64242]_ ,
    \new_[64243]_ , \new_[64244]_ , \new_[64247]_ , \new_[64250]_ ,
    \new_[64251]_ , \new_[64254]_ , \new_[64257]_ , \new_[64258]_ ,
    \new_[64259]_ , \new_[64262]_ , \new_[64265]_ , \new_[64266]_ ,
    \new_[64269]_ , \new_[64273]_ , \new_[64274]_ , \new_[64275]_ ,
    \new_[64276]_ , \new_[64279]_ , \new_[64282]_ , \new_[64283]_ ,
    \new_[64286]_ , \new_[64289]_ , \new_[64290]_ , \new_[64291]_ ,
    \new_[64294]_ , \new_[64297]_ , \new_[64298]_ , \new_[64301]_ ,
    \new_[64305]_ , \new_[64306]_ , \new_[64307]_ , \new_[64308]_ ,
    \new_[64311]_ , \new_[64314]_ , \new_[64315]_ , \new_[64318]_ ,
    \new_[64321]_ , \new_[64322]_ , \new_[64323]_ , \new_[64326]_ ,
    \new_[64329]_ , \new_[64330]_ , \new_[64333]_ , \new_[64337]_ ,
    \new_[64338]_ , \new_[64339]_ , \new_[64340]_ , \new_[64343]_ ,
    \new_[64346]_ , \new_[64347]_ , \new_[64350]_ , \new_[64353]_ ,
    \new_[64354]_ , \new_[64355]_ , \new_[64358]_ , \new_[64361]_ ,
    \new_[64362]_ , \new_[64365]_ , \new_[64369]_ , \new_[64370]_ ,
    \new_[64371]_ , \new_[64372]_ , \new_[64375]_ , \new_[64378]_ ,
    \new_[64379]_ , \new_[64382]_ , \new_[64385]_ , \new_[64386]_ ,
    \new_[64387]_ , \new_[64390]_ , \new_[64393]_ , \new_[64394]_ ,
    \new_[64397]_ , \new_[64401]_ , \new_[64402]_ , \new_[64403]_ ,
    \new_[64404]_ , \new_[64407]_ , \new_[64410]_ , \new_[64411]_ ,
    \new_[64414]_ , \new_[64417]_ , \new_[64418]_ , \new_[64419]_ ,
    \new_[64422]_ , \new_[64425]_ , \new_[64426]_ , \new_[64429]_ ,
    \new_[64433]_ , \new_[64434]_ , \new_[64435]_ , \new_[64436]_ ,
    \new_[64439]_ , \new_[64442]_ , \new_[64443]_ , \new_[64446]_ ,
    \new_[64449]_ , \new_[64450]_ , \new_[64451]_ , \new_[64454]_ ,
    \new_[64457]_ , \new_[64458]_ , \new_[64461]_ , \new_[64465]_ ,
    \new_[64466]_ , \new_[64467]_ , \new_[64468]_ , \new_[64471]_ ,
    \new_[64474]_ , \new_[64475]_ , \new_[64478]_ , \new_[64481]_ ,
    \new_[64482]_ , \new_[64483]_ , \new_[64486]_ , \new_[64489]_ ,
    \new_[64490]_ , \new_[64493]_ , \new_[64497]_ , \new_[64498]_ ,
    \new_[64499]_ , \new_[64500]_ , \new_[64503]_ , \new_[64506]_ ,
    \new_[64507]_ , \new_[64510]_ , \new_[64513]_ , \new_[64514]_ ,
    \new_[64515]_ , \new_[64518]_ , \new_[64521]_ , \new_[64522]_ ,
    \new_[64525]_ , \new_[64529]_ , \new_[64530]_ , \new_[64531]_ ,
    \new_[64532]_ , \new_[64535]_ , \new_[64538]_ , \new_[64539]_ ,
    \new_[64542]_ , \new_[64545]_ , \new_[64546]_ , \new_[64547]_ ,
    \new_[64550]_ , \new_[64553]_ , \new_[64554]_ , \new_[64557]_ ,
    \new_[64561]_ , \new_[64562]_ , \new_[64563]_ , \new_[64564]_ ,
    \new_[64567]_ , \new_[64570]_ , \new_[64571]_ , \new_[64574]_ ,
    \new_[64577]_ , \new_[64578]_ , \new_[64579]_ , \new_[64582]_ ,
    \new_[64585]_ , \new_[64586]_ , \new_[64589]_ , \new_[64593]_ ,
    \new_[64594]_ , \new_[64595]_ , \new_[64596]_ , \new_[64599]_ ,
    \new_[64602]_ , \new_[64603]_ , \new_[64606]_ , \new_[64609]_ ,
    \new_[64610]_ , \new_[64611]_ , \new_[64614]_ , \new_[64617]_ ,
    \new_[64618]_ , \new_[64621]_ , \new_[64625]_ , \new_[64626]_ ,
    \new_[64627]_ , \new_[64628]_ , \new_[64631]_ , \new_[64634]_ ,
    \new_[64635]_ , \new_[64638]_ , \new_[64641]_ , \new_[64642]_ ,
    \new_[64643]_ , \new_[64646]_ , \new_[64649]_ , \new_[64650]_ ,
    \new_[64653]_ , \new_[64657]_ , \new_[64658]_ , \new_[64659]_ ,
    \new_[64660]_ , \new_[64663]_ , \new_[64666]_ , \new_[64667]_ ,
    \new_[64670]_ , \new_[64673]_ , \new_[64674]_ , \new_[64675]_ ,
    \new_[64678]_ , \new_[64681]_ , \new_[64682]_ , \new_[64685]_ ,
    \new_[64689]_ , \new_[64690]_ , \new_[64691]_ , \new_[64692]_ ,
    \new_[64695]_ , \new_[64698]_ , \new_[64699]_ , \new_[64702]_ ,
    \new_[64705]_ , \new_[64706]_ , \new_[64707]_ , \new_[64710]_ ,
    \new_[64713]_ , \new_[64714]_ , \new_[64717]_ , \new_[64721]_ ,
    \new_[64722]_ , \new_[64723]_ , \new_[64724]_ , \new_[64727]_ ,
    \new_[64730]_ , \new_[64731]_ , \new_[64734]_ , \new_[64737]_ ,
    \new_[64738]_ , \new_[64739]_ , \new_[64742]_ , \new_[64745]_ ,
    \new_[64746]_ , \new_[64749]_ , \new_[64753]_ , \new_[64754]_ ,
    \new_[64755]_ , \new_[64756]_ , \new_[64759]_ , \new_[64762]_ ,
    \new_[64763]_ , \new_[64766]_ , \new_[64769]_ , \new_[64770]_ ,
    \new_[64771]_ , \new_[64774]_ , \new_[64777]_ , \new_[64778]_ ,
    \new_[64781]_ , \new_[64785]_ , \new_[64786]_ , \new_[64787]_ ,
    \new_[64788]_ , \new_[64791]_ , \new_[64794]_ , \new_[64795]_ ,
    \new_[64798]_ , \new_[64801]_ , \new_[64802]_ , \new_[64803]_ ,
    \new_[64806]_ , \new_[64809]_ , \new_[64810]_ , \new_[64813]_ ,
    \new_[64817]_ , \new_[64818]_ , \new_[64819]_ , \new_[64820]_ ,
    \new_[64823]_ , \new_[64826]_ , \new_[64827]_ , \new_[64830]_ ,
    \new_[64833]_ , \new_[64834]_ , \new_[64835]_ , \new_[64838]_ ,
    \new_[64841]_ , \new_[64842]_ , \new_[64845]_ , \new_[64849]_ ,
    \new_[64850]_ , \new_[64851]_ , \new_[64852]_ , \new_[64855]_ ,
    \new_[64858]_ , \new_[64859]_ , \new_[64862]_ , \new_[64865]_ ,
    \new_[64866]_ , \new_[64867]_ , \new_[64870]_ , \new_[64873]_ ,
    \new_[64874]_ , \new_[64877]_ , \new_[64881]_ , \new_[64882]_ ,
    \new_[64883]_ , \new_[64884]_ , \new_[64887]_ , \new_[64890]_ ,
    \new_[64891]_ , \new_[64894]_ , \new_[64897]_ , \new_[64898]_ ,
    \new_[64899]_ , \new_[64902]_ , \new_[64905]_ , \new_[64906]_ ,
    \new_[64909]_ , \new_[64913]_ , \new_[64914]_ , \new_[64915]_ ,
    \new_[64916]_ , \new_[64919]_ , \new_[64922]_ , \new_[64923]_ ,
    \new_[64926]_ , \new_[64929]_ , \new_[64930]_ , \new_[64931]_ ,
    \new_[64934]_ , \new_[64937]_ , \new_[64938]_ , \new_[64941]_ ,
    \new_[64945]_ , \new_[64946]_ , \new_[64947]_ , \new_[64948]_ ,
    \new_[64951]_ , \new_[64954]_ , \new_[64955]_ , \new_[64958]_ ,
    \new_[64961]_ , \new_[64962]_ , \new_[64963]_ , \new_[64966]_ ,
    \new_[64969]_ , \new_[64970]_ , \new_[64973]_ , \new_[64977]_ ,
    \new_[64978]_ , \new_[64979]_ , \new_[64980]_ , \new_[64983]_ ,
    \new_[64986]_ , \new_[64987]_ , \new_[64990]_ , \new_[64993]_ ,
    \new_[64994]_ , \new_[64995]_ , \new_[64998]_ , \new_[65001]_ ,
    \new_[65002]_ , \new_[65005]_ , \new_[65009]_ , \new_[65010]_ ,
    \new_[65011]_ , \new_[65012]_ , \new_[65015]_ , \new_[65018]_ ,
    \new_[65019]_ , \new_[65022]_ , \new_[65025]_ , \new_[65026]_ ,
    \new_[65027]_ , \new_[65030]_ , \new_[65033]_ , \new_[65034]_ ,
    \new_[65037]_ , \new_[65041]_ , \new_[65042]_ , \new_[65043]_ ,
    \new_[65044]_ , \new_[65047]_ , \new_[65050]_ , \new_[65051]_ ,
    \new_[65054]_ , \new_[65057]_ , \new_[65058]_ , \new_[65059]_ ,
    \new_[65062]_ , \new_[65065]_ , \new_[65066]_ , \new_[65069]_ ,
    \new_[65073]_ , \new_[65074]_ , \new_[65075]_ , \new_[65076]_ ,
    \new_[65079]_ , \new_[65082]_ , \new_[65083]_ , \new_[65086]_ ,
    \new_[65089]_ , \new_[65090]_ , \new_[65091]_ , \new_[65094]_ ,
    \new_[65097]_ , \new_[65098]_ , \new_[65101]_ , \new_[65105]_ ,
    \new_[65106]_ , \new_[65107]_ , \new_[65108]_ , \new_[65111]_ ,
    \new_[65114]_ , \new_[65115]_ , \new_[65118]_ , \new_[65121]_ ,
    \new_[65122]_ , \new_[65123]_ , \new_[65126]_ , \new_[65129]_ ,
    \new_[65130]_ , \new_[65133]_ , \new_[65137]_ , \new_[65138]_ ,
    \new_[65139]_ , \new_[65140]_ , \new_[65143]_ , \new_[65146]_ ,
    \new_[65147]_ , \new_[65150]_ , \new_[65153]_ , \new_[65154]_ ,
    \new_[65155]_ , \new_[65158]_ , \new_[65161]_ , \new_[65162]_ ,
    \new_[65165]_ , \new_[65169]_ , \new_[65170]_ , \new_[65171]_ ,
    \new_[65172]_ , \new_[65175]_ , \new_[65178]_ , \new_[65179]_ ,
    \new_[65182]_ , \new_[65185]_ , \new_[65186]_ , \new_[65187]_ ,
    \new_[65190]_ , \new_[65193]_ , \new_[65194]_ , \new_[65197]_ ,
    \new_[65201]_ , \new_[65202]_ , \new_[65203]_ , \new_[65204]_ ,
    \new_[65207]_ , \new_[65210]_ , \new_[65211]_ , \new_[65214]_ ,
    \new_[65217]_ , \new_[65218]_ , \new_[65219]_ , \new_[65222]_ ,
    \new_[65225]_ , \new_[65226]_ , \new_[65229]_ , \new_[65233]_ ,
    \new_[65234]_ , \new_[65235]_ , \new_[65236]_ , \new_[65239]_ ,
    \new_[65242]_ , \new_[65243]_ , \new_[65246]_ , \new_[65249]_ ,
    \new_[65250]_ , \new_[65251]_ , \new_[65254]_ , \new_[65257]_ ,
    \new_[65258]_ , \new_[65261]_ , \new_[65265]_ , \new_[65266]_ ,
    \new_[65267]_ , \new_[65268]_ , \new_[65271]_ , \new_[65274]_ ,
    \new_[65275]_ , \new_[65278]_ , \new_[65281]_ , \new_[65282]_ ,
    \new_[65283]_ , \new_[65286]_ , \new_[65289]_ , \new_[65290]_ ,
    \new_[65293]_ , \new_[65297]_ , \new_[65298]_ , \new_[65299]_ ,
    \new_[65300]_ , \new_[65303]_ , \new_[65306]_ , \new_[65307]_ ,
    \new_[65310]_ , \new_[65313]_ , \new_[65314]_ , \new_[65315]_ ,
    \new_[65318]_ , \new_[65321]_ , \new_[65322]_ , \new_[65325]_ ,
    \new_[65329]_ , \new_[65330]_ , \new_[65331]_ , \new_[65332]_ ,
    \new_[65335]_ , \new_[65338]_ , \new_[65339]_ , \new_[65342]_ ,
    \new_[65345]_ , \new_[65346]_ , \new_[65347]_ , \new_[65350]_ ,
    \new_[65353]_ , \new_[65354]_ , \new_[65357]_ , \new_[65361]_ ,
    \new_[65362]_ , \new_[65363]_ , \new_[65364]_ , \new_[65367]_ ,
    \new_[65370]_ , \new_[65371]_ , \new_[65374]_ , \new_[65377]_ ,
    \new_[65378]_ , \new_[65379]_ , \new_[65382]_ , \new_[65385]_ ,
    \new_[65386]_ , \new_[65389]_ , \new_[65393]_ , \new_[65394]_ ,
    \new_[65395]_ , \new_[65396]_ , \new_[65399]_ , \new_[65402]_ ,
    \new_[65403]_ , \new_[65406]_ , \new_[65409]_ , \new_[65410]_ ,
    \new_[65411]_ , \new_[65414]_ , \new_[65417]_ , \new_[65418]_ ,
    \new_[65421]_ , \new_[65425]_ , \new_[65426]_ , \new_[65427]_ ,
    \new_[65428]_ , \new_[65431]_ , \new_[65434]_ , \new_[65435]_ ,
    \new_[65438]_ , \new_[65441]_ , \new_[65442]_ , \new_[65443]_ ,
    \new_[65446]_ , \new_[65449]_ , \new_[65450]_ , \new_[65453]_ ,
    \new_[65457]_ , \new_[65458]_ , \new_[65459]_ , \new_[65460]_ ,
    \new_[65463]_ , \new_[65466]_ , \new_[65467]_ , \new_[65470]_ ,
    \new_[65473]_ , \new_[65474]_ , \new_[65475]_ , \new_[65478]_ ,
    \new_[65481]_ , \new_[65482]_ , \new_[65485]_ , \new_[65489]_ ,
    \new_[65490]_ , \new_[65491]_ , \new_[65492]_ , \new_[65495]_ ,
    \new_[65498]_ , \new_[65499]_ , \new_[65502]_ , \new_[65505]_ ,
    \new_[65506]_ , \new_[65507]_ , \new_[65510]_ , \new_[65513]_ ,
    \new_[65514]_ , \new_[65517]_ , \new_[65521]_ , \new_[65522]_ ,
    \new_[65523]_ , \new_[65524]_ , \new_[65527]_ , \new_[65530]_ ,
    \new_[65531]_ , \new_[65534]_ , \new_[65537]_ , \new_[65538]_ ,
    \new_[65539]_ , \new_[65542]_ , \new_[65545]_ , \new_[65546]_ ,
    \new_[65549]_ , \new_[65553]_ , \new_[65554]_ , \new_[65555]_ ,
    \new_[65556]_ , \new_[65559]_ , \new_[65562]_ , \new_[65563]_ ,
    \new_[65566]_ , \new_[65569]_ , \new_[65570]_ , \new_[65571]_ ,
    \new_[65574]_ , \new_[65577]_ , \new_[65578]_ , \new_[65581]_ ,
    \new_[65585]_ , \new_[65586]_ , \new_[65587]_ , \new_[65588]_ ,
    \new_[65591]_ , \new_[65594]_ , \new_[65595]_ , \new_[65598]_ ,
    \new_[65601]_ , \new_[65602]_ , \new_[65603]_ , \new_[65606]_ ,
    \new_[65609]_ , \new_[65610]_ , \new_[65613]_ , \new_[65617]_ ,
    \new_[65618]_ , \new_[65619]_ , \new_[65620]_ , \new_[65623]_ ,
    \new_[65626]_ , \new_[65627]_ , \new_[65630]_ , \new_[65633]_ ,
    \new_[65634]_ , \new_[65635]_ , \new_[65638]_ , \new_[65641]_ ,
    \new_[65642]_ , \new_[65645]_ , \new_[65649]_ , \new_[65650]_ ,
    \new_[65651]_ , \new_[65652]_ , \new_[65655]_ , \new_[65658]_ ,
    \new_[65659]_ , \new_[65662]_ , \new_[65665]_ , \new_[65666]_ ,
    \new_[65667]_ , \new_[65670]_ , \new_[65673]_ , \new_[65674]_ ,
    \new_[65677]_ , \new_[65681]_ , \new_[65682]_ , \new_[65683]_ ,
    \new_[65684]_ , \new_[65687]_ , \new_[65690]_ , \new_[65691]_ ,
    \new_[65694]_ , \new_[65697]_ , \new_[65698]_ , \new_[65699]_ ,
    \new_[65702]_ , \new_[65705]_ , \new_[65706]_ , \new_[65709]_ ,
    \new_[65713]_ , \new_[65714]_ , \new_[65715]_ , \new_[65716]_ ,
    \new_[65719]_ , \new_[65722]_ , \new_[65723]_ , \new_[65726]_ ,
    \new_[65729]_ , \new_[65730]_ , \new_[65731]_ , \new_[65734]_ ,
    \new_[65737]_ , \new_[65738]_ , \new_[65741]_ , \new_[65745]_ ,
    \new_[65746]_ , \new_[65747]_ , \new_[65748]_ , \new_[65751]_ ,
    \new_[65754]_ , \new_[65755]_ , \new_[65758]_ , \new_[65761]_ ,
    \new_[65762]_ , \new_[65763]_ , \new_[65766]_ , \new_[65769]_ ,
    \new_[65770]_ , \new_[65773]_ , \new_[65777]_ , \new_[65778]_ ,
    \new_[65779]_ , \new_[65780]_ , \new_[65783]_ , \new_[65786]_ ,
    \new_[65787]_ , \new_[65790]_ , \new_[65793]_ , \new_[65794]_ ,
    \new_[65795]_ , \new_[65798]_ , \new_[65801]_ , \new_[65802]_ ,
    \new_[65805]_ , \new_[65809]_ , \new_[65810]_ , \new_[65811]_ ,
    \new_[65812]_ , \new_[65815]_ , \new_[65818]_ , \new_[65819]_ ,
    \new_[65822]_ , \new_[65825]_ , \new_[65826]_ , \new_[65827]_ ,
    \new_[65830]_ , \new_[65833]_ , \new_[65834]_ , \new_[65837]_ ,
    \new_[65841]_ , \new_[65842]_ , \new_[65843]_ , \new_[65844]_ ,
    \new_[65847]_ , \new_[65850]_ , \new_[65851]_ , \new_[65854]_ ,
    \new_[65857]_ , \new_[65858]_ , \new_[65859]_ , \new_[65862]_ ,
    \new_[65865]_ , \new_[65866]_ , \new_[65869]_ , \new_[65873]_ ,
    \new_[65874]_ , \new_[65875]_ , \new_[65876]_ , \new_[65879]_ ,
    \new_[65882]_ , \new_[65883]_ , \new_[65886]_ , \new_[65889]_ ,
    \new_[65890]_ , \new_[65891]_ , \new_[65894]_ , \new_[65897]_ ,
    \new_[65898]_ , \new_[65901]_ , \new_[65905]_ , \new_[65906]_ ,
    \new_[65907]_ , \new_[65908]_ , \new_[65911]_ , \new_[65914]_ ,
    \new_[65915]_ , \new_[65918]_ , \new_[65921]_ , \new_[65922]_ ,
    \new_[65923]_ , \new_[65926]_ , \new_[65929]_ , \new_[65930]_ ,
    \new_[65933]_ , \new_[65937]_ , \new_[65938]_ , \new_[65939]_ ,
    \new_[65940]_ , \new_[65943]_ , \new_[65946]_ , \new_[65947]_ ,
    \new_[65950]_ , \new_[65953]_ , \new_[65954]_ , \new_[65955]_ ,
    \new_[65958]_ , \new_[65961]_ , \new_[65962]_ , \new_[65965]_ ,
    \new_[65969]_ , \new_[65970]_ , \new_[65971]_ , \new_[65972]_ ,
    \new_[65975]_ , \new_[65978]_ , \new_[65979]_ , \new_[65982]_ ,
    \new_[65985]_ , \new_[65986]_ , \new_[65987]_ , \new_[65990]_ ,
    \new_[65993]_ , \new_[65994]_ , \new_[65997]_ , \new_[66001]_ ,
    \new_[66002]_ , \new_[66003]_ , \new_[66004]_ , \new_[66007]_ ,
    \new_[66010]_ , \new_[66011]_ , \new_[66014]_ , \new_[66017]_ ,
    \new_[66018]_ , \new_[66019]_ , \new_[66022]_ , \new_[66025]_ ,
    \new_[66026]_ , \new_[66029]_ , \new_[66033]_ , \new_[66034]_ ,
    \new_[66035]_ , \new_[66036]_ , \new_[66039]_ , \new_[66042]_ ,
    \new_[66043]_ , \new_[66046]_ , \new_[66049]_ , \new_[66050]_ ,
    \new_[66051]_ , \new_[66054]_ , \new_[66057]_ , \new_[66058]_ ,
    \new_[66061]_ , \new_[66065]_ , \new_[66066]_ , \new_[66067]_ ,
    \new_[66068]_ , \new_[66071]_ , \new_[66074]_ , \new_[66075]_ ,
    \new_[66078]_ , \new_[66081]_ , \new_[66082]_ , \new_[66083]_ ,
    \new_[66086]_ , \new_[66089]_ , \new_[66090]_ , \new_[66093]_ ,
    \new_[66097]_ , \new_[66098]_ , \new_[66099]_ , \new_[66100]_ ,
    \new_[66103]_ , \new_[66106]_ , \new_[66107]_ , \new_[66110]_ ,
    \new_[66113]_ , \new_[66114]_ , \new_[66115]_ , \new_[66118]_ ,
    \new_[66121]_ , \new_[66122]_ , \new_[66125]_ , \new_[66129]_ ,
    \new_[66130]_ , \new_[66131]_ , \new_[66132]_ , \new_[66135]_ ,
    \new_[66138]_ , \new_[66139]_ , \new_[66142]_ , \new_[66145]_ ,
    \new_[66146]_ , \new_[66147]_ , \new_[66150]_ , \new_[66153]_ ,
    \new_[66154]_ , \new_[66157]_ , \new_[66161]_ , \new_[66162]_ ,
    \new_[66163]_ , \new_[66164]_ , \new_[66167]_ , \new_[66170]_ ,
    \new_[66171]_ , \new_[66174]_ , \new_[66177]_ , \new_[66178]_ ,
    \new_[66179]_ , \new_[66182]_ , \new_[66185]_ , \new_[66186]_ ,
    \new_[66189]_ , \new_[66193]_ , \new_[66194]_ , \new_[66195]_ ,
    \new_[66196]_ , \new_[66199]_ , \new_[66202]_ , \new_[66203]_ ,
    \new_[66206]_ , \new_[66209]_ , \new_[66210]_ , \new_[66211]_ ,
    \new_[66214]_ , \new_[66217]_ , \new_[66218]_ , \new_[66221]_ ,
    \new_[66225]_ , \new_[66226]_ , \new_[66227]_ , \new_[66228]_ ,
    \new_[66231]_ , \new_[66234]_ , \new_[66235]_ , \new_[66238]_ ,
    \new_[66241]_ , \new_[66242]_ , \new_[66243]_ , \new_[66246]_ ,
    \new_[66249]_ , \new_[66250]_ , \new_[66253]_ , \new_[66257]_ ,
    \new_[66258]_ , \new_[66259]_ , \new_[66260]_ , \new_[66263]_ ,
    \new_[66266]_ , \new_[66267]_ , \new_[66270]_ , \new_[66273]_ ,
    \new_[66274]_ , \new_[66275]_ , \new_[66278]_ , \new_[66281]_ ,
    \new_[66282]_ , \new_[66285]_ , \new_[66289]_ , \new_[66290]_ ,
    \new_[66291]_ , \new_[66292]_ , \new_[66295]_ , \new_[66298]_ ,
    \new_[66299]_ , \new_[66302]_ , \new_[66305]_ , \new_[66306]_ ,
    \new_[66307]_ , \new_[66310]_ , \new_[66313]_ , \new_[66314]_ ,
    \new_[66317]_ , \new_[66321]_ , \new_[66322]_ , \new_[66323]_ ,
    \new_[66324]_ , \new_[66327]_ , \new_[66330]_ , \new_[66331]_ ,
    \new_[66334]_ , \new_[66337]_ , \new_[66338]_ , \new_[66339]_ ,
    \new_[66342]_ , \new_[66345]_ , \new_[66346]_ , \new_[66349]_ ,
    \new_[66353]_ , \new_[66354]_ , \new_[66355]_ , \new_[66356]_ ,
    \new_[66359]_ , \new_[66362]_ , \new_[66363]_ , \new_[66366]_ ,
    \new_[66369]_ , \new_[66370]_ , \new_[66371]_ , \new_[66374]_ ,
    \new_[66377]_ , \new_[66378]_ , \new_[66381]_ , \new_[66385]_ ,
    \new_[66386]_ , \new_[66387]_ , \new_[66388]_ , \new_[66391]_ ,
    \new_[66394]_ , \new_[66395]_ , \new_[66398]_ , \new_[66401]_ ,
    \new_[66402]_ , \new_[66403]_ , \new_[66406]_ , \new_[66409]_ ,
    \new_[66410]_ , \new_[66413]_ , \new_[66417]_ , \new_[66418]_ ,
    \new_[66419]_ , \new_[66420]_ , \new_[66423]_ , \new_[66426]_ ,
    \new_[66427]_ , \new_[66430]_ , \new_[66433]_ , \new_[66434]_ ,
    \new_[66435]_ , \new_[66438]_ , \new_[66441]_ , \new_[66442]_ ,
    \new_[66445]_ , \new_[66449]_ , \new_[66450]_ , \new_[66451]_ ,
    \new_[66452]_ , \new_[66455]_ , \new_[66458]_ , \new_[66459]_ ,
    \new_[66462]_ , \new_[66465]_ , \new_[66466]_ , \new_[66467]_ ,
    \new_[66470]_ , \new_[66473]_ , \new_[66474]_ , \new_[66477]_ ,
    \new_[66481]_ , \new_[66482]_ , \new_[66483]_ , \new_[66484]_ ,
    \new_[66487]_ , \new_[66490]_ , \new_[66491]_ , \new_[66494]_ ,
    \new_[66497]_ , \new_[66498]_ , \new_[66499]_ , \new_[66502]_ ,
    \new_[66505]_ , \new_[66506]_ , \new_[66509]_ , \new_[66513]_ ,
    \new_[66514]_ , \new_[66515]_ , \new_[66516]_ , \new_[66519]_ ,
    \new_[66522]_ , \new_[66523]_ , \new_[66526]_ , \new_[66529]_ ,
    \new_[66530]_ , \new_[66531]_ , \new_[66534]_ , \new_[66537]_ ,
    \new_[66538]_ , \new_[66541]_ , \new_[66545]_ , \new_[66546]_ ,
    \new_[66547]_ , \new_[66548]_ , \new_[66551]_ , \new_[66554]_ ,
    \new_[66555]_ , \new_[66558]_ , \new_[66561]_ , \new_[66562]_ ,
    \new_[66563]_ , \new_[66566]_ , \new_[66569]_ , \new_[66570]_ ,
    \new_[66573]_ , \new_[66577]_ , \new_[66578]_ , \new_[66579]_ ,
    \new_[66580]_ , \new_[66583]_ , \new_[66586]_ , \new_[66587]_ ,
    \new_[66590]_ , \new_[66593]_ , \new_[66594]_ , \new_[66595]_ ,
    \new_[66598]_ , \new_[66601]_ , \new_[66602]_ , \new_[66605]_ ,
    \new_[66609]_ , \new_[66610]_ , \new_[66611]_ , \new_[66612]_ ,
    \new_[66615]_ , \new_[66618]_ , \new_[66619]_ , \new_[66622]_ ,
    \new_[66625]_ , \new_[66626]_ , \new_[66627]_ , \new_[66630]_ ,
    \new_[66633]_ , \new_[66634]_ , \new_[66637]_ , \new_[66641]_ ,
    \new_[66642]_ , \new_[66643]_ , \new_[66644]_ , \new_[66647]_ ,
    \new_[66650]_ , \new_[66651]_ , \new_[66654]_ , \new_[66657]_ ,
    \new_[66658]_ , \new_[66659]_ , \new_[66662]_ , \new_[66665]_ ,
    \new_[66666]_ , \new_[66669]_ , \new_[66673]_ , \new_[66674]_ ,
    \new_[66675]_ , \new_[66676]_ , \new_[66679]_ , \new_[66682]_ ,
    \new_[66683]_ , \new_[66686]_ , \new_[66689]_ , \new_[66690]_ ,
    \new_[66691]_ , \new_[66694]_ , \new_[66697]_ , \new_[66698]_ ,
    \new_[66701]_ , \new_[66705]_ , \new_[66706]_ , \new_[66707]_ ,
    \new_[66708]_ , \new_[66711]_ , \new_[66714]_ , \new_[66715]_ ,
    \new_[66718]_ , \new_[66721]_ , \new_[66722]_ , \new_[66723]_ ,
    \new_[66726]_ , \new_[66729]_ , \new_[66730]_ , \new_[66733]_ ,
    \new_[66737]_ , \new_[66738]_ , \new_[66739]_ , \new_[66740]_ ,
    \new_[66743]_ , \new_[66746]_ , \new_[66747]_ , \new_[66750]_ ,
    \new_[66753]_ , \new_[66754]_ , \new_[66755]_ , \new_[66758]_ ,
    \new_[66761]_ , \new_[66762]_ , \new_[66765]_ , \new_[66769]_ ,
    \new_[66770]_ , \new_[66771]_ , \new_[66772]_ , \new_[66775]_ ,
    \new_[66778]_ , \new_[66779]_ , \new_[66782]_ , \new_[66785]_ ,
    \new_[66786]_ , \new_[66787]_ , \new_[66790]_ , \new_[66793]_ ,
    \new_[66794]_ , \new_[66797]_ , \new_[66801]_ , \new_[66802]_ ,
    \new_[66803]_ , \new_[66804]_ , \new_[66807]_ , \new_[66810]_ ,
    \new_[66811]_ , \new_[66814]_ , \new_[66817]_ , \new_[66818]_ ,
    \new_[66819]_ , \new_[66822]_ , \new_[66825]_ , \new_[66826]_ ,
    \new_[66829]_ , \new_[66833]_ , \new_[66834]_ , \new_[66835]_ ,
    \new_[66836]_ , \new_[66839]_ , \new_[66842]_ , \new_[66843]_ ,
    \new_[66846]_ , \new_[66849]_ , \new_[66850]_ , \new_[66851]_ ,
    \new_[66854]_ , \new_[66857]_ , \new_[66858]_ , \new_[66861]_ ,
    \new_[66865]_ , \new_[66866]_ , \new_[66867]_ , \new_[66868]_ ,
    \new_[66871]_ , \new_[66874]_ , \new_[66875]_ , \new_[66878]_ ,
    \new_[66881]_ , \new_[66882]_ , \new_[66883]_ , \new_[66886]_ ,
    \new_[66889]_ , \new_[66890]_ , \new_[66893]_ , \new_[66897]_ ,
    \new_[66898]_ , \new_[66899]_ , \new_[66900]_ , \new_[66903]_ ,
    \new_[66906]_ , \new_[66907]_ , \new_[66910]_ , \new_[66913]_ ,
    \new_[66914]_ , \new_[66915]_ , \new_[66918]_ , \new_[66921]_ ,
    \new_[66922]_ , \new_[66925]_ , \new_[66929]_ , \new_[66930]_ ,
    \new_[66931]_ , \new_[66932]_ , \new_[66935]_ , \new_[66938]_ ,
    \new_[66939]_ , \new_[66942]_ , \new_[66945]_ , \new_[66946]_ ,
    \new_[66947]_ , \new_[66950]_ , \new_[66953]_ , \new_[66954]_ ,
    \new_[66957]_ , \new_[66961]_ , \new_[66962]_ , \new_[66963]_ ,
    \new_[66964]_ , \new_[66967]_ , \new_[66970]_ , \new_[66971]_ ,
    \new_[66974]_ , \new_[66977]_ , \new_[66978]_ , \new_[66979]_ ,
    \new_[66982]_ , \new_[66985]_ , \new_[66986]_ , \new_[66989]_ ,
    \new_[66993]_ , \new_[66994]_ , \new_[66995]_ , \new_[66996]_ ,
    \new_[66999]_ , \new_[67002]_ , \new_[67003]_ , \new_[67006]_ ,
    \new_[67009]_ , \new_[67010]_ , \new_[67011]_ , \new_[67014]_ ,
    \new_[67017]_ , \new_[67018]_ , \new_[67021]_ , \new_[67025]_ ,
    \new_[67026]_ , \new_[67027]_ , \new_[67028]_ , \new_[67031]_ ,
    \new_[67034]_ , \new_[67035]_ , \new_[67038]_ , \new_[67041]_ ,
    \new_[67042]_ , \new_[67043]_ , \new_[67046]_ , \new_[67049]_ ,
    \new_[67050]_ , \new_[67053]_ , \new_[67057]_ , \new_[67058]_ ,
    \new_[67059]_ , \new_[67060]_ , \new_[67063]_ , \new_[67066]_ ,
    \new_[67067]_ , \new_[67070]_ , \new_[67073]_ , \new_[67074]_ ,
    \new_[67075]_ , \new_[67078]_ , \new_[67081]_ , \new_[67082]_ ,
    \new_[67085]_ , \new_[67089]_ , \new_[67090]_ , \new_[67091]_ ,
    \new_[67092]_ , \new_[67095]_ , \new_[67098]_ , \new_[67099]_ ,
    \new_[67102]_ , \new_[67105]_ , \new_[67106]_ , \new_[67107]_ ,
    \new_[67110]_ , \new_[67113]_ , \new_[67114]_ , \new_[67117]_ ,
    \new_[67121]_ , \new_[67122]_ , \new_[67123]_ , \new_[67124]_ ,
    \new_[67127]_ , \new_[67130]_ , \new_[67131]_ , \new_[67134]_ ,
    \new_[67137]_ , \new_[67138]_ , \new_[67139]_ , \new_[67142]_ ,
    \new_[67145]_ , \new_[67146]_ , \new_[67149]_ , \new_[67153]_ ,
    \new_[67154]_ , \new_[67155]_ , \new_[67156]_ , \new_[67159]_ ,
    \new_[67162]_ , \new_[67163]_ , \new_[67166]_ , \new_[67169]_ ,
    \new_[67170]_ , \new_[67171]_ , \new_[67174]_ , \new_[67177]_ ,
    \new_[67178]_ , \new_[67181]_ , \new_[67185]_ , \new_[67186]_ ,
    \new_[67187]_ , \new_[67188]_ , \new_[67191]_ , \new_[67194]_ ,
    \new_[67195]_ , \new_[67198]_ , \new_[67201]_ , \new_[67202]_ ,
    \new_[67203]_ , \new_[67206]_ , \new_[67209]_ , \new_[67210]_ ,
    \new_[67213]_ , \new_[67217]_ , \new_[67218]_ , \new_[67219]_ ,
    \new_[67220]_ , \new_[67223]_ , \new_[67226]_ , \new_[67227]_ ,
    \new_[67230]_ , \new_[67233]_ , \new_[67234]_ , \new_[67235]_ ,
    \new_[67238]_ , \new_[67241]_ , \new_[67242]_ , \new_[67245]_ ,
    \new_[67249]_ , \new_[67250]_ , \new_[67251]_ , \new_[67252]_ ,
    \new_[67255]_ , \new_[67258]_ , \new_[67259]_ , \new_[67262]_ ,
    \new_[67265]_ , \new_[67266]_ , \new_[67267]_ , \new_[67270]_ ,
    \new_[67273]_ , \new_[67274]_ , \new_[67277]_ , \new_[67281]_ ,
    \new_[67282]_ , \new_[67283]_ , \new_[67284]_ , \new_[67287]_ ,
    \new_[67290]_ , \new_[67291]_ , \new_[67294]_ , \new_[67297]_ ,
    \new_[67298]_ , \new_[67299]_ , \new_[67302]_ , \new_[67305]_ ,
    \new_[67306]_ , \new_[67309]_ , \new_[67313]_ , \new_[67314]_ ,
    \new_[67315]_ , \new_[67316]_ , \new_[67319]_ , \new_[67322]_ ,
    \new_[67323]_ , \new_[67326]_ , \new_[67329]_ , \new_[67330]_ ,
    \new_[67331]_ , \new_[67334]_ , \new_[67337]_ , \new_[67338]_ ,
    \new_[67341]_ , \new_[67345]_ , \new_[67346]_ , \new_[67347]_ ,
    \new_[67348]_ , \new_[67351]_ , \new_[67354]_ , \new_[67355]_ ,
    \new_[67358]_ , \new_[67361]_ , \new_[67362]_ , \new_[67363]_ ,
    \new_[67366]_ , \new_[67369]_ , \new_[67370]_ , \new_[67373]_ ,
    \new_[67377]_ , \new_[67378]_ , \new_[67379]_ , \new_[67380]_ ,
    \new_[67383]_ , \new_[67386]_ , \new_[67387]_ , \new_[67390]_ ,
    \new_[67393]_ , \new_[67394]_ , \new_[67395]_ , \new_[67398]_ ,
    \new_[67401]_ , \new_[67402]_ , \new_[67405]_ , \new_[67409]_ ,
    \new_[67410]_ , \new_[67411]_ , \new_[67412]_ , \new_[67415]_ ,
    \new_[67418]_ , \new_[67419]_ , \new_[67422]_ , \new_[67425]_ ,
    \new_[67426]_ , \new_[67427]_ , \new_[67430]_ , \new_[67433]_ ,
    \new_[67434]_ , \new_[67437]_ , \new_[67441]_ , \new_[67442]_ ,
    \new_[67443]_ , \new_[67444]_ , \new_[67447]_ , \new_[67450]_ ,
    \new_[67451]_ , \new_[67454]_ , \new_[67457]_ , \new_[67458]_ ,
    \new_[67459]_ , \new_[67462]_ , \new_[67465]_ , \new_[67466]_ ,
    \new_[67469]_ , \new_[67473]_ , \new_[67474]_ , \new_[67475]_ ,
    \new_[67476]_ , \new_[67479]_ , \new_[67482]_ , \new_[67483]_ ,
    \new_[67486]_ , \new_[67489]_ , \new_[67490]_ , \new_[67491]_ ,
    \new_[67494]_ , \new_[67497]_ , \new_[67498]_ , \new_[67501]_ ,
    \new_[67505]_ , \new_[67506]_ , \new_[67507]_ , \new_[67508]_ ,
    \new_[67511]_ , \new_[67514]_ , \new_[67515]_ , \new_[67518]_ ,
    \new_[67521]_ , \new_[67522]_ , \new_[67523]_ , \new_[67526]_ ,
    \new_[67529]_ , \new_[67530]_ , \new_[67533]_ , \new_[67537]_ ,
    \new_[67538]_ , \new_[67539]_ , \new_[67540]_ , \new_[67543]_ ,
    \new_[67546]_ , \new_[67547]_ , \new_[67550]_ , \new_[67553]_ ,
    \new_[67554]_ , \new_[67555]_ , \new_[67558]_ , \new_[67561]_ ,
    \new_[67562]_ , \new_[67565]_ , \new_[67569]_ , \new_[67570]_ ,
    \new_[67571]_ , \new_[67572]_ , \new_[67575]_ , \new_[67578]_ ,
    \new_[67579]_ , \new_[67582]_ , \new_[67585]_ , \new_[67586]_ ,
    \new_[67587]_ , \new_[67590]_ , \new_[67593]_ , \new_[67594]_ ,
    \new_[67597]_ , \new_[67601]_ , \new_[67602]_ , \new_[67603]_ ,
    \new_[67604]_ , \new_[67607]_ , \new_[67610]_ , \new_[67611]_ ,
    \new_[67614]_ , \new_[67617]_ , \new_[67618]_ , \new_[67619]_ ,
    \new_[67622]_ , \new_[67625]_ , \new_[67626]_ , \new_[67629]_ ,
    \new_[67633]_ , \new_[67634]_ , \new_[67635]_ , \new_[67636]_ ,
    \new_[67639]_ , \new_[67642]_ , \new_[67643]_ , \new_[67646]_ ,
    \new_[67649]_ , \new_[67650]_ , \new_[67651]_ , \new_[67654]_ ,
    \new_[67657]_ , \new_[67658]_ , \new_[67661]_ , \new_[67665]_ ,
    \new_[67666]_ , \new_[67667]_ , \new_[67668]_ , \new_[67671]_ ,
    \new_[67674]_ , \new_[67675]_ , \new_[67678]_ , \new_[67681]_ ,
    \new_[67682]_ , \new_[67683]_ , \new_[67686]_ , \new_[67689]_ ,
    \new_[67690]_ , \new_[67693]_ , \new_[67697]_ , \new_[67698]_ ,
    \new_[67699]_ , \new_[67700]_ , \new_[67703]_ , \new_[67706]_ ,
    \new_[67707]_ , \new_[67710]_ , \new_[67714]_ , \new_[67715]_ ,
    \new_[67716]_ , \new_[67717]_ , \new_[67720]_ , \new_[67723]_ ,
    \new_[67724]_ , \new_[67727]_ , \new_[67731]_ , \new_[67732]_ ,
    \new_[67733]_ , \new_[67734]_ , \new_[67737]_ , \new_[67740]_ ,
    \new_[67741]_ , \new_[67744]_ , \new_[67748]_ , \new_[67749]_ ,
    \new_[67750]_ , \new_[67751]_ , \new_[67754]_ , \new_[67757]_ ,
    \new_[67758]_ , \new_[67761]_ , \new_[67765]_ , \new_[67766]_ ,
    \new_[67767]_ , \new_[67768]_ , \new_[67771]_ , \new_[67774]_ ,
    \new_[67775]_ , \new_[67778]_ , \new_[67782]_ , \new_[67783]_ ,
    \new_[67784]_ , \new_[67785]_ , \new_[67788]_ , \new_[67791]_ ,
    \new_[67792]_ , \new_[67795]_ , \new_[67799]_ , \new_[67800]_ ,
    \new_[67801]_ , \new_[67802]_ , \new_[67805]_ , \new_[67808]_ ,
    \new_[67809]_ , \new_[67812]_ , \new_[67816]_ , \new_[67817]_ ,
    \new_[67818]_ , \new_[67819]_ , \new_[67822]_ , \new_[67825]_ ,
    \new_[67826]_ , \new_[67829]_ , \new_[67833]_ , \new_[67834]_ ,
    \new_[67835]_ , \new_[67836]_ , \new_[67839]_ , \new_[67842]_ ,
    \new_[67843]_ , \new_[67846]_ , \new_[67850]_ , \new_[67851]_ ,
    \new_[67852]_ , \new_[67853]_ , \new_[67856]_ , \new_[67859]_ ,
    \new_[67860]_ , \new_[67863]_ , \new_[67867]_ , \new_[67868]_ ,
    \new_[67869]_ , \new_[67870]_ , \new_[67873]_ , \new_[67876]_ ,
    \new_[67877]_ , \new_[67880]_ , \new_[67884]_ , \new_[67885]_ ,
    \new_[67886]_ , \new_[67887]_ , \new_[67890]_ , \new_[67893]_ ,
    \new_[67894]_ , \new_[67897]_ , \new_[67901]_ , \new_[67902]_ ,
    \new_[67903]_ , \new_[67904]_ , \new_[67907]_ , \new_[67910]_ ,
    \new_[67911]_ , \new_[67914]_ , \new_[67918]_ , \new_[67919]_ ,
    \new_[67920]_ , \new_[67921]_ , \new_[67924]_ , \new_[67927]_ ,
    \new_[67928]_ , \new_[67931]_ , \new_[67935]_ , \new_[67936]_ ,
    \new_[67937]_ , \new_[67938]_ , \new_[67941]_ , \new_[67944]_ ,
    \new_[67945]_ , \new_[67948]_ , \new_[67952]_ , \new_[67953]_ ,
    \new_[67954]_ , \new_[67955]_ , \new_[67958]_ , \new_[67961]_ ,
    \new_[67962]_ , \new_[67965]_ , \new_[67969]_ , \new_[67970]_ ,
    \new_[67971]_ , \new_[67972]_ , \new_[67975]_ , \new_[67978]_ ,
    \new_[67979]_ , \new_[67982]_ , \new_[67986]_ , \new_[67987]_ ,
    \new_[67988]_ , \new_[67989]_ , \new_[67992]_ , \new_[67995]_ ,
    \new_[67996]_ , \new_[67999]_ , \new_[68003]_ , \new_[68004]_ ,
    \new_[68005]_ , \new_[68006]_ , \new_[68009]_ , \new_[68012]_ ,
    \new_[68013]_ , \new_[68016]_ , \new_[68020]_ , \new_[68021]_ ,
    \new_[68022]_ , \new_[68023]_ , \new_[68026]_ , \new_[68029]_ ,
    \new_[68030]_ , \new_[68033]_ , \new_[68037]_ , \new_[68038]_ ,
    \new_[68039]_ , \new_[68040]_ , \new_[68043]_ , \new_[68046]_ ,
    \new_[68047]_ , \new_[68050]_ , \new_[68054]_ , \new_[68055]_ ,
    \new_[68056]_ , \new_[68057]_ , \new_[68060]_ , \new_[68063]_ ,
    \new_[68064]_ , \new_[68067]_ , \new_[68071]_ , \new_[68072]_ ,
    \new_[68073]_ , \new_[68074]_ , \new_[68077]_ , \new_[68080]_ ,
    \new_[68081]_ , \new_[68084]_ , \new_[68088]_ , \new_[68089]_ ,
    \new_[68090]_ , \new_[68091]_ , \new_[68094]_ , \new_[68097]_ ,
    \new_[68098]_ , \new_[68101]_ , \new_[68105]_ , \new_[68106]_ ,
    \new_[68107]_ , \new_[68108]_ , \new_[68111]_ , \new_[68114]_ ,
    \new_[68115]_ , \new_[68118]_ , \new_[68122]_ , \new_[68123]_ ,
    \new_[68124]_ , \new_[68125]_ , \new_[68128]_ , \new_[68131]_ ,
    \new_[68132]_ , \new_[68135]_ , \new_[68139]_ , \new_[68140]_ ,
    \new_[68141]_ , \new_[68142]_ , \new_[68145]_ , \new_[68148]_ ,
    \new_[68149]_ , \new_[68152]_ , \new_[68156]_ , \new_[68157]_ ,
    \new_[68158]_ , \new_[68159]_ , \new_[68162]_ , \new_[68165]_ ,
    \new_[68166]_ , \new_[68169]_ , \new_[68173]_ , \new_[68174]_ ,
    \new_[68175]_ , \new_[68176]_ , \new_[68179]_ , \new_[68182]_ ,
    \new_[68183]_ , \new_[68186]_ , \new_[68190]_ , \new_[68191]_ ,
    \new_[68192]_ , \new_[68193]_ , \new_[68196]_ , \new_[68199]_ ,
    \new_[68200]_ , \new_[68203]_ , \new_[68207]_ , \new_[68208]_ ,
    \new_[68209]_ , \new_[68210]_ , \new_[68213]_ , \new_[68216]_ ,
    \new_[68217]_ , \new_[68220]_ , \new_[68224]_ , \new_[68225]_ ,
    \new_[68226]_ , \new_[68227]_ , \new_[68230]_ , \new_[68233]_ ,
    \new_[68234]_ , \new_[68237]_ , \new_[68241]_ , \new_[68242]_ ,
    \new_[68243]_ , \new_[68244]_ ;
  assign A9 = \new_[6568]_  | \new_[4379]_ ;
  assign \new_[1]_  = \new_[68244]_  & \new_[68227]_ ;
  assign \new_[2]_  = \new_[68210]_  & \new_[68193]_ ;
  assign \new_[3]_  = \new_[68176]_  & \new_[68159]_ ;
  assign \new_[4]_  = \new_[68142]_  & \new_[68125]_ ;
  assign \new_[5]_  = \new_[68108]_  & \new_[68091]_ ;
  assign \new_[6]_  = \new_[68074]_  & \new_[68057]_ ;
  assign \new_[7]_  = \new_[68040]_  & \new_[68023]_ ;
  assign \new_[8]_  = \new_[68006]_  & \new_[67989]_ ;
  assign \new_[9]_  = \new_[67972]_  & \new_[67955]_ ;
  assign \new_[10]_  = \new_[67938]_  & \new_[67921]_ ;
  assign \new_[11]_  = \new_[67904]_  & \new_[67887]_ ;
  assign \new_[12]_  = \new_[67870]_  & \new_[67853]_ ;
  assign \new_[13]_  = \new_[67836]_  & \new_[67819]_ ;
  assign \new_[14]_  = \new_[67802]_  & \new_[67785]_ ;
  assign \new_[15]_  = \new_[67768]_  & \new_[67751]_ ;
  assign \new_[16]_  = \new_[67734]_  & \new_[67717]_ ;
  assign \new_[17]_  = \new_[67700]_  & \new_[67683]_ ;
  assign \new_[18]_  = \new_[67668]_  & \new_[67651]_ ;
  assign \new_[19]_  = \new_[67636]_  & \new_[67619]_ ;
  assign \new_[20]_  = \new_[67604]_  & \new_[67587]_ ;
  assign \new_[21]_  = \new_[67572]_  & \new_[67555]_ ;
  assign \new_[22]_  = \new_[67540]_  & \new_[67523]_ ;
  assign \new_[23]_  = \new_[67508]_  & \new_[67491]_ ;
  assign \new_[24]_  = \new_[67476]_  & \new_[67459]_ ;
  assign \new_[25]_  = \new_[67444]_  & \new_[67427]_ ;
  assign \new_[26]_  = \new_[67412]_  & \new_[67395]_ ;
  assign \new_[27]_  = \new_[67380]_  & \new_[67363]_ ;
  assign \new_[28]_  = \new_[67348]_  & \new_[67331]_ ;
  assign \new_[29]_  = \new_[67316]_  & \new_[67299]_ ;
  assign \new_[30]_  = \new_[67284]_  & \new_[67267]_ ;
  assign \new_[31]_  = \new_[67252]_  & \new_[67235]_ ;
  assign \new_[32]_  = \new_[67220]_  & \new_[67203]_ ;
  assign \new_[33]_  = \new_[67188]_  & \new_[67171]_ ;
  assign \new_[34]_  = \new_[67156]_  & \new_[67139]_ ;
  assign \new_[35]_  = \new_[67124]_  & \new_[67107]_ ;
  assign \new_[36]_  = \new_[67092]_  & \new_[67075]_ ;
  assign \new_[37]_  = \new_[67060]_  & \new_[67043]_ ;
  assign \new_[38]_  = \new_[67028]_  & \new_[67011]_ ;
  assign \new_[39]_  = \new_[66996]_  & \new_[66979]_ ;
  assign \new_[40]_  = \new_[66964]_  & \new_[66947]_ ;
  assign \new_[41]_  = \new_[66932]_  & \new_[66915]_ ;
  assign \new_[42]_  = \new_[66900]_  & \new_[66883]_ ;
  assign \new_[43]_  = \new_[66868]_  & \new_[66851]_ ;
  assign \new_[44]_  = \new_[66836]_  & \new_[66819]_ ;
  assign \new_[45]_  = \new_[66804]_  & \new_[66787]_ ;
  assign \new_[46]_  = \new_[66772]_  & \new_[66755]_ ;
  assign \new_[47]_  = \new_[66740]_  & \new_[66723]_ ;
  assign \new_[48]_  = \new_[66708]_  & \new_[66691]_ ;
  assign \new_[49]_  = \new_[66676]_  & \new_[66659]_ ;
  assign \new_[50]_  = \new_[66644]_  & \new_[66627]_ ;
  assign \new_[51]_  = \new_[66612]_  & \new_[66595]_ ;
  assign \new_[52]_  = \new_[66580]_  & \new_[66563]_ ;
  assign \new_[53]_  = \new_[66548]_  & \new_[66531]_ ;
  assign \new_[54]_  = \new_[66516]_  & \new_[66499]_ ;
  assign \new_[55]_  = \new_[66484]_  & \new_[66467]_ ;
  assign \new_[56]_  = \new_[66452]_  & \new_[66435]_ ;
  assign \new_[57]_  = \new_[66420]_  & \new_[66403]_ ;
  assign \new_[58]_  = \new_[66388]_  & \new_[66371]_ ;
  assign \new_[59]_  = \new_[66356]_  & \new_[66339]_ ;
  assign \new_[60]_  = \new_[66324]_  & \new_[66307]_ ;
  assign \new_[61]_  = \new_[66292]_  & \new_[66275]_ ;
  assign \new_[62]_  = \new_[66260]_  & \new_[66243]_ ;
  assign \new_[63]_  = \new_[66228]_  & \new_[66211]_ ;
  assign \new_[64]_  = \new_[66196]_  & \new_[66179]_ ;
  assign \new_[65]_  = \new_[66164]_  & \new_[66147]_ ;
  assign \new_[66]_  = \new_[66132]_  & \new_[66115]_ ;
  assign \new_[67]_  = \new_[66100]_  & \new_[66083]_ ;
  assign \new_[68]_  = \new_[66068]_  & \new_[66051]_ ;
  assign \new_[69]_  = \new_[66036]_  & \new_[66019]_ ;
  assign \new_[70]_  = \new_[66004]_  & \new_[65987]_ ;
  assign \new_[71]_  = \new_[65972]_  & \new_[65955]_ ;
  assign \new_[72]_  = \new_[65940]_  & \new_[65923]_ ;
  assign \new_[73]_  = \new_[65908]_  & \new_[65891]_ ;
  assign \new_[74]_  = \new_[65876]_  & \new_[65859]_ ;
  assign \new_[75]_  = \new_[65844]_  & \new_[65827]_ ;
  assign \new_[76]_  = \new_[65812]_  & \new_[65795]_ ;
  assign \new_[77]_  = \new_[65780]_  & \new_[65763]_ ;
  assign \new_[78]_  = \new_[65748]_  & \new_[65731]_ ;
  assign \new_[79]_  = \new_[65716]_  & \new_[65699]_ ;
  assign \new_[80]_  = \new_[65684]_  & \new_[65667]_ ;
  assign \new_[81]_  = \new_[65652]_  & \new_[65635]_ ;
  assign \new_[82]_  = \new_[65620]_  & \new_[65603]_ ;
  assign \new_[83]_  = \new_[65588]_  & \new_[65571]_ ;
  assign \new_[84]_  = \new_[65556]_  & \new_[65539]_ ;
  assign \new_[85]_  = \new_[65524]_  & \new_[65507]_ ;
  assign \new_[86]_  = \new_[65492]_  & \new_[65475]_ ;
  assign \new_[87]_  = \new_[65460]_  & \new_[65443]_ ;
  assign \new_[88]_  = \new_[65428]_  & \new_[65411]_ ;
  assign \new_[89]_  = \new_[65396]_  & \new_[65379]_ ;
  assign \new_[90]_  = \new_[65364]_  & \new_[65347]_ ;
  assign \new_[91]_  = \new_[65332]_  & \new_[65315]_ ;
  assign \new_[92]_  = \new_[65300]_  & \new_[65283]_ ;
  assign \new_[93]_  = \new_[65268]_  & \new_[65251]_ ;
  assign \new_[94]_  = \new_[65236]_  & \new_[65219]_ ;
  assign \new_[95]_  = \new_[65204]_  & \new_[65187]_ ;
  assign \new_[96]_  = \new_[65172]_  & \new_[65155]_ ;
  assign \new_[97]_  = \new_[65140]_  & \new_[65123]_ ;
  assign \new_[98]_  = \new_[65108]_  & \new_[65091]_ ;
  assign \new_[99]_  = \new_[65076]_  & \new_[65059]_ ;
  assign \new_[100]_  = \new_[65044]_  & \new_[65027]_ ;
  assign \new_[101]_  = \new_[65012]_  & \new_[64995]_ ;
  assign \new_[102]_  = \new_[64980]_  & \new_[64963]_ ;
  assign \new_[103]_  = \new_[64948]_  & \new_[64931]_ ;
  assign \new_[104]_  = \new_[64916]_  & \new_[64899]_ ;
  assign \new_[105]_  = \new_[64884]_  & \new_[64867]_ ;
  assign \new_[106]_  = \new_[64852]_  & \new_[64835]_ ;
  assign \new_[107]_  = \new_[64820]_  & \new_[64803]_ ;
  assign \new_[108]_  = \new_[64788]_  & \new_[64771]_ ;
  assign \new_[109]_  = \new_[64756]_  & \new_[64739]_ ;
  assign \new_[110]_  = \new_[64724]_  & \new_[64707]_ ;
  assign \new_[111]_  = \new_[64692]_  & \new_[64675]_ ;
  assign \new_[112]_  = \new_[64660]_  & \new_[64643]_ ;
  assign \new_[113]_  = \new_[64628]_  & \new_[64611]_ ;
  assign \new_[114]_  = \new_[64596]_  & \new_[64579]_ ;
  assign \new_[115]_  = \new_[64564]_  & \new_[64547]_ ;
  assign \new_[116]_  = \new_[64532]_  & \new_[64515]_ ;
  assign \new_[117]_  = \new_[64500]_  & \new_[64483]_ ;
  assign \new_[118]_  = \new_[64468]_  & \new_[64451]_ ;
  assign \new_[119]_  = \new_[64436]_  & \new_[64419]_ ;
  assign \new_[120]_  = \new_[64404]_  & \new_[64387]_ ;
  assign \new_[121]_  = \new_[64372]_  & \new_[64355]_ ;
  assign \new_[122]_  = \new_[64340]_  & \new_[64323]_ ;
  assign \new_[123]_  = \new_[64308]_  & \new_[64291]_ ;
  assign \new_[124]_  = \new_[64276]_  & \new_[64259]_ ;
  assign \new_[125]_  = \new_[64244]_  & \new_[64227]_ ;
  assign \new_[126]_  = \new_[64212]_  & \new_[64195]_ ;
  assign \new_[127]_  = \new_[64180]_  & \new_[64163]_ ;
  assign \new_[128]_  = \new_[64148]_  & \new_[64131]_ ;
  assign \new_[129]_  = \new_[64116]_  & \new_[64099]_ ;
  assign \new_[130]_  = \new_[64084]_  & \new_[64067]_ ;
  assign \new_[131]_  = \new_[64052]_  & \new_[64035]_ ;
  assign \new_[132]_  = \new_[64020]_  & \new_[64003]_ ;
  assign \new_[133]_  = \new_[63988]_  & \new_[63971]_ ;
  assign \new_[134]_  = \new_[63956]_  & \new_[63939]_ ;
  assign \new_[135]_  = \new_[63924]_  & \new_[63907]_ ;
  assign \new_[136]_  = \new_[63892]_  & \new_[63875]_ ;
  assign \new_[137]_  = \new_[63860]_  & \new_[63843]_ ;
  assign \new_[138]_  = \new_[63828]_  & \new_[63811]_ ;
  assign \new_[139]_  = \new_[63796]_  & \new_[63779]_ ;
  assign \new_[140]_  = \new_[63764]_  & \new_[63747]_ ;
  assign \new_[141]_  = \new_[63732]_  & \new_[63715]_ ;
  assign \new_[142]_  = \new_[63700]_  & \new_[63683]_ ;
  assign \new_[143]_  = \new_[63668]_  & \new_[63651]_ ;
  assign \new_[144]_  = \new_[63636]_  & \new_[63619]_ ;
  assign \new_[145]_  = \new_[63604]_  & \new_[63587]_ ;
  assign \new_[146]_  = \new_[63572]_  & \new_[63555]_ ;
  assign \new_[147]_  = \new_[63540]_  & \new_[63523]_ ;
  assign \new_[148]_  = \new_[63508]_  & \new_[63491]_ ;
  assign \new_[149]_  = \new_[63476]_  & \new_[63459]_ ;
  assign \new_[150]_  = \new_[63444]_  & \new_[63427]_ ;
  assign \new_[151]_  = \new_[63412]_  & \new_[63395]_ ;
  assign \new_[152]_  = \new_[63380]_  & \new_[63363]_ ;
  assign \new_[153]_  = \new_[63348]_  & \new_[63331]_ ;
  assign \new_[154]_  = \new_[63316]_  & \new_[63299]_ ;
  assign \new_[155]_  = \new_[63284]_  & \new_[63267]_ ;
  assign \new_[156]_  = \new_[63252]_  & \new_[63235]_ ;
  assign \new_[157]_  = \new_[63220]_  & \new_[63203]_ ;
  assign \new_[158]_  = \new_[63188]_  & \new_[63171]_ ;
  assign \new_[159]_  = \new_[63156]_  & \new_[63139]_ ;
  assign \new_[160]_  = \new_[63124]_  & \new_[63107]_ ;
  assign \new_[161]_  = \new_[63092]_  & \new_[63075]_ ;
  assign \new_[162]_  = \new_[63060]_  & \new_[63043]_ ;
  assign \new_[163]_  = \new_[63028]_  & \new_[63011]_ ;
  assign \new_[164]_  = \new_[62996]_  & \new_[62979]_ ;
  assign \new_[165]_  = \new_[62964]_  & \new_[62947]_ ;
  assign \new_[166]_  = \new_[62932]_  & \new_[62915]_ ;
  assign \new_[167]_  = \new_[62900]_  & \new_[62883]_ ;
  assign \new_[168]_  = \new_[62868]_  & \new_[62851]_ ;
  assign \new_[169]_  = \new_[62836]_  & \new_[62819]_ ;
  assign \new_[170]_  = \new_[62804]_  & \new_[62787]_ ;
  assign \new_[171]_  = \new_[62772]_  & \new_[62755]_ ;
  assign \new_[172]_  = \new_[62740]_  & \new_[62723]_ ;
  assign \new_[173]_  = \new_[62708]_  & \new_[62691]_ ;
  assign \new_[174]_  = \new_[62676]_  & \new_[62659]_ ;
  assign \new_[175]_  = \new_[62644]_  & \new_[62627]_ ;
  assign \new_[176]_  = \new_[62612]_  & \new_[62595]_ ;
  assign \new_[177]_  = \new_[62580]_  & \new_[62565]_ ;
  assign \new_[178]_  = \new_[62550]_  & \new_[62535]_ ;
  assign \new_[179]_  = \new_[62520]_  & \new_[62505]_ ;
  assign \new_[180]_  = \new_[62490]_  & \new_[62475]_ ;
  assign \new_[181]_  = \new_[62460]_  & \new_[62445]_ ;
  assign \new_[182]_  = \new_[62430]_  & \new_[62415]_ ;
  assign \new_[183]_  = \new_[62400]_  & \new_[62385]_ ;
  assign \new_[184]_  = \new_[62370]_  & \new_[62355]_ ;
  assign \new_[185]_  = \new_[62340]_  & \new_[62325]_ ;
  assign \new_[186]_  = \new_[62310]_  & \new_[62295]_ ;
  assign \new_[187]_  = \new_[62280]_  & \new_[62265]_ ;
  assign \new_[188]_  = \new_[62250]_  & \new_[62235]_ ;
  assign \new_[189]_  = \new_[62220]_  & \new_[62205]_ ;
  assign \new_[190]_  = \new_[62190]_  & \new_[62175]_ ;
  assign \new_[191]_  = \new_[62160]_  & \new_[62145]_ ;
  assign \new_[192]_  = \new_[62130]_  & \new_[62115]_ ;
  assign \new_[193]_  = \new_[62100]_  & \new_[62085]_ ;
  assign \new_[194]_  = \new_[62070]_  & \new_[62055]_ ;
  assign \new_[195]_  = \new_[62040]_  & \new_[62025]_ ;
  assign \new_[196]_  = \new_[62010]_  & \new_[61995]_ ;
  assign \new_[197]_  = \new_[61980]_  & \new_[61965]_ ;
  assign \new_[198]_  = \new_[61950]_  & \new_[61935]_ ;
  assign \new_[199]_  = \new_[61920]_  & \new_[61905]_ ;
  assign \new_[200]_  = \new_[61890]_  & \new_[61875]_ ;
  assign \new_[201]_  = \new_[61860]_  & \new_[61845]_ ;
  assign \new_[202]_  = \new_[61830]_  & \new_[61815]_ ;
  assign \new_[203]_  = \new_[61800]_  & \new_[61785]_ ;
  assign \new_[204]_  = \new_[61770]_  & \new_[61755]_ ;
  assign \new_[205]_  = \new_[61740]_  & \new_[61725]_ ;
  assign \new_[206]_  = \new_[61710]_  & \new_[61695]_ ;
  assign \new_[207]_  = \new_[61680]_  & \new_[61665]_ ;
  assign \new_[208]_  = \new_[61650]_  & \new_[61635]_ ;
  assign \new_[209]_  = \new_[61620]_  & \new_[61605]_ ;
  assign \new_[210]_  = \new_[61590]_  & \new_[61575]_ ;
  assign \new_[211]_  = \new_[61560]_  & \new_[61545]_ ;
  assign \new_[212]_  = \new_[61530]_  & \new_[61515]_ ;
  assign \new_[213]_  = \new_[61500]_  & \new_[61485]_ ;
  assign \new_[214]_  = \new_[61470]_  & \new_[61455]_ ;
  assign \new_[215]_  = \new_[61440]_  & \new_[61425]_ ;
  assign \new_[216]_  = \new_[61410]_  & \new_[61395]_ ;
  assign \new_[217]_  = \new_[61380]_  & \new_[61365]_ ;
  assign \new_[218]_  = \new_[61350]_  & \new_[61335]_ ;
  assign \new_[219]_  = \new_[61320]_  & \new_[61305]_ ;
  assign \new_[220]_  = \new_[61290]_  & \new_[61275]_ ;
  assign \new_[221]_  = \new_[61260]_  & \new_[61245]_ ;
  assign \new_[222]_  = \new_[61230]_  & \new_[61215]_ ;
  assign \new_[223]_  = \new_[61200]_  & \new_[61185]_ ;
  assign \new_[224]_  = \new_[61170]_  & \new_[61155]_ ;
  assign \new_[225]_  = \new_[61140]_  & \new_[61125]_ ;
  assign \new_[226]_  = \new_[61110]_  & \new_[61095]_ ;
  assign \new_[227]_  = \new_[61080]_  & \new_[61065]_ ;
  assign \new_[228]_  = \new_[61050]_  & \new_[61035]_ ;
  assign \new_[229]_  = \new_[61020]_  & \new_[61005]_ ;
  assign \new_[230]_  = \new_[60990]_  & \new_[60975]_ ;
  assign \new_[231]_  = \new_[60960]_  & \new_[60945]_ ;
  assign \new_[232]_  = \new_[60930]_  & \new_[60915]_ ;
  assign \new_[233]_  = \new_[60900]_  & \new_[60885]_ ;
  assign \new_[234]_  = \new_[60870]_  & \new_[60855]_ ;
  assign \new_[235]_  = \new_[60840]_  & \new_[60825]_ ;
  assign \new_[236]_  = \new_[60810]_  & \new_[60795]_ ;
  assign \new_[237]_  = \new_[60780]_  & \new_[60765]_ ;
  assign \new_[238]_  = \new_[60750]_  & \new_[60735]_ ;
  assign \new_[239]_  = \new_[60720]_  & \new_[60705]_ ;
  assign \new_[240]_  = \new_[60690]_  & \new_[60675]_ ;
  assign \new_[241]_  = \new_[60660]_  & \new_[60645]_ ;
  assign \new_[242]_  = \new_[60630]_  & \new_[60615]_ ;
  assign \new_[243]_  = \new_[60600]_  & \new_[60585]_ ;
  assign \new_[244]_  = \new_[60570]_  & \new_[60555]_ ;
  assign \new_[245]_  = \new_[60540]_  & \new_[60525]_ ;
  assign \new_[246]_  = \new_[60510]_  & \new_[60495]_ ;
  assign \new_[247]_  = \new_[60480]_  & \new_[60465]_ ;
  assign \new_[248]_  = \new_[60450]_  & \new_[60435]_ ;
  assign \new_[249]_  = \new_[60420]_  & \new_[60405]_ ;
  assign \new_[250]_  = \new_[60390]_  & \new_[60375]_ ;
  assign \new_[251]_  = \new_[60360]_  & \new_[60345]_ ;
  assign \new_[252]_  = \new_[60330]_  & \new_[60315]_ ;
  assign \new_[253]_  = \new_[60300]_  & \new_[60285]_ ;
  assign \new_[254]_  = \new_[60270]_  & \new_[60255]_ ;
  assign \new_[255]_  = \new_[60240]_  & \new_[60225]_ ;
  assign \new_[256]_  = \new_[60210]_  & \new_[60195]_ ;
  assign \new_[257]_  = \new_[60180]_  & \new_[60165]_ ;
  assign \new_[258]_  = \new_[60150]_  & \new_[60135]_ ;
  assign \new_[259]_  = \new_[60120]_  & \new_[60105]_ ;
  assign \new_[260]_  = \new_[60090]_  & \new_[60075]_ ;
  assign \new_[261]_  = \new_[60060]_  & \new_[60045]_ ;
  assign \new_[262]_  = \new_[60030]_  & \new_[60015]_ ;
  assign \new_[263]_  = \new_[60000]_  & \new_[59985]_ ;
  assign \new_[264]_  = \new_[59970]_  & \new_[59955]_ ;
  assign \new_[265]_  = \new_[59940]_  & \new_[59925]_ ;
  assign \new_[266]_  = \new_[59910]_  & \new_[59895]_ ;
  assign \new_[267]_  = \new_[59880]_  & \new_[59865]_ ;
  assign \new_[268]_  = \new_[59850]_  & \new_[59835]_ ;
  assign \new_[269]_  = \new_[59820]_  & \new_[59805]_ ;
  assign \new_[270]_  = \new_[59790]_  & \new_[59775]_ ;
  assign \new_[271]_  = \new_[59760]_  & \new_[59745]_ ;
  assign \new_[272]_  = \new_[59730]_  & \new_[59715]_ ;
  assign \new_[273]_  = \new_[59700]_  & \new_[59685]_ ;
  assign \new_[274]_  = \new_[59670]_  & \new_[59655]_ ;
  assign \new_[275]_  = \new_[59640]_  & \new_[59625]_ ;
  assign \new_[276]_  = \new_[59610]_  & \new_[59595]_ ;
  assign \new_[277]_  = \new_[59580]_  & \new_[59565]_ ;
  assign \new_[278]_  = \new_[59550]_  & \new_[59535]_ ;
  assign \new_[279]_  = \new_[59520]_  & \new_[59505]_ ;
  assign \new_[280]_  = \new_[59490]_  & \new_[59475]_ ;
  assign \new_[281]_  = \new_[59460]_  & \new_[59445]_ ;
  assign \new_[282]_  = \new_[59430]_  & \new_[59415]_ ;
  assign \new_[283]_  = \new_[59400]_  & \new_[59385]_ ;
  assign \new_[284]_  = \new_[59370]_  & \new_[59355]_ ;
  assign \new_[285]_  = \new_[59340]_  & \new_[59325]_ ;
  assign \new_[286]_  = \new_[59310]_  & \new_[59295]_ ;
  assign \new_[287]_  = \new_[59280]_  & \new_[59265]_ ;
  assign \new_[288]_  = \new_[59250]_  & \new_[59235]_ ;
  assign \new_[289]_  = \new_[59220]_  & \new_[59205]_ ;
  assign \new_[290]_  = \new_[59190]_  & \new_[59175]_ ;
  assign \new_[291]_  = \new_[59160]_  & \new_[59145]_ ;
  assign \new_[292]_  = \new_[59130]_  & \new_[59115]_ ;
  assign \new_[293]_  = \new_[59100]_  & \new_[59085]_ ;
  assign \new_[294]_  = \new_[59070]_  & \new_[59055]_ ;
  assign \new_[295]_  = \new_[59040]_  & \new_[59025]_ ;
  assign \new_[296]_  = \new_[59010]_  & \new_[58995]_ ;
  assign \new_[297]_  = \new_[58980]_  & \new_[58965]_ ;
  assign \new_[298]_  = \new_[58950]_  & \new_[58935]_ ;
  assign \new_[299]_  = \new_[58920]_  & \new_[58905]_ ;
  assign \new_[300]_  = \new_[58890]_  & \new_[58875]_ ;
  assign \new_[301]_  = \new_[58860]_  & \new_[58845]_ ;
  assign \new_[302]_  = \new_[58830]_  & \new_[58815]_ ;
  assign \new_[303]_  = \new_[58800]_  & \new_[58785]_ ;
  assign \new_[304]_  = \new_[58770]_  & \new_[58755]_ ;
  assign \new_[305]_  = \new_[58740]_  & \new_[58725]_ ;
  assign \new_[306]_  = \new_[58710]_  & \new_[58695]_ ;
  assign \new_[307]_  = \new_[58680]_  & \new_[58665]_ ;
  assign \new_[308]_  = \new_[58650]_  & \new_[58635]_ ;
  assign \new_[309]_  = \new_[58620]_  & \new_[58605]_ ;
  assign \new_[310]_  = \new_[58590]_  & \new_[58575]_ ;
  assign \new_[311]_  = \new_[58560]_  & \new_[58545]_ ;
  assign \new_[312]_  = \new_[58530]_  & \new_[58515]_ ;
  assign \new_[313]_  = \new_[58500]_  & \new_[58485]_ ;
  assign \new_[314]_  = \new_[58470]_  & \new_[58455]_ ;
  assign \new_[315]_  = \new_[58440]_  & \new_[58425]_ ;
  assign \new_[316]_  = \new_[58410]_  & \new_[58395]_ ;
  assign \new_[317]_  = \new_[58380]_  & \new_[58365]_ ;
  assign \new_[318]_  = \new_[58350]_  & \new_[58335]_ ;
  assign \new_[319]_  = \new_[58320]_  & \new_[58305]_ ;
  assign \new_[320]_  = \new_[58290]_  & \new_[58275]_ ;
  assign \new_[321]_  = \new_[58260]_  & \new_[58245]_ ;
  assign \new_[322]_  = \new_[58230]_  & \new_[58215]_ ;
  assign \new_[323]_  = \new_[58200]_  & \new_[58185]_ ;
  assign \new_[324]_  = \new_[58170]_  & \new_[58155]_ ;
  assign \new_[325]_  = \new_[58140]_  & \new_[58125]_ ;
  assign \new_[326]_  = \new_[58110]_  & \new_[58095]_ ;
  assign \new_[327]_  = \new_[58080]_  & \new_[58065]_ ;
  assign \new_[328]_  = \new_[58050]_  & \new_[58035]_ ;
  assign \new_[329]_  = \new_[58020]_  & \new_[58005]_ ;
  assign \new_[330]_  = \new_[57990]_  & \new_[57975]_ ;
  assign \new_[331]_  = \new_[57960]_  & \new_[57945]_ ;
  assign \new_[332]_  = \new_[57930]_  & \new_[57915]_ ;
  assign \new_[333]_  = \new_[57900]_  & \new_[57885]_ ;
  assign \new_[334]_  = \new_[57870]_  & \new_[57855]_ ;
  assign \new_[335]_  = \new_[57840]_  & \new_[57825]_ ;
  assign \new_[336]_  = \new_[57810]_  & \new_[57795]_ ;
  assign \new_[337]_  = \new_[57780]_  & \new_[57765]_ ;
  assign \new_[338]_  = \new_[57750]_  & \new_[57735]_ ;
  assign \new_[339]_  = \new_[57720]_  & \new_[57705]_ ;
  assign \new_[340]_  = \new_[57690]_  & \new_[57675]_ ;
  assign \new_[341]_  = \new_[57660]_  & \new_[57645]_ ;
  assign \new_[342]_  = \new_[57630]_  & \new_[57615]_ ;
  assign \new_[343]_  = \new_[57600]_  & \new_[57585]_ ;
  assign \new_[344]_  = \new_[57570]_  & \new_[57555]_ ;
  assign \new_[345]_  = \new_[57540]_  & \new_[57525]_ ;
  assign \new_[346]_  = \new_[57510]_  & \new_[57495]_ ;
  assign \new_[347]_  = \new_[57480]_  & \new_[57465]_ ;
  assign \new_[348]_  = \new_[57450]_  & \new_[57435]_ ;
  assign \new_[349]_  = \new_[57420]_  & \new_[57405]_ ;
  assign \new_[350]_  = \new_[57390]_  & \new_[57375]_ ;
  assign \new_[351]_  = \new_[57360]_  & \new_[57345]_ ;
  assign \new_[352]_  = \new_[57330]_  & \new_[57315]_ ;
  assign \new_[353]_  = \new_[57300]_  & \new_[57285]_ ;
  assign \new_[354]_  = \new_[57270]_  & \new_[57255]_ ;
  assign \new_[355]_  = \new_[57240]_  & \new_[57225]_ ;
  assign \new_[356]_  = \new_[57210]_  & \new_[57195]_ ;
  assign \new_[357]_  = \new_[57180]_  & \new_[57165]_ ;
  assign \new_[358]_  = \new_[57150]_  & \new_[57135]_ ;
  assign \new_[359]_  = \new_[57120]_  & \new_[57105]_ ;
  assign \new_[360]_  = \new_[57090]_  & \new_[57075]_ ;
  assign \new_[361]_  = \new_[57060]_  & \new_[57045]_ ;
  assign \new_[362]_  = \new_[57030]_  & \new_[57015]_ ;
  assign \new_[363]_  = \new_[57000]_  & \new_[56985]_ ;
  assign \new_[364]_  = \new_[56970]_  & \new_[56955]_ ;
  assign \new_[365]_  = \new_[56940]_  & \new_[56925]_ ;
  assign \new_[366]_  = \new_[56910]_  & \new_[56895]_ ;
  assign \new_[367]_  = \new_[56880]_  & \new_[56865]_ ;
  assign \new_[368]_  = \new_[56850]_  & \new_[56835]_ ;
  assign \new_[369]_  = \new_[56820]_  & \new_[56805]_ ;
  assign \new_[370]_  = \new_[56790]_  & \new_[56775]_ ;
  assign \new_[371]_  = \new_[56760]_  & \new_[56745]_ ;
  assign \new_[372]_  = \new_[56730]_  & \new_[56715]_ ;
  assign \new_[373]_  = \new_[56700]_  & \new_[56685]_ ;
  assign \new_[374]_  = \new_[56670]_  & \new_[56655]_ ;
  assign \new_[375]_  = \new_[56640]_  & \new_[56625]_ ;
  assign \new_[376]_  = \new_[56610]_  & \new_[56595]_ ;
  assign \new_[377]_  = \new_[56580]_  & \new_[56565]_ ;
  assign \new_[378]_  = \new_[56550]_  & \new_[56535]_ ;
  assign \new_[379]_  = \new_[56520]_  & \new_[56505]_ ;
  assign \new_[380]_  = \new_[56490]_  & \new_[56475]_ ;
  assign \new_[381]_  = \new_[56460]_  & \new_[56445]_ ;
  assign \new_[382]_  = \new_[56430]_  & \new_[56415]_ ;
  assign \new_[383]_  = \new_[56400]_  & \new_[56385]_ ;
  assign \new_[384]_  = \new_[56370]_  & \new_[56355]_ ;
  assign \new_[385]_  = \new_[56340]_  & \new_[56325]_ ;
  assign \new_[386]_  = \new_[56310]_  & \new_[56295]_ ;
  assign \new_[387]_  = \new_[56280]_  & \new_[56265]_ ;
  assign \new_[388]_  = \new_[56250]_  & \new_[56235]_ ;
  assign \new_[389]_  = \new_[56220]_  & \new_[56205]_ ;
  assign \new_[390]_  = \new_[56190]_  & \new_[56175]_ ;
  assign \new_[391]_  = \new_[56160]_  & \new_[56145]_ ;
  assign \new_[392]_  = \new_[56130]_  & \new_[56115]_ ;
  assign \new_[393]_  = \new_[56100]_  & \new_[56085]_ ;
  assign \new_[394]_  = \new_[56070]_  & \new_[56055]_ ;
  assign \new_[395]_  = \new_[56040]_  & \new_[56025]_ ;
  assign \new_[396]_  = \new_[56010]_  & \new_[55995]_ ;
  assign \new_[397]_  = \new_[55980]_  & \new_[55965]_ ;
  assign \new_[398]_  = \new_[55950]_  & \new_[55935]_ ;
  assign \new_[399]_  = \new_[55920]_  & \new_[55905]_ ;
  assign \new_[400]_  = \new_[55890]_  & \new_[55875]_ ;
  assign \new_[401]_  = \new_[55860]_  & \new_[55845]_ ;
  assign \new_[402]_  = \new_[55830]_  & \new_[55815]_ ;
  assign \new_[403]_  = \new_[55800]_  & \new_[55785]_ ;
  assign \new_[404]_  = \new_[55770]_  & \new_[55755]_ ;
  assign \new_[405]_  = \new_[55740]_  & \new_[55725]_ ;
  assign \new_[406]_  = \new_[55710]_  & \new_[55695]_ ;
  assign \new_[407]_  = \new_[55680]_  & \new_[55665]_ ;
  assign \new_[408]_  = \new_[55650]_  & \new_[55635]_ ;
  assign \new_[409]_  = \new_[55620]_  & \new_[55605]_ ;
  assign \new_[410]_  = \new_[55590]_  & \new_[55575]_ ;
  assign \new_[411]_  = \new_[55560]_  & \new_[55545]_ ;
  assign \new_[412]_  = \new_[55530]_  & \new_[55515]_ ;
  assign \new_[413]_  = \new_[55500]_  & \new_[55485]_ ;
  assign \new_[414]_  = \new_[55470]_  & \new_[55455]_ ;
  assign \new_[415]_  = \new_[55440]_  & \new_[55425]_ ;
  assign \new_[416]_  = \new_[55410]_  & \new_[55395]_ ;
  assign \new_[417]_  = \new_[55380]_  & \new_[55365]_ ;
  assign \new_[418]_  = \new_[55350]_  & \new_[55335]_ ;
  assign \new_[419]_  = \new_[55320]_  & \new_[55305]_ ;
  assign \new_[420]_  = \new_[55290]_  & \new_[55275]_ ;
  assign \new_[421]_  = \new_[55260]_  & \new_[55245]_ ;
  assign \new_[422]_  = \new_[55230]_  & \new_[55215]_ ;
  assign \new_[423]_  = \new_[55200]_  & \new_[55185]_ ;
  assign \new_[424]_  = \new_[55170]_  & \new_[55155]_ ;
  assign \new_[425]_  = \new_[55140]_  & \new_[55125]_ ;
  assign \new_[426]_  = \new_[55110]_  & \new_[55095]_ ;
  assign \new_[427]_  = \new_[55080]_  & \new_[55065]_ ;
  assign \new_[428]_  = \new_[55050]_  & \new_[55035]_ ;
  assign \new_[429]_  = \new_[55020]_  & \new_[55005]_ ;
  assign \new_[430]_  = \new_[54990]_  & \new_[54975]_ ;
  assign \new_[431]_  = \new_[54960]_  & \new_[54945]_ ;
  assign \new_[432]_  = \new_[54930]_  & \new_[54915]_ ;
  assign \new_[433]_  = \new_[54900]_  & \new_[54885]_ ;
  assign \new_[434]_  = \new_[54870]_  & \new_[54855]_ ;
  assign \new_[435]_  = \new_[54840]_  & \new_[54825]_ ;
  assign \new_[436]_  = \new_[54810]_  & \new_[54795]_ ;
  assign \new_[437]_  = \new_[54780]_  & \new_[54765]_ ;
  assign \new_[438]_  = \new_[54750]_  & \new_[54735]_ ;
  assign \new_[439]_  = \new_[54720]_  & \new_[54705]_ ;
  assign \new_[440]_  = \new_[54690]_  & \new_[54675]_ ;
  assign \new_[441]_  = \new_[54660]_  & \new_[54645]_ ;
  assign \new_[442]_  = \new_[54630]_  & \new_[54615]_ ;
  assign \new_[443]_  = \new_[54600]_  & \new_[54585]_ ;
  assign \new_[444]_  = \new_[54570]_  & \new_[54555]_ ;
  assign \new_[445]_  = \new_[54540]_  & \new_[54525]_ ;
  assign \new_[446]_  = \new_[54510]_  & \new_[54495]_ ;
  assign \new_[447]_  = \new_[54480]_  & \new_[54465]_ ;
  assign \new_[448]_  = \new_[54450]_  & \new_[54435]_ ;
  assign \new_[449]_  = \new_[54420]_  & \new_[54405]_ ;
  assign \new_[450]_  = \new_[54390]_  & \new_[54375]_ ;
  assign \new_[451]_  = \new_[54360]_  & \new_[54345]_ ;
  assign \new_[452]_  = \new_[54330]_  & \new_[54315]_ ;
  assign \new_[453]_  = \new_[54300]_  & \new_[54285]_ ;
  assign \new_[454]_  = \new_[54270]_  & \new_[54255]_ ;
  assign \new_[455]_  = \new_[54240]_  & \new_[54225]_ ;
  assign \new_[456]_  = \new_[54210]_  & \new_[54195]_ ;
  assign \new_[457]_  = \new_[54180]_  & \new_[54165]_ ;
  assign \new_[458]_  = \new_[54150]_  & \new_[54135]_ ;
  assign \new_[459]_  = \new_[54120]_  & \new_[54105]_ ;
  assign \new_[460]_  = \new_[54090]_  & \new_[54075]_ ;
  assign \new_[461]_  = \new_[54060]_  & \new_[54045]_ ;
  assign \new_[462]_  = \new_[54030]_  & \new_[54015]_ ;
  assign \new_[463]_  = \new_[54000]_  & \new_[53985]_ ;
  assign \new_[464]_  = \new_[53970]_  & \new_[53955]_ ;
  assign \new_[465]_  = \new_[53940]_  & \new_[53925]_ ;
  assign \new_[466]_  = \new_[53910]_  & \new_[53895]_ ;
  assign \new_[467]_  = \new_[53880]_  & \new_[53865]_ ;
  assign \new_[468]_  = \new_[53850]_  & \new_[53835]_ ;
  assign \new_[469]_  = \new_[53820]_  & \new_[53805]_ ;
  assign \new_[470]_  = \new_[53790]_  & \new_[53775]_ ;
  assign \new_[471]_  = \new_[53760]_  & \new_[53745]_ ;
  assign \new_[472]_  = \new_[53730]_  & \new_[53715]_ ;
  assign \new_[473]_  = \new_[53700]_  & \new_[53685]_ ;
  assign \new_[474]_  = \new_[53670]_  & \new_[53655]_ ;
  assign \new_[475]_  = \new_[53640]_  & \new_[53625]_ ;
  assign \new_[476]_  = \new_[53610]_  & \new_[53595]_ ;
  assign \new_[477]_  = \new_[53580]_  & \new_[53565]_ ;
  assign \new_[478]_  = \new_[53550]_  & \new_[53535]_ ;
  assign \new_[479]_  = \new_[53520]_  & \new_[53505]_ ;
  assign \new_[480]_  = \new_[53490]_  & \new_[53475]_ ;
  assign \new_[481]_  = \new_[53460]_  & \new_[53445]_ ;
  assign \new_[482]_  = \new_[53430]_  & \new_[53415]_ ;
  assign \new_[483]_  = \new_[53400]_  & \new_[53385]_ ;
  assign \new_[484]_  = \new_[53370]_  & \new_[53355]_ ;
  assign \new_[485]_  = \new_[53340]_  & \new_[53325]_ ;
  assign \new_[486]_  = \new_[53310]_  & \new_[53295]_ ;
  assign \new_[487]_  = \new_[53280]_  & \new_[53265]_ ;
  assign \new_[488]_  = \new_[53250]_  & \new_[53235]_ ;
  assign \new_[489]_  = \new_[53220]_  & \new_[53205]_ ;
  assign \new_[490]_  = \new_[53190]_  & \new_[53175]_ ;
  assign \new_[491]_  = \new_[53160]_  & \new_[53145]_ ;
  assign \new_[492]_  = \new_[53130]_  & \new_[53115]_ ;
  assign \new_[493]_  = \new_[53100]_  & \new_[53085]_ ;
  assign \new_[494]_  = \new_[53070]_  & \new_[53055]_ ;
  assign \new_[495]_  = \new_[53040]_  & \new_[53025]_ ;
  assign \new_[496]_  = \new_[53010]_  & \new_[52995]_ ;
  assign \new_[497]_  = \new_[52980]_  & \new_[52965]_ ;
  assign \new_[498]_  = \new_[52950]_  & \new_[52935]_ ;
  assign \new_[499]_  = \new_[52920]_  & \new_[52905]_ ;
  assign \new_[500]_  = \new_[52890]_  & \new_[52875]_ ;
  assign \new_[501]_  = \new_[52860]_  & \new_[52845]_ ;
  assign \new_[502]_  = \new_[52830]_  & \new_[52815]_ ;
  assign \new_[503]_  = \new_[52800]_  & \new_[52785]_ ;
  assign \new_[504]_  = \new_[52770]_  & \new_[52755]_ ;
  assign \new_[505]_  = \new_[52740]_  & \new_[52725]_ ;
  assign \new_[506]_  = \new_[52710]_  & \new_[52695]_ ;
  assign \new_[507]_  = \new_[52680]_  & \new_[52665]_ ;
  assign \new_[508]_  = \new_[52650]_  & \new_[52635]_ ;
  assign \new_[509]_  = \new_[52620]_  & \new_[52605]_ ;
  assign \new_[510]_  = \new_[52590]_  & \new_[52575]_ ;
  assign \new_[511]_  = \new_[52560]_  & \new_[52545]_ ;
  assign \new_[512]_  = \new_[52530]_  & \new_[52515]_ ;
  assign \new_[513]_  = \new_[52500]_  & \new_[52485]_ ;
  assign \new_[514]_  = \new_[52470]_  & \new_[52455]_ ;
  assign \new_[515]_  = \new_[52440]_  & \new_[52425]_ ;
  assign \new_[516]_  = \new_[52410]_  & \new_[52395]_ ;
  assign \new_[517]_  = \new_[52380]_  & \new_[52365]_ ;
  assign \new_[518]_  = \new_[52350]_  & \new_[52335]_ ;
  assign \new_[519]_  = \new_[52320]_  & \new_[52305]_ ;
  assign \new_[520]_  = \new_[52290]_  & \new_[52275]_ ;
  assign \new_[521]_  = \new_[52260]_  & \new_[52245]_ ;
  assign \new_[522]_  = \new_[52230]_  & \new_[52215]_ ;
  assign \new_[523]_  = \new_[52200]_  & \new_[52185]_ ;
  assign \new_[524]_  = \new_[52170]_  & \new_[52155]_ ;
  assign \new_[525]_  = \new_[52140]_  & \new_[52125]_ ;
  assign \new_[526]_  = \new_[52110]_  & \new_[52095]_ ;
  assign \new_[527]_  = \new_[52080]_  & \new_[52065]_ ;
  assign \new_[528]_  = \new_[52050]_  & \new_[52035]_ ;
  assign \new_[529]_  = \new_[52020]_  & \new_[52005]_ ;
  assign \new_[530]_  = \new_[51990]_  & \new_[51975]_ ;
  assign \new_[531]_  = \new_[51960]_  & \new_[51945]_ ;
  assign \new_[532]_  = \new_[51930]_  & \new_[51915]_ ;
  assign \new_[533]_  = \new_[51900]_  & \new_[51885]_ ;
  assign \new_[534]_  = \new_[51870]_  & \new_[51855]_ ;
  assign \new_[535]_  = \new_[51840]_  & \new_[51825]_ ;
  assign \new_[536]_  = \new_[51810]_  & \new_[51795]_ ;
  assign \new_[537]_  = \new_[51780]_  & \new_[51765]_ ;
  assign \new_[538]_  = \new_[51750]_  & \new_[51735]_ ;
  assign \new_[539]_  = \new_[51720]_  & \new_[51705]_ ;
  assign \new_[540]_  = \new_[51690]_  & \new_[51675]_ ;
  assign \new_[541]_  = \new_[51660]_  & \new_[51645]_ ;
  assign \new_[542]_  = \new_[51630]_  & \new_[51615]_ ;
  assign \new_[543]_  = \new_[51600]_  & \new_[51585]_ ;
  assign \new_[544]_  = \new_[51570]_  & \new_[51555]_ ;
  assign \new_[545]_  = \new_[51540]_  & \new_[51525]_ ;
  assign \new_[546]_  = \new_[51510]_  & \new_[51495]_ ;
  assign \new_[547]_  = \new_[51480]_  & \new_[51465]_ ;
  assign \new_[548]_  = \new_[51450]_  & \new_[51435]_ ;
  assign \new_[549]_  = \new_[51420]_  & \new_[51405]_ ;
  assign \new_[550]_  = \new_[51390]_  & \new_[51375]_ ;
  assign \new_[551]_  = \new_[51360]_  & \new_[51345]_ ;
  assign \new_[552]_  = \new_[51330]_  & \new_[51315]_ ;
  assign \new_[553]_  = \new_[51300]_  & \new_[51285]_ ;
  assign \new_[554]_  = \new_[51270]_  & \new_[51255]_ ;
  assign \new_[555]_  = \new_[51240]_  & \new_[51225]_ ;
  assign \new_[556]_  = \new_[51210]_  & \new_[51195]_ ;
  assign \new_[557]_  = \new_[51180]_  & \new_[51165]_ ;
  assign \new_[558]_  = \new_[51150]_  & \new_[51135]_ ;
  assign \new_[559]_  = \new_[51120]_  & \new_[51105]_ ;
  assign \new_[560]_  = \new_[51090]_  & \new_[51075]_ ;
  assign \new_[561]_  = \new_[51060]_  & \new_[51045]_ ;
  assign \new_[562]_  = \new_[51030]_  & \new_[51015]_ ;
  assign \new_[563]_  = \new_[51000]_  & \new_[50985]_ ;
  assign \new_[564]_  = \new_[50970]_  & \new_[50955]_ ;
  assign \new_[565]_  = \new_[50940]_  & \new_[50925]_ ;
  assign \new_[566]_  = \new_[50910]_  & \new_[50895]_ ;
  assign \new_[567]_  = \new_[50880]_  & \new_[50865]_ ;
  assign \new_[568]_  = \new_[50850]_  & \new_[50835]_ ;
  assign \new_[569]_  = \new_[50820]_  & \new_[50805]_ ;
  assign \new_[570]_  = \new_[50790]_  & \new_[50775]_ ;
  assign \new_[571]_  = \new_[50760]_  & \new_[50745]_ ;
  assign \new_[572]_  = \new_[50730]_  & \new_[50715]_ ;
  assign \new_[573]_  = \new_[50700]_  & \new_[50685]_ ;
  assign \new_[574]_  = \new_[50670]_  & \new_[50655]_ ;
  assign \new_[575]_  = \new_[50640]_  & \new_[50625]_ ;
  assign \new_[576]_  = \new_[50610]_  & \new_[50595]_ ;
  assign \new_[577]_  = \new_[50580]_  & \new_[50565]_ ;
  assign \new_[578]_  = \new_[50550]_  & \new_[50535]_ ;
  assign \new_[579]_  = \new_[50520]_  & \new_[50505]_ ;
  assign \new_[580]_  = \new_[50490]_  & \new_[50475]_ ;
  assign \new_[581]_  = \new_[50460]_  & \new_[50445]_ ;
  assign \new_[582]_  = \new_[50430]_  & \new_[50415]_ ;
  assign \new_[583]_  = \new_[50400]_  & \new_[50385]_ ;
  assign \new_[584]_  = \new_[50370]_  & \new_[50355]_ ;
  assign \new_[585]_  = \new_[50340]_  & \new_[50325]_ ;
  assign \new_[586]_  = \new_[50310]_  & \new_[50295]_ ;
  assign \new_[587]_  = \new_[50280]_  & \new_[50265]_ ;
  assign \new_[588]_  = \new_[50250]_  & \new_[50235]_ ;
  assign \new_[589]_  = \new_[50220]_  & \new_[50205]_ ;
  assign \new_[590]_  = \new_[50190]_  & \new_[50175]_ ;
  assign \new_[591]_  = \new_[50160]_  & \new_[50145]_ ;
  assign \new_[592]_  = \new_[50130]_  & \new_[50115]_ ;
  assign \new_[593]_  = \new_[50100]_  & \new_[50085]_ ;
  assign \new_[594]_  = \new_[50070]_  & \new_[50055]_ ;
  assign \new_[595]_  = \new_[50040]_  & \new_[50025]_ ;
  assign \new_[596]_  = \new_[50010]_  & \new_[49995]_ ;
  assign \new_[597]_  = \new_[49980]_  & \new_[49965]_ ;
  assign \new_[598]_  = \new_[49950]_  & \new_[49935]_ ;
  assign \new_[599]_  = \new_[49920]_  & \new_[49905]_ ;
  assign \new_[600]_  = \new_[49890]_  & \new_[49875]_ ;
  assign \new_[601]_  = \new_[49860]_  & \new_[49845]_ ;
  assign \new_[602]_  = \new_[49830]_  & \new_[49815]_ ;
  assign \new_[603]_  = \new_[49800]_  & \new_[49785]_ ;
  assign \new_[604]_  = \new_[49770]_  & \new_[49755]_ ;
  assign \new_[605]_  = \new_[49740]_  & \new_[49725]_ ;
  assign \new_[606]_  = \new_[49710]_  & \new_[49695]_ ;
  assign \new_[607]_  = \new_[49680]_  & \new_[49665]_ ;
  assign \new_[608]_  = \new_[49650]_  & \new_[49635]_ ;
  assign \new_[609]_  = \new_[49620]_  & \new_[49605]_ ;
  assign \new_[610]_  = \new_[49590]_  & \new_[49575]_ ;
  assign \new_[611]_  = \new_[49560]_  & \new_[49545]_ ;
  assign \new_[612]_  = \new_[49530]_  & \new_[49515]_ ;
  assign \new_[613]_  = \new_[49500]_  & \new_[49485]_ ;
  assign \new_[614]_  = \new_[49470]_  & \new_[49455]_ ;
  assign \new_[615]_  = \new_[49440]_  & \new_[49425]_ ;
  assign \new_[616]_  = \new_[49410]_  & \new_[49395]_ ;
  assign \new_[617]_  = \new_[49380]_  & \new_[49365]_ ;
  assign \new_[618]_  = \new_[49350]_  & \new_[49335]_ ;
  assign \new_[619]_  = \new_[49320]_  & \new_[49305]_ ;
  assign \new_[620]_  = \new_[49290]_  & \new_[49275]_ ;
  assign \new_[621]_  = \new_[49260]_  & \new_[49245]_ ;
  assign \new_[622]_  = \new_[49230]_  & \new_[49215]_ ;
  assign \new_[623]_  = \new_[49200]_  & \new_[49185]_ ;
  assign \new_[624]_  = \new_[49170]_  & \new_[49155]_ ;
  assign \new_[625]_  = \new_[49140]_  & \new_[49125]_ ;
  assign \new_[626]_  = \new_[49110]_  & \new_[49095]_ ;
  assign \new_[627]_  = \new_[49080]_  & \new_[49065]_ ;
  assign \new_[628]_  = \new_[49050]_  & \new_[49035]_ ;
  assign \new_[629]_  = \new_[49020]_  & \new_[49005]_ ;
  assign \new_[630]_  = \new_[48990]_  & \new_[48975]_ ;
  assign \new_[631]_  = \new_[48960]_  & \new_[48945]_ ;
  assign \new_[632]_  = \new_[48930]_  & \new_[48915]_ ;
  assign \new_[633]_  = \new_[48900]_  & \new_[48885]_ ;
  assign \new_[634]_  = \new_[48870]_  & \new_[48855]_ ;
  assign \new_[635]_  = \new_[48840]_  & \new_[48825]_ ;
  assign \new_[636]_  = \new_[48810]_  & \new_[48795]_ ;
  assign \new_[637]_  = \new_[48780]_  & \new_[48765]_ ;
  assign \new_[638]_  = \new_[48750]_  & \new_[48735]_ ;
  assign \new_[639]_  = \new_[48720]_  & \new_[48705]_ ;
  assign \new_[640]_  = \new_[48690]_  & \new_[48675]_ ;
  assign \new_[641]_  = \new_[48660]_  & \new_[48645]_ ;
  assign \new_[642]_  = \new_[48630]_  & \new_[48615]_ ;
  assign \new_[643]_  = \new_[48600]_  & \new_[48585]_ ;
  assign \new_[644]_  = \new_[48570]_  & \new_[48555]_ ;
  assign \new_[645]_  = \new_[48540]_  & \new_[48525]_ ;
  assign \new_[646]_  = \new_[48510]_  & \new_[48495]_ ;
  assign \new_[647]_  = \new_[48480]_  & \new_[48465]_ ;
  assign \new_[648]_  = \new_[48450]_  & \new_[48435]_ ;
  assign \new_[649]_  = \new_[48420]_  & \new_[48405]_ ;
  assign \new_[650]_  = \new_[48390]_  & \new_[48375]_ ;
  assign \new_[651]_  = \new_[48360]_  & \new_[48345]_ ;
  assign \new_[652]_  = \new_[48330]_  & \new_[48315]_ ;
  assign \new_[653]_  = \new_[48300]_  & \new_[48285]_ ;
  assign \new_[654]_  = \new_[48270]_  & \new_[48255]_ ;
  assign \new_[655]_  = \new_[48240]_  & \new_[48225]_ ;
  assign \new_[656]_  = \new_[48210]_  & \new_[48195]_ ;
  assign \new_[657]_  = \new_[48180]_  & \new_[48165]_ ;
  assign \new_[658]_  = \new_[48150]_  & \new_[48135]_ ;
  assign \new_[659]_  = \new_[48120]_  & \new_[48105]_ ;
  assign \new_[660]_  = \new_[48090]_  & \new_[48075]_ ;
  assign \new_[661]_  = \new_[48060]_  & \new_[48045]_ ;
  assign \new_[662]_  = \new_[48030]_  & \new_[48015]_ ;
  assign \new_[663]_  = \new_[48000]_  & \new_[47985]_ ;
  assign \new_[664]_  = \new_[47970]_  & \new_[47955]_ ;
  assign \new_[665]_  = \new_[47940]_  & \new_[47925]_ ;
  assign \new_[666]_  = \new_[47910]_  & \new_[47895]_ ;
  assign \new_[667]_  = \new_[47880]_  & \new_[47865]_ ;
  assign \new_[668]_  = \new_[47850]_  & \new_[47835]_ ;
  assign \new_[669]_  = \new_[47820]_  & \new_[47805]_ ;
  assign \new_[670]_  = \new_[47790]_  & \new_[47775]_ ;
  assign \new_[671]_  = \new_[47760]_  & \new_[47745]_ ;
  assign \new_[672]_  = \new_[47730]_  & \new_[47715]_ ;
  assign \new_[673]_  = \new_[47700]_  & \new_[47685]_ ;
  assign \new_[674]_  = \new_[47670]_  & \new_[47655]_ ;
  assign \new_[675]_  = \new_[47640]_  & \new_[47625]_ ;
  assign \new_[676]_  = \new_[47610]_  & \new_[47595]_ ;
  assign \new_[677]_  = \new_[47580]_  & \new_[47565]_ ;
  assign \new_[678]_  = \new_[47550]_  & \new_[47535]_ ;
  assign \new_[679]_  = \new_[47520]_  & \new_[47505]_ ;
  assign \new_[680]_  = \new_[47490]_  & \new_[47475]_ ;
  assign \new_[681]_  = \new_[47460]_  & \new_[47445]_ ;
  assign \new_[682]_  = \new_[47430]_  & \new_[47415]_ ;
  assign \new_[683]_  = \new_[47400]_  & \new_[47385]_ ;
  assign \new_[684]_  = \new_[47370]_  & \new_[47355]_ ;
  assign \new_[685]_  = \new_[47340]_  & \new_[47325]_ ;
  assign \new_[686]_  = \new_[47310]_  & \new_[47295]_ ;
  assign \new_[687]_  = \new_[47280]_  & \new_[47265]_ ;
  assign \new_[688]_  = \new_[47250]_  & \new_[47235]_ ;
  assign \new_[689]_  = \new_[47220]_  & \new_[47205]_ ;
  assign \new_[690]_  = \new_[47190]_  & \new_[47175]_ ;
  assign \new_[691]_  = \new_[47160]_  & \new_[47145]_ ;
  assign \new_[692]_  = \new_[47130]_  & \new_[47115]_ ;
  assign \new_[693]_  = \new_[47100]_  & \new_[47085]_ ;
  assign \new_[694]_  = \new_[47070]_  & \new_[47055]_ ;
  assign \new_[695]_  = \new_[47040]_  & \new_[47025]_ ;
  assign \new_[696]_  = \new_[47010]_  & \new_[46995]_ ;
  assign \new_[697]_  = \new_[46980]_  & \new_[46965]_ ;
  assign \new_[698]_  = \new_[46950]_  & \new_[46935]_ ;
  assign \new_[699]_  = \new_[46920]_  & \new_[46905]_ ;
  assign \new_[700]_  = \new_[46890]_  & \new_[46875]_ ;
  assign \new_[701]_  = \new_[46860]_  & \new_[46845]_ ;
  assign \new_[702]_  = \new_[46830]_  & \new_[46815]_ ;
  assign \new_[703]_  = \new_[46800]_  & \new_[46785]_ ;
  assign \new_[704]_  = \new_[46770]_  & \new_[46755]_ ;
  assign \new_[705]_  = \new_[46740]_  & \new_[46725]_ ;
  assign \new_[706]_  = \new_[46710]_  & \new_[46695]_ ;
  assign \new_[707]_  = \new_[46680]_  & \new_[46665]_ ;
  assign \new_[708]_  = \new_[46650]_  & \new_[46635]_ ;
  assign \new_[709]_  = \new_[46620]_  & \new_[46605]_ ;
  assign \new_[710]_  = \new_[46590]_  & \new_[46575]_ ;
  assign \new_[711]_  = \new_[46560]_  & \new_[46545]_ ;
  assign \new_[712]_  = \new_[46530]_  & \new_[46515]_ ;
  assign \new_[713]_  = \new_[46500]_  & \new_[46485]_ ;
  assign \new_[714]_  = \new_[46470]_  & \new_[46455]_ ;
  assign \new_[715]_  = \new_[46440]_  & \new_[46425]_ ;
  assign \new_[716]_  = \new_[46410]_  & \new_[46395]_ ;
  assign \new_[717]_  = \new_[46380]_  & \new_[46365]_ ;
  assign \new_[718]_  = \new_[46350]_  & \new_[46335]_ ;
  assign \new_[719]_  = \new_[46320]_  & \new_[46305]_ ;
  assign \new_[720]_  = \new_[46290]_  & \new_[46275]_ ;
  assign \new_[721]_  = \new_[46260]_  & \new_[46245]_ ;
  assign \new_[722]_  = \new_[46230]_  & \new_[46215]_ ;
  assign \new_[723]_  = \new_[46200]_  & \new_[46185]_ ;
  assign \new_[724]_  = \new_[46170]_  & \new_[46155]_ ;
  assign \new_[725]_  = \new_[46140]_  & \new_[46125]_ ;
  assign \new_[726]_  = \new_[46110]_  & \new_[46095]_ ;
  assign \new_[727]_  = \new_[46080]_  & \new_[46065]_ ;
  assign \new_[728]_  = \new_[46050]_  & \new_[46035]_ ;
  assign \new_[729]_  = \new_[46020]_  & \new_[46005]_ ;
  assign \new_[730]_  = \new_[45990]_  & \new_[45975]_ ;
  assign \new_[731]_  = \new_[45960]_  & \new_[45945]_ ;
  assign \new_[732]_  = \new_[45930]_  & \new_[45915]_ ;
  assign \new_[733]_  = \new_[45900]_  & \new_[45885]_ ;
  assign \new_[734]_  = \new_[45870]_  & \new_[45855]_ ;
  assign \new_[735]_  = \new_[45840]_  & \new_[45825]_ ;
  assign \new_[736]_  = \new_[45810]_  & \new_[45795]_ ;
  assign \new_[737]_  = \new_[45780]_  & \new_[45765]_ ;
  assign \new_[738]_  = \new_[45750]_  & \new_[45735]_ ;
  assign \new_[739]_  = \new_[45720]_  & \new_[45705]_ ;
  assign \new_[740]_  = \new_[45690]_  & \new_[45675]_ ;
  assign \new_[741]_  = \new_[45660]_  & \new_[45645]_ ;
  assign \new_[742]_  = \new_[45630]_  & \new_[45615]_ ;
  assign \new_[743]_  = \new_[45600]_  & \new_[45585]_ ;
  assign \new_[744]_  = \new_[45570]_  & \new_[45555]_ ;
  assign \new_[745]_  = \new_[45540]_  & \new_[45525]_ ;
  assign \new_[746]_  = \new_[45510]_  & \new_[45495]_ ;
  assign \new_[747]_  = \new_[45480]_  & \new_[45465]_ ;
  assign \new_[748]_  = \new_[45450]_  & \new_[45435]_ ;
  assign \new_[749]_  = \new_[45420]_  & \new_[45405]_ ;
  assign \new_[750]_  = \new_[45390]_  & \new_[45375]_ ;
  assign \new_[751]_  = \new_[45360]_  & \new_[45345]_ ;
  assign \new_[752]_  = \new_[45330]_  & \new_[45315]_ ;
  assign \new_[753]_  = \new_[45300]_  & \new_[45285]_ ;
  assign \new_[754]_  = \new_[45272]_  & \new_[45257]_ ;
  assign \new_[755]_  = \new_[45244]_  & \new_[45229]_ ;
  assign \new_[756]_  = \new_[45216]_  & \new_[45201]_ ;
  assign \new_[757]_  = \new_[45188]_  & \new_[45173]_ ;
  assign \new_[758]_  = \new_[45160]_  & \new_[45145]_ ;
  assign \new_[759]_  = \new_[45132]_  & \new_[45117]_ ;
  assign \new_[760]_  = \new_[45104]_  & \new_[45089]_ ;
  assign \new_[761]_  = \new_[45076]_  & \new_[45061]_ ;
  assign \new_[762]_  = \new_[45048]_  & \new_[45033]_ ;
  assign \new_[763]_  = \new_[45020]_  & \new_[45005]_ ;
  assign \new_[764]_  = \new_[44992]_  & \new_[44977]_ ;
  assign \new_[765]_  = \new_[44964]_  & \new_[44949]_ ;
  assign \new_[766]_  = \new_[44936]_  & \new_[44921]_ ;
  assign \new_[767]_  = \new_[44908]_  & \new_[44893]_ ;
  assign \new_[768]_  = \new_[44880]_  & \new_[44865]_ ;
  assign \new_[769]_  = \new_[44852]_  & \new_[44837]_ ;
  assign \new_[770]_  = \new_[44824]_  & \new_[44809]_ ;
  assign \new_[771]_  = \new_[44796]_  & \new_[44781]_ ;
  assign \new_[772]_  = \new_[44768]_  & \new_[44753]_ ;
  assign \new_[773]_  = \new_[44740]_  & \new_[44725]_ ;
  assign \new_[774]_  = \new_[44712]_  & \new_[44697]_ ;
  assign \new_[775]_  = \new_[44684]_  & \new_[44669]_ ;
  assign \new_[776]_  = \new_[44656]_  & \new_[44641]_ ;
  assign \new_[777]_  = \new_[44628]_  & \new_[44613]_ ;
  assign \new_[778]_  = \new_[44600]_  & \new_[44585]_ ;
  assign \new_[779]_  = \new_[44572]_  & \new_[44557]_ ;
  assign \new_[780]_  = \new_[44544]_  & \new_[44529]_ ;
  assign \new_[781]_  = \new_[44516]_  & \new_[44501]_ ;
  assign \new_[782]_  = \new_[44488]_  & \new_[44473]_ ;
  assign \new_[783]_  = \new_[44460]_  & \new_[44445]_ ;
  assign \new_[784]_  = \new_[44432]_  & \new_[44417]_ ;
  assign \new_[785]_  = \new_[44404]_  & \new_[44389]_ ;
  assign \new_[786]_  = \new_[44376]_  & \new_[44361]_ ;
  assign \new_[787]_  = \new_[44348]_  & \new_[44333]_ ;
  assign \new_[788]_  = \new_[44320]_  & \new_[44305]_ ;
  assign \new_[789]_  = \new_[44292]_  & \new_[44277]_ ;
  assign \new_[790]_  = \new_[44264]_  & \new_[44249]_ ;
  assign \new_[791]_  = \new_[44236]_  & \new_[44221]_ ;
  assign \new_[792]_  = \new_[44208]_  & \new_[44193]_ ;
  assign \new_[793]_  = \new_[44180]_  & \new_[44165]_ ;
  assign \new_[794]_  = \new_[44152]_  & \new_[44137]_ ;
  assign \new_[795]_  = \new_[44124]_  & \new_[44109]_ ;
  assign \new_[796]_  = \new_[44096]_  & \new_[44081]_ ;
  assign \new_[797]_  = \new_[44068]_  & \new_[44053]_ ;
  assign \new_[798]_  = \new_[44040]_  & \new_[44025]_ ;
  assign \new_[799]_  = \new_[44012]_  & \new_[43997]_ ;
  assign \new_[800]_  = \new_[43984]_  & \new_[43969]_ ;
  assign \new_[801]_  = \new_[43956]_  & \new_[43941]_ ;
  assign \new_[802]_  = \new_[43928]_  & \new_[43913]_ ;
  assign \new_[803]_  = \new_[43900]_  & \new_[43885]_ ;
  assign \new_[804]_  = \new_[43872]_  & \new_[43857]_ ;
  assign \new_[805]_  = \new_[43844]_  & \new_[43829]_ ;
  assign \new_[806]_  = \new_[43816]_  & \new_[43801]_ ;
  assign \new_[807]_  = \new_[43788]_  & \new_[43773]_ ;
  assign \new_[808]_  = \new_[43760]_  & \new_[43745]_ ;
  assign \new_[809]_  = \new_[43732]_  & \new_[43717]_ ;
  assign \new_[810]_  = \new_[43704]_  & \new_[43689]_ ;
  assign \new_[811]_  = \new_[43676]_  & \new_[43661]_ ;
  assign \new_[812]_  = \new_[43648]_  & \new_[43633]_ ;
  assign \new_[813]_  = \new_[43620]_  & \new_[43605]_ ;
  assign \new_[814]_  = \new_[43592]_  & \new_[43577]_ ;
  assign \new_[815]_  = \new_[43564]_  & \new_[43549]_ ;
  assign \new_[816]_  = \new_[43536]_  & \new_[43521]_ ;
  assign \new_[817]_  = \new_[43508]_  & \new_[43493]_ ;
  assign \new_[818]_  = \new_[43480]_  & \new_[43465]_ ;
  assign \new_[819]_  = \new_[43452]_  & \new_[43437]_ ;
  assign \new_[820]_  = \new_[43424]_  & \new_[43409]_ ;
  assign \new_[821]_  = \new_[43396]_  & \new_[43381]_ ;
  assign \new_[822]_  = \new_[43368]_  & \new_[43353]_ ;
  assign \new_[823]_  = \new_[43340]_  & \new_[43325]_ ;
  assign \new_[824]_  = \new_[43312]_  & \new_[43297]_ ;
  assign \new_[825]_  = \new_[43284]_  & \new_[43269]_ ;
  assign \new_[826]_  = \new_[43256]_  & \new_[43241]_ ;
  assign \new_[827]_  = \new_[43228]_  & \new_[43213]_ ;
  assign \new_[828]_  = \new_[43200]_  & \new_[43185]_ ;
  assign \new_[829]_  = \new_[43172]_  & \new_[43157]_ ;
  assign \new_[830]_  = \new_[43144]_  & \new_[43129]_ ;
  assign \new_[831]_  = \new_[43116]_  & \new_[43101]_ ;
  assign \new_[832]_  = \new_[43088]_  & \new_[43073]_ ;
  assign \new_[833]_  = \new_[43060]_  & \new_[43045]_ ;
  assign \new_[834]_  = \new_[43032]_  & \new_[43017]_ ;
  assign \new_[835]_  = \new_[43004]_  & \new_[42989]_ ;
  assign \new_[836]_  = \new_[42976]_  & \new_[42961]_ ;
  assign \new_[837]_  = \new_[42948]_  & \new_[42933]_ ;
  assign \new_[838]_  = \new_[42920]_  & \new_[42905]_ ;
  assign \new_[839]_  = \new_[42892]_  & \new_[42877]_ ;
  assign \new_[840]_  = \new_[42864]_  & \new_[42849]_ ;
  assign \new_[841]_  = \new_[42836]_  & \new_[42821]_ ;
  assign \new_[842]_  = \new_[42808]_  & \new_[42793]_ ;
  assign \new_[843]_  = \new_[42780]_  & \new_[42765]_ ;
  assign \new_[844]_  = \new_[42752]_  & \new_[42737]_ ;
  assign \new_[845]_  = \new_[42724]_  & \new_[42709]_ ;
  assign \new_[846]_  = \new_[42696]_  & \new_[42681]_ ;
  assign \new_[847]_  = \new_[42668]_  & \new_[42653]_ ;
  assign \new_[848]_  = \new_[42640]_  & \new_[42625]_ ;
  assign \new_[849]_  = \new_[42612]_  & \new_[42597]_ ;
  assign \new_[850]_  = \new_[42584]_  & \new_[42569]_ ;
  assign \new_[851]_  = \new_[42556]_  & \new_[42541]_ ;
  assign \new_[852]_  = \new_[42528]_  & \new_[42513]_ ;
  assign \new_[853]_  = \new_[42500]_  & \new_[42485]_ ;
  assign \new_[854]_  = \new_[42472]_  & \new_[42457]_ ;
  assign \new_[855]_  = \new_[42444]_  & \new_[42429]_ ;
  assign \new_[856]_  = \new_[42416]_  & \new_[42401]_ ;
  assign \new_[857]_  = \new_[42388]_  & \new_[42373]_ ;
  assign \new_[858]_  = \new_[42360]_  & \new_[42345]_ ;
  assign \new_[859]_  = \new_[42332]_  & \new_[42317]_ ;
  assign \new_[860]_  = \new_[42304]_  & \new_[42289]_ ;
  assign \new_[861]_  = \new_[42276]_  & \new_[42261]_ ;
  assign \new_[862]_  = \new_[42248]_  & \new_[42233]_ ;
  assign \new_[863]_  = \new_[42220]_  & \new_[42205]_ ;
  assign \new_[864]_  = \new_[42192]_  & \new_[42177]_ ;
  assign \new_[865]_  = \new_[42164]_  & \new_[42149]_ ;
  assign \new_[866]_  = \new_[42136]_  & \new_[42121]_ ;
  assign \new_[867]_  = \new_[42108]_  & \new_[42093]_ ;
  assign \new_[868]_  = \new_[42080]_  & \new_[42065]_ ;
  assign \new_[869]_  = \new_[42052]_  & \new_[42037]_ ;
  assign \new_[870]_  = \new_[42024]_  & \new_[42009]_ ;
  assign \new_[871]_  = \new_[41996]_  & \new_[41981]_ ;
  assign \new_[872]_  = \new_[41968]_  & \new_[41953]_ ;
  assign \new_[873]_  = \new_[41940]_  & \new_[41925]_ ;
  assign \new_[874]_  = \new_[41912]_  & \new_[41897]_ ;
  assign \new_[875]_  = \new_[41884]_  & \new_[41869]_ ;
  assign \new_[876]_  = \new_[41856]_  & \new_[41841]_ ;
  assign \new_[877]_  = \new_[41828]_  & \new_[41813]_ ;
  assign \new_[878]_  = \new_[41800]_  & \new_[41785]_ ;
  assign \new_[879]_  = \new_[41772]_  & \new_[41757]_ ;
  assign \new_[880]_  = \new_[41744]_  & \new_[41729]_ ;
  assign \new_[881]_  = \new_[41716]_  & \new_[41701]_ ;
  assign \new_[882]_  = \new_[41688]_  & \new_[41673]_ ;
  assign \new_[883]_  = \new_[41660]_  & \new_[41645]_ ;
  assign \new_[884]_  = \new_[41632]_  & \new_[41617]_ ;
  assign \new_[885]_  = \new_[41604]_  & \new_[41589]_ ;
  assign \new_[886]_  = \new_[41576]_  & \new_[41561]_ ;
  assign \new_[887]_  = \new_[41548]_  & \new_[41533]_ ;
  assign \new_[888]_  = \new_[41520]_  & \new_[41505]_ ;
  assign \new_[889]_  = \new_[41492]_  & \new_[41477]_ ;
  assign \new_[890]_  = \new_[41464]_  & \new_[41449]_ ;
  assign \new_[891]_  = \new_[41436]_  & \new_[41421]_ ;
  assign \new_[892]_  = \new_[41408]_  & \new_[41393]_ ;
  assign \new_[893]_  = \new_[41380]_  & \new_[41365]_ ;
  assign \new_[894]_  = \new_[41352]_  & \new_[41337]_ ;
  assign \new_[895]_  = \new_[41324]_  & \new_[41309]_ ;
  assign \new_[896]_  = \new_[41296]_  & \new_[41281]_ ;
  assign \new_[897]_  = \new_[41268]_  & \new_[41253]_ ;
  assign \new_[898]_  = \new_[41240]_  & \new_[41225]_ ;
  assign \new_[899]_  = \new_[41212]_  & \new_[41197]_ ;
  assign \new_[900]_  = \new_[41184]_  & \new_[41169]_ ;
  assign \new_[901]_  = \new_[41156]_  & \new_[41141]_ ;
  assign \new_[902]_  = \new_[41128]_  & \new_[41113]_ ;
  assign \new_[903]_  = \new_[41100]_  & \new_[41085]_ ;
  assign \new_[904]_  = \new_[41072]_  & \new_[41057]_ ;
  assign \new_[905]_  = \new_[41044]_  & \new_[41029]_ ;
  assign \new_[906]_  = \new_[41016]_  & \new_[41001]_ ;
  assign \new_[907]_  = \new_[40988]_  & \new_[40973]_ ;
  assign \new_[908]_  = \new_[40960]_  & \new_[40945]_ ;
  assign \new_[909]_  = \new_[40932]_  & \new_[40917]_ ;
  assign \new_[910]_  = \new_[40904]_  & \new_[40889]_ ;
  assign \new_[911]_  = \new_[40876]_  & \new_[40861]_ ;
  assign \new_[912]_  = \new_[40848]_  & \new_[40833]_ ;
  assign \new_[913]_  = \new_[40820]_  & \new_[40805]_ ;
  assign \new_[914]_  = \new_[40792]_  & \new_[40777]_ ;
  assign \new_[915]_  = \new_[40764]_  & \new_[40749]_ ;
  assign \new_[916]_  = \new_[40736]_  & \new_[40721]_ ;
  assign \new_[917]_  = \new_[40708]_  & \new_[40693]_ ;
  assign \new_[918]_  = \new_[40680]_  & \new_[40665]_ ;
  assign \new_[919]_  = \new_[40652]_  & \new_[40637]_ ;
  assign \new_[920]_  = \new_[40624]_  & \new_[40609]_ ;
  assign \new_[921]_  = \new_[40596]_  & \new_[40581]_ ;
  assign \new_[922]_  = \new_[40568]_  & \new_[40553]_ ;
  assign \new_[923]_  = \new_[40540]_  & \new_[40525]_ ;
  assign \new_[924]_  = \new_[40512]_  & \new_[40497]_ ;
  assign \new_[925]_  = \new_[40484]_  & \new_[40469]_ ;
  assign \new_[926]_  = \new_[40456]_  & \new_[40441]_ ;
  assign \new_[927]_  = \new_[40428]_  & \new_[40413]_ ;
  assign \new_[928]_  = \new_[40400]_  & \new_[40385]_ ;
  assign \new_[929]_  = \new_[40372]_  & \new_[40357]_ ;
  assign \new_[930]_  = \new_[40344]_  & \new_[40329]_ ;
  assign \new_[931]_  = \new_[40316]_  & \new_[40301]_ ;
  assign \new_[932]_  = \new_[40288]_  & \new_[40273]_ ;
  assign \new_[933]_  = \new_[40260]_  & \new_[40245]_ ;
  assign \new_[934]_  = \new_[40232]_  & \new_[40217]_ ;
  assign \new_[935]_  = \new_[40204]_  & \new_[40189]_ ;
  assign \new_[936]_  = \new_[40176]_  & \new_[40161]_ ;
  assign \new_[937]_  = \new_[40148]_  & \new_[40133]_ ;
  assign \new_[938]_  = \new_[40120]_  & \new_[40105]_ ;
  assign \new_[939]_  = \new_[40092]_  & \new_[40077]_ ;
  assign \new_[940]_  = \new_[40064]_  & \new_[40049]_ ;
  assign \new_[941]_  = \new_[40036]_  & \new_[40021]_ ;
  assign \new_[942]_  = \new_[40008]_  & \new_[39993]_ ;
  assign \new_[943]_  = \new_[39980]_  & \new_[39965]_ ;
  assign \new_[944]_  = \new_[39952]_  & \new_[39937]_ ;
  assign \new_[945]_  = \new_[39924]_  & \new_[39909]_ ;
  assign \new_[946]_  = \new_[39896]_  & \new_[39881]_ ;
  assign \new_[947]_  = \new_[39868]_  & \new_[39853]_ ;
  assign \new_[948]_  = \new_[39840]_  & \new_[39825]_ ;
  assign \new_[949]_  = \new_[39812]_  & \new_[39797]_ ;
  assign \new_[950]_  = \new_[39784]_  & \new_[39769]_ ;
  assign \new_[951]_  = \new_[39756]_  & \new_[39741]_ ;
  assign \new_[952]_  = \new_[39728]_  & \new_[39713]_ ;
  assign \new_[953]_  = \new_[39700]_  & \new_[39685]_ ;
  assign \new_[954]_  = \new_[39672]_  & \new_[39657]_ ;
  assign \new_[955]_  = \new_[39644]_  & \new_[39629]_ ;
  assign \new_[956]_  = \new_[39616]_  & \new_[39601]_ ;
  assign \new_[957]_  = \new_[39588]_  & \new_[39573]_ ;
  assign \new_[958]_  = \new_[39560]_  & \new_[39545]_ ;
  assign \new_[959]_  = \new_[39532]_  & \new_[39517]_ ;
  assign \new_[960]_  = \new_[39504]_  & \new_[39489]_ ;
  assign \new_[961]_  = \new_[39476]_  & \new_[39461]_ ;
  assign \new_[962]_  = \new_[39448]_  & \new_[39433]_ ;
  assign \new_[963]_  = \new_[39420]_  & \new_[39405]_ ;
  assign \new_[964]_  = \new_[39392]_  & \new_[39377]_ ;
  assign \new_[965]_  = \new_[39364]_  & \new_[39349]_ ;
  assign \new_[966]_  = \new_[39336]_  & \new_[39321]_ ;
  assign \new_[967]_  = \new_[39308]_  & \new_[39293]_ ;
  assign \new_[968]_  = \new_[39280]_  & \new_[39265]_ ;
  assign \new_[969]_  = \new_[39252]_  & \new_[39237]_ ;
  assign \new_[970]_  = \new_[39224]_  & \new_[39209]_ ;
  assign \new_[971]_  = \new_[39196]_  & \new_[39181]_ ;
  assign \new_[972]_  = \new_[39168]_  & \new_[39153]_ ;
  assign \new_[973]_  = \new_[39140]_  & \new_[39125]_ ;
  assign \new_[974]_  = \new_[39112]_  & \new_[39097]_ ;
  assign \new_[975]_  = \new_[39084]_  & \new_[39069]_ ;
  assign \new_[976]_  = \new_[39056]_  & \new_[39041]_ ;
  assign \new_[977]_  = \new_[39028]_  & \new_[39013]_ ;
  assign \new_[978]_  = \new_[39000]_  & \new_[38985]_ ;
  assign \new_[979]_  = \new_[38972]_  & \new_[38957]_ ;
  assign \new_[980]_  = \new_[38944]_  & \new_[38929]_ ;
  assign \new_[981]_  = \new_[38916]_  & \new_[38901]_ ;
  assign \new_[982]_  = \new_[38888]_  & \new_[38873]_ ;
  assign \new_[983]_  = \new_[38860]_  & \new_[38845]_ ;
  assign \new_[984]_  = \new_[38832]_  & \new_[38817]_ ;
  assign \new_[985]_  = \new_[38804]_  & \new_[38789]_ ;
  assign \new_[986]_  = \new_[38776]_  & \new_[38761]_ ;
  assign \new_[987]_  = \new_[38748]_  & \new_[38733]_ ;
  assign \new_[988]_  = \new_[38720]_  & \new_[38705]_ ;
  assign \new_[989]_  = \new_[38692]_  & \new_[38677]_ ;
  assign \new_[990]_  = \new_[38664]_  & \new_[38649]_ ;
  assign \new_[991]_  = \new_[38636]_  & \new_[38621]_ ;
  assign \new_[992]_  = \new_[38608]_  & \new_[38593]_ ;
  assign \new_[993]_  = \new_[38580]_  & \new_[38565]_ ;
  assign \new_[994]_  = \new_[38552]_  & \new_[38537]_ ;
  assign \new_[995]_  = \new_[38524]_  & \new_[38509]_ ;
  assign \new_[996]_  = \new_[38496]_  & \new_[38481]_ ;
  assign \new_[997]_  = \new_[38468]_  & \new_[38453]_ ;
  assign \new_[998]_  = \new_[38440]_  & \new_[38425]_ ;
  assign \new_[999]_  = \new_[38412]_  & \new_[38397]_ ;
  assign \new_[1000]_  = \new_[38384]_  & \new_[38369]_ ;
  assign \new_[1001]_  = \new_[38356]_  & \new_[38341]_ ;
  assign \new_[1002]_  = \new_[38328]_  & \new_[38313]_ ;
  assign \new_[1003]_  = \new_[38300]_  & \new_[38285]_ ;
  assign \new_[1004]_  = \new_[38272]_  & \new_[38257]_ ;
  assign \new_[1005]_  = \new_[38244]_  & \new_[38229]_ ;
  assign \new_[1006]_  = \new_[38216]_  & \new_[38201]_ ;
  assign \new_[1007]_  = \new_[38188]_  & \new_[38173]_ ;
  assign \new_[1008]_  = \new_[38160]_  & \new_[38145]_ ;
  assign \new_[1009]_  = \new_[38132]_  & \new_[38117]_ ;
  assign \new_[1010]_  = \new_[38104]_  & \new_[38089]_ ;
  assign \new_[1011]_  = \new_[38076]_  & \new_[38061]_ ;
  assign \new_[1012]_  = \new_[38048]_  & \new_[38033]_ ;
  assign \new_[1013]_  = \new_[38020]_  & \new_[38005]_ ;
  assign \new_[1014]_  = \new_[37992]_  & \new_[37977]_ ;
  assign \new_[1015]_  = \new_[37964]_  & \new_[37949]_ ;
  assign \new_[1016]_  = \new_[37936]_  & \new_[37921]_ ;
  assign \new_[1017]_  = \new_[37908]_  & \new_[37893]_ ;
  assign \new_[1018]_  = \new_[37880]_  & \new_[37865]_ ;
  assign \new_[1019]_  = \new_[37852]_  & \new_[37837]_ ;
  assign \new_[1020]_  = \new_[37824]_  & \new_[37809]_ ;
  assign \new_[1021]_  = \new_[37796]_  & \new_[37781]_ ;
  assign \new_[1022]_  = \new_[37768]_  & \new_[37753]_ ;
  assign \new_[1023]_  = \new_[37740]_  & \new_[37725]_ ;
  assign \new_[1024]_  = \new_[37712]_  & \new_[37697]_ ;
  assign \new_[1025]_  = \new_[37684]_  & \new_[37669]_ ;
  assign \new_[1026]_  = \new_[37656]_  & \new_[37641]_ ;
  assign \new_[1027]_  = \new_[37628]_  & \new_[37613]_ ;
  assign \new_[1028]_  = \new_[37600]_  & \new_[37585]_ ;
  assign \new_[1029]_  = \new_[37572]_  & \new_[37557]_ ;
  assign \new_[1030]_  = \new_[37544]_  & \new_[37529]_ ;
  assign \new_[1031]_  = \new_[37516]_  & \new_[37501]_ ;
  assign \new_[1032]_  = \new_[37488]_  & \new_[37473]_ ;
  assign \new_[1033]_  = \new_[37460]_  & \new_[37445]_ ;
  assign \new_[1034]_  = \new_[37432]_  & \new_[37417]_ ;
  assign \new_[1035]_  = \new_[37404]_  & \new_[37389]_ ;
  assign \new_[1036]_  = \new_[37376]_  & \new_[37361]_ ;
  assign \new_[1037]_  = \new_[37348]_  & \new_[37333]_ ;
  assign \new_[1038]_  = \new_[37320]_  & \new_[37305]_ ;
  assign \new_[1039]_  = \new_[37292]_  & \new_[37277]_ ;
  assign \new_[1040]_  = \new_[37264]_  & \new_[37249]_ ;
  assign \new_[1041]_  = \new_[37236]_  & \new_[37221]_ ;
  assign \new_[1042]_  = \new_[37208]_  & \new_[37193]_ ;
  assign \new_[1043]_  = \new_[37180]_  & \new_[37165]_ ;
  assign \new_[1044]_  = \new_[37152]_  & \new_[37137]_ ;
  assign \new_[1045]_  = \new_[37124]_  & \new_[37109]_ ;
  assign \new_[1046]_  = \new_[37096]_  & \new_[37081]_ ;
  assign \new_[1047]_  = \new_[37068]_  & \new_[37053]_ ;
  assign \new_[1048]_  = \new_[37040]_  & \new_[37025]_ ;
  assign \new_[1049]_  = \new_[37012]_  & \new_[36997]_ ;
  assign \new_[1050]_  = \new_[36984]_  & \new_[36969]_ ;
  assign \new_[1051]_  = \new_[36956]_  & \new_[36941]_ ;
  assign \new_[1052]_  = \new_[36928]_  & \new_[36913]_ ;
  assign \new_[1053]_  = \new_[36900]_  & \new_[36885]_ ;
  assign \new_[1054]_  = \new_[36872]_  & \new_[36857]_ ;
  assign \new_[1055]_  = \new_[36844]_  & \new_[36829]_ ;
  assign \new_[1056]_  = \new_[36816]_  & \new_[36801]_ ;
  assign \new_[1057]_  = \new_[36788]_  & \new_[36773]_ ;
  assign \new_[1058]_  = \new_[36760]_  & \new_[36745]_ ;
  assign \new_[1059]_  = \new_[36732]_  & \new_[36717]_ ;
  assign \new_[1060]_  = \new_[36704]_  & \new_[36689]_ ;
  assign \new_[1061]_  = \new_[36676]_  & \new_[36661]_ ;
  assign \new_[1062]_  = \new_[36648]_  & \new_[36633]_ ;
  assign \new_[1063]_  = \new_[36620]_  & \new_[36605]_ ;
  assign \new_[1064]_  = \new_[36592]_  & \new_[36577]_ ;
  assign \new_[1065]_  = \new_[36564]_  & \new_[36549]_ ;
  assign \new_[1066]_  = \new_[36536]_  & \new_[36521]_ ;
  assign \new_[1067]_  = \new_[36508]_  & \new_[36493]_ ;
  assign \new_[1068]_  = \new_[36480]_  & \new_[36465]_ ;
  assign \new_[1069]_  = \new_[36452]_  & \new_[36437]_ ;
  assign \new_[1070]_  = \new_[36424]_  & \new_[36409]_ ;
  assign \new_[1071]_  = \new_[36396]_  & \new_[36381]_ ;
  assign \new_[1072]_  = \new_[36368]_  & \new_[36353]_ ;
  assign \new_[1073]_  = \new_[36340]_  & \new_[36325]_ ;
  assign \new_[1074]_  = \new_[36312]_  & \new_[36297]_ ;
  assign \new_[1075]_  = \new_[36284]_  & \new_[36269]_ ;
  assign \new_[1076]_  = \new_[36256]_  & \new_[36241]_ ;
  assign \new_[1077]_  = \new_[36228]_  & \new_[36213]_ ;
  assign \new_[1078]_  = \new_[36200]_  & \new_[36185]_ ;
  assign \new_[1079]_  = \new_[36172]_  & \new_[36157]_ ;
  assign \new_[1080]_  = \new_[36144]_  & \new_[36129]_ ;
  assign \new_[1081]_  = \new_[36116]_  & \new_[36101]_ ;
  assign \new_[1082]_  = \new_[36088]_  & \new_[36073]_ ;
  assign \new_[1083]_  = \new_[36060]_  & \new_[36045]_ ;
  assign \new_[1084]_  = \new_[36032]_  & \new_[36017]_ ;
  assign \new_[1085]_  = \new_[36004]_  & \new_[35989]_ ;
  assign \new_[1086]_  = \new_[35976]_  & \new_[35961]_ ;
  assign \new_[1087]_  = \new_[35948]_  & \new_[35933]_ ;
  assign \new_[1088]_  = \new_[35920]_  & \new_[35905]_ ;
  assign \new_[1089]_  = \new_[35892]_  & \new_[35877]_ ;
  assign \new_[1090]_  = \new_[35864]_  & \new_[35849]_ ;
  assign \new_[1091]_  = \new_[35836]_  & \new_[35821]_ ;
  assign \new_[1092]_  = \new_[35808]_  & \new_[35793]_ ;
  assign \new_[1093]_  = \new_[35780]_  & \new_[35765]_ ;
  assign \new_[1094]_  = \new_[35752]_  & \new_[35737]_ ;
  assign \new_[1095]_  = \new_[35724]_  & \new_[35709]_ ;
  assign \new_[1096]_  = \new_[35696]_  & \new_[35681]_ ;
  assign \new_[1097]_  = \new_[35668]_  & \new_[35653]_ ;
  assign \new_[1098]_  = \new_[35640]_  & \new_[35625]_ ;
  assign \new_[1099]_  = \new_[35612]_  & \new_[35597]_ ;
  assign \new_[1100]_  = \new_[35584]_  & \new_[35569]_ ;
  assign \new_[1101]_  = \new_[35556]_  & \new_[35541]_ ;
  assign \new_[1102]_  = \new_[35528]_  & \new_[35513]_ ;
  assign \new_[1103]_  = \new_[35500]_  & \new_[35485]_ ;
  assign \new_[1104]_  = \new_[35472]_  & \new_[35457]_ ;
  assign \new_[1105]_  = \new_[35444]_  & \new_[35429]_ ;
  assign \new_[1106]_  = \new_[35416]_  & \new_[35401]_ ;
  assign \new_[1107]_  = \new_[35388]_  & \new_[35373]_ ;
  assign \new_[1108]_  = \new_[35360]_  & \new_[35345]_ ;
  assign \new_[1109]_  = \new_[35332]_  & \new_[35317]_ ;
  assign \new_[1110]_  = \new_[35304]_  & \new_[35289]_ ;
  assign \new_[1111]_  = \new_[35276]_  & \new_[35261]_ ;
  assign \new_[1112]_  = \new_[35248]_  & \new_[35233]_ ;
  assign \new_[1113]_  = \new_[35220]_  & \new_[35205]_ ;
  assign \new_[1114]_  = \new_[35192]_  & \new_[35177]_ ;
  assign \new_[1115]_  = \new_[35164]_  & \new_[35149]_ ;
  assign \new_[1116]_  = \new_[35136]_  & \new_[35121]_ ;
  assign \new_[1117]_  = \new_[35108]_  & \new_[35093]_ ;
  assign \new_[1118]_  = \new_[35080]_  & \new_[35065]_ ;
  assign \new_[1119]_  = \new_[35052]_  & \new_[35037]_ ;
  assign \new_[1120]_  = \new_[35024]_  & \new_[35009]_ ;
  assign \new_[1121]_  = \new_[34996]_  & \new_[34981]_ ;
  assign \new_[1122]_  = \new_[34968]_  & \new_[34953]_ ;
  assign \new_[1123]_  = \new_[34940]_  & \new_[34925]_ ;
  assign \new_[1124]_  = \new_[34912]_  & \new_[34897]_ ;
  assign \new_[1125]_  = \new_[34884]_  & \new_[34869]_ ;
  assign \new_[1126]_  = \new_[34856]_  & \new_[34841]_ ;
  assign \new_[1127]_  = \new_[34828]_  & \new_[34813]_ ;
  assign \new_[1128]_  = \new_[34800]_  & \new_[34785]_ ;
  assign \new_[1129]_  = \new_[34772]_  & \new_[34757]_ ;
  assign \new_[1130]_  = \new_[34744]_  & \new_[34729]_ ;
  assign \new_[1131]_  = \new_[34716]_  & \new_[34701]_ ;
  assign \new_[1132]_  = \new_[34688]_  & \new_[34673]_ ;
  assign \new_[1133]_  = \new_[34660]_  & \new_[34645]_ ;
  assign \new_[1134]_  = \new_[34632]_  & \new_[34617]_ ;
  assign \new_[1135]_  = \new_[34604]_  & \new_[34589]_ ;
  assign \new_[1136]_  = \new_[34576]_  & \new_[34561]_ ;
  assign \new_[1137]_  = \new_[34548]_  & \new_[34533]_ ;
  assign \new_[1138]_  = \new_[34520]_  & \new_[34505]_ ;
  assign \new_[1139]_  = \new_[34492]_  & \new_[34477]_ ;
  assign \new_[1140]_  = \new_[34464]_  & \new_[34449]_ ;
  assign \new_[1141]_  = \new_[34436]_  & \new_[34421]_ ;
  assign \new_[1142]_  = \new_[34408]_  & \new_[34393]_ ;
  assign \new_[1143]_  = \new_[34380]_  & \new_[34365]_ ;
  assign \new_[1144]_  = \new_[34352]_  & \new_[34337]_ ;
  assign \new_[1145]_  = \new_[34324]_  & \new_[34309]_ ;
  assign \new_[1146]_  = \new_[34296]_  & \new_[34281]_ ;
  assign \new_[1147]_  = \new_[34268]_  & \new_[34253]_ ;
  assign \new_[1148]_  = \new_[34240]_  & \new_[34225]_ ;
  assign \new_[1149]_  = \new_[34212]_  & \new_[34197]_ ;
  assign \new_[1150]_  = \new_[34184]_  & \new_[34169]_ ;
  assign \new_[1151]_  = \new_[34156]_  & \new_[34141]_ ;
  assign \new_[1152]_  = \new_[34128]_  & \new_[34113]_ ;
  assign \new_[1153]_  = \new_[34100]_  & \new_[34085]_ ;
  assign \new_[1154]_  = \new_[34072]_  & \new_[34057]_ ;
  assign \new_[1155]_  = \new_[34044]_  & \new_[34029]_ ;
  assign \new_[1156]_  = \new_[34016]_  & \new_[34001]_ ;
  assign \new_[1157]_  = \new_[33988]_  & \new_[33973]_ ;
  assign \new_[1158]_  = \new_[33960]_  & \new_[33945]_ ;
  assign \new_[1159]_  = \new_[33932]_  & \new_[33917]_ ;
  assign \new_[1160]_  = \new_[33904]_  & \new_[33889]_ ;
  assign \new_[1161]_  = \new_[33876]_  & \new_[33861]_ ;
  assign \new_[1162]_  = \new_[33848]_  & \new_[33833]_ ;
  assign \new_[1163]_  = \new_[33820]_  & \new_[33805]_ ;
  assign \new_[1164]_  = \new_[33792]_  & \new_[33777]_ ;
  assign \new_[1165]_  = \new_[33764]_  & \new_[33749]_ ;
  assign \new_[1166]_  = \new_[33736]_  & \new_[33721]_ ;
  assign \new_[1167]_  = \new_[33708]_  & \new_[33693]_ ;
  assign \new_[1168]_  = \new_[33680]_  & \new_[33665]_ ;
  assign \new_[1169]_  = \new_[33652]_  & \new_[33637]_ ;
  assign \new_[1170]_  = \new_[33624]_  & \new_[33609]_ ;
  assign \new_[1171]_  = \new_[33596]_  & \new_[33581]_ ;
  assign \new_[1172]_  = \new_[33568]_  & \new_[33553]_ ;
  assign \new_[1173]_  = \new_[33540]_  & \new_[33525]_ ;
  assign \new_[1174]_  = \new_[33512]_  & \new_[33497]_ ;
  assign \new_[1175]_  = \new_[33484]_  & \new_[33469]_ ;
  assign \new_[1176]_  = \new_[33456]_  & \new_[33441]_ ;
  assign \new_[1177]_  = \new_[33428]_  & \new_[33413]_ ;
  assign \new_[1178]_  = \new_[33400]_  & \new_[33385]_ ;
  assign \new_[1179]_  = \new_[33372]_  & \new_[33357]_ ;
  assign \new_[1180]_  = \new_[33344]_  & \new_[33329]_ ;
  assign \new_[1181]_  = \new_[33316]_  & \new_[33301]_ ;
  assign \new_[1182]_  = \new_[33288]_  & \new_[33273]_ ;
  assign \new_[1183]_  = \new_[33260]_  & \new_[33245]_ ;
  assign \new_[1184]_  = \new_[33232]_  & \new_[33217]_ ;
  assign \new_[1185]_  = \new_[33204]_  & \new_[33189]_ ;
  assign \new_[1186]_  = \new_[33176]_  & \new_[33161]_ ;
  assign \new_[1187]_  = \new_[33148]_  & \new_[33133]_ ;
  assign \new_[1188]_  = \new_[33120]_  & \new_[33105]_ ;
  assign \new_[1189]_  = \new_[33092]_  & \new_[33077]_ ;
  assign \new_[1190]_  = \new_[33064]_  & \new_[33049]_ ;
  assign \new_[1191]_  = \new_[33036]_  & \new_[33021]_ ;
  assign \new_[1192]_  = \new_[33008]_  & \new_[32993]_ ;
  assign \new_[1193]_  = \new_[32980]_  & \new_[32965]_ ;
  assign \new_[1194]_  = \new_[32952]_  & \new_[32937]_ ;
  assign \new_[1195]_  = \new_[32924]_  & \new_[32909]_ ;
  assign \new_[1196]_  = \new_[32896]_  & \new_[32881]_ ;
  assign \new_[1197]_  = \new_[32868]_  & \new_[32853]_ ;
  assign \new_[1198]_  = \new_[32840]_  & \new_[32825]_ ;
  assign \new_[1199]_  = \new_[32812]_  & \new_[32797]_ ;
  assign \new_[1200]_  = \new_[32784]_  & \new_[32769]_ ;
  assign \new_[1201]_  = \new_[32756]_  & \new_[32741]_ ;
  assign \new_[1202]_  = \new_[32728]_  & \new_[32713]_ ;
  assign \new_[1203]_  = \new_[32700]_  & \new_[32685]_ ;
  assign \new_[1204]_  = \new_[32672]_  & \new_[32657]_ ;
  assign \new_[1205]_  = \new_[32644]_  & \new_[32629]_ ;
  assign \new_[1206]_  = \new_[32616]_  & \new_[32601]_ ;
  assign \new_[1207]_  = \new_[32588]_  & \new_[32573]_ ;
  assign \new_[1208]_  = \new_[32560]_  & \new_[32545]_ ;
  assign \new_[1209]_  = \new_[32532]_  & \new_[32517]_ ;
  assign \new_[1210]_  = \new_[32504]_  & \new_[32489]_ ;
  assign \new_[1211]_  = \new_[32476]_  & \new_[32461]_ ;
  assign \new_[1212]_  = \new_[32448]_  & \new_[32433]_ ;
  assign \new_[1213]_  = \new_[32420]_  & \new_[32405]_ ;
  assign \new_[1214]_  = \new_[32392]_  & \new_[32377]_ ;
  assign \new_[1215]_  = \new_[32364]_  & \new_[32349]_ ;
  assign \new_[1216]_  = \new_[32336]_  & \new_[32321]_ ;
  assign \new_[1217]_  = \new_[32308]_  & \new_[32293]_ ;
  assign \new_[1218]_  = \new_[32280]_  & \new_[32265]_ ;
  assign \new_[1219]_  = \new_[32252]_  & \new_[32237]_ ;
  assign \new_[1220]_  = \new_[32224]_  & \new_[32209]_ ;
  assign \new_[1221]_  = \new_[32196]_  & \new_[32181]_ ;
  assign \new_[1222]_  = \new_[32168]_  & \new_[32153]_ ;
  assign \new_[1223]_  = \new_[32140]_  & \new_[32125]_ ;
  assign \new_[1224]_  = \new_[32112]_  & \new_[32097]_ ;
  assign \new_[1225]_  = \new_[32084]_  & \new_[32069]_ ;
  assign \new_[1226]_  = \new_[32056]_  & \new_[32041]_ ;
  assign \new_[1227]_  = \new_[32028]_  & \new_[32013]_ ;
  assign \new_[1228]_  = \new_[32000]_  & \new_[31985]_ ;
  assign \new_[1229]_  = \new_[31972]_  & \new_[31957]_ ;
  assign \new_[1230]_  = \new_[31944]_  & \new_[31929]_ ;
  assign \new_[1231]_  = \new_[31916]_  & \new_[31901]_ ;
  assign \new_[1232]_  = \new_[31888]_  & \new_[31873]_ ;
  assign \new_[1233]_  = \new_[31860]_  & \new_[31845]_ ;
  assign \new_[1234]_  = \new_[31832]_  & \new_[31817]_ ;
  assign \new_[1235]_  = \new_[31804]_  & \new_[31789]_ ;
  assign \new_[1236]_  = \new_[31776]_  & \new_[31761]_ ;
  assign \new_[1237]_  = \new_[31748]_  & \new_[31733]_ ;
  assign \new_[1238]_  = \new_[31720]_  & \new_[31705]_ ;
  assign \new_[1239]_  = \new_[31692]_  & \new_[31677]_ ;
  assign \new_[1240]_  = \new_[31664]_  & \new_[31649]_ ;
  assign \new_[1241]_  = \new_[31636]_  & \new_[31621]_ ;
  assign \new_[1242]_  = \new_[31608]_  & \new_[31593]_ ;
  assign \new_[1243]_  = \new_[31580]_  & \new_[31565]_ ;
  assign \new_[1244]_  = \new_[31552]_  & \new_[31537]_ ;
  assign \new_[1245]_  = \new_[31524]_  & \new_[31509]_ ;
  assign \new_[1246]_  = \new_[31496]_  & \new_[31481]_ ;
  assign \new_[1247]_  = \new_[31468]_  & \new_[31453]_ ;
  assign \new_[1248]_  = \new_[31440]_  & \new_[31425]_ ;
  assign \new_[1249]_  = \new_[31412]_  & \new_[31397]_ ;
  assign \new_[1250]_  = \new_[31384]_  & \new_[31369]_ ;
  assign \new_[1251]_  = \new_[31356]_  & \new_[31341]_ ;
  assign \new_[1252]_  = \new_[31328]_  & \new_[31313]_ ;
  assign \new_[1253]_  = \new_[31300]_  & \new_[31285]_ ;
  assign \new_[1254]_  = \new_[31272]_  & \new_[31257]_ ;
  assign \new_[1255]_  = \new_[31244]_  & \new_[31229]_ ;
  assign \new_[1256]_  = \new_[31216]_  & \new_[31201]_ ;
  assign \new_[1257]_  = \new_[31188]_  & \new_[31173]_ ;
  assign \new_[1258]_  = \new_[31160]_  & \new_[31145]_ ;
  assign \new_[1259]_  = \new_[31132]_  & \new_[31117]_ ;
  assign \new_[1260]_  = \new_[31104]_  & \new_[31089]_ ;
  assign \new_[1261]_  = \new_[31076]_  & \new_[31061]_ ;
  assign \new_[1262]_  = \new_[31048]_  & \new_[31033]_ ;
  assign \new_[1263]_  = \new_[31020]_  & \new_[31005]_ ;
  assign \new_[1264]_  = \new_[30992]_  & \new_[30977]_ ;
  assign \new_[1265]_  = \new_[30964]_  & \new_[30949]_ ;
  assign \new_[1266]_  = \new_[30936]_  & \new_[30921]_ ;
  assign \new_[1267]_  = \new_[30908]_  & \new_[30893]_ ;
  assign \new_[1268]_  = \new_[30880]_  & \new_[30865]_ ;
  assign \new_[1269]_  = \new_[30852]_  & \new_[30837]_ ;
  assign \new_[1270]_  = \new_[30824]_  & \new_[30809]_ ;
  assign \new_[1271]_  = \new_[30796]_  & \new_[30781]_ ;
  assign \new_[1272]_  = \new_[30768]_  & \new_[30753]_ ;
  assign \new_[1273]_  = \new_[30740]_  & \new_[30725]_ ;
  assign \new_[1274]_  = \new_[30712]_  & \new_[30697]_ ;
  assign \new_[1275]_  = \new_[30684]_  & \new_[30669]_ ;
  assign \new_[1276]_  = \new_[30656]_  & \new_[30641]_ ;
  assign \new_[1277]_  = \new_[30628]_  & \new_[30613]_ ;
  assign \new_[1278]_  = \new_[30600]_  & \new_[30585]_ ;
  assign \new_[1279]_  = \new_[30572]_  & \new_[30557]_ ;
  assign \new_[1280]_  = \new_[30544]_  & \new_[30529]_ ;
  assign \new_[1281]_  = \new_[30516]_  & \new_[30501]_ ;
  assign \new_[1282]_  = \new_[30488]_  & \new_[30473]_ ;
  assign \new_[1283]_  = \new_[30460]_  & \new_[30445]_ ;
  assign \new_[1284]_  = \new_[30432]_  & \new_[30417]_ ;
  assign \new_[1285]_  = \new_[30404]_  & \new_[30389]_ ;
  assign \new_[1286]_  = \new_[30376]_  & \new_[30361]_ ;
  assign \new_[1287]_  = \new_[30348]_  & \new_[30333]_ ;
  assign \new_[1288]_  = \new_[30320]_  & \new_[30305]_ ;
  assign \new_[1289]_  = \new_[30292]_  & \new_[30277]_ ;
  assign \new_[1290]_  = \new_[30264]_  & \new_[30249]_ ;
  assign \new_[1291]_  = \new_[30236]_  & \new_[30221]_ ;
  assign \new_[1292]_  = \new_[30208]_  & \new_[30193]_ ;
  assign \new_[1293]_  = \new_[30180]_  & \new_[30165]_ ;
  assign \new_[1294]_  = \new_[30152]_  & \new_[30137]_ ;
  assign \new_[1295]_  = \new_[30124]_  & \new_[30109]_ ;
  assign \new_[1296]_  = \new_[30096]_  & \new_[30081]_ ;
  assign \new_[1297]_  = \new_[30068]_  & \new_[30053]_ ;
  assign \new_[1298]_  = \new_[30040]_  & \new_[30025]_ ;
  assign \new_[1299]_  = \new_[30012]_  & \new_[29997]_ ;
  assign \new_[1300]_  = \new_[29984]_  & \new_[29969]_ ;
  assign \new_[1301]_  = \new_[29956]_  & \new_[29941]_ ;
  assign \new_[1302]_  = \new_[29928]_  & \new_[29913]_ ;
  assign \new_[1303]_  = \new_[29900]_  & \new_[29885]_ ;
  assign \new_[1304]_  = \new_[29872]_  & \new_[29857]_ ;
  assign \new_[1305]_  = \new_[29844]_  & \new_[29829]_ ;
  assign \new_[1306]_  = \new_[29816]_  & \new_[29801]_ ;
  assign \new_[1307]_  = \new_[29788]_  & \new_[29773]_ ;
  assign \new_[1308]_  = \new_[29760]_  & \new_[29745]_ ;
  assign \new_[1309]_  = \new_[29732]_  & \new_[29717]_ ;
  assign \new_[1310]_  = \new_[29704]_  & \new_[29689]_ ;
  assign \new_[1311]_  = \new_[29676]_  & \new_[29661]_ ;
  assign \new_[1312]_  = \new_[29648]_  & \new_[29633]_ ;
  assign \new_[1313]_  = \new_[29620]_  & \new_[29605]_ ;
  assign \new_[1314]_  = \new_[29592]_  & \new_[29577]_ ;
  assign \new_[1315]_  = \new_[29564]_  & \new_[29549]_ ;
  assign \new_[1316]_  = \new_[29536]_  & \new_[29521]_ ;
  assign \new_[1317]_  = \new_[29508]_  & \new_[29493]_ ;
  assign \new_[1318]_  = \new_[29480]_  & \new_[29465]_ ;
  assign \new_[1319]_  = \new_[29452]_  & \new_[29437]_ ;
  assign \new_[1320]_  = \new_[29424]_  & \new_[29409]_ ;
  assign \new_[1321]_  = \new_[29396]_  & \new_[29381]_ ;
  assign \new_[1322]_  = \new_[29368]_  & \new_[29353]_ ;
  assign \new_[1323]_  = \new_[29340]_  & \new_[29325]_ ;
  assign \new_[1324]_  = \new_[29312]_  & \new_[29297]_ ;
  assign \new_[1325]_  = \new_[29284]_  & \new_[29269]_ ;
  assign \new_[1326]_  = \new_[29256]_  & \new_[29241]_ ;
  assign \new_[1327]_  = \new_[29228]_  & \new_[29213]_ ;
  assign \new_[1328]_  = \new_[29200]_  & \new_[29185]_ ;
  assign \new_[1329]_  = \new_[29172]_  & \new_[29157]_ ;
  assign \new_[1330]_  = \new_[29144]_  & \new_[29129]_ ;
  assign \new_[1331]_  = \new_[29116]_  & \new_[29101]_ ;
  assign \new_[1332]_  = \new_[29088]_  & \new_[29073]_ ;
  assign \new_[1333]_  = \new_[29060]_  & \new_[29045]_ ;
  assign \new_[1334]_  = \new_[29032]_  & \new_[29017]_ ;
  assign \new_[1335]_  = \new_[29004]_  & \new_[28989]_ ;
  assign \new_[1336]_  = \new_[28976]_  & \new_[28961]_ ;
  assign \new_[1337]_  = \new_[28948]_  & \new_[28933]_ ;
  assign \new_[1338]_  = \new_[28920]_  & \new_[28905]_ ;
  assign \new_[1339]_  = \new_[28892]_  & \new_[28877]_ ;
  assign \new_[1340]_  = \new_[28864]_  & \new_[28849]_ ;
  assign \new_[1341]_  = \new_[28836]_  & \new_[28821]_ ;
  assign \new_[1342]_  = \new_[28808]_  & \new_[28793]_ ;
  assign \new_[1343]_  = \new_[28780]_  & \new_[28765]_ ;
  assign \new_[1344]_  = \new_[28752]_  & \new_[28737]_ ;
  assign \new_[1345]_  = \new_[28724]_  & \new_[28709]_ ;
  assign \new_[1346]_  = \new_[28696]_  & \new_[28681]_ ;
  assign \new_[1347]_  = \new_[28668]_  & \new_[28653]_ ;
  assign \new_[1348]_  = \new_[28640]_  & \new_[28625]_ ;
  assign \new_[1349]_  = \new_[28612]_  & \new_[28597]_ ;
  assign \new_[1350]_  = \new_[28584]_  & \new_[28569]_ ;
  assign \new_[1351]_  = \new_[28556]_  & \new_[28541]_ ;
  assign \new_[1352]_  = \new_[28528]_  & \new_[28513]_ ;
  assign \new_[1353]_  = \new_[28500]_  & \new_[28485]_ ;
  assign \new_[1354]_  = \new_[28472]_  & \new_[28457]_ ;
  assign \new_[1355]_  = \new_[28444]_  & \new_[28429]_ ;
  assign \new_[1356]_  = \new_[28416]_  & \new_[28401]_ ;
  assign \new_[1357]_  = \new_[28388]_  & \new_[28373]_ ;
  assign \new_[1358]_  = \new_[28360]_  & \new_[28345]_ ;
  assign \new_[1359]_  = \new_[28332]_  & \new_[28317]_ ;
  assign \new_[1360]_  = \new_[28304]_  & \new_[28289]_ ;
  assign \new_[1361]_  = \new_[28276]_  & \new_[28261]_ ;
  assign \new_[1362]_  = \new_[28248]_  & \new_[28233]_ ;
  assign \new_[1363]_  = \new_[28220]_  & \new_[28205]_ ;
  assign \new_[1364]_  = \new_[28192]_  & \new_[28177]_ ;
  assign \new_[1365]_  = \new_[28164]_  & \new_[28149]_ ;
  assign \new_[1366]_  = \new_[28136]_  & \new_[28121]_ ;
  assign \new_[1367]_  = \new_[28108]_  & \new_[28093]_ ;
  assign \new_[1368]_  = \new_[28080]_  & \new_[28065]_ ;
  assign \new_[1369]_  = \new_[28052]_  & \new_[28037]_ ;
  assign \new_[1370]_  = \new_[28024]_  & \new_[28009]_ ;
  assign \new_[1371]_  = \new_[27996]_  & \new_[27981]_ ;
  assign \new_[1372]_  = \new_[27968]_  & \new_[27953]_ ;
  assign \new_[1373]_  = \new_[27940]_  & \new_[27925]_ ;
  assign \new_[1374]_  = \new_[27912]_  & \new_[27897]_ ;
  assign \new_[1375]_  = \new_[27884]_  & \new_[27869]_ ;
  assign \new_[1376]_  = \new_[27856]_  & \new_[27841]_ ;
  assign \new_[1377]_  = \new_[27828]_  & \new_[27813]_ ;
  assign \new_[1378]_  = \new_[27800]_  & \new_[27785]_ ;
  assign \new_[1379]_  = \new_[27772]_  & \new_[27757]_ ;
  assign \new_[1380]_  = \new_[27744]_  & \new_[27729]_ ;
  assign \new_[1381]_  = \new_[27716]_  & \new_[27701]_ ;
  assign \new_[1382]_  = \new_[27688]_  & \new_[27673]_ ;
  assign \new_[1383]_  = \new_[27660]_  & \new_[27645]_ ;
  assign \new_[1384]_  = \new_[27632]_  & \new_[27617]_ ;
  assign \new_[1385]_  = \new_[27604]_  & \new_[27589]_ ;
  assign \new_[1386]_  = \new_[27576]_  & \new_[27561]_ ;
  assign \new_[1387]_  = \new_[27548]_  & \new_[27533]_ ;
  assign \new_[1388]_  = \new_[27520]_  & \new_[27505]_ ;
  assign \new_[1389]_  = \new_[27492]_  & \new_[27477]_ ;
  assign \new_[1390]_  = \new_[27464]_  & \new_[27449]_ ;
  assign \new_[1391]_  = \new_[27436]_  & \new_[27421]_ ;
  assign \new_[1392]_  = \new_[27408]_  & \new_[27393]_ ;
  assign \new_[1393]_  = \new_[27380]_  & \new_[27365]_ ;
  assign \new_[1394]_  = \new_[27352]_  & \new_[27337]_ ;
  assign \new_[1395]_  = \new_[27324]_  & \new_[27309]_ ;
  assign \new_[1396]_  = \new_[27296]_  & \new_[27281]_ ;
  assign \new_[1397]_  = \new_[27268]_  & \new_[27253]_ ;
  assign \new_[1398]_  = \new_[27240]_  & \new_[27225]_ ;
  assign \new_[1399]_  = \new_[27212]_  & \new_[27197]_ ;
  assign \new_[1400]_  = \new_[27184]_  & \new_[27169]_ ;
  assign \new_[1401]_  = \new_[27156]_  & \new_[27141]_ ;
  assign \new_[1402]_  = \new_[27128]_  & \new_[27113]_ ;
  assign \new_[1403]_  = \new_[27100]_  & \new_[27085]_ ;
  assign \new_[1404]_  = \new_[27072]_  & \new_[27057]_ ;
  assign \new_[1405]_  = \new_[27044]_  & \new_[27029]_ ;
  assign \new_[1406]_  = \new_[27016]_  & \new_[27001]_ ;
  assign \new_[1407]_  = \new_[26988]_  & \new_[26973]_ ;
  assign \new_[1408]_  = \new_[26960]_  & \new_[26945]_ ;
  assign \new_[1409]_  = \new_[26932]_  & \new_[26917]_ ;
  assign \new_[1410]_  = \new_[26904]_  & \new_[26889]_ ;
  assign \new_[1411]_  = \new_[26876]_  & \new_[26861]_ ;
  assign \new_[1412]_  = \new_[26848]_  & \new_[26833]_ ;
  assign \new_[1413]_  = \new_[26820]_  & \new_[26805]_ ;
  assign \new_[1414]_  = \new_[26792]_  & \new_[26777]_ ;
  assign \new_[1415]_  = \new_[26764]_  & \new_[26749]_ ;
  assign \new_[1416]_  = \new_[26736]_  & \new_[26721]_ ;
  assign \new_[1417]_  = \new_[26708]_  & \new_[26693]_ ;
  assign \new_[1418]_  = \new_[26680]_  & \new_[26665]_ ;
  assign \new_[1419]_  = \new_[26652]_  & \new_[26637]_ ;
  assign \new_[1420]_  = \new_[26624]_  & \new_[26609]_ ;
  assign \new_[1421]_  = \new_[26596]_  & \new_[26581]_ ;
  assign \new_[1422]_  = \new_[26568]_  & \new_[26553]_ ;
  assign \new_[1423]_  = \new_[26540]_  & \new_[26525]_ ;
  assign \new_[1424]_  = \new_[26512]_  & \new_[26497]_ ;
  assign \new_[1425]_  = \new_[26484]_  & \new_[26469]_ ;
  assign \new_[1426]_  = \new_[26456]_  & \new_[26441]_ ;
  assign \new_[1427]_  = \new_[26428]_  & \new_[26413]_ ;
  assign \new_[1428]_  = \new_[26400]_  & \new_[26385]_ ;
  assign \new_[1429]_  = \new_[26372]_  & \new_[26357]_ ;
  assign \new_[1430]_  = \new_[26344]_  & \new_[26329]_ ;
  assign \new_[1431]_  = \new_[26316]_  & \new_[26301]_ ;
  assign \new_[1432]_  = \new_[26288]_  & \new_[26273]_ ;
  assign \new_[1433]_  = \new_[26260]_  & \new_[26245]_ ;
  assign \new_[1434]_  = \new_[26232]_  & \new_[26217]_ ;
  assign \new_[1435]_  = \new_[26204]_  & \new_[26189]_ ;
  assign \new_[1436]_  = \new_[26176]_  & \new_[26161]_ ;
  assign \new_[1437]_  = \new_[26148]_  & \new_[26133]_ ;
  assign \new_[1438]_  = \new_[26120]_  & \new_[26105]_ ;
  assign \new_[1439]_  = \new_[26092]_  & \new_[26077]_ ;
  assign \new_[1440]_  = \new_[26064]_  & \new_[26049]_ ;
  assign \new_[1441]_  = \new_[26036]_  & \new_[26021]_ ;
  assign \new_[1442]_  = \new_[26008]_  & \new_[25993]_ ;
  assign \new_[1443]_  = \new_[25980]_  & \new_[25965]_ ;
  assign \new_[1444]_  = \new_[25952]_  & \new_[25937]_ ;
  assign \new_[1445]_  = \new_[25924]_  & \new_[25909]_ ;
  assign \new_[1446]_  = \new_[25896]_  & \new_[25881]_ ;
  assign \new_[1447]_  = \new_[25868]_  & \new_[25853]_ ;
  assign \new_[1448]_  = \new_[25840]_  & \new_[25825]_ ;
  assign \new_[1449]_  = \new_[25812]_  & \new_[25797]_ ;
  assign \new_[1450]_  = \new_[25784]_  & \new_[25769]_ ;
  assign \new_[1451]_  = \new_[25756]_  & \new_[25741]_ ;
  assign \new_[1452]_  = \new_[25728]_  & \new_[25713]_ ;
  assign \new_[1453]_  = \new_[25700]_  & \new_[25685]_ ;
  assign \new_[1454]_  = \new_[25672]_  & \new_[25657]_ ;
  assign \new_[1455]_  = \new_[25644]_  & \new_[25629]_ ;
  assign \new_[1456]_  = \new_[25616]_  & \new_[25601]_ ;
  assign \new_[1457]_  = \new_[25588]_  & \new_[25573]_ ;
  assign \new_[1458]_  = \new_[25560]_  & \new_[25545]_ ;
  assign \new_[1459]_  = \new_[25532]_  & \new_[25517]_ ;
  assign \new_[1460]_  = \new_[25504]_  & \new_[25489]_ ;
  assign \new_[1461]_  = \new_[25476]_  & \new_[25461]_ ;
  assign \new_[1462]_  = \new_[25448]_  & \new_[25433]_ ;
  assign \new_[1463]_  = \new_[25420]_  & \new_[25405]_ ;
  assign \new_[1464]_  = \new_[25392]_  & \new_[25377]_ ;
  assign \new_[1465]_  = \new_[25364]_  & \new_[25349]_ ;
  assign \new_[1466]_  = \new_[25336]_  & \new_[25321]_ ;
  assign \new_[1467]_  = \new_[25308]_  & \new_[25293]_ ;
  assign \new_[1468]_  = \new_[25280]_  & \new_[25265]_ ;
  assign \new_[1469]_  = \new_[25252]_  & \new_[25237]_ ;
  assign \new_[1470]_  = \new_[25224]_  & \new_[25209]_ ;
  assign \new_[1471]_  = \new_[25196]_  & \new_[25181]_ ;
  assign \new_[1472]_  = \new_[25168]_  & \new_[25153]_ ;
  assign \new_[1473]_  = \new_[25140]_  & \new_[25125]_ ;
  assign \new_[1474]_  = \new_[25112]_  & \new_[25097]_ ;
  assign \new_[1475]_  = \new_[25084]_  & \new_[25069]_ ;
  assign \new_[1476]_  = \new_[25056]_  & \new_[25041]_ ;
  assign \new_[1477]_  = \new_[25028]_  & \new_[25013]_ ;
  assign \new_[1478]_  = \new_[25000]_  & \new_[24985]_ ;
  assign \new_[1479]_  = \new_[24972]_  & \new_[24957]_ ;
  assign \new_[1480]_  = \new_[24944]_  & \new_[24929]_ ;
  assign \new_[1481]_  = \new_[24916]_  & \new_[24901]_ ;
  assign \new_[1482]_  = \new_[24888]_  & \new_[24873]_ ;
  assign \new_[1483]_  = \new_[24860]_  & \new_[24845]_ ;
  assign \new_[1484]_  = \new_[24832]_  & \new_[24817]_ ;
  assign \new_[1485]_  = \new_[24804]_  & \new_[24789]_ ;
  assign \new_[1486]_  = \new_[24776]_  & \new_[24761]_ ;
  assign \new_[1487]_  = \new_[24748]_  & \new_[24733]_ ;
  assign \new_[1488]_  = \new_[24720]_  & \new_[24705]_ ;
  assign \new_[1489]_  = \new_[24692]_  & \new_[24677]_ ;
  assign \new_[1490]_  = \new_[24664]_  & \new_[24649]_ ;
  assign \new_[1491]_  = \new_[24636]_  & \new_[24621]_ ;
  assign \new_[1492]_  = \new_[24608]_  & \new_[24593]_ ;
  assign \new_[1493]_  = \new_[24580]_  & \new_[24565]_ ;
  assign \new_[1494]_  = \new_[24552]_  & \new_[24537]_ ;
  assign \new_[1495]_  = \new_[24524]_  & \new_[24509]_ ;
  assign \new_[1496]_  = \new_[24496]_  & \new_[24481]_ ;
  assign \new_[1497]_  = \new_[24468]_  & \new_[24453]_ ;
  assign \new_[1498]_  = \new_[24440]_  & \new_[24425]_ ;
  assign \new_[1499]_  = \new_[24412]_  & \new_[24397]_ ;
  assign \new_[1500]_  = \new_[24384]_  & \new_[24369]_ ;
  assign \new_[1501]_  = \new_[24356]_  & \new_[24341]_ ;
  assign \new_[1502]_  = \new_[24328]_  & \new_[24313]_ ;
  assign \new_[1503]_  = \new_[24300]_  & \new_[24285]_ ;
  assign \new_[1504]_  = \new_[24272]_  & \new_[24257]_ ;
  assign \new_[1505]_  = \new_[24244]_  & \new_[24229]_ ;
  assign \new_[1506]_  = \new_[24216]_  & \new_[24201]_ ;
  assign \new_[1507]_  = \new_[24188]_  & \new_[24173]_ ;
  assign \new_[1508]_  = \new_[24160]_  & \new_[24145]_ ;
  assign \new_[1509]_  = \new_[24132]_  & \new_[24117]_ ;
  assign \new_[1510]_  = \new_[24104]_  & \new_[24089]_ ;
  assign \new_[1511]_  = \new_[24076]_  & \new_[24061]_ ;
  assign \new_[1512]_  = \new_[24048]_  & \new_[24033]_ ;
  assign \new_[1513]_  = \new_[24020]_  & \new_[24005]_ ;
  assign \new_[1514]_  = \new_[23992]_  & \new_[23977]_ ;
  assign \new_[1515]_  = \new_[23964]_  & \new_[23949]_ ;
  assign \new_[1516]_  = \new_[23936]_  & \new_[23921]_ ;
  assign \new_[1517]_  = \new_[23908]_  & \new_[23893]_ ;
  assign \new_[1518]_  = \new_[23880]_  & \new_[23865]_ ;
  assign \new_[1519]_  = \new_[23852]_  & \new_[23837]_ ;
  assign \new_[1520]_  = \new_[23824]_  & \new_[23809]_ ;
  assign \new_[1521]_  = \new_[23796]_  & \new_[23781]_ ;
  assign \new_[1522]_  = \new_[23768]_  & \new_[23753]_ ;
  assign \new_[1523]_  = \new_[23740]_  & \new_[23725]_ ;
  assign \new_[1524]_  = \new_[23712]_  & \new_[23697]_ ;
  assign \new_[1525]_  = \new_[23684]_  & \new_[23669]_ ;
  assign \new_[1526]_  = \new_[23656]_  & \new_[23641]_ ;
  assign \new_[1527]_  = \new_[23628]_  & \new_[23613]_ ;
  assign \new_[1528]_  = \new_[23600]_  & \new_[23585]_ ;
  assign \new_[1529]_  = \new_[23572]_  & \new_[23557]_ ;
  assign \new_[1530]_  = \new_[23544]_  & \new_[23529]_ ;
  assign \new_[1531]_  = \new_[23516]_  & \new_[23501]_ ;
  assign \new_[1532]_  = \new_[23488]_  & \new_[23473]_ ;
  assign \new_[1533]_  = \new_[23460]_  & \new_[23445]_ ;
  assign \new_[1534]_  = \new_[23432]_  & \new_[23417]_ ;
  assign \new_[1535]_  = \new_[23404]_  & \new_[23389]_ ;
  assign \new_[1536]_  = \new_[23376]_  & \new_[23361]_ ;
  assign \new_[1537]_  = \new_[23348]_  & \new_[23333]_ ;
  assign \new_[1538]_  = \new_[23320]_  & \new_[23305]_ ;
  assign \new_[1539]_  = \new_[23292]_  & \new_[23277]_ ;
  assign \new_[1540]_  = \new_[23264]_  & \new_[23249]_ ;
  assign \new_[1541]_  = \new_[23236]_  & \new_[23221]_ ;
  assign \new_[1542]_  = \new_[23208]_  & \new_[23193]_ ;
  assign \new_[1543]_  = \new_[23180]_  & \new_[23165]_ ;
  assign \new_[1544]_  = \new_[23152]_  & \new_[23137]_ ;
  assign \new_[1545]_  = \new_[23124]_  & \new_[23109]_ ;
  assign \new_[1546]_  = \new_[23096]_  & \new_[23081]_ ;
  assign \new_[1547]_  = \new_[23068]_  & \new_[23053]_ ;
  assign \new_[1548]_  = \new_[23040]_  & \new_[23025]_ ;
  assign \new_[1549]_  = \new_[23012]_  & \new_[22997]_ ;
  assign \new_[1550]_  = \new_[22984]_  & \new_[22969]_ ;
  assign \new_[1551]_  = \new_[22956]_  & \new_[22941]_ ;
  assign \new_[1552]_  = \new_[22928]_  & \new_[22913]_ ;
  assign \new_[1553]_  = \new_[22900]_  & \new_[22885]_ ;
  assign \new_[1554]_  = \new_[22872]_  & \new_[22857]_ ;
  assign \new_[1555]_  = \new_[22844]_  & \new_[22829]_ ;
  assign \new_[1556]_  = \new_[22816]_  & \new_[22801]_ ;
  assign \new_[1557]_  = \new_[22788]_  & \new_[22773]_ ;
  assign \new_[1558]_  = \new_[22760]_  & \new_[22745]_ ;
  assign \new_[1559]_  = \new_[22732]_  & \new_[22717]_ ;
  assign \new_[1560]_  = \new_[22704]_  & \new_[22689]_ ;
  assign \new_[1561]_  = \new_[22676]_  & \new_[22661]_ ;
  assign \new_[1562]_  = \new_[22648]_  & \new_[22633]_ ;
  assign \new_[1563]_  = \new_[22620]_  & \new_[22605]_ ;
  assign \new_[1564]_  = \new_[22592]_  & \new_[22577]_ ;
  assign \new_[1565]_  = \new_[22564]_  & \new_[22549]_ ;
  assign \new_[1566]_  = \new_[22536]_  & \new_[22521]_ ;
  assign \new_[1567]_  = \new_[22508]_  & \new_[22493]_ ;
  assign \new_[1568]_  = \new_[22480]_  & \new_[22465]_ ;
  assign \new_[1569]_  = \new_[22452]_  & \new_[22437]_ ;
  assign \new_[1570]_  = \new_[22424]_  & \new_[22409]_ ;
  assign \new_[1571]_  = \new_[22396]_  & \new_[22381]_ ;
  assign \new_[1572]_  = \new_[22368]_  & \new_[22353]_ ;
  assign \new_[1573]_  = \new_[22340]_  & \new_[22325]_ ;
  assign \new_[1574]_  = \new_[22312]_  & \new_[22297]_ ;
  assign \new_[1575]_  = \new_[22284]_  & \new_[22269]_ ;
  assign \new_[1576]_  = \new_[22256]_  & \new_[22241]_ ;
  assign \new_[1577]_  = \new_[22228]_  & \new_[22213]_ ;
  assign \new_[1578]_  = \new_[22200]_  & \new_[22185]_ ;
  assign \new_[1579]_  = \new_[22172]_  & \new_[22157]_ ;
  assign \new_[1580]_  = \new_[22144]_  & \new_[22129]_ ;
  assign \new_[1581]_  = \new_[22116]_  & \new_[22101]_ ;
  assign \new_[1582]_  = \new_[22088]_  & \new_[22073]_ ;
  assign \new_[1583]_  = \new_[22060]_  & \new_[22045]_ ;
  assign \new_[1584]_  = \new_[22032]_  & \new_[22017]_ ;
  assign \new_[1585]_  = \new_[22004]_  & \new_[21989]_ ;
  assign \new_[1586]_  = \new_[21976]_  & \new_[21961]_ ;
  assign \new_[1587]_  = \new_[21948]_  & \new_[21933]_ ;
  assign \new_[1588]_  = \new_[21920]_  & \new_[21905]_ ;
  assign \new_[1589]_  = \new_[21892]_  & \new_[21877]_ ;
  assign \new_[1590]_  = \new_[21864]_  & \new_[21849]_ ;
  assign \new_[1591]_  = \new_[21836]_  & \new_[21821]_ ;
  assign \new_[1592]_  = \new_[21808]_  & \new_[21793]_ ;
  assign \new_[1593]_  = \new_[21780]_  & \new_[21765]_ ;
  assign \new_[1594]_  = \new_[21752]_  & \new_[21737]_ ;
  assign \new_[1595]_  = \new_[21724]_  & \new_[21709]_ ;
  assign \new_[1596]_  = \new_[21696]_  & \new_[21681]_ ;
  assign \new_[1597]_  = \new_[21668]_  & \new_[21653]_ ;
  assign \new_[1598]_  = \new_[21640]_  & \new_[21625]_ ;
  assign \new_[1599]_  = \new_[21612]_  & \new_[21597]_ ;
  assign \new_[1600]_  = \new_[21584]_  & \new_[21569]_ ;
  assign \new_[1601]_  = \new_[21556]_  & \new_[21541]_ ;
  assign \new_[1602]_  = \new_[21528]_  & \new_[21513]_ ;
  assign \new_[1603]_  = \new_[21500]_  & \new_[21485]_ ;
  assign \new_[1604]_  = \new_[21472]_  & \new_[21457]_ ;
  assign \new_[1605]_  = \new_[21444]_  & \new_[21429]_ ;
  assign \new_[1606]_  = \new_[21416]_  & \new_[21401]_ ;
  assign \new_[1607]_  = \new_[21388]_  & \new_[21373]_ ;
  assign \new_[1608]_  = \new_[21360]_  & \new_[21345]_ ;
  assign \new_[1609]_  = \new_[21332]_  & \new_[21317]_ ;
  assign \new_[1610]_  = \new_[21304]_  & \new_[21289]_ ;
  assign \new_[1611]_  = \new_[21276]_  & \new_[21261]_ ;
  assign \new_[1612]_  = \new_[21248]_  & \new_[21233]_ ;
  assign \new_[1613]_  = \new_[21220]_  & \new_[21205]_ ;
  assign \new_[1614]_  = \new_[21192]_  & \new_[21177]_ ;
  assign \new_[1615]_  = \new_[21164]_  & \new_[21149]_ ;
  assign \new_[1616]_  = \new_[21136]_  & \new_[21121]_ ;
  assign \new_[1617]_  = \new_[21108]_  & \new_[21093]_ ;
  assign \new_[1618]_  = \new_[21080]_  & \new_[21065]_ ;
  assign \new_[1619]_  = \new_[21052]_  & \new_[21037]_ ;
  assign \new_[1620]_  = \new_[21024]_  & \new_[21009]_ ;
  assign \new_[1621]_  = \new_[20996]_  & \new_[20981]_ ;
  assign \new_[1622]_  = \new_[20968]_  & \new_[20953]_ ;
  assign \new_[1623]_  = \new_[20940]_  & \new_[20925]_ ;
  assign \new_[1624]_  = \new_[20912]_  & \new_[20897]_ ;
  assign \new_[1625]_  = \new_[20884]_  & \new_[20869]_ ;
  assign \new_[1626]_  = \new_[20856]_  & \new_[20841]_ ;
  assign \new_[1627]_  = \new_[20828]_  & \new_[20813]_ ;
  assign \new_[1628]_  = \new_[20800]_  & \new_[20785]_ ;
  assign \new_[1629]_  = \new_[20772]_  & \new_[20757]_ ;
  assign \new_[1630]_  = \new_[20744]_  & \new_[20729]_ ;
  assign \new_[1631]_  = \new_[20716]_  & \new_[20701]_ ;
  assign \new_[1632]_  = \new_[20688]_  & \new_[20673]_ ;
  assign \new_[1633]_  = \new_[20660]_  & \new_[20645]_ ;
  assign \new_[1634]_  = \new_[20632]_  & \new_[20617]_ ;
  assign \new_[1635]_  = \new_[20604]_  & \new_[20589]_ ;
  assign \new_[1636]_  = \new_[20576]_  & \new_[20561]_ ;
  assign \new_[1637]_  = \new_[20548]_  & \new_[20533]_ ;
  assign \new_[1638]_  = \new_[20520]_  & \new_[20505]_ ;
  assign \new_[1639]_  = \new_[20492]_  & \new_[20477]_ ;
  assign \new_[1640]_  = \new_[20464]_  & \new_[20449]_ ;
  assign \new_[1641]_  = \new_[20436]_  & \new_[20421]_ ;
  assign \new_[1642]_  = \new_[20408]_  & \new_[20393]_ ;
  assign \new_[1643]_  = \new_[20380]_  & \new_[20365]_ ;
  assign \new_[1644]_  = \new_[20352]_  & \new_[20337]_ ;
  assign \new_[1645]_  = \new_[20324]_  & \new_[20309]_ ;
  assign \new_[1646]_  = \new_[20296]_  & \new_[20281]_ ;
  assign \new_[1647]_  = \new_[20268]_  & \new_[20253]_ ;
  assign \new_[1648]_  = \new_[20240]_  & \new_[20225]_ ;
  assign \new_[1649]_  = \new_[20212]_  & \new_[20199]_ ;
  assign \new_[1650]_  = \new_[20186]_  & \new_[20173]_ ;
  assign \new_[1651]_  = \new_[20160]_  & \new_[20147]_ ;
  assign \new_[1652]_  = \new_[20134]_  & \new_[20121]_ ;
  assign \new_[1653]_  = \new_[20108]_  & \new_[20095]_ ;
  assign \new_[1654]_  = \new_[20082]_  & \new_[20069]_ ;
  assign \new_[1655]_  = \new_[20056]_  & \new_[20043]_ ;
  assign \new_[1656]_  = \new_[20030]_  & \new_[20017]_ ;
  assign \new_[1657]_  = \new_[20004]_  & \new_[19991]_ ;
  assign \new_[1658]_  = \new_[19978]_  & \new_[19965]_ ;
  assign \new_[1659]_  = \new_[19952]_  & \new_[19939]_ ;
  assign \new_[1660]_  = \new_[19926]_  & \new_[19913]_ ;
  assign \new_[1661]_  = \new_[19900]_  & \new_[19887]_ ;
  assign \new_[1662]_  = \new_[19874]_  & \new_[19861]_ ;
  assign \new_[1663]_  = \new_[19848]_  & \new_[19835]_ ;
  assign \new_[1664]_  = \new_[19822]_  & \new_[19809]_ ;
  assign \new_[1665]_  = \new_[19796]_  & \new_[19783]_ ;
  assign \new_[1666]_  = \new_[19770]_  & \new_[19757]_ ;
  assign \new_[1667]_  = \new_[19744]_  & \new_[19731]_ ;
  assign \new_[1668]_  = \new_[19718]_  & \new_[19705]_ ;
  assign \new_[1669]_  = \new_[19692]_  & \new_[19679]_ ;
  assign \new_[1670]_  = \new_[19666]_  & \new_[19653]_ ;
  assign \new_[1671]_  = \new_[19640]_  & \new_[19627]_ ;
  assign \new_[1672]_  = \new_[19614]_  & \new_[19601]_ ;
  assign \new_[1673]_  = \new_[19588]_  & \new_[19575]_ ;
  assign \new_[1674]_  = \new_[19562]_  & \new_[19549]_ ;
  assign \new_[1675]_  = \new_[19536]_  & \new_[19523]_ ;
  assign \new_[1676]_  = \new_[19510]_  & \new_[19497]_ ;
  assign \new_[1677]_  = \new_[19484]_  & \new_[19471]_ ;
  assign \new_[1678]_  = \new_[19458]_  & \new_[19445]_ ;
  assign \new_[1679]_  = \new_[19432]_  & \new_[19419]_ ;
  assign \new_[1680]_  = \new_[19406]_  & \new_[19393]_ ;
  assign \new_[1681]_  = \new_[19380]_  & \new_[19367]_ ;
  assign \new_[1682]_  = \new_[19354]_  & \new_[19341]_ ;
  assign \new_[1683]_  = \new_[19328]_  & \new_[19315]_ ;
  assign \new_[1684]_  = \new_[19302]_  & \new_[19289]_ ;
  assign \new_[1685]_  = \new_[19276]_  & \new_[19263]_ ;
  assign \new_[1686]_  = \new_[19250]_  & \new_[19237]_ ;
  assign \new_[1687]_  = \new_[19224]_  & \new_[19211]_ ;
  assign \new_[1688]_  = \new_[19198]_  & \new_[19185]_ ;
  assign \new_[1689]_  = \new_[19172]_  & \new_[19159]_ ;
  assign \new_[1690]_  = \new_[19146]_  & \new_[19133]_ ;
  assign \new_[1691]_  = \new_[19120]_  & \new_[19107]_ ;
  assign \new_[1692]_  = \new_[19094]_  & \new_[19081]_ ;
  assign \new_[1693]_  = \new_[19068]_  & \new_[19055]_ ;
  assign \new_[1694]_  = \new_[19042]_  & \new_[19029]_ ;
  assign \new_[1695]_  = \new_[19016]_  & \new_[19003]_ ;
  assign \new_[1696]_  = \new_[18990]_  & \new_[18977]_ ;
  assign \new_[1697]_  = \new_[18964]_  & \new_[18951]_ ;
  assign \new_[1698]_  = \new_[18938]_  & \new_[18925]_ ;
  assign \new_[1699]_  = \new_[18912]_  & \new_[18899]_ ;
  assign \new_[1700]_  = \new_[18886]_  & \new_[18873]_ ;
  assign \new_[1701]_  = \new_[18860]_  & \new_[18847]_ ;
  assign \new_[1702]_  = \new_[18834]_  & \new_[18821]_ ;
  assign \new_[1703]_  = \new_[18808]_  & \new_[18795]_ ;
  assign \new_[1704]_  = \new_[18782]_  & \new_[18769]_ ;
  assign \new_[1705]_  = \new_[18756]_  & \new_[18743]_ ;
  assign \new_[1706]_  = \new_[18730]_  & \new_[18717]_ ;
  assign \new_[1707]_  = \new_[18704]_  & \new_[18691]_ ;
  assign \new_[1708]_  = \new_[18678]_  & \new_[18665]_ ;
  assign \new_[1709]_  = \new_[18652]_  & \new_[18639]_ ;
  assign \new_[1710]_  = \new_[18626]_  & \new_[18613]_ ;
  assign \new_[1711]_  = \new_[18600]_  & \new_[18587]_ ;
  assign \new_[1712]_  = \new_[18574]_  & \new_[18561]_ ;
  assign \new_[1713]_  = \new_[18548]_  & \new_[18535]_ ;
  assign \new_[1714]_  = \new_[18522]_  & \new_[18509]_ ;
  assign \new_[1715]_  = \new_[18496]_  & \new_[18483]_ ;
  assign \new_[1716]_  = \new_[18470]_  & \new_[18457]_ ;
  assign \new_[1717]_  = \new_[18444]_  & \new_[18431]_ ;
  assign \new_[1718]_  = \new_[18418]_  & \new_[18405]_ ;
  assign \new_[1719]_  = \new_[18392]_  & \new_[18379]_ ;
  assign \new_[1720]_  = \new_[18366]_  & \new_[18353]_ ;
  assign \new_[1721]_  = \new_[18340]_  & \new_[18327]_ ;
  assign \new_[1722]_  = \new_[18314]_  & \new_[18301]_ ;
  assign \new_[1723]_  = \new_[18288]_  & \new_[18275]_ ;
  assign \new_[1724]_  = \new_[18262]_  & \new_[18249]_ ;
  assign \new_[1725]_  = \new_[18236]_  & \new_[18223]_ ;
  assign \new_[1726]_  = \new_[18210]_  & \new_[18197]_ ;
  assign \new_[1727]_  = \new_[18184]_  & \new_[18171]_ ;
  assign \new_[1728]_  = \new_[18158]_  & \new_[18145]_ ;
  assign \new_[1729]_  = \new_[18132]_  & \new_[18119]_ ;
  assign \new_[1730]_  = \new_[18106]_  & \new_[18093]_ ;
  assign \new_[1731]_  = \new_[18080]_  & \new_[18067]_ ;
  assign \new_[1732]_  = \new_[18054]_  & \new_[18041]_ ;
  assign \new_[1733]_  = \new_[18028]_  & \new_[18015]_ ;
  assign \new_[1734]_  = \new_[18002]_  & \new_[17989]_ ;
  assign \new_[1735]_  = \new_[17976]_  & \new_[17963]_ ;
  assign \new_[1736]_  = \new_[17950]_  & \new_[17937]_ ;
  assign \new_[1737]_  = \new_[17924]_  & \new_[17911]_ ;
  assign \new_[1738]_  = \new_[17898]_  & \new_[17885]_ ;
  assign \new_[1739]_  = \new_[17872]_  & \new_[17859]_ ;
  assign \new_[1740]_  = \new_[17846]_  & \new_[17833]_ ;
  assign \new_[1741]_  = \new_[17820]_  & \new_[17807]_ ;
  assign \new_[1742]_  = \new_[17794]_  & \new_[17781]_ ;
  assign \new_[1743]_  = \new_[17768]_  & \new_[17755]_ ;
  assign \new_[1744]_  = \new_[17742]_  & \new_[17729]_ ;
  assign \new_[1745]_  = \new_[17716]_  & \new_[17703]_ ;
  assign \new_[1746]_  = \new_[17690]_  & \new_[17677]_ ;
  assign \new_[1747]_  = \new_[17664]_  & \new_[17651]_ ;
  assign \new_[1748]_  = \new_[17638]_  & \new_[17625]_ ;
  assign \new_[1749]_  = \new_[17612]_  & \new_[17599]_ ;
  assign \new_[1750]_  = \new_[17586]_  & \new_[17573]_ ;
  assign \new_[1751]_  = \new_[17560]_  & \new_[17547]_ ;
  assign \new_[1752]_  = \new_[17534]_  & \new_[17521]_ ;
  assign \new_[1753]_  = \new_[17508]_  & \new_[17495]_ ;
  assign \new_[1754]_  = \new_[17482]_  & \new_[17469]_ ;
  assign \new_[1755]_  = \new_[17456]_  & \new_[17443]_ ;
  assign \new_[1756]_  = \new_[17430]_  & \new_[17417]_ ;
  assign \new_[1757]_  = \new_[17404]_  & \new_[17391]_ ;
  assign \new_[1758]_  = \new_[17378]_  & \new_[17365]_ ;
  assign \new_[1759]_  = \new_[17352]_  & \new_[17339]_ ;
  assign \new_[1760]_  = \new_[17326]_  & \new_[17313]_ ;
  assign \new_[1761]_  = \new_[17300]_  & \new_[17287]_ ;
  assign \new_[1762]_  = \new_[17274]_  & \new_[17261]_ ;
  assign \new_[1763]_  = \new_[17248]_  & \new_[17235]_ ;
  assign \new_[1764]_  = \new_[17222]_  & \new_[17209]_ ;
  assign \new_[1765]_  = \new_[17196]_  & \new_[17183]_ ;
  assign \new_[1766]_  = \new_[17170]_  & \new_[17157]_ ;
  assign \new_[1767]_  = \new_[17144]_  & \new_[17131]_ ;
  assign \new_[1768]_  = \new_[17118]_  & \new_[17105]_ ;
  assign \new_[1769]_  = \new_[17092]_  & \new_[17079]_ ;
  assign \new_[1770]_  = \new_[17066]_  & \new_[17053]_ ;
  assign \new_[1771]_  = \new_[17040]_  & \new_[17027]_ ;
  assign \new_[1772]_  = \new_[17014]_  & \new_[17001]_ ;
  assign \new_[1773]_  = \new_[16988]_  & \new_[16975]_ ;
  assign \new_[1774]_  = \new_[16962]_  & \new_[16949]_ ;
  assign \new_[1775]_  = \new_[16936]_  & \new_[16923]_ ;
  assign \new_[1776]_  = \new_[16910]_  & \new_[16897]_ ;
  assign \new_[1777]_  = \new_[16884]_  & \new_[16871]_ ;
  assign \new_[1778]_  = \new_[16858]_  & \new_[16845]_ ;
  assign \new_[1779]_  = \new_[16832]_  & \new_[16819]_ ;
  assign \new_[1780]_  = \new_[16806]_  & \new_[16793]_ ;
  assign \new_[1781]_  = \new_[16780]_  & \new_[16767]_ ;
  assign \new_[1782]_  = \new_[16754]_  & \new_[16741]_ ;
  assign \new_[1783]_  = \new_[16728]_  & \new_[16715]_ ;
  assign \new_[1784]_  = \new_[16702]_  & \new_[16689]_ ;
  assign \new_[1785]_  = \new_[16676]_  & \new_[16663]_ ;
  assign \new_[1786]_  = \new_[16650]_  & \new_[16637]_ ;
  assign \new_[1787]_  = \new_[16624]_  & \new_[16611]_ ;
  assign \new_[1788]_  = \new_[16598]_  & \new_[16585]_ ;
  assign \new_[1789]_  = \new_[16572]_  & \new_[16559]_ ;
  assign \new_[1790]_  = \new_[16546]_  & \new_[16533]_ ;
  assign \new_[1791]_  = \new_[16520]_  & \new_[16507]_ ;
  assign \new_[1792]_  = \new_[16494]_  & \new_[16481]_ ;
  assign \new_[1793]_  = \new_[16468]_  & \new_[16455]_ ;
  assign \new_[1794]_  = \new_[16442]_  & \new_[16429]_ ;
  assign \new_[1795]_  = \new_[16416]_  & \new_[16403]_ ;
  assign \new_[1796]_  = \new_[16390]_  & \new_[16377]_ ;
  assign \new_[1797]_  = \new_[16364]_  & \new_[16351]_ ;
  assign \new_[1798]_  = \new_[16338]_  & \new_[16325]_ ;
  assign \new_[1799]_  = \new_[16312]_  & \new_[16299]_ ;
  assign \new_[1800]_  = \new_[16286]_  & \new_[16273]_ ;
  assign \new_[1801]_  = \new_[16260]_  & \new_[16247]_ ;
  assign \new_[1802]_  = \new_[16234]_  & \new_[16221]_ ;
  assign \new_[1803]_  = \new_[16208]_  & \new_[16195]_ ;
  assign \new_[1804]_  = \new_[16182]_  & \new_[16169]_ ;
  assign \new_[1805]_  = \new_[16156]_  & \new_[16143]_ ;
  assign \new_[1806]_  = \new_[16130]_  & \new_[16117]_ ;
  assign \new_[1807]_  = \new_[16104]_  & \new_[16091]_ ;
  assign \new_[1808]_  = \new_[16078]_  & \new_[16065]_ ;
  assign \new_[1809]_  = \new_[16052]_  & \new_[16039]_ ;
  assign \new_[1810]_  = \new_[16026]_  & \new_[16013]_ ;
  assign \new_[1811]_  = \new_[16000]_  & \new_[15987]_ ;
  assign \new_[1812]_  = \new_[15974]_  & \new_[15961]_ ;
  assign \new_[1813]_  = \new_[15948]_  & \new_[15935]_ ;
  assign \new_[1814]_  = \new_[15922]_  & \new_[15909]_ ;
  assign \new_[1815]_  = \new_[15896]_  & \new_[15883]_ ;
  assign \new_[1816]_  = \new_[15870]_  & \new_[15857]_ ;
  assign \new_[1817]_  = \new_[15844]_  & \new_[15831]_ ;
  assign \new_[1818]_  = \new_[15818]_  & \new_[15805]_ ;
  assign \new_[1819]_  = \new_[15792]_  & \new_[15779]_ ;
  assign \new_[1820]_  = \new_[15766]_  & \new_[15753]_ ;
  assign \new_[1821]_  = \new_[15740]_  & \new_[15727]_ ;
  assign \new_[1822]_  = \new_[15714]_  & \new_[15701]_ ;
  assign \new_[1823]_  = \new_[15688]_  & \new_[15675]_ ;
  assign \new_[1824]_  = \new_[15662]_  & \new_[15649]_ ;
  assign \new_[1825]_  = \new_[15636]_  & \new_[15623]_ ;
  assign \new_[1826]_  = \new_[15610]_  & \new_[15597]_ ;
  assign \new_[1827]_  = \new_[15584]_  & \new_[15571]_ ;
  assign \new_[1828]_  = \new_[15558]_  & \new_[15545]_ ;
  assign \new_[1829]_  = \new_[15532]_  & \new_[15519]_ ;
  assign \new_[1830]_  = \new_[15506]_  & \new_[15493]_ ;
  assign \new_[1831]_  = \new_[15480]_  & \new_[15467]_ ;
  assign \new_[1832]_  = \new_[15454]_  & \new_[15441]_ ;
  assign \new_[1833]_  = \new_[15428]_  & \new_[15415]_ ;
  assign \new_[1834]_  = \new_[15402]_  & \new_[15389]_ ;
  assign \new_[1835]_  = \new_[15376]_  & \new_[15363]_ ;
  assign \new_[1836]_  = \new_[15350]_  & \new_[15337]_ ;
  assign \new_[1837]_  = \new_[15324]_  & \new_[15311]_ ;
  assign \new_[1838]_  = \new_[15298]_  & \new_[15285]_ ;
  assign \new_[1839]_  = \new_[15272]_  & \new_[15259]_ ;
  assign \new_[1840]_  = \new_[15246]_  & \new_[15233]_ ;
  assign \new_[1841]_  = \new_[15220]_  & \new_[15207]_ ;
  assign \new_[1842]_  = \new_[15194]_  & \new_[15181]_ ;
  assign \new_[1843]_  = \new_[15168]_  & \new_[15155]_ ;
  assign \new_[1844]_  = \new_[15142]_  & \new_[15129]_ ;
  assign \new_[1845]_  = \new_[15116]_  & \new_[15103]_ ;
  assign \new_[1846]_  = \new_[15090]_  & \new_[15077]_ ;
  assign \new_[1847]_  = \new_[15064]_  & \new_[15051]_ ;
  assign \new_[1848]_  = \new_[15038]_  & \new_[15025]_ ;
  assign \new_[1849]_  = \new_[15012]_  & \new_[14999]_ ;
  assign \new_[1850]_  = \new_[14986]_  & \new_[14973]_ ;
  assign \new_[1851]_  = \new_[14960]_  & \new_[14947]_ ;
  assign \new_[1852]_  = \new_[14934]_  & \new_[14921]_ ;
  assign \new_[1853]_  = \new_[14908]_  & \new_[14895]_ ;
  assign \new_[1854]_  = \new_[14882]_  & \new_[14869]_ ;
  assign \new_[1855]_  = \new_[14856]_  & \new_[14843]_ ;
  assign \new_[1856]_  = \new_[14830]_  & \new_[14817]_ ;
  assign \new_[1857]_  = \new_[14804]_  & \new_[14791]_ ;
  assign \new_[1858]_  = \new_[14778]_  & \new_[14765]_ ;
  assign \new_[1859]_  = \new_[14752]_  & \new_[14739]_ ;
  assign \new_[1860]_  = \new_[14726]_  & \new_[14713]_ ;
  assign \new_[1861]_  = \new_[14700]_  & \new_[14687]_ ;
  assign \new_[1862]_  = \new_[14674]_  & \new_[14661]_ ;
  assign \new_[1863]_  = \new_[14648]_  & \new_[14635]_ ;
  assign \new_[1864]_  = \new_[14622]_  & \new_[14609]_ ;
  assign \new_[1865]_  = \new_[14596]_  & \new_[14583]_ ;
  assign \new_[1866]_  = \new_[14570]_  & \new_[14557]_ ;
  assign \new_[1867]_  = \new_[14544]_  & \new_[14531]_ ;
  assign \new_[1868]_  = \new_[14518]_  & \new_[14505]_ ;
  assign \new_[1869]_  = \new_[14492]_  & \new_[14479]_ ;
  assign \new_[1870]_  = \new_[14466]_  & \new_[14453]_ ;
  assign \new_[1871]_  = \new_[14440]_  & \new_[14427]_ ;
  assign \new_[1872]_  = \new_[14414]_  & \new_[14401]_ ;
  assign \new_[1873]_  = \new_[14388]_  & \new_[14375]_ ;
  assign \new_[1874]_  = \new_[14362]_  & \new_[14349]_ ;
  assign \new_[1875]_  = \new_[14336]_  & \new_[14323]_ ;
  assign \new_[1876]_  = \new_[14310]_  & \new_[14297]_ ;
  assign \new_[1877]_  = \new_[14284]_  & \new_[14271]_ ;
  assign \new_[1878]_  = \new_[14258]_  & \new_[14245]_ ;
  assign \new_[1879]_  = \new_[14232]_  & \new_[14219]_ ;
  assign \new_[1880]_  = \new_[14206]_  & \new_[14193]_ ;
  assign \new_[1881]_  = \new_[14180]_  & \new_[14167]_ ;
  assign \new_[1882]_  = \new_[14154]_  & \new_[14141]_ ;
  assign \new_[1883]_  = \new_[14128]_  & \new_[14115]_ ;
  assign \new_[1884]_  = \new_[14102]_  & \new_[14089]_ ;
  assign \new_[1885]_  = \new_[14076]_  & \new_[14063]_ ;
  assign \new_[1886]_  = \new_[14050]_  & \new_[14037]_ ;
  assign \new_[1887]_  = \new_[14024]_  & \new_[14011]_ ;
  assign \new_[1888]_  = \new_[13998]_  & \new_[13985]_ ;
  assign \new_[1889]_  = \new_[13972]_  & \new_[13959]_ ;
  assign \new_[1890]_  = \new_[13946]_  & \new_[13933]_ ;
  assign \new_[1891]_  = \new_[13920]_  & \new_[13907]_ ;
  assign \new_[1892]_  = \new_[13894]_  & \new_[13881]_ ;
  assign \new_[1893]_  = \new_[13868]_  & \new_[13855]_ ;
  assign \new_[1894]_  = \new_[13842]_  & \new_[13829]_ ;
  assign \new_[1895]_  = \new_[13816]_  & \new_[13803]_ ;
  assign \new_[1896]_  = \new_[13790]_  & \new_[13777]_ ;
  assign \new_[1897]_  = \new_[13764]_  & \new_[13751]_ ;
  assign \new_[1898]_  = \new_[13738]_  & \new_[13725]_ ;
  assign \new_[1899]_  = \new_[13712]_  & \new_[13699]_ ;
  assign \new_[1900]_  = \new_[13686]_  & \new_[13673]_ ;
  assign \new_[1901]_  = \new_[13660]_  & \new_[13647]_ ;
  assign \new_[1902]_  = \new_[13634]_  & \new_[13621]_ ;
  assign \new_[1903]_  = \new_[13608]_  & \new_[13595]_ ;
  assign \new_[1904]_  = \new_[13582]_  & \new_[13569]_ ;
  assign \new_[1905]_  = \new_[13556]_  & \new_[13543]_ ;
  assign \new_[1906]_  = \new_[13530]_  & \new_[13517]_ ;
  assign \new_[1907]_  = \new_[13504]_  & \new_[13491]_ ;
  assign \new_[1908]_  = \new_[13478]_  & \new_[13465]_ ;
  assign \new_[1909]_  = \new_[13452]_  & \new_[13439]_ ;
  assign \new_[1910]_  = \new_[13426]_  & \new_[13413]_ ;
  assign \new_[1911]_  = \new_[13400]_  & \new_[13387]_ ;
  assign \new_[1912]_  = \new_[13374]_  & \new_[13361]_ ;
  assign \new_[1913]_  = \new_[13348]_  & \new_[13335]_ ;
  assign \new_[1914]_  = \new_[13322]_  & \new_[13309]_ ;
  assign \new_[1915]_  = \new_[13296]_  & \new_[13283]_ ;
  assign \new_[1916]_  = \new_[13270]_  & \new_[13257]_ ;
  assign \new_[1917]_  = \new_[13244]_  & \new_[13231]_ ;
  assign \new_[1918]_  = \new_[13218]_  & \new_[13205]_ ;
  assign \new_[1919]_  = \new_[13192]_  & \new_[13179]_ ;
  assign \new_[1920]_  = \new_[13166]_  & \new_[13153]_ ;
  assign \new_[1921]_  = \new_[13140]_  & \new_[13127]_ ;
  assign \new_[1922]_  = \new_[13114]_  & \new_[13101]_ ;
  assign \new_[1923]_  = \new_[13088]_  & \new_[13075]_ ;
  assign \new_[1924]_  = \new_[13062]_  & \new_[13049]_ ;
  assign \new_[1925]_  = \new_[13036]_  & \new_[13023]_ ;
  assign \new_[1926]_  = \new_[13010]_  & \new_[12997]_ ;
  assign \new_[1927]_  = \new_[12984]_  & \new_[12971]_ ;
  assign \new_[1928]_  = \new_[12958]_  & \new_[12945]_ ;
  assign \new_[1929]_  = \new_[12932]_  & \new_[12919]_ ;
  assign \new_[1930]_  = \new_[12906]_  & \new_[12893]_ ;
  assign \new_[1931]_  = \new_[12880]_  & \new_[12867]_ ;
  assign \new_[1932]_  = \new_[12854]_  & \new_[12841]_ ;
  assign \new_[1933]_  = \new_[12828]_  & \new_[12815]_ ;
  assign \new_[1934]_  = \new_[12802]_  & \new_[12789]_ ;
  assign \new_[1935]_  = \new_[12776]_  & \new_[12763]_ ;
  assign \new_[1936]_  = \new_[12750]_  & \new_[12737]_ ;
  assign \new_[1937]_  = \new_[12724]_  & \new_[12711]_ ;
  assign \new_[1938]_  = \new_[12698]_  & \new_[12685]_ ;
  assign \new_[1939]_  = \new_[12672]_  & \new_[12659]_ ;
  assign \new_[1940]_  = \new_[12646]_  & \new_[12633]_ ;
  assign \new_[1941]_  = \new_[12620]_  & \new_[12607]_ ;
  assign \new_[1942]_  = \new_[12594]_  & \new_[12581]_ ;
  assign \new_[1943]_  = \new_[12568]_  & \new_[12555]_ ;
  assign \new_[1944]_  = \new_[12542]_  & \new_[12529]_ ;
  assign \new_[1945]_  = \new_[12516]_  & \new_[12503]_ ;
  assign \new_[1946]_  = \new_[12490]_  & \new_[12477]_ ;
  assign \new_[1947]_  = \new_[12464]_  & \new_[12451]_ ;
  assign \new_[1948]_  = \new_[12438]_  & \new_[12425]_ ;
  assign \new_[1949]_  = \new_[12412]_  & \new_[12399]_ ;
  assign \new_[1950]_  = \new_[12386]_  & \new_[12373]_ ;
  assign \new_[1951]_  = \new_[12360]_  & \new_[12347]_ ;
  assign \new_[1952]_  = \new_[12334]_  & \new_[12321]_ ;
  assign \new_[1953]_  = \new_[12308]_  & \new_[12295]_ ;
  assign \new_[1954]_  = \new_[12282]_  & \new_[12269]_ ;
  assign \new_[1955]_  = \new_[12256]_  & \new_[12243]_ ;
  assign \new_[1956]_  = \new_[12230]_  & \new_[12217]_ ;
  assign \new_[1957]_  = \new_[12204]_  & \new_[12191]_ ;
  assign \new_[1958]_  = \new_[12178]_  & \new_[12165]_ ;
  assign \new_[1959]_  = \new_[12152]_  & \new_[12139]_ ;
  assign \new_[1960]_  = \new_[12126]_  & \new_[12113]_ ;
  assign \new_[1961]_  = \new_[12100]_  & \new_[12087]_ ;
  assign \new_[1962]_  = \new_[12074]_  & \new_[12061]_ ;
  assign \new_[1963]_  = \new_[12048]_  & \new_[12035]_ ;
  assign \new_[1964]_  = \new_[12022]_  & \new_[12009]_ ;
  assign \new_[1965]_  = \new_[11996]_  & \new_[11983]_ ;
  assign \new_[1966]_  = \new_[11970]_  & \new_[11957]_ ;
  assign \new_[1967]_  = \new_[11944]_  & \new_[11931]_ ;
  assign \new_[1968]_  = \new_[11918]_  & \new_[11905]_ ;
  assign \new_[1969]_  = \new_[11892]_  & \new_[11879]_ ;
  assign \new_[1970]_  = \new_[11866]_  & \new_[11853]_ ;
  assign \new_[1971]_  = \new_[11840]_  & \new_[11827]_ ;
  assign \new_[1972]_  = \new_[11814]_  & \new_[11801]_ ;
  assign \new_[1973]_  = \new_[11788]_  & \new_[11775]_ ;
  assign \new_[1974]_  = \new_[11762]_  & \new_[11749]_ ;
  assign \new_[1975]_  = \new_[11736]_  & \new_[11723]_ ;
  assign \new_[1976]_  = \new_[11710]_  & \new_[11697]_ ;
  assign \new_[1977]_  = \new_[11684]_  & \new_[11671]_ ;
  assign \new_[1978]_  = \new_[11658]_  & \new_[11645]_ ;
  assign \new_[1979]_  = \new_[11632]_  & \new_[11619]_ ;
  assign \new_[1980]_  = \new_[11606]_  & \new_[11593]_ ;
  assign \new_[1981]_  = \new_[11580]_  & \new_[11567]_ ;
  assign \new_[1982]_  = \new_[11554]_  & \new_[11541]_ ;
  assign \new_[1983]_  = \new_[11528]_  & \new_[11515]_ ;
  assign \new_[1984]_  = \new_[11502]_  & \new_[11489]_ ;
  assign \new_[1985]_  = \new_[11476]_  & \new_[11463]_ ;
  assign \new_[1986]_  = \new_[11450]_  & \new_[11437]_ ;
  assign \new_[1987]_  = \new_[11424]_  & \new_[11411]_ ;
  assign \new_[1988]_  = \new_[11398]_  & \new_[11385]_ ;
  assign \new_[1989]_  = \new_[11372]_  & \new_[11359]_ ;
  assign \new_[1990]_  = \new_[11346]_  & \new_[11333]_ ;
  assign \new_[1991]_  = \new_[11320]_  & \new_[11307]_ ;
  assign \new_[1992]_  = \new_[11294]_  & \new_[11281]_ ;
  assign \new_[1993]_  = \new_[11268]_  & \new_[11255]_ ;
  assign \new_[1994]_  = \new_[11242]_  & \new_[11229]_ ;
  assign \new_[1995]_  = \new_[11216]_  & \new_[11203]_ ;
  assign \new_[1996]_  = \new_[11190]_  & \new_[11177]_ ;
  assign \new_[1997]_  = \new_[11164]_  & \new_[11151]_ ;
  assign \new_[1998]_  = \new_[11138]_  & \new_[11125]_ ;
  assign \new_[1999]_  = \new_[11112]_  & \new_[11099]_ ;
  assign \new_[2000]_  = \new_[11086]_  & \new_[11073]_ ;
  assign \new_[2001]_  = \new_[11060]_  & \new_[11047]_ ;
  assign \new_[2002]_  = \new_[11034]_  & \new_[11021]_ ;
  assign \new_[2003]_  = \new_[11008]_  & \new_[10995]_ ;
  assign \new_[2004]_  = \new_[10982]_  & \new_[10969]_ ;
  assign \new_[2005]_  = \new_[10956]_  & \new_[10943]_ ;
  assign \new_[2006]_  = \new_[10930]_  & \new_[10917]_ ;
  assign \new_[2007]_  = \new_[10904]_  & \new_[10891]_ ;
  assign \new_[2008]_  = \new_[10878]_  & \new_[10865]_ ;
  assign \new_[2009]_  = \new_[10852]_  & \new_[10839]_ ;
  assign \new_[2010]_  = \new_[10826]_  & \new_[10813]_ ;
  assign \new_[2011]_  = \new_[10800]_  & \new_[10787]_ ;
  assign \new_[2012]_  = \new_[10774]_  & \new_[10761]_ ;
  assign \new_[2013]_  = \new_[10748]_  & \new_[10735]_ ;
  assign \new_[2014]_  = \new_[10722]_  & \new_[10709]_ ;
  assign \new_[2015]_  = \new_[10696]_  & \new_[10683]_ ;
  assign \new_[2016]_  = \new_[10670]_  & \new_[10657]_ ;
  assign \new_[2017]_  = \new_[10644]_  & \new_[10631]_ ;
  assign \new_[2018]_  = \new_[10618]_  & \new_[10605]_ ;
  assign \new_[2019]_  = \new_[10592]_  & \new_[10579]_ ;
  assign \new_[2020]_  = \new_[10566]_  & \new_[10553]_ ;
  assign \new_[2021]_  = \new_[10540]_  & \new_[10527]_ ;
  assign \new_[2022]_  = \new_[10514]_  & \new_[10501]_ ;
  assign \new_[2023]_  = \new_[10488]_  & \new_[10475]_ ;
  assign \new_[2024]_  = \new_[10462]_  & \new_[10449]_ ;
  assign \new_[2025]_  = \new_[10436]_  & \new_[10423]_ ;
  assign \new_[2026]_  = \new_[10410]_  & \new_[10397]_ ;
  assign \new_[2027]_  = \new_[10384]_  & \new_[10371]_ ;
  assign \new_[2028]_  = \new_[10358]_  & \new_[10345]_ ;
  assign \new_[2029]_  = \new_[10332]_  & \new_[10319]_ ;
  assign \new_[2030]_  = \new_[10306]_  & \new_[10293]_ ;
  assign \new_[2031]_  = \new_[10280]_  & \new_[10267]_ ;
  assign \new_[2032]_  = \new_[10254]_  & \new_[10241]_ ;
  assign \new_[2033]_  = \new_[10228]_  & \new_[10215]_ ;
  assign \new_[2034]_  = \new_[10202]_  & \new_[10189]_ ;
  assign \new_[2035]_  = \new_[10176]_  & \new_[10163]_ ;
  assign \new_[2036]_  = \new_[10150]_  & \new_[10137]_ ;
  assign \new_[2037]_  = \new_[10124]_  & \new_[10111]_ ;
  assign \new_[2038]_  = \new_[10098]_  & \new_[10085]_ ;
  assign \new_[2039]_  = \new_[10072]_  & \new_[10059]_ ;
  assign \new_[2040]_  = \new_[10046]_  & \new_[10033]_ ;
  assign \new_[2041]_  = \new_[10020]_  & \new_[10007]_ ;
  assign \new_[2042]_  = \new_[9994]_  & \new_[9981]_ ;
  assign \new_[2043]_  = \new_[9968]_  & \new_[9955]_ ;
  assign \new_[2044]_  = \new_[9942]_  & \new_[9929]_ ;
  assign \new_[2045]_  = \new_[9916]_  & \new_[9903]_ ;
  assign \new_[2046]_  = \new_[9890]_  & \new_[9877]_ ;
  assign \new_[2047]_  = \new_[9864]_  & \new_[9851]_ ;
  assign \new_[2048]_  = \new_[9838]_  & \new_[9825]_ ;
  assign \new_[2049]_  = \new_[9812]_  & \new_[9799]_ ;
  assign \new_[2050]_  = \new_[9786]_  & \new_[9773]_ ;
  assign \new_[2051]_  = \new_[9760]_  & \new_[9747]_ ;
  assign \new_[2052]_  = \new_[9734]_  & \new_[9721]_ ;
  assign \new_[2053]_  = \new_[9708]_  & \new_[9695]_ ;
  assign \new_[2054]_  = \new_[9682]_  & \new_[9669]_ ;
  assign \new_[2055]_  = \new_[9656]_  & \new_[9643]_ ;
  assign \new_[2056]_  = \new_[9630]_  & \new_[9617]_ ;
  assign \new_[2057]_  = \new_[9604]_  & \new_[9591]_ ;
  assign \new_[2058]_  = \new_[9578]_  & \new_[9565]_ ;
  assign \new_[2059]_  = \new_[9552]_  & \new_[9539]_ ;
  assign \new_[2060]_  = \new_[9526]_  & \new_[9513]_ ;
  assign \new_[2061]_  = \new_[9500]_  & \new_[9487]_ ;
  assign \new_[2062]_  = \new_[9474]_  & \new_[9461]_ ;
  assign \new_[2063]_  = \new_[9448]_  & \new_[9435]_ ;
  assign \new_[2064]_  = \new_[9422]_  & \new_[9409]_ ;
  assign \new_[2065]_  = \new_[9396]_  & \new_[9383]_ ;
  assign \new_[2066]_  = \new_[9370]_  & \new_[9357]_ ;
  assign \new_[2067]_  = \new_[9344]_  & \new_[9331]_ ;
  assign \new_[2068]_  = \new_[9318]_  & \new_[9305]_ ;
  assign \new_[2069]_  = \new_[9292]_  & \new_[9279]_ ;
  assign \new_[2070]_  = \new_[9266]_  & \new_[9253]_ ;
  assign \new_[2071]_  = \new_[9240]_  & \new_[9227]_ ;
  assign \new_[2072]_  = \new_[9214]_  & \new_[9201]_ ;
  assign \new_[2073]_  = \new_[9188]_  & \new_[9175]_ ;
  assign \new_[2074]_  = \new_[9162]_  & \new_[9149]_ ;
  assign \new_[2075]_  = \new_[9136]_  & \new_[9123]_ ;
  assign \new_[2076]_  = \new_[9110]_  & \new_[9097]_ ;
  assign \new_[2077]_  = \new_[9084]_  & \new_[9071]_ ;
  assign \new_[2078]_  = \new_[9058]_  & \new_[9045]_ ;
  assign \new_[2079]_  = \new_[9032]_  & \new_[9019]_ ;
  assign \new_[2080]_  = \new_[9006]_  & \new_[8993]_ ;
  assign \new_[2081]_  = \new_[8980]_  & \new_[8967]_ ;
  assign \new_[2082]_  = \new_[8954]_  & \new_[8941]_ ;
  assign \new_[2083]_  = \new_[8928]_  & \new_[8915]_ ;
  assign \new_[2084]_  = \new_[8902]_  & \new_[8889]_ ;
  assign \new_[2085]_  = \new_[8876]_  & \new_[8863]_ ;
  assign \new_[2086]_  = \new_[8850]_  & \new_[8837]_ ;
  assign \new_[2087]_  = \new_[8824]_  & \new_[8811]_ ;
  assign \new_[2088]_  = \new_[8798]_  & \new_[8785]_ ;
  assign \new_[2089]_  = \new_[8772]_  & \new_[8759]_ ;
  assign \new_[2090]_  = \new_[8746]_  & \new_[8733]_ ;
  assign \new_[2091]_  = \new_[8720]_  & \new_[8707]_ ;
  assign \new_[2092]_  = \new_[8694]_  & \new_[8681]_ ;
  assign \new_[2093]_  = \new_[8668]_  & \new_[8655]_ ;
  assign \new_[2094]_  = \new_[8642]_  & \new_[8629]_ ;
  assign \new_[2095]_  = \new_[8616]_  & \new_[8603]_ ;
  assign \new_[2096]_  = \new_[8590]_  & \new_[8577]_ ;
  assign \new_[2097]_  = \new_[8564]_  & \new_[8551]_ ;
  assign \new_[2098]_  = \new_[8538]_  & \new_[8525]_ ;
  assign \new_[2099]_  = \new_[8512]_  & \new_[8499]_ ;
  assign \new_[2100]_  = \new_[8486]_  & \new_[8473]_ ;
  assign \new_[2101]_  = \new_[8460]_  & \new_[8447]_ ;
  assign \new_[2102]_  = \new_[8434]_  & \new_[8421]_ ;
  assign \new_[2103]_  = \new_[8408]_  & \new_[8395]_ ;
  assign \new_[2104]_  = \new_[8382]_  & \new_[8369]_ ;
  assign \new_[2105]_  = \new_[8356]_  & \new_[8343]_ ;
  assign \new_[2106]_  = \new_[8330]_  & \new_[8317]_ ;
  assign \new_[2107]_  = \new_[8304]_  & \new_[8291]_ ;
  assign \new_[2108]_  = \new_[8278]_  & \new_[8265]_ ;
  assign \new_[2109]_  = \new_[8252]_  & \new_[8239]_ ;
  assign \new_[2110]_  = \new_[8226]_  & \new_[8213]_ ;
  assign \new_[2111]_  = \new_[8200]_  & \new_[8187]_ ;
  assign \new_[2112]_  = \new_[8174]_  & \new_[8161]_ ;
  assign \new_[2113]_  = \new_[8148]_  & \new_[8135]_ ;
  assign \new_[2114]_  = \new_[8122]_  & \new_[8109]_ ;
  assign \new_[2115]_  = \new_[8096]_  & \new_[8083]_ ;
  assign \new_[2116]_  = \new_[8070]_  & \new_[8057]_ ;
  assign \new_[2117]_  = \new_[8044]_  & \new_[8031]_ ;
  assign \new_[2118]_  = \new_[8018]_  & \new_[8005]_ ;
  assign \new_[2119]_  = \new_[7992]_  & \new_[7979]_ ;
  assign \new_[2120]_  = \new_[7966]_  & \new_[7953]_ ;
  assign \new_[2121]_  = \new_[7940]_  & \new_[7927]_ ;
  assign \new_[2122]_  = \new_[7914]_  & \new_[7901]_ ;
  assign \new_[2123]_  = \new_[7888]_  & \new_[7875]_ ;
  assign \new_[2124]_  = \new_[7862]_  & \new_[7849]_ ;
  assign \new_[2125]_  = \new_[7836]_  & \new_[7823]_ ;
  assign \new_[2126]_  = \new_[7810]_  & \new_[7797]_ ;
  assign \new_[2127]_  = \new_[7784]_  & \new_[7771]_ ;
  assign \new_[2128]_  = \new_[7758]_  & \new_[7745]_ ;
  assign \new_[2129]_  = \new_[7732]_  & \new_[7719]_ ;
  assign \new_[2130]_  = \new_[7706]_  & \new_[7693]_ ;
  assign \new_[2131]_  = \new_[7680]_  & \new_[7667]_ ;
  assign \new_[2132]_  = \new_[7654]_  & \new_[7641]_ ;
  assign \new_[2133]_  = \new_[7628]_  & \new_[7615]_ ;
  assign \new_[2134]_  = \new_[7602]_  & \new_[7589]_ ;
  assign \new_[2135]_  = \new_[7576]_  & \new_[7563]_ ;
  assign \new_[2136]_  = \new_[7550]_  & \new_[7537]_ ;
  assign \new_[2137]_  = \new_[7524]_  & \new_[7511]_ ;
  assign \new_[2138]_  = \new_[7498]_  & \new_[7485]_ ;
  assign \new_[2139]_  = \new_[7472]_  & \new_[7459]_ ;
  assign \new_[2140]_  = \new_[7446]_  & \new_[7433]_ ;
  assign \new_[2141]_  = \new_[7420]_  & \new_[7407]_ ;
  assign \new_[2142]_  = \new_[7394]_  & \new_[7381]_ ;
  assign \new_[2143]_  = \new_[7368]_  & \new_[7355]_ ;
  assign \new_[2144]_  = \new_[7342]_  & \new_[7329]_ ;
  assign \new_[2145]_  = \new_[7316]_  & \new_[7303]_ ;
  assign \new_[2146]_  = \new_[7290]_  & \new_[7277]_ ;
  assign \new_[2147]_  = \new_[7264]_  & \new_[7251]_ ;
  assign \new_[2148]_  = \new_[7238]_  & \new_[7225]_ ;
  assign \new_[2149]_  = \new_[7212]_  & \new_[7199]_ ;
  assign \new_[2150]_  = \new_[7186]_  & \new_[7173]_ ;
  assign \new_[2151]_  = \new_[7160]_  & \new_[7147]_ ;
  assign \new_[2152]_  = \new_[7134]_  & \new_[7121]_ ;
  assign \new_[2153]_  = \new_[7108]_  & \new_[7095]_ ;
  assign \new_[2154]_  = \new_[7082]_  & \new_[7069]_ ;
  assign \new_[2155]_  = \new_[7056]_  & \new_[7043]_ ;
  assign \new_[2156]_  = \new_[7030]_  & \new_[7017]_ ;
  assign \new_[2157]_  = \new_[7004]_  & \new_[6991]_ ;
  assign \new_[2158]_  = \new_[6978]_  & \new_[6965]_ ;
  assign \new_[2159]_  = \new_[6952]_  & \new_[6939]_ ;
  assign \new_[2160]_  = \new_[6926]_  & \new_[6913]_ ;
  assign \new_[2161]_  = \new_[6900]_  & \new_[6893]_ ;
  assign \new_[2162]_  = \new_[6886]_  & \new_[6879]_ ;
  assign \new_[2163]_  = \new_[6872]_  & \new_[6865]_ ;
  assign \new_[2164]_  = \new_[6860]_  & \new_[6853]_ ;
  assign \new_[2165]_  = \new_[6848]_  & \new_[6841]_ ;
  assign \new_[2166]_  = \new_[6836]_  & \new_[6829]_ ;
  assign \new_[2167]_  = \new_[6824]_  & \new_[6817]_ ;
  assign \new_[2168]_  = \new_[6812]_  & \new_[6805]_ ;
  assign \new_[2169]_  = \new_[6800]_  & \new_[6793]_ ;
  assign \new_[2170]_  = \new_[6788]_  & \new_[6781]_ ;
  assign \new_[2171]_  = \new_[6776]_  & \new_[6769]_ ;
  assign \new_[2172]_  = \new_[6764]_  & \new_[6757]_ ;
  assign \new_[2173]_  = \new_[6752]_  & \new_[6745]_ ;
  assign \new_[2174]_  = \new_[6740]_  & \new_[6733]_ ;
  assign \new_[2175]_  = \new_[6728]_  & \new_[6723]_ ;
  assign \new_[2176]_  = \new_[6718]_  & \new_[6713]_ ;
  assign \new_[2177]_  = \new_[6708]_  & \new_[6703]_ ;
  assign \new_[2178]_  = \new_[6698]_  & \new_[6693]_ ;
  assign \new_[2179]_  = \new_[6688]_  & \new_[6683]_ ;
  assign \new_[2180]_  = \new_[6678]_  & \new_[6673]_ ;
  assign \new_[2181]_  = \new_[6668]_  & \new_[6663]_ ;
  assign \new_[2182]_  = \new_[6658]_  & \new_[6653]_ ;
  assign \new_[2183]_  = \new_[6648]_  & \new_[6643]_ ;
  assign \new_[2184]_  = \new_[6638]_  & \new_[6633]_ ;
  assign \new_[2185]_  = \new_[6628]_  & \new_[6623]_ ;
  assign \new_[2186]_  = \new_[6618]_  & \new_[6613]_ ;
  assign \new_[2187]_  = \new_[6608]_  & \new_[6603]_ ;
  assign \new_[2188]_  = \new_[6598]_  & \new_[6593]_ ;
  assign \new_[2189]_  = \new_[6588]_  & \new_[6583]_ ;
  assign \new_[2190]_  = \new_[6578]_  & \new_[6573]_ ;
  assign \new_[2193]_  = \new_[2189]_  | \new_[2190]_ ;
  assign \new_[2196]_  = \new_[2187]_  | \new_[2188]_ ;
  assign \new_[2197]_  = \new_[2196]_  | \new_[2193]_ ;
  assign \new_[2200]_  = \new_[2185]_  | \new_[2186]_ ;
  assign \new_[2203]_  = \new_[2183]_  | \new_[2184]_ ;
  assign \new_[2204]_  = \new_[2203]_  | \new_[2200]_ ;
  assign \new_[2205]_  = \new_[2204]_  | \new_[2197]_ ;
  assign \new_[2208]_  = \new_[2181]_  | \new_[2182]_ ;
  assign \new_[2211]_  = \new_[2179]_  | \new_[2180]_ ;
  assign \new_[2212]_  = \new_[2211]_  | \new_[2208]_ ;
  assign \new_[2215]_  = \new_[2177]_  | \new_[2178]_ ;
  assign \new_[2219]_  = \new_[2174]_  | \new_[2175]_ ;
  assign \new_[2220]_  = \new_[2176]_  | \new_[2219]_ ;
  assign \new_[2221]_  = \new_[2220]_  | \new_[2215]_ ;
  assign \new_[2222]_  = \new_[2221]_  | \new_[2212]_ ;
  assign \new_[2223]_  = \new_[2222]_  | \new_[2205]_ ;
  assign \new_[2226]_  = \new_[2172]_  | \new_[2173]_ ;
  assign \new_[2229]_  = \new_[2170]_  | \new_[2171]_ ;
  assign \new_[2230]_  = \new_[2229]_  | \new_[2226]_ ;
  assign \new_[2233]_  = \new_[2168]_  | \new_[2169]_ ;
  assign \new_[2236]_  = \new_[2166]_  | \new_[2167]_ ;
  assign \new_[2237]_  = \new_[2236]_  | \new_[2233]_ ;
  assign \new_[2238]_  = \new_[2237]_  | \new_[2230]_ ;
  assign \new_[2241]_  = \new_[2164]_  | \new_[2165]_ ;
  assign \new_[2244]_  = \new_[2162]_  | \new_[2163]_ ;
  assign \new_[2245]_  = \new_[2244]_  | \new_[2241]_ ;
  assign \new_[2248]_  = \new_[2160]_  | \new_[2161]_ ;
  assign \new_[2252]_  = \new_[2157]_  | \new_[2158]_ ;
  assign \new_[2253]_  = \new_[2159]_  | \new_[2252]_ ;
  assign \new_[2254]_  = \new_[2253]_  | \new_[2248]_ ;
  assign \new_[2255]_  = \new_[2254]_  | \new_[2245]_ ;
  assign \new_[2256]_  = \new_[2255]_  | \new_[2238]_ ;
  assign \new_[2257]_  = \new_[2256]_  | \new_[2223]_ ;
  assign \new_[2260]_  = \new_[2155]_  | \new_[2156]_ ;
  assign \new_[2263]_  = \new_[2153]_  | \new_[2154]_ ;
  assign \new_[2264]_  = \new_[2263]_  | \new_[2260]_ ;
  assign \new_[2267]_  = \new_[2151]_  | \new_[2152]_ ;
  assign \new_[2270]_  = \new_[2149]_  | \new_[2150]_ ;
  assign \new_[2271]_  = \new_[2270]_  | \new_[2267]_ ;
  assign \new_[2272]_  = \new_[2271]_  | \new_[2264]_ ;
  assign \new_[2275]_  = \new_[2147]_  | \new_[2148]_ ;
  assign \new_[2278]_  = \new_[2145]_  | \new_[2146]_ ;
  assign \new_[2279]_  = \new_[2278]_  | \new_[2275]_ ;
  assign \new_[2282]_  = \new_[2143]_  | \new_[2144]_ ;
  assign \new_[2286]_  = \new_[2140]_  | \new_[2141]_ ;
  assign \new_[2287]_  = \new_[2142]_  | \new_[2286]_ ;
  assign \new_[2288]_  = \new_[2287]_  | \new_[2282]_ ;
  assign \new_[2289]_  = \new_[2288]_  | \new_[2279]_ ;
  assign \new_[2290]_  = \new_[2289]_  | \new_[2272]_ ;
  assign \new_[2293]_  = \new_[2138]_  | \new_[2139]_ ;
  assign \new_[2296]_  = \new_[2136]_  | \new_[2137]_ ;
  assign \new_[2297]_  = \new_[2296]_  | \new_[2293]_ ;
  assign \new_[2300]_  = \new_[2134]_  | \new_[2135]_ ;
  assign \new_[2303]_  = \new_[2132]_  | \new_[2133]_ ;
  assign \new_[2304]_  = \new_[2303]_  | \new_[2300]_ ;
  assign \new_[2305]_  = \new_[2304]_  | \new_[2297]_ ;
  assign \new_[2308]_  = \new_[2130]_  | \new_[2131]_ ;
  assign \new_[2311]_  = \new_[2128]_  | \new_[2129]_ ;
  assign \new_[2312]_  = \new_[2311]_  | \new_[2308]_ ;
  assign \new_[2315]_  = \new_[2126]_  | \new_[2127]_ ;
  assign \new_[2319]_  = \new_[2123]_  | \new_[2124]_ ;
  assign \new_[2320]_  = \new_[2125]_  | \new_[2319]_ ;
  assign \new_[2321]_  = \new_[2320]_  | \new_[2315]_ ;
  assign \new_[2322]_  = \new_[2321]_  | \new_[2312]_ ;
  assign \new_[2323]_  = \new_[2322]_  | \new_[2305]_ ;
  assign \new_[2324]_  = \new_[2323]_  | \new_[2290]_ ;
  assign \new_[2325]_  = \new_[2324]_  | \new_[2257]_ ;
  assign \new_[2328]_  = \new_[2121]_  | \new_[2122]_ ;
  assign \new_[2331]_  = \new_[2119]_  | \new_[2120]_ ;
  assign \new_[2332]_  = \new_[2331]_  | \new_[2328]_ ;
  assign \new_[2335]_  = \new_[2117]_  | \new_[2118]_ ;
  assign \new_[2338]_  = \new_[2115]_  | \new_[2116]_ ;
  assign \new_[2339]_  = \new_[2338]_  | \new_[2335]_ ;
  assign \new_[2340]_  = \new_[2339]_  | \new_[2332]_ ;
  assign \new_[2343]_  = \new_[2113]_  | \new_[2114]_ ;
  assign \new_[2346]_  = \new_[2111]_  | \new_[2112]_ ;
  assign \new_[2347]_  = \new_[2346]_  | \new_[2343]_ ;
  assign \new_[2350]_  = \new_[2109]_  | \new_[2110]_ ;
  assign \new_[2354]_  = \new_[2106]_  | \new_[2107]_ ;
  assign \new_[2355]_  = \new_[2108]_  | \new_[2354]_ ;
  assign \new_[2356]_  = \new_[2355]_  | \new_[2350]_ ;
  assign \new_[2357]_  = \new_[2356]_  | \new_[2347]_ ;
  assign \new_[2358]_  = \new_[2357]_  | \new_[2340]_ ;
  assign \new_[2361]_  = \new_[2104]_  | \new_[2105]_ ;
  assign \new_[2364]_  = \new_[2102]_  | \new_[2103]_ ;
  assign \new_[2365]_  = \new_[2364]_  | \new_[2361]_ ;
  assign \new_[2368]_  = \new_[2100]_  | \new_[2101]_ ;
  assign \new_[2371]_  = \new_[2098]_  | \new_[2099]_ ;
  assign \new_[2372]_  = \new_[2371]_  | \new_[2368]_ ;
  assign \new_[2373]_  = \new_[2372]_  | \new_[2365]_ ;
  assign \new_[2376]_  = \new_[2096]_  | \new_[2097]_ ;
  assign \new_[2379]_  = \new_[2094]_  | \new_[2095]_ ;
  assign \new_[2380]_  = \new_[2379]_  | \new_[2376]_ ;
  assign \new_[2383]_  = \new_[2092]_  | \new_[2093]_ ;
  assign \new_[2387]_  = \new_[2089]_  | \new_[2090]_ ;
  assign \new_[2388]_  = \new_[2091]_  | \new_[2387]_ ;
  assign \new_[2389]_  = \new_[2388]_  | \new_[2383]_ ;
  assign \new_[2390]_  = \new_[2389]_  | \new_[2380]_ ;
  assign \new_[2391]_  = \new_[2390]_  | \new_[2373]_ ;
  assign \new_[2392]_  = \new_[2391]_  | \new_[2358]_ ;
  assign \new_[2395]_  = \new_[2087]_  | \new_[2088]_ ;
  assign \new_[2398]_  = \new_[2085]_  | \new_[2086]_ ;
  assign \new_[2399]_  = \new_[2398]_  | \new_[2395]_ ;
  assign \new_[2402]_  = \new_[2083]_  | \new_[2084]_ ;
  assign \new_[2405]_  = \new_[2081]_  | \new_[2082]_ ;
  assign \new_[2406]_  = \new_[2405]_  | \new_[2402]_ ;
  assign \new_[2407]_  = \new_[2406]_  | \new_[2399]_ ;
  assign \new_[2410]_  = \new_[2079]_  | \new_[2080]_ ;
  assign \new_[2413]_  = \new_[2077]_  | \new_[2078]_ ;
  assign \new_[2414]_  = \new_[2413]_  | \new_[2410]_ ;
  assign \new_[2417]_  = \new_[2075]_  | \new_[2076]_ ;
  assign \new_[2421]_  = \new_[2072]_  | \new_[2073]_ ;
  assign \new_[2422]_  = \new_[2074]_  | \new_[2421]_ ;
  assign \new_[2423]_  = \new_[2422]_  | \new_[2417]_ ;
  assign \new_[2424]_  = \new_[2423]_  | \new_[2414]_ ;
  assign \new_[2425]_  = \new_[2424]_  | \new_[2407]_ ;
  assign \new_[2428]_  = \new_[2070]_  | \new_[2071]_ ;
  assign \new_[2431]_  = \new_[2068]_  | \new_[2069]_ ;
  assign \new_[2432]_  = \new_[2431]_  | \new_[2428]_ ;
  assign \new_[2435]_  = \new_[2066]_  | \new_[2067]_ ;
  assign \new_[2438]_  = \new_[2064]_  | \new_[2065]_ ;
  assign \new_[2439]_  = \new_[2438]_  | \new_[2435]_ ;
  assign \new_[2440]_  = \new_[2439]_  | \new_[2432]_ ;
  assign \new_[2443]_  = \new_[2062]_  | \new_[2063]_ ;
  assign \new_[2446]_  = \new_[2060]_  | \new_[2061]_ ;
  assign \new_[2447]_  = \new_[2446]_  | \new_[2443]_ ;
  assign \new_[2450]_  = \new_[2058]_  | \new_[2059]_ ;
  assign \new_[2454]_  = \new_[2055]_  | \new_[2056]_ ;
  assign \new_[2455]_  = \new_[2057]_  | \new_[2454]_ ;
  assign \new_[2456]_  = \new_[2455]_  | \new_[2450]_ ;
  assign \new_[2457]_  = \new_[2456]_  | \new_[2447]_ ;
  assign \new_[2458]_  = \new_[2457]_  | \new_[2440]_ ;
  assign \new_[2459]_  = \new_[2458]_  | \new_[2425]_ ;
  assign \new_[2460]_  = \new_[2459]_  | \new_[2392]_ ;
  assign \new_[2461]_  = \new_[2460]_  | \new_[2325]_ ;
  assign \new_[2464]_  = \new_[2053]_  | \new_[2054]_ ;
  assign \new_[2467]_  = \new_[2051]_  | \new_[2052]_ ;
  assign \new_[2468]_  = \new_[2467]_  | \new_[2464]_ ;
  assign \new_[2471]_  = \new_[2049]_  | \new_[2050]_ ;
  assign \new_[2474]_  = \new_[2047]_  | \new_[2048]_ ;
  assign \new_[2475]_  = \new_[2474]_  | \new_[2471]_ ;
  assign \new_[2476]_  = \new_[2475]_  | \new_[2468]_ ;
  assign \new_[2479]_  = \new_[2045]_  | \new_[2046]_ ;
  assign \new_[2482]_  = \new_[2043]_  | \new_[2044]_ ;
  assign \new_[2483]_  = \new_[2482]_  | \new_[2479]_ ;
  assign \new_[2486]_  = \new_[2041]_  | \new_[2042]_ ;
  assign \new_[2490]_  = \new_[2038]_  | \new_[2039]_ ;
  assign \new_[2491]_  = \new_[2040]_  | \new_[2490]_ ;
  assign \new_[2492]_  = \new_[2491]_  | \new_[2486]_ ;
  assign \new_[2493]_  = \new_[2492]_  | \new_[2483]_ ;
  assign \new_[2494]_  = \new_[2493]_  | \new_[2476]_ ;
  assign \new_[2497]_  = \new_[2036]_  | \new_[2037]_ ;
  assign \new_[2500]_  = \new_[2034]_  | \new_[2035]_ ;
  assign \new_[2501]_  = \new_[2500]_  | \new_[2497]_ ;
  assign \new_[2504]_  = \new_[2032]_  | \new_[2033]_ ;
  assign \new_[2507]_  = \new_[2030]_  | \new_[2031]_ ;
  assign \new_[2508]_  = \new_[2507]_  | \new_[2504]_ ;
  assign \new_[2509]_  = \new_[2508]_  | \new_[2501]_ ;
  assign \new_[2512]_  = \new_[2028]_  | \new_[2029]_ ;
  assign \new_[2515]_  = \new_[2026]_  | \new_[2027]_ ;
  assign \new_[2516]_  = \new_[2515]_  | \new_[2512]_ ;
  assign \new_[2519]_  = \new_[2024]_  | \new_[2025]_ ;
  assign \new_[2523]_  = \new_[2021]_  | \new_[2022]_ ;
  assign \new_[2524]_  = \new_[2023]_  | \new_[2523]_ ;
  assign \new_[2525]_  = \new_[2524]_  | \new_[2519]_ ;
  assign \new_[2526]_  = \new_[2525]_  | \new_[2516]_ ;
  assign \new_[2527]_  = \new_[2526]_  | \new_[2509]_ ;
  assign \new_[2528]_  = \new_[2527]_  | \new_[2494]_ ;
  assign \new_[2531]_  = \new_[2019]_  | \new_[2020]_ ;
  assign \new_[2534]_  = \new_[2017]_  | \new_[2018]_ ;
  assign \new_[2535]_  = \new_[2534]_  | \new_[2531]_ ;
  assign \new_[2538]_  = \new_[2015]_  | \new_[2016]_ ;
  assign \new_[2541]_  = \new_[2013]_  | \new_[2014]_ ;
  assign \new_[2542]_  = \new_[2541]_  | \new_[2538]_ ;
  assign \new_[2543]_  = \new_[2542]_  | \new_[2535]_ ;
  assign \new_[2546]_  = \new_[2011]_  | \new_[2012]_ ;
  assign \new_[2549]_  = \new_[2009]_  | \new_[2010]_ ;
  assign \new_[2550]_  = \new_[2549]_  | \new_[2546]_ ;
  assign \new_[2553]_  = \new_[2007]_  | \new_[2008]_ ;
  assign \new_[2557]_  = \new_[2004]_  | \new_[2005]_ ;
  assign \new_[2558]_  = \new_[2006]_  | \new_[2557]_ ;
  assign \new_[2559]_  = \new_[2558]_  | \new_[2553]_ ;
  assign \new_[2560]_  = \new_[2559]_  | \new_[2550]_ ;
  assign \new_[2561]_  = \new_[2560]_  | \new_[2543]_ ;
  assign \new_[2564]_  = \new_[2002]_  | \new_[2003]_ ;
  assign \new_[2567]_  = \new_[2000]_  | \new_[2001]_ ;
  assign \new_[2568]_  = \new_[2567]_  | \new_[2564]_ ;
  assign \new_[2571]_  = \new_[1998]_  | \new_[1999]_ ;
  assign \new_[2574]_  = \new_[1996]_  | \new_[1997]_ ;
  assign \new_[2575]_  = \new_[2574]_  | \new_[2571]_ ;
  assign \new_[2576]_  = \new_[2575]_  | \new_[2568]_ ;
  assign \new_[2579]_  = \new_[1994]_  | \new_[1995]_ ;
  assign \new_[2582]_  = \new_[1992]_  | \new_[1993]_ ;
  assign \new_[2583]_  = \new_[2582]_  | \new_[2579]_ ;
  assign \new_[2586]_  = \new_[1990]_  | \new_[1991]_ ;
  assign \new_[2590]_  = \new_[1987]_  | \new_[1988]_ ;
  assign \new_[2591]_  = \new_[1989]_  | \new_[2590]_ ;
  assign \new_[2592]_  = \new_[2591]_  | \new_[2586]_ ;
  assign \new_[2593]_  = \new_[2592]_  | \new_[2583]_ ;
  assign \new_[2594]_  = \new_[2593]_  | \new_[2576]_ ;
  assign \new_[2595]_  = \new_[2594]_  | \new_[2561]_ ;
  assign \new_[2596]_  = \new_[2595]_  | \new_[2528]_ ;
  assign \new_[2599]_  = \new_[1985]_  | \new_[1986]_ ;
  assign \new_[2602]_  = \new_[1983]_  | \new_[1984]_ ;
  assign \new_[2603]_  = \new_[2602]_  | \new_[2599]_ ;
  assign \new_[2606]_  = \new_[1981]_  | \new_[1982]_ ;
  assign \new_[2609]_  = \new_[1979]_  | \new_[1980]_ ;
  assign \new_[2610]_  = \new_[2609]_  | \new_[2606]_ ;
  assign \new_[2611]_  = \new_[2610]_  | \new_[2603]_ ;
  assign \new_[2614]_  = \new_[1977]_  | \new_[1978]_ ;
  assign \new_[2617]_  = \new_[1975]_  | \new_[1976]_ ;
  assign \new_[2618]_  = \new_[2617]_  | \new_[2614]_ ;
  assign \new_[2621]_  = \new_[1973]_  | \new_[1974]_ ;
  assign \new_[2625]_  = \new_[1970]_  | \new_[1971]_ ;
  assign \new_[2626]_  = \new_[1972]_  | \new_[2625]_ ;
  assign \new_[2627]_  = \new_[2626]_  | \new_[2621]_ ;
  assign \new_[2628]_  = \new_[2627]_  | \new_[2618]_ ;
  assign \new_[2629]_  = \new_[2628]_  | \new_[2611]_ ;
  assign \new_[2632]_  = \new_[1968]_  | \new_[1969]_ ;
  assign \new_[2635]_  = \new_[1966]_  | \new_[1967]_ ;
  assign \new_[2636]_  = \new_[2635]_  | \new_[2632]_ ;
  assign \new_[2639]_  = \new_[1964]_  | \new_[1965]_ ;
  assign \new_[2642]_  = \new_[1962]_  | \new_[1963]_ ;
  assign \new_[2643]_  = \new_[2642]_  | \new_[2639]_ ;
  assign \new_[2644]_  = \new_[2643]_  | \new_[2636]_ ;
  assign \new_[2647]_  = \new_[1960]_  | \new_[1961]_ ;
  assign \new_[2650]_  = \new_[1958]_  | \new_[1959]_ ;
  assign \new_[2651]_  = \new_[2650]_  | \new_[2647]_ ;
  assign \new_[2654]_  = \new_[1956]_  | \new_[1957]_ ;
  assign \new_[2658]_  = \new_[1953]_  | \new_[1954]_ ;
  assign \new_[2659]_  = \new_[1955]_  | \new_[2658]_ ;
  assign \new_[2660]_  = \new_[2659]_  | \new_[2654]_ ;
  assign \new_[2661]_  = \new_[2660]_  | \new_[2651]_ ;
  assign \new_[2662]_  = \new_[2661]_  | \new_[2644]_ ;
  assign \new_[2663]_  = \new_[2662]_  | \new_[2629]_ ;
  assign \new_[2666]_  = \new_[1951]_  | \new_[1952]_ ;
  assign \new_[2669]_  = \new_[1949]_  | \new_[1950]_ ;
  assign \new_[2670]_  = \new_[2669]_  | \new_[2666]_ ;
  assign \new_[2673]_  = \new_[1947]_  | \new_[1948]_ ;
  assign \new_[2676]_  = \new_[1945]_  | \new_[1946]_ ;
  assign \new_[2677]_  = \new_[2676]_  | \new_[2673]_ ;
  assign \new_[2678]_  = \new_[2677]_  | \new_[2670]_ ;
  assign \new_[2681]_  = \new_[1943]_  | \new_[1944]_ ;
  assign \new_[2684]_  = \new_[1941]_  | \new_[1942]_ ;
  assign \new_[2685]_  = \new_[2684]_  | \new_[2681]_ ;
  assign \new_[2688]_  = \new_[1939]_  | \new_[1940]_ ;
  assign \new_[2692]_  = \new_[1936]_  | \new_[1937]_ ;
  assign \new_[2693]_  = \new_[1938]_  | \new_[2692]_ ;
  assign \new_[2694]_  = \new_[2693]_  | \new_[2688]_ ;
  assign \new_[2695]_  = \new_[2694]_  | \new_[2685]_ ;
  assign \new_[2696]_  = \new_[2695]_  | \new_[2678]_ ;
  assign \new_[2699]_  = \new_[1934]_  | \new_[1935]_ ;
  assign \new_[2702]_  = \new_[1932]_  | \new_[1933]_ ;
  assign \new_[2703]_  = \new_[2702]_  | \new_[2699]_ ;
  assign \new_[2706]_  = \new_[1930]_  | \new_[1931]_ ;
  assign \new_[2710]_  = \new_[1927]_  | \new_[1928]_ ;
  assign \new_[2711]_  = \new_[1929]_  | \new_[2710]_ ;
  assign \new_[2712]_  = \new_[2711]_  | \new_[2706]_ ;
  assign \new_[2713]_  = \new_[2712]_  | \new_[2703]_ ;
  assign \new_[2716]_  = \new_[1925]_  | \new_[1926]_ ;
  assign \new_[2719]_  = \new_[1923]_  | \new_[1924]_ ;
  assign \new_[2720]_  = \new_[2719]_  | \new_[2716]_ ;
  assign \new_[2723]_  = \new_[1921]_  | \new_[1922]_ ;
  assign \new_[2727]_  = \new_[1918]_  | \new_[1919]_ ;
  assign \new_[2728]_  = \new_[1920]_  | \new_[2727]_ ;
  assign \new_[2729]_  = \new_[2728]_  | \new_[2723]_ ;
  assign \new_[2730]_  = \new_[2729]_  | \new_[2720]_ ;
  assign \new_[2731]_  = \new_[2730]_  | \new_[2713]_ ;
  assign \new_[2732]_  = \new_[2731]_  | \new_[2696]_ ;
  assign \new_[2733]_  = \new_[2732]_  | \new_[2663]_ ;
  assign \new_[2734]_  = \new_[2733]_  | \new_[2596]_ ;
  assign \new_[2735]_  = \new_[2734]_  | \new_[2461]_ ;
  assign \new_[2738]_  = \new_[1916]_  | \new_[1917]_ ;
  assign \new_[2741]_  = \new_[1914]_  | \new_[1915]_ ;
  assign \new_[2742]_  = \new_[2741]_  | \new_[2738]_ ;
  assign \new_[2745]_  = \new_[1912]_  | \new_[1913]_ ;
  assign \new_[2748]_  = \new_[1910]_  | \new_[1911]_ ;
  assign \new_[2749]_  = \new_[2748]_  | \new_[2745]_ ;
  assign \new_[2750]_  = \new_[2749]_  | \new_[2742]_ ;
  assign \new_[2753]_  = \new_[1908]_  | \new_[1909]_ ;
  assign \new_[2756]_  = \new_[1906]_  | \new_[1907]_ ;
  assign \new_[2757]_  = \new_[2756]_  | \new_[2753]_ ;
  assign \new_[2760]_  = \new_[1904]_  | \new_[1905]_ ;
  assign \new_[2764]_  = \new_[1901]_  | \new_[1902]_ ;
  assign \new_[2765]_  = \new_[1903]_  | \new_[2764]_ ;
  assign \new_[2766]_  = \new_[2765]_  | \new_[2760]_ ;
  assign \new_[2767]_  = \new_[2766]_  | \new_[2757]_ ;
  assign \new_[2768]_  = \new_[2767]_  | \new_[2750]_ ;
  assign \new_[2771]_  = \new_[1899]_  | \new_[1900]_ ;
  assign \new_[2774]_  = \new_[1897]_  | \new_[1898]_ ;
  assign \new_[2775]_  = \new_[2774]_  | \new_[2771]_ ;
  assign \new_[2778]_  = \new_[1895]_  | \new_[1896]_ ;
  assign \new_[2781]_  = \new_[1893]_  | \new_[1894]_ ;
  assign \new_[2782]_  = \new_[2781]_  | \new_[2778]_ ;
  assign \new_[2783]_  = \new_[2782]_  | \new_[2775]_ ;
  assign \new_[2786]_  = \new_[1891]_  | \new_[1892]_ ;
  assign \new_[2789]_  = \new_[1889]_  | \new_[1890]_ ;
  assign \new_[2790]_  = \new_[2789]_  | \new_[2786]_ ;
  assign \new_[2793]_  = \new_[1887]_  | \new_[1888]_ ;
  assign \new_[2797]_  = \new_[1884]_  | \new_[1885]_ ;
  assign \new_[2798]_  = \new_[1886]_  | \new_[2797]_ ;
  assign \new_[2799]_  = \new_[2798]_  | \new_[2793]_ ;
  assign \new_[2800]_  = \new_[2799]_  | \new_[2790]_ ;
  assign \new_[2801]_  = \new_[2800]_  | \new_[2783]_ ;
  assign \new_[2802]_  = \new_[2801]_  | \new_[2768]_ ;
  assign \new_[2805]_  = \new_[1882]_  | \new_[1883]_ ;
  assign \new_[2808]_  = \new_[1880]_  | \new_[1881]_ ;
  assign \new_[2809]_  = \new_[2808]_  | \new_[2805]_ ;
  assign \new_[2812]_  = \new_[1878]_  | \new_[1879]_ ;
  assign \new_[2815]_  = \new_[1876]_  | \new_[1877]_ ;
  assign \new_[2816]_  = \new_[2815]_  | \new_[2812]_ ;
  assign \new_[2817]_  = \new_[2816]_  | \new_[2809]_ ;
  assign \new_[2820]_  = \new_[1874]_  | \new_[1875]_ ;
  assign \new_[2823]_  = \new_[1872]_  | \new_[1873]_ ;
  assign \new_[2824]_  = \new_[2823]_  | \new_[2820]_ ;
  assign \new_[2827]_  = \new_[1870]_  | \new_[1871]_ ;
  assign \new_[2831]_  = \new_[1867]_  | \new_[1868]_ ;
  assign \new_[2832]_  = \new_[1869]_  | \new_[2831]_ ;
  assign \new_[2833]_  = \new_[2832]_  | \new_[2827]_ ;
  assign \new_[2834]_  = \new_[2833]_  | \new_[2824]_ ;
  assign \new_[2835]_  = \new_[2834]_  | \new_[2817]_ ;
  assign \new_[2838]_  = \new_[1865]_  | \new_[1866]_ ;
  assign \new_[2841]_  = \new_[1863]_  | \new_[1864]_ ;
  assign \new_[2842]_  = \new_[2841]_  | \new_[2838]_ ;
  assign \new_[2845]_  = \new_[1861]_  | \new_[1862]_ ;
  assign \new_[2848]_  = \new_[1859]_  | \new_[1860]_ ;
  assign \new_[2849]_  = \new_[2848]_  | \new_[2845]_ ;
  assign \new_[2850]_  = \new_[2849]_  | \new_[2842]_ ;
  assign \new_[2853]_  = \new_[1857]_  | \new_[1858]_ ;
  assign \new_[2856]_  = \new_[1855]_  | \new_[1856]_ ;
  assign \new_[2857]_  = \new_[2856]_  | \new_[2853]_ ;
  assign \new_[2860]_  = \new_[1853]_  | \new_[1854]_ ;
  assign \new_[2864]_  = \new_[1850]_  | \new_[1851]_ ;
  assign \new_[2865]_  = \new_[1852]_  | \new_[2864]_ ;
  assign \new_[2866]_  = \new_[2865]_  | \new_[2860]_ ;
  assign \new_[2867]_  = \new_[2866]_  | \new_[2857]_ ;
  assign \new_[2868]_  = \new_[2867]_  | \new_[2850]_ ;
  assign \new_[2869]_  = \new_[2868]_  | \new_[2835]_ ;
  assign \new_[2870]_  = \new_[2869]_  | \new_[2802]_ ;
  assign \new_[2873]_  = \new_[1848]_  | \new_[1849]_ ;
  assign \new_[2876]_  = \new_[1846]_  | \new_[1847]_ ;
  assign \new_[2877]_  = \new_[2876]_  | \new_[2873]_ ;
  assign \new_[2880]_  = \new_[1844]_  | \new_[1845]_ ;
  assign \new_[2883]_  = \new_[1842]_  | \new_[1843]_ ;
  assign \new_[2884]_  = \new_[2883]_  | \new_[2880]_ ;
  assign \new_[2885]_  = \new_[2884]_  | \new_[2877]_ ;
  assign \new_[2888]_  = \new_[1840]_  | \new_[1841]_ ;
  assign \new_[2891]_  = \new_[1838]_  | \new_[1839]_ ;
  assign \new_[2892]_  = \new_[2891]_  | \new_[2888]_ ;
  assign \new_[2895]_  = \new_[1836]_  | \new_[1837]_ ;
  assign \new_[2899]_  = \new_[1833]_  | \new_[1834]_ ;
  assign \new_[2900]_  = \new_[1835]_  | \new_[2899]_ ;
  assign \new_[2901]_  = \new_[2900]_  | \new_[2895]_ ;
  assign \new_[2902]_  = \new_[2901]_  | \new_[2892]_ ;
  assign \new_[2903]_  = \new_[2902]_  | \new_[2885]_ ;
  assign \new_[2906]_  = \new_[1831]_  | \new_[1832]_ ;
  assign \new_[2909]_  = \new_[1829]_  | \new_[1830]_ ;
  assign \new_[2910]_  = \new_[2909]_  | \new_[2906]_ ;
  assign \new_[2913]_  = \new_[1827]_  | \new_[1828]_ ;
  assign \new_[2916]_  = \new_[1825]_  | \new_[1826]_ ;
  assign \new_[2917]_  = \new_[2916]_  | \new_[2913]_ ;
  assign \new_[2918]_  = \new_[2917]_  | \new_[2910]_ ;
  assign \new_[2921]_  = \new_[1823]_  | \new_[1824]_ ;
  assign \new_[2924]_  = \new_[1821]_  | \new_[1822]_ ;
  assign \new_[2925]_  = \new_[2924]_  | \new_[2921]_ ;
  assign \new_[2928]_  = \new_[1819]_  | \new_[1820]_ ;
  assign \new_[2932]_  = \new_[1816]_  | \new_[1817]_ ;
  assign \new_[2933]_  = \new_[1818]_  | \new_[2932]_ ;
  assign \new_[2934]_  = \new_[2933]_  | \new_[2928]_ ;
  assign \new_[2935]_  = \new_[2934]_  | \new_[2925]_ ;
  assign \new_[2936]_  = \new_[2935]_  | \new_[2918]_ ;
  assign \new_[2937]_  = \new_[2936]_  | \new_[2903]_ ;
  assign \new_[2940]_  = \new_[1814]_  | \new_[1815]_ ;
  assign \new_[2943]_  = \new_[1812]_  | \new_[1813]_ ;
  assign \new_[2944]_  = \new_[2943]_  | \new_[2940]_ ;
  assign \new_[2947]_  = \new_[1810]_  | \new_[1811]_ ;
  assign \new_[2950]_  = \new_[1808]_  | \new_[1809]_ ;
  assign \new_[2951]_  = \new_[2950]_  | \new_[2947]_ ;
  assign \new_[2952]_  = \new_[2951]_  | \new_[2944]_ ;
  assign \new_[2955]_  = \new_[1806]_  | \new_[1807]_ ;
  assign \new_[2958]_  = \new_[1804]_  | \new_[1805]_ ;
  assign \new_[2959]_  = \new_[2958]_  | \new_[2955]_ ;
  assign \new_[2962]_  = \new_[1802]_  | \new_[1803]_ ;
  assign \new_[2966]_  = \new_[1799]_  | \new_[1800]_ ;
  assign \new_[2967]_  = \new_[1801]_  | \new_[2966]_ ;
  assign \new_[2968]_  = \new_[2967]_  | \new_[2962]_ ;
  assign \new_[2969]_  = \new_[2968]_  | \new_[2959]_ ;
  assign \new_[2970]_  = \new_[2969]_  | \new_[2952]_ ;
  assign \new_[2973]_  = \new_[1797]_  | \new_[1798]_ ;
  assign \new_[2976]_  = \new_[1795]_  | \new_[1796]_ ;
  assign \new_[2977]_  = \new_[2976]_  | \new_[2973]_ ;
  assign \new_[2980]_  = \new_[1793]_  | \new_[1794]_ ;
  assign \new_[2984]_  = \new_[1790]_  | \new_[1791]_ ;
  assign \new_[2985]_  = \new_[1792]_  | \new_[2984]_ ;
  assign \new_[2986]_  = \new_[2985]_  | \new_[2980]_ ;
  assign \new_[2987]_  = \new_[2986]_  | \new_[2977]_ ;
  assign \new_[2990]_  = \new_[1788]_  | \new_[1789]_ ;
  assign \new_[2993]_  = \new_[1786]_  | \new_[1787]_ ;
  assign \new_[2994]_  = \new_[2993]_  | \new_[2990]_ ;
  assign \new_[2997]_  = \new_[1784]_  | \new_[1785]_ ;
  assign \new_[3001]_  = \new_[1781]_  | \new_[1782]_ ;
  assign \new_[3002]_  = \new_[1783]_  | \new_[3001]_ ;
  assign \new_[3003]_  = \new_[3002]_  | \new_[2997]_ ;
  assign \new_[3004]_  = \new_[3003]_  | \new_[2994]_ ;
  assign \new_[3005]_  = \new_[3004]_  | \new_[2987]_ ;
  assign \new_[3006]_  = \new_[3005]_  | \new_[2970]_ ;
  assign \new_[3007]_  = \new_[3006]_  | \new_[2937]_ ;
  assign \new_[3008]_  = \new_[3007]_  | \new_[2870]_ ;
  assign \new_[3011]_  = \new_[1779]_  | \new_[1780]_ ;
  assign \new_[3014]_  = \new_[1777]_  | \new_[1778]_ ;
  assign \new_[3015]_  = \new_[3014]_  | \new_[3011]_ ;
  assign \new_[3018]_  = \new_[1775]_  | \new_[1776]_ ;
  assign \new_[3021]_  = \new_[1773]_  | \new_[1774]_ ;
  assign \new_[3022]_  = \new_[3021]_  | \new_[3018]_ ;
  assign \new_[3023]_  = \new_[3022]_  | \new_[3015]_ ;
  assign \new_[3026]_  = \new_[1771]_  | \new_[1772]_ ;
  assign \new_[3029]_  = \new_[1769]_  | \new_[1770]_ ;
  assign \new_[3030]_  = \new_[3029]_  | \new_[3026]_ ;
  assign \new_[3033]_  = \new_[1767]_  | \new_[1768]_ ;
  assign \new_[3037]_  = \new_[1764]_  | \new_[1765]_ ;
  assign \new_[3038]_  = \new_[1766]_  | \new_[3037]_ ;
  assign \new_[3039]_  = \new_[3038]_  | \new_[3033]_ ;
  assign \new_[3040]_  = \new_[3039]_  | \new_[3030]_ ;
  assign \new_[3041]_  = \new_[3040]_  | \new_[3023]_ ;
  assign \new_[3044]_  = \new_[1762]_  | \new_[1763]_ ;
  assign \new_[3047]_  = \new_[1760]_  | \new_[1761]_ ;
  assign \new_[3048]_  = \new_[3047]_  | \new_[3044]_ ;
  assign \new_[3051]_  = \new_[1758]_  | \new_[1759]_ ;
  assign \new_[3054]_  = \new_[1756]_  | \new_[1757]_ ;
  assign \new_[3055]_  = \new_[3054]_  | \new_[3051]_ ;
  assign \new_[3056]_  = \new_[3055]_  | \new_[3048]_ ;
  assign \new_[3059]_  = \new_[1754]_  | \new_[1755]_ ;
  assign \new_[3062]_  = \new_[1752]_  | \new_[1753]_ ;
  assign \new_[3063]_  = \new_[3062]_  | \new_[3059]_ ;
  assign \new_[3066]_  = \new_[1750]_  | \new_[1751]_ ;
  assign \new_[3070]_  = \new_[1747]_  | \new_[1748]_ ;
  assign \new_[3071]_  = \new_[1749]_  | \new_[3070]_ ;
  assign \new_[3072]_  = \new_[3071]_  | \new_[3066]_ ;
  assign \new_[3073]_  = \new_[3072]_  | \new_[3063]_ ;
  assign \new_[3074]_  = \new_[3073]_  | \new_[3056]_ ;
  assign \new_[3075]_  = \new_[3074]_  | \new_[3041]_ ;
  assign \new_[3078]_  = \new_[1745]_  | \new_[1746]_ ;
  assign \new_[3081]_  = \new_[1743]_  | \new_[1744]_ ;
  assign \new_[3082]_  = \new_[3081]_  | \new_[3078]_ ;
  assign \new_[3085]_  = \new_[1741]_  | \new_[1742]_ ;
  assign \new_[3088]_  = \new_[1739]_  | \new_[1740]_ ;
  assign \new_[3089]_  = \new_[3088]_  | \new_[3085]_ ;
  assign \new_[3090]_  = \new_[3089]_  | \new_[3082]_ ;
  assign \new_[3093]_  = \new_[1737]_  | \new_[1738]_ ;
  assign \new_[3096]_  = \new_[1735]_  | \new_[1736]_ ;
  assign \new_[3097]_  = \new_[3096]_  | \new_[3093]_ ;
  assign \new_[3100]_  = \new_[1733]_  | \new_[1734]_ ;
  assign \new_[3104]_  = \new_[1730]_  | \new_[1731]_ ;
  assign \new_[3105]_  = \new_[1732]_  | \new_[3104]_ ;
  assign \new_[3106]_  = \new_[3105]_  | \new_[3100]_ ;
  assign \new_[3107]_  = \new_[3106]_  | \new_[3097]_ ;
  assign \new_[3108]_  = \new_[3107]_  | \new_[3090]_ ;
  assign \new_[3111]_  = \new_[1728]_  | \new_[1729]_ ;
  assign \new_[3114]_  = \new_[1726]_  | \new_[1727]_ ;
  assign \new_[3115]_  = \new_[3114]_  | \new_[3111]_ ;
  assign \new_[3118]_  = \new_[1724]_  | \new_[1725]_ ;
  assign \new_[3121]_  = \new_[1722]_  | \new_[1723]_ ;
  assign \new_[3122]_  = \new_[3121]_  | \new_[3118]_ ;
  assign \new_[3123]_  = \new_[3122]_  | \new_[3115]_ ;
  assign \new_[3126]_  = \new_[1720]_  | \new_[1721]_ ;
  assign \new_[3129]_  = \new_[1718]_  | \new_[1719]_ ;
  assign \new_[3130]_  = \new_[3129]_  | \new_[3126]_ ;
  assign \new_[3133]_  = \new_[1716]_  | \new_[1717]_ ;
  assign \new_[3137]_  = \new_[1713]_  | \new_[1714]_ ;
  assign \new_[3138]_  = \new_[1715]_  | \new_[3137]_ ;
  assign \new_[3139]_  = \new_[3138]_  | \new_[3133]_ ;
  assign \new_[3140]_  = \new_[3139]_  | \new_[3130]_ ;
  assign \new_[3141]_  = \new_[3140]_  | \new_[3123]_ ;
  assign \new_[3142]_  = \new_[3141]_  | \new_[3108]_ ;
  assign \new_[3143]_  = \new_[3142]_  | \new_[3075]_ ;
  assign \new_[3146]_  = \new_[1711]_  | \new_[1712]_ ;
  assign \new_[3149]_  = \new_[1709]_  | \new_[1710]_ ;
  assign \new_[3150]_  = \new_[3149]_  | \new_[3146]_ ;
  assign \new_[3153]_  = \new_[1707]_  | \new_[1708]_ ;
  assign \new_[3156]_  = \new_[1705]_  | \new_[1706]_ ;
  assign \new_[3157]_  = \new_[3156]_  | \new_[3153]_ ;
  assign \new_[3158]_  = \new_[3157]_  | \new_[3150]_ ;
  assign \new_[3161]_  = \new_[1703]_  | \new_[1704]_ ;
  assign \new_[3164]_  = \new_[1701]_  | \new_[1702]_ ;
  assign \new_[3165]_  = \new_[3164]_  | \new_[3161]_ ;
  assign \new_[3168]_  = \new_[1699]_  | \new_[1700]_ ;
  assign \new_[3172]_  = \new_[1696]_  | \new_[1697]_ ;
  assign \new_[3173]_  = \new_[1698]_  | \new_[3172]_ ;
  assign \new_[3174]_  = \new_[3173]_  | \new_[3168]_ ;
  assign \new_[3175]_  = \new_[3174]_  | \new_[3165]_ ;
  assign \new_[3176]_  = \new_[3175]_  | \new_[3158]_ ;
  assign \new_[3179]_  = \new_[1694]_  | \new_[1695]_ ;
  assign \new_[3182]_  = \new_[1692]_  | \new_[1693]_ ;
  assign \new_[3183]_  = \new_[3182]_  | \new_[3179]_ ;
  assign \new_[3186]_  = \new_[1690]_  | \new_[1691]_ ;
  assign \new_[3189]_  = \new_[1688]_  | \new_[1689]_ ;
  assign \new_[3190]_  = \new_[3189]_  | \new_[3186]_ ;
  assign \new_[3191]_  = \new_[3190]_  | \new_[3183]_ ;
  assign \new_[3194]_  = \new_[1686]_  | \new_[1687]_ ;
  assign \new_[3197]_  = \new_[1684]_  | \new_[1685]_ ;
  assign \new_[3198]_  = \new_[3197]_  | \new_[3194]_ ;
  assign \new_[3201]_  = \new_[1682]_  | \new_[1683]_ ;
  assign \new_[3205]_  = \new_[1679]_  | \new_[1680]_ ;
  assign \new_[3206]_  = \new_[1681]_  | \new_[3205]_ ;
  assign \new_[3207]_  = \new_[3206]_  | \new_[3201]_ ;
  assign \new_[3208]_  = \new_[3207]_  | \new_[3198]_ ;
  assign \new_[3209]_  = \new_[3208]_  | \new_[3191]_ ;
  assign \new_[3210]_  = \new_[3209]_  | \new_[3176]_ ;
  assign \new_[3213]_  = \new_[1677]_  | \new_[1678]_ ;
  assign \new_[3216]_  = \new_[1675]_  | \new_[1676]_ ;
  assign \new_[3217]_  = \new_[3216]_  | \new_[3213]_ ;
  assign \new_[3220]_  = \new_[1673]_  | \new_[1674]_ ;
  assign \new_[3223]_  = \new_[1671]_  | \new_[1672]_ ;
  assign \new_[3224]_  = \new_[3223]_  | \new_[3220]_ ;
  assign \new_[3225]_  = \new_[3224]_  | \new_[3217]_ ;
  assign \new_[3228]_  = \new_[1669]_  | \new_[1670]_ ;
  assign \new_[3231]_  = \new_[1667]_  | \new_[1668]_ ;
  assign \new_[3232]_  = \new_[3231]_  | \new_[3228]_ ;
  assign \new_[3235]_  = \new_[1665]_  | \new_[1666]_ ;
  assign \new_[3239]_  = \new_[1662]_  | \new_[1663]_ ;
  assign \new_[3240]_  = \new_[1664]_  | \new_[3239]_ ;
  assign \new_[3241]_  = \new_[3240]_  | \new_[3235]_ ;
  assign \new_[3242]_  = \new_[3241]_  | \new_[3232]_ ;
  assign \new_[3243]_  = \new_[3242]_  | \new_[3225]_ ;
  assign \new_[3246]_  = \new_[1660]_  | \new_[1661]_ ;
  assign \new_[3249]_  = \new_[1658]_  | \new_[1659]_ ;
  assign \new_[3250]_  = \new_[3249]_  | \new_[3246]_ ;
  assign \new_[3253]_  = \new_[1656]_  | \new_[1657]_ ;
  assign \new_[3257]_  = \new_[1653]_  | \new_[1654]_ ;
  assign \new_[3258]_  = \new_[1655]_  | \new_[3257]_ ;
  assign \new_[3259]_  = \new_[3258]_  | \new_[3253]_ ;
  assign \new_[3260]_  = \new_[3259]_  | \new_[3250]_ ;
  assign \new_[3263]_  = \new_[1651]_  | \new_[1652]_ ;
  assign \new_[3266]_  = \new_[1649]_  | \new_[1650]_ ;
  assign \new_[3267]_  = \new_[3266]_  | \new_[3263]_ ;
  assign \new_[3270]_  = \new_[1647]_  | \new_[1648]_ ;
  assign \new_[3274]_  = \new_[1644]_  | \new_[1645]_ ;
  assign \new_[3275]_  = \new_[1646]_  | \new_[3274]_ ;
  assign \new_[3276]_  = \new_[3275]_  | \new_[3270]_ ;
  assign \new_[3277]_  = \new_[3276]_  | \new_[3267]_ ;
  assign \new_[3278]_  = \new_[3277]_  | \new_[3260]_ ;
  assign \new_[3279]_  = \new_[3278]_  | \new_[3243]_ ;
  assign \new_[3280]_  = \new_[3279]_  | \new_[3210]_ ;
  assign \new_[3281]_  = \new_[3280]_  | \new_[3143]_ ;
  assign \new_[3282]_  = \new_[3281]_  | \new_[3008]_ ;
  assign \new_[3283]_  = \new_[3282]_  | \new_[2735]_ ;
  assign \new_[3286]_  = \new_[1642]_  | \new_[1643]_ ;
  assign \new_[3289]_  = \new_[1640]_  | \new_[1641]_ ;
  assign \new_[3290]_  = \new_[3289]_  | \new_[3286]_ ;
  assign \new_[3293]_  = \new_[1638]_  | \new_[1639]_ ;
  assign \new_[3296]_  = \new_[1636]_  | \new_[1637]_ ;
  assign \new_[3297]_  = \new_[3296]_  | \new_[3293]_ ;
  assign \new_[3298]_  = \new_[3297]_  | \new_[3290]_ ;
  assign \new_[3301]_  = \new_[1634]_  | \new_[1635]_ ;
  assign \new_[3304]_  = \new_[1632]_  | \new_[1633]_ ;
  assign \new_[3305]_  = \new_[3304]_  | \new_[3301]_ ;
  assign \new_[3308]_  = \new_[1630]_  | \new_[1631]_ ;
  assign \new_[3312]_  = \new_[1627]_  | \new_[1628]_ ;
  assign \new_[3313]_  = \new_[1629]_  | \new_[3312]_ ;
  assign \new_[3314]_  = \new_[3313]_  | \new_[3308]_ ;
  assign \new_[3315]_  = \new_[3314]_  | \new_[3305]_ ;
  assign \new_[3316]_  = \new_[3315]_  | \new_[3298]_ ;
  assign \new_[3319]_  = \new_[1625]_  | \new_[1626]_ ;
  assign \new_[3322]_  = \new_[1623]_  | \new_[1624]_ ;
  assign \new_[3323]_  = \new_[3322]_  | \new_[3319]_ ;
  assign \new_[3326]_  = \new_[1621]_  | \new_[1622]_ ;
  assign \new_[3329]_  = \new_[1619]_  | \new_[1620]_ ;
  assign \new_[3330]_  = \new_[3329]_  | \new_[3326]_ ;
  assign \new_[3331]_  = \new_[3330]_  | \new_[3323]_ ;
  assign \new_[3334]_  = \new_[1617]_  | \new_[1618]_ ;
  assign \new_[3337]_  = \new_[1615]_  | \new_[1616]_ ;
  assign \new_[3338]_  = \new_[3337]_  | \new_[3334]_ ;
  assign \new_[3341]_  = \new_[1613]_  | \new_[1614]_ ;
  assign \new_[3345]_  = \new_[1610]_  | \new_[1611]_ ;
  assign \new_[3346]_  = \new_[1612]_  | \new_[3345]_ ;
  assign \new_[3347]_  = \new_[3346]_  | \new_[3341]_ ;
  assign \new_[3348]_  = \new_[3347]_  | \new_[3338]_ ;
  assign \new_[3349]_  = \new_[3348]_  | \new_[3331]_ ;
  assign \new_[3350]_  = \new_[3349]_  | \new_[3316]_ ;
  assign \new_[3353]_  = \new_[1608]_  | \new_[1609]_ ;
  assign \new_[3356]_  = \new_[1606]_  | \new_[1607]_ ;
  assign \new_[3357]_  = \new_[3356]_  | \new_[3353]_ ;
  assign \new_[3360]_  = \new_[1604]_  | \new_[1605]_ ;
  assign \new_[3363]_  = \new_[1602]_  | \new_[1603]_ ;
  assign \new_[3364]_  = \new_[3363]_  | \new_[3360]_ ;
  assign \new_[3365]_  = \new_[3364]_  | \new_[3357]_ ;
  assign \new_[3368]_  = \new_[1600]_  | \new_[1601]_ ;
  assign \new_[3371]_  = \new_[1598]_  | \new_[1599]_ ;
  assign \new_[3372]_  = \new_[3371]_  | \new_[3368]_ ;
  assign \new_[3375]_  = \new_[1596]_  | \new_[1597]_ ;
  assign \new_[3379]_  = \new_[1593]_  | \new_[1594]_ ;
  assign \new_[3380]_  = \new_[1595]_  | \new_[3379]_ ;
  assign \new_[3381]_  = \new_[3380]_  | \new_[3375]_ ;
  assign \new_[3382]_  = \new_[3381]_  | \new_[3372]_ ;
  assign \new_[3383]_  = \new_[3382]_  | \new_[3365]_ ;
  assign \new_[3386]_  = \new_[1591]_  | \new_[1592]_ ;
  assign \new_[3389]_  = \new_[1589]_  | \new_[1590]_ ;
  assign \new_[3390]_  = \new_[3389]_  | \new_[3386]_ ;
  assign \new_[3393]_  = \new_[1587]_  | \new_[1588]_ ;
  assign \new_[3396]_  = \new_[1585]_  | \new_[1586]_ ;
  assign \new_[3397]_  = \new_[3396]_  | \new_[3393]_ ;
  assign \new_[3398]_  = \new_[3397]_  | \new_[3390]_ ;
  assign \new_[3401]_  = \new_[1583]_  | \new_[1584]_ ;
  assign \new_[3404]_  = \new_[1581]_  | \new_[1582]_ ;
  assign \new_[3405]_  = \new_[3404]_  | \new_[3401]_ ;
  assign \new_[3408]_  = \new_[1579]_  | \new_[1580]_ ;
  assign \new_[3412]_  = \new_[1576]_  | \new_[1577]_ ;
  assign \new_[3413]_  = \new_[1578]_  | \new_[3412]_ ;
  assign \new_[3414]_  = \new_[3413]_  | \new_[3408]_ ;
  assign \new_[3415]_  = \new_[3414]_  | \new_[3405]_ ;
  assign \new_[3416]_  = \new_[3415]_  | \new_[3398]_ ;
  assign \new_[3417]_  = \new_[3416]_  | \new_[3383]_ ;
  assign \new_[3418]_  = \new_[3417]_  | \new_[3350]_ ;
  assign \new_[3421]_  = \new_[1574]_  | \new_[1575]_ ;
  assign \new_[3424]_  = \new_[1572]_  | \new_[1573]_ ;
  assign \new_[3425]_  = \new_[3424]_  | \new_[3421]_ ;
  assign \new_[3428]_  = \new_[1570]_  | \new_[1571]_ ;
  assign \new_[3431]_  = \new_[1568]_  | \new_[1569]_ ;
  assign \new_[3432]_  = \new_[3431]_  | \new_[3428]_ ;
  assign \new_[3433]_  = \new_[3432]_  | \new_[3425]_ ;
  assign \new_[3436]_  = \new_[1566]_  | \new_[1567]_ ;
  assign \new_[3439]_  = \new_[1564]_  | \new_[1565]_ ;
  assign \new_[3440]_  = \new_[3439]_  | \new_[3436]_ ;
  assign \new_[3443]_  = \new_[1562]_  | \new_[1563]_ ;
  assign \new_[3447]_  = \new_[1559]_  | \new_[1560]_ ;
  assign \new_[3448]_  = \new_[1561]_  | \new_[3447]_ ;
  assign \new_[3449]_  = \new_[3448]_  | \new_[3443]_ ;
  assign \new_[3450]_  = \new_[3449]_  | \new_[3440]_ ;
  assign \new_[3451]_  = \new_[3450]_  | \new_[3433]_ ;
  assign \new_[3454]_  = \new_[1557]_  | \new_[1558]_ ;
  assign \new_[3457]_  = \new_[1555]_  | \new_[1556]_ ;
  assign \new_[3458]_  = \new_[3457]_  | \new_[3454]_ ;
  assign \new_[3461]_  = \new_[1553]_  | \new_[1554]_ ;
  assign \new_[3464]_  = \new_[1551]_  | \new_[1552]_ ;
  assign \new_[3465]_  = \new_[3464]_  | \new_[3461]_ ;
  assign \new_[3466]_  = \new_[3465]_  | \new_[3458]_ ;
  assign \new_[3469]_  = \new_[1549]_  | \new_[1550]_ ;
  assign \new_[3472]_  = \new_[1547]_  | \new_[1548]_ ;
  assign \new_[3473]_  = \new_[3472]_  | \new_[3469]_ ;
  assign \new_[3476]_  = \new_[1545]_  | \new_[1546]_ ;
  assign \new_[3480]_  = \new_[1542]_  | \new_[1543]_ ;
  assign \new_[3481]_  = \new_[1544]_  | \new_[3480]_ ;
  assign \new_[3482]_  = \new_[3481]_  | \new_[3476]_ ;
  assign \new_[3483]_  = \new_[3482]_  | \new_[3473]_ ;
  assign \new_[3484]_  = \new_[3483]_  | \new_[3466]_ ;
  assign \new_[3485]_  = \new_[3484]_  | \new_[3451]_ ;
  assign \new_[3488]_  = \new_[1540]_  | \new_[1541]_ ;
  assign \new_[3491]_  = \new_[1538]_  | \new_[1539]_ ;
  assign \new_[3492]_  = \new_[3491]_  | \new_[3488]_ ;
  assign \new_[3495]_  = \new_[1536]_  | \new_[1537]_ ;
  assign \new_[3498]_  = \new_[1534]_  | \new_[1535]_ ;
  assign \new_[3499]_  = \new_[3498]_  | \new_[3495]_ ;
  assign \new_[3500]_  = \new_[3499]_  | \new_[3492]_ ;
  assign \new_[3503]_  = \new_[1532]_  | \new_[1533]_ ;
  assign \new_[3506]_  = \new_[1530]_  | \new_[1531]_ ;
  assign \new_[3507]_  = \new_[3506]_  | \new_[3503]_ ;
  assign \new_[3510]_  = \new_[1528]_  | \new_[1529]_ ;
  assign \new_[3514]_  = \new_[1525]_  | \new_[1526]_ ;
  assign \new_[3515]_  = \new_[1527]_  | \new_[3514]_ ;
  assign \new_[3516]_  = \new_[3515]_  | \new_[3510]_ ;
  assign \new_[3517]_  = \new_[3516]_  | \new_[3507]_ ;
  assign \new_[3518]_  = \new_[3517]_  | \new_[3500]_ ;
  assign \new_[3521]_  = \new_[1523]_  | \new_[1524]_ ;
  assign \new_[3524]_  = \new_[1521]_  | \new_[1522]_ ;
  assign \new_[3525]_  = \new_[3524]_  | \new_[3521]_ ;
  assign \new_[3528]_  = \new_[1519]_  | \new_[1520]_ ;
  assign \new_[3532]_  = \new_[1516]_  | \new_[1517]_ ;
  assign \new_[3533]_  = \new_[1518]_  | \new_[3532]_ ;
  assign \new_[3534]_  = \new_[3533]_  | \new_[3528]_ ;
  assign \new_[3535]_  = \new_[3534]_  | \new_[3525]_ ;
  assign \new_[3538]_  = \new_[1514]_  | \new_[1515]_ ;
  assign \new_[3541]_  = \new_[1512]_  | \new_[1513]_ ;
  assign \new_[3542]_  = \new_[3541]_  | \new_[3538]_ ;
  assign \new_[3545]_  = \new_[1510]_  | \new_[1511]_ ;
  assign \new_[3549]_  = \new_[1507]_  | \new_[1508]_ ;
  assign \new_[3550]_  = \new_[1509]_  | \new_[3549]_ ;
  assign \new_[3551]_  = \new_[3550]_  | \new_[3545]_ ;
  assign \new_[3552]_  = \new_[3551]_  | \new_[3542]_ ;
  assign \new_[3553]_  = \new_[3552]_  | \new_[3535]_ ;
  assign \new_[3554]_  = \new_[3553]_  | \new_[3518]_ ;
  assign \new_[3555]_  = \new_[3554]_  | \new_[3485]_ ;
  assign \new_[3556]_  = \new_[3555]_  | \new_[3418]_ ;
  assign \new_[3559]_  = \new_[1505]_  | \new_[1506]_ ;
  assign \new_[3562]_  = \new_[1503]_  | \new_[1504]_ ;
  assign \new_[3563]_  = \new_[3562]_  | \new_[3559]_ ;
  assign \new_[3566]_  = \new_[1501]_  | \new_[1502]_ ;
  assign \new_[3569]_  = \new_[1499]_  | \new_[1500]_ ;
  assign \new_[3570]_  = \new_[3569]_  | \new_[3566]_ ;
  assign \new_[3571]_  = \new_[3570]_  | \new_[3563]_ ;
  assign \new_[3574]_  = \new_[1497]_  | \new_[1498]_ ;
  assign \new_[3577]_  = \new_[1495]_  | \new_[1496]_ ;
  assign \new_[3578]_  = \new_[3577]_  | \new_[3574]_ ;
  assign \new_[3581]_  = \new_[1493]_  | \new_[1494]_ ;
  assign \new_[3585]_  = \new_[1490]_  | \new_[1491]_ ;
  assign \new_[3586]_  = \new_[1492]_  | \new_[3585]_ ;
  assign \new_[3587]_  = \new_[3586]_  | \new_[3581]_ ;
  assign \new_[3588]_  = \new_[3587]_  | \new_[3578]_ ;
  assign \new_[3589]_  = \new_[3588]_  | \new_[3571]_ ;
  assign \new_[3592]_  = \new_[1488]_  | \new_[1489]_ ;
  assign \new_[3595]_  = \new_[1486]_  | \new_[1487]_ ;
  assign \new_[3596]_  = \new_[3595]_  | \new_[3592]_ ;
  assign \new_[3599]_  = \new_[1484]_  | \new_[1485]_ ;
  assign \new_[3602]_  = \new_[1482]_  | \new_[1483]_ ;
  assign \new_[3603]_  = \new_[3602]_  | \new_[3599]_ ;
  assign \new_[3604]_  = \new_[3603]_  | \new_[3596]_ ;
  assign \new_[3607]_  = \new_[1480]_  | \new_[1481]_ ;
  assign \new_[3610]_  = \new_[1478]_  | \new_[1479]_ ;
  assign \new_[3611]_  = \new_[3610]_  | \new_[3607]_ ;
  assign \new_[3614]_  = \new_[1476]_  | \new_[1477]_ ;
  assign \new_[3618]_  = \new_[1473]_  | \new_[1474]_ ;
  assign \new_[3619]_  = \new_[1475]_  | \new_[3618]_ ;
  assign \new_[3620]_  = \new_[3619]_  | \new_[3614]_ ;
  assign \new_[3621]_  = \new_[3620]_  | \new_[3611]_ ;
  assign \new_[3622]_  = \new_[3621]_  | \new_[3604]_ ;
  assign \new_[3623]_  = \new_[3622]_  | \new_[3589]_ ;
  assign \new_[3626]_  = \new_[1471]_  | \new_[1472]_ ;
  assign \new_[3629]_  = \new_[1469]_  | \new_[1470]_ ;
  assign \new_[3630]_  = \new_[3629]_  | \new_[3626]_ ;
  assign \new_[3633]_  = \new_[1467]_  | \new_[1468]_ ;
  assign \new_[3636]_  = \new_[1465]_  | \new_[1466]_ ;
  assign \new_[3637]_  = \new_[3636]_  | \new_[3633]_ ;
  assign \new_[3638]_  = \new_[3637]_  | \new_[3630]_ ;
  assign \new_[3641]_  = \new_[1463]_  | \new_[1464]_ ;
  assign \new_[3644]_  = \new_[1461]_  | \new_[1462]_ ;
  assign \new_[3645]_  = \new_[3644]_  | \new_[3641]_ ;
  assign \new_[3648]_  = \new_[1459]_  | \new_[1460]_ ;
  assign \new_[3652]_  = \new_[1456]_  | \new_[1457]_ ;
  assign \new_[3653]_  = \new_[1458]_  | \new_[3652]_ ;
  assign \new_[3654]_  = \new_[3653]_  | \new_[3648]_ ;
  assign \new_[3655]_  = \new_[3654]_  | \new_[3645]_ ;
  assign \new_[3656]_  = \new_[3655]_  | \new_[3638]_ ;
  assign \new_[3659]_  = \new_[1454]_  | \new_[1455]_ ;
  assign \new_[3662]_  = \new_[1452]_  | \new_[1453]_ ;
  assign \new_[3663]_  = \new_[3662]_  | \new_[3659]_ ;
  assign \new_[3666]_  = \new_[1450]_  | \new_[1451]_ ;
  assign \new_[3669]_  = \new_[1448]_  | \new_[1449]_ ;
  assign \new_[3670]_  = \new_[3669]_  | \new_[3666]_ ;
  assign \new_[3671]_  = \new_[3670]_  | \new_[3663]_ ;
  assign \new_[3674]_  = \new_[1446]_  | \new_[1447]_ ;
  assign \new_[3677]_  = \new_[1444]_  | \new_[1445]_ ;
  assign \new_[3678]_  = \new_[3677]_  | \new_[3674]_ ;
  assign \new_[3681]_  = \new_[1442]_  | \new_[1443]_ ;
  assign \new_[3685]_  = \new_[1439]_  | \new_[1440]_ ;
  assign \new_[3686]_  = \new_[1441]_  | \new_[3685]_ ;
  assign \new_[3687]_  = \new_[3686]_  | \new_[3681]_ ;
  assign \new_[3688]_  = \new_[3687]_  | \new_[3678]_ ;
  assign \new_[3689]_  = \new_[3688]_  | \new_[3671]_ ;
  assign \new_[3690]_  = \new_[3689]_  | \new_[3656]_ ;
  assign \new_[3691]_  = \new_[3690]_  | \new_[3623]_ ;
  assign \new_[3694]_  = \new_[1437]_  | \new_[1438]_ ;
  assign \new_[3697]_  = \new_[1435]_  | \new_[1436]_ ;
  assign \new_[3698]_  = \new_[3697]_  | \new_[3694]_ ;
  assign \new_[3701]_  = \new_[1433]_  | \new_[1434]_ ;
  assign \new_[3704]_  = \new_[1431]_  | \new_[1432]_ ;
  assign \new_[3705]_  = \new_[3704]_  | \new_[3701]_ ;
  assign \new_[3706]_  = \new_[3705]_  | \new_[3698]_ ;
  assign \new_[3709]_  = \new_[1429]_  | \new_[1430]_ ;
  assign \new_[3712]_  = \new_[1427]_  | \new_[1428]_ ;
  assign \new_[3713]_  = \new_[3712]_  | \new_[3709]_ ;
  assign \new_[3716]_  = \new_[1425]_  | \new_[1426]_ ;
  assign \new_[3720]_  = \new_[1422]_  | \new_[1423]_ ;
  assign \new_[3721]_  = \new_[1424]_  | \new_[3720]_ ;
  assign \new_[3722]_  = \new_[3721]_  | \new_[3716]_ ;
  assign \new_[3723]_  = \new_[3722]_  | \new_[3713]_ ;
  assign \new_[3724]_  = \new_[3723]_  | \new_[3706]_ ;
  assign \new_[3727]_  = \new_[1420]_  | \new_[1421]_ ;
  assign \new_[3730]_  = \new_[1418]_  | \new_[1419]_ ;
  assign \new_[3731]_  = \new_[3730]_  | \new_[3727]_ ;
  assign \new_[3734]_  = \new_[1416]_  | \new_[1417]_ ;
  assign \new_[3737]_  = \new_[1414]_  | \new_[1415]_ ;
  assign \new_[3738]_  = \new_[3737]_  | \new_[3734]_ ;
  assign \new_[3739]_  = \new_[3738]_  | \new_[3731]_ ;
  assign \new_[3742]_  = \new_[1412]_  | \new_[1413]_ ;
  assign \new_[3745]_  = \new_[1410]_  | \new_[1411]_ ;
  assign \new_[3746]_  = \new_[3745]_  | \new_[3742]_ ;
  assign \new_[3749]_  = \new_[1408]_  | \new_[1409]_ ;
  assign \new_[3753]_  = \new_[1405]_  | \new_[1406]_ ;
  assign \new_[3754]_  = \new_[1407]_  | \new_[3753]_ ;
  assign \new_[3755]_  = \new_[3754]_  | \new_[3749]_ ;
  assign \new_[3756]_  = \new_[3755]_  | \new_[3746]_ ;
  assign \new_[3757]_  = \new_[3756]_  | \new_[3739]_ ;
  assign \new_[3758]_  = \new_[3757]_  | \new_[3724]_ ;
  assign \new_[3761]_  = \new_[1403]_  | \new_[1404]_ ;
  assign \new_[3764]_  = \new_[1401]_  | \new_[1402]_ ;
  assign \new_[3765]_  = \new_[3764]_  | \new_[3761]_ ;
  assign \new_[3768]_  = \new_[1399]_  | \new_[1400]_ ;
  assign \new_[3771]_  = \new_[1397]_  | \new_[1398]_ ;
  assign \new_[3772]_  = \new_[3771]_  | \new_[3768]_ ;
  assign \new_[3773]_  = \new_[3772]_  | \new_[3765]_ ;
  assign \new_[3776]_  = \new_[1395]_  | \new_[1396]_ ;
  assign \new_[3779]_  = \new_[1393]_  | \new_[1394]_ ;
  assign \new_[3780]_  = \new_[3779]_  | \new_[3776]_ ;
  assign \new_[3783]_  = \new_[1391]_  | \new_[1392]_ ;
  assign \new_[3787]_  = \new_[1388]_  | \new_[1389]_ ;
  assign \new_[3788]_  = \new_[1390]_  | \new_[3787]_ ;
  assign \new_[3789]_  = \new_[3788]_  | \new_[3783]_ ;
  assign \new_[3790]_  = \new_[3789]_  | \new_[3780]_ ;
  assign \new_[3791]_  = \new_[3790]_  | \new_[3773]_ ;
  assign \new_[3794]_  = \new_[1386]_  | \new_[1387]_ ;
  assign \new_[3797]_  = \new_[1384]_  | \new_[1385]_ ;
  assign \new_[3798]_  = \new_[3797]_  | \new_[3794]_ ;
  assign \new_[3801]_  = \new_[1382]_  | \new_[1383]_ ;
  assign \new_[3805]_  = \new_[1379]_  | \new_[1380]_ ;
  assign \new_[3806]_  = \new_[1381]_  | \new_[3805]_ ;
  assign \new_[3807]_  = \new_[3806]_  | \new_[3801]_ ;
  assign \new_[3808]_  = \new_[3807]_  | \new_[3798]_ ;
  assign \new_[3811]_  = \new_[1377]_  | \new_[1378]_ ;
  assign \new_[3814]_  = \new_[1375]_  | \new_[1376]_ ;
  assign \new_[3815]_  = \new_[3814]_  | \new_[3811]_ ;
  assign \new_[3818]_  = \new_[1373]_  | \new_[1374]_ ;
  assign \new_[3822]_  = \new_[1370]_  | \new_[1371]_ ;
  assign \new_[3823]_  = \new_[1372]_  | \new_[3822]_ ;
  assign \new_[3824]_  = \new_[3823]_  | \new_[3818]_ ;
  assign \new_[3825]_  = \new_[3824]_  | \new_[3815]_ ;
  assign \new_[3826]_  = \new_[3825]_  | \new_[3808]_ ;
  assign \new_[3827]_  = \new_[3826]_  | \new_[3791]_ ;
  assign \new_[3828]_  = \new_[3827]_  | \new_[3758]_ ;
  assign \new_[3829]_  = \new_[3828]_  | \new_[3691]_ ;
  assign \new_[3830]_  = \new_[3829]_  | \new_[3556]_ ;
  assign \new_[3833]_  = \new_[1368]_  | \new_[1369]_ ;
  assign \new_[3836]_  = \new_[1366]_  | \new_[1367]_ ;
  assign \new_[3837]_  = \new_[3836]_  | \new_[3833]_ ;
  assign \new_[3840]_  = \new_[1364]_  | \new_[1365]_ ;
  assign \new_[3843]_  = \new_[1362]_  | \new_[1363]_ ;
  assign \new_[3844]_  = \new_[3843]_  | \new_[3840]_ ;
  assign \new_[3845]_  = \new_[3844]_  | \new_[3837]_ ;
  assign \new_[3848]_  = \new_[1360]_  | \new_[1361]_ ;
  assign \new_[3851]_  = \new_[1358]_  | \new_[1359]_ ;
  assign \new_[3852]_  = \new_[3851]_  | \new_[3848]_ ;
  assign \new_[3855]_  = \new_[1356]_  | \new_[1357]_ ;
  assign \new_[3859]_  = \new_[1353]_  | \new_[1354]_ ;
  assign \new_[3860]_  = \new_[1355]_  | \new_[3859]_ ;
  assign \new_[3861]_  = \new_[3860]_  | \new_[3855]_ ;
  assign \new_[3862]_  = \new_[3861]_  | \new_[3852]_ ;
  assign \new_[3863]_  = \new_[3862]_  | \new_[3845]_ ;
  assign \new_[3866]_  = \new_[1351]_  | \new_[1352]_ ;
  assign \new_[3869]_  = \new_[1349]_  | \new_[1350]_ ;
  assign \new_[3870]_  = \new_[3869]_  | \new_[3866]_ ;
  assign \new_[3873]_  = \new_[1347]_  | \new_[1348]_ ;
  assign \new_[3876]_  = \new_[1345]_  | \new_[1346]_ ;
  assign \new_[3877]_  = \new_[3876]_  | \new_[3873]_ ;
  assign \new_[3878]_  = \new_[3877]_  | \new_[3870]_ ;
  assign \new_[3881]_  = \new_[1343]_  | \new_[1344]_ ;
  assign \new_[3884]_  = \new_[1341]_  | \new_[1342]_ ;
  assign \new_[3885]_  = \new_[3884]_  | \new_[3881]_ ;
  assign \new_[3888]_  = \new_[1339]_  | \new_[1340]_ ;
  assign \new_[3892]_  = \new_[1336]_  | \new_[1337]_ ;
  assign \new_[3893]_  = \new_[1338]_  | \new_[3892]_ ;
  assign \new_[3894]_  = \new_[3893]_  | \new_[3888]_ ;
  assign \new_[3895]_  = \new_[3894]_  | \new_[3885]_ ;
  assign \new_[3896]_  = \new_[3895]_  | \new_[3878]_ ;
  assign \new_[3897]_  = \new_[3896]_  | \new_[3863]_ ;
  assign \new_[3900]_  = \new_[1334]_  | \new_[1335]_ ;
  assign \new_[3903]_  = \new_[1332]_  | \new_[1333]_ ;
  assign \new_[3904]_  = \new_[3903]_  | \new_[3900]_ ;
  assign \new_[3907]_  = \new_[1330]_  | \new_[1331]_ ;
  assign \new_[3910]_  = \new_[1328]_  | \new_[1329]_ ;
  assign \new_[3911]_  = \new_[3910]_  | \new_[3907]_ ;
  assign \new_[3912]_  = \new_[3911]_  | \new_[3904]_ ;
  assign \new_[3915]_  = \new_[1326]_  | \new_[1327]_ ;
  assign \new_[3918]_  = \new_[1324]_  | \new_[1325]_ ;
  assign \new_[3919]_  = \new_[3918]_  | \new_[3915]_ ;
  assign \new_[3922]_  = \new_[1322]_  | \new_[1323]_ ;
  assign \new_[3926]_  = \new_[1319]_  | \new_[1320]_ ;
  assign \new_[3927]_  = \new_[1321]_  | \new_[3926]_ ;
  assign \new_[3928]_  = \new_[3927]_  | \new_[3922]_ ;
  assign \new_[3929]_  = \new_[3928]_  | \new_[3919]_ ;
  assign \new_[3930]_  = \new_[3929]_  | \new_[3912]_ ;
  assign \new_[3933]_  = \new_[1317]_  | \new_[1318]_ ;
  assign \new_[3936]_  = \new_[1315]_  | \new_[1316]_ ;
  assign \new_[3937]_  = \new_[3936]_  | \new_[3933]_ ;
  assign \new_[3940]_  = \new_[1313]_  | \new_[1314]_ ;
  assign \new_[3943]_  = \new_[1311]_  | \new_[1312]_ ;
  assign \new_[3944]_  = \new_[3943]_  | \new_[3940]_ ;
  assign \new_[3945]_  = \new_[3944]_  | \new_[3937]_ ;
  assign \new_[3948]_  = \new_[1309]_  | \new_[1310]_ ;
  assign \new_[3951]_  = \new_[1307]_  | \new_[1308]_ ;
  assign \new_[3952]_  = \new_[3951]_  | \new_[3948]_ ;
  assign \new_[3955]_  = \new_[1305]_  | \new_[1306]_ ;
  assign \new_[3959]_  = \new_[1302]_  | \new_[1303]_ ;
  assign \new_[3960]_  = \new_[1304]_  | \new_[3959]_ ;
  assign \new_[3961]_  = \new_[3960]_  | \new_[3955]_ ;
  assign \new_[3962]_  = \new_[3961]_  | \new_[3952]_ ;
  assign \new_[3963]_  = \new_[3962]_  | \new_[3945]_ ;
  assign \new_[3964]_  = \new_[3963]_  | \new_[3930]_ ;
  assign \new_[3965]_  = \new_[3964]_  | \new_[3897]_ ;
  assign \new_[3968]_  = \new_[1300]_  | \new_[1301]_ ;
  assign \new_[3971]_  = \new_[1298]_  | \new_[1299]_ ;
  assign \new_[3972]_  = \new_[3971]_  | \new_[3968]_ ;
  assign \new_[3975]_  = \new_[1296]_  | \new_[1297]_ ;
  assign \new_[3978]_  = \new_[1294]_  | \new_[1295]_ ;
  assign \new_[3979]_  = \new_[3978]_  | \new_[3975]_ ;
  assign \new_[3980]_  = \new_[3979]_  | \new_[3972]_ ;
  assign \new_[3983]_  = \new_[1292]_  | \new_[1293]_ ;
  assign \new_[3986]_  = \new_[1290]_  | \new_[1291]_ ;
  assign \new_[3987]_  = \new_[3986]_  | \new_[3983]_ ;
  assign \new_[3990]_  = \new_[1288]_  | \new_[1289]_ ;
  assign \new_[3994]_  = \new_[1285]_  | \new_[1286]_ ;
  assign \new_[3995]_  = \new_[1287]_  | \new_[3994]_ ;
  assign \new_[3996]_  = \new_[3995]_  | \new_[3990]_ ;
  assign \new_[3997]_  = \new_[3996]_  | \new_[3987]_ ;
  assign \new_[3998]_  = \new_[3997]_  | \new_[3980]_ ;
  assign \new_[4001]_  = \new_[1283]_  | \new_[1284]_ ;
  assign \new_[4004]_  = \new_[1281]_  | \new_[1282]_ ;
  assign \new_[4005]_  = \new_[4004]_  | \new_[4001]_ ;
  assign \new_[4008]_  = \new_[1279]_  | \new_[1280]_ ;
  assign \new_[4011]_  = \new_[1277]_  | \new_[1278]_ ;
  assign \new_[4012]_  = \new_[4011]_  | \new_[4008]_ ;
  assign \new_[4013]_  = \new_[4012]_  | \new_[4005]_ ;
  assign \new_[4016]_  = \new_[1275]_  | \new_[1276]_ ;
  assign \new_[4019]_  = \new_[1273]_  | \new_[1274]_ ;
  assign \new_[4020]_  = \new_[4019]_  | \new_[4016]_ ;
  assign \new_[4023]_  = \new_[1271]_  | \new_[1272]_ ;
  assign \new_[4027]_  = \new_[1268]_  | \new_[1269]_ ;
  assign \new_[4028]_  = \new_[1270]_  | \new_[4027]_ ;
  assign \new_[4029]_  = \new_[4028]_  | \new_[4023]_ ;
  assign \new_[4030]_  = \new_[4029]_  | \new_[4020]_ ;
  assign \new_[4031]_  = \new_[4030]_  | \new_[4013]_ ;
  assign \new_[4032]_  = \new_[4031]_  | \new_[3998]_ ;
  assign \new_[4035]_  = \new_[1266]_  | \new_[1267]_ ;
  assign \new_[4038]_  = \new_[1264]_  | \new_[1265]_ ;
  assign \new_[4039]_  = \new_[4038]_  | \new_[4035]_ ;
  assign \new_[4042]_  = \new_[1262]_  | \new_[1263]_ ;
  assign \new_[4045]_  = \new_[1260]_  | \new_[1261]_ ;
  assign \new_[4046]_  = \new_[4045]_  | \new_[4042]_ ;
  assign \new_[4047]_  = \new_[4046]_  | \new_[4039]_ ;
  assign \new_[4050]_  = \new_[1258]_  | \new_[1259]_ ;
  assign \new_[4053]_  = \new_[1256]_  | \new_[1257]_ ;
  assign \new_[4054]_  = \new_[4053]_  | \new_[4050]_ ;
  assign \new_[4057]_  = \new_[1254]_  | \new_[1255]_ ;
  assign \new_[4061]_  = \new_[1251]_  | \new_[1252]_ ;
  assign \new_[4062]_  = \new_[1253]_  | \new_[4061]_ ;
  assign \new_[4063]_  = \new_[4062]_  | \new_[4057]_ ;
  assign \new_[4064]_  = \new_[4063]_  | \new_[4054]_ ;
  assign \new_[4065]_  = \new_[4064]_  | \new_[4047]_ ;
  assign \new_[4068]_  = \new_[1249]_  | \new_[1250]_ ;
  assign \new_[4071]_  = \new_[1247]_  | \new_[1248]_ ;
  assign \new_[4072]_  = \new_[4071]_  | \new_[4068]_ ;
  assign \new_[4075]_  = \new_[1245]_  | \new_[1246]_ ;
  assign \new_[4079]_  = \new_[1242]_  | \new_[1243]_ ;
  assign \new_[4080]_  = \new_[1244]_  | \new_[4079]_ ;
  assign \new_[4081]_  = \new_[4080]_  | \new_[4075]_ ;
  assign \new_[4082]_  = \new_[4081]_  | \new_[4072]_ ;
  assign \new_[4085]_  = \new_[1240]_  | \new_[1241]_ ;
  assign \new_[4088]_  = \new_[1238]_  | \new_[1239]_ ;
  assign \new_[4089]_  = \new_[4088]_  | \new_[4085]_ ;
  assign \new_[4092]_  = \new_[1236]_  | \new_[1237]_ ;
  assign \new_[4096]_  = \new_[1233]_  | \new_[1234]_ ;
  assign \new_[4097]_  = \new_[1235]_  | \new_[4096]_ ;
  assign \new_[4098]_  = \new_[4097]_  | \new_[4092]_ ;
  assign \new_[4099]_  = \new_[4098]_  | \new_[4089]_ ;
  assign \new_[4100]_  = \new_[4099]_  | \new_[4082]_ ;
  assign \new_[4101]_  = \new_[4100]_  | \new_[4065]_ ;
  assign \new_[4102]_  = \new_[4101]_  | \new_[4032]_ ;
  assign \new_[4103]_  = \new_[4102]_  | \new_[3965]_ ;
  assign \new_[4106]_  = \new_[1231]_  | \new_[1232]_ ;
  assign \new_[4109]_  = \new_[1229]_  | \new_[1230]_ ;
  assign \new_[4110]_  = \new_[4109]_  | \new_[4106]_ ;
  assign \new_[4113]_  = \new_[1227]_  | \new_[1228]_ ;
  assign \new_[4116]_  = \new_[1225]_  | \new_[1226]_ ;
  assign \new_[4117]_  = \new_[4116]_  | \new_[4113]_ ;
  assign \new_[4118]_  = \new_[4117]_  | \new_[4110]_ ;
  assign \new_[4121]_  = \new_[1223]_  | \new_[1224]_ ;
  assign \new_[4124]_  = \new_[1221]_  | \new_[1222]_ ;
  assign \new_[4125]_  = \new_[4124]_  | \new_[4121]_ ;
  assign \new_[4128]_  = \new_[1219]_  | \new_[1220]_ ;
  assign \new_[4132]_  = \new_[1216]_  | \new_[1217]_ ;
  assign \new_[4133]_  = \new_[1218]_  | \new_[4132]_ ;
  assign \new_[4134]_  = \new_[4133]_  | \new_[4128]_ ;
  assign \new_[4135]_  = \new_[4134]_  | \new_[4125]_ ;
  assign \new_[4136]_  = \new_[4135]_  | \new_[4118]_ ;
  assign \new_[4139]_  = \new_[1214]_  | \new_[1215]_ ;
  assign \new_[4142]_  = \new_[1212]_  | \new_[1213]_ ;
  assign \new_[4143]_  = \new_[4142]_  | \new_[4139]_ ;
  assign \new_[4146]_  = \new_[1210]_  | \new_[1211]_ ;
  assign \new_[4149]_  = \new_[1208]_  | \new_[1209]_ ;
  assign \new_[4150]_  = \new_[4149]_  | \new_[4146]_ ;
  assign \new_[4151]_  = \new_[4150]_  | \new_[4143]_ ;
  assign \new_[4154]_  = \new_[1206]_  | \new_[1207]_ ;
  assign \new_[4157]_  = \new_[1204]_  | \new_[1205]_ ;
  assign \new_[4158]_  = \new_[4157]_  | \new_[4154]_ ;
  assign \new_[4161]_  = \new_[1202]_  | \new_[1203]_ ;
  assign \new_[4165]_  = \new_[1199]_  | \new_[1200]_ ;
  assign \new_[4166]_  = \new_[1201]_  | \new_[4165]_ ;
  assign \new_[4167]_  = \new_[4166]_  | \new_[4161]_ ;
  assign \new_[4168]_  = \new_[4167]_  | \new_[4158]_ ;
  assign \new_[4169]_  = \new_[4168]_  | \new_[4151]_ ;
  assign \new_[4170]_  = \new_[4169]_  | \new_[4136]_ ;
  assign \new_[4173]_  = \new_[1197]_  | \new_[1198]_ ;
  assign \new_[4176]_  = \new_[1195]_  | \new_[1196]_ ;
  assign \new_[4177]_  = \new_[4176]_  | \new_[4173]_ ;
  assign \new_[4180]_  = \new_[1193]_  | \new_[1194]_ ;
  assign \new_[4183]_  = \new_[1191]_  | \new_[1192]_ ;
  assign \new_[4184]_  = \new_[4183]_  | \new_[4180]_ ;
  assign \new_[4185]_  = \new_[4184]_  | \new_[4177]_ ;
  assign \new_[4188]_  = \new_[1189]_  | \new_[1190]_ ;
  assign \new_[4191]_  = \new_[1187]_  | \new_[1188]_ ;
  assign \new_[4192]_  = \new_[4191]_  | \new_[4188]_ ;
  assign \new_[4195]_  = \new_[1185]_  | \new_[1186]_ ;
  assign \new_[4199]_  = \new_[1182]_  | \new_[1183]_ ;
  assign \new_[4200]_  = \new_[1184]_  | \new_[4199]_ ;
  assign \new_[4201]_  = \new_[4200]_  | \new_[4195]_ ;
  assign \new_[4202]_  = \new_[4201]_  | \new_[4192]_ ;
  assign \new_[4203]_  = \new_[4202]_  | \new_[4185]_ ;
  assign \new_[4206]_  = \new_[1180]_  | \new_[1181]_ ;
  assign \new_[4209]_  = \new_[1178]_  | \new_[1179]_ ;
  assign \new_[4210]_  = \new_[4209]_  | \new_[4206]_ ;
  assign \new_[4213]_  = \new_[1176]_  | \new_[1177]_ ;
  assign \new_[4216]_  = \new_[1174]_  | \new_[1175]_ ;
  assign \new_[4217]_  = \new_[4216]_  | \new_[4213]_ ;
  assign \new_[4218]_  = \new_[4217]_  | \new_[4210]_ ;
  assign \new_[4221]_  = \new_[1172]_  | \new_[1173]_ ;
  assign \new_[4224]_  = \new_[1170]_  | \new_[1171]_ ;
  assign \new_[4225]_  = \new_[4224]_  | \new_[4221]_ ;
  assign \new_[4228]_  = \new_[1168]_  | \new_[1169]_ ;
  assign \new_[4232]_  = \new_[1165]_  | \new_[1166]_ ;
  assign \new_[4233]_  = \new_[1167]_  | \new_[4232]_ ;
  assign \new_[4234]_  = \new_[4233]_  | \new_[4228]_ ;
  assign \new_[4235]_  = \new_[4234]_  | \new_[4225]_ ;
  assign \new_[4236]_  = \new_[4235]_  | \new_[4218]_ ;
  assign \new_[4237]_  = \new_[4236]_  | \new_[4203]_ ;
  assign \new_[4238]_  = \new_[4237]_  | \new_[4170]_ ;
  assign \new_[4241]_  = \new_[1163]_  | \new_[1164]_ ;
  assign \new_[4244]_  = \new_[1161]_  | \new_[1162]_ ;
  assign \new_[4245]_  = \new_[4244]_  | \new_[4241]_ ;
  assign \new_[4248]_  = \new_[1159]_  | \new_[1160]_ ;
  assign \new_[4251]_  = \new_[1157]_  | \new_[1158]_ ;
  assign \new_[4252]_  = \new_[4251]_  | \new_[4248]_ ;
  assign \new_[4253]_  = \new_[4252]_  | \new_[4245]_ ;
  assign \new_[4256]_  = \new_[1155]_  | \new_[1156]_ ;
  assign \new_[4259]_  = \new_[1153]_  | \new_[1154]_ ;
  assign \new_[4260]_  = \new_[4259]_  | \new_[4256]_ ;
  assign \new_[4263]_  = \new_[1151]_  | \new_[1152]_ ;
  assign \new_[4267]_  = \new_[1148]_  | \new_[1149]_ ;
  assign \new_[4268]_  = \new_[1150]_  | \new_[4267]_ ;
  assign \new_[4269]_  = \new_[4268]_  | \new_[4263]_ ;
  assign \new_[4270]_  = \new_[4269]_  | \new_[4260]_ ;
  assign \new_[4271]_  = \new_[4270]_  | \new_[4253]_ ;
  assign \new_[4274]_  = \new_[1146]_  | \new_[1147]_ ;
  assign \new_[4277]_  = \new_[1144]_  | \new_[1145]_ ;
  assign \new_[4278]_  = \new_[4277]_  | \new_[4274]_ ;
  assign \new_[4281]_  = \new_[1142]_  | \new_[1143]_ ;
  assign \new_[4284]_  = \new_[1140]_  | \new_[1141]_ ;
  assign \new_[4285]_  = \new_[4284]_  | \new_[4281]_ ;
  assign \new_[4286]_  = \new_[4285]_  | \new_[4278]_ ;
  assign \new_[4289]_  = \new_[1138]_  | \new_[1139]_ ;
  assign \new_[4292]_  = \new_[1136]_  | \new_[1137]_ ;
  assign \new_[4293]_  = \new_[4292]_  | \new_[4289]_ ;
  assign \new_[4296]_  = \new_[1134]_  | \new_[1135]_ ;
  assign \new_[4300]_  = \new_[1131]_  | \new_[1132]_ ;
  assign \new_[4301]_  = \new_[1133]_  | \new_[4300]_ ;
  assign \new_[4302]_  = \new_[4301]_  | \new_[4296]_ ;
  assign \new_[4303]_  = \new_[4302]_  | \new_[4293]_ ;
  assign \new_[4304]_  = \new_[4303]_  | \new_[4286]_ ;
  assign \new_[4305]_  = \new_[4304]_  | \new_[4271]_ ;
  assign \new_[4308]_  = \new_[1129]_  | \new_[1130]_ ;
  assign \new_[4311]_  = \new_[1127]_  | \new_[1128]_ ;
  assign \new_[4312]_  = \new_[4311]_  | \new_[4308]_ ;
  assign \new_[4315]_  = \new_[1125]_  | \new_[1126]_ ;
  assign \new_[4318]_  = \new_[1123]_  | \new_[1124]_ ;
  assign \new_[4319]_  = \new_[4318]_  | \new_[4315]_ ;
  assign \new_[4320]_  = \new_[4319]_  | \new_[4312]_ ;
  assign \new_[4323]_  = \new_[1121]_  | \new_[1122]_ ;
  assign \new_[4326]_  = \new_[1119]_  | \new_[1120]_ ;
  assign \new_[4327]_  = \new_[4326]_  | \new_[4323]_ ;
  assign \new_[4330]_  = \new_[1117]_  | \new_[1118]_ ;
  assign \new_[4334]_  = \new_[1114]_  | \new_[1115]_ ;
  assign \new_[4335]_  = \new_[1116]_  | \new_[4334]_ ;
  assign \new_[4336]_  = \new_[4335]_  | \new_[4330]_ ;
  assign \new_[4337]_  = \new_[4336]_  | \new_[4327]_ ;
  assign \new_[4338]_  = \new_[4337]_  | \new_[4320]_ ;
  assign \new_[4341]_  = \new_[1112]_  | \new_[1113]_ ;
  assign \new_[4344]_  = \new_[1110]_  | \new_[1111]_ ;
  assign \new_[4345]_  = \new_[4344]_  | \new_[4341]_ ;
  assign \new_[4348]_  = \new_[1108]_  | \new_[1109]_ ;
  assign \new_[4352]_  = \new_[1105]_  | \new_[1106]_ ;
  assign \new_[4353]_  = \new_[1107]_  | \new_[4352]_ ;
  assign \new_[4354]_  = \new_[4353]_  | \new_[4348]_ ;
  assign \new_[4355]_  = \new_[4354]_  | \new_[4345]_ ;
  assign \new_[4358]_  = \new_[1103]_  | \new_[1104]_ ;
  assign \new_[4361]_  = \new_[1101]_  | \new_[1102]_ ;
  assign \new_[4362]_  = \new_[4361]_  | \new_[4358]_ ;
  assign \new_[4365]_  = \new_[1099]_  | \new_[1100]_ ;
  assign \new_[4369]_  = \new_[1096]_  | \new_[1097]_ ;
  assign \new_[4370]_  = \new_[1098]_  | \new_[4369]_ ;
  assign \new_[4371]_  = \new_[4370]_  | \new_[4365]_ ;
  assign \new_[4372]_  = \new_[4371]_  | \new_[4362]_ ;
  assign \new_[4373]_  = \new_[4372]_  | \new_[4355]_ ;
  assign \new_[4374]_  = \new_[4373]_  | \new_[4338]_ ;
  assign \new_[4375]_  = \new_[4374]_  | \new_[4305]_ ;
  assign \new_[4376]_  = \new_[4375]_  | \new_[4238]_ ;
  assign \new_[4377]_  = \new_[4376]_  | \new_[4103]_ ;
  assign \new_[4378]_  = \new_[4377]_  | \new_[3830]_ ;
  assign \new_[4379]_  = \new_[4378]_  | \new_[3283]_ ;
  assign \new_[4382]_  = \new_[1094]_  | \new_[1095]_ ;
  assign \new_[4385]_  = \new_[1092]_  | \new_[1093]_ ;
  assign \new_[4386]_  = \new_[4385]_  | \new_[4382]_ ;
  assign \new_[4389]_  = \new_[1090]_  | \new_[1091]_ ;
  assign \new_[4392]_  = \new_[1088]_  | \new_[1089]_ ;
  assign \new_[4393]_  = \new_[4392]_  | \new_[4389]_ ;
  assign \new_[4394]_  = \new_[4393]_  | \new_[4386]_ ;
  assign \new_[4397]_  = \new_[1086]_  | \new_[1087]_ ;
  assign \new_[4400]_  = \new_[1084]_  | \new_[1085]_ ;
  assign \new_[4401]_  = \new_[4400]_  | \new_[4397]_ ;
  assign \new_[4404]_  = \new_[1082]_  | \new_[1083]_ ;
  assign \new_[4408]_  = \new_[1079]_  | \new_[1080]_ ;
  assign \new_[4409]_  = \new_[1081]_  | \new_[4408]_ ;
  assign \new_[4410]_  = \new_[4409]_  | \new_[4404]_ ;
  assign \new_[4411]_  = \new_[4410]_  | \new_[4401]_ ;
  assign \new_[4412]_  = \new_[4411]_  | \new_[4394]_ ;
  assign \new_[4415]_  = \new_[1077]_  | \new_[1078]_ ;
  assign \new_[4418]_  = \new_[1075]_  | \new_[1076]_ ;
  assign \new_[4419]_  = \new_[4418]_  | \new_[4415]_ ;
  assign \new_[4422]_  = \new_[1073]_  | \new_[1074]_ ;
  assign \new_[4425]_  = \new_[1071]_  | \new_[1072]_ ;
  assign \new_[4426]_  = \new_[4425]_  | \new_[4422]_ ;
  assign \new_[4427]_  = \new_[4426]_  | \new_[4419]_ ;
  assign \new_[4430]_  = \new_[1069]_  | \new_[1070]_ ;
  assign \new_[4433]_  = \new_[1067]_  | \new_[1068]_ ;
  assign \new_[4434]_  = \new_[4433]_  | \new_[4430]_ ;
  assign \new_[4437]_  = \new_[1065]_  | \new_[1066]_ ;
  assign \new_[4441]_  = \new_[1062]_  | \new_[1063]_ ;
  assign \new_[4442]_  = \new_[1064]_  | \new_[4441]_ ;
  assign \new_[4443]_  = \new_[4442]_  | \new_[4437]_ ;
  assign \new_[4444]_  = \new_[4443]_  | \new_[4434]_ ;
  assign \new_[4445]_  = \new_[4444]_  | \new_[4427]_ ;
  assign \new_[4446]_  = \new_[4445]_  | \new_[4412]_ ;
  assign \new_[4449]_  = \new_[1060]_  | \new_[1061]_ ;
  assign \new_[4452]_  = \new_[1058]_  | \new_[1059]_ ;
  assign \new_[4453]_  = \new_[4452]_  | \new_[4449]_ ;
  assign \new_[4456]_  = \new_[1056]_  | \new_[1057]_ ;
  assign \new_[4459]_  = \new_[1054]_  | \new_[1055]_ ;
  assign \new_[4460]_  = \new_[4459]_  | \new_[4456]_ ;
  assign \new_[4461]_  = \new_[4460]_  | \new_[4453]_ ;
  assign \new_[4464]_  = \new_[1052]_  | \new_[1053]_ ;
  assign \new_[4467]_  = \new_[1050]_  | \new_[1051]_ ;
  assign \new_[4468]_  = \new_[4467]_  | \new_[4464]_ ;
  assign \new_[4471]_  = \new_[1048]_  | \new_[1049]_ ;
  assign \new_[4475]_  = \new_[1045]_  | \new_[1046]_ ;
  assign \new_[4476]_  = \new_[1047]_  | \new_[4475]_ ;
  assign \new_[4477]_  = \new_[4476]_  | \new_[4471]_ ;
  assign \new_[4478]_  = \new_[4477]_  | \new_[4468]_ ;
  assign \new_[4479]_  = \new_[4478]_  | \new_[4461]_ ;
  assign \new_[4482]_  = \new_[1043]_  | \new_[1044]_ ;
  assign \new_[4485]_  = \new_[1041]_  | \new_[1042]_ ;
  assign \new_[4486]_  = \new_[4485]_  | \new_[4482]_ ;
  assign \new_[4489]_  = \new_[1039]_  | \new_[1040]_ ;
  assign \new_[4492]_  = \new_[1037]_  | \new_[1038]_ ;
  assign \new_[4493]_  = \new_[4492]_  | \new_[4489]_ ;
  assign \new_[4494]_  = \new_[4493]_  | \new_[4486]_ ;
  assign \new_[4497]_  = \new_[1035]_  | \new_[1036]_ ;
  assign \new_[4500]_  = \new_[1033]_  | \new_[1034]_ ;
  assign \new_[4501]_  = \new_[4500]_  | \new_[4497]_ ;
  assign \new_[4504]_  = \new_[1031]_  | \new_[1032]_ ;
  assign \new_[4508]_  = \new_[1028]_  | \new_[1029]_ ;
  assign \new_[4509]_  = \new_[1030]_  | \new_[4508]_ ;
  assign \new_[4510]_  = \new_[4509]_  | \new_[4504]_ ;
  assign \new_[4511]_  = \new_[4510]_  | \new_[4501]_ ;
  assign \new_[4512]_  = \new_[4511]_  | \new_[4494]_ ;
  assign \new_[4513]_  = \new_[4512]_  | \new_[4479]_ ;
  assign \new_[4514]_  = \new_[4513]_  | \new_[4446]_ ;
  assign \new_[4517]_  = \new_[1026]_  | \new_[1027]_ ;
  assign \new_[4520]_  = \new_[1024]_  | \new_[1025]_ ;
  assign \new_[4521]_  = \new_[4520]_  | \new_[4517]_ ;
  assign \new_[4524]_  = \new_[1022]_  | \new_[1023]_ ;
  assign \new_[4527]_  = \new_[1020]_  | \new_[1021]_ ;
  assign \new_[4528]_  = \new_[4527]_  | \new_[4524]_ ;
  assign \new_[4529]_  = \new_[4528]_  | \new_[4521]_ ;
  assign \new_[4532]_  = \new_[1018]_  | \new_[1019]_ ;
  assign \new_[4535]_  = \new_[1016]_  | \new_[1017]_ ;
  assign \new_[4536]_  = \new_[4535]_  | \new_[4532]_ ;
  assign \new_[4539]_  = \new_[1014]_  | \new_[1015]_ ;
  assign \new_[4543]_  = \new_[1011]_  | \new_[1012]_ ;
  assign \new_[4544]_  = \new_[1013]_  | \new_[4543]_ ;
  assign \new_[4545]_  = \new_[4544]_  | \new_[4539]_ ;
  assign \new_[4546]_  = \new_[4545]_  | \new_[4536]_ ;
  assign \new_[4547]_  = \new_[4546]_  | \new_[4529]_ ;
  assign \new_[4550]_  = \new_[1009]_  | \new_[1010]_ ;
  assign \new_[4553]_  = \new_[1007]_  | \new_[1008]_ ;
  assign \new_[4554]_  = \new_[4553]_  | \new_[4550]_ ;
  assign \new_[4557]_  = \new_[1005]_  | \new_[1006]_ ;
  assign \new_[4560]_  = \new_[1003]_  | \new_[1004]_ ;
  assign \new_[4561]_  = \new_[4560]_  | \new_[4557]_ ;
  assign \new_[4562]_  = \new_[4561]_  | \new_[4554]_ ;
  assign \new_[4565]_  = \new_[1001]_  | \new_[1002]_ ;
  assign \new_[4568]_  = \new_[999]_  | \new_[1000]_ ;
  assign \new_[4569]_  = \new_[4568]_  | \new_[4565]_ ;
  assign \new_[4572]_  = \new_[997]_  | \new_[998]_ ;
  assign \new_[4576]_  = \new_[994]_  | \new_[995]_ ;
  assign \new_[4577]_  = \new_[996]_  | \new_[4576]_ ;
  assign \new_[4578]_  = \new_[4577]_  | \new_[4572]_ ;
  assign \new_[4579]_  = \new_[4578]_  | \new_[4569]_ ;
  assign \new_[4580]_  = \new_[4579]_  | \new_[4562]_ ;
  assign \new_[4581]_  = \new_[4580]_  | \new_[4547]_ ;
  assign \new_[4584]_  = \new_[992]_  | \new_[993]_ ;
  assign \new_[4587]_  = \new_[990]_  | \new_[991]_ ;
  assign \new_[4588]_  = \new_[4587]_  | \new_[4584]_ ;
  assign \new_[4591]_  = \new_[988]_  | \new_[989]_ ;
  assign \new_[4594]_  = \new_[986]_  | \new_[987]_ ;
  assign \new_[4595]_  = \new_[4594]_  | \new_[4591]_ ;
  assign \new_[4596]_  = \new_[4595]_  | \new_[4588]_ ;
  assign \new_[4599]_  = \new_[984]_  | \new_[985]_ ;
  assign \new_[4602]_  = \new_[982]_  | \new_[983]_ ;
  assign \new_[4603]_  = \new_[4602]_  | \new_[4599]_ ;
  assign \new_[4606]_  = \new_[980]_  | \new_[981]_ ;
  assign \new_[4610]_  = \new_[977]_  | \new_[978]_ ;
  assign \new_[4611]_  = \new_[979]_  | \new_[4610]_ ;
  assign \new_[4612]_  = \new_[4611]_  | \new_[4606]_ ;
  assign \new_[4613]_  = \new_[4612]_  | \new_[4603]_ ;
  assign \new_[4614]_  = \new_[4613]_  | \new_[4596]_ ;
  assign \new_[4617]_  = \new_[975]_  | \new_[976]_ ;
  assign \new_[4620]_  = \new_[973]_  | \new_[974]_ ;
  assign \new_[4621]_  = \new_[4620]_  | \new_[4617]_ ;
  assign \new_[4624]_  = \new_[971]_  | \new_[972]_ ;
  assign \new_[4627]_  = \new_[969]_  | \new_[970]_ ;
  assign \new_[4628]_  = \new_[4627]_  | \new_[4624]_ ;
  assign \new_[4629]_  = \new_[4628]_  | \new_[4621]_ ;
  assign \new_[4632]_  = \new_[967]_  | \new_[968]_ ;
  assign \new_[4635]_  = \new_[965]_  | \new_[966]_ ;
  assign \new_[4636]_  = \new_[4635]_  | \new_[4632]_ ;
  assign \new_[4639]_  = \new_[963]_  | \new_[964]_ ;
  assign \new_[4643]_  = \new_[960]_  | \new_[961]_ ;
  assign \new_[4644]_  = \new_[962]_  | \new_[4643]_ ;
  assign \new_[4645]_  = \new_[4644]_  | \new_[4639]_ ;
  assign \new_[4646]_  = \new_[4645]_  | \new_[4636]_ ;
  assign \new_[4647]_  = \new_[4646]_  | \new_[4629]_ ;
  assign \new_[4648]_  = \new_[4647]_  | \new_[4614]_ ;
  assign \new_[4649]_  = \new_[4648]_  | \new_[4581]_ ;
  assign \new_[4650]_  = \new_[4649]_  | \new_[4514]_ ;
  assign \new_[4653]_  = \new_[958]_  | \new_[959]_ ;
  assign \new_[4656]_  = \new_[956]_  | \new_[957]_ ;
  assign \new_[4657]_  = \new_[4656]_  | \new_[4653]_ ;
  assign \new_[4660]_  = \new_[954]_  | \new_[955]_ ;
  assign \new_[4663]_  = \new_[952]_  | \new_[953]_ ;
  assign \new_[4664]_  = \new_[4663]_  | \new_[4660]_ ;
  assign \new_[4665]_  = \new_[4664]_  | \new_[4657]_ ;
  assign \new_[4668]_  = \new_[950]_  | \new_[951]_ ;
  assign \new_[4671]_  = \new_[948]_  | \new_[949]_ ;
  assign \new_[4672]_  = \new_[4671]_  | \new_[4668]_ ;
  assign \new_[4675]_  = \new_[946]_  | \new_[947]_ ;
  assign \new_[4679]_  = \new_[943]_  | \new_[944]_ ;
  assign \new_[4680]_  = \new_[945]_  | \new_[4679]_ ;
  assign \new_[4681]_  = \new_[4680]_  | \new_[4675]_ ;
  assign \new_[4682]_  = \new_[4681]_  | \new_[4672]_ ;
  assign \new_[4683]_  = \new_[4682]_  | \new_[4665]_ ;
  assign \new_[4686]_  = \new_[941]_  | \new_[942]_ ;
  assign \new_[4689]_  = \new_[939]_  | \new_[940]_ ;
  assign \new_[4690]_  = \new_[4689]_  | \new_[4686]_ ;
  assign \new_[4693]_  = \new_[937]_  | \new_[938]_ ;
  assign \new_[4696]_  = \new_[935]_  | \new_[936]_ ;
  assign \new_[4697]_  = \new_[4696]_  | \new_[4693]_ ;
  assign \new_[4698]_  = \new_[4697]_  | \new_[4690]_ ;
  assign \new_[4701]_  = \new_[933]_  | \new_[934]_ ;
  assign \new_[4704]_  = \new_[931]_  | \new_[932]_ ;
  assign \new_[4705]_  = \new_[4704]_  | \new_[4701]_ ;
  assign \new_[4708]_  = \new_[929]_  | \new_[930]_ ;
  assign \new_[4712]_  = \new_[926]_  | \new_[927]_ ;
  assign \new_[4713]_  = \new_[928]_  | \new_[4712]_ ;
  assign \new_[4714]_  = \new_[4713]_  | \new_[4708]_ ;
  assign \new_[4715]_  = \new_[4714]_  | \new_[4705]_ ;
  assign \new_[4716]_  = \new_[4715]_  | \new_[4698]_ ;
  assign \new_[4717]_  = \new_[4716]_  | \new_[4683]_ ;
  assign \new_[4720]_  = \new_[924]_  | \new_[925]_ ;
  assign \new_[4723]_  = \new_[922]_  | \new_[923]_ ;
  assign \new_[4724]_  = \new_[4723]_  | \new_[4720]_ ;
  assign \new_[4727]_  = \new_[920]_  | \new_[921]_ ;
  assign \new_[4730]_  = \new_[918]_  | \new_[919]_ ;
  assign \new_[4731]_  = \new_[4730]_  | \new_[4727]_ ;
  assign \new_[4732]_  = \new_[4731]_  | \new_[4724]_ ;
  assign \new_[4735]_  = \new_[916]_  | \new_[917]_ ;
  assign \new_[4738]_  = \new_[914]_  | \new_[915]_ ;
  assign \new_[4739]_  = \new_[4738]_  | \new_[4735]_ ;
  assign \new_[4742]_  = \new_[912]_  | \new_[913]_ ;
  assign \new_[4746]_  = \new_[909]_  | \new_[910]_ ;
  assign \new_[4747]_  = \new_[911]_  | \new_[4746]_ ;
  assign \new_[4748]_  = \new_[4747]_  | \new_[4742]_ ;
  assign \new_[4749]_  = \new_[4748]_  | \new_[4739]_ ;
  assign \new_[4750]_  = \new_[4749]_  | \new_[4732]_ ;
  assign \new_[4753]_  = \new_[907]_  | \new_[908]_ ;
  assign \new_[4756]_  = \new_[905]_  | \new_[906]_ ;
  assign \new_[4757]_  = \new_[4756]_  | \new_[4753]_ ;
  assign \new_[4760]_  = \new_[903]_  | \new_[904]_ ;
  assign \new_[4763]_  = \new_[901]_  | \new_[902]_ ;
  assign \new_[4764]_  = \new_[4763]_  | \new_[4760]_ ;
  assign \new_[4765]_  = \new_[4764]_  | \new_[4757]_ ;
  assign \new_[4768]_  = \new_[899]_  | \new_[900]_ ;
  assign \new_[4771]_  = \new_[897]_  | \new_[898]_ ;
  assign \new_[4772]_  = \new_[4771]_  | \new_[4768]_ ;
  assign \new_[4775]_  = \new_[895]_  | \new_[896]_ ;
  assign \new_[4779]_  = \new_[892]_  | \new_[893]_ ;
  assign \new_[4780]_  = \new_[894]_  | \new_[4779]_ ;
  assign \new_[4781]_  = \new_[4780]_  | \new_[4775]_ ;
  assign \new_[4782]_  = \new_[4781]_  | \new_[4772]_ ;
  assign \new_[4783]_  = \new_[4782]_  | \new_[4765]_ ;
  assign \new_[4784]_  = \new_[4783]_  | \new_[4750]_ ;
  assign \new_[4785]_  = \new_[4784]_  | \new_[4717]_ ;
  assign \new_[4788]_  = \new_[890]_  | \new_[891]_ ;
  assign \new_[4791]_  = \new_[888]_  | \new_[889]_ ;
  assign \new_[4792]_  = \new_[4791]_  | \new_[4788]_ ;
  assign \new_[4795]_  = \new_[886]_  | \new_[887]_ ;
  assign \new_[4798]_  = \new_[884]_  | \new_[885]_ ;
  assign \new_[4799]_  = \new_[4798]_  | \new_[4795]_ ;
  assign \new_[4800]_  = \new_[4799]_  | \new_[4792]_ ;
  assign \new_[4803]_  = \new_[882]_  | \new_[883]_ ;
  assign \new_[4806]_  = \new_[880]_  | \new_[881]_ ;
  assign \new_[4807]_  = \new_[4806]_  | \new_[4803]_ ;
  assign \new_[4810]_  = \new_[878]_  | \new_[879]_ ;
  assign \new_[4814]_  = \new_[875]_  | \new_[876]_ ;
  assign \new_[4815]_  = \new_[877]_  | \new_[4814]_ ;
  assign \new_[4816]_  = \new_[4815]_  | \new_[4810]_ ;
  assign \new_[4817]_  = \new_[4816]_  | \new_[4807]_ ;
  assign \new_[4818]_  = \new_[4817]_  | \new_[4800]_ ;
  assign \new_[4821]_  = \new_[873]_  | \new_[874]_ ;
  assign \new_[4824]_  = \new_[871]_  | \new_[872]_ ;
  assign \new_[4825]_  = \new_[4824]_  | \new_[4821]_ ;
  assign \new_[4828]_  = \new_[869]_  | \new_[870]_ ;
  assign \new_[4831]_  = \new_[867]_  | \new_[868]_ ;
  assign \new_[4832]_  = \new_[4831]_  | \new_[4828]_ ;
  assign \new_[4833]_  = \new_[4832]_  | \new_[4825]_ ;
  assign \new_[4836]_  = \new_[865]_  | \new_[866]_ ;
  assign \new_[4839]_  = \new_[863]_  | \new_[864]_ ;
  assign \new_[4840]_  = \new_[4839]_  | \new_[4836]_ ;
  assign \new_[4843]_  = \new_[861]_  | \new_[862]_ ;
  assign \new_[4847]_  = \new_[858]_  | \new_[859]_ ;
  assign \new_[4848]_  = \new_[860]_  | \new_[4847]_ ;
  assign \new_[4849]_  = \new_[4848]_  | \new_[4843]_ ;
  assign \new_[4850]_  = \new_[4849]_  | \new_[4840]_ ;
  assign \new_[4851]_  = \new_[4850]_  | \new_[4833]_ ;
  assign \new_[4852]_  = \new_[4851]_  | \new_[4818]_ ;
  assign \new_[4855]_  = \new_[856]_  | \new_[857]_ ;
  assign \new_[4858]_  = \new_[854]_  | \new_[855]_ ;
  assign \new_[4859]_  = \new_[4858]_  | \new_[4855]_ ;
  assign \new_[4862]_  = \new_[852]_  | \new_[853]_ ;
  assign \new_[4865]_  = \new_[850]_  | \new_[851]_ ;
  assign \new_[4866]_  = \new_[4865]_  | \new_[4862]_ ;
  assign \new_[4867]_  = \new_[4866]_  | \new_[4859]_ ;
  assign \new_[4870]_  = \new_[848]_  | \new_[849]_ ;
  assign \new_[4873]_  = \new_[846]_  | \new_[847]_ ;
  assign \new_[4874]_  = \new_[4873]_  | \new_[4870]_ ;
  assign \new_[4877]_  = \new_[844]_  | \new_[845]_ ;
  assign \new_[4881]_  = \new_[841]_  | \new_[842]_ ;
  assign \new_[4882]_  = \new_[843]_  | \new_[4881]_ ;
  assign \new_[4883]_  = \new_[4882]_  | \new_[4877]_ ;
  assign \new_[4884]_  = \new_[4883]_  | \new_[4874]_ ;
  assign \new_[4885]_  = \new_[4884]_  | \new_[4867]_ ;
  assign \new_[4888]_  = \new_[839]_  | \new_[840]_ ;
  assign \new_[4891]_  = \new_[837]_  | \new_[838]_ ;
  assign \new_[4892]_  = \new_[4891]_  | \new_[4888]_ ;
  assign \new_[4895]_  = \new_[835]_  | \new_[836]_ ;
  assign \new_[4899]_  = \new_[832]_  | \new_[833]_ ;
  assign \new_[4900]_  = \new_[834]_  | \new_[4899]_ ;
  assign \new_[4901]_  = \new_[4900]_  | \new_[4895]_ ;
  assign \new_[4902]_  = \new_[4901]_  | \new_[4892]_ ;
  assign \new_[4905]_  = \new_[830]_  | \new_[831]_ ;
  assign \new_[4908]_  = \new_[828]_  | \new_[829]_ ;
  assign \new_[4909]_  = \new_[4908]_  | \new_[4905]_ ;
  assign \new_[4912]_  = \new_[826]_  | \new_[827]_ ;
  assign \new_[4916]_  = \new_[823]_  | \new_[824]_ ;
  assign \new_[4917]_  = \new_[825]_  | \new_[4916]_ ;
  assign \new_[4918]_  = \new_[4917]_  | \new_[4912]_ ;
  assign \new_[4919]_  = \new_[4918]_  | \new_[4909]_ ;
  assign \new_[4920]_  = \new_[4919]_  | \new_[4902]_ ;
  assign \new_[4921]_  = \new_[4920]_  | \new_[4885]_ ;
  assign \new_[4922]_  = \new_[4921]_  | \new_[4852]_ ;
  assign \new_[4923]_  = \new_[4922]_  | \new_[4785]_ ;
  assign \new_[4924]_  = \new_[4923]_  | \new_[4650]_ ;
  assign \new_[4927]_  = \new_[821]_  | \new_[822]_ ;
  assign \new_[4930]_  = \new_[819]_  | \new_[820]_ ;
  assign \new_[4931]_  = \new_[4930]_  | \new_[4927]_ ;
  assign \new_[4934]_  = \new_[817]_  | \new_[818]_ ;
  assign \new_[4937]_  = \new_[815]_  | \new_[816]_ ;
  assign \new_[4938]_  = \new_[4937]_  | \new_[4934]_ ;
  assign \new_[4939]_  = \new_[4938]_  | \new_[4931]_ ;
  assign \new_[4942]_  = \new_[813]_  | \new_[814]_ ;
  assign \new_[4945]_  = \new_[811]_  | \new_[812]_ ;
  assign \new_[4946]_  = \new_[4945]_  | \new_[4942]_ ;
  assign \new_[4949]_  = \new_[809]_  | \new_[810]_ ;
  assign \new_[4953]_  = \new_[806]_  | \new_[807]_ ;
  assign \new_[4954]_  = \new_[808]_  | \new_[4953]_ ;
  assign \new_[4955]_  = \new_[4954]_  | \new_[4949]_ ;
  assign \new_[4956]_  = \new_[4955]_  | \new_[4946]_ ;
  assign \new_[4957]_  = \new_[4956]_  | \new_[4939]_ ;
  assign \new_[4960]_  = \new_[804]_  | \new_[805]_ ;
  assign \new_[4963]_  = \new_[802]_  | \new_[803]_ ;
  assign \new_[4964]_  = \new_[4963]_  | \new_[4960]_ ;
  assign \new_[4967]_  = \new_[800]_  | \new_[801]_ ;
  assign \new_[4970]_  = \new_[798]_  | \new_[799]_ ;
  assign \new_[4971]_  = \new_[4970]_  | \new_[4967]_ ;
  assign \new_[4972]_  = \new_[4971]_  | \new_[4964]_ ;
  assign \new_[4975]_  = \new_[796]_  | \new_[797]_ ;
  assign \new_[4978]_  = \new_[794]_  | \new_[795]_ ;
  assign \new_[4979]_  = \new_[4978]_  | \new_[4975]_ ;
  assign \new_[4982]_  = \new_[792]_  | \new_[793]_ ;
  assign \new_[4986]_  = \new_[789]_  | \new_[790]_ ;
  assign \new_[4987]_  = \new_[791]_  | \new_[4986]_ ;
  assign \new_[4988]_  = \new_[4987]_  | \new_[4982]_ ;
  assign \new_[4989]_  = \new_[4988]_  | \new_[4979]_ ;
  assign \new_[4990]_  = \new_[4989]_  | \new_[4972]_ ;
  assign \new_[4991]_  = \new_[4990]_  | \new_[4957]_ ;
  assign \new_[4994]_  = \new_[787]_  | \new_[788]_ ;
  assign \new_[4997]_  = \new_[785]_  | \new_[786]_ ;
  assign \new_[4998]_  = \new_[4997]_  | \new_[4994]_ ;
  assign \new_[5001]_  = \new_[783]_  | \new_[784]_ ;
  assign \new_[5004]_  = \new_[781]_  | \new_[782]_ ;
  assign \new_[5005]_  = \new_[5004]_  | \new_[5001]_ ;
  assign \new_[5006]_  = \new_[5005]_  | \new_[4998]_ ;
  assign \new_[5009]_  = \new_[779]_  | \new_[780]_ ;
  assign \new_[5012]_  = \new_[777]_  | \new_[778]_ ;
  assign \new_[5013]_  = \new_[5012]_  | \new_[5009]_ ;
  assign \new_[5016]_  = \new_[775]_  | \new_[776]_ ;
  assign \new_[5020]_  = \new_[772]_  | \new_[773]_ ;
  assign \new_[5021]_  = \new_[774]_  | \new_[5020]_ ;
  assign \new_[5022]_  = \new_[5021]_  | \new_[5016]_ ;
  assign \new_[5023]_  = \new_[5022]_  | \new_[5013]_ ;
  assign \new_[5024]_  = \new_[5023]_  | \new_[5006]_ ;
  assign \new_[5027]_  = \new_[770]_  | \new_[771]_ ;
  assign \new_[5030]_  = \new_[768]_  | \new_[769]_ ;
  assign \new_[5031]_  = \new_[5030]_  | \new_[5027]_ ;
  assign \new_[5034]_  = \new_[766]_  | \new_[767]_ ;
  assign \new_[5037]_  = \new_[764]_  | \new_[765]_ ;
  assign \new_[5038]_  = \new_[5037]_  | \new_[5034]_ ;
  assign \new_[5039]_  = \new_[5038]_  | \new_[5031]_ ;
  assign \new_[5042]_  = \new_[762]_  | \new_[763]_ ;
  assign \new_[5045]_  = \new_[760]_  | \new_[761]_ ;
  assign \new_[5046]_  = \new_[5045]_  | \new_[5042]_ ;
  assign \new_[5049]_  = \new_[758]_  | \new_[759]_ ;
  assign \new_[5053]_  = \new_[755]_  | \new_[756]_ ;
  assign \new_[5054]_  = \new_[757]_  | \new_[5053]_ ;
  assign \new_[5055]_  = \new_[5054]_  | \new_[5049]_ ;
  assign \new_[5056]_  = \new_[5055]_  | \new_[5046]_ ;
  assign \new_[5057]_  = \new_[5056]_  | \new_[5039]_ ;
  assign \new_[5058]_  = \new_[5057]_  | \new_[5024]_ ;
  assign \new_[5059]_  = \new_[5058]_  | \new_[4991]_ ;
  assign \new_[5062]_  = \new_[753]_  | \new_[754]_ ;
  assign \new_[5065]_  = \new_[751]_  | \new_[752]_ ;
  assign \new_[5066]_  = \new_[5065]_  | \new_[5062]_ ;
  assign \new_[5069]_  = \new_[749]_  | \new_[750]_ ;
  assign \new_[5072]_  = \new_[747]_  | \new_[748]_ ;
  assign \new_[5073]_  = \new_[5072]_  | \new_[5069]_ ;
  assign \new_[5074]_  = \new_[5073]_  | \new_[5066]_ ;
  assign \new_[5077]_  = \new_[745]_  | \new_[746]_ ;
  assign \new_[5080]_  = \new_[743]_  | \new_[744]_ ;
  assign \new_[5081]_  = \new_[5080]_  | \new_[5077]_ ;
  assign \new_[5084]_  = \new_[741]_  | \new_[742]_ ;
  assign \new_[5088]_  = \new_[738]_  | \new_[739]_ ;
  assign \new_[5089]_  = \new_[740]_  | \new_[5088]_ ;
  assign \new_[5090]_  = \new_[5089]_  | \new_[5084]_ ;
  assign \new_[5091]_  = \new_[5090]_  | \new_[5081]_ ;
  assign \new_[5092]_  = \new_[5091]_  | \new_[5074]_ ;
  assign \new_[5095]_  = \new_[736]_  | \new_[737]_ ;
  assign \new_[5098]_  = \new_[734]_  | \new_[735]_ ;
  assign \new_[5099]_  = \new_[5098]_  | \new_[5095]_ ;
  assign \new_[5102]_  = \new_[732]_  | \new_[733]_ ;
  assign \new_[5105]_  = \new_[730]_  | \new_[731]_ ;
  assign \new_[5106]_  = \new_[5105]_  | \new_[5102]_ ;
  assign \new_[5107]_  = \new_[5106]_  | \new_[5099]_ ;
  assign \new_[5110]_  = \new_[728]_  | \new_[729]_ ;
  assign \new_[5113]_  = \new_[726]_  | \new_[727]_ ;
  assign \new_[5114]_  = \new_[5113]_  | \new_[5110]_ ;
  assign \new_[5117]_  = \new_[724]_  | \new_[725]_ ;
  assign \new_[5121]_  = \new_[721]_  | \new_[722]_ ;
  assign \new_[5122]_  = \new_[723]_  | \new_[5121]_ ;
  assign \new_[5123]_  = \new_[5122]_  | \new_[5117]_ ;
  assign \new_[5124]_  = \new_[5123]_  | \new_[5114]_ ;
  assign \new_[5125]_  = \new_[5124]_  | \new_[5107]_ ;
  assign \new_[5126]_  = \new_[5125]_  | \new_[5092]_ ;
  assign \new_[5129]_  = \new_[719]_  | \new_[720]_ ;
  assign \new_[5132]_  = \new_[717]_  | \new_[718]_ ;
  assign \new_[5133]_  = \new_[5132]_  | \new_[5129]_ ;
  assign \new_[5136]_  = \new_[715]_  | \new_[716]_ ;
  assign \new_[5139]_  = \new_[713]_  | \new_[714]_ ;
  assign \new_[5140]_  = \new_[5139]_  | \new_[5136]_ ;
  assign \new_[5141]_  = \new_[5140]_  | \new_[5133]_ ;
  assign \new_[5144]_  = \new_[711]_  | \new_[712]_ ;
  assign \new_[5147]_  = \new_[709]_  | \new_[710]_ ;
  assign \new_[5148]_  = \new_[5147]_  | \new_[5144]_ ;
  assign \new_[5151]_  = \new_[707]_  | \new_[708]_ ;
  assign \new_[5155]_  = \new_[704]_  | \new_[705]_ ;
  assign \new_[5156]_  = \new_[706]_  | \new_[5155]_ ;
  assign \new_[5157]_  = \new_[5156]_  | \new_[5151]_ ;
  assign \new_[5158]_  = \new_[5157]_  | \new_[5148]_ ;
  assign \new_[5159]_  = \new_[5158]_  | \new_[5141]_ ;
  assign \new_[5162]_  = \new_[702]_  | \new_[703]_ ;
  assign \new_[5165]_  = \new_[700]_  | \new_[701]_ ;
  assign \new_[5166]_  = \new_[5165]_  | \new_[5162]_ ;
  assign \new_[5169]_  = \new_[698]_  | \new_[699]_ ;
  assign \new_[5173]_  = \new_[695]_  | \new_[696]_ ;
  assign \new_[5174]_  = \new_[697]_  | \new_[5173]_ ;
  assign \new_[5175]_  = \new_[5174]_  | \new_[5169]_ ;
  assign \new_[5176]_  = \new_[5175]_  | \new_[5166]_ ;
  assign \new_[5179]_  = \new_[693]_  | \new_[694]_ ;
  assign \new_[5182]_  = \new_[691]_  | \new_[692]_ ;
  assign \new_[5183]_  = \new_[5182]_  | \new_[5179]_ ;
  assign \new_[5186]_  = \new_[689]_  | \new_[690]_ ;
  assign \new_[5190]_  = \new_[686]_  | \new_[687]_ ;
  assign \new_[5191]_  = \new_[688]_  | \new_[5190]_ ;
  assign \new_[5192]_  = \new_[5191]_  | \new_[5186]_ ;
  assign \new_[5193]_  = \new_[5192]_  | \new_[5183]_ ;
  assign \new_[5194]_  = \new_[5193]_  | \new_[5176]_ ;
  assign \new_[5195]_  = \new_[5194]_  | \new_[5159]_ ;
  assign \new_[5196]_  = \new_[5195]_  | \new_[5126]_ ;
  assign \new_[5197]_  = \new_[5196]_  | \new_[5059]_ ;
  assign \new_[5200]_  = \new_[684]_  | \new_[685]_ ;
  assign \new_[5203]_  = \new_[682]_  | \new_[683]_ ;
  assign \new_[5204]_  = \new_[5203]_  | \new_[5200]_ ;
  assign \new_[5207]_  = \new_[680]_  | \new_[681]_ ;
  assign \new_[5210]_  = \new_[678]_  | \new_[679]_ ;
  assign \new_[5211]_  = \new_[5210]_  | \new_[5207]_ ;
  assign \new_[5212]_  = \new_[5211]_  | \new_[5204]_ ;
  assign \new_[5215]_  = \new_[676]_  | \new_[677]_ ;
  assign \new_[5218]_  = \new_[674]_  | \new_[675]_ ;
  assign \new_[5219]_  = \new_[5218]_  | \new_[5215]_ ;
  assign \new_[5222]_  = \new_[672]_  | \new_[673]_ ;
  assign \new_[5226]_  = \new_[669]_  | \new_[670]_ ;
  assign \new_[5227]_  = \new_[671]_  | \new_[5226]_ ;
  assign \new_[5228]_  = \new_[5227]_  | \new_[5222]_ ;
  assign \new_[5229]_  = \new_[5228]_  | \new_[5219]_ ;
  assign \new_[5230]_  = \new_[5229]_  | \new_[5212]_ ;
  assign \new_[5233]_  = \new_[667]_  | \new_[668]_ ;
  assign \new_[5236]_  = \new_[665]_  | \new_[666]_ ;
  assign \new_[5237]_  = \new_[5236]_  | \new_[5233]_ ;
  assign \new_[5240]_  = \new_[663]_  | \new_[664]_ ;
  assign \new_[5243]_  = \new_[661]_  | \new_[662]_ ;
  assign \new_[5244]_  = \new_[5243]_  | \new_[5240]_ ;
  assign \new_[5245]_  = \new_[5244]_  | \new_[5237]_ ;
  assign \new_[5248]_  = \new_[659]_  | \new_[660]_ ;
  assign \new_[5251]_  = \new_[657]_  | \new_[658]_ ;
  assign \new_[5252]_  = \new_[5251]_  | \new_[5248]_ ;
  assign \new_[5255]_  = \new_[655]_  | \new_[656]_ ;
  assign \new_[5259]_  = \new_[652]_  | \new_[653]_ ;
  assign \new_[5260]_  = \new_[654]_  | \new_[5259]_ ;
  assign \new_[5261]_  = \new_[5260]_  | \new_[5255]_ ;
  assign \new_[5262]_  = \new_[5261]_  | \new_[5252]_ ;
  assign \new_[5263]_  = \new_[5262]_  | \new_[5245]_ ;
  assign \new_[5264]_  = \new_[5263]_  | \new_[5230]_ ;
  assign \new_[5267]_  = \new_[650]_  | \new_[651]_ ;
  assign \new_[5270]_  = \new_[648]_  | \new_[649]_ ;
  assign \new_[5271]_  = \new_[5270]_  | \new_[5267]_ ;
  assign \new_[5274]_  = \new_[646]_  | \new_[647]_ ;
  assign \new_[5277]_  = \new_[644]_  | \new_[645]_ ;
  assign \new_[5278]_  = \new_[5277]_  | \new_[5274]_ ;
  assign \new_[5279]_  = \new_[5278]_  | \new_[5271]_ ;
  assign \new_[5282]_  = \new_[642]_  | \new_[643]_ ;
  assign \new_[5285]_  = \new_[640]_  | \new_[641]_ ;
  assign \new_[5286]_  = \new_[5285]_  | \new_[5282]_ ;
  assign \new_[5289]_  = \new_[638]_  | \new_[639]_ ;
  assign \new_[5293]_  = \new_[635]_  | \new_[636]_ ;
  assign \new_[5294]_  = \new_[637]_  | \new_[5293]_ ;
  assign \new_[5295]_  = \new_[5294]_  | \new_[5289]_ ;
  assign \new_[5296]_  = \new_[5295]_  | \new_[5286]_ ;
  assign \new_[5297]_  = \new_[5296]_  | \new_[5279]_ ;
  assign \new_[5300]_  = \new_[633]_  | \new_[634]_ ;
  assign \new_[5303]_  = \new_[631]_  | \new_[632]_ ;
  assign \new_[5304]_  = \new_[5303]_  | \new_[5300]_ ;
  assign \new_[5307]_  = \new_[629]_  | \new_[630]_ ;
  assign \new_[5310]_  = \new_[627]_  | \new_[628]_ ;
  assign \new_[5311]_  = \new_[5310]_  | \new_[5307]_ ;
  assign \new_[5312]_  = \new_[5311]_  | \new_[5304]_ ;
  assign \new_[5315]_  = \new_[625]_  | \new_[626]_ ;
  assign \new_[5318]_  = \new_[623]_  | \new_[624]_ ;
  assign \new_[5319]_  = \new_[5318]_  | \new_[5315]_ ;
  assign \new_[5322]_  = \new_[621]_  | \new_[622]_ ;
  assign \new_[5326]_  = \new_[618]_  | \new_[619]_ ;
  assign \new_[5327]_  = \new_[620]_  | \new_[5326]_ ;
  assign \new_[5328]_  = \new_[5327]_  | \new_[5322]_ ;
  assign \new_[5329]_  = \new_[5328]_  | \new_[5319]_ ;
  assign \new_[5330]_  = \new_[5329]_  | \new_[5312]_ ;
  assign \new_[5331]_  = \new_[5330]_  | \new_[5297]_ ;
  assign \new_[5332]_  = \new_[5331]_  | \new_[5264]_ ;
  assign \new_[5335]_  = \new_[616]_  | \new_[617]_ ;
  assign \new_[5338]_  = \new_[614]_  | \new_[615]_ ;
  assign \new_[5339]_  = \new_[5338]_  | \new_[5335]_ ;
  assign \new_[5342]_  = \new_[612]_  | \new_[613]_ ;
  assign \new_[5345]_  = \new_[610]_  | \new_[611]_ ;
  assign \new_[5346]_  = \new_[5345]_  | \new_[5342]_ ;
  assign \new_[5347]_  = \new_[5346]_  | \new_[5339]_ ;
  assign \new_[5350]_  = \new_[608]_  | \new_[609]_ ;
  assign \new_[5353]_  = \new_[606]_  | \new_[607]_ ;
  assign \new_[5354]_  = \new_[5353]_  | \new_[5350]_ ;
  assign \new_[5357]_  = \new_[604]_  | \new_[605]_ ;
  assign \new_[5361]_  = \new_[601]_  | \new_[602]_ ;
  assign \new_[5362]_  = \new_[603]_  | \new_[5361]_ ;
  assign \new_[5363]_  = \new_[5362]_  | \new_[5357]_ ;
  assign \new_[5364]_  = \new_[5363]_  | \new_[5354]_ ;
  assign \new_[5365]_  = \new_[5364]_  | \new_[5347]_ ;
  assign \new_[5368]_  = \new_[599]_  | \new_[600]_ ;
  assign \new_[5371]_  = \new_[597]_  | \new_[598]_ ;
  assign \new_[5372]_  = \new_[5371]_  | \new_[5368]_ ;
  assign \new_[5375]_  = \new_[595]_  | \new_[596]_ ;
  assign \new_[5378]_  = \new_[593]_  | \new_[594]_ ;
  assign \new_[5379]_  = \new_[5378]_  | \new_[5375]_ ;
  assign \new_[5380]_  = \new_[5379]_  | \new_[5372]_ ;
  assign \new_[5383]_  = \new_[591]_  | \new_[592]_ ;
  assign \new_[5386]_  = \new_[589]_  | \new_[590]_ ;
  assign \new_[5387]_  = \new_[5386]_  | \new_[5383]_ ;
  assign \new_[5390]_  = \new_[587]_  | \new_[588]_ ;
  assign \new_[5394]_  = \new_[584]_  | \new_[585]_ ;
  assign \new_[5395]_  = \new_[586]_  | \new_[5394]_ ;
  assign \new_[5396]_  = \new_[5395]_  | \new_[5390]_ ;
  assign \new_[5397]_  = \new_[5396]_  | \new_[5387]_ ;
  assign \new_[5398]_  = \new_[5397]_  | \new_[5380]_ ;
  assign \new_[5399]_  = \new_[5398]_  | \new_[5365]_ ;
  assign \new_[5402]_  = \new_[582]_  | \new_[583]_ ;
  assign \new_[5405]_  = \new_[580]_  | \new_[581]_ ;
  assign \new_[5406]_  = \new_[5405]_  | \new_[5402]_ ;
  assign \new_[5409]_  = \new_[578]_  | \new_[579]_ ;
  assign \new_[5412]_  = \new_[576]_  | \new_[577]_ ;
  assign \new_[5413]_  = \new_[5412]_  | \new_[5409]_ ;
  assign \new_[5414]_  = \new_[5413]_  | \new_[5406]_ ;
  assign \new_[5417]_  = \new_[574]_  | \new_[575]_ ;
  assign \new_[5420]_  = \new_[572]_  | \new_[573]_ ;
  assign \new_[5421]_  = \new_[5420]_  | \new_[5417]_ ;
  assign \new_[5424]_  = \new_[570]_  | \new_[571]_ ;
  assign \new_[5428]_  = \new_[567]_  | \new_[568]_ ;
  assign \new_[5429]_  = \new_[569]_  | \new_[5428]_ ;
  assign \new_[5430]_  = \new_[5429]_  | \new_[5424]_ ;
  assign \new_[5431]_  = \new_[5430]_  | \new_[5421]_ ;
  assign \new_[5432]_  = \new_[5431]_  | \new_[5414]_ ;
  assign \new_[5435]_  = \new_[565]_  | \new_[566]_ ;
  assign \new_[5438]_  = \new_[563]_  | \new_[564]_ ;
  assign \new_[5439]_  = \new_[5438]_  | \new_[5435]_ ;
  assign \new_[5442]_  = \new_[561]_  | \new_[562]_ ;
  assign \new_[5446]_  = \new_[558]_  | \new_[559]_ ;
  assign \new_[5447]_  = \new_[560]_  | \new_[5446]_ ;
  assign \new_[5448]_  = \new_[5447]_  | \new_[5442]_ ;
  assign \new_[5449]_  = \new_[5448]_  | \new_[5439]_ ;
  assign \new_[5452]_  = \new_[556]_  | \new_[557]_ ;
  assign \new_[5455]_  = \new_[554]_  | \new_[555]_ ;
  assign \new_[5456]_  = \new_[5455]_  | \new_[5452]_ ;
  assign \new_[5459]_  = \new_[552]_  | \new_[553]_ ;
  assign \new_[5463]_  = \new_[549]_  | \new_[550]_ ;
  assign \new_[5464]_  = \new_[551]_  | \new_[5463]_ ;
  assign \new_[5465]_  = \new_[5464]_  | \new_[5459]_ ;
  assign \new_[5466]_  = \new_[5465]_  | \new_[5456]_ ;
  assign \new_[5467]_  = \new_[5466]_  | \new_[5449]_ ;
  assign \new_[5468]_  = \new_[5467]_  | \new_[5432]_ ;
  assign \new_[5469]_  = \new_[5468]_  | \new_[5399]_ ;
  assign \new_[5470]_  = \new_[5469]_  | \new_[5332]_ ;
  assign \new_[5471]_  = \new_[5470]_  | \new_[5197]_ ;
  assign \new_[5472]_  = \new_[5471]_  | \new_[4924]_ ;
  assign \new_[5475]_  = \new_[547]_  | \new_[548]_ ;
  assign \new_[5478]_  = \new_[545]_  | \new_[546]_ ;
  assign \new_[5479]_  = \new_[5478]_  | \new_[5475]_ ;
  assign \new_[5482]_  = \new_[543]_  | \new_[544]_ ;
  assign \new_[5485]_  = \new_[541]_  | \new_[542]_ ;
  assign \new_[5486]_  = \new_[5485]_  | \new_[5482]_ ;
  assign \new_[5487]_  = \new_[5486]_  | \new_[5479]_ ;
  assign \new_[5490]_  = \new_[539]_  | \new_[540]_ ;
  assign \new_[5493]_  = \new_[537]_  | \new_[538]_ ;
  assign \new_[5494]_  = \new_[5493]_  | \new_[5490]_ ;
  assign \new_[5497]_  = \new_[535]_  | \new_[536]_ ;
  assign \new_[5501]_  = \new_[532]_  | \new_[533]_ ;
  assign \new_[5502]_  = \new_[534]_  | \new_[5501]_ ;
  assign \new_[5503]_  = \new_[5502]_  | \new_[5497]_ ;
  assign \new_[5504]_  = \new_[5503]_  | \new_[5494]_ ;
  assign \new_[5505]_  = \new_[5504]_  | \new_[5487]_ ;
  assign \new_[5508]_  = \new_[530]_  | \new_[531]_ ;
  assign \new_[5511]_  = \new_[528]_  | \new_[529]_ ;
  assign \new_[5512]_  = \new_[5511]_  | \new_[5508]_ ;
  assign \new_[5515]_  = \new_[526]_  | \new_[527]_ ;
  assign \new_[5518]_  = \new_[524]_  | \new_[525]_ ;
  assign \new_[5519]_  = \new_[5518]_  | \new_[5515]_ ;
  assign \new_[5520]_  = \new_[5519]_  | \new_[5512]_ ;
  assign \new_[5523]_  = \new_[522]_  | \new_[523]_ ;
  assign \new_[5526]_  = \new_[520]_  | \new_[521]_ ;
  assign \new_[5527]_  = \new_[5526]_  | \new_[5523]_ ;
  assign \new_[5530]_  = \new_[518]_  | \new_[519]_ ;
  assign \new_[5534]_  = \new_[515]_  | \new_[516]_ ;
  assign \new_[5535]_  = \new_[517]_  | \new_[5534]_ ;
  assign \new_[5536]_  = \new_[5535]_  | \new_[5530]_ ;
  assign \new_[5537]_  = \new_[5536]_  | \new_[5527]_ ;
  assign \new_[5538]_  = \new_[5537]_  | \new_[5520]_ ;
  assign \new_[5539]_  = \new_[5538]_  | \new_[5505]_ ;
  assign \new_[5542]_  = \new_[513]_  | \new_[514]_ ;
  assign \new_[5545]_  = \new_[511]_  | \new_[512]_ ;
  assign \new_[5546]_  = \new_[5545]_  | \new_[5542]_ ;
  assign \new_[5549]_  = \new_[509]_  | \new_[510]_ ;
  assign \new_[5552]_  = \new_[507]_  | \new_[508]_ ;
  assign \new_[5553]_  = \new_[5552]_  | \new_[5549]_ ;
  assign \new_[5554]_  = \new_[5553]_  | \new_[5546]_ ;
  assign \new_[5557]_  = \new_[505]_  | \new_[506]_ ;
  assign \new_[5560]_  = \new_[503]_  | \new_[504]_ ;
  assign \new_[5561]_  = \new_[5560]_  | \new_[5557]_ ;
  assign \new_[5564]_  = \new_[501]_  | \new_[502]_ ;
  assign \new_[5568]_  = \new_[498]_  | \new_[499]_ ;
  assign \new_[5569]_  = \new_[500]_  | \new_[5568]_ ;
  assign \new_[5570]_  = \new_[5569]_  | \new_[5564]_ ;
  assign \new_[5571]_  = \new_[5570]_  | \new_[5561]_ ;
  assign \new_[5572]_  = \new_[5571]_  | \new_[5554]_ ;
  assign \new_[5575]_  = \new_[496]_  | \new_[497]_ ;
  assign \new_[5578]_  = \new_[494]_  | \new_[495]_ ;
  assign \new_[5579]_  = \new_[5578]_  | \new_[5575]_ ;
  assign \new_[5582]_  = \new_[492]_  | \new_[493]_ ;
  assign \new_[5585]_  = \new_[490]_  | \new_[491]_ ;
  assign \new_[5586]_  = \new_[5585]_  | \new_[5582]_ ;
  assign \new_[5587]_  = \new_[5586]_  | \new_[5579]_ ;
  assign \new_[5590]_  = \new_[488]_  | \new_[489]_ ;
  assign \new_[5593]_  = \new_[486]_  | \new_[487]_ ;
  assign \new_[5594]_  = \new_[5593]_  | \new_[5590]_ ;
  assign \new_[5597]_  = \new_[484]_  | \new_[485]_ ;
  assign \new_[5601]_  = \new_[481]_  | \new_[482]_ ;
  assign \new_[5602]_  = \new_[483]_  | \new_[5601]_ ;
  assign \new_[5603]_  = \new_[5602]_  | \new_[5597]_ ;
  assign \new_[5604]_  = \new_[5603]_  | \new_[5594]_ ;
  assign \new_[5605]_  = \new_[5604]_  | \new_[5587]_ ;
  assign \new_[5606]_  = \new_[5605]_  | \new_[5572]_ ;
  assign \new_[5607]_  = \new_[5606]_  | \new_[5539]_ ;
  assign \new_[5610]_  = \new_[479]_  | \new_[480]_ ;
  assign \new_[5613]_  = \new_[477]_  | \new_[478]_ ;
  assign \new_[5614]_  = \new_[5613]_  | \new_[5610]_ ;
  assign \new_[5617]_  = \new_[475]_  | \new_[476]_ ;
  assign \new_[5620]_  = \new_[473]_  | \new_[474]_ ;
  assign \new_[5621]_  = \new_[5620]_  | \new_[5617]_ ;
  assign \new_[5622]_  = \new_[5621]_  | \new_[5614]_ ;
  assign \new_[5625]_  = \new_[471]_  | \new_[472]_ ;
  assign \new_[5628]_  = \new_[469]_  | \new_[470]_ ;
  assign \new_[5629]_  = \new_[5628]_  | \new_[5625]_ ;
  assign \new_[5632]_  = \new_[467]_  | \new_[468]_ ;
  assign \new_[5636]_  = \new_[464]_  | \new_[465]_ ;
  assign \new_[5637]_  = \new_[466]_  | \new_[5636]_ ;
  assign \new_[5638]_  = \new_[5637]_  | \new_[5632]_ ;
  assign \new_[5639]_  = \new_[5638]_  | \new_[5629]_ ;
  assign \new_[5640]_  = \new_[5639]_  | \new_[5622]_ ;
  assign \new_[5643]_  = \new_[462]_  | \new_[463]_ ;
  assign \new_[5646]_  = \new_[460]_  | \new_[461]_ ;
  assign \new_[5647]_  = \new_[5646]_  | \new_[5643]_ ;
  assign \new_[5650]_  = \new_[458]_  | \new_[459]_ ;
  assign \new_[5653]_  = \new_[456]_  | \new_[457]_ ;
  assign \new_[5654]_  = \new_[5653]_  | \new_[5650]_ ;
  assign \new_[5655]_  = \new_[5654]_  | \new_[5647]_ ;
  assign \new_[5658]_  = \new_[454]_  | \new_[455]_ ;
  assign \new_[5661]_  = \new_[452]_  | \new_[453]_ ;
  assign \new_[5662]_  = \new_[5661]_  | \new_[5658]_ ;
  assign \new_[5665]_  = \new_[450]_  | \new_[451]_ ;
  assign \new_[5669]_  = \new_[447]_  | \new_[448]_ ;
  assign \new_[5670]_  = \new_[449]_  | \new_[5669]_ ;
  assign \new_[5671]_  = \new_[5670]_  | \new_[5665]_ ;
  assign \new_[5672]_  = \new_[5671]_  | \new_[5662]_ ;
  assign \new_[5673]_  = \new_[5672]_  | \new_[5655]_ ;
  assign \new_[5674]_  = \new_[5673]_  | \new_[5640]_ ;
  assign \new_[5677]_  = \new_[445]_  | \new_[446]_ ;
  assign \new_[5680]_  = \new_[443]_  | \new_[444]_ ;
  assign \new_[5681]_  = \new_[5680]_  | \new_[5677]_ ;
  assign \new_[5684]_  = \new_[441]_  | \new_[442]_ ;
  assign \new_[5687]_  = \new_[439]_  | \new_[440]_ ;
  assign \new_[5688]_  = \new_[5687]_  | \new_[5684]_ ;
  assign \new_[5689]_  = \new_[5688]_  | \new_[5681]_ ;
  assign \new_[5692]_  = \new_[437]_  | \new_[438]_ ;
  assign \new_[5695]_  = \new_[435]_  | \new_[436]_ ;
  assign \new_[5696]_  = \new_[5695]_  | \new_[5692]_ ;
  assign \new_[5699]_  = \new_[433]_  | \new_[434]_ ;
  assign \new_[5703]_  = \new_[430]_  | \new_[431]_ ;
  assign \new_[5704]_  = \new_[432]_  | \new_[5703]_ ;
  assign \new_[5705]_  = \new_[5704]_  | \new_[5699]_ ;
  assign \new_[5706]_  = \new_[5705]_  | \new_[5696]_ ;
  assign \new_[5707]_  = \new_[5706]_  | \new_[5689]_ ;
  assign \new_[5710]_  = \new_[428]_  | \new_[429]_ ;
  assign \new_[5713]_  = \new_[426]_  | \new_[427]_ ;
  assign \new_[5714]_  = \new_[5713]_  | \new_[5710]_ ;
  assign \new_[5717]_  = \new_[424]_  | \new_[425]_ ;
  assign \new_[5721]_  = \new_[421]_  | \new_[422]_ ;
  assign \new_[5722]_  = \new_[423]_  | \new_[5721]_ ;
  assign \new_[5723]_  = \new_[5722]_  | \new_[5717]_ ;
  assign \new_[5724]_  = \new_[5723]_  | \new_[5714]_ ;
  assign \new_[5727]_  = \new_[419]_  | \new_[420]_ ;
  assign \new_[5730]_  = \new_[417]_  | \new_[418]_ ;
  assign \new_[5731]_  = \new_[5730]_  | \new_[5727]_ ;
  assign \new_[5734]_  = \new_[415]_  | \new_[416]_ ;
  assign \new_[5738]_  = \new_[412]_  | \new_[413]_ ;
  assign \new_[5739]_  = \new_[414]_  | \new_[5738]_ ;
  assign \new_[5740]_  = \new_[5739]_  | \new_[5734]_ ;
  assign \new_[5741]_  = \new_[5740]_  | \new_[5731]_ ;
  assign \new_[5742]_  = \new_[5741]_  | \new_[5724]_ ;
  assign \new_[5743]_  = \new_[5742]_  | \new_[5707]_ ;
  assign \new_[5744]_  = \new_[5743]_  | \new_[5674]_ ;
  assign \new_[5745]_  = \new_[5744]_  | \new_[5607]_ ;
  assign \new_[5748]_  = \new_[410]_  | \new_[411]_ ;
  assign \new_[5751]_  = \new_[408]_  | \new_[409]_ ;
  assign \new_[5752]_  = \new_[5751]_  | \new_[5748]_ ;
  assign \new_[5755]_  = \new_[406]_  | \new_[407]_ ;
  assign \new_[5758]_  = \new_[404]_  | \new_[405]_ ;
  assign \new_[5759]_  = \new_[5758]_  | \new_[5755]_ ;
  assign \new_[5760]_  = \new_[5759]_  | \new_[5752]_ ;
  assign \new_[5763]_  = \new_[402]_  | \new_[403]_ ;
  assign \new_[5766]_  = \new_[400]_  | \new_[401]_ ;
  assign \new_[5767]_  = \new_[5766]_  | \new_[5763]_ ;
  assign \new_[5770]_  = \new_[398]_  | \new_[399]_ ;
  assign \new_[5774]_  = \new_[395]_  | \new_[396]_ ;
  assign \new_[5775]_  = \new_[397]_  | \new_[5774]_ ;
  assign \new_[5776]_  = \new_[5775]_  | \new_[5770]_ ;
  assign \new_[5777]_  = \new_[5776]_  | \new_[5767]_ ;
  assign \new_[5778]_  = \new_[5777]_  | \new_[5760]_ ;
  assign \new_[5781]_  = \new_[393]_  | \new_[394]_ ;
  assign \new_[5784]_  = \new_[391]_  | \new_[392]_ ;
  assign \new_[5785]_  = \new_[5784]_  | \new_[5781]_ ;
  assign \new_[5788]_  = \new_[389]_  | \new_[390]_ ;
  assign \new_[5791]_  = \new_[387]_  | \new_[388]_ ;
  assign \new_[5792]_  = \new_[5791]_  | \new_[5788]_ ;
  assign \new_[5793]_  = \new_[5792]_  | \new_[5785]_ ;
  assign \new_[5796]_  = \new_[385]_  | \new_[386]_ ;
  assign \new_[5799]_  = \new_[383]_  | \new_[384]_ ;
  assign \new_[5800]_  = \new_[5799]_  | \new_[5796]_ ;
  assign \new_[5803]_  = \new_[381]_  | \new_[382]_ ;
  assign \new_[5807]_  = \new_[378]_  | \new_[379]_ ;
  assign \new_[5808]_  = \new_[380]_  | \new_[5807]_ ;
  assign \new_[5809]_  = \new_[5808]_  | \new_[5803]_ ;
  assign \new_[5810]_  = \new_[5809]_  | \new_[5800]_ ;
  assign \new_[5811]_  = \new_[5810]_  | \new_[5793]_ ;
  assign \new_[5812]_  = \new_[5811]_  | \new_[5778]_ ;
  assign \new_[5815]_  = \new_[376]_  | \new_[377]_ ;
  assign \new_[5818]_  = \new_[374]_  | \new_[375]_ ;
  assign \new_[5819]_  = \new_[5818]_  | \new_[5815]_ ;
  assign \new_[5822]_  = \new_[372]_  | \new_[373]_ ;
  assign \new_[5825]_  = \new_[370]_  | \new_[371]_ ;
  assign \new_[5826]_  = \new_[5825]_  | \new_[5822]_ ;
  assign \new_[5827]_  = \new_[5826]_  | \new_[5819]_ ;
  assign \new_[5830]_  = \new_[368]_  | \new_[369]_ ;
  assign \new_[5833]_  = \new_[366]_  | \new_[367]_ ;
  assign \new_[5834]_  = \new_[5833]_  | \new_[5830]_ ;
  assign \new_[5837]_  = \new_[364]_  | \new_[365]_ ;
  assign \new_[5841]_  = \new_[361]_  | \new_[362]_ ;
  assign \new_[5842]_  = \new_[363]_  | \new_[5841]_ ;
  assign \new_[5843]_  = \new_[5842]_  | \new_[5837]_ ;
  assign \new_[5844]_  = \new_[5843]_  | \new_[5834]_ ;
  assign \new_[5845]_  = \new_[5844]_  | \new_[5827]_ ;
  assign \new_[5848]_  = \new_[359]_  | \new_[360]_ ;
  assign \new_[5851]_  = \new_[357]_  | \new_[358]_ ;
  assign \new_[5852]_  = \new_[5851]_  | \new_[5848]_ ;
  assign \new_[5855]_  = \new_[355]_  | \new_[356]_ ;
  assign \new_[5858]_  = \new_[353]_  | \new_[354]_ ;
  assign \new_[5859]_  = \new_[5858]_  | \new_[5855]_ ;
  assign \new_[5860]_  = \new_[5859]_  | \new_[5852]_ ;
  assign \new_[5863]_  = \new_[351]_  | \new_[352]_ ;
  assign \new_[5866]_  = \new_[349]_  | \new_[350]_ ;
  assign \new_[5867]_  = \new_[5866]_  | \new_[5863]_ ;
  assign \new_[5870]_  = \new_[347]_  | \new_[348]_ ;
  assign \new_[5874]_  = \new_[344]_  | \new_[345]_ ;
  assign \new_[5875]_  = \new_[346]_  | \new_[5874]_ ;
  assign \new_[5876]_  = \new_[5875]_  | \new_[5870]_ ;
  assign \new_[5877]_  = \new_[5876]_  | \new_[5867]_ ;
  assign \new_[5878]_  = \new_[5877]_  | \new_[5860]_ ;
  assign \new_[5879]_  = \new_[5878]_  | \new_[5845]_ ;
  assign \new_[5880]_  = \new_[5879]_  | \new_[5812]_ ;
  assign \new_[5883]_  = \new_[342]_  | \new_[343]_ ;
  assign \new_[5886]_  = \new_[340]_  | \new_[341]_ ;
  assign \new_[5887]_  = \new_[5886]_  | \new_[5883]_ ;
  assign \new_[5890]_  = \new_[338]_  | \new_[339]_ ;
  assign \new_[5893]_  = \new_[336]_  | \new_[337]_ ;
  assign \new_[5894]_  = \new_[5893]_  | \new_[5890]_ ;
  assign \new_[5895]_  = \new_[5894]_  | \new_[5887]_ ;
  assign \new_[5898]_  = \new_[334]_  | \new_[335]_ ;
  assign \new_[5901]_  = \new_[332]_  | \new_[333]_ ;
  assign \new_[5902]_  = \new_[5901]_  | \new_[5898]_ ;
  assign \new_[5905]_  = \new_[330]_  | \new_[331]_ ;
  assign \new_[5909]_  = \new_[327]_  | \new_[328]_ ;
  assign \new_[5910]_  = \new_[329]_  | \new_[5909]_ ;
  assign \new_[5911]_  = \new_[5910]_  | \new_[5905]_ ;
  assign \new_[5912]_  = \new_[5911]_  | \new_[5902]_ ;
  assign \new_[5913]_  = \new_[5912]_  | \new_[5895]_ ;
  assign \new_[5916]_  = \new_[325]_  | \new_[326]_ ;
  assign \new_[5919]_  = \new_[323]_  | \new_[324]_ ;
  assign \new_[5920]_  = \new_[5919]_  | \new_[5916]_ ;
  assign \new_[5923]_  = \new_[321]_  | \new_[322]_ ;
  assign \new_[5926]_  = \new_[319]_  | \new_[320]_ ;
  assign \new_[5927]_  = \new_[5926]_  | \new_[5923]_ ;
  assign \new_[5928]_  = \new_[5927]_  | \new_[5920]_ ;
  assign \new_[5931]_  = \new_[317]_  | \new_[318]_ ;
  assign \new_[5934]_  = \new_[315]_  | \new_[316]_ ;
  assign \new_[5935]_  = \new_[5934]_  | \new_[5931]_ ;
  assign \new_[5938]_  = \new_[313]_  | \new_[314]_ ;
  assign \new_[5942]_  = \new_[310]_  | \new_[311]_ ;
  assign \new_[5943]_  = \new_[312]_  | \new_[5942]_ ;
  assign \new_[5944]_  = \new_[5943]_  | \new_[5938]_ ;
  assign \new_[5945]_  = \new_[5944]_  | \new_[5935]_ ;
  assign \new_[5946]_  = \new_[5945]_  | \new_[5928]_ ;
  assign \new_[5947]_  = \new_[5946]_  | \new_[5913]_ ;
  assign \new_[5950]_  = \new_[308]_  | \new_[309]_ ;
  assign \new_[5953]_  = \new_[306]_  | \new_[307]_ ;
  assign \new_[5954]_  = \new_[5953]_  | \new_[5950]_ ;
  assign \new_[5957]_  = \new_[304]_  | \new_[305]_ ;
  assign \new_[5960]_  = \new_[302]_  | \new_[303]_ ;
  assign \new_[5961]_  = \new_[5960]_  | \new_[5957]_ ;
  assign \new_[5962]_  = \new_[5961]_  | \new_[5954]_ ;
  assign \new_[5965]_  = \new_[300]_  | \new_[301]_ ;
  assign \new_[5968]_  = \new_[298]_  | \new_[299]_ ;
  assign \new_[5969]_  = \new_[5968]_  | \new_[5965]_ ;
  assign \new_[5972]_  = \new_[296]_  | \new_[297]_ ;
  assign \new_[5976]_  = \new_[293]_  | \new_[294]_ ;
  assign \new_[5977]_  = \new_[295]_  | \new_[5976]_ ;
  assign \new_[5978]_  = \new_[5977]_  | \new_[5972]_ ;
  assign \new_[5979]_  = \new_[5978]_  | \new_[5969]_ ;
  assign \new_[5980]_  = \new_[5979]_  | \new_[5962]_ ;
  assign \new_[5983]_  = \new_[291]_  | \new_[292]_ ;
  assign \new_[5986]_  = \new_[289]_  | \new_[290]_ ;
  assign \new_[5987]_  = \new_[5986]_  | \new_[5983]_ ;
  assign \new_[5990]_  = \new_[287]_  | \new_[288]_ ;
  assign \new_[5994]_  = \new_[284]_  | \new_[285]_ ;
  assign \new_[5995]_  = \new_[286]_  | \new_[5994]_ ;
  assign \new_[5996]_  = \new_[5995]_  | \new_[5990]_ ;
  assign \new_[5997]_  = \new_[5996]_  | \new_[5987]_ ;
  assign \new_[6000]_  = \new_[282]_  | \new_[283]_ ;
  assign \new_[6003]_  = \new_[280]_  | \new_[281]_ ;
  assign \new_[6004]_  = \new_[6003]_  | \new_[6000]_ ;
  assign \new_[6007]_  = \new_[278]_  | \new_[279]_ ;
  assign \new_[6011]_  = \new_[275]_  | \new_[276]_ ;
  assign \new_[6012]_  = \new_[277]_  | \new_[6011]_ ;
  assign \new_[6013]_  = \new_[6012]_  | \new_[6007]_ ;
  assign \new_[6014]_  = \new_[6013]_  | \new_[6004]_ ;
  assign \new_[6015]_  = \new_[6014]_  | \new_[5997]_ ;
  assign \new_[6016]_  = \new_[6015]_  | \new_[5980]_ ;
  assign \new_[6017]_  = \new_[6016]_  | \new_[5947]_ ;
  assign \new_[6018]_  = \new_[6017]_  | \new_[5880]_ ;
  assign \new_[6019]_  = \new_[6018]_  | \new_[5745]_ ;
  assign \new_[6022]_  = \new_[273]_  | \new_[274]_ ;
  assign \new_[6025]_  = \new_[271]_  | \new_[272]_ ;
  assign \new_[6026]_  = \new_[6025]_  | \new_[6022]_ ;
  assign \new_[6029]_  = \new_[269]_  | \new_[270]_ ;
  assign \new_[6032]_  = \new_[267]_  | \new_[268]_ ;
  assign \new_[6033]_  = \new_[6032]_  | \new_[6029]_ ;
  assign \new_[6034]_  = \new_[6033]_  | \new_[6026]_ ;
  assign \new_[6037]_  = \new_[265]_  | \new_[266]_ ;
  assign \new_[6040]_  = \new_[263]_  | \new_[264]_ ;
  assign \new_[6041]_  = \new_[6040]_  | \new_[6037]_ ;
  assign \new_[6044]_  = \new_[261]_  | \new_[262]_ ;
  assign \new_[6048]_  = \new_[258]_  | \new_[259]_ ;
  assign \new_[6049]_  = \new_[260]_  | \new_[6048]_ ;
  assign \new_[6050]_  = \new_[6049]_  | \new_[6044]_ ;
  assign \new_[6051]_  = \new_[6050]_  | \new_[6041]_ ;
  assign \new_[6052]_  = \new_[6051]_  | \new_[6034]_ ;
  assign \new_[6055]_  = \new_[256]_  | \new_[257]_ ;
  assign \new_[6058]_  = \new_[254]_  | \new_[255]_ ;
  assign \new_[6059]_  = \new_[6058]_  | \new_[6055]_ ;
  assign \new_[6062]_  = \new_[252]_  | \new_[253]_ ;
  assign \new_[6065]_  = \new_[250]_  | \new_[251]_ ;
  assign \new_[6066]_  = \new_[6065]_  | \new_[6062]_ ;
  assign \new_[6067]_  = \new_[6066]_  | \new_[6059]_ ;
  assign \new_[6070]_  = \new_[248]_  | \new_[249]_ ;
  assign \new_[6073]_  = \new_[246]_  | \new_[247]_ ;
  assign \new_[6074]_  = \new_[6073]_  | \new_[6070]_ ;
  assign \new_[6077]_  = \new_[244]_  | \new_[245]_ ;
  assign \new_[6081]_  = \new_[241]_  | \new_[242]_ ;
  assign \new_[6082]_  = \new_[243]_  | \new_[6081]_ ;
  assign \new_[6083]_  = \new_[6082]_  | \new_[6077]_ ;
  assign \new_[6084]_  = \new_[6083]_  | \new_[6074]_ ;
  assign \new_[6085]_  = \new_[6084]_  | \new_[6067]_ ;
  assign \new_[6086]_  = \new_[6085]_  | \new_[6052]_ ;
  assign \new_[6089]_  = \new_[239]_  | \new_[240]_ ;
  assign \new_[6092]_  = \new_[237]_  | \new_[238]_ ;
  assign \new_[6093]_  = \new_[6092]_  | \new_[6089]_ ;
  assign \new_[6096]_  = \new_[235]_  | \new_[236]_ ;
  assign \new_[6099]_  = \new_[233]_  | \new_[234]_ ;
  assign \new_[6100]_  = \new_[6099]_  | \new_[6096]_ ;
  assign \new_[6101]_  = \new_[6100]_  | \new_[6093]_ ;
  assign \new_[6104]_  = \new_[231]_  | \new_[232]_ ;
  assign \new_[6107]_  = \new_[229]_  | \new_[230]_ ;
  assign \new_[6108]_  = \new_[6107]_  | \new_[6104]_ ;
  assign \new_[6111]_  = \new_[227]_  | \new_[228]_ ;
  assign \new_[6115]_  = \new_[224]_  | \new_[225]_ ;
  assign \new_[6116]_  = \new_[226]_  | \new_[6115]_ ;
  assign \new_[6117]_  = \new_[6116]_  | \new_[6111]_ ;
  assign \new_[6118]_  = \new_[6117]_  | \new_[6108]_ ;
  assign \new_[6119]_  = \new_[6118]_  | \new_[6101]_ ;
  assign \new_[6122]_  = \new_[222]_  | \new_[223]_ ;
  assign \new_[6125]_  = \new_[220]_  | \new_[221]_ ;
  assign \new_[6126]_  = \new_[6125]_  | \new_[6122]_ ;
  assign \new_[6129]_  = \new_[218]_  | \new_[219]_ ;
  assign \new_[6132]_  = \new_[216]_  | \new_[217]_ ;
  assign \new_[6133]_  = \new_[6132]_  | \new_[6129]_ ;
  assign \new_[6134]_  = \new_[6133]_  | \new_[6126]_ ;
  assign \new_[6137]_  = \new_[214]_  | \new_[215]_ ;
  assign \new_[6140]_  = \new_[212]_  | \new_[213]_ ;
  assign \new_[6141]_  = \new_[6140]_  | \new_[6137]_ ;
  assign \new_[6144]_  = \new_[210]_  | \new_[211]_ ;
  assign \new_[6148]_  = \new_[207]_  | \new_[208]_ ;
  assign \new_[6149]_  = \new_[209]_  | \new_[6148]_ ;
  assign \new_[6150]_  = \new_[6149]_  | \new_[6144]_ ;
  assign \new_[6151]_  = \new_[6150]_  | \new_[6141]_ ;
  assign \new_[6152]_  = \new_[6151]_  | \new_[6134]_ ;
  assign \new_[6153]_  = \new_[6152]_  | \new_[6119]_ ;
  assign \new_[6154]_  = \new_[6153]_  | \new_[6086]_ ;
  assign \new_[6157]_  = \new_[205]_  | \new_[206]_ ;
  assign \new_[6160]_  = \new_[203]_  | \new_[204]_ ;
  assign \new_[6161]_  = \new_[6160]_  | \new_[6157]_ ;
  assign \new_[6164]_  = \new_[201]_  | \new_[202]_ ;
  assign \new_[6167]_  = \new_[199]_  | \new_[200]_ ;
  assign \new_[6168]_  = \new_[6167]_  | \new_[6164]_ ;
  assign \new_[6169]_  = \new_[6168]_  | \new_[6161]_ ;
  assign \new_[6172]_  = \new_[197]_  | \new_[198]_ ;
  assign \new_[6175]_  = \new_[195]_  | \new_[196]_ ;
  assign \new_[6176]_  = \new_[6175]_  | \new_[6172]_ ;
  assign \new_[6179]_  = \new_[193]_  | \new_[194]_ ;
  assign \new_[6183]_  = \new_[190]_  | \new_[191]_ ;
  assign \new_[6184]_  = \new_[192]_  | \new_[6183]_ ;
  assign \new_[6185]_  = \new_[6184]_  | \new_[6179]_ ;
  assign \new_[6186]_  = \new_[6185]_  | \new_[6176]_ ;
  assign \new_[6187]_  = \new_[6186]_  | \new_[6169]_ ;
  assign \new_[6190]_  = \new_[188]_  | \new_[189]_ ;
  assign \new_[6193]_  = \new_[186]_  | \new_[187]_ ;
  assign \new_[6194]_  = \new_[6193]_  | \new_[6190]_ ;
  assign \new_[6197]_  = \new_[184]_  | \new_[185]_ ;
  assign \new_[6200]_  = \new_[182]_  | \new_[183]_ ;
  assign \new_[6201]_  = \new_[6200]_  | \new_[6197]_ ;
  assign \new_[6202]_  = \new_[6201]_  | \new_[6194]_ ;
  assign \new_[6205]_  = \new_[180]_  | \new_[181]_ ;
  assign \new_[6208]_  = \new_[178]_  | \new_[179]_ ;
  assign \new_[6209]_  = \new_[6208]_  | \new_[6205]_ ;
  assign \new_[6212]_  = \new_[176]_  | \new_[177]_ ;
  assign \new_[6216]_  = \new_[173]_  | \new_[174]_ ;
  assign \new_[6217]_  = \new_[175]_  | \new_[6216]_ ;
  assign \new_[6218]_  = \new_[6217]_  | \new_[6212]_ ;
  assign \new_[6219]_  = \new_[6218]_  | \new_[6209]_ ;
  assign \new_[6220]_  = \new_[6219]_  | \new_[6202]_ ;
  assign \new_[6221]_  = \new_[6220]_  | \new_[6187]_ ;
  assign \new_[6224]_  = \new_[171]_  | \new_[172]_ ;
  assign \new_[6227]_  = \new_[169]_  | \new_[170]_ ;
  assign \new_[6228]_  = \new_[6227]_  | \new_[6224]_ ;
  assign \new_[6231]_  = \new_[167]_  | \new_[168]_ ;
  assign \new_[6234]_  = \new_[165]_  | \new_[166]_ ;
  assign \new_[6235]_  = \new_[6234]_  | \new_[6231]_ ;
  assign \new_[6236]_  = \new_[6235]_  | \new_[6228]_ ;
  assign \new_[6239]_  = \new_[163]_  | \new_[164]_ ;
  assign \new_[6242]_  = \new_[161]_  | \new_[162]_ ;
  assign \new_[6243]_  = \new_[6242]_  | \new_[6239]_ ;
  assign \new_[6246]_  = \new_[159]_  | \new_[160]_ ;
  assign \new_[6250]_  = \new_[156]_  | \new_[157]_ ;
  assign \new_[6251]_  = \new_[158]_  | \new_[6250]_ ;
  assign \new_[6252]_  = \new_[6251]_  | \new_[6246]_ ;
  assign \new_[6253]_  = \new_[6252]_  | \new_[6243]_ ;
  assign \new_[6254]_  = \new_[6253]_  | \new_[6236]_ ;
  assign \new_[6257]_  = \new_[154]_  | \new_[155]_ ;
  assign \new_[6260]_  = \new_[152]_  | \new_[153]_ ;
  assign \new_[6261]_  = \new_[6260]_  | \new_[6257]_ ;
  assign \new_[6264]_  = \new_[150]_  | \new_[151]_ ;
  assign \new_[6268]_  = \new_[147]_  | \new_[148]_ ;
  assign \new_[6269]_  = \new_[149]_  | \new_[6268]_ ;
  assign \new_[6270]_  = \new_[6269]_  | \new_[6264]_ ;
  assign \new_[6271]_  = \new_[6270]_  | \new_[6261]_ ;
  assign \new_[6274]_  = \new_[145]_  | \new_[146]_ ;
  assign \new_[6277]_  = \new_[143]_  | \new_[144]_ ;
  assign \new_[6278]_  = \new_[6277]_  | \new_[6274]_ ;
  assign \new_[6281]_  = \new_[141]_  | \new_[142]_ ;
  assign \new_[6285]_  = \new_[138]_  | \new_[139]_ ;
  assign \new_[6286]_  = \new_[140]_  | \new_[6285]_ ;
  assign \new_[6287]_  = \new_[6286]_  | \new_[6281]_ ;
  assign \new_[6288]_  = \new_[6287]_  | \new_[6278]_ ;
  assign \new_[6289]_  = \new_[6288]_  | \new_[6271]_ ;
  assign \new_[6290]_  = \new_[6289]_  | \new_[6254]_ ;
  assign \new_[6291]_  = \new_[6290]_  | \new_[6221]_ ;
  assign \new_[6292]_  = \new_[6291]_  | \new_[6154]_ ;
  assign \new_[6295]_  = \new_[136]_  | \new_[137]_ ;
  assign \new_[6298]_  = \new_[134]_  | \new_[135]_ ;
  assign \new_[6299]_  = \new_[6298]_  | \new_[6295]_ ;
  assign \new_[6302]_  = \new_[132]_  | \new_[133]_ ;
  assign \new_[6305]_  = \new_[130]_  | \new_[131]_ ;
  assign \new_[6306]_  = \new_[6305]_  | \new_[6302]_ ;
  assign \new_[6307]_  = \new_[6306]_  | \new_[6299]_ ;
  assign \new_[6310]_  = \new_[128]_  | \new_[129]_ ;
  assign \new_[6313]_  = \new_[126]_  | \new_[127]_ ;
  assign \new_[6314]_  = \new_[6313]_  | \new_[6310]_ ;
  assign \new_[6317]_  = \new_[124]_  | \new_[125]_ ;
  assign \new_[6321]_  = \new_[121]_  | \new_[122]_ ;
  assign \new_[6322]_  = \new_[123]_  | \new_[6321]_ ;
  assign \new_[6323]_  = \new_[6322]_  | \new_[6317]_ ;
  assign \new_[6324]_  = \new_[6323]_  | \new_[6314]_ ;
  assign \new_[6325]_  = \new_[6324]_  | \new_[6307]_ ;
  assign \new_[6328]_  = \new_[119]_  | \new_[120]_ ;
  assign \new_[6331]_  = \new_[117]_  | \new_[118]_ ;
  assign \new_[6332]_  = \new_[6331]_  | \new_[6328]_ ;
  assign \new_[6335]_  = \new_[115]_  | \new_[116]_ ;
  assign \new_[6338]_  = \new_[113]_  | \new_[114]_ ;
  assign \new_[6339]_  = \new_[6338]_  | \new_[6335]_ ;
  assign \new_[6340]_  = \new_[6339]_  | \new_[6332]_ ;
  assign \new_[6343]_  = \new_[111]_  | \new_[112]_ ;
  assign \new_[6346]_  = \new_[109]_  | \new_[110]_ ;
  assign \new_[6347]_  = \new_[6346]_  | \new_[6343]_ ;
  assign \new_[6350]_  = \new_[107]_  | \new_[108]_ ;
  assign \new_[6354]_  = \new_[104]_  | \new_[105]_ ;
  assign \new_[6355]_  = \new_[106]_  | \new_[6354]_ ;
  assign \new_[6356]_  = \new_[6355]_  | \new_[6350]_ ;
  assign \new_[6357]_  = \new_[6356]_  | \new_[6347]_ ;
  assign \new_[6358]_  = \new_[6357]_  | \new_[6340]_ ;
  assign \new_[6359]_  = \new_[6358]_  | \new_[6325]_ ;
  assign \new_[6362]_  = \new_[102]_  | \new_[103]_ ;
  assign \new_[6365]_  = \new_[100]_  | \new_[101]_ ;
  assign \new_[6366]_  = \new_[6365]_  | \new_[6362]_ ;
  assign \new_[6369]_  = \new_[98]_  | \new_[99]_ ;
  assign \new_[6372]_  = \new_[96]_  | \new_[97]_ ;
  assign \new_[6373]_  = \new_[6372]_  | \new_[6369]_ ;
  assign \new_[6374]_  = \new_[6373]_  | \new_[6366]_ ;
  assign \new_[6377]_  = \new_[94]_  | \new_[95]_ ;
  assign \new_[6380]_  = \new_[92]_  | \new_[93]_ ;
  assign \new_[6381]_  = \new_[6380]_  | \new_[6377]_ ;
  assign \new_[6384]_  = \new_[90]_  | \new_[91]_ ;
  assign \new_[6388]_  = \new_[87]_  | \new_[88]_ ;
  assign \new_[6389]_  = \new_[89]_  | \new_[6388]_ ;
  assign \new_[6390]_  = \new_[6389]_  | \new_[6384]_ ;
  assign \new_[6391]_  = \new_[6390]_  | \new_[6381]_ ;
  assign \new_[6392]_  = \new_[6391]_  | \new_[6374]_ ;
  assign \new_[6395]_  = \new_[85]_  | \new_[86]_ ;
  assign \new_[6398]_  = \new_[83]_  | \new_[84]_ ;
  assign \new_[6399]_  = \new_[6398]_  | \new_[6395]_ ;
  assign \new_[6402]_  = \new_[81]_  | \new_[82]_ ;
  assign \new_[6405]_  = \new_[79]_  | \new_[80]_ ;
  assign \new_[6406]_  = \new_[6405]_  | \new_[6402]_ ;
  assign \new_[6407]_  = \new_[6406]_  | \new_[6399]_ ;
  assign \new_[6410]_  = \new_[77]_  | \new_[78]_ ;
  assign \new_[6413]_  = \new_[75]_  | \new_[76]_ ;
  assign \new_[6414]_  = \new_[6413]_  | \new_[6410]_ ;
  assign \new_[6417]_  = \new_[73]_  | \new_[74]_ ;
  assign \new_[6421]_  = \new_[70]_  | \new_[71]_ ;
  assign \new_[6422]_  = \new_[72]_  | \new_[6421]_ ;
  assign \new_[6423]_  = \new_[6422]_  | \new_[6417]_ ;
  assign \new_[6424]_  = \new_[6423]_  | \new_[6414]_ ;
  assign \new_[6425]_  = \new_[6424]_  | \new_[6407]_ ;
  assign \new_[6426]_  = \new_[6425]_  | \new_[6392]_ ;
  assign \new_[6427]_  = \new_[6426]_  | \new_[6359]_ ;
  assign \new_[6430]_  = \new_[68]_  | \new_[69]_ ;
  assign \new_[6433]_  = \new_[66]_  | \new_[67]_ ;
  assign \new_[6434]_  = \new_[6433]_  | \new_[6430]_ ;
  assign \new_[6437]_  = \new_[64]_  | \new_[65]_ ;
  assign \new_[6440]_  = \new_[62]_  | \new_[63]_ ;
  assign \new_[6441]_  = \new_[6440]_  | \new_[6437]_ ;
  assign \new_[6442]_  = \new_[6441]_  | \new_[6434]_ ;
  assign \new_[6445]_  = \new_[60]_  | \new_[61]_ ;
  assign \new_[6448]_  = \new_[58]_  | \new_[59]_ ;
  assign \new_[6449]_  = \new_[6448]_  | \new_[6445]_ ;
  assign \new_[6452]_  = \new_[56]_  | \new_[57]_ ;
  assign \new_[6456]_  = \new_[53]_  | \new_[54]_ ;
  assign \new_[6457]_  = \new_[55]_  | \new_[6456]_ ;
  assign \new_[6458]_  = \new_[6457]_  | \new_[6452]_ ;
  assign \new_[6459]_  = \new_[6458]_  | \new_[6449]_ ;
  assign \new_[6460]_  = \new_[6459]_  | \new_[6442]_ ;
  assign \new_[6463]_  = \new_[51]_  | \new_[52]_ ;
  assign \new_[6466]_  = \new_[49]_  | \new_[50]_ ;
  assign \new_[6467]_  = \new_[6466]_  | \new_[6463]_ ;
  assign \new_[6470]_  = \new_[47]_  | \new_[48]_ ;
  assign \new_[6473]_  = \new_[45]_  | \new_[46]_ ;
  assign \new_[6474]_  = \new_[6473]_  | \new_[6470]_ ;
  assign \new_[6475]_  = \new_[6474]_  | \new_[6467]_ ;
  assign \new_[6478]_  = \new_[43]_  | \new_[44]_ ;
  assign \new_[6481]_  = \new_[41]_  | \new_[42]_ ;
  assign \new_[6482]_  = \new_[6481]_  | \new_[6478]_ ;
  assign \new_[6485]_  = \new_[39]_  | \new_[40]_ ;
  assign \new_[6489]_  = \new_[36]_  | \new_[37]_ ;
  assign \new_[6490]_  = \new_[38]_  | \new_[6489]_ ;
  assign \new_[6491]_  = \new_[6490]_  | \new_[6485]_ ;
  assign \new_[6492]_  = \new_[6491]_  | \new_[6482]_ ;
  assign \new_[6493]_  = \new_[6492]_  | \new_[6475]_ ;
  assign \new_[6494]_  = \new_[6493]_  | \new_[6460]_ ;
  assign \new_[6497]_  = \new_[34]_  | \new_[35]_ ;
  assign \new_[6500]_  = \new_[32]_  | \new_[33]_ ;
  assign \new_[6501]_  = \new_[6500]_  | \new_[6497]_ ;
  assign \new_[6504]_  = \new_[30]_  | \new_[31]_ ;
  assign \new_[6507]_  = \new_[28]_  | \new_[29]_ ;
  assign \new_[6508]_  = \new_[6507]_  | \new_[6504]_ ;
  assign \new_[6509]_  = \new_[6508]_  | \new_[6501]_ ;
  assign \new_[6512]_  = \new_[26]_  | \new_[27]_ ;
  assign \new_[6515]_  = \new_[24]_  | \new_[25]_ ;
  assign \new_[6516]_  = \new_[6515]_  | \new_[6512]_ ;
  assign \new_[6519]_  = \new_[22]_  | \new_[23]_ ;
  assign \new_[6523]_  = \new_[19]_  | \new_[20]_ ;
  assign \new_[6524]_  = \new_[21]_  | \new_[6523]_ ;
  assign \new_[6525]_  = \new_[6524]_  | \new_[6519]_ ;
  assign \new_[6526]_  = \new_[6525]_  | \new_[6516]_ ;
  assign \new_[6527]_  = \new_[6526]_  | \new_[6509]_ ;
  assign \new_[6530]_  = \new_[17]_  | \new_[18]_ ;
  assign \new_[6533]_  = \new_[15]_  | \new_[16]_ ;
  assign \new_[6534]_  = \new_[6533]_  | \new_[6530]_ ;
  assign \new_[6537]_  = \new_[13]_  | \new_[14]_ ;
  assign \new_[6541]_  = \new_[10]_  | \new_[11]_ ;
  assign \new_[6542]_  = \new_[12]_  | \new_[6541]_ ;
  assign \new_[6543]_  = \new_[6542]_  | \new_[6537]_ ;
  assign \new_[6544]_  = \new_[6543]_  | \new_[6534]_ ;
  assign \new_[6547]_  = \new_[8]_  | \new_[9]_ ;
  assign \new_[6550]_  = \new_[6]_  | \new_[7]_ ;
  assign \new_[6551]_  = \new_[6550]_  | \new_[6547]_ ;
  assign \new_[6554]_  = \new_[4]_  | \new_[5]_ ;
  assign \new_[6558]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[6559]_  = \new_[3]_  | \new_[6558]_ ;
  assign \new_[6560]_  = \new_[6559]_  | \new_[6554]_ ;
  assign \new_[6561]_  = \new_[6560]_  | \new_[6551]_ ;
  assign \new_[6562]_  = \new_[6561]_  | \new_[6544]_ ;
  assign \new_[6563]_  = \new_[6562]_  | \new_[6527]_ ;
  assign \new_[6564]_  = \new_[6563]_  | \new_[6494]_ ;
  assign \new_[6565]_  = \new_[6564]_  | \new_[6427]_ ;
  assign \new_[6566]_  = \new_[6565]_  | \new_[6292]_ ;
  assign \new_[6567]_  = \new_[6566]_  | \new_[6019]_ ;
  assign \new_[6568]_  = \new_[6567]_  | \new_[5472]_ ;
  assign \new_[6572]_  = A267 & A266;
  assign \new_[6573]_  = ~A265 & \new_[6572]_ ;
  assign \new_[6577]_  = A301 & ~A300;
  assign \new_[6578]_  = A268 & \new_[6577]_ ;
  assign \new_[6582]_  = A267 & A266;
  assign \new_[6583]_  = ~A265 & \new_[6582]_ ;
  assign \new_[6587]_  = ~A302 & ~A300;
  assign \new_[6588]_  = A268 & \new_[6587]_ ;
  assign \new_[6592]_  = A267 & A266;
  assign \new_[6593]_  = ~A265 & \new_[6592]_ ;
  assign \new_[6597]_  = A299 & A298;
  assign \new_[6598]_  = A268 & \new_[6597]_ ;
  assign \new_[6602]_  = A267 & A266;
  assign \new_[6603]_  = ~A265 & \new_[6602]_ ;
  assign \new_[6607]_  = ~A299 & ~A298;
  assign \new_[6608]_  = A268 & \new_[6607]_ ;
  assign \new_[6612]_  = A267 & A266;
  assign \new_[6613]_  = ~A265 & \new_[6612]_ ;
  assign \new_[6617]_  = A301 & ~A300;
  assign \new_[6618]_  = ~A269 & \new_[6617]_ ;
  assign \new_[6622]_  = A267 & A266;
  assign \new_[6623]_  = ~A265 & \new_[6622]_ ;
  assign \new_[6627]_  = ~A302 & ~A300;
  assign \new_[6628]_  = ~A269 & \new_[6627]_ ;
  assign \new_[6632]_  = A267 & A266;
  assign \new_[6633]_  = ~A265 & \new_[6632]_ ;
  assign \new_[6637]_  = A299 & A298;
  assign \new_[6638]_  = ~A269 & \new_[6637]_ ;
  assign \new_[6642]_  = A267 & A266;
  assign \new_[6643]_  = ~A265 & \new_[6642]_ ;
  assign \new_[6647]_  = ~A299 & ~A298;
  assign \new_[6648]_  = ~A269 & \new_[6647]_ ;
  assign \new_[6652]_  = A267 & ~A266;
  assign \new_[6653]_  = A265 & \new_[6652]_ ;
  assign \new_[6657]_  = A301 & ~A300;
  assign \new_[6658]_  = A268 & \new_[6657]_ ;
  assign \new_[6662]_  = A267 & ~A266;
  assign \new_[6663]_  = A265 & \new_[6662]_ ;
  assign \new_[6667]_  = ~A302 & ~A300;
  assign \new_[6668]_  = A268 & \new_[6667]_ ;
  assign \new_[6672]_  = A267 & ~A266;
  assign \new_[6673]_  = A265 & \new_[6672]_ ;
  assign \new_[6677]_  = A299 & A298;
  assign \new_[6678]_  = A268 & \new_[6677]_ ;
  assign \new_[6682]_  = A267 & ~A266;
  assign \new_[6683]_  = A265 & \new_[6682]_ ;
  assign \new_[6687]_  = ~A299 & ~A298;
  assign \new_[6688]_  = A268 & \new_[6687]_ ;
  assign \new_[6692]_  = A267 & ~A266;
  assign \new_[6693]_  = A265 & \new_[6692]_ ;
  assign \new_[6697]_  = A301 & ~A300;
  assign \new_[6698]_  = ~A269 & \new_[6697]_ ;
  assign \new_[6702]_  = A267 & ~A266;
  assign \new_[6703]_  = A265 & \new_[6702]_ ;
  assign \new_[6707]_  = ~A302 & ~A300;
  assign \new_[6708]_  = ~A269 & \new_[6707]_ ;
  assign \new_[6712]_  = A267 & ~A266;
  assign \new_[6713]_  = A265 & \new_[6712]_ ;
  assign \new_[6717]_  = A299 & A298;
  assign \new_[6718]_  = ~A269 & \new_[6717]_ ;
  assign \new_[6722]_  = A267 & ~A266;
  assign \new_[6723]_  = A265 & \new_[6722]_ ;
  assign \new_[6727]_  = ~A299 & ~A298;
  assign \new_[6728]_  = ~A269 & \new_[6727]_ ;
  assign \new_[6732]_  = A267 & A266;
  assign \new_[6733]_  = ~A265 & \new_[6732]_ ;
  assign \new_[6736]_  = A300 & A268;
  assign \new_[6739]_  = A302 & ~A301;
  assign \new_[6740]_  = \new_[6739]_  & \new_[6736]_ ;
  assign \new_[6744]_  = A267 & A266;
  assign \new_[6745]_  = ~A265 & \new_[6744]_ ;
  assign \new_[6748]_  = A300 & ~A269;
  assign \new_[6751]_  = A302 & ~A301;
  assign \new_[6752]_  = \new_[6751]_  & \new_[6748]_ ;
  assign \new_[6756]_  = ~A267 & A266;
  assign \new_[6757]_  = ~A265 & \new_[6756]_ ;
  assign \new_[6760]_  = A269 & ~A268;
  assign \new_[6763]_  = A301 & ~A300;
  assign \new_[6764]_  = \new_[6763]_  & \new_[6760]_ ;
  assign \new_[6768]_  = ~A267 & A266;
  assign \new_[6769]_  = ~A265 & \new_[6768]_ ;
  assign \new_[6772]_  = A269 & ~A268;
  assign \new_[6775]_  = ~A302 & ~A300;
  assign \new_[6776]_  = \new_[6775]_  & \new_[6772]_ ;
  assign \new_[6780]_  = ~A267 & A266;
  assign \new_[6781]_  = ~A265 & \new_[6780]_ ;
  assign \new_[6784]_  = A269 & ~A268;
  assign \new_[6787]_  = A299 & A298;
  assign \new_[6788]_  = \new_[6787]_  & \new_[6784]_ ;
  assign \new_[6792]_  = ~A267 & A266;
  assign \new_[6793]_  = ~A265 & \new_[6792]_ ;
  assign \new_[6796]_  = A269 & ~A268;
  assign \new_[6799]_  = ~A299 & ~A298;
  assign \new_[6800]_  = \new_[6799]_  & \new_[6796]_ ;
  assign \new_[6804]_  = A267 & ~A266;
  assign \new_[6805]_  = A265 & \new_[6804]_ ;
  assign \new_[6808]_  = A300 & A268;
  assign \new_[6811]_  = A302 & ~A301;
  assign \new_[6812]_  = \new_[6811]_  & \new_[6808]_ ;
  assign \new_[6816]_  = A267 & ~A266;
  assign \new_[6817]_  = A265 & \new_[6816]_ ;
  assign \new_[6820]_  = A300 & ~A269;
  assign \new_[6823]_  = A302 & ~A301;
  assign \new_[6824]_  = \new_[6823]_  & \new_[6820]_ ;
  assign \new_[6828]_  = ~A267 & ~A266;
  assign \new_[6829]_  = A265 & \new_[6828]_ ;
  assign \new_[6832]_  = A269 & ~A268;
  assign \new_[6835]_  = A301 & ~A300;
  assign \new_[6836]_  = \new_[6835]_  & \new_[6832]_ ;
  assign \new_[6840]_  = ~A267 & ~A266;
  assign \new_[6841]_  = A265 & \new_[6840]_ ;
  assign \new_[6844]_  = A269 & ~A268;
  assign \new_[6847]_  = ~A302 & ~A300;
  assign \new_[6848]_  = \new_[6847]_  & \new_[6844]_ ;
  assign \new_[6852]_  = ~A267 & ~A266;
  assign \new_[6853]_  = A265 & \new_[6852]_ ;
  assign \new_[6856]_  = A269 & ~A268;
  assign \new_[6859]_  = A299 & A298;
  assign \new_[6860]_  = \new_[6859]_  & \new_[6856]_ ;
  assign \new_[6864]_  = ~A267 & ~A266;
  assign \new_[6865]_  = A265 & \new_[6864]_ ;
  assign \new_[6868]_  = A269 & ~A268;
  assign \new_[6871]_  = ~A299 & ~A298;
  assign \new_[6872]_  = \new_[6871]_  & \new_[6868]_ ;
  assign \new_[6875]_  = A266 & ~A265;
  assign \new_[6878]_  = ~A268 & ~A267;
  assign \new_[6879]_  = \new_[6878]_  & \new_[6875]_ ;
  assign \new_[6882]_  = A300 & A269;
  assign \new_[6885]_  = A302 & ~A301;
  assign \new_[6886]_  = \new_[6885]_  & \new_[6882]_ ;
  assign \new_[6889]_  = ~A266 & A265;
  assign \new_[6892]_  = ~A268 & ~A267;
  assign \new_[6893]_  = \new_[6892]_  & \new_[6889]_ ;
  assign \new_[6896]_  = A300 & A269;
  assign \new_[6899]_  = A302 & ~A301;
  assign \new_[6900]_  = \new_[6899]_  & \new_[6896]_ ;
  assign \new_[6904]_  = A201 & A200;
  assign \new_[6905]_  = ~A199 & \new_[6904]_ ;
  assign \new_[6908]_  = ~A232 & A202;
  assign \new_[6911]_  = A234 & A233;
  assign \new_[6912]_  = \new_[6911]_  & \new_[6908]_ ;
  assign \new_[6913]_  = \new_[6912]_  & \new_[6905]_ ;
  assign \new_[6917]_  = A268 & ~A267;
  assign \new_[6918]_  = A235 & \new_[6917]_ ;
  assign \new_[6921]_  = ~A299 & A298;
  assign \new_[6924]_  = A301 & A300;
  assign \new_[6925]_  = \new_[6924]_  & \new_[6921]_ ;
  assign \new_[6926]_  = \new_[6925]_  & \new_[6918]_ ;
  assign \new_[6930]_  = A201 & A200;
  assign \new_[6931]_  = ~A199 & \new_[6930]_ ;
  assign \new_[6934]_  = ~A232 & A202;
  assign \new_[6937]_  = A234 & A233;
  assign \new_[6938]_  = \new_[6937]_  & \new_[6934]_ ;
  assign \new_[6939]_  = \new_[6938]_  & \new_[6931]_ ;
  assign \new_[6943]_  = A268 & ~A267;
  assign \new_[6944]_  = A235 & \new_[6943]_ ;
  assign \new_[6947]_  = ~A299 & A298;
  assign \new_[6950]_  = ~A302 & A300;
  assign \new_[6951]_  = \new_[6950]_  & \new_[6947]_ ;
  assign \new_[6952]_  = \new_[6951]_  & \new_[6944]_ ;
  assign \new_[6956]_  = A201 & A200;
  assign \new_[6957]_  = ~A199 & \new_[6956]_ ;
  assign \new_[6960]_  = ~A232 & A202;
  assign \new_[6963]_  = A234 & A233;
  assign \new_[6964]_  = \new_[6963]_  & \new_[6960]_ ;
  assign \new_[6965]_  = \new_[6964]_  & \new_[6957]_ ;
  assign \new_[6969]_  = A268 & ~A267;
  assign \new_[6970]_  = A235 & \new_[6969]_ ;
  assign \new_[6973]_  = A299 & ~A298;
  assign \new_[6976]_  = A301 & A300;
  assign \new_[6977]_  = \new_[6976]_  & \new_[6973]_ ;
  assign \new_[6978]_  = \new_[6977]_  & \new_[6970]_ ;
  assign \new_[6982]_  = A201 & A200;
  assign \new_[6983]_  = ~A199 & \new_[6982]_ ;
  assign \new_[6986]_  = ~A232 & A202;
  assign \new_[6989]_  = A234 & A233;
  assign \new_[6990]_  = \new_[6989]_  & \new_[6986]_ ;
  assign \new_[6991]_  = \new_[6990]_  & \new_[6983]_ ;
  assign \new_[6995]_  = A268 & ~A267;
  assign \new_[6996]_  = A235 & \new_[6995]_ ;
  assign \new_[6999]_  = A299 & ~A298;
  assign \new_[7002]_  = ~A302 & A300;
  assign \new_[7003]_  = \new_[7002]_  & \new_[6999]_ ;
  assign \new_[7004]_  = \new_[7003]_  & \new_[6996]_ ;
  assign \new_[7008]_  = A201 & A200;
  assign \new_[7009]_  = ~A199 & \new_[7008]_ ;
  assign \new_[7012]_  = ~A232 & A202;
  assign \new_[7015]_  = A234 & A233;
  assign \new_[7016]_  = \new_[7015]_  & \new_[7012]_ ;
  assign \new_[7017]_  = \new_[7016]_  & \new_[7009]_ ;
  assign \new_[7021]_  = ~A269 & ~A267;
  assign \new_[7022]_  = A235 & \new_[7021]_ ;
  assign \new_[7025]_  = ~A299 & A298;
  assign \new_[7028]_  = A301 & A300;
  assign \new_[7029]_  = \new_[7028]_  & \new_[7025]_ ;
  assign \new_[7030]_  = \new_[7029]_  & \new_[7022]_ ;
  assign \new_[7034]_  = A201 & A200;
  assign \new_[7035]_  = ~A199 & \new_[7034]_ ;
  assign \new_[7038]_  = ~A232 & A202;
  assign \new_[7041]_  = A234 & A233;
  assign \new_[7042]_  = \new_[7041]_  & \new_[7038]_ ;
  assign \new_[7043]_  = \new_[7042]_  & \new_[7035]_ ;
  assign \new_[7047]_  = ~A269 & ~A267;
  assign \new_[7048]_  = A235 & \new_[7047]_ ;
  assign \new_[7051]_  = ~A299 & A298;
  assign \new_[7054]_  = ~A302 & A300;
  assign \new_[7055]_  = \new_[7054]_  & \new_[7051]_ ;
  assign \new_[7056]_  = \new_[7055]_  & \new_[7048]_ ;
  assign \new_[7060]_  = A201 & A200;
  assign \new_[7061]_  = ~A199 & \new_[7060]_ ;
  assign \new_[7064]_  = ~A232 & A202;
  assign \new_[7067]_  = A234 & A233;
  assign \new_[7068]_  = \new_[7067]_  & \new_[7064]_ ;
  assign \new_[7069]_  = \new_[7068]_  & \new_[7061]_ ;
  assign \new_[7073]_  = ~A269 & ~A267;
  assign \new_[7074]_  = A235 & \new_[7073]_ ;
  assign \new_[7077]_  = A299 & ~A298;
  assign \new_[7080]_  = A301 & A300;
  assign \new_[7081]_  = \new_[7080]_  & \new_[7077]_ ;
  assign \new_[7082]_  = \new_[7081]_  & \new_[7074]_ ;
  assign \new_[7086]_  = A201 & A200;
  assign \new_[7087]_  = ~A199 & \new_[7086]_ ;
  assign \new_[7090]_  = ~A232 & A202;
  assign \new_[7093]_  = A234 & A233;
  assign \new_[7094]_  = \new_[7093]_  & \new_[7090]_ ;
  assign \new_[7095]_  = \new_[7094]_  & \new_[7087]_ ;
  assign \new_[7099]_  = ~A269 & ~A267;
  assign \new_[7100]_  = A235 & \new_[7099]_ ;
  assign \new_[7103]_  = A299 & ~A298;
  assign \new_[7106]_  = ~A302 & A300;
  assign \new_[7107]_  = \new_[7106]_  & \new_[7103]_ ;
  assign \new_[7108]_  = \new_[7107]_  & \new_[7100]_ ;
  assign \new_[7112]_  = A201 & A200;
  assign \new_[7113]_  = ~A199 & \new_[7112]_ ;
  assign \new_[7116]_  = ~A232 & A202;
  assign \new_[7119]_  = A234 & A233;
  assign \new_[7120]_  = \new_[7119]_  & \new_[7116]_ ;
  assign \new_[7121]_  = \new_[7120]_  & \new_[7113]_ ;
  assign \new_[7125]_  = A266 & A265;
  assign \new_[7126]_  = A235 & \new_[7125]_ ;
  assign \new_[7129]_  = ~A299 & A298;
  assign \new_[7132]_  = A301 & A300;
  assign \new_[7133]_  = \new_[7132]_  & \new_[7129]_ ;
  assign \new_[7134]_  = \new_[7133]_  & \new_[7126]_ ;
  assign \new_[7138]_  = A201 & A200;
  assign \new_[7139]_  = ~A199 & \new_[7138]_ ;
  assign \new_[7142]_  = ~A232 & A202;
  assign \new_[7145]_  = A234 & A233;
  assign \new_[7146]_  = \new_[7145]_  & \new_[7142]_ ;
  assign \new_[7147]_  = \new_[7146]_  & \new_[7139]_ ;
  assign \new_[7151]_  = A266 & A265;
  assign \new_[7152]_  = A235 & \new_[7151]_ ;
  assign \new_[7155]_  = ~A299 & A298;
  assign \new_[7158]_  = ~A302 & A300;
  assign \new_[7159]_  = \new_[7158]_  & \new_[7155]_ ;
  assign \new_[7160]_  = \new_[7159]_  & \new_[7152]_ ;
  assign \new_[7164]_  = A201 & A200;
  assign \new_[7165]_  = ~A199 & \new_[7164]_ ;
  assign \new_[7168]_  = ~A232 & A202;
  assign \new_[7171]_  = A234 & A233;
  assign \new_[7172]_  = \new_[7171]_  & \new_[7168]_ ;
  assign \new_[7173]_  = \new_[7172]_  & \new_[7165]_ ;
  assign \new_[7177]_  = A266 & A265;
  assign \new_[7178]_  = A235 & \new_[7177]_ ;
  assign \new_[7181]_  = A299 & ~A298;
  assign \new_[7184]_  = A301 & A300;
  assign \new_[7185]_  = \new_[7184]_  & \new_[7181]_ ;
  assign \new_[7186]_  = \new_[7185]_  & \new_[7178]_ ;
  assign \new_[7190]_  = A201 & A200;
  assign \new_[7191]_  = ~A199 & \new_[7190]_ ;
  assign \new_[7194]_  = ~A232 & A202;
  assign \new_[7197]_  = A234 & A233;
  assign \new_[7198]_  = \new_[7197]_  & \new_[7194]_ ;
  assign \new_[7199]_  = \new_[7198]_  & \new_[7191]_ ;
  assign \new_[7203]_  = A266 & A265;
  assign \new_[7204]_  = A235 & \new_[7203]_ ;
  assign \new_[7207]_  = A299 & ~A298;
  assign \new_[7210]_  = ~A302 & A300;
  assign \new_[7211]_  = \new_[7210]_  & \new_[7207]_ ;
  assign \new_[7212]_  = \new_[7211]_  & \new_[7204]_ ;
  assign \new_[7216]_  = A201 & A200;
  assign \new_[7217]_  = ~A199 & \new_[7216]_ ;
  assign \new_[7220]_  = ~A232 & A202;
  assign \new_[7223]_  = A234 & A233;
  assign \new_[7224]_  = \new_[7223]_  & \new_[7220]_ ;
  assign \new_[7225]_  = \new_[7224]_  & \new_[7217]_ ;
  assign \new_[7229]_  = ~A266 & ~A265;
  assign \new_[7230]_  = A235 & \new_[7229]_ ;
  assign \new_[7233]_  = ~A299 & A298;
  assign \new_[7236]_  = A301 & A300;
  assign \new_[7237]_  = \new_[7236]_  & \new_[7233]_ ;
  assign \new_[7238]_  = \new_[7237]_  & \new_[7230]_ ;
  assign \new_[7242]_  = A201 & A200;
  assign \new_[7243]_  = ~A199 & \new_[7242]_ ;
  assign \new_[7246]_  = ~A232 & A202;
  assign \new_[7249]_  = A234 & A233;
  assign \new_[7250]_  = \new_[7249]_  & \new_[7246]_ ;
  assign \new_[7251]_  = \new_[7250]_  & \new_[7243]_ ;
  assign \new_[7255]_  = ~A266 & ~A265;
  assign \new_[7256]_  = A235 & \new_[7255]_ ;
  assign \new_[7259]_  = ~A299 & A298;
  assign \new_[7262]_  = ~A302 & A300;
  assign \new_[7263]_  = \new_[7262]_  & \new_[7259]_ ;
  assign \new_[7264]_  = \new_[7263]_  & \new_[7256]_ ;
  assign \new_[7268]_  = A201 & A200;
  assign \new_[7269]_  = ~A199 & \new_[7268]_ ;
  assign \new_[7272]_  = ~A232 & A202;
  assign \new_[7275]_  = A234 & A233;
  assign \new_[7276]_  = \new_[7275]_  & \new_[7272]_ ;
  assign \new_[7277]_  = \new_[7276]_  & \new_[7269]_ ;
  assign \new_[7281]_  = ~A266 & ~A265;
  assign \new_[7282]_  = A235 & \new_[7281]_ ;
  assign \new_[7285]_  = A299 & ~A298;
  assign \new_[7288]_  = A301 & A300;
  assign \new_[7289]_  = \new_[7288]_  & \new_[7285]_ ;
  assign \new_[7290]_  = \new_[7289]_  & \new_[7282]_ ;
  assign \new_[7294]_  = A201 & A200;
  assign \new_[7295]_  = ~A199 & \new_[7294]_ ;
  assign \new_[7298]_  = ~A232 & A202;
  assign \new_[7301]_  = A234 & A233;
  assign \new_[7302]_  = \new_[7301]_  & \new_[7298]_ ;
  assign \new_[7303]_  = \new_[7302]_  & \new_[7295]_ ;
  assign \new_[7307]_  = ~A266 & ~A265;
  assign \new_[7308]_  = A235 & \new_[7307]_ ;
  assign \new_[7311]_  = A299 & ~A298;
  assign \new_[7314]_  = ~A302 & A300;
  assign \new_[7315]_  = \new_[7314]_  & \new_[7311]_ ;
  assign \new_[7316]_  = \new_[7315]_  & \new_[7308]_ ;
  assign \new_[7320]_  = A201 & A200;
  assign \new_[7321]_  = ~A199 & \new_[7320]_ ;
  assign \new_[7324]_  = ~A232 & A202;
  assign \new_[7327]_  = A234 & A233;
  assign \new_[7328]_  = \new_[7327]_  & \new_[7324]_ ;
  assign \new_[7329]_  = \new_[7328]_  & \new_[7321]_ ;
  assign \new_[7333]_  = A268 & ~A267;
  assign \new_[7334]_  = ~A236 & \new_[7333]_ ;
  assign \new_[7337]_  = ~A299 & A298;
  assign \new_[7340]_  = A301 & A300;
  assign \new_[7341]_  = \new_[7340]_  & \new_[7337]_ ;
  assign \new_[7342]_  = \new_[7341]_  & \new_[7334]_ ;
  assign \new_[7346]_  = A201 & A200;
  assign \new_[7347]_  = ~A199 & \new_[7346]_ ;
  assign \new_[7350]_  = ~A232 & A202;
  assign \new_[7353]_  = A234 & A233;
  assign \new_[7354]_  = \new_[7353]_  & \new_[7350]_ ;
  assign \new_[7355]_  = \new_[7354]_  & \new_[7347]_ ;
  assign \new_[7359]_  = A268 & ~A267;
  assign \new_[7360]_  = ~A236 & \new_[7359]_ ;
  assign \new_[7363]_  = ~A299 & A298;
  assign \new_[7366]_  = ~A302 & A300;
  assign \new_[7367]_  = \new_[7366]_  & \new_[7363]_ ;
  assign \new_[7368]_  = \new_[7367]_  & \new_[7360]_ ;
  assign \new_[7372]_  = A201 & A200;
  assign \new_[7373]_  = ~A199 & \new_[7372]_ ;
  assign \new_[7376]_  = ~A232 & A202;
  assign \new_[7379]_  = A234 & A233;
  assign \new_[7380]_  = \new_[7379]_  & \new_[7376]_ ;
  assign \new_[7381]_  = \new_[7380]_  & \new_[7373]_ ;
  assign \new_[7385]_  = A268 & ~A267;
  assign \new_[7386]_  = ~A236 & \new_[7385]_ ;
  assign \new_[7389]_  = A299 & ~A298;
  assign \new_[7392]_  = A301 & A300;
  assign \new_[7393]_  = \new_[7392]_  & \new_[7389]_ ;
  assign \new_[7394]_  = \new_[7393]_  & \new_[7386]_ ;
  assign \new_[7398]_  = A201 & A200;
  assign \new_[7399]_  = ~A199 & \new_[7398]_ ;
  assign \new_[7402]_  = ~A232 & A202;
  assign \new_[7405]_  = A234 & A233;
  assign \new_[7406]_  = \new_[7405]_  & \new_[7402]_ ;
  assign \new_[7407]_  = \new_[7406]_  & \new_[7399]_ ;
  assign \new_[7411]_  = A268 & ~A267;
  assign \new_[7412]_  = ~A236 & \new_[7411]_ ;
  assign \new_[7415]_  = A299 & ~A298;
  assign \new_[7418]_  = ~A302 & A300;
  assign \new_[7419]_  = \new_[7418]_  & \new_[7415]_ ;
  assign \new_[7420]_  = \new_[7419]_  & \new_[7412]_ ;
  assign \new_[7424]_  = A201 & A200;
  assign \new_[7425]_  = ~A199 & \new_[7424]_ ;
  assign \new_[7428]_  = ~A232 & A202;
  assign \new_[7431]_  = A234 & A233;
  assign \new_[7432]_  = \new_[7431]_  & \new_[7428]_ ;
  assign \new_[7433]_  = \new_[7432]_  & \new_[7425]_ ;
  assign \new_[7437]_  = ~A269 & ~A267;
  assign \new_[7438]_  = ~A236 & \new_[7437]_ ;
  assign \new_[7441]_  = ~A299 & A298;
  assign \new_[7444]_  = A301 & A300;
  assign \new_[7445]_  = \new_[7444]_  & \new_[7441]_ ;
  assign \new_[7446]_  = \new_[7445]_  & \new_[7438]_ ;
  assign \new_[7450]_  = A201 & A200;
  assign \new_[7451]_  = ~A199 & \new_[7450]_ ;
  assign \new_[7454]_  = ~A232 & A202;
  assign \new_[7457]_  = A234 & A233;
  assign \new_[7458]_  = \new_[7457]_  & \new_[7454]_ ;
  assign \new_[7459]_  = \new_[7458]_  & \new_[7451]_ ;
  assign \new_[7463]_  = ~A269 & ~A267;
  assign \new_[7464]_  = ~A236 & \new_[7463]_ ;
  assign \new_[7467]_  = ~A299 & A298;
  assign \new_[7470]_  = ~A302 & A300;
  assign \new_[7471]_  = \new_[7470]_  & \new_[7467]_ ;
  assign \new_[7472]_  = \new_[7471]_  & \new_[7464]_ ;
  assign \new_[7476]_  = A201 & A200;
  assign \new_[7477]_  = ~A199 & \new_[7476]_ ;
  assign \new_[7480]_  = ~A232 & A202;
  assign \new_[7483]_  = A234 & A233;
  assign \new_[7484]_  = \new_[7483]_  & \new_[7480]_ ;
  assign \new_[7485]_  = \new_[7484]_  & \new_[7477]_ ;
  assign \new_[7489]_  = ~A269 & ~A267;
  assign \new_[7490]_  = ~A236 & \new_[7489]_ ;
  assign \new_[7493]_  = A299 & ~A298;
  assign \new_[7496]_  = A301 & A300;
  assign \new_[7497]_  = \new_[7496]_  & \new_[7493]_ ;
  assign \new_[7498]_  = \new_[7497]_  & \new_[7490]_ ;
  assign \new_[7502]_  = A201 & A200;
  assign \new_[7503]_  = ~A199 & \new_[7502]_ ;
  assign \new_[7506]_  = ~A232 & A202;
  assign \new_[7509]_  = A234 & A233;
  assign \new_[7510]_  = \new_[7509]_  & \new_[7506]_ ;
  assign \new_[7511]_  = \new_[7510]_  & \new_[7503]_ ;
  assign \new_[7515]_  = ~A269 & ~A267;
  assign \new_[7516]_  = ~A236 & \new_[7515]_ ;
  assign \new_[7519]_  = A299 & ~A298;
  assign \new_[7522]_  = ~A302 & A300;
  assign \new_[7523]_  = \new_[7522]_  & \new_[7519]_ ;
  assign \new_[7524]_  = \new_[7523]_  & \new_[7516]_ ;
  assign \new_[7528]_  = A201 & A200;
  assign \new_[7529]_  = ~A199 & \new_[7528]_ ;
  assign \new_[7532]_  = ~A232 & A202;
  assign \new_[7535]_  = A234 & A233;
  assign \new_[7536]_  = \new_[7535]_  & \new_[7532]_ ;
  assign \new_[7537]_  = \new_[7536]_  & \new_[7529]_ ;
  assign \new_[7541]_  = A266 & A265;
  assign \new_[7542]_  = ~A236 & \new_[7541]_ ;
  assign \new_[7545]_  = ~A299 & A298;
  assign \new_[7548]_  = A301 & A300;
  assign \new_[7549]_  = \new_[7548]_  & \new_[7545]_ ;
  assign \new_[7550]_  = \new_[7549]_  & \new_[7542]_ ;
  assign \new_[7554]_  = A201 & A200;
  assign \new_[7555]_  = ~A199 & \new_[7554]_ ;
  assign \new_[7558]_  = ~A232 & A202;
  assign \new_[7561]_  = A234 & A233;
  assign \new_[7562]_  = \new_[7561]_  & \new_[7558]_ ;
  assign \new_[7563]_  = \new_[7562]_  & \new_[7555]_ ;
  assign \new_[7567]_  = A266 & A265;
  assign \new_[7568]_  = ~A236 & \new_[7567]_ ;
  assign \new_[7571]_  = ~A299 & A298;
  assign \new_[7574]_  = ~A302 & A300;
  assign \new_[7575]_  = \new_[7574]_  & \new_[7571]_ ;
  assign \new_[7576]_  = \new_[7575]_  & \new_[7568]_ ;
  assign \new_[7580]_  = A201 & A200;
  assign \new_[7581]_  = ~A199 & \new_[7580]_ ;
  assign \new_[7584]_  = ~A232 & A202;
  assign \new_[7587]_  = A234 & A233;
  assign \new_[7588]_  = \new_[7587]_  & \new_[7584]_ ;
  assign \new_[7589]_  = \new_[7588]_  & \new_[7581]_ ;
  assign \new_[7593]_  = A266 & A265;
  assign \new_[7594]_  = ~A236 & \new_[7593]_ ;
  assign \new_[7597]_  = A299 & ~A298;
  assign \new_[7600]_  = A301 & A300;
  assign \new_[7601]_  = \new_[7600]_  & \new_[7597]_ ;
  assign \new_[7602]_  = \new_[7601]_  & \new_[7594]_ ;
  assign \new_[7606]_  = A201 & A200;
  assign \new_[7607]_  = ~A199 & \new_[7606]_ ;
  assign \new_[7610]_  = ~A232 & A202;
  assign \new_[7613]_  = A234 & A233;
  assign \new_[7614]_  = \new_[7613]_  & \new_[7610]_ ;
  assign \new_[7615]_  = \new_[7614]_  & \new_[7607]_ ;
  assign \new_[7619]_  = A266 & A265;
  assign \new_[7620]_  = ~A236 & \new_[7619]_ ;
  assign \new_[7623]_  = A299 & ~A298;
  assign \new_[7626]_  = ~A302 & A300;
  assign \new_[7627]_  = \new_[7626]_  & \new_[7623]_ ;
  assign \new_[7628]_  = \new_[7627]_  & \new_[7620]_ ;
  assign \new_[7632]_  = A201 & A200;
  assign \new_[7633]_  = ~A199 & \new_[7632]_ ;
  assign \new_[7636]_  = ~A232 & A202;
  assign \new_[7639]_  = A234 & A233;
  assign \new_[7640]_  = \new_[7639]_  & \new_[7636]_ ;
  assign \new_[7641]_  = \new_[7640]_  & \new_[7633]_ ;
  assign \new_[7645]_  = ~A266 & ~A265;
  assign \new_[7646]_  = ~A236 & \new_[7645]_ ;
  assign \new_[7649]_  = ~A299 & A298;
  assign \new_[7652]_  = A301 & A300;
  assign \new_[7653]_  = \new_[7652]_  & \new_[7649]_ ;
  assign \new_[7654]_  = \new_[7653]_  & \new_[7646]_ ;
  assign \new_[7658]_  = A201 & A200;
  assign \new_[7659]_  = ~A199 & \new_[7658]_ ;
  assign \new_[7662]_  = ~A232 & A202;
  assign \new_[7665]_  = A234 & A233;
  assign \new_[7666]_  = \new_[7665]_  & \new_[7662]_ ;
  assign \new_[7667]_  = \new_[7666]_  & \new_[7659]_ ;
  assign \new_[7671]_  = ~A266 & ~A265;
  assign \new_[7672]_  = ~A236 & \new_[7671]_ ;
  assign \new_[7675]_  = ~A299 & A298;
  assign \new_[7678]_  = ~A302 & A300;
  assign \new_[7679]_  = \new_[7678]_  & \new_[7675]_ ;
  assign \new_[7680]_  = \new_[7679]_  & \new_[7672]_ ;
  assign \new_[7684]_  = A201 & A200;
  assign \new_[7685]_  = ~A199 & \new_[7684]_ ;
  assign \new_[7688]_  = ~A232 & A202;
  assign \new_[7691]_  = A234 & A233;
  assign \new_[7692]_  = \new_[7691]_  & \new_[7688]_ ;
  assign \new_[7693]_  = \new_[7692]_  & \new_[7685]_ ;
  assign \new_[7697]_  = ~A266 & ~A265;
  assign \new_[7698]_  = ~A236 & \new_[7697]_ ;
  assign \new_[7701]_  = A299 & ~A298;
  assign \new_[7704]_  = A301 & A300;
  assign \new_[7705]_  = \new_[7704]_  & \new_[7701]_ ;
  assign \new_[7706]_  = \new_[7705]_  & \new_[7698]_ ;
  assign \new_[7710]_  = A201 & A200;
  assign \new_[7711]_  = ~A199 & \new_[7710]_ ;
  assign \new_[7714]_  = ~A232 & A202;
  assign \new_[7717]_  = A234 & A233;
  assign \new_[7718]_  = \new_[7717]_  & \new_[7714]_ ;
  assign \new_[7719]_  = \new_[7718]_  & \new_[7711]_ ;
  assign \new_[7723]_  = ~A266 & ~A265;
  assign \new_[7724]_  = ~A236 & \new_[7723]_ ;
  assign \new_[7727]_  = A299 & ~A298;
  assign \new_[7730]_  = ~A302 & A300;
  assign \new_[7731]_  = \new_[7730]_  & \new_[7727]_ ;
  assign \new_[7732]_  = \new_[7731]_  & \new_[7724]_ ;
  assign \new_[7736]_  = A201 & A200;
  assign \new_[7737]_  = ~A199 & \new_[7736]_ ;
  assign \new_[7740]_  = A232 & A202;
  assign \new_[7743]_  = A234 & ~A233;
  assign \new_[7744]_  = \new_[7743]_  & \new_[7740]_ ;
  assign \new_[7745]_  = \new_[7744]_  & \new_[7737]_ ;
  assign \new_[7749]_  = A268 & ~A267;
  assign \new_[7750]_  = A235 & \new_[7749]_ ;
  assign \new_[7753]_  = ~A299 & A298;
  assign \new_[7756]_  = A301 & A300;
  assign \new_[7757]_  = \new_[7756]_  & \new_[7753]_ ;
  assign \new_[7758]_  = \new_[7757]_  & \new_[7750]_ ;
  assign \new_[7762]_  = A201 & A200;
  assign \new_[7763]_  = ~A199 & \new_[7762]_ ;
  assign \new_[7766]_  = A232 & A202;
  assign \new_[7769]_  = A234 & ~A233;
  assign \new_[7770]_  = \new_[7769]_  & \new_[7766]_ ;
  assign \new_[7771]_  = \new_[7770]_  & \new_[7763]_ ;
  assign \new_[7775]_  = A268 & ~A267;
  assign \new_[7776]_  = A235 & \new_[7775]_ ;
  assign \new_[7779]_  = ~A299 & A298;
  assign \new_[7782]_  = ~A302 & A300;
  assign \new_[7783]_  = \new_[7782]_  & \new_[7779]_ ;
  assign \new_[7784]_  = \new_[7783]_  & \new_[7776]_ ;
  assign \new_[7788]_  = A201 & A200;
  assign \new_[7789]_  = ~A199 & \new_[7788]_ ;
  assign \new_[7792]_  = A232 & A202;
  assign \new_[7795]_  = A234 & ~A233;
  assign \new_[7796]_  = \new_[7795]_  & \new_[7792]_ ;
  assign \new_[7797]_  = \new_[7796]_  & \new_[7789]_ ;
  assign \new_[7801]_  = A268 & ~A267;
  assign \new_[7802]_  = A235 & \new_[7801]_ ;
  assign \new_[7805]_  = A299 & ~A298;
  assign \new_[7808]_  = A301 & A300;
  assign \new_[7809]_  = \new_[7808]_  & \new_[7805]_ ;
  assign \new_[7810]_  = \new_[7809]_  & \new_[7802]_ ;
  assign \new_[7814]_  = A201 & A200;
  assign \new_[7815]_  = ~A199 & \new_[7814]_ ;
  assign \new_[7818]_  = A232 & A202;
  assign \new_[7821]_  = A234 & ~A233;
  assign \new_[7822]_  = \new_[7821]_  & \new_[7818]_ ;
  assign \new_[7823]_  = \new_[7822]_  & \new_[7815]_ ;
  assign \new_[7827]_  = A268 & ~A267;
  assign \new_[7828]_  = A235 & \new_[7827]_ ;
  assign \new_[7831]_  = A299 & ~A298;
  assign \new_[7834]_  = ~A302 & A300;
  assign \new_[7835]_  = \new_[7834]_  & \new_[7831]_ ;
  assign \new_[7836]_  = \new_[7835]_  & \new_[7828]_ ;
  assign \new_[7840]_  = A201 & A200;
  assign \new_[7841]_  = ~A199 & \new_[7840]_ ;
  assign \new_[7844]_  = A232 & A202;
  assign \new_[7847]_  = A234 & ~A233;
  assign \new_[7848]_  = \new_[7847]_  & \new_[7844]_ ;
  assign \new_[7849]_  = \new_[7848]_  & \new_[7841]_ ;
  assign \new_[7853]_  = ~A269 & ~A267;
  assign \new_[7854]_  = A235 & \new_[7853]_ ;
  assign \new_[7857]_  = ~A299 & A298;
  assign \new_[7860]_  = A301 & A300;
  assign \new_[7861]_  = \new_[7860]_  & \new_[7857]_ ;
  assign \new_[7862]_  = \new_[7861]_  & \new_[7854]_ ;
  assign \new_[7866]_  = A201 & A200;
  assign \new_[7867]_  = ~A199 & \new_[7866]_ ;
  assign \new_[7870]_  = A232 & A202;
  assign \new_[7873]_  = A234 & ~A233;
  assign \new_[7874]_  = \new_[7873]_  & \new_[7870]_ ;
  assign \new_[7875]_  = \new_[7874]_  & \new_[7867]_ ;
  assign \new_[7879]_  = ~A269 & ~A267;
  assign \new_[7880]_  = A235 & \new_[7879]_ ;
  assign \new_[7883]_  = ~A299 & A298;
  assign \new_[7886]_  = ~A302 & A300;
  assign \new_[7887]_  = \new_[7886]_  & \new_[7883]_ ;
  assign \new_[7888]_  = \new_[7887]_  & \new_[7880]_ ;
  assign \new_[7892]_  = A201 & A200;
  assign \new_[7893]_  = ~A199 & \new_[7892]_ ;
  assign \new_[7896]_  = A232 & A202;
  assign \new_[7899]_  = A234 & ~A233;
  assign \new_[7900]_  = \new_[7899]_  & \new_[7896]_ ;
  assign \new_[7901]_  = \new_[7900]_  & \new_[7893]_ ;
  assign \new_[7905]_  = ~A269 & ~A267;
  assign \new_[7906]_  = A235 & \new_[7905]_ ;
  assign \new_[7909]_  = A299 & ~A298;
  assign \new_[7912]_  = A301 & A300;
  assign \new_[7913]_  = \new_[7912]_  & \new_[7909]_ ;
  assign \new_[7914]_  = \new_[7913]_  & \new_[7906]_ ;
  assign \new_[7918]_  = A201 & A200;
  assign \new_[7919]_  = ~A199 & \new_[7918]_ ;
  assign \new_[7922]_  = A232 & A202;
  assign \new_[7925]_  = A234 & ~A233;
  assign \new_[7926]_  = \new_[7925]_  & \new_[7922]_ ;
  assign \new_[7927]_  = \new_[7926]_  & \new_[7919]_ ;
  assign \new_[7931]_  = ~A269 & ~A267;
  assign \new_[7932]_  = A235 & \new_[7931]_ ;
  assign \new_[7935]_  = A299 & ~A298;
  assign \new_[7938]_  = ~A302 & A300;
  assign \new_[7939]_  = \new_[7938]_  & \new_[7935]_ ;
  assign \new_[7940]_  = \new_[7939]_  & \new_[7932]_ ;
  assign \new_[7944]_  = A201 & A200;
  assign \new_[7945]_  = ~A199 & \new_[7944]_ ;
  assign \new_[7948]_  = A232 & A202;
  assign \new_[7951]_  = A234 & ~A233;
  assign \new_[7952]_  = \new_[7951]_  & \new_[7948]_ ;
  assign \new_[7953]_  = \new_[7952]_  & \new_[7945]_ ;
  assign \new_[7957]_  = A266 & A265;
  assign \new_[7958]_  = A235 & \new_[7957]_ ;
  assign \new_[7961]_  = ~A299 & A298;
  assign \new_[7964]_  = A301 & A300;
  assign \new_[7965]_  = \new_[7964]_  & \new_[7961]_ ;
  assign \new_[7966]_  = \new_[7965]_  & \new_[7958]_ ;
  assign \new_[7970]_  = A201 & A200;
  assign \new_[7971]_  = ~A199 & \new_[7970]_ ;
  assign \new_[7974]_  = A232 & A202;
  assign \new_[7977]_  = A234 & ~A233;
  assign \new_[7978]_  = \new_[7977]_  & \new_[7974]_ ;
  assign \new_[7979]_  = \new_[7978]_  & \new_[7971]_ ;
  assign \new_[7983]_  = A266 & A265;
  assign \new_[7984]_  = A235 & \new_[7983]_ ;
  assign \new_[7987]_  = ~A299 & A298;
  assign \new_[7990]_  = ~A302 & A300;
  assign \new_[7991]_  = \new_[7990]_  & \new_[7987]_ ;
  assign \new_[7992]_  = \new_[7991]_  & \new_[7984]_ ;
  assign \new_[7996]_  = A201 & A200;
  assign \new_[7997]_  = ~A199 & \new_[7996]_ ;
  assign \new_[8000]_  = A232 & A202;
  assign \new_[8003]_  = A234 & ~A233;
  assign \new_[8004]_  = \new_[8003]_  & \new_[8000]_ ;
  assign \new_[8005]_  = \new_[8004]_  & \new_[7997]_ ;
  assign \new_[8009]_  = A266 & A265;
  assign \new_[8010]_  = A235 & \new_[8009]_ ;
  assign \new_[8013]_  = A299 & ~A298;
  assign \new_[8016]_  = A301 & A300;
  assign \new_[8017]_  = \new_[8016]_  & \new_[8013]_ ;
  assign \new_[8018]_  = \new_[8017]_  & \new_[8010]_ ;
  assign \new_[8022]_  = A201 & A200;
  assign \new_[8023]_  = ~A199 & \new_[8022]_ ;
  assign \new_[8026]_  = A232 & A202;
  assign \new_[8029]_  = A234 & ~A233;
  assign \new_[8030]_  = \new_[8029]_  & \new_[8026]_ ;
  assign \new_[8031]_  = \new_[8030]_  & \new_[8023]_ ;
  assign \new_[8035]_  = A266 & A265;
  assign \new_[8036]_  = A235 & \new_[8035]_ ;
  assign \new_[8039]_  = A299 & ~A298;
  assign \new_[8042]_  = ~A302 & A300;
  assign \new_[8043]_  = \new_[8042]_  & \new_[8039]_ ;
  assign \new_[8044]_  = \new_[8043]_  & \new_[8036]_ ;
  assign \new_[8048]_  = A201 & A200;
  assign \new_[8049]_  = ~A199 & \new_[8048]_ ;
  assign \new_[8052]_  = A232 & A202;
  assign \new_[8055]_  = A234 & ~A233;
  assign \new_[8056]_  = \new_[8055]_  & \new_[8052]_ ;
  assign \new_[8057]_  = \new_[8056]_  & \new_[8049]_ ;
  assign \new_[8061]_  = ~A266 & ~A265;
  assign \new_[8062]_  = A235 & \new_[8061]_ ;
  assign \new_[8065]_  = ~A299 & A298;
  assign \new_[8068]_  = A301 & A300;
  assign \new_[8069]_  = \new_[8068]_  & \new_[8065]_ ;
  assign \new_[8070]_  = \new_[8069]_  & \new_[8062]_ ;
  assign \new_[8074]_  = A201 & A200;
  assign \new_[8075]_  = ~A199 & \new_[8074]_ ;
  assign \new_[8078]_  = A232 & A202;
  assign \new_[8081]_  = A234 & ~A233;
  assign \new_[8082]_  = \new_[8081]_  & \new_[8078]_ ;
  assign \new_[8083]_  = \new_[8082]_  & \new_[8075]_ ;
  assign \new_[8087]_  = ~A266 & ~A265;
  assign \new_[8088]_  = A235 & \new_[8087]_ ;
  assign \new_[8091]_  = ~A299 & A298;
  assign \new_[8094]_  = ~A302 & A300;
  assign \new_[8095]_  = \new_[8094]_  & \new_[8091]_ ;
  assign \new_[8096]_  = \new_[8095]_  & \new_[8088]_ ;
  assign \new_[8100]_  = A201 & A200;
  assign \new_[8101]_  = ~A199 & \new_[8100]_ ;
  assign \new_[8104]_  = A232 & A202;
  assign \new_[8107]_  = A234 & ~A233;
  assign \new_[8108]_  = \new_[8107]_  & \new_[8104]_ ;
  assign \new_[8109]_  = \new_[8108]_  & \new_[8101]_ ;
  assign \new_[8113]_  = ~A266 & ~A265;
  assign \new_[8114]_  = A235 & \new_[8113]_ ;
  assign \new_[8117]_  = A299 & ~A298;
  assign \new_[8120]_  = A301 & A300;
  assign \new_[8121]_  = \new_[8120]_  & \new_[8117]_ ;
  assign \new_[8122]_  = \new_[8121]_  & \new_[8114]_ ;
  assign \new_[8126]_  = A201 & A200;
  assign \new_[8127]_  = ~A199 & \new_[8126]_ ;
  assign \new_[8130]_  = A232 & A202;
  assign \new_[8133]_  = A234 & ~A233;
  assign \new_[8134]_  = \new_[8133]_  & \new_[8130]_ ;
  assign \new_[8135]_  = \new_[8134]_  & \new_[8127]_ ;
  assign \new_[8139]_  = ~A266 & ~A265;
  assign \new_[8140]_  = A235 & \new_[8139]_ ;
  assign \new_[8143]_  = A299 & ~A298;
  assign \new_[8146]_  = ~A302 & A300;
  assign \new_[8147]_  = \new_[8146]_  & \new_[8143]_ ;
  assign \new_[8148]_  = \new_[8147]_  & \new_[8140]_ ;
  assign \new_[8152]_  = A201 & A200;
  assign \new_[8153]_  = ~A199 & \new_[8152]_ ;
  assign \new_[8156]_  = A232 & A202;
  assign \new_[8159]_  = A234 & ~A233;
  assign \new_[8160]_  = \new_[8159]_  & \new_[8156]_ ;
  assign \new_[8161]_  = \new_[8160]_  & \new_[8153]_ ;
  assign \new_[8165]_  = A268 & ~A267;
  assign \new_[8166]_  = ~A236 & \new_[8165]_ ;
  assign \new_[8169]_  = ~A299 & A298;
  assign \new_[8172]_  = A301 & A300;
  assign \new_[8173]_  = \new_[8172]_  & \new_[8169]_ ;
  assign \new_[8174]_  = \new_[8173]_  & \new_[8166]_ ;
  assign \new_[8178]_  = A201 & A200;
  assign \new_[8179]_  = ~A199 & \new_[8178]_ ;
  assign \new_[8182]_  = A232 & A202;
  assign \new_[8185]_  = A234 & ~A233;
  assign \new_[8186]_  = \new_[8185]_  & \new_[8182]_ ;
  assign \new_[8187]_  = \new_[8186]_  & \new_[8179]_ ;
  assign \new_[8191]_  = A268 & ~A267;
  assign \new_[8192]_  = ~A236 & \new_[8191]_ ;
  assign \new_[8195]_  = ~A299 & A298;
  assign \new_[8198]_  = ~A302 & A300;
  assign \new_[8199]_  = \new_[8198]_  & \new_[8195]_ ;
  assign \new_[8200]_  = \new_[8199]_  & \new_[8192]_ ;
  assign \new_[8204]_  = A201 & A200;
  assign \new_[8205]_  = ~A199 & \new_[8204]_ ;
  assign \new_[8208]_  = A232 & A202;
  assign \new_[8211]_  = A234 & ~A233;
  assign \new_[8212]_  = \new_[8211]_  & \new_[8208]_ ;
  assign \new_[8213]_  = \new_[8212]_  & \new_[8205]_ ;
  assign \new_[8217]_  = A268 & ~A267;
  assign \new_[8218]_  = ~A236 & \new_[8217]_ ;
  assign \new_[8221]_  = A299 & ~A298;
  assign \new_[8224]_  = A301 & A300;
  assign \new_[8225]_  = \new_[8224]_  & \new_[8221]_ ;
  assign \new_[8226]_  = \new_[8225]_  & \new_[8218]_ ;
  assign \new_[8230]_  = A201 & A200;
  assign \new_[8231]_  = ~A199 & \new_[8230]_ ;
  assign \new_[8234]_  = A232 & A202;
  assign \new_[8237]_  = A234 & ~A233;
  assign \new_[8238]_  = \new_[8237]_  & \new_[8234]_ ;
  assign \new_[8239]_  = \new_[8238]_  & \new_[8231]_ ;
  assign \new_[8243]_  = A268 & ~A267;
  assign \new_[8244]_  = ~A236 & \new_[8243]_ ;
  assign \new_[8247]_  = A299 & ~A298;
  assign \new_[8250]_  = ~A302 & A300;
  assign \new_[8251]_  = \new_[8250]_  & \new_[8247]_ ;
  assign \new_[8252]_  = \new_[8251]_  & \new_[8244]_ ;
  assign \new_[8256]_  = A201 & A200;
  assign \new_[8257]_  = ~A199 & \new_[8256]_ ;
  assign \new_[8260]_  = A232 & A202;
  assign \new_[8263]_  = A234 & ~A233;
  assign \new_[8264]_  = \new_[8263]_  & \new_[8260]_ ;
  assign \new_[8265]_  = \new_[8264]_  & \new_[8257]_ ;
  assign \new_[8269]_  = ~A269 & ~A267;
  assign \new_[8270]_  = ~A236 & \new_[8269]_ ;
  assign \new_[8273]_  = ~A299 & A298;
  assign \new_[8276]_  = A301 & A300;
  assign \new_[8277]_  = \new_[8276]_  & \new_[8273]_ ;
  assign \new_[8278]_  = \new_[8277]_  & \new_[8270]_ ;
  assign \new_[8282]_  = A201 & A200;
  assign \new_[8283]_  = ~A199 & \new_[8282]_ ;
  assign \new_[8286]_  = A232 & A202;
  assign \new_[8289]_  = A234 & ~A233;
  assign \new_[8290]_  = \new_[8289]_  & \new_[8286]_ ;
  assign \new_[8291]_  = \new_[8290]_  & \new_[8283]_ ;
  assign \new_[8295]_  = ~A269 & ~A267;
  assign \new_[8296]_  = ~A236 & \new_[8295]_ ;
  assign \new_[8299]_  = ~A299 & A298;
  assign \new_[8302]_  = ~A302 & A300;
  assign \new_[8303]_  = \new_[8302]_  & \new_[8299]_ ;
  assign \new_[8304]_  = \new_[8303]_  & \new_[8296]_ ;
  assign \new_[8308]_  = A201 & A200;
  assign \new_[8309]_  = ~A199 & \new_[8308]_ ;
  assign \new_[8312]_  = A232 & A202;
  assign \new_[8315]_  = A234 & ~A233;
  assign \new_[8316]_  = \new_[8315]_  & \new_[8312]_ ;
  assign \new_[8317]_  = \new_[8316]_  & \new_[8309]_ ;
  assign \new_[8321]_  = ~A269 & ~A267;
  assign \new_[8322]_  = ~A236 & \new_[8321]_ ;
  assign \new_[8325]_  = A299 & ~A298;
  assign \new_[8328]_  = A301 & A300;
  assign \new_[8329]_  = \new_[8328]_  & \new_[8325]_ ;
  assign \new_[8330]_  = \new_[8329]_  & \new_[8322]_ ;
  assign \new_[8334]_  = A201 & A200;
  assign \new_[8335]_  = ~A199 & \new_[8334]_ ;
  assign \new_[8338]_  = A232 & A202;
  assign \new_[8341]_  = A234 & ~A233;
  assign \new_[8342]_  = \new_[8341]_  & \new_[8338]_ ;
  assign \new_[8343]_  = \new_[8342]_  & \new_[8335]_ ;
  assign \new_[8347]_  = ~A269 & ~A267;
  assign \new_[8348]_  = ~A236 & \new_[8347]_ ;
  assign \new_[8351]_  = A299 & ~A298;
  assign \new_[8354]_  = ~A302 & A300;
  assign \new_[8355]_  = \new_[8354]_  & \new_[8351]_ ;
  assign \new_[8356]_  = \new_[8355]_  & \new_[8348]_ ;
  assign \new_[8360]_  = A201 & A200;
  assign \new_[8361]_  = ~A199 & \new_[8360]_ ;
  assign \new_[8364]_  = A232 & A202;
  assign \new_[8367]_  = A234 & ~A233;
  assign \new_[8368]_  = \new_[8367]_  & \new_[8364]_ ;
  assign \new_[8369]_  = \new_[8368]_  & \new_[8361]_ ;
  assign \new_[8373]_  = A266 & A265;
  assign \new_[8374]_  = ~A236 & \new_[8373]_ ;
  assign \new_[8377]_  = ~A299 & A298;
  assign \new_[8380]_  = A301 & A300;
  assign \new_[8381]_  = \new_[8380]_  & \new_[8377]_ ;
  assign \new_[8382]_  = \new_[8381]_  & \new_[8374]_ ;
  assign \new_[8386]_  = A201 & A200;
  assign \new_[8387]_  = ~A199 & \new_[8386]_ ;
  assign \new_[8390]_  = A232 & A202;
  assign \new_[8393]_  = A234 & ~A233;
  assign \new_[8394]_  = \new_[8393]_  & \new_[8390]_ ;
  assign \new_[8395]_  = \new_[8394]_  & \new_[8387]_ ;
  assign \new_[8399]_  = A266 & A265;
  assign \new_[8400]_  = ~A236 & \new_[8399]_ ;
  assign \new_[8403]_  = ~A299 & A298;
  assign \new_[8406]_  = ~A302 & A300;
  assign \new_[8407]_  = \new_[8406]_  & \new_[8403]_ ;
  assign \new_[8408]_  = \new_[8407]_  & \new_[8400]_ ;
  assign \new_[8412]_  = A201 & A200;
  assign \new_[8413]_  = ~A199 & \new_[8412]_ ;
  assign \new_[8416]_  = A232 & A202;
  assign \new_[8419]_  = A234 & ~A233;
  assign \new_[8420]_  = \new_[8419]_  & \new_[8416]_ ;
  assign \new_[8421]_  = \new_[8420]_  & \new_[8413]_ ;
  assign \new_[8425]_  = A266 & A265;
  assign \new_[8426]_  = ~A236 & \new_[8425]_ ;
  assign \new_[8429]_  = A299 & ~A298;
  assign \new_[8432]_  = A301 & A300;
  assign \new_[8433]_  = \new_[8432]_  & \new_[8429]_ ;
  assign \new_[8434]_  = \new_[8433]_  & \new_[8426]_ ;
  assign \new_[8438]_  = A201 & A200;
  assign \new_[8439]_  = ~A199 & \new_[8438]_ ;
  assign \new_[8442]_  = A232 & A202;
  assign \new_[8445]_  = A234 & ~A233;
  assign \new_[8446]_  = \new_[8445]_  & \new_[8442]_ ;
  assign \new_[8447]_  = \new_[8446]_  & \new_[8439]_ ;
  assign \new_[8451]_  = A266 & A265;
  assign \new_[8452]_  = ~A236 & \new_[8451]_ ;
  assign \new_[8455]_  = A299 & ~A298;
  assign \new_[8458]_  = ~A302 & A300;
  assign \new_[8459]_  = \new_[8458]_  & \new_[8455]_ ;
  assign \new_[8460]_  = \new_[8459]_  & \new_[8452]_ ;
  assign \new_[8464]_  = A201 & A200;
  assign \new_[8465]_  = ~A199 & \new_[8464]_ ;
  assign \new_[8468]_  = A232 & A202;
  assign \new_[8471]_  = A234 & ~A233;
  assign \new_[8472]_  = \new_[8471]_  & \new_[8468]_ ;
  assign \new_[8473]_  = \new_[8472]_  & \new_[8465]_ ;
  assign \new_[8477]_  = ~A266 & ~A265;
  assign \new_[8478]_  = ~A236 & \new_[8477]_ ;
  assign \new_[8481]_  = ~A299 & A298;
  assign \new_[8484]_  = A301 & A300;
  assign \new_[8485]_  = \new_[8484]_  & \new_[8481]_ ;
  assign \new_[8486]_  = \new_[8485]_  & \new_[8478]_ ;
  assign \new_[8490]_  = A201 & A200;
  assign \new_[8491]_  = ~A199 & \new_[8490]_ ;
  assign \new_[8494]_  = A232 & A202;
  assign \new_[8497]_  = A234 & ~A233;
  assign \new_[8498]_  = \new_[8497]_  & \new_[8494]_ ;
  assign \new_[8499]_  = \new_[8498]_  & \new_[8491]_ ;
  assign \new_[8503]_  = ~A266 & ~A265;
  assign \new_[8504]_  = ~A236 & \new_[8503]_ ;
  assign \new_[8507]_  = ~A299 & A298;
  assign \new_[8510]_  = ~A302 & A300;
  assign \new_[8511]_  = \new_[8510]_  & \new_[8507]_ ;
  assign \new_[8512]_  = \new_[8511]_  & \new_[8504]_ ;
  assign \new_[8516]_  = A201 & A200;
  assign \new_[8517]_  = ~A199 & \new_[8516]_ ;
  assign \new_[8520]_  = A232 & A202;
  assign \new_[8523]_  = A234 & ~A233;
  assign \new_[8524]_  = \new_[8523]_  & \new_[8520]_ ;
  assign \new_[8525]_  = \new_[8524]_  & \new_[8517]_ ;
  assign \new_[8529]_  = ~A266 & ~A265;
  assign \new_[8530]_  = ~A236 & \new_[8529]_ ;
  assign \new_[8533]_  = A299 & ~A298;
  assign \new_[8536]_  = A301 & A300;
  assign \new_[8537]_  = \new_[8536]_  & \new_[8533]_ ;
  assign \new_[8538]_  = \new_[8537]_  & \new_[8530]_ ;
  assign \new_[8542]_  = A201 & A200;
  assign \new_[8543]_  = ~A199 & \new_[8542]_ ;
  assign \new_[8546]_  = A232 & A202;
  assign \new_[8549]_  = A234 & ~A233;
  assign \new_[8550]_  = \new_[8549]_  & \new_[8546]_ ;
  assign \new_[8551]_  = \new_[8550]_  & \new_[8543]_ ;
  assign \new_[8555]_  = ~A266 & ~A265;
  assign \new_[8556]_  = ~A236 & \new_[8555]_ ;
  assign \new_[8559]_  = A299 & ~A298;
  assign \new_[8562]_  = ~A302 & A300;
  assign \new_[8563]_  = \new_[8562]_  & \new_[8559]_ ;
  assign \new_[8564]_  = \new_[8563]_  & \new_[8556]_ ;
  assign \new_[8568]_  = A201 & A200;
  assign \new_[8569]_  = ~A199 & \new_[8568]_ ;
  assign \new_[8572]_  = ~A232 & ~A203;
  assign \new_[8575]_  = A234 & A233;
  assign \new_[8576]_  = \new_[8575]_  & \new_[8572]_ ;
  assign \new_[8577]_  = \new_[8576]_  & \new_[8569]_ ;
  assign \new_[8581]_  = A268 & ~A267;
  assign \new_[8582]_  = A235 & \new_[8581]_ ;
  assign \new_[8585]_  = ~A299 & A298;
  assign \new_[8588]_  = A301 & A300;
  assign \new_[8589]_  = \new_[8588]_  & \new_[8585]_ ;
  assign \new_[8590]_  = \new_[8589]_  & \new_[8582]_ ;
  assign \new_[8594]_  = A201 & A200;
  assign \new_[8595]_  = ~A199 & \new_[8594]_ ;
  assign \new_[8598]_  = ~A232 & ~A203;
  assign \new_[8601]_  = A234 & A233;
  assign \new_[8602]_  = \new_[8601]_  & \new_[8598]_ ;
  assign \new_[8603]_  = \new_[8602]_  & \new_[8595]_ ;
  assign \new_[8607]_  = A268 & ~A267;
  assign \new_[8608]_  = A235 & \new_[8607]_ ;
  assign \new_[8611]_  = ~A299 & A298;
  assign \new_[8614]_  = ~A302 & A300;
  assign \new_[8615]_  = \new_[8614]_  & \new_[8611]_ ;
  assign \new_[8616]_  = \new_[8615]_  & \new_[8608]_ ;
  assign \new_[8620]_  = A201 & A200;
  assign \new_[8621]_  = ~A199 & \new_[8620]_ ;
  assign \new_[8624]_  = ~A232 & ~A203;
  assign \new_[8627]_  = A234 & A233;
  assign \new_[8628]_  = \new_[8627]_  & \new_[8624]_ ;
  assign \new_[8629]_  = \new_[8628]_  & \new_[8621]_ ;
  assign \new_[8633]_  = A268 & ~A267;
  assign \new_[8634]_  = A235 & \new_[8633]_ ;
  assign \new_[8637]_  = A299 & ~A298;
  assign \new_[8640]_  = A301 & A300;
  assign \new_[8641]_  = \new_[8640]_  & \new_[8637]_ ;
  assign \new_[8642]_  = \new_[8641]_  & \new_[8634]_ ;
  assign \new_[8646]_  = A201 & A200;
  assign \new_[8647]_  = ~A199 & \new_[8646]_ ;
  assign \new_[8650]_  = ~A232 & ~A203;
  assign \new_[8653]_  = A234 & A233;
  assign \new_[8654]_  = \new_[8653]_  & \new_[8650]_ ;
  assign \new_[8655]_  = \new_[8654]_  & \new_[8647]_ ;
  assign \new_[8659]_  = A268 & ~A267;
  assign \new_[8660]_  = A235 & \new_[8659]_ ;
  assign \new_[8663]_  = A299 & ~A298;
  assign \new_[8666]_  = ~A302 & A300;
  assign \new_[8667]_  = \new_[8666]_  & \new_[8663]_ ;
  assign \new_[8668]_  = \new_[8667]_  & \new_[8660]_ ;
  assign \new_[8672]_  = A201 & A200;
  assign \new_[8673]_  = ~A199 & \new_[8672]_ ;
  assign \new_[8676]_  = ~A232 & ~A203;
  assign \new_[8679]_  = A234 & A233;
  assign \new_[8680]_  = \new_[8679]_  & \new_[8676]_ ;
  assign \new_[8681]_  = \new_[8680]_  & \new_[8673]_ ;
  assign \new_[8685]_  = ~A269 & ~A267;
  assign \new_[8686]_  = A235 & \new_[8685]_ ;
  assign \new_[8689]_  = ~A299 & A298;
  assign \new_[8692]_  = A301 & A300;
  assign \new_[8693]_  = \new_[8692]_  & \new_[8689]_ ;
  assign \new_[8694]_  = \new_[8693]_  & \new_[8686]_ ;
  assign \new_[8698]_  = A201 & A200;
  assign \new_[8699]_  = ~A199 & \new_[8698]_ ;
  assign \new_[8702]_  = ~A232 & ~A203;
  assign \new_[8705]_  = A234 & A233;
  assign \new_[8706]_  = \new_[8705]_  & \new_[8702]_ ;
  assign \new_[8707]_  = \new_[8706]_  & \new_[8699]_ ;
  assign \new_[8711]_  = ~A269 & ~A267;
  assign \new_[8712]_  = A235 & \new_[8711]_ ;
  assign \new_[8715]_  = ~A299 & A298;
  assign \new_[8718]_  = ~A302 & A300;
  assign \new_[8719]_  = \new_[8718]_  & \new_[8715]_ ;
  assign \new_[8720]_  = \new_[8719]_  & \new_[8712]_ ;
  assign \new_[8724]_  = A201 & A200;
  assign \new_[8725]_  = ~A199 & \new_[8724]_ ;
  assign \new_[8728]_  = ~A232 & ~A203;
  assign \new_[8731]_  = A234 & A233;
  assign \new_[8732]_  = \new_[8731]_  & \new_[8728]_ ;
  assign \new_[8733]_  = \new_[8732]_  & \new_[8725]_ ;
  assign \new_[8737]_  = ~A269 & ~A267;
  assign \new_[8738]_  = A235 & \new_[8737]_ ;
  assign \new_[8741]_  = A299 & ~A298;
  assign \new_[8744]_  = A301 & A300;
  assign \new_[8745]_  = \new_[8744]_  & \new_[8741]_ ;
  assign \new_[8746]_  = \new_[8745]_  & \new_[8738]_ ;
  assign \new_[8750]_  = A201 & A200;
  assign \new_[8751]_  = ~A199 & \new_[8750]_ ;
  assign \new_[8754]_  = ~A232 & ~A203;
  assign \new_[8757]_  = A234 & A233;
  assign \new_[8758]_  = \new_[8757]_  & \new_[8754]_ ;
  assign \new_[8759]_  = \new_[8758]_  & \new_[8751]_ ;
  assign \new_[8763]_  = ~A269 & ~A267;
  assign \new_[8764]_  = A235 & \new_[8763]_ ;
  assign \new_[8767]_  = A299 & ~A298;
  assign \new_[8770]_  = ~A302 & A300;
  assign \new_[8771]_  = \new_[8770]_  & \new_[8767]_ ;
  assign \new_[8772]_  = \new_[8771]_  & \new_[8764]_ ;
  assign \new_[8776]_  = A201 & A200;
  assign \new_[8777]_  = ~A199 & \new_[8776]_ ;
  assign \new_[8780]_  = ~A232 & ~A203;
  assign \new_[8783]_  = A234 & A233;
  assign \new_[8784]_  = \new_[8783]_  & \new_[8780]_ ;
  assign \new_[8785]_  = \new_[8784]_  & \new_[8777]_ ;
  assign \new_[8789]_  = A266 & A265;
  assign \new_[8790]_  = A235 & \new_[8789]_ ;
  assign \new_[8793]_  = ~A299 & A298;
  assign \new_[8796]_  = A301 & A300;
  assign \new_[8797]_  = \new_[8796]_  & \new_[8793]_ ;
  assign \new_[8798]_  = \new_[8797]_  & \new_[8790]_ ;
  assign \new_[8802]_  = A201 & A200;
  assign \new_[8803]_  = ~A199 & \new_[8802]_ ;
  assign \new_[8806]_  = ~A232 & ~A203;
  assign \new_[8809]_  = A234 & A233;
  assign \new_[8810]_  = \new_[8809]_  & \new_[8806]_ ;
  assign \new_[8811]_  = \new_[8810]_  & \new_[8803]_ ;
  assign \new_[8815]_  = A266 & A265;
  assign \new_[8816]_  = A235 & \new_[8815]_ ;
  assign \new_[8819]_  = ~A299 & A298;
  assign \new_[8822]_  = ~A302 & A300;
  assign \new_[8823]_  = \new_[8822]_  & \new_[8819]_ ;
  assign \new_[8824]_  = \new_[8823]_  & \new_[8816]_ ;
  assign \new_[8828]_  = A201 & A200;
  assign \new_[8829]_  = ~A199 & \new_[8828]_ ;
  assign \new_[8832]_  = ~A232 & ~A203;
  assign \new_[8835]_  = A234 & A233;
  assign \new_[8836]_  = \new_[8835]_  & \new_[8832]_ ;
  assign \new_[8837]_  = \new_[8836]_  & \new_[8829]_ ;
  assign \new_[8841]_  = A266 & A265;
  assign \new_[8842]_  = A235 & \new_[8841]_ ;
  assign \new_[8845]_  = A299 & ~A298;
  assign \new_[8848]_  = A301 & A300;
  assign \new_[8849]_  = \new_[8848]_  & \new_[8845]_ ;
  assign \new_[8850]_  = \new_[8849]_  & \new_[8842]_ ;
  assign \new_[8854]_  = A201 & A200;
  assign \new_[8855]_  = ~A199 & \new_[8854]_ ;
  assign \new_[8858]_  = ~A232 & ~A203;
  assign \new_[8861]_  = A234 & A233;
  assign \new_[8862]_  = \new_[8861]_  & \new_[8858]_ ;
  assign \new_[8863]_  = \new_[8862]_  & \new_[8855]_ ;
  assign \new_[8867]_  = A266 & A265;
  assign \new_[8868]_  = A235 & \new_[8867]_ ;
  assign \new_[8871]_  = A299 & ~A298;
  assign \new_[8874]_  = ~A302 & A300;
  assign \new_[8875]_  = \new_[8874]_  & \new_[8871]_ ;
  assign \new_[8876]_  = \new_[8875]_  & \new_[8868]_ ;
  assign \new_[8880]_  = A201 & A200;
  assign \new_[8881]_  = ~A199 & \new_[8880]_ ;
  assign \new_[8884]_  = ~A232 & ~A203;
  assign \new_[8887]_  = A234 & A233;
  assign \new_[8888]_  = \new_[8887]_  & \new_[8884]_ ;
  assign \new_[8889]_  = \new_[8888]_  & \new_[8881]_ ;
  assign \new_[8893]_  = ~A266 & ~A265;
  assign \new_[8894]_  = A235 & \new_[8893]_ ;
  assign \new_[8897]_  = ~A299 & A298;
  assign \new_[8900]_  = A301 & A300;
  assign \new_[8901]_  = \new_[8900]_  & \new_[8897]_ ;
  assign \new_[8902]_  = \new_[8901]_  & \new_[8894]_ ;
  assign \new_[8906]_  = A201 & A200;
  assign \new_[8907]_  = ~A199 & \new_[8906]_ ;
  assign \new_[8910]_  = ~A232 & ~A203;
  assign \new_[8913]_  = A234 & A233;
  assign \new_[8914]_  = \new_[8913]_  & \new_[8910]_ ;
  assign \new_[8915]_  = \new_[8914]_  & \new_[8907]_ ;
  assign \new_[8919]_  = ~A266 & ~A265;
  assign \new_[8920]_  = A235 & \new_[8919]_ ;
  assign \new_[8923]_  = ~A299 & A298;
  assign \new_[8926]_  = ~A302 & A300;
  assign \new_[8927]_  = \new_[8926]_  & \new_[8923]_ ;
  assign \new_[8928]_  = \new_[8927]_  & \new_[8920]_ ;
  assign \new_[8932]_  = A201 & A200;
  assign \new_[8933]_  = ~A199 & \new_[8932]_ ;
  assign \new_[8936]_  = ~A232 & ~A203;
  assign \new_[8939]_  = A234 & A233;
  assign \new_[8940]_  = \new_[8939]_  & \new_[8936]_ ;
  assign \new_[8941]_  = \new_[8940]_  & \new_[8933]_ ;
  assign \new_[8945]_  = ~A266 & ~A265;
  assign \new_[8946]_  = A235 & \new_[8945]_ ;
  assign \new_[8949]_  = A299 & ~A298;
  assign \new_[8952]_  = A301 & A300;
  assign \new_[8953]_  = \new_[8952]_  & \new_[8949]_ ;
  assign \new_[8954]_  = \new_[8953]_  & \new_[8946]_ ;
  assign \new_[8958]_  = A201 & A200;
  assign \new_[8959]_  = ~A199 & \new_[8958]_ ;
  assign \new_[8962]_  = ~A232 & ~A203;
  assign \new_[8965]_  = A234 & A233;
  assign \new_[8966]_  = \new_[8965]_  & \new_[8962]_ ;
  assign \new_[8967]_  = \new_[8966]_  & \new_[8959]_ ;
  assign \new_[8971]_  = ~A266 & ~A265;
  assign \new_[8972]_  = A235 & \new_[8971]_ ;
  assign \new_[8975]_  = A299 & ~A298;
  assign \new_[8978]_  = ~A302 & A300;
  assign \new_[8979]_  = \new_[8978]_  & \new_[8975]_ ;
  assign \new_[8980]_  = \new_[8979]_  & \new_[8972]_ ;
  assign \new_[8984]_  = A201 & A200;
  assign \new_[8985]_  = ~A199 & \new_[8984]_ ;
  assign \new_[8988]_  = ~A232 & ~A203;
  assign \new_[8991]_  = A234 & A233;
  assign \new_[8992]_  = \new_[8991]_  & \new_[8988]_ ;
  assign \new_[8993]_  = \new_[8992]_  & \new_[8985]_ ;
  assign \new_[8997]_  = A268 & ~A267;
  assign \new_[8998]_  = ~A236 & \new_[8997]_ ;
  assign \new_[9001]_  = ~A299 & A298;
  assign \new_[9004]_  = A301 & A300;
  assign \new_[9005]_  = \new_[9004]_  & \new_[9001]_ ;
  assign \new_[9006]_  = \new_[9005]_  & \new_[8998]_ ;
  assign \new_[9010]_  = A201 & A200;
  assign \new_[9011]_  = ~A199 & \new_[9010]_ ;
  assign \new_[9014]_  = ~A232 & ~A203;
  assign \new_[9017]_  = A234 & A233;
  assign \new_[9018]_  = \new_[9017]_  & \new_[9014]_ ;
  assign \new_[9019]_  = \new_[9018]_  & \new_[9011]_ ;
  assign \new_[9023]_  = A268 & ~A267;
  assign \new_[9024]_  = ~A236 & \new_[9023]_ ;
  assign \new_[9027]_  = ~A299 & A298;
  assign \new_[9030]_  = ~A302 & A300;
  assign \new_[9031]_  = \new_[9030]_  & \new_[9027]_ ;
  assign \new_[9032]_  = \new_[9031]_  & \new_[9024]_ ;
  assign \new_[9036]_  = A201 & A200;
  assign \new_[9037]_  = ~A199 & \new_[9036]_ ;
  assign \new_[9040]_  = ~A232 & ~A203;
  assign \new_[9043]_  = A234 & A233;
  assign \new_[9044]_  = \new_[9043]_  & \new_[9040]_ ;
  assign \new_[9045]_  = \new_[9044]_  & \new_[9037]_ ;
  assign \new_[9049]_  = A268 & ~A267;
  assign \new_[9050]_  = ~A236 & \new_[9049]_ ;
  assign \new_[9053]_  = A299 & ~A298;
  assign \new_[9056]_  = A301 & A300;
  assign \new_[9057]_  = \new_[9056]_  & \new_[9053]_ ;
  assign \new_[9058]_  = \new_[9057]_  & \new_[9050]_ ;
  assign \new_[9062]_  = A201 & A200;
  assign \new_[9063]_  = ~A199 & \new_[9062]_ ;
  assign \new_[9066]_  = ~A232 & ~A203;
  assign \new_[9069]_  = A234 & A233;
  assign \new_[9070]_  = \new_[9069]_  & \new_[9066]_ ;
  assign \new_[9071]_  = \new_[9070]_  & \new_[9063]_ ;
  assign \new_[9075]_  = A268 & ~A267;
  assign \new_[9076]_  = ~A236 & \new_[9075]_ ;
  assign \new_[9079]_  = A299 & ~A298;
  assign \new_[9082]_  = ~A302 & A300;
  assign \new_[9083]_  = \new_[9082]_  & \new_[9079]_ ;
  assign \new_[9084]_  = \new_[9083]_  & \new_[9076]_ ;
  assign \new_[9088]_  = A201 & A200;
  assign \new_[9089]_  = ~A199 & \new_[9088]_ ;
  assign \new_[9092]_  = ~A232 & ~A203;
  assign \new_[9095]_  = A234 & A233;
  assign \new_[9096]_  = \new_[9095]_  & \new_[9092]_ ;
  assign \new_[9097]_  = \new_[9096]_  & \new_[9089]_ ;
  assign \new_[9101]_  = ~A269 & ~A267;
  assign \new_[9102]_  = ~A236 & \new_[9101]_ ;
  assign \new_[9105]_  = ~A299 & A298;
  assign \new_[9108]_  = A301 & A300;
  assign \new_[9109]_  = \new_[9108]_  & \new_[9105]_ ;
  assign \new_[9110]_  = \new_[9109]_  & \new_[9102]_ ;
  assign \new_[9114]_  = A201 & A200;
  assign \new_[9115]_  = ~A199 & \new_[9114]_ ;
  assign \new_[9118]_  = ~A232 & ~A203;
  assign \new_[9121]_  = A234 & A233;
  assign \new_[9122]_  = \new_[9121]_  & \new_[9118]_ ;
  assign \new_[9123]_  = \new_[9122]_  & \new_[9115]_ ;
  assign \new_[9127]_  = ~A269 & ~A267;
  assign \new_[9128]_  = ~A236 & \new_[9127]_ ;
  assign \new_[9131]_  = ~A299 & A298;
  assign \new_[9134]_  = ~A302 & A300;
  assign \new_[9135]_  = \new_[9134]_  & \new_[9131]_ ;
  assign \new_[9136]_  = \new_[9135]_  & \new_[9128]_ ;
  assign \new_[9140]_  = A201 & A200;
  assign \new_[9141]_  = ~A199 & \new_[9140]_ ;
  assign \new_[9144]_  = ~A232 & ~A203;
  assign \new_[9147]_  = A234 & A233;
  assign \new_[9148]_  = \new_[9147]_  & \new_[9144]_ ;
  assign \new_[9149]_  = \new_[9148]_  & \new_[9141]_ ;
  assign \new_[9153]_  = ~A269 & ~A267;
  assign \new_[9154]_  = ~A236 & \new_[9153]_ ;
  assign \new_[9157]_  = A299 & ~A298;
  assign \new_[9160]_  = A301 & A300;
  assign \new_[9161]_  = \new_[9160]_  & \new_[9157]_ ;
  assign \new_[9162]_  = \new_[9161]_  & \new_[9154]_ ;
  assign \new_[9166]_  = A201 & A200;
  assign \new_[9167]_  = ~A199 & \new_[9166]_ ;
  assign \new_[9170]_  = ~A232 & ~A203;
  assign \new_[9173]_  = A234 & A233;
  assign \new_[9174]_  = \new_[9173]_  & \new_[9170]_ ;
  assign \new_[9175]_  = \new_[9174]_  & \new_[9167]_ ;
  assign \new_[9179]_  = ~A269 & ~A267;
  assign \new_[9180]_  = ~A236 & \new_[9179]_ ;
  assign \new_[9183]_  = A299 & ~A298;
  assign \new_[9186]_  = ~A302 & A300;
  assign \new_[9187]_  = \new_[9186]_  & \new_[9183]_ ;
  assign \new_[9188]_  = \new_[9187]_  & \new_[9180]_ ;
  assign \new_[9192]_  = A201 & A200;
  assign \new_[9193]_  = ~A199 & \new_[9192]_ ;
  assign \new_[9196]_  = ~A232 & ~A203;
  assign \new_[9199]_  = A234 & A233;
  assign \new_[9200]_  = \new_[9199]_  & \new_[9196]_ ;
  assign \new_[9201]_  = \new_[9200]_  & \new_[9193]_ ;
  assign \new_[9205]_  = A266 & A265;
  assign \new_[9206]_  = ~A236 & \new_[9205]_ ;
  assign \new_[9209]_  = ~A299 & A298;
  assign \new_[9212]_  = A301 & A300;
  assign \new_[9213]_  = \new_[9212]_  & \new_[9209]_ ;
  assign \new_[9214]_  = \new_[9213]_  & \new_[9206]_ ;
  assign \new_[9218]_  = A201 & A200;
  assign \new_[9219]_  = ~A199 & \new_[9218]_ ;
  assign \new_[9222]_  = ~A232 & ~A203;
  assign \new_[9225]_  = A234 & A233;
  assign \new_[9226]_  = \new_[9225]_  & \new_[9222]_ ;
  assign \new_[9227]_  = \new_[9226]_  & \new_[9219]_ ;
  assign \new_[9231]_  = A266 & A265;
  assign \new_[9232]_  = ~A236 & \new_[9231]_ ;
  assign \new_[9235]_  = ~A299 & A298;
  assign \new_[9238]_  = ~A302 & A300;
  assign \new_[9239]_  = \new_[9238]_  & \new_[9235]_ ;
  assign \new_[9240]_  = \new_[9239]_  & \new_[9232]_ ;
  assign \new_[9244]_  = A201 & A200;
  assign \new_[9245]_  = ~A199 & \new_[9244]_ ;
  assign \new_[9248]_  = ~A232 & ~A203;
  assign \new_[9251]_  = A234 & A233;
  assign \new_[9252]_  = \new_[9251]_  & \new_[9248]_ ;
  assign \new_[9253]_  = \new_[9252]_  & \new_[9245]_ ;
  assign \new_[9257]_  = A266 & A265;
  assign \new_[9258]_  = ~A236 & \new_[9257]_ ;
  assign \new_[9261]_  = A299 & ~A298;
  assign \new_[9264]_  = A301 & A300;
  assign \new_[9265]_  = \new_[9264]_  & \new_[9261]_ ;
  assign \new_[9266]_  = \new_[9265]_  & \new_[9258]_ ;
  assign \new_[9270]_  = A201 & A200;
  assign \new_[9271]_  = ~A199 & \new_[9270]_ ;
  assign \new_[9274]_  = ~A232 & ~A203;
  assign \new_[9277]_  = A234 & A233;
  assign \new_[9278]_  = \new_[9277]_  & \new_[9274]_ ;
  assign \new_[9279]_  = \new_[9278]_  & \new_[9271]_ ;
  assign \new_[9283]_  = A266 & A265;
  assign \new_[9284]_  = ~A236 & \new_[9283]_ ;
  assign \new_[9287]_  = A299 & ~A298;
  assign \new_[9290]_  = ~A302 & A300;
  assign \new_[9291]_  = \new_[9290]_  & \new_[9287]_ ;
  assign \new_[9292]_  = \new_[9291]_  & \new_[9284]_ ;
  assign \new_[9296]_  = A201 & A200;
  assign \new_[9297]_  = ~A199 & \new_[9296]_ ;
  assign \new_[9300]_  = ~A232 & ~A203;
  assign \new_[9303]_  = A234 & A233;
  assign \new_[9304]_  = \new_[9303]_  & \new_[9300]_ ;
  assign \new_[9305]_  = \new_[9304]_  & \new_[9297]_ ;
  assign \new_[9309]_  = ~A266 & ~A265;
  assign \new_[9310]_  = ~A236 & \new_[9309]_ ;
  assign \new_[9313]_  = ~A299 & A298;
  assign \new_[9316]_  = A301 & A300;
  assign \new_[9317]_  = \new_[9316]_  & \new_[9313]_ ;
  assign \new_[9318]_  = \new_[9317]_  & \new_[9310]_ ;
  assign \new_[9322]_  = A201 & A200;
  assign \new_[9323]_  = ~A199 & \new_[9322]_ ;
  assign \new_[9326]_  = ~A232 & ~A203;
  assign \new_[9329]_  = A234 & A233;
  assign \new_[9330]_  = \new_[9329]_  & \new_[9326]_ ;
  assign \new_[9331]_  = \new_[9330]_  & \new_[9323]_ ;
  assign \new_[9335]_  = ~A266 & ~A265;
  assign \new_[9336]_  = ~A236 & \new_[9335]_ ;
  assign \new_[9339]_  = ~A299 & A298;
  assign \new_[9342]_  = ~A302 & A300;
  assign \new_[9343]_  = \new_[9342]_  & \new_[9339]_ ;
  assign \new_[9344]_  = \new_[9343]_  & \new_[9336]_ ;
  assign \new_[9348]_  = A201 & A200;
  assign \new_[9349]_  = ~A199 & \new_[9348]_ ;
  assign \new_[9352]_  = ~A232 & ~A203;
  assign \new_[9355]_  = A234 & A233;
  assign \new_[9356]_  = \new_[9355]_  & \new_[9352]_ ;
  assign \new_[9357]_  = \new_[9356]_  & \new_[9349]_ ;
  assign \new_[9361]_  = ~A266 & ~A265;
  assign \new_[9362]_  = ~A236 & \new_[9361]_ ;
  assign \new_[9365]_  = A299 & ~A298;
  assign \new_[9368]_  = A301 & A300;
  assign \new_[9369]_  = \new_[9368]_  & \new_[9365]_ ;
  assign \new_[9370]_  = \new_[9369]_  & \new_[9362]_ ;
  assign \new_[9374]_  = A201 & A200;
  assign \new_[9375]_  = ~A199 & \new_[9374]_ ;
  assign \new_[9378]_  = ~A232 & ~A203;
  assign \new_[9381]_  = A234 & A233;
  assign \new_[9382]_  = \new_[9381]_  & \new_[9378]_ ;
  assign \new_[9383]_  = \new_[9382]_  & \new_[9375]_ ;
  assign \new_[9387]_  = ~A266 & ~A265;
  assign \new_[9388]_  = ~A236 & \new_[9387]_ ;
  assign \new_[9391]_  = A299 & ~A298;
  assign \new_[9394]_  = ~A302 & A300;
  assign \new_[9395]_  = \new_[9394]_  & \new_[9391]_ ;
  assign \new_[9396]_  = \new_[9395]_  & \new_[9388]_ ;
  assign \new_[9400]_  = A201 & A200;
  assign \new_[9401]_  = ~A199 & \new_[9400]_ ;
  assign \new_[9404]_  = A232 & ~A203;
  assign \new_[9407]_  = A234 & ~A233;
  assign \new_[9408]_  = \new_[9407]_  & \new_[9404]_ ;
  assign \new_[9409]_  = \new_[9408]_  & \new_[9401]_ ;
  assign \new_[9413]_  = A268 & ~A267;
  assign \new_[9414]_  = A235 & \new_[9413]_ ;
  assign \new_[9417]_  = ~A299 & A298;
  assign \new_[9420]_  = A301 & A300;
  assign \new_[9421]_  = \new_[9420]_  & \new_[9417]_ ;
  assign \new_[9422]_  = \new_[9421]_  & \new_[9414]_ ;
  assign \new_[9426]_  = A201 & A200;
  assign \new_[9427]_  = ~A199 & \new_[9426]_ ;
  assign \new_[9430]_  = A232 & ~A203;
  assign \new_[9433]_  = A234 & ~A233;
  assign \new_[9434]_  = \new_[9433]_  & \new_[9430]_ ;
  assign \new_[9435]_  = \new_[9434]_  & \new_[9427]_ ;
  assign \new_[9439]_  = A268 & ~A267;
  assign \new_[9440]_  = A235 & \new_[9439]_ ;
  assign \new_[9443]_  = ~A299 & A298;
  assign \new_[9446]_  = ~A302 & A300;
  assign \new_[9447]_  = \new_[9446]_  & \new_[9443]_ ;
  assign \new_[9448]_  = \new_[9447]_  & \new_[9440]_ ;
  assign \new_[9452]_  = A201 & A200;
  assign \new_[9453]_  = ~A199 & \new_[9452]_ ;
  assign \new_[9456]_  = A232 & ~A203;
  assign \new_[9459]_  = A234 & ~A233;
  assign \new_[9460]_  = \new_[9459]_  & \new_[9456]_ ;
  assign \new_[9461]_  = \new_[9460]_  & \new_[9453]_ ;
  assign \new_[9465]_  = A268 & ~A267;
  assign \new_[9466]_  = A235 & \new_[9465]_ ;
  assign \new_[9469]_  = A299 & ~A298;
  assign \new_[9472]_  = A301 & A300;
  assign \new_[9473]_  = \new_[9472]_  & \new_[9469]_ ;
  assign \new_[9474]_  = \new_[9473]_  & \new_[9466]_ ;
  assign \new_[9478]_  = A201 & A200;
  assign \new_[9479]_  = ~A199 & \new_[9478]_ ;
  assign \new_[9482]_  = A232 & ~A203;
  assign \new_[9485]_  = A234 & ~A233;
  assign \new_[9486]_  = \new_[9485]_  & \new_[9482]_ ;
  assign \new_[9487]_  = \new_[9486]_  & \new_[9479]_ ;
  assign \new_[9491]_  = A268 & ~A267;
  assign \new_[9492]_  = A235 & \new_[9491]_ ;
  assign \new_[9495]_  = A299 & ~A298;
  assign \new_[9498]_  = ~A302 & A300;
  assign \new_[9499]_  = \new_[9498]_  & \new_[9495]_ ;
  assign \new_[9500]_  = \new_[9499]_  & \new_[9492]_ ;
  assign \new_[9504]_  = A201 & A200;
  assign \new_[9505]_  = ~A199 & \new_[9504]_ ;
  assign \new_[9508]_  = A232 & ~A203;
  assign \new_[9511]_  = A234 & ~A233;
  assign \new_[9512]_  = \new_[9511]_  & \new_[9508]_ ;
  assign \new_[9513]_  = \new_[9512]_  & \new_[9505]_ ;
  assign \new_[9517]_  = ~A269 & ~A267;
  assign \new_[9518]_  = A235 & \new_[9517]_ ;
  assign \new_[9521]_  = ~A299 & A298;
  assign \new_[9524]_  = A301 & A300;
  assign \new_[9525]_  = \new_[9524]_  & \new_[9521]_ ;
  assign \new_[9526]_  = \new_[9525]_  & \new_[9518]_ ;
  assign \new_[9530]_  = A201 & A200;
  assign \new_[9531]_  = ~A199 & \new_[9530]_ ;
  assign \new_[9534]_  = A232 & ~A203;
  assign \new_[9537]_  = A234 & ~A233;
  assign \new_[9538]_  = \new_[9537]_  & \new_[9534]_ ;
  assign \new_[9539]_  = \new_[9538]_  & \new_[9531]_ ;
  assign \new_[9543]_  = ~A269 & ~A267;
  assign \new_[9544]_  = A235 & \new_[9543]_ ;
  assign \new_[9547]_  = ~A299 & A298;
  assign \new_[9550]_  = ~A302 & A300;
  assign \new_[9551]_  = \new_[9550]_  & \new_[9547]_ ;
  assign \new_[9552]_  = \new_[9551]_  & \new_[9544]_ ;
  assign \new_[9556]_  = A201 & A200;
  assign \new_[9557]_  = ~A199 & \new_[9556]_ ;
  assign \new_[9560]_  = A232 & ~A203;
  assign \new_[9563]_  = A234 & ~A233;
  assign \new_[9564]_  = \new_[9563]_  & \new_[9560]_ ;
  assign \new_[9565]_  = \new_[9564]_  & \new_[9557]_ ;
  assign \new_[9569]_  = ~A269 & ~A267;
  assign \new_[9570]_  = A235 & \new_[9569]_ ;
  assign \new_[9573]_  = A299 & ~A298;
  assign \new_[9576]_  = A301 & A300;
  assign \new_[9577]_  = \new_[9576]_  & \new_[9573]_ ;
  assign \new_[9578]_  = \new_[9577]_  & \new_[9570]_ ;
  assign \new_[9582]_  = A201 & A200;
  assign \new_[9583]_  = ~A199 & \new_[9582]_ ;
  assign \new_[9586]_  = A232 & ~A203;
  assign \new_[9589]_  = A234 & ~A233;
  assign \new_[9590]_  = \new_[9589]_  & \new_[9586]_ ;
  assign \new_[9591]_  = \new_[9590]_  & \new_[9583]_ ;
  assign \new_[9595]_  = ~A269 & ~A267;
  assign \new_[9596]_  = A235 & \new_[9595]_ ;
  assign \new_[9599]_  = A299 & ~A298;
  assign \new_[9602]_  = ~A302 & A300;
  assign \new_[9603]_  = \new_[9602]_  & \new_[9599]_ ;
  assign \new_[9604]_  = \new_[9603]_  & \new_[9596]_ ;
  assign \new_[9608]_  = A201 & A200;
  assign \new_[9609]_  = ~A199 & \new_[9608]_ ;
  assign \new_[9612]_  = A232 & ~A203;
  assign \new_[9615]_  = A234 & ~A233;
  assign \new_[9616]_  = \new_[9615]_  & \new_[9612]_ ;
  assign \new_[9617]_  = \new_[9616]_  & \new_[9609]_ ;
  assign \new_[9621]_  = A266 & A265;
  assign \new_[9622]_  = A235 & \new_[9621]_ ;
  assign \new_[9625]_  = ~A299 & A298;
  assign \new_[9628]_  = A301 & A300;
  assign \new_[9629]_  = \new_[9628]_  & \new_[9625]_ ;
  assign \new_[9630]_  = \new_[9629]_  & \new_[9622]_ ;
  assign \new_[9634]_  = A201 & A200;
  assign \new_[9635]_  = ~A199 & \new_[9634]_ ;
  assign \new_[9638]_  = A232 & ~A203;
  assign \new_[9641]_  = A234 & ~A233;
  assign \new_[9642]_  = \new_[9641]_  & \new_[9638]_ ;
  assign \new_[9643]_  = \new_[9642]_  & \new_[9635]_ ;
  assign \new_[9647]_  = A266 & A265;
  assign \new_[9648]_  = A235 & \new_[9647]_ ;
  assign \new_[9651]_  = ~A299 & A298;
  assign \new_[9654]_  = ~A302 & A300;
  assign \new_[9655]_  = \new_[9654]_  & \new_[9651]_ ;
  assign \new_[9656]_  = \new_[9655]_  & \new_[9648]_ ;
  assign \new_[9660]_  = A201 & A200;
  assign \new_[9661]_  = ~A199 & \new_[9660]_ ;
  assign \new_[9664]_  = A232 & ~A203;
  assign \new_[9667]_  = A234 & ~A233;
  assign \new_[9668]_  = \new_[9667]_  & \new_[9664]_ ;
  assign \new_[9669]_  = \new_[9668]_  & \new_[9661]_ ;
  assign \new_[9673]_  = A266 & A265;
  assign \new_[9674]_  = A235 & \new_[9673]_ ;
  assign \new_[9677]_  = A299 & ~A298;
  assign \new_[9680]_  = A301 & A300;
  assign \new_[9681]_  = \new_[9680]_  & \new_[9677]_ ;
  assign \new_[9682]_  = \new_[9681]_  & \new_[9674]_ ;
  assign \new_[9686]_  = A201 & A200;
  assign \new_[9687]_  = ~A199 & \new_[9686]_ ;
  assign \new_[9690]_  = A232 & ~A203;
  assign \new_[9693]_  = A234 & ~A233;
  assign \new_[9694]_  = \new_[9693]_  & \new_[9690]_ ;
  assign \new_[9695]_  = \new_[9694]_  & \new_[9687]_ ;
  assign \new_[9699]_  = A266 & A265;
  assign \new_[9700]_  = A235 & \new_[9699]_ ;
  assign \new_[9703]_  = A299 & ~A298;
  assign \new_[9706]_  = ~A302 & A300;
  assign \new_[9707]_  = \new_[9706]_  & \new_[9703]_ ;
  assign \new_[9708]_  = \new_[9707]_  & \new_[9700]_ ;
  assign \new_[9712]_  = A201 & A200;
  assign \new_[9713]_  = ~A199 & \new_[9712]_ ;
  assign \new_[9716]_  = A232 & ~A203;
  assign \new_[9719]_  = A234 & ~A233;
  assign \new_[9720]_  = \new_[9719]_  & \new_[9716]_ ;
  assign \new_[9721]_  = \new_[9720]_  & \new_[9713]_ ;
  assign \new_[9725]_  = ~A266 & ~A265;
  assign \new_[9726]_  = A235 & \new_[9725]_ ;
  assign \new_[9729]_  = ~A299 & A298;
  assign \new_[9732]_  = A301 & A300;
  assign \new_[9733]_  = \new_[9732]_  & \new_[9729]_ ;
  assign \new_[9734]_  = \new_[9733]_  & \new_[9726]_ ;
  assign \new_[9738]_  = A201 & A200;
  assign \new_[9739]_  = ~A199 & \new_[9738]_ ;
  assign \new_[9742]_  = A232 & ~A203;
  assign \new_[9745]_  = A234 & ~A233;
  assign \new_[9746]_  = \new_[9745]_  & \new_[9742]_ ;
  assign \new_[9747]_  = \new_[9746]_  & \new_[9739]_ ;
  assign \new_[9751]_  = ~A266 & ~A265;
  assign \new_[9752]_  = A235 & \new_[9751]_ ;
  assign \new_[9755]_  = ~A299 & A298;
  assign \new_[9758]_  = ~A302 & A300;
  assign \new_[9759]_  = \new_[9758]_  & \new_[9755]_ ;
  assign \new_[9760]_  = \new_[9759]_  & \new_[9752]_ ;
  assign \new_[9764]_  = A201 & A200;
  assign \new_[9765]_  = ~A199 & \new_[9764]_ ;
  assign \new_[9768]_  = A232 & ~A203;
  assign \new_[9771]_  = A234 & ~A233;
  assign \new_[9772]_  = \new_[9771]_  & \new_[9768]_ ;
  assign \new_[9773]_  = \new_[9772]_  & \new_[9765]_ ;
  assign \new_[9777]_  = ~A266 & ~A265;
  assign \new_[9778]_  = A235 & \new_[9777]_ ;
  assign \new_[9781]_  = A299 & ~A298;
  assign \new_[9784]_  = A301 & A300;
  assign \new_[9785]_  = \new_[9784]_  & \new_[9781]_ ;
  assign \new_[9786]_  = \new_[9785]_  & \new_[9778]_ ;
  assign \new_[9790]_  = A201 & A200;
  assign \new_[9791]_  = ~A199 & \new_[9790]_ ;
  assign \new_[9794]_  = A232 & ~A203;
  assign \new_[9797]_  = A234 & ~A233;
  assign \new_[9798]_  = \new_[9797]_  & \new_[9794]_ ;
  assign \new_[9799]_  = \new_[9798]_  & \new_[9791]_ ;
  assign \new_[9803]_  = ~A266 & ~A265;
  assign \new_[9804]_  = A235 & \new_[9803]_ ;
  assign \new_[9807]_  = A299 & ~A298;
  assign \new_[9810]_  = ~A302 & A300;
  assign \new_[9811]_  = \new_[9810]_  & \new_[9807]_ ;
  assign \new_[9812]_  = \new_[9811]_  & \new_[9804]_ ;
  assign \new_[9816]_  = A201 & A200;
  assign \new_[9817]_  = ~A199 & \new_[9816]_ ;
  assign \new_[9820]_  = A232 & ~A203;
  assign \new_[9823]_  = A234 & ~A233;
  assign \new_[9824]_  = \new_[9823]_  & \new_[9820]_ ;
  assign \new_[9825]_  = \new_[9824]_  & \new_[9817]_ ;
  assign \new_[9829]_  = A268 & ~A267;
  assign \new_[9830]_  = ~A236 & \new_[9829]_ ;
  assign \new_[9833]_  = ~A299 & A298;
  assign \new_[9836]_  = A301 & A300;
  assign \new_[9837]_  = \new_[9836]_  & \new_[9833]_ ;
  assign \new_[9838]_  = \new_[9837]_  & \new_[9830]_ ;
  assign \new_[9842]_  = A201 & A200;
  assign \new_[9843]_  = ~A199 & \new_[9842]_ ;
  assign \new_[9846]_  = A232 & ~A203;
  assign \new_[9849]_  = A234 & ~A233;
  assign \new_[9850]_  = \new_[9849]_  & \new_[9846]_ ;
  assign \new_[9851]_  = \new_[9850]_  & \new_[9843]_ ;
  assign \new_[9855]_  = A268 & ~A267;
  assign \new_[9856]_  = ~A236 & \new_[9855]_ ;
  assign \new_[9859]_  = ~A299 & A298;
  assign \new_[9862]_  = ~A302 & A300;
  assign \new_[9863]_  = \new_[9862]_  & \new_[9859]_ ;
  assign \new_[9864]_  = \new_[9863]_  & \new_[9856]_ ;
  assign \new_[9868]_  = A201 & A200;
  assign \new_[9869]_  = ~A199 & \new_[9868]_ ;
  assign \new_[9872]_  = A232 & ~A203;
  assign \new_[9875]_  = A234 & ~A233;
  assign \new_[9876]_  = \new_[9875]_  & \new_[9872]_ ;
  assign \new_[9877]_  = \new_[9876]_  & \new_[9869]_ ;
  assign \new_[9881]_  = A268 & ~A267;
  assign \new_[9882]_  = ~A236 & \new_[9881]_ ;
  assign \new_[9885]_  = A299 & ~A298;
  assign \new_[9888]_  = A301 & A300;
  assign \new_[9889]_  = \new_[9888]_  & \new_[9885]_ ;
  assign \new_[9890]_  = \new_[9889]_  & \new_[9882]_ ;
  assign \new_[9894]_  = A201 & A200;
  assign \new_[9895]_  = ~A199 & \new_[9894]_ ;
  assign \new_[9898]_  = A232 & ~A203;
  assign \new_[9901]_  = A234 & ~A233;
  assign \new_[9902]_  = \new_[9901]_  & \new_[9898]_ ;
  assign \new_[9903]_  = \new_[9902]_  & \new_[9895]_ ;
  assign \new_[9907]_  = A268 & ~A267;
  assign \new_[9908]_  = ~A236 & \new_[9907]_ ;
  assign \new_[9911]_  = A299 & ~A298;
  assign \new_[9914]_  = ~A302 & A300;
  assign \new_[9915]_  = \new_[9914]_  & \new_[9911]_ ;
  assign \new_[9916]_  = \new_[9915]_  & \new_[9908]_ ;
  assign \new_[9920]_  = A201 & A200;
  assign \new_[9921]_  = ~A199 & \new_[9920]_ ;
  assign \new_[9924]_  = A232 & ~A203;
  assign \new_[9927]_  = A234 & ~A233;
  assign \new_[9928]_  = \new_[9927]_  & \new_[9924]_ ;
  assign \new_[9929]_  = \new_[9928]_  & \new_[9921]_ ;
  assign \new_[9933]_  = ~A269 & ~A267;
  assign \new_[9934]_  = ~A236 & \new_[9933]_ ;
  assign \new_[9937]_  = ~A299 & A298;
  assign \new_[9940]_  = A301 & A300;
  assign \new_[9941]_  = \new_[9940]_  & \new_[9937]_ ;
  assign \new_[9942]_  = \new_[9941]_  & \new_[9934]_ ;
  assign \new_[9946]_  = A201 & A200;
  assign \new_[9947]_  = ~A199 & \new_[9946]_ ;
  assign \new_[9950]_  = A232 & ~A203;
  assign \new_[9953]_  = A234 & ~A233;
  assign \new_[9954]_  = \new_[9953]_  & \new_[9950]_ ;
  assign \new_[9955]_  = \new_[9954]_  & \new_[9947]_ ;
  assign \new_[9959]_  = ~A269 & ~A267;
  assign \new_[9960]_  = ~A236 & \new_[9959]_ ;
  assign \new_[9963]_  = ~A299 & A298;
  assign \new_[9966]_  = ~A302 & A300;
  assign \new_[9967]_  = \new_[9966]_  & \new_[9963]_ ;
  assign \new_[9968]_  = \new_[9967]_  & \new_[9960]_ ;
  assign \new_[9972]_  = A201 & A200;
  assign \new_[9973]_  = ~A199 & \new_[9972]_ ;
  assign \new_[9976]_  = A232 & ~A203;
  assign \new_[9979]_  = A234 & ~A233;
  assign \new_[9980]_  = \new_[9979]_  & \new_[9976]_ ;
  assign \new_[9981]_  = \new_[9980]_  & \new_[9973]_ ;
  assign \new_[9985]_  = ~A269 & ~A267;
  assign \new_[9986]_  = ~A236 & \new_[9985]_ ;
  assign \new_[9989]_  = A299 & ~A298;
  assign \new_[9992]_  = A301 & A300;
  assign \new_[9993]_  = \new_[9992]_  & \new_[9989]_ ;
  assign \new_[9994]_  = \new_[9993]_  & \new_[9986]_ ;
  assign \new_[9998]_  = A201 & A200;
  assign \new_[9999]_  = ~A199 & \new_[9998]_ ;
  assign \new_[10002]_  = A232 & ~A203;
  assign \new_[10005]_  = A234 & ~A233;
  assign \new_[10006]_  = \new_[10005]_  & \new_[10002]_ ;
  assign \new_[10007]_  = \new_[10006]_  & \new_[9999]_ ;
  assign \new_[10011]_  = ~A269 & ~A267;
  assign \new_[10012]_  = ~A236 & \new_[10011]_ ;
  assign \new_[10015]_  = A299 & ~A298;
  assign \new_[10018]_  = ~A302 & A300;
  assign \new_[10019]_  = \new_[10018]_  & \new_[10015]_ ;
  assign \new_[10020]_  = \new_[10019]_  & \new_[10012]_ ;
  assign \new_[10024]_  = A201 & A200;
  assign \new_[10025]_  = ~A199 & \new_[10024]_ ;
  assign \new_[10028]_  = A232 & ~A203;
  assign \new_[10031]_  = A234 & ~A233;
  assign \new_[10032]_  = \new_[10031]_  & \new_[10028]_ ;
  assign \new_[10033]_  = \new_[10032]_  & \new_[10025]_ ;
  assign \new_[10037]_  = A266 & A265;
  assign \new_[10038]_  = ~A236 & \new_[10037]_ ;
  assign \new_[10041]_  = ~A299 & A298;
  assign \new_[10044]_  = A301 & A300;
  assign \new_[10045]_  = \new_[10044]_  & \new_[10041]_ ;
  assign \new_[10046]_  = \new_[10045]_  & \new_[10038]_ ;
  assign \new_[10050]_  = A201 & A200;
  assign \new_[10051]_  = ~A199 & \new_[10050]_ ;
  assign \new_[10054]_  = A232 & ~A203;
  assign \new_[10057]_  = A234 & ~A233;
  assign \new_[10058]_  = \new_[10057]_  & \new_[10054]_ ;
  assign \new_[10059]_  = \new_[10058]_  & \new_[10051]_ ;
  assign \new_[10063]_  = A266 & A265;
  assign \new_[10064]_  = ~A236 & \new_[10063]_ ;
  assign \new_[10067]_  = ~A299 & A298;
  assign \new_[10070]_  = ~A302 & A300;
  assign \new_[10071]_  = \new_[10070]_  & \new_[10067]_ ;
  assign \new_[10072]_  = \new_[10071]_  & \new_[10064]_ ;
  assign \new_[10076]_  = A201 & A200;
  assign \new_[10077]_  = ~A199 & \new_[10076]_ ;
  assign \new_[10080]_  = A232 & ~A203;
  assign \new_[10083]_  = A234 & ~A233;
  assign \new_[10084]_  = \new_[10083]_  & \new_[10080]_ ;
  assign \new_[10085]_  = \new_[10084]_  & \new_[10077]_ ;
  assign \new_[10089]_  = A266 & A265;
  assign \new_[10090]_  = ~A236 & \new_[10089]_ ;
  assign \new_[10093]_  = A299 & ~A298;
  assign \new_[10096]_  = A301 & A300;
  assign \new_[10097]_  = \new_[10096]_  & \new_[10093]_ ;
  assign \new_[10098]_  = \new_[10097]_  & \new_[10090]_ ;
  assign \new_[10102]_  = A201 & A200;
  assign \new_[10103]_  = ~A199 & \new_[10102]_ ;
  assign \new_[10106]_  = A232 & ~A203;
  assign \new_[10109]_  = A234 & ~A233;
  assign \new_[10110]_  = \new_[10109]_  & \new_[10106]_ ;
  assign \new_[10111]_  = \new_[10110]_  & \new_[10103]_ ;
  assign \new_[10115]_  = A266 & A265;
  assign \new_[10116]_  = ~A236 & \new_[10115]_ ;
  assign \new_[10119]_  = A299 & ~A298;
  assign \new_[10122]_  = ~A302 & A300;
  assign \new_[10123]_  = \new_[10122]_  & \new_[10119]_ ;
  assign \new_[10124]_  = \new_[10123]_  & \new_[10116]_ ;
  assign \new_[10128]_  = A201 & A200;
  assign \new_[10129]_  = ~A199 & \new_[10128]_ ;
  assign \new_[10132]_  = A232 & ~A203;
  assign \new_[10135]_  = A234 & ~A233;
  assign \new_[10136]_  = \new_[10135]_  & \new_[10132]_ ;
  assign \new_[10137]_  = \new_[10136]_  & \new_[10129]_ ;
  assign \new_[10141]_  = ~A266 & ~A265;
  assign \new_[10142]_  = ~A236 & \new_[10141]_ ;
  assign \new_[10145]_  = ~A299 & A298;
  assign \new_[10148]_  = A301 & A300;
  assign \new_[10149]_  = \new_[10148]_  & \new_[10145]_ ;
  assign \new_[10150]_  = \new_[10149]_  & \new_[10142]_ ;
  assign \new_[10154]_  = A201 & A200;
  assign \new_[10155]_  = ~A199 & \new_[10154]_ ;
  assign \new_[10158]_  = A232 & ~A203;
  assign \new_[10161]_  = A234 & ~A233;
  assign \new_[10162]_  = \new_[10161]_  & \new_[10158]_ ;
  assign \new_[10163]_  = \new_[10162]_  & \new_[10155]_ ;
  assign \new_[10167]_  = ~A266 & ~A265;
  assign \new_[10168]_  = ~A236 & \new_[10167]_ ;
  assign \new_[10171]_  = ~A299 & A298;
  assign \new_[10174]_  = ~A302 & A300;
  assign \new_[10175]_  = \new_[10174]_  & \new_[10171]_ ;
  assign \new_[10176]_  = \new_[10175]_  & \new_[10168]_ ;
  assign \new_[10180]_  = A201 & A200;
  assign \new_[10181]_  = ~A199 & \new_[10180]_ ;
  assign \new_[10184]_  = A232 & ~A203;
  assign \new_[10187]_  = A234 & ~A233;
  assign \new_[10188]_  = \new_[10187]_  & \new_[10184]_ ;
  assign \new_[10189]_  = \new_[10188]_  & \new_[10181]_ ;
  assign \new_[10193]_  = ~A266 & ~A265;
  assign \new_[10194]_  = ~A236 & \new_[10193]_ ;
  assign \new_[10197]_  = A299 & ~A298;
  assign \new_[10200]_  = A301 & A300;
  assign \new_[10201]_  = \new_[10200]_  & \new_[10197]_ ;
  assign \new_[10202]_  = \new_[10201]_  & \new_[10194]_ ;
  assign \new_[10206]_  = A201 & A200;
  assign \new_[10207]_  = ~A199 & \new_[10206]_ ;
  assign \new_[10210]_  = A232 & ~A203;
  assign \new_[10213]_  = A234 & ~A233;
  assign \new_[10214]_  = \new_[10213]_  & \new_[10210]_ ;
  assign \new_[10215]_  = \new_[10214]_  & \new_[10207]_ ;
  assign \new_[10219]_  = ~A266 & ~A265;
  assign \new_[10220]_  = ~A236 & \new_[10219]_ ;
  assign \new_[10223]_  = A299 & ~A298;
  assign \new_[10226]_  = ~A302 & A300;
  assign \new_[10227]_  = \new_[10226]_  & \new_[10223]_ ;
  assign \new_[10228]_  = \new_[10227]_  & \new_[10220]_ ;
  assign \new_[10232]_  = A201 & ~A200;
  assign \new_[10233]_  = A199 & \new_[10232]_ ;
  assign \new_[10236]_  = ~A232 & A202;
  assign \new_[10239]_  = A234 & A233;
  assign \new_[10240]_  = \new_[10239]_  & \new_[10236]_ ;
  assign \new_[10241]_  = \new_[10240]_  & \new_[10233]_ ;
  assign \new_[10245]_  = A268 & ~A267;
  assign \new_[10246]_  = A235 & \new_[10245]_ ;
  assign \new_[10249]_  = ~A299 & A298;
  assign \new_[10252]_  = A301 & A300;
  assign \new_[10253]_  = \new_[10252]_  & \new_[10249]_ ;
  assign \new_[10254]_  = \new_[10253]_  & \new_[10246]_ ;
  assign \new_[10258]_  = A201 & ~A200;
  assign \new_[10259]_  = A199 & \new_[10258]_ ;
  assign \new_[10262]_  = ~A232 & A202;
  assign \new_[10265]_  = A234 & A233;
  assign \new_[10266]_  = \new_[10265]_  & \new_[10262]_ ;
  assign \new_[10267]_  = \new_[10266]_  & \new_[10259]_ ;
  assign \new_[10271]_  = A268 & ~A267;
  assign \new_[10272]_  = A235 & \new_[10271]_ ;
  assign \new_[10275]_  = ~A299 & A298;
  assign \new_[10278]_  = ~A302 & A300;
  assign \new_[10279]_  = \new_[10278]_  & \new_[10275]_ ;
  assign \new_[10280]_  = \new_[10279]_  & \new_[10272]_ ;
  assign \new_[10284]_  = A201 & ~A200;
  assign \new_[10285]_  = A199 & \new_[10284]_ ;
  assign \new_[10288]_  = ~A232 & A202;
  assign \new_[10291]_  = A234 & A233;
  assign \new_[10292]_  = \new_[10291]_  & \new_[10288]_ ;
  assign \new_[10293]_  = \new_[10292]_  & \new_[10285]_ ;
  assign \new_[10297]_  = A268 & ~A267;
  assign \new_[10298]_  = A235 & \new_[10297]_ ;
  assign \new_[10301]_  = A299 & ~A298;
  assign \new_[10304]_  = A301 & A300;
  assign \new_[10305]_  = \new_[10304]_  & \new_[10301]_ ;
  assign \new_[10306]_  = \new_[10305]_  & \new_[10298]_ ;
  assign \new_[10310]_  = A201 & ~A200;
  assign \new_[10311]_  = A199 & \new_[10310]_ ;
  assign \new_[10314]_  = ~A232 & A202;
  assign \new_[10317]_  = A234 & A233;
  assign \new_[10318]_  = \new_[10317]_  & \new_[10314]_ ;
  assign \new_[10319]_  = \new_[10318]_  & \new_[10311]_ ;
  assign \new_[10323]_  = A268 & ~A267;
  assign \new_[10324]_  = A235 & \new_[10323]_ ;
  assign \new_[10327]_  = A299 & ~A298;
  assign \new_[10330]_  = ~A302 & A300;
  assign \new_[10331]_  = \new_[10330]_  & \new_[10327]_ ;
  assign \new_[10332]_  = \new_[10331]_  & \new_[10324]_ ;
  assign \new_[10336]_  = A201 & ~A200;
  assign \new_[10337]_  = A199 & \new_[10336]_ ;
  assign \new_[10340]_  = ~A232 & A202;
  assign \new_[10343]_  = A234 & A233;
  assign \new_[10344]_  = \new_[10343]_  & \new_[10340]_ ;
  assign \new_[10345]_  = \new_[10344]_  & \new_[10337]_ ;
  assign \new_[10349]_  = ~A269 & ~A267;
  assign \new_[10350]_  = A235 & \new_[10349]_ ;
  assign \new_[10353]_  = ~A299 & A298;
  assign \new_[10356]_  = A301 & A300;
  assign \new_[10357]_  = \new_[10356]_  & \new_[10353]_ ;
  assign \new_[10358]_  = \new_[10357]_  & \new_[10350]_ ;
  assign \new_[10362]_  = A201 & ~A200;
  assign \new_[10363]_  = A199 & \new_[10362]_ ;
  assign \new_[10366]_  = ~A232 & A202;
  assign \new_[10369]_  = A234 & A233;
  assign \new_[10370]_  = \new_[10369]_  & \new_[10366]_ ;
  assign \new_[10371]_  = \new_[10370]_  & \new_[10363]_ ;
  assign \new_[10375]_  = ~A269 & ~A267;
  assign \new_[10376]_  = A235 & \new_[10375]_ ;
  assign \new_[10379]_  = ~A299 & A298;
  assign \new_[10382]_  = ~A302 & A300;
  assign \new_[10383]_  = \new_[10382]_  & \new_[10379]_ ;
  assign \new_[10384]_  = \new_[10383]_  & \new_[10376]_ ;
  assign \new_[10388]_  = A201 & ~A200;
  assign \new_[10389]_  = A199 & \new_[10388]_ ;
  assign \new_[10392]_  = ~A232 & A202;
  assign \new_[10395]_  = A234 & A233;
  assign \new_[10396]_  = \new_[10395]_  & \new_[10392]_ ;
  assign \new_[10397]_  = \new_[10396]_  & \new_[10389]_ ;
  assign \new_[10401]_  = ~A269 & ~A267;
  assign \new_[10402]_  = A235 & \new_[10401]_ ;
  assign \new_[10405]_  = A299 & ~A298;
  assign \new_[10408]_  = A301 & A300;
  assign \new_[10409]_  = \new_[10408]_  & \new_[10405]_ ;
  assign \new_[10410]_  = \new_[10409]_  & \new_[10402]_ ;
  assign \new_[10414]_  = A201 & ~A200;
  assign \new_[10415]_  = A199 & \new_[10414]_ ;
  assign \new_[10418]_  = ~A232 & A202;
  assign \new_[10421]_  = A234 & A233;
  assign \new_[10422]_  = \new_[10421]_  & \new_[10418]_ ;
  assign \new_[10423]_  = \new_[10422]_  & \new_[10415]_ ;
  assign \new_[10427]_  = ~A269 & ~A267;
  assign \new_[10428]_  = A235 & \new_[10427]_ ;
  assign \new_[10431]_  = A299 & ~A298;
  assign \new_[10434]_  = ~A302 & A300;
  assign \new_[10435]_  = \new_[10434]_  & \new_[10431]_ ;
  assign \new_[10436]_  = \new_[10435]_  & \new_[10428]_ ;
  assign \new_[10440]_  = A201 & ~A200;
  assign \new_[10441]_  = A199 & \new_[10440]_ ;
  assign \new_[10444]_  = ~A232 & A202;
  assign \new_[10447]_  = A234 & A233;
  assign \new_[10448]_  = \new_[10447]_  & \new_[10444]_ ;
  assign \new_[10449]_  = \new_[10448]_  & \new_[10441]_ ;
  assign \new_[10453]_  = A266 & A265;
  assign \new_[10454]_  = A235 & \new_[10453]_ ;
  assign \new_[10457]_  = ~A299 & A298;
  assign \new_[10460]_  = A301 & A300;
  assign \new_[10461]_  = \new_[10460]_  & \new_[10457]_ ;
  assign \new_[10462]_  = \new_[10461]_  & \new_[10454]_ ;
  assign \new_[10466]_  = A201 & ~A200;
  assign \new_[10467]_  = A199 & \new_[10466]_ ;
  assign \new_[10470]_  = ~A232 & A202;
  assign \new_[10473]_  = A234 & A233;
  assign \new_[10474]_  = \new_[10473]_  & \new_[10470]_ ;
  assign \new_[10475]_  = \new_[10474]_  & \new_[10467]_ ;
  assign \new_[10479]_  = A266 & A265;
  assign \new_[10480]_  = A235 & \new_[10479]_ ;
  assign \new_[10483]_  = ~A299 & A298;
  assign \new_[10486]_  = ~A302 & A300;
  assign \new_[10487]_  = \new_[10486]_  & \new_[10483]_ ;
  assign \new_[10488]_  = \new_[10487]_  & \new_[10480]_ ;
  assign \new_[10492]_  = A201 & ~A200;
  assign \new_[10493]_  = A199 & \new_[10492]_ ;
  assign \new_[10496]_  = ~A232 & A202;
  assign \new_[10499]_  = A234 & A233;
  assign \new_[10500]_  = \new_[10499]_  & \new_[10496]_ ;
  assign \new_[10501]_  = \new_[10500]_  & \new_[10493]_ ;
  assign \new_[10505]_  = A266 & A265;
  assign \new_[10506]_  = A235 & \new_[10505]_ ;
  assign \new_[10509]_  = A299 & ~A298;
  assign \new_[10512]_  = A301 & A300;
  assign \new_[10513]_  = \new_[10512]_  & \new_[10509]_ ;
  assign \new_[10514]_  = \new_[10513]_  & \new_[10506]_ ;
  assign \new_[10518]_  = A201 & ~A200;
  assign \new_[10519]_  = A199 & \new_[10518]_ ;
  assign \new_[10522]_  = ~A232 & A202;
  assign \new_[10525]_  = A234 & A233;
  assign \new_[10526]_  = \new_[10525]_  & \new_[10522]_ ;
  assign \new_[10527]_  = \new_[10526]_  & \new_[10519]_ ;
  assign \new_[10531]_  = A266 & A265;
  assign \new_[10532]_  = A235 & \new_[10531]_ ;
  assign \new_[10535]_  = A299 & ~A298;
  assign \new_[10538]_  = ~A302 & A300;
  assign \new_[10539]_  = \new_[10538]_  & \new_[10535]_ ;
  assign \new_[10540]_  = \new_[10539]_  & \new_[10532]_ ;
  assign \new_[10544]_  = A201 & ~A200;
  assign \new_[10545]_  = A199 & \new_[10544]_ ;
  assign \new_[10548]_  = ~A232 & A202;
  assign \new_[10551]_  = A234 & A233;
  assign \new_[10552]_  = \new_[10551]_  & \new_[10548]_ ;
  assign \new_[10553]_  = \new_[10552]_  & \new_[10545]_ ;
  assign \new_[10557]_  = ~A266 & ~A265;
  assign \new_[10558]_  = A235 & \new_[10557]_ ;
  assign \new_[10561]_  = ~A299 & A298;
  assign \new_[10564]_  = A301 & A300;
  assign \new_[10565]_  = \new_[10564]_  & \new_[10561]_ ;
  assign \new_[10566]_  = \new_[10565]_  & \new_[10558]_ ;
  assign \new_[10570]_  = A201 & ~A200;
  assign \new_[10571]_  = A199 & \new_[10570]_ ;
  assign \new_[10574]_  = ~A232 & A202;
  assign \new_[10577]_  = A234 & A233;
  assign \new_[10578]_  = \new_[10577]_  & \new_[10574]_ ;
  assign \new_[10579]_  = \new_[10578]_  & \new_[10571]_ ;
  assign \new_[10583]_  = ~A266 & ~A265;
  assign \new_[10584]_  = A235 & \new_[10583]_ ;
  assign \new_[10587]_  = ~A299 & A298;
  assign \new_[10590]_  = ~A302 & A300;
  assign \new_[10591]_  = \new_[10590]_  & \new_[10587]_ ;
  assign \new_[10592]_  = \new_[10591]_  & \new_[10584]_ ;
  assign \new_[10596]_  = A201 & ~A200;
  assign \new_[10597]_  = A199 & \new_[10596]_ ;
  assign \new_[10600]_  = ~A232 & A202;
  assign \new_[10603]_  = A234 & A233;
  assign \new_[10604]_  = \new_[10603]_  & \new_[10600]_ ;
  assign \new_[10605]_  = \new_[10604]_  & \new_[10597]_ ;
  assign \new_[10609]_  = ~A266 & ~A265;
  assign \new_[10610]_  = A235 & \new_[10609]_ ;
  assign \new_[10613]_  = A299 & ~A298;
  assign \new_[10616]_  = A301 & A300;
  assign \new_[10617]_  = \new_[10616]_  & \new_[10613]_ ;
  assign \new_[10618]_  = \new_[10617]_  & \new_[10610]_ ;
  assign \new_[10622]_  = A201 & ~A200;
  assign \new_[10623]_  = A199 & \new_[10622]_ ;
  assign \new_[10626]_  = ~A232 & A202;
  assign \new_[10629]_  = A234 & A233;
  assign \new_[10630]_  = \new_[10629]_  & \new_[10626]_ ;
  assign \new_[10631]_  = \new_[10630]_  & \new_[10623]_ ;
  assign \new_[10635]_  = ~A266 & ~A265;
  assign \new_[10636]_  = A235 & \new_[10635]_ ;
  assign \new_[10639]_  = A299 & ~A298;
  assign \new_[10642]_  = ~A302 & A300;
  assign \new_[10643]_  = \new_[10642]_  & \new_[10639]_ ;
  assign \new_[10644]_  = \new_[10643]_  & \new_[10636]_ ;
  assign \new_[10648]_  = A201 & ~A200;
  assign \new_[10649]_  = A199 & \new_[10648]_ ;
  assign \new_[10652]_  = ~A232 & A202;
  assign \new_[10655]_  = A234 & A233;
  assign \new_[10656]_  = \new_[10655]_  & \new_[10652]_ ;
  assign \new_[10657]_  = \new_[10656]_  & \new_[10649]_ ;
  assign \new_[10661]_  = A268 & ~A267;
  assign \new_[10662]_  = ~A236 & \new_[10661]_ ;
  assign \new_[10665]_  = ~A299 & A298;
  assign \new_[10668]_  = A301 & A300;
  assign \new_[10669]_  = \new_[10668]_  & \new_[10665]_ ;
  assign \new_[10670]_  = \new_[10669]_  & \new_[10662]_ ;
  assign \new_[10674]_  = A201 & ~A200;
  assign \new_[10675]_  = A199 & \new_[10674]_ ;
  assign \new_[10678]_  = ~A232 & A202;
  assign \new_[10681]_  = A234 & A233;
  assign \new_[10682]_  = \new_[10681]_  & \new_[10678]_ ;
  assign \new_[10683]_  = \new_[10682]_  & \new_[10675]_ ;
  assign \new_[10687]_  = A268 & ~A267;
  assign \new_[10688]_  = ~A236 & \new_[10687]_ ;
  assign \new_[10691]_  = ~A299 & A298;
  assign \new_[10694]_  = ~A302 & A300;
  assign \new_[10695]_  = \new_[10694]_  & \new_[10691]_ ;
  assign \new_[10696]_  = \new_[10695]_  & \new_[10688]_ ;
  assign \new_[10700]_  = A201 & ~A200;
  assign \new_[10701]_  = A199 & \new_[10700]_ ;
  assign \new_[10704]_  = ~A232 & A202;
  assign \new_[10707]_  = A234 & A233;
  assign \new_[10708]_  = \new_[10707]_  & \new_[10704]_ ;
  assign \new_[10709]_  = \new_[10708]_  & \new_[10701]_ ;
  assign \new_[10713]_  = A268 & ~A267;
  assign \new_[10714]_  = ~A236 & \new_[10713]_ ;
  assign \new_[10717]_  = A299 & ~A298;
  assign \new_[10720]_  = A301 & A300;
  assign \new_[10721]_  = \new_[10720]_  & \new_[10717]_ ;
  assign \new_[10722]_  = \new_[10721]_  & \new_[10714]_ ;
  assign \new_[10726]_  = A201 & ~A200;
  assign \new_[10727]_  = A199 & \new_[10726]_ ;
  assign \new_[10730]_  = ~A232 & A202;
  assign \new_[10733]_  = A234 & A233;
  assign \new_[10734]_  = \new_[10733]_  & \new_[10730]_ ;
  assign \new_[10735]_  = \new_[10734]_  & \new_[10727]_ ;
  assign \new_[10739]_  = A268 & ~A267;
  assign \new_[10740]_  = ~A236 & \new_[10739]_ ;
  assign \new_[10743]_  = A299 & ~A298;
  assign \new_[10746]_  = ~A302 & A300;
  assign \new_[10747]_  = \new_[10746]_  & \new_[10743]_ ;
  assign \new_[10748]_  = \new_[10747]_  & \new_[10740]_ ;
  assign \new_[10752]_  = A201 & ~A200;
  assign \new_[10753]_  = A199 & \new_[10752]_ ;
  assign \new_[10756]_  = ~A232 & A202;
  assign \new_[10759]_  = A234 & A233;
  assign \new_[10760]_  = \new_[10759]_  & \new_[10756]_ ;
  assign \new_[10761]_  = \new_[10760]_  & \new_[10753]_ ;
  assign \new_[10765]_  = ~A269 & ~A267;
  assign \new_[10766]_  = ~A236 & \new_[10765]_ ;
  assign \new_[10769]_  = ~A299 & A298;
  assign \new_[10772]_  = A301 & A300;
  assign \new_[10773]_  = \new_[10772]_  & \new_[10769]_ ;
  assign \new_[10774]_  = \new_[10773]_  & \new_[10766]_ ;
  assign \new_[10778]_  = A201 & ~A200;
  assign \new_[10779]_  = A199 & \new_[10778]_ ;
  assign \new_[10782]_  = ~A232 & A202;
  assign \new_[10785]_  = A234 & A233;
  assign \new_[10786]_  = \new_[10785]_  & \new_[10782]_ ;
  assign \new_[10787]_  = \new_[10786]_  & \new_[10779]_ ;
  assign \new_[10791]_  = ~A269 & ~A267;
  assign \new_[10792]_  = ~A236 & \new_[10791]_ ;
  assign \new_[10795]_  = ~A299 & A298;
  assign \new_[10798]_  = ~A302 & A300;
  assign \new_[10799]_  = \new_[10798]_  & \new_[10795]_ ;
  assign \new_[10800]_  = \new_[10799]_  & \new_[10792]_ ;
  assign \new_[10804]_  = A201 & ~A200;
  assign \new_[10805]_  = A199 & \new_[10804]_ ;
  assign \new_[10808]_  = ~A232 & A202;
  assign \new_[10811]_  = A234 & A233;
  assign \new_[10812]_  = \new_[10811]_  & \new_[10808]_ ;
  assign \new_[10813]_  = \new_[10812]_  & \new_[10805]_ ;
  assign \new_[10817]_  = ~A269 & ~A267;
  assign \new_[10818]_  = ~A236 & \new_[10817]_ ;
  assign \new_[10821]_  = A299 & ~A298;
  assign \new_[10824]_  = A301 & A300;
  assign \new_[10825]_  = \new_[10824]_  & \new_[10821]_ ;
  assign \new_[10826]_  = \new_[10825]_  & \new_[10818]_ ;
  assign \new_[10830]_  = A201 & ~A200;
  assign \new_[10831]_  = A199 & \new_[10830]_ ;
  assign \new_[10834]_  = ~A232 & A202;
  assign \new_[10837]_  = A234 & A233;
  assign \new_[10838]_  = \new_[10837]_  & \new_[10834]_ ;
  assign \new_[10839]_  = \new_[10838]_  & \new_[10831]_ ;
  assign \new_[10843]_  = ~A269 & ~A267;
  assign \new_[10844]_  = ~A236 & \new_[10843]_ ;
  assign \new_[10847]_  = A299 & ~A298;
  assign \new_[10850]_  = ~A302 & A300;
  assign \new_[10851]_  = \new_[10850]_  & \new_[10847]_ ;
  assign \new_[10852]_  = \new_[10851]_  & \new_[10844]_ ;
  assign \new_[10856]_  = A201 & ~A200;
  assign \new_[10857]_  = A199 & \new_[10856]_ ;
  assign \new_[10860]_  = ~A232 & A202;
  assign \new_[10863]_  = A234 & A233;
  assign \new_[10864]_  = \new_[10863]_  & \new_[10860]_ ;
  assign \new_[10865]_  = \new_[10864]_  & \new_[10857]_ ;
  assign \new_[10869]_  = A266 & A265;
  assign \new_[10870]_  = ~A236 & \new_[10869]_ ;
  assign \new_[10873]_  = ~A299 & A298;
  assign \new_[10876]_  = A301 & A300;
  assign \new_[10877]_  = \new_[10876]_  & \new_[10873]_ ;
  assign \new_[10878]_  = \new_[10877]_  & \new_[10870]_ ;
  assign \new_[10882]_  = A201 & ~A200;
  assign \new_[10883]_  = A199 & \new_[10882]_ ;
  assign \new_[10886]_  = ~A232 & A202;
  assign \new_[10889]_  = A234 & A233;
  assign \new_[10890]_  = \new_[10889]_  & \new_[10886]_ ;
  assign \new_[10891]_  = \new_[10890]_  & \new_[10883]_ ;
  assign \new_[10895]_  = A266 & A265;
  assign \new_[10896]_  = ~A236 & \new_[10895]_ ;
  assign \new_[10899]_  = ~A299 & A298;
  assign \new_[10902]_  = ~A302 & A300;
  assign \new_[10903]_  = \new_[10902]_  & \new_[10899]_ ;
  assign \new_[10904]_  = \new_[10903]_  & \new_[10896]_ ;
  assign \new_[10908]_  = A201 & ~A200;
  assign \new_[10909]_  = A199 & \new_[10908]_ ;
  assign \new_[10912]_  = ~A232 & A202;
  assign \new_[10915]_  = A234 & A233;
  assign \new_[10916]_  = \new_[10915]_  & \new_[10912]_ ;
  assign \new_[10917]_  = \new_[10916]_  & \new_[10909]_ ;
  assign \new_[10921]_  = A266 & A265;
  assign \new_[10922]_  = ~A236 & \new_[10921]_ ;
  assign \new_[10925]_  = A299 & ~A298;
  assign \new_[10928]_  = A301 & A300;
  assign \new_[10929]_  = \new_[10928]_  & \new_[10925]_ ;
  assign \new_[10930]_  = \new_[10929]_  & \new_[10922]_ ;
  assign \new_[10934]_  = A201 & ~A200;
  assign \new_[10935]_  = A199 & \new_[10934]_ ;
  assign \new_[10938]_  = ~A232 & A202;
  assign \new_[10941]_  = A234 & A233;
  assign \new_[10942]_  = \new_[10941]_  & \new_[10938]_ ;
  assign \new_[10943]_  = \new_[10942]_  & \new_[10935]_ ;
  assign \new_[10947]_  = A266 & A265;
  assign \new_[10948]_  = ~A236 & \new_[10947]_ ;
  assign \new_[10951]_  = A299 & ~A298;
  assign \new_[10954]_  = ~A302 & A300;
  assign \new_[10955]_  = \new_[10954]_  & \new_[10951]_ ;
  assign \new_[10956]_  = \new_[10955]_  & \new_[10948]_ ;
  assign \new_[10960]_  = A201 & ~A200;
  assign \new_[10961]_  = A199 & \new_[10960]_ ;
  assign \new_[10964]_  = ~A232 & A202;
  assign \new_[10967]_  = A234 & A233;
  assign \new_[10968]_  = \new_[10967]_  & \new_[10964]_ ;
  assign \new_[10969]_  = \new_[10968]_  & \new_[10961]_ ;
  assign \new_[10973]_  = ~A266 & ~A265;
  assign \new_[10974]_  = ~A236 & \new_[10973]_ ;
  assign \new_[10977]_  = ~A299 & A298;
  assign \new_[10980]_  = A301 & A300;
  assign \new_[10981]_  = \new_[10980]_  & \new_[10977]_ ;
  assign \new_[10982]_  = \new_[10981]_  & \new_[10974]_ ;
  assign \new_[10986]_  = A201 & ~A200;
  assign \new_[10987]_  = A199 & \new_[10986]_ ;
  assign \new_[10990]_  = ~A232 & A202;
  assign \new_[10993]_  = A234 & A233;
  assign \new_[10994]_  = \new_[10993]_  & \new_[10990]_ ;
  assign \new_[10995]_  = \new_[10994]_  & \new_[10987]_ ;
  assign \new_[10999]_  = ~A266 & ~A265;
  assign \new_[11000]_  = ~A236 & \new_[10999]_ ;
  assign \new_[11003]_  = ~A299 & A298;
  assign \new_[11006]_  = ~A302 & A300;
  assign \new_[11007]_  = \new_[11006]_  & \new_[11003]_ ;
  assign \new_[11008]_  = \new_[11007]_  & \new_[11000]_ ;
  assign \new_[11012]_  = A201 & ~A200;
  assign \new_[11013]_  = A199 & \new_[11012]_ ;
  assign \new_[11016]_  = ~A232 & A202;
  assign \new_[11019]_  = A234 & A233;
  assign \new_[11020]_  = \new_[11019]_  & \new_[11016]_ ;
  assign \new_[11021]_  = \new_[11020]_  & \new_[11013]_ ;
  assign \new_[11025]_  = ~A266 & ~A265;
  assign \new_[11026]_  = ~A236 & \new_[11025]_ ;
  assign \new_[11029]_  = A299 & ~A298;
  assign \new_[11032]_  = A301 & A300;
  assign \new_[11033]_  = \new_[11032]_  & \new_[11029]_ ;
  assign \new_[11034]_  = \new_[11033]_  & \new_[11026]_ ;
  assign \new_[11038]_  = A201 & ~A200;
  assign \new_[11039]_  = A199 & \new_[11038]_ ;
  assign \new_[11042]_  = ~A232 & A202;
  assign \new_[11045]_  = A234 & A233;
  assign \new_[11046]_  = \new_[11045]_  & \new_[11042]_ ;
  assign \new_[11047]_  = \new_[11046]_  & \new_[11039]_ ;
  assign \new_[11051]_  = ~A266 & ~A265;
  assign \new_[11052]_  = ~A236 & \new_[11051]_ ;
  assign \new_[11055]_  = A299 & ~A298;
  assign \new_[11058]_  = ~A302 & A300;
  assign \new_[11059]_  = \new_[11058]_  & \new_[11055]_ ;
  assign \new_[11060]_  = \new_[11059]_  & \new_[11052]_ ;
  assign \new_[11064]_  = A201 & ~A200;
  assign \new_[11065]_  = A199 & \new_[11064]_ ;
  assign \new_[11068]_  = A232 & A202;
  assign \new_[11071]_  = A234 & ~A233;
  assign \new_[11072]_  = \new_[11071]_  & \new_[11068]_ ;
  assign \new_[11073]_  = \new_[11072]_  & \new_[11065]_ ;
  assign \new_[11077]_  = A268 & ~A267;
  assign \new_[11078]_  = A235 & \new_[11077]_ ;
  assign \new_[11081]_  = ~A299 & A298;
  assign \new_[11084]_  = A301 & A300;
  assign \new_[11085]_  = \new_[11084]_  & \new_[11081]_ ;
  assign \new_[11086]_  = \new_[11085]_  & \new_[11078]_ ;
  assign \new_[11090]_  = A201 & ~A200;
  assign \new_[11091]_  = A199 & \new_[11090]_ ;
  assign \new_[11094]_  = A232 & A202;
  assign \new_[11097]_  = A234 & ~A233;
  assign \new_[11098]_  = \new_[11097]_  & \new_[11094]_ ;
  assign \new_[11099]_  = \new_[11098]_  & \new_[11091]_ ;
  assign \new_[11103]_  = A268 & ~A267;
  assign \new_[11104]_  = A235 & \new_[11103]_ ;
  assign \new_[11107]_  = ~A299 & A298;
  assign \new_[11110]_  = ~A302 & A300;
  assign \new_[11111]_  = \new_[11110]_  & \new_[11107]_ ;
  assign \new_[11112]_  = \new_[11111]_  & \new_[11104]_ ;
  assign \new_[11116]_  = A201 & ~A200;
  assign \new_[11117]_  = A199 & \new_[11116]_ ;
  assign \new_[11120]_  = A232 & A202;
  assign \new_[11123]_  = A234 & ~A233;
  assign \new_[11124]_  = \new_[11123]_  & \new_[11120]_ ;
  assign \new_[11125]_  = \new_[11124]_  & \new_[11117]_ ;
  assign \new_[11129]_  = A268 & ~A267;
  assign \new_[11130]_  = A235 & \new_[11129]_ ;
  assign \new_[11133]_  = A299 & ~A298;
  assign \new_[11136]_  = A301 & A300;
  assign \new_[11137]_  = \new_[11136]_  & \new_[11133]_ ;
  assign \new_[11138]_  = \new_[11137]_  & \new_[11130]_ ;
  assign \new_[11142]_  = A201 & ~A200;
  assign \new_[11143]_  = A199 & \new_[11142]_ ;
  assign \new_[11146]_  = A232 & A202;
  assign \new_[11149]_  = A234 & ~A233;
  assign \new_[11150]_  = \new_[11149]_  & \new_[11146]_ ;
  assign \new_[11151]_  = \new_[11150]_  & \new_[11143]_ ;
  assign \new_[11155]_  = A268 & ~A267;
  assign \new_[11156]_  = A235 & \new_[11155]_ ;
  assign \new_[11159]_  = A299 & ~A298;
  assign \new_[11162]_  = ~A302 & A300;
  assign \new_[11163]_  = \new_[11162]_  & \new_[11159]_ ;
  assign \new_[11164]_  = \new_[11163]_  & \new_[11156]_ ;
  assign \new_[11168]_  = A201 & ~A200;
  assign \new_[11169]_  = A199 & \new_[11168]_ ;
  assign \new_[11172]_  = A232 & A202;
  assign \new_[11175]_  = A234 & ~A233;
  assign \new_[11176]_  = \new_[11175]_  & \new_[11172]_ ;
  assign \new_[11177]_  = \new_[11176]_  & \new_[11169]_ ;
  assign \new_[11181]_  = ~A269 & ~A267;
  assign \new_[11182]_  = A235 & \new_[11181]_ ;
  assign \new_[11185]_  = ~A299 & A298;
  assign \new_[11188]_  = A301 & A300;
  assign \new_[11189]_  = \new_[11188]_  & \new_[11185]_ ;
  assign \new_[11190]_  = \new_[11189]_  & \new_[11182]_ ;
  assign \new_[11194]_  = A201 & ~A200;
  assign \new_[11195]_  = A199 & \new_[11194]_ ;
  assign \new_[11198]_  = A232 & A202;
  assign \new_[11201]_  = A234 & ~A233;
  assign \new_[11202]_  = \new_[11201]_  & \new_[11198]_ ;
  assign \new_[11203]_  = \new_[11202]_  & \new_[11195]_ ;
  assign \new_[11207]_  = ~A269 & ~A267;
  assign \new_[11208]_  = A235 & \new_[11207]_ ;
  assign \new_[11211]_  = ~A299 & A298;
  assign \new_[11214]_  = ~A302 & A300;
  assign \new_[11215]_  = \new_[11214]_  & \new_[11211]_ ;
  assign \new_[11216]_  = \new_[11215]_  & \new_[11208]_ ;
  assign \new_[11220]_  = A201 & ~A200;
  assign \new_[11221]_  = A199 & \new_[11220]_ ;
  assign \new_[11224]_  = A232 & A202;
  assign \new_[11227]_  = A234 & ~A233;
  assign \new_[11228]_  = \new_[11227]_  & \new_[11224]_ ;
  assign \new_[11229]_  = \new_[11228]_  & \new_[11221]_ ;
  assign \new_[11233]_  = ~A269 & ~A267;
  assign \new_[11234]_  = A235 & \new_[11233]_ ;
  assign \new_[11237]_  = A299 & ~A298;
  assign \new_[11240]_  = A301 & A300;
  assign \new_[11241]_  = \new_[11240]_  & \new_[11237]_ ;
  assign \new_[11242]_  = \new_[11241]_  & \new_[11234]_ ;
  assign \new_[11246]_  = A201 & ~A200;
  assign \new_[11247]_  = A199 & \new_[11246]_ ;
  assign \new_[11250]_  = A232 & A202;
  assign \new_[11253]_  = A234 & ~A233;
  assign \new_[11254]_  = \new_[11253]_  & \new_[11250]_ ;
  assign \new_[11255]_  = \new_[11254]_  & \new_[11247]_ ;
  assign \new_[11259]_  = ~A269 & ~A267;
  assign \new_[11260]_  = A235 & \new_[11259]_ ;
  assign \new_[11263]_  = A299 & ~A298;
  assign \new_[11266]_  = ~A302 & A300;
  assign \new_[11267]_  = \new_[11266]_  & \new_[11263]_ ;
  assign \new_[11268]_  = \new_[11267]_  & \new_[11260]_ ;
  assign \new_[11272]_  = A201 & ~A200;
  assign \new_[11273]_  = A199 & \new_[11272]_ ;
  assign \new_[11276]_  = A232 & A202;
  assign \new_[11279]_  = A234 & ~A233;
  assign \new_[11280]_  = \new_[11279]_  & \new_[11276]_ ;
  assign \new_[11281]_  = \new_[11280]_  & \new_[11273]_ ;
  assign \new_[11285]_  = A266 & A265;
  assign \new_[11286]_  = A235 & \new_[11285]_ ;
  assign \new_[11289]_  = ~A299 & A298;
  assign \new_[11292]_  = A301 & A300;
  assign \new_[11293]_  = \new_[11292]_  & \new_[11289]_ ;
  assign \new_[11294]_  = \new_[11293]_  & \new_[11286]_ ;
  assign \new_[11298]_  = A201 & ~A200;
  assign \new_[11299]_  = A199 & \new_[11298]_ ;
  assign \new_[11302]_  = A232 & A202;
  assign \new_[11305]_  = A234 & ~A233;
  assign \new_[11306]_  = \new_[11305]_  & \new_[11302]_ ;
  assign \new_[11307]_  = \new_[11306]_  & \new_[11299]_ ;
  assign \new_[11311]_  = A266 & A265;
  assign \new_[11312]_  = A235 & \new_[11311]_ ;
  assign \new_[11315]_  = ~A299 & A298;
  assign \new_[11318]_  = ~A302 & A300;
  assign \new_[11319]_  = \new_[11318]_  & \new_[11315]_ ;
  assign \new_[11320]_  = \new_[11319]_  & \new_[11312]_ ;
  assign \new_[11324]_  = A201 & ~A200;
  assign \new_[11325]_  = A199 & \new_[11324]_ ;
  assign \new_[11328]_  = A232 & A202;
  assign \new_[11331]_  = A234 & ~A233;
  assign \new_[11332]_  = \new_[11331]_  & \new_[11328]_ ;
  assign \new_[11333]_  = \new_[11332]_  & \new_[11325]_ ;
  assign \new_[11337]_  = A266 & A265;
  assign \new_[11338]_  = A235 & \new_[11337]_ ;
  assign \new_[11341]_  = A299 & ~A298;
  assign \new_[11344]_  = A301 & A300;
  assign \new_[11345]_  = \new_[11344]_  & \new_[11341]_ ;
  assign \new_[11346]_  = \new_[11345]_  & \new_[11338]_ ;
  assign \new_[11350]_  = A201 & ~A200;
  assign \new_[11351]_  = A199 & \new_[11350]_ ;
  assign \new_[11354]_  = A232 & A202;
  assign \new_[11357]_  = A234 & ~A233;
  assign \new_[11358]_  = \new_[11357]_  & \new_[11354]_ ;
  assign \new_[11359]_  = \new_[11358]_  & \new_[11351]_ ;
  assign \new_[11363]_  = A266 & A265;
  assign \new_[11364]_  = A235 & \new_[11363]_ ;
  assign \new_[11367]_  = A299 & ~A298;
  assign \new_[11370]_  = ~A302 & A300;
  assign \new_[11371]_  = \new_[11370]_  & \new_[11367]_ ;
  assign \new_[11372]_  = \new_[11371]_  & \new_[11364]_ ;
  assign \new_[11376]_  = A201 & ~A200;
  assign \new_[11377]_  = A199 & \new_[11376]_ ;
  assign \new_[11380]_  = A232 & A202;
  assign \new_[11383]_  = A234 & ~A233;
  assign \new_[11384]_  = \new_[11383]_  & \new_[11380]_ ;
  assign \new_[11385]_  = \new_[11384]_  & \new_[11377]_ ;
  assign \new_[11389]_  = ~A266 & ~A265;
  assign \new_[11390]_  = A235 & \new_[11389]_ ;
  assign \new_[11393]_  = ~A299 & A298;
  assign \new_[11396]_  = A301 & A300;
  assign \new_[11397]_  = \new_[11396]_  & \new_[11393]_ ;
  assign \new_[11398]_  = \new_[11397]_  & \new_[11390]_ ;
  assign \new_[11402]_  = A201 & ~A200;
  assign \new_[11403]_  = A199 & \new_[11402]_ ;
  assign \new_[11406]_  = A232 & A202;
  assign \new_[11409]_  = A234 & ~A233;
  assign \new_[11410]_  = \new_[11409]_  & \new_[11406]_ ;
  assign \new_[11411]_  = \new_[11410]_  & \new_[11403]_ ;
  assign \new_[11415]_  = ~A266 & ~A265;
  assign \new_[11416]_  = A235 & \new_[11415]_ ;
  assign \new_[11419]_  = ~A299 & A298;
  assign \new_[11422]_  = ~A302 & A300;
  assign \new_[11423]_  = \new_[11422]_  & \new_[11419]_ ;
  assign \new_[11424]_  = \new_[11423]_  & \new_[11416]_ ;
  assign \new_[11428]_  = A201 & ~A200;
  assign \new_[11429]_  = A199 & \new_[11428]_ ;
  assign \new_[11432]_  = A232 & A202;
  assign \new_[11435]_  = A234 & ~A233;
  assign \new_[11436]_  = \new_[11435]_  & \new_[11432]_ ;
  assign \new_[11437]_  = \new_[11436]_  & \new_[11429]_ ;
  assign \new_[11441]_  = ~A266 & ~A265;
  assign \new_[11442]_  = A235 & \new_[11441]_ ;
  assign \new_[11445]_  = A299 & ~A298;
  assign \new_[11448]_  = A301 & A300;
  assign \new_[11449]_  = \new_[11448]_  & \new_[11445]_ ;
  assign \new_[11450]_  = \new_[11449]_  & \new_[11442]_ ;
  assign \new_[11454]_  = A201 & ~A200;
  assign \new_[11455]_  = A199 & \new_[11454]_ ;
  assign \new_[11458]_  = A232 & A202;
  assign \new_[11461]_  = A234 & ~A233;
  assign \new_[11462]_  = \new_[11461]_  & \new_[11458]_ ;
  assign \new_[11463]_  = \new_[11462]_  & \new_[11455]_ ;
  assign \new_[11467]_  = ~A266 & ~A265;
  assign \new_[11468]_  = A235 & \new_[11467]_ ;
  assign \new_[11471]_  = A299 & ~A298;
  assign \new_[11474]_  = ~A302 & A300;
  assign \new_[11475]_  = \new_[11474]_  & \new_[11471]_ ;
  assign \new_[11476]_  = \new_[11475]_  & \new_[11468]_ ;
  assign \new_[11480]_  = A201 & ~A200;
  assign \new_[11481]_  = A199 & \new_[11480]_ ;
  assign \new_[11484]_  = A232 & A202;
  assign \new_[11487]_  = A234 & ~A233;
  assign \new_[11488]_  = \new_[11487]_  & \new_[11484]_ ;
  assign \new_[11489]_  = \new_[11488]_  & \new_[11481]_ ;
  assign \new_[11493]_  = A268 & ~A267;
  assign \new_[11494]_  = ~A236 & \new_[11493]_ ;
  assign \new_[11497]_  = ~A299 & A298;
  assign \new_[11500]_  = A301 & A300;
  assign \new_[11501]_  = \new_[11500]_  & \new_[11497]_ ;
  assign \new_[11502]_  = \new_[11501]_  & \new_[11494]_ ;
  assign \new_[11506]_  = A201 & ~A200;
  assign \new_[11507]_  = A199 & \new_[11506]_ ;
  assign \new_[11510]_  = A232 & A202;
  assign \new_[11513]_  = A234 & ~A233;
  assign \new_[11514]_  = \new_[11513]_  & \new_[11510]_ ;
  assign \new_[11515]_  = \new_[11514]_  & \new_[11507]_ ;
  assign \new_[11519]_  = A268 & ~A267;
  assign \new_[11520]_  = ~A236 & \new_[11519]_ ;
  assign \new_[11523]_  = ~A299 & A298;
  assign \new_[11526]_  = ~A302 & A300;
  assign \new_[11527]_  = \new_[11526]_  & \new_[11523]_ ;
  assign \new_[11528]_  = \new_[11527]_  & \new_[11520]_ ;
  assign \new_[11532]_  = A201 & ~A200;
  assign \new_[11533]_  = A199 & \new_[11532]_ ;
  assign \new_[11536]_  = A232 & A202;
  assign \new_[11539]_  = A234 & ~A233;
  assign \new_[11540]_  = \new_[11539]_  & \new_[11536]_ ;
  assign \new_[11541]_  = \new_[11540]_  & \new_[11533]_ ;
  assign \new_[11545]_  = A268 & ~A267;
  assign \new_[11546]_  = ~A236 & \new_[11545]_ ;
  assign \new_[11549]_  = A299 & ~A298;
  assign \new_[11552]_  = A301 & A300;
  assign \new_[11553]_  = \new_[11552]_  & \new_[11549]_ ;
  assign \new_[11554]_  = \new_[11553]_  & \new_[11546]_ ;
  assign \new_[11558]_  = A201 & ~A200;
  assign \new_[11559]_  = A199 & \new_[11558]_ ;
  assign \new_[11562]_  = A232 & A202;
  assign \new_[11565]_  = A234 & ~A233;
  assign \new_[11566]_  = \new_[11565]_  & \new_[11562]_ ;
  assign \new_[11567]_  = \new_[11566]_  & \new_[11559]_ ;
  assign \new_[11571]_  = A268 & ~A267;
  assign \new_[11572]_  = ~A236 & \new_[11571]_ ;
  assign \new_[11575]_  = A299 & ~A298;
  assign \new_[11578]_  = ~A302 & A300;
  assign \new_[11579]_  = \new_[11578]_  & \new_[11575]_ ;
  assign \new_[11580]_  = \new_[11579]_  & \new_[11572]_ ;
  assign \new_[11584]_  = A201 & ~A200;
  assign \new_[11585]_  = A199 & \new_[11584]_ ;
  assign \new_[11588]_  = A232 & A202;
  assign \new_[11591]_  = A234 & ~A233;
  assign \new_[11592]_  = \new_[11591]_  & \new_[11588]_ ;
  assign \new_[11593]_  = \new_[11592]_  & \new_[11585]_ ;
  assign \new_[11597]_  = ~A269 & ~A267;
  assign \new_[11598]_  = ~A236 & \new_[11597]_ ;
  assign \new_[11601]_  = ~A299 & A298;
  assign \new_[11604]_  = A301 & A300;
  assign \new_[11605]_  = \new_[11604]_  & \new_[11601]_ ;
  assign \new_[11606]_  = \new_[11605]_  & \new_[11598]_ ;
  assign \new_[11610]_  = A201 & ~A200;
  assign \new_[11611]_  = A199 & \new_[11610]_ ;
  assign \new_[11614]_  = A232 & A202;
  assign \new_[11617]_  = A234 & ~A233;
  assign \new_[11618]_  = \new_[11617]_  & \new_[11614]_ ;
  assign \new_[11619]_  = \new_[11618]_  & \new_[11611]_ ;
  assign \new_[11623]_  = ~A269 & ~A267;
  assign \new_[11624]_  = ~A236 & \new_[11623]_ ;
  assign \new_[11627]_  = ~A299 & A298;
  assign \new_[11630]_  = ~A302 & A300;
  assign \new_[11631]_  = \new_[11630]_  & \new_[11627]_ ;
  assign \new_[11632]_  = \new_[11631]_  & \new_[11624]_ ;
  assign \new_[11636]_  = A201 & ~A200;
  assign \new_[11637]_  = A199 & \new_[11636]_ ;
  assign \new_[11640]_  = A232 & A202;
  assign \new_[11643]_  = A234 & ~A233;
  assign \new_[11644]_  = \new_[11643]_  & \new_[11640]_ ;
  assign \new_[11645]_  = \new_[11644]_  & \new_[11637]_ ;
  assign \new_[11649]_  = ~A269 & ~A267;
  assign \new_[11650]_  = ~A236 & \new_[11649]_ ;
  assign \new_[11653]_  = A299 & ~A298;
  assign \new_[11656]_  = A301 & A300;
  assign \new_[11657]_  = \new_[11656]_  & \new_[11653]_ ;
  assign \new_[11658]_  = \new_[11657]_  & \new_[11650]_ ;
  assign \new_[11662]_  = A201 & ~A200;
  assign \new_[11663]_  = A199 & \new_[11662]_ ;
  assign \new_[11666]_  = A232 & A202;
  assign \new_[11669]_  = A234 & ~A233;
  assign \new_[11670]_  = \new_[11669]_  & \new_[11666]_ ;
  assign \new_[11671]_  = \new_[11670]_  & \new_[11663]_ ;
  assign \new_[11675]_  = ~A269 & ~A267;
  assign \new_[11676]_  = ~A236 & \new_[11675]_ ;
  assign \new_[11679]_  = A299 & ~A298;
  assign \new_[11682]_  = ~A302 & A300;
  assign \new_[11683]_  = \new_[11682]_  & \new_[11679]_ ;
  assign \new_[11684]_  = \new_[11683]_  & \new_[11676]_ ;
  assign \new_[11688]_  = A201 & ~A200;
  assign \new_[11689]_  = A199 & \new_[11688]_ ;
  assign \new_[11692]_  = A232 & A202;
  assign \new_[11695]_  = A234 & ~A233;
  assign \new_[11696]_  = \new_[11695]_  & \new_[11692]_ ;
  assign \new_[11697]_  = \new_[11696]_  & \new_[11689]_ ;
  assign \new_[11701]_  = A266 & A265;
  assign \new_[11702]_  = ~A236 & \new_[11701]_ ;
  assign \new_[11705]_  = ~A299 & A298;
  assign \new_[11708]_  = A301 & A300;
  assign \new_[11709]_  = \new_[11708]_  & \new_[11705]_ ;
  assign \new_[11710]_  = \new_[11709]_  & \new_[11702]_ ;
  assign \new_[11714]_  = A201 & ~A200;
  assign \new_[11715]_  = A199 & \new_[11714]_ ;
  assign \new_[11718]_  = A232 & A202;
  assign \new_[11721]_  = A234 & ~A233;
  assign \new_[11722]_  = \new_[11721]_  & \new_[11718]_ ;
  assign \new_[11723]_  = \new_[11722]_  & \new_[11715]_ ;
  assign \new_[11727]_  = A266 & A265;
  assign \new_[11728]_  = ~A236 & \new_[11727]_ ;
  assign \new_[11731]_  = ~A299 & A298;
  assign \new_[11734]_  = ~A302 & A300;
  assign \new_[11735]_  = \new_[11734]_  & \new_[11731]_ ;
  assign \new_[11736]_  = \new_[11735]_  & \new_[11728]_ ;
  assign \new_[11740]_  = A201 & ~A200;
  assign \new_[11741]_  = A199 & \new_[11740]_ ;
  assign \new_[11744]_  = A232 & A202;
  assign \new_[11747]_  = A234 & ~A233;
  assign \new_[11748]_  = \new_[11747]_  & \new_[11744]_ ;
  assign \new_[11749]_  = \new_[11748]_  & \new_[11741]_ ;
  assign \new_[11753]_  = A266 & A265;
  assign \new_[11754]_  = ~A236 & \new_[11753]_ ;
  assign \new_[11757]_  = A299 & ~A298;
  assign \new_[11760]_  = A301 & A300;
  assign \new_[11761]_  = \new_[11760]_  & \new_[11757]_ ;
  assign \new_[11762]_  = \new_[11761]_  & \new_[11754]_ ;
  assign \new_[11766]_  = A201 & ~A200;
  assign \new_[11767]_  = A199 & \new_[11766]_ ;
  assign \new_[11770]_  = A232 & A202;
  assign \new_[11773]_  = A234 & ~A233;
  assign \new_[11774]_  = \new_[11773]_  & \new_[11770]_ ;
  assign \new_[11775]_  = \new_[11774]_  & \new_[11767]_ ;
  assign \new_[11779]_  = A266 & A265;
  assign \new_[11780]_  = ~A236 & \new_[11779]_ ;
  assign \new_[11783]_  = A299 & ~A298;
  assign \new_[11786]_  = ~A302 & A300;
  assign \new_[11787]_  = \new_[11786]_  & \new_[11783]_ ;
  assign \new_[11788]_  = \new_[11787]_  & \new_[11780]_ ;
  assign \new_[11792]_  = A201 & ~A200;
  assign \new_[11793]_  = A199 & \new_[11792]_ ;
  assign \new_[11796]_  = A232 & A202;
  assign \new_[11799]_  = A234 & ~A233;
  assign \new_[11800]_  = \new_[11799]_  & \new_[11796]_ ;
  assign \new_[11801]_  = \new_[11800]_  & \new_[11793]_ ;
  assign \new_[11805]_  = ~A266 & ~A265;
  assign \new_[11806]_  = ~A236 & \new_[11805]_ ;
  assign \new_[11809]_  = ~A299 & A298;
  assign \new_[11812]_  = A301 & A300;
  assign \new_[11813]_  = \new_[11812]_  & \new_[11809]_ ;
  assign \new_[11814]_  = \new_[11813]_  & \new_[11806]_ ;
  assign \new_[11818]_  = A201 & ~A200;
  assign \new_[11819]_  = A199 & \new_[11818]_ ;
  assign \new_[11822]_  = A232 & A202;
  assign \new_[11825]_  = A234 & ~A233;
  assign \new_[11826]_  = \new_[11825]_  & \new_[11822]_ ;
  assign \new_[11827]_  = \new_[11826]_  & \new_[11819]_ ;
  assign \new_[11831]_  = ~A266 & ~A265;
  assign \new_[11832]_  = ~A236 & \new_[11831]_ ;
  assign \new_[11835]_  = ~A299 & A298;
  assign \new_[11838]_  = ~A302 & A300;
  assign \new_[11839]_  = \new_[11838]_  & \new_[11835]_ ;
  assign \new_[11840]_  = \new_[11839]_  & \new_[11832]_ ;
  assign \new_[11844]_  = A201 & ~A200;
  assign \new_[11845]_  = A199 & \new_[11844]_ ;
  assign \new_[11848]_  = A232 & A202;
  assign \new_[11851]_  = A234 & ~A233;
  assign \new_[11852]_  = \new_[11851]_  & \new_[11848]_ ;
  assign \new_[11853]_  = \new_[11852]_  & \new_[11845]_ ;
  assign \new_[11857]_  = ~A266 & ~A265;
  assign \new_[11858]_  = ~A236 & \new_[11857]_ ;
  assign \new_[11861]_  = A299 & ~A298;
  assign \new_[11864]_  = A301 & A300;
  assign \new_[11865]_  = \new_[11864]_  & \new_[11861]_ ;
  assign \new_[11866]_  = \new_[11865]_  & \new_[11858]_ ;
  assign \new_[11870]_  = A201 & ~A200;
  assign \new_[11871]_  = A199 & \new_[11870]_ ;
  assign \new_[11874]_  = A232 & A202;
  assign \new_[11877]_  = A234 & ~A233;
  assign \new_[11878]_  = \new_[11877]_  & \new_[11874]_ ;
  assign \new_[11879]_  = \new_[11878]_  & \new_[11871]_ ;
  assign \new_[11883]_  = ~A266 & ~A265;
  assign \new_[11884]_  = ~A236 & \new_[11883]_ ;
  assign \new_[11887]_  = A299 & ~A298;
  assign \new_[11890]_  = ~A302 & A300;
  assign \new_[11891]_  = \new_[11890]_  & \new_[11887]_ ;
  assign \new_[11892]_  = \new_[11891]_  & \new_[11884]_ ;
  assign \new_[11896]_  = A201 & ~A200;
  assign \new_[11897]_  = A199 & \new_[11896]_ ;
  assign \new_[11900]_  = ~A232 & ~A203;
  assign \new_[11903]_  = A234 & A233;
  assign \new_[11904]_  = \new_[11903]_  & \new_[11900]_ ;
  assign \new_[11905]_  = \new_[11904]_  & \new_[11897]_ ;
  assign \new_[11909]_  = A268 & ~A267;
  assign \new_[11910]_  = A235 & \new_[11909]_ ;
  assign \new_[11913]_  = ~A299 & A298;
  assign \new_[11916]_  = A301 & A300;
  assign \new_[11917]_  = \new_[11916]_  & \new_[11913]_ ;
  assign \new_[11918]_  = \new_[11917]_  & \new_[11910]_ ;
  assign \new_[11922]_  = A201 & ~A200;
  assign \new_[11923]_  = A199 & \new_[11922]_ ;
  assign \new_[11926]_  = ~A232 & ~A203;
  assign \new_[11929]_  = A234 & A233;
  assign \new_[11930]_  = \new_[11929]_  & \new_[11926]_ ;
  assign \new_[11931]_  = \new_[11930]_  & \new_[11923]_ ;
  assign \new_[11935]_  = A268 & ~A267;
  assign \new_[11936]_  = A235 & \new_[11935]_ ;
  assign \new_[11939]_  = ~A299 & A298;
  assign \new_[11942]_  = ~A302 & A300;
  assign \new_[11943]_  = \new_[11942]_  & \new_[11939]_ ;
  assign \new_[11944]_  = \new_[11943]_  & \new_[11936]_ ;
  assign \new_[11948]_  = A201 & ~A200;
  assign \new_[11949]_  = A199 & \new_[11948]_ ;
  assign \new_[11952]_  = ~A232 & ~A203;
  assign \new_[11955]_  = A234 & A233;
  assign \new_[11956]_  = \new_[11955]_  & \new_[11952]_ ;
  assign \new_[11957]_  = \new_[11956]_  & \new_[11949]_ ;
  assign \new_[11961]_  = A268 & ~A267;
  assign \new_[11962]_  = A235 & \new_[11961]_ ;
  assign \new_[11965]_  = A299 & ~A298;
  assign \new_[11968]_  = A301 & A300;
  assign \new_[11969]_  = \new_[11968]_  & \new_[11965]_ ;
  assign \new_[11970]_  = \new_[11969]_  & \new_[11962]_ ;
  assign \new_[11974]_  = A201 & ~A200;
  assign \new_[11975]_  = A199 & \new_[11974]_ ;
  assign \new_[11978]_  = ~A232 & ~A203;
  assign \new_[11981]_  = A234 & A233;
  assign \new_[11982]_  = \new_[11981]_  & \new_[11978]_ ;
  assign \new_[11983]_  = \new_[11982]_  & \new_[11975]_ ;
  assign \new_[11987]_  = A268 & ~A267;
  assign \new_[11988]_  = A235 & \new_[11987]_ ;
  assign \new_[11991]_  = A299 & ~A298;
  assign \new_[11994]_  = ~A302 & A300;
  assign \new_[11995]_  = \new_[11994]_  & \new_[11991]_ ;
  assign \new_[11996]_  = \new_[11995]_  & \new_[11988]_ ;
  assign \new_[12000]_  = A201 & ~A200;
  assign \new_[12001]_  = A199 & \new_[12000]_ ;
  assign \new_[12004]_  = ~A232 & ~A203;
  assign \new_[12007]_  = A234 & A233;
  assign \new_[12008]_  = \new_[12007]_  & \new_[12004]_ ;
  assign \new_[12009]_  = \new_[12008]_  & \new_[12001]_ ;
  assign \new_[12013]_  = ~A269 & ~A267;
  assign \new_[12014]_  = A235 & \new_[12013]_ ;
  assign \new_[12017]_  = ~A299 & A298;
  assign \new_[12020]_  = A301 & A300;
  assign \new_[12021]_  = \new_[12020]_  & \new_[12017]_ ;
  assign \new_[12022]_  = \new_[12021]_  & \new_[12014]_ ;
  assign \new_[12026]_  = A201 & ~A200;
  assign \new_[12027]_  = A199 & \new_[12026]_ ;
  assign \new_[12030]_  = ~A232 & ~A203;
  assign \new_[12033]_  = A234 & A233;
  assign \new_[12034]_  = \new_[12033]_  & \new_[12030]_ ;
  assign \new_[12035]_  = \new_[12034]_  & \new_[12027]_ ;
  assign \new_[12039]_  = ~A269 & ~A267;
  assign \new_[12040]_  = A235 & \new_[12039]_ ;
  assign \new_[12043]_  = ~A299 & A298;
  assign \new_[12046]_  = ~A302 & A300;
  assign \new_[12047]_  = \new_[12046]_  & \new_[12043]_ ;
  assign \new_[12048]_  = \new_[12047]_  & \new_[12040]_ ;
  assign \new_[12052]_  = A201 & ~A200;
  assign \new_[12053]_  = A199 & \new_[12052]_ ;
  assign \new_[12056]_  = ~A232 & ~A203;
  assign \new_[12059]_  = A234 & A233;
  assign \new_[12060]_  = \new_[12059]_  & \new_[12056]_ ;
  assign \new_[12061]_  = \new_[12060]_  & \new_[12053]_ ;
  assign \new_[12065]_  = ~A269 & ~A267;
  assign \new_[12066]_  = A235 & \new_[12065]_ ;
  assign \new_[12069]_  = A299 & ~A298;
  assign \new_[12072]_  = A301 & A300;
  assign \new_[12073]_  = \new_[12072]_  & \new_[12069]_ ;
  assign \new_[12074]_  = \new_[12073]_  & \new_[12066]_ ;
  assign \new_[12078]_  = A201 & ~A200;
  assign \new_[12079]_  = A199 & \new_[12078]_ ;
  assign \new_[12082]_  = ~A232 & ~A203;
  assign \new_[12085]_  = A234 & A233;
  assign \new_[12086]_  = \new_[12085]_  & \new_[12082]_ ;
  assign \new_[12087]_  = \new_[12086]_  & \new_[12079]_ ;
  assign \new_[12091]_  = ~A269 & ~A267;
  assign \new_[12092]_  = A235 & \new_[12091]_ ;
  assign \new_[12095]_  = A299 & ~A298;
  assign \new_[12098]_  = ~A302 & A300;
  assign \new_[12099]_  = \new_[12098]_  & \new_[12095]_ ;
  assign \new_[12100]_  = \new_[12099]_  & \new_[12092]_ ;
  assign \new_[12104]_  = A201 & ~A200;
  assign \new_[12105]_  = A199 & \new_[12104]_ ;
  assign \new_[12108]_  = ~A232 & ~A203;
  assign \new_[12111]_  = A234 & A233;
  assign \new_[12112]_  = \new_[12111]_  & \new_[12108]_ ;
  assign \new_[12113]_  = \new_[12112]_  & \new_[12105]_ ;
  assign \new_[12117]_  = A266 & A265;
  assign \new_[12118]_  = A235 & \new_[12117]_ ;
  assign \new_[12121]_  = ~A299 & A298;
  assign \new_[12124]_  = A301 & A300;
  assign \new_[12125]_  = \new_[12124]_  & \new_[12121]_ ;
  assign \new_[12126]_  = \new_[12125]_  & \new_[12118]_ ;
  assign \new_[12130]_  = A201 & ~A200;
  assign \new_[12131]_  = A199 & \new_[12130]_ ;
  assign \new_[12134]_  = ~A232 & ~A203;
  assign \new_[12137]_  = A234 & A233;
  assign \new_[12138]_  = \new_[12137]_  & \new_[12134]_ ;
  assign \new_[12139]_  = \new_[12138]_  & \new_[12131]_ ;
  assign \new_[12143]_  = A266 & A265;
  assign \new_[12144]_  = A235 & \new_[12143]_ ;
  assign \new_[12147]_  = ~A299 & A298;
  assign \new_[12150]_  = ~A302 & A300;
  assign \new_[12151]_  = \new_[12150]_  & \new_[12147]_ ;
  assign \new_[12152]_  = \new_[12151]_  & \new_[12144]_ ;
  assign \new_[12156]_  = A201 & ~A200;
  assign \new_[12157]_  = A199 & \new_[12156]_ ;
  assign \new_[12160]_  = ~A232 & ~A203;
  assign \new_[12163]_  = A234 & A233;
  assign \new_[12164]_  = \new_[12163]_  & \new_[12160]_ ;
  assign \new_[12165]_  = \new_[12164]_  & \new_[12157]_ ;
  assign \new_[12169]_  = A266 & A265;
  assign \new_[12170]_  = A235 & \new_[12169]_ ;
  assign \new_[12173]_  = A299 & ~A298;
  assign \new_[12176]_  = A301 & A300;
  assign \new_[12177]_  = \new_[12176]_  & \new_[12173]_ ;
  assign \new_[12178]_  = \new_[12177]_  & \new_[12170]_ ;
  assign \new_[12182]_  = A201 & ~A200;
  assign \new_[12183]_  = A199 & \new_[12182]_ ;
  assign \new_[12186]_  = ~A232 & ~A203;
  assign \new_[12189]_  = A234 & A233;
  assign \new_[12190]_  = \new_[12189]_  & \new_[12186]_ ;
  assign \new_[12191]_  = \new_[12190]_  & \new_[12183]_ ;
  assign \new_[12195]_  = A266 & A265;
  assign \new_[12196]_  = A235 & \new_[12195]_ ;
  assign \new_[12199]_  = A299 & ~A298;
  assign \new_[12202]_  = ~A302 & A300;
  assign \new_[12203]_  = \new_[12202]_  & \new_[12199]_ ;
  assign \new_[12204]_  = \new_[12203]_  & \new_[12196]_ ;
  assign \new_[12208]_  = A201 & ~A200;
  assign \new_[12209]_  = A199 & \new_[12208]_ ;
  assign \new_[12212]_  = ~A232 & ~A203;
  assign \new_[12215]_  = A234 & A233;
  assign \new_[12216]_  = \new_[12215]_  & \new_[12212]_ ;
  assign \new_[12217]_  = \new_[12216]_  & \new_[12209]_ ;
  assign \new_[12221]_  = ~A266 & ~A265;
  assign \new_[12222]_  = A235 & \new_[12221]_ ;
  assign \new_[12225]_  = ~A299 & A298;
  assign \new_[12228]_  = A301 & A300;
  assign \new_[12229]_  = \new_[12228]_  & \new_[12225]_ ;
  assign \new_[12230]_  = \new_[12229]_  & \new_[12222]_ ;
  assign \new_[12234]_  = A201 & ~A200;
  assign \new_[12235]_  = A199 & \new_[12234]_ ;
  assign \new_[12238]_  = ~A232 & ~A203;
  assign \new_[12241]_  = A234 & A233;
  assign \new_[12242]_  = \new_[12241]_  & \new_[12238]_ ;
  assign \new_[12243]_  = \new_[12242]_  & \new_[12235]_ ;
  assign \new_[12247]_  = ~A266 & ~A265;
  assign \new_[12248]_  = A235 & \new_[12247]_ ;
  assign \new_[12251]_  = ~A299 & A298;
  assign \new_[12254]_  = ~A302 & A300;
  assign \new_[12255]_  = \new_[12254]_  & \new_[12251]_ ;
  assign \new_[12256]_  = \new_[12255]_  & \new_[12248]_ ;
  assign \new_[12260]_  = A201 & ~A200;
  assign \new_[12261]_  = A199 & \new_[12260]_ ;
  assign \new_[12264]_  = ~A232 & ~A203;
  assign \new_[12267]_  = A234 & A233;
  assign \new_[12268]_  = \new_[12267]_  & \new_[12264]_ ;
  assign \new_[12269]_  = \new_[12268]_  & \new_[12261]_ ;
  assign \new_[12273]_  = ~A266 & ~A265;
  assign \new_[12274]_  = A235 & \new_[12273]_ ;
  assign \new_[12277]_  = A299 & ~A298;
  assign \new_[12280]_  = A301 & A300;
  assign \new_[12281]_  = \new_[12280]_  & \new_[12277]_ ;
  assign \new_[12282]_  = \new_[12281]_  & \new_[12274]_ ;
  assign \new_[12286]_  = A201 & ~A200;
  assign \new_[12287]_  = A199 & \new_[12286]_ ;
  assign \new_[12290]_  = ~A232 & ~A203;
  assign \new_[12293]_  = A234 & A233;
  assign \new_[12294]_  = \new_[12293]_  & \new_[12290]_ ;
  assign \new_[12295]_  = \new_[12294]_  & \new_[12287]_ ;
  assign \new_[12299]_  = ~A266 & ~A265;
  assign \new_[12300]_  = A235 & \new_[12299]_ ;
  assign \new_[12303]_  = A299 & ~A298;
  assign \new_[12306]_  = ~A302 & A300;
  assign \new_[12307]_  = \new_[12306]_  & \new_[12303]_ ;
  assign \new_[12308]_  = \new_[12307]_  & \new_[12300]_ ;
  assign \new_[12312]_  = A201 & ~A200;
  assign \new_[12313]_  = A199 & \new_[12312]_ ;
  assign \new_[12316]_  = ~A232 & ~A203;
  assign \new_[12319]_  = A234 & A233;
  assign \new_[12320]_  = \new_[12319]_  & \new_[12316]_ ;
  assign \new_[12321]_  = \new_[12320]_  & \new_[12313]_ ;
  assign \new_[12325]_  = A268 & ~A267;
  assign \new_[12326]_  = ~A236 & \new_[12325]_ ;
  assign \new_[12329]_  = ~A299 & A298;
  assign \new_[12332]_  = A301 & A300;
  assign \new_[12333]_  = \new_[12332]_  & \new_[12329]_ ;
  assign \new_[12334]_  = \new_[12333]_  & \new_[12326]_ ;
  assign \new_[12338]_  = A201 & ~A200;
  assign \new_[12339]_  = A199 & \new_[12338]_ ;
  assign \new_[12342]_  = ~A232 & ~A203;
  assign \new_[12345]_  = A234 & A233;
  assign \new_[12346]_  = \new_[12345]_  & \new_[12342]_ ;
  assign \new_[12347]_  = \new_[12346]_  & \new_[12339]_ ;
  assign \new_[12351]_  = A268 & ~A267;
  assign \new_[12352]_  = ~A236 & \new_[12351]_ ;
  assign \new_[12355]_  = ~A299 & A298;
  assign \new_[12358]_  = ~A302 & A300;
  assign \new_[12359]_  = \new_[12358]_  & \new_[12355]_ ;
  assign \new_[12360]_  = \new_[12359]_  & \new_[12352]_ ;
  assign \new_[12364]_  = A201 & ~A200;
  assign \new_[12365]_  = A199 & \new_[12364]_ ;
  assign \new_[12368]_  = ~A232 & ~A203;
  assign \new_[12371]_  = A234 & A233;
  assign \new_[12372]_  = \new_[12371]_  & \new_[12368]_ ;
  assign \new_[12373]_  = \new_[12372]_  & \new_[12365]_ ;
  assign \new_[12377]_  = A268 & ~A267;
  assign \new_[12378]_  = ~A236 & \new_[12377]_ ;
  assign \new_[12381]_  = A299 & ~A298;
  assign \new_[12384]_  = A301 & A300;
  assign \new_[12385]_  = \new_[12384]_  & \new_[12381]_ ;
  assign \new_[12386]_  = \new_[12385]_  & \new_[12378]_ ;
  assign \new_[12390]_  = A201 & ~A200;
  assign \new_[12391]_  = A199 & \new_[12390]_ ;
  assign \new_[12394]_  = ~A232 & ~A203;
  assign \new_[12397]_  = A234 & A233;
  assign \new_[12398]_  = \new_[12397]_  & \new_[12394]_ ;
  assign \new_[12399]_  = \new_[12398]_  & \new_[12391]_ ;
  assign \new_[12403]_  = A268 & ~A267;
  assign \new_[12404]_  = ~A236 & \new_[12403]_ ;
  assign \new_[12407]_  = A299 & ~A298;
  assign \new_[12410]_  = ~A302 & A300;
  assign \new_[12411]_  = \new_[12410]_  & \new_[12407]_ ;
  assign \new_[12412]_  = \new_[12411]_  & \new_[12404]_ ;
  assign \new_[12416]_  = A201 & ~A200;
  assign \new_[12417]_  = A199 & \new_[12416]_ ;
  assign \new_[12420]_  = ~A232 & ~A203;
  assign \new_[12423]_  = A234 & A233;
  assign \new_[12424]_  = \new_[12423]_  & \new_[12420]_ ;
  assign \new_[12425]_  = \new_[12424]_  & \new_[12417]_ ;
  assign \new_[12429]_  = ~A269 & ~A267;
  assign \new_[12430]_  = ~A236 & \new_[12429]_ ;
  assign \new_[12433]_  = ~A299 & A298;
  assign \new_[12436]_  = A301 & A300;
  assign \new_[12437]_  = \new_[12436]_  & \new_[12433]_ ;
  assign \new_[12438]_  = \new_[12437]_  & \new_[12430]_ ;
  assign \new_[12442]_  = A201 & ~A200;
  assign \new_[12443]_  = A199 & \new_[12442]_ ;
  assign \new_[12446]_  = ~A232 & ~A203;
  assign \new_[12449]_  = A234 & A233;
  assign \new_[12450]_  = \new_[12449]_  & \new_[12446]_ ;
  assign \new_[12451]_  = \new_[12450]_  & \new_[12443]_ ;
  assign \new_[12455]_  = ~A269 & ~A267;
  assign \new_[12456]_  = ~A236 & \new_[12455]_ ;
  assign \new_[12459]_  = ~A299 & A298;
  assign \new_[12462]_  = ~A302 & A300;
  assign \new_[12463]_  = \new_[12462]_  & \new_[12459]_ ;
  assign \new_[12464]_  = \new_[12463]_  & \new_[12456]_ ;
  assign \new_[12468]_  = A201 & ~A200;
  assign \new_[12469]_  = A199 & \new_[12468]_ ;
  assign \new_[12472]_  = ~A232 & ~A203;
  assign \new_[12475]_  = A234 & A233;
  assign \new_[12476]_  = \new_[12475]_  & \new_[12472]_ ;
  assign \new_[12477]_  = \new_[12476]_  & \new_[12469]_ ;
  assign \new_[12481]_  = ~A269 & ~A267;
  assign \new_[12482]_  = ~A236 & \new_[12481]_ ;
  assign \new_[12485]_  = A299 & ~A298;
  assign \new_[12488]_  = A301 & A300;
  assign \new_[12489]_  = \new_[12488]_  & \new_[12485]_ ;
  assign \new_[12490]_  = \new_[12489]_  & \new_[12482]_ ;
  assign \new_[12494]_  = A201 & ~A200;
  assign \new_[12495]_  = A199 & \new_[12494]_ ;
  assign \new_[12498]_  = ~A232 & ~A203;
  assign \new_[12501]_  = A234 & A233;
  assign \new_[12502]_  = \new_[12501]_  & \new_[12498]_ ;
  assign \new_[12503]_  = \new_[12502]_  & \new_[12495]_ ;
  assign \new_[12507]_  = ~A269 & ~A267;
  assign \new_[12508]_  = ~A236 & \new_[12507]_ ;
  assign \new_[12511]_  = A299 & ~A298;
  assign \new_[12514]_  = ~A302 & A300;
  assign \new_[12515]_  = \new_[12514]_  & \new_[12511]_ ;
  assign \new_[12516]_  = \new_[12515]_  & \new_[12508]_ ;
  assign \new_[12520]_  = A201 & ~A200;
  assign \new_[12521]_  = A199 & \new_[12520]_ ;
  assign \new_[12524]_  = ~A232 & ~A203;
  assign \new_[12527]_  = A234 & A233;
  assign \new_[12528]_  = \new_[12527]_  & \new_[12524]_ ;
  assign \new_[12529]_  = \new_[12528]_  & \new_[12521]_ ;
  assign \new_[12533]_  = A266 & A265;
  assign \new_[12534]_  = ~A236 & \new_[12533]_ ;
  assign \new_[12537]_  = ~A299 & A298;
  assign \new_[12540]_  = A301 & A300;
  assign \new_[12541]_  = \new_[12540]_  & \new_[12537]_ ;
  assign \new_[12542]_  = \new_[12541]_  & \new_[12534]_ ;
  assign \new_[12546]_  = A201 & ~A200;
  assign \new_[12547]_  = A199 & \new_[12546]_ ;
  assign \new_[12550]_  = ~A232 & ~A203;
  assign \new_[12553]_  = A234 & A233;
  assign \new_[12554]_  = \new_[12553]_  & \new_[12550]_ ;
  assign \new_[12555]_  = \new_[12554]_  & \new_[12547]_ ;
  assign \new_[12559]_  = A266 & A265;
  assign \new_[12560]_  = ~A236 & \new_[12559]_ ;
  assign \new_[12563]_  = ~A299 & A298;
  assign \new_[12566]_  = ~A302 & A300;
  assign \new_[12567]_  = \new_[12566]_  & \new_[12563]_ ;
  assign \new_[12568]_  = \new_[12567]_  & \new_[12560]_ ;
  assign \new_[12572]_  = A201 & ~A200;
  assign \new_[12573]_  = A199 & \new_[12572]_ ;
  assign \new_[12576]_  = ~A232 & ~A203;
  assign \new_[12579]_  = A234 & A233;
  assign \new_[12580]_  = \new_[12579]_  & \new_[12576]_ ;
  assign \new_[12581]_  = \new_[12580]_  & \new_[12573]_ ;
  assign \new_[12585]_  = A266 & A265;
  assign \new_[12586]_  = ~A236 & \new_[12585]_ ;
  assign \new_[12589]_  = A299 & ~A298;
  assign \new_[12592]_  = A301 & A300;
  assign \new_[12593]_  = \new_[12592]_  & \new_[12589]_ ;
  assign \new_[12594]_  = \new_[12593]_  & \new_[12586]_ ;
  assign \new_[12598]_  = A201 & ~A200;
  assign \new_[12599]_  = A199 & \new_[12598]_ ;
  assign \new_[12602]_  = ~A232 & ~A203;
  assign \new_[12605]_  = A234 & A233;
  assign \new_[12606]_  = \new_[12605]_  & \new_[12602]_ ;
  assign \new_[12607]_  = \new_[12606]_  & \new_[12599]_ ;
  assign \new_[12611]_  = A266 & A265;
  assign \new_[12612]_  = ~A236 & \new_[12611]_ ;
  assign \new_[12615]_  = A299 & ~A298;
  assign \new_[12618]_  = ~A302 & A300;
  assign \new_[12619]_  = \new_[12618]_  & \new_[12615]_ ;
  assign \new_[12620]_  = \new_[12619]_  & \new_[12612]_ ;
  assign \new_[12624]_  = A201 & ~A200;
  assign \new_[12625]_  = A199 & \new_[12624]_ ;
  assign \new_[12628]_  = ~A232 & ~A203;
  assign \new_[12631]_  = A234 & A233;
  assign \new_[12632]_  = \new_[12631]_  & \new_[12628]_ ;
  assign \new_[12633]_  = \new_[12632]_  & \new_[12625]_ ;
  assign \new_[12637]_  = ~A266 & ~A265;
  assign \new_[12638]_  = ~A236 & \new_[12637]_ ;
  assign \new_[12641]_  = ~A299 & A298;
  assign \new_[12644]_  = A301 & A300;
  assign \new_[12645]_  = \new_[12644]_  & \new_[12641]_ ;
  assign \new_[12646]_  = \new_[12645]_  & \new_[12638]_ ;
  assign \new_[12650]_  = A201 & ~A200;
  assign \new_[12651]_  = A199 & \new_[12650]_ ;
  assign \new_[12654]_  = ~A232 & ~A203;
  assign \new_[12657]_  = A234 & A233;
  assign \new_[12658]_  = \new_[12657]_  & \new_[12654]_ ;
  assign \new_[12659]_  = \new_[12658]_  & \new_[12651]_ ;
  assign \new_[12663]_  = ~A266 & ~A265;
  assign \new_[12664]_  = ~A236 & \new_[12663]_ ;
  assign \new_[12667]_  = ~A299 & A298;
  assign \new_[12670]_  = ~A302 & A300;
  assign \new_[12671]_  = \new_[12670]_  & \new_[12667]_ ;
  assign \new_[12672]_  = \new_[12671]_  & \new_[12664]_ ;
  assign \new_[12676]_  = A201 & ~A200;
  assign \new_[12677]_  = A199 & \new_[12676]_ ;
  assign \new_[12680]_  = ~A232 & ~A203;
  assign \new_[12683]_  = A234 & A233;
  assign \new_[12684]_  = \new_[12683]_  & \new_[12680]_ ;
  assign \new_[12685]_  = \new_[12684]_  & \new_[12677]_ ;
  assign \new_[12689]_  = ~A266 & ~A265;
  assign \new_[12690]_  = ~A236 & \new_[12689]_ ;
  assign \new_[12693]_  = A299 & ~A298;
  assign \new_[12696]_  = A301 & A300;
  assign \new_[12697]_  = \new_[12696]_  & \new_[12693]_ ;
  assign \new_[12698]_  = \new_[12697]_  & \new_[12690]_ ;
  assign \new_[12702]_  = A201 & ~A200;
  assign \new_[12703]_  = A199 & \new_[12702]_ ;
  assign \new_[12706]_  = ~A232 & ~A203;
  assign \new_[12709]_  = A234 & A233;
  assign \new_[12710]_  = \new_[12709]_  & \new_[12706]_ ;
  assign \new_[12711]_  = \new_[12710]_  & \new_[12703]_ ;
  assign \new_[12715]_  = ~A266 & ~A265;
  assign \new_[12716]_  = ~A236 & \new_[12715]_ ;
  assign \new_[12719]_  = A299 & ~A298;
  assign \new_[12722]_  = ~A302 & A300;
  assign \new_[12723]_  = \new_[12722]_  & \new_[12719]_ ;
  assign \new_[12724]_  = \new_[12723]_  & \new_[12716]_ ;
  assign \new_[12728]_  = A201 & ~A200;
  assign \new_[12729]_  = A199 & \new_[12728]_ ;
  assign \new_[12732]_  = A232 & ~A203;
  assign \new_[12735]_  = A234 & ~A233;
  assign \new_[12736]_  = \new_[12735]_  & \new_[12732]_ ;
  assign \new_[12737]_  = \new_[12736]_  & \new_[12729]_ ;
  assign \new_[12741]_  = A268 & ~A267;
  assign \new_[12742]_  = A235 & \new_[12741]_ ;
  assign \new_[12745]_  = ~A299 & A298;
  assign \new_[12748]_  = A301 & A300;
  assign \new_[12749]_  = \new_[12748]_  & \new_[12745]_ ;
  assign \new_[12750]_  = \new_[12749]_  & \new_[12742]_ ;
  assign \new_[12754]_  = A201 & ~A200;
  assign \new_[12755]_  = A199 & \new_[12754]_ ;
  assign \new_[12758]_  = A232 & ~A203;
  assign \new_[12761]_  = A234 & ~A233;
  assign \new_[12762]_  = \new_[12761]_  & \new_[12758]_ ;
  assign \new_[12763]_  = \new_[12762]_  & \new_[12755]_ ;
  assign \new_[12767]_  = A268 & ~A267;
  assign \new_[12768]_  = A235 & \new_[12767]_ ;
  assign \new_[12771]_  = ~A299 & A298;
  assign \new_[12774]_  = ~A302 & A300;
  assign \new_[12775]_  = \new_[12774]_  & \new_[12771]_ ;
  assign \new_[12776]_  = \new_[12775]_  & \new_[12768]_ ;
  assign \new_[12780]_  = A201 & ~A200;
  assign \new_[12781]_  = A199 & \new_[12780]_ ;
  assign \new_[12784]_  = A232 & ~A203;
  assign \new_[12787]_  = A234 & ~A233;
  assign \new_[12788]_  = \new_[12787]_  & \new_[12784]_ ;
  assign \new_[12789]_  = \new_[12788]_  & \new_[12781]_ ;
  assign \new_[12793]_  = A268 & ~A267;
  assign \new_[12794]_  = A235 & \new_[12793]_ ;
  assign \new_[12797]_  = A299 & ~A298;
  assign \new_[12800]_  = A301 & A300;
  assign \new_[12801]_  = \new_[12800]_  & \new_[12797]_ ;
  assign \new_[12802]_  = \new_[12801]_  & \new_[12794]_ ;
  assign \new_[12806]_  = A201 & ~A200;
  assign \new_[12807]_  = A199 & \new_[12806]_ ;
  assign \new_[12810]_  = A232 & ~A203;
  assign \new_[12813]_  = A234 & ~A233;
  assign \new_[12814]_  = \new_[12813]_  & \new_[12810]_ ;
  assign \new_[12815]_  = \new_[12814]_  & \new_[12807]_ ;
  assign \new_[12819]_  = A268 & ~A267;
  assign \new_[12820]_  = A235 & \new_[12819]_ ;
  assign \new_[12823]_  = A299 & ~A298;
  assign \new_[12826]_  = ~A302 & A300;
  assign \new_[12827]_  = \new_[12826]_  & \new_[12823]_ ;
  assign \new_[12828]_  = \new_[12827]_  & \new_[12820]_ ;
  assign \new_[12832]_  = A201 & ~A200;
  assign \new_[12833]_  = A199 & \new_[12832]_ ;
  assign \new_[12836]_  = A232 & ~A203;
  assign \new_[12839]_  = A234 & ~A233;
  assign \new_[12840]_  = \new_[12839]_  & \new_[12836]_ ;
  assign \new_[12841]_  = \new_[12840]_  & \new_[12833]_ ;
  assign \new_[12845]_  = ~A269 & ~A267;
  assign \new_[12846]_  = A235 & \new_[12845]_ ;
  assign \new_[12849]_  = ~A299 & A298;
  assign \new_[12852]_  = A301 & A300;
  assign \new_[12853]_  = \new_[12852]_  & \new_[12849]_ ;
  assign \new_[12854]_  = \new_[12853]_  & \new_[12846]_ ;
  assign \new_[12858]_  = A201 & ~A200;
  assign \new_[12859]_  = A199 & \new_[12858]_ ;
  assign \new_[12862]_  = A232 & ~A203;
  assign \new_[12865]_  = A234 & ~A233;
  assign \new_[12866]_  = \new_[12865]_  & \new_[12862]_ ;
  assign \new_[12867]_  = \new_[12866]_  & \new_[12859]_ ;
  assign \new_[12871]_  = ~A269 & ~A267;
  assign \new_[12872]_  = A235 & \new_[12871]_ ;
  assign \new_[12875]_  = ~A299 & A298;
  assign \new_[12878]_  = ~A302 & A300;
  assign \new_[12879]_  = \new_[12878]_  & \new_[12875]_ ;
  assign \new_[12880]_  = \new_[12879]_  & \new_[12872]_ ;
  assign \new_[12884]_  = A201 & ~A200;
  assign \new_[12885]_  = A199 & \new_[12884]_ ;
  assign \new_[12888]_  = A232 & ~A203;
  assign \new_[12891]_  = A234 & ~A233;
  assign \new_[12892]_  = \new_[12891]_  & \new_[12888]_ ;
  assign \new_[12893]_  = \new_[12892]_  & \new_[12885]_ ;
  assign \new_[12897]_  = ~A269 & ~A267;
  assign \new_[12898]_  = A235 & \new_[12897]_ ;
  assign \new_[12901]_  = A299 & ~A298;
  assign \new_[12904]_  = A301 & A300;
  assign \new_[12905]_  = \new_[12904]_  & \new_[12901]_ ;
  assign \new_[12906]_  = \new_[12905]_  & \new_[12898]_ ;
  assign \new_[12910]_  = A201 & ~A200;
  assign \new_[12911]_  = A199 & \new_[12910]_ ;
  assign \new_[12914]_  = A232 & ~A203;
  assign \new_[12917]_  = A234 & ~A233;
  assign \new_[12918]_  = \new_[12917]_  & \new_[12914]_ ;
  assign \new_[12919]_  = \new_[12918]_  & \new_[12911]_ ;
  assign \new_[12923]_  = ~A269 & ~A267;
  assign \new_[12924]_  = A235 & \new_[12923]_ ;
  assign \new_[12927]_  = A299 & ~A298;
  assign \new_[12930]_  = ~A302 & A300;
  assign \new_[12931]_  = \new_[12930]_  & \new_[12927]_ ;
  assign \new_[12932]_  = \new_[12931]_  & \new_[12924]_ ;
  assign \new_[12936]_  = A201 & ~A200;
  assign \new_[12937]_  = A199 & \new_[12936]_ ;
  assign \new_[12940]_  = A232 & ~A203;
  assign \new_[12943]_  = A234 & ~A233;
  assign \new_[12944]_  = \new_[12943]_  & \new_[12940]_ ;
  assign \new_[12945]_  = \new_[12944]_  & \new_[12937]_ ;
  assign \new_[12949]_  = A266 & A265;
  assign \new_[12950]_  = A235 & \new_[12949]_ ;
  assign \new_[12953]_  = ~A299 & A298;
  assign \new_[12956]_  = A301 & A300;
  assign \new_[12957]_  = \new_[12956]_  & \new_[12953]_ ;
  assign \new_[12958]_  = \new_[12957]_  & \new_[12950]_ ;
  assign \new_[12962]_  = A201 & ~A200;
  assign \new_[12963]_  = A199 & \new_[12962]_ ;
  assign \new_[12966]_  = A232 & ~A203;
  assign \new_[12969]_  = A234 & ~A233;
  assign \new_[12970]_  = \new_[12969]_  & \new_[12966]_ ;
  assign \new_[12971]_  = \new_[12970]_  & \new_[12963]_ ;
  assign \new_[12975]_  = A266 & A265;
  assign \new_[12976]_  = A235 & \new_[12975]_ ;
  assign \new_[12979]_  = ~A299 & A298;
  assign \new_[12982]_  = ~A302 & A300;
  assign \new_[12983]_  = \new_[12982]_  & \new_[12979]_ ;
  assign \new_[12984]_  = \new_[12983]_  & \new_[12976]_ ;
  assign \new_[12988]_  = A201 & ~A200;
  assign \new_[12989]_  = A199 & \new_[12988]_ ;
  assign \new_[12992]_  = A232 & ~A203;
  assign \new_[12995]_  = A234 & ~A233;
  assign \new_[12996]_  = \new_[12995]_  & \new_[12992]_ ;
  assign \new_[12997]_  = \new_[12996]_  & \new_[12989]_ ;
  assign \new_[13001]_  = A266 & A265;
  assign \new_[13002]_  = A235 & \new_[13001]_ ;
  assign \new_[13005]_  = A299 & ~A298;
  assign \new_[13008]_  = A301 & A300;
  assign \new_[13009]_  = \new_[13008]_  & \new_[13005]_ ;
  assign \new_[13010]_  = \new_[13009]_  & \new_[13002]_ ;
  assign \new_[13014]_  = A201 & ~A200;
  assign \new_[13015]_  = A199 & \new_[13014]_ ;
  assign \new_[13018]_  = A232 & ~A203;
  assign \new_[13021]_  = A234 & ~A233;
  assign \new_[13022]_  = \new_[13021]_  & \new_[13018]_ ;
  assign \new_[13023]_  = \new_[13022]_  & \new_[13015]_ ;
  assign \new_[13027]_  = A266 & A265;
  assign \new_[13028]_  = A235 & \new_[13027]_ ;
  assign \new_[13031]_  = A299 & ~A298;
  assign \new_[13034]_  = ~A302 & A300;
  assign \new_[13035]_  = \new_[13034]_  & \new_[13031]_ ;
  assign \new_[13036]_  = \new_[13035]_  & \new_[13028]_ ;
  assign \new_[13040]_  = A201 & ~A200;
  assign \new_[13041]_  = A199 & \new_[13040]_ ;
  assign \new_[13044]_  = A232 & ~A203;
  assign \new_[13047]_  = A234 & ~A233;
  assign \new_[13048]_  = \new_[13047]_  & \new_[13044]_ ;
  assign \new_[13049]_  = \new_[13048]_  & \new_[13041]_ ;
  assign \new_[13053]_  = ~A266 & ~A265;
  assign \new_[13054]_  = A235 & \new_[13053]_ ;
  assign \new_[13057]_  = ~A299 & A298;
  assign \new_[13060]_  = A301 & A300;
  assign \new_[13061]_  = \new_[13060]_  & \new_[13057]_ ;
  assign \new_[13062]_  = \new_[13061]_  & \new_[13054]_ ;
  assign \new_[13066]_  = A201 & ~A200;
  assign \new_[13067]_  = A199 & \new_[13066]_ ;
  assign \new_[13070]_  = A232 & ~A203;
  assign \new_[13073]_  = A234 & ~A233;
  assign \new_[13074]_  = \new_[13073]_  & \new_[13070]_ ;
  assign \new_[13075]_  = \new_[13074]_  & \new_[13067]_ ;
  assign \new_[13079]_  = ~A266 & ~A265;
  assign \new_[13080]_  = A235 & \new_[13079]_ ;
  assign \new_[13083]_  = ~A299 & A298;
  assign \new_[13086]_  = ~A302 & A300;
  assign \new_[13087]_  = \new_[13086]_  & \new_[13083]_ ;
  assign \new_[13088]_  = \new_[13087]_  & \new_[13080]_ ;
  assign \new_[13092]_  = A201 & ~A200;
  assign \new_[13093]_  = A199 & \new_[13092]_ ;
  assign \new_[13096]_  = A232 & ~A203;
  assign \new_[13099]_  = A234 & ~A233;
  assign \new_[13100]_  = \new_[13099]_  & \new_[13096]_ ;
  assign \new_[13101]_  = \new_[13100]_  & \new_[13093]_ ;
  assign \new_[13105]_  = ~A266 & ~A265;
  assign \new_[13106]_  = A235 & \new_[13105]_ ;
  assign \new_[13109]_  = A299 & ~A298;
  assign \new_[13112]_  = A301 & A300;
  assign \new_[13113]_  = \new_[13112]_  & \new_[13109]_ ;
  assign \new_[13114]_  = \new_[13113]_  & \new_[13106]_ ;
  assign \new_[13118]_  = A201 & ~A200;
  assign \new_[13119]_  = A199 & \new_[13118]_ ;
  assign \new_[13122]_  = A232 & ~A203;
  assign \new_[13125]_  = A234 & ~A233;
  assign \new_[13126]_  = \new_[13125]_  & \new_[13122]_ ;
  assign \new_[13127]_  = \new_[13126]_  & \new_[13119]_ ;
  assign \new_[13131]_  = ~A266 & ~A265;
  assign \new_[13132]_  = A235 & \new_[13131]_ ;
  assign \new_[13135]_  = A299 & ~A298;
  assign \new_[13138]_  = ~A302 & A300;
  assign \new_[13139]_  = \new_[13138]_  & \new_[13135]_ ;
  assign \new_[13140]_  = \new_[13139]_  & \new_[13132]_ ;
  assign \new_[13144]_  = A201 & ~A200;
  assign \new_[13145]_  = A199 & \new_[13144]_ ;
  assign \new_[13148]_  = A232 & ~A203;
  assign \new_[13151]_  = A234 & ~A233;
  assign \new_[13152]_  = \new_[13151]_  & \new_[13148]_ ;
  assign \new_[13153]_  = \new_[13152]_  & \new_[13145]_ ;
  assign \new_[13157]_  = A268 & ~A267;
  assign \new_[13158]_  = ~A236 & \new_[13157]_ ;
  assign \new_[13161]_  = ~A299 & A298;
  assign \new_[13164]_  = A301 & A300;
  assign \new_[13165]_  = \new_[13164]_  & \new_[13161]_ ;
  assign \new_[13166]_  = \new_[13165]_  & \new_[13158]_ ;
  assign \new_[13170]_  = A201 & ~A200;
  assign \new_[13171]_  = A199 & \new_[13170]_ ;
  assign \new_[13174]_  = A232 & ~A203;
  assign \new_[13177]_  = A234 & ~A233;
  assign \new_[13178]_  = \new_[13177]_  & \new_[13174]_ ;
  assign \new_[13179]_  = \new_[13178]_  & \new_[13171]_ ;
  assign \new_[13183]_  = A268 & ~A267;
  assign \new_[13184]_  = ~A236 & \new_[13183]_ ;
  assign \new_[13187]_  = ~A299 & A298;
  assign \new_[13190]_  = ~A302 & A300;
  assign \new_[13191]_  = \new_[13190]_  & \new_[13187]_ ;
  assign \new_[13192]_  = \new_[13191]_  & \new_[13184]_ ;
  assign \new_[13196]_  = A201 & ~A200;
  assign \new_[13197]_  = A199 & \new_[13196]_ ;
  assign \new_[13200]_  = A232 & ~A203;
  assign \new_[13203]_  = A234 & ~A233;
  assign \new_[13204]_  = \new_[13203]_  & \new_[13200]_ ;
  assign \new_[13205]_  = \new_[13204]_  & \new_[13197]_ ;
  assign \new_[13209]_  = A268 & ~A267;
  assign \new_[13210]_  = ~A236 & \new_[13209]_ ;
  assign \new_[13213]_  = A299 & ~A298;
  assign \new_[13216]_  = A301 & A300;
  assign \new_[13217]_  = \new_[13216]_  & \new_[13213]_ ;
  assign \new_[13218]_  = \new_[13217]_  & \new_[13210]_ ;
  assign \new_[13222]_  = A201 & ~A200;
  assign \new_[13223]_  = A199 & \new_[13222]_ ;
  assign \new_[13226]_  = A232 & ~A203;
  assign \new_[13229]_  = A234 & ~A233;
  assign \new_[13230]_  = \new_[13229]_  & \new_[13226]_ ;
  assign \new_[13231]_  = \new_[13230]_  & \new_[13223]_ ;
  assign \new_[13235]_  = A268 & ~A267;
  assign \new_[13236]_  = ~A236 & \new_[13235]_ ;
  assign \new_[13239]_  = A299 & ~A298;
  assign \new_[13242]_  = ~A302 & A300;
  assign \new_[13243]_  = \new_[13242]_  & \new_[13239]_ ;
  assign \new_[13244]_  = \new_[13243]_  & \new_[13236]_ ;
  assign \new_[13248]_  = A201 & ~A200;
  assign \new_[13249]_  = A199 & \new_[13248]_ ;
  assign \new_[13252]_  = A232 & ~A203;
  assign \new_[13255]_  = A234 & ~A233;
  assign \new_[13256]_  = \new_[13255]_  & \new_[13252]_ ;
  assign \new_[13257]_  = \new_[13256]_  & \new_[13249]_ ;
  assign \new_[13261]_  = ~A269 & ~A267;
  assign \new_[13262]_  = ~A236 & \new_[13261]_ ;
  assign \new_[13265]_  = ~A299 & A298;
  assign \new_[13268]_  = A301 & A300;
  assign \new_[13269]_  = \new_[13268]_  & \new_[13265]_ ;
  assign \new_[13270]_  = \new_[13269]_  & \new_[13262]_ ;
  assign \new_[13274]_  = A201 & ~A200;
  assign \new_[13275]_  = A199 & \new_[13274]_ ;
  assign \new_[13278]_  = A232 & ~A203;
  assign \new_[13281]_  = A234 & ~A233;
  assign \new_[13282]_  = \new_[13281]_  & \new_[13278]_ ;
  assign \new_[13283]_  = \new_[13282]_  & \new_[13275]_ ;
  assign \new_[13287]_  = ~A269 & ~A267;
  assign \new_[13288]_  = ~A236 & \new_[13287]_ ;
  assign \new_[13291]_  = ~A299 & A298;
  assign \new_[13294]_  = ~A302 & A300;
  assign \new_[13295]_  = \new_[13294]_  & \new_[13291]_ ;
  assign \new_[13296]_  = \new_[13295]_  & \new_[13288]_ ;
  assign \new_[13300]_  = A201 & ~A200;
  assign \new_[13301]_  = A199 & \new_[13300]_ ;
  assign \new_[13304]_  = A232 & ~A203;
  assign \new_[13307]_  = A234 & ~A233;
  assign \new_[13308]_  = \new_[13307]_  & \new_[13304]_ ;
  assign \new_[13309]_  = \new_[13308]_  & \new_[13301]_ ;
  assign \new_[13313]_  = ~A269 & ~A267;
  assign \new_[13314]_  = ~A236 & \new_[13313]_ ;
  assign \new_[13317]_  = A299 & ~A298;
  assign \new_[13320]_  = A301 & A300;
  assign \new_[13321]_  = \new_[13320]_  & \new_[13317]_ ;
  assign \new_[13322]_  = \new_[13321]_  & \new_[13314]_ ;
  assign \new_[13326]_  = A201 & ~A200;
  assign \new_[13327]_  = A199 & \new_[13326]_ ;
  assign \new_[13330]_  = A232 & ~A203;
  assign \new_[13333]_  = A234 & ~A233;
  assign \new_[13334]_  = \new_[13333]_  & \new_[13330]_ ;
  assign \new_[13335]_  = \new_[13334]_  & \new_[13327]_ ;
  assign \new_[13339]_  = ~A269 & ~A267;
  assign \new_[13340]_  = ~A236 & \new_[13339]_ ;
  assign \new_[13343]_  = A299 & ~A298;
  assign \new_[13346]_  = ~A302 & A300;
  assign \new_[13347]_  = \new_[13346]_  & \new_[13343]_ ;
  assign \new_[13348]_  = \new_[13347]_  & \new_[13340]_ ;
  assign \new_[13352]_  = A201 & ~A200;
  assign \new_[13353]_  = A199 & \new_[13352]_ ;
  assign \new_[13356]_  = A232 & ~A203;
  assign \new_[13359]_  = A234 & ~A233;
  assign \new_[13360]_  = \new_[13359]_  & \new_[13356]_ ;
  assign \new_[13361]_  = \new_[13360]_  & \new_[13353]_ ;
  assign \new_[13365]_  = A266 & A265;
  assign \new_[13366]_  = ~A236 & \new_[13365]_ ;
  assign \new_[13369]_  = ~A299 & A298;
  assign \new_[13372]_  = A301 & A300;
  assign \new_[13373]_  = \new_[13372]_  & \new_[13369]_ ;
  assign \new_[13374]_  = \new_[13373]_  & \new_[13366]_ ;
  assign \new_[13378]_  = A201 & ~A200;
  assign \new_[13379]_  = A199 & \new_[13378]_ ;
  assign \new_[13382]_  = A232 & ~A203;
  assign \new_[13385]_  = A234 & ~A233;
  assign \new_[13386]_  = \new_[13385]_  & \new_[13382]_ ;
  assign \new_[13387]_  = \new_[13386]_  & \new_[13379]_ ;
  assign \new_[13391]_  = A266 & A265;
  assign \new_[13392]_  = ~A236 & \new_[13391]_ ;
  assign \new_[13395]_  = ~A299 & A298;
  assign \new_[13398]_  = ~A302 & A300;
  assign \new_[13399]_  = \new_[13398]_  & \new_[13395]_ ;
  assign \new_[13400]_  = \new_[13399]_  & \new_[13392]_ ;
  assign \new_[13404]_  = A201 & ~A200;
  assign \new_[13405]_  = A199 & \new_[13404]_ ;
  assign \new_[13408]_  = A232 & ~A203;
  assign \new_[13411]_  = A234 & ~A233;
  assign \new_[13412]_  = \new_[13411]_  & \new_[13408]_ ;
  assign \new_[13413]_  = \new_[13412]_  & \new_[13405]_ ;
  assign \new_[13417]_  = A266 & A265;
  assign \new_[13418]_  = ~A236 & \new_[13417]_ ;
  assign \new_[13421]_  = A299 & ~A298;
  assign \new_[13424]_  = A301 & A300;
  assign \new_[13425]_  = \new_[13424]_  & \new_[13421]_ ;
  assign \new_[13426]_  = \new_[13425]_  & \new_[13418]_ ;
  assign \new_[13430]_  = A201 & ~A200;
  assign \new_[13431]_  = A199 & \new_[13430]_ ;
  assign \new_[13434]_  = A232 & ~A203;
  assign \new_[13437]_  = A234 & ~A233;
  assign \new_[13438]_  = \new_[13437]_  & \new_[13434]_ ;
  assign \new_[13439]_  = \new_[13438]_  & \new_[13431]_ ;
  assign \new_[13443]_  = A266 & A265;
  assign \new_[13444]_  = ~A236 & \new_[13443]_ ;
  assign \new_[13447]_  = A299 & ~A298;
  assign \new_[13450]_  = ~A302 & A300;
  assign \new_[13451]_  = \new_[13450]_  & \new_[13447]_ ;
  assign \new_[13452]_  = \new_[13451]_  & \new_[13444]_ ;
  assign \new_[13456]_  = A201 & ~A200;
  assign \new_[13457]_  = A199 & \new_[13456]_ ;
  assign \new_[13460]_  = A232 & ~A203;
  assign \new_[13463]_  = A234 & ~A233;
  assign \new_[13464]_  = \new_[13463]_  & \new_[13460]_ ;
  assign \new_[13465]_  = \new_[13464]_  & \new_[13457]_ ;
  assign \new_[13469]_  = ~A266 & ~A265;
  assign \new_[13470]_  = ~A236 & \new_[13469]_ ;
  assign \new_[13473]_  = ~A299 & A298;
  assign \new_[13476]_  = A301 & A300;
  assign \new_[13477]_  = \new_[13476]_  & \new_[13473]_ ;
  assign \new_[13478]_  = \new_[13477]_  & \new_[13470]_ ;
  assign \new_[13482]_  = A201 & ~A200;
  assign \new_[13483]_  = A199 & \new_[13482]_ ;
  assign \new_[13486]_  = A232 & ~A203;
  assign \new_[13489]_  = A234 & ~A233;
  assign \new_[13490]_  = \new_[13489]_  & \new_[13486]_ ;
  assign \new_[13491]_  = \new_[13490]_  & \new_[13483]_ ;
  assign \new_[13495]_  = ~A266 & ~A265;
  assign \new_[13496]_  = ~A236 & \new_[13495]_ ;
  assign \new_[13499]_  = ~A299 & A298;
  assign \new_[13502]_  = ~A302 & A300;
  assign \new_[13503]_  = \new_[13502]_  & \new_[13499]_ ;
  assign \new_[13504]_  = \new_[13503]_  & \new_[13496]_ ;
  assign \new_[13508]_  = A201 & ~A200;
  assign \new_[13509]_  = A199 & \new_[13508]_ ;
  assign \new_[13512]_  = A232 & ~A203;
  assign \new_[13515]_  = A234 & ~A233;
  assign \new_[13516]_  = \new_[13515]_  & \new_[13512]_ ;
  assign \new_[13517]_  = \new_[13516]_  & \new_[13509]_ ;
  assign \new_[13521]_  = ~A266 & ~A265;
  assign \new_[13522]_  = ~A236 & \new_[13521]_ ;
  assign \new_[13525]_  = A299 & ~A298;
  assign \new_[13528]_  = A301 & A300;
  assign \new_[13529]_  = \new_[13528]_  & \new_[13525]_ ;
  assign \new_[13530]_  = \new_[13529]_  & \new_[13522]_ ;
  assign \new_[13534]_  = A201 & ~A200;
  assign \new_[13535]_  = A199 & \new_[13534]_ ;
  assign \new_[13538]_  = A232 & ~A203;
  assign \new_[13541]_  = A234 & ~A233;
  assign \new_[13542]_  = \new_[13541]_  & \new_[13538]_ ;
  assign \new_[13543]_  = \new_[13542]_  & \new_[13535]_ ;
  assign \new_[13547]_  = ~A266 & ~A265;
  assign \new_[13548]_  = ~A236 & \new_[13547]_ ;
  assign \new_[13551]_  = A299 & ~A298;
  assign \new_[13554]_  = ~A302 & A300;
  assign \new_[13555]_  = \new_[13554]_  & \new_[13551]_ ;
  assign \new_[13556]_  = \new_[13555]_  & \new_[13548]_ ;
  assign \new_[13560]_  = A167 & A168;
  assign \new_[13561]_  = A170 & \new_[13560]_ ;
  assign \new_[13564]_  = ~A232 & ~A166;
  assign \new_[13567]_  = A234 & A233;
  assign \new_[13568]_  = \new_[13567]_  & \new_[13564]_ ;
  assign \new_[13569]_  = \new_[13568]_  & \new_[13561]_ ;
  assign \new_[13573]_  = A268 & ~A267;
  assign \new_[13574]_  = A235 & \new_[13573]_ ;
  assign \new_[13577]_  = ~A299 & A298;
  assign \new_[13580]_  = A301 & A300;
  assign \new_[13581]_  = \new_[13580]_  & \new_[13577]_ ;
  assign \new_[13582]_  = \new_[13581]_  & \new_[13574]_ ;
  assign \new_[13586]_  = A167 & A168;
  assign \new_[13587]_  = A170 & \new_[13586]_ ;
  assign \new_[13590]_  = ~A232 & ~A166;
  assign \new_[13593]_  = A234 & A233;
  assign \new_[13594]_  = \new_[13593]_  & \new_[13590]_ ;
  assign \new_[13595]_  = \new_[13594]_  & \new_[13587]_ ;
  assign \new_[13599]_  = A268 & ~A267;
  assign \new_[13600]_  = A235 & \new_[13599]_ ;
  assign \new_[13603]_  = ~A299 & A298;
  assign \new_[13606]_  = ~A302 & A300;
  assign \new_[13607]_  = \new_[13606]_  & \new_[13603]_ ;
  assign \new_[13608]_  = \new_[13607]_  & \new_[13600]_ ;
  assign \new_[13612]_  = A167 & A168;
  assign \new_[13613]_  = A170 & \new_[13612]_ ;
  assign \new_[13616]_  = ~A232 & ~A166;
  assign \new_[13619]_  = A234 & A233;
  assign \new_[13620]_  = \new_[13619]_  & \new_[13616]_ ;
  assign \new_[13621]_  = \new_[13620]_  & \new_[13613]_ ;
  assign \new_[13625]_  = A268 & ~A267;
  assign \new_[13626]_  = A235 & \new_[13625]_ ;
  assign \new_[13629]_  = A299 & ~A298;
  assign \new_[13632]_  = A301 & A300;
  assign \new_[13633]_  = \new_[13632]_  & \new_[13629]_ ;
  assign \new_[13634]_  = \new_[13633]_  & \new_[13626]_ ;
  assign \new_[13638]_  = A167 & A168;
  assign \new_[13639]_  = A170 & \new_[13638]_ ;
  assign \new_[13642]_  = ~A232 & ~A166;
  assign \new_[13645]_  = A234 & A233;
  assign \new_[13646]_  = \new_[13645]_  & \new_[13642]_ ;
  assign \new_[13647]_  = \new_[13646]_  & \new_[13639]_ ;
  assign \new_[13651]_  = A268 & ~A267;
  assign \new_[13652]_  = A235 & \new_[13651]_ ;
  assign \new_[13655]_  = A299 & ~A298;
  assign \new_[13658]_  = ~A302 & A300;
  assign \new_[13659]_  = \new_[13658]_  & \new_[13655]_ ;
  assign \new_[13660]_  = \new_[13659]_  & \new_[13652]_ ;
  assign \new_[13664]_  = A167 & A168;
  assign \new_[13665]_  = A170 & \new_[13664]_ ;
  assign \new_[13668]_  = ~A232 & ~A166;
  assign \new_[13671]_  = A234 & A233;
  assign \new_[13672]_  = \new_[13671]_  & \new_[13668]_ ;
  assign \new_[13673]_  = \new_[13672]_  & \new_[13665]_ ;
  assign \new_[13677]_  = ~A269 & ~A267;
  assign \new_[13678]_  = A235 & \new_[13677]_ ;
  assign \new_[13681]_  = ~A299 & A298;
  assign \new_[13684]_  = A301 & A300;
  assign \new_[13685]_  = \new_[13684]_  & \new_[13681]_ ;
  assign \new_[13686]_  = \new_[13685]_  & \new_[13678]_ ;
  assign \new_[13690]_  = A167 & A168;
  assign \new_[13691]_  = A170 & \new_[13690]_ ;
  assign \new_[13694]_  = ~A232 & ~A166;
  assign \new_[13697]_  = A234 & A233;
  assign \new_[13698]_  = \new_[13697]_  & \new_[13694]_ ;
  assign \new_[13699]_  = \new_[13698]_  & \new_[13691]_ ;
  assign \new_[13703]_  = ~A269 & ~A267;
  assign \new_[13704]_  = A235 & \new_[13703]_ ;
  assign \new_[13707]_  = ~A299 & A298;
  assign \new_[13710]_  = ~A302 & A300;
  assign \new_[13711]_  = \new_[13710]_  & \new_[13707]_ ;
  assign \new_[13712]_  = \new_[13711]_  & \new_[13704]_ ;
  assign \new_[13716]_  = A167 & A168;
  assign \new_[13717]_  = A170 & \new_[13716]_ ;
  assign \new_[13720]_  = ~A232 & ~A166;
  assign \new_[13723]_  = A234 & A233;
  assign \new_[13724]_  = \new_[13723]_  & \new_[13720]_ ;
  assign \new_[13725]_  = \new_[13724]_  & \new_[13717]_ ;
  assign \new_[13729]_  = ~A269 & ~A267;
  assign \new_[13730]_  = A235 & \new_[13729]_ ;
  assign \new_[13733]_  = A299 & ~A298;
  assign \new_[13736]_  = A301 & A300;
  assign \new_[13737]_  = \new_[13736]_  & \new_[13733]_ ;
  assign \new_[13738]_  = \new_[13737]_  & \new_[13730]_ ;
  assign \new_[13742]_  = A167 & A168;
  assign \new_[13743]_  = A170 & \new_[13742]_ ;
  assign \new_[13746]_  = ~A232 & ~A166;
  assign \new_[13749]_  = A234 & A233;
  assign \new_[13750]_  = \new_[13749]_  & \new_[13746]_ ;
  assign \new_[13751]_  = \new_[13750]_  & \new_[13743]_ ;
  assign \new_[13755]_  = ~A269 & ~A267;
  assign \new_[13756]_  = A235 & \new_[13755]_ ;
  assign \new_[13759]_  = A299 & ~A298;
  assign \new_[13762]_  = ~A302 & A300;
  assign \new_[13763]_  = \new_[13762]_  & \new_[13759]_ ;
  assign \new_[13764]_  = \new_[13763]_  & \new_[13756]_ ;
  assign \new_[13768]_  = A167 & A168;
  assign \new_[13769]_  = A170 & \new_[13768]_ ;
  assign \new_[13772]_  = ~A232 & ~A166;
  assign \new_[13775]_  = A234 & A233;
  assign \new_[13776]_  = \new_[13775]_  & \new_[13772]_ ;
  assign \new_[13777]_  = \new_[13776]_  & \new_[13769]_ ;
  assign \new_[13781]_  = A266 & A265;
  assign \new_[13782]_  = A235 & \new_[13781]_ ;
  assign \new_[13785]_  = ~A299 & A298;
  assign \new_[13788]_  = A301 & A300;
  assign \new_[13789]_  = \new_[13788]_  & \new_[13785]_ ;
  assign \new_[13790]_  = \new_[13789]_  & \new_[13782]_ ;
  assign \new_[13794]_  = A167 & A168;
  assign \new_[13795]_  = A170 & \new_[13794]_ ;
  assign \new_[13798]_  = ~A232 & ~A166;
  assign \new_[13801]_  = A234 & A233;
  assign \new_[13802]_  = \new_[13801]_  & \new_[13798]_ ;
  assign \new_[13803]_  = \new_[13802]_  & \new_[13795]_ ;
  assign \new_[13807]_  = A266 & A265;
  assign \new_[13808]_  = A235 & \new_[13807]_ ;
  assign \new_[13811]_  = ~A299 & A298;
  assign \new_[13814]_  = ~A302 & A300;
  assign \new_[13815]_  = \new_[13814]_  & \new_[13811]_ ;
  assign \new_[13816]_  = \new_[13815]_  & \new_[13808]_ ;
  assign \new_[13820]_  = A167 & A168;
  assign \new_[13821]_  = A170 & \new_[13820]_ ;
  assign \new_[13824]_  = ~A232 & ~A166;
  assign \new_[13827]_  = A234 & A233;
  assign \new_[13828]_  = \new_[13827]_  & \new_[13824]_ ;
  assign \new_[13829]_  = \new_[13828]_  & \new_[13821]_ ;
  assign \new_[13833]_  = A266 & A265;
  assign \new_[13834]_  = A235 & \new_[13833]_ ;
  assign \new_[13837]_  = A299 & ~A298;
  assign \new_[13840]_  = A301 & A300;
  assign \new_[13841]_  = \new_[13840]_  & \new_[13837]_ ;
  assign \new_[13842]_  = \new_[13841]_  & \new_[13834]_ ;
  assign \new_[13846]_  = A167 & A168;
  assign \new_[13847]_  = A170 & \new_[13846]_ ;
  assign \new_[13850]_  = ~A232 & ~A166;
  assign \new_[13853]_  = A234 & A233;
  assign \new_[13854]_  = \new_[13853]_  & \new_[13850]_ ;
  assign \new_[13855]_  = \new_[13854]_  & \new_[13847]_ ;
  assign \new_[13859]_  = A266 & A265;
  assign \new_[13860]_  = A235 & \new_[13859]_ ;
  assign \new_[13863]_  = A299 & ~A298;
  assign \new_[13866]_  = ~A302 & A300;
  assign \new_[13867]_  = \new_[13866]_  & \new_[13863]_ ;
  assign \new_[13868]_  = \new_[13867]_  & \new_[13860]_ ;
  assign \new_[13872]_  = A167 & A168;
  assign \new_[13873]_  = A170 & \new_[13872]_ ;
  assign \new_[13876]_  = ~A232 & ~A166;
  assign \new_[13879]_  = A234 & A233;
  assign \new_[13880]_  = \new_[13879]_  & \new_[13876]_ ;
  assign \new_[13881]_  = \new_[13880]_  & \new_[13873]_ ;
  assign \new_[13885]_  = ~A266 & ~A265;
  assign \new_[13886]_  = A235 & \new_[13885]_ ;
  assign \new_[13889]_  = ~A299 & A298;
  assign \new_[13892]_  = A301 & A300;
  assign \new_[13893]_  = \new_[13892]_  & \new_[13889]_ ;
  assign \new_[13894]_  = \new_[13893]_  & \new_[13886]_ ;
  assign \new_[13898]_  = A167 & A168;
  assign \new_[13899]_  = A170 & \new_[13898]_ ;
  assign \new_[13902]_  = ~A232 & ~A166;
  assign \new_[13905]_  = A234 & A233;
  assign \new_[13906]_  = \new_[13905]_  & \new_[13902]_ ;
  assign \new_[13907]_  = \new_[13906]_  & \new_[13899]_ ;
  assign \new_[13911]_  = ~A266 & ~A265;
  assign \new_[13912]_  = A235 & \new_[13911]_ ;
  assign \new_[13915]_  = ~A299 & A298;
  assign \new_[13918]_  = ~A302 & A300;
  assign \new_[13919]_  = \new_[13918]_  & \new_[13915]_ ;
  assign \new_[13920]_  = \new_[13919]_  & \new_[13912]_ ;
  assign \new_[13924]_  = A167 & A168;
  assign \new_[13925]_  = A170 & \new_[13924]_ ;
  assign \new_[13928]_  = ~A232 & ~A166;
  assign \new_[13931]_  = A234 & A233;
  assign \new_[13932]_  = \new_[13931]_  & \new_[13928]_ ;
  assign \new_[13933]_  = \new_[13932]_  & \new_[13925]_ ;
  assign \new_[13937]_  = ~A266 & ~A265;
  assign \new_[13938]_  = A235 & \new_[13937]_ ;
  assign \new_[13941]_  = A299 & ~A298;
  assign \new_[13944]_  = A301 & A300;
  assign \new_[13945]_  = \new_[13944]_  & \new_[13941]_ ;
  assign \new_[13946]_  = \new_[13945]_  & \new_[13938]_ ;
  assign \new_[13950]_  = A167 & A168;
  assign \new_[13951]_  = A170 & \new_[13950]_ ;
  assign \new_[13954]_  = ~A232 & ~A166;
  assign \new_[13957]_  = A234 & A233;
  assign \new_[13958]_  = \new_[13957]_  & \new_[13954]_ ;
  assign \new_[13959]_  = \new_[13958]_  & \new_[13951]_ ;
  assign \new_[13963]_  = ~A266 & ~A265;
  assign \new_[13964]_  = A235 & \new_[13963]_ ;
  assign \new_[13967]_  = A299 & ~A298;
  assign \new_[13970]_  = ~A302 & A300;
  assign \new_[13971]_  = \new_[13970]_  & \new_[13967]_ ;
  assign \new_[13972]_  = \new_[13971]_  & \new_[13964]_ ;
  assign \new_[13976]_  = A167 & A168;
  assign \new_[13977]_  = A170 & \new_[13976]_ ;
  assign \new_[13980]_  = ~A232 & ~A166;
  assign \new_[13983]_  = A234 & A233;
  assign \new_[13984]_  = \new_[13983]_  & \new_[13980]_ ;
  assign \new_[13985]_  = \new_[13984]_  & \new_[13977]_ ;
  assign \new_[13989]_  = A268 & ~A267;
  assign \new_[13990]_  = ~A236 & \new_[13989]_ ;
  assign \new_[13993]_  = ~A299 & A298;
  assign \new_[13996]_  = A301 & A300;
  assign \new_[13997]_  = \new_[13996]_  & \new_[13993]_ ;
  assign \new_[13998]_  = \new_[13997]_  & \new_[13990]_ ;
  assign \new_[14002]_  = A167 & A168;
  assign \new_[14003]_  = A170 & \new_[14002]_ ;
  assign \new_[14006]_  = ~A232 & ~A166;
  assign \new_[14009]_  = A234 & A233;
  assign \new_[14010]_  = \new_[14009]_  & \new_[14006]_ ;
  assign \new_[14011]_  = \new_[14010]_  & \new_[14003]_ ;
  assign \new_[14015]_  = A268 & ~A267;
  assign \new_[14016]_  = ~A236 & \new_[14015]_ ;
  assign \new_[14019]_  = ~A299 & A298;
  assign \new_[14022]_  = ~A302 & A300;
  assign \new_[14023]_  = \new_[14022]_  & \new_[14019]_ ;
  assign \new_[14024]_  = \new_[14023]_  & \new_[14016]_ ;
  assign \new_[14028]_  = A167 & A168;
  assign \new_[14029]_  = A170 & \new_[14028]_ ;
  assign \new_[14032]_  = ~A232 & ~A166;
  assign \new_[14035]_  = A234 & A233;
  assign \new_[14036]_  = \new_[14035]_  & \new_[14032]_ ;
  assign \new_[14037]_  = \new_[14036]_  & \new_[14029]_ ;
  assign \new_[14041]_  = A268 & ~A267;
  assign \new_[14042]_  = ~A236 & \new_[14041]_ ;
  assign \new_[14045]_  = A299 & ~A298;
  assign \new_[14048]_  = A301 & A300;
  assign \new_[14049]_  = \new_[14048]_  & \new_[14045]_ ;
  assign \new_[14050]_  = \new_[14049]_  & \new_[14042]_ ;
  assign \new_[14054]_  = A167 & A168;
  assign \new_[14055]_  = A170 & \new_[14054]_ ;
  assign \new_[14058]_  = ~A232 & ~A166;
  assign \new_[14061]_  = A234 & A233;
  assign \new_[14062]_  = \new_[14061]_  & \new_[14058]_ ;
  assign \new_[14063]_  = \new_[14062]_  & \new_[14055]_ ;
  assign \new_[14067]_  = A268 & ~A267;
  assign \new_[14068]_  = ~A236 & \new_[14067]_ ;
  assign \new_[14071]_  = A299 & ~A298;
  assign \new_[14074]_  = ~A302 & A300;
  assign \new_[14075]_  = \new_[14074]_  & \new_[14071]_ ;
  assign \new_[14076]_  = \new_[14075]_  & \new_[14068]_ ;
  assign \new_[14080]_  = A167 & A168;
  assign \new_[14081]_  = A170 & \new_[14080]_ ;
  assign \new_[14084]_  = ~A232 & ~A166;
  assign \new_[14087]_  = A234 & A233;
  assign \new_[14088]_  = \new_[14087]_  & \new_[14084]_ ;
  assign \new_[14089]_  = \new_[14088]_  & \new_[14081]_ ;
  assign \new_[14093]_  = ~A269 & ~A267;
  assign \new_[14094]_  = ~A236 & \new_[14093]_ ;
  assign \new_[14097]_  = ~A299 & A298;
  assign \new_[14100]_  = A301 & A300;
  assign \new_[14101]_  = \new_[14100]_  & \new_[14097]_ ;
  assign \new_[14102]_  = \new_[14101]_  & \new_[14094]_ ;
  assign \new_[14106]_  = A167 & A168;
  assign \new_[14107]_  = A170 & \new_[14106]_ ;
  assign \new_[14110]_  = ~A232 & ~A166;
  assign \new_[14113]_  = A234 & A233;
  assign \new_[14114]_  = \new_[14113]_  & \new_[14110]_ ;
  assign \new_[14115]_  = \new_[14114]_  & \new_[14107]_ ;
  assign \new_[14119]_  = ~A269 & ~A267;
  assign \new_[14120]_  = ~A236 & \new_[14119]_ ;
  assign \new_[14123]_  = ~A299 & A298;
  assign \new_[14126]_  = ~A302 & A300;
  assign \new_[14127]_  = \new_[14126]_  & \new_[14123]_ ;
  assign \new_[14128]_  = \new_[14127]_  & \new_[14120]_ ;
  assign \new_[14132]_  = A167 & A168;
  assign \new_[14133]_  = A170 & \new_[14132]_ ;
  assign \new_[14136]_  = ~A232 & ~A166;
  assign \new_[14139]_  = A234 & A233;
  assign \new_[14140]_  = \new_[14139]_  & \new_[14136]_ ;
  assign \new_[14141]_  = \new_[14140]_  & \new_[14133]_ ;
  assign \new_[14145]_  = ~A269 & ~A267;
  assign \new_[14146]_  = ~A236 & \new_[14145]_ ;
  assign \new_[14149]_  = A299 & ~A298;
  assign \new_[14152]_  = A301 & A300;
  assign \new_[14153]_  = \new_[14152]_  & \new_[14149]_ ;
  assign \new_[14154]_  = \new_[14153]_  & \new_[14146]_ ;
  assign \new_[14158]_  = A167 & A168;
  assign \new_[14159]_  = A170 & \new_[14158]_ ;
  assign \new_[14162]_  = ~A232 & ~A166;
  assign \new_[14165]_  = A234 & A233;
  assign \new_[14166]_  = \new_[14165]_  & \new_[14162]_ ;
  assign \new_[14167]_  = \new_[14166]_  & \new_[14159]_ ;
  assign \new_[14171]_  = ~A269 & ~A267;
  assign \new_[14172]_  = ~A236 & \new_[14171]_ ;
  assign \new_[14175]_  = A299 & ~A298;
  assign \new_[14178]_  = ~A302 & A300;
  assign \new_[14179]_  = \new_[14178]_  & \new_[14175]_ ;
  assign \new_[14180]_  = \new_[14179]_  & \new_[14172]_ ;
  assign \new_[14184]_  = A167 & A168;
  assign \new_[14185]_  = A170 & \new_[14184]_ ;
  assign \new_[14188]_  = ~A232 & ~A166;
  assign \new_[14191]_  = A234 & A233;
  assign \new_[14192]_  = \new_[14191]_  & \new_[14188]_ ;
  assign \new_[14193]_  = \new_[14192]_  & \new_[14185]_ ;
  assign \new_[14197]_  = A266 & A265;
  assign \new_[14198]_  = ~A236 & \new_[14197]_ ;
  assign \new_[14201]_  = ~A299 & A298;
  assign \new_[14204]_  = A301 & A300;
  assign \new_[14205]_  = \new_[14204]_  & \new_[14201]_ ;
  assign \new_[14206]_  = \new_[14205]_  & \new_[14198]_ ;
  assign \new_[14210]_  = A167 & A168;
  assign \new_[14211]_  = A170 & \new_[14210]_ ;
  assign \new_[14214]_  = ~A232 & ~A166;
  assign \new_[14217]_  = A234 & A233;
  assign \new_[14218]_  = \new_[14217]_  & \new_[14214]_ ;
  assign \new_[14219]_  = \new_[14218]_  & \new_[14211]_ ;
  assign \new_[14223]_  = A266 & A265;
  assign \new_[14224]_  = ~A236 & \new_[14223]_ ;
  assign \new_[14227]_  = ~A299 & A298;
  assign \new_[14230]_  = ~A302 & A300;
  assign \new_[14231]_  = \new_[14230]_  & \new_[14227]_ ;
  assign \new_[14232]_  = \new_[14231]_  & \new_[14224]_ ;
  assign \new_[14236]_  = A167 & A168;
  assign \new_[14237]_  = A170 & \new_[14236]_ ;
  assign \new_[14240]_  = ~A232 & ~A166;
  assign \new_[14243]_  = A234 & A233;
  assign \new_[14244]_  = \new_[14243]_  & \new_[14240]_ ;
  assign \new_[14245]_  = \new_[14244]_  & \new_[14237]_ ;
  assign \new_[14249]_  = A266 & A265;
  assign \new_[14250]_  = ~A236 & \new_[14249]_ ;
  assign \new_[14253]_  = A299 & ~A298;
  assign \new_[14256]_  = A301 & A300;
  assign \new_[14257]_  = \new_[14256]_  & \new_[14253]_ ;
  assign \new_[14258]_  = \new_[14257]_  & \new_[14250]_ ;
  assign \new_[14262]_  = A167 & A168;
  assign \new_[14263]_  = A170 & \new_[14262]_ ;
  assign \new_[14266]_  = ~A232 & ~A166;
  assign \new_[14269]_  = A234 & A233;
  assign \new_[14270]_  = \new_[14269]_  & \new_[14266]_ ;
  assign \new_[14271]_  = \new_[14270]_  & \new_[14263]_ ;
  assign \new_[14275]_  = A266 & A265;
  assign \new_[14276]_  = ~A236 & \new_[14275]_ ;
  assign \new_[14279]_  = A299 & ~A298;
  assign \new_[14282]_  = ~A302 & A300;
  assign \new_[14283]_  = \new_[14282]_  & \new_[14279]_ ;
  assign \new_[14284]_  = \new_[14283]_  & \new_[14276]_ ;
  assign \new_[14288]_  = A167 & A168;
  assign \new_[14289]_  = A170 & \new_[14288]_ ;
  assign \new_[14292]_  = ~A232 & ~A166;
  assign \new_[14295]_  = A234 & A233;
  assign \new_[14296]_  = \new_[14295]_  & \new_[14292]_ ;
  assign \new_[14297]_  = \new_[14296]_  & \new_[14289]_ ;
  assign \new_[14301]_  = ~A266 & ~A265;
  assign \new_[14302]_  = ~A236 & \new_[14301]_ ;
  assign \new_[14305]_  = ~A299 & A298;
  assign \new_[14308]_  = A301 & A300;
  assign \new_[14309]_  = \new_[14308]_  & \new_[14305]_ ;
  assign \new_[14310]_  = \new_[14309]_  & \new_[14302]_ ;
  assign \new_[14314]_  = A167 & A168;
  assign \new_[14315]_  = A170 & \new_[14314]_ ;
  assign \new_[14318]_  = ~A232 & ~A166;
  assign \new_[14321]_  = A234 & A233;
  assign \new_[14322]_  = \new_[14321]_  & \new_[14318]_ ;
  assign \new_[14323]_  = \new_[14322]_  & \new_[14315]_ ;
  assign \new_[14327]_  = ~A266 & ~A265;
  assign \new_[14328]_  = ~A236 & \new_[14327]_ ;
  assign \new_[14331]_  = ~A299 & A298;
  assign \new_[14334]_  = ~A302 & A300;
  assign \new_[14335]_  = \new_[14334]_  & \new_[14331]_ ;
  assign \new_[14336]_  = \new_[14335]_  & \new_[14328]_ ;
  assign \new_[14340]_  = A167 & A168;
  assign \new_[14341]_  = A170 & \new_[14340]_ ;
  assign \new_[14344]_  = ~A232 & ~A166;
  assign \new_[14347]_  = A234 & A233;
  assign \new_[14348]_  = \new_[14347]_  & \new_[14344]_ ;
  assign \new_[14349]_  = \new_[14348]_  & \new_[14341]_ ;
  assign \new_[14353]_  = ~A266 & ~A265;
  assign \new_[14354]_  = ~A236 & \new_[14353]_ ;
  assign \new_[14357]_  = A299 & ~A298;
  assign \new_[14360]_  = A301 & A300;
  assign \new_[14361]_  = \new_[14360]_  & \new_[14357]_ ;
  assign \new_[14362]_  = \new_[14361]_  & \new_[14354]_ ;
  assign \new_[14366]_  = A167 & A168;
  assign \new_[14367]_  = A170 & \new_[14366]_ ;
  assign \new_[14370]_  = ~A232 & ~A166;
  assign \new_[14373]_  = A234 & A233;
  assign \new_[14374]_  = \new_[14373]_  & \new_[14370]_ ;
  assign \new_[14375]_  = \new_[14374]_  & \new_[14367]_ ;
  assign \new_[14379]_  = ~A266 & ~A265;
  assign \new_[14380]_  = ~A236 & \new_[14379]_ ;
  assign \new_[14383]_  = A299 & ~A298;
  assign \new_[14386]_  = ~A302 & A300;
  assign \new_[14387]_  = \new_[14386]_  & \new_[14383]_ ;
  assign \new_[14388]_  = \new_[14387]_  & \new_[14380]_ ;
  assign \new_[14392]_  = A167 & A168;
  assign \new_[14393]_  = A170 & \new_[14392]_ ;
  assign \new_[14396]_  = A232 & ~A166;
  assign \new_[14399]_  = A234 & ~A233;
  assign \new_[14400]_  = \new_[14399]_  & \new_[14396]_ ;
  assign \new_[14401]_  = \new_[14400]_  & \new_[14393]_ ;
  assign \new_[14405]_  = A268 & ~A267;
  assign \new_[14406]_  = A235 & \new_[14405]_ ;
  assign \new_[14409]_  = ~A299 & A298;
  assign \new_[14412]_  = A301 & A300;
  assign \new_[14413]_  = \new_[14412]_  & \new_[14409]_ ;
  assign \new_[14414]_  = \new_[14413]_  & \new_[14406]_ ;
  assign \new_[14418]_  = A167 & A168;
  assign \new_[14419]_  = A170 & \new_[14418]_ ;
  assign \new_[14422]_  = A232 & ~A166;
  assign \new_[14425]_  = A234 & ~A233;
  assign \new_[14426]_  = \new_[14425]_  & \new_[14422]_ ;
  assign \new_[14427]_  = \new_[14426]_  & \new_[14419]_ ;
  assign \new_[14431]_  = A268 & ~A267;
  assign \new_[14432]_  = A235 & \new_[14431]_ ;
  assign \new_[14435]_  = ~A299 & A298;
  assign \new_[14438]_  = ~A302 & A300;
  assign \new_[14439]_  = \new_[14438]_  & \new_[14435]_ ;
  assign \new_[14440]_  = \new_[14439]_  & \new_[14432]_ ;
  assign \new_[14444]_  = A167 & A168;
  assign \new_[14445]_  = A170 & \new_[14444]_ ;
  assign \new_[14448]_  = A232 & ~A166;
  assign \new_[14451]_  = A234 & ~A233;
  assign \new_[14452]_  = \new_[14451]_  & \new_[14448]_ ;
  assign \new_[14453]_  = \new_[14452]_  & \new_[14445]_ ;
  assign \new_[14457]_  = A268 & ~A267;
  assign \new_[14458]_  = A235 & \new_[14457]_ ;
  assign \new_[14461]_  = A299 & ~A298;
  assign \new_[14464]_  = A301 & A300;
  assign \new_[14465]_  = \new_[14464]_  & \new_[14461]_ ;
  assign \new_[14466]_  = \new_[14465]_  & \new_[14458]_ ;
  assign \new_[14470]_  = A167 & A168;
  assign \new_[14471]_  = A170 & \new_[14470]_ ;
  assign \new_[14474]_  = A232 & ~A166;
  assign \new_[14477]_  = A234 & ~A233;
  assign \new_[14478]_  = \new_[14477]_  & \new_[14474]_ ;
  assign \new_[14479]_  = \new_[14478]_  & \new_[14471]_ ;
  assign \new_[14483]_  = A268 & ~A267;
  assign \new_[14484]_  = A235 & \new_[14483]_ ;
  assign \new_[14487]_  = A299 & ~A298;
  assign \new_[14490]_  = ~A302 & A300;
  assign \new_[14491]_  = \new_[14490]_  & \new_[14487]_ ;
  assign \new_[14492]_  = \new_[14491]_  & \new_[14484]_ ;
  assign \new_[14496]_  = A167 & A168;
  assign \new_[14497]_  = A170 & \new_[14496]_ ;
  assign \new_[14500]_  = A232 & ~A166;
  assign \new_[14503]_  = A234 & ~A233;
  assign \new_[14504]_  = \new_[14503]_  & \new_[14500]_ ;
  assign \new_[14505]_  = \new_[14504]_  & \new_[14497]_ ;
  assign \new_[14509]_  = ~A269 & ~A267;
  assign \new_[14510]_  = A235 & \new_[14509]_ ;
  assign \new_[14513]_  = ~A299 & A298;
  assign \new_[14516]_  = A301 & A300;
  assign \new_[14517]_  = \new_[14516]_  & \new_[14513]_ ;
  assign \new_[14518]_  = \new_[14517]_  & \new_[14510]_ ;
  assign \new_[14522]_  = A167 & A168;
  assign \new_[14523]_  = A170 & \new_[14522]_ ;
  assign \new_[14526]_  = A232 & ~A166;
  assign \new_[14529]_  = A234 & ~A233;
  assign \new_[14530]_  = \new_[14529]_  & \new_[14526]_ ;
  assign \new_[14531]_  = \new_[14530]_  & \new_[14523]_ ;
  assign \new_[14535]_  = ~A269 & ~A267;
  assign \new_[14536]_  = A235 & \new_[14535]_ ;
  assign \new_[14539]_  = ~A299 & A298;
  assign \new_[14542]_  = ~A302 & A300;
  assign \new_[14543]_  = \new_[14542]_  & \new_[14539]_ ;
  assign \new_[14544]_  = \new_[14543]_  & \new_[14536]_ ;
  assign \new_[14548]_  = A167 & A168;
  assign \new_[14549]_  = A170 & \new_[14548]_ ;
  assign \new_[14552]_  = A232 & ~A166;
  assign \new_[14555]_  = A234 & ~A233;
  assign \new_[14556]_  = \new_[14555]_  & \new_[14552]_ ;
  assign \new_[14557]_  = \new_[14556]_  & \new_[14549]_ ;
  assign \new_[14561]_  = ~A269 & ~A267;
  assign \new_[14562]_  = A235 & \new_[14561]_ ;
  assign \new_[14565]_  = A299 & ~A298;
  assign \new_[14568]_  = A301 & A300;
  assign \new_[14569]_  = \new_[14568]_  & \new_[14565]_ ;
  assign \new_[14570]_  = \new_[14569]_  & \new_[14562]_ ;
  assign \new_[14574]_  = A167 & A168;
  assign \new_[14575]_  = A170 & \new_[14574]_ ;
  assign \new_[14578]_  = A232 & ~A166;
  assign \new_[14581]_  = A234 & ~A233;
  assign \new_[14582]_  = \new_[14581]_  & \new_[14578]_ ;
  assign \new_[14583]_  = \new_[14582]_  & \new_[14575]_ ;
  assign \new_[14587]_  = ~A269 & ~A267;
  assign \new_[14588]_  = A235 & \new_[14587]_ ;
  assign \new_[14591]_  = A299 & ~A298;
  assign \new_[14594]_  = ~A302 & A300;
  assign \new_[14595]_  = \new_[14594]_  & \new_[14591]_ ;
  assign \new_[14596]_  = \new_[14595]_  & \new_[14588]_ ;
  assign \new_[14600]_  = A167 & A168;
  assign \new_[14601]_  = A170 & \new_[14600]_ ;
  assign \new_[14604]_  = A232 & ~A166;
  assign \new_[14607]_  = A234 & ~A233;
  assign \new_[14608]_  = \new_[14607]_  & \new_[14604]_ ;
  assign \new_[14609]_  = \new_[14608]_  & \new_[14601]_ ;
  assign \new_[14613]_  = A266 & A265;
  assign \new_[14614]_  = A235 & \new_[14613]_ ;
  assign \new_[14617]_  = ~A299 & A298;
  assign \new_[14620]_  = A301 & A300;
  assign \new_[14621]_  = \new_[14620]_  & \new_[14617]_ ;
  assign \new_[14622]_  = \new_[14621]_  & \new_[14614]_ ;
  assign \new_[14626]_  = A167 & A168;
  assign \new_[14627]_  = A170 & \new_[14626]_ ;
  assign \new_[14630]_  = A232 & ~A166;
  assign \new_[14633]_  = A234 & ~A233;
  assign \new_[14634]_  = \new_[14633]_  & \new_[14630]_ ;
  assign \new_[14635]_  = \new_[14634]_  & \new_[14627]_ ;
  assign \new_[14639]_  = A266 & A265;
  assign \new_[14640]_  = A235 & \new_[14639]_ ;
  assign \new_[14643]_  = ~A299 & A298;
  assign \new_[14646]_  = ~A302 & A300;
  assign \new_[14647]_  = \new_[14646]_  & \new_[14643]_ ;
  assign \new_[14648]_  = \new_[14647]_  & \new_[14640]_ ;
  assign \new_[14652]_  = A167 & A168;
  assign \new_[14653]_  = A170 & \new_[14652]_ ;
  assign \new_[14656]_  = A232 & ~A166;
  assign \new_[14659]_  = A234 & ~A233;
  assign \new_[14660]_  = \new_[14659]_  & \new_[14656]_ ;
  assign \new_[14661]_  = \new_[14660]_  & \new_[14653]_ ;
  assign \new_[14665]_  = A266 & A265;
  assign \new_[14666]_  = A235 & \new_[14665]_ ;
  assign \new_[14669]_  = A299 & ~A298;
  assign \new_[14672]_  = A301 & A300;
  assign \new_[14673]_  = \new_[14672]_  & \new_[14669]_ ;
  assign \new_[14674]_  = \new_[14673]_  & \new_[14666]_ ;
  assign \new_[14678]_  = A167 & A168;
  assign \new_[14679]_  = A170 & \new_[14678]_ ;
  assign \new_[14682]_  = A232 & ~A166;
  assign \new_[14685]_  = A234 & ~A233;
  assign \new_[14686]_  = \new_[14685]_  & \new_[14682]_ ;
  assign \new_[14687]_  = \new_[14686]_  & \new_[14679]_ ;
  assign \new_[14691]_  = A266 & A265;
  assign \new_[14692]_  = A235 & \new_[14691]_ ;
  assign \new_[14695]_  = A299 & ~A298;
  assign \new_[14698]_  = ~A302 & A300;
  assign \new_[14699]_  = \new_[14698]_  & \new_[14695]_ ;
  assign \new_[14700]_  = \new_[14699]_  & \new_[14692]_ ;
  assign \new_[14704]_  = A167 & A168;
  assign \new_[14705]_  = A170 & \new_[14704]_ ;
  assign \new_[14708]_  = A232 & ~A166;
  assign \new_[14711]_  = A234 & ~A233;
  assign \new_[14712]_  = \new_[14711]_  & \new_[14708]_ ;
  assign \new_[14713]_  = \new_[14712]_  & \new_[14705]_ ;
  assign \new_[14717]_  = ~A266 & ~A265;
  assign \new_[14718]_  = A235 & \new_[14717]_ ;
  assign \new_[14721]_  = ~A299 & A298;
  assign \new_[14724]_  = A301 & A300;
  assign \new_[14725]_  = \new_[14724]_  & \new_[14721]_ ;
  assign \new_[14726]_  = \new_[14725]_  & \new_[14718]_ ;
  assign \new_[14730]_  = A167 & A168;
  assign \new_[14731]_  = A170 & \new_[14730]_ ;
  assign \new_[14734]_  = A232 & ~A166;
  assign \new_[14737]_  = A234 & ~A233;
  assign \new_[14738]_  = \new_[14737]_  & \new_[14734]_ ;
  assign \new_[14739]_  = \new_[14738]_  & \new_[14731]_ ;
  assign \new_[14743]_  = ~A266 & ~A265;
  assign \new_[14744]_  = A235 & \new_[14743]_ ;
  assign \new_[14747]_  = ~A299 & A298;
  assign \new_[14750]_  = ~A302 & A300;
  assign \new_[14751]_  = \new_[14750]_  & \new_[14747]_ ;
  assign \new_[14752]_  = \new_[14751]_  & \new_[14744]_ ;
  assign \new_[14756]_  = A167 & A168;
  assign \new_[14757]_  = A170 & \new_[14756]_ ;
  assign \new_[14760]_  = A232 & ~A166;
  assign \new_[14763]_  = A234 & ~A233;
  assign \new_[14764]_  = \new_[14763]_  & \new_[14760]_ ;
  assign \new_[14765]_  = \new_[14764]_  & \new_[14757]_ ;
  assign \new_[14769]_  = ~A266 & ~A265;
  assign \new_[14770]_  = A235 & \new_[14769]_ ;
  assign \new_[14773]_  = A299 & ~A298;
  assign \new_[14776]_  = A301 & A300;
  assign \new_[14777]_  = \new_[14776]_  & \new_[14773]_ ;
  assign \new_[14778]_  = \new_[14777]_  & \new_[14770]_ ;
  assign \new_[14782]_  = A167 & A168;
  assign \new_[14783]_  = A170 & \new_[14782]_ ;
  assign \new_[14786]_  = A232 & ~A166;
  assign \new_[14789]_  = A234 & ~A233;
  assign \new_[14790]_  = \new_[14789]_  & \new_[14786]_ ;
  assign \new_[14791]_  = \new_[14790]_  & \new_[14783]_ ;
  assign \new_[14795]_  = ~A266 & ~A265;
  assign \new_[14796]_  = A235 & \new_[14795]_ ;
  assign \new_[14799]_  = A299 & ~A298;
  assign \new_[14802]_  = ~A302 & A300;
  assign \new_[14803]_  = \new_[14802]_  & \new_[14799]_ ;
  assign \new_[14804]_  = \new_[14803]_  & \new_[14796]_ ;
  assign \new_[14808]_  = A167 & A168;
  assign \new_[14809]_  = A170 & \new_[14808]_ ;
  assign \new_[14812]_  = A232 & ~A166;
  assign \new_[14815]_  = A234 & ~A233;
  assign \new_[14816]_  = \new_[14815]_  & \new_[14812]_ ;
  assign \new_[14817]_  = \new_[14816]_  & \new_[14809]_ ;
  assign \new_[14821]_  = A268 & ~A267;
  assign \new_[14822]_  = ~A236 & \new_[14821]_ ;
  assign \new_[14825]_  = ~A299 & A298;
  assign \new_[14828]_  = A301 & A300;
  assign \new_[14829]_  = \new_[14828]_  & \new_[14825]_ ;
  assign \new_[14830]_  = \new_[14829]_  & \new_[14822]_ ;
  assign \new_[14834]_  = A167 & A168;
  assign \new_[14835]_  = A170 & \new_[14834]_ ;
  assign \new_[14838]_  = A232 & ~A166;
  assign \new_[14841]_  = A234 & ~A233;
  assign \new_[14842]_  = \new_[14841]_  & \new_[14838]_ ;
  assign \new_[14843]_  = \new_[14842]_  & \new_[14835]_ ;
  assign \new_[14847]_  = A268 & ~A267;
  assign \new_[14848]_  = ~A236 & \new_[14847]_ ;
  assign \new_[14851]_  = ~A299 & A298;
  assign \new_[14854]_  = ~A302 & A300;
  assign \new_[14855]_  = \new_[14854]_  & \new_[14851]_ ;
  assign \new_[14856]_  = \new_[14855]_  & \new_[14848]_ ;
  assign \new_[14860]_  = A167 & A168;
  assign \new_[14861]_  = A170 & \new_[14860]_ ;
  assign \new_[14864]_  = A232 & ~A166;
  assign \new_[14867]_  = A234 & ~A233;
  assign \new_[14868]_  = \new_[14867]_  & \new_[14864]_ ;
  assign \new_[14869]_  = \new_[14868]_  & \new_[14861]_ ;
  assign \new_[14873]_  = A268 & ~A267;
  assign \new_[14874]_  = ~A236 & \new_[14873]_ ;
  assign \new_[14877]_  = A299 & ~A298;
  assign \new_[14880]_  = A301 & A300;
  assign \new_[14881]_  = \new_[14880]_  & \new_[14877]_ ;
  assign \new_[14882]_  = \new_[14881]_  & \new_[14874]_ ;
  assign \new_[14886]_  = A167 & A168;
  assign \new_[14887]_  = A170 & \new_[14886]_ ;
  assign \new_[14890]_  = A232 & ~A166;
  assign \new_[14893]_  = A234 & ~A233;
  assign \new_[14894]_  = \new_[14893]_  & \new_[14890]_ ;
  assign \new_[14895]_  = \new_[14894]_  & \new_[14887]_ ;
  assign \new_[14899]_  = A268 & ~A267;
  assign \new_[14900]_  = ~A236 & \new_[14899]_ ;
  assign \new_[14903]_  = A299 & ~A298;
  assign \new_[14906]_  = ~A302 & A300;
  assign \new_[14907]_  = \new_[14906]_  & \new_[14903]_ ;
  assign \new_[14908]_  = \new_[14907]_  & \new_[14900]_ ;
  assign \new_[14912]_  = A167 & A168;
  assign \new_[14913]_  = A170 & \new_[14912]_ ;
  assign \new_[14916]_  = A232 & ~A166;
  assign \new_[14919]_  = A234 & ~A233;
  assign \new_[14920]_  = \new_[14919]_  & \new_[14916]_ ;
  assign \new_[14921]_  = \new_[14920]_  & \new_[14913]_ ;
  assign \new_[14925]_  = ~A269 & ~A267;
  assign \new_[14926]_  = ~A236 & \new_[14925]_ ;
  assign \new_[14929]_  = ~A299 & A298;
  assign \new_[14932]_  = A301 & A300;
  assign \new_[14933]_  = \new_[14932]_  & \new_[14929]_ ;
  assign \new_[14934]_  = \new_[14933]_  & \new_[14926]_ ;
  assign \new_[14938]_  = A167 & A168;
  assign \new_[14939]_  = A170 & \new_[14938]_ ;
  assign \new_[14942]_  = A232 & ~A166;
  assign \new_[14945]_  = A234 & ~A233;
  assign \new_[14946]_  = \new_[14945]_  & \new_[14942]_ ;
  assign \new_[14947]_  = \new_[14946]_  & \new_[14939]_ ;
  assign \new_[14951]_  = ~A269 & ~A267;
  assign \new_[14952]_  = ~A236 & \new_[14951]_ ;
  assign \new_[14955]_  = ~A299 & A298;
  assign \new_[14958]_  = ~A302 & A300;
  assign \new_[14959]_  = \new_[14958]_  & \new_[14955]_ ;
  assign \new_[14960]_  = \new_[14959]_  & \new_[14952]_ ;
  assign \new_[14964]_  = A167 & A168;
  assign \new_[14965]_  = A170 & \new_[14964]_ ;
  assign \new_[14968]_  = A232 & ~A166;
  assign \new_[14971]_  = A234 & ~A233;
  assign \new_[14972]_  = \new_[14971]_  & \new_[14968]_ ;
  assign \new_[14973]_  = \new_[14972]_  & \new_[14965]_ ;
  assign \new_[14977]_  = ~A269 & ~A267;
  assign \new_[14978]_  = ~A236 & \new_[14977]_ ;
  assign \new_[14981]_  = A299 & ~A298;
  assign \new_[14984]_  = A301 & A300;
  assign \new_[14985]_  = \new_[14984]_  & \new_[14981]_ ;
  assign \new_[14986]_  = \new_[14985]_  & \new_[14978]_ ;
  assign \new_[14990]_  = A167 & A168;
  assign \new_[14991]_  = A170 & \new_[14990]_ ;
  assign \new_[14994]_  = A232 & ~A166;
  assign \new_[14997]_  = A234 & ~A233;
  assign \new_[14998]_  = \new_[14997]_  & \new_[14994]_ ;
  assign \new_[14999]_  = \new_[14998]_  & \new_[14991]_ ;
  assign \new_[15003]_  = ~A269 & ~A267;
  assign \new_[15004]_  = ~A236 & \new_[15003]_ ;
  assign \new_[15007]_  = A299 & ~A298;
  assign \new_[15010]_  = ~A302 & A300;
  assign \new_[15011]_  = \new_[15010]_  & \new_[15007]_ ;
  assign \new_[15012]_  = \new_[15011]_  & \new_[15004]_ ;
  assign \new_[15016]_  = A167 & A168;
  assign \new_[15017]_  = A170 & \new_[15016]_ ;
  assign \new_[15020]_  = A232 & ~A166;
  assign \new_[15023]_  = A234 & ~A233;
  assign \new_[15024]_  = \new_[15023]_  & \new_[15020]_ ;
  assign \new_[15025]_  = \new_[15024]_  & \new_[15017]_ ;
  assign \new_[15029]_  = A266 & A265;
  assign \new_[15030]_  = ~A236 & \new_[15029]_ ;
  assign \new_[15033]_  = ~A299 & A298;
  assign \new_[15036]_  = A301 & A300;
  assign \new_[15037]_  = \new_[15036]_  & \new_[15033]_ ;
  assign \new_[15038]_  = \new_[15037]_  & \new_[15030]_ ;
  assign \new_[15042]_  = A167 & A168;
  assign \new_[15043]_  = A170 & \new_[15042]_ ;
  assign \new_[15046]_  = A232 & ~A166;
  assign \new_[15049]_  = A234 & ~A233;
  assign \new_[15050]_  = \new_[15049]_  & \new_[15046]_ ;
  assign \new_[15051]_  = \new_[15050]_  & \new_[15043]_ ;
  assign \new_[15055]_  = A266 & A265;
  assign \new_[15056]_  = ~A236 & \new_[15055]_ ;
  assign \new_[15059]_  = ~A299 & A298;
  assign \new_[15062]_  = ~A302 & A300;
  assign \new_[15063]_  = \new_[15062]_  & \new_[15059]_ ;
  assign \new_[15064]_  = \new_[15063]_  & \new_[15056]_ ;
  assign \new_[15068]_  = A167 & A168;
  assign \new_[15069]_  = A170 & \new_[15068]_ ;
  assign \new_[15072]_  = A232 & ~A166;
  assign \new_[15075]_  = A234 & ~A233;
  assign \new_[15076]_  = \new_[15075]_  & \new_[15072]_ ;
  assign \new_[15077]_  = \new_[15076]_  & \new_[15069]_ ;
  assign \new_[15081]_  = A266 & A265;
  assign \new_[15082]_  = ~A236 & \new_[15081]_ ;
  assign \new_[15085]_  = A299 & ~A298;
  assign \new_[15088]_  = A301 & A300;
  assign \new_[15089]_  = \new_[15088]_  & \new_[15085]_ ;
  assign \new_[15090]_  = \new_[15089]_  & \new_[15082]_ ;
  assign \new_[15094]_  = A167 & A168;
  assign \new_[15095]_  = A170 & \new_[15094]_ ;
  assign \new_[15098]_  = A232 & ~A166;
  assign \new_[15101]_  = A234 & ~A233;
  assign \new_[15102]_  = \new_[15101]_  & \new_[15098]_ ;
  assign \new_[15103]_  = \new_[15102]_  & \new_[15095]_ ;
  assign \new_[15107]_  = A266 & A265;
  assign \new_[15108]_  = ~A236 & \new_[15107]_ ;
  assign \new_[15111]_  = A299 & ~A298;
  assign \new_[15114]_  = ~A302 & A300;
  assign \new_[15115]_  = \new_[15114]_  & \new_[15111]_ ;
  assign \new_[15116]_  = \new_[15115]_  & \new_[15108]_ ;
  assign \new_[15120]_  = A167 & A168;
  assign \new_[15121]_  = A170 & \new_[15120]_ ;
  assign \new_[15124]_  = A232 & ~A166;
  assign \new_[15127]_  = A234 & ~A233;
  assign \new_[15128]_  = \new_[15127]_  & \new_[15124]_ ;
  assign \new_[15129]_  = \new_[15128]_  & \new_[15121]_ ;
  assign \new_[15133]_  = ~A266 & ~A265;
  assign \new_[15134]_  = ~A236 & \new_[15133]_ ;
  assign \new_[15137]_  = ~A299 & A298;
  assign \new_[15140]_  = A301 & A300;
  assign \new_[15141]_  = \new_[15140]_  & \new_[15137]_ ;
  assign \new_[15142]_  = \new_[15141]_  & \new_[15134]_ ;
  assign \new_[15146]_  = A167 & A168;
  assign \new_[15147]_  = A170 & \new_[15146]_ ;
  assign \new_[15150]_  = A232 & ~A166;
  assign \new_[15153]_  = A234 & ~A233;
  assign \new_[15154]_  = \new_[15153]_  & \new_[15150]_ ;
  assign \new_[15155]_  = \new_[15154]_  & \new_[15147]_ ;
  assign \new_[15159]_  = ~A266 & ~A265;
  assign \new_[15160]_  = ~A236 & \new_[15159]_ ;
  assign \new_[15163]_  = ~A299 & A298;
  assign \new_[15166]_  = ~A302 & A300;
  assign \new_[15167]_  = \new_[15166]_  & \new_[15163]_ ;
  assign \new_[15168]_  = \new_[15167]_  & \new_[15160]_ ;
  assign \new_[15172]_  = A167 & A168;
  assign \new_[15173]_  = A170 & \new_[15172]_ ;
  assign \new_[15176]_  = A232 & ~A166;
  assign \new_[15179]_  = A234 & ~A233;
  assign \new_[15180]_  = \new_[15179]_  & \new_[15176]_ ;
  assign \new_[15181]_  = \new_[15180]_  & \new_[15173]_ ;
  assign \new_[15185]_  = ~A266 & ~A265;
  assign \new_[15186]_  = ~A236 & \new_[15185]_ ;
  assign \new_[15189]_  = A299 & ~A298;
  assign \new_[15192]_  = A301 & A300;
  assign \new_[15193]_  = \new_[15192]_  & \new_[15189]_ ;
  assign \new_[15194]_  = \new_[15193]_  & \new_[15186]_ ;
  assign \new_[15198]_  = A167 & A168;
  assign \new_[15199]_  = A170 & \new_[15198]_ ;
  assign \new_[15202]_  = A232 & ~A166;
  assign \new_[15205]_  = A234 & ~A233;
  assign \new_[15206]_  = \new_[15205]_  & \new_[15202]_ ;
  assign \new_[15207]_  = \new_[15206]_  & \new_[15199]_ ;
  assign \new_[15211]_  = ~A266 & ~A265;
  assign \new_[15212]_  = ~A236 & \new_[15211]_ ;
  assign \new_[15215]_  = A299 & ~A298;
  assign \new_[15218]_  = ~A302 & A300;
  assign \new_[15219]_  = \new_[15218]_  & \new_[15215]_ ;
  assign \new_[15220]_  = \new_[15219]_  & \new_[15212]_ ;
  assign \new_[15224]_  = ~A167 & A168;
  assign \new_[15225]_  = A170 & \new_[15224]_ ;
  assign \new_[15228]_  = ~A232 & A166;
  assign \new_[15231]_  = A234 & A233;
  assign \new_[15232]_  = \new_[15231]_  & \new_[15228]_ ;
  assign \new_[15233]_  = \new_[15232]_  & \new_[15225]_ ;
  assign \new_[15237]_  = A268 & ~A267;
  assign \new_[15238]_  = A235 & \new_[15237]_ ;
  assign \new_[15241]_  = ~A299 & A298;
  assign \new_[15244]_  = A301 & A300;
  assign \new_[15245]_  = \new_[15244]_  & \new_[15241]_ ;
  assign \new_[15246]_  = \new_[15245]_  & \new_[15238]_ ;
  assign \new_[15250]_  = ~A167 & A168;
  assign \new_[15251]_  = A170 & \new_[15250]_ ;
  assign \new_[15254]_  = ~A232 & A166;
  assign \new_[15257]_  = A234 & A233;
  assign \new_[15258]_  = \new_[15257]_  & \new_[15254]_ ;
  assign \new_[15259]_  = \new_[15258]_  & \new_[15251]_ ;
  assign \new_[15263]_  = A268 & ~A267;
  assign \new_[15264]_  = A235 & \new_[15263]_ ;
  assign \new_[15267]_  = ~A299 & A298;
  assign \new_[15270]_  = ~A302 & A300;
  assign \new_[15271]_  = \new_[15270]_  & \new_[15267]_ ;
  assign \new_[15272]_  = \new_[15271]_  & \new_[15264]_ ;
  assign \new_[15276]_  = ~A167 & A168;
  assign \new_[15277]_  = A170 & \new_[15276]_ ;
  assign \new_[15280]_  = ~A232 & A166;
  assign \new_[15283]_  = A234 & A233;
  assign \new_[15284]_  = \new_[15283]_  & \new_[15280]_ ;
  assign \new_[15285]_  = \new_[15284]_  & \new_[15277]_ ;
  assign \new_[15289]_  = A268 & ~A267;
  assign \new_[15290]_  = A235 & \new_[15289]_ ;
  assign \new_[15293]_  = A299 & ~A298;
  assign \new_[15296]_  = A301 & A300;
  assign \new_[15297]_  = \new_[15296]_  & \new_[15293]_ ;
  assign \new_[15298]_  = \new_[15297]_  & \new_[15290]_ ;
  assign \new_[15302]_  = ~A167 & A168;
  assign \new_[15303]_  = A170 & \new_[15302]_ ;
  assign \new_[15306]_  = ~A232 & A166;
  assign \new_[15309]_  = A234 & A233;
  assign \new_[15310]_  = \new_[15309]_  & \new_[15306]_ ;
  assign \new_[15311]_  = \new_[15310]_  & \new_[15303]_ ;
  assign \new_[15315]_  = A268 & ~A267;
  assign \new_[15316]_  = A235 & \new_[15315]_ ;
  assign \new_[15319]_  = A299 & ~A298;
  assign \new_[15322]_  = ~A302 & A300;
  assign \new_[15323]_  = \new_[15322]_  & \new_[15319]_ ;
  assign \new_[15324]_  = \new_[15323]_  & \new_[15316]_ ;
  assign \new_[15328]_  = ~A167 & A168;
  assign \new_[15329]_  = A170 & \new_[15328]_ ;
  assign \new_[15332]_  = ~A232 & A166;
  assign \new_[15335]_  = A234 & A233;
  assign \new_[15336]_  = \new_[15335]_  & \new_[15332]_ ;
  assign \new_[15337]_  = \new_[15336]_  & \new_[15329]_ ;
  assign \new_[15341]_  = ~A269 & ~A267;
  assign \new_[15342]_  = A235 & \new_[15341]_ ;
  assign \new_[15345]_  = ~A299 & A298;
  assign \new_[15348]_  = A301 & A300;
  assign \new_[15349]_  = \new_[15348]_  & \new_[15345]_ ;
  assign \new_[15350]_  = \new_[15349]_  & \new_[15342]_ ;
  assign \new_[15354]_  = ~A167 & A168;
  assign \new_[15355]_  = A170 & \new_[15354]_ ;
  assign \new_[15358]_  = ~A232 & A166;
  assign \new_[15361]_  = A234 & A233;
  assign \new_[15362]_  = \new_[15361]_  & \new_[15358]_ ;
  assign \new_[15363]_  = \new_[15362]_  & \new_[15355]_ ;
  assign \new_[15367]_  = ~A269 & ~A267;
  assign \new_[15368]_  = A235 & \new_[15367]_ ;
  assign \new_[15371]_  = ~A299 & A298;
  assign \new_[15374]_  = ~A302 & A300;
  assign \new_[15375]_  = \new_[15374]_  & \new_[15371]_ ;
  assign \new_[15376]_  = \new_[15375]_  & \new_[15368]_ ;
  assign \new_[15380]_  = ~A167 & A168;
  assign \new_[15381]_  = A170 & \new_[15380]_ ;
  assign \new_[15384]_  = ~A232 & A166;
  assign \new_[15387]_  = A234 & A233;
  assign \new_[15388]_  = \new_[15387]_  & \new_[15384]_ ;
  assign \new_[15389]_  = \new_[15388]_  & \new_[15381]_ ;
  assign \new_[15393]_  = ~A269 & ~A267;
  assign \new_[15394]_  = A235 & \new_[15393]_ ;
  assign \new_[15397]_  = A299 & ~A298;
  assign \new_[15400]_  = A301 & A300;
  assign \new_[15401]_  = \new_[15400]_  & \new_[15397]_ ;
  assign \new_[15402]_  = \new_[15401]_  & \new_[15394]_ ;
  assign \new_[15406]_  = ~A167 & A168;
  assign \new_[15407]_  = A170 & \new_[15406]_ ;
  assign \new_[15410]_  = ~A232 & A166;
  assign \new_[15413]_  = A234 & A233;
  assign \new_[15414]_  = \new_[15413]_  & \new_[15410]_ ;
  assign \new_[15415]_  = \new_[15414]_  & \new_[15407]_ ;
  assign \new_[15419]_  = ~A269 & ~A267;
  assign \new_[15420]_  = A235 & \new_[15419]_ ;
  assign \new_[15423]_  = A299 & ~A298;
  assign \new_[15426]_  = ~A302 & A300;
  assign \new_[15427]_  = \new_[15426]_  & \new_[15423]_ ;
  assign \new_[15428]_  = \new_[15427]_  & \new_[15420]_ ;
  assign \new_[15432]_  = ~A167 & A168;
  assign \new_[15433]_  = A170 & \new_[15432]_ ;
  assign \new_[15436]_  = ~A232 & A166;
  assign \new_[15439]_  = A234 & A233;
  assign \new_[15440]_  = \new_[15439]_  & \new_[15436]_ ;
  assign \new_[15441]_  = \new_[15440]_  & \new_[15433]_ ;
  assign \new_[15445]_  = A266 & A265;
  assign \new_[15446]_  = A235 & \new_[15445]_ ;
  assign \new_[15449]_  = ~A299 & A298;
  assign \new_[15452]_  = A301 & A300;
  assign \new_[15453]_  = \new_[15452]_  & \new_[15449]_ ;
  assign \new_[15454]_  = \new_[15453]_  & \new_[15446]_ ;
  assign \new_[15458]_  = ~A167 & A168;
  assign \new_[15459]_  = A170 & \new_[15458]_ ;
  assign \new_[15462]_  = ~A232 & A166;
  assign \new_[15465]_  = A234 & A233;
  assign \new_[15466]_  = \new_[15465]_  & \new_[15462]_ ;
  assign \new_[15467]_  = \new_[15466]_  & \new_[15459]_ ;
  assign \new_[15471]_  = A266 & A265;
  assign \new_[15472]_  = A235 & \new_[15471]_ ;
  assign \new_[15475]_  = ~A299 & A298;
  assign \new_[15478]_  = ~A302 & A300;
  assign \new_[15479]_  = \new_[15478]_  & \new_[15475]_ ;
  assign \new_[15480]_  = \new_[15479]_  & \new_[15472]_ ;
  assign \new_[15484]_  = ~A167 & A168;
  assign \new_[15485]_  = A170 & \new_[15484]_ ;
  assign \new_[15488]_  = ~A232 & A166;
  assign \new_[15491]_  = A234 & A233;
  assign \new_[15492]_  = \new_[15491]_  & \new_[15488]_ ;
  assign \new_[15493]_  = \new_[15492]_  & \new_[15485]_ ;
  assign \new_[15497]_  = A266 & A265;
  assign \new_[15498]_  = A235 & \new_[15497]_ ;
  assign \new_[15501]_  = A299 & ~A298;
  assign \new_[15504]_  = A301 & A300;
  assign \new_[15505]_  = \new_[15504]_  & \new_[15501]_ ;
  assign \new_[15506]_  = \new_[15505]_  & \new_[15498]_ ;
  assign \new_[15510]_  = ~A167 & A168;
  assign \new_[15511]_  = A170 & \new_[15510]_ ;
  assign \new_[15514]_  = ~A232 & A166;
  assign \new_[15517]_  = A234 & A233;
  assign \new_[15518]_  = \new_[15517]_  & \new_[15514]_ ;
  assign \new_[15519]_  = \new_[15518]_  & \new_[15511]_ ;
  assign \new_[15523]_  = A266 & A265;
  assign \new_[15524]_  = A235 & \new_[15523]_ ;
  assign \new_[15527]_  = A299 & ~A298;
  assign \new_[15530]_  = ~A302 & A300;
  assign \new_[15531]_  = \new_[15530]_  & \new_[15527]_ ;
  assign \new_[15532]_  = \new_[15531]_  & \new_[15524]_ ;
  assign \new_[15536]_  = ~A167 & A168;
  assign \new_[15537]_  = A170 & \new_[15536]_ ;
  assign \new_[15540]_  = ~A232 & A166;
  assign \new_[15543]_  = A234 & A233;
  assign \new_[15544]_  = \new_[15543]_  & \new_[15540]_ ;
  assign \new_[15545]_  = \new_[15544]_  & \new_[15537]_ ;
  assign \new_[15549]_  = ~A266 & ~A265;
  assign \new_[15550]_  = A235 & \new_[15549]_ ;
  assign \new_[15553]_  = ~A299 & A298;
  assign \new_[15556]_  = A301 & A300;
  assign \new_[15557]_  = \new_[15556]_  & \new_[15553]_ ;
  assign \new_[15558]_  = \new_[15557]_  & \new_[15550]_ ;
  assign \new_[15562]_  = ~A167 & A168;
  assign \new_[15563]_  = A170 & \new_[15562]_ ;
  assign \new_[15566]_  = ~A232 & A166;
  assign \new_[15569]_  = A234 & A233;
  assign \new_[15570]_  = \new_[15569]_  & \new_[15566]_ ;
  assign \new_[15571]_  = \new_[15570]_  & \new_[15563]_ ;
  assign \new_[15575]_  = ~A266 & ~A265;
  assign \new_[15576]_  = A235 & \new_[15575]_ ;
  assign \new_[15579]_  = ~A299 & A298;
  assign \new_[15582]_  = ~A302 & A300;
  assign \new_[15583]_  = \new_[15582]_  & \new_[15579]_ ;
  assign \new_[15584]_  = \new_[15583]_  & \new_[15576]_ ;
  assign \new_[15588]_  = ~A167 & A168;
  assign \new_[15589]_  = A170 & \new_[15588]_ ;
  assign \new_[15592]_  = ~A232 & A166;
  assign \new_[15595]_  = A234 & A233;
  assign \new_[15596]_  = \new_[15595]_  & \new_[15592]_ ;
  assign \new_[15597]_  = \new_[15596]_  & \new_[15589]_ ;
  assign \new_[15601]_  = ~A266 & ~A265;
  assign \new_[15602]_  = A235 & \new_[15601]_ ;
  assign \new_[15605]_  = A299 & ~A298;
  assign \new_[15608]_  = A301 & A300;
  assign \new_[15609]_  = \new_[15608]_  & \new_[15605]_ ;
  assign \new_[15610]_  = \new_[15609]_  & \new_[15602]_ ;
  assign \new_[15614]_  = ~A167 & A168;
  assign \new_[15615]_  = A170 & \new_[15614]_ ;
  assign \new_[15618]_  = ~A232 & A166;
  assign \new_[15621]_  = A234 & A233;
  assign \new_[15622]_  = \new_[15621]_  & \new_[15618]_ ;
  assign \new_[15623]_  = \new_[15622]_  & \new_[15615]_ ;
  assign \new_[15627]_  = ~A266 & ~A265;
  assign \new_[15628]_  = A235 & \new_[15627]_ ;
  assign \new_[15631]_  = A299 & ~A298;
  assign \new_[15634]_  = ~A302 & A300;
  assign \new_[15635]_  = \new_[15634]_  & \new_[15631]_ ;
  assign \new_[15636]_  = \new_[15635]_  & \new_[15628]_ ;
  assign \new_[15640]_  = ~A167 & A168;
  assign \new_[15641]_  = A170 & \new_[15640]_ ;
  assign \new_[15644]_  = ~A232 & A166;
  assign \new_[15647]_  = A234 & A233;
  assign \new_[15648]_  = \new_[15647]_  & \new_[15644]_ ;
  assign \new_[15649]_  = \new_[15648]_  & \new_[15641]_ ;
  assign \new_[15653]_  = A268 & ~A267;
  assign \new_[15654]_  = ~A236 & \new_[15653]_ ;
  assign \new_[15657]_  = ~A299 & A298;
  assign \new_[15660]_  = A301 & A300;
  assign \new_[15661]_  = \new_[15660]_  & \new_[15657]_ ;
  assign \new_[15662]_  = \new_[15661]_  & \new_[15654]_ ;
  assign \new_[15666]_  = ~A167 & A168;
  assign \new_[15667]_  = A170 & \new_[15666]_ ;
  assign \new_[15670]_  = ~A232 & A166;
  assign \new_[15673]_  = A234 & A233;
  assign \new_[15674]_  = \new_[15673]_  & \new_[15670]_ ;
  assign \new_[15675]_  = \new_[15674]_  & \new_[15667]_ ;
  assign \new_[15679]_  = A268 & ~A267;
  assign \new_[15680]_  = ~A236 & \new_[15679]_ ;
  assign \new_[15683]_  = ~A299 & A298;
  assign \new_[15686]_  = ~A302 & A300;
  assign \new_[15687]_  = \new_[15686]_  & \new_[15683]_ ;
  assign \new_[15688]_  = \new_[15687]_  & \new_[15680]_ ;
  assign \new_[15692]_  = ~A167 & A168;
  assign \new_[15693]_  = A170 & \new_[15692]_ ;
  assign \new_[15696]_  = ~A232 & A166;
  assign \new_[15699]_  = A234 & A233;
  assign \new_[15700]_  = \new_[15699]_  & \new_[15696]_ ;
  assign \new_[15701]_  = \new_[15700]_  & \new_[15693]_ ;
  assign \new_[15705]_  = A268 & ~A267;
  assign \new_[15706]_  = ~A236 & \new_[15705]_ ;
  assign \new_[15709]_  = A299 & ~A298;
  assign \new_[15712]_  = A301 & A300;
  assign \new_[15713]_  = \new_[15712]_  & \new_[15709]_ ;
  assign \new_[15714]_  = \new_[15713]_  & \new_[15706]_ ;
  assign \new_[15718]_  = ~A167 & A168;
  assign \new_[15719]_  = A170 & \new_[15718]_ ;
  assign \new_[15722]_  = ~A232 & A166;
  assign \new_[15725]_  = A234 & A233;
  assign \new_[15726]_  = \new_[15725]_  & \new_[15722]_ ;
  assign \new_[15727]_  = \new_[15726]_  & \new_[15719]_ ;
  assign \new_[15731]_  = A268 & ~A267;
  assign \new_[15732]_  = ~A236 & \new_[15731]_ ;
  assign \new_[15735]_  = A299 & ~A298;
  assign \new_[15738]_  = ~A302 & A300;
  assign \new_[15739]_  = \new_[15738]_  & \new_[15735]_ ;
  assign \new_[15740]_  = \new_[15739]_  & \new_[15732]_ ;
  assign \new_[15744]_  = ~A167 & A168;
  assign \new_[15745]_  = A170 & \new_[15744]_ ;
  assign \new_[15748]_  = ~A232 & A166;
  assign \new_[15751]_  = A234 & A233;
  assign \new_[15752]_  = \new_[15751]_  & \new_[15748]_ ;
  assign \new_[15753]_  = \new_[15752]_  & \new_[15745]_ ;
  assign \new_[15757]_  = ~A269 & ~A267;
  assign \new_[15758]_  = ~A236 & \new_[15757]_ ;
  assign \new_[15761]_  = ~A299 & A298;
  assign \new_[15764]_  = A301 & A300;
  assign \new_[15765]_  = \new_[15764]_  & \new_[15761]_ ;
  assign \new_[15766]_  = \new_[15765]_  & \new_[15758]_ ;
  assign \new_[15770]_  = ~A167 & A168;
  assign \new_[15771]_  = A170 & \new_[15770]_ ;
  assign \new_[15774]_  = ~A232 & A166;
  assign \new_[15777]_  = A234 & A233;
  assign \new_[15778]_  = \new_[15777]_  & \new_[15774]_ ;
  assign \new_[15779]_  = \new_[15778]_  & \new_[15771]_ ;
  assign \new_[15783]_  = ~A269 & ~A267;
  assign \new_[15784]_  = ~A236 & \new_[15783]_ ;
  assign \new_[15787]_  = ~A299 & A298;
  assign \new_[15790]_  = ~A302 & A300;
  assign \new_[15791]_  = \new_[15790]_  & \new_[15787]_ ;
  assign \new_[15792]_  = \new_[15791]_  & \new_[15784]_ ;
  assign \new_[15796]_  = ~A167 & A168;
  assign \new_[15797]_  = A170 & \new_[15796]_ ;
  assign \new_[15800]_  = ~A232 & A166;
  assign \new_[15803]_  = A234 & A233;
  assign \new_[15804]_  = \new_[15803]_  & \new_[15800]_ ;
  assign \new_[15805]_  = \new_[15804]_  & \new_[15797]_ ;
  assign \new_[15809]_  = ~A269 & ~A267;
  assign \new_[15810]_  = ~A236 & \new_[15809]_ ;
  assign \new_[15813]_  = A299 & ~A298;
  assign \new_[15816]_  = A301 & A300;
  assign \new_[15817]_  = \new_[15816]_  & \new_[15813]_ ;
  assign \new_[15818]_  = \new_[15817]_  & \new_[15810]_ ;
  assign \new_[15822]_  = ~A167 & A168;
  assign \new_[15823]_  = A170 & \new_[15822]_ ;
  assign \new_[15826]_  = ~A232 & A166;
  assign \new_[15829]_  = A234 & A233;
  assign \new_[15830]_  = \new_[15829]_  & \new_[15826]_ ;
  assign \new_[15831]_  = \new_[15830]_  & \new_[15823]_ ;
  assign \new_[15835]_  = ~A269 & ~A267;
  assign \new_[15836]_  = ~A236 & \new_[15835]_ ;
  assign \new_[15839]_  = A299 & ~A298;
  assign \new_[15842]_  = ~A302 & A300;
  assign \new_[15843]_  = \new_[15842]_  & \new_[15839]_ ;
  assign \new_[15844]_  = \new_[15843]_  & \new_[15836]_ ;
  assign \new_[15848]_  = ~A167 & A168;
  assign \new_[15849]_  = A170 & \new_[15848]_ ;
  assign \new_[15852]_  = ~A232 & A166;
  assign \new_[15855]_  = A234 & A233;
  assign \new_[15856]_  = \new_[15855]_  & \new_[15852]_ ;
  assign \new_[15857]_  = \new_[15856]_  & \new_[15849]_ ;
  assign \new_[15861]_  = A266 & A265;
  assign \new_[15862]_  = ~A236 & \new_[15861]_ ;
  assign \new_[15865]_  = ~A299 & A298;
  assign \new_[15868]_  = A301 & A300;
  assign \new_[15869]_  = \new_[15868]_  & \new_[15865]_ ;
  assign \new_[15870]_  = \new_[15869]_  & \new_[15862]_ ;
  assign \new_[15874]_  = ~A167 & A168;
  assign \new_[15875]_  = A170 & \new_[15874]_ ;
  assign \new_[15878]_  = ~A232 & A166;
  assign \new_[15881]_  = A234 & A233;
  assign \new_[15882]_  = \new_[15881]_  & \new_[15878]_ ;
  assign \new_[15883]_  = \new_[15882]_  & \new_[15875]_ ;
  assign \new_[15887]_  = A266 & A265;
  assign \new_[15888]_  = ~A236 & \new_[15887]_ ;
  assign \new_[15891]_  = ~A299 & A298;
  assign \new_[15894]_  = ~A302 & A300;
  assign \new_[15895]_  = \new_[15894]_  & \new_[15891]_ ;
  assign \new_[15896]_  = \new_[15895]_  & \new_[15888]_ ;
  assign \new_[15900]_  = ~A167 & A168;
  assign \new_[15901]_  = A170 & \new_[15900]_ ;
  assign \new_[15904]_  = ~A232 & A166;
  assign \new_[15907]_  = A234 & A233;
  assign \new_[15908]_  = \new_[15907]_  & \new_[15904]_ ;
  assign \new_[15909]_  = \new_[15908]_  & \new_[15901]_ ;
  assign \new_[15913]_  = A266 & A265;
  assign \new_[15914]_  = ~A236 & \new_[15913]_ ;
  assign \new_[15917]_  = A299 & ~A298;
  assign \new_[15920]_  = A301 & A300;
  assign \new_[15921]_  = \new_[15920]_  & \new_[15917]_ ;
  assign \new_[15922]_  = \new_[15921]_  & \new_[15914]_ ;
  assign \new_[15926]_  = ~A167 & A168;
  assign \new_[15927]_  = A170 & \new_[15926]_ ;
  assign \new_[15930]_  = ~A232 & A166;
  assign \new_[15933]_  = A234 & A233;
  assign \new_[15934]_  = \new_[15933]_  & \new_[15930]_ ;
  assign \new_[15935]_  = \new_[15934]_  & \new_[15927]_ ;
  assign \new_[15939]_  = A266 & A265;
  assign \new_[15940]_  = ~A236 & \new_[15939]_ ;
  assign \new_[15943]_  = A299 & ~A298;
  assign \new_[15946]_  = ~A302 & A300;
  assign \new_[15947]_  = \new_[15946]_  & \new_[15943]_ ;
  assign \new_[15948]_  = \new_[15947]_  & \new_[15940]_ ;
  assign \new_[15952]_  = ~A167 & A168;
  assign \new_[15953]_  = A170 & \new_[15952]_ ;
  assign \new_[15956]_  = ~A232 & A166;
  assign \new_[15959]_  = A234 & A233;
  assign \new_[15960]_  = \new_[15959]_  & \new_[15956]_ ;
  assign \new_[15961]_  = \new_[15960]_  & \new_[15953]_ ;
  assign \new_[15965]_  = ~A266 & ~A265;
  assign \new_[15966]_  = ~A236 & \new_[15965]_ ;
  assign \new_[15969]_  = ~A299 & A298;
  assign \new_[15972]_  = A301 & A300;
  assign \new_[15973]_  = \new_[15972]_  & \new_[15969]_ ;
  assign \new_[15974]_  = \new_[15973]_  & \new_[15966]_ ;
  assign \new_[15978]_  = ~A167 & A168;
  assign \new_[15979]_  = A170 & \new_[15978]_ ;
  assign \new_[15982]_  = ~A232 & A166;
  assign \new_[15985]_  = A234 & A233;
  assign \new_[15986]_  = \new_[15985]_  & \new_[15982]_ ;
  assign \new_[15987]_  = \new_[15986]_  & \new_[15979]_ ;
  assign \new_[15991]_  = ~A266 & ~A265;
  assign \new_[15992]_  = ~A236 & \new_[15991]_ ;
  assign \new_[15995]_  = ~A299 & A298;
  assign \new_[15998]_  = ~A302 & A300;
  assign \new_[15999]_  = \new_[15998]_  & \new_[15995]_ ;
  assign \new_[16000]_  = \new_[15999]_  & \new_[15992]_ ;
  assign \new_[16004]_  = ~A167 & A168;
  assign \new_[16005]_  = A170 & \new_[16004]_ ;
  assign \new_[16008]_  = ~A232 & A166;
  assign \new_[16011]_  = A234 & A233;
  assign \new_[16012]_  = \new_[16011]_  & \new_[16008]_ ;
  assign \new_[16013]_  = \new_[16012]_  & \new_[16005]_ ;
  assign \new_[16017]_  = ~A266 & ~A265;
  assign \new_[16018]_  = ~A236 & \new_[16017]_ ;
  assign \new_[16021]_  = A299 & ~A298;
  assign \new_[16024]_  = A301 & A300;
  assign \new_[16025]_  = \new_[16024]_  & \new_[16021]_ ;
  assign \new_[16026]_  = \new_[16025]_  & \new_[16018]_ ;
  assign \new_[16030]_  = ~A167 & A168;
  assign \new_[16031]_  = A170 & \new_[16030]_ ;
  assign \new_[16034]_  = ~A232 & A166;
  assign \new_[16037]_  = A234 & A233;
  assign \new_[16038]_  = \new_[16037]_  & \new_[16034]_ ;
  assign \new_[16039]_  = \new_[16038]_  & \new_[16031]_ ;
  assign \new_[16043]_  = ~A266 & ~A265;
  assign \new_[16044]_  = ~A236 & \new_[16043]_ ;
  assign \new_[16047]_  = A299 & ~A298;
  assign \new_[16050]_  = ~A302 & A300;
  assign \new_[16051]_  = \new_[16050]_  & \new_[16047]_ ;
  assign \new_[16052]_  = \new_[16051]_  & \new_[16044]_ ;
  assign \new_[16056]_  = ~A167 & A168;
  assign \new_[16057]_  = A170 & \new_[16056]_ ;
  assign \new_[16060]_  = A232 & A166;
  assign \new_[16063]_  = A234 & ~A233;
  assign \new_[16064]_  = \new_[16063]_  & \new_[16060]_ ;
  assign \new_[16065]_  = \new_[16064]_  & \new_[16057]_ ;
  assign \new_[16069]_  = A268 & ~A267;
  assign \new_[16070]_  = A235 & \new_[16069]_ ;
  assign \new_[16073]_  = ~A299 & A298;
  assign \new_[16076]_  = A301 & A300;
  assign \new_[16077]_  = \new_[16076]_  & \new_[16073]_ ;
  assign \new_[16078]_  = \new_[16077]_  & \new_[16070]_ ;
  assign \new_[16082]_  = ~A167 & A168;
  assign \new_[16083]_  = A170 & \new_[16082]_ ;
  assign \new_[16086]_  = A232 & A166;
  assign \new_[16089]_  = A234 & ~A233;
  assign \new_[16090]_  = \new_[16089]_  & \new_[16086]_ ;
  assign \new_[16091]_  = \new_[16090]_  & \new_[16083]_ ;
  assign \new_[16095]_  = A268 & ~A267;
  assign \new_[16096]_  = A235 & \new_[16095]_ ;
  assign \new_[16099]_  = ~A299 & A298;
  assign \new_[16102]_  = ~A302 & A300;
  assign \new_[16103]_  = \new_[16102]_  & \new_[16099]_ ;
  assign \new_[16104]_  = \new_[16103]_  & \new_[16096]_ ;
  assign \new_[16108]_  = ~A167 & A168;
  assign \new_[16109]_  = A170 & \new_[16108]_ ;
  assign \new_[16112]_  = A232 & A166;
  assign \new_[16115]_  = A234 & ~A233;
  assign \new_[16116]_  = \new_[16115]_  & \new_[16112]_ ;
  assign \new_[16117]_  = \new_[16116]_  & \new_[16109]_ ;
  assign \new_[16121]_  = A268 & ~A267;
  assign \new_[16122]_  = A235 & \new_[16121]_ ;
  assign \new_[16125]_  = A299 & ~A298;
  assign \new_[16128]_  = A301 & A300;
  assign \new_[16129]_  = \new_[16128]_  & \new_[16125]_ ;
  assign \new_[16130]_  = \new_[16129]_  & \new_[16122]_ ;
  assign \new_[16134]_  = ~A167 & A168;
  assign \new_[16135]_  = A170 & \new_[16134]_ ;
  assign \new_[16138]_  = A232 & A166;
  assign \new_[16141]_  = A234 & ~A233;
  assign \new_[16142]_  = \new_[16141]_  & \new_[16138]_ ;
  assign \new_[16143]_  = \new_[16142]_  & \new_[16135]_ ;
  assign \new_[16147]_  = A268 & ~A267;
  assign \new_[16148]_  = A235 & \new_[16147]_ ;
  assign \new_[16151]_  = A299 & ~A298;
  assign \new_[16154]_  = ~A302 & A300;
  assign \new_[16155]_  = \new_[16154]_  & \new_[16151]_ ;
  assign \new_[16156]_  = \new_[16155]_  & \new_[16148]_ ;
  assign \new_[16160]_  = ~A167 & A168;
  assign \new_[16161]_  = A170 & \new_[16160]_ ;
  assign \new_[16164]_  = A232 & A166;
  assign \new_[16167]_  = A234 & ~A233;
  assign \new_[16168]_  = \new_[16167]_  & \new_[16164]_ ;
  assign \new_[16169]_  = \new_[16168]_  & \new_[16161]_ ;
  assign \new_[16173]_  = ~A269 & ~A267;
  assign \new_[16174]_  = A235 & \new_[16173]_ ;
  assign \new_[16177]_  = ~A299 & A298;
  assign \new_[16180]_  = A301 & A300;
  assign \new_[16181]_  = \new_[16180]_  & \new_[16177]_ ;
  assign \new_[16182]_  = \new_[16181]_  & \new_[16174]_ ;
  assign \new_[16186]_  = ~A167 & A168;
  assign \new_[16187]_  = A170 & \new_[16186]_ ;
  assign \new_[16190]_  = A232 & A166;
  assign \new_[16193]_  = A234 & ~A233;
  assign \new_[16194]_  = \new_[16193]_  & \new_[16190]_ ;
  assign \new_[16195]_  = \new_[16194]_  & \new_[16187]_ ;
  assign \new_[16199]_  = ~A269 & ~A267;
  assign \new_[16200]_  = A235 & \new_[16199]_ ;
  assign \new_[16203]_  = ~A299 & A298;
  assign \new_[16206]_  = ~A302 & A300;
  assign \new_[16207]_  = \new_[16206]_  & \new_[16203]_ ;
  assign \new_[16208]_  = \new_[16207]_  & \new_[16200]_ ;
  assign \new_[16212]_  = ~A167 & A168;
  assign \new_[16213]_  = A170 & \new_[16212]_ ;
  assign \new_[16216]_  = A232 & A166;
  assign \new_[16219]_  = A234 & ~A233;
  assign \new_[16220]_  = \new_[16219]_  & \new_[16216]_ ;
  assign \new_[16221]_  = \new_[16220]_  & \new_[16213]_ ;
  assign \new_[16225]_  = ~A269 & ~A267;
  assign \new_[16226]_  = A235 & \new_[16225]_ ;
  assign \new_[16229]_  = A299 & ~A298;
  assign \new_[16232]_  = A301 & A300;
  assign \new_[16233]_  = \new_[16232]_  & \new_[16229]_ ;
  assign \new_[16234]_  = \new_[16233]_  & \new_[16226]_ ;
  assign \new_[16238]_  = ~A167 & A168;
  assign \new_[16239]_  = A170 & \new_[16238]_ ;
  assign \new_[16242]_  = A232 & A166;
  assign \new_[16245]_  = A234 & ~A233;
  assign \new_[16246]_  = \new_[16245]_  & \new_[16242]_ ;
  assign \new_[16247]_  = \new_[16246]_  & \new_[16239]_ ;
  assign \new_[16251]_  = ~A269 & ~A267;
  assign \new_[16252]_  = A235 & \new_[16251]_ ;
  assign \new_[16255]_  = A299 & ~A298;
  assign \new_[16258]_  = ~A302 & A300;
  assign \new_[16259]_  = \new_[16258]_  & \new_[16255]_ ;
  assign \new_[16260]_  = \new_[16259]_  & \new_[16252]_ ;
  assign \new_[16264]_  = ~A167 & A168;
  assign \new_[16265]_  = A170 & \new_[16264]_ ;
  assign \new_[16268]_  = A232 & A166;
  assign \new_[16271]_  = A234 & ~A233;
  assign \new_[16272]_  = \new_[16271]_  & \new_[16268]_ ;
  assign \new_[16273]_  = \new_[16272]_  & \new_[16265]_ ;
  assign \new_[16277]_  = A266 & A265;
  assign \new_[16278]_  = A235 & \new_[16277]_ ;
  assign \new_[16281]_  = ~A299 & A298;
  assign \new_[16284]_  = A301 & A300;
  assign \new_[16285]_  = \new_[16284]_  & \new_[16281]_ ;
  assign \new_[16286]_  = \new_[16285]_  & \new_[16278]_ ;
  assign \new_[16290]_  = ~A167 & A168;
  assign \new_[16291]_  = A170 & \new_[16290]_ ;
  assign \new_[16294]_  = A232 & A166;
  assign \new_[16297]_  = A234 & ~A233;
  assign \new_[16298]_  = \new_[16297]_  & \new_[16294]_ ;
  assign \new_[16299]_  = \new_[16298]_  & \new_[16291]_ ;
  assign \new_[16303]_  = A266 & A265;
  assign \new_[16304]_  = A235 & \new_[16303]_ ;
  assign \new_[16307]_  = ~A299 & A298;
  assign \new_[16310]_  = ~A302 & A300;
  assign \new_[16311]_  = \new_[16310]_  & \new_[16307]_ ;
  assign \new_[16312]_  = \new_[16311]_  & \new_[16304]_ ;
  assign \new_[16316]_  = ~A167 & A168;
  assign \new_[16317]_  = A170 & \new_[16316]_ ;
  assign \new_[16320]_  = A232 & A166;
  assign \new_[16323]_  = A234 & ~A233;
  assign \new_[16324]_  = \new_[16323]_  & \new_[16320]_ ;
  assign \new_[16325]_  = \new_[16324]_  & \new_[16317]_ ;
  assign \new_[16329]_  = A266 & A265;
  assign \new_[16330]_  = A235 & \new_[16329]_ ;
  assign \new_[16333]_  = A299 & ~A298;
  assign \new_[16336]_  = A301 & A300;
  assign \new_[16337]_  = \new_[16336]_  & \new_[16333]_ ;
  assign \new_[16338]_  = \new_[16337]_  & \new_[16330]_ ;
  assign \new_[16342]_  = ~A167 & A168;
  assign \new_[16343]_  = A170 & \new_[16342]_ ;
  assign \new_[16346]_  = A232 & A166;
  assign \new_[16349]_  = A234 & ~A233;
  assign \new_[16350]_  = \new_[16349]_  & \new_[16346]_ ;
  assign \new_[16351]_  = \new_[16350]_  & \new_[16343]_ ;
  assign \new_[16355]_  = A266 & A265;
  assign \new_[16356]_  = A235 & \new_[16355]_ ;
  assign \new_[16359]_  = A299 & ~A298;
  assign \new_[16362]_  = ~A302 & A300;
  assign \new_[16363]_  = \new_[16362]_  & \new_[16359]_ ;
  assign \new_[16364]_  = \new_[16363]_  & \new_[16356]_ ;
  assign \new_[16368]_  = ~A167 & A168;
  assign \new_[16369]_  = A170 & \new_[16368]_ ;
  assign \new_[16372]_  = A232 & A166;
  assign \new_[16375]_  = A234 & ~A233;
  assign \new_[16376]_  = \new_[16375]_  & \new_[16372]_ ;
  assign \new_[16377]_  = \new_[16376]_  & \new_[16369]_ ;
  assign \new_[16381]_  = ~A266 & ~A265;
  assign \new_[16382]_  = A235 & \new_[16381]_ ;
  assign \new_[16385]_  = ~A299 & A298;
  assign \new_[16388]_  = A301 & A300;
  assign \new_[16389]_  = \new_[16388]_  & \new_[16385]_ ;
  assign \new_[16390]_  = \new_[16389]_  & \new_[16382]_ ;
  assign \new_[16394]_  = ~A167 & A168;
  assign \new_[16395]_  = A170 & \new_[16394]_ ;
  assign \new_[16398]_  = A232 & A166;
  assign \new_[16401]_  = A234 & ~A233;
  assign \new_[16402]_  = \new_[16401]_  & \new_[16398]_ ;
  assign \new_[16403]_  = \new_[16402]_  & \new_[16395]_ ;
  assign \new_[16407]_  = ~A266 & ~A265;
  assign \new_[16408]_  = A235 & \new_[16407]_ ;
  assign \new_[16411]_  = ~A299 & A298;
  assign \new_[16414]_  = ~A302 & A300;
  assign \new_[16415]_  = \new_[16414]_  & \new_[16411]_ ;
  assign \new_[16416]_  = \new_[16415]_  & \new_[16408]_ ;
  assign \new_[16420]_  = ~A167 & A168;
  assign \new_[16421]_  = A170 & \new_[16420]_ ;
  assign \new_[16424]_  = A232 & A166;
  assign \new_[16427]_  = A234 & ~A233;
  assign \new_[16428]_  = \new_[16427]_  & \new_[16424]_ ;
  assign \new_[16429]_  = \new_[16428]_  & \new_[16421]_ ;
  assign \new_[16433]_  = ~A266 & ~A265;
  assign \new_[16434]_  = A235 & \new_[16433]_ ;
  assign \new_[16437]_  = A299 & ~A298;
  assign \new_[16440]_  = A301 & A300;
  assign \new_[16441]_  = \new_[16440]_  & \new_[16437]_ ;
  assign \new_[16442]_  = \new_[16441]_  & \new_[16434]_ ;
  assign \new_[16446]_  = ~A167 & A168;
  assign \new_[16447]_  = A170 & \new_[16446]_ ;
  assign \new_[16450]_  = A232 & A166;
  assign \new_[16453]_  = A234 & ~A233;
  assign \new_[16454]_  = \new_[16453]_  & \new_[16450]_ ;
  assign \new_[16455]_  = \new_[16454]_  & \new_[16447]_ ;
  assign \new_[16459]_  = ~A266 & ~A265;
  assign \new_[16460]_  = A235 & \new_[16459]_ ;
  assign \new_[16463]_  = A299 & ~A298;
  assign \new_[16466]_  = ~A302 & A300;
  assign \new_[16467]_  = \new_[16466]_  & \new_[16463]_ ;
  assign \new_[16468]_  = \new_[16467]_  & \new_[16460]_ ;
  assign \new_[16472]_  = ~A167 & A168;
  assign \new_[16473]_  = A170 & \new_[16472]_ ;
  assign \new_[16476]_  = A232 & A166;
  assign \new_[16479]_  = A234 & ~A233;
  assign \new_[16480]_  = \new_[16479]_  & \new_[16476]_ ;
  assign \new_[16481]_  = \new_[16480]_  & \new_[16473]_ ;
  assign \new_[16485]_  = A268 & ~A267;
  assign \new_[16486]_  = ~A236 & \new_[16485]_ ;
  assign \new_[16489]_  = ~A299 & A298;
  assign \new_[16492]_  = A301 & A300;
  assign \new_[16493]_  = \new_[16492]_  & \new_[16489]_ ;
  assign \new_[16494]_  = \new_[16493]_  & \new_[16486]_ ;
  assign \new_[16498]_  = ~A167 & A168;
  assign \new_[16499]_  = A170 & \new_[16498]_ ;
  assign \new_[16502]_  = A232 & A166;
  assign \new_[16505]_  = A234 & ~A233;
  assign \new_[16506]_  = \new_[16505]_  & \new_[16502]_ ;
  assign \new_[16507]_  = \new_[16506]_  & \new_[16499]_ ;
  assign \new_[16511]_  = A268 & ~A267;
  assign \new_[16512]_  = ~A236 & \new_[16511]_ ;
  assign \new_[16515]_  = ~A299 & A298;
  assign \new_[16518]_  = ~A302 & A300;
  assign \new_[16519]_  = \new_[16518]_  & \new_[16515]_ ;
  assign \new_[16520]_  = \new_[16519]_  & \new_[16512]_ ;
  assign \new_[16524]_  = ~A167 & A168;
  assign \new_[16525]_  = A170 & \new_[16524]_ ;
  assign \new_[16528]_  = A232 & A166;
  assign \new_[16531]_  = A234 & ~A233;
  assign \new_[16532]_  = \new_[16531]_  & \new_[16528]_ ;
  assign \new_[16533]_  = \new_[16532]_  & \new_[16525]_ ;
  assign \new_[16537]_  = A268 & ~A267;
  assign \new_[16538]_  = ~A236 & \new_[16537]_ ;
  assign \new_[16541]_  = A299 & ~A298;
  assign \new_[16544]_  = A301 & A300;
  assign \new_[16545]_  = \new_[16544]_  & \new_[16541]_ ;
  assign \new_[16546]_  = \new_[16545]_  & \new_[16538]_ ;
  assign \new_[16550]_  = ~A167 & A168;
  assign \new_[16551]_  = A170 & \new_[16550]_ ;
  assign \new_[16554]_  = A232 & A166;
  assign \new_[16557]_  = A234 & ~A233;
  assign \new_[16558]_  = \new_[16557]_  & \new_[16554]_ ;
  assign \new_[16559]_  = \new_[16558]_  & \new_[16551]_ ;
  assign \new_[16563]_  = A268 & ~A267;
  assign \new_[16564]_  = ~A236 & \new_[16563]_ ;
  assign \new_[16567]_  = A299 & ~A298;
  assign \new_[16570]_  = ~A302 & A300;
  assign \new_[16571]_  = \new_[16570]_  & \new_[16567]_ ;
  assign \new_[16572]_  = \new_[16571]_  & \new_[16564]_ ;
  assign \new_[16576]_  = ~A167 & A168;
  assign \new_[16577]_  = A170 & \new_[16576]_ ;
  assign \new_[16580]_  = A232 & A166;
  assign \new_[16583]_  = A234 & ~A233;
  assign \new_[16584]_  = \new_[16583]_  & \new_[16580]_ ;
  assign \new_[16585]_  = \new_[16584]_  & \new_[16577]_ ;
  assign \new_[16589]_  = ~A269 & ~A267;
  assign \new_[16590]_  = ~A236 & \new_[16589]_ ;
  assign \new_[16593]_  = ~A299 & A298;
  assign \new_[16596]_  = A301 & A300;
  assign \new_[16597]_  = \new_[16596]_  & \new_[16593]_ ;
  assign \new_[16598]_  = \new_[16597]_  & \new_[16590]_ ;
  assign \new_[16602]_  = ~A167 & A168;
  assign \new_[16603]_  = A170 & \new_[16602]_ ;
  assign \new_[16606]_  = A232 & A166;
  assign \new_[16609]_  = A234 & ~A233;
  assign \new_[16610]_  = \new_[16609]_  & \new_[16606]_ ;
  assign \new_[16611]_  = \new_[16610]_  & \new_[16603]_ ;
  assign \new_[16615]_  = ~A269 & ~A267;
  assign \new_[16616]_  = ~A236 & \new_[16615]_ ;
  assign \new_[16619]_  = ~A299 & A298;
  assign \new_[16622]_  = ~A302 & A300;
  assign \new_[16623]_  = \new_[16622]_  & \new_[16619]_ ;
  assign \new_[16624]_  = \new_[16623]_  & \new_[16616]_ ;
  assign \new_[16628]_  = ~A167 & A168;
  assign \new_[16629]_  = A170 & \new_[16628]_ ;
  assign \new_[16632]_  = A232 & A166;
  assign \new_[16635]_  = A234 & ~A233;
  assign \new_[16636]_  = \new_[16635]_  & \new_[16632]_ ;
  assign \new_[16637]_  = \new_[16636]_  & \new_[16629]_ ;
  assign \new_[16641]_  = ~A269 & ~A267;
  assign \new_[16642]_  = ~A236 & \new_[16641]_ ;
  assign \new_[16645]_  = A299 & ~A298;
  assign \new_[16648]_  = A301 & A300;
  assign \new_[16649]_  = \new_[16648]_  & \new_[16645]_ ;
  assign \new_[16650]_  = \new_[16649]_  & \new_[16642]_ ;
  assign \new_[16654]_  = ~A167 & A168;
  assign \new_[16655]_  = A170 & \new_[16654]_ ;
  assign \new_[16658]_  = A232 & A166;
  assign \new_[16661]_  = A234 & ~A233;
  assign \new_[16662]_  = \new_[16661]_  & \new_[16658]_ ;
  assign \new_[16663]_  = \new_[16662]_  & \new_[16655]_ ;
  assign \new_[16667]_  = ~A269 & ~A267;
  assign \new_[16668]_  = ~A236 & \new_[16667]_ ;
  assign \new_[16671]_  = A299 & ~A298;
  assign \new_[16674]_  = ~A302 & A300;
  assign \new_[16675]_  = \new_[16674]_  & \new_[16671]_ ;
  assign \new_[16676]_  = \new_[16675]_  & \new_[16668]_ ;
  assign \new_[16680]_  = ~A167 & A168;
  assign \new_[16681]_  = A170 & \new_[16680]_ ;
  assign \new_[16684]_  = A232 & A166;
  assign \new_[16687]_  = A234 & ~A233;
  assign \new_[16688]_  = \new_[16687]_  & \new_[16684]_ ;
  assign \new_[16689]_  = \new_[16688]_  & \new_[16681]_ ;
  assign \new_[16693]_  = A266 & A265;
  assign \new_[16694]_  = ~A236 & \new_[16693]_ ;
  assign \new_[16697]_  = ~A299 & A298;
  assign \new_[16700]_  = A301 & A300;
  assign \new_[16701]_  = \new_[16700]_  & \new_[16697]_ ;
  assign \new_[16702]_  = \new_[16701]_  & \new_[16694]_ ;
  assign \new_[16706]_  = ~A167 & A168;
  assign \new_[16707]_  = A170 & \new_[16706]_ ;
  assign \new_[16710]_  = A232 & A166;
  assign \new_[16713]_  = A234 & ~A233;
  assign \new_[16714]_  = \new_[16713]_  & \new_[16710]_ ;
  assign \new_[16715]_  = \new_[16714]_  & \new_[16707]_ ;
  assign \new_[16719]_  = A266 & A265;
  assign \new_[16720]_  = ~A236 & \new_[16719]_ ;
  assign \new_[16723]_  = ~A299 & A298;
  assign \new_[16726]_  = ~A302 & A300;
  assign \new_[16727]_  = \new_[16726]_  & \new_[16723]_ ;
  assign \new_[16728]_  = \new_[16727]_  & \new_[16720]_ ;
  assign \new_[16732]_  = ~A167 & A168;
  assign \new_[16733]_  = A170 & \new_[16732]_ ;
  assign \new_[16736]_  = A232 & A166;
  assign \new_[16739]_  = A234 & ~A233;
  assign \new_[16740]_  = \new_[16739]_  & \new_[16736]_ ;
  assign \new_[16741]_  = \new_[16740]_  & \new_[16733]_ ;
  assign \new_[16745]_  = A266 & A265;
  assign \new_[16746]_  = ~A236 & \new_[16745]_ ;
  assign \new_[16749]_  = A299 & ~A298;
  assign \new_[16752]_  = A301 & A300;
  assign \new_[16753]_  = \new_[16752]_  & \new_[16749]_ ;
  assign \new_[16754]_  = \new_[16753]_  & \new_[16746]_ ;
  assign \new_[16758]_  = ~A167 & A168;
  assign \new_[16759]_  = A170 & \new_[16758]_ ;
  assign \new_[16762]_  = A232 & A166;
  assign \new_[16765]_  = A234 & ~A233;
  assign \new_[16766]_  = \new_[16765]_  & \new_[16762]_ ;
  assign \new_[16767]_  = \new_[16766]_  & \new_[16759]_ ;
  assign \new_[16771]_  = A266 & A265;
  assign \new_[16772]_  = ~A236 & \new_[16771]_ ;
  assign \new_[16775]_  = A299 & ~A298;
  assign \new_[16778]_  = ~A302 & A300;
  assign \new_[16779]_  = \new_[16778]_  & \new_[16775]_ ;
  assign \new_[16780]_  = \new_[16779]_  & \new_[16772]_ ;
  assign \new_[16784]_  = ~A167 & A168;
  assign \new_[16785]_  = A170 & \new_[16784]_ ;
  assign \new_[16788]_  = A232 & A166;
  assign \new_[16791]_  = A234 & ~A233;
  assign \new_[16792]_  = \new_[16791]_  & \new_[16788]_ ;
  assign \new_[16793]_  = \new_[16792]_  & \new_[16785]_ ;
  assign \new_[16797]_  = ~A266 & ~A265;
  assign \new_[16798]_  = ~A236 & \new_[16797]_ ;
  assign \new_[16801]_  = ~A299 & A298;
  assign \new_[16804]_  = A301 & A300;
  assign \new_[16805]_  = \new_[16804]_  & \new_[16801]_ ;
  assign \new_[16806]_  = \new_[16805]_  & \new_[16798]_ ;
  assign \new_[16810]_  = ~A167 & A168;
  assign \new_[16811]_  = A170 & \new_[16810]_ ;
  assign \new_[16814]_  = A232 & A166;
  assign \new_[16817]_  = A234 & ~A233;
  assign \new_[16818]_  = \new_[16817]_  & \new_[16814]_ ;
  assign \new_[16819]_  = \new_[16818]_  & \new_[16811]_ ;
  assign \new_[16823]_  = ~A266 & ~A265;
  assign \new_[16824]_  = ~A236 & \new_[16823]_ ;
  assign \new_[16827]_  = ~A299 & A298;
  assign \new_[16830]_  = ~A302 & A300;
  assign \new_[16831]_  = \new_[16830]_  & \new_[16827]_ ;
  assign \new_[16832]_  = \new_[16831]_  & \new_[16824]_ ;
  assign \new_[16836]_  = ~A167 & A168;
  assign \new_[16837]_  = A170 & \new_[16836]_ ;
  assign \new_[16840]_  = A232 & A166;
  assign \new_[16843]_  = A234 & ~A233;
  assign \new_[16844]_  = \new_[16843]_  & \new_[16840]_ ;
  assign \new_[16845]_  = \new_[16844]_  & \new_[16837]_ ;
  assign \new_[16849]_  = ~A266 & ~A265;
  assign \new_[16850]_  = ~A236 & \new_[16849]_ ;
  assign \new_[16853]_  = A299 & ~A298;
  assign \new_[16856]_  = A301 & A300;
  assign \new_[16857]_  = \new_[16856]_  & \new_[16853]_ ;
  assign \new_[16858]_  = \new_[16857]_  & \new_[16850]_ ;
  assign \new_[16862]_  = ~A167 & A168;
  assign \new_[16863]_  = A170 & \new_[16862]_ ;
  assign \new_[16866]_  = A232 & A166;
  assign \new_[16869]_  = A234 & ~A233;
  assign \new_[16870]_  = \new_[16869]_  & \new_[16866]_ ;
  assign \new_[16871]_  = \new_[16870]_  & \new_[16863]_ ;
  assign \new_[16875]_  = ~A266 & ~A265;
  assign \new_[16876]_  = ~A236 & \new_[16875]_ ;
  assign \new_[16879]_  = A299 & ~A298;
  assign \new_[16882]_  = ~A302 & A300;
  assign \new_[16883]_  = \new_[16882]_  & \new_[16879]_ ;
  assign \new_[16884]_  = \new_[16883]_  & \new_[16876]_ ;
  assign \new_[16888]_  = A167 & A168;
  assign \new_[16889]_  = A169 & \new_[16888]_ ;
  assign \new_[16892]_  = ~A232 & ~A166;
  assign \new_[16895]_  = A234 & A233;
  assign \new_[16896]_  = \new_[16895]_  & \new_[16892]_ ;
  assign \new_[16897]_  = \new_[16896]_  & \new_[16889]_ ;
  assign \new_[16901]_  = A268 & ~A267;
  assign \new_[16902]_  = A235 & \new_[16901]_ ;
  assign \new_[16905]_  = ~A299 & A298;
  assign \new_[16908]_  = A301 & A300;
  assign \new_[16909]_  = \new_[16908]_  & \new_[16905]_ ;
  assign \new_[16910]_  = \new_[16909]_  & \new_[16902]_ ;
  assign \new_[16914]_  = A167 & A168;
  assign \new_[16915]_  = A169 & \new_[16914]_ ;
  assign \new_[16918]_  = ~A232 & ~A166;
  assign \new_[16921]_  = A234 & A233;
  assign \new_[16922]_  = \new_[16921]_  & \new_[16918]_ ;
  assign \new_[16923]_  = \new_[16922]_  & \new_[16915]_ ;
  assign \new_[16927]_  = A268 & ~A267;
  assign \new_[16928]_  = A235 & \new_[16927]_ ;
  assign \new_[16931]_  = ~A299 & A298;
  assign \new_[16934]_  = ~A302 & A300;
  assign \new_[16935]_  = \new_[16934]_  & \new_[16931]_ ;
  assign \new_[16936]_  = \new_[16935]_  & \new_[16928]_ ;
  assign \new_[16940]_  = A167 & A168;
  assign \new_[16941]_  = A169 & \new_[16940]_ ;
  assign \new_[16944]_  = ~A232 & ~A166;
  assign \new_[16947]_  = A234 & A233;
  assign \new_[16948]_  = \new_[16947]_  & \new_[16944]_ ;
  assign \new_[16949]_  = \new_[16948]_  & \new_[16941]_ ;
  assign \new_[16953]_  = A268 & ~A267;
  assign \new_[16954]_  = A235 & \new_[16953]_ ;
  assign \new_[16957]_  = A299 & ~A298;
  assign \new_[16960]_  = A301 & A300;
  assign \new_[16961]_  = \new_[16960]_  & \new_[16957]_ ;
  assign \new_[16962]_  = \new_[16961]_  & \new_[16954]_ ;
  assign \new_[16966]_  = A167 & A168;
  assign \new_[16967]_  = A169 & \new_[16966]_ ;
  assign \new_[16970]_  = ~A232 & ~A166;
  assign \new_[16973]_  = A234 & A233;
  assign \new_[16974]_  = \new_[16973]_  & \new_[16970]_ ;
  assign \new_[16975]_  = \new_[16974]_  & \new_[16967]_ ;
  assign \new_[16979]_  = A268 & ~A267;
  assign \new_[16980]_  = A235 & \new_[16979]_ ;
  assign \new_[16983]_  = A299 & ~A298;
  assign \new_[16986]_  = ~A302 & A300;
  assign \new_[16987]_  = \new_[16986]_  & \new_[16983]_ ;
  assign \new_[16988]_  = \new_[16987]_  & \new_[16980]_ ;
  assign \new_[16992]_  = A167 & A168;
  assign \new_[16993]_  = A169 & \new_[16992]_ ;
  assign \new_[16996]_  = ~A232 & ~A166;
  assign \new_[16999]_  = A234 & A233;
  assign \new_[17000]_  = \new_[16999]_  & \new_[16996]_ ;
  assign \new_[17001]_  = \new_[17000]_  & \new_[16993]_ ;
  assign \new_[17005]_  = ~A269 & ~A267;
  assign \new_[17006]_  = A235 & \new_[17005]_ ;
  assign \new_[17009]_  = ~A299 & A298;
  assign \new_[17012]_  = A301 & A300;
  assign \new_[17013]_  = \new_[17012]_  & \new_[17009]_ ;
  assign \new_[17014]_  = \new_[17013]_  & \new_[17006]_ ;
  assign \new_[17018]_  = A167 & A168;
  assign \new_[17019]_  = A169 & \new_[17018]_ ;
  assign \new_[17022]_  = ~A232 & ~A166;
  assign \new_[17025]_  = A234 & A233;
  assign \new_[17026]_  = \new_[17025]_  & \new_[17022]_ ;
  assign \new_[17027]_  = \new_[17026]_  & \new_[17019]_ ;
  assign \new_[17031]_  = ~A269 & ~A267;
  assign \new_[17032]_  = A235 & \new_[17031]_ ;
  assign \new_[17035]_  = ~A299 & A298;
  assign \new_[17038]_  = ~A302 & A300;
  assign \new_[17039]_  = \new_[17038]_  & \new_[17035]_ ;
  assign \new_[17040]_  = \new_[17039]_  & \new_[17032]_ ;
  assign \new_[17044]_  = A167 & A168;
  assign \new_[17045]_  = A169 & \new_[17044]_ ;
  assign \new_[17048]_  = ~A232 & ~A166;
  assign \new_[17051]_  = A234 & A233;
  assign \new_[17052]_  = \new_[17051]_  & \new_[17048]_ ;
  assign \new_[17053]_  = \new_[17052]_  & \new_[17045]_ ;
  assign \new_[17057]_  = ~A269 & ~A267;
  assign \new_[17058]_  = A235 & \new_[17057]_ ;
  assign \new_[17061]_  = A299 & ~A298;
  assign \new_[17064]_  = A301 & A300;
  assign \new_[17065]_  = \new_[17064]_  & \new_[17061]_ ;
  assign \new_[17066]_  = \new_[17065]_  & \new_[17058]_ ;
  assign \new_[17070]_  = A167 & A168;
  assign \new_[17071]_  = A169 & \new_[17070]_ ;
  assign \new_[17074]_  = ~A232 & ~A166;
  assign \new_[17077]_  = A234 & A233;
  assign \new_[17078]_  = \new_[17077]_  & \new_[17074]_ ;
  assign \new_[17079]_  = \new_[17078]_  & \new_[17071]_ ;
  assign \new_[17083]_  = ~A269 & ~A267;
  assign \new_[17084]_  = A235 & \new_[17083]_ ;
  assign \new_[17087]_  = A299 & ~A298;
  assign \new_[17090]_  = ~A302 & A300;
  assign \new_[17091]_  = \new_[17090]_  & \new_[17087]_ ;
  assign \new_[17092]_  = \new_[17091]_  & \new_[17084]_ ;
  assign \new_[17096]_  = A167 & A168;
  assign \new_[17097]_  = A169 & \new_[17096]_ ;
  assign \new_[17100]_  = ~A232 & ~A166;
  assign \new_[17103]_  = A234 & A233;
  assign \new_[17104]_  = \new_[17103]_  & \new_[17100]_ ;
  assign \new_[17105]_  = \new_[17104]_  & \new_[17097]_ ;
  assign \new_[17109]_  = A266 & A265;
  assign \new_[17110]_  = A235 & \new_[17109]_ ;
  assign \new_[17113]_  = ~A299 & A298;
  assign \new_[17116]_  = A301 & A300;
  assign \new_[17117]_  = \new_[17116]_  & \new_[17113]_ ;
  assign \new_[17118]_  = \new_[17117]_  & \new_[17110]_ ;
  assign \new_[17122]_  = A167 & A168;
  assign \new_[17123]_  = A169 & \new_[17122]_ ;
  assign \new_[17126]_  = ~A232 & ~A166;
  assign \new_[17129]_  = A234 & A233;
  assign \new_[17130]_  = \new_[17129]_  & \new_[17126]_ ;
  assign \new_[17131]_  = \new_[17130]_  & \new_[17123]_ ;
  assign \new_[17135]_  = A266 & A265;
  assign \new_[17136]_  = A235 & \new_[17135]_ ;
  assign \new_[17139]_  = ~A299 & A298;
  assign \new_[17142]_  = ~A302 & A300;
  assign \new_[17143]_  = \new_[17142]_  & \new_[17139]_ ;
  assign \new_[17144]_  = \new_[17143]_  & \new_[17136]_ ;
  assign \new_[17148]_  = A167 & A168;
  assign \new_[17149]_  = A169 & \new_[17148]_ ;
  assign \new_[17152]_  = ~A232 & ~A166;
  assign \new_[17155]_  = A234 & A233;
  assign \new_[17156]_  = \new_[17155]_  & \new_[17152]_ ;
  assign \new_[17157]_  = \new_[17156]_  & \new_[17149]_ ;
  assign \new_[17161]_  = A266 & A265;
  assign \new_[17162]_  = A235 & \new_[17161]_ ;
  assign \new_[17165]_  = A299 & ~A298;
  assign \new_[17168]_  = A301 & A300;
  assign \new_[17169]_  = \new_[17168]_  & \new_[17165]_ ;
  assign \new_[17170]_  = \new_[17169]_  & \new_[17162]_ ;
  assign \new_[17174]_  = A167 & A168;
  assign \new_[17175]_  = A169 & \new_[17174]_ ;
  assign \new_[17178]_  = ~A232 & ~A166;
  assign \new_[17181]_  = A234 & A233;
  assign \new_[17182]_  = \new_[17181]_  & \new_[17178]_ ;
  assign \new_[17183]_  = \new_[17182]_  & \new_[17175]_ ;
  assign \new_[17187]_  = A266 & A265;
  assign \new_[17188]_  = A235 & \new_[17187]_ ;
  assign \new_[17191]_  = A299 & ~A298;
  assign \new_[17194]_  = ~A302 & A300;
  assign \new_[17195]_  = \new_[17194]_  & \new_[17191]_ ;
  assign \new_[17196]_  = \new_[17195]_  & \new_[17188]_ ;
  assign \new_[17200]_  = A167 & A168;
  assign \new_[17201]_  = A169 & \new_[17200]_ ;
  assign \new_[17204]_  = ~A232 & ~A166;
  assign \new_[17207]_  = A234 & A233;
  assign \new_[17208]_  = \new_[17207]_  & \new_[17204]_ ;
  assign \new_[17209]_  = \new_[17208]_  & \new_[17201]_ ;
  assign \new_[17213]_  = ~A266 & ~A265;
  assign \new_[17214]_  = A235 & \new_[17213]_ ;
  assign \new_[17217]_  = ~A299 & A298;
  assign \new_[17220]_  = A301 & A300;
  assign \new_[17221]_  = \new_[17220]_  & \new_[17217]_ ;
  assign \new_[17222]_  = \new_[17221]_  & \new_[17214]_ ;
  assign \new_[17226]_  = A167 & A168;
  assign \new_[17227]_  = A169 & \new_[17226]_ ;
  assign \new_[17230]_  = ~A232 & ~A166;
  assign \new_[17233]_  = A234 & A233;
  assign \new_[17234]_  = \new_[17233]_  & \new_[17230]_ ;
  assign \new_[17235]_  = \new_[17234]_  & \new_[17227]_ ;
  assign \new_[17239]_  = ~A266 & ~A265;
  assign \new_[17240]_  = A235 & \new_[17239]_ ;
  assign \new_[17243]_  = ~A299 & A298;
  assign \new_[17246]_  = ~A302 & A300;
  assign \new_[17247]_  = \new_[17246]_  & \new_[17243]_ ;
  assign \new_[17248]_  = \new_[17247]_  & \new_[17240]_ ;
  assign \new_[17252]_  = A167 & A168;
  assign \new_[17253]_  = A169 & \new_[17252]_ ;
  assign \new_[17256]_  = ~A232 & ~A166;
  assign \new_[17259]_  = A234 & A233;
  assign \new_[17260]_  = \new_[17259]_  & \new_[17256]_ ;
  assign \new_[17261]_  = \new_[17260]_  & \new_[17253]_ ;
  assign \new_[17265]_  = ~A266 & ~A265;
  assign \new_[17266]_  = A235 & \new_[17265]_ ;
  assign \new_[17269]_  = A299 & ~A298;
  assign \new_[17272]_  = A301 & A300;
  assign \new_[17273]_  = \new_[17272]_  & \new_[17269]_ ;
  assign \new_[17274]_  = \new_[17273]_  & \new_[17266]_ ;
  assign \new_[17278]_  = A167 & A168;
  assign \new_[17279]_  = A169 & \new_[17278]_ ;
  assign \new_[17282]_  = ~A232 & ~A166;
  assign \new_[17285]_  = A234 & A233;
  assign \new_[17286]_  = \new_[17285]_  & \new_[17282]_ ;
  assign \new_[17287]_  = \new_[17286]_  & \new_[17279]_ ;
  assign \new_[17291]_  = ~A266 & ~A265;
  assign \new_[17292]_  = A235 & \new_[17291]_ ;
  assign \new_[17295]_  = A299 & ~A298;
  assign \new_[17298]_  = ~A302 & A300;
  assign \new_[17299]_  = \new_[17298]_  & \new_[17295]_ ;
  assign \new_[17300]_  = \new_[17299]_  & \new_[17292]_ ;
  assign \new_[17304]_  = A167 & A168;
  assign \new_[17305]_  = A169 & \new_[17304]_ ;
  assign \new_[17308]_  = ~A232 & ~A166;
  assign \new_[17311]_  = A234 & A233;
  assign \new_[17312]_  = \new_[17311]_  & \new_[17308]_ ;
  assign \new_[17313]_  = \new_[17312]_  & \new_[17305]_ ;
  assign \new_[17317]_  = A268 & ~A267;
  assign \new_[17318]_  = ~A236 & \new_[17317]_ ;
  assign \new_[17321]_  = ~A299 & A298;
  assign \new_[17324]_  = A301 & A300;
  assign \new_[17325]_  = \new_[17324]_  & \new_[17321]_ ;
  assign \new_[17326]_  = \new_[17325]_  & \new_[17318]_ ;
  assign \new_[17330]_  = A167 & A168;
  assign \new_[17331]_  = A169 & \new_[17330]_ ;
  assign \new_[17334]_  = ~A232 & ~A166;
  assign \new_[17337]_  = A234 & A233;
  assign \new_[17338]_  = \new_[17337]_  & \new_[17334]_ ;
  assign \new_[17339]_  = \new_[17338]_  & \new_[17331]_ ;
  assign \new_[17343]_  = A268 & ~A267;
  assign \new_[17344]_  = ~A236 & \new_[17343]_ ;
  assign \new_[17347]_  = ~A299 & A298;
  assign \new_[17350]_  = ~A302 & A300;
  assign \new_[17351]_  = \new_[17350]_  & \new_[17347]_ ;
  assign \new_[17352]_  = \new_[17351]_  & \new_[17344]_ ;
  assign \new_[17356]_  = A167 & A168;
  assign \new_[17357]_  = A169 & \new_[17356]_ ;
  assign \new_[17360]_  = ~A232 & ~A166;
  assign \new_[17363]_  = A234 & A233;
  assign \new_[17364]_  = \new_[17363]_  & \new_[17360]_ ;
  assign \new_[17365]_  = \new_[17364]_  & \new_[17357]_ ;
  assign \new_[17369]_  = A268 & ~A267;
  assign \new_[17370]_  = ~A236 & \new_[17369]_ ;
  assign \new_[17373]_  = A299 & ~A298;
  assign \new_[17376]_  = A301 & A300;
  assign \new_[17377]_  = \new_[17376]_  & \new_[17373]_ ;
  assign \new_[17378]_  = \new_[17377]_  & \new_[17370]_ ;
  assign \new_[17382]_  = A167 & A168;
  assign \new_[17383]_  = A169 & \new_[17382]_ ;
  assign \new_[17386]_  = ~A232 & ~A166;
  assign \new_[17389]_  = A234 & A233;
  assign \new_[17390]_  = \new_[17389]_  & \new_[17386]_ ;
  assign \new_[17391]_  = \new_[17390]_  & \new_[17383]_ ;
  assign \new_[17395]_  = A268 & ~A267;
  assign \new_[17396]_  = ~A236 & \new_[17395]_ ;
  assign \new_[17399]_  = A299 & ~A298;
  assign \new_[17402]_  = ~A302 & A300;
  assign \new_[17403]_  = \new_[17402]_  & \new_[17399]_ ;
  assign \new_[17404]_  = \new_[17403]_  & \new_[17396]_ ;
  assign \new_[17408]_  = A167 & A168;
  assign \new_[17409]_  = A169 & \new_[17408]_ ;
  assign \new_[17412]_  = ~A232 & ~A166;
  assign \new_[17415]_  = A234 & A233;
  assign \new_[17416]_  = \new_[17415]_  & \new_[17412]_ ;
  assign \new_[17417]_  = \new_[17416]_  & \new_[17409]_ ;
  assign \new_[17421]_  = ~A269 & ~A267;
  assign \new_[17422]_  = ~A236 & \new_[17421]_ ;
  assign \new_[17425]_  = ~A299 & A298;
  assign \new_[17428]_  = A301 & A300;
  assign \new_[17429]_  = \new_[17428]_  & \new_[17425]_ ;
  assign \new_[17430]_  = \new_[17429]_  & \new_[17422]_ ;
  assign \new_[17434]_  = A167 & A168;
  assign \new_[17435]_  = A169 & \new_[17434]_ ;
  assign \new_[17438]_  = ~A232 & ~A166;
  assign \new_[17441]_  = A234 & A233;
  assign \new_[17442]_  = \new_[17441]_  & \new_[17438]_ ;
  assign \new_[17443]_  = \new_[17442]_  & \new_[17435]_ ;
  assign \new_[17447]_  = ~A269 & ~A267;
  assign \new_[17448]_  = ~A236 & \new_[17447]_ ;
  assign \new_[17451]_  = ~A299 & A298;
  assign \new_[17454]_  = ~A302 & A300;
  assign \new_[17455]_  = \new_[17454]_  & \new_[17451]_ ;
  assign \new_[17456]_  = \new_[17455]_  & \new_[17448]_ ;
  assign \new_[17460]_  = A167 & A168;
  assign \new_[17461]_  = A169 & \new_[17460]_ ;
  assign \new_[17464]_  = ~A232 & ~A166;
  assign \new_[17467]_  = A234 & A233;
  assign \new_[17468]_  = \new_[17467]_  & \new_[17464]_ ;
  assign \new_[17469]_  = \new_[17468]_  & \new_[17461]_ ;
  assign \new_[17473]_  = ~A269 & ~A267;
  assign \new_[17474]_  = ~A236 & \new_[17473]_ ;
  assign \new_[17477]_  = A299 & ~A298;
  assign \new_[17480]_  = A301 & A300;
  assign \new_[17481]_  = \new_[17480]_  & \new_[17477]_ ;
  assign \new_[17482]_  = \new_[17481]_  & \new_[17474]_ ;
  assign \new_[17486]_  = A167 & A168;
  assign \new_[17487]_  = A169 & \new_[17486]_ ;
  assign \new_[17490]_  = ~A232 & ~A166;
  assign \new_[17493]_  = A234 & A233;
  assign \new_[17494]_  = \new_[17493]_  & \new_[17490]_ ;
  assign \new_[17495]_  = \new_[17494]_  & \new_[17487]_ ;
  assign \new_[17499]_  = ~A269 & ~A267;
  assign \new_[17500]_  = ~A236 & \new_[17499]_ ;
  assign \new_[17503]_  = A299 & ~A298;
  assign \new_[17506]_  = ~A302 & A300;
  assign \new_[17507]_  = \new_[17506]_  & \new_[17503]_ ;
  assign \new_[17508]_  = \new_[17507]_  & \new_[17500]_ ;
  assign \new_[17512]_  = A167 & A168;
  assign \new_[17513]_  = A169 & \new_[17512]_ ;
  assign \new_[17516]_  = ~A232 & ~A166;
  assign \new_[17519]_  = A234 & A233;
  assign \new_[17520]_  = \new_[17519]_  & \new_[17516]_ ;
  assign \new_[17521]_  = \new_[17520]_  & \new_[17513]_ ;
  assign \new_[17525]_  = A266 & A265;
  assign \new_[17526]_  = ~A236 & \new_[17525]_ ;
  assign \new_[17529]_  = ~A299 & A298;
  assign \new_[17532]_  = A301 & A300;
  assign \new_[17533]_  = \new_[17532]_  & \new_[17529]_ ;
  assign \new_[17534]_  = \new_[17533]_  & \new_[17526]_ ;
  assign \new_[17538]_  = A167 & A168;
  assign \new_[17539]_  = A169 & \new_[17538]_ ;
  assign \new_[17542]_  = ~A232 & ~A166;
  assign \new_[17545]_  = A234 & A233;
  assign \new_[17546]_  = \new_[17545]_  & \new_[17542]_ ;
  assign \new_[17547]_  = \new_[17546]_  & \new_[17539]_ ;
  assign \new_[17551]_  = A266 & A265;
  assign \new_[17552]_  = ~A236 & \new_[17551]_ ;
  assign \new_[17555]_  = ~A299 & A298;
  assign \new_[17558]_  = ~A302 & A300;
  assign \new_[17559]_  = \new_[17558]_  & \new_[17555]_ ;
  assign \new_[17560]_  = \new_[17559]_  & \new_[17552]_ ;
  assign \new_[17564]_  = A167 & A168;
  assign \new_[17565]_  = A169 & \new_[17564]_ ;
  assign \new_[17568]_  = ~A232 & ~A166;
  assign \new_[17571]_  = A234 & A233;
  assign \new_[17572]_  = \new_[17571]_  & \new_[17568]_ ;
  assign \new_[17573]_  = \new_[17572]_  & \new_[17565]_ ;
  assign \new_[17577]_  = A266 & A265;
  assign \new_[17578]_  = ~A236 & \new_[17577]_ ;
  assign \new_[17581]_  = A299 & ~A298;
  assign \new_[17584]_  = A301 & A300;
  assign \new_[17585]_  = \new_[17584]_  & \new_[17581]_ ;
  assign \new_[17586]_  = \new_[17585]_  & \new_[17578]_ ;
  assign \new_[17590]_  = A167 & A168;
  assign \new_[17591]_  = A169 & \new_[17590]_ ;
  assign \new_[17594]_  = ~A232 & ~A166;
  assign \new_[17597]_  = A234 & A233;
  assign \new_[17598]_  = \new_[17597]_  & \new_[17594]_ ;
  assign \new_[17599]_  = \new_[17598]_  & \new_[17591]_ ;
  assign \new_[17603]_  = A266 & A265;
  assign \new_[17604]_  = ~A236 & \new_[17603]_ ;
  assign \new_[17607]_  = A299 & ~A298;
  assign \new_[17610]_  = ~A302 & A300;
  assign \new_[17611]_  = \new_[17610]_  & \new_[17607]_ ;
  assign \new_[17612]_  = \new_[17611]_  & \new_[17604]_ ;
  assign \new_[17616]_  = A167 & A168;
  assign \new_[17617]_  = A169 & \new_[17616]_ ;
  assign \new_[17620]_  = ~A232 & ~A166;
  assign \new_[17623]_  = A234 & A233;
  assign \new_[17624]_  = \new_[17623]_  & \new_[17620]_ ;
  assign \new_[17625]_  = \new_[17624]_  & \new_[17617]_ ;
  assign \new_[17629]_  = ~A266 & ~A265;
  assign \new_[17630]_  = ~A236 & \new_[17629]_ ;
  assign \new_[17633]_  = ~A299 & A298;
  assign \new_[17636]_  = A301 & A300;
  assign \new_[17637]_  = \new_[17636]_  & \new_[17633]_ ;
  assign \new_[17638]_  = \new_[17637]_  & \new_[17630]_ ;
  assign \new_[17642]_  = A167 & A168;
  assign \new_[17643]_  = A169 & \new_[17642]_ ;
  assign \new_[17646]_  = ~A232 & ~A166;
  assign \new_[17649]_  = A234 & A233;
  assign \new_[17650]_  = \new_[17649]_  & \new_[17646]_ ;
  assign \new_[17651]_  = \new_[17650]_  & \new_[17643]_ ;
  assign \new_[17655]_  = ~A266 & ~A265;
  assign \new_[17656]_  = ~A236 & \new_[17655]_ ;
  assign \new_[17659]_  = ~A299 & A298;
  assign \new_[17662]_  = ~A302 & A300;
  assign \new_[17663]_  = \new_[17662]_  & \new_[17659]_ ;
  assign \new_[17664]_  = \new_[17663]_  & \new_[17656]_ ;
  assign \new_[17668]_  = A167 & A168;
  assign \new_[17669]_  = A169 & \new_[17668]_ ;
  assign \new_[17672]_  = ~A232 & ~A166;
  assign \new_[17675]_  = A234 & A233;
  assign \new_[17676]_  = \new_[17675]_  & \new_[17672]_ ;
  assign \new_[17677]_  = \new_[17676]_  & \new_[17669]_ ;
  assign \new_[17681]_  = ~A266 & ~A265;
  assign \new_[17682]_  = ~A236 & \new_[17681]_ ;
  assign \new_[17685]_  = A299 & ~A298;
  assign \new_[17688]_  = A301 & A300;
  assign \new_[17689]_  = \new_[17688]_  & \new_[17685]_ ;
  assign \new_[17690]_  = \new_[17689]_  & \new_[17682]_ ;
  assign \new_[17694]_  = A167 & A168;
  assign \new_[17695]_  = A169 & \new_[17694]_ ;
  assign \new_[17698]_  = ~A232 & ~A166;
  assign \new_[17701]_  = A234 & A233;
  assign \new_[17702]_  = \new_[17701]_  & \new_[17698]_ ;
  assign \new_[17703]_  = \new_[17702]_  & \new_[17695]_ ;
  assign \new_[17707]_  = ~A266 & ~A265;
  assign \new_[17708]_  = ~A236 & \new_[17707]_ ;
  assign \new_[17711]_  = A299 & ~A298;
  assign \new_[17714]_  = ~A302 & A300;
  assign \new_[17715]_  = \new_[17714]_  & \new_[17711]_ ;
  assign \new_[17716]_  = \new_[17715]_  & \new_[17708]_ ;
  assign \new_[17720]_  = A167 & A168;
  assign \new_[17721]_  = A169 & \new_[17720]_ ;
  assign \new_[17724]_  = A232 & ~A166;
  assign \new_[17727]_  = A234 & ~A233;
  assign \new_[17728]_  = \new_[17727]_  & \new_[17724]_ ;
  assign \new_[17729]_  = \new_[17728]_  & \new_[17721]_ ;
  assign \new_[17733]_  = A268 & ~A267;
  assign \new_[17734]_  = A235 & \new_[17733]_ ;
  assign \new_[17737]_  = ~A299 & A298;
  assign \new_[17740]_  = A301 & A300;
  assign \new_[17741]_  = \new_[17740]_  & \new_[17737]_ ;
  assign \new_[17742]_  = \new_[17741]_  & \new_[17734]_ ;
  assign \new_[17746]_  = A167 & A168;
  assign \new_[17747]_  = A169 & \new_[17746]_ ;
  assign \new_[17750]_  = A232 & ~A166;
  assign \new_[17753]_  = A234 & ~A233;
  assign \new_[17754]_  = \new_[17753]_  & \new_[17750]_ ;
  assign \new_[17755]_  = \new_[17754]_  & \new_[17747]_ ;
  assign \new_[17759]_  = A268 & ~A267;
  assign \new_[17760]_  = A235 & \new_[17759]_ ;
  assign \new_[17763]_  = ~A299 & A298;
  assign \new_[17766]_  = ~A302 & A300;
  assign \new_[17767]_  = \new_[17766]_  & \new_[17763]_ ;
  assign \new_[17768]_  = \new_[17767]_  & \new_[17760]_ ;
  assign \new_[17772]_  = A167 & A168;
  assign \new_[17773]_  = A169 & \new_[17772]_ ;
  assign \new_[17776]_  = A232 & ~A166;
  assign \new_[17779]_  = A234 & ~A233;
  assign \new_[17780]_  = \new_[17779]_  & \new_[17776]_ ;
  assign \new_[17781]_  = \new_[17780]_  & \new_[17773]_ ;
  assign \new_[17785]_  = A268 & ~A267;
  assign \new_[17786]_  = A235 & \new_[17785]_ ;
  assign \new_[17789]_  = A299 & ~A298;
  assign \new_[17792]_  = A301 & A300;
  assign \new_[17793]_  = \new_[17792]_  & \new_[17789]_ ;
  assign \new_[17794]_  = \new_[17793]_  & \new_[17786]_ ;
  assign \new_[17798]_  = A167 & A168;
  assign \new_[17799]_  = A169 & \new_[17798]_ ;
  assign \new_[17802]_  = A232 & ~A166;
  assign \new_[17805]_  = A234 & ~A233;
  assign \new_[17806]_  = \new_[17805]_  & \new_[17802]_ ;
  assign \new_[17807]_  = \new_[17806]_  & \new_[17799]_ ;
  assign \new_[17811]_  = A268 & ~A267;
  assign \new_[17812]_  = A235 & \new_[17811]_ ;
  assign \new_[17815]_  = A299 & ~A298;
  assign \new_[17818]_  = ~A302 & A300;
  assign \new_[17819]_  = \new_[17818]_  & \new_[17815]_ ;
  assign \new_[17820]_  = \new_[17819]_  & \new_[17812]_ ;
  assign \new_[17824]_  = A167 & A168;
  assign \new_[17825]_  = A169 & \new_[17824]_ ;
  assign \new_[17828]_  = A232 & ~A166;
  assign \new_[17831]_  = A234 & ~A233;
  assign \new_[17832]_  = \new_[17831]_  & \new_[17828]_ ;
  assign \new_[17833]_  = \new_[17832]_  & \new_[17825]_ ;
  assign \new_[17837]_  = ~A269 & ~A267;
  assign \new_[17838]_  = A235 & \new_[17837]_ ;
  assign \new_[17841]_  = ~A299 & A298;
  assign \new_[17844]_  = A301 & A300;
  assign \new_[17845]_  = \new_[17844]_  & \new_[17841]_ ;
  assign \new_[17846]_  = \new_[17845]_  & \new_[17838]_ ;
  assign \new_[17850]_  = A167 & A168;
  assign \new_[17851]_  = A169 & \new_[17850]_ ;
  assign \new_[17854]_  = A232 & ~A166;
  assign \new_[17857]_  = A234 & ~A233;
  assign \new_[17858]_  = \new_[17857]_  & \new_[17854]_ ;
  assign \new_[17859]_  = \new_[17858]_  & \new_[17851]_ ;
  assign \new_[17863]_  = ~A269 & ~A267;
  assign \new_[17864]_  = A235 & \new_[17863]_ ;
  assign \new_[17867]_  = ~A299 & A298;
  assign \new_[17870]_  = ~A302 & A300;
  assign \new_[17871]_  = \new_[17870]_  & \new_[17867]_ ;
  assign \new_[17872]_  = \new_[17871]_  & \new_[17864]_ ;
  assign \new_[17876]_  = A167 & A168;
  assign \new_[17877]_  = A169 & \new_[17876]_ ;
  assign \new_[17880]_  = A232 & ~A166;
  assign \new_[17883]_  = A234 & ~A233;
  assign \new_[17884]_  = \new_[17883]_  & \new_[17880]_ ;
  assign \new_[17885]_  = \new_[17884]_  & \new_[17877]_ ;
  assign \new_[17889]_  = ~A269 & ~A267;
  assign \new_[17890]_  = A235 & \new_[17889]_ ;
  assign \new_[17893]_  = A299 & ~A298;
  assign \new_[17896]_  = A301 & A300;
  assign \new_[17897]_  = \new_[17896]_  & \new_[17893]_ ;
  assign \new_[17898]_  = \new_[17897]_  & \new_[17890]_ ;
  assign \new_[17902]_  = A167 & A168;
  assign \new_[17903]_  = A169 & \new_[17902]_ ;
  assign \new_[17906]_  = A232 & ~A166;
  assign \new_[17909]_  = A234 & ~A233;
  assign \new_[17910]_  = \new_[17909]_  & \new_[17906]_ ;
  assign \new_[17911]_  = \new_[17910]_  & \new_[17903]_ ;
  assign \new_[17915]_  = ~A269 & ~A267;
  assign \new_[17916]_  = A235 & \new_[17915]_ ;
  assign \new_[17919]_  = A299 & ~A298;
  assign \new_[17922]_  = ~A302 & A300;
  assign \new_[17923]_  = \new_[17922]_  & \new_[17919]_ ;
  assign \new_[17924]_  = \new_[17923]_  & \new_[17916]_ ;
  assign \new_[17928]_  = A167 & A168;
  assign \new_[17929]_  = A169 & \new_[17928]_ ;
  assign \new_[17932]_  = A232 & ~A166;
  assign \new_[17935]_  = A234 & ~A233;
  assign \new_[17936]_  = \new_[17935]_  & \new_[17932]_ ;
  assign \new_[17937]_  = \new_[17936]_  & \new_[17929]_ ;
  assign \new_[17941]_  = A266 & A265;
  assign \new_[17942]_  = A235 & \new_[17941]_ ;
  assign \new_[17945]_  = ~A299 & A298;
  assign \new_[17948]_  = A301 & A300;
  assign \new_[17949]_  = \new_[17948]_  & \new_[17945]_ ;
  assign \new_[17950]_  = \new_[17949]_  & \new_[17942]_ ;
  assign \new_[17954]_  = A167 & A168;
  assign \new_[17955]_  = A169 & \new_[17954]_ ;
  assign \new_[17958]_  = A232 & ~A166;
  assign \new_[17961]_  = A234 & ~A233;
  assign \new_[17962]_  = \new_[17961]_  & \new_[17958]_ ;
  assign \new_[17963]_  = \new_[17962]_  & \new_[17955]_ ;
  assign \new_[17967]_  = A266 & A265;
  assign \new_[17968]_  = A235 & \new_[17967]_ ;
  assign \new_[17971]_  = ~A299 & A298;
  assign \new_[17974]_  = ~A302 & A300;
  assign \new_[17975]_  = \new_[17974]_  & \new_[17971]_ ;
  assign \new_[17976]_  = \new_[17975]_  & \new_[17968]_ ;
  assign \new_[17980]_  = A167 & A168;
  assign \new_[17981]_  = A169 & \new_[17980]_ ;
  assign \new_[17984]_  = A232 & ~A166;
  assign \new_[17987]_  = A234 & ~A233;
  assign \new_[17988]_  = \new_[17987]_  & \new_[17984]_ ;
  assign \new_[17989]_  = \new_[17988]_  & \new_[17981]_ ;
  assign \new_[17993]_  = A266 & A265;
  assign \new_[17994]_  = A235 & \new_[17993]_ ;
  assign \new_[17997]_  = A299 & ~A298;
  assign \new_[18000]_  = A301 & A300;
  assign \new_[18001]_  = \new_[18000]_  & \new_[17997]_ ;
  assign \new_[18002]_  = \new_[18001]_  & \new_[17994]_ ;
  assign \new_[18006]_  = A167 & A168;
  assign \new_[18007]_  = A169 & \new_[18006]_ ;
  assign \new_[18010]_  = A232 & ~A166;
  assign \new_[18013]_  = A234 & ~A233;
  assign \new_[18014]_  = \new_[18013]_  & \new_[18010]_ ;
  assign \new_[18015]_  = \new_[18014]_  & \new_[18007]_ ;
  assign \new_[18019]_  = A266 & A265;
  assign \new_[18020]_  = A235 & \new_[18019]_ ;
  assign \new_[18023]_  = A299 & ~A298;
  assign \new_[18026]_  = ~A302 & A300;
  assign \new_[18027]_  = \new_[18026]_  & \new_[18023]_ ;
  assign \new_[18028]_  = \new_[18027]_  & \new_[18020]_ ;
  assign \new_[18032]_  = A167 & A168;
  assign \new_[18033]_  = A169 & \new_[18032]_ ;
  assign \new_[18036]_  = A232 & ~A166;
  assign \new_[18039]_  = A234 & ~A233;
  assign \new_[18040]_  = \new_[18039]_  & \new_[18036]_ ;
  assign \new_[18041]_  = \new_[18040]_  & \new_[18033]_ ;
  assign \new_[18045]_  = ~A266 & ~A265;
  assign \new_[18046]_  = A235 & \new_[18045]_ ;
  assign \new_[18049]_  = ~A299 & A298;
  assign \new_[18052]_  = A301 & A300;
  assign \new_[18053]_  = \new_[18052]_  & \new_[18049]_ ;
  assign \new_[18054]_  = \new_[18053]_  & \new_[18046]_ ;
  assign \new_[18058]_  = A167 & A168;
  assign \new_[18059]_  = A169 & \new_[18058]_ ;
  assign \new_[18062]_  = A232 & ~A166;
  assign \new_[18065]_  = A234 & ~A233;
  assign \new_[18066]_  = \new_[18065]_  & \new_[18062]_ ;
  assign \new_[18067]_  = \new_[18066]_  & \new_[18059]_ ;
  assign \new_[18071]_  = ~A266 & ~A265;
  assign \new_[18072]_  = A235 & \new_[18071]_ ;
  assign \new_[18075]_  = ~A299 & A298;
  assign \new_[18078]_  = ~A302 & A300;
  assign \new_[18079]_  = \new_[18078]_  & \new_[18075]_ ;
  assign \new_[18080]_  = \new_[18079]_  & \new_[18072]_ ;
  assign \new_[18084]_  = A167 & A168;
  assign \new_[18085]_  = A169 & \new_[18084]_ ;
  assign \new_[18088]_  = A232 & ~A166;
  assign \new_[18091]_  = A234 & ~A233;
  assign \new_[18092]_  = \new_[18091]_  & \new_[18088]_ ;
  assign \new_[18093]_  = \new_[18092]_  & \new_[18085]_ ;
  assign \new_[18097]_  = ~A266 & ~A265;
  assign \new_[18098]_  = A235 & \new_[18097]_ ;
  assign \new_[18101]_  = A299 & ~A298;
  assign \new_[18104]_  = A301 & A300;
  assign \new_[18105]_  = \new_[18104]_  & \new_[18101]_ ;
  assign \new_[18106]_  = \new_[18105]_  & \new_[18098]_ ;
  assign \new_[18110]_  = A167 & A168;
  assign \new_[18111]_  = A169 & \new_[18110]_ ;
  assign \new_[18114]_  = A232 & ~A166;
  assign \new_[18117]_  = A234 & ~A233;
  assign \new_[18118]_  = \new_[18117]_  & \new_[18114]_ ;
  assign \new_[18119]_  = \new_[18118]_  & \new_[18111]_ ;
  assign \new_[18123]_  = ~A266 & ~A265;
  assign \new_[18124]_  = A235 & \new_[18123]_ ;
  assign \new_[18127]_  = A299 & ~A298;
  assign \new_[18130]_  = ~A302 & A300;
  assign \new_[18131]_  = \new_[18130]_  & \new_[18127]_ ;
  assign \new_[18132]_  = \new_[18131]_  & \new_[18124]_ ;
  assign \new_[18136]_  = A167 & A168;
  assign \new_[18137]_  = A169 & \new_[18136]_ ;
  assign \new_[18140]_  = A232 & ~A166;
  assign \new_[18143]_  = A234 & ~A233;
  assign \new_[18144]_  = \new_[18143]_  & \new_[18140]_ ;
  assign \new_[18145]_  = \new_[18144]_  & \new_[18137]_ ;
  assign \new_[18149]_  = A268 & ~A267;
  assign \new_[18150]_  = ~A236 & \new_[18149]_ ;
  assign \new_[18153]_  = ~A299 & A298;
  assign \new_[18156]_  = A301 & A300;
  assign \new_[18157]_  = \new_[18156]_  & \new_[18153]_ ;
  assign \new_[18158]_  = \new_[18157]_  & \new_[18150]_ ;
  assign \new_[18162]_  = A167 & A168;
  assign \new_[18163]_  = A169 & \new_[18162]_ ;
  assign \new_[18166]_  = A232 & ~A166;
  assign \new_[18169]_  = A234 & ~A233;
  assign \new_[18170]_  = \new_[18169]_  & \new_[18166]_ ;
  assign \new_[18171]_  = \new_[18170]_  & \new_[18163]_ ;
  assign \new_[18175]_  = A268 & ~A267;
  assign \new_[18176]_  = ~A236 & \new_[18175]_ ;
  assign \new_[18179]_  = ~A299 & A298;
  assign \new_[18182]_  = ~A302 & A300;
  assign \new_[18183]_  = \new_[18182]_  & \new_[18179]_ ;
  assign \new_[18184]_  = \new_[18183]_  & \new_[18176]_ ;
  assign \new_[18188]_  = A167 & A168;
  assign \new_[18189]_  = A169 & \new_[18188]_ ;
  assign \new_[18192]_  = A232 & ~A166;
  assign \new_[18195]_  = A234 & ~A233;
  assign \new_[18196]_  = \new_[18195]_  & \new_[18192]_ ;
  assign \new_[18197]_  = \new_[18196]_  & \new_[18189]_ ;
  assign \new_[18201]_  = A268 & ~A267;
  assign \new_[18202]_  = ~A236 & \new_[18201]_ ;
  assign \new_[18205]_  = A299 & ~A298;
  assign \new_[18208]_  = A301 & A300;
  assign \new_[18209]_  = \new_[18208]_  & \new_[18205]_ ;
  assign \new_[18210]_  = \new_[18209]_  & \new_[18202]_ ;
  assign \new_[18214]_  = A167 & A168;
  assign \new_[18215]_  = A169 & \new_[18214]_ ;
  assign \new_[18218]_  = A232 & ~A166;
  assign \new_[18221]_  = A234 & ~A233;
  assign \new_[18222]_  = \new_[18221]_  & \new_[18218]_ ;
  assign \new_[18223]_  = \new_[18222]_  & \new_[18215]_ ;
  assign \new_[18227]_  = A268 & ~A267;
  assign \new_[18228]_  = ~A236 & \new_[18227]_ ;
  assign \new_[18231]_  = A299 & ~A298;
  assign \new_[18234]_  = ~A302 & A300;
  assign \new_[18235]_  = \new_[18234]_  & \new_[18231]_ ;
  assign \new_[18236]_  = \new_[18235]_  & \new_[18228]_ ;
  assign \new_[18240]_  = A167 & A168;
  assign \new_[18241]_  = A169 & \new_[18240]_ ;
  assign \new_[18244]_  = A232 & ~A166;
  assign \new_[18247]_  = A234 & ~A233;
  assign \new_[18248]_  = \new_[18247]_  & \new_[18244]_ ;
  assign \new_[18249]_  = \new_[18248]_  & \new_[18241]_ ;
  assign \new_[18253]_  = ~A269 & ~A267;
  assign \new_[18254]_  = ~A236 & \new_[18253]_ ;
  assign \new_[18257]_  = ~A299 & A298;
  assign \new_[18260]_  = A301 & A300;
  assign \new_[18261]_  = \new_[18260]_  & \new_[18257]_ ;
  assign \new_[18262]_  = \new_[18261]_  & \new_[18254]_ ;
  assign \new_[18266]_  = A167 & A168;
  assign \new_[18267]_  = A169 & \new_[18266]_ ;
  assign \new_[18270]_  = A232 & ~A166;
  assign \new_[18273]_  = A234 & ~A233;
  assign \new_[18274]_  = \new_[18273]_  & \new_[18270]_ ;
  assign \new_[18275]_  = \new_[18274]_  & \new_[18267]_ ;
  assign \new_[18279]_  = ~A269 & ~A267;
  assign \new_[18280]_  = ~A236 & \new_[18279]_ ;
  assign \new_[18283]_  = ~A299 & A298;
  assign \new_[18286]_  = ~A302 & A300;
  assign \new_[18287]_  = \new_[18286]_  & \new_[18283]_ ;
  assign \new_[18288]_  = \new_[18287]_  & \new_[18280]_ ;
  assign \new_[18292]_  = A167 & A168;
  assign \new_[18293]_  = A169 & \new_[18292]_ ;
  assign \new_[18296]_  = A232 & ~A166;
  assign \new_[18299]_  = A234 & ~A233;
  assign \new_[18300]_  = \new_[18299]_  & \new_[18296]_ ;
  assign \new_[18301]_  = \new_[18300]_  & \new_[18293]_ ;
  assign \new_[18305]_  = ~A269 & ~A267;
  assign \new_[18306]_  = ~A236 & \new_[18305]_ ;
  assign \new_[18309]_  = A299 & ~A298;
  assign \new_[18312]_  = A301 & A300;
  assign \new_[18313]_  = \new_[18312]_  & \new_[18309]_ ;
  assign \new_[18314]_  = \new_[18313]_  & \new_[18306]_ ;
  assign \new_[18318]_  = A167 & A168;
  assign \new_[18319]_  = A169 & \new_[18318]_ ;
  assign \new_[18322]_  = A232 & ~A166;
  assign \new_[18325]_  = A234 & ~A233;
  assign \new_[18326]_  = \new_[18325]_  & \new_[18322]_ ;
  assign \new_[18327]_  = \new_[18326]_  & \new_[18319]_ ;
  assign \new_[18331]_  = ~A269 & ~A267;
  assign \new_[18332]_  = ~A236 & \new_[18331]_ ;
  assign \new_[18335]_  = A299 & ~A298;
  assign \new_[18338]_  = ~A302 & A300;
  assign \new_[18339]_  = \new_[18338]_  & \new_[18335]_ ;
  assign \new_[18340]_  = \new_[18339]_  & \new_[18332]_ ;
  assign \new_[18344]_  = A167 & A168;
  assign \new_[18345]_  = A169 & \new_[18344]_ ;
  assign \new_[18348]_  = A232 & ~A166;
  assign \new_[18351]_  = A234 & ~A233;
  assign \new_[18352]_  = \new_[18351]_  & \new_[18348]_ ;
  assign \new_[18353]_  = \new_[18352]_  & \new_[18345]_ ;
  assign \new_[18357]_  = A266 & A265;
  assign \new_[18358]_  = ~A236 & \new_[18357]_ ;
  assign \new_[18361]_  = ~A299 & A298;
  assign \new_[18364]_  = A301 & A300;
  assign \new_[18365]_  = \new_[18364]_  & \new_[18361]_ ;
  assign \new_[18366]_  = \new_[18365]_  & \new_[18358]_ ;
  assign \new_[18370]_  = A167 & A168;
  assign \new_[18371]_  = A169 & \new_[18370]_ ;
  assign \new_[18374]_  = A232 & ~A166;
  assign \new_[18377]_  = A234 & ~A233;
  assign \new_[18378]_  = \new_[18377]_  & \new_[18374]_ ;
  assign \new_[18379]_  = \new_[18378]_  & \new_[18371]_ ;
  assign \new_[18383]_  = A266 & A265;
  assign \new_[18384]_  = ~A236 & \new_[18383]_ ;
  assign \new_[18387]_  = ~A299 & A298;
  assign \new_[18390]_  = ~A302 & A300;
  assign \new_[18391]_  = \new_[18390]_  & \new_[18387]_ ;
  assign \new_[18392]_  = \new_[18391]_  & \new_[18384]_ ;
  assign \new_[18396]_  = A167 & A168;
  assign \new_[18397]_  = A169 & \new_[18396]_ ;
  assign \new_[18400]_  = A232 & ~A166;
  assign \new_[18403]_  = A234 & ~A233;
  assign \new_[18404]_  = \new_[18403]_  & \new_[18400]_ ;
  assign \new_[18405]_  = \new_[18404]_  & \new_[18397]_ ;
  assign \new_[18409]_  = A266 & A265;
  assign \new_[18410]_  = ~A236 & \new_[18409]_ ;
  assign \new_[18413]_  = A299 & ~A298;
  assign \new_[18416]_  = A301 & A300;
  assign \new_[18417]_  = \new_[18416]_  & \new_[18413]_ ;
  assign \new_[18418]_  = \new_[18417]_  & \new_[18410]_ ;
  assign \new_[18422]_  = A167 & A168;
  assign \new_[18423]_  = A169 & \new_[18422]_ ;
  assign \new_[18426]_  = A232 & ~A166;
  assign \new_[18429]_  = A234 & ~A233;
  assign \new_[18430]_  = \new_[18429]_  & \new_[18426]_ ;
  assign \new_[18431]_  = \new_[18430]_  & \new_[18423]_ ;
  assign \new_[18435]_  = A266 & A265;
  assign \new_[18436]_  = ~A236 & \new_[18435]_ ;
  assign \new_[18439]_  = A299 & ~A298;
  assign \new_[18442]_  = ~A302 & A300;
  assign \new_[18443]_  = \new_[18442]_  & \new_[18439]_ ;
  assign \new_[18444]_  = \new_[18443]_  & \new_[18436]_ ;
  assign \new_[18448]_  = A167 & A168;
  assign \new_[18449]_  = A169 & \new_[18448]_ ;
  assign \new_[18452]_  = A232 & ~A166;
  assign \new_[18455]_  = A234 & ~A233;
  assign \new_[18456]_  = \new_[18455]_  & \new_[18452]_ ;
  assign \new_[18457]_  = \new_[18456]_  & \new_[18449]_ ;
  assign \new_[18461]_  = ~A266 & ~A265;
  assign \new_[18462]_  = ~A236 & \new_[18461]_ ;
  assign \new_[18465]_  = ~A299 & A298;
  assign \new_[18468]_  = A301 & A300;
  assign \new_[18469]_  = \new_[18468]_  & \new_[18465]_ ;
  assign \new_[18470]_  = \new_[18469]_  & \new_[18462]_ ;
  assign \new_[18474]_  = A167 & A168;
  assign \new_[18475]_  = A169 & \new_[18474]_ ;
  assign \new_[18478]_  = A232 & ~A166;
  assign \new_[18481]_  = A234 & ~A233;
  assign \new_[18482]_  = \new_[18481]_  & \new_[18478]_ ;
  assign \new_[18483]_  = \new_[18482]_  & \new_[18475]_ ;
  assign \new_[18487]_  = ~A266 & ~A265;
  assign \new_[18488]_  = ~A236 & \new_[18487]_ ;
  assign \new_[18491]_  = ~A299 & A298;
  assign \new_[18494]_  = ~A302 & A300;
  assign \new_[18495]_  = \new_[18494]_  & \new_[18491]_ ;
  assign \new_[18496]_  = \new_[18495]_  & \new_[18488]_ ;
  assign \new_[18500]_  = A167 & A168;
  assign \new_[18501]_  = A169 & \new_[18500]_ ;
  assign \new_[18504]_  = A232 & ~A166;
  assign \new_[18507]_  = A234 & ~A233;
  assign \new_[18508]_  = \new_[18507]_  & \new_[18504]_ ;
  assign \new_[18509]_  = \new_[18508]_  & \new_[18501]_ ;
  assign \new_[18513]_  = ~A266 & ~A265;
  assign \new_[18514]_  = ~A236 & \new_[18513]_ ;
  assign \new_[18517]_  = A299 & ~A298;
  assign \new_[18520]_  = A301 & A300;
  assign \new_[18521]_  = \new_[18520]_  & \new_[18517]_ ;
  assign \new_[18522]_  = \new_[18521]_  & \new_[18514]_ ;
  assign \new_[18526]_  = A167 & A168;
  assign \new_[18527]_  = A169 & \new_[18526]_ ;
  assign \new_[18530]_  = A232 & ~A166;
  assign \new_[18533]_  = A234 & ~A233;
  assign \new_[18534]_  = \new_[18533]_  & \new_[18530]_ ;
  assign \new_[18535]_  = \new_[18534]_  & \new_[18527]_ ;
  assign \new_[18539]_  = ~A266 & ~A265;
  assign \new_[18540]_  = ~A236 & \new_[18539]_ ;
  assign \new_[18543]_  = A299 & ~A298;
  assign \new_[18546]_  = ~A302 & A300;
  assign \new_[18547]_  = \new_[18546]_  & \new_[18543]_ ;
  assign \new_[18548]_  = \new_[18547]_  & \new_[18540]_ ;
  assign \new_[18552]_  = ~A167 & A168;
  assign \new_[18553]_  = A169 & \new_[18552]_ ;
  assign \new_[18556]_  = ~A232 & A166;
  assign \new_[18559]_  = A234 & A233;
  assign \new_[18560]_  = \new_[18559]_  & \new_[18556]_ ;
  assign \new_[18561]_  = \new_[18560]_  & \new_[18553]_ ;
  assign \new_[18565]_  = A268 & ~A267;
  assign \new_[18566]_  = A235 & \new_[18565]_ ;
  assign \new_[18569]_  = ~A299 & A298;
  assign \new_[18572]_  = A301 & A300;
  assign \new_[18573]_  = \new_[18572]_  & \new_[18569]_ ;
  assign \new_[18574]_  = \new_[18573]_  & \new_[18566]_ ;
  assign \new_[18578]_  = ~A167 & A168;
  assign \new_[18579]_  = A169 & \new_[18578]_ ;
  assign \new_[18582]_  = ~A232 & A166;
  assign \new_[18585]_  = A234 & A233;
  assign \new_[18586]_  = \new_[18585]_  & \new_[18582]_ ;
  assign \new_[18587]_  = \new_[18586]_  & \new_[18579]_ ;
  assign \new_[18591]_  = A268 & ~A267;
  assign \new_[18592]_  = A235 & \new_[18591]_ ;
  assign \new_[18595]_  = ~A299 & A298;
  assign \new_[18598]_  = ~A302 & A300;
  assign \new_[18599]_  = \new_[18598]_  & \new_[18595]_ ;
  assign \new_[18600]_  = \new_[18599]_  & \new_[18592]_ ;
  assign \new_[18604]_  = ~A167 & A168;
  assign \new_[18605]_  = A169 & \new_[18604]_ ;
  assign \new_[18608]_  = ~A232 & A166;
  assign \new_[18611]_  = A234 & A233;
  assign \new_[18612]_  = \new_[18611]_  & \new_[18608]_ ;
  assign \new_[18613]_  = \new_[18612]_  & \new_[18605]_ ;
  assign \new_[18617]_  = A268 & ~A267;
  assign \new_[18618]_  = A235 & \new_[18617]_ ;
  assign \new_[18621]_  = A299 & ~A298;
  assign \new_[18624]_  = A301 & A300;
  assign \new_[18625]_  = \new_[18624]_  & \new_[18621]_ ;
  assign \new_[18626]_  = \new_[18625]_  & \new_[18618]_ ;
  assign \new_[18630]_  = ~A167 & A168;
  assign \new_[18631]_  = A169 & \new_[18630]_ ;
  assign \new_[18634]_  = ~A232 & A166;
  assign \new_[18637]_  = A234 & A233;
  assign \new_[18638]_  = \new_[18637]_  & \new_[18634]_ ;
  assign \new_[18639]_  = \new_[18638]_  & \new_[18631]_ ;
  assign \new_[18643]_  = A268 & ~A267;
  assign \new_[18644]_  = A235 & \new_[18643]_ ;
  assign \new_[18647]_  = A299 & ~A298;
  assign \new_[18650]_  = ~A302 & A300;
  assign \new_[18651]_  = \new_[18650]_  & \new_[18647]_ ;
  assign \new_[18652]_  = \new_[18651]_  & \new_[18644]_ ;
  assign \new_[18656]_  = ~A167 & A168;
  assign \new_[18657]_  = A169 & \new_[18656]_ ;
  assign \new_[18660]_  = ~A232 & A166;
  assign \new_[18663]_  = A234 & A233;
  assign \new_[18664]_  = \new_[18663]_  & \new_[18660]_ ;
  assign \new_[18665]_  = \new_[18664]_  & \new_[18657]_ ;
  assign \new_[18669]_  = ~A269 & ~A267;
  assign \new_[18670]_  = A235 & \new_[18669]_ ;
  assign \new_[18673]_  = ~A299 & A298;
  assign \new_[18676]_  = A301 & A300;
  assign \new_[18677]_  = \new_[18676]_  & \new_[18673]_ ;
  assign \new_[18678]_  = \new_[18677]_  & \new_[18670]_ ;
  assign \new_[18682]_  = ~A167 & A168;
  assign \new_[18683]_  = A169 & \new_[18682]_ ;
  assign \new_[18686]_  = ~A232 & A166;
  assign \new_[18689]_  = A234 & A233;
  assign \new_[18690]_  = \new_[18689]_  & \new_[18686]_ ;
  assign \new_[18691]_  = \new_[18690]_  & \new_[18683]_ ;
  assign \new_[18695]_  = ~A269 & ~A267;
  assign \new_[18696]_  = A235 & \new_[18695]_ ;
  assign \new_[18699]_  = ~A299 & A298;
  assign \new_[18702]_  = ~A302 & A300;
  assign \new_[18703]_  = \new_[18702]_  & \new_[18699]_ ;
  assign \new_[18704]_  = \new_[18703]_  & \new_[18696]_ ;
  assign \new_[18708]_  = ~A167 & A168;
  assign \new_[18709]_  = A169 & \new_[18708]_ ;
  assign \new_[18712]_  = ~A232 & A166;
  assign \new_[18715]_  = A234 & A233;
  assign \new_[18716]_  = \new_[18715]_  & \new_[18712]_ ;
  assign \new_[18717]_  = \new_[18716]_  & \new_[18709]_ ;
  assign \new_[18721]_  = ~A269 & ~A267;
  assign \new_[18722]_  = A235 & \new_[18721]_ ;
  assign \new_[18725]_  = A299 & ~A298;
  assign \new_[18728]_  = A301 & A300;
  assign \new_[18729]_  = \new_[18728]_  & \new_[18725]_ ;
  assign \new_[18730]_  = \new_[18729]_  & \new_[18722]_ ;
  assign \new_[18734]_  = ~A167 & A168;
  assign \new_[18735]_  = A169 & \new_[18734]_ ;
  assign \new_[18738]_  = ~A232 & A166;
  assign \new_[18741]_  = A234 & A233;
  assign \new_[18742]_  = \new_[18741]_  & \new_[18738]_ ;
  assign \new_[18743]_  = \new_[18742]_  & \new_[18735]_ ;
  assign \new_[18747]_  = ~A269 & ~A267;
  assign \new_[18748]_  = A235 & \new_[18747]_ ;
  assign \new_[18751]_  = A299 & ~A298;
  assign \new_[18754]_  = ~A302 & A300;
  assign \new_[18755]_  = \new_[18754]_  & \new_[18751]_ ;
  assign \new_[18756]_  = \new_[18755]_  & \new_[18748]_ ;
  assign \new_[18760]_  = ~A167 & A168;
  assign \new_[18761]_  = A169 & \new_[18760]_ ;
  assign \new_[18764]_  = ~A232 & A166;
  assign \new_[18767]_  = A234 & A233;
  assign \new_[18768]_  = \new_[18767]_  & \new_[18764]_ ;
  assign \new_[18769]_  = \new_[18768]_  & \new_[18761]_ ;
  assign \new_[18773]_  = A266 & A265;
  assign \new_[18774]_  = A235 & \new_[18773]_ ;
  assign \new_[18777]_  = ~A299 & A298;
  assign \new_[18780]_  = A301 & A300;
  assign \new_[18781]_  = \new_[18780]_  & \new_[18777]_ ;
  assign \new_[18782]_  = \new_[18781]_  & \new_[18774]_ ;
  assign \new_[18786]_  = ~A167 & A168;
  assign \new_[18787]_  = A169 & \new_[18786]_ ;
  assign \new_[18790]_  = ~A232 & A166;
  assign \new_[18793]_  = A234 & A233;
  assign \new_[18794]_  = \new_[18793]_  & \new_[18790]_ ;
  assign \new_[18795]_  = \new_[18794]_  & \new_[18787]_ ;
  assign \new_[18799]_  = A266 & A265;
  assign \new_[18800]_  = A235 & \new_[18799]_ ;
  assign \new_[18803]_  = ~A299 & A298;
  assign \new_[18806]_  = ~A302 & A300;
  assign \new_[18807]_  = \new_[18806]_  & \new_[18803]_ ;
  assign \new_[18808]_  = \new_[18807]_  & \new_[18800]_ ;
  assign \new_[18812]_  = ~A167 & A168;
  assign \new_[18813]_  = A169 & \new_[18812]_ ;
  assign \new_[18816]_  = ~A232 & A166;
  assign \new_[18819]_  = A234 & A233;
  assign \new_[18820]_  = \new_[18819]_  & \new_[18816]_ ;
  assign \new_[18821]_  = \new_[18820]_  & \new_[18813]_ ;
  assign \new_[18825]_  = A266 & A265;
  assign \new_[18826]_  = A235 & \new_[18825]_ ;
  assign \new_[18829]_  = A299 & ~A298;
  assign \new_[18832]_  = A301 & A300;
  assign \new_[18833]_  = \new_[18832]_  & \new_[18829]_ ;
  assign \new_[18834]_  = \new_[18833]_  & \new_[18826]_ ;
  assign \new_[18838]_  = ~A167 & A168;
  assign \new_[18839]_  = A169 & \new_[18838]_ ;
  assign \new_[18842]_  = ~A232 & A166;
  assign \new_[18845]_  = A234 & A233;
  assign \new_[18846]_  = \new_[18845]_  & \new_[18842]_ ;
  assign \new_[18847]_  = \new_[18846]_  & \new_[18839]_ ;
  assign \new_[18851]_  = A266 & A265;
  assign \new_[18852]_  = A235 & \new_[18851]_ ;
  assign \new_[18855]_  = A299 & ~A298;
  assign \new_[18858]_  = ~A302 & A300;
  assign \new_[18859]_  = \new_[18858]_  & \new_[18855]_ ;
  assign \new_[18860]_  = \new_[18859]_  & \new_[18852]_ ;
  assign \new_[18864]_  = ~A167 & A168;
  assign \new_[18865]_  = A169 & \new_[18864]_ ;
  assign \new_[18868]_  = ~A232 & A166;
  assign \new_[18871]_  = A234 & A233;
  assign \new_[18872]_  = \new_[18871]_  & \new_[18868]_ ;
  assign \new_[18873]_  = \new_[18872]_  & \new_[18865]_ ;
  assign \new_[18877]_  = ~A266 & ~A265;
  assign \new_[18878]_  = A235 & \new_[18877]_ ;
  assign \new_[18881]_  = ~A299 & A298;
  assign \new_[18884]_  = A301 & A300;
  assign \new_[18885]_  = \new_[18884]_  & \new_[18881]_ ;
  assign \new_[18886]_  = \new_[18885]_  & \new_[18878]_ ;
  assign \new_[18890]_  = ~A167 & A168;
  assign \new_[18891]_  = A169 & \new_[18890]_ ;
  assign \new_[18894]_  = ~A232 & A166;
  assign \new_[18897]_  = A234 & A233;
  assign \new_[18898]_  = \new_[18897]_  & \new_[18894]_ ;
  assign \new_[18899]_  = \new_[18898]_  & \new_[18891]_ ;
  assign \new_[18903]_  = ~A266 & ~A265;
  assign \new_[18904]_  = A235 & \new_[18903]_ ;
  assign \new_[18907]_  = ~A299 & A298;
  assign \new_[18910]_  = ~A302 & A300;
  assign \new_[18911]_  = \new_[18910]_  & \new_[18907]_ ;
  assign \new_[18912]_  = \new_[18911]_  & \new_[18904]_ ;
  assign \new_[18916]_  = ~A167 & A168;
  assign \new_[18917]_  = A169 & \new_[18916]_ ;
  assign \new_[18920]_  = ~A232 & A166;
  assign \new_[18923]_  = A234 & A233;
  assign \new_[18924]_  = \new_[18923]_  & \new_[18920]_ ;
  assign \new_[18925]_  = \new_[18924]_  & \new_[18917]_ ;
  assign \new_[18929]_  = ~A266 & ~A265;
  assign \new_[18930]_  = A235 & \new_[18929]_ ;
  assign \new_[18933]_  = A299 & ~A298;
  assign \new_[18936]_  = A301 & A300;
  assign \new_[18937]_  = \new_[18936]_  & \new_[18933]_ ;
  assign \new_[18938]_  = \new_[18937]_  & \new_[18930]_ ;
  assign \new_[18942]_  = ~A167 & A168;
  assign \new_[18943]_  = A169 & \new_[18942]_ ;
  assign \new_[18946]_  = ~A232 & A166;
  assign \new_[18949]_  = A234 & A233;
  assign \new_[18950]_  = \new_[18949]_  & \new_[18946]_ ;
  assign \new_[18951]_  = \new_[18950]_  & \new_[18943]_ ;
  assign \new_[18955]_  = ~A266 & ~A265;
  assign \new_[18956]_  = A235 & \new_[18955]_ ;
  assign \new_[18959]_  = A299 & ~A298;
  assign \new_[18962]_  = ~A302 & A300;
  assign \new_[18963]_  = \new_[18962]_  & \new_[18959]_ ;
  assign \new_[18964]_  = \new_[18963]_  & \new_[18956]_ ;
  assign \new_[18968]_  = ~A167 & A168;
  assign \new_[18969]_  = A169 & \new_[18968]_ ;
  assign \new_[18972]_  = ~A232 & A166;
  assign \new_[18975]_  = A234 & A233;
  assign \new_[18976]_  = \new_[18975]_  & \new_[18972]_ ;
  assign \new_[18977]_  = \new_[18976]_  & \new_[18969]_ ;
  assign \new_[18981]_  = A268 & ~A267;
  assign \new_[18982]_  = ~A236 & \new_[18981]_ ;
  assign \new_[18985]_  = ~A299 & A298;
  assign \new_[18988]_  = A301 & A300;
  assign \new_[18989]_  = \new_[18988]_  & \new_[18985]_ ;
  assign \new_[18990]_  = \new_[18989]_  & \new_[18982]_ ;
  assign \new_[18994]_  = ~A167 & A168;
  assign \new_[18995]_  = A169 & \new_[18994]_ ;
  assign \new_[18998]_  = ~A232 & A166;
  assign \new_[19001]_  = A234 & A233;
  assign \new_[19002]_  = \new_[19001]_  & \new_[18998]_ ;
  assign \new_[19003]_  = \new_[19002]_  & \new_[18995]_ ;
  assign \new_[19007]_  = A268 & ~A267;
  assign \new_[19008]_  = ~A236 & \new_[19007]_ ;
  assign \new_[19011]_  = ~A299 & A298;
  assign \new_[19014]_  = ~A302 & A300;
  assign \new_[19015]_  = \new_[19014]_  & \new_[19011]_ ;
  assign \new_[19016]_  = \new_[19015]_  & \new_[19008]_ ;
  assign \new_[19020]_  = ~A167 & A168;
  assign \new_[19021]_  = A169 & \new_[19020]_ ;
  assign \new_[19024]_  = ~A232 & A166;
  assign \new_[19027]_  = A234 & A233;
  assign \new_[19028]_  = \new_[19027]_  & \new_[19024]_ ;
  assign \new_[19029]_  = \new_[19028]_  & \new_[19021]_ ;
  assign \new_[19033]_  = A268 & ~A267;
  assign \new_[19034]_  = ~A236 & \new_[19033]_ ;
  assign \new_[19037]_  = A299 & ~A298;
  assign \new_[19040]_  = A301 & A300;
  assign \new_[19041]_  = \new_[19040]_  & \new_[19037]_ ;
  assign \new_[19042]_  = \new_[19041]_  & \new_[19034]_ ;
  assign \new_[19046]_  = ~A167 & A168;
  assign \new_[19047]_  = A169 & \new_[19046]_ ;
  assign \new_[19050]_  = ~A232 & A166;
  assign \new_[19053]_  = A234 & A233;
  assign \new_[19054]_  = \new_[19053]_  & \new_[19050]_ ;
  assign \new_[19055]_  = \new_[19054]_  & \new_[19047]_ ;
  assign \new_[19059]_  = A268 & ~A267;
  assign \new_[19060]_  = ~A236 & \new_[19059]_ ;
  assign \new_[19063]_  = A299 & ~A298;
  assign \new_[19066]_  = ~A302 & A300;
  assign \new_[19067]_  = \new_[19066]_  & \new_[19063]_ ;
  assign \new_[19068]_  = \new_[19067]_  & \new_[19060]_ ;
  assign \new_[19072]_  = ~A167 & A168;
  assign \new_[19073]_  = A169 & \new_[19072]_ ;
  assign \new_[19076]_  = ~A232 & A166;
  assign \new_[19079]_  = A234 & A233;
  assign \new_[19080]_  = \new_[19079]_  & \new_[19076]_ ;
  assign \new_[19081]_  = \new_[19080]_  & \new_[19073]_ ;
  assign \new_[19085]_  = ~A269 & ~A267;
  assign \new_[19086]_  = ~A236 & \new_[19085]_ ;
  assign \new_[19089]_  = ~A299 & A298;
  assign \new_[19092]_  = A301 & A300;
  assign \new_[19093]_  = \new_[19092]_  & \new_[19089]_ ;
  assign \new_[19094]_  = \new_[19093]_  & \new_[19086]_ ;
  assign \new_[19098]_  = ~A167 & A168;
  assign \new_[19099]_  = A169 & \new_[19098]_ ;
  assign \new_[19102]_  = ~A232 & A166;
  assign \new_[19105]_  = A234 & A233;
  assign \new_[19106]_  = \new_[19105]_  & \new_[19102]_ ;
  assign \new_[19107]_  = \new_[19106]_  & \new_[19099]_ ;
  assign \new_[19111]_  = ~A269 & ~A267;
  assign \new_[19112]_  = ~A236 & \new_[19111]_ ;
  assign \new_[19115]_  = ~A299 & A298;
  assign \new_[19118]_  = ~A302 & A300;
  assign \new_[19119]_  = \new_[19118]_  & \new_[19115]_ ;
  assign \new_[19120]_  = \new_[19119]_  & \new_[19112]_ ;
  assign \new_[19124]_  = ~A167 & A168;
  assign \new_[19125]_  = A169 & \new_[19124]_ ;
  assign \new_[19128]_  = ~A232 & A166;
  assign \new_[19131]_  = A234 & A233;
  assign \new_[19132]_  = \new_[19131]_  & \new_[19128]_ ;
  assign \new_[19133]_  = \new_[19132]_  & \new_[19125]_ ;
  assign \new_[19137]_  = ~A269 & ~A267;
  assign \new_[19138]_  = ~A236 & \new_[19137]_ ;
  assign \new_[19141]_  = A299 & ~A298;
  assign \new_[19144]_  = A301 & A300;
  assign \new_[19145]_  = \new_[19144]_  & \new_[19141]_ ;
  assign \new_[19146]_  = \new_[19145]_  & \new_[19138]_ ;
  assign \new_[19150]_  = ~A167 & A168;
  assign \new_[19151]_  = A169 & \new_[19150]_ ;
  assign \new_[19154]_  = ~A232 & A166;
  assign \new_[19157]_  = A234 & A233;
  assign \new_[19158]_  = \new_[19157]_  & \new_[19154]_ ;
  assign \new_[19159]_  = \new_[19158]_  & \new_[19151]_ ;
  assign \new_[19163]_  = ~A269 & ~A267;
  assign \new_[19164]_  = ~A236 & \new_[19163]_ ;
  assign \new_[19167]_  = A299 & ~A298;
  assign \new_[19170]_  = ~A302 & A300;
  assign \new_[19171]_  = \new_[19170]_  & \new_[19167]_ ;
  assign \new_[19172]_  = \new_[19171]_  & \new_[19164]_ ;
  assign \new_[19176]_  = ~A167 & A168;
  assign \new_[19177]_  = A169 & \new_[19176]_ ;
  assign \new_[19180]_  = ~A232 & A166;
  assign \new_[19183]_  = A234 & A233;
  assign \new_[19184]_  = \new_[19183]_  & \new_[19180]_ ;
  assign \new_[19185]_  = \new_[19184]_  & \new_[19177]_ ;
  assign \new_[19189]_  = A266 & A265;
  assign \new_[19190]_  = ~A236 & \new_[19189]_ ;
  assign \new_[19193]_  = ~A299 & A298;
  assign \new_[19196]_  = A301 & A300;
  assign \new_[19197]_  = \new_[19196]_  & \new_[19193]_ ;
  assign \new_[19198]_  = \new_[19197]_  & \new_[19190]_ ;
  assign \new_[19202]_  = ~A167 & A168;
  assign \new_[19203]_  = A169 & \new_[19202]_ ;
  assign \new_[19206]_  = ~A232 & A166;
  assign \new_[19209]_  = A234 & A233;
  assign \new_[19210]_  = \new_[19209]_  & \new_[19206]_ ;
  assign \new_[19211]_  = \new_[19210]_  & \new_[19203]_ ;
  assign \new_[19215]_  = A266 & A265;
  assign \new_[19216]_  = ~A236 & \new_[19215]_ ;
  assign \new_[19219]_  = ~A299 & A298;
  assign \new_[19222]_  = ~A302 & A300;
  assign \new_[19223]_  = \new_[19222]_  & \new_[19219]_ ;
  assign \new_[19224]_  = \new_[19223]_  & \new_[19216]_ ;
  assign \new_[19228]_  = ~A167 & A168;
  assign \new_[19229]_  = A169 & \new_[19228]_ ;
  assign \new_[19232]_  = ~A232 & A166;
  assign \new_[19235]_  = A234 & A233;
  assign \new_[19236]_  = \new_[19235]_  & \new_[19232]_ ;
  assign \new_[19237]_  = \new_[19236]_  & \new_[19229]_ ;
  assign \new_[19241]_  = A266 & A265;
  assign \new_[19242]_  = ~A236 & \new_[19241]_ ;
  assign \new_[19245]_  = A299 & ~A298;
  assign \new_[19248]_  = A301 & A300;
  assign \new_[19249]_  = \new_[19248]_  & \new_[19245]_ ;
  assign \new_[19250]_  = \new_[19249]_  & \new_[19242]_ ;
  assign \new_[19254]_  = ~A167 & A168;
  assign \new_[19255]_  = A169 & \new_[19254]_ ;
  assign \new_[19258]_  = ~A232 & A166;
  assign \new_[19261]_  = A234 & A233;
  assign \new_[19262]_  = \new_[19261]_  & \new_[19258]_ ;
  assign \new_[19263]_  = \new_[19262]_  & \new_[19255]_ ;
  assign \new_[19267]_  = A266 & A265;
  assign \new_[19268]_  = ~A236 & \new_[19267]_ ;
  assign \new_[19271]_  = A299 & ~A298;
  assign \new_[19274]_  = ~A302 & A300;
  assign \new_[19275]_  = \new_[19274]_  & \new_[19271]_ ;
  assign \new_[19276]_  = \new_[19275]_  & \new_[19268]_ ;
  assign \new_[19280]_  = ~A167 & A168;
  assign \new_[19281]_  = A169 & \new_[19280]_ ;
  assign \new_[19284]_  = ~A232 & A166;
  assign \new_[19287]_  = A234 & A233;
  assign \new_[19288]_  = \new_[19287]_  & \new_[19284]_ ;
  assign \new_[19289]_  = \new_[19288]_  & \new_[19281]_ ;
  assign \new_[19293]_  = ~A266 & ~A265;
  assign \new_[19294]_  = ~A236 & \new_[19293]_ ;
  assign \new_[19297]_  = ~A299 & A298;
  assign \new_[19300]_  = A301 & A300;
  assign \new_[19301]_  = \new_[19300]_  & \new_[19297]_ ;
  assign \new_[19302]_  = \new_[19301]_  & \new_[19294]_ ;
  assign \new_[19306]_  = ~A167 & A168;
  assign \new_[19307]_  = A169 & \new_[19306]_ ;
  assign \new_[19310]_  = ~A232 & A166;
  assign \new_[19313]_  = A234 & A233;
  assign \new_[19314]_  = \new_[19313]_  & \new_[19310]_ ;
  assign \new_[19315]_  = \new_[19314]_  & \new_[19307]_ ;
  assign \new_[19319]_  = ~A266 & ~A265;
  assign \new_[19320]_  = ~A236 & \new_[19319]_ ;
  assign \new_[19323]_  = ~A299 & A298;
  assign \new_[19326]_  = ~A302 & A300;
  assign \new_[19327]_  = \new_[19326]_  & \new_[19323]_ ;
  assign \new_[19328]_  = \new_[19327]_  & \new_[19320]_ ;
  assign \new_[19332]_  = ~A167 & A168;
  assign \new_[19333]_  = A169 & \new_[19332]_ ;
  assign \new_[19336]_  = ~A232 & A166;
  assign \new_[19339]_  = A234 & A233;
  assign \new_[19340]_  = \new_[19339]_  & \new_[19336]_ ;
  assign \new_[19341]_  = \new_[19340]_  & \new_[19333]_ ;
  assign \new_[19345]_  = ~A266 & ~A265;
  assign \new_[19346]_  = ~A236 & \new_[19345]_ ;
  assign \new_[19349]_  = A299 & ~A298;
  assign \new_[19352]_  = A301 & A300;
  assign \new_[19353]_  = \new_[19352]_  & \new_[19349]_ ;
  assign \new_[19354]_  = \new_[19353]_  & \new_[19346]_ ;
  assign \new_[19358]_  = ~A167 & A168;
  assign \new_[19359]_  = A169 & \new_[19358]_ ;
  assign \new_[19362]_  = ~A232 & A166;
  assign \new_[19365]_  = A234 & A233;
  assign \new_[19366]_  = \new_[19365]_  & \new_[19362]_ ;
  assign \new_[19367]_  = \new_[19366]_  & \new_[19359]_ ;
  assign \new_[19371]_  = ~A266 & ~A265;
  assign \new_[19372]_  = ~A236 & \new_[19371]_ ;
  assign \new_[19375]_  = A299 & ~A298;
  assign \new_[19378]_  = ~A302 & A300;
  assign \new_[19379]_  = \new_[19378]_  & \new_[19375]_ ;
  assign \new_[19380]_  = \new_[19379]_  & \new_[19372]_ ;
  assign \new_[19384]_  = ~A167 & A168;
  assign \new_[19385]_  = A169 & \new_[19384]_ ;
  assign \new_[19388]_  = A232 & A166;
  assign \new_[19391]_  = A234 & ~A233;
  assign \new_[19392]_  = \new_[19391]_  & \new_[19388]_ ;
  assign \new_[19393]_  = \new_[19392]_  & \new_[19385]_ ;
  assign \new_[19397]_  = A268 & ~A267;
  assign \new_[19398]_  = A235 & \new_[19397]_ ;
  assign \new_[19401]_  = ~A299 & A298;
  assign \new_[19404]_  = A301 & A300;
  assign \new_[19405]_  = \new_[19404]_  & \new_[19401]_ ;
  assign \new_[19406]_  = \new_[19405]_  & \new_[19398]_ ;
  assign \new_[19410]_  = ~A167 & A168;
  assign \new_[19411]_  = A169 & \new_[19410]_ ;
  assign \new_[19414]_  = A232 & A166;
  assign \new_[19417]_  = A234 & ~A233;
  assign \new_[19418]_  = \new_[19417]_  & \new_[19414]_ ;
  assign \new_[19419]_  = \new_[19418]_  & \new_[19411]_ ;
  assign \new_[19423]_  = A268 & ~A267;
  assign \new_[19424]_  = A235 & \new_[19423]_ ;
  assign \new_[19427]_  = ~A299 & A298;
  assign \new_[19430]_  = ~A302 & A300;
  assign \new_[19431]_  = \new_[19430]_  & \new_[19427]_ ;
  assign \new_[19432]_  = \new_[19431]_  & \new_[19424]_ ;
  assign \new_[19436]_  = ~A167 & A168;
  assign \new_[19437]_  = A169 & \new_[19436]_ ;
  assign \new_[19440]_  = A232 & A166;
  assign \new_[19443]_  = A234 & ~A233;
  assign \new_[19444]_  = \new_[19443]_  & \new_[19440]_ ;
  assign \new_[19445]_  = \new_[19444]_  & \new_[19437]_ ;
  assign \new_[19449]_  = A268 & ~A267;
  assign \new_[19450]_  = A235 & \new_[19449]_ ;
  assign \new_[19453]_  = A299 & ~A298;
  assign \new_[19456]_  = A301 & A300;
  assign \new_[19457]_  = \new_[19456]_  & \new_[19453]_ ;
  assign \new_[19458]_  = \new_[19457]_  & \new_[19450]_ ;
  assign \new_[19462]_  = ~A167 & A168;
  assign \new_[19463]_  = A169 & \new_[19462]_ ;
  assign \new_[19466]_  = A232 & A166;
  assign \new_[19469]_  = A234 & ~A233;
  assign \new_[19470]_  = \new_[19469]_  & \new_[19466]_ ;
  assign \new_[19471]_  = \new_[19470]_  & \new_[19463]_ ;
  assign \new_[19475]_  = A268 & ~A267;
  assign \new_[19476]_  = A235 & \new_[19475]_ ;
  assign \new_[19479]_  = A299 & ~A298;
  assign \new_[19482]_  = ~A302 & A300;
  assign \new_[19483]_  = \new_[19482]_  & \new_[19479]_ ;
  assign \new_[19484]_  = \new_[19483]_  & \new_[19476]_ ;
  assign \new_[19488]_  = ~A167 & A168;
  assign \new_[19489]_  = A169 & \new_[19488]_ ;
  assign \new_[19492]_  = A232 & A166;
  assign \new_[19495]_  = A234 & ~A233;
  assign \new_[19496]_  = \new_[19495]_  & \new_[19492]_ ;
  assign \new_[19497]_  = \new_[19496]_  & \new_[19489]_ ;
  assign \new_[19501]_  = ~A269 & ~A267;
  assign \new_[19502]_  = A235 & \new_[19501]_ ;
  assign \new_[19505]_  = ~A299 & A298;
  assign \new_[19508]_  = A301 & A300;
  assign \new_[19509]_  = \new_[19508]_  & \new_[19505]_ ;
  assign \new_[19510]_  = \new_[19509]_  & \new_[19502]_ ;
  assign \new_[19514]_  = ~A167 & A168;
  assign \new_[19515]_  = A169 & \new_[19514]_ ;
  assign \new_[19518]_  = A232 & A166;
  assign \new_[19521]_  = A234 & ~A233;
  assign \new_[19522]_  = \new_[19521]_  & \new_[19518]_ ;
  assign \new_[19523]_  = \new_[19522]_  & \new_[19515]_ ;
  assign \new_[19527]_  = ~A269 & ~A267;
  assign \new_[19528]_  = A235 & \new_[19527]_ ;
  assign \new_[19531]_  = ~A299 & A298;
  assign \new_[19534]_  = ~A302 & A300;
  assign \new_[19535]_  = \new_[19534]_  & \new_[19531]_ ;
  assign \new_[19536]_  = \new_[19535]_  & \new_[19528]_ ;
  assign \new_[19540]_  = ~A167 & A168;
  assign \new_[19541]_  = A169 & \new_[19540]_ ;
  assign \new_[19544]_  = A232 & A166;
  assign \new_[19547]_  = A234 & ~A233;
  assign \new_[19548]_  = \new_[19547]_  & \new_[19544]_ ;
  assign \new_[19549]_  = \new_[19548]_  & \new_[19541]_ ;
  assign \new_[19553]_  = ~A269 & ~A267;
  assign \new_[19554]_  = A235 & \new_[19553]_ ;
  assign \new_[19557]_  = A299 & ~A298;
  assign \new_[19560]_  = A301 & A300;
  assign \new_[19561]_  = \new_[19560]_  & \new_[19557]_ ;
  assign \new_[19562]_  = \new_[19561]_  & \new_[19554]_ ;
  assign \new_[19566]_  = ~A167 & A168;
  assign \new_[19567]_  = A169 & \new_[19566]_ ;
  assign \new_[19570]_  = A232 & A166;
  assign \new_[19573]_  = A234 & ~A233;
  assign \new_[19574]_  = \new_[19573]_  & \new_[19570]_ ;
  assign \new_[19575]_  = \new_[19574]_  & \new_[19567]_ ;
  assign \new_[19579]_  = ~A269 & ~A267;
  assign \new_[19580]_  = A235 & \new_[19579]_ ;
  assign \new_[19583]_  = A299 & ~A298;
  assign \new_[19586]_  = ~A302 & A300;
  assign \new_[19587]_  = \new_[19586]_  & \new_[19583]_ ;
  assign \new_[19588]_  = \new_[19587]_  & \new_[19580]_ ;
  assign \new_[19592]_  = ~A167 & A168;
  assign \new_[19593]_  = A169 & \new_[19592]_ ;
  assign \new_[19596]_  = A232 & A166;
  assign \new_[19599]_  = A234 & ~A233;
  assign \new_[19600]_  = \new_[19599]_  & \new_[19596]_ ;
  assign \new_[19601]_  = \new_[19600]_  & \new_[19593]_ ;
  assign \new_[19605]_  = A266 & A265;
  assign \new_[19606]_  = A235 & \new_[19605]_ ;
  assign \new_[19609]_  = ~A299 & A298;
  assign \new_[19612]_  = A301 & A300;
  assign \new_[19613]_  = \new_[19612]_  & \new_[19609]_ ;
  assign \new_[19614]_  = \new_[19613]_  & \new_[19606]_ ;
  assign \new_[19618]_  = ~A167 & A168;
  assign \new_[19619]_  = A169 & \new_[19618]_ ;
  assign \new_[19622]_  = A232 & A166;
  assign \new_[19625]_  = A234 & ~A233;
  assign \new_[19626]_  = \new_[19625]_  & \new_[19622]_ ;
  assign \new_[19627]_  = \new_[19626]_  & \new_[19619]_ ;
  assign \new_[19631]_  = A266 & A265;
  assign \new_[19632]_  = A235 & \new_[19631]_ ;
  assign \new_[19635]_  = ~A299 & A298;
  assign \new_[19638]_  = ~A302 & A300;
  assign \new_[19639]_  = \new_[19638]_  & \new_[19635]_ ;
  assign \new_[19640]_  = \new_[19639]_  & \new_[19632]_ ;
  assign \new_[19644]_  = ~A167 & A168;
  assign \new_[19645]_  = A169 & \new_[19644]_ ;
  assign \new_[19648]_  = A232 & A166;
  assign \new_[19651]_  = A234 & ~A233;
  assign \new_[19652]_  = \new_[19651]_  & \new_[19648]_ ;
  assign \new_[19653]_  = \new_[19652]_  & \new_[19645]_ ;
  assign \new_[19657]_  = A266 & A265;
  assign \new_[19658]_  = A235 & \new_[19657]_ ;
  assign \new_[19661]_  = A299 & ~A298;
  assign \new_[19664]_  = A301 & A300;
  assign \new_[19665]_  = \new_[19664]_  & \new_[19661]_ ;
  assign \new_[19666]_  = \new_[19665]_  & \new_[19658]_ ;
  assign \new_[19670]_  = ~A167 & A168;
  assign \new_[19671]_  = A169 & \new_[19670]_ ;
  assign \new_[19674]_  = A232 & A166;
  assign \new_[19677]_  = A234 & ~A233;
  assign \new_[19678]_  = \new_[19677]_  & \new_[19674]_ ;
  assign \new_[19679]_  = \new_[19678]_  & \new_[19671]_ ;
  assign \new_[19683]_  = A266 & A265;
  assign \new_[19684]_  = A235 & \new_[19683]_ ;
  assign \new_[19687]_  = A299 & ~A298;
  assign \new_[19690]_  = ~A302 & A300;
  assign \new_[19691]_  = \new_[19690]_  & \new_[19687]_ ;
  assign \new_[19692]_  = \new_[19691]_  & \new_[19684]_ ;
  assign \new_[19696]_  = ~A167 & A168;
  assign \new_[19697]_  = A169 & \new_[19696]_ ;
  assign \new_[19700]_  = A232 & A166;
  assign \new_[19703]_  = A234 & ~A233;
  assign \new_[19704]_  = \new_[19703]_  & \new_[19700]_ ;
  assign \new_[19705]_  = \new_[19704]_  & \new_[19697]_ ;
  assign \new_[19709]_  = ~A266 & ~A265;
  assign \new_[19710]_  = A235 & \new_[19709]_ ;
  assign \new_[19713]_  = ~A299 & A298;
  assign \new_[19716]_  = A301 & A300;
  assign \new_[19717]_  = \new_[19716]_  & \new_[19713]_ ;
  assign \new_[19718]_  = \new_[19717]_  & \new_[19710]_ ;
  assign \new_[19722]_  = ~A167 & A168;
  assign \new_[19723]_  = A169 & \new_[19722]_ ;
  assign \new_[19726]_  = A232 & A166;
  assign \new_[19729]_  = A234 & ~A233;
  assign \new_[19730]_  = \new_[19729]_  & \new_[19726]_ ;
  assign \new_[19731]_  = \new_[19730]_  & \new_[19723]_ ;
  assign \new_[19735]_  = ~A266 & ~A265;
  assign \new_[19736]_  = A235 & \new_[19735]_ ;
  assign \new_[19739]_  = ~A299 & A298;
  assign \new_[19742]_  = ~A302 & A300;
  assign \new_[19743]_  = \new_[19742]_  & \new_[19739]_ ;
  assign \new_[19744]_  = \new_[19743]_  & \new_[19736]_ ;
  assign \new_[19748]_  = ~A167 & A168;
  assign \new_[19749]_  = A169 & \new_[19748]_ ;
  assign \new_[19752]_  = A232 & A166;
  assign \new_[19755]_  = A234 & ~A233;
  assign \new_[19756]_  = \new_[19755]_  & \new_[19752]_ ;
  assign \new_[19757]_  = \new_[19756]_  & \new_[19749]_ ;
  assign \new_[19761]_  = ~A266 & ~A265;
  assign \new_[19762]_  = A235 & \new_[19761]_ ;
  assign \new_[19765]_  = A299 & ~A298;
  assign \new_[19768]_  = A301 & A300;
  assign \new_[19769]_  = \new_[19768]_  & \new_[19765]_ ;
  assign \new_[19770]_  = \new_[19769]_  & \new_[19762]_ ;
  assign \new_[19774]_  = ~A167 & A168;
  assign \new_[19775]_  = A169 & \new_[19774]_ ;
  assign \new_[19778]_  = A232 & A166;
  assign \new_[19781]_  = A234 & ~A233;
  assign \new_[19782]_  = \new_[19781]_  & \new_[19778]_ ;
  assign \new_[19783]_  = \new_[19782]_  & \new_[19775]_ ;
  assign \new_[19787]_  = ~A266 & ~A265;
  assign \new_[19788]_  = A235 & \new_[19787]_ ;
  assign \new_[19791]_  = A299 & ~A298;
  assign \new_[19794]_  = ~A302 & A300;
  assign \new_[19795]_  = \new_[19794]_  & \new_[19791]_ ;
  assign \new_[19796]_  = \new_[19795]_  & \new_[19788]_ ;
  assign \new_[19800]_  = ~A167 & A168;
  assign \new_[19801]_  = A169 & \new_[19800]_ ;
  assign \new_[19804]_  = A232 & A166;
  assign \new_[19807]_  = A234 & ~A233;
  assign \new_[19808]_  = \new_[19807]_  & \new_[19804]_ ;
  assign \new_[19809]_  = \new_[19808]_  & \new_[19801]_ ;
  assign \new_[19813]_  = A268 & ~A267;
  assign \new_[19814]_  = ~A236 & \new_[19813]_ ;
  assign \new_[19817]_  = ~A299 & A298;
  assign \new_[19820]_  = A301 & A300;
  assign \new_[19821]_  = \new_[19820]_  & \new_[19817]_ ;
  assign \new_[19822]_  = \new_[19821]_  & \new_[19814]_ ;
  assign \new_[19826]_  = ~A167 & A168;
  assign \new_[19827]_  = A169 & \new_[19826]_ ;
  assign \new_[19830]_  = A232 & A166;
  assign \new_[19833]_  = A234 & ~A233;
  assign \new_[19834]_  = \new_[19833]_  & \new_[19830]_ ;
  assign \new_[19835]_  = \new_[19834]_  & \new_[19827]_ ;
  assign \new_[19839]_  = A268 & ~A267;
  assign \new_[19840]_  = ~A236 & \new_[19839]_ ;
  assign \new_[19843]_  = ~A299 & A298;
  assign \new_[19846]_  = ~A302 & A300;
  assign \new_[19847]_  = \new_[19846]_  & \new_[19843]_ ;
  assign \new_[19848]_  = \new_[19847]_  & \new_[19840]_ ;
  assign \new_[19852]_  = ~A167 & A168;
  assign \new_[19853]_  = A169 & \new_[19852]_ ;
  assign \new_[19856]_  = A232 & A166;
  assign \new_[19859]_  = A234 & ~A233;
  assign \new_[19860]_  = \new_[19859]_  & \new_[19856]_ ;
  assign \new_[19861]_  = \new_[19860]_  & \new_[19853]_ ;
  assign \new_[19865]_  = A268 & ~A267;
  assign \new_[19866]_  = ~A236 & \new_[19865]_ ;
  assign \new_[19869]_  = A299 & ~A298;
  assign \new_[19872]_  = A301 & A300;
  assign \new_[19873]_  = \new_[19872]_  & \new_[19869]_ ;
  assign \new_[19874]_  = \new_[19873]_  & \new_[19866]_ ;
  assign \new_[19878]_  = ~A167 & A168;
  assign \new_[19879]_  = A169 & \new_[19878]_ ;
  assign \new_[19882]_  = A232 & A166;
  assign \new_[19885]_  = A234 & ~A233;
  assign \new_[19886]_  = \new_[19885]_  & \new_[19882]_ ;
  assign \new_[19887]_  = \new_[19886]_  & \new_[19879]_ ;
  assign \new_[19891]_  = A268 & ~A267;
  assign \new_[19892]_  = ~A236 & \new_[19891]_ ;
  assign \new_[19895]_  = A299 & ~A298;
  assign \new_[19898]_  = ~A302 & A300;
  assign \new_[19899]_  = \new_[19898]_  & \new_[19895]_ ;
  assign \new_[19900]_  = \new_[19899]_  & \new_[19892]_ ;
  assign \new_[19904]_  = ~A167 & A168;
  assign \new_[19905]_  = A169 & \new_[19904]_ ;
  assign \new_[19908]_  = A232 & A166;
  assign \new_[19911]_  = A234 & ~A233;
  assign \new_[19912]_  = \new_[19911]_  & \new_[19908]_ ;
  assign \new_[19913]_  = \new_[19912]_  & \new_[19905]_ ;
  assign \new_[19917]_  = ~A269 & ~A267;
  assign \new_[19918]_  = ~A236 & \new_[19917]_ ;
  assign \new_[19921]_  = ~A299 & A298;
  assign \new_[19924]_  = A301 & A300;
  assign \new_[19925]_  = \new_[19924]_  & \new_[19921]_ ;
  assign \new_[19926]_  = \new_[19925]_  & \new_[19918]_ ;
  assign \new_[19930]_  = ~A167 & A168;
  assign \new_[19931]_  = A169 & \new_[19930]_ ;
  assign \new_[19934]_  = A232 & A166;
  assign \new_[19937]_  = A234 & ~A233;
  assign \new_[19938]_  = \new_[19937]_  & \new_[19934]_ ;
  assign \new_[19939]_  = \new_[19938]_  & \new_[19931]_ ;
  assign \new_[19943]_  = ~A269 & ~A267;
  assign \new_[19944]_  = ~A236 & \new_[19943]_ ;
  assign \new_[19947]_  = ~A299 & A298;
  assign \new_[19950]_  = ~A302 & A300;
  assign \new_[19951]_  = \new_[19950]_  & \new_[19947]_ ;
  assign \new_[19952]_  = \new_[19951]_  & \new_[19944]_ ;
  assign \new_[19956]_  = ~A167 & A168;
  assign \new_[19957]_  = A169 & \new_[19956]_ ;
  assign \new_[19960]_  = A232 & A166;
  assign \new_[19963]_  = A234 & ~A233;
  assign \new_[19964]_  = \new_[19963]_  & \new_[19960]_ ;
  assign \new_[19965]_  = \new_[19964]_  & \new_[19957]_ ;
  assign \new_[19969]_  = ~A269 & ~A267;
  assign \new_[19970]_  = ~A236 & \new_[19969]_ ;
  assign \new_[19973]_  = A299 & ~A298;
  assign \new_[19976]_  = A301 & A300;
  assign \new_[19977]_  = \new_[19976]_  & \new_[19973]_ ;
  assign \new_[19978]_  = \new_[19977]_  & \new_[19970]_ ;
  assign \new_[19982]_  = ~A167 & A168;
  assign \new_[19983]_  = A169 & \new_[19982]_ ;
  assign \new_[19986]_  = A232 & A166;
  assign \new_[19989]_  = A234 & ~A233;
  assign \new_[19990]_  = \new_[19989]_  & \new_[19986]_ ;
  assign \new_[19991]_  = \new_[19990]_  & \new_[19983]_ ;
  assign \new_[19995]_  = ~A269 & ~A267;
  assign \new_[19996]_  = ~A236 & \new_[19995]_ ;
  assign \new_[19999]_  = A299 & ~A298;
  assign \new_[20002]_  = ~A302 & A300;
  assign \new_[20003]_  = \new_[20002]_  & \new_[19999]_ ;
  assign \new_[20004]_  = \new_[20003]_  & \new_[19996]_ ;
  assign \new_[20008]_  = ~A167 & A168;
  assign \new_[20009]_  = A169 & \new_[20008]_ ;
  assign \new_[20012]_  = A232 & A166;
  assign \new_[20015]_  = A234 & ~A233;
  assign \new_[20016]_  = \new_[20015]_  & \new_[20012]_ ;
  assign \new_[20017]_  = \new_[20016]_  & \new_[20009]_ ;
  assign \new_[20021]_  = A266 & A265;
  assign \new_[20022]_  = ~A236 & \new_[20021]_ ;
  assign \new_[20025]_  = ~A299 & A298;
  assign \new_[20028]_  = A301 & A300;
  assign \new_[20029]_  = \new_[20028]_  & \new_[20025]_ ;
  assign \new_[20030]_  = \new_[20029]_  & \new_[20022]_ ;
  assign \new_[20034]_  = ~A167 & A168;
  assign \new_[20035]_  = A169 & \new_[20034]_ ;
  assign \new_[20038]_  = A232 & A166;
  assign \new_[20041]_  = A234 & ~A233;
  assign \new_[20042]_  = \new_[20041]_  & \new_[20038]_ ;
  assign \new_[20043]_  = \new_[20042]_  & \new_[20035]_ ;
  assign \new_[20047]_  = A266 & A265;
  assign \new_[20048]_  = ~A236 & \new_[20047]_ ;
  assign \new_[20051]_  = ~A299 & A298;
  assign \new_[20054]_  = ~A302 & A300;
  assign \new_[20055]_  = \new_[20054]_  & \new_[20051]_ ;
  assign \new_[20056]_  = \new_[20055]_  & \new_[20048]_ ;
  assign \new_[20060]_  = ~A167 & A168;
  assign \new_[20061]_  = A169 & \new_[20060]_ ;
  assign \new_[20064]_  = A232 & A166;
  assign \new_[20067]_  = A234 & ~A233;
  assign \new_[20068]_  = \new_[20067]_  & \new_[20064]_ ;
  assign \new_[20069]_  = \new_[20068]_  & \new_[20061]_ ;
  assign \new_[20073]_  = A266 & A265;
  assign \new_[20074]_  = ~A236 & \new_[20073]_ ;
  assign \new_[20077]_  = A299 & ~A298;
  assign \new_[20080]_  = A301 & A300;
  assign \new_[20081]_  = \new_[20080]_  & \new_[20077]_ ;
  assign \new_[20082]_  = \new_[20081]_  & \new_[20074]_ ;
  assign \new_[20086]_  = ~A167 & A168;
  assign \new_[20087]_  = A169 & \new_[20086]_ ;
  assign \new_[20090]_  = A232 & A166;
  assign \new_[20093]_  = A234 & ~A233;
  assign \new_[20094]_  = \new_[20093]_  & \new_[20090]_ ;
  assign \new_[20095]_  = \new_[20094]_  & \new_[20087]_ ;
  assign \new_[20099]_  = A266 & A265;
  assign \new_[20100]_  = ~A236 & \new_[20099]_ ;
  assign \new_[20103]_  = A299 & ~A298;
  assign \new_[20106]_  = ~A302 & A300;
  assign \new_[20107]_  = \new_[20106]_  & \new_[20103]_ ;
  assign \new_[20108]_  = \new_[20107]_  & \new_[20100]_ ;
  assign \new_[20112]_  = ~A167 & A168;
  assign \new_[20113]_  = A169 & \new_[20112]_ ;
  assign \new_[20116]_  = A232 & A166;
  assign \new_[20119]_  = A234 & ~A233;
  assign \new_[20120]_  = \new_[20119]_  & \new_[20116]_ ;
  assign \new_[20121]_  = \new_[20120]_  & \new_[20113]_ ;
  assign \new_[20125]_  = ~A266 & ~A265;
  assign \new_[20126]_  = ~A236 & \new_[20125]_ ;
  assign \new_[20129]_  = ~A299 & A298;
  assign \new_[20132]_  = A301 & A300;
  assign \new_[20133]_  = \new_[20132]_  & \new_[20129]_ ;
  assign \new_[20134]_  = \new_[20133]_  & \new_[20126]_ ;
  assign \new_[20138]_  = ~A167 & A168;
  assign \new_[20139]_  = A169 & \new_[20138]_ ;
  assign \new_[20142]_  = A232 & A166;
  assign \new_[20145]_  = A234 & ~A233;
  assign \new_[20146]_  = \new_[20145]_  & \new_[20142]_ ;
  assign \new_[20147]_  = \new_[20146]_  & \new_[20139]_ ;
  assign \new_[20151]_  = ~A266 & ~A265;
  assign \new_[20152]_  = ~A236 & \new_[20151]_ ;
  assign \new_[20155]_  = ~A299 & A298;
  assign \new_[20158]_  = ~A302 & A300;
  assign \new_[20159]_  = \new_[20158]_  & \new_[20155]_ ;
  assign \new_[20160]_  = \new_[20159]_  & \new_[20152]_ ;
  assign \new_[20164]_  = ~A167 & A168;
  assign \new_[20165]_  = A169 & \new_[20164]_ ;
  assign \new_[20168]_  = A232 & A166;
  assign \new_[20171]_  = A234 & ~A233;
  assign \new_[20172]_  = \new_[20171]_  & \new_[20168]_ ;
  assign \new_[20173]_  = \new_[20172]_  & \new_[20165]_ ;
  assign \new_[20177]_  = ~A266 & ~A265;
  assign \new_[20178]_  = ~A236 & \new_[20177]_ ;
  assign \new_[20181]_  = A299 & ~A298;
  assign \new_[20184]_  = A301 & A300;
  assign \new_[20185]_  = \new_[20184]_  & \new_[20181]_ ;
  assign \new_[20186]_  = \new_[20185]_  & \new_[20178]_ ;
  assign \new_[20190]_  = ~A167 & A168;
  assign \new_[20191]_  = A169 & \new_[20190]_ ;
  assign \new_[20194]_  = A232 & A166;
  assign \new_[20197]_  = A234 & ~A233;
  assign \new_[20198]_  = \new_[20197]_  & \new_[20194]_ ;
  assign \new_[20199]_  = \new_[20198]_  & \new_[20191]_ ;
  assign \new_[20203]_  = ~A266 & ~A265;
  assign \new_[20204]_  = ~A236 & \new_[20203]_ ;
  assign \new_[20207]_  = A299 & ~A298;
  assign \new_[20210]_  = ~A302 & A300;
  assign \new_[20211]_  = \new_[20210]_  & \new_[20207]_ ;
  assign \new_[20212]_  = \new_[20211]_  & \new_[20204]_ ;
  assign \new_[20216]_  = A201 & A200;
  assign \new_[20217]_  = ~A199 & \new_[20216]_ ;
  assign \new_[20220]_  = ~A232 & A202;
  assign \new_[20223]_  = A234 & A233;
  assign \new_[20224]_  = \new_[20223]_  & \new_[20220]_ ;
  assign \new_[20225]_  = \new_[20224]_  & \new_[20217]_ ;
  assign \new_[20228]_  = A267 & A235;
  assign \new_[20231]_  = A269 & ~A268;
  assign \new_[20232]_  = \new_[20231]_  & \new_[20228]_ ;
  assign \new_[20235]_  = ~A299 & A298;
  assign \new_[20238]_  = A301 & A300;
  assign \new_[20239]_  = \new_[20238]_  & \new_[20235]_ ;
  assign \new_[20240]_  = \new_[20239]_  & \new_[20232]_ ;
  assign \new_[20244]_  = A201 & A200;
  assign \new_[20245]_  = ~A199 & \new_[20244]_ ;
  assign \new_[20248]_  = ~A232 & A202;
  assign \new_[20251]_  = A234 & A233;
  assign \new_[20252]_  = \new_[20251]_  & \new_[20248]_ ;
  assign \new_[20253]_  = \new_[20252]_  & \new_[20245]_ ;
  assign \new_[20256]_  = A267 & A235;
  assign \new_[20259]_  = A269 & ~A268;
  assign \new_[20260]_  = \new_[20259]_  & \new_[20256]_ ;
  assign \new_[20263]_  = ~A299 & A298;
  assign \new_[20266]_  = ~A302 & A300;
  assign \new_[20267]_  = \new_[20266]_  & \new_[20263]_ ;
  assign \new_[20268]_  = \new_[20267]_  & \new_[20260]_ ;
  assign \new_[20272]_  = A201 & A200;
  assign \new_[20273]_  = ~A199 & \new_[20272]_ ;
  assign \new_[20276]_  = ~A232 & A202;
  assign \new_[20279]_  = A234 & A233;
  assign \new_[20280]_  = \new_[20279]_  & \new_[20276]_ ;
  assign \new_[20281]_  = \new_[20280]_  & \new_[20273]_ ;
  assign \new_[20284]_  = A267 & A235;
  assign \new_[20287]_  = A269 & ~A268;
  assign \new_[20288]_  = \new_[20287]_  & \new_[20284]_ ;
  assign \new_[20291]_  = A299 & ~A298;
  assign \new_[20294]_  = A301 & A300;
  assign \new_[20295]_  = \new_[20294]_  & \new_[20291]_ ;
  assign \new_[20296]_  = \new_[20295]_  & \new_[20288]_ ;
  assign \new_[20300]_  = A201 & A200;
  assign \new_[20301]_  = ~A199 & \new_[20300]_ ;
  assign \new_[20304]_  = ~A232 & A202;
  assign \new_[20307]_  = A234 & A233;
  assign \new_[20308]_  = \new_[20307]_  & \new_[20304]_ ;
  assign \new_[20309]_  = \new_[20308]_  & \new_[20301]_ ;
  assign \new_[20312]_  = A267 & A235;
  assign \new_[20315]_  = A269 & ~A268;
  assign \new_[20316]_  = \new_[20315]_  & \new_[20312]_ ;
  assign \new_[20319]_  = A299 & ~A298;
  assign \new_[20322]_  = ~A302 & A300;
  assign \new_[20323]_  = \new_[20322]_  & \new_[20319]_ ;
  assign \new_[20324]_  = \new_[20323]_  & \new_[20316]_ ;
  assign \new_[20328]_  = A201 & A200;
  assign \new_[20329]_  = ~A199 & \new_[20328]_ ;
  assign \new_[20332]_  = ~A232 & A202;
  assign \new_[20335]_  = A234 & A233;
  assign \new_[20336]_  = \new_[20335]_  & \new_[20332]_ ;
  assign \new_[20337]_  = \new_[20336]_  & \new_[20329]_ ;
  assign \new_[20340]_  = ~A267 & A235;
  assign \new_[20343]_  = A298 & A268;
  assign \new_[20344]_  = \new_[20343]_  & \new_[20340]_ ;
  assign \new_[20347]_  = ~A300 & ~A299;
  assign \new_[20350]_  = A302 & ~A301;
  assign \new_[20351]_  = \new_[20350]_  & \new_[20347]_ ;
  assign \new_[20352]_  = \new_[20351]_  & \new_[20344]_ ;
  assign \new_[20356]_  = A201 & A200;
  assign \new_[20357]_  = ~A199 & \new_[20356]_ ;
  assign \new_[20360]_  = ~A232 & A202;
  assign \new_[20363]_  = A234 & A233;
  assign \new_[20364]_  = \new_[20363]_  & \new_[20360]_ ;
  assign \new_[20365]_  = \new_[20364]_  & \new_[20357]_ ;
  assign \new_[20368]_  = ~A267 & A235;
  assign \new_[20371]_  = ~A298 & A268;
  assign \new_[20372]_  = \new_[20371]_  & \new_[20368]_ ;
  assign \new_[20375]_  = ~A300 & A299;
  assign \new_[20378]_  = A302 & ~A301;
  assign \new_[20379]_  = \new_[20378]_  & \new_[20375]_ ;
  assign \new_[20380]_  = \new_[20379]_  & \new_[20372]_ ;
  assign \new_[20384]_  = A201 & A200;
  assign \new_[20385]_  = ~A199 & \new_[20384]_ ;
  assign \new_[20388]_  = ~A232 & A202;
  assign \new_[20391]_  = A234 & A233;
  assign \new_[20392]_  = \new_[20391]_  & \new_[20388]_ ;
  assign \new_[20393]_  = \new_[20392]_  & \new_[20385]_ ;
  assign \new_[20396]_  = ~A267 & A235;
  assign \new_[20399]_  = A298 & ~A269;
  assign \new_[20400]_  = \new_[20399]_  & \new_[20396]_ ;
  assign \new_[20403]_  = ~A300 & ~A299;
  assign \new_[20406]_  = A302 & ~A301;
  assign \new_[20407]_  = \new_[20406]_  & \new_[20403]_ ;
  assign \new_[20408]_  = \new_[20407]_  & \new_[20400]_ ;
  assign \new_[20412]_  = A201 & A200;
  assign \new_[20413]_  = ~A199 & \new_[20412]_ ;
  assign \new_[20416]_  = ~A232 & A202;
  assign \new_[20419]_  = A234 & A233;
  assign \new_[20420]_  = \new_[20419]_  & \new_[20416]_ ;
  assign \new_[20421]_  = \new_[20420]_  & \new_[20413]_ ;
  assign \new_[20424]_  = ~A267 & A235;
  assign \new_[20427]_  = ~A298 & ~A269;
  assign \new_[20428]_  = \new_[20427]_  & \new_[20424]_ ;
  assign \new_[20431]_  = ~A300 & A299;
  assign \new_[20434]_  = A302 & ~A301;
  assign \new_[20435]_  = \new_[20434]_  & \new_[20431]_ ;
  assign \new_[20436]_  = \new_[20435]_  & \new_[20428]_ ;
  assign \new_[20440]_  = A201 & A200;
  assign \new_[20441]_  = ~A199 & \new_[20440]_ ;
  assign \new_[20444]_  = ~A232 & A202;
  assign \new_[20447]_  = A234 & A233;
  assign \new_[20448]_  = \new_[20447]_  & \new_[20444]_ ;
  assign \new_[20449]_  = \new_[20448]_  & \new_[20441]_ ;
  assign \new_[20452]_  = A265 & A235;
  assign \new_[20455]_  = A298 & A266;
  assign \new_[20456]_  = \new_[20455]_  & \new_[20452]_ ;
  assign \new_[20459]_  = ~A300 & ~A299;
  assign \new_[20462]_  = A302 & ~A301;
  assign \new_[20463]_  = \new_[20462]_  & \new_[20459]_ ;
  assign \new_[20464]_  = \new_[20463]_  & \new_[20456]_ ;
  assign \new_[20468]_  = A201 & A200;
  assign \new_[20469]_  = ~A199 & \new_[20468]_ ;
  assign \new_[20472]_  = ~A232 & A202;
  assign \new_[20475]_  = A234 & A233;
  assign \new_[20476]_  = \new_[20475]_  & \new_[20472]_ ;
  assign \new_[20477]_  = \new_[20476]_  & \new_[20469]_ ;
  assign \new_[20480]_  = A265 & A235;
  assign \new_[20483]_  = ~A298 & A266;
  assign \new_[20484]_  = \new_[20483]_  & \new_[20480]_ ;
  assign \new_[20487]_  = ~A300 & A299;
  assign \new_[20490]_  = A302 & ~A301;
  assign \new_[20491]_  = \new_[20490]_  & \new_[20487]_ ;
  assign \new_[20492]_  = \new_[20491]_  & \new_[20484]_ ;
  assign \new_[20496]_  = A201 & A200;
  assign \new_[20497]_  = ~A199 & \new_[20496]_ ;
  assign \new_[20500]_  = ~A232 & A202;
  assign \new_[20503]_  = A234 & A233;
  assign \new_[20504]_  = \new_[20503]_  & \new_[20500]_ ;
  assign \new_[20505]_  = \new_[20504]_  & \new_[20497]_ ;
  assign \new_[20508]_  = ~A265 & A235;
  assign \new_[20511]_  = A298 & ~A266;
  assign \new_[20512]_  = \new_[20511]_  & \new_[20508]_ ;
  assign \new_[20515]_  = ~A300 & ~A299;
  assign \new_[20518]_  = A302 & ~A301;
  assign \new_[20519]_  = \new_[20518]_  & \new_[20515]_ ;
  assign \new_[20520]_  = \new_[20519]_  & \new_[20512]_ ;
  assign \new_[20524]_  = A201 & A200;
  assign \new_[20525]_  = ~A199 & \new_[20524]_ ;
  assign \new_[20528]_  = ~A232 & A202;
  assign \new_[20531]_  = A234 & A233;
  assign \new_[20532]_  = \new_[20531]_  & \new_[20528]_ ;
  assign \new_[20533]_  = \new_[20532]_  & \new_[20525]_ ;
  assign \new_[20536]_  = ~A265 & A235;
  assign \new_[20539]_  = ~A298 & ~A266;
  assign \new_[20540]_  = \new_[20539]_  & \new_[20536]_ ;
  assign \new_[20543]_  = ~A300 & A299;
  assign \new_[20546]_  = A302 & ~A301;
  assign \new_[20547]_  = \new_[20546]_  & \new_[20543]_ ;
  assign \new_[20548]_  = \new_[20547]_  & \new_[20540]_ ;
  assign \new_[20552]_  = A201 & A200;
  assign \new_[20553]_  = ~A199 & \new_[20552]_ ;
  assign \new_[20556]_  = ~A232 & A202;
  assign \new_[20559]_  = A234 & A233;
  assign \new_[20560]_  = \new_[20559]_  & \new_[20556]_ ;
  assign \new_[20561]_  = \new_[20560]_  & \new_[20553]_ ;
  assign \new_[20564]_  = A267 & ~A236;
  assign \new_[20567]_  = A269 & ~A268;
  assign \new_[20568]_  = \new_[20567]_  & \new_[20564]_ ;
  assign \new_[20571]_  = ~A299 & A298;
  assign \new_[20574]_  = A301 & A300;
  assign \new_[20575]_  = \new_[20574]_  & \new_[20571]_ ;
  assign \new_[20576]_  = \new_[20575]_  & \new_[20568]_ ;
  assign \new_[20580]_  = A201 & A200;
  assign \new_[20581]_  = ~A199 & \new_[20580]_ ;
  assign \new_[20584]_  = ~A232 & A202;
  assign \new_[20587]_  = A234 & A233;
  assign \new_[20588]_  = \new_[20587]_  & \new_[20584]_ ;
  assign \new_[20589]_  = \new_[20588]_  & \new_[20581]_ ;
  assign \new_[20592]_  = A267 & ~A236;
  assign \new_[20595]_  = A269 & ~A268;
  assign \new_[20596]_  = \new_[20595]_  & \new_[20592]_ ;
  assign \new_[20599]_  = ~A299 & A298;
  assign \new_[20602]_  = ~A302 & A300;
  assign \new_[20603]_  = \new_[20602]_  & \new_[20599]_ ;
  assign \new_[20604]_  = \new_[20603]_  & \new_[20596]_ ;
  assign \new_[20608]_  = A201 & A200;
  assign \new_[20609]_  = ~A199 & \new_[20608]_ ;
  assign \new_[20612]_  = ~A232 & A202;
  assign \new_[20615]_  = A234 & A233;
  assign \new_[20616]_  = \new_[20615]_  & \new_[20612]_ ;
  assign \new_[20617]_  = \new_[20616]_  & \new_[20609]_ ;
  assign \new_[20620]_  = A267 & ~A236;
  assign \new_[20623]_  = A269 & ~A268;
  assign \new_[20624]_  = \new_[20623]_  & \new_[20620]_ ;
  assign \new_[20627]_  = A299 & ~A298;
  assign \new_[20630]_  = A301 & A300;
  assign \new_[20631]_  = \new_[20630]_  & \new_[20627]_ ;
  assign \new_[20632]_  = \new_[20631]_  & \new_[20624]_ ;
  assign \new_[20636]_  = A201 & A200;
  assign \new_[20637]_  = ~A199 & \new_[20636]_ ;
  assign \new_[20640]_  = ~A232 & A202;
  assign \new_[20643]_  = A234 & A233;
  assign \new_[20644]_  = \new_[20643]_  & \new_[20640]_ ;
  assign \new_[20645]_  = \new_[20644]_  & \new_[20637]_ ;
  assign \new_[20648]_  = A267 & ~A236;
  assign \new_[20651]_  = A269 & ~A268;
  assign \new_[20652]_  = \new_[20651]_  & \new_[20648]_ ;
  assign \new_[20655]_  = A299 & ~A298;
  assign \new_[20658]_  = ~A302 & A300;
  assign \new_[20659]_  = \new_[20658]_  & \new_[20655]_ ;
  assign \new_[20660]_  = \new_[20659]_  & \new_[20652]_ ;
  assign \new_[20664]_  = A201 & A200;
  assign \new_[20665]_  = ~A199 & \new_[20664]_ ;
  assign \new_[20668]_  = ~A232 & A202;
  assign \new_[20671]_  = A234 & A233;
  assign \new_[20672]_  = \new_[20671]_  & \new_[20668]_ ;
  assign \new_[20673]_  = \new_[20672]_  & \new_[20665]_ ;
  assign \new_[20676]_  = ~A267 & ~A236;
  assign \new_[20679]_  = A298 & A268;
  assign \new_[20680]_  = \new_[20679]_  & \new_[20676]_ ;
  assign \new_[20683]_  = ~A300 & ~A299;
  assign \new_[20686]_  = A302 & ~A301;
  assign \new_[20687]_  = \new_[20686]_  & \new_[20683]_ ;
  assign \new_[20688]_  = \new_[20687]_  & \new_[20680]_ ;
  assign \new_[20692]_  = A201 & A200;
  assign \new_[20693]_  = ~A199 & \new_[20692]_ ;
  assign \new_[20696]_  = ~A232 & A202;
  assign \new_[20699]_  = A234 & A233;
  assign \new_[20700]_  = \new_[20699]_  & \new_[20696]_ ;
  assign \new_[20701]_  = \new_[20700]_  & \new_[20693]_ ;
  assign \new_[20704]_  = ~A267 & ~A236;
  assign \new_[20707]_  = ~A298 & A268;
  assign \new_[20708]_  = \new_[20707]_  & \new_[20704]_ ;
  assign \new_[20711]_  = ~A300 & A299;
  assign \new_[20714]_  = A302 & ~A301;
  assign \new_[20715]_  = \new_[20714]_  & \new_[20711]_ ;
  assign \new_[20716]_  = \new_[20715]_  & \new_[20708]_ ;
  assign \new_[20720]_  = A201 & A200;
  assign \new_[20721]_  = ~A199 & \new_[20720]_ ;
  assign \new_[20724]_  = ~A232 & A202;
  assign \new_[20727]_  = A234 & A233;
  assign \new_[20728]_  = \new_[20727]_  & \new_[20724]_ ;
  assign \new_[20729]_  = \new_[20728]_  & \new_[20721]_ ;
  assign \new_[20732]_  = ~A267 & ~A236;
  assign \new_[20735]_  = A298 & ~A269;
  assign \new_[20736]_  = \new_[20735]_  & \new_[20732]_ ;
  assign \new_[20739]_  = ~A300 & ~A299;
  assign \new_[20742]_  = A302 & ~A301;
  assign \new_[20743]_  = \new_[20742]_  & \new_[20739]_ ;
  assign \new_[20744]_  = \new_[20743]_  & \new_[20736]_ ;
  assign \new_[20748]_  = A201 & A200;
  assign \new_[20749]_  = ~A199 & \new_[20748]_ ;
  assign \new_[20752]_  = ~A232 & A202;
  assign \new_[20755]_  = A234 & A233;
  assign \new_[20756]_  = \new_[20755]_  & \new_[20752]_ ;
  assign \new_[20757]_  = \new_[20756]_  & \new_[20749]_ ;
  assign \new_[20760]_  = ~A267 & ~A236;
  assign \new_[20763]_  = ~A298 & ~A269;
  assign \new_[20764]_  = \new_[20763]_  & \new_[20760]_ ;
  assign \new_[20767]_  = ~A300 & A299;
  assign \new_[20770]_  = A302 & ~A301;
  assign \new_[20771]_  = \new_[20770]_  & \new_[20767]_ ;
  assign \new_[20772]_  = \new_[20771]_  & \new_[20764]_ ;
  assign \new_[20776]_  = A201 & A200;
  assign \new_[20777]_  = ~A199 & \new_[20776]_ ;
  assign \new_[20780]_  = ~A232 & A202;
  assign \new_[20783]_  = A234 & A233;
  assign \new_[20784]_  = \new_[20783]_  & \new_[20780]_ ;
  assign \new_[20785]_  = \new_[20784]_  & \new_[20777]_ ;
  assign \new_[20788]_  = A265 & ~A236;
  assign \new_[20791]_  = A298 & A266;
  assign \new_[20792]_  = \new_[20791]_  & \new_[20788]_ ;
  assign \new_[20795]_  = ~A300 & ~A299;
  assign \new_[20798]_  = A302 & ~A301;
  assign \new_[20799]_  = \new_[20798]_  & \new_[20795]_ ;
  assign \new_[20800]_  = \new_[20799]_  & \new_[20792]_ ;
  assign \new_[20804]_  = A201 & A200;
  assign \new_[20805]_  = ~A199 & \new_[20804]_ ;
  assign \new_[20808]_  = ~A232 & A202;
  assign \new_[20811]_  = A234 & A233;
  assign \new_[20812]_  = \new_[20811]_  & \new_[20808]_ ;
  assign \new_[20813]_  = \new_[20812]_  & \new_[20805]_ ;
  assign \new_[20816]_  = A265 & ~A236;
  assign \new_[20819]_  = ~A298 & A266;
  assign \new_[20820]_  = \new_[20819]_  & \new_[20816]_ ;
  assign \new_[20823]_  = ~A300 & A299;
  assign \new_[20826]_  = A302 & ~A301;
  assign \new_[20827]_  = \new_[20826]_  & \new_[20823]_ ;
  assign \new_[20828]_  = \new_[20827]_  & \new_[20820]_ ;
  assign \new_[20832]_  = A201 & A200;
  assign \new_[20833]_  = ~A199 & \new_[20832]_ ;
  assign \new_[20836]_  = ~A232 & A202;
  assign \new_[20839]_  = A234 & A233;
  assign \new_[20840]_  = \new_[20839]_  & \new_[20836]_ ;
  assign \new_[20841]_  = \new_[20840]_  & \new_[20833]_ ;
  assign \new_[20844]_  = ~A265 & ~A236;
  assign \new_[20847]_  = A298 & ~A266;
  assign \new_[20848]_  = \new_[20847]_  & \new_[20844]_ ;
  assign \new_[20851]_  = ~A300 & ~A299;
  assign \new_[20854]_  = A302 & ~A301;
  assign \new_[20855]_  = \new_[20854]_  & \new_[20851]_ ;
  assign \new_[20856]_  = \new_[20855]_  & \new_[20848]_ ;
  assign \new_[20860]_  = A201 & A200;
  assign \new_[20861]_  = ~A199 & \new_[20860]_ ;
  assign \new_[20864]_  = ~A232 & A202;
  assign \new_[20867]_  = A234 & A233;
  assign \new_[20868]_  = \new_[20867]_  & \new_[20864]_ ;
  assign \new_[20869]_  = \new_[20868]_  & \new_[20861]_ ;
  assign \new_[20872]_  = ~A265 & ~A236;
  assign \new_[20875]_  = ~A298 & ~A266;
  assign \new_[20876]_  = \new_[20875]_  & \new_[20872]_ ;
  assign \new_[20879]_  = ~A300 & A299;
  assign \new_[20882]_  = A302 & ~A301;
  assign \new_[20883]_  = \new_[20882]_  & \new_[20879]_ ;
  assign \new_[20884]_  = \new_[20883]_  & \new_[20876]_ ;
  assign \new_[20888]_  = A201 & A200;
  assign \new_[20889]_  = ~A199 & \new_[20888]_ ;
  assign \new_[20892]_  = ~A232 & A202;
  assign \new_[20895]_  = ~A234 & A233;
  assign \new_[20896]_  = \new_[20895]_  & \new_[20892]_ ;
  assign \new_[20897]_  = \new_[20896]_  & \new_[20889]_ ;
  assign \new_[20900]_  = A236 & ~A235;
  assign \new_[20903]_  = A268 & ~A267;
  assign \new_[20904]_  = \new_[20903]_  & \new_[20900]_ ;
  assign \new_[20907]_  = ~A299 & A298;
  assign \new_[20910]_  = A301 & A300;
  assign \new_[20911]_  = \new_[20910]_  & \new_[20907]_ ;
  assign \new_[20912]_  = \new_[20911]_  & \new_[20904]_ ;
  assign \new_[20916]_  = A201 & A200;
  assign \new_[20917]_  = ~A199 & \new_[20916]_ ;
  assign \new_[20920]_  = ~A232 & A202;
  assign \new_[20923]_  = ~A234 & A233;
  assign \new_[20924]_  = \new_[20923]_  & \new_[20920]_ ;
  assign \new_[20925]_  = \new_[20924]_  & \new_[20917]_ ;
  assign \new_[20928]_  = A236 & ~A235;
  assign \new_[20931]_  = A268 & ~A267;
  assign \new_[20932]_  = \new_[20931]_  & \new_[20928]_ ;
  assign \new_[20935]_  = ~A299 & A298;
  assign \new_[20938]_  = ~A302 & A300;
  assign \new_[20939]_  = \new_[20938]_  & \new_[20935]_ ;
  assign \new_[20940]_  = \new_[20939]_  & \new_[20932]_ ;
  assign \new_[20944]_  = A201 & A200;
  assign \new_[20945]_  = ~A199 & \new_[20944]_ ;
  assign \new_[20948]_  = ~A232 & A202;
  assign \new_[20951]_  = ~A234 & A233;
  assign \new_[20952]_  = \new_[20951]_  & \new_[20948]_ ;
  assign \new_[20953]_  = \new_[20952]_  & \new_[20945]_ ;
  assign \new_[20956]_  = A236 & ~A235;
  assign \new_[20959]_  = A268 & ~A267;
  assign \new_[20960]_  = \new_[20959]_  & \new_[20956]_ ;
  assign \new_[20963]_  = A299 & ~A298;
  assign \new_[20966]_  = A301 & A300;
  assign \new_[20967]_  = \new_[20966]_  & \new_[20963]_ ;
  assign \new_[20968]_  = \new_[20967]_  & \new_[20960]_ ;
  assign \new_[20972]_  = A201 & A200;
  assign \new_[20973]_  = ~A199 & \new_[20972]_ ;
  assign \new_[20976]_  = ~A232 & A202;
  assign \new_[20979]_  = ~A234 & A233;
  assign \new_[20980]_  = \new_[20979]_  & \new_[20976]_ ;
  assign \new_[20981]_  = \new_[20980]_  & \new_[20973]_ ;
  assign \new_[20984]_  = A236 & ~A235;
  assign \new_[20987]_  = A268 & ~A267;
  assign \new_[20988]_  = \new_[20987]_  & \new_[20984]_ ;
  assign \new_[20991]_  = A299 & ~A298;
  assign \new_[20994]_  = ~A302 & A300;
  assign \new_[20995]_  = \new_[20994]_  & \new_[20991]_ ;
  assign \new_[20996]_  = \new_[20995]_  & \new_[20988]_ ;
  assign \new_[21000]_  = A201 & A200;
  assign \new_[21001]_  = ~A199 & \new_[21000]_ ;
  assign \new_[21004]_  = ~A232 & A202;
  assign \new_[21007]_  = ~A234 & A233;
  assign \new_[21008]_  = \new_[21007]_  & \new_[21004]_ ;
  assign \new_[21009]_  = \new_[21008]_  & \new_[21001]_ ;
  assign \new_[21012]_  = A236 & ~A235;
  assign \new_[21015]_  = ~A269 & ~A267;
  assign \new_[21016]_  = \new_[21015]_  & \new_[21012]_ ;
  assign \new_[21019]_  = ~A299 & A298;
  assign \new_[21022]_  = A301 & A300;
  assign \new_[21023]_  = \new_[21022]_  & \new_[21019]_ ;
  assign \new_[21024]_  = \new_[21023]_  & \new_[21016]_ ;
  assign \new_[21028]_  = A201 & A200;
  assign \new_[21029]_  = ~A199 & \new_[21028]_ ;
  assign \new_[21032]_  = ~A232 & A202;
  assign \new_[21035]_  = ~A234 & A233;
  assign \new_[21036]_  = \new_[21035]_  & \new_[21032]_ ;
  assign \new_[21037]_  = \new_[21036]_  & \new_[21029]_ ;
  assign \new_[21040]_  = A236 & ~A235;
  assign \new_[21043]_  = ~A269 & ~A267;
  assign \new_[21044]_  = \new_[21043]_  & \new_[21040]_ ;
  assign \new_[21047]_  = ~A299 & A298;
  assign \new_[21050]_  = ~A302 & A300;
  assign \new_[21051]_  = \new_[21050]_  & \new_[21047]_ ;
  assign \new_[21052]_  = \new_[21051]_  & \new_[21044]_ ;
  assign \new_[21056]_  = A201 & A200;
  assign \new_[21057]_  = ~A199 & \new_[21056]_ ;
  assign \new_[21060]_  = ~A232 & A202;
  assign \new_[21063]_  = ~A234 & A233;
  assign \new_[21064]_  = \new_[21063]_  & \new_[21060]_ ;
  assign \new_[21065]_  = \new_[21064]_  & \new_[21057]_ ;
  assign \new_[21068]_  = A236 & ~A235;
  assign \new_[21071]_  = ~A269 & ~A267;
  assign \new_[21072]_  = \new_[21071]_  & \new_[21068]_ ;
  assign \new_[21075]_  = A299 & ~A298;
  assign \new_[21078]_  = A301 & A300;
  assign \new_[21079]_  = \new_[21078]_  & \new_[21075]_ ;
  assign \new_[21080]_  = \new_[21079]_  & \new_[21072]_ ;
  assign \new_[21084]_  = A201 & A200;
  assign \new_[21085]_  = ~A199 & \new_[21084]_ ;
  assign \new_[21088]_  = ~A232 & A202;
  assign \new_[21091]_  = ~A234 & A233;
  assign \new_[21092]_  = \new_[21091]_  & \new_[21088]_ ;
  assign \new_[21093]_  = \new_[21092]_  & \new_[21085]_ ;
  assign \new_[21096]_  = A236 & ~A235;
  assign \new_[21099]_  = ~A269 & ~A267;
  assign \new_[21100]_  = \new_[21099]_  & \new_[21096]_ ;
  assign \new_[21103]_  = A299 & ~A298;
  assign \new_[21106]_  = ~A302 & A300;
  assign \new_[21107]_  = \new_[21106]_  & \new_[21103]_ ;
  assign \new_[21108]_  = \new_[21107]_  & \new_[21100]_ ;
  assign \new_[21112]_  = A201 & A200;
  assign \new_[21113]_  = ~A199 & \new_[21112]_ ;
  assign \new_[21116]_  = ~A232 & A202;
  assign \new_[21119]_  = ~A234 & A233;
  assign \new_[21120]_  = \new_[21119]_  & \new_[21116]_ ;
  assign \new_[21121]_  = \new_[21120]_  & \new_[21113]_ ;
  assign \new_[21124]_  = A236 & ~A235;
  assign \new_[21127]_  = A266 & A265;
  assign \new_[21128]_  = \new_[21127]_  & \new_[21124]_ ;
  assign \new_[21131]_  = ~A299 & A298;
  assign \new_[21134]_  = A301 & A300;
  assign \new_[21135]_  = \new_[21134]_  & \new_[21131]_ ;
  assign \new_[21136]_  = \new_[21135]_  & \new_[21128]_ ;
  assign \new_[21140]_  = A201 & A200;
  assign \new_[21141]_  = ~A199 & \new_[21140]_ ;
  assign \new_[21144]_  = ~A232 & A202;
  assign \new_[21147]_  = ~A234 & A233;
  assign \new_[21148]_  = \new_[21147]_  & \new_[21144]_ ;
  assign \new_[21149]_  = \new_[21148]_  & \new_[21141]_ ;
  assign \new_[21152]_  = A236 & ~A235;
  assign \new_[21155]_  = A266 & A265;
  assign \new_[21156]_  = \new_[21155]_  & \new_[21152]_ ;
  assign \new_[21159]_  = ~A299 & A298;
  assign \new_[21162]_  = ~A302 & A300;
  assign \new_[21163]_  = \new_[21162]_  & \new_[21159]_ ;
  assign \new_[21164]_  = \new_[21163]_  & \new_[21156]_ ;
  assign \new_[21168]_  = A201 & A200;
  assign \new_[21169]_  = ~A199 & \new_[21168]_ ;
  assign \new_[21172]_  = ~A232 & A202;
  assign \new_[21175]_  = ~A234 & A233;
  assign \new_[21176]_  = \new_[21175]_  & \new_[21172]_ ;
  assign \new_[21177]_  = \new_[21176]_  & \new_[21169]_ ;
  assign \new_[21180]_  = A236 & ~A235;
  assign \new_[21183]_  = A266 & A265;
  assign \new_[21184]_  = \new_[21183]_  & \new_[21180]_ ;
  assign \new_[21187]_  = A299 & ~A298;
  assign \new_[21190]_  = A301 & A300;
  assign \new_[21191]_  = \new_[21190]_  & \new_[21187]_ ;
  assign \new_[21192]_  = \new_[21191]_  & \new_[21184]_ ;
  assign \new_[21196]_  = A201 & A200;
  assign \new_[21197]_  = ~A199 & \new_[21196]_ ;
  assign \new_[21200]_  = ~A232 & A202;
  assign \new_[21203]_  = ~A234 & A233;
  assign \new_[21204]_  = \new_[21203]_  & \new_[21200]_ ;
  assign \new_[21205]_  = \new_[21204]_  & \new_[21197]_ ;
  assign \new_[21208]_  = A236 & ~A235;
  assign \new_[21211]_  = A266 & A265;
  assign \new_[21212]_  = \new_[21211]_  & \new_[21208]_ ;
  assign \new_[21215]_  = A299 & ~A298;
  assign \new_[21218]_  = ~A302 & A300;
  assign \new_[21219]_  = \new_[21218]_  & \new_[21215]_ ;
  assign \new_[21220]_  = \new_[21219]_  & \new_[21212]_ ;
  assign \new_[21224]_  = A201 & A200;
  assign \new_[21225]_  = ~A199 & \new_[21224]_ ;
  assign \new_[21228]_  = ~A232 & A202;
  assign \new_[21231]_  = ~A234 & A233;
  assign \new_[21232]_  = \new_[21231]_  & \new_[21228]_ ;
  assign \new_[21233]_  = \new_[21232]_  & \new_[21225]_ ;
  assign \new_[21236]_  = A236 & ~A235;
  assign \new_[21239]_  = ~A266 & ~A265;
  assign \new_[21240]_  = \new_[21239]_  & \new_[21236]_ ;
  assign \new_[21243]_  = ~A299 & A298;
  assign \new_[21246]_  = A301 & A300;
  assign \new_[21247]_  = \new_[21246]_  & \new_[21243]_ ;
  assign \new_[21248]_  = \new_[21247]_  & \new_[21240]_ ;
  assign \new_[21252]_  = A201 & A200;
  assign \new_[21253]_  = ~A199 & \new_[21252]_ ;
  assign \new_[21256]_  = ~A232 & A202;
  assign \new_[21259]_  = ~A234 & A233;
  assign \new_[21260]_  = \new_[21259]_  & \new_[21256]_ ;
  assign \new_[21261]_  = \new_[21260]_  & \new_[21253]_ ;
  assign \new_[21264]_  = A236 & ~A235;
  assign \new_[21267]_  = ~A266 & ~A265;
  assign \new_[21268]_  = \new_[21267]_  & \new_[21264]_ ;
  assign \new_[21271]_  = ~A299 & A298;
  assign \new_[21274]_  = ~A302 & A300;
  assign \new_[21275]_  = \new_[21274]_  & \new_[21271]_ ;
  assign \new_[21276]_  = \new_[21275]_  & \new_[21268]_ ;
  assign \new_[21280]_  = A201 & A200;
  assign \new_[21281]_  = ~A199 & \new_[21280]_ ;
  assign \new_[21284]_  = ~A232 & A202;
  assign \new_[21287]_  = ~A234 & A233;
  assign \new_[21288]_  = \new_[21287]_  & \new_[21284]_ ;
  assign \new_[21289]_  = \new_[21288]_  & \new_[21281]_ ;
  assign \new_[21292]_  = A236 & ~A235;
  assign \new_[21295]_  = ~A266 & ~A265;
  assign \new_[21296]_  = \new_[21295]_  & \new_[21292]_ ;
  assign \new_[21299]_  = A299 & ~A298;
  assign \new_[21302]_  = A301 & A300;
  assign \new_[21303]_  = \new_[21302]_  & \new_[21299]_ ;
  assign \new_[21304]_  = \new_[21303]_  & \new_[21296]_ ;
  assign \new_[21308]_  = A201 & A200;
  assign \new_[21309]_  = ~A199 & \new_[21308]_ ;
  assign \new_[21312]_  = ~A232 & A202;
  assign \new_[21315]_  = ~A234 & A233;
  assign \new_[21316]_  = \new_[21315]_  & \new_[21312]_ ;
  assign \new_[21317]_  = \new_[21316]_  & \new_[21309]_ ;
  assign \new_[21320]_  = A236 & ~A235;
  assign \new_[21323]_  = ~A266 & ~A265;
  assign \new_[21324]_  = \new_[21323]_  & \new_[21320]_ ;
  assign \new_[21327]_  = A299 & ~A298;
  assign \new_[21330]_  = ~A302 & A300;
  assign \new_[21331]_  = \new_[21330]_  & \new_[21327]_ ;
  assign \new_[21332]_  = \new_[21331]_  & \new_[21324]_ ;
  assign \new_[21336]_  = A201 & A200;
  assign \new_[21337]_  = ~A199 & \new_[21336]_ ;
  assign \new_[21340]_  = A232 & A202;
  assign \new_[21343]_  = A234 & ~A233;
  assign \new_[21344]_  = \new_[21343]_  & \new_[21340]_ ;
  assign \new_[21345]_  = \new_[21344]_  & \new_[21337]_ ;
  assign \new_[21348]_  = A267 & A235;
  assign \new_[21351]_  = A269 & ~A268;
  assign \new_[21352]_  = \new_[21351]_  & \new_[21348]_ ;
  assign \new_[21355]_  = ~A299 & A298;
  assign \new_[21358]_  = A301 & A300;
  assign \new_[21359]_  = \new_[21358]_  & \new_[21355]_ ;
  assign \new_[21360]_  = \new_[21359]_  & \new_[21352]_ ;
  assign \new_[21364]_  = A201 & A200;
  assign \new_[21365]_  = ~A199 & \new_[21364]_ ;
  assign \new_[21368]_  = A232 & A202;
  assign \new_[21371]_  = A234 & ~A233;
  assign \new_[21372]_  = \new_[21371]_  & \new_[21368]_ ;
  assign \new_[21373]_  = \new_[21372]_  & \new_[21365]_ ;
  assign \new_[21376]_  = A267 & A235;
  assign \new_[21379]_  = A269 & ~A268;
  assign \new_[21380]_  = \new_[21379]_  & \new_[21376]_ ;
  assign \new_[21383]_  = ~A299 & A298;
  assign \new_[21386]_  = ~A302 & A300;
  assign \new_[21387]_  = \new_[21386]_  & \new_[21383]_ ;
  assign \new_[21388]_  = \new_[21387]_  & \new_[21380]_ ;
  assign \new_[21392]_  = A201 & A200;
  assign \new_[21393]_  = ~A199 & \new_[21392]_ ;
  assign \new_[21396]_  = A232 & A202;
  assign \new_[21399]_  = A234 & ~A233;
  assign \new_[21400]_  = \new_[21399]_  & \new_[21396]_ ;
  assign \new_[21401]_  = \new_[21400]_  & \new_[21393]_ ;
  assign \new_[21404]_  = A267 & A235;
  assign \new_[21407]_  = A269 & ~A268;
  assign \new_[21408]_  = \new_[21407]_  & \new_[21404]_ ;
  assign \new_[21411]_  = A299 & ~A298;
  assign \new_[21414]_  = A301 & A300;
  assign \new_[21415]_  = \new_[21414]_  & \new_[21411]_ ;
  assign \new_[21416]_  = \new_[21415]_  & \new_[21408]_ ;
  assign \new_[21420]_  = A201 & A200;
  assign \new_[21421]_  = ~A199 & \new_[21420]_ ;
  assign \new_[21424]_  = A232 & A202;
  assign \new_[21427]_  = A234 & ~A233;
  assign \new_[21428]_  = \new_[21427]_  & \new_[21424]_ ;
  assign \new_[21429]_  = \new_[21428]_  & \new_[21421]_ ;
  assign \new_[21432]_  = A267 & A235;
  assign \new_[21435]_  = A269 & ~A268;
  assign \new_[21436]_  = \new_[21435]_  & \new_[21432]_ ;
  assign \new_[21439]_  = A299 & ~A298;
  assign \new_[21442]_  = ~A302 & A300;
  assign \new_[21443]_  = \new_[21442]_  & \new_[21439]_ ;
  assign \new_[21444]_  = \new_[21443]_  & \new_[21436]_ ;
  assign \new_[21448]_  = A201 & A200;
  assign \new_[21449]_  = ~A199 & \new_[21448]_ ;
  assign \new_[21452]_  = A232 & A202;
  assign \new_[21455]_  = A234 & ~A233;
  assign \new_[21456]_  = \new_[21455]_  & \new_[21452]_ ;
  assign \new_[21457]_  = \new_[21456]_  & \new_[21449]_ ;
  assign \new_[21460]_  = ~A267 & A235;
  assign \new_[21463]_  = A298 & A268;
  assign \new_[21464]_  = \new_[21463]_  & \new_[21460]_ ;
  assign \new_[21467]_  = ~A300 & ~A299;
  assign \new_[21470]_  = A302 & ~A301;
  assign \new_[21471]_  = \new_[21470]_  & \new_[21467]_ ;
  assign \new_[21472]_  = \new_[21471]_  & \new_[21464]_ ;
  assign \new_[21476]_  = A201 & A200;
  assign \new_[21477]_  = ~A199 & \new_[21476]_ ;
  assign \new_[21480]_  = A232 & A202;
  assign \new_[21483]_  = A234 & ~A233;
  assign \new_[21484]_  = \new_[21483]_  & \new_[21480]_ ;
  assign \new_[21485]_  = \new_[21484]_  & \new_[21477]_ ;
  assign \new_[21488]_  = ~A267 & A235;
  assign \new_[21491]_  = ~A298 & A268;
  assign \new_[21492]_  = \new_[21491]_  & \new_[21488]_ ;
  assign \new_[21495]_  = ~A300 & A299;
  assign \new_[21498]_  = A302 & ~A301;
  assign \new_[21499]_  = \new_[21498]_  & \new_[21495]_ ;
  assign \new_[21500]_  = \new_[21499]_  & \new_[21492]_ ;
  assign \new_[21504]_  = A201 & A200;
  assign \new_[21505]_  = ~A199 & \new_[21504]_ ;
  assign \new_[21508]_  = A232 & A202;
  assign \new_[21511]_  = A234 & ~A233;
  assign \new_[21512]_  = \new_[21511]_  & \new_[21508]_ ;
  assign \new_[21513]_  = \new_[21512]_  & \new_[21505]_ ;
  assign \new_[21516]_  = ~A267 & A235;
  assign \new_[21519]_  = A298 & ~A269;
  assign \new_[21520]_  = \new_[21519]_  & \new_[21516]_ ;
  assign \new_[21523]_  = ~A300 & ~A299;
  assign \new_[21526]_  = A302 & ~A301;
  assign \new_[21527]_  = \new_[21526]_  & \new_[21523]_ ;
  assign \new_[21528]_  = \new_[21527]_  & \new_[21520]_ ;
  assign \new_[21532]_  = A201 & A200;
  assign \new_[21533]_  = ~A199 & \new_[21532]_ ;
  assign \new_[21536]_  = A232 & A202;
  assign \new_[21539]_  = A234 & ~A233;
  assign \new_[21540]_  = \new_[21539]_  & \new_[21536]_ ;
  assign \new_[21541]_  = \new_[21540]_  & \new_[21533]_ ;
  assign \new_[21544]_  = ~A267 & A235;
  assign \new_[21547]_  = ~A298 & ~A269;
  assign \new_[21548]_  = \new_[21547]_  & \new_[21544]_ ;
  assign \new_[21551]_  = ~A300 & A299;
  assign \new_[21554]_  = A302 & ~A301;
  assign \new_[21555]_  = \new_[21554]_  & \new_[21551]_ ;
  assign \new_[21556]_  = \new_[21555]_  & \new_[21548]_ ;
  assign \new_[21560]_  = A201 & A200;
  assign \new_[21561]_  = ~A199 & \new_[21560]_ ;
  assign \new_[21564]_  = A232 & A202;
  assign \new_[21567]_  = A234 & ~A233;
  assign \new_[21568]_  = \new_[21567]_  & \new_[21564]_ ;
  assign \new_[21569]_  = \new_[21568]_  & \new_[21561]_ ;
  assign \new_[21572]_  = A265 & A235;
  assign \new_[21575]_  = A298 & A266;
  assign \new_[21576]_  = \new_[21575]_  & \new_[21572]_ ;
  assign \new_[21579]_  = ~A300 & ~A299;
  assign \new_[21582]_  = A302 & ~A301;
  assign \new_[21583]_  = \new_[21582]_  & \new_[21579]_ ;
  assign \new_[21584]_  = \new_[21583]_  & \new_[21576]_ ;
  assign \new_[21588]_  = A201 & A200;
  assign \new_[21589]_  = ~A199 & \new_[21588]_ ;
  assign \new_[21592]_  = A232 & A202;
  assign \new_[21595]_  = A234 & ~A233;
  assign \new_[21596]_  = \new_[21595]_  & \new_[21592]_ ;
  assign \new_[21597]_  = \new_[21596]_  & \new_[21589]_ ;
  assign \new_[21600]_  = A265 & A235;
  assign \new_[21603]_  = ~A298 & A266;
  assign \new_[21604]_  = \new_[21603]_  & \new_[21600]_ ;
  assign \new_[21607]_  = ~A300 & A299;
  assign \new_[21610]_  = A302 & ~A301;
  assign \new_[21611]_  = \new_[21610]_  & \new_[21607]_ ;
  assign \new_[21612]_  = \new_[21611]_  & \new_[21604]_ ;
  assign \new_[21616]_  = A201 & A200;
  assign \new_[21617]_  = ~A199 & \new_[21616]_ ;
  assign \new_[21620]_  = A232 & A202;
  assign \new_[21623]_  = A234 & ~A233;
  assign \new_[21624]_  = \new_[21623]_  & \new_[21620]_ ;
  assign \new_[21625]_  = \new_[21624]_  & \new_[21617]_ ;
  assign \new_[21628]_  = ~A265 & A235;
  assign \new_[21631]_  = A298 & ~A266;
  assign \new_[21632]_  = \new_[21631]_  & \new_[21628]_ ;
  assign \new_[21635]_  = ~A300 & ~A299;
  assign \new_[21638]_  = A302 & ~A301;
  assign \new_[21639]_  = \new_[21638]_  & \new_[21635]_ ;
  assign \new_[21640]_  = \new_[21639]_  & \new_[21632]_ ;
  assign \new_[21644]_  = A201 & A200;
  assign \new_[21645]_  = ~A199 & \new_[21644]_ ;
  assign \new_[21648]_  = A232 & A202;
  assign \new_[21651]_  = A234 & ~A233;
  assign \new_[21652]_  = \new_[21651]_  & \new_[21648]_ ;
  assign \new_[21653]_  = \new_[21652]_  & \new_[21645]_ ;
  assign \new_[21656]_  = ~A265 & A235;
  assign \new_[21659]_  = ~A298 & ~A266;
  assign \new_[21660]_  = \new_[21659]_  & \new_[21656]_ ;
  assign \new_[21663]_  = ~A300 & A299;
  assign \new_[21666]_  = A302 & ~A301;
  assign \new_[21667]_  = \new_[21666]_  & \new_[21663]_ ;
  assign \new_[21668]_  = \new_[21667]_  & \new_[21660]_ ;
  assign \new_[21672]_  = A201 & A200;
  assign \new_[21673]_  = ~A199 & \new_[21672]_ ;
  assign \new_[21676]_  = A232 & A202;
  assign \new_[21679]_  = A234 & ~A233;
  assign \new_[21680]_  = \new_[21679]_  & \new_[21676]_ ;
  assign \new_[21681]_  = \new_[21680]_  & \new_[21673]_ ;
  assign \new_[21684]_  = A267 & ~A236;
  assign \new_[21687]_  = A269 & ~A268;
  assign \new_[21688]_  = \new_[21687]_  & \new_[21684]_ ;
  assign \new_[21691]_  = ~A299 & A298;
  assign \new_[21694]_  = A301 & A300;
  assign \new_[21695]_  = \new_[21694]_  & \new_[21691]_ ;
  assign \new_[21696]_  = \new_[21695]_  & \new_[21688]_ ;
  assign \new_[21700]_  = A201 & A200;
  assign \new_[21701]_  = ~A199 & \new_[21700]_ ;
  assign \new_[21704]_  = A232 & A202;
  assign \new_[21707]_  = A234 & ~A233;
  assign \new_[21708]_  = \new_[21707]_  & \new_[21704]_ ;
  assign \new_[21709]_  = \new_[21708]_  & \new_[21701]_ ;
  assign \new_[21712]_  = A267 & ~A236;
  assign \new_[21715]_  = A269 & ~A268;
  assign \new_[21716]_  = \new_[21715]_  & \new_[21712]_ ;
  assign \new_[21719]_  = ~A299 & A298;
  assign \new_[21722]_  = ~A302 & A300;
  assign \new_[21723]_  = \new_[21722]_  & \new_[21719]_ ;
  assign \new_[21724]_  = \new_[21723]_  & \new_[21716]_ ;
  assign \new_[21728]_  = A201 & A200;
  assign \new_[21729]_  = ~A199 & \new_[21728]_ ;
  assign \new_[21732]_  = A232 & A202;
  assign \new_[21735]_  = A234 & ~A233;
  assign \new_[21736]_  = \new_[21735]_  & \new_[21732]_ ;
  assign \new_[21737]_  = \new_[21736]_  & \new_[21729]_ ;
  assign \new_[21740]_  = A267 & ~A236;
  assign \new_[21743]_  = A269 & ~A268;
  assign \new_[21744]_  = \new_[21743]_  & \new_[21740]_ ;
  assign \new_[21747]_  = A299 & ~A298;
  assign \new_[21750]_  = A301 & A300;
  assign \new_[21751]_  = \new_[21750]_  & \new_[21747]_ ;
  assign \new_[21752]_  = \new_[21751]_  & \new_[21744]_ ;
  assign \new_[21756]_  = A201 & A200;
  assign \new_[21757]_  = ~A199 & \new_[21756]_ ;
  assign \new_[21760]_  = A232 & A202;
  assign \new_[21763]_  = A234 & ~A233;
  assign \new_[21764]_  = \new_[21763]_  & \new_[21760]_ ;
  assign \new_[21765]_  = \new_[21764]_  & \new_[21757]_ ;
  assign \new_[21768]_  = A267 & ~A236;
  assign \new_[21771]_  = A269 & ~A268;
  assign \new_[21772]_  = \new_[21771]_  & \new_[21768]_ ;
  assign \new_[21775]_  = A299 & ~A298;
  assign \new_[21778]_  = ~A302 & A300;
  assign \new_[21779]_  = \new_[21778]_  & \new_[21775]_ ;
  assign \new_[21780]_  = \new_[21779]_  & \new_[21772]_ ;
  assign \new_[21784]_  = A201 & A200;
  assign \new_[21785]_  = ~A199 & \new_[21784]_ ;
  assign \new_[21788]_  = A232 & A202;
  assign \new_[21791]_  = A234 & ~A233;
  assign \new_[21792]_  = \new_[21791]_  & \new_[21788]_ ;
  assign \new_[21793]_  = \new_[21792]_  & \new_[21785]_ ;
  assign \new_[21796]_  = ~A267 & ~A236;
  assign \new_[21799]_  = A298 & A268;
  assign \new_[21800]_  = \new_[21799]_  & \new_[21796]_ ;
  assign \new_[21803]_  = ~A300 & ~A299;
  assign \new_[21806]_  = A302 & ~A301;
  assign \new_[21807]_  = \new_[21806]_  & \new_[21803]_ ;
  assign \new_[21808]_  = \new_[21807]_  & \new_[21800]_ ;
  assign \new_[21812]_  = A201 & A200;
  assign \new_[21813]_  = ~A199 & \new_[21812]_ ;
  assign \new_[21816]_  = A232 & A202;
  assign \new_[21819]_  = A234 & ~A233;
  assign \new_[21820]_  = \new_[21819]_  & \new_[21816]_ ;
  assign \new_[21821]_  = \new_[21820]_  & \new_[21813]_ ;
  assign \new_[21824]_  = ~A267 & ~A236;
  assign \new_[21827]_  = ~A298 & A268;
  assign \new_[21828]_  = \new_[21827]_  & \new_[21824]_ ;
  assign \new_[21831]_  = ~A300 & A299;
  assign \new_[21834]_  = A302 & ~A301;
  assign \new_[21835]_  = \new_[21834]_  & \new_[21831]_ ;
  assign \new_[21836]_  = \new_[21835]_  & \new_[21828]_ ;
  assign \new_[21840]_  = A201 & A200;
  assign \new_[21841]_  = ~A199 & \new_[21840]_ ;
  assign \new_[21844]_  = A232 & A202;
  assign \new_[21847]_  = A234 & ~A233;
  assign \new_[21848]_  = \new_[21847]_  & \new_[21844]_ ;
  assign \new_[21849]_  = \new_[21848]_  & \new_[21841]_ ;
  assign \new_[21852]_  = ~A267 & ~A236;
  assign \new_[21855]_  = A298 & ~A269;
  assign \new_[21856]_  = \new_[21855]_  & \new_[21852]_ ;
  assign \new_[21859]_  = ~A300 & ~A299;
  assign \new_[21862]_  = A302 & ~A301;
  assign \new_[21863]_  = \new_[21862]_  & \new_[21859]_ ;
  assign \new_[21864]_  = \new_[21863]_  & \new_[21856]_ ;
  assign \new_[21868]_  = A201 & A200;
  assign \new_[21869]_  = ~A199 & \new_[21868]_ ;
  assign \new_[21872]_  = A232 & A202;
  assign \new_[21875]_  = A234 & ~A233;
  assign \new_[21876]_  = \new_[21875]_  & \new_[21872]_ ;
  assign \new_[21877]_  = \new_[21876]_  & \new_[21869]_ ;
  assign \new_[21880]_  = ~A267 & ~A236;
  assign \new_[21883]_  = ~A298 & ~A269;
  assign \new_[21884]_  = \new_[21883]_  & \new_[21880]_ ;
  assign \new_[21887]_  = ~A300 & A299;
  assign \new_[21890]_  = A302 & ~A301;
  assign \new_[21891]_  = \new_[21890]_  & \new_[21887]_ ;
  assign \new_[21892]_  = \new_[21891]_  & \new_[21884]_ ;
  assign \new_[21896]_  = A201 & A200;
  assign \new_[21897]_  = ~A199 & \new_[21896]_ ;
  assign \new_[21900]_  = A232 & A202;
  assign \new_[21903]_  = A234 & ~A233;
  assign \new_[21904]_  = \new_[21903]_  & \new_[21900]_ ;
  assign \new_[21905]_  = \new_[21904]_  & \new_[21897]_ ;
  assign \new_[21908]_  = A265 & ~A236;
  assign \new_[21911]_  = A298 & A266;
  assign \new_[21912]_  = \new_[21911]_  & \new_[21908]_ ;
  assign \new_[21915]_  = ~A300 & ~A299;
  assign \new_[21918]_  = A302 & ~A301;
  assign \new_[21919]_  = \new_[21918]_  & \new_[21915]_ ;
  assign \new_[21920]_  = \new_[21919]_  & \new_[21912]_ ;
  assign \new_[21924]_  = A201 & A200;
  assign \new_[21925]_  = ~A199 & \new_[21924]_ ;
  assign \new_[21928]_  = A232 & A202;
  assign \new_[21931]_  = A234 & ~A233;
  assign \new_[21932]_  = \new_[21931]_  & \new_[21928]_ ;
  assign \new_[21933]_  = \new_[21932]_  & \new_[21925]_ ;
  assign \new_[21936]_  = A265 & ~A236;
  assign \new_[21939]_  = ~A298 & A266;
  assign \new_[21940]_  = \new_[21939]_  & \new_[21936]_ ;
  assign \new_[21943]_  = ~A300 & A299;
  assign \new_[21946]_  = A302 & ~A301;
  assign \new_[21947]_  = \new_[21946]_  & \new_[21943]_ ;
  assign \new_[21948]_  = \new_[21947]_  & \new_[21940]_ ;
  assign \new_[21952]_  = A201 & A200;
  assign \new_[21953]_  = ~A199 & \new_[21952]_ ;
  assign \new_[21956]_  = A232 & A202;
  assign \new_[21959]_  = A234 & ~A233;
  assign \new_[21960]_  = \new_[21959]_  & \new_[21956]_ ;
  assign \new_[21961]_  = \new_[21960]_  & \new_[21953]_ ;
  assign \new_[21964]_  = ~A265 & ~A236;
  assign \new_[21967]_  = A298 & ~A266;
  assign \new_[21968]_  = \new_[21967]_  & \new_[21964]_ ;
  assign \new_[21971]_  = ~A300 & ~A299;
  assign \new_[21974]_  = A302 & ~A301;
  assign \new_[21975]_  = \new_[21974]_  & \new_[21971]_ ;
  assign \new_[21976]_  = \new_[21975]_  & \new_[21968]_ ;
  assign \new_[21980]_  = A201 & A200;
  assign \new_[21981]_  = ~A199 & \new_[21980]_ ;
  assign \new_[21984]_  = A232 & A202;
  assign \new_[21987]_  = A234 & ~A233;
  assign \new_[21988]_  = \new_[21987]_  & \new_[21984]_ ;
  assign \new_[21989]_  = \new_[21988]_  & \new_[21981]_ ;
  assign \new_[21992]_  = ~A265 & ~A236;
  assign \new_[21995]_  = ~A298 & ~A266;
  assign \new_[21996]_  = \new_[21995]_  & \new_[21992]_ ;
  assign \new_[21999]_  = ~A300 & A299;
  assign \new_[22002]_  = A302 & ~A301;
  assign \new_[22003]_  = \new_[22002]_  & \new_[21999]_ ;
  assign \new_[22004]_  = \new_[22003]_  & \new_[21996]_ ;
  assign \new_[22008]_  = A201 & A200;
  assign \new_[22009]_  = ~A199 & \new_[22008]_ ;
  assign \new_[22012]_  = A232 & A202;
  assign \new_[22015]_  = ~A234 & ~A233;
  assign \new_[22016]_  = \new_[22015]_  & \new_[22012]_ ;
  assign \new_[22017]_  = \new_[22016]_  & \new_[22009]_ ;
  assign \new_[22020]_  = A236 & ~A235;
  assign \new_[22023]_  = A268 & ~A267;
  assign \new_[22024]_  = \new_[22023]_  & \new_[22020]_ ;
  assign \new_[22027]_  = ~A299 & A298;
  assign \new_[22030]_  = A301 & A300;
  assign \new_[22031]_  = \new_[22030]_  & \new_[22027]_ ;
  assign \new_[22032]_  = \new_[22031]_  & \new_[22024]_ ;
  assign \new_[22036]_  = A201 & A200;
  assign \new_[22037]_  = ~A199 & \new_[22036]_ ;
  assign \new_[22040]_  = A232 & A202;
  assign \new_[22043]_  = ~A234 & ~A233;
  assign \new_[22044]_  = \new_[22043]_  & \new_[22040]_ ;
  assign \new_[22045]_  = \new_[22044]_  & \new_[22037]_ ;
  assign \new_[22048]_  = A236 & ~A235;
  assign \new_[22051]_  = A268 & ~A267;
  assign \new_[22052]_  = \new_[22051]_  & \new_[22048]_ ;
  assign \new_[22055]_  = ~A299 & A298;
  assign \new_[22058]_  = ~A302 & A300;
  assign \new_[22059]_  = \new_[22058]_  & \new_[22055]_ ;
  assign \new_[22060]_  = \new_[22059]_  & \new_[22052]_ ;
  assign \new_[22064]_  = A201 & A200;
  assign \new_[22065]_  = ~A199 & \new_[22064]_ ;
  assign \new_[22068]_  = A232 & A202;
  assign \new_[22071]_  = ~A234 & ~A233;
  assign \new_[22072]_  = \new_[22071]_  & \new_[22068]_ ;
  assign \new_[22073]_  = \new_[22072]_  & \new_[22065]_ ;
  assign \new_[22076]_  = A236 & ~A235;
  assign \new_[22079]_  = A268 & ~A267;
  assign \new_[22080]_  = \new_[22079]_  & \new_[22076]_ ;
  assign \new_[22083]_  = A299 & ~A298;
  assign \new_[22086]_  = A301 & A300;
  assign \new_[22087]_  = \new_[22086]_  & \new_[22083]_ ;
  assign \new_[22088]_  = \new_[22087]_  & \new_[22080]_ ;
  assign \new_[22092]_  = A201 & A200;
  assign \new_[22093]_  = ~A199 & \new_[22092]_ ;
  assign \new_[22096]_  = A232 & A202;
  assign \new_[22099]_  = ~A234 & ~A233;
  assign \new_[22100]_  = \new_[22099]_  & \new_[22096]_ ;
  assign \new_[22101]_  = \new_[22100]_  & \new_[22093]_ ;
  assign \new_[22104]_  = A236 & ~A235;
  assign \new_[22107]_  = A268 & ~A267;
  assign \new_[22108]_  = \new_[22107]_  & \new_[22104]_ ;
  assign \new_[22111]_  = A299 & ~A298;
  assign \new_[22114]_  = ~A302 & A300;
  assign \new_[22115]_  = \new_[22114]_  & \new_[22111]_ ;
  assign \new_[22116]_  = \new_[22115]_  & \new_[22108]_ ;
  assign \new_[22120]_  = A201 & A200;
  assign \new_[22121]_  = ~A199 & \new_[22120]_ ;
  assign \new_[22124]_  = A232 & A202;
  assign \new_[22127]_  = ~A234 & ~A233;
  assign \new_[22128]_  = \new_[22127]_  & \new_[22124]_ ;
  assign \new_[22129]_  = \new_[22128]_  & \new_[22121]_ ;
  assign \new_[22132]_  = A236 & ~A235;
  assign \new_[22135]_  = ~A269 & ~A267;
  assign \new_[22136]_  = \new_[22135]_  & \new_[22132]_ ;
  assign \new_[22139]_  = ~A299 & A298;
  assign \new_[22142]_  = A301 & A300;
  assign \new_[22143]_  = \new_[22142]_  & \new_[22139]_ ;
  assign \new_[22144]_  = \new_[22143]_  & \new_[22136]_ ;
  assign \new_[22148]_  = A201 & A200;
  assign \new_[22149]_  = ~A199 & \new_[22148]_ ;
  assign \new_[22152]_  = A232 & A202;
  assign \new_[22155]_  = ~A234 & ~A233;
  assign \new_[22156]_  = \new_[22155]_  & \new_[22152]_ ;
  assign \new_[22157]_  = \new_[22156]_  & \new_[22149]_ ;
  assign \new_[22160]_  = A236 & ~A235;
  assign \new_[22163]_  = ~A269 & ~A267;
  assign \new_[22164]_  = \new_[22163]_  & \new_[22160]_ ;
  assign \new_[22167]_  = ~A299 & A298;
  assign \new_[22170]_  = ~A302 & A300;
  assign \new_[22171]_  = \new_[22170]_  & \new_[22167]_ ;
  assign \new_[22172]_  = \new_[22171]_  & \new_[22164]_ ;
  assign \new_[22176]_  = A201 & A200;
  assign \new_[22177]_  = ~A199 & \new_[22176]_ ;
  assign \new_[22180]_  = A232 & A202;
  assign \new_[22183]_  = ~A234 & ~A233;
  assign \new_[22184]_  = \new_[22183]_  & \new_[22180]_ ;
  assign \new_[22185]_  = \new_[22184]_  & \new_[22177]_ ;
  assign \new_[22188]_  = A236 & ~A235;
  assign \new_[22191]_  = ~A269 & ~A267;
  assign \new_[22192]_  = \new_[22191]_  & \new_[22188]_ ;
  assign \new_[22195]_  = A299 & ~A298;
  assign \new_[22198]_  = A301 & A300;
  assign \new_[22199]_  = \new_[22198]_  & \new_[22195]_ ;
  assign \new_[22200]_  = \new_[22199]_  & \new_[22192]_ ;
  assign \new_[22204]_  = A201 & A200;
  assign \new_[22205]_  = ~A199 & \new_[22204]_ ;
  assign \new_[22208]_  = A232 & A202;
  assign \new_[22211]_  = ~A234 & ~A233;
  assign \new_[22212]_  = \new_[22211]_  & \new_[22208]_ ;
  assign \new_[22213]_  = \new_[22212]_  & \new_[22205]_ ;
  assign \new_[22216]_  = A236 & ~A235;
  assign \new_[22219]_  = ~A269 & ~A267;
  assign \new_[22220]_  = \new_[22219]_  & \new_[22216]_ ;
  assign \new_[22223]_  = A299 & ~A298;
  assign \new_[22226]_  = ~A302 & A300;
  assign \new_[22227]_  = \new_[22226]_  & \new_[22223]_ ;
  assign \new_[22228]_  = \new_[22227]_  & \new_[22220]_ ;
  assign \new_[22232]_  = A201 & A200;
  assign \new_[22233]_  = ~A199 & \new_[22232]_ ;
  assign \new_[22236]_  = A232 & A202;
  assign \new_[22239]_  = ~A234 & ~A233;
  assign \new_[22240]_  = \new_[22239]_  & \new_[22236]_ ;
  assign \new_[22241]_  = \new_[22240]_  & \new_[22233]_ ;
  assign \new_[22244]_  = A236 & ~A235;
  assign \new_[22247]_  = A266 & A265;
  assign \new_[22248]_  = \new_[22247]_  & \new_[22244]_ ;
  assign \new_[22251]_  = ~A299 & A298;
  assign \new_[22254]_  = A301 & A300;
  assign \new_[22255]_  = \new_[22254]_  & \new_[22251]_ ;
  assign \new_[22256]_  = \new_[22255]_  & \new_[22248]_ ;
  assign \new_[22260]_  = A201 & A200;
  assign \new_[22261]_  = ~A199 & \new_[22260]_ ;
  assign \new_[22264]_  = A232 & A202;
  assign \new_[22267]_  = ~A234 & ~A233;
  assign \new_[22268]_  = \new_[22267]_  & \new_[22264]_ ;
  assign \new_[22269]_  = \new_[22268]_  & \new_[22261]_ ;
  assign \new_[22272]_  = A236 & ~A235;
  assign \new_[22275]_  = A266 & A265;
  assign \new_[22276]_  = \new_[22275]_  & \new_[22272]_ ;
  assign \new_[22279]_  = ~A299 & A298;
  assign \new_[22282]_  = ~A302 & A300;
  assign \new_[22283]_  = \new_[22282]_  & \new_[22279]_ ;
  assign \new_[22284]_  = \new_[22283]_  & \new_[22276]_ ;
  assign \new_[22288]_  = A201 & A200;
  assign \new_[22289]_  = ~A199 & \new_[22288]_ ;
  assign \new_[22292]_  = A232 & A202;
  assign \new_[22295]_  = ~A234 & ~A233;
  assign \new_[22296]_  = \new_[22295]_  & \new_[22292]_ ;
  assign \new_[22297]_  = \new_[22296]_  & \new_[22289]_ ;
  assign \new_[22300]_  = A236 & ~A235;
  assign \new_[22303]_  = A266 & A265;
  assign \new_[22304]_  = \new_[22303]_  & \new_[22300]_ ;
  assign \new_[22307]_  = A299 & ~A298;
  assign \new_[22310]_  = A301 & A300;
  assign \new_[22311]_  = \new_[22310]_  & \new_[22307]_ ;
  assign \new_[22312]_  = \new_[22311]_  & \new_[22304]_ ;
  assign \new_[22316]_  = A201 & A200;
  assign \new_[22317]_  = ~A199 & \new_[22316]_ ;
  assign \new_[22320]_  = A232 & A202;
  assign \new_[22323]_  = ~A234 & ~A233;
  assign \new_[22324]_  = \new_[22323]_  & \new_[22320]_ ;
  assign \new_[22325]_  = \new_[22324]_  & \new_[22317]_ ;
  assign \new_[22328]_  = A236 & ~A235;
  assign \new_[22331]_  = A266 & A265;
  assign \new_[22332]_  = \new_[22331]_  & \new_[22328]_ ;
  assign \new_[22335]_  = A299 & ~A298;
  assign \new_[22338]_  = ~A302 & A300;
  assign \new_[22339]_  = \new_[22338]_  & \new_[22335]_ ;
  assign \new_[22340]_  = \new_[22339]_  & \new_[22332]_ ;
  assign \new_[22344]_  = A201 & A200;
  assign \new_[22345]_  = ~A199 & \new_[22344]_ ;
  assign \new_[22348]_  = A232 & A202;
  assign \new_[22351]_  = ~A234 & ~A233;
  assign \new_[22352]_  = \new_[22351]_  & \new_[22348]_ ;
  assign \new_[22353]_  = \new_[22352]_  & \new_[22345]_ ;
  assign \new_[22356]_  = A236 & ~A235;
  assign \new_[22359]_  = ~A266 & ~A265;
  assign \new_[22360]_  = \new_[22359]_  & \new_[22356]_ ;
  assign \new_[22363]_  = ~A299 & A298;
  assign \new_[22366]_  = A301 & A300;
  assign \new_[22367]_  = \new_[22366]_  & \new_[22363]_ ;
  assign \new_[22368]_  = \new_[22367]_  & \new_[22360]_ ;
  assign \new_[22372]_  = A201 & A200;
  assign \new_[22373]_  = ~A199 & \new_[22372]_ ;
  assign \new_[22376]_  = A232 & A202;
  assign \new_[22379]_  = ~A234 & ~A233;
  assign \new_[22380]_  = \new_[22379]_  & \new_[22376]_ ;
  assign \new_[22381]_  = \new_[22380]_  & \new_[22373]_ ;
  assign \new_[22384]_  = A236 & ~A235;
  assign \new_[22387]_  = ~A266 & ~A265;
  assign \new_[22388]_  = \new_[22387]_  & \new_[22384]_ ;
  assign \new_[22391]_  = ~A299 & A298;
  assign \new_[22394]_  = ~A302 & A300;
  assign \new_[22395]_  = \new_[22394]_  & \new_[22391]_ ;
  assign \new_[22396]_  = \new_[22395]_  & \new_[22388]_ ;
  assign \new_[22400]_  = A201 & A200;
  assign \new_[22401]_  = ~A199 & \new_[22400]_ ;
  assign \new_[22404]_  = A232 & A202;
  assign \new_[22407]_  = ~A234 & ~A233;
  assign \new_[22408]_  = \new_[22407]_  & \new_[22404]_ ;
  assign \new_[22409]_  = \new_[22408]_  & \new_[22401]_ ;
  assign \new_[22412]_  = A236 & ~A235;
  assign \new_[22415]_  = ~A266 & ~A265;
  assign \new_[22416]_  = \new_[22415]_  & \new_[22412]_ ;
  assign \new_[22419]_  = A299 & ~A298;
  assign \new_[22422]_  = A301 & A300;
  assign \new_[22423]_  = \new_[22422]_  & \new_[22419]_ ;
  assign \new_[22424]_  = \new_[22423]_  & \new_[22416]_ ;
  assign \new_[22428]_  = A201 & A200;
  assign \new_[22429]_  = ~A199 & \new_[22428]_ ;
  assign \new_[22432]_  = A232 & A202;
  assign \new_[22435]_  = ~A234 & ~A233;
  assign \new_[22436]_  = \new_[22435]_  & \new_[22432]_ ;
  assign \new_[22437]_  = \new_[22436]_  & \new_[22429]_ ;
  assign \new_[22440]_  = A236 & ~A235;
  assign \new_[22443]_  = ~A266 & ~A265;
  assign \new_[22444]_  = \new_[22443]_  & \new_[22440]_ ;
  assign \new_[22447]_  = A299 & ~A298;
  assign \new_[22450]_  = ~A302 & A300;
  assign \new_[22451]_  = \new_[22450]_  & \new_[22447]_ ;
  assign \new_[22452]_  = \new_[22451]_  & \new_[22444]_ ;
  assign \new_[22456]_  = A201 & A200;
  assign \new_[22457]_  = ~A199 & \new_[22456]_ ;
  assign \new_[22460]_  = ~A232 & ~A203;
  assign \new_[22463]_  = A234 & A233;
  assign \new_[22464]_  = \new_[22463]_  & \new_[22460]_ ;
  assign \new_[22465]_  = \new_[22464]_  & \new_[22457]_ ;
  assign \new_[22468]_  = A267 & A235;
  assign \new_[22471]_  = A269 & ~A268;
  assign \new_[22472]_  = \new_[22471]_  & \new_[22468]_ ;
  assign \new_[22475]_  = ~A299 & A298;
  assign \new_[22478]_  = A301 & A300;
  assign \new_[22479]_  = \new_[22478]_  & \new_[22475]_ ;
  assign \new_[22480]_  = \new_[22479]_  & \new_[22472]_ ;
  assign \new_[22484]_  = A201 & A200;
  assign \new_[22485]_  = ~A199 & \new_[22484]_ ;
  assign \new_[22488]_  = ~A232 & ~A203;
  assign \new_[22491]_  = A234 & A233;
  assign \new_[22492]_  = \new_[22491]_  & \new_[22488]_ ;
  assign \new_[22493]_  = \new_[22492]_  & \new_[22485]_ ;
  assign \new_[22496]_  = A267 & A235;
  assign \new_[22499]_  = A269 & ~A268;
  assign \new_[22500]_  = \new_[22499]_  & \new_[22496]_ ;
  assign \new_[22503]_  = ~A299 & A298;
  assign \new_[22506]_  = ~A302 & A300;
  assign \new_[22507]_  = \new_[22506]_  & \new_[22503]_ ;
  assign \new_[22508]_  = \new_[22507]_  & \new_[22500]_ ;
  assign \new_[22512]_  = A201 & A200;
  assign \new_[22513]_  = ~A199 & \new_[22512]_ ;
  assign \new_[22516]_  = ~A232 & ~A203;
  assign \new_[22519]_  = A234 & A233;
  assign \new_[22520]_  = \new_[22519]_  & \new_[22516]_ ;
  assign \new_[22521]_  = \new_[22520]_  & \new_[22513]_ ;
  assign \new_[22524]_  = A267 & A235;
  assign \new_[22527]_  = A269 & ~A268;
  assign \new_[22528]_  = \new_[22527]_  & \new_[22524]_ ;
  assign \new_[22531]_  = A299 & ~A298;
  assign \new_[22534]_  = A301 & A300;
  assign \new_[22535]_  = \new_[22534]_  & \new_[22531]_ ;
  assign \new_[22536]_  = \new_[22535]_  & \new_[22528]_ ;
  assign \new_[22540]_  = A201 & A200;
  assign \new_[22541]_  = ~A199 & \new_[22540]_ ;
  assign \new_[22544]_  = ~A232 & ~A203;
  assign \new_[22547]_  = A234 & A233;
  assign \new_[22548]_  = \new_[22547]_  & \new_[22544]_ ;
  assign \new_[22549]_  = \new_[22548]_  & \new_[22541]_ ;
  assign \new_[22552]_  = A267 & A235;
  assign \new_[22555]_  = A269 & ~A268;
  assign \new_[22556]_  = \new_[22555]_  & \new_[22552]_ ;
  assign \new_[22559]_  = A299 & ~A298;
  assign \new_[22562]_  = ~A302 & A300;
  assign \new_[22563]_  = \new_[22562]_  & \new_[22559]_ ;
  assign \new_[22564]_  = \new_[22563]_  & \new_[22556]_ ;
  assign \new_[22568]_  = A201 & A200;
  assign \new_[22569]_  = ~A199 & \new_[22568]_ ;
  assign \new_[22572]_  = ~A232 & ~A203;
  assign \new_[22575]_  = A234 & A233;
  assign \new_[22576]_  = \new_[22575]_  & \new_[22572]_ ;
  assign \new_[22577]_  = \new_[22576]_  & \new_[22569]_ ;
  assign \new_[22580]_  = ~A267 & A235;
  assign \new_[22583]_  = A298 & A268;
  assign \new_[22584]_  = \new_[22583]_  & \new_[22580]_ ;
  assign \new_[22587]_  = ~A300 & ~A299;
  assign \new_[22590]_  = A302 & ~A301;
  assign \new_[22591]_  = \new_[22590]_  & \new_[22587]_ ;
  assign \new_[22592]_  = \new_[22591]_  & \new_[22584]_ ;
  assign \new_[22596]_  = A201 & A200;
  assign \new_[22597]_  = ~A199 & \new_[22596]_ ;
  assign \new_[22600]_  = ~A232 & ~A203;
  assign \new_[22603]_  = A234 & A233;
  assign \new_[22604]_  = \new_[22603]_  & \new_[22600]_ ;
  assign \new_[22605]_  = \new_[22604]_  & \new_[22597]_ ;
  assign \new_[22608]_  = ~A267 & A235;
  assign \new_[22611]_  = ~A298 & A268;
  assign \new_[22612]_  = \new_[22611]_  & \new_[22608]_ ;
  assign \new_[22615]_  = ~A300 & A299;
  assign \new_[22618]_  = A302 & ~A301;
  assign \new_[22619]_  = \new_[22618]_  & \new_[22615]_ ;
  assign \new_[22620]_  = \new_[22619]_  & \new_[22612]_ ;
  assign \new_[22624]_  = A201 & A200;
  assign \new_[22625]_  = ~A199 & \new_[22624]_ ;
  assign \new_[22628]_  = ~A232 & ~A203;
  assign \new_[22631]_  = A234 & A233;
  assign \new_[22632]_  = \new_[22631]_  & \new_[22628]_ ;
  assign \new_[22633]_  = \new_[22632]_  & \new_[22625]_ ;
  assign \new_[22636]_  = ~A267 & A235;
  assign \new_[22639]_  = A298 & ~A269;
  assign \new_[22640]_  = \new_[22639]_  & \new_[22636]_ ;
  assign \new_[22643]_  = ~A300 & ~A299;
  assign \new_[22646]_  = A302 & ~A301;
  assign \new_[22647]_  = \new_[22646]_  & \new_[22643]_ ;
  assign \new_[22648]_  = \new_[22647]_  & \new_[22640]_ ;
  assign \new_[22652]_  = A201 & A200;
  assign \new_[22653]_  = ~A199 & \new_[22652]_ ;
  assign \new_[22656]_  = ~A232 & ~A203;
  assign \new_[22659]_  = A234 & A233;
  assign \new_[22660]_  = \new_[22659]_  & \new_[22656]_ ;
  assign \new_[22661]_  = \new_[22660]_  & \new_[22653]_ ;
  assign \new_[22664]_  = ~A267 & A235;
  assign \new_[22667]_  = ~A298 & ~A269;
  assign \new_[22668]_  = \new_[22667]_  & \new_[22664]_ ;
  assign \new_[22671]_  = ~A300 & A299;
  assign \new_[22674]_  = A302 & ~A301;
  assign \new_[22675]_  = \new_[22674]_  & \new_[22671]_ ;
  assign \new_[22676]_  = \new_[22675]_  & \new_[22668]_ ;
  assign \new_[22680]_  = A201 & A200;
  assign \new_[22681]_  = ~A199 & \new_[22680]_ ;
  assign \new_[22684]_  = ~A232 & ~A203;
  assign \new_[22687]_  = A234 & A233;
  assign \new_[22688]_  = \new_[22687]_  & \new_[22684]_ ;
  assign \new_[22689]_  = \new_[22688]_  & \new_[22681]_ ;
  assign \new_[22692]_  = A265 & A235;
  assign \new_[22695]_  = A298 & A266;
  assign \new_[22696]_  = \new_[22695]_  & \new_[22692]_ ;
  assign \new_[22699]_  = ~A300 & ~A299;
  assign \new_[22702]_  = A302 & ~A301;
  assign \new_[22703]_  = \new_[22702]_  & \new_[22699]_ ;
  assign \new_[22704]_  = \new_[22703]_  & \new_[22696]_ ;
  assign \new_[22708]_  = A201 & A200;
  assign \new_[22709]_  = ~A199 & \new_[22708]_ ;
  assign \new_[22712]_  = ~A232 & ~A203;
  assign \new_[22715]_  = A234 & A233;
  assign \new_[22716]_  = \new_[22715]_  & \new_[22712]_ ;
  assign \new_[22717]_  = \new_[22716]_  & \new_[22709]_ ;
  assign \new_[22720]_  = A265 & A235;
  assign \new_[22723]_  = ~A298 & A266;
  assign \new_[22724]_  = \new_[22723]_  & \new_[22720]_ ;
  assign \new_[22727]_  = ~A300 & A299;
  assign \new_[22730]_  = A302 & ~A301;
  assign \new_[22731]_  = \new_[22730]_  & \new_[22727]_ ;
  assign \new_[22732]_  = \new_[22731]_  & \new_[22724]_ ;
  assign \new_[22736]_  = A201 & A200;
  assign \new_[22737]_  = ~A199 & \new_[22736]_ ;
  assign \new_[22740]_  = ~A232 & ~A203;
  assign \new_[22743]_  = A234 & A233;
  assign \new_[22744]_  = \new_[22743]_  & \new_[22740]_ ;
  assign \new_[22745]_  = \new_[22744]_  & \new_[22737]_ ;
  assign \new_[22748]_  = ~A265 & A235;
  assign \new_[22751]_  = A298 & ~A266;
  assign \new_[22752]_  = \new_[22751]_  & \new_[22748]_ ;
  assign \new_[22755]_  = ~A300 & ~A299;
  assign \new_[22758]_  = A302 & ~A301;
  assign \new_[22759]_  = \new_[22758]_  & \new_[22755]_ ;
  assign \new_[22760]_  = \new_[22759]_  & \new_[22752]_ ;
  assign \new_[22764]_  = A201 & A200;
  assign \new_[22765]_  = ~A199 & \new_[22764]_ ;
  assign \new_[22768]_  = ~A232 & ~A203;
  assign \new_[22771]_  = A234 & A233;
  assign \new_[22772]_  = \new_[22771]_  & \new_[22768]_ ;
  assign \new_[22773]_  = \new_[22772]_  & \new_[22765]_ ;
  assign \new_[22776]_  = ~A265 & A235;
  assign \new_[22779]_  = ~A298 & ~A266;
  assign \new_[22780]_  = \new_[22779]_  & \new_[22776]_ ;
  assign \new_[22783]_  = ~A300 & A299;
  assign \new_[22786]_  = A302 & ~A301;
  assign \new_[22787]_  = \new_[22786]_  & \new_[22783]_ ;
  assign \new_[22788]_  = \new_[22787]_  & \new_[22780]_ ;
  assign \new_[22792]_  = A201 & A200;
  assign \new_[22793]_  = ~A199 & \new_[22792]_ ;
  assign \new_[22796]_  = ~A232 & ~A203;
  assign \new_[22799]_  = A234 & A233;
  assign \new_[22800]_  = \new_[22799]_  & \new_[22796]_ ;
  assign \new_[22801]_  = \new_[22800]_  & \new_[22793]_ ;
  assign \new_[22804]_  = A267 & ~A236;
  assign \new_[22807]_  = A269 & ~A268;
  assign \new_[22808]_  = \new_[22807]_  & \new_[22804]_ ;
  assign \new_[22811]_  = ~A299 & A298;
  assign \new_[22814]_  = A301 & A300;
  assign \new_[22815]_  = \new_[22814]_  & \new_[22811]_ ;
  assign \new_[22816]_  = \new_[22815]_  & \new_[22808]_ ;
  assign \new_[22820]_  = A201 & A200;
  assign \new_[22821]_  = ~A199 & \new_[22820]_ ;
  assign \new_[22824]_  = ~A232 & ~A203;
  assign \new_[22827]_  = A234 & A233;
  assign \new_[22828]_  = \new_[22827]_  & \new_[22824]_ ;
  assign \new_[22829]_  = \new_[22828]_  & \new_[22821]_ ;
  assign \new_[22832]_  = A267 & ~A236;
  assign \new_[22835]_  = A269 & ~A268;
  assign \new_[22836]_  = \new_[22835]_  & \new_[22832]_ ;
  assign \new_[22839]_  = ~A299 & A298;
  assign \new_[22842]_  = ~A302 & A300;
  assign \new_[22843]_  = \new_[22842]_  & \new_[22839]_ ;
  assign \new_[22844]_  = \new_[22843]_  & \new_[22836]_ ;
  assign \new_[22848]_  = A201 & A200;
  assign \new_[22849]_  = ~A199 & \new_[22848]_ ;
  assign \new_[22852]_  = ~A232 & ~A203;
  assign \new_[22855]_  = A234 & A233;
  assign \new_[22856]_  = \new_[22855]_  & \new_[22852]_ ;
  assign \new_[22857]_  = \new_[22856]_  & \new_[22849]_ ;
  assign \new_[22860]_  = A267 & ~A236;
  assign \new_[22863]_  = A269 & ~A268;
  assign \new_[22864]_  = \new_[22863]_  & \new_[22860]_ ;
  assign \new_[22867]_  = A299 & ~A298;
  assign \new_[22870]_  = A301 & A300;
  assign \new_[22871]_  = \new_[22870]_  & \new_[22867]_ ;
  assign \new_[22872]_  = \new_[22871]_  & \new_[22864]_ ;
  assign \new_[22876]_  = A201 & A200;
  assign \new_[22877]_  = ~A199 & \new_[22876]_ ;
  assign \new_[22880]_  = ~A232 & ~A203;
  assign \new_[22883]_  = A234 & A233;
  assign \new_[22884]_  = \new_[22883]_  & \new_[22880]_ ;
  assign \new_[22885]_  = \new_[22884]_  & \new_[22877]_ ;
  assign \new_[22888]_  = A267 & ~A236;
  assign \new_[22891]_  = A269 & ~A268;
  assign \new_[22892]_  = \new_[22891]_  & \new_[22888]_ ;
  assign \new_[22895]_  = A299 & ~A298;
  assign \new_[22898]_  = ~A302 & A300;
  assign \new_[22899]_  = \new_[22898]_  & \new_[22895]_ ;
  assign \new_[22900]_  = \new_[22899]_  & \new_[22892]_ ;
  assign \new_[22904]_  = A201 & A200;
  assign \new_[22905]_  = ~A199 & \new_[22904]_ ;
  assign \new_[22908]_  = ~A232 & ~A203;
  assign \new_[22911]_  = A234 & A233;
  assign \new_[22912]_  = \new_[22911]_  & \new_[22908]_ ;
  assign \new_[22913]_  = \new_[22912]_  & \new_[22905]_ ;
  assign \new_[22916]_  = ~A267 & ~A236;
  assign \new_[22919]_  = A298 & A268;
  assign \new_[22920]_  = \new_[22919]_  & \new_[22916]_ ;
  assign \new_[22923]_  = ~A300 & ~A299;
  assign \new_[22926]_  = A302 & ~A301;
  assign \new_[22927]_  = \new_[22926]_  & \new_[22923]_ ;
  assign \new_[22928]_  = \new_[22927]_  & \new_[22920]_ ;
  assign \new_[22932]_  = A201 & A200;
  assign \new_[22933]_  = ~A199 & \new_[22932]_ ;
  assign \new_[22936]_  = ~A232 & ~A203;
  assign \new_[22939]_  = A234 & A233;
  assign \new_[22940]_  = \new_[22939]_  & \new_[22936]_ ;
  assign \new_[22941]_  = \new_[22940]_  & \new_[22933]_ ;
  assign \new_[22944]_  = ~A267 & ~A236;
  assign \new_[22947]_  = ~A298 & A268;
  assign \new_[22948]_  = \new_[22947]_  & \new_[22944]_ ;
  assign \new_[22951]_  = ~A300 & A299;
  assign \new_[22954]_  = A302 & ~A301;
  assign \new_[22955]_  = \new_[22954]_  & \new_[22951]_ ;
  assign \new_[22956]_  = \new_[22955]_  & \new_[22948]_ ;
  assign \new_[22960]_  = A201 & A200;
  assign \new_[22961]_  = ~A199 & \new_[22960]_ ;
  assign \new_[22964]_  = ~A232 & ~A203;
  assign \new_[22967]_  = A234 & A233;
  assign \new_[22968]_  = \new_[22967]_  & \new_[22964]_ ;
  assign \new_[22969]_  = \new_[22968]_  & \new_[22961]_ ;
  assign \new_[22972]_  = ~A267 & ~A236;
  assign \new_[22975]_  = A298 & ~A269;
  assign \new_[22976]_  = \new_[22975]_  & \new_[22972]_ ;
  assign \new_[22979]_  = ~A300 & ~A299;
  assign \new_[22982]_  = A302 & ~A301;
  assign \new_[22983]_  = \new_[22982]_  & \new_[22979]_ ;
  assign \new_[22984]_  = \new_[22983]_  & \new_[22976]_ ;
  assign \new_[22988]_  = A201 & A200;
  assign \new_[22989]_  = ~A199 & \new_[22988]_ ;
  assign \new_[22992]_  = ~A232 & ~A203;
  assign \new_[22995]_  = A234 & A233;
  assign \new_[22996]_  = \new_[22995]_  & \new_[22992]_ ;
  assign \new_[22997]_  = \new_[22996]_  & \new_[22989]_ ;
  assign \new_[23000]_  = ~A267 & ~A236;
  assign \new_[23003]_  = ~A298 & ~A269;
  assign \new_[23004]_  = \new_[23003]_  & \new_[23000]_ ;
  assign \new_[23007]_  = ~A300 & A299;
  assign \new_[23010]_  = A302 & ~A301;
  assign \new_[23011]_  = \new_[23010]_  & \new_[23007]_ ;
  assign \new_[23012]_  = \new_[23011]_  & \new_[23004]_ ;
  assign \new_[23016]_  = A201 & A200;
  assign \new_[23017]_  = ~A199 & \new_[23016]_ ;
  assign \new_[23020]_  = ~A232 & ~A203;
  assign \new_[23023]_  = A234 & A233;
  assign \new_[23024]_  = \new_[23023]_  & \new_[23020]_ ;
  assign \new_[23025]_  = \new_[23024]_  & \new_[23017]_ ;
  assign \new_[23028]_  = A265 & ~A236;
  assign \new_[23031]_  = A298 & A266;
  assign \new_[23032]_  = \new_[23031]_  & \new_[23028]_ ;
  assign \new_[23035]_  = ~A300 & ~A299;
  assign \new_[23038]_  = A302 & ~A301;
  assign \new_[23039]_  = \new_[23038]_  & \new_[23035]_ ;
  assign \new_[23040]_  = \new_[23039]_  & \new_[23032]_ ;
  assign \new_[23044]_  = A201 & A200;
  assign \new_[23045]_  = ~A199 & \new_[23044]_ ;
  assign \new_[23048]_  = ~A232 & ~A203;
  assign \new_[23051]_  = A234 & A233;
  assign \new_[23052]_  = \new_[23051]_  & \new_[23048]_ ;
  assign \new_[23053]_  = \new_[23052]_  & \new_[23045]_ ;
  assign \new_[23056]_  = A265 & ~A236;
  assign \new_[23059]_  = ~A298 & A266;
  assign \new_[23060]_  = \new_[23059]_  & \new_[23056]_ ;
  assign \new_[23063]_  = ~A300 & A299;
  assign \new_[23066]_  = A302 & ~A301;
  assign \new_[23067]_  = \new_[23066]_  & \new_[23063]_ ;
  assign \new_[23068]_  = \new_[23067]_  & \new_[23060]_ ;
  assign \new_[23072]_  = A201 & A200;
  assign \new_[23073]_  = ~A199 & \new_[23072]_ ;
  assign \new_[23076]_  = ~A232 & ~A203;
  assign \new_[23079]_  = A234 & A233;
  assign \new_[23080]_  = \new_[23079]_  & \new_[23076]_ ;
  assign \new_[23081]_  = \new_[23080]_  & \new_[23073]_ ;
  assign \new_[23084]_  = ~A265 & ~A236;
  assign \new_[23087]_  = A298 & ~A266;
  assign \new_[23088]_  = \new_[23087]_  & \new_[23084]_ ;
  assign \new_[23091]_  = ~A300 & ~A299;
  assign \new_[23094]_  = A302 & ~A301;
  assign \new_[23095]_  = \new_[23094]_  & \new_[23091]_ ;
  assign \new_[23096]_  = \new_[23095]_  & \new_[23088]_ ;
  assign \new_[23100]_  = A201 & A200;
  assign \new_[23101]_  = ~A199 & \new_[23100]_ ;
  assign \new_[23104]_  = ~A232 & ~A203;
  assign \new_[23107]_  = A234 & A233;
  assign \new_[23108]_  = \new_[23107]_  & \new_[23104]_ ;
  assign \new_[23109]_  = \new_[23108]_  & \new_[23101]_ ;
  assign \new_[23112]_  = ~A265 & ~A236;
  assign \new_[23115]_  = ~A298 & ~A266;
  assign \new_[23116]_  = \new_[23115]_  & \new_[23112]_ ;
  assign \new_[23119]_  = ~A300 & A299;
  assign \new_[23122]_  = A302 & ~A301;
  assign \new_[23123]_  = \new_[23122]_  & \new_[23119]_ ;
  assign \new_[23124]_  = \new_[23123]_  & \new_[23116]_ ;
  assign \new_[23128]_  = A201 & A200;
  assign \new_[23129]_  = ~A199 & \new_[23128]_ ;
  assign \new_[23132]_  = ~A232 & ~A203;
  assign \new_[23135]_  = ~A234 & A233;
  assign \new_[23136]_  = \new_[23135]_  & \new_[23132]_ ;
  assign \new_[23137]_  = \new_[23136]_  & \new_[23129]_ ;
  assign \new_[23140]_  = A236 & ~A235;
  assign \new_[23143]_  = A268 & ~A267;
  assign \new_[23144]_  = \new_[23143]_  & \new_[23140]_ ;
  assign \new_[23147]_  = ~A299 & A298;
  assign \new_[23150]_  = A301 & A300;
  assign \new_[23151]_  = \new_[23150]_  & \new_[23147]_ ;
  assign \new_[23152]_  = \new_[23151]_  & \new_[23144]_ ;
  assign \new_[23156]_  = A201 & A200;
  assign \new_[23157]_  = ~A199 & \new_[23156]_ ;
  assign \new_[23160]_  = ~A232 & ~A203;
  assign \new_[23163]_  = ~A234 & A233;
  assign \new_[23164]_  = \new_[23163]_  & \new_[23160]_ ;
  assign \new_[23165]_  = \new_[23164]_  & \new_[23157]_ ;
  assign \new_[23168]_  = A236 & ~A235;
  assign \new_[23171]_  = A268 & ~A267;
  assign \new_[23172]_  = \new_[23171]_  & \new_[23168]_ ;
  assign \new_[23175]_  = ~A299 & A298;
  assign \new_[23178]_  = ~A302 & A300;
  assign \new_[23179]_  = \new_[23178]_  & \new_[23175]_ ;
  assign \new_[23180]_  = \new_[23179]_  & \new_[23172]_ ;
  assign \new_[23184]_  = A201 & A200;
  assign \new_[23185]_  = ~A199 & \new_[23184]_ ;
  assign \new_[23188]_  = ~A232 & ~A203;
  assign \new_[23191]_  = ~A234 & A233;
  assign \new_[23192]_  = \new_[23191]_  & \new_[23188]_ ;
  assign \new_[23193]_  = \new_[23192]_  & \new_[23185]_ ;
  assign \new_[23196]_  = A236 & ~A235;
  assign \new_[23199]_  = A268 & ~A267;
  assign \new_[23200]_  = \new_[23199]_  & \new_[23196]_ ;
  assign \new_[23203]_  = A299 & ~A298;
  assign \new_[23206]_  = A301 & A300;
  assign \new_[23207]_  = \new_[23206]_  & \new_[23203]_ ;
  assign \new_[23208]_  = \new_[23207]_  & \new_[23200]_ ;
  assign \new_[23212]_  = A201 & A200;
  assign \new_[23213]_  = ~A199 & \new_[23212]_ ;
  assign \new_[23216]_  = ~A232 & ~A203;
  assign \new_[23219]_  = ~A234 & A233;
  assign \new_[23220]_  = \new_[23219]_  & \new_[23216]_ ;
  assign \new_[23221]_  = \new_[23220]_  & \new_[23213]_ ;
  assign \new_[23224]_  = A236 & ~A235;
  assign \new_[23227]_  = A268 & ~A267;
  assign \new_[23228]_  = \new_[23227]_  & \new_[23224]_ ;
  assign \new_[23231]_  = A299 & ~A298;
  assign \new_[23234]_  = ~A302 & A300;
  assign \new_[23235]_  = \new_[23234]_  & \new_[23231]_ ;
  assign \new_[23236]_  = \new_[23235]_  & \new_[23228]_ ;
  assign \new_[23240]_  = A201 & A200;
  assign \new_[23241]_  = ~A199 & \new_[23240]_ ;
  assign \new_[23244]_  = ~A232 & ~A203;
  assign \new_[23247]_  = ~A234 & A233;
  assign \new_[23248]_  = \new_[23247]_  & \new_[23244]_ ;
  assign \new_[23249]_  = \new_[23248]_  & \new_[23241]_ ;
  assign \new_[23252]_  = A236 & ~A235;
  assign \new_[23255]_  = ~A269 & ~A267;
  assign \new_[23256]_  = \new_[23255]_  & \new_[23252]_ ;
  assign \new_[23259]_  = ~A299 & A298;
  assign \new_[23262]_  = A301 & A300;
  assign \new_[23263]_  = \new_[23262]_  & \new_[23259]_ ;
  assign \new_[23264]_  = \new_[23263]_  & \new_[23256]_ ;
  assign \new_[23268]_  = A201 & A200;
  assign \new_[23269]_  = ~A199 & \new_[23268]_ ;
  assign \new_[23272]_  = ~A232 & ~A203;
  assign \new_[23275]_  = ~A234 & A233;
  assign \new_[23276]_  = \new_[23275]_  & \new_[23272]_ ;
  assign \new_[23277]_  = \new_[23276]_  & \new_[23269]_ ;
  assign \new_[23280]_  = A236 & ~A235;
  assign \new_[23283]_  = ~A269 & ~A267;
  assign \new_[23284]_  = \new_[23283]_  & \new_[23280]_ ;
  assign \new_[23287]_  = ~A299 & A298;
  assign \new_[23290]_  = ~A302 & A300;
  assign \new_[23291]_  = \new_[23290]_  & \new_[23287]_ ;
  assign \new_[23292]_  = \new_[23291]_  & \new_[23284]_ ;
  assign \new_[23296]_  = A201 & A200;
  assign \new_[23297]_  = ~A199 & \new_[23296]_ ;
  assign \new_[23300]_  = ~A232 & ~A203;
  assign \new_[23303]_  = ~A234 & A233;
  assign \new_[23304]_  = \new_[23303]_  & \new_[23300]_ ;
  assign \new_[23305]_  = \new_[23304]_  & \new_[23297]_ ;
  assign \new_[23308]_  = A236 & ~A235;
  assign \new_[23311]_  = ~A269 & ~A267;
  assign \new_[23312]_  = \new_[23311]_  & \new_[23308]_ ;
  assign \new_[23315]_  = A299 & ~A298;
  assign \new_[23318]_  = A301 & A300;
  assign \new_[23319]_  = \new_[23318]_  & \new_[23315]_ ;
  assign \new_[23320]_  = \new_[23319]_  & \new_[23312]_ ;
  assign \new_[23324]_  = A201 & A200;
  assign \new_[23325]_  = ~A199 & \new_[23324]_ ;
  assign \new_[23328]_  = ~A232 & ~A203;
  assign \new_[23331]_  = ~A234 & A233;
  assign \new_[23332]_  = \new_[23331]_  & \new_[23328]_ ;
  assign \new_[23333]_  = \new_[23332]_  & \new_[23325]_ ;
  assign \new_[23336]_  = A236 & ~A235;
  assign \new_[23339]_  = ~A269 & ~A267;
  assign \new_[23340]_  = \new_[23339]_  & \new_[23336]_ ;
  assign \new_[23343]_  = A299 & ~A298;
  assign \new_[23346]_  = ~A302 & A300;
  assign \new_[23347]_  = \new_[23346]_  & \new_[23343]_ ;
  assign \new_[23348]_  = \new_[23347]_  & \new_[23340]_ ;
  assign \new_[23352]_  = A201 & A200;
  assign \new_[23353]_  = ~A199 & \new_[23352]_ ;
  assign \new_[23356]_  = ~A232 & ~A203;
  assign \new_[23359]_  = ~A234 & A233;
  assign \new_[23360]_  = \new_[23359]_  & \new_[23356]_ ;
  assign \new_[23361]_  = \new_[23360]_  & \new_[23353]_ ;
  assign \new_[23364]_  = A236 & ~A235;
  assign \new_[23367]_  = A266 & A265;
  assign \new_[23368]_  = \new_[23367]_  & \new_[23364]_ ;
  assign \new_[23371]_  = ~A299 & A298;
  assign \new_[23374]_  = A301 & A300;
  assign \new_[23375]_  = \new_[23374]_  & \new_[23371]_ ;
  assign \new_[23376]_  = \new_[23375]_  & \new_[23368]_ ;
  assign \new_[23380]_  = A201 & A200;
  assign \new_[23381]_  = ~A199 & \new_[23380]_ ;
  assign \new_[23384]_  = ~A232 & ~A203;
  assign \new_[23387]_  = ~A234 & A233;
  assign \new_[23388]_  = \new_[23387]_  & \new_[23384]_ ;
  assign \new_[23389]_  = \new_[23388]_  & \new_[23381]_ ;
  assign \new_[23392]_  = A236 & ~A235;
  assign \new_[23395]_  = A266 & A265;
  assign \new_[23396]_  = \new_[23395]_  & \new_[23392]_ ;
  assign \new_[23399]_  = ~A299 & A298;
  assign \new_[23402]_  = ~A302 & A300;
  assign \new_[23403]_  = \new_[23402]_  & \new_[23399]_ ;
  assign \new_[23404]_  = \new_[23403]_  & \new_[23396]_ ;
  assign \new_[23408]_  = A201 & A200;
  assign \new_[23409]_  = ~A199 & \new_[23408]_ ;
  assign \new_[23412]_  = ~A232 & ~A203;
  assign \new_[23415]_  = ~A234 & A233;
  assign \new_[23416]_  = \new_[23415]_  & \new_[23412]_ ;
  assign \new_[23417]_  = \new_[23416]_  & \new_[23409]_ ;
  assign \new_[23420]_  = A236 & ~A235;
  assign \new_[23423]_  = A266 & A265;
  assign \new_[23424]_  = \new_[23423]_  & \new_[23420]_ ;
  assign \new_[23427]_  = A299 & ~A298;
  assign \new_[23430]_  = A301 & A300;
  assign \new_[23431]_  = \new_[23430]_  & \new_[23427]_ ;
  assign \new_[23432]_  = \new_[23431]_  & \new_[23424]_ ;
  assign \new_[23436]_  = A201 & A200;
  assign \new_[23437]_  = ~A199 & \new_[23436]_ ;
  assign \new_[23440]_  = ~A232 & ~A203;
  assign \new_[23443]_  = ~A234 & A233;
  assign \new_[23444]_  = \new_[23443]_  & \new_[23440]_ ;
  assign \new_[23445]_  = \new_[23444]_  & \new_[23437]_ ;
  assign \new_[23448]_  = A236 & ~A235;
  assign \new_[23451]_  = A266 & A265;
  assign \new_[23452]_  = \new_[23451]_  & \new_[23448]_ ;
  assign \new_[23455]_  = A299 & ~A298;
  assign \new_[23458]_  = ~A302 & A300;
  assign \new_[23459]_  = \new_[23458]_  & \new_[23455]_ ;
  assign \new_[23460]_  = \new_[23459]_  & \new_[23452]_ ;
  assign \new_[23464]_  = A201 & A200;
  assign \new_[23465]_  = ~A199 & \new_[23464]_ ;
  assign \new_[23468]_  = ~A232 & ~A203;
  assign \new_[23471]_  = ~A234 & A233;
  assign \new_[23472]_  = \new_[23471]_  & \new_[23468]_ ;
  assign \new_[23473]_  = \new_[23472]_  & \new_[23465]_ ;
  assign \new_[23476]_  = A236 & ~A235;
  assign \new_[23479]_  = ~A266 & ~A265;
  assign \new_[23480]_  = \new_[23479]_  & \new_[23476]_ ;
  assign \new_[23483]_  = ~A299 & A298;
  assign \new_[23486]_  = A301 & A300;
  assign \new_[23487]_  = \new_[23486]_  & \new_[23483]_ ;
  assign \new_[23488]_  = \new_[23487]_  & \new_[23480]_ ;
  assign \new_[23492]_  = A201 & A200;
  assign \new_[23493]_  = ~A199 & \new_[23492]_ ;
  assign \new_[23496]_  = ~A232 & ~A203;
  assign \new_[23499]_  = ~A234 & A233;
  assign \new_[23500]_  = \new_[23499]_  & \new_[23496]_ ;
  assign \new_[23501]_  = \new_[23500]_  & \new_[23493]_ ;
  assign \new_[23504]_  = A236 & ~A235;
  assign \new_[23507]_  = ~A266 & ~A265;
  assign \new_[23508]_  = \new_[23507]_  & \new_[23504]_ ;
  assign \new_[23511]_  = ~A299 & A298;
  assign \new_[23514]_  = ~A302 & A300;
  assign \new_[23515]_  = \new_[23514]_  & \new_[23511]_ ;
  assign \new_[23516]_  = \new_[23515]_  & \new_[23508]_ ;
  assign \new_[23520]_  = A201 & A200;
  assign \new_[23521]_  = ~A199 & \new_[23520]_ ;
  assign \new_[23524]_  = ~A232 & ~A203;
  assign \new_[23527]_  = ~A234 & A233;
  assign \new_[23528]_  = \new_[23527]_  & \new_[23524]_ ;
  assign \new_[23529]_  = \new_[23528]_  & \new_[23521]_ ;
  assign \new_[23532]_  = A236 & ~A235;
  assign \new_[23535]_  = ~A266 & ~A265;
  assign \new_[23536]_  = \new_[23535]_  & \new_[23532]_ ;
  assign \new_[23539]_  = A299 & ~A298;
  assign \new_[23542]_  = A301 & A300;
  assign \new_[23543]_  = \new_[23542]_  & \new_[23539]_ ;
  assign \new_[23544]_  = \new_[23543]_  & \new_[23536]_ ;
  assign \new_[23548]_  = A201 & A200;
  assign \new_[23549]_  = ~A199 & \new_[23548]_ ;
  assign \new_[23552]_  = ~A232 & ~A203;
  assign \new_[23555]_  = ~A234 & A233;
  assign \new_[23556]_  = \new_[23555]_  & \new_[23552]_ ;
  assign \new_[23557]_  = \new_[23556]_  & \new_[23549]_ ;
  assign \new_[23560]_  = A236 & ~A235;
  assign \new_[23563]_  = ~A266 & ~A265;
  assign \new_[23564]_  = \new_[23563]_  & \new_[23560]_ ;
  assign \new_[23567]_  = A299 & ~A298;
  assign \new_[23570]_  = ~A302 & A300;
  assign \new_[23571]_  = \new_[23570]_  & \new_[23567]_ ;
  assign \new_[23572]_  = \new_[23571]_  & \new_[23564]_ ;
  assign \new_[23576]_  = A201 & A200;
  assign \new_[23577]_  = ~A199 & \new_[23576]_ ;
  assign \new_[23580]_  = A232 & ~A203;
  assign \new_[23583]_  = A234 & ~A233;
  assign \new_[23584]_  = \new_[23583]_  & \new_[23580]_ ;
  assign \new_[23585]_  = \new_[23584]_  & \new_[23577]_ ;
  assign \new_[23588]_  = A267 & A235;
  assign \new_[23591]_  = A269 & ~A268;
  assign \new_[23592]_  = \new_[23591]_  & \new_[23588]_ ;
  assign \new_[23595]_  = ~A299 & A298;
  assign \new_[23598]_  = A301 & A300;
  assign \new_[23599]_  = \new_[23598]_  & \new_[23595]_ ;
  assign \new_[23600]_  = \new_[23599]_  & \new_[23592]_ ;
  assign \new_[23604]_  = A201 & A200;
  assign \new_[23605]_  = ~A199 & \new_[23604]_ ;
  assign \new_[23608]_  = A232 & ~A203;
  assign \new_[23611]_  = A234 & ~A233;
  assign \new_[23612]_  = \new_[23611]_  & \new_[23608]_ ;
  assign \new_[23613]_  = \new_[23612]_  & \new_[23605]_ ;
  assign \new_[23616]_  = A267 & A235;
  assign \new_[23619]_  = A269 & ~A268;
  assign \new_[23620]_  = \new_[23619]_  & \new_[23616]_ ;
  assign \new_[23623]_  = ~A299 & A298;
  assign \new_[23626]_  = ~A302 & A300;
  assign \new_[23627]_  = \new_[23626]_  & \new_[23623]_ ;
  assign \new_[23628]_  = \new_[23627]_  & \new_[23620]_ ;
  assign \new_[23632]_  = A201 & A200;
  assign \new_[23633]_  = ~A199 & \new_[23632]_ ;
  assign \new_[23636]_  = A232 & ~A203;
  assign \new_[23639]_  = A234 & ~A233;
  assign \new_[23640]_  = \new_[23639]_  & \new_[23636]_ ;
  assign \new_[23641]_  = \new_[23640]_  & \new_[23633]_ ;
  assign \new_[23644]_  = A267 & A235;
  assign \new_[23647]_  = A269 & ~A268;
  assign \new_[23648]_  = \new_[23647]_  & \new_[23644]_ ;
  assign \new_[23651]_  = A299 & ~A298;
  assign \new_[23654]_  = A301 & A300;
  assign \new_[23655]_  = \new_[23654]_  & \new_[23651]_ ;
  assign \new_[23656]_  = \new_[23655]_  & \new_[23648]_ ;
  assign \new_[23660]_  = A201 & A200;
  assign \new_[23661]_  = ~A199 & \new_[23660]_ ;
  assign \new_[23664]_  = A232 & ~A203;
  assign \new_[23667]_  = A234 & ~A233;
  assign \new_[23668]_  = \new_[23667]_  & \new_[23664]_ ;
  assign \new_[23669]_  = \new_[23668]_  & \new_[23661]_ ;
  assign \new_[23672]_  = A267 & A235;
  assign \new_[23675]_  = A269 & ~A268;
  assign \new_[23676]_  = \new_[23675]_  & \new_[23672]_ ;
  assign \new_[23679]_  = A299 & ~A298;
  assign \new_[23682]_  = ~A302 & A300;
  assign \new_[23683]_  = \new_[23682]_  & \new_[23679]_ ;
  assign \new_[23684]_  = \new_[23683]_  & \new_[23676]_ ;
  assign \new_[23688]_  = A201 & A200;
  assign \new_[23689]_  = ~A199 & \new_[23688]_ ;
  assign \new_[23692]_  = A232 & ~A203;
  assign \new_[23695]_  = A234 & ~A233;
  assign \new_[23696]_  = \new_[23695]_  & \new_[23692]_ ;
  assign \new_[23697]_  = \new_[23696]_  & \new_[23689]_ ;
  assign \new_[23700]_  = ~A267 & A235;
  assign \new_[23703]_  = A298 & A268;
  assign \new_[23704]_  = \new_[23703]_  & \new_[23700]_ ;
  assign \new_[23707]_  = ~A300 & ~A299;
  assign \new_[23710]_  = A302 & ~A301;
  assign \new_[23711]_  = \new_[23710]_  & \new_[23707]_ ;
  assign \new_[23712]_  = \new_[23711]_  & \new_[23704]_ ;
  assign \new_[23716]_  = A201 & A200;
  assign \new_[23717]_  = ~A199 & \new_[23716]_ ;
  assign \new_[23720]_  = A232 & ~A203;
  assign \new_[23723]_  = A234 & ~A233;
  assign \new_[23724]_  = \new_[23723]_  & \new_[23720]_ ;
  assign \new_[23725]_  = \new_[23724]_  & \new_[23717]_ ;
  assign \new_[23728]_  = ~A267 & A235;
  assign \new_[23731]_  = ~A298 & A268;
  assign \new_[23732]_  = \new_[23731]_  & \new_[23728]_ ;
  assign \new_[23735]_  = ~A300 & A299;
  assign \new_[23738]_  = A302 & ~A301;
  assign \new_[23739]_  = \new_[23738]_  & \new_[23735]_ ;
  assign \new_[23740]_  = \new_[23739]_  & \new_[23732]_ ;
  assign \new_[23744]_  = A201 & A200;
  assign \new_[23745]_  = ~A199 & \new_[23744]_ ;
  assign \new_[23748]_  = A232 & ~A203;
  assign \new_[23751]_  = A234 & ~A233;
  assign \new_[23752]_  = \new_[23751]_  & \new_[23748]_ ;
  assign \new_[23753]_  = \new_[23752]_  & \new_[23745]_ ;
  assign \new_[23756]_  = ~A267 & A235;
  assign \new_[23759]_  = A298 & ~A269;
  assign \new_[23760]_  = \new_[23759]_  & \new_[23756]_ ;
  assign \new_[23763]_  = ~A300 & ~A299;
  assign \new_[23766]_  = A302 & ~A301;
  assign \new_[23767]_  = \new_[23766]_  & \new_[23763]_ ;
  assign \new_[23768]_  = \new_[23767]_  & \new_[23760]_ ;
  assign \new_[23772]_  = A201 & A200;
  assign \new_[23773]_  = ~A199 & \new_[23772]_ ;
  assign \new_[23776]_  = A232 & ~A203;
  assign \new_[23779]_  = A234 & ~A233;
  assign \new_[23780]_  = \new_[23779]_  & \new_[23776]_ ;
  assign \new_[23781]_  = \new_[23780]_  & \new_[23773]_ ;
  assign \new_[23784]_  = ~A267 & A235;
  assign \new_[23787]_  = ~A298 & ~A269;
  assign \new_[23788]_  = \new_[23787]_  & \new_[23784]_ ;
  assign \new_[23791]_  = ~A300 & A299;
  assign \new_[23794]_  = A302 & ~A301;
  assign \new_[23795]_  = \new_[23794]_  & \new_[23791]_ ;
  assign \new_[23796]_  = \new_[23795]_  & \new_[23788]_ ;
  assign \new_[23800]_  = A201 & A200;
  assign \new_[23801]_  = ~A199 & \new_[23800]_ ;
  assign \new_[23804]_  = A232 & ~A203;
  assign \new_[23807]_  = A234 & ~A233;
  assign \new_[23808]_  = \new_[23807]_  & \new_[23804]_ ;
  assign \new_[23809]_  = \new_[23808]_  & \new_[23801]_ ;
  assign \new_[23812]_  = A265 & A235;
  assign \new_[23815]_  = A298 & A266;
  assign \new_[23816]_  = \new_[23815]_  & \new_[23812]_ ;
  assign \new_[23819]_  = ~A300 & ~A299;
  assign \new_[23822]_  = A302 & ~A301;
  assign \new_[23823]_  = \new_[23822]_  & \new_[23819]_ ;
  assign \new_[23824]_  = \new_[23823]_  & \new_[23816]_ ;
  assign \new_[23828]_  = A201 & A200;
  assign \new_[23829]_  = ~A199 & \new_[23828]_ ;
  assign \new_[23832]_  = A232 & ~A203;
  assign \new_[23835]_  = A234 & ~A233;
  assign \new_[23836]_  = \new_[23835]_  & \new_[23832]_ ;
  assign \new_[23837]_  = \new_[23836]_  & \new_[23829]_ ;
  assign \new_[23840]_  = A265 & A235;
  assign \new_[23843]_  = ~A298 & A266;
  assign \new_[23844]_  = \new_[23843]_  & \new_[23840]_ ;
  assign \new_[23847]_  = ~A300 & A299;
  assign \new_[23850]_  = A302 & ~A301;
  assign \new_[23851]_  = \new_[23850]_  & \new_[23847]_ ;
  assign \new_[23852]_  = \new_[23851]_  & \new_[23844]_ ;
  assign \new_[23856]_  = A201 & A200;
  assign \new_[23857]_  = ~A199 & \new_[23856]_ ;
  assign \new_[23860]_  = A232 & ~A203;
  assign \new_[23863]_  = A234 & ~A233;
  assign \new_[23864]_  = \new_[23863]_  & \new_[23860]_ ;
  assign \new_[23865]_  = \new_[23864]_  & \new_[23857]_ ;
  assign \new_[23868]_  = ~A265 & A235;
  assign \new_[23871]_  = A298 & ~A266;
  assign \new_[23872]_  = \new_[23871]_  & \new_[23868]_ ;
  assign \new_[23875]_  = ~A300 & ~A299;
  assign \new_[23878]_  = A302 & ~A301;
  assign \new_[23879]_  = \new_[23878]_  & \new_[23875]_ ;
  assign \new_[23880]_  = \new_[23879]_  & \new_[23872]_ ;
  assign \new_[23884]_  = A201 & A200;
  assign \new_[23885]_  = ~A199 & \new_[23884]_ ;
  assign \new_[23888]_  = A232 & ~A203;
  assign \new_[23891]_  = A234 & ~A233;
  assign \new_[23892]_  = \new_[23891]_  & \new_[23888]_ ;
  assign \new_[23893]_  = \new_[23892]_  & \new_[23885]_ ;
  assign \new_[23896]_  = ~A265 & A235;
  assign \new_[23899]_  = ~A298 & ~A266;
  assign \new_[23900]_  = \new_[23899]_  & \new_[23896]_ ;
  assign \new_[23903]_  = ~A300 & A299;
  assign \new_[23906]_  = A302 & ~A301;
  assign \new_[23907]_  = \new_[23906]_  & \new_[23903]_ ;
  assign \new_[23908]_  = \new_[23907]_  & \new_[23900]_ ;
  assign \new_[23912]_  = A201 & A200;
  assign \new_[23913]_  = ~A199 & \new_[23912]_ ;
  assign \new_[23916]_  = A232 & ~A203;
  assign \new_[23919]_  = A234 & ~A233;
  assign \new_[23920]_  = \new_[23919]_  & \new_[23916]_ ;
  assign \new_[23921]_  = \new_[23920]_  & \new_[23913]_ ;
  assign \new_[23924]_  = A267 & ~A236;
  assign \new_[23927]_  = A269 & ~A268;
  assign \new_[23928]_  = \new_[23927]_  & \new_[23924]_ ;
  assign \new_[23931]_  = ~A299 & A298;
  assign \new_[23934]_  = A301 & A300;
  assign \new_[23935]_  = \new_[23934]_  & \new_[23931]_ ;
  assign \new_[23936]_  = \new_[23935]_  & \new_[23928]_ ;
  assign \new_[23940]_  = A201 & A200;
  assign \new_[23941]_  = ~A199 & \new_[23940]_ ;
  assign \new_[23944]_  = A232 & ~A203;
  assign \new_[23947]_  = A234 & ~A233;
  assign \new_[23948]_  = \new_[23947]_  & \new_[23944]_ ;
  assign \new_[23949]_  = \new_[23948]_  & \new_[23941]_ ;
  assign \new_[23952]_  = A267 & ~A236;
  assign \new_[23955]_  = A269 & ~A268;
  assign \new_[23956]_  = \new_[23955]_  & \new_[23952]_ ;
  assign \new_[23959]_  = ~A299 & A298;
  assign \new_[23962]_  = ~A302 & A300;
  assign \new_[23963]_  = \new_[23962]_  & \new_[23959]_ ;
  assign \new_[23964]_  = \new_[23963]_  & \new_[23956]_ ;
  assign \new_[23968]_  = A201 & A200;
  assign \new_[23969]_  = ~A199 & \new_[23968]_ ;
  assign \new_[23972]_  = A232 & ~A203;
  assign \new_[23975]_  = A234 & ~A233;
  assign \new_[23976]_  = \new_[23975]_  & \new_[23972]_ ;
  assign \new_[23977]_  = \new_[23976]_  & \new_[23969]_ ;
  assign \new_[23980]_  = A267 & ~A236;
  assign \new_[23983]_  = A269 & ~A268;
  assign \new_[23984]_  = \new_[23983]_  & \new_[23980]_ ;
  assign \new_[23987]_  = A299 & ~A298;
  assign \new_[23990]_  = A301 & A300;
  assign \new_[23991]_  = \new_[23990]_  & \new_[23987]_ ;
  assign \new_[23992]_  = \new_[23991]_  & \new_[23984]_ ;
  assign \new_[23996]_  = A201 & A200;
  assign \new_[23997]_  = ~A199 & \new_[23996]_ ;
  assign \new_[24000]_  = A232 & ~A203;
  assign \new_[24003]_  = A234 & ~A233;
  assign \new_[24004]_  = \new_[24003]_  & \new_[24000]_ ;
  assign \new_[24005]_  = \new_[24004]_  & \new_[23997]_ ;
  assign \new_[24008]_  = A267 & ~A236;
  assign \new_[24011]_  = A269 & ~A268;
  assign \new_[24012]_  = \new_[24011]_  & \new_[24008]_ ;
  assign \new_[24015]_  = A299 & ~A298;
  assign \new_[24018]_  = ~A302 & A300;
  assign \new_[24019]_  = \new_[24018]_  & \new_[24015]_ ;
  assign \new_[24020]_  = \new_[24019]_  & \new_[24012]_ ;
  assign \new_[24024]_  = A201 & A200;
  assign \new_[24025]_  = ~A199 & \new_[24024]_ ;
  assign \new_[24028]_  = A232 & ~A203;
  assign \new_[24031]_  = A234 & ~A233;
  assign \new_[24032]_  = \new_[24031]_  & \new_[24028]_ ;
  assign \new_[24033]_  = \new_[24032]_  & \new_[24025]_ ;
  assign \new_[24036]_  = ~A267 & ~A236;
  assign \new_[24039]_  = A298 & A268;
  assign \new_[24040]_  = \new_[24039]_  & \new_[24036]_ ;
  assign \new_[24043]_  = ~A300 & ~A299;
  assign \new_[24046]_  = A302 & ~A301;
  assign \new_[24047]_  = \new_[24046]_  & \new_[24043]_ ;
  assign \new_[24048]_  = \new_[24047]_  & \new_[24040]_ ;
  assign \new_[24052]_  = A201 & A200;
  assign \new_[24053]_  = ~A199 & \new_[24052]_ ;
  assign \new_[24056]_  = A232 & ~A203;
  assign \new_[24059]_  = A234 & ~A233;
  assign \new_[24060]_  = \new_[24059]_  & \new_[24056]_ ;
  assign \new_[24061]_  = \new_[24060]_  & \new_[24053]_ ;
  assign \new_[24064]_  = ~A267 & ~A236;
  assign \new_[24067]_  = ~A298 & A268;
  assign \new_[24068]_  = \new_[24067]_  & \new_[24064]_ ;
  assign \new_[24071]_  = ~A300 & A299;
  assign \new_[24074]_  = A302 & ~A301;
  assign \new_[24075]_  = \new_[24074]_  & \new_[24071]_ ;
  assign \new_[24076]_  = \new_[24075]_  & \new_[24068]_ ;
  assign \new_[24080]_  = A201 & A200;
  assign \new_[24081]_  = ~A199 & \new_[24080]_ ;
  assign \new_[24084]_  = A232 & ~A203;
  assign \new_[24087]_  = A234 & ~A233;
  assign \new_[24088]_  = \new_[24087]_  & \new_[24084]_ ;
  assign \new_[24089]_  = \new_[24088]_  & \new_[24081]_ ;
  assign \new_[24092]_  = ~A267 & ~A236;
  assign \new_[24095]_  = A298 & ~A269;
  assign \new_[24096]_  = \new_[24095]_  & \new_[24092]_ ;
  assign \new_[24099]_  = ~A300 & ~A299;
  assign \new_[24102]_  = A302 & ~A301;
  assign \new_[24103]_  = \new_[24102]_  & \new_[24099]_ ;
  assign \new_[24104]_  = \new_[24103]_  & \new_[24096]_ ;
  assign \new_[24108]_  = A201 & A200;
  assign \new_[24109]_  = ~A199 & \new_[24108]_ ;
  assign \new_[24112]_  = A232 & ~A203;
  assign \new_[24115]_  = A234 & ~A233;
  assign \new_[24116]_  = \new_[24115]_  & \new_[24112]_ ;
  assign \new_[24117]_  = \new_[24116]_  & \new_[24109]_ ;
  assign \new_[24120]_  = ~A267 & ~A236;
  assign \new_[24123]_  = ~A298 & ~A269;
  assign \new_[24124]_  = \new_[24123]_  & \new_[24120]_ ;
  assign \new_[24127]_  = ~A300 & A299;
  assign \new_[24130]_  = A302 & ~A301;
  assign \new_[24131]_  = \new_[24130]_  & \new_[24127]_ ;
  assign \new_[24132]_  = \new_[24131]_  & \new_[24124]_ ;
  assign \new_[24136]_  = A201 & A200;
  assign \new_[24137]_  = ~A199 & \new_[24136]_ ;
  assign \new_[24140]_  = A232 & ~A203;
  assign \new_[24143]_  = A234 & ~A233;
  assign \new_[24144]_  = \new_[24143]_  & \new_[24140]_ ;
  assign \new_[24145]_  = \new_[24144]_  & \new_[24137]_ ;
  assign \new_[24148]_  = A265 & ~A236;
  assign \new_[24151]_  = A298 & A266;
  assign \new_[24152]_  = \new_[24151]_  & \new_[24148]_ ;
  assign \new_[24155]_  = ~A300 & ~A299;
  assign \new_[24158]_  = A302 & ~A301;
  assign \new_[24159]_  = \new_[24158]_  & \new_[24155]_ ;
  assign \new_[24160]_  = \new_[24159]_  & \new_[24152]_ ;
  assign \new_[24164]_  = A201 & A200;
  assign \new_[24165]_  = ~A199 & \new_[24164]_ ;
  assign \new_[24168]_  = A232 & ~A203;
  assign \new_[24171]_  = A234 & ~A233;
  assign \new_[24172]_  = \new_[24171]_  & \new_[24168]_ ;
  assign \new_[24173]_  = \new_[24172]_  & \new_[24165]_ ;
  assign \new_[24176]_  = A265 & ~A236;
  assign \new_[24179]_  = ~A298 & A266;
  assign \new_[24180]_  = \new_[24179]_  & \new_[24176]_ ;
  assign \new_[24183]_  = ~A300 & A299;
  assign \new_[24186]_  = A302 & ~A301;
  assign \new_[24187]_  = \new_[24186]_  & \new_[24183]_ ;
  assign \new_[24188]_  = \new_[24187]_  & \new_[24180]_ ;
  assign \new_[24192]_  = A201 & A200;
  assign \new_[24193]_  = ~A199 & \new_[24192]_ ;
  assign \new_[24196]_  = A232 & ~A203;
  assign \new_[24199]_  = A234 & ~A233;
  assign \new_[24200]_  = \new_[24199]_  & \new_[24196]_ ;
  assign \new_[24201]_  = \new_[24200]_  & \new_[24193]_ ;
  assign \new_[24204]_  = ~A265 & ~A236;
  assign \new_[24207]_  = A298 & ~A266;
  assign \new_[24208]_  = \new_[24207]_  & \new_[24204]_ ;
  assign \new_[24211]_  = ~A300 & ~A299;
  assign \new_[24214]_  = A302 & ~A301;
  assign \new_[24215]_  = \new_[24214]_  & \new_[24211]_ ;
  assign \new_[24216]_  = \new_[24215]_  & \new_[24208]_ ;
  assign \new_[24220]_  = A201 & A200;
  assign \new_[24221]_  = ~A199 & \new_[24220]_ ;
  assign \new_[24224]_  = A232 & ~A203;
  assign \new_[24227]_  = A234 & ~A233;
  assign \new_[24228]_  = \new_[24227]_  & \new_[24224]_ ;
  assign \new_[24229]_  = \new_[24228]_  & \new_[24221]_ ;
  assign \new_[24232]_  = ~A265 & ~A236;
  assign \new_[24235]_  = ~A298 & ~A266;
  assign \new_[24236]_  = \new_[24235]_  & \new_[24232]_ ;
  assign \new_[24239]_  = ~A300 & A299;
  assign \new_[24242]_  = A302 & ~A301;
  assign \new_[24243]_  = \new_[24242]_  & \new_[24239]_ ;
  assign \new_[24244]_  = \new_[24243]_  & \new_[24236]_ ;
  assign \new_[24248]_  = A201 & A200;
  assign \new_[24249]_  = ~A199 & \new_[24248]_ ;
  assign \new_[24252]_  = A232 & ~A203;
  assign \new_[24255]_  = ~A234 & ~A233;
  assign \new_[24256]_  = \new_[24255]_  & \new_[24252]_ ;
  assign \new_[24257]_  = \new_[24256]_  & \new_[24249]_ ;
  assign \new_[24260]_  = A236 & ~A235;
  assign \new_[24263]_  = A268 & ~A267;
  assign \new_[24264]_  = \new_[24263]_  & \new_[24260]_ ;
  assign \new_[24267]_  = ~A299 & A298;
  assign \new_[24270]_  = A301 & A300;
  assign \new_[24271]_  = \new_[24270]_  & \new_[24267]_ ;
  assign \new_[24272]_  = \new_[24271]_  & \new_[24264]_ ;
  assign \new_[24276]_  = A201 & A200;
  assign \new_[24277]_  = ~A199 & \new_[24276]_ ;
  assign \new_[24280]_  = A232 & ~A203;
  assign \new_[24283]_  = ~A234 & ~A233;
  assign \new_[24284]_  = \new_[24283]_  & \new_[24280]_ ;
  assign \new_[24285]_  = \new_[24284]_  & \new_[24277]_ ;
  assign \new_[24288]_  = A236 & ~A235;
  assign \new_[24291]_  = A268 & ~A267;
  assign \new_[24292]_  = \new_[24291]_  & \new_[24288]_ ;
  assign \new_[24295]_  = ~A299 & A298;
  assign \new_[24298]_  = ~A302 & A300;
  assign \new_[24299]_  = \new_[24298]_  & \new_[24295]_ ;
  assign \new_[24300]_  = \new_[24299]_  & \new_[24292]_ ;
  assign \new_[24304]_  = A201 & A200;
  assign \new_[24305]_  = ~A199 & \new_[24304]_ ;
  assign \new_[24308]_  = A232 & ~A203;
  assign \new_[24311]_  = ~A234 & ~A233;
  assign \new_[24312]_  = \new_[24311]_  & \new_[24308]_ ;
  assign \new_[24313]_  = \new_[24312]_  & \new_[24305]_ ;
  assign \new_[24316]_  = A236 & ~A235;
  assign \new_[24319]_  = A268 & ~A267;
  assign \new_[24320]_  = \new_[24319]_  & \new_[24316]_ ;
  assign \new_[24323]_  = A299 & ~A298;
  assign \new_[24326]_  = A301 & A300;
  assign \new_[24327]_  = \new_[24326]_  & \new_[24323]_ ;
  assign \new_[24328]_  = \new_[24327]_  & \new_[24320]_ ;
  assign \new_[24332]_  = A201 & A200;
  assign \new_[24333]_  = ~A199 & \new_[24332]_ ;
  assign \new_[24336]_  = A232 & ~A203;
  assign \new_[24339]_  = ~A234 & ~A233;
  assign \new_[24340]_  = \new_[24339]_  & \new_[24336]_ ;
  assign \new_[24341]_  = \new_[24340]_  & \new_[24333]_ ;
  assign \new_[24344]_  = A236 & ~A235;
  assign \new_[24347]_  = A268 & ~A267;
  assign \new_[24348]_  = \new_[24347]_  & \new_[24344]_ ;
  assign \new_[24351]_  = A299 & ~A298;
  assign \new_[24354]_  = ~A302 & A300;
  assign \new_[24355]_  = \new_[24354]_  & \new_[24351]_ ;
  assign \new_[24356]_  = \new_[24355]_  & \new_[24348]_ ;
  assign \new_[24360]_  = A201 & A200;
  assign \new_[24361]_  = ~A199 & \new_[24360]_ ;
  assign \new_[24364]_  = A232 & ~A203;
  assign \new_[24367]_  = ~A234 & ~A233;
  assign \new_[24368]_  = \new_[24367]_  & \new_[24364]_ ;
  assign \new_[24369]_  = \new_[24368]_  & \new_[24361]_ ;
  assign \new_[24372]_  = A236 & ~A235;
  assign \new_[24375]_  = ~A269 & ~A267;
  assign \new_[24376]_  = \new_[24375]_  & \new_[24372]_ ;
  assign \new_[24379]_  = ~A299 & A298;
  assign \new_[24382]_  = A301 & A300;
  assign \new_[24383]_  = \new_[24382]_  & \new_[24379]_ ;
  assign \new_[24384]_  = \new_[24383]_  & \new_[24376]_ ;
  assign \new_[24388]_  = A201 & A200;
  assign \new_[24389]_  = ~A199 & \new_[24388]_ ;
  assign \new_[24392]_  = A232 & ~A203;
  assign \new_[24395]_  = ~A234 & ~A233;
  assign \new_[24396]_  = \new_[24395]_  & \new_[24392]_ ;
  assign \new_[24397]_  = \new_[24396]_  & \new_[24389]_ ;
  assign \new_[24400]_  = A236 & ~A235;
  assign \new_[24403]_  = ~A269 & ~A267;
  assign \new_[24404]_  = \new_[24403]_  & \new_[24400]_ ;
  assign \new_[24407]_  = ~A299 & A298;
  assign \new_[24410]_  = ~A302 & A300;
  assign \new_[24411]_  = \new_[24410]_  & \new_[24407]_ ;
  assign \new_[24412]_  = \new_[24411]_  & \new_[24404]_ ;
  assign \new_[24416]_  = A201 & A200;
  assign \new_[24417]_  = ~A199 & \new_[24416]_ ;
  assign \new_[24420]_  = A232 & ~A203;
  assign \new_[24423]_  = ~A234 & ~A233;
  assign \new_[24424]_  = \new_[24423]_  & \new_[24420]_ ;
  assign \new_[24425]_  = \new_[24424]_  & \new_[24417]_ ;
  assign \new_[24428]_  = A236 & ~A235;
  assign \new_[24431]_  = ~A269 & ~A267;
  assign \new_[24432]_  = \new_[24431]_  & \new_[24428]_ ;
  assign \new_[24435]_  = A299 & ~A298;
  assign \new_[24438]_  = A301 & A300;
  assign \new_[24439]_  = \new_[24438]_  & \new_[24435]_ ;
  assign \new_[24440]_  = \new_[24439]_  & \new_[24432]_ ;
  assign \new_[24444]_  = A201 & A200;
  assign \new_[24445]_  = ~A199 & \new_[24444]_ ;
  assign \new_[24448]_  = A232 & ~A203;
  assign \new_[24451]_  = ~A234 & ~A233;
  assign \new_[24452]_  = \new_[24451]_  & \new_[24448]_ ;
  assign \new_[24453]_  = \new_[24452]_  & \new_[24445]_ ;
  assign \new_[24456]_  = A236 & ~A235;
  assign \new_[24459]_  = ~A269 & ~A267;
  assign \new_[24460]_  = \new_[24459]_  & \new_[24456]_ ;
  assign \new_[24463]_  = A299 & ~A298;
  assign \new_[24466]_  = ~A302 & A300;
  assign \new_[24467]_  = \new_[24466]_  & \new_[24463]_ ;
  assign \new_[24468]_  = \new_[24467]_  & \new_[24460]_ ;
  assign \new_[24472]_  = A201 & A200;
  assign \new_[24473]_  = ~A199 & \new_[24472]_ ;
  assign \new_[24476]_  = A232 & ~A203;
  assign \new_[24479]_  = ~A234 & ~A233;
  assign \new_[24480]_  = \new_[24479]_  & \new_[24476]_ ;
  assign \new_[24481]_  = \new_[24480]_  & \new_[24473]_ ;
  assign \new_[24484]_  = A236 & ~A235;
  assign \new_[24487]_  = A266 & A265;
  assign \new_[24488]_  = \new_[24487]_  & \new_[24484]_ ;
  assign \new_[24491]_  = ~A299 & A298;
  assign \new_[24494]_  = A301 & A300;
  assign \new_[24495]_  = \new_[24494]_  & \new_[24491]_ ;
  assign \new_[24496]_  = \new_[24495]_  & \new_[24488]_ ;
  assign \new_[24500]_  = A201 & A200;
  assign \new_[24501]_  = ~A199 & \new_[24500]_ ;
  assign \new_[24504]_  = A232 & ~A203;
  assign \new_[24507]_  = ~A234 & ~A233;
  assign \new_[24508]_  = \new_[24507]_  & \new_[24504]_ ;
  assign \new_[24509]_  = \new_[24508]_  & \new_[24501]_ ;
  assign \new_[24512]_  = A236 & ~A235;
  assign \new_[24515]_  = A266 & A265;
  assign \new_[24516]_  = \new_[24515]_  & \new_[24512]_ ;
  assign \new_[24519]_  = ~A299 & A298;
  assign \new_[24522]_  = ~A302 & A300;
  assign \new_[24523]_  = \new_[24522]_  & \new_[24519]_ ;
  assign \new_[24524]_  = \new_[24523]_  & \new_[24516]_ ;
  assign \new_[24528]_  = A201 & A200;
  assign \new_[24529]_  = ~A199 & \new_[24528]_ ;
  assign \new_[24532]_  = A232 & ~A203;
  assign \new_[24535]_  = ~A234 & ~A233;
  assign \new_[24536]_  = \new_[24535]_  & \new_[24532]_ ;
  assign \new_[24537]_  = \new_[24536]_  & \new_[24529]_ ;
  assign \new_[24540]_  = A236 & ~A235;
  assign \new_[24543]_  = A266 & A265;
  assign \new_[24544]_  = \new_[24543]_  & \new_[24540]_ ;
  assign \new_[24547]_  = A299 & ~A298;
  assign \new_[24550]_  = A301 & A300;
  assign \new_[24551]_  = \new_[24550]_  & \new_[24547]_ ;
  assign \new_[24552]_  = \new_[24551]_  & \new_[24544]_ ;
  assign \new_[24556]_  = A201 & A200;
  assign \new_[24557]_  = ~A199 & \new_[24556]_ ;
  assign \new_[24560]_  = A232 & ~A203;
  assign \new_[24563]_  = ~A234 & ~A233;
  assign \new_[24564]_  = \new_[24563]_  & \new_[24560]_ ;
  assign \new_[24565]_  = \new_[24564]_  & \new_[24557]_ ;
  assign \new_[24568]_  = A236 & ~A235;
  assign \new_[24571]_  = A266 & A265;
  assign \new_[24572]_  = \new_[24571]_  & \new_[24568]_ ;
  assign \new_[24575]_  = A299 & ~A298;
  assign \new_[24578]_  = ~A302 & A300;
  assign \new_[24579]_  = \new_[24578]_  & \new_[24575]_ ;
  assign \new_[24580]_  = \new_[24579]_  & \new_[24572]_ ;
  assign \new_[24584]_  = A201 & A200;
  assign \new_[24585]_  = ~A199 & \new_[24584]_ ;
  assign \new_[24588]_  = A232 & ~A203;
  assign \new_[24591]_  = ~A234 & ~A233;
  assign \new_[24592]_  = \new_[24591]_  & \new_[24588]_ ;
  assign \new_[24593]_  = \new_[24592]_  & \new_[24585]_ ;
  assign \new_[24596]_  = A236 & ~A235;
  assign \new_[24599]_  = ~A266 & ~A265;
  assign \new_[24600]_  = \new_[24599]_  & \new_[24596]_ ;
  assign \new_[24603]_  = ~A299 & A298;
  assign \new_[24606]_  = A301 & A300;
  assign \new_[24607]_  = \new_[24606]_  & \new_[24603]_ ;
  assign \new_[24608]_  = \new_[24607]_  & \new_[24600]_ ;
  assign \new_[24612]_  = A201 & A200;
  assign \new_[24613]_  = ~A199 & \new_[24612]_ ;
  assign \new_[24616]_  = A232 & ~A203;
  assign \new_[24619]_  = ~A234 & ~A233;
  assign \new_[24620]_  = \new_[24619]_  & \new_[24616]_ ;
  assign \new_[24621]_  = \new_[24620]_  & \new_[24613]_ ;
  assign \new_[24624]_  = A236 & ~A235;
  assign \new_[24627]_  = ~A266 & ~A265;
  assign \new_[24628]_  = \new_[24627]_  & \new_[24624]_ ;
  assign \new_[24631]_  = ~A299 & A298;
  assign \new_[24634]_  = ~A302 & A300;
  assign \new_[24635]_  = \new_[24634]_  & \new_[24631]_ ;
  assign \new_[24636]_  = \new_[24635]_  & \new_[24628]_ ;
  assign \new_[24640]_  = A201 & A200;
  assign \new_[24641]_  = ~A199 & \new_[24640]_ ;
  assign \new_[24644]_  = A232 & ~A203;
  assign \new_[24647]_  = ~A234 & ~A233;
  assign \new_[24648]_  = \new_[24647]_  & \new_[24644]_ ;
  assign \new_[24649]_  = \new_[24648]_  & \new_[24641]_ ;
  assign \new_[24652]_  = A236 & ~A235;
  assign \new_[24655]_  = ~A266 & ~A265;
  assign \new_[24656]_  = \new_[24655]_  & \new_[24652]_ ;
  assign \new_[24659]_  = A299 & ~A298;
  assign \new_[24662]_  = A301 & A300;
  assign \new_[24663]_  = \new_[24662]_  & \new_[24659]_ ;
  assign \new_[24664]_  = \new_[24663]_  & \new_[24656]_ ;
  assign \new_[24668]_  = A201 & A200;
  assign \new_[24669]_  = ~A199 & \new_[24668]_ ;
  assign \new_[24672]_  = A232 & ~A203;
  assign \new_[24675]_  = ~A234 & ~A233;
  assign \new_[24676]_  = \new_[24675]_  & \new_[24672]_ ;
  assign \new_[24677]_  = \new_[24676]_  & \new_[24669]_ ;
  assign \new_[24680]_  = A236 & ~A235;
  assign \new_[24683]_  = ~A266 & ~A265;
  assign \new_[24684]_  = \new_[24683]_  & \new_[24680]_ ;
  assign \new_[24687]_  = A299 & ~A298;
  assign \new_[24690]_  = ~A302 & A300;
  assign \new_[24691]_  = \new_[24690]_  & \new_[24687]_ ;
  assign \new_[24692]_  = \new_[24691]_  & \new_[24684]_ ;
  assign \new_[24696]_  = ~A201 & A200;
  assign \new_[24697]_  = ~A199 & \new_[24696]_ ;
  assign \new_[24700]_  = A203 & ~A202;
  assign \new_[24703]_  = A233 & ~A232;
  assign \new_[24704]_  = \new_[24703]_  & \new_[24700]_ ;
  assign \new_[24705]_  = \new_[24704]_  & \new_[24697]_ ;
  assign \new_[24708]_  = A235 & A234;
  assign \new_[24711]_  = A268 & ~A267;
  assign \new_[24712]_  = \new_[24711]_  & \new_[24708]_ ;
  assign \new_[24715]_  = ~A299 & A298;
  assign \new_[24718]_  = A301 & A300;
  assign \new_[24719]_  = \new_[24718]_  & \new_[24715]_ ;
  assign \new_[24720]_  = \new_[24719]_  & \new_[24712]_ ;
  assign \new_[24724]_  = ~A201 & A200;
  assign \new_[24725]_  = ~A199 & \new_[24724]_ ;
  assign \new_[24728]_  = A203 & ~A202;
  assign \new_[24731]_  = A233 & ~A232;
  assign \new_[24732]_  = \new_[24731]_  & \new_[24728]_ ;
  assign \new_[24733]_  = \new_[24732]_  & \new_[24725]_ ;
  assign \new_[24736]_  = A235 & A234;
  assign \new_[24739]_  = A268 & ~A267;
  assign \new_[24740]_  = \new_[24739]_  & \new_[24736]_ ;
  assign \new_[24743]_  = ~A299 & A298;
  assign \new_[24746]_  = ~A302 & A300;
  assign \new_[24747]_  = \new_[24746]_  & \new_[24743]_ ;
  assign \new_[24748]_  = \new_[24747]_  & \new_[24740]_ ;
  assign \new_[24752]_  = ~A201 & A200;
  assign \new_[24753]_  = ~A199 & \new_[24752]_ ;
  assign \new_[24756]_  = A203 & ~A202;
  assign \new_[24759]_  = A233 & ~A232;
  assign \new_[24760]_  = \new_[24759]_  & \new_[24756]_ ;
  assign \new_[24761]_  = \new_[24760]_  & \new_[24753]_ ;
  assign \new_[24764]_  = A235 & A234;
  assign \new_[24767]_  = A268 & ~A267;
  assign \new_[24768]_  = \new_[24767]_  & \new_[24764]_ ;
  assign \new_[24771]_  = A299 & ~A298;
  assign \new_[24774]_  = A301 & A300;
  assign \new_[24775]_  = \new_[24774]_  & \new_[24771]_ ;
  assign \new_[24776]_  = \new_[24775]_  & \new_[24768]_ ;
  assign \new_[24780]_  = ~A201 & A200;
  assign \new_[24781]_  = ~A199 & \new_[24780]_ ;
  assign \new_[24784]_  = A203 & ~A202;
  assign \new_[24787]_  = A233 & ~A232;
  assign \new_[24788]_  = \new_[24787]_  & \new_[24784]_ ;
  assign \new_[24789]_  = \new_[24788]_  & \new_[24781]_ ;
  assign \new_[24792]_  = A235 & A234;
  assign \new_[24795]_  = A268 & ~A267;
  assign \new_[24796]_  = \new_[24795]_  & \new_[24792]_ ;
  assign \new_[24799]_  = A299 & ~A298;
  assign \new_[24802]_  = ~A302 & A300;
  assign \new_[24803]_  = \new_[24802]_  & \new_[24799]_ ;
  assign \new_[24804]_  = \new_[24803]_  & \new_[24796]_ ;
  assign \new_[24808]_  = ~A201 & A200;
  assign \new_[24809]_  = ~A199 & \new_[24808]_ ;
  assign \new_[24812]_  = A203 & ~A202;
  assign \new_[24815]_  = A233 & ~A232;
  assign \new_[24816]_  = \new_[24815]_  & \new_[24812]_ ;
  assign \new_[24817]_  = \new_[24816]_  & \new_[24809]_ ;
  assign \new_[24820]_  = A235 & A234;
  assign \new_[24823]_  = ~A269 & ~A267;
  assign \new_[24824]_  = \new_[24823]_  & \new_[24820]_ ;
  assign \new_[24827]_  = ~A299 & A298;
  assign \new_[24830]_  = A301 & A300;
  assign \new_[24831]_  = \new_[24830]_  & \new_[24827]_ ;
  assign \new_[24832]_  = \new_[24831]_  & \new_[24824]_ ;
  assign \new_[24836]_  = ~A201 & A200;
  assign \new_[24837]_  = ~A199 & \new_[24836]_ ;
  assign \new_[24840]_  = A203 & ~A202;
  assign \new_[24843]_  = A233 & ~A232;
  assign \new_[24844]_  = \new_[24843]_  & \new_[24840]_ ;
  assign \new_[24845]_  = \new_[24844]_  & \new_[24837]_ ;
  assign \new_[24848]_  = A235 & A234;
  assign \new_[24851]_  = ~A269 & ~A267;
  assign \new_[24852]_  = \new_[24851]_  & \new_[24848]_ ;
  assign \new_[24855]_  = ~A299 & A298;
  assign \new_[24858]_  = ~A302 & A300;
  assign \new_[24859]_  = \new_[24858]_  & \new_[24855]_ ;
  assign \new_[24860]_  = \new_[24859]_  & \new_[24852]_ ;
  assign \new_[24864]_  = ~A201 & A200;
  assign \new_[24865]_  = ~A199 & \new_[24864]_ ;
  assign \new_[24868]_  = A203 & ~A202;
  assign \new_[24871]_  = A233 & ~A232;
  assign \new_[24872]_  = \new_[24871]_  & \new_[24868]_ ;
  assign \new_[24873]_  = \new_[24872]_  & \new_[24865]_ ;
  assign \new_[24876]_  = A235 & A234;
  assign \new_[24879]_  = ~A269 & ~A267;
  assign \new_[24880]_  = \new_[24879]_  & \new_[24876]_ ;
  assign \new_[24883]_  = A299 & ~A298;
  assign \new_[24886]_  = A301 & A300;
  assign \new_[24887]_  = \new_[24886]_  & \new_[24883]_ ;
  assign \new_[24888]_  = \new_[24887]_  & \new_[24880]_ ;
  assign \new_[24892]_  = ~A201 & A200;
  assign \new_[24893]_  = ~A199 & \new_[24892]_ ;
  assign \new_[24896]_  = A203 & ~A202;
  assign \new_[24899]_  = A233 & ~A232;
  assign \new_[24900]_  = \new_[24899]_  & \new_[24896]_ ;
  assign \new_[24901]_  = \new_[24900]_  & \new_[24893]_ ;
  assign \new_[24904]_  = A235 & A234;
  assign \new_[24907]_  = ~A269 & ~A267;
  assign \new_[24908]_  = \new_[24907]_  & \new_[24904]_ ;
  assign \new_[24911]_  = A299 & ~A298;
  assign \new_[24914]_  = ~A302 & A300;
  assign \new_[24915]_  = \new_[24914]_  & \new_[24911]_ ;
  assign \new_[24916]_  = \new_[24915]_  & \new_[24908]_ ;
  assign \new_[24920]_  = ~A201 & A200;
  assign \new_[24921]_  = ~A199 & \new_[24920]_ ;
  assign \new_[24924]_  = A203 & ~A202;
  assign \new_[24927]_  = A233 & ~A232;
  assign \new_[24928]_  = \new_[24927]_  & \new_[24924]_ ;
  assign \new_[24929]_  = \new_[24928]_  & \new_[24921]_ ;
  assign \new_[24932]_  = A235 & A234;
  assign \new_[24935]_  = A266 & A265;
  assign \new_[24936]_  = \new_[24935]_  & \new_[24932]_ ;
  assign \new_[24939]_  = ~A299 & A298;
  assign \new_[24942]_  = A301 & A300;
  assign \new_[24943]_  = \new_[24942]_  & \new_[24939]_ ;
  assign \new_[24944]_  = \new_[24943]_  & \new_[24936]_ ;
  assign \new_[24948]_  = ~A201 & A200;
  assign \new_[24949]_  = ~A199 & \new_[24948]_ ;
  assign \new_[24952]_  = A203 & ~A202;
  assign \new_[24955]_  = A233 & ~A232;
  assign \new_[24956]_  = \new_[24955]_  & \new_[24952]_ ;
  assign \new_[24957]_  = \new_[24956]_  & \new_[24949]_ ;
  assign \new_[24960]_  = A235 & A234;
  assign \new_[24963]_  = A266 & A265;
  assign \new_[24964]_  = \new_[24963]_  & \new_[24960]_ ;
  assign \new_[24967]_  = ~A299 & A298;
  assign \new_[24970]_  = ~A302 & A300;
  assign \new_[24971]_  = \new_[24970]_  & \new_[24967]_ ;
  assign \new_[24972]_  = \new_[24971]_  & \new_[24964]_ ;
  assign \new_[24976]_  = ~A201 & A200;
  assign \new_[24977]_  = ~A199 & \new_[24976]_ ;
  assign \new_[24980]_  = A203 & ~A202;
  assign \new_[24983]_  = A233 & ~A232;
  assign \new_[24984]_  = \new_[24983]_  & \new_[24980]_ ;
  assign \new_[24985]_  = \new_[24984]_  & \new_[24977]_ ;
  assign \new_[24988]_  = A235 & A234;
  assign \new_[24991]_  = A266 & A265;
  assign \new_[24992]_  = \new_[24991]_  & \new_[24988]_ ;
  assign \new_[24995]_  = A299 & ~A298;
  assign \new_[24998]_  = A301 & A300;
  assign \new_[24999]_  = \new_[24998]_  & \new_[24995]_ ;
  assign \new_[25000]_  = \new_[24999]_  & \new_[24992]_ ;
  assign \new_[25004]_  = ~A201 & A200;
  assign \new_[25005]_  = ~A199 & \new_[25004]_ ;
  assign \new_[25008]_  = A203 & ~A202;
  assign \new_[25011]_  = A233 & ~A232;
  assign \new_[25012]_  = \new_[25011]_  & \new_[25008]_ ;
  assign \new_[25013]_  = \new_[25012]_  & \new_[25005]_ ;
  assign \new_[25016]_  = A235 & A234;
  assign \new_[25019]_  = A266 & A265;
  assign \new_[25020]_  = \new_[25019]_  & \new_[25016]_ ;
  assign \new_[25023]_  = A299 & ~A298;
  assign \new_[25026]_  = ~A302 & A300;
  assign \new_[25027]_  = \new_[25026]_  & \new_[25023]_ ;
  assign \new_[25028]_  = \new_[25027]_  & \new_[25020]_ ;
  assign \new_[25032]_  = ~A201 & A200;
  assign \new_[25033]_  = ~A199 & \new_[25032]_ ;
  assign \new_[25036]_  = A203 & ~A202;
  assign \new_[25039]_  = A233 & ~A232;
  assign \new_[25040]_  = \new_[25039]_  & \new_[25036]_ ;
  assign \new_[25041]_  = \new_[25040]_  & \new_[25033]_ ;
  assign \new_[25044]_  = A235 & A234;
  assign \new_[25047]_  = ~A266 & ~A265;
  assign \new_[25048]_  = \new_[25047]_  & \new_[25044]_ ;
  assign \new_[25051]_  = ~A299 & A298;
  assign \new_[25054]_  = A301 & A300;
  assign \new_[25055]_  = \new_[25054]_  & \new_[25051]_ ;
  assign \new_[25056]_  = \new_[25055]_  & \new_[25048]_ ;
  assign \new_[25060]_  = ~A201 & A200;
  assign \new_[25061]_  = ~A199 & \new_[25060]_ ;
  assign \new_[25064]_  = A203 & ~A202;
  assign \new_[25067]_  = A233 & ~A232;
  assign \new_[25068]_  = \new_[25067]_  & \new_[25064]_ ;
  assign \new_[25069]_  = \new_[25068]_  & \new_[25061]_ ;
  assign \new_[25072]_  = A235 & A234;
  assign \new_[25075]_  = ~A266 & ~A265;
  assign \new_[25076]_  = \new_[25075]_  & \new_[25072]_ ;
  assign \new_[25079]_  = ~A299 & A298;
  assign \new_[25082]_  = ~A302 & A300;
  assign \new_[25083]_  = \new_[25082]_  & \new_[25079]_ ;
  assign \new_[25084]_  = \new_[25083]_  & \new_[25076]_ ;
  assign \new_[25088]_  = ~A201 & A200;
  assign \new_[25089]_  = ~A199 & \new_[25088]_ ;
  assign \new_[25092]_  = A203 & ~A202;
  assign \new_[25095]_  = A233 & ~A232;
  assign \new_[25096]_  = \new_[25095]_  & \new_[25092]_ ;
  assign \new_[25097]_  = \new_[25096]_  & \new_[25089]_ ;
  assign \new_[25100]_  = A235 & A234;
  assign \new_[25103]_  = ~A266 & ~A265;
  assign \new_[25104]_  = \new_[25103]_  & \new_[25100]_ ;
  assign \new_[25107]_  = A299 & ~A298;
  assign \new_[25110]_  = A301 & A300;
  assign \new_[25111]_  = \new_[25110]_  & \new_[25107]_ ;
  assign \new_[25112]_  = \new_[25111]_  & \new_[25104]_ ;
  assign \new_[25116]_  = ~A201 & A200;
  assign \new_[25117]_  = ~A199 & \new_[25116]_ ;
  assign \new_[25120]_  = A203 & ~A202;
  assign \new_[25123]_  = A233 & ~A232;
  assign \new_[25124]_  = \new_[25123]_  & \new_[25120]_ ;
  assign \new_[25125]_  = \new_[25124]_  & \new_[25117]_ ;
  assign \new_[25128]_  = A235 & A234;
  assign \new_[25131]_  = ~A266 & ~A265;
  assign \new_[25132]_  = \new_[25131]_  & \new_[25128]_ ;
  assign \new_[25135]_  = A299 & ~A298;
  assign \new_[25138]_  = ~A302 & A300;
  assign \new_[25139]_  = \new_[25138]_  & \new_[25135]_ ;
  assign \new_[25140]_  = \new_[25139]_  & \new_[25132]_ ;
  assign \new_[25144]_  = ~A201 & A200;
  assign \new_[25145]_  = ~A199 & \new_[25144]_ ;
  assign \new_[25148]_  = A203 & ~A202;
  assign \new_[25151]_  = A233 & ~A232;
  assign \new_[25152]_  = \new_[25151]_  & \new_[25148]_ ;
  assign \new_[25153]_  = \new_[25152]_  & \new_[25145]_ ;
  assign \new_[25156]_  = ~A236 & A234;
  assign \new_[25159]_  = A268 & ~A267;
  assign \new_[25160]_  = \new_[25159]_  & \new_[25156]_ ;
  assign \new_[25163]_  = ~A299 & A298;
  assign \new_[25166]_  = A301 & A300;
  assign \new_[25167]_  = \new_[25166]_  & \new_[25163]_ ;
  assign \new_[25168]_  = \new_[25167]_  & \new_[25160]_ ;
  assign \new_[25172]_  = ~A201 & A200;
  assign \new_[25173]_  = ~A199 & \new_[25172]_ ;
  assign \new_[25176]_  = A203 & ~A202;
  assign \new_[25179]_  = A233 & ~A232;
  assign \new_[25180]_  = \new_[25179]_  & \new_[25176]_ ;
  assign \new_[25181]_  = \new_[25180]_  & \new_[25173]_ ;
  assign \new_[25184]_  = ~A236 & A234;
  assign \new_[25187]_  = A268 & ~A267;
  assign \new_[25188]_  = \new_[25187]_  & \new_[25184]_ ;
  assign \new_[25191]_  = ~A299 & A298;
  assign \new_[25194]_  = ~A302 & A300;
  assign \new_[25195]_  = \new_[25194]_  & \new_[25191]_ ;
  assign \new_[25196]_  = \new_[25195]_  & \new_[25188]_ ;
  assign \new_[25200]_  = ~A201 & A200;
  assign \new_[25201]_  = ~A199 & \new_[25200]_ ;
  assign \new_[25204]_  = A203 & ~A202;
  assign \new_[25207]_  = A233 & ~A232;
  assign \new_[25208]_  = \new_[25207]_  & \new_[25204]_ ;
  assign \new_[25209]_  = \new_[25208]_  & \new_[25201]_ ;
  assign \new_[25212]_  = ~A236 & A234;
  assign \new_[25215]_  = A268 & ~A267;
  assign \new_[25216]_  = \new_[25215]_  & \new_[25212]_ ;
  assign \new_[25219]_  = A299 & ~A298;
  assign \new_[25222]_  = A301 & A300;
  assign \new_[25223]_  = \new_[25222]_  & \new_[25219]_ ;
  assign \new_[25224]_  = \new_[25223]_  & \new_[25216]_ ;
  assign \new_[25228]_  = ~A201 & A200;
  assign \new_[25229]_  = ~A199 & \new_[25228]_ ;
  assign \new_[25232]_  = A203 & ~A202;
  assign \new_[25235]_  = A233 & ~A232;
  assign \new_[25236]_  = \new_[25235]_  & \new_[25232]_ ;
  assign \new_[25237]_  = \new_[25236]_  & \new_[25229]_ ;
  assign \new_[25240]_  = ~A236 & A234;
  assign \new_[25243]_  = A268 & ~A267;
  assign \new_[25244]_  = \new_[25243]_  & \new_[25240]_ ;
  assign \new_[25247]_  = A299 & ~A298;
  assign \new_[25250]_  = ~A302 & A300;
  assign \new_[25251]_  = \new_[25250]_  & \new_[25247]_ ;
  assign \new_[25252]_  = \new_[25251]_  & \new_[25244]_ ;
  assign \new_[25256]_  = ~A201 & A200;
  assign \new_[25257]_  = ~A199 & \new_[25256]_ ;
  assign \new_[25260]_  = A203 & ~A202;
  assign \new_[25263]_  = A233 & ~A232;
  assign \new_[25264]_  = \new_[25263]_  & \new_[25260]_ ;
  assign \new_[25265]_  = \new_[25264]_  & \new_[25257]_ ;
  assign \new_[25268]_  = ~A236 & A234;
  assign \new_[25271]_  = ~A269 & ~A267;
  assign \new_[25272]_  = \new_[25271]_  & \new_[25268]_ ;
  assign \new_[25275]_  = ~A299 & A298;
  assign \new_[25278]_  = A301 & A300;
  assign \new_[25279]_  = \new_[25278]_  & \new_[25275]_ ;
  assign \new_[25280]_  = \new_[25279]_  & \new_[25272]_ ;
  assign \new_[25284]_  = ~A201 & A200;
  assign \new_[25285]_  = ~A199 & \new_[25284]_ ;
  assign \new_[25288]_  = A203 & ~A202;
  assign \new_[25291]_  = A233 & ~A232;
  assign \new_[25292]_  = \new_[25291]_  & \new_[25288]_ ;
  assign \new_[25293]_  = \new_[25292]_  & \new_[25285]_ ;
  assign \new_[25296]_  = ~A236 & A234;
  assign \new_[25299]_  = ~A269 & ~A267;
  assign \new_[25300]_  = \new_[25299]_  & \new_[25296]_ ;
  assign \new_[25303]_  = ~A299 & A298;
  assign \new_[25306]_  = ~A302 & A300;
  assign \new_[25307]_  = \new_[25306]_  & \new_[25303]_ ;
  assign \new_[25308]_  = \new_[25307]_  & \new_[25300]_ ;
  assign \new_[25312]_  = ~A201 & A200;
  assign \new_[25313]_  = ~A199 & \new_[25312]_ ;
  assign \new_[25316]_  = A203 & ~A202;
  assign \new_[25319]_  = A233 & ~A232;
  assign \new_[25320]_  = \new_[25319]_  & \new_[25316]_ ;
  assign \new_[25321]_  = \new_[25320]_  & \new_[25313]_ ;
  assign \new_[25324]_  = ~A236 & A234;
  assign \new_[25327]_  = ~A269 & ~A267;
  assign \new_[25328]_  = \new_[25327]_  & \new_[25324]_ ;
  assign \new_[25331]_  = A299 & ~A298;
  assign \new_[25334]_  = A301 & A300;
  assign \new_[25335]_  = \new_[25334]_  & \new_[25331]_ ;
  assign \new_[25336]_  = \new_[25335]_  & \new_[25328]_ ;
  assign \new_[25340]_  = ~A201 & A200;
  assign \new_[25341]_  = ~A199 & \new_[25340]_ ;
  assign \new_[25344]_  = A203 & ~A202;
  assign \new_[25347]_  = A233 & ~A232;
  assign \new_[25348]_  = \new_[25347]_  & \new_[25344]_ ;
  assign \new_[25349]_  = \new_[25348]_  & \new_[25341]_ ;
  assign \new_[25352]_  = ~A236 & A234;
  assign \new_[25355]_  = ~A269 & ~A267;
  assign \new_[25356]_  = \new_[25355]_  & \new_[25352]_ ;
  assign \new_[25359]_  = A299 & ~A298;
  assign \new_[25362]_  = ~A302 & A300;
  assign \new_[25363]_  = \new_[25362]_  & \new_[25359]_ ;
  assign \new_[25364]_  = \new_[25363]_  & \new_[25356]_ ;
  assign \new_[25368]_  = ~A201 & A200;
  assign \new_[25369]_  = ~A199 & \new_[25368]_ ;
  assign \new_[25372]_  = A203 & ~A202;
  assign \new_[25375]_  = A233 & ~A232;
  assign \new_[25376]_  = \new_[25375]_  & \new_[25372]_ ;
  assign \new_[25377]_  = \new_[25376]_  & \new_[25369]_ ;
  assign \new_[25380]_  = ~A236 & A234;
  assign \new_[25383]_  = A266 & A265;
  assign \new_[25384]_  = \new_[25383]_  & \new_[25380]_ ;
  assign \new_[25387]_  = ~A299 & A298;
  assign \new_[25390]_  = A301 & A300;
  assign \new_[25391]_  = \new_[25390]_  & \new_[25387]_ ;
  assign \new_[25392]_  = \new_[25391]_  & \new_[25384]_ ;
  assign \new_[25396]_  = ~A201 & A200;
  assign \new_[25397]_  = ~A199 & \new_[25396]_ ;
  assign \new_[25400]_  = A203 & ~A202;
  assign \new_[25403]_  = A233 & ~A232;
  assign \new_[25404]_  = \new_[25403]_  & \new_[25400]_ ;
  assign \new_[25405]_  = \new_[25404]_  & \new_[25397]_ ;
  assign \new_[25408]_  = ~A236 & A234;
  assign \new_[25411]_  = A266 & A265;
  assign \new_[25412]_  = \new_[25411]_  & \new_[25408]_ ;
  assign \new_[25415]_  = ~A299 & A298;
  assign \new_[25418]_  = ~A302 & A300;
  assign \new_[25419]_  = \new_[25418]_  & \new_[25415]_ ;
  assign \new_[25420]_  = \new_[25419]_  & \new_[25412]_ ;
  assign \new_[25424]_  = ~A201 & A200;
  assign \new_[25425]_  = ~A199 & \new_[25424]_ ;
  assign \new_[25428]_  = A203 & ~A202;
  assign \new_[25431]_  = A233 & ~A232;
  assign \new_[25432]_  = \new_[25431]_  & \new_[25428]_ ;
  assign \new_[25433]_  = \new_[25432]_  & \new_[25425]_ ;
  assign \new_[25436]_  = ~A236 & A234;
  assign \new_[25439]_  = A266 & A265;
  assign \new_[25440]_  = \new_[25439]_  & \new_[25436]_ ;
  assign \new_[25443]_  = A299 & ~A298;
  assign \new_[25446]_  = A301 & A300;
  assign \new_[25447]_  = \new_[25446]_  & \new_[25443]_ ;
  assign \new_[25448]_  = \new_[25447]_  & \new_[25440]_ ;
  assign \new_[25452]_  = ~A201 & A200;
  assign \new_[25453]_  = ~A199 & \new_[25452]_ ;
  assign \new_[25456]_  = A203 & ~A202;
  assign \new_[25459]_  = A233 & ~A232;
  assign \new_[25460]_  = \new_[25459]_  & \new_[25456]_ ;
  assign \new_[25461]_  = \new_[25460]_  & \new_[25453]_ ;
  assign \new_[25464]_  = ~A236 & A234;
  assign \new_[25467]_  = A266 & A265;
  assign \new_[25468]_  = \new_[25467]_  & \new_[25464]_ ;
  assign \new_[25471]_  = A299 & ~A298;
  assign \new_[25474]_  = ~A302 & A300;
  assign \new_[25475]_  = \new_[25474]_  & \new_[25471]_ ;
  assign \new_[25476]_  = \new_[25475]_  & \new_[25468]_ ;
  assign \new_[25480]_  = ~A201 & A200;
  assign \new_[25481]_  = ~A199 & \new_[25480]_ ;
  assign \new_[25484]_  = A203 & ~A202;
  assign \new_[25487]_  = A233 & ~A232;
  assign \new_[25488]_  = \new_[25487]_  & \new_[25484]_ ;
  assign \new_[25489]_  = \new_[25488]_  & \new_[25481]_ ;
  assign \new_[25492]_  = ~A236 & A234;
  assign \new_[25495]_  = ~A266 & ~A265;
  assign \new_[25496]_  = \new_[25495]_  & \new_[25492]_ ;
  assign \new_[25499]_  = ~A299 & A298;
  assign \new_[25502]_  = A301 & A300;
  assign \new_[25503]_  = \new_[25502]_  & \new_[25499]_ ;
  assign \new_[25504]_  = \new_[25503]_  & \new_[25496]_ ;
  assign \new_[25508]_  = ~A201 & A200;
  assign \new_[25509]_  = ~A199 & \new_[25508]_ ;
  assign \new_[25512]_  = A203 & ~A202;
  assign \new_[25515]_  = A233 & ~A232;
  assign \new_[25516]_  = \new_[25515]_  & \new_[25512]_ ;
  assign \new_[25517]_  = \new_[25516]_  & \new_[25509]_ ;
  assign \new_[25520]_  = ~A236 & A234;
  assign \new_[25523]_  = ~A266 & ~A265;
  assign \new_[25524]_  = \new_[25523]_  & \new_[25520]_ ;
  assign \new_[25527]_  = ~A299 & A298;
  assign \new_[25530]_  = ~A302 & A300;
  assign \new_[25531]_  = \new_[25530]_  & \new_[25527]_ ;
  assign \new_[25532]_  = \new_[25531]_  & \new_[25524]_ ;
  assign \new_[25536]_  = ~A201 & A200;
  assign \new_[25537]_  = ~A199 & \new_[25536]_ ;
  assign \new_[25540]_  = A203 & ~A202;
  assign \new_[25543]_  = A233 & ~A232;
  assign \new_[25544]_  = \new_[25543]_  & \new_[25540]_ ;
  assign \new_[25545]_  = \new_[25544]_  & \new_[25537]_ ;
  assign \new_[25548]_  = ~A236 & A234;
  assign \new_[25551]_  = ~A266 & ~A265;
  assign \new_[25552]_  = \new_[25551]_  & \new_[25548]_ ;
  assign \new_[25555]_  = A299 & ~A298;
  assign \new_[25558]_  = A301 & A300;
  assign \new_[25559]_  = \new_[25558]_  & \new_[25555]_ ;
  assign \new_[25560]_  = \new_[25559]_  & \new_[25552]_ ;
  assign \new_[25564]_  = ~A201 & A200;
  assign \new_[25565]_  = ~A199 & \new_[25564]_ ;
  assign \new_[25568]_  = A203 & ~A202;
  assign \new_[25571]_  = A233 & ~A232;
  assign \new_[25572]_  = \new_[25571]_  & \new_[25568]_ ;
  assign \new_[25573]_  = \new_[25572]_  & \new_[25565]_ ;
  assign \new_[25576]_  = ~A236 & A234;
  assign \new_[25579]_  = ~A266 & ~A265;
  assign \new_[25580]_  = \new_[25579]_  & \new_[25576]_ ;
  assign \new_[25583]_  = A299 & ~A298;
  assign \new_[25586]_  = ~A302 & A300;
  assign \new_[25587]_  = \new_[25586]_  & \new_[25583]_ ;
  assign \new_[25588]_  = \new_[25587]_  & \new_[25580]_ ;
  assign \new_[25592]_  = ~A201 & A200;
  assign \new_[25593]_  = ~A199 & \new_[25592]_ ;
  assign \new_[25596]_  = A203 & ~A202;
  assign \new_[25599]_  = ~A233 & A232;
  assign \new_[25600]_  = \new_[25599]_  & \new_[25596]_ ;
  assign \new_[25601]_  = \new_[25600]_  & \new_[25593]_ ;
  assign \new_[25604]_  = A235 & A234;
  assign \new_[25607]_  = A268 & ~A267;
  assign \new_[25608]_  = \new_[25607]_  & \new_[25604]_ ;
  assign \new_[25611]_  = ~A299 & A298;
  assign \new_[25614]_  = A301 & A300;
  assign \new_[25615]_  = \new_[25614]_  & \new_[25611]_ ;
  assign \new_[25616]_  = \new_[25615]_  & \new_[25608]_ ;
  assign \new_[25620]_  = ~A201 & A200;
  assign \new_[25621]_  = ~A199 & \new_[25620]_ ;
  assign \new_[25624]_  = A203 & ~A202;
  assign \new_[25627]_  = ~A233 & A232;
  assign \new_[25628]_  = \new_[25627]_  & \new_[25624]_ ;
  assign \new_[25629]_  = \new_[25628]_  & \new_[25621]_ ;
  assign \new_[25632]_  = A235 & A234;
  assign \new_[25635]_  = A268 & ~A267;
  assign \new_[25636]_  = \new_[25635]_  & \new_[25632]_ ;
  assign \new_[25639]_  = ~A299 & A298;
  assign \new_[25642]_  = ~A302 & A300;
  assign \new_[25643]_  = \new_[25642]_  & \new_[25639]_ ;
  assign \new_[25644]_  = \new_[25643]_  & \new_[25636]_ ;
  assign \new_[25648]_  = ~A201 & A200;
  assign \new_[25649]_  = ~A199 & \new_[25648]_ ;
  assign \new_[25652]_  = A203 & ~A202;
  assign \new_[25655]_  = ~A233 & A232;
  assign \new_[25656]_  = \new_[25655]_  & \new_[25652]_ ;
  assign \new_[25657]_  = \new_[25656]_  & \new_[25649]_ ;
  assign \new_[25660]_  = A235 & A234;
  assign \new_[25663]_  = A268 & ~A267;
  assign \new_[25664]_  = \new_[25663]_  & \new_[25660]_ ;
  assign \new_[25667]_  = A299 & ~A298;
  assign \new_[25670]_  = A301 & A300;
  assign \new_[25671]_  = \new_[25670]_  & \new_[25667]_ ;
  assign \new_[25672]_  = \new_[25671]_  & \new_[25664]_ ;
  assign \new_[25676]_  = ~A201 & A200;
  assign \new_[25677]_  = ~A199 & \new_[25676]_ ;
  assign \new_[25680]_  = A203 & ~A202;
  assign \new_[25683]_  = ~A233 & A232;
  assign \new_[25684]_  = \new_[25683]_  & \new_[25680]_ ;
  assign \new_[25685]_  = \new_[25684]_  & \new_[25677]_ ;
  assign \new_[25688]_  = A235 & A234;
  assign \new_[25691]_  = A268 & ~A267;
  assign \new_[25692]_  = \new_[25691]_  & \new_[25688]_ ;
  assign \new_[25695]_  = A299 & ~A298;
  assign \new_[25698]_  = ~A302 & A300;
  assign \new_[25699]_  = \new_[25698]_  & \new_[25695]_ ;
  assign \new_[25700]_  = \new_[25699]_  & \new_[25692]_ ;
  assign \new_[25704]_  = ~A201 & A200;
  assign \new_[25705]_  = ~A199 & \new_[25704]_ ;
  assign \new_[25708]_  = A203 & ~A202;
  assign \new_[25711]_  = ~A233 & A232;
  assign \new_[25712]_  = \new_[25711]_  & \new_[25708]_ ;
  assign \new_[25713]_  = \new_[25712]_  & \new_[25705]_ ;
  assign \new_[25716]_  = A235 & A234;
  assign \new_[25719]_  = ~A269 & ~A267;
  assign \new_[25720]_  = \new_[25719]_  & \new_[25716]_ ;
  assign \new_[25723]_  = ~A299 & A298;
  assign \new_[25726]_  = A301 & A300;
  assign \new_[25727]_  = \new_[25726]_  & \new_[25723]_ ;
  assign \new_[25728]_  = \new_[25727]_  & \new_[25720]_ ;
  assign \new_[25732]_  = ~A201 & A200;
  assign \new_[25733]_  = ~A199 & \new_[25732]_ ;
  assign \new_[25736]_  = A203 & ~A202;
  assign \new_[25739]_  = ~A233 & A232;
  assign \new_[25740]_  = \new_[25739]_  & \new_[25736]_ ;
  assign \new_[25741]_  = \new_[25740]_  & \new_[25733]_ ;
  assign \new_[25744]_  = A235 & A234;
  assign \new_[25747]_  = ~A269 & ~A267;
  assign \new_[25748]_  = \new_[25747]_  & \new_[25744]_ ;
  assign \new_[25751]_  = ~A299 & A298;
  assign \new_[25754]_  = ~A302 & A300;
  assign \new_[25755]_  = \new_[25754]_  & \new_[25751]_ ;
  assign \new_[25756]_  = \new_[25755]_  & \new_[25748]_ ;
  assign \new_[25760]_  = ~A201 & A200;
  assign \new_[25761]_  = ~A199 & \new_[25760]_ ;
  assign \new_[25764]_  = A203 & ~A202;
  assign \new_[25767]_  = ~A233 & A232;
  assign \new_[25768]_  = \new_[25767]_  & \new_[25764]_ ;
  assign \new_[25769]_  = \new_[25768]_  & \new_[25761]_ ;
  assign \new_[25772]_  = A235 & A234;
  assign \new_[25775]_  = ~A269 & ~A267;
  assign \new_[25776]_  = \new_[25775]_  & \new_[25772]_ ;
  assign \new_[25779]_  = A299 & ~A298;
  assign \new_[25782]_  = A301 & A300;
  assign \new_[25783]_  = \new_[25782]_  & \new_[25779]_ ;
  assign \new_[25784]_  = \new_[25783]_  & \new_[25776]_ ;
  assign \new_[25788]_  = ~A201 & A200;
  assign \new_[25789]_  = ~A199 & \new_[25788]_ ;
  assign \new_[25792]_  = A203 & ~A202;
  assign \new_[25795]_  = ~A233 & A232;
  assign \new_[25796]_  = \new_[25795]_  & \new_[25792]_ ;
  assign \new_[25797]_  = \new_[25796]_  & \new_[25789]_ ;
  assign \new_[25800]_  = A235 & A234;
  assign \new_[25803]_  = ~A269 & ~A267;
  assign \new_[25804]_  = \new_[25803]_  & \new_[25800]_ ;
  assign \new_[25807]_  = A299 & ~A298;
  assign \new_[25810]_  = ~A302 & A300;
  assign \new_[25811]_  = \new_[25810]_  & \new_[25807]_ ;
  assign \new_[25812]_  = \new_[25811]_  & \new_[25804]_ ;
  assign \new_[25816]_  = ~A201 & A200;
  assign \new_[25817]_  = ~A199 & \new_[25816]_ ;
  assign \new_[25820]_  = A203 & ~A202;
  assign \new_[25823]_  = ~A233 & A232;
  assign \new_[25824]_  = \new_[25823]_  & \new_[25820]_ ;
  assign \new_[25825]_  = \new_[25824]_  & \new_[25817]_ ;
  assign \new_[25828]_  = A235 & A234;
  assign \new_[25831]_  = A266 & A265;
  assign \new_[25832]_  = \new_[25831]_  & \new_[25828]_ ;
  assign \new_[25835]_  = ~A299 & A298;
  assign \new_[25838]_  = A301 & A300;
  assign \new_[25839]_  = \new_[25838]_  & \new_[25835]_ ;
  assign \new_[25840]_  = \new_[25839]_  & \new_[25832]_ ;
  assign \new_[25844]_  = ~A201 & A200;
  assign \new_[25845]_  = ~A199 & \new_[25844]_ ;
  assign \new_[25848]_  = A203 & ~A202;
  assign \new_[25851]_  = ~A233 & A232;
  assign \new_[25852]_  = \new_[25851]_  & \new_[25848]_ ;
  assign \new_[25853]_  = \new_[25852]_  & \new_[25845]_ ;
  assign \new_[25856]_  = A235 & A234;
  assign \new_[25859]_  = A266 & A265;
  assign \new_[25860]_  = \new_[25859]_  & \new_[25856]_ ;
  assign \new_[25863]_  = ~A299 & A298;
  assign \new_[25866]_  = ~A302 & A300;
  assign \new_[25867]_  = \new_[25866]_  & \new_[25863]_ ;
  assign \new_[25868]_  = \new_[25867]_  & \new_[25860]_ ;
  assign \new_[25872]_  = ~A201 & A200;
  assign \new_[25873]_  = ~A199 & \new_[25872]_ ;
  assign \new_[25876]_  = A203 & ~A202;
  assign \new_[25879]_  = ~A233 & A232;
  assign \new_[25880]_  = \new_[25879]_  & \new_[25876]_ ;
  assign \new_[25881]_  = \new_[25880]_  & \new_[25873]_ ;
  assign \new_[25884]_  = A235 & A234;
  assign \new_[25887]_  = A266 & A265;
  assign \new_[25888]_  = \new_[25887]_  & \new_[25884]_ ;
  assign \new_[25891]_  = A299 & ~A298;
  assign \new_[25894]_  = A301 & A300;
  assign \new_[25895]_  = \new_[25894]_  & \new_[25891]_ ;
  assign \new_[25896]_  = \new_[25895]_  & \new_[25888]_ ;
  assign \new_[25900]_  = ~A201 & A200;
  assign \new_[25901]_  = ~A199 & \new_[25900]_ ;
  assign \new_[25904]_  = A203 & ~A202;
  assign \new_[25907]_  = ~A233 & A232;
  assign \new_[25908]_  = \new_[25907]_  & \new_[25904]_ ;
  assign \new_[25909]_  = \new_[25908]_  & \new_[25901]_ ;
  assign \new_[25912]_  = A235 & A234;
  assign \new_[25915]_  = A266 & A265;
  assign \new_[25916]_  = \new_[25915]_  & \new_[25912]_ ;
  assign \new_[25919]_  = A299 & ~A298;
  assign \new_[25922]_  = ~A302 & A300;
  assign \new_[25923]_  = \new_[25922]_  & \new_[25919]_ ;
  assign \new_[25924]_  = \new_[25923]_  & \new_[25916]_ ;
  assign \new_[25928]_  = ~A201 & A200;
  assign \new_[25929]_  = ~A199 & \new_[25928]_ ;
  assign \new_[25932]_  = A203 & ~A202;
  assign \new_[25935]_  = ~A233 & A232;
  assign \new_[25936]_  = \new_[25935]_  & \new_[25932]_ ;
  assign \new_[25937]_  = \new_[25936]_  & \new_[25929]_ ;
  assign \new_[25940]_  = A235 & A234;
  assign \new_[25943]_  = ~A266 & ~A265;
  assign \new_[25944]_  = \new_[25943]_  & \new_[25940]_ ;
  assign \new_[25947]_  = ~A299 & A298;
  assign \new_[25950]_  = A301 & A300;
  assign \new_[25951]_  = \new_[25950]_  & \new_[25947]_ ;
  assign \new_[25952]_  = \new_[25951]_  & \new_[25944]_ ;
  assign \new_[25956]_  = ~A201 & A200;
  assign \new_[25957]_  = ~A199 & \new_[25956]_ ;
  assign \new_[25960]_  = A203 & ~A202;
  assign \new_[25963]_  = ~A233 & A232;
  assign \new_[25964]_  = \new_[25963]_  & \new_[25960]_ ;
  assign \new_[25965]_  = \new_[25964]_  & \new_[25957]_ ;
  assign \new_[25968]_  = A235 & A234;
  assign \new_[25971]_  = ~A266 & ~A265;
  assign \new_[25972]_  = \new_[25971]_  & \new_[25968]_ ;
  assign \new_[25975]_  = ~A299 & A298;
  assign \new_[25978]_  = ~A302 & A300;
  assign \new_[25979]_  = \new_[25978]_  & \new_[25975]_ ;
  assign \new_[25980]_  = \new_[25979]_  & \new_[25972]_ ;
  assign \new_[25984]_  = ~A201 & A200;
  assign \new_[25985]_  = ~A199 & \new_[25984]_ ;
  assign \new_[25988]_  = A203 & ~A202;
  assign \new_[25991]_  = ~A233 & A232;
  assign \new_[25992]_  = \new_[25991]_  & \new_[25988]_ ;
  assign \new_[25993]_  = \new_[25992]_  & \new_[25985]_ ;
  assign \new_[25996]_  = A235 & A234;
  assign \new_[25999]_  = ~A266 & ~A265;
  assign \new_[26000]_  = \new_[25999]_  & \new_[25996]_ ;
  assign \new_[26003]_  = A299 & ~A298;
  assign \new_[26006]_  = A301 & A300;
  assign \new_[26007]_  = \new_[26006]_  & \new_[26003]_ ;
  assign \new_[26008]_  = \new_[26007]_  & \new_[26000]_ ;
  assign \new_[26012]_  = ~A201 & A200;
  assign \new_[26013]_  = ~A199 & \new_[26012]_ ;
  assign \new_[26016]_  = A203 & ~A202;
  assign \new_[26019]_  = ~A233 & A232;
  assign \new_[26020]_  = \new_[26019]_  & \new_[26016]_ ;
  assign \new_[26021]_  = \new_[26020]_  & \new_[26013]_ ;
  assign \new_[26024]_  = A235 & A234;
  assign \new_[26027]_  = ~A266 & ~A265;
  assign \new_[26028]_  = \new_[26027]_  & \new_[26024]_ ;
  assign \new_[26031]_  = A299 & ~A298;
  assign \new_[26034]_  = ~A302 & A300;
  assign \new_[26035]_  = \new_[26034]_  & \new_[26031]_ ;
  assign \new_[26036]_  = \new_[26035]_  & \new_[26028]_ ;
  assign \new_[26040]_  = ~A201 & A200;
  assign \new_[26041]_  = ~A199 & \new_[26040]_ ;
  assign \new_[26044]_  = A203 & ~A202;
  assign \new_[26047]_  = ~A233 & A232;
  assign \new_[26048]_  = \new_[26047]_  & \new_[26044]_ ;
  assign \new_[26049]_  = \new_[26048]_  & \new_[26041]_ ;
  assign \new_[26052]_  = ~A236 & A234;
  assign \new_[26055]_  = A268 & ~A267;
  assign \new_[26056]_  = \new_[26055]_  & \new_[26052]_ ;
  assign \new_[26059]_  = ~A299 & A298;
  assign \new_[26062]_  = A301 & A300;
  assign \new_[26063]_  = \new_[26062]_  & \new_[26059]_ ;
  assign \new_[26064]_  = \new_[26063]_  & \new_[26056]_ ;
  assign \new_[26068]_  = ~A201 & A200;
  assign \new_[26069]_  = ~A199 & \new_[26068]_ ;
  assign \new_[26072]_  = A203 & ~A202;
  assign \new_[26075]_  = ~A233 & A232;
  assign \new_[26076]_  = \new_[26075]_  & \new_[26072]_ ;
  assign \new_[26077]_  = \new_[26076]_  & \new_[26069]_ ;
  assign \new_[26080]_  = ~A236 & A234;
  assign \new_[26083]_  = A268 & ~A267;
  assign \new_[26084]_  = \new_[26083]_  & \new_[26080]_ ;
  assign \new_[26087]_  = ~A299 & A298;
  assign \new_[26090]_  = ~A302 & A300;
  assign \new_[26091]_  = \new_[26090]_  & \new_[26087]_ ;
  assign \new_[26092]_  = \new_[26091]_  & \new_[26084]_ ;
  assign \new_[26096]_  = ~A201 & A200;
  assign \new_[26097]_  = ~A199 & \new_[26096]_ ;
  assign \new_[26100]_  = A203 & ~A202;
  assign \new_[26103]_  = ~A233 & A232;
  assign \new_[26104]_  = \new_[26103]_  & \new_[26100]_ ;
  assign \new_[26105]_  = \new_[26104]_  & \new_[26097]_ ;
  assign \new_[26108]_  = ~A236 & A234;
  assign \new_[26111]_  = A268 & ~A267;
  assign \new_[26112]_  = \new_[26111]_  & \new_[26108]_ ;
  assign \new_[26115]_  = A299 & ~A298;
  assign \new_[26118]_  = A301 & A300;
  assign \new_[26119]_  = \new_[26118]_  & \new_[26115]_ ;
  assign \new_[26120]_  = \new_[26119]_  & \new_[26112]_ ;
  assign \new_[26124]_  = ~A201 & A200;
  assign \new_[26125]_  = ~A199 & \new_[26124]_ ;
  assign \new_[26128]_  = A203 & ~A202;
  assign \new_[26131]_  = ~A233 & A232;
  assign \new_[26132]_  = \new_[26131]_  & \new_[26128]_ ;
  assign \new_[26133]_  = \new_[26132]_  & \new_[26125]_ ;
  assign \new_[26136]_  = ~A236 & A234;
  assign \new_[26139]_  = A268 & ~A267;
  assign \new_[26140]_  = \new_[26139]_  & \new_[26136]_ ;
  assign \new_[26143]_  = A299 & ~A298;
  assign \new_[26146]_  = ~A302 & A300;
  assign \new_[26147]_  = \new_[26146]_  & \new_[26143]_ ;
  assign \new_[26148]_  = \new_[26147]_  & \new_[26140]_ ;
  assign \new_[26152]_  = ~A201 & A200;
  assign \new_[26153]_  = ~A199 & \new_[26152]_ ;
  assign \new_[26156]_  = A203 & ~A202;
  assign \new_[26159]_  = ~A233 & A232;
  assign \new_[26160]_  = \new_[26159]_  & \new_[26156]_ ;
  assign \new_[26161]_  = \new_[26160]_  & \new_[26153]_ ;
  assign \new_[26164]_  = ~A236 & A234;
  assign \new_[26167]_  = ~A269 & ~A267;
  assign \new_[26168]_  = \new_[26167]_  & \new_[26164]_ ;
  assign \new_[26171]_  = ~A299 & A298;
  assign \new_[26174]_  = A301 & A300;
  assign \new_[26175]_  = \new_[26174]_  & \new_[26171]_ ;
  assign \new_[26176]_  = \new_[26175]_  & \new_[26168]_ ;
  assign \new_[26180]_  = ~A201 & A200;
  assign \new_[26181]_  = ~A199 & \new_[26180]_ ;
  assign \new_[26184]_  = A203 & ~A202;
  assign \new_[26187]_  = ~A233 & A232;
  assign \new_[26188]_  = \new_[26187]_  & \new_[26184]_ ;
  assign \new_[26189]_  = \new_[26188]_  & \new_[26181]_ ;
  assign \new_[26192]_  = ~A236 & A234;
  assign \new_[26195]_  = ~A269 & ~A267;
  assign \new_[26196]_  = \new_[26195]_  & \new_[26192]_ ;
  assign \new_[26199]_  = ~A299 & A298;
  assign \new_[26202]_  = ~A302 & A300;
  assign \new_[26203]_  = \new_[26202]_  & \new_[26199]_ ;
  assign \new_[26204]_  = \new_[26203]_  & \new_[26196]_ ;
  assign \new_[26208]_  = ~A201 & A200;
  assign \new_[26209]_  = ~A199 & \new_[26208]_ ;
  assign \new_[26212]_  = A203 & ~A202;
  assign \new_[26215]_  = ~A233 & A232;
  assign \new_[26216]_  = \new_[26215]_  & \new_[26212]_ ;
  assign \new_[26217]_  = \new_[26216]_  & \new_[26209]_ ;
  assign \new_[26220]_  = ~A236 & A234;
  assign \new_[26223]_  = ~A269 & ~A267;
  assign \new_[26224]_  = \new_[26223]_  & \new_[26220]_ ;
  assign \new_[26227]_  = A299 & ~A298;
  assign \new_[26230]_  = A301 & A300;
  assign \new_[26231]_  = \new_[26230]_  & \new_[26227]_ ;
  assign \new_[26232]_  = \new_[26231]_  & \new_[26224]_ ;
  assign \new_[26236]_  = ~A201 & A200;
  assign \new_[26237]_  = ~A199 & \new_[26236]_ ;
  assign \new_[26240]_  = A203 & ~A202;
  assign \new_[26243]_  = ~A233 & A232;
  assign \new_[26244]_  = \new_[26243]_  & \new_[26240]_ ;
  assign \new_[26245]_  = \new_[26244]_  & \new_[26237]_ ;
  assign \new_[26248]_  = ~A236 & A234;
  assign \new_[26251]_  = ~A269 & ~A267;
  assign \new_[26252]_  = \new_[26251]_  & \new_[26248]_ ;
  assign \new_[26255]_  = A299 & ~A298;
  assign \new_[26258]_  = ~A302 & A300;
  assign \new_[26259]_  = \new_[26258]_  & \new_[26255]_ ;
  assign \new_[26260]_  = \new_[26259]_  & \new_[26252]_ ;
  assign \new_[26264]_  = ~A201 & A200;
  assign \new_[26265]_  = ~A199 & \new_[26264]_ ;
  assign \new_[26268]_  = A203 & ~A202;
  assign \new_[26271]_  = ~A233 & A232;
  assign \new_[26272]_  = \new_[26271]_  & \new_[26268]_ ;
  assign \new_[26273]_  = \new_[26272]_  & \new_[26265]_ ;
  assign \new_[26276]_  = ~A236 & A234;
  assign \new_[26279]_  = A266 & A265;
  assign \new_[26280]_  = \new_[26279]_  & \new_[26276]_ ;
  assign \new_[26283]_  = ~A299 & A298;
  assign \new_[26286]_  = A301 & A300;
  assign \new_[26287]_  = \new_[26286]_  & \new_[26283]_ ;
  assign \new_[26288]_  = \new_[26287]_  & \new_[26280]_ ;
  assign \new_[26292]_  = ~A201 & A200;
  assign \new_[26293]_  = ~A199 & \new_[26292]_ ;
  assign \new_[26296]_  = A203 & ~A202;
  assign \new_[26299]_  = ~A233 & A232;
  assign \new_[26300]_  = \new_[26299]_  & \new_[26296]_ ;
  assign \new_[26301]_  = \new_[26300]_  & \new_[26293]_ ;
  assign \new_[26304]_  = ~A236 & A234;
  assign \new_[26307]_  = A266 & A265;
  assign \new_[26308]_  = \new_[26307]_  & \new_[26304]_ ;
  assign \new_[26311]_  = ~A299 & A298;
  assign \new_[26314]_  = ~A302 & A300;
  assign \new_[26315]_  = \new_[26314]_  & \new_[26311]_ ;
  assign \new_[26316]_  = \new_[26315]_  & \new_[26308]_ ;
  assign \new_[26320]_  = ~A201 & A200;
  assign \new_[26321]_  = ~A199 & \new_[26320]_ ;
  assign \new_[26324]_  = A203 & ~A202;
  assign \new_[26327]_  = ~A233 & A232;
  assign \new_[26328]_  = \new_[26327]_  & \new_[26324]_ ;
  assign \new_[26329]_  = \new_[26328]_  & \new_[26321]_ ;
  assign \new_[26332]_  = ~A236 & A234;
  assign \new_[26335]_  = A266 & A265;
  assign \new_[26336]_  = \new_[26335]_  & \new_[26332]_ ;
  assign \new_[26339]_  = A299 & ~A298;
  assign \new_[26342]_  = A301 & A300;
  assign \new_[26343]_  = \new_[26342]_  & \new_[26339]_ ;
  assign \new_[26344]_  = \new_[26343]_  & \new_[26336]_ ;
  assign \new_[26348]_  = ~A201 & A200;
  assign \new_[26349]_  = ~A199 & \new_[26348]_ ;
  assign \new_[26352]_  = A203 & ~A202;
  assign \new_[26355]_  = ~A233 & A232;
  assign \new_[26356]_  = \new_[26355]_  & \new_[26352]_ ;
  assign \new_[26357]_  = \new_[26356]_  & \new_[26349]_ ;
  assign \new_[26360]_  = ~A236 & A234;
  assign \new_[26363]_  = A266 & A265;
  assign \new_[26364]_  = \new_[26363]_  & \new_[26360]_ ;
  assign \new_[26367]_  = A299 & ~A298;
  assign \new_[26370]_  = ~A302 & A300;
  assign \new_[26371]_  = \new_[26370]_  & \new_[26367]_ ;
  assign \new_[26372]_  = \new_[26371]_  & \new_[26364]_ ;
  assign \new_[26376]_  = ~A201 & A200;
  assign \new_[26377]_  = ~A199 & \new_[26376]_ ;
  assign \new_[26380]_  = A203 & ~A202;
  assign \new_[26383]_  = ~A233 & A232;
  assign \new_[26384]_  = \new_[26383]_  & \new_[26380]_ ;
  assign \new_[26385]_  = \new_[26384]_  & \new_[26377]_ ;
  assign \new_[26388]_  = ~A236 & A234;
  assign \new_[26391]_  = ~A266 & ~A265;
  assign \new_[26392]_  = \new_[26391]_  & \new_[26388]_ ;
  assign \new_[26395]_  = ~A299 & A298;
  assign \new_[26398]_  = A301 & A300;
  assign \new_[26399]_  = \new_[26398]_  & \new_[26395]_ ;
  assign \new_[26400]_  = \new_[26399]_  & \new_[26392]_ ;
  assign \new_[26404]_  = ~A201 & A200;
  assign \new_[26405]_  = ~A199 & \new_[26404]_ ;
  assign \new_[26408]_  = A203 & ~A202;
  assign \new_[26411]_  = ~A233 & A232;
  assign \new_[26412]_  = \new_[26411]_  & \new_[26408]_ ;
  assign \new_[26413]_  = \new_[26412]_  & \new_[26405]_ ;
  assign \new_[26416]_  = ~A236 & A234;
  assign \new_[26419]_  = ~A266 & ~A265;
  assign \new_[26420]_  = \new_[26419]_  & \new_[26416]_ ;
  assign \new_[26423]_  = ~A299 & A298;
  assign \new_[26426]_  = ~A302 & A300;
  assign \new_[26427]_  = \new_[26426]_  & \new_[26423]_ ;
  assign \new_[26428]_  = \new_[26427]_  & \new_[26420]_ ;
  assign \new_[26432]_  = ~A201 & A200;
  assign \new_[26433]_  = ~A199 & \new_[26432]_ ;
  assign \new_[26436]_  = A203 & ~A202;
  assign \new_[26439]_  = ~A233 & A232;
  assign \new_[26440]_  = \new_[26439]_  & \new_[26436]_ ;
  assign \new_[26441]_  = \new_[26440]_  & \new_[26433]_ ;
  assign \new_[26444]_  = ~A236 & A234;
  assign \new_[26447]_  = ~A266 & ~A265;
  assign \new_[26448]_  = \new_[26447]_  & \new_[26444]_ ;
  assign \new_[26451]_  = A299 & ~A298;
  assign \new_[26454]_  = A301 & A300;
  assign \new_[26455]_  = \new_[26454]_  & \new_[26451]_ ;
  assign \new_[26456]_  = \new_[26455]_  & \new_[26448]_ ;
  assign \new_[26460]_  = ~A201 & A200;
  assign \new_[26461]_  = ~A199 & \new_[26460]_ ;
  assign \new_[26464]_  = A203 & ~A202;
  assign \new_[26467]_  = ~A233 & A232;
  assign \new_[26468]_  = \new_[26467]_  & \new_[26464]_ ;
  assign \new_[26469]_  = \new_[26468]_  & \new_[26461]_ ;
  assign \new_[26472]_  = ~A236 & A234;
  assign \new_[26475]_  = ~A266 & ~A265;
  assign \new_[26476]_  = \new_[26475]_  & \new_[26472]_ ;
  assign \new_[26479]_  = A299 & ~A298;
  assign \new_[26482]_  = ~A302 & A300;
  assign \new_[26483]_  = \new_[26482]_  & \new_[26479]_ ;
  assign \new_[26484]_  = \new_[26483]_  & \new_[26476]_ ;
  assign \new_[26488]_  = A201 & ~A200;
  assign \new_[26489]_  = A199 & \new_[26488]_ ;
  assign \new_[26492]_  = ~A232 & A202;
  assign \new_[26495]_  = A234 & A233;
  assign \new_[26496]_  = \new_[26495]_  & \new_[26492]_ ;
  assign \new_[26497]_  = \new_[26496]_  & \new_[26489]_ ;
  assign \new_[26500]_  = A267 & A235;
  assign \new_[26503]_  = A269 & ~A268;
  assign \new_[26504]_  = \new_[26503]_  & \new_[26500]_ ;
  assign \new_[26507]_  = ~A299 & A298;
  assign \new_[26510]_  = A301 & A300;
  assign \new_[26511]_  = \new_[26510]_  & \new_[26507]_ ;
  assign \new_[26512]_  = \new_[26511]_  & \new_[26504]_ ;
  assign \new_[26516]_  = A201 & ~A200;
  assign \new_[26517]_  = A199 & \new_[26516]_ ;
  assign \new_[26520]_  = ~A232 & A202;
  assign \new_[26523]_  = A234 & A233;
  assign \new_[26524]_  = \new_[26523]_  & \new_[26520]_ ;
  assign \new_[26525]_  = \new_[26524]_  & \new_[26517]_ ;
  assign \new_[26528]_  = A267 & A235;
  assign \new_[26531]_  = A269 & ~A268;
  assign \new_[26532]_  = \new_[26531]_  & \new_[26528]_ ;
  assign \new_[26535]_  = ~A299 & A298;
  assign \new_[26538]_  = ~A302 & A300;
  assign \new_[26539]_  = \new_[26538]_  & \new_[26535]_ ;
  assign \new_[26540]_  = \new_[26539]_  & \new_[26532]_ ;
  assign \new_[26544]_  = A201 & ~A200;
  assign \new_[26545]_  = A199 & \new_[26544]_ ;
  assign \new_[26548]_  = ~A232 & A202;
  assign \new_[26551]_  = A234 & A233;
  assign \new_[26552]_  = \new_[26551]_  & \new_[26548]_ ;
  assign \new_[26553]_  = \new_[26552]_  & \new_[26545]_ ;
  assign \new_[26556]_  = A267 & A235;
  assign \new_[26559]_  = A269 & ~A268;
  assign \new_[26560]_  = \new_[26559]_  & \new_[26556]_ ;
  assign \new_[26563]_  = A299 & ~A298;
  assign \new_[26566]_  = A301 & A300;
  assign \new_[26567]_  = \new_[26566]_  & \new_[26563]_ ;
  assign \new_[26568]_  = \new_[26567]_  & \new_[26560]_ ;
  assign \new_[26572]_  = A201 & ~A200;
  assign \new_[26573]_  = A199 & \new_[26572]_ ;
  assign \new_[26576]_  = ~A232 & A202;
  assign \new_[26579]_  = A234 & A233;
  assign \new_[26580]_  = \new_[26579]_  & \new_[26576]_ ;
  assign \new_[26581]_  = \new_[26580]_  & \new_[26573]_ ;
  assign \new_[26584]_  = A267 & A235;
  assign \new_[26587]_  = A269 & ~A268;
  assign \new_[26588]_  = \new_[26587]_  & \new_[26584]_ ;
  assign \new_[26591]_  = A299 & ~A298;
  assign \new_[26594]_  = ~A302 & A300;
  assign \new_[26595]_  = \new_[26594]_  & \new_[26591]_ ;
  assign \new_[26596]_  = \new_[26595]_  & \new_[26588]_ ;
  assign \new_[26600]_  = A201 & ~A200;
  assign \new_[26601]_  = A199 & \new_[26600]_ ;
  assign \new_[26604]_  = ~A232 & A202;
  assign \new_[26607]_  = A234 & A233;
  assign \new_[26608]_  = \new_[26607]_  & \new_[26604]_ ;
  assign \new_[26609]_  = \new_[26608]_  & \new_[26601]_ ;
  assign \new_[26612]_  = ~A267 & A235;
  assign \new_[26615]_  = A298 & A268;
  assign \new_[26616]_  = \new_[26615]_  & \new_[26612]_ ;
  assign \new_[26619]_  = ~A300 & ~A299;
  assign \new_[26622]_  = A302 & ~A301;
  assign \new_[26623]_  = \new_[26622]_  & \new_[26619]_ ;
  assign \new_[26624]_  = \new_[26623]_  & \new_[26616]_ ;
  assign \new_[26628]_  = A201 & ~A200;
  assign \new_[26629]_  = A199 & \new_[26628]_ ;
  assign \new_[26632]_  = ~A232 & A202;
  assign \new_[26635]_  = A234 & A233;
  assign \new_[26636]_  = \new_[26635]_  & \new_[26632]_ ;
  assign \new_[26637]_  = \new_[26636]_  & \new_[26629]_ ;
  assign \new_[26640]_  = ~A267 & A235;
  assign \new_[26643]_  = ~A298 & A268;
  assign \new_[26644]_  = \new_[26643]_  & \new_[26640]_ ;
  assign \new_[26647]_  = ~A300 & A299;
  assign \new_[26650]_  = A302 & ~A301;
  assign \new_[26651]_  = \new_[26650]_  & \new_[26647]_ ;
  assign \new_[26652]_  = \new_[26651]_  & \new_[26644]_ ;
  assign \new_[26656]_  = A201 & ~A200;
  assign \new_[26657]_  = A199 & \new_[26656]_ ;
  assign \new_[26660]_  = ~A232 & A202;
  assign \new_[26663]_  = A234 & A233;
  assign \new_[26664]_  = \new_[26663]_  & \new_[26660]_ ;
  assign \new_[26665]_  = \new_[26664]_  & \new_[26657]_ ;
  assign \new_[26668]_  = ~A267 & A235;
  assign \new_[26671]_  = A298 & ~A269;
  assign \new_[26672]_  = \new_[26671]_  & \new_[26668]_ ;
  assign \new_[26675]_  = ~A300 & ~A299;
  assign \new_[26678]_  = A302 & ~A301;
  assign \new_[26679]_  = \new_[26678]_  & \new_[26675]_ ;
  assign \new_[26680]_  = \new_[26679]_  & \new_[26672]_ ;
  assign \new_[26684]_  = A201 & ~A200;
  assign \new_[26685]_  = A199 & \new_[26684]_ ;
  assign \new_[26688]_  = ~A232 & A202;
  assign \new_[26691]_  = A234 & A233;
  assign \new_[26692]_  = \new_[26691]_  & \new_[26688]_ ;
  assign \new_[26693]_  = \new_[26692]_  & \new_[26685]_ ;
  assign \new_[26696]_  = ~A267 & A235;
  assign \new_[26699]_  = ~A298 & ~A269;
  assign \new_[26700]_  = \new_[26699]_  & \new_[26696]_ ;
  assign \new_[26703]_  = ~A300 & A299;
  assign \new_[26706]_  = A302 & ~A301;
  assign \new_[26707]_  = \new_[26706]_  & \new_[26703]_ ;
  assign \new_[26708]_  = \new_[26707]_  & \new_[26700]_ ;
  assign \new_[26712]_  = A201 & ~A200;
  assign \new_[26713]_  = A199 & \new_[26712]_ ;
  assign \new_[26716]_  = ~A232 & A202;
  assign \new_[26719]_  = A234 & A233;
  assign \new_[26720]_  = \new_[26719]_  & \new_[26716]_ ;
  assign \new_[26721]_  = \new_[26720]_  & \new_[26713]_ ;
  assign \new_[26724]_  = A265 & A235;
  assign \new_[26727]_  = A298 & A266;
  assign \new_[26728]_  = \new_[26727]_  & \new_[26724]_ ;
  assign \new_[26731]_  = ~A300 & ~A299;
  assign \new_[26734]_  = A302 & ~A301;
  assign \new_[26735]_  = \new_[26734]_  & \new_[26731]_ ;
  assign \new_[26736]_  = \new_[26735]_  & \new_[26728]_ ;
  assign \new_[26740]_  = A201 & ~A200;
  assign \new_[26741]_  = A199 & \new_[26740]_ ;
  assign \new_[26744]_  = ~A232 & A202;
  assign \new_[26747]_  = A234 & A233;
  assign \new_[26748]_  = \new_[26747]_  & \new_[26744]_ ;
  assign \new_[26749]_  = \new_[26748]_  & \new_[26741]_ ;
  assign \new_[26752]_  = A265 & A235;
  assign \new_[26755]_  = ~A298 & A266;
  assign \new_[26756]_  = \new_[26755]_  & \new_[26752]_ ;
  assign \new_[26759]_  = ~A300 & A299;
  assign \new_[26762]_  = A302 & ~A301;
  assign \new_[26763]_  = \new_[26762]_  & \new_[26759]_ ;
  assign \new_[26764]_  = \new_[26763]_  & \new_[26756]_ ;
  assign \new_[26768]_  = A201 & ~A200;
  assign \new_[26769]_  = A199 & \new_[26768]_ ;
  assign \new_[26772]_  = ~A232 & A202;
  assign \new_[26775]_  = A234 & A233;
  assign \new_[26776]_  = \new_[26775]_  & \new_[26772]_ ;
  assign \new_[26777]_  = \new_[26776]_  & \new_[26769]_ ;
  assign \new_[26780]_  = ~A265 & A235;
  assign \new_[26783]_  = A298 & ~A266;
  assign \new_[26784]_  = \new_[26783]_  & \new_[26780]_ ;
  assign \new_[26787]_  = ~A300 & ~A299;
  assign \new_[26790]_  = A302 & ~A301;
  assign \new_[26791]_  = \new_[26790]_  & \new_[26787]_ ;
  assign \new_[26792]_  = \new_[26791]_  & \new_[26784]_ ;
  assign \new_[26796]_  = A201 & ~A200;
  assign \new_[26797]_  = A199 & \new_[26796]_ ;
  assign \new_[26800]_  = ~A232 & A202;
  assign \new_[26803]_  = A234 & A233;
  assign \new_[26804]_  = \new_[26803]_  & \new_[26800]_ ;
  assign \new_[26805]_  = \new_[26804]_  & \new_[26797]_ ;
  assign \new_[26808]_  = ~A265 & A235;
  assign \new_[26811]_  = ~A298 & ~A266;
  assign \new_[26812]_  = \new_[26811]_  & \new_[26808]_ ;
  assign \new_[26815]_  = ~A300 & A299;
  assign \new_[26818]_  = A302 & ~A301;
  assign \new_[26819]_  = \new_[26818]_  & \new_[26815]_ ;
  assign \new_[26820]_  = \new_[26819]_  & \new_[26812]_ ;
  assign \new_[26824]_  = A201 & ~A200;
  assign \new_[26825]_  = A199 & \new_[26824]_ ;
  assign \new_[26828]_  = ~A232 & A202;
  assign \new_[26831]_  = A234 & A233;
  assign \new_[26832]_  = \new_[26831]_  & \new_[26828]_ ;
  assign \new_[26833]_  = \new_[26832]_  & \new_[26825]_ ;
  assign \new_[26836]_  = A267 & ~A236;
  assign \new_[26839]_  = A269 & ~A268;
  assign \new_[26840]_  = \new_[26839]_  & \new_[26836]_ ;
  assign \new_[26843]_  = ~A299 & A298;
  assign \new_[26846]_  = A301 & A300;
  assign \new_[26847]_  = \new_[26846]_  & \new_[26843]_ ;
  assign \new_[26848]_  = \new_[26847]_  & \new_[26840]_ ;
  assign \new_[26852]_  = A201 & ~A200;
  assign \new_[26853]_  = A199 & \new_[26852]_ ;
  assign \new_[26856]_  = ~A232 & A202;
  assign \new_[26859]_  = A234 & A233;
  assign \new_[26860]_  = \new_[26859]_  & \new_[26856]_ ;
  assign \new_[26861]_  = \new_[26860]_  & \new_[26853]_ ;
  assign \new_[26864]_  = A267 & ~A236;
  assign \new_[26867]_  = A269 & ~A268;
  assign \new_[26868]_  = \new_[26867]_  & \new_[26864]_ ;
  assign \new_[26871]_  = ~A299 & A298;
  assign \new_[26874]_  = ~A302 & A300;
  assign \new_[26875]_  = \new_[26874]_  & \new_[26871]_ ;
  assign \new_[26876]_  = \new_[26875]_  & \new_[26868]_ ;
  assign \new_[26880]_  = A201 & ~A200;
  assign \new_[26881]_  = A199 & \new_[26880]_ ;
  assign \new_[26884]_  = ~A232 & A202;
  assign \new_[26887]_  = A234 & A233;
  assign \new_[26888]_  = \new_[26887]_  & \new_[26884]_ ;
  assign \new_[26889]_  = \new_[26888]_  & \new_[26881]_ ;
  assign \new_[26892]_  = A267 & ~A236;
  assign \new_[26895]_  = A269 & ~A268;
  assign \new_[26896]_  = \new_[26895]_  & \new_[26892]_ ;
  assign \new_[26899]_  = A299 & ~A298;
  assign \new_[26902]_  = A301 & A300;
  assign \new_[26903]_  = \new_[26902]_  & \new_[26899]_ ;
  assign \new_[26904]_  = \new_[26903]_  & \new_[26896]_ ;
  assign \new_[26908]_  = A201 & ~A200;
  assign \new_[26909]_  = A199 & \new_[26908]_ ;
  assign \new_[26912]_  = ~A232 & A202;
  assign \new_[26915]_  = A234 & A233;
  assign \new_[26916]_  = \new_[26915]_  & \new_[26912]_ ;
  assign \new_[26917]_  = \new_[26916]_  & \new_[26909]_ ;
  assign \new_[26920]_  = A267 & ~A236;
  assign \new_[26923]_  = A269 & ~A268;
  assign \new_[26924]_  = \new_[26923]_  & \new_[26920]_ ;
  assign \new_[26927]_  = A299 & ~A298;
  assign \new_[26930]_  = ~A302 & A300;
  assign \new_[26931]_  = \new_[26930]_  & \new_[26927]_ ;
  assign \new_[26932]_  = \new_[26931]_  & \new_[26924]_ ;
  assign \new_[26936]_  = A201 & ~A200;
  assign \new_[26937]_  = A199 & \new_[26936]_ ;
  assign \new_[26940]_  = ~A232 & A202;
  assign \new_[26943]_  = A234 & A233;
  assign \new_[26944]_  = \new_[26943]_  & \new_[26940]_ ;
  assign \new_[26945]_  = \new_[26944]_  & \new_[26937]_ ;
  assign \new_[26948]_  = ~A267 & ~A236;
  assign \new_[26951]_  = A298 & A268;
  assign \new_[26952]_  = \new_[26951]_  & \new_[26948]_ ;
  assign \new_[26955]_  = ~A300 & ~A299;
  assign \new_[26958]_  = A302 & ~A301;
  assign \new_[26959]_  = \new_[26958]_  & \new_[26955]_ ;
  assign \new_[26960]_  = \new_[26959]_  & \new_[26952]_ ;
  assign \new_[26964]_  = A201 & ~A200;
  assign \new_[26965]_  = A199 & \new_[26964]_ ;
  assign \new_[26968]_  = ~A232 & A202;
  assign \new_[26971]_  = A234 & A233;
  assign \new_[26972]_  = \new_[26971]_  & \new_[26968]_ ;
  assign \new_[26973]_  = \new_[26972]_  & \new_[26965]_ ;
  assign \new_[26976]_  = ~A267 & ~A236;
  assign \new_[26979]_  = ~A298 & A268;
  assign \new_[26980]_  = \new_[26979]_  & \new_[26976]_ ;
  assign \new_[26983]_  = ~A300 & A299;
  assign \new_[26986]_  = A302 & ~A301;
  assign \new_[26987]_  = \new_[26986]_  & \new_[26983]_ ;
  assign \new_[26988]_  = \new_[26987]_  & \new_[26980]_ ;
  assign \new_[26992]_  = A201 & ~A200;
  assign \new_[26993]_  = A199 & \new_[26992]_ ;
  assign \new_[26996]_  = ~A232 & A202;
  assign \new_[26999]_  = A234 & A233;
  assign \new_[27000]_  = \new_[26999]_  & \new_[26996]_ ;
  assign \new_[27001]_  = \new_[27000]_  & \new_[26993]_ ;
  assign \new_[27004]_  = ~A267 & ~A236;
  assign \new_[27007]_  = A298 & ~A269;
  assign \new_[27008]_  = \new_[27007]_  & \new_[27004]_ ;
  assign \new_[27011]_  = ~A300 & ~A299;
  assign \new_[27014]_  = A302 & ~A301;
  assign \new_[27015]_  = \new_[27014]_  & \new_[27011]_ ;
  assign \new_[27016]_  = \new_[27015]_  & \new_[27008]_ ;
  assign \new_[27020]_  = A201 & ~A200;
  assign \new_[27021]_  = A199 & \new_[27020]_ ;
  assign \new_[27024]_  = ~A232 & A202;
  assign \new_[27027]_  = A234 & A233;
  assign \new_[27028]_  = \new_[27027]_  & \new_[27024]_ ;
  assign \new_[27029]_  = \new_[27028]_  & \new_[27021]_ ;
  assign \new_[27032]_  = ~A267 & ~A236;
  assign \new_[27035]_  = ~A298 & ~A269;
  assign \new_[27036]_  = \new_[27035]_  & \new_[27032]_ ;
  assign \new_[27039]_  = ~A300 & A299;
  assign \new_[27042]_  = A302 & ~A301;
  assign \new_[27043]_  = \new_[27042]_  & \new_[27039]_ ;
  assign \new_[27044]_  = \new_[27043]_  & \new_[27036]_ ;
  assign \new_[27048]_  = A201 & ~A200;
  assign \new_[27049]_  = A199 & \new_[27048]_ ;
  assign \new_[27052]_  = ~A232 & A202;
  assign \new_[27055]_  = A234 & A233;
  assign \new_[27056]_  = \new_[27055]_  & \new_[27052]_ ;
  assign \new_[27057]_  = \new_[27056]_  & \new_[27049]_ ;
  assign \new_[27060]_  = A265 & ~A236;
  assign \new_[27063]_  = A298 & A266;
  assign \new_[27064]_  = \new_[27063]_  & \new_[27060]_ ;
  assign \new_[27067]_  = ~A300 & ~A299;
  assign \new_[27070]_  = A302 & ~A301;
  assign \new_[27071]_  = \new_[27070]_  & \new_[27067]_ ;
  assign \new_[27072]_  = \new_[27071]_  & \new_[27064]_ ;
  assign \new_[27076]_  = A201 & ~A200;
  assign \new_[27077]_  = A199 & \new_[27076]_ ;
  assign \new_[27080]_  = ~A232 & A202;
  assign \new_[27083]_  = A234 & A233;
  assign \new_[27084]_  = \new_[27083]_  & \new_[27080]_ ;
  assign \new_[27085]_  = \new_[27084]_  & \new_[27077]_ ;
  assign \new_[27088]_  = A265 & ~A236;
  assign \new_[27091]_  = ~A298 & A266;
  assign \new_[27092]_  = \new_[27091]_  & \new_[27088]_ ;
  assign \new_[27095]_  = ~A300 & A299;
  assign \new_[27098]_  = A302 & ~A301;
  assign \new_[27099]_  = \new_[27098]_  & \new_[27095]_ ;
  assign \new_[27100]_  = \new_[27099]_  & \new_[27092]_ ;
  assign \new_[27104]_  = A201 & ~A200;
  assign \new_[27105]_  = A199 & \new_[27104]_ ;
  assign \new_[27108]_  = ~A232 & A202;
  assign \new_[27111]_  = A234 & A233;
  assign \new_[27112]_  = \new_[27111]_  & \new_[27108]_ ;
  assign \new_[27113]_  = \new_[27112]_  & \new_[27105]_ ;
  assign \new_[27116]_  = ~A265 & ~A236;
  assign \new_[27119]_  = A298 & ~A266;
  assign \new_[27120]_  = \new_[27119]_  & \new_[27116]_ ;
  assign \new_[27123]_  = ~A300 & ~A299;
  assign \new_[27126]_  = A302 & ~A301;
  assign \new_[27127]_  = \new_[27126]_  & \new_[27123]_ ;
  assign \new_[27128]_  = \new_[27127]_  & \new_[27120]_ ;
  assign \new_[27132]_  = A201 & ~A200;
  assign \new_[27133]_  = A199 & \new_[27132]_ ;
  assign \new_[27136]_  = ~A232 & A202;
  assign \new_[27139]_  = A234 & A233;
  assign \new_[27140]_  = \new_[27139]_  & \new_[27136]_ ;
  assign \new_[27141]_  = \new_[27140]_  & \new_[27133]_ ;
  assign \new_[27144]_  = ~A265 & ~A236;
  assign \new_[27147]_  = ~A298 & ~A266;
  assign \new_[27148]_  = \new_[27147]_  & \new_[27144]_ ;
  assign \new_[27151]_  = ~A300 & A299;
  assign \new_[27154]_  = A302 & ~A301;
  assign \new_[27155]_  = \new_[27154]_  & \new_[27151]_ ;
  assign \new_[27156]_  = \new_[27155]_  & \new_[27148]_ ;
  assign \new_[27160]_  = A201 & ~A200;
  assign \new_[27161]_  = A199 & \new_[27160]_ ;
  assign \new_[27164]_  = ~A232 & A202;
  assign \new_[27167]_  = ~A234 & A233;
  assign \new_[27168]_  = \new_[27167]_  & \new_[27164]_ ;
  assign \new_[27169]_  = \new_[27168]_  & \new_[27161]_ ;
  assign \new_[27172]_  = A236 & ~A235;
  assign \new_[27175]_  = A268 & ~A267;
  assign \new_[27176]_  = \new_[27175]_  & \new_[27172]_ ;
  assign \new_[27179]_  = ~A299 & A298;
  assign \new_[27182]_  = A301 & A300;
  assign \new_[27183]_  = \new_[27182]_  & \new_[27179]_ ;
  assign \new_[27184]_  = \new_[27183]_  & \new_[27176]_ ;
  assign \new_[27188]_  = A201 & ~A200;
  assign \new_[27189]_  = A199 & \new_[27188]_ ;
  assign \new_[27192]_  = ~A232 & A202;
  assign \new_[27195]_  = ~A234 & A233;
  assign \new_[27196]_  = \new_[27195]_  & \new_[27192]_ ;
  assign \new_[27197]_  = \new_[27196]_  & \new_[27189]_ ;
  assign \new_[27200]_  = A236 & ~A235;
  assign \new_[27203]_  = A268 & ~A267;
  assign \new_[27204]_  = \new_[27203]_  & \new_[27200]_ ;
  assign \new_[27207]_  = ~A299 & A298;
  assign \new_[27210]_  = ~A302 & A300;
  assign \new_[27211]_  = \new_[27210]_  & \new_[27207]_ ;
  assign \new_[27212]_  = \new_[27211]_  & \new_[27204]_ ;
  assign \new_[27216]_  = A201 & ~A200;
  assign \new_[27217]_  = A199 & \new_[27216]_ ;
  assign \new_[27220]_  = ~A232 & A202;
  assign \new_[27223]_  = ~A234 & A233;
  assign \new_[27224]_  = \new_[27223]_  & \new_[27220]_ ;
  assign \new_[27225]_  = \new_[27224]_  & \new_[27217]_ ;
  assign \new_[27228]_  = A236 & ~A235;
  assign \new_[27231]_  = A268 & ~A267;
  assign \new_[27232]_  = \new_[27231]_  & \new_[27228]_ ;
  assign \new_[27235]_  = A299 & ~A298;
  assign \new_[27238]_  = A301 & A300;
  assign \new_[27239]_  = \new_[27238]_  & \new_[27235]_ ;
  assign \new_[27240]_  = \new_[27239]_  & \new_[27232]_ ;
  assign \new_[27244]_  = A201 & ~A200;
  assign \new_[27245]_  = A199 & \new_[27244]_ ;
  assign \new_[27248]_  = ~A232 & A202;
  assign \new_[27251]_  = ~A234 & A233;
  assign \new_[27252]_  = \new_[27251]_  & \new_[27248]_ ;
  assign \new_[27253]_  = \new_[27252]_  & \new_[27245]_ ;
  assign \new_[27256]_  = A236 & ~A235;
  assign \new_[27259]_  = A268 & ~A267;
  assign \new_[27260]_  = \new_[27259]_  & \new_[27256]_ ;
  assign \new_[27263]_  = A299 & ~A298;
  assign \new_[27266]_  = ~A302 & A300;
  assign \new_[27267]_  = \new_[27266]_  & \new_[27263]_ ;
  assign \new_[27268]_  = \new_[27267]_  & \new_[27260]_ ;
  assign \new_[27272]_  = A201 & ~A200;
  assign \new_[27273]_  = A199 & \new_[27272]_ ;
  assign \new_[27276]_  = ~A232 & A202;
  assign \new_[27279]_  = ~A234 & A233;
  assign \new_[27280]_  = \new_[27279]_  & \new_[27276]_ ;
  assign \new_[27281]_  = \new_[27280]_  & \new_[27273]_ ;
  assign \new_[27284]_  = A236 & ~A235;
  assign \new_[27287]_  = ~A269 & ~A267;
  assign \new_[27288]_  = \new_[27287]_  & \new_[27284]_ ;
  assign \new_[27291]_  = ~A299 & A298;
  assign \new_[27294]_  = A301 & A300;
  assign \new_[27295]_  = \new_[27294]_  & \new_[27291]_ ;
  assign \new_[27296]_  = \new_[27295]_  & \new_[27288]_ ;
  assign \new_[27300]_  = A201 & ~A200;
  assign \new_[27301]_  = A199 & \new_[27300]_ ;
  assign \new_[27304]_  = ~A232 & A202;
  assign \new_[27307]_  = ~A234 & A233;
  assign \new_[27308]_  = \new_[27307]_  & \new_[27304]_ ;
  assign \new_[27309]_  = \new_[27308]_  & \new_[27301]_ ;
  assign \new_[27312]_  = A236 & ~A235;
  assign \new_[27315]_  = ~A269 & ~A267;
  assign \new_[27316]_  = \new_[27315]_  & \new_[27312]_ ;
  assign \new_[27319]_  = ~A299 & A298;
  assign \new_[27322]_  = ~A302 & A300;
  assign \new_[27323]_  = \new_[27322]_  & \new_[27319]_ ;
  assign \new_[27324]_  = \new_[27323]_  & \new_[27316]_ ;
  assign \new_[27328]_  = A201 & ~A200;
  assign \new_[27329]_  = A199 & \new_[27328]_ ;
  assign \new_[27332]_  = ~A232 & A202;
  assign \new_[27335]_  = ~A234 & A233;
  assign \new_[27336]_  = \new_[27335]_  & \new_[27332]_ ;
  assign \new_[27337]_  = \new_[27336]_  & \new_[27329]_ ;
  assign \new_[27340]_  = A236 & ~A235;
  assign \new_[27343]_  = ~A269 & ~A267;
  assign \new_[27344]_  = \new_[27343]_  & \new_[27340]_ ;
  assign \new_[27347]_  = A299 & ~A298;
  assign \new_[27350]_  = A301 & A300;
  assign \new_[27351]_  = \new_[27350]_  & \new_[27347]_ ;
  assign \new_[27352]_  = \new_[27351]_  & \new_[27344]_ ;
  assign \new_[27356]_  = A201 & ~A200;
  assign \new_[27357]_  = A199 & \new_[27356]_ ;
  assign \new_[27360]_  = ~A232 & A202;
  assign \new_[27363]_  = ~A234 & A233;
  assign \new_[27364]_  = \new_[27363]_  & \new_[27360]_ ;
  assign \new_[27365]_  = \new_[27364]_  & \new_[27357]_ ;
  assign \new_[27368]_  = A236 & ~A235;
  assign \new_[27371]_  = ~A269 & ~A267;
  assign \new_[27372]_  = \new_[27371]_  & \new_[27368]_ ;
  assign \new_[27375]_  = A299 & ~A298;
  assign \new_[27378]_  = ~A302 & A300;
  assign \new_[27379]_  = \new_[27378]_  & \new_[27375]_ ;
  assign \new_[27380]_  = \new_[27379]_  & \new_[27372]_ ;
  assign \new_[27384]_  = A201 & ~A200;
  assign \new_[27385]_  = A199 & \new_[27384]_ ;
  assign \new_[27388]_  = ~A232 & A202;
  assign \new_[27391]_  = ~A234 & A233;
  assign \new_[27392]_  = \new_[27391]_  & \new_[27388]_ ;
  assign \new_[27393]_  = \new_[27392]_  & \new_[27385]_ ;
  assign \new_[27396]_  = A236 & ~A235;
  assign \new_[27399]_  = A266 & A265;
  assign \new_[27400]_  = \new_[27399]_  & \new_[27396]_ ;
  assign \new_[27403]_  = ~A299 & A298;
  assign \new_[27406]_  = A301 & A300;
  assign \new_[27407]_  = \new_[27406]_  & \new_[27403]_ ;
  assign \new_[27408]_  = \new_[27407]_  & \new_[27400]_ ;
  assign \new_[27412]_  = A201 & ~A200;
  assign \new_[27413]_  = A199 & \new_[27412]_ ;
  assign \new_[27416]_  = ~A232 & A202;
  assign \new_[27419]_  = ~A234 & A233;
  assign \new_[27420]_  = \new_[27419]_  & \new_[27416]_ ;
  assign \new_[27421]_  = \new_[27420]_  & \new_[27413]_ ;
  assign \new_[27424]_  = A236 & ~A235;
  assign \new_[27427]_  = A266 & A265;
  assign \new_[27428]_  = \new_[27427]_  & \new_[27424]_ ;
  assign \new_[27431]_  = ~A299 & A298;
  assign \new_[27434]_  = ~A302 & A300;
  assign \new_[27435]_  = \new_[27434]_  & \new_[27431]_ ;
  assign \new_[27436]_  = \new_[27435]_  & \new_[27428]_ ;
  assign \new_[27440]_  = A201 & ~A200;
  assign \new_[27441]_  = A199 & \new_[27440]_ ;
  assign \new_[27444]_  = ~A232 & A202;
  assign \new_[27447]_  = ~A234 & A233;
  assign \new_[27448]_  = \new_[27447]_  & \new_[27444]_ ;
  assign \new_[27449]_  = \new_[27448]_  & \new_[27441]_ ;
  assign \new_[27452]_  = A236 & ~A235;
  assign \new_[27455]_  = A266 & A265;
  assign \new_[27456]_  = \new_[27455]_  & \new_[27452]_ ;
  assign \new_[27459]_  = A299 & ~A298;
  assign \new_[27462]_  = A301 & A300;
  assign \new_[27463]_  = \new_[27462]_  & \new_[27459]_ ;
  assign \new_[27464]_  = \new_[27463]_  & \new_[27456]_ ;
  assign \new_[27468]_  = A201 & ~A200;
  assign \new_[27469]_  = A199 & \new_[27468]_ ;
  assign \new_[27472]_  = ~A232 & A202;
  assign \new_[27475]_  = ~A234 & A233;
  assign \new_[27476]_  = \new_[27475]_  & \new_[27472]_ ;
  assign \new_[27477]_  = \new_[27476]_  & \new_[27469]_ ;
  assign \new_[27480]_  = A236 & ~A235;
  assign \new_[27483]_  = A266 & A265;
  assign \new_[27484]_  = \new_[27483]_  & \new_[27480]_ ;
  assign \new_[27487]_  = A299 & ~A298;
  assign \new_[27490]_  = ~A302 & A300;
  assign \new_[27491]_  = \new_[27490]_  & \new_[27487]_ ;
  assign \new_[27492]_  = \new_[27491]_  & \new_[27484]_ ;
  assign \new_[27496]_  = A201 & ~A200;
  assign \new_[27497]_  = A199 & \new_[27496]_ ;
  assign \new_[27500]_  = ~A232 & A202;
  assign \new_[27503]_  = ~A234 & A233;
  assign \new_[27504]_  = \new_[27503]_  & \new_[27500]_ ;
  assign \new_[27505]_  = \new_[27504]_  & \new_[27497]_ ;
  assign \new_[27508]_  = A236 & ~A235;
  assign \new_[27511]_  = ~A266 & ~A265;
  assign \new_[27512]_  = \new_[27511]_  & \new_[27508]_ ;
  assign \new_[27515]_  = ~A299 & A298;
  assign \new_[27518]_  = A301 & A300;
  assign \new_[27519]_  = \new_[27518]_  & \new_[27515]_ ;
  assign \new_[27520]_  = \new_[27519]_  & \new_[27512]_ ;
  assign \new_[27524]_  = A201 & ~A200;
  assign \new_[27525]_  = A199 & \new_[27524]_ ;
  assign \new_[27528]_  = ~A232 & A202;
  assign \new_[27531]_  = ~A234 & A233;
  assign \new_[27532]_  = \new_[27531]_  & \new_[27528]_ ;
  assign \new_[27533]_  = \new_[27532]_  & \new_[27525]_ ;
  assign \new_[27536]_  = A236 & ~A235;
  assign \new_[27539]_  = ~A266 & ~A265;
  assign \new_[27540]_  = \new_[27539]_  & \new_[27536]_ ;
  assign \new_[27543]_  = ~A299 & A298;
  assign \new_[27546]_  = ~A302 & A300;
  assign \new_[27547]_  = \new_[27546]_  & \new_[27543]_ ;
  assign \new_[27548]_  = \new_[27547]_  & \new_[27540]_ ;
  assign \new_[27552]_  = A201 & ~A200;
  assign \new_[27553]_  = A199 & \new_[27552]_ ;
  assign \new_[27556]_  = ~A232 & A202;
  assign \new_[27559]_  = ~A234 & A233;
  assign \new_[27560]_  = \new_[27559]_  & \new_[27556]_ ;
  assign \new_[27561]_  = \new_[27560]_  & \new_[27553]_ ;
  assign \new_[27564]_  = A236 & ~A235;
  assign \new_[27567]_  = ~A266 & ~A265;
  assign \new_[27568]_  = \new_[27567]_  & \new_[27564]_ ;
  assign \new_[27571]_  = A299 & ~A298;
  assign \new_[27574]_  = A301 & A300;
  assign \new_[27575]_  = \new_[27574]_  & \new_[27571]_ ;
  assign \new_[27576]_  = \new_[27575]_  & \new_[27568]_ ;
  assign \new_[27580]_  = A201 & ~A200;
  assign \new_[27581]_  = A199 & \new_[27580]_ ;
  assign \new_[27584]_  = ~A232 & A202;
  assign \new_[27587]_  = ~A234 & A233;
  assign \new_[27588]_  = \new_[27587]_  & \new_[27584]_ ;
  assign \new_[27589]_  = \new_[27588]_  & \new_[27581]_ ;
  assign \new_[27592]_  = A236 & ~A235;
  assign \new_[27595]_  = ~A266 & ~A265;
  assign \new_[27596]_  = \new_[27595]_  & \new_[27592]_ ;
  assign \new_[27599]_  = A299 & ~A298;
  assign \new_[27602]_  = ~A302 & A300;
  assign \new_[27603]_  = \new_[27602]_  & \new_[27599]_ ;
  assign \new_[27604]_  = \new_[27603]_  & \new_[27596]_ ;
  assign \new_[27608]_  = A201 & ~A200;
  assign \new_[27609]_  = A199 & \new_[27608]_ ;
  assign \new_[27612]_  = A232 & A202;
  assign \new_[27615]_  = A234 & ~A233;
  assign \new_[27616]_  = \new_[27615]_  & \new_[27612]_ ;
  assign \new_[27617]_  = \new_[27616]_  & \new_[27609]_ ;
  assign \new_[27620]_  = A267 & A235;
  assign \new_[27623]_  = A269 & ~A268;
  assign \new_[27624]_  = \new_[27623]_  & \new_[27620]_ ;
  assign \new_[27627]_  = ~A299 & A298;
  assign \new_[27630]_  = A301 & A300;
  assign \new_[27631]_  = \new_[27630]_  & \new_[27627]_ ;
  assign \new_[27632]_  = \new_[27631]_  & \new_[27624]_ ;
  assign \new_[27636]_  = A201 & ~A200;
  assign \new_[27637]_  = A199 & \new_[27636]_ ;
  assign \new_[27640]_  = A232 & A202;
  assign \new_[27643]_  = A234 & ~A233;
  assign \new_[27644]_  = \new_[27643]_  & \new_[27640]_ ;
  assign \new_[27645]_  = \new_[27644]_  & \new_[27637]_ ;
  assign \new_[27648]_  = A267 & A235;
  assign \new_[27651]_  = A269 & ~A268;
  assign \new_[27652]_  = \new_[27651]_  & \new_[27648]_ ;
  assign \new_[27655]_  = ~A299 & A298;
  assign \new_[27658]_  = ~A302 & A300;
  assign \new_[27659]_  = \new_[27658]_  & \new_[27655]_ ;
  assign \new_[27660]_  = \new_[27659]_  & \new_[27652]_ ;
  assign \new_[27664]_  = A201 & ~A200;
  assign \new_[27665]_  = A199 & \new_[27664]_ ;
  assign \new_[27668]_  = A232 & A202;
  assign \new_[27671]_  = A234 & ~A233;
  assign \new_[27672]_  = \new_[27671]_  & \new_[27668]_ ;
  assign \new_[27673]_  = \new_[27672]_  & \new_[27665]_ ;
  assign \new_[27676]_  = A267 & A235;
  assign \new_[27679]_  = A269 & ~A268;
  assign \new_[27680]_  = \new_[27679]_  & \new_[27676]_ ;
  assign \new_[27683]_  = A299 & ~A298;
  assign \new_[27686]_  = A301 & A300;
  assign \new_[27687]_  = \new_[27686]_  & \new_[27683]_ ;
  assign \new_[27688]_  = \new_[27687]_  & \new_[27680]_ ;
  assign \new_[27692]_  = A201 & ~A200;
  assign \new_[27693]_  = A199 & \new_[27692]_ ;
  assign \new_[27696]_  = A232 & A202;
  assign \new_[27699]_  = A234 & ~A233;
  assign \new_[27700]_  = \new_[27699]_  & \new_[27696]_ ;
  assign \new_[27701]_  = \new_[27700]_  & \new_[27693]_ ;
  assign \new_[27704]_  = A267 & A235;
  assign \new_[27707]_  = A269 & ~A268;
  assign \new_[27708]_  = \new_[27707]_  & \new_[27704]_ ;
  assign \new_[27711]_  = A299 & ~A298;
  assign \new_[27714]_  = ~A302 & A300;
  assign \new_[27715]_  = \new_[27714]_  & \new_[27711]_ ;
  assign \new_[27716]_  = \new_[27715]_  & \new_[27708]_ ;
  assign \new_[27720]_  = A201 & ~A200;
  assign \new_[27721]_  = A199 & \new_[27720]_ ;
  assign \new_[27724]_  = A232 & A202;
  assign \new_[27727]_  = A234 & ~A233;
  assign \new_[27728]_  = \new_[27727]_  & \new_[27724]_ ;
  assign \new_[27729]_  = \new_[27728]_  & \new_[27721]_ ;
  assign \new_[27732]_  = ~A267 & A235;
  assign \new_[27735]_  = A298 & A268;
  assign \new_[27736]_  = \new_[27735]_  & \new_[27732]_ ;
  assign \new_[27739]_  = ~A300 & ~A299;
  assign \new_[27742]_  = A302 & ~A301;
  assign \new_[27743]_  = \new_[27742]_  & \new_[27739]_ ;
  assign \new_[27744]_  = \new_[27743]_  & \new_[27736]_ ;
  assign \new_[27748]_  = A201 & ~A200;
  assign \new_[27749]_  = A199 & \new_[27748]_ ;
  assign \new_[27752]_  = A232 & A202;
  assign \new_[27755]_  = A234 & ~A233;
  assign \new_[27756]_  = \new_[27755]_  & \new_[27752]_ ;
  assign \new_[27757]_  = \new_[27756]_  & \new_[27749]_ ;
  assign \new_[27760]_  = ~A267 & A235;
  assign \new_[27763]_  = ~A298 & A268;
  assign \new_[27764]_  = \new_[27763]_  & \new_[27760]_ ;
  assign \new_[27767]_  = ~A300 & A299;
  assign \new_[27770]_  = A302 & ~A301;
  assign \new_[27771]_  = \new_[27770]_  & \new_[27767]_ ;
  assign \new_[27772]_  = \new_[27771]_  & \new_[27764]_ ;
  assign \new_[27776]_  = A201 & ~A200;
  assign \new_[27777]_  = A199 & \new_[27776]_ ;
  assign \new_[27780]_  = A232 & A202;
  assign \new_[27783]_  = A234 & ~A233;
  assign \new_[27784]_  = \new_[27783]_  & \new_[27780]_ ;
  assign \new_[27785]_  = \new_[27784]_  & \new_[27777]_ ;
  assign \new_[27788]_  = ~A267 & A235;
  assign \new_[27791]_  = A298 & ~A269;
  assign \new_[27792]_  = \new_[27791]_  & \new_[27788]_ ;
  assign \new_[27795]_  = ~A300 & ~A299;
  assign \new_[27798]_  = A302 & ~A301;
  assign \new_[27799]_  = \new_[27798]_  & \new_[27795]_ ;
  assign \new_[27800]_  = \new_[27799]_  & \new_[27792]_ ;
  assign \new_[27804]_  = A201 & ~A200;
  assign \new_[27805]_  = A199 & \new_[27804]_ ;
  assign \new_[27808]_  = A232 & A202;
  assign \new_[27811]_  = A234 & ~A233;
  assign \new_[27812]_  = \new_[27811]_  & \new_[27808]_ ;
  assign \new_[27813]_  = \new_[27812]_  & \new_[27805]_ ;
  assign \new_[27816]_  = ~A267 & A235;
  assign \new_[27819]_  = ~A298 & ~A269;
  assign \new_[27820]_  = \new_[27819]_  & \new_[27816]_ ;
  assign \new_[27823]_  = ~A300 & A299;
  assign \new_[27826]_  = A302 & ~A301;
  assign \new_[27827]_  = \new_[27826]_  & \new_[27823]_ ;
  assign \new_[27828]_  = \new_[27827]_  & \new_[27820]_ ;
  assign \new_[27832]_  = A201 & ~A200;
  assign \new_[27833]_  = A199 & \new_[27832]_ ;
  assign \new_[27836]_  = A232 & A202;
  assign \new_[27839]_  = A234 & ~A233;
  assign \new_[27840]_  = \new_[27839]_  & \new_[27836]_ ;
  assign \new_[27841]_  = \new_[27840]_  & \new_[27833]_ ;
  assign \new_[27844]_  = A265 & A235;
  assign \new_[27847]_  = A298 & A266;
  assign \new_[27848]_  = \new_[27847]_  & \new_[27844]_ ;
  assign \new_[27851]_  = ~A300 & ~A299;
  assign \new_[27854]_  = A302 & ~A301;
  assign \new_[27855]_  = \new_[27854]_  & \new_[27851]_ ;
  assign \new_[27856]_  = \new_[27855]_  & \new_[27848]_ ;
  assign \new_[27860]_  = A201 & ~A200;
  assign \new_[27861]_  = A199 & \new_[27860]_ ;
  assign \new_[27864]_  = A232 & A202;
  assign \new_[27867]_  = A234 & ~A233;
  assign \new_[27868]_  = \new_[27867]_  & \new_[27864]_ ;
  assign \new_[27869]_  = \new_[27868]_  & \new_[27861]_ ;
  assign \new_[27872]_  = A265 & A235;
  assign \new_[27875]_  = ~A298 & A266;
  assign \new_[27876]_  = \new_[27875]_  & \new_[27872]_ ;
  assign \new_[27879]_  = ~A300 & A299;
  assign \new_[27882]_  = A302 & ~A301;
  assign \new_[27883]_  = \new_[27882]_  & \new_[27879]_ ;
  assign \new_[27884]_  = \new_[27883]_  & \new_[27876]_ ;
  assign \new_[27888]_  = A201 & ~A200;
  assign \new_[27889]_  = A199 & \new_[27888]_ ;
  assign \new_[27892]_  = A232 & A202;
  assign \new_[27895]_  = A234 & ~A233;
  assign \new_[27896]_  = \new_[27895]_  & \new_[27892]_ ;
  assign \new_[27897]_  = \new_[27896]_  & \new_[27889]_ ;
  assign \new_[27900]_  = ~A265 & A235;
  assign \new_[27903]_  = A298 & ~A266;
  assign \new_[27904]_  = \new_[27903]_  & \new_[27900]_ ;
  assign \new_[27907]_  = ~A300 & ~A299;
  assign \new_[27910]_  = A302 & ~A301;
  assign \new_[27911]_  = \new_[27910]_  & \new_[27907]_ ;
  assign \new_[27912]_  = \new_[27911]_  & \new_[27904]_ ;
  assign \new_[27916]_  = A201 & ~A200;
  assign \new_[27917]_  = A199 & \new_[27916]_ ;
  assign \new_[27920]_  = A232 & A202;
  assign \new_[27923]_  = A234 & ~A233;
  assign \new_[27924]_  = \new_[27923]_  & \new_[27920]_ ;
  assign \new_[27925]_  = \new_[27924]_  & \new_[27917]_ ;
  assign \new_[27928]_  = ~A265 & A235;
  assign \new_[27931]_  = ~A298 & ~A266;
  assign \new_[27932]_  = \new_[27931]_  & \new_[27928]_ ;
  assign \new_[27935]_  = ~A300 & A299;
  assign \new_[27938]_  = A302 & ~A301;
  assign \new_[27939]_  = \new_[27938]_  & \new_[27935]_ ;
  assign \new_[27940]_  = \new_[27939]_  & \new_[27932]_ ;
  assign \new_[27944]_  = A201 & ~A200;
  assign \new_[27945]_  = A199 & \new_[27944]_ ;
  assign \new_[27948]_  = A232 & A202;
  assign \new_[27951]_  = A234 & ~A233;
  assign \new_[27952]_  = \new_[27951]_  & \new_[27948]_ ;
  assign \new_[27953]_  = \new_[27952]_  & \new_[27945]_ ;
  assign \new_[27956]_  = A267 & ~A236;
  assign \new_[27959]_  = A269 & ~A268;
  assign \new_[27960]_  = \new_[27959]_  & \new_[27956]_ ;
  assign \new_[27963]_  = ~A299 & A298;
  assign \new_[27966]_  = A301 & A300;
  assign \new_[27967]_  = \new_[27966]_  & \new_[27963]_ ;
  assign \new_[27968]_  = \new_[27967]_  & \new_[27960]_ ;
  assign \new_[27972]_  = A201 & ~A200;
  assign \new_[27973]_  = A199 & \new_[27972]_ ;
  assign \new_[27976]_  = A232 & A202;
  assign \new_[27979]_  = A234 & ~A233;
  assign \new_[27980]_  = \new_[27979]_  & \new_[27976]_ ;
  assign \new_[27981]_  = \new_[27980]_  & \new_[27973]_ ;
  assign \new_[27984]_  = A267 & ~A236;
  assign \new_[27987]_  = A269 & ~A268;
  assign \new_[27988]_  = \new_[27987]_  & \new_[27984]_ ;
  assign \new_[27991]_  = ~A299 & A298;
  assign \new_[27994]_  = ~A302 & A300;
  assign \new_[27995]_  = \new_[27994]_  & \new_[27991]_ ;
  assign \new_[27996]_  = \new_[27995]_  & \new_[27988]_ ;
  assign \new_[28000]_  = A201 & ~A200;
  assign \new_[28001]_  = A199 & \new_[28000]_ ;
  assign \new_[28004]_  = A232 & A202;
  assign \new_[28007]_  = A234 & ~A233;
  assign \new_[28008]_  = \new_[28007]_  & \new_[28004]_ ;
  assign \new_[28009]_  = \new_[28008]_  & \new_[28001]_ ;
  assign \new_[28012]_  = A267 & ~A236;
  assign \new_[28015]_  = A269 & ~A268;
  assign \new_[28016]_  = \new_[28015]_  & \new_[28012]_ ;
  assign \new_[28019]_  = A299 & ~A298;
  assign \new_[28022]_  = A301 & A300;
  assign \new_[28023]_  = \new_[28022]_  & \new_[28019]_ ;
  assign \new_[28024]_  = \new_[28023]_  & \new_[28016]_ ;
  assign \new_[28028]_  = A201 & ~A200;
  assign \new_[28029]_  = A199 & \new_[28028]_ ;
  assign \new_[28032]_  = A232 & A202;
  assign \new_[28035]_  = A234 & ~A233;
  assign \new_[28036]_  = \new_[28035]_  & \new_[28032]_ ;
  assign \new_[28037]_  = \new_[28036]_  & \new_[28029]_ ;
  assign \new_[28040]_  = A267 & ~A236;
  assign \new_[28043]_  = A269 & ~A268;
  assign \new_[28044]_  = \new_[28043]_  & \new_[28040]_ ;
  assign \new_[28047]_  = A299 & ~A298;
  assign \new_[28050]_  = ~A302 & A300;
  assign \new_[28051]_  = \new_[28050]_  & \new_[28047]_ ;
  assign \new_[28052]_  = \new_[28051]_  & \new_[28044]_ ;
  assign \new_[28056]_  = A201 & ~A200;
  assign \new_[28057]_  = A199 & \new_[28056]_ ;
  assign \new_[28060]_  = A232 & A202;
  assign \new_[28063]_  = A234 & ~A233;
  assign \new_[28064]_  = \new_[28063]_  & \new_[28060]_ ;
  assign \new_[28065]_  = \new_[28064]_  & \new_[28057]_ ;
  assign \new_[28068]_  = ~A267 & ~A236;
  assign \new_[28071]_  = A298 & A268;
  assign \new_[28072]_  = \new_[28071]_  & \new_[28068]_ ;
  assign \new_[28075]_  = ~A300 & ~A299;
  assign \new_[28078]_  = A302 & ~A301;
  assign \new_[28079]_  = \new_[28078]_  & \new_[28075]_ ;
  assign \new_[28080]_  = \new_[28079]_  & \new_[28072]_ ;
  assign \new_[28084]_  = A201 & ~A200;
  assign \new_[28085]_  = A199 & \new_[28084]_ ;
  assign \new_[28088]_  = A232 & A202;
  assign \new_[28091]_  = A234 & ~A233;
  assign \new_[28092]_  = \new_[28091]_  & \new_[28088]_ ;
  assign \new_[28093]_  = \new_[28092]_  & \new_[28085]_ ;
  assign \new_[28096]_  = ~A267 & ~A236;
  assign \new_[28099]_  = ~A298 & A268;
  assign \new_[28100]_  = \new_[28099]_  & \new_[28096]_ ;
  assign \new_[28103]_  = ~A300 & A299;
  assign \new_[28106]_  = A302 & ~A301;
  assign \new_[28107]_  = \new_[28106]_  & \new_[28103]_ ;
  assign \new_[28108]_  = \new_[28107]_  & \new_[28100]_ ;
  assign \new_[28112]_  = A201 & ~A200;
  assign \new_[28113]_  = A199 & \new_[28112]_ ;
  assign \new_[28116]_  = A232 & A202;
  assign \new_[28119]_  = A234 & ~A233;
  assign \new_[28120]_  = \new_[28119]_  & \new_[28116]_ ;
  assign \new_[28121]_  = \new_[28120]_  & \new_[28113]_ ;
  assign \new_[28124]_  = ~A267 & ~A236;
  assign \new_[28127]_  = A298 & ~A269;
  assign \new_[28128]_  = \new_[28127]_  & \new_[28124]_ ;
  assign \new_[28131]_  = ~A300 & ~A299;
  assign \new_[28134]_  = A302 & ~A301;
  assign \new_[28135]_  = \new_[28134]_  & \new_[28131]_ ;
  assign \new_[28136]_  = \new_[28135]_  & \new_[28128]_ ;
  assign \new_[28140]_  = A201 & ~A200;
  assign \new_[28141]_  = A199 & \new_[28140]_ ;
  assign \new_[28144]_  = A232 & A202;
  assign \new_[28147]_  = A234 & ~A233;
  assign \new_[28148]_  = \new_[28147]_  & \new_[28144]_ ;
  assign \new_[28149]_  = \new_[28148]_  & \new_[28141]_ ;
  assign \new_[28152]_  = ~A267 & ~A236;
  assign \new_[28155]_  = ~A298 & ~A269;
  assign \new_[28156]_  = \new_[28155]_  & \new_[28152]_ ;
  assign \new_[28159]_  = ~A300 & A299;
  assign \new_[28162]_  = A302 & ~A301;
  assign \new_[28163]_  = \new_[28162]_  & \new_[28159]_ ;
  assign \new_[28164]_  = \new_[28163]_  & \new_[28156]_ ;
  assign \new_[28168]_  = A201 & ~A200;
  assign \new_[28169]_  = A199 & \new_[28168]_ ;
  assign \new_[28172]_  = A232 & A202;
  assign \new_[28175]_  = A234 & ~A233;
  assign \new_[28176]_  = \new_[28175]_  & \new_[28172]_ ;
  assign \new_[28177]_  = \new_[28176]_  & \new_[28169]_ ;
  assign \new_[28180]_  = A265 & ~A236;
  assign \new_[28183]_  = A298 & A266;
  assign \new_[28184]_  = \new_[28183]_  & \new_[28180]_ ;
  assign \new_[28187]_  = ~A300 & ~A299;
  assign \new_[28190]_  = A302 & ~A301;
  assign \new_[28191]_  = \new_[28190]_  & \new_[28187]_ ;
  assign \new_[28192]_  = \new_[28191]_  & \new_[28184]_ ;
  assign \new_[28196]_  = A201 & ~A200;
  assign \new_[28197]_  = A199 & \new_[28196]_ ;
  assign \new_[28200]_  = A232 & A202;
  assign \new_[28203]_  = A234 & ~A233;
  assign \new_[28204]_  = \new_[28203]_  & \new_[28200]_ ;
  assign \new_[28205]_  = \new_[28204]_  & \new_[28197]_ ;
  assign \new_[28208]_  = A265 & ~A236;
  assign \new_[28211]_  = ~A298 & A266;
  assign \new_[28212]_  = \new_[28211]_  & \new_[28208]_ ;
  assign \new_[28215]_  = ~A300 & A299;
  assign \new_[28218]_  = A302 & ~A301;
  assign \new_[28219]_  = \new_[28218]_  & \new_[28215]_ ;
  assign \new_[28220]_  = \new_[28219]_  & \new_[28212]_ ;
  assign \new_[28224]_  = A201 & ~A200;
  assign \new_[28225]_  = A199 & \new_[28224]_ ;
  assign \new_[28228]_  = A232 & A202;
  assign \new_[28231]_  = A234 & ~A233;
  assign \new_[28232]_  = \new_[28231]_  & \new_[28228]_ ;
  assign \new_[28233]_  = \new_[28232]_  & \new_[28225]_ ;
  assign \new_[28236]_  = ~A265 & ~A236;
  assign \new_[28239]_  = A298 & ~A266;
  assign \new_[28240]_  = \new_[28239]_  & \new_[28236]_ ;
  assign \new_[28243]_  = ~A300 & ~A299;
  assign \new_[28246]_  = A302 & ~A301;
  assign \new_[28247]_  = \new_[28246]_  & \new_[28243]_ ;
  assign \new_[28248]_  = \new_[28247]_  & \new_[28240]_ ;
  assign \new_[28252]_  = A201 & ~A200;
  assign \new_[28253]_  = A199 & \new_[28252]_ ;
  assign \new_[28256]_  = A232 & A202;
  assign \new_[28259]_  = A234 & ~A233;
  assign \new_[28260]_  = \new_[28259]_  & \new_[28256]_ ;
  assign \new_[28261]_  = \new_[28260]_  & \new_[28253]_ ;
  assign \new_[28264]_  = ~A265 & ~A236;
  assign \new_[28267]_  = ~A298 & ~A266;
  assign \new_[28268]_  = \new_[28267]_  & \new_[28264]_ ;
  assign \new_[28271]_  = ~A300 & A299;
  assign \new_[28274]_  = A302 & ~A301;
  assign \new_[28275]_  = \new_[28274]_  & \new_[28271]_ ;
  assign \new_[28276]_  = \new_[28275]_  & \new_[28268]_ ;
  assign \new_[28280]_  = A201 & ~A200;
  assign \new_[28281]_  = A199 & \new_[28280]_ ;
  assign \new_[28284]_  = A232 & A202;
  assign \new_[28287]_  = ~A234 & ~A233;
  assign \new_[28288]_  = \new_[28287]_  & \new_[28284]_ ;
  assign \new_[28289]_  = \new_[28288]_  & \new_[28281]_ ;
  assign \new_[28292]_  = A236 & ~A235;
  assign \new_[28295]_  = A268 & ~A267;
  assign \new_[28296]_  = \new_[28295]_  & \new_[28292]_ ;
  assign \new_[28299]_  = ~A299 & A298;
  assign \new_[28302]_  = A301 & A300;
  assign \new_[28303]_  = \new_[28302]_  & \new_[28299]_ ;
  assign \new_[28304]_  = \new_[28303]_  & \new_[28296]_ ;
  assign \new_[28308]_  = A201 & ~A200;
  assign \new_[28309]_  = A199 & \new_[28308]_ ;
  assign \new_[28312]_  = A232 & A202;
  assign \new_[28315]_  = ~A234 & ~A233;
  assign \new_[28316]_  = \new_[28315]_  & \new_[28312]_ ;
  assign \new_[28317]_  = \new_[28316]_  & \new_[28309]_ ;
  assign \new_[28320]_  = A236 & ~A235;
  assign \new_[28323]_  = A268 & ~A267;
  assign \new_[28324]_  = \new_[28323]_  & \new_[28320]_ ;
  assign \new_[28327]_  = ~A299 & A298;
  assign \new_[28330]_  = ~A302 & A300;
  assign \new_[28331]_  = \new_[28330]_  & \new_[28327]_ ;
  assign \new_[28332]_  = \new_[28331]_  & \new_[28324]_ ;
  assign \new_[28336]_  = A201 & ~A200;
  assign \new_[28337]_  = A199 & \new_[28336]_ ;
  assign \new_[28340]_  = A232 & A202;
  assign \new_[28343]_  = ~A234 & ~A233;
  assign \new_[28344]_  = \new_[28343]_  & \new_[28340]_ ;
  assign \new_[28345]_  = \new_[28344]_  & \new_[28337]_ ;
  assign \new_[28348]_  = A236 & ~A235;
  assign \new_[28351]_  = A268 & ~A267;
  assign \new_[28352]_  = \new_[28351]_  & \new_[28348]_ ;
  assign \new_[28355]_  = A299 & ~A298;
  assign \new_[28358]_  = A301 & A300;
  assign \new_[28359]_  = \new_[28358]_  & \new_[28355]_ ;
  assign \new_[28360]_  = \new_[28359]_  & \new_[28352]_ ;
  assign \new_[28364]_  = A201 & ~A200;
  assign \new_[28365]_  = A199 & \new_[28364]_ ;
  assign \new_[28368]_  = A232 & A202;
  assign \new_[28371]_  = ~A234 & ~A233;
  assign \new_[28372]_  = \new_[28371]_  & \new_[28368]_ ;
  assign \new_[28373]_  = \new_[28372]_  & \new_[28365]_ ;
  assign \new_[28376]_  = A236 & ~A235;
  assign \new_[28379]_  = A268 & ~A267;
  assign \new_[28380]_  = \new_[28379]_  & \new_[28376]_ ;
  assign \new_[28383]_  = A299 & ~A298;
  assign \new_[28386]_  = ~A302 & A300;
  assign \new_[28387]_  = \new_[28386]_  & \new_[28383]_ ;
  assign \new_[28388]_  = \new_[28387]_  & \new_[28380]_ ;
  assign \new_[28392]_  = A201 & ~A200;
  assign \new_[28393]_  = A199 & \new_[28392]_ ;
  assign \new_[28396]_  = A232 & A202;
  assign \new_[28399]_  = ~A234 & ~A233;
  assign \new_[28400]_  = \new_[28399]_  & \new_[28396]_ ;
  assign \new_[28401]_  = \new_[28400]_  & \new_[28393]_ ;
  assign \new_[28404]_  = A236 & ~A235;
  assign \new_[28407]_  = ~A269 & ~A267;
  assign \new_[28408]_  = \new_[28407]_  & \new_[28404]_ ;
  assign \new_[28411]_  = ~A299 & A298;
  assign \new_[28414]_  = A301 & A300;
  assign \new_[28415]_  = \new_[28414]_  & \new_[28411]_ ;
  assign \new_[28416]_  = \new_[28415]_  & \new_[28408]_ ;
  assign \new_[28420]_  = A201 & ~A200;
  assign \new_[28421]_  = A199 & \new_[28420]_ ;
  assign \new_[28424]_  = A232 & A202;
  assign \new_[28427]_  = ~A234 & ~A233;
  assign \new_[28428]_  = \new_[28427]_  & \new_[28424]_ ;
  assign \new_[28429]_  = \new_[28428]_  & \new_[28421]_ ;
  assign \new_[28432]_  = A236 & ~A235;
  assign \new_[28435]_  = ~A269 & ~A267;
  assign \new_[28436]_  = \new_[28435]_  & \new_[28432]_ ;
  assign \new_[28439]_  = ~A299 & A298;
  assign \new_[28442]_  = ~A302 & A300;
  assign \new_[28443]_  = \new_[28442]_  & \new_[28439]_ ;
  assign \new_[28444]_  = \new_[28443]_  & \new_[28436]_ ;
  assign \new_[28448]_  = A201 & ~A200;
  assign \new_[28449]_  = A199 & \new_[28448]_ ;
  assign \new_[28452]_  = A232 & A202;
  assign \new_[28455]_  = ~A234 & ~A233;
  assign \new_[28456]_  = \new_[28455]_  & \new_[28452]_ ;
  assign \new_[28457]_  = \new_[28456]_  & \new_[28449]_ ;
  assign \new_[28460]_  = A236 & ~A235;
  assign \new_[28463]_  = ~A269 & ~A267;
  assign \new_[28464]_  = \new_[28463]_  & \new_[28460]_ ;
  assign \new_[28467]_  = A299 & ~A298;
  assign \new_[28470]_  = A301 & A300;
  assign \new_[28471]_  = \new_[28470]_  & \new_[28467]_ ;
  assign \new_[28472]_  = \new_[28471]_  & \new_[28464]_ ;
  assign \new_[28476]_  = A201 & ~A200;
  assign \new_[28477]_  = A199 & \new_[28476]_ ;
  assign \new_[28480]_  = A232 & A202;
  assign \new_[28483]_  = ~A234 & ~A233;
  assign \new_[28484]_  = \new_[28483]_  & \new_[28480]_ ;
  assign \new_[28485]_  = \new_[28484]_  & \new_[28477]_ ;
  assign \new_[28488]_  = A236 & ~A235;
  assign \new_[28491]_  = ~A269 & ~A267;
  assign \new_[28492]_  = \new_[28491]_  & \new_[28488]_ ;
  assign \new_[28495]_  = A299 & ~A298;
  assign \new_[28498]_  = ~A302 & A300;
  assign \new_[28499]_  = \new_[28498]_  & \new_[28495]_ ;
  assign \new_[28500]_  = \new_[28499]_  & \new_[28492]_ ;
  assign \new_[28504]_  = A201 & ~A200;
  assign \new_[28505]_  = A199 & \new_[28504]_ ;
  assign \new_[28508]_  = A232 & A202;
  assign \new_[28511]_  = ~A234 & ~A233;
  assign \new_[28512]_  = \new_[28511]_  & \new_[28508]_ ;
  assign \new_[28513]_  = \new_[28512]_  & \new_[28505]_ ;
  assign \new_[28516]_  = A236 & ~A235;
  assign \new_[28519]_  = A266 & A265;
  assign \new_[28520]_  = \new_[28519]_  & \new_[28516]_ ;
  assign \new_[28523]_  = ~A299 & A298;
  assign \new_[28526]_  = A301 & A300;
  assign \new_[28527]_  = \new_[28526]_  & \new_[28523]_ ;
  assign \new_[28528]_  = \new_[28527]_  & \new_[28520]_ ;
  assign \new_[28532]_  = A201 & ~A200;
  assign \new_[28533]_  = A199 & \new_[28532]_ ;
  assign \new_[28536]_  = A232 & A202;
  assign \new_[28539]_  = ~A234 & ~A233;
  assign \new_[28540]_  = \new_[28539]_  & \new_[28536]_ ;
  assign \new_[28541]_  = \new_[28540]_  & \new_[28533]_ ;
  assign \new_[28544]_  = A236 & ~A235;
  assign \new_[28547]_  = A266 & A265;
  assign \new_[28548]_  = \new_[28547]_  & \new_[28544]_ ;
  assign \new_[28551]_  = ~A299 & A298;
  assign \new_[28554]_  = ~A302 & A300;
  assign \new_[28555]_  = \new_[28554]_  & \new_[28551]_ ;
  assign \new_[28556]_  = \new_[28555]_  & \new_[28548]_ ;
  assign \new_[28560]_  = A201 & ~A200;
  assign \new_[28561]_  = A199 & \new_[28560]_ ;
  assign \new_[28564]_  = A232 & A202;
  assign \new_[28567]_  = ~A234 & ~A233;
  assign \new_[28568]_  = \new_[28567]_  & \new_[28564]_ ;
  assign \new_[28569]_  = \new_[28568]_  & \new_[28561]_ ;
  assign \new_[28572]_  = A236 & ~A235;
  assign \new_[28575]_  = A266 & A265;
  assign \new_[28576]_  = \new_[28575]_  & \new_[28572]_ ;
  assign \new_[28579]_  = A299 & ~A298;
  assign \new_[28582]_  = A301 & A300;
  assign \new_[28583]_  = \new_[28582]_  & \new_[28579]_ ;
  assign \new_[28584]_  = \new_[28583]_  & \new_[28576]_ ;
  assign \new_[28588]_  = A201 & ~A200;
  assign \new_[28589]_  = A199 & \new_[28588]_ ;
  assign \new_[28592]_  = A232 & A202;
  assign \new_[28595]_  = ~A234 & ~A233;
  assign \new_[28596]_  = \new_[28595]_  & \new_[28592]_ ;
  assign \new_[28597]_  = \new_[28596]_  & \new_[28589]_ ;
  assign \new_[28600]_  = A236 & ~A235;
  assign \new_[28603]_  = A266 & A265;
  assign \new_[28604]_  = \new_[28603]_  & \new_[28600]_ ;
  assign \new_[28607]_  = A299 & ~A298;
  assign \new_[28610]_  = ~A302 & A300;
  assign \new_[28611]_  = \new_[28610]_  & \new_[28607]_ ;
  assign \new_[28612]_  = \new_[28611]_  & \new_[28604]_ ;
  assign \new_[28616]_  = A201 & ~A200;
  assign \new_[28617]_  = A199 & \new_[28616]_ ;
  assign \new_[28620]_  = A232 & A202;
  assign \new_[28623]_  = ~A234 & ~A233;
  assign \new_[28624]_  = \new_[28623]_  & \new_[28620]_ ;
  assign \new_[28625]_  = \new_[28624]_  & \new_[28617]_ ;
  assign \new_[28628]_  = A236 & ~A235;
  assign \new_[28631]_  = ~A266 & ~A265;
  assign \new_[28632]_  = \new_[28631]_  & \new_[28628]_ ;
  assign \new_[28635]_  = ~A299 & A298;
  assign \new_[28638]_  = A301 & A300;
  assign \new_[28639]_  = \new_[28638]_  & \new_[28635]_ ;
  assign \new_[28640]_  = \new_[28639]_  & \new_[28632]_ ;
  assign \new_[28644]_  = A201 & ~A200;
  assign \new_[28645]_  = A199 & \new_[28644]_ ;
  assign \new_[28648]_  = A232 & A202;
  assign \new_[28651]_  = ~A234 & ~A233;
  assign \new_[28652]_  = \new_[28651]_  & \new_[28648]_ ;
  assign \new_[28653]_  = \new_[28652]_  & \new_[28645]_ ;
  assign \new_[28656]_  = A236 & ~A235;
  assign \new_[28659]_  = ~A266 & ~A265;
  assign \new_[28660]_  = \new_[28659]_  & \new_[28656]_ ;
  assign \new_[28663]_  = ~A299 & A298;
  assign \new_[28666]_  = ~A302 & A300;
  assign \new_[28667]_  = \new_[28666]_  & \new_[28663]_ ;
  assign \new_[28668]_  = \new_[28667]_  & \new_[28660]_ ;
  assign \new_[28672]_  = A201 & ~A200;
  assign \new_[28673]_  = A199 & \new_[28672]_ ;
  assign \new_[28676]_  = A232 & A202;
  assign \new_[28679]_  = ~A234 & ~A233;
  assign \new_[28680]_  = \new_[28679]_  & \new_[28676]_ ;
  assign \new_[28681]_  = \new_[28680]_  & \new_[28673]_ ;
  assign \new_[28684]_  = A236 & ~A235;
  assign \new_[28687]_  = ~A266 & ~A265;
  assign \new_[28688]_  = \new_[28687]_  & \new_[28684]_ ;
  assign \new_[28691]_  = A299 & ~A298;
  assign \new_[28694]_  = A301 & A300;
  assign \new_[28695]_  = \new_[28694]_  & \new_[28691]_ ;
  assign \new_[28696]_  = \new_[28695]_  & \new_[28688]_ ;
  assign \new_[28700]_  = A201 & ~A200;
  assign \new_[28701]_  = A199 & \new_[28700]_ ;
  assign \new_[28704]_  = A232 & A202;
  assign \new_[28707]_  = ~A234 & ~A233;
  assign \new_[28708]_  = \new_[28707]_  & \new_[28704]_ ;
  assign \new_[28709]_  = \new_[28708]_  & \new_[28701]_ ;
  assign \new_[28712]_  = A236 & ~A235;
  assign \new_[28715]_  = ~A266 & ~A265;
  assign \new_[28716]_  = \new_[28715]_  & \new_[28712]_ ;
  assign \new_[28719]_  = A299 & ~A298;
  assign \new_[28722]_  = ~A302 & A300;
  assign \new_[28723]_  = \new_[28722]_  & \new_[28719]_ ;
  assign \new_[28724]_  = \new_[28723]_  & \new_[28716]_ ;
  assign \new_[28728]_  = A201 & ~A200;
  assign \new_[28729]_  = A199 & \new_[28728]_ ;
  assign \new_[28732]_  = ~A232 & ~A203;
  assign \new_[28735]_  = A234 & A233;
  assign \new_[28736]_  = \new_[28735]_  & \new_[28732]_ ;
  assign \new_[28737]_  = \new_[28736]_  & \new_[28729]_ ;
  assign \new_[28740]_  = A267 & A235;
  assign \new_[28743]_  = A269 & ~A268;
  assign \new_[28744]_  = \new_[28743]_  & \new_[28740]_ ;
  assign \new_[28747]_  = ~A299 & A298;
  assign \new_[28750]_  = A301 & A300;
  assign \new_[28751]_  = \new_[28750]_  & \new_[28747]_ ;
  assign \new_[28752]_  = \new_[28751]_  & \new_[28744]_ ;
  assign \new_[28756]_  = A201 & ~A200;
  assign \new_[28757]_  = A199 & \new_[28756]_ ;
  assign \new_[28760]_  = ~A232 & ~A203;
  assign \new_[28763]_  = A234 & A233;
  assign \new_[28764]_  = \new_[28763]_  & \new_[28760]_ ;
  assign \new_[28765]_  = \new_[28764]_  & \new_[28757]_ ;
  assign \new_[28768]_  = A267 & A235;
  assign \new_[28771]_  = A269 & ~A268;
  assign \new_[28772]_  = \new_[28771]_  & \new_[28768]_ ;
  assign \new_[28775]_  = ~A299 & A298;
  assign \new_[28778]_  = ~A302 & A300;
  assign \new_[28779]_  = \new_[28778]_  & \new_[28775]_ ;
  assign \new_[28780]_  = \new_[28779]_  & \new_[28772]_ ;
  assign \new_[28784]_  = A201 & ~A200;
  assign \new_[28785]_  = A199 & \new_[28784]_ ;
  assign \new_[28788]_  = ~A232 & ~A203;
  assign \new_[28791]_  = A234 & A233;
  assign \new_[28792]_  = \new_[28791]_  & \new_[28788]_ ;
  assign \new_[28793]_  = \new_[28792]_  & \new_[28785]_ ;
  assign \new_[28796]_  = A267 & A235;
  assign \new_[28799]_  = A269 & ~A268;
  assign \new_[28800]_  = \new_[28799]_  & \new_[28796]_ ;
  assign \new_[28803]_  = A299 & ~A298;
  assign \new_[28806]_  = A301 & A300;
  assign \new_[28807]_  = \new_[28806]_  & \new_[28803]_ ;
  assign \new_[28808]_  = \new_[28807]_  & \new_[28800]_ ;
  assign \new_[28812]_  = A201 & ~A200;
  assign \new_[28813]_  = A199 & \new_[28812]_ ;
  assign \new_[28816]_  = ~A232 & ~A203;
  assign \new_[28819]_  = A234 & A233;
  assign \new_[28820]_  = \new_[28819]_  & \new_[28816]_ ;
  assign \new_[28821]_  = \new_[28820]_  & \new_[28813]_ ;
  assign \new_[28824]_  = A267 & A235;
  assign \new_[28827]_  = A269 & ~A268;
  assign \new_[28828]_  = \new_[28827]_  & \new_[28824]_ ;
  assign \new_[28831]_  = A299 & ~A298;
  assign \new_[28834]_  = ~A302 & A300;
  assign \new_[28835]_  = \new_[28834]_  & \new_[28831]_ ;
  assign \new_[28836]_  = \new_[28835]_  & \new_[28828]_ ;
  assign \new_[28840]_  = A201 & ~A200;
  assign \new_[28841]_  = A199 & \new_[28840]_ ;
  assign \new_[28844]_  = ~A232 & ~A203;
  assign \new_[28847]_  = A234 & A233;
  assign \new_[28848]_  = \new_[28847]_  & \new_[28844]_ ;
  assign \new_[28849]_  = \new_[28848]_  & \new_[28841]_ ;
  assign \new_[28852]_  = ~A267 & A235;
  assign \new_[28855]_  = A298 & A268;
  assign \new_[28856]_  = \new_[28855]_  & \new_[28852]_ ;
  assign \new_[28859]_  = ~A300 & ~A299;
  assign \new_[28862]_  = A302 & ~A301;
  assign \new_[28863]_  = \new_[28862]_  & \new_[28859]_ ;
  assign \new_[28864]_  = \new_[28863]_  & \new_[28856]_ ;
  assign \new_[28868]_  = A201 & ~A200;
  assign \new_[28869]_  = A199 & \new_[28868]_ ;
  assign \new_[28872]_  = ~A232 & ~A203;
  assign \new_[28875]_  = A234 & A233;
  assign \new_[28876]_  = \new_[28875]_  & \new_[28872]_ ;
  assign \new_[28877]_  = \new_[28876]_  & \new_[28869]_ ;
  assign \new_[28880]_  = ~A267 & A235;
  assign \new_[28883]_  = ~A298 & A268;
  assign \new_[28884]_  = \new_[28883]_  & \new_[28880]_ ;
  assign \new_[28887]_  = ~A300 & A299;
  assign \new_[28890]_  = A302 & ~A301;
  assign \new_[28891]_  = \new_[28890]_  & \new_[28887]_ ;
  assign \new_[28892]_  = \new_[28891]_  & \new_[28884]_ ;
  assign \new_[28896]_  = A201 & ~A200;
  assign \new_[28897]_  = A199 & \new_[28896]_ ;
  assign \new_[28900]_  = ~A232 & ~A203;
  assign \new_[28903]_  = A234 & A233;
  assign \new_[28904]_  = \new_[28903]_  & \new_[28900]_ ;
  assign \new_[28905]_  = \new_[28904]_  & \new_[28897]_ ;
  assign \new_[28908]_  = ~A267 & A235;
  assign \new_[28911]_  = A298 & ~A269;
  assign \new_[28912]_  = \new_[28911]_  & \new_[28908]_ ;
  assign \new_[28915]_  = ~A300 & ~A299;
  assign \new_[28918]_  = A302 & ~A301;
  assign \new_[28919]_  = \new_[28918]_  & \new_[28915]_ ;
  assign \new_[28920]_  = \new_[28919]_  & \new_[28912]_ ;
  assign \new_[28924]_  = A201 & ~A200;
  assign \new_[28925]_  = A199 & \new_[28924]_ ;
  assign \new_[28928]_  = ~A232 & ~A203;
  assign \new_[28931]_  = A234 & A233;
  assign \new_[28932]_  = \new_[28931]_  & \new_[28928]_ ;
  assign \new_[28933]_  = \new_[28932]_  & \new_[28925]_ ;
  assign \new_[28936]_  = ~A267 & A235;
  assign \new_[28939]_  = ~A298 & ~A269;
  assign \new_[28940]_  = \new_[28939]_  & \new_[28936]_ ;
  assign \new_[28943]_  = ~A300 & A299;
  assign \new_[28946]_  = A302 & ~A301;
  assign \new_[28947]_  = \new_[28946]_  & \new_[28943]_ ;
  assign \new_[28948]_  = \new_[28947]_  & \new_[28940]_ ;
  assign \new_[28952]_  = A201 & ~A200;
  assign \new_[28953]_  = A199 & \new_[28952]_ ;
  assign \new_[28956]_  = ~A232 & ~A203;
  assign \new_[28959]_  = A234 & A233;
  assign \new_[28960]_  = \new_[28959]_  & \new_[28956]_ ;
  assign \new_[28961]_  = \new_[28960]_  & \new_[28953]_ ;
  assign \new_[28964]_  = A265 & A235;
  assign \new_[28967]_  = A298 & A266;
  assign \new_[28968]_  = \new_[28967]_  & \new_[28964]_ ;
  assign \new_[28971]_  = ~A300 & ~A299;
  assign \new_[28974]_  = A302 & ~A301;
  assign \new_[28975]_  = \new_[28974]_  & \new_[28971]_ ;
  assign \new_[28976]_  = \new_[28975]_  & \new_[28968]_ ;
  assign \new_[28980]_  = A201 & ~A200;
  assign \new_[28981]_  = A199 & \new_[28980]_ ;
  assign \new_[28984]_  = ~A232 & ~A203;
  assign \new_[28987]_  = A234 & A233;
  assign \new_[28988]_  = \new_[28987]_  & \new_[28984]_ ;
  assign \new_[28989]_  = \new_[28988]_  & \new_[28981]_ ;
  assign \new_[28992]_  = A265 & A235;
  assign \new_[28995]_  = ~A298 & A266;
  assign \new_[28996]_  = \new_[28995]_  & \new_[28992]_ ;
  assign \new_[28999]_  = ~A300 & A299;
  assign \new_[29002]_  = A302 & ~A301;
  assign \new_[29003]_  = \new_[29002]_  & \new_[28999]_ ;
  assign \new_[29004]_  = \new_[29003]_  & \new_[28996]_ ;
  assign \new_[29008]_  = A201 & ~A200;
  assign \new_[29009]_  = A199 & \new_[29008]_ ;
  assign \new_[29012]_  = ~A232 & ~A203;
  assign \new_[29015]_  = A234 & A233;
  assign \new_[29016]_  = \new_[29015]_  & \new_[29012]_ ;
  assign \new_[29017]_  = \new_[29016]_  & \new_[29009]_ ;
  assign \new_[29020]_  = ~A265 & A235;
  assign \new_[29023]_  = A298 & ~A266;
  assign \new_[29024]_  = \new_[29023]_  & \new_[29020]_ ;
  assign \new_[29027]_  = ~A300 & ~A299;
  assign \new_[29030]_  = A302 & ~A301;
  assign \new_[29031]_  = \new_[29030]_  & \new_[29027]_ ;
  assign \new_[29032]_  = \new_[29031]_  & \new_[29024]_ ;
  assign \new_[29036]_  = A201 & ~A200;
  assign \new_[29037]_  = A199 & \new_[29036]_ ;
  assign \new_[29040]_  = ~A232 & ~A203;
  assign \new_[29043]_  = A234 & A233;
  assign \new_[29044]_  = \new_[29043]_  & \new_[29040]_ ;
  assign \new_[29045]_  = \new_[29044]_  & \new_[29037]_ ;
  assign \new_[29048]_  = ~A265 & A235;
  assign \new_[29051]_  = ~A298 & ~A266;
  assign \new_[29052]_  = \new_[29051]_  & \new_[29048]_ ;
  assign \new_[29055]_  = ~A300 & A299;
  assign \new_[29058]_  = A302 & ~A301;
  assign \new_[29059]_  = \new_[29058]_  & \new_[29055]_ ;
  assign \new_[29060]_  = \new_[29059]_  & \new_[29052]_ ;
  assign \new_[29064]_  = A201 & ~A200;
  assign \new_[29065]_  = A199 & \new_[29064]_ ;
  assign \new_[29068]_  = ~A232 & ~A203;
  assign \new_[29071]_  = A234 & A233;
  assign \new_[29072]_  = \new_[29071]_  & \new_[29068]_ ;
  assign \new_[29073]_  = \new_[29072]_  & \new_[29065]_ ;
  assign \new_[29076]_  = A267 & ~A236;
  assign \new_[29079]_  = A269 & ~A268;
  assign \new_[29080]_  = \new_[29079]_  & \new_[29076]_ ;
  assign \new_[29083]_  = ~A299 & A298;
  assign \new_[29086]_  = A301 & A300;
  assign \new_[29087]_  = \new_[29086]_  & \new_[29083]_ ;
  assign \new_[29088]_  = \new_[29087]_  & \new_[29080]_ ;
  assign \new_[29092]_  = A201 & ~A200;
  assign \new_[29093]_  = A199 & \new_[29092]_ ;
  assign \new_[29096]_  = ~A232 & ~A203;
  assign \new_[29099]_  = A234 & A233;
  assign \new_[29100]_  = \new_[29099]_  & \new_[29096]_ ;
  assign \new_[29101]_  = \new_[29100]_  & \new_[29093]_ ;
  assign \new_[29104]_  = A267 & ~A236;
  assign \new_[29107]_  = A269 & ~A268;
  assign \new_[29108]_  = \new_[29107]_  & \new_[29104]_ ;
  assign \new_[29111]_  = ~A299 & A298;
  assign \new_[29114]_  = ~A302 & A300;
  assign \new_[29115]_  = \new_[29114]_  & \new_[29111]_ ;
  assign \new_[29116]_  = \new_[29115]_  & \new_[29108]_ ;
  assign \new_[29120]_  = A201 & ~A200;
  assign \new_[29121]_  = A199 & \new_[29120]_ ;
  assign \new_[29124]_  = ~A232 & ~A203;
  assign \new_[29127]_  = A234 & A233;
  assign \new_[29128]_  = \new_[29127]_  & \new_[29124]_ ;
  assign \new_[29129]_  = \new_[29128]_  & \new_[29121]_ ;
  assign \new_[29132]_  = A267 & ~A236;
  assign \new_[29135]_  = A269 & ~A268;
  assign \new_[29136]_  = \new_[29135]_  & \new_[29132]_ ;
  assign \new_[29139]_  = A299 & ~A298;
  assign \new_[29142]_  = A301 & A300;
  assign \new_[29143]_  = \new_[29142]_  & \new_[29139]_ ;
  assign \new_[29144]_  = \new_[29143]_  & \new_[29136]_ ;
  assign \new_[29148]_  = A201 & ~A200;
  assign \new_[29149]_  = A199 & \new_[29148]_ ;
  assign \new_[29152]_  = ~A232 & ~A203;
  assign \new_[29155]_  = A234 & A233;
  assign \new_[29156]_  = \new_[29155]_  & \new_[29152]_ ;
  assign \new_[29157]_  = \new_[29156]_  & \new_[29149]_ ;
  assign \new_[29160]_  = A267 & ~A236;
  assign \new_[29163]_  = A269 & ~A268;
  assign \new_[29164]_  = \new_[29163]_  & \new_[29160]_ ;
  assign \new_[29167]_  = A299 & ~A298;
  assign \new_[29170]_  = ~A302 & A300;
  assign \new_[29171]_  = \new_[29170]_  & \new_[29167]_ ;
  assign \new_[29172]_  = \new_[29171]_  & \new_[29164]_ ;
  assign \new_[29176]_  = A201 & ~A200;
  assign \new_[29177]_  = A199 & \new_[29176]_ ;
  assign \new_[29180]_  = ~A232 & ~A203;
  assign \new_[29183]_  = A234 & A233;
  assign \new_[29184]_  = \new_[29183]_  & \new_[29180]_ ;
  assign \new_[29185]_  = \new_[29184]_  & \new_[29177]_ ;
  assign \new_[29188]_  = ~A267 & ~A236;
  assign \new_[29191]_  = A298 & A268;
  assign \new_[29192]_  = \new_[29191]_  & \new_[29188]_ ;
  assign \new_[29195]_  = ~A300 & ~A299;
  assign \new_[29198]_  = A302 & ~A301;
  assign \new_[29199]_  = \new_[29198]_  & \new_[29195]_ ;
  assign \new_[29200]_  = \new_[29199]_  & \new_[29192]_ ;
  assign \new_[29204]_  = A201 & ~A200;
  assign \new_[29205]_  = A199 & \new_[29204]_ ;
  assign \new_[29208]_  = ~A232 & ~A203;
  assign \new_[29211]_  = A234 & A233;
  assign \new_[29212]_  = \new_[29211]_  & \new_[29208]_ ;
  assign \new_[29213]_  = \new_[29212]_  & \new_[29205]_ ;
  assign \new_[29216]_  = ~A267 & ~A236;
  assign \new_[29219]_  = ~A298 & A268;
  assign \new_[29220]_  = \new_[29219]_  & \new_[29216]_ ;
  assign \new_[29223]_  = ~A300 & A299;
  assign \new_[29226]_  = A302 & ~A301;
  assign \new_[29227]_  = \new_[29226]_  & \new_[29223]_ ;
  assign \new_[29228]_  = \new_[29227]_  & \new_[29220]_ ;
  assign \new_[29232]_  = A201 & ~A200;
  assign \new_[29233]_  = A199 & \new_[29232]_ ;
  assign \new_[29236]_  = ~A232 & ~A203;
  assign \new_[29239]_  = A234 & A233;
  assign \new_[29240]_  = \new_[29239]_  & \new_[29236]_ ;
  assign \new_[29241]_  = \new_[29240]_  & \new_[29233]_ ;
  assign \new_[29244]_  = ~A267 & ~A236;
  assign \new_[29247]_  = A298 & ~A269;
  assign \new_[29248]_  = \new_[29247]_  & \new_[29244]_ ;
  assign \new_[29251]_  = ~A300 & ~A299;
  assign \new_[29254]_  = A302 & ~A301;
  assign \new_[29255]_  = \new_[29254]_  & \new_[29251]_ ;
  assign \new_[29256]_  = \new_[29255]_  & \new_[29248]_ ;
  assign \new_[29260]_  = A201 & ~A200;
  assign \new_[29261]_  = A199 & \new_[29260]_ ;
  assign \new_[29264]_  = ~A232 & ~A203;
  assign \new_[29267]_  = A234 & A233;
  assign \new_[29268]_  = \new_[29267]_  & \new_[29264]_ ;
  assign \new_[29269]_  = \new_[29268]_  & \new_[29261]_ ;
  assign \new_[29272]_  = ~A267 & ~A236;
  assign \new_[29275]_  = ~A298 & ~A269;
  assign \new_[29276]_  = \new_[29275]_  & \new_[29272]_ ;
  assign \new_[29279]_  = ~A300 & A299;
  assign \new_[29282]_  = A302 & ~A301;
  assign \new_[29283]_  = \new_[29282]_  & \new_[29279]_ ;
  assign \new_[29284]_  = \new_[29283]_  & \new_[29276]_ ;
  assign \new_[29288]_  = A201 & ~A200;
  assign \new_[29289]_  = A199 & \new_[29288]_ ;
  assign \new_[29292]_  = ~A232 & ~A203;
  assign \new_[29295]_  = A234 & A233;
  assign \new_[29296]_  = \new_[29295]_  & \new_[29292]_ ;
  assign \new_[29297]_  = \new_[29296]_  & \new_[29289]_ ;
  assign \new_[29300]_  = A265 & ~A236;
  assign \new_[29303]_  = A298 & A266;
  assign \new_[29304]_  = \new_[29303]_  & \new_[29300]_ ;
  assign \new_[29307]_  = ~A300 & ~A299;
  assign \new_[29310]_  = A302 & ~A301;
  assign \new_[29311]_  = \new_[29310]_  & \new_[29307]_ ;
  assign \new_[29312]_  = \new_[29311]_  & \new_[29304]_ ;
  assign \new_[29316]_  = A201 & ~A200;
  assign \new_[29317]_  = A199 & \new_[29316]_ ;
  assign \new_[29320]_  = ~A232 & ~A203;
  assign \new_[29323]_  = A234 & A233;
  assign \new_[29324]_  = \new_[29323]_  & \new_[29320]_ ;
  assign \new_[29325]_  = \new_[29324]_  & \new_[29317]_ ;
  assign \new_[29328]_  = A265 & ~A236;
  assign \new_[29331]_  = ~A298 & A266;
  assign \new_[29332]_  = \new_[29331]_  & \new_[29328]_ ;
  assign \new_[29335]_  = ~A300 & A299;
  assign \new_[29338]_  = A302 & ~A301;
  assign \new_[29339]_  = \new_[29338]_  & \new_[29335]_ ;
  assign \new_[29340]_  = \new_[29339]_  & \new_[29332]_ ;
  assign \new_[29344]_  = A201 & ~A200;
  assign \new_[29345]_  = A199 & \new_[29344]_ ;
  assign \new_[29348]_  = ~A232 & ~A203;
  assign \new_[29351]_  = A234 & A233;
  assign \new_[29352]_  = \new_[29351]_  & \new_[29348]_ ;
  assign \new_[29353]_  = \new_[29352]_  & \new_[29345]_ ;
  assign \new_[29356]_  = ~A265 & ~A236;
  assign \new_[29359]_  = A298 & ~A266;
  assign \new_[29360]_  = \new_[29359]_  & \new_[29356]_ ;
  assign \new_[29363]_  = ~A300 & ~A299;
  assign \new_[29366]_  = A302 & ~A301;
  assign \new_[29367]_  = \new_[29366]_  & \new_[29363]_ ;
  assign \new_[29368]_  = \new_[29367]_  & \new_[29360]_ ;
  assign \new_[29372]_  = A201 & ~A200;
  assign \new_[29373]_  = A199 & \new_[29372]_ ;
  assign \new_[29376]_  = ~A232 & ~A203;
  assign \new_[29379]_  = A234 & A233;
  assign \new_[29380]_  = \new_[29379]_  & \new_[29376]_ ;
  assign \new_[29381]_  = \new_[29380]_  & \new_[29373]_ ;
  assign \new_[29384]_  = ~A265 & ~A236;
  assign \new_[29387]_  = ~A298 & ~A266;
  assign \new_[29388]_  = \new_[29387]_  & \new_[29384]_ ;
  assign \new_[29391]_  = ~A300 & A299;
  assign \new_[29394]_  = A302 & ~A301;
  assign \new_[29395]_  = \new_[29394]_  & \new_[29391]_ ;
  assign \new_[29396]_  = \new_[29395]_  & \new_[29388]_ ;
  assign \new_[29400]_  = A201 & ~A200;
  assign \new_[29401]_  = A199 & \new_[29400]_ ;
  assign \new_[29404]_  = ~A232 & ~A203;
  assign \new_[29407]_  = ~A234 & A233;
  assign \new_[29408]_  = \new_[29407]_  & \new_[29404]_ ;
  assign \new_[29409]_  = \new_[29408]_  & \new_[29401]_ ;
  assign \new_[29412]_  = A236 & ~A235;
  assign \new_[29415]_  = A268 & ~A267;
  assign \new_[29416]_  = \new_[29415]_  & \new_[29412]_ ;
  assign \new_[29419]_  = ~A299 & A298;
  assign \new_[29422]_  = A301 & A300;
  assign \new_[29423]_  = \new_[29422]_  & \new_[29419]_ ;
  assign \new_[29424]_  = \new_[29423]_  & \new_[29416]_ ;
  assign \new_[29428]_  = A201 & ~A200;
  assign \new_[29429]_  = A199 & \new_[29428]_ ;
  assign \new_[29432]_  = ~A232 & ~A203;
  assign \new_[29435]_  = ~A234 & A233;
  assign \new_[29436]_  = \new_[29435]_  & \new_[29432]_ ;
  assign \new_[29437]_  = \new_[29436]_  & \new_[29429]_ ;
  assign \new_[29440]_  = A236 & ~A235;
  assign \new_[29443]_  = A268 & ~A267;
  assign \new_[29444]_  = \new_[29443]_  & \new_[29440]_ ;
  assign \new_[29447]_  = ~A299 & A298;
  assign \new_[29450]_  = ~A302 & A300;
  assign \new_[29451]_  = \new_[29450]_  & \new_[29447]_ ;
  assign \new_[29452]_  = \new_[29451]_  & \new_[29444]_ ;
  assign \new_[29456]_  = A201 & ~A200;
  assign \new_[29457]_  = A199 & \new_[29456]_ ;
  assign \new_[29460]_  = ~A232 & ~A203;
  assign \new_[29463]_  = ~A234 & A233;
  assign \new_[29464]_  = \new_[29463]_  & \new_[29460]_ ;
  assign \new_[29465]_  = \new_[29464]_  & \new_[29457]_ ;
  assign \new_[29468]_  = A236 & ~A235;
  assign \new_[29471]_  = A268 & ~A267;
  assign \new_[29472]_  = \new_[29471]_  & \new_[29468]_ ;
  assign \new_[29475]_  = A299 & ~A298;
  assign \new_[29478]_  = A301 & A300;
  assign \new_[29479]_  = \new_[29478]_  & \new_[29475]_ ;
  assign \new_[29480]_  = \new_[29479]_  & \new_[29472]_ ;
  assign \new_[29484]_  = A201 & ~A200;
  assign \new_[29485]_  = A199 & \new_[29484]_ ;
  assign \new_[29488]_  = ~A232 & ~A203;
  assign \new_[29491]_  = ~A234 & A233;
  assign \new_[29492]_  = \new_[29491]_  & \new_[29488]_ ;
  assign \new_[29493]_  = \new_[29492]_  & \new_[29485]_ ;
  assign \new_[29496]_  = A236 & ~A235;
  assign \new_[29499]_  = A268 & ~A267;
  assign \new_[29500]_  = \new_[29499]_  & \new_[29496]_ ;
  assign \new_[29503]_  = A299 & ~A298;
  assign \new_[29506]_  = ~A302 & A300;
  assign \new_[29507]_  = \new_[29506]_  & \new_[29503]_ ;
  assign \new_[29508]_  = \new_[29507]_  & \new_[29500]_ ;
  assign \new_[29512]_  = A201 & ~A200;
  assign \new_[29513]_  = A199 & \new_[29512]_ ;
  assign \new_[29516]_  = ~A232 & ~A203;
  assign \new_[29519]_  = ~A234 & A233;
  assign \new_[29520]_  = \new_[29519]_  & \new_[29516]_ ;
  assign \new_[29521]_  = \new_[29520]_  & \new_[29513]_ ;
  assign \new_[29524]_  = A236 & ~A235;
  assign \new_[29527]_  = ~A269 & ~A267;
  assign \new_[29528]_  = \new_[29527]_  & \new_[29524]_ ;
  assign \new_[29531]_  = ~A299 & A298;
  assign \new_[29534]_  = A301 & A300;
  assign \new_[29535]_  = \new_[29534]_  & \new_[29531]_ ;
  assign \new_[29536]_  = \new_[29535]_  & \new_[29528]_ ;
  assign \new_[29540]_  = A201 & ~A200;
  assign \new_[29541]_  = A199 & \new_[29540]_ ;
  assign \new_[29544]_  = ~A232 & ~A203;
  assign \new_[29547]_  = ~A234 & A233;
  assign \new_[29548]_  = \new_[29547]_  & \new_[29544]_ ;
  assign \new_[29549]_  = \new_[29548]_  & \new_[29541]_ ;
  assign \new_[29552]_  = A236 & ~A235;
  assign \new_[29555]_  = ~A269 & ~A267;
  assign \new_[29556]_  = \new_[29555]_  & \new_[29552]_ ;
  assign \new_[29559]_  = ~A299 & A298;
  assign \new_[29562]_  = ~A302 & A300;
  assign \new_[29563]_  = \new_[29562]_  & \new_[29559]_ ;
  assign \new_[29564]_  = \new_[29563]_  & \new_[29556]_ ;
  assign \new_[29568]_  = A201 & ~A200;
  assign \new_[29569]_  = A199 & \new_[29568]_ ;
  assign \new_[29572]_  = ~A232 & ~A203;
  assign \new_[29575]_  = ~A234 & A233;
  assign \new_[29576]_  = \new_[29575]_  & \new_[29572]_ ;
  assign \new_[29577]_  = \new_[29576]_  & \new_[29569]_ ;
  assign \new_[29580]_  = A236 & ~A235;
  assign \new_[29583]_  = ~A269 & ~A267;
  assign \new_[29584]_  = \new_[29583]_  & \new_[29580]_ ;
  assign \new_[29587]_  = A299 & ~A298;
  assign \new_[29590]_  = A301 & A300;
  assign \new_[29591]_  = \new_[29590]_  & \new_[29587]_ ;
  assign \new_[29592]_  = \new_[29591]_  & \new_[29584]_ ;
  assign \new_[29596]_  = A201 & ~A200;
  assign \new_[29597]_  = A199 & \new_[29596]_ ;
  assign \new_[29600]_  = ~A232 & ~A203;
  assign \new_[29603]_  = ~A234 & A233;
  assign \new_[29604]_  = \new_[29603]_  & \new_[29600]_ ;
  assign \new_[29605]_  = \new_[29604]_  & \new_[29597]_ ;
  assign \new_[29608]_  = A236 & ~A235;
  assign \new_[29611]_  = ~A269 & ~A267;
  assign \new_[29612]_  = \new_[29611]_  & \new_[29608]_ ;
  assign \new_[29615]_  = A299 & ~A298;
  assign \new_[29618]_  = ~A302 & A300;
  assign \new_[29619]_  = \new_[29618]_  & \new_[29615]_ ;
  assign \new_[29620]_  = \new_[29619]_  & \new_[29612]_ ;
  assign \new_[29624]_  = A201 & ~A200;
  assign \new_[29625]_  = A199 & \new_[29624]_ ;
  assign \new_[29628]_  = ~A232 & ~A203;
  assign \new_[29631]_  = ~A234 & A233;
  assign \new_[29632]_  = \new_[29631]_  & \new_[29628]_ ;
  assign \new_[29633]_  = \new_[29632]_  & \new_[29625]_ ;
  assign \new_[29636]_  = A236 & ~A235;
  assign \new_[29639]_  = A266 & A265;
  assign \new_[29640]_  = \new_[29639]_  & \new_[29636]_ ;
  assign \new_[29643]_  = ~A299 & A298;
  assign \new_[29646]_  = A301 & A300;
  assign \new_[29647]_  = \new_[29646]_  & \new_[29643]_ ;
  assign \new_[29648]_  = \new_[29647]_  & \new_[29640]_ ;
  assign \new_[29652]_  = A201 & ~A200;
  assign \new_[29653]_  = A199 & \new_[29652]_ ;
  assign \new_[29656]_  = ~A232 & ~A203;
  assign \new_[29659]_  = ~A234 & A233;
  assign \new_[29660]_  = \new_[29659]_  & \new_[29656]_ ;
  assign \new_[29661]_  = \new_[29660]_  & \new_[29653]_ ;
  assign \new_[29664]_  = A236 & ~A235;
  assign \new_[29667]_  = A266 & A265;
  assign \new_[29668]_  = \new_[29667]_  & \new_[29664]_ ;
  assign \new_[29671]_  = ~A299 & A298;
  assign \new_[29674]_  = ~A302 & A300;
  assign \new_[29675]_  = \new_[29674]_  & \new_[29671]_ ;
  assign \new_[29676]_  = \new_[29675]_  & \new_[29668]_ ;
  assign \new_[29680]_  = A201 & ~A200;
  assign \new_[29681]_  = A199 & \new_[29680]_ ;
  assign \new_[29684]_  = ~A232 & ~A203;
  assign \new_[29687]_  = ~A234 & A233;
  assign \new_[29688]_  = \new_[29687]_  & \new_[29684]_ ;
  assign \new_[29689]_  = \new_[29688]_  & \new_[29681]_ ;
  assign \new_[29692]_  = A236 & ~A235;
  assign \new_[29695]_  = A266 & A265;
  assign \new_[29696]_  = \new_[29695]_  & \new_[29692]_ ;
  assign \new_[29699]_  = A299 & ~A298;
  assign \new_[29702]_  = A301 & A300;
  assign \new_[29703]_  = \new_[29702]_  & \new_[29699]_ ;
  assign \new_[29704]_  = \new_[29703]_  & \new_[29696]_ ;
  assign \new_[29708]_  = A201 & ~A200;
  assign \new_[29709]_  = A199 & \new_[29708]_ ;
  assign \new_[29712]_  = ~A232 & ~A203;
  assign \new_[29715]_  = ~A234 & A233;
  assign \new_[29716]_  = \new_[29715]_  & \new_[29712]_ ;
  assign \new_[29717]_  = \new_[29716]_  & \new_[29709]_ ;
  assign \new_[29720]_  = A236 & ~A235;
  assign \new_[29723]_  = A266 & A265;
  assign \new_[29724]_  = \new_[29723]_  & \new_[29720]_ ;
  assign \new_[29727]_  = A299 & ~A298;
  assign \new_[29730]_  = ~A302 & A300;
  assign \new_[29731]_  = \new_[29730]_  & \new_[29727]_ ;
  assign \new_[29732]_  = \new_[29731]_  & \new_[29724]_ ;
  assign \new_[29736]_  = A201 & ~A200;
  assign \new_[29737]_  = A199 & \new_[29736]_ ;
  assign \new_[29740]_  = ~A232 & ~A203;
  assign \new_[29743]_  = ~A234 & A233;
  assign \new_[29744]_  = \new_[29743]_  & \new_[29740]_ ;
  assign \new_[29745]_  = \new_[29744]_  & \new_[29737]_ ;
  assign \new_[29748]_  = A236 & ~A235;
  assign \new_[29751]_  = ~A266 & ~A265;
  assign \new_[29752]_  = \new_[29751]_  & \new_[29748]_ ;
  assign \new_[29755]_  = ~A299 & A298;
  assign \new_[29758]_  = A301 & A300;
  assign \new_[29759]_  = \new_[29758]_  & \new_[29755]_ ;
  assign \new_[29760]_  = \new_[29759]_  & \new_[29752]_ ;
  assign \new_[29764]_  = A201 & ~A200;
  assign \new_[29765]_  = A199 & \new_[29764]_ ;
  assign \new_[29768]_  = ~A232 & ~A203;
  assign \new_[29771]_  = ~A234 & A233;
  assign \new_[29772]_  = \new_[29771]_  & \new_[29768]_ ;
  assign \new_[29773]_  = \new_[29772]_  & \new_[29765]_ ;
  assign \new_[29776]_  = A236 & ~A235;
  assign \new_[29779]_  = ~A266 & ~A265;
  assign \new_[29780]_  = \new_[29779]_  & \new_[29776]_ ;
  assign \new_[29783]_  = ~A299 & A298;
  assign \new_[29786]_  = ~A302 & A300;
  assign \new_[29787]_  = \new_[29786]_  & \new_[29783]_ ;
  assign \new_[29788]_  = \new_[29787]_  & \new_[29780]_ ;
  assign \new_[29792]_  = A201 & ~A200;
  assign \new_[29793]_  = A199 & \new_[29792]_ ;
  assign \new_[29796]_  = ~A232 & ~A203;
  assign \new_[29799]_  = ~A234 & A233;
  assign \new_[29800]_  = \new_[29799]_  & \new_[29796]_ ;
  assign \new_[29801]_  = \new_[29800]_  & \new_[29793]_ ;
  assign \new_[29804]_  = A236 & ~A235;
  assign \new_[29807]_  = ~A266 & ~A265;
  assign \new_[29808]_  = \new_[29807]_  & \new_[29804]_ ;
  assign \new_[29811]_  = A299 & ~A298;
  assign \new_[29814]_  = A301 & A300;
  assign \new_[29815]_  = \new_[29814]_  & \new_[29811]_ ;
  assign \new_[29816]_  = \new_[29815]_  & \new_[29808]_ ;
  assign \new_[29820]_  = A201 & ~A200;
  assign \new_[29821]_  = A199 & \new_[29820]_ ;
  assign \new_[29824]_  = ~A232 & ~A203;
  assign \new_[29827]_  = ~A234 & A233;
  assign \new_[29828]_  = \new_[29827]_  & \new_[29824]_ ;
  assign \new_[29829]_  = \new_[29828]_  & \new_[29821]_ ;
  assign \new_[29832]_  = A236 & ~A235;
  assign \new_[29835]_  = ~A266 & ~A265;
  assign \new_[29836]_  = \new_[29835]_  & \new_[29832]_ ;
  assign \new_[29839]_  = A299 & ~A298;
  assign \new_[29842]_  = ~A302 & A300;
  assign \new_[29843]_  = \new_[29842]_  & \new_[29839]_ ;
  assign \new_[29844]_  = \new_[29843]_  & \new_[29836]_ ;
  assign \new_[29848]_  = A201 & ~A200;
  assign \new_[29849]_  = A199 & \new_[29848]_ ;
  assign \new_[29852]_  = A232 & ~A203;
  assign \new_[29855]_  = A234 & ~A233;
  assign \new_[29856]_  = \new_[29855]_  & \new_[29852]_ ;
  assign \new_[29857]_  = \new_[29856]_  & \new_[29849]_ ;
  assign \new_[29860]_  = A267 & A235;
  assign \new_[29863]_  = A269 & ~A268;
  assign \new_[29864]_  = \new_[29863]_  & \new_[29860]_ ;
  assign \new_[29867]_  = ~A299 & A298;
  assign \new_[29870]_  = A301 & A300;
  assign \new_[29871]_  = \new_[29870]_  & \new_[29867]_ ;
  assign \new_[29872]_  = \new_[29871]_  & \new_[29864]_ ;
  assign \new_[29876]_  = A201 & ~A200;
  assign \new_[29877]_  = A199 & \new_[29876]_ ;
  assign \new_[29880]_  = A232 & ~A203;
  assign \new_[29883]_  = A234 & ~A233;
  assign \new_[29884]_  = \new_[29883]_  & \new_[29880]_ ;
  assign \new_[29885]_  = \new_[29884]_  & \new_[29877]_ ;
  assign \new_[29888]_  = A267 & A235;
  assign \new_[29891]_  = A269 & ~A268;
  assign \new_[29892]_  = \new_[29891]_  & \new_[29888]_ ;
  assign \new_[29895]_  = ~A299 & A298;
  assign \new_[29898]_  = ~A302 & A300;
  assign \new_[29899]_  = \new_[29898]_  & \new_[29895]_ ;
  assign \new_[29900]_  = \new_[29899]_  & \new_[29892]_ ;
  assign \new_[29904]_  = A201 & ~A200;
  assign \new_[29905]_  = A199 & \new_[29904]_ ;
  assign \new_[29908]_  = A232 & ~A203;
  assign \new_[29911]_  = A234 & ~A233;
  assign \new_[29912]_  = \new_[29911]_  & \new_[29908]_ ;
  assign \new_[29913]_  = \new_[29912]_  & \new_[29905]_ ;
  assign \new_[29916]_  = A267 & A235;
  assign \new_[29919]_  = A269 & ~A268;
  assign \new_[29920]_  = \new_[29919]_  & \new_[29916]_ ;
  assign \new_[29923]_  = A299 & ~A298;
  assign \new_[29926]_  = A301 & A300;
  assign \new_[29927]_  = \new_[29926]_  & \new_[29923]_ ;
  assign \new_[29928]_  = \new_[29927]_  & \new_[29920]_ ;
  assign \new_[29932]_  = A201 & ~A200;
  assign \new_[29933]_  = A199 & \new_[29932]_ ;
  assign \new_[29936]_  = A232 & ~A203;
  assign \new_[29939]_  = A234 & ~A233;
  assign \new_[29940]_  = \new_[29939]_  & \new_[29936]_ ;
  assign \new_[29941]_  = \new_[29940]_  & \new_[29933]_ ;
  assign \new_[29944]_  = A267 & A235;
  assign \new_[29947]_  = A269 & ~A268;
  assign \new_[29948]_  = \new_[29947]_  & \new_[29944]_ ;
  assign \new_[29951]_  = A299 & ~A298;
  assign \new_[29954]_  = ~A302 & A300;
  assign \new_[29955]_  = \new_[29954]_  & \new_[29951]_ ;
  assign \new_[29956]_  = \new_[29955]_  & \new_[29948]_ ;
  assign \new_[29960]_  = A201 & ~A200;
  assign \new_[29961]_  = A199 & \new_[29960]_ ;
  assign \new_[29964]_  = A232 & ~A203;
  assign \new_[29967]_  = A234 & ~A233;
  assign \new_[29968]_  = \new_[29967]_  & \new_[29964]_ ;
  assign \new_[29969]_  = \new_[29968]_  & \new_[29961]_ ;
  assign \new_[29972]_  = ~A267 & A235;
  assign \new_[29975]_  = A298 & A268;
  assign \new_[29976]_  = \new_[29975]_  & \new_[29972]_ ;
  assign \new_[29979]_  = ~A300 & ~A299;
  assign \new_[29982]_  = A302 & ~A301;
  assign \new_[29983]_  = \new_[29982]_  & \new_[29979]_ ;
  assign \new_[29984]_  = \new_[29983]_  & \new_[29976]_ ;
  assign \new_[29988]_  = A201 & ~A200;
  assign \new_[29989]_  = A199 & \new_[29988]_ ;
  assign \new_[29992]_  = A232 & ~A203;
  assign \new_[29995]_  = A234 & ~A233;
  assign \new_[29996]_  = \new_[29995]_  & \new_[29992]_ ;
  assign \new_[29997]_  = \new_[29996]_  & \new_[29989]_ ;
  assign \new_[30000]_  = ~A267 & A235;
  assign \new_[30003]_  = ~A298 & A268;
  assign \new_[30004]_  = \new_[30003]_  & \new_[30000]_ ;
  assign \new_[30007]_  = ~A300 & A299;
  assign \new_[30010]_  = A302 & ~A301;
  assign \new_[30011]_  = \new_[30010]_  & \new_[30007]_ ;
  assign \new_[30012]_  = \new_[30011]_  & \new_[30004]_ ;
  assign \new_[30016]_  = A201 & ~A200;
  assign \new_[30017]_  = A199 & \new_[30016]_ ;
  assign \new_[30020]_  = A232 & ~A203;
  assign \new_[30023]_  = A234 & ~A233;
  assign \new_[30024]_  = \new_[30023]_  & \new_[30020]_ ;
  assign \new_[30025]_  = \new_[30024]_  & \new_[30017]_ ;
  assign \new_[30028]_  = ~A267 & A235;
  assign \new_[30031]_  = A298 & ~A269;
  assign \new_[30032]_  = \new_[30031]_  & \new_[30028]_ ;
  assign \new_[30035]_  = ~A300 & ~A299;
  assign \new_[30038]_  = A302 & ~A301;
  assign \new_[30039]_  = \new_[30038]_  & \new_[30035]_ ;
  assign \new_[30040]_  = \new_[30039]_  & \new_[30032]_ ;
  assign \new_[30044]_  = A201 & ~A200;
  assign \new_[30045]_  = A199 & \new_[30044]_ ;
  assign \new_[30048]_  = A232 & ~A203;
  assign \new_[30051]_  = A234 & ~A233;
  assign \new_[30052]_  = \new_[30051]_  & \new_[30048]_ ;
  assign \new_[30053]_  = \new_[30052]_  & \new_[30045]_ ;
  assign \new_[30056]_  = ~A267 & A235;
  assign \new_[30059]_  = ~A298 & ~A269;
  assign \new_[30060]_  = \new_[30059]_  & \new_[30056]_ ;
  assign \new_[30063]_  = ~A300 & A299;
  assign \new_[30066]_  = A302 & ~A301;
  assign \new_[30067]_  = \new_[30066]_  & \new_[30063]_ ;
  assign \new_[30068]_  = \new_[30067]_  & \new_[30060]_ ;
  assign \new_[30072]_  = A201 & ~A200;
  assign \new_[30073]_  = A199 & \new_[30072]_ ;
  assign \new_[30076]_  = A232 & ~A203;
  assign \new_[30079]_  = A234 & ~A233;
  assign \new_[30080]_  = \new_[30079]_  & \new_[30076]_ ;
  assign \new_[30081]_  = \new_[30080]_  & \new_[30073]_ ;
  assign \new_[30084]_  = A265 & A235;
  assign \new_[30087]_  = A298 & A266;
  assign \new_[30088]_  = \new_[30087]_  & \new_[30084]_ ;
  assign \new_[30091]_  = ~A300 & ~A299;
  assign \new_[30094]_  = A302 & ~A301;
  assign \new_[30095]_  = \new_[30094]_  & \new_[30091]_ ;
  assign \new_[30096]_  = \new_[30095]_  & \new_[30088]_ ;
  assign \new_[30100]_  = A201 & ~A200;
  assign \new_[30101]_  = A199 & \new_[30100]_ ;
  assign \new_[30104]_  = A232 & ~A203;
  assign \new_[30107]_  = A234 & ~A233;
  assign \new_[30108]_  = \new_[30107]_  & \new_[30104]_ ;
  assign \new_[30109]_  = \new_[30108]_  & \new_[30101]_ ;
  assign \new_[30112]_  = A265 & A235;
  assign \new_[30115]_  = ~A298 & A266;
  assign \new_[30116]_  = \new_[30115]_  & \new_[30112]_ ;
  assign \new_[30119]_  = ~A300 & A299;
  assign \new_[30122]_  = A302 & ~A301;
  assign \new_[30123]_  = \new_[30122]_  & \new_[30119]_ ;
  assign \new_[30124]_  = \new_[30123]_  & \new_[30116]_ ;
  assign \new_[30128]_  = A201 & ~A200;
  assign \new_[30129]_  = A199 & \new_[30128]_ ;
  assign \new_[30132]_  = A232 & ~A203;
  assign \new_[30135]_  = A234 & ~A233;
  assign \new_[30136]_  = \new_[30135]_  & \new_[30132]_ ;
  assign \new_[30137]_  = \new_[30136]_  & \new_[30129]_ ;
  assign \new_[30140]_  = ~A265 & A235;
  assign \new_[30143]_  = A298 & ~A266;
  assign \new_[30144]_  = \new_[30143]_  & \new_[30140]_ ;
  assign \new_[30147]_  = ~A300 & ~A299;
  assign \new_[30150]_  = A302 & ~A301;
  assign \new_[30151]_  = \new_[30150]_  & \new_[30147]_ ;
  assign \new_[30152]_  = \new_[30151]_  & \new_[30144]_ ;
  assign \new_[30156]_  = A201 & ~A200;
  assign \new_[30157]_  = A199 & \new_[30156]_ ;
  assign \new_[30160]_  = A232 & ~A203;
  assign \new_[30163]_  = A234 & ~A233;
  assign \new_[30164]_  = \new_[30163]_  & \new_[30160]_ ;
  assign \new_[30165]_  = \new_[30164]_  & \new_[30157]_ ;
  assign \new_[30168]_  = ~A265 & A235;
  assign \new_[30171]_  = ~A298 & ~A266;
  assign \new_[30172]_  = \new_[30171]_  & \new_[30168]_ ;
  assign \new_[30175]_  = ~A300 & A299;
  assign \new_[30178]_  = A302 & ~A301;
  assign \new_[30179]_  = \new_[30178]_  & \new_[30175]_ ;
  assign \new_[30180]_  = \new_[30179]_  & \new_[30172]_ ;
  assign \new_[30184]_  = A201 & ~A200;
  assign \new_[30185]_  = A199 & \new_[30184]_ ;
  assign \new_[30188]_  = A232 & ~A203;
  assign \new_[30191]_  = A234 & ~A233;
  assign \new_[30192]_  = \new_[30191]_  & \new_[30188]_ ;
  assign \new_[30193]_  = \new_[30192]_  & \new_[30185]_ ;
  assign \new_[30196]_  = A267 & ~A236;
  assign \new_[30199]_  = A269 & ~A268;
  assign \new_[30200]_  = \new_[30199]_  & \new_[30196]_ ;
  assign \new_[30203]_  = ~A299 & A298;
  assign \new_[30206]_  = A301 & A300;
  assign \new_[30207]_  = \new_[30206]_  & \new_[30203]_ ;
  assign \new_[30208]_  = \new_[30207]_  & \new_[30200]_ ;
  assign \new_[30212]_  = A201 & ~A200;
  assign \new_[30213]_  = A199 & \new_[30212]_ ;
  assign \new_[30216]_  = A232 & ~A203;
  assign \new_[30219]_  = A234 & ~A233;
  assign \new_[30220]_  = \new_[30219]_  & \new_[30216]_ ;
  assign \new_[30221]_  = \new_[30220]_  & \new_[30213]_ ;
  assign \new_[30224]_  = A267 & ~A236;
  assign \new_[30227]_  = A269 & ~A268;
  assign \new_[30228]_  = \new_[30227]_  & \new_[30224]_ ;
  assign \new_[30231]_  = ~A299 & A298;
  assign \new_[30234]_  = ~A302 & A300;
  assign \new_[30235]_  = \new_[30234]_  & \new_[30231]_ ;
  assign \new_[30236]_  = \new_[30235]_  & \new_[30228]_ ;
  assign \new_[30240]_  = A201 & ~A200;
  assign \new_[30241]_  = A199 & \new_[30240]_ ;
  assign \new_[30244]_  = A232 & ~A203;
  assign \new_[30247]_  = A234 & ~A233;
  assign \new_[30248]_  = \new_[30247]_  & \new_[30244]_ ;
  assign \new_[30249]_  = \new_[30248]_  & \new_[30241]_ ;
  assign \new_[30252]_  = A267 & ~A236;
  assign \new_[30255]_  = A269 & ~A268;
  assign \new_[30256]_  = \new_[30255]_  & \new_[30252]_ ;
  assign \new_[30259]_  = A299 & ~A298;
  assign \new_[30262]_  = A301 & A300;
  assign \new_[30263]_  = \new_[30262]_  & \new_[30259]_ ;
  assign \new_[30264]_  = \new_[30263]_  & \new_[30256]_ ;
  assign \new_[30268]_  = A201 & ~A200;
  assign \new_[30269]_  = A199 & \new_[30268]_ ;
  assign \new_[30272]_  = A232 & ~A203;
  assign \new_[30275]_  = A234 & ~A233;
  assign \new_[30276]_  = \new_[30275]_  & \new_[30272]_ ;
  assign \new_[30277]_  = \new_[30276]_  & \new_[30269]_ ;
  assign \new_[30280]_  = A267 & ~A236;
  assign \new_[30283]_  = A269 & ~A268;
  assign \new_[30284]_  = \new_[30283]_  & \new_[30280]_ ;
  assign \new_[30287]_  = A299 & ~A298;
  assign \new_[30290]_  = ~A302 & A300;
  assign \new_[30291]_  = \new_[30290]_  & \new_[30287]_ ;
  assign \new_[30292]_  = \new_[30291]_  & \new_[30284]_ ;
  assign \new_[30296]_  = A201 & ~A200;
  assign \new_[30297]_  = A199 & \new_[30296]_ ;
  assign \new_[30300]_  = A232 & ~A203;
  assign \new_[30303]_  = A234 & ~A233;
  assign \new_[30304]_  = \new_[30303]_  & \new_[30300]_ ;
  assign \new_[30305]_  = \new_[30304]_  & \new_[30297]_ ;
  assign \new_[30308]_  = ~A267 & ~A236;
  assign \new_[30311]_  = A298 & A268;
  assign \new_[30312]_  = \new_[30311]_  & \new_[30308]_ ;
  assign \new_[30315]_  = ~A300 & ~A299;
  assign \new_[30318]_  = A302 & ~A301;
  assign \new_[30319]_  = \new_[30318]_  & \new_[30315]_ ;
  assign \new_[30320]_  = \new_[30319]_  & \new_[30312]_ ;
  assign \new_[30324]_  = A201 & ~A200;
  assign \new_[30325]_  = A199 & \new_[30324]_ ;
  assign \new_[30328]_  = A232 & ~A203;
  assign \new_[30331]_  = A234 & ~A233;
  assign \new_[30332]_  = \new_[30331]_  & \new_[30328]_ ;
  assign \new_[30333]_  = \new_[30332]_  & \new_[30325]_ ;
  assign \new_[30336]_  = ~A267 & ~A236;
  assign \new_[30339]_  = ~A298 & A268;
  assign \new_[30340]_  = \new_[30339]_  & \new_[30336]_ ;
  assign \new_[30343]_  = ~A300 & A299;
  assign \new_[30346]_  = A302 & ~A301;
  assign \new_[30347]_  = \new_[30346]_  & \new_[30343]_ ;
  assign \new_[30348]_  = \new_[30347]_  & \new_[30340]_ ;
  assign \new_[30352]_  = A201 & ~A200;
  assign \new_[30353]_  = A199 & \new_[30352]_ ;
  assign \new_[30356]_  = A232 & ~A203;
  assign \new_[30359]_  = A234 & ~A233;
  assign \new_[30360]_  = \new_[30359]_  & \new_[30356]_ ;
  assign \new_[30361]_  = \new_[30360]_  & \new_[30353]_ ;
  assign \new_[30364]_  = ~A267 & ~A236;
  assign \new_[30367]_  = A298 & ~A269;
  assign \new_[30368]_  = \new_[30367]_  & \new_[30364]_ ;
  assign \new_[30371]_  = ~A300 & ~A299;
  assign \new_[30374]_  = A302 & ~A301;
  assign \new_[30375]_  = \new_[30374]_  & \new_[30371]_ ;
  assign \new_[30376]_  = \new_[30375]_  & \new_[30368]_ ;
  assign \new_[30380]_  = A201 & ~A200;
  assign \new_[30381]_  = A199 & \new_[30380]_ ;
  assign \new_[30384]_  = A232 & ~A203;
  assign \new_[30387]_  = A234 & ~A233;
  assign \new_[30388]_  = \new_[30387]_  & \new_[30384]_ ;
  assign \new_[30389]_  = \new_[30388]_  & \new_[30381]_ ;
  assign \new_[30392]_  = ~A267 & ~A236;
  assign \new_[30395]_  = ~A298 & ~A269;
  assign \new_[30396]_  = \new_[30395]_  & \new_[30392]_ ;
  assign \new_[30399]_  = ~A300 & A299;
  assign \new_[30402]_  = A302 & ~A301;
  assign \new_[30403]_  = \new_[30402]_  & \new_[30399]_ ;
  assign \new_[30404]_  = \new_[30403]_  & \new_[30396]_ ;
  assign \new_[30408]_  = A201 & ~A200;
  assign \new_[30409]_  = A199 & \new_[30408]_ ;
  assign \new_[30412]_  = A232 & ~A203;
  assign \new_[30415]_  = A234 & ~A233;
  assign \new_[30416]_  = \new_[30415]_  & \new_[30412]_ ;
  assign \new_[30417]_  = \new_[30416]_  & \new_[30409]_ ;
  assign \new_[30420]_  = A265 & ~A236;
  assign \new_[30423]_  = A298 & A266;
  assign \new_[30424]_  = \new_[30423]_  & \new_[30420]_ ;
  assign \new_[30427]_  = ~A300 & ~A299;
  assign \new_[30430]_  = A302 & ~A301;
  assign \new_[30431]_  = \new_[30430]_  & \new_[30427]_ ;
  assign \new_[30432]_  = \new_[30431]_  & \new_[30424]_ ;
  assign \new_[30436]_  = A201 & ~A200;
  assign \new_[30437]_  = A199 & \new_[30436]_ ;
  assign \new_[30440]_  = A232 & ~A203;
  assign \new_[30443]_  = A234 & ~A233;
  assign \new_[30444]_  = \new_[30443]_  & \new_[30440]_ ;
  assign \new_[30445]_  = \new_[30444]_  & \new_[30437]_ ;
  assign \new_[30448]_  = A265 & ~A236;
  assign \new_[30451]_  = ~A298 & A266;
  assign \new_[30452]_  = \new_[30451]_  & \new_[30448]_ ;
  assign \new_[30455]_  = ~A300 & A299;
  assign \new_[30458]_  = A302 & ~A301;
  assign \new_[30459]_  = \new_[30458]_  & \new_[30455]_ ;
  assign \new_[30460]_  = \new_[30459]_  & \new_[30452]_ ;
  assign \new_[30464]_  = A201 & ~A200;
  assign \new_[30465]_  = A199 & \new_[30464]_ ;
  assign \new_[30468]_  = A232 & ~A203;
  assign \new_[30471]_  = A234 & ~A233;
  assign \new_[30472]_  = \new_[30471]_  & \new_[30468]_ ;
  assign \new_[30473]_  = \new_[30472]_  & \new_[30465]_ ;
  assign \new_[30476]_  = ~A265 & ~A236;
  assign \new_[30479]_  = A298 & ~A266;
  assign \new_[30480]_  = \new_[30479]_  & \new_[30476]_ ;
  assign \new_[30483]_  = ~A300 & ~A299;
  assign \new_[30486]_  = A302 & ~A301;
  assign \new_[30487]_  = \new_[30486]_  & \new_[30483]_ ;
  assign \new_[30488]_  = \new_[30487]_  & \new_[30480]_ ;
  assign \new_[30492]_  = A201 & ~A200;
  assign \new_[30493]_  = A199 & \new_[30492]_ ;
  assign \new_[30496]_  = A232 & ~A203;
  assign \new_[30499]_  = A234 & ~A233;
  assign \new_[30500]_  = \new_[30499]_  & \new_[30496]_ ;
  assign \new_[30501]_  = \new_[30500]_  & \new_[30493]_ ;
  assign \new_[30504]_  = ~A265 & ~A236;
  assign \new_[30507]_  = ~A298 & ~A266;
  assign \new_[30508]_  = \new_[30507]_  & \new_[30504]_ ;
  assign \new_[30511]_  = ~A300 & A299;
  assign \new_[30514]_  = A302 & ~A301;
  assign \new_[30515]_  = \new_[30514]_  & \new_[30511]_ ;
  assign \new_[30516]_  = \new_[30515]_  & \new_[30508]_ ;
  assign \new_[30520]_  = A201 & ~A200;
  assign \new_[30521]_  = A199 & \new_[30520]_ ;
  assign \new_[30524]_  = A232 & ~A203;
  assign \new_[30527]_  = ~A234 & ~A233;
  assign \new_[30528]_  = \new_[30527]_  & \new_[30524]_ ;
  assign \new_[30529]_  = \new_[30528]_  & \new_[30521]_ ;
  assign \new_[30532]_  = A236 & ~A235;
  assign \new_[30535]_  = A268 & ~A267;
  assign \new_[30536]_  = \new_[30535]_  & \new_[30532]_ ;
  assign \new_[30539]_  = ~A299 & A298;
  assign \new_[30542]_  = A301 & A300;
  assign \new_[30543]_  = \new_[30542]_  & \new_[30539]_ ;
  assign \new_[30544]_  = \new_[30543]_  & \new_[30536]_ ;
  assign \new_[30548]_  = A201 & ~A200;
  assign \new_[30549]_  = A199 & \new_[30548]_ ;
  assign \new_[30552]_  = A232 & ~A203;
  assign \new_[30555]_  = ~A234 & ~A233;
  assign \new_[30556]_  = \new_[30555]_  & \new_[30552]_ ;
  assign \new_[30557]_  = \new_[30556]_  & \new_[30549]_ ;
  assign \new_[30560]_  = A236 & ~A235;
  assign \new_[30563]_  = A268 & ~A267;
  assign \new_[30564]_  = \new_[30563]_  & \new_[30560]_ ;
  assign \new_[30567]_  = ~A299 & A298;
  assign \new_[30570]_  = ~A302 & A300;
  assign \new_[30571]_  = \new_[30570]_  & \new_[30567]_ ;
  assign \new_[30572]_  = \new_[30571]_  & \new_[30564]_ ;
  assign \new_[30576]_  = A201 & ~A200;
  assign \new_[30577]_  = A199 & \new_[30576]_ ;
  assign \new_[30580]_  = A232 & ~A203;
  assign \new_[30583]_  = ~A234 & ~A233;
  assign \new_[30584]_  = \new_[30583]_  & \new_[30580]_ ;
  assign \new_[30585]_  = \new_[30584]_  & \new_[30577]_ ;
  assign \new_[30588]_  = A236 & ~A235;
  assign \new_[30591]_  = A268 & ~A267;
  assign \new_[30592]_  = \new_[30591]_  & \new_[30588]_ ;
  assign \new_[30595]_  = A299 & ~A298;
  assign \new_[30598]_  = A301 & A300;
  assign \new_[30599]_  = \new_[30598]_  & \new_[30595]_ ;
  assign \new_[30600]_  = \new_[30599]_  & \new_[30592]_ ;
  assign \new_[30604]_  = A201 & ~A200;
  assign \new_[30605]_  = A199 & \new_[30604]_ ;
  assign \new_[30608]_  = A232 & ~A203;
  assign \new_[30611]_  = ~A234 & ~A233;
  assign \new_[30612]_  = \new_[30611]_  & \new_[30608]_ ;
  assign \new_[30613]_  = \new_[30612]_  & \new_[30605]_ ;
  assign \new_[30616]_  = A236 & ~A235;
  assign \new_[30619]_  = A268 & ~A267;
  assign \new_[30620]_  = \new_[30619]_  & \new_[30616]_ ;
  assign \new_[30623]_  = A299 & ~A298;
  assign \new_[30626]_  = ~A302 & A300;
  assign \new_[30627]_  = \new_[30626]_  & \new_[30623]_ ;
  assign \new_[30628]_  = \new_[30627]_  & \new_[30620]_ ;
  assign \new_[30632]_  = A201 & ~A200;
  assign \new_[30633]_  = A199 & \new_[30632]_ ;
  assign \new_[30636]_  = A232 & ~A203;
  assign \new_[30639]_  = ~A234 & ~A233;
  assign \new_[30640]_  = \new_[30639]_  & \new_[30636]_ ;
  assign \new_[30641]_  = \new_[30640]_  & \new_[30633]_ ;
  assign \new_[30644]_  = A236 & ~A235;
  assign \new_[30647]_  = ~A269 & ~A267;
  assign \new_[30648]_  = \new_[30647]_  & \new_[30644]_ ;
  assign \new_[30651]_  = ~A299 & A298;
  assign \new_[30654]_  = A301 & A300;
  assign \new_[30655]_  = \new_[30654]_  & \new_[30651]_ ;
  assign \new_[30656]_  = \new_[30655]_  & \new_[30648]_ ;
  assign \new_[30660]_  = A201 & ~A200;
  assign \new_[30661]_  = A199 & \new_[30660]_ ;
  assign \new_[30664]_  = A232 & ~A203;
  assign \new_[30667]_  = ~A234 & ~A233;
  assign \new_[30668]_  = \new_[30667]_  & \new_[30664]_ ;
  assign \new_[30669]_  = \new_[30668]_  & \new_[30661]_ ;
  assign \new_[30672]_  = A236 & ~A235;
  assign \new_[30675]_  = ~A269 & ~A267;
  assign \new_[30676]_  = \new_[30675]_  & \new_[30672]_ ;
  assign \new_[30679]_  = ~A299 & A298;
  assign \new_[30682]_  = ~A302 & A300;
  assign \new_[30683]_  = \new_[30682]_  & \new_[30679]_ ;
  assign \new_[30684]_  = \new_[30683]_  & \new_[30676]_ ;
  assign \new_[30688]_  = A201 & ~A200;
  assign \new_[30689]_  = A199 & \new_[30688]_ ;
  assign \new_[30692]_  = A232 & ~A203;
  assign \new_[30695]_  = ~A234 & ~A233;
  assign \new_[30696]_  = \new_[30695]_  & \new_[30692]_ ;
  assign \new_[30697]_  = \new_[30696]_  & \new_[30689]_ ;
  assign \new_[30700]_  = A236 & ~A235;
  assign \new_[30703]_  = ~A269 & ~A267;
  assign \new_[30704]_  = \new_[30703]_  & \new_[30700]_ ;
  assign \new_[30707]_  = A299 & ~A298;
  assign \new_[30710]_  = A301 & A300;
  assign \new_[30711]_  = \new_[30710]_  & \new_[30707]_ ;
  assign \new_[30712]_  = \new_[30711]_  & \new_[30704]_ ;
  assign \new_[30716]_  = A201 & ~A200;
  assign \new_[30717]_  = A199 & \new_[30716]_ ;
  assign \new_[30720]_  = A232 & ~A203;
  assign \new_[30723]_  = ~A234 & ~A233;
  assign \new_[30724]_  = \new_[30723]_  & \new_[30720]_ ;
  assign \new_[30725]_  = \new_[30724]_  & \new_[30717]_ ;
  assign \new_[30728]_  = A236 & ~A235;
  assign \new_[30731]_  = ~A269 & ~A267;
  assign \new_[30732]_  = \new_[30731]_  & \new_[30728]_ ;
  assign \new_[30735]_  = A299 & ~A298;
  assign \new_[30738]_  = ~A302 & A300;
  assign \new_[30739]_  = \new_[30738]_  & \new_[30735]_ ;
  assign \new_[30740]_  = \new_[30739]_  & \new_[30732]_ ;
  assign \new_[30744]_  = A201 & ~A200;
  assign \new_[30745]_  = A199 & \new_[30744]_ ;
  assign \new_[30748]_  = A232 & ~A203;
  assign \new_[30751]_  = ~A234 & ~A233;
  assign \new_[30752]_  = \new_[30751]_  & \new_[30748]_ ;
  assign \new_[30753]_  = \new_[30752]_  & \new_[30745]_ ;
  assign \new_[30756]_  = A236 & ~A235;
  assign \new_[30759]_  = A266 & A265;
  assign \new_[30760]_  = \new_[30759]_  & \new_[30756]_ ;
  assign \new_[30763]_  = ~A299 & A298;
  assign \new_[30766]_  = A301 & A300;
  assign \new_[30767]_  = \new_[30766]_  & \new_[30763]_ ;
  assign \new_[30768]_  = \new_[30767]_  & \new_[30760]_ ;
  assign \new_[30772]_  = A201 & ~A200;
  assign \new_[30773]_  = A199 & \new_[30772]_ ;
  assign \new_[30776]_  = A232 & ~A203;
  assign \new_[30779]_  = ~A234 & ~A233;
  assign \new_[30780]_  = \new_[30779]_  & \new_[30776]_ ;
  assign \new_[30781]_  = \new_[30780]_  & \new_[30773]_ ;
  assign \new_[30784]_  = A236 & ~A235;
  assign \new_[30787]_  = A266 & A265;
  assign \new_[30788]_  = \new_[30787]_  & \new_[30784]_ ;
  assign \new_[30791]_  = ~A299 & A298;
  assign \new_[30794]_  = ~A302 & A300;
  assign \new_[30795]_  = \new_[30794]_  & \new_[30791]_ ;
  assign \new_[30796]_  = \new_[30795]_  & \new_[30788]_ ;
  assign \new_[30800]_  = A201 & ~A200;
  assign \new_[30801]_  = A199 & \new_[30800]_ ;
  assign \new_[30804]_  = A232 & ~A203;
  assign \new_[30807]_  = ~A234 & ~A233;
  assign \new_[30808]_  = \new_[30807]_  & \new_[30804]_ ;
  assign \new_[30809]_  = \new_[30808]_  & \new_[30801]_ ;
  assign \new_[30812]_  = A236 & ~A235;
  assign \new_[30815]_  = A266 & A265;
  assign \new_[30816]_  = \new_[30815]_  & \new_[30812]_ ;
  assign \new_[30819]_  = A299 & ~A298;
  assign \new_[30822]_  = A301 & A300;
  assign \new_[30823]_  = \new_[30822]_  & \new_[30819]_ ;
  assign \new_[30824]_  = \new_[30823]_  & \new_[30816]_ ;
  assign \new_[30828]_  = A201 & ~A200;
  assign \new_[30829]_  = A199 & \new_[30828]_ ;
  assign \new_[30832]_  = A232 & ~A203;
  assign \new_[30835]_  = ~A234 & ~A233;
  assign \new_[30836]_  = \new_[30835]_  & \new_[30832]_ ;
  assign \new_[30837]_  = \new_[30836]_  & \new_[30829]_ ;
  assign \new_[30840]_  = A236 & ~A235;
  assign \new_[30843]_  = A266 & A265;
  assign \new_[30844]_  = \new_[30843]_  & \new_[30840]_ ;
  assign \new_[30847]_  = A299 & ~A298;
  assign \new_[30850]_  = ~A302 & A300;
  assign \new_[30851]_  = \new_[30850]_  & \new_[30847]_ ;
  assign \new_[30852]_  = \new_[30851]_  & \new_[30844]_ ;
  assign \new_[30856]_  = A201 & ~A200;
  assign \new_[30857]_  = A199 & \new_[30856]_ ;
  assign \new_[30860]_  = A232 & ~A203;
  assign \new_[30863]_  = ~A234 & ~A233;
  assign \new_[30864]_  = \new_[30863]_  & \new_[30860]_ ;
  assign \new_[30865]_  = \new_[30864]_  & \new_[30857]_ ;
  assign \new_[30868]_  = A236 & ~A235;
  assign \new_[30871]_  = ~A266 & ~A265;
  assign \new_[30872]_  = \new_[30871]_  & \new_[30868]_ ;
  assign \new_[30875]_  = ~A299 & A298;
  assign \new_[30878]_  = A301 & A300;
  assign \new_[30879]_  = \new_[30878]_  & \new_[30875]_ ;
  assign \new_[30880]_  = \new_[30879]_  & \new_[30872]_ ;
  assign \new_[30884]_  = A201 & ~A200;
  assign \new_[30885]_  = A199 & \new_[30884]_ ;
  assign \new_[30888]_  = A232 & ~A203;
  assign \new_[30891]_  = ~A234 & ~A233;
  assign \new_[30892]_  = \new_[30891]_  & \new_[30888]_ ;
  assign \new_[30893]_  = \new_[30892]_  & \new_[30885]_ ;
  assign \new_[30896]_  = A236 & ~A235;
  assign \new_[30899]_  = ~A266 & ~A265;
  assign \new_[30900]_  = \new_[30899]_  & \new_[30896]_ ;
  assign \new_[30903]_  = ~A299 & A298;
  assign \new_[30906]_  = ~A302 & A300;
  assign \new_[30907]_  = \new_[30906]_  & \new_[30903]_ ;
  assign \new_[30908]_  = \new_[30907]_  & \new_[30900]_ ;
  assign \new_[30912]_  = A201 & ~A200;
  assign \new_[30913]_  = A199 & \new_[30912]_ ;
  assign \new_[30916]_  = A232 & ~A203;
  assign \new_[30919]_  = ~A234 & ~A233;
  assign \new_[30920]_  = \new_[30919]_  & \new_[30916]_ ;
  assign \new_[30921]_  = \new_[30920]_  & \new_[30913]_ ;
  assign \new_[30924]_  = A236 & ~A235;
  assign \new_[30927]_  = ~A266 & ~A265;
  assign \new_[30928]_  = \new_[30927]_  & \new_[30924]_ ;
  assign \new_[30931]_  = A299 & ~A298;
  assign \new_[30934]_  = A301 & A300;
  assign \new_[30935]_  = \new_[30934]_  & \new_[30931]_ ;
  assign \new_[30936]_  = \new_[30935]_  & \new_[30928]_ ;
  assign \new_[30940]_  = A201 & ~A200;
  assign \new_[30941]_  = A199 & \new_[30940]_ ;
  assign \new_[30944]_  = A232 & ~A203;
  assign \new_[30947]_  = ~A234 & ~A233;
  assign \new_[30948]_  = \new_[30947]_  & \new_[30944]_ ;
  assign \new_[30949]_  = \new_[30948]_  & \new_[30941]_ ;
  assign \new_[30952]_  = A236 & ~A235;
  assign \new_[30955]_  = ~A266 & ~A265;
  assign \new_[30956]_  = \new_[30955]_  & \new_[30952]_ ;
  assign \new_[30959]_  = A299 & ~A298;
  assign \new_[30962]_  = ~A302 & A300;
  assign \new_[30963]_  = \new_[30962]_  & \new_[30959]_ ;
  assign \new_[30964]_  = \new_[30963]_  & \new_[30956]_ ;
  assign \new_[30968]_  = ~A201 & ~A200;
  assign \new_[30969]_  = A199 & \new_[30968]_ ;
  assign \new_[30972]_  = A203 & ~A202;
  assign \new_[30975]_  = A233 & ~A232;
  assign \new_[30976]_  = \new_[30975]_  & \new_[30972]_ ;
  assign \new_[30977]_  = \new_[30976]_  & \new_[30969]_ ;
  assign \new_[30980]_  = A235 & A234;
  assign \new_[30983]_  = A268 & ~A267;
  assign \new_[30984]_  = \new_[30983]_  & \new_[30980]_ ;
  assign \new_[30987]_  = ~A299 & A298;
  assign \new_[30990]_  = A301 & A300;
  assign \new_[30991]_  = \new_[30990]_  & \new_[30987]_ ;
  assign \new_[30992]_  = \new_[30991]_  & \new_[30984]_ ;
  assign \new_[30996]_  = ~A201 & ~A200;
  assign \new_[30997]_  = A199 & \new_[30996]_ ;
  assign \new_[31000]_  = A203 & ~A202;
  assign \new_[31003]_  = A233 & ~A232;
  assign \new_[31004]_  = \new_[31003]_  & \new_[31000]_ ;
  assign \new_[31005]_  = \new_[31004]_  & \new_[30997]_ ;
  assign \new_[31008]_  = A235 & A234;
  assign \new_[31011]_  = A268 & ~A267;
  assign \new_[31012]_  = \new_[31011]_  & \new_[31008]_ ;
  assign \new_[31015]_  = ~A299 & A298;
  assign \new_[31018]_  = ~A302 & A300;
  assign \new_[31019]_  = \new_[31018]_  & \new_[31015]_ ;
  assign \new_[31020]_  = \new_[31019]_  & \new_[31012]_ ;
  assign \new_[31024]_  = ~A201 & ~A200;
  assign \new_[31025]_  = A199 & \new_[31024]_ ;
  assign \new_[31028]_  = A203 & ~A202;
  assign \new_[31031]_  = A233 & ~A232;
  assign \new_[31032]_  = \new_[31031]_  & \new_[31028]_ ;
  assign \new_[31033]_  = \new_[31032]_  & \new_[31025]_ ;
  assign \new_[31036]_  = A235 & A234;
  assign \new_[31039]_  = A268 & ~A267;
  assign \new_[31040]_  = \new_[31039]_  & \new_[31036]_ ;
  assign \new_[31043]_  = A299 & ~A298;
  assign \new_[31046]_  = A301 & A300;
  assign \new_[31047]_  = \new_[31046]_  & \new_[31043]_ ;
  assign \new_[31048]_  = \new_[31047]_  & \new_[31040]_ ;
  assign \new_[31052]_  = ~A201 & ~A200;
  assign \new_[31053]_  = A199 & \new_[31052]_ ;
  assign \new_[31056]_  = A203 & ~A202;
  assign \new_[31059]_  = A233 & ~A232;
  assign \new_[31060]_  = \new_[31059]_  & \new_[31056]_ ;
  assign \new_[31061]_  = \new_[31060]_  & \new_[31053]_ ;
  assign \new_[31064]_  = A235 & A234;
  assign \new_[31067]_  = A268 & ~A267;
  assign \new_[31068]_  = \new_[31067]_  & \new_[31064]_ ;
  assign \new_[31071]_  = A299 & ~A298;
  assign \new_[31074]_  = ~A302 & A300;
  assign \new_[31075]_  = \new_[31074]_  & \new_[31071]_ ;
  assign \new_[31076]_  = \new_[31075]_  & \new_[31068]_ ;
  assign \new_[31080]_  = ~A201 & ~A200;
  assign \new_[31081]_  = A199 & \new_[31080]_ ;
  assign \new_[31084]_  = A203 & ~A202;
  assign \new_[31087]_  = A233 & ~A232;
  assign \new_[31088]_  = \new_[31087]_  & \new_[31084]_ ;
  assign \new_[31089]_  = \new_[31088]_  & \new_[31081]_ ;
  assign \new_[31092]_  = A235 & A234;
  assign \new_[31095]_  = ~A269 & ~A267;
  assign \new_[31096]_  = \new_[31095]_  & \new_[31092]_ ;
  assign \new_[31099]_  = ~A299 & A298;
  assign \new_[31102]_  = A301 & A300;
  assign \new_[31103]_  = \new_[31102]_  & \new_[31099]_ ;
  assign \new_[31104]_  = \new_[31103]_  & \new_[31096]_ ;
  assign \new_[31108]_  = ~A201 & ~A200;
  assign \new_[31109]_  = A199 & \new_[31108]_ ;
  assign \new_[31112]_  = A203 & ~A202;
  assign \new_[31115]_  = A233 & ~A232;
  assign \new_[31116]_  = \new_[31115]_  & \new_[31112]_ ;
  assign \new_[31117]_  = \new_[31116]_  & \new_[31109]_ ;
  assign \new_[31120]_  = A235 & A234;
  assign \new_[31123]_  = ~A269 & ~A267;
  assign \new_[31124]_  = \new_[31123]_  & \new_[31120]_ ;
  assign \new_[31127]_  = ~A299 & A298;
  assign \new_[31130]_  = ~A302 & A300;
  assign \new_[31131]_  = \new_[31130]_  & \new_[31127]_ ;
  assign \new_[31132]_  = \new_[31131]_  & \new_[31124]_ ;
  assign \new_[31136]_  = ~A201 & ~A200;
  assign \new_[31137]_  = A199 & \new_[31136]_ ;
  assign \new_[31140]_  = A203 & ~A202;
  assign \new_[31143]_  = A233 & ~A232;
  assign \new_[31144]_  = \new_[31143]_  & \new_[31140]_ ;
  assign \new_[31145]_  = \new_[31144]_  & \new_[31137]_ ;
  assign \new_[31148]_  = A235 & A234;
  assign \new_[31151]_  = ~A269 & ~A267;
  assign \new_[31152]_  = \new_[31151]_  & \new_[31148]_ ;
  assign \new_[31155]_  = A299 & ~A298;
  assign \new_[31158]_  = A301 & A300;
  assign \new_[31159]_  = \new_[31158]_  & \new_[31155]_ ;
  assign \new_[31160]_  = \new_[31159]_  & \new_[31152]_ ;
  assign \new_[31164]_  = ~A201 & ~A200;
  assign \new_[31165]_  = A199 & \new_[31164]_ ;
  assign \new_[31168]_  = A203 & ~A202;
  assign \new_[31171]_  = A233 & ~A232;
  assign \new_[31172]_  = \new_[31171]_  & \new_[31168]_ ;
  assign \new_[31173]_  = \new_[31172]_  & \new_[31165]_ ;
  assign \new_[31176]_  = A235 & A234;
  assign \new_[31179]_  = ~A269 & ~A267;
  assign \new_[31180]_  = \new_[31179]_  & \new_[31176]_ ;
  assign \new_[31183]_  = A299 & ~A298;
  assign \new_[31186]_  = ~A302 & A300;
  assign \new_[31187]_  = \new_[31186]_  & \new_[31183]_ ;
  assign \new_[31188]_  = \new_[31187]_  & \new_[31180]_ ;
  assign \new_[31192]_  = ~A201 & ~A200;
  assign \new_[31193]_  = A199 & \new_[31192]_ ;
  assign \new_[31196]_  = A203 & ~A202;
  assign \new_[31199]_  = A233 & ~A232;
  assign \new_[31200]_  = \new_[31199]_  & \new_[31196]_ ;
  assign \new_[31201]_  = \new_[31200]_  & \new_[31193]_ ;
  assign \new_[31204]_  = A235 & A234;
  assign \new_[31207]_  = A266 & A265;
  assign \new_[31208]_  = \new_[31207]_  & \new_[31204]_ ;
  assign \new_[31211]_  = ~A299 & A298;
  assign \new_[31214]_  = A301 & A300;
  assign \new_[31215]_  = \new_[31214]_  & \new_[31211]_ ;
  assign \new_[31216]_  = \new_[31215]_  & \new_[31208]_ ;
  assign \new_[31220]_  = ~A201 & ~A200;
  assign \new_[31221]_  = A199 & \new_[31220]_ ;
  assign \new_[31224]_  = A203 & ~A202;
  assign \new_[31227]_  = A233 & ~A232;
  assign \new_[31228]_  = \new_[31227]_  & \new_[31224]_ ;
  assign \new_[31229]_  = \new_[31228]_  & \new_[31221]_ ;
  assign \new_[31232]_  = A235 & A234;
  assign \new_[31235]_  = A266 & A265;
  assign \new_[31236]_  = \new_[31235]_  & \new_[31232]_ ;
  assign \new_[31239]_  = ~A299 & A298;
  assign \new_[31242]_  = ~A302 & A300;
  assign \new_[31243]_  = \new_[31242]_  & \new_[31239]_ ;
  assign \new_[31244]_  = \new_[31243]_  & \new_[31236]_ ;
  assign \new_[31248]_  = ~A201 & ~A200;
  assign \new_[31249]_  = A199 & \new_[31248]_ ;
  assign \new_[31252]_  = A203 & ~A202;
  assign \new_[31255]_  = A233 & ~A232;
  assign \new_[31256]_  = \new_[31255]_  & \new_[31252]_ ;
  assign \new_[31257]_  = \new_[31256]_  & \new_[31249]_ ;
  assign \new_[31260]_  = A235 & A234;
  assign \new_[31263]_  = A266 & A265;
  assign \new_[31264]_  = \new_[31263]_  & \new_[31260]_ ;
  assign \new_[31267]_  = A299 & ~A298;
  assign \new_[31270]_  = A301 & A300;
  assign \new_[31271]_  = \new_[31270]_  & \new_[31267]_ ;
  assign \new_[31272]_  = \new_[31271]_  & \new_[31264]_ ;
  assign \new_[31276]_  = ~A201 & ~A200;
  assign \new_[31277]_  = A199 & \new_[31276]_ ;
  assign \new_[31280]_  = A203 & ~A202;
  assign \new_[31283]_  = A233 & ~A232;
  assign \new_[31284]_  = \new_[31283]_  & \new_[31280]_ ;
  assign \new_[31285]_  = \new_[31284]_  & \new_[31277]_ ;
  assign \new_[31288]_  = A235 & A234;
  assign \new_[31291]_  = A266 & A265;
  assign \new_[31292]_  = \new_[31291]_  & \new_[31288]_ ;
  assign \new_[31295]_  = A299 & ~A298;
  assign \new_[31298]_  = ~A302 & A300;
  assign \new_[31299]_  = \new_[31298]_  & \new_[31295]_ ;
  assign \new_[31300]_  = \new_[31299]_  & \new_[31292]_ ;
  assign \new_[31304]_  = ~A201 & ~A200;
  assign \new_[31305]_  = A199 & \new_[31304]_ ;
  assign \new_[31308]_  = A203 & ~A202;
  assign \new_[31311]_  = A233 & ~A232;
  assign \new_[31312]_  = \new_[31311]_  & \new_[31308]_ ;
  assign \new_[31313]_  = \new_[31312]_  & \new_[31305]_ ;
  assign \new_[31316]_  = A235 & A234;
  assign \new_[31319]_  = ~A266 & ~A265;
  assign \new_[31320]_  = \new_[31319]_  & \new_[31316]_ ;
  assign \new_[31323]_  = ~A299 & A298;
  assign \new_[31326]_  = A301 & A300;
  assign \new_[31327]_  = \new_[31326]_  & \new_[31323]_ ;
  assign \new_[31328]_  = \new_[31327]_  & \new_[31320]_ ;
  assign \new_[31332]_  = ~A201 & ~A200;
  assign \new_[31333]_  = A199 & \new_[31332]_ ;
  assign \new_[31336]_  = A203 & ~A202;
  assign \new_[31339]_  = A233 & ~A232;
  assign \new_[31340]_  = \new_[31339]_  & \new_[31336]_ ;
  assign \new_[31341]_  = \new_[31340]_  & \new_[31333]_ ;
  assign \new_[31344]_  = A235 & A234;
  assign \new_[31347]_  = ~A266 & ~A265;
  assign \new_[31348]_  = \new_[31347]_  & \new_[31344]_ ;
  assign \new_[31351]_  = ~A299 & A298;
  assign \new_[31354]_  = ~A302 & A300;
  assign \new_[31355]_  = \new_[31354]_  & \new_[31351]_ ;
  assign \new_[31356]_  = \new_[31355]_  & \new_[31348]_ ;
  assign \new_[31360]_  = ~A201 & ~A200;
  assign \new_[31361]_  = A199 & \new_[31360]_ ;
  assign \new_[31364]_  = A203 & ~A202;
  assign \new_[31367]_  = A233 & ~A232;
  assign \new_[31368]_  = \new_[31367]_  & \new_[31364]_ ;
  assign \new_[31369]_  = \new_[31368]_  & \new_[31361]_ ;
  assign \new_[31372]_  = A235 & A234;
  assign \new_[31375]_  = ~A266 & ~A265;
  assign \new_[31376]_  = \new_[31375]_  & \new_[31372]_ ;
  assign \new_[31379]_  = A299 & ~A298;
  assign \new_[31382]_  = A301 & A300;
  assign \new_[31383]_  = \new_[31382]_  & \new_[31379]_ ;
  assign \new_[31384]_  = \new_[31383]_  & \new_[31376]_ ;
  assign \new_[31388]_  = ~A201 & ~A200;
  assign \new_[31389]_  = A199 & \new_[31388]_ ;
  assign \new_[31392]_  = A203 & ~A202;
  assign \new_[31395]_  = A233 & ~A232;
  assign \new_[31396]_  = \new_[31395]_  & \new_[31392]_ ;
  assign \new_[31397]_  = \new_[31396]_  & \new_[31389]_ ;
  assign \new_[31400]_  = A235 & A234;
  assign \new_[31403]_  = ~A266 & ~A265;
  assign \new_[31404]_  = \new_[31403]_  & \new_[31400]_ ;
  assign \new_[31407]_  = A299 & ~A298;
  assign \new_[31410]_  = ~A302 & A300;
  assign \new_[31411]_  = \new_[31410]_  & \new_[31407]_ ;
  assign \new_[31412]_  = \new_[31411]_  & \new_[31404]_ ;
  assign \new_[31416]_  = ~A201 & ~A200;
  assign \new_[31417]_  = A199 & \new_[31416]_ ;
  assign \new_[31420]_  = A203 & ~A202;
  assign \new_[31423]_  = A233 & ~A232;
  assign \new_[31424]_  = \new_[31423]_  & \new_[31420]_ ;
  assign \new_[31425]_  = \new_[31424]_  & \new_[31417]_ ;
  assign \new_[31428]_  = ~A236 & A234;
  assign \new_[31431]_  = A268 & ~A267;
  assign \new_[31432]_  = \new_[31431]_  & \new_[31428]_ ;
  assign \new_[31435]_  = ~A299 & A298;
  assign \new_[31438]_  = A301 & A300;
  assign \new_[31439]_  = \new_[31438]_  & \new_[31435]_ ;
  assign \new_[31440]_  = \new_[31439]_  & \new_[31432]_ ;
  assign \new_[31444]_  = ~A201 & ~A200;
  assign \new_[31445]_  = A199 & \new_[31444]_ ;
  assign \new_[31448]_  = A203 & ~A202;
  assign \new_[31451]_  = A233 & ~A232;
  assign \new_[31452]_  = \new_[31451]_  & \new_[31448]_ ;
  assign \new_[31453]_  = \new_[31452]_  & \new_[31445]_ ;
  assign \new_[31456]_  = ~A236 & A234;
  assign \new_[31459]_  = A268 & ~A267;
  assign \new_[31460]_  = \new_[31459]_  & \new_[31456]_ ;
  assign \new_[31463]_  = ~A299 & A298;
  assign \new_[31466]_  = ~A302 & A300;
  assign \new_[31467]_  = \new_[31466]_  & \new_[31463]_ ;
  assign \new_[31468]_  = \new_[31467]_  & \new_[31460]_ ;
  assign \new_[31472]_  = ~A201 & ~A200;
  assign \new_[31473]_  = A199 & \new_[31472]_ ;
  assign \new_[31476]_  = A203 & ~A202;
  assign \new_[31479]_  = A233 & ~A232;
  assign \new_[31480]_  = \new_[31479]_  & \new_[31476]_ ;
  assign \new_[31481]_  = \new_[31480]_  & \new_[31473]_ ;
  assign \new_[31484]_  = ~A236 & A234;
  assign \new_[31487]_  = A268 & ~A267;
  assign \new_[31488]_  = \new_[31487]_  & \new_[31484]_ ;
  assign \new_[31491]_  = A299 & ~A298;
  assign \new_[31494]_  = A301 & A300;
  assign \new_[31495]_  = \new_[31494]_  & \new_[31491]_ ;
  assign \new_[31496]_  = \new_[31495]_  & \new_[31488]_ ;
  assign \new_[31500]_  = ~A201 & ~A200;
  assign \new_[31501]_  = A199 & \new_[31500]_ ;
  assign \new_[31504]_  = A203 & ~A202;
  assign \new_[31507]_  = A233 & ~A232;
  assign \new_[31508]_  = \new_[31507]_  & \new_[31504]_ ;
  assign \new_[31509]_  = \new_[31508]_  & \new_[31501]_ ;
  assign \new_[31512]_  = ~A236 & A234;
  assign \new_[31515]_  = A268 & ~A267;
  assign \new_[31516]_  = \new_[31515]_  & \new_[31512]_ ;
  assign \new_[31519]_  = A299 & ~A298;
  assign \new_[31522]_  = ~A302 & A300;
  assign \new_[31523]_  = \new_[31522]_  & \new_[31519]_ ;
  assign \new_[31524]_  = \new_[31523]_  & \new_[31516]_ ;
  assign \new_[31528]_  = ~A201 & ~A200;
  assign \new_[31529]_  = A199 & \new_[31528]_ ;
  assign \new_[31532]_  = A203 & ~A202;
  assign \new_[31535]_  = A233 & ~A232;
  assign \new_[31536]_  = \new_[31535]_  & \new_[31532]_ ;
  assign \new_[31537]_  = \new_[31536]_  & \new_[31529]_ ;
  assign \new_[31540]_  = ~A236 & A234;
  assign \new_[31543]_  = ~A269 & ~A267;
  assign \new_[31544]_  = \new_[31543]_  & \new_[31540]_ ;
  assign \new_[31547]_  = ~A299 & A298;
  assign \new_[31550]_  = A301 & A300;
  assign \new_[31551]_  = \new_[31550]_  & \new_[31547]_ ;
  assign \new_[31552]_  = \new_[31551]_  & \new_[31544]_ ;
  assign \new_[31556]_  = ~A201 & ~A200;
  assign \new_[31557]_  = A199 & \new_[31556]_ ;
  assign \new_[31560]_  = A203 & ~A202;
  assign \new_[31563]_  = A233 & ~A232;
  assign \new_[31564]_  = \new_[31563]_  & \new_[31560]_ ;
  assign \new_[31565]_  = \new_[31564]_  & \new_[31557]_ ;
  assign \new_[31568]_  = ~A236 & A234;
  assign \new_[31571]_  = ~A269 & ~A267;
  assign \new_[31572]_  = \new_[31571]_  & \new_[31568]_ ;
  assign \new_[31575]_  = ~A299 & A298;
  assign \new_[31578]_  = ~A302 & A300;
  assign \new_[31579]_  = \new_[31578]_  & \new_[31575]_ ;
  assign \new_[31580]_  = \new_[31579]_  & \new_[31572]_ ;
  assign \new_[31584]_  = ~A201 & ~A200;
  assign \new_[31585]_  = A199 & \new_[31584]_ ;
  assign \new_[31588]_  = A203 & ~A202;
  assign \new_[31591]_  = A233 & ~A232;
  assign \new_[31592]_  = \new_[31591]_  & \new_[31588]_ ;
  assign \new_[31593]_  = \new_[31592]_  & \new_[31585]_ ;
  assign \new_[31596]_  = ~A236 & A234;
  assign \new_[31599]_  = ~A269 & ~A267;
  assign \new_[31600]_  = \new_[31599]_  & \new_[31596]_ ;
  assign \new_[31603]_  = A299 & ~A298;
  assign \new_[31606]_  = A301 & A300;
  assign \new_[31607]_  = \new_[31606]_  & \new_[31603]_ ;
  assign \new_[31608]_  = \new_[31607]_  & \new_[31600]_ ;
  assign \new_[31612]_  = ~A201 & ~A200;
  assign \new_[31613]_  = A199 & \new_[31612]_ ;
  assign \new_[31616]_  = A203 & ~A202;
  assign \new_[31619]_  = A233 & ~A232;
  assign \new_[31620]_  = \new_[31619]_  & \new_[31616]_ ;
  assign \new_[31621]_  = \new_[31620]_  & \new_[31613]_ ;
  assign \new_[31624]_  = ~A236 & A234;
  assign \new_[31627]_  = ~A269 & ~A267;
  assign \new_[31628]_  = \new_[31627]_  & \new_[31624]_ ;
  assign \new_[31631]_  = A299 & ~A298;
  assign \new_[31634]_  = ~A302 & A300;
  assign \new_[31635]_  = \new_[31634]_  & \new_[31631]_ ;
  assign \new_[31636]_  = \new_[31635]_  & \new_[31628]_ ;
  assign \new_[31640]_  = ~A201 & ~A200;
  assign \new_[31641]_  = A199 & \new_[31640]_ ;
  assign \new_[31644]_  = A203 & ~A202;
  assign \new_[31647]_  = A233 & ~A232;
  assign \new_[31648]_  = \new_[31647]_  & \new_[31644]_ ;
  assign \new_[31649]_  = \new_[31648]_  & \new_[31641]_ ;
  assign \new_[31652]_  = ~A236 & A234;
  assign \new_[31655]_  = A266 & A265;
  assign \new_[31656]_  = \new_[31655]_  & \new_[31652]_ ;
  assign \new_[31659]_  = ~A299 & A298;
  assign \new_[31662]_  = A301 & A300;
  assign \new_[31663]_  = \new_[31662]_  & \new_[31659]_ ;
  assign \new_[31664]_  = \new_[31663]_  & \new_[31656]_ ;
  assign \new_[31668]_  = ~A201 & ~A200;
  assign \new_[31669]_  = A199 & \new_[31668]_ ;
  assign \new_[31672]_  = A203 & ~A202;
  assign \new_[31675]_  = A233 & ~A232;
  assign \new_[31676]_  = \new_[31675]_  & \new_[31672]_ ;
  assign \new_[31677]_  = \new_[31676]_  & \new_[31669]_ ;
  assign \new_[31680]_  = ~A236 & A234;
  assign \new_[31683]_  = A266 & A265;
  assign \new_[31684]_  = \new_[31683]_  & \new_[31680]_ ;
  assign \new_[31687]_  = ~A299 & A298;
  assign \new_[31690]_  = ~A302 & A300;
  assign \new_[31691]_  = \new_[31690]_  & \new_[31687]_ ;
  assign \new_[31692]_  = \new_[31691]_  & \new_[31684]_ ;
  assign \new_[31696]_  = ~A201 & ~A200;
  assign \new_[31697]_  = A199 & \new_[31696]_ ;
  assign \new_[31700]_  = A203 & ~A202;
  assign \new_[31703]_  = A233 & ~A232;
  assign \new_[31704]_  = \new_[31703]_  & \new_[31700]_ ;
  assign \new_[31705]_  = \new_[31704]_  & \new_[31697]_ ;
  assign \new_[31708]_  = ~A236 & A234;
  assign \new_[31711]_  = A266 & A265;
  assign \new_[31712]_  = \new_[31711]_  & \new_[31708]_ ;
  assign \new_[31715]_  = A299 & ~A298;
  assign \new_[31718]_  = A301 & A300;
  assign \new_[31719]_  = \new_[31718]_  & \new_[31715]_ ;
  assign \new_[31720]_  = \new_[31719]_  & \new_[31712]_ ;
  assign \new_[31724]_  = ~A201 & ~A200;
  assign \new_[31725]_  = A199 & \new_[31724]_ ;
  assign \new_[31728]_  = A203 & ~A202;
  assign \new_[31731]_  = A233 & ~A232;
  assign \new_[31732]_  = \new_[31731]_  & \new_[31728]_ ;
  assign \new_[31733]_  = \new_[31732]_  & \new_[31725]_ ;
  assign \new_[31736]_  = ~A236 & A234;
  assign \new_[31739]_  = A266 & A265;
  assign \new_[31740]_  = \new_[31739]_  & \new_[31736]_ ;
  assign \new_[31743]_  = A299 & ~A298;
  assign \new_[31746]_  = ~A302 & A300;
  assign \new_[31747]_  = \new_[31746]_  & \new_[31743]_ ;
  assign \new_[31748]_  = \new_[31747]_  & \new_[31740]_ ;
  assign \new_[31752]_  = ~A201 & ~A200;
  assign \new_[31753]_  = A199 & \new_[31752]_ ;
  assign \new_[31756]_  = A203 & ~A202;
  assign \new_[31759]_  = A233 & ~A232;
  assign \new_[31760]_  = \new_[31759]_  & \new_[31756]_ ;
  assign \new_[31761]_  = \new_[31760]_  & \new_[31753]_ ;
  assign \new_[31764]_  = ~A236 & A234;
  assign \new_[31767]_  = ~A266 & ~A265;
  assign \new_[31768]_  = \new_[31767]_  & \new_[31764]_ ;
  assign \new_[31771]_  = ~A299 & A298;
  assign \new_[31774]_  = A301 & A300;
  assign \new_[31775]_  = \new_[31774]_  & \new_[31771]_ ;
  assign \new_[31776]_  = \new_[31775]_  & \new_[31768]_ ;
  assign \new_[31780]_  = ~A201 & ~A200;
  assign \new_[31781]_  = A199 & \new_[31780]_ ;
  assign \new_[31784]_  = A203 & ~A202;
  assign \new_[31787]_  = A233 & ~A232;
  assign \new_[31788]_  = \new_[31787]_  & \new_[31784]_ ;
  assign \new_[31789]_  = \new_[31788]_  & \new_[31781]_ ;
  assign \new_[31792]_  = ~A236 & A234;
  assign \new_[31795]_  = ~A266 & ~A265;
  assign \new_[31796]_  = \new_[31795]_  & \new_[31792]_ ;
  assign \new_[31799]_  = ~A299 & A298;
  assign \new_[31802]_  = ~A302 & A300;
  assign \new_[31803]_  = \new_[31802]_  & \new_[31799]_ ;
  assign \new_[31804]_  = \new_[31803]_  & \new_[31796]_ ;
  assign \new_[31808]_  = ~A201 & ~A200;
  assign \new_[31809]_  = A199 & \new_[31808]_ ;
  assign \new_[31812]_  = A203 & ~A202;
  assign \new_[31815]_  = A233 & ~A232;
  assign \new_[31816]_  = \new_[31815]_  & \new_[31812]_ ;
  assign \new_[31817]_  = \new_[31816]_  & \new_[31809]_ ;
  assign \new_[31820]_  = ~A236 & A234;
  assign \new_[31823]_  = ~A266 & ~A265;
  assign \new_[31824]_  = \new_[31823]_  & \new_[31820]_ ;
  assign \new_[31827]_  = A299 & ~A298;
  assign \new_[31830]_  = A301 & A300;
  assign \new_[31831]_  = \new_[31830]_  & \new_[31827]_ ;
  assign \new_[31832]_  = \new_[31831]_  & \new_[31824]_ ;
  assign \new_[31836]_  = ~A201 & ~A200;
  assign \new_[31837]_  = A199 & \new_[31836]_ ;
  assign \new_[31840]_  = A203 & ~A202;
  assign \new_[31843]_  = A233 & ~A232;
  assign \new_[31844]_  = \new_[31843]_  & \new_[31840]_ ;
  assign \new_[31845]_  = \new_[31844]_  & \new_[31837]_ ;
  assign \new_[31848]_  = ~A236 & A234;
  assign \new_[31851]_  = ~A266 & ~A265;
  assign \new_[31852]_  = \new_[31851]_  & \new_[31848]_ ;
  assign \new_[31855]_  = A299 & ~A298;
  assign \new_[31858]_  = ~A302 & A300;
  assign \new_[31859]_  = \new_[31858]_  & \new_[31855]_ ;
  assign \new_[31860]_  = \new_[31859]_  & \new_[31852]_ ;
  assign \new_[31864]_  = ~A201 & ~A200;
  assign \new_[31865]_  = A199 & \new_[31864]_ ;
  assign \new_[31868]_  = A203 & ~A202;
  assign \new_[31871]_  = ~A233 & A232;
  assign \new_[31872]_  = \new_[31871]_  & \new_[31868]_ ;
  assign \new_[31873]_  = \new_[31872]_  & \new_[31865]_ ;
  assign \new_[31876]_  = A235 & A234;
  assign \new_[31879]_  = A268 & ~A267;
  assign \new_[31880]_  = \new_[31879]_  & \new_[31876]_ ;
  assign \new_[31883]_  = ~A299 & A298;
  assign \new_[31886]_  = A301 & A300;
  assign \new_[31887]_  = \new_[31886]_  & \new_[31883]_ ;
  assign \new_[31888]_  = \new_[31887]_  & \new_[31880]_ ;
  assign \new_[31892]_  = ~A201 & ~A200;
  assign \new_[31893]_  = A199 & \new_[31892]_ ;
  assign \new_[31896]_  = A203 & ~A202;
  assign \new_[31899]_  = ~A233 & A232;
  assign \new_[31900]_  = \new_[31899]_  & \new_[31896]_ ;
  assign \new_[31901]_  = \new_[31900]_  & \new_[31893]_ ;
  assign \new_[31904]_  = A235 & A234;
  assign \new_[31907]_  = A268 & ~A267;
  assign \new_[31908]_  = \new_[31907]_  & \new_[31904]_ ;
  assign \new_[31911]_  = ~A299 & A298;
  assign \new_[31914]_  = ~A302 & A300;
  assign \new_[31915]_  = \new_[31914]_  & \new_[31911]_ ;
  assign \new_[31916]_  = \new_[31915]_  & \new_[31908]_ ;
  assign \new_[31920]_  = ~A201 & ~A200;
  assign \new_[31921]_  = A199 & \new_[31920]_ ;
  assign \new_[31924]_  = A203 & ~A202;
  assign \new_[31927]_  = ~A233 & A232;
  assign \new_[31928]_  = \new_[31927]_  & \new_[31924]_ ;
  assign \new_[31929]_  = \new_[31928]_  & \new_[31921]_ ;
  assign \new_[31932]_  = A235 & A234;
  assign \new_[31935]_  = A268 & ~A267;
  assign \new_[31936]_  = \new_[31935]_  & \new_[31932]_ ;
  assign \new_[31939]_  = A299 & ~A298;
  assign \new_[31942]_  = A301 & A300;
  assign \new_[31943]_  = \new_[31942]_  & \new_[31939]_ ;
  assign \new_[31944]_  = \new_[31943]_  & \new_[31936]_ ;
  assign \new_[31948]_  = ~A201 & ~A200;
  assign \new_[31949]_  = A199 & \new_[31948]_ ;
  assign \new_[31952]_  = A203 & ~A202;
  assign \new_[31955]_  = ~A233 & A232;
  assign \new_[31956]_  = \new_[31955]_  & \new_[31952]_ ;
  assign \new_[31957]_  = \new_[31956]_  & \new_[31949]_ ;
  assign \new_[31960]_  = A235 & A234;
  assign \new_[31963]_  = A268 & ~A267;
  assign \new_[31964]_  = \new_[31963]_  & \new_[31960]_ ;
  assign \new_[31967]_  = A299 & ~A298;
  assign \new_[31970]_  = ~A302 & A300;
  assign \new_[31971]_  = \new_[31970]_  & \new_[31967]_ ;
  assign \new_[31972]_  = \new_[31971]_  & \new_[31964]_ ;
  assign \new_[31976]_  = ~A201 & ~A200;
  assign \new_[31977]_  = A199 & \new_[31976]_ ;
  assign \new_[31980]_  = A203 & ~A202;
  assign \new_[31983]_  = ~A233 & A232;
  assign \new_[31984]_  = \new_[31983]_  & \new_[31980]_ ;
  assign \new_[31985]_  = \new_[31984]_  & \new_[31977]_ ;
  assign \new_[31988]_  = A235 & A234;
  assign \new_[31991]_  = ~A269 & ~A267;
  assign \new_[31992]_  = \new_[31991]_  & \new_[31988]_ ;
  assign \new_[31995]_  = ~A299 & A298;
  assign \new_[31998]_  = A301 & A300;
  assign \new_[31999]_  = \new_[31998]_  & \new_[31995]_ ;
  assign \new_[32000]_  = \new_[31999]_  & \new_[31992]_ ;
  assign \new_[32004]_  = ~A201 & ~A200;
  assign \new_[32005]_  = A199 & \new_[32004]_ ;
  assign \new_[32008]_  = A203 & ~A202;
  assign \new_[32011]_  = ~A233 & A232;
  assign \new_[32012]_  = \new_[32011]_  & \new_[32008]_ ;
  assign \new_[32013]_  = \new_[32012]_  & \new_[32005]_ ;
  assign \new_[32016]_  = A235 & A234;
  assign \new_[32019]_  = ~A269 & ~A267;
  assign \new_[32020]_  = \new_[32019]_  & \new_[32016]_ ;
  assign \new_[32023]_  = ~A299 & A298;
  assign \new_[32026]_  = ~A302 & A300;
  assign \new_[32027]_  = \new_[32026]_  & \new_[32023]_ ;
  assign \new_[32028]_  = \new_[32027]_  & \new_[32020]_ ;
  assign \new_[32032]_  = ~A201 & ~A200;
  assign \new_[32033]_  = A199 & \new_[32032]_ ;
  assign \new_[32036]_  = A203 & ~A202;
  assign \new_[32039]_  = ~A233 & A232;
  assign \new_[32040]_  = \new_[32039]_  & \new_[32036]_ ;
  assign \new_[32041]_  = \new_[32040]_  & \new_[32033]_ ;
  assign \new_[32044]_  = A235 & A234;
  assign \new_[32047]_  = ~A269 & ~A267;
  assign \new_[32048]_  = \new_[32047]_  & \new_[32044]_ ;
  assign \new_[32051]_  = A299 & ~A298;
  assign \new_[32054]_  = A301 & A300;
  assign \new_[32055]_  = \new_[32054]_  & \new_[32051]_ ;
  assign \new_[32056]_  = \new_[32055]_  & \new_[32048]_ ;
  assign \new_[32060]_  = ~A201 & ~A200;
  assign \new_[32061]_  = A199 & \new_[32060]_ ;
  assign \new_[32064]_  = A203 & ~A202;
  assign \new_[32067]_  = ~A233 & A232;
  assign \new_[32068]_  = \new_[32067]_  & \new_[32064]_ ;
  assign \new_[32069]_  = \new_[32068]_  & \new_[32061]_ ;
  assign \new_[32072]_  = A235 & A234;
  assign \new_[32075]_  = ~A269 & ~A267;
  assign \new_[32076]_  = \new_[32075]_  & \new_[32072]_ ;
  assign \new_[32079]_  = A299 & ~A298;
  assign \new_[32082]_  = ~A302 & A300;
  assign \new_[32083]_  = \new_[32082]_  & \new_[32079]_ ;
  assign \new_[32084]_  = \new_[32083]_  & \new_[32076]_ ;
  assign \new_[32088]_  = ~A201 & ~A200;
  assign \new_[32089]_  = A199 & \new_[32088]_ ;
  assign \new_[32092]_  = A203 & ~A202;
  assign \new_[32095]_  = ~A233 & A232;
  assign \new_[32096]_  = \new_[32095]_  & \new_[32092]_ ;
  assign \new_[32097]_  = \new_[32096]_  & \new_[32089]_ ;
  assign \new_[32100]_  = A235 & A234;
  assign \new_[32103]_  = A266 & A265;
  assign \new_[32104]_  = \new_[32103]_  & \new_[32100]_ ;
  assign \new_[32107]_  = ~A299 & A298;
  assign \new_[32110]_  = A301 & A300;
  assign \new_[32111]_  = \new_[32110]_  & \new_[32107]_ ;
  assign \new_[32112]_  = \new_[32111]_  & \new_[32104]_ ;
  assign \new_[32116]_  = ~A201 & ~A200;
  assign \new_[32117]_  = A199 & \new_[32116]_ ;
  assign \new_[32120]_  = A203 & ~A202;
  assign \new_[32123]_  = ~A233 & A232;
  assign \new_[32124]_  = \new_[32123]_  & \new_[32120]_ ;
  assign \new_[32125]_  = \new_[32124]_  & \new_[32117]_ ;
  assign \new_[32128]_  = A235 & A234;
  assign \new_[32131]_  = A266 & A265;
  assign \new_[32132]_  = \new_[32131]_  & \new_[32128]_ ;
  assign \new_[32135]_  = ~A299 & A298;
  assign \new_[32138]_  = ~A302 & A300;
  assign \new_[32139]_  = \new_[32138]_  & \new_[32135]_ ;
  assign \new_[32140]_  = \new_[32139]_  & \new_[32132]_ ;
  assign \new_[32144]_  = ~A201 & ~A200;
  assign \new_[32145]_  = A199 & \new_[32144]_ ;
  assign \new_[32148]_  = A203 & ~A202;
  assign \new_[32151]_  = ~A233 & A232;
  assign \new_[32152]_  = \new_[32151]_  & \new_[32148]_ ;
  assign \new_[32153]_  = \new_[32152]_  & \new_[32145]_ ;
  assign \new_[32156]_  = A235 & A234;
  assign \new_[32159]_  = A266 & A265;
  assign \new_[32160]_  = \new_[32159]_  & \new_[32156]_ ;
  assign \new_[32163]_  = A299 & ~A298;
  assign \new_[32166]_  = A301 & A300;
  assign \new_[32167]_  = \new_[32166]_  & \new_[32163]_ ;
  assign \new_[32168]_  = \new_[32167]_  & \new_[32160]_ ;
  assign \new_[32172]_  = ~A201 & ~A200;
  assign \new_[32173]_  = A199 & \new_[32172]_ ;
  assign \new_[32176]_  = A203 & ~A202;
  assign \new_[32179]_  = ~A233 & A232;
  assign \new_[32180]_  = \new_[32179]_  & \new_[32176]_ ;
  assign \new_[32181]_  = \new_[32180]_  & \new_[32173]_ ;
  assign \new_[32184]_  = A235 & A234;
  assign \new_[32187]_  = A266 & A265;
  assign \new_[32188]_  = \new_[32187]_  & \new_[32184]_ ;
  assign \new_[32191]_  = A299 & ~A298;
  assign \new_[32194]_  = ~A302 & A300;
  assign \new_[32195]_  = \new_[32194]_  & \new_[32191]_ ;
  assign \new_[32196]_  = \new_[32195]_  & \new_[32188]_ ;
  assign \new_[32200]_  = ~A201 & ~A200;
  assign \new_[32201]_  = A199 & \new_[32200]_ ;
  assign \new_[32204]_  = A203 & ~A202;
  assign \new_[32207]_  = ~A233 & A232;
  assign \new_[32208]_  = \new_[32207]_  & \new_[32204]_ ;
  assign \new_[32209]_  = \new_[32208]_  & \new_[32201]_ ;
  assign \new_[32212]_  = A235 & A234;
  assign \new_[32215]_  = ~A266 & ~A265;
  assign \new_[32216]_  = \new_[32215]_  & \new_[32212]_ ;
  assign \new_[32219]_  = ~A299 & A298;
  assign \new_[32222]_  = A301 & A300;
  assign \new_[32223]_  = \new_[32222]_  & \new_[32219]_ ;
  assign \new_[32224]_  = \new_[32223]_  & \new_[32216]_ ;
  assign \new_[32228]_  = ~A201 & ~A200;
  assign \new_[32229]_  = A199 & \new_[32228]_ ;
  assign \new_[32232]_  = A203 & ~A202;
  assign \new_[32235]_  = ~A233 & A232;
  assign \new_[32236]_  = \new_[32235]_  & \new_[32232]_ ;
  assign \new_[32237]_  = \new_[32236]_  & \new_[32229]_ ;
  assign \new_[32240]_  = A235 & A234;
  assign \new_[32243]_  = ~A266 & ~A265;
  assign \new_[32244]_  = \new_[32243]_  & \new_[32240]_ ;
  assign \new_[32247]_  = ~A299 & A298;
  assign \new_[32250]_  = ~A302 & A300;
  assign \new_[32251]_  = \new_[32250]_  & \new_[32247]_ ;
  assign \new_[32252]_  = \new_[32251]_  & \new_[32244]_ ;
  assign \new_[32256]_  = ~A201 & ~A200;
  assign \new_[32257]_  = A199 & \new_[32256]_ ;
  assign \new_[32260]_  = A203 & ~A202;
  assign \new_[32263]_  = ~A233 & A232;
  assign \new_[32264]_  = \new_[32263]_  & \new_[32260]_ ;
  assign \new_[32265]_  = \new_[32264]_  & \new_[32257]_ ;
  assign \new_[32268]_  = A235 & A234;
  assign \new_[32271]_  = ~A266 & ~A265;
  assign \new_[32272]_  = \new_[32271]_  & \new_[32268]_ ;
  assign \new_[32275]_  = A299 & ~A298;
  assign \new_[32278]_  = A301 & A300;
  assign \new_[32279]_  = \new_[32278]_  & \new_[32275]_ ;
  assign \new_[32280]_  = \new_[32279]_  & \new_[32272]_ ;
  assign \new_[32284]_  = ~A201 & ~A200;
  assign \new_[32285]_  = A199 & \new_[32284]_ ;
  assign \new_[32288]_  = A203 & ~A202;
  assign \new_[32291]_  = ~A233 & A232;
  assign \new_[32292]_  = \new_[32291]_  & \new_[32288]_ ;
  assign \new_[32293]_  = \new_[32292]_  & \new_[32285]_ ;
  assign \new_[32296]_  = A235 & A234;
  assign \new_[32299]_  = ~A266 & ~A265;
  assign \new_[32300]_  = \new_[32299]_  & \new_[32296]_ ;
  assign \new_[32303]_  = A299 & ~A298;
  assign \new_[32306]_  = ~A302 & A300;
  assign \new_[32307]_  = \new_[32306]_  & \new_[32303]_ ;
  assign \new_[32308]_  = \new_[32307]_  & \new_[32300]_ ;
  assign \new_[32312]_  = ~A201 & ~A200;
  assign \new_[32313]_  = A199 & \new_[32312]_ ;
  assign \new_[32316]_  = A203 & ~A202;
  assign \new_[32319]_  = ~A233 & A232;
  assign \new_[32320]_  = \new_[32319]_  & \new_[32316]_ ;
  assign \new_[32321]_  = \new_[32320]_  & \new_[32313]_ ;
  assign \new_[32324]_  = ~A236 & A234;
  assign \new_[32327]_  = A268 & ~A267;
  assign \new_[32328]_  = \new_[32327]_  & \new_[32324]_ ;
  assign \new_[32331]_  = ~A299 & A298;
  assign \new_[32334]_  = A301 & A300;
  assign \new_[32335]_  = \new_[32334]_  & \new_[32331]_ ;
  assign \new_[32336]_  = \new_[32335]_  & \new_[32328]_ ;
  assign \new_[32340]_  = ~A201 & ~A200;
  assign \new_[32341]_  = A199 & \new_[32340]_ ;
  assign \new_[32344]_  = A203 & ~A202;
  assign \new_[32347]_  = ~A233 & A232;
  assign \new_[32348]_  = \new_[32347]_  & \new_[32344]_ ;
  assign \new_[32349]_  = \new_[32348]_  & \new_[32341]_ ;
  assign \new_[32352]_  = ~A236 & A234;
  assign \new_[32355]_  = A268 & ~A267;
  assign \new_[32356]_  = \new_[32355]_  & \new_[32352]_ ;
  assign \new_[32359]_  = ~A299 & A298;
  assign \new_[32362]_  = ~A302 & A300;
  assign \new_[32363]_  = \new_[32362]_  & \new_[32359]_ ;
  assign \new_[32364]_  = \new_[32363]_  & \new_[32356]_ ;
  assign \new_[32368]_  = ~A201 & ~A200;
  assign \new_[32369]_  = A199 & \new_[32368]_ ;
  assign \new_[32372]_  = A203 & ~A202;
  assign \new_[32375]_  = ~A233 & A232;
  assign \new_[32376]_  = \new_[32375]_  & \new_[32372]_ ;
  assign \new_[32377]_  = \new_[32376]_  & \new_[32369]_ ;
  assign \new_[32380]_  = ~A236 & A234;
  assign \new_[32383]_  = A268 & ~A267;
  assign \new_[32384]_  = \new_[32383]_  & \new_[32380]_ ;
  assign \new_[32387]_  = A299 & ~A298;
  assign \new_[32390]_  = A301 & A300;
  assign \new_[32391]_  = \new_[32390]_  & \new_[32387]_ ;
  assign \new_[32392]_  = \new_[32391]_  & \new_[32384]_ ;
  assign \new_[32396]_  = ~A201 & ~A200;
  assign \new_[32397]_  = A199 & \new_[32396]_ ;
  assign \new_[32400]_  = A203 & ~A202;
  assign \new_[32403]_  = ~A233 & A232;
  assign \new_[32404]_  = \new_[32403]_  & \new_[32400]_ ;
  assign \new_[32405]_  = \new_[32404]_  & \new_[32397]_ ;
  assign \new_[32408]_  = ~A236 & A234;
  assign \new_[32411]_  = A268 & ~A267;
  assign \new_[32412]_  = \new_[32411]_  & \new_[32408]_ ;
  assign \new_[32415]_  = A299 & ~A298;
  assign \new_[32418]_  = ~A302 & A300;
  assign \new_[32419]_  = \new_[32418]_  & \new_[32415]_ ;
  assign \new_[32420]_  = \new_[32419]_  & \new_[32412]_ ;
  assign \new_[32424]_  = ~A201 & ~A200;
  assign \new_[32425]_  = A199 & \new_[32424]_ ;
  assign \new_[32428]_  = A203 & ~A202;
  assign \new_[32431]_  = ~A233 & A232;
  assign \new_[32432]_  = \new_[32431]_  & \new_[32428]_ ;
  assign \new_[32433]_  = \new_[32432]_  & \new_[32425]_ ;
  assign \new_[32436]_  = ~A236 & A234;
  assign \new_[32439]_  = ~A269 & ~A267;
  assign \new_[32440]_  = \new_[32439]_  & \new_[32436]_ ;
  assign \new_[32443]_  = ~A299 & A298;
  assign \new_[32446]_  = A301 & A300;
  assign \new_[32447]_  = \new_[32446]_  & \new_[32443]_ ;
  assign \new_[32448]_  = \new_[32447]_  & \new_[32440]_ ;
  assign \new_[32452]_  = ~A201 & ~A200;
  assign \new_[32453]_  = A199 & \new_[32452]_ ;
  assign \new_[32456]_  = A203 & ~A202;
  assign \new_[32459]_  = ~A233 & A232;
  assign \new_[32460]_  = \new_[32459]_  & \new_[32456]_ ;
  assign \new_[32461]_  = \new_[32460]_  & \new_[32453]_ ;
  assign \new_[32464]_  = ~A236 & A234;
  assign \new_[32467]_  = ~A269 & ~A267;
  assign \new_[32468]_  = \new_[32467]_  & \new_[32464]_ ;
  assign \new_[32471]_  = ~A299 & A298;
  assign \new_[32474]_  = ~A302 & A300;
  assign \new_[32475]_  = \new_[32474]_  & \new_[32471]_ ;
  assign \new_[32476]_  = \new_[32475]_  & \new_[32468]_ ;
  assign \new_[32480]_  = ~A201 & ~A200;
  assign \new_[32481]_  = A199 & \new_[32480]_ ;
  assign \new_[32484]_  = A203 & ~A202;
  assign \new_[32487]_  = ~A233 & A232;
  assign \new_[32488]_  = \new_[32487]_  & \new_[32484]_ ;
  assign \new_[32489]_  = \new_[32488]_  & \new_[32481]_ ;
  assign \new_[32492]_  = ~A236 & A234;
  assign \new_[32495]_  = ~A269 & ~A267;
  assign \new_[32496]_  = \new_[32495]_  & \new_[32492]_ ;
  assign \new_[32499]_  = A299 & ~A298;
  assign \new_[32502]_  = A301 & A300;
  assign \new_[32503]_  = \new_[32502]_  & \new_[32499]_ ;
  assign \new_[32504]_  = \new_[32503]_  & \new_[32496]_ ;
  assign \new_[32508]_  = ~A201 & ~A200;
  assign \new_[32509]_  = A199 & \new_[32508]_ ;
  assign \new_[32512]_  = A203 & ~A202;
  assign \new_[32515]_  = ~A233 & A232;
  assign \new_[32516]_  = \new_[32515]_  & \new_[32512]_ ;
  assign \new_[32517]_  = \new_[32516]_  & \new_[32509]_ ;
  assign \new_[32520]_  = ~A236 & A234;
  assign \new_[32523]_  = ~A269 & ~A267;
  assign \new_[32524]_  = \new_[32523]_  & \new_[32520]_ ;
  assign \new_[32527]_  = A299 & ~A298;
  assign \new_[32530]_  = ~A302 & A300;
  assign \new_[32531]_  = \new_[32530]_  & \new_[32527]_ ;
  assign \new_[32532]_  = \new_[32531]_  & \new_[32524]_ ;
  assign \new_[32536]_  = ~A201 & ~A200;
  assign \new_[32537]_  = A199 & \new_[32536]_ ;
  assign \new_[32540]_  = A203 & ~A202;
  assign \new_[32543]_  = ~A233 & A232;
  assign \new_[32544]_  = \new_[32543]_  & \new_[32540]_ ;
  assign \new_[32545]_  = \new_[32544]_  & \new_[32537]_ ;
  assign \new_[32548]_  = ~A236 & A234;
  assign \new_[32551]_  = A266 & A265;
  assign \new_[32552]_  = \new_[32551]_  & \new_[32548]_ ;
  assign \new_[32555]_  = ~A299 & A298;
  assign \new_[32558]_  = A301 & A300;
  assign \new_[32559]_  = \new_[32558]_  & \new_[32555]_ ;
  assign \new_[32560]_  = \new_[32559]_  & \new_[32552]_ ;
  assign \new_[32564]_  = ~A201 & ~A200;
  assign \new_[32565]_  = A199 & \new_[32564]_ ;
  assign \new_[32568]_  = A203 & ~A202;
  assign \new_[32571]_  = ~A233 & A232;
  assign \new_[32572]_  = \new_[32571]_  & \new_[32568]_ ;
  assign \new_[32573]_  = \new_[32572]_  & \new_[32565]_ ;
  assign \new_[32576]_  = ~A236 & A234;
  assign \new_[32579]_  = A266 & A265;
  assign \new_[32580]_  = \new_[32579]_  & \new_[32576]_ ;
  assign \new_[32583]_  = ~A299 & A298;
  assign \new_[32586]_  = ~A302 & A300;
  assign \new_[32587]_  = \new_[32586]_  & \new_[32583]_ ;
  assign \new_[32588]_  = \new_[32587]_  & \new_[32580]_ ;
  assign \new_[32592]_  = ~A201 & ~A200;
  assign \new_[32593]_  = A199 & \new_[32592]_ ;
  assign \new_[32596]_  = A203 & ~A202;
  assign \new_[32599]_  = ~A233 & A232;
  assign \new_[32600]_  = \new_[32599]_  & \new_[32596]_ ;
  assign \new_[32601]_  = \new_[32600]_  & \new_[32593]_ ;
  assign \new_[32604]_  = ~A236 & A234;
  assign \new_[32607]_  = A266 & A265;
  assign \new_[32608]_  = \new_[32607]_  & \new_[32604]_ ;
  assign \new_[32611]_  = A299 & ~A298;
  assign \new_[32614]_  = A301 & A300;
  assign \new_[32615]_  = \new_[32614]_  & \new_[32611]_ ;
  assign \new_[32616]_  = \new_[32615]_  & \new_[32608]_ ;
  assign \new_[32620]_  = ~A201 & ~A200;
  assign \new_[32621]_  = A199 & \new_[32620]_ ;
  assign \new_[32624]_  = A203 & ~A202;
  assign \new_[32627]_  = ~A233 & A232;
  assign \new_[32628]_  = \new_[32627]_  & \new_[32624]_ ;
  assign \new_[32629]_  = \new_[32628]_  & \new_[32621]_ ;
  assign \new_[32632]_  = ~A236 & A234;
  assign \new_[32635]_  = A266 & A265;
  assign \new_[32636]_  = \new_[32635]_  & \new_[32632]_ ;
  assign \new_[32639]_  = A299 & ~A298;
  assign \new_[32642]_  = ~A302 & A300;
  assign \new_[32643]_  = \new_[32642]_  & \new_[32639]_ ;
  assign \new_[32644]_  = \new_[32643]_  & \new_[32636]_ ;
  assign \new_[32648]_  = ~A201 & ~A200;
  assign \new_[32649]_  = A199 & \new_[32648]_ ;
  assign \new_[32652]_  = A203 & ~A202;
  assign \new_[32655]_  = ~A233 & A232;
  assign \new_[32656]_  = \new_[32655]_  & \new_[32652]_ ;
  assign \new_[32657]_  = \new_[32656]_  & \new_[32649]_ ;
  assign \new_[32660]_  = ~A236 & A234;
  assign \new_[32663]_  = ~A266 & ~A265;
  assign \new_[32664]_  = \new_[32663]_  & \new_[32660]_ ;
  assign \new_[32667]_  = ~A299 & A298;
  assign \new_[32670]_  = A301 & A300;
  assign \new_[32671]_  = \new_[32670]_  & \new_[32667]_ ;
  assign \new_[32672]_  = \new_[32671]_  & \new_[32664]_ ;
  assign \new_[32676]_  = ~A201 & ~A200;
  assign \new_[32677]_  = A199 & \new_[32676]_ ;
  assign \new_[32680]_  = A203 & ~A202;
  assign \new_[32683]_  = ~A233 & A232;
  assign \new_[32684]_  = \new_[32683]_  & \new_[32680]_ ;
  assign \new_[32685]_  = \new_[32684]_  & \new_[32677]_ ;
  assign \new_[32688]_  = ~A236 & A234;
  assign \new_[32691]_  = ~A266 & ~A265;
  assign \new_[32692]_  = \new_[32691]_  & \new_[32688]_ ;
  assign \new_[32695]_  = ~A299 & A298;
  assign \new_[32698]_  = ~A302 & A300;
  assign \new_[32699]_  = \new_[32698]_  & \new_[32695]_ ;
  assign \new_[32700]_  = \new_[32699]_  & \new_[32692]_ ;
  assign \new_[32704]_  = ~A201 & ~A200;
  assign \new_[32705]_  = A199 & \new_[32704]_ ;
  assign \new_[32708]_  = A203 & ~A202;
  assign \new_[32711]_  = ~A233 & A232;
  assign \new_[32712]_  = \new_[32711]_  & \new_[32708]_ ;
  assign \new_[32713]_  = \new_[32712]_  & \new_[32705]_ ;
  assign \new_[32716]_  = ~A236 & A234;
  assign \new_[32719]_  = ~A266 & ~A265;
  assign \new_[32720]_  = \new_[32719]_  & \new_[32716]_ ;
  assign \new_[32723]_  = A299 & ~A298;
  assign \new_[32726]_  = A301 & A300;
  assign \new_[32727]_  = \new_[32726]_  & \new_[32723]_ ;
  assign \new_[32728]_  = \new_[32727]_  & \new_[32720]_ ;
  assign \new_[32732]_  = ~A201 & ~A200;
  assign \new_[32733]_  = A199 & \new_[32732]_ ;
  assign \new_[32736]_  = A203 & ~A202;
  assign \new_[32739]_  = ~A233 & A232;
  assign \new_[32740]_  = \new_[32739]_  & \new_[32736]_ ;
  assign \new_[32741]_  = \new_[32740]_  & \new_[32733]_ ;
  assign \new_[32744]_  = ~A236 & A234;
  assign \new_[32747]_  = ~A266 & ~A265;
  assign \new_[32748]_  = \new_[32747]_  & \new_[32744]_ ;
  assign \new_[32751]_  = A299 & ~A298;
  assign \new_[32754]_  = ~A302 & A300;
  assign \new_[32755]_  = \new_[32754]_  & \new_[32751]_ ;
  assign \new_[32756]_  = \new_[32755]_  & \new_[32748]_ ;
  assign \new_[32760]_  = A167 & A168;
  assign \new_[32761]_  = A170 & \new_[32760]_ ;
  assign \new_[32764]_  = ~A232 & ~A166;
  assign \new_[32767]_  = A234 & A233;
  assign \new_[32768]_  = \new_[32767]_  & \new_[32764]_ ;
  assign \new_[32769]_  = \new_[32768]_  & \new_[32761]_ ;
  assign \new_[32772]_  = A267 & A235;
  assign \new_[32775]_  = A269 & ~A268;
  assign \new_[32776]_  = \new_[32775]_  & \new_[32772]_ ;
  assign \new_[32779]_  = ~A299 & A298;
  assign \new_[32782]_  = A301 & A300;
  assign \new_[32783]_  = \new_[32782]_  & \new_[32779]_ ;
  assign \new_[32784]_  = \new_[32783]_  & \new_[32776]_ ;
  assign \new_[32788]_  = A167 & A168;
  assign \new_[32789]_  = A170 & \new_[32788]_ ;
  assign \new_[32792]_  = ~A232 & ~A166;
  assign \new_[32795]_  = A234 & A233;
  assign \new_[32796]_  = \new_[32795]_  & \new_[32792]_ ;
  assign \new_[32797]_  = \new_[32796]_  & \new_[32789]_ ;
  assign \new_[32800]_  = A267 & A235;
  assign \new_[32803]_  = A269 & ~A268;
  assign \new_[32804]_  = \new_[32803]_  & \new_[32800]_ ;
  assign \new_[32807]_  = ~A299 & A298;
  assign \new_[32810]_  = ~A302 & A300;
  assign \new_[32811]_  = \new_[32810]_  & \new_[32807]_ ;
  assign \new_[32812]_  = \new_[32811]_  & \new_[32804]_ ;
  assign \new_[32816]_  = A167 & A168;
  assign \new_[32817]_  = A170 & \new_[32816]_ ;
  assign \new_[32820]_  = ~A232 & ~A166;
  assign \new_[32823]_  = A234 & A233;
  assign \new_[32824]_  = \new_[32823]_  & \new_[32820]_ ;
  assign \new_[32825]_  = \new_[32824]_  & \new_[32817]_ ;
  assign \new_[32828]_  = A267 & A235;
  assign \new_[32831]_  = A269 & ~A268;
  assign \new_[32832]_  = \new_[32831]_  & \new_[32828]_ ;
  assign \new_[32835]_  = A299 & ~A298;
  assign \new_[32838]_  = A301 & A300;
  assign \new_[32839]_  = \new_[32838]_  & \new_[32835]_ ;
  assign \new_[32840]_  = \new_[32839]_  & \new_[32832]_ ;
  assign \new_[32844]_  = A167 & A168;
  assign \new_[32845]_  = A170 & \new_[32844]_ ;
  assign \new_[32848]_  = ~A232 & ~A166;
  assign \new_[32851]_  = A234 & A233;
  assign \new_[32852]_  = \new_[32851]_  & \new_[32848]_ ;
  assign \new_[32853]_  = \new_[32852]_  & \new_[32845]_ ;
  assign \new_[32856]_  = A267 & A235;
  assign \new_[32859]_  = A269 & ~A268;
  assign \new_[32860]_  = \new_[32859]_  & \new_[32856]_ ;
  assign \new_[32863]_  = A299 & ~A298;
  assign \new_[32866]_  = ~A302 & A300;
  assign \new_[32867]_  = \new_[32866]_  & \new_[32863]_ ;
  assign \new_[32868]_  = \new_[32867]_  & \new_[32860]_ ;
  assign \new_[32872]_  = A167 & A168;
  assign \new_[32873]_  = A170 & \new_[32872]_ ;
  assign \new_[32876]_  = ~A232 & ~A166;
  assign \new_[32879]_  = A234 & A233;
  assign \new_[32880]_  = \new_[32879]_  & \new_[32876]_ ;
  assign \new_[32881]_  = \new_[32880]_  & \new_[32873]_ ;
  assign \new_[32884]_  = ~A267 & A235;
  assign \new_[32887]_  = A298 & A268;
  assign \new_[32888]_  = \new_[32887]_  & \new_[32884]_ ;
  assign \new_[32891]_  = ~A300 & ~A299;
  assign \new_[32894]_  = A302 & ~A301;
  assign \new_[32895]_  = \new_[32894]_  & \new_[32891]_ ;
  assign \new_[32896]_  = \new_[32895]_  & \new_[32888]_ ;
  assign \new_[32900]_  = A167 & A168;
  assign \new_[32901]_  = A170 & \new_[32900]_ ;
  assign \new_[32904]_  = ~A232 & ~A166;
  assign \new_[32907]_  = A234 & A233;
  assign \new_[32908]_  = \new_[32907]_  & \new_[32904]_ ;
  assign \new_[32909]_  = \new_[32908]_  & \new_[32901]_ ;
  assign \new_[32912]_  = ~A267 & A235;
  assign \new_[32915]_  = ~A298 & A268;
  assign \new_[32916]_  = \new_[32915]_  & \new_[32912]_ ;
  assign \new_[32919]_  = ~A300 & A299;
  assign \new_[32922]_  = A302 & ~A301;
  assign \new_[32923]_  = \new_[32922]_  & \new_[32919]_ ;
  assign \new_[32924]_  = \new_[32923]_  & \new_[32916]_ ;
  assign \new_[32928]_  = A167 & A168;
  assign \new_[32929]_  = A170 & \new_[32928]_ ;
  assign \new_[32932]_  = ~A232 & ~A166;
  assign \new_[32935]_  = A234 & A233;
  assign \new_[32936]_  = \new_[32935]_  & \new_[32932]_ ;
  assign \new_[32937]_  = \new_[32936]_  & \new_[32929]_ ;
  assign \new_[32940]_  = ~A267 & A235;
  assign \new_[32943]_  = A298 & ~A269;
  assign \new_[32944]_  = \new_[32943]_  & \new_[32940]_ ;
  assign \new_[32947]_  = ~A300 & ~A299;
  assign \new_[32950]_  = A302 & ~A301;
  assign \new_[32951]_  = \new_[32950]_  & \new_[32947]_ ;
  assign \new_[32952]_  = \new_[32951]_  & \new_[32944]_ ;
  assign \new_[32956]_  = A167 & A168;
  assign \new_[32957]_  = A170 & \new_[32956]_ ;
  assign \new_[32960]_  = ~A232 & ~A166;
  assign \new_[32963]_  = A234 & A233;
  assign \new_[32964]_  = \new_[32963]_  & \new_[32960]_ ;
  assign \new_[32965]_  = \new_[32964]_  & \new_[32957]_ ;
  assign \new_[32968]_  = ~A267 & A235;
  assign \new_[32971]_  = ~A298 & ~A269;
  assign \new_[32972]_  = \new_[32971]_  & \new_[32968]_ ;
  assign \new_[32975]_  = ~A300 & A299;
  assign \new_[32978]_  = A302 & ~A301;
  assign \new_[32979]_  = \new_[32978]_  & \new_[32975]_ ;
  assign \new_[32980]_  = \new_[32979]_  & \new_[32972]_ ;
  assign \new_[32984]_  = A167 & A168;
  assign \new_[32985]_  = A170 & \new_[32984]_ ;
  assign \new_[32988]_  = ~A232 & ~A166;
  assign \new_[32991]_  = A234 & A233;
  assign \new_[32992]_  = \new_[32991]_  & \new_[32988]_ ;
  assign \new_[32993]_  = \new_[32992]_  & \new_[32985]_ ;
  assign \new_[32996]_  = A265 & A235;
  assign \new_[32999]_  = A298 & A266;
  assign \new_[33000]_  = \new_[32999]_  & \new_[32996]_ ;
  assign \new_[33003]_  = ~A300 & ~A299;
  assign \new_[33006]_  = A302 & ~A301;
  assign \new_[33007]_  = \new_[33006]_  & \new_[33003]_ ;
  assign \new_[33008]_  = \new_[33007]_  & \new_[33000]_ ;
  assign \new_[33012]_  = A167 & A168;
  assign \new_[33013]_  = A170 & \new_[33012]_ ;
  assign \new_[33016]_  = ~A232 & ~A166;
  assign \new_[33019]_  = A234 & A233;
  assign \new_[33020]_  = \new_[33019]_  & \new_[33016]_ ;
  assign \new_[33021]_  = \new_[33020]_  & \new_[33013]_ ;
  assign \new_[33024]_  = A265 & A235;
  assign \new_[33027]_  = ~A298 & A266;
  assign \new_[33028]_  = \new_[33027]_  & \new_[33024]_ ;
  assign \new_[33031]_  = ~A300 & A299;
  assign \new_[33034]_  = A302 & ~A301;
  assign \new_[33035]_  = \new_[33034]_  & \new_[33031]_ ;
  assign \new_[33036]_  = \new_[33035]_  & \new_[33028]_ ;
  assign \new_[33040]_  = A167 & A168;
  assign \new_[33041]_  = A170 & \new_[33040]_ ;
  assign \new_[33044]_  = ~A232 & ~A166;
  assign \new_[33047]_  = A234 & A233;
  assign \new_[33048]_  = \new_[33047]_  & \new_[33044]_ ;
  assign \new_[33049]_  = \new_[33048]_  & \new_[33041]_ ;
  assign \new_[33052]_  = ~A265 & A235;
  assign \new_[33055]_  = A298 & ~A266;
  assign \new_[33056]_  = \new_[33055]_  & \new_[33052]_ ;
  assign \new_[33059]_  = ~A300 & ~A299;
  assign \new_[33062]_  = A302 & ~A301;
  assign \new_[33063]_  = \new_[33062]_  & \new_[33059]_ ;
  assign \new_[33064]_  = \new_[33063]_  & \new_[33056]_ ;
  assign \new_[33068]_  = A167 & A168;
  assign \new_[33069]_  = A170 & \new_[33068]_ ;
  assign \new_[33072]_  = ~A232 & ~A166;
  assign \new_[33075]_  = A234 & A233;
  assign \new_[33076]_  = \new_[33075]_  & \new_[33072]_ ;
  assign \new_[33077]_  = \new_[33076]_  & \new_[33069]_ ;
  assign \new_[33080]_  = ~A265 & A235;
  assign \new_[33083]_  = ~A298 & ~A266;
  assign \new_[33084]_  = \new_[33083]_  & \new_[33080]_ ;
  assign \new_[33087]_  = ~A300 & A299;
  assign \new_[33090]_  = A302 & ~A301;
  assign \new_[33091]_  = \new_[33090]_  & \new_[33087]_ ;
  assign \new_[33092]_  = \new_[33091]_  & \new_[33084]_ ;
  assign \new_[33096]_  = A167 & A168;
  assign \new_[33097]_  = A170 & \new_[33096]_ ;
  assign \new_[33100]_  = ~A232 & ~A166;
  assign \new_[33103]_  = A234 & A233;
  assign \new_[33104]_  = \new_[33103]_  & \new_[33100]_ ;
  assign \new_[33105]_  = \new_[33104]_  & \new_[33097]_ ;
  assign \new_[33108]_  = A267 & ~A236;
  assign \new_[33111]_  = A269 & ~A268;
  assign \new_[33112]_  = \new_[33111]_  & \new_[33108]_ ;
  assign \new_[33115]_  = ~A299 & A298;
  assign \new_[33118]_  = A301 & A300;
  assign \new_[33119]_  = \new_[33118]_  & \new_[33115]_ ;
  assign \new_[33120]_  = \new_[33119]_  & \new_[33112]_ ;
  assign \new_[33124]_  = A167 & A168;
  assign \new_[33125]_  = A170 & \new_[33124]_ ;
  assign \new_[33128]_  = ~A232 & ~A166;
  assign \new_[33131]_  = A234 & A233;
  assign \new_[33132]_  = \new_[33131]_  & \new_[33128]_ ;
  assign \new_[33133]_  = \new_[33132]_  & \new_[33125]_ ;
  assign \new_[33136]_  = A267 & ~A236;
  assign \new_[33139]_  = A269 & ~A268;
  assign \new_[33140]_  = \new_[33139]_  & \new_[33136]_ ;
  assign \new_[33143]_  = ~A299 & A298;
  assign \new_[33146]_  = ~A302 & A300;
  assign \new_[33147]_  = \new_[33146]_  & \new_[33143]_ ;
  assign \new_[33148]_  = \new_[33147]_  & \new_[33140]_ ;
  assign \new_[33152]_  = A167 & A168;
  assign \new_[33153]_  = A170 & \new_[33152]_ ;
  assign \new_[33156]_  = ~A232 & ~A166;
  assign \new_[33159]_  = A234 & A233;
  assign \new_[33160]_  = \new_[33159]_  & \new_[33156]_ ;
  assign \new_[33161]_  = \new_[33160]_  & \new_[33153]_ ;
  assign \new_[33164]_  = A267 & ~A236;
  assign \new_[33167]_  = A269 & ~A268;
  assign \new_[33168]_  = \new_[33167]_  & \new_[33164]_ ;
  assign \new_[33171]_  = A299 & ~A298;
  assign \new_[33174]_  = A301 & A300;
  assign \new_[33175]_  = \new_[33174]_  & \new_[33171]_ ;
  assign \new_[33176]_  = \new_[33175]_  & \new_[33168]_ ;
  assign \new_[33180]_  = A167 & A168;
  assign \new_[33181]_  = A170 & \new_[33180]_ ;
  assign \new_[33184]_  = ~A232 & ~A166;
  assign \new_[33187]_  = A234 & A233;
  assign \new_[33188]_  = \new_[33187]_  & \new_[33184]_ ;
  assign \new_[33189]_  = \new_[33188]_  & \new_[33181]_ ;
  assign \new_[33192]_  = A267 & ~A236;
  assign \new_[33195]_  = A269 & ~A268;
  assign \new_[33196]_  = \new_[33195]_  & \new_[33192]_ ;
  assign \new_[33199]_  = A299 & ~A298;
  assign \new_[33202]_  = ~A302 & A300;
  assign \new_[33203]_  = \new_[33202]_  & \new_[33199]_ ;
  assign \new_[33204]_  = \new_[33203]_  & \new_[33196]_ ;
  assign \new_[33208]_  = A167 & A168;
  assign \new_[33209]_  = A170 & \new_[33208]_ ;
  assign \new_[33212]_  = ~A232 & ~A166;
  assign \new_[33215]_  = A234 & A233;
  assign \new_[33216]_  = \new_[33215]_  & \new_[33212]_ ;
  assign \new_[33217]_  = \new_[33216]_  & \new_[33209]_ ;
  assign \new_[33220]_  = ~A267 & ~A236;
  assign \new_[33223]_  = A298 & A268;
  assign \new_[33224]_  = \new_[33223]_  & \new_[33220]_ ;
  assign \new_[33227]_  = ~A300 & ~A299;
  assign \new_[33230]_  = A302 & ~A301;
  assign \new_[33231]_  = \new_[33230]_  & \new_[33227]_ ;
  assign \new_[33232]_  = \new_[33231]_  & \new_[33224]_ ;
  assign \new_[33236]_  = A167 & A168;
  assign \new_[33237]_  = A170 & \new_[33236]_ ;
  assign \new_[33240]_  = ~A232 & ~A166;
  assign \new_[33243]_  = A234 & A233;
  assign \new_[33244]_  = \new_[33243]_  & \new_[33240]_ ;
  assign \new_[33245]_  = \new_[33244]_  & \new_[33237]_ ;
  assign \new_[33248]_  = ~A267 & ~A236;
  assign \new_[33251]_  = ~A298 & A268;
  assign \new_[33252]_  = \new_[33251]_  & \new_[33248]_ ;
  assign \new_[33255]_  = ~A300 & A299;
  assign \new_[33258]_  = A302 & ~A301;
  assign \new_[33259]_  = \new_[33258]_  & \new_[33255]_ ;
  assign \new_[33260]_  = \new_[33259]_  & \new_[33252]_ ;
  assign \new_[33264]_  = A167 & A168;
  assign \new_[33265]_  = A170 & \new_[33264]_ ;
  assign \new_[33268]_  = ~A232 & ~A166;
  assign \new_[33271]_  = A234 & A233;
  assign \new_[33272]_  = \new_[33271]_  & \new_[33268]_ ;
  assign \new_[33273]_  = \new_[33272]_  & \new_[33265]_ ;
  assign \new_[33276]_  = ~A267 & ~A236;
  assign \new_[33279]_  = A298 & ~A269;
  assign \new_[33280]_  = \new_[33279]_  & \new_[33276]_ ;
  assign \new_[33283]_  = ~A300 & ~A299;
  assign \new_[33286]_  = A302 & ~A301;
  assign \new_[33287]_  = \new_[33286]_  & \new_[33283]_ ;
  assign \new_[33288]_  = \new_[33287]_  & \new_[33280]_ ;
  assign \new_[33292]_  = A167 & A168;
  assign \new_[33293]_  = A170 & \new_[33292]_ ;
  assign \new_[33296]_  = ~A232 & ~A166;
  assign \new_[33299]_  = A234 & A233;
  assign \new_[33300]_  = \new_[33299]_  & \new_[33296]_ ;
  assign \new_[33301]_  = \new_[33300]_  & \new_[33293]_ ;
  assign \new_[33304]_  = ~A267 & ~A236;
  assign \new_[33307]_  = ~A298 & ~A269;
  assign \new_[33308]_  = \new_[33307]_  & \new_[33304]_ ;
  assign \new_[33311]_  = ~A300 & A299;
  assign \new_[33314]_  = A302 & ~A301;
  assign \new_[33315]_  = \new_[33314]_  & \new_[33311]_ ;
  assign \new_[33316]_  = \new_[33315]_  & \new_[33308]_ ;
  assign \new_[33320]_  = A167 & A168;
  assign \new_[33321]_  = A170 & \new_[33320]_ ;
  assign \new_[33324]_  = ~A232 & ~A166;
  assign \new_[33327]_  = A234 & A233;
  assign \new_[33328]_  = \new_[33327]_  & \new_[33324]_ ;
  assign \new_[33329]_  = \new_[33328]_  & \new_[33321]_ ;
  assign \new_[33332]_  = A265 & ~A236;
  assign \new_[33335]_  = A298 & A266;
  assign \new_[33336]_  = \new_[33335]_  & \new_[33332]_ ;
  assign \new_[33339]_  = ~A300 & ~A299;
  assign \new_[33342]_  = A302 & ~A301;
  assign \new_[33343]_  = \new_[33342]_  & \new_[33339]_ ;
  assign \new_[33344]_  = \new_[33343]_  & \new_[33336]_ ;
  assign \new_[33348]_  = A167 & A168;
  assign \new_[33349]_  = A170 & \new_[33348]_ ;
  assign \new_[33352]_  = ~A232 & ~A166;
  assign \new_[33355]_  = A234 & A233;
  assign \new_[33356]_  = \new_[33355]_  & \new_[33352]_ ;
  assign \new_[33357]_  = \new_[33356]_  & \new_[33349]_ ;
  assign \new_[33360]_  = A265 & ~A236;
  assign \new_[33363]_  = ~A298 & A266;
  assign \new_[33364]_  = \new_[33363]_  & \new_[33360]_ ;
  assign \new_[33367]_  = ~A300 & A299;
  assign \new_[33370]_  = A302 & ~A301;
  assign \new_[33371]_  = \new_[33370]_  & \new_[33367]_ ;
  assign \new_[33372]_  = \new_[33371]_  & \new_[33364]_ ;
  assign \new_[33376]_  = A167 & A168;
  assign \new_[33377]_  = A170 & \new_[33376]_ ;
  assign \new_[33380]_  = ~A232 & ~A166;
  assign \new_[33383]_  = A234 & A233;
  assign \new_[33384]_  = \new_[33383]_  & \new_[33380]_ ;
  assign \new_[33385]_  = \new_[33384]_  & \new_[33377]_ ;
  assign \new_[33388]_  = ~A265 & ~A236;
  assign \new_[33391]_  = A298 & ~A266;
  assign \new_[33392]_  = \new_[33391]_  & \new_[33388]_ ;
  assign \new_[33395]_  = ~A300 & ~A299;
  assign \new_[33398]_  = A302 & ~A301;
  assign \new_[33399]_  = \new_[33398]_  & \new_[33395]_ ;
  assign \new_[33400]_  = \new_[33399]_  & \new_[33392]_ ;
  assign \new_[33404]_  = A167 & A168;
  assign \new_[33405]_  = A170 & \new_[33404]_ ;
  assign \new_[33408]_  = ~A232 & ~A166;
  assign \new_[33411]_  = A234 & A233;
  assign \new_[33412]_  = \new_[33411]_  & \new_[33408]_ ;
  assign \new_[33413]_  = \new_[33412]_  & \new_[33405]_ ;
  assign \new_[33416]_  = ~A265 & ~A236;
  assign \new_[33419]_  = ~A298 & ~A266;
  assign \new_[33420]_  = \new_[33419]_  & \new_[33416]_ ;
  assign \new_[33423]_  = ~A300 & A299;
  assign \new_[33426]_  = A302 & ~A301;
  assign \new_[33427]_  = \new_[33426]_  & \new_[33423]_ ;
  assign \new_[33428]_  = \new_[33427]_  & \new_[33420]_ ;
  assign \new_[33432]_  = A167 & A168;
  assign \new_[33433]_  = A170 & \new_[33432]_ ;
  assign \new_[33436]_  = ~A232 & ~A166;
  assign \new_[33439]_  = ~A234 & A233;
  assign \new_[33440]_  = \new_[33439]_  & \new_[33436]_ ;
  assign \new_[33441]_  = \new_[33440]_  & \new_[33433]_ ;
  assign \new_[33444]_  = A236 & ~A235;
  assign \new_[33447]_  = A268 & ~A267;
  assign \new_[33448]_  = \new_[33447]_  & \new_[33444]_ ;
  assign \new_[33451]_  = ~A299 & A298;
  assign \new_[33454]_  = A301 & A300;
  assign \new_[33455]_  = \new_[33454]_  & \new_[33451]_ ;
  assign \new_[33456]_  = \new_[33455]_  & \new_[33448]_ ;
  assign \new_[33460]_  = A167 & A168;
  assign \new_[33461]_  = A170 & \new_[33460]_ ;
  assign \new_[33464]_  = ~A232 & ~A166;
  assign \new_[33467]_  = ~A234 & A233;
  assign \new_[33468]_  = \new_[33467]_  & \new_[33464]_ ;
  assign \new_[33469]_  = \new_[33468]_  & \new_[33461]_ ;
  assign \new_[33472]_  = A236 & ~A235;
  assign \new_[33475]_  = A268 & ~A267;
  assign \new_[33476]_  = \new_[33475]_  & \new_[33472]_ ;
  assign \new_[33479]_  = ~A299 & A298;
  assign \new_[33482]_  = ~A302 & A300;
  assign \new_[33483]_  = \new_[33482]_  & \new_[33479]_ ;
  assign \new_[33484]_  = \new_[33483]_  & \new_[33476]_ ;
  assign \new_[33488]_  = A167 & A168;
  assign \new_[33489]_  = A170 & \new_[33488]_ ;
  assign \new_[33492]_  = ~A232 & ~A166;
  assign \new_[33495]_  = ~A234 & A233;
  assign \new_[33496]_  = \new_[33495]_  & \new_[33492]_ ;
  assign \new_[33497]_  = \new_[33496]_  & \new_[33489]_ ;
  assign \new_[33500]_  = A236 & ~A235;
  assign \new_[33503]_  = A268 & ~A267;
  assign \new_[33504]_  = \new_[33503]_  & \new_[33500]_ ;
  assign \new_[33507]_  = A299 & ~A298;
  assign \new_[33510]_  = A301 & A300;
  assign \new_[33511]_  = \new_[33510]_  & \new_[33507]_ ;
  assign \new_[33512]_  = \new_[33511]_  & \new_[33504]_ ;
  assign \new_[33516]_  = A167 & A168;
  assign \new_[33517]_  = A170 & \new_[33516]_ ;
  assign \new_[33520]_  = ~A232 & ~A166;
  assign \new_[33523]_  = ~A234 & A233;
  assign \new_[33524]_  = \new_[33523]_  & \new_[33520]_ ;
  assign \new_[33525]_  = \new_[33524]_  & \new_[33517]_ ;
  assign \new_[33528]_  = A236 & ~A235;
  assign \new_[33531]_  = A268 & ~A267;
  assign \new_[33532]_  = \new_[33531]_  & \new_[33528]_ ;
  assign \new_[33535]_  = A299 & ~A298;
  assign \new_[33538]_  = ~A302 & A300;
  assign \new_[33539]_  = \new_[33538]_  & \new_[33535]_ ;
  assign \new_[33540]_  = \new_[33539]_  & \new_[33532]_ ;
  assign \new_[33544]_  = A167 & A168;
  assign \new_[33545]_  = A170 & \new_[33544]_ ;
  assign \new_[33548]_  = ~A232 & ~A166;
  assign \new_[33551]_  = ~A234 & A233;
  assign \new_[33552]_  = \new_[33551]_  & \new_[33548]_ ;
  assign \new_[33553]_  = \new_[33552]_  & \new_[33545]_ ;
  assign \new_[33556]_  = A236 & ~A235;
  assign \new_[33559]_  = ~A269 & ~A267;
  assign \new_[33560]_  = \new_[33559]_  & \new_[33556]_ ;
  assign \new_[33563]_  = ~A299 & A298;
  assign \new_[33566]_  = A301 & A300;
  assign \new_[33567]_  = \new_[33566]_  & \new_[33563]_ ;
  assign \new_[33568]_  = \new_[33567]_  & \new_[33560]_ ;
  assign \new_[33572]_  = A167 & A168;
  assign \new_[33573]_  = A170 & \new_[33572]_ ;
  assign \new_[33576]_  = ~A232 & ~A166;
  assign \new_[33579]_  = ~A234 & A233;
  assign \new_[33580]_  = \new_[33579]_  & \new_[33576]_ ;
  assign \new_[33581]_  = \new_[33580]_  & \new_[33573]_ ;
  assign \new_[33584]_  = A236 & ~A235;
  assign \new_[33587]_  = ~A269 & ~A267;
  assign \new_[33588]_  = \new_[33587]_  & \new_[33584]_ ;
  assign \new_[33591]_  = ~A299 & A298;
  assign \new_[33594]_  = ~A302 & A300;
  assign \new_[33595]_  = \new_[33594]_  & \new_[33591]_ ;
  assign \new_[33596]_  = \new_[33595]_  & \new_[33588]_ ;
  assign \new_[33600]_  = A167 & A168;
  assign \new_[33601]_  = A170 & \new_[33600]_ ;
  assign \new_[33604]_  = ~A232 & ~A166;
  assign \new_[33607]_  = ~A234 & A233;
  assign \new_[33608]_  = \new_[33607]_  & \new_[33604]_ ;
  assign \new_[33609]_  = \new_[33608]_  & \new_[33601]_ ;
  assign \new_[33612]_  = A236 & ~A235;
  assign \new_[33615]_  = ~A269 & ~A267;
  assign \new_[33616]_  = \new_[33615]_  & \new_[33612]_ ;
  assign \new_[33619]_  = A299 & ~A298;
  assign \new_[33622]_  = A301 & A300;
  assign \new_[33623]_  = \new_[33622]_  & \new_[33619]_ ;
  assign \new_[33624]_  = \new_[33623]_  & \new_[33616]_ ;
  assign \new_[33628]_  = A167 & A168;
  assign \new_[33629]_  = A170 & \new_[33628]_ ;
  assign \new_[33632]_  = ~A232 & ~A166;
  assign \new_[33635]_  = ~A234 & A233;
  assign \new_[33636]_  = \new_[33635]_  & \new_[33632]_ ;
  assign \new_[33637]_  = \new_[33636]_  & \new_[33629]_ ;
  assign \new_[33640]_  = A236 & ~A235;
  assign \new_[33643]_  = ~A269 & ~A267;
  assign \new_[33644]_  = \new_[33643]_  & \new_[33640]_ ;
  assign \new_[33647]_  = A299 & ~A298;
  assign \new_[33650]_  = ~A302 & A300;
  assign \new_[33651]_  = \new_[33650]_  & \new_[33647]_ ;
  assign \new_[33652]_  = \new_[33651]_  & \new_[33644]_ ;
  assign \new_[33656]_  = A167 & A168;
  assign \new_[33657]_  = A170 & \new_[33656]_ ;
  assign \new_[33660]_  = ~A232 & ~A166;
  assign \new_[33663]_  = ~A234 & A233;
  assign \new_[33664]_  = \new_[33663]_  & \new_[33660]_ ;
  assign \new_[33665]_  = \new_[33664]_  & \new_[33657]_ ;
  assign \new_[33668]_  = A236 & ~A235;
  assign \new_[33671]_  = A266 & A265;
  assign \new_[33672]_  = \new_[33671]_  & \new_[33668]_ ;
  assign \new_[33675]_  = ~A299 & A298;
  assign \new_[33678]_  = A301 & A300;
  assign \new_[33679]_  = \new_[33678]_  & \new_[33675]_ ;
  assign \new_[33680]_  = \new_[33679]_  & \new_[33672]_ ;
  assign \new_[33684]_  = A167 & A168;
  assign \new_[33685]_  = A170 & \new_[33684]_ ;
  assign \new_[33688]_  = ~A232 & ~A166;
  assign \new_[33691]_  = ~A234 & A233;
  assign \new_[33692]_  = \new_[33691]_  & \new_[33688]_ ;
  assign \new_[33693]_  = \new_[33692]_  & \new_[33685]_ ;
  assign \new_[33696]_  = A236 & ~A235;
  assign \new_[33699]_  = A266 & A265;
  assign \new_[33700]_  = \new_[33699]_  & \new_[33696]_ ;
  assign \new_[33703]_  = ~A299 & A298;
  assign \new_[33706]_  = ~A302 & A300;
  assign \new_[33707]_  = \new_[33706]_  & \new_[33703]_ ;
  assign \new_[33708]_  = \new_[33707]_  & \new_[33700]_ ;
  assign \new_[33712]_  = A167 & A168;
  assign \new_[33713]_  = A170 & \new_[33712]_ ;
  assign \new_[33716]_  = ~A232 & ~A166;
  assign \new_[33719]_  = ~A234 & A233;
  assign \new_[33720]_  = \new_[33719]_  & \new_[33716]_ ;
  assign \new_[33721]_  = \new_[33720]_  & \new_[33713]_ ;
  assign \new_[33724]_  = A236 & ~A235;
  assign \new_[33727]_  = A266 & A265;
  assign \new_[33728]_  = \new_[33727]_  & \new_[33724]_ ;
  assign \new_[33731]_  = A299 & ~A298;
  assign \new_[33734]_  = A301 & A300;
  assign \new_[33735]_  = \new_[33734]_  & \new_[33731]_ ;
  assign \new_[33736]_  = \new_[33735]_  & \new_[33728]_ ;
  assign \new_[33740]_  = A167 & A168;
  assign \new_[33741]_  = A170 & \new_[33740]_ ;
  assign \new_[33744]_  = ~A232 & ~A166;
  assign \new_[33747]_  = ~A234 & A233;
  assign \new_[33748]_  = \new_[33747]_  & \new_[33744]_ ;
  assign \new_[33749]_  = \new_[33748]_  & \new_[33741]_ ;
  assign \new_[33752]_  = A236 & ~A235;
  assign \new_[33755]_  = A266 & A265;
  assign \new_[33756]_  = \new_[33755]_  & \new_[33752]_ ;
  assign \new_[33759]_  = A299 & ~A298;
  assign \new_[33762]_  = ~A302 & A300;
  assign \new_[33763]_  = \new_[33762]_  & \new_[33759]_ ;
  assign \new_[33764]_  = \new_[33763]_  & \new_[33756]_ ;
  assign \new_[33768]_  = A167 & A168;
  assign \new_[33769]_  = A170 & \new_[33768]_ ;
  assign \new_[33772]_  = ~A232 & ~A166;
  assign \new_[33775]_  = ~A234 & A233;
  assign \new_[33776]_  = \new_[33775]_  & \new_[33772]_ ;
  assign \new_[33777]_  = \new_[33776]_  & \new_[33769]_ ;
  assign \new_[33780]_  = A236 & ~A235;
  assign \new_[33783]_  = ~A266 & ~A265;
  assign \new_[33784]_  = \new_[33783]_  & \new_[33780]_ ;
  assign \new_[33787]_  = ~A299 & A298;
  assign \new_[33790]_  = A301 & A300;
  assign \new_[33791]_  = \new_[33790]_  & \new_[33787]_ ;
  assign \new_[33792]_  = \new_[33791]_  & \new_[33784]_ ;
  assign \new_[33796]_  = A167 & A168;
  assign \new_[33797]_  = A170 & \new_[33796]_ ;
  assign \new_[33800]_  = ~A232 & ~A166;
  assign \new_[33803]_  = ~A234 & A233;
  assign \new_[33804]_  = \new_[33803]_  & \new_[33800]_ ;
  assign \new_[33805]_  = \new_[33804]_  & \new_[33797]_ ;
  assign \new_[33808]_  = A236 & ~A235;
  assign \new_[33811]_  = ~A266 & ~A265;
  assign \new_[33812]_  = \new_[33811]_  & \new_[33808]_ ;
  assign \new_[33815]_  = ~A299 & A298;
  assign \new_[33818]_  = ~A302 & A300;
  assign \new_[33819]_  = \new_[33818]_  & \new_[33815]_ ;
  assign \new_[33820]_  = \new_[33819]_  & \new_[33812]_ ;
  assign \new_[33824]_  = A167 & A168;
  assign \new_[33825]_  = A170 & \new_[33824]_ ;
  assign \new_[33828]_  = ~A232 & ~A166;
  assign \new_[33831]_  = ~A234 & A233;
  assign \new_[33832]_  = \new_[33831]_  & \new_[33828]_ ;
  assign \new_[33833]_  = \new_[33832]_  & \new_[33825]_ ;
  assign \new_[33836]_  = A236 & ~A235;
  assign \new_[33839]_  = ~A266 & ~A265;
  assign \new_[33840]_  = \new_[33839]_  & \new_[33836]_ ;
  assign \new_[33843]_  = A299 & ~A298;
  assign \new_[33846]_  = A301 & A300;
  assign \new_[33847]_  = \new_[33846]_  & \new_[33843]_ ;
  assign \new_[33848]_  = \new_[33847]_  & \new_[33840]_ ;
  assign \new_[33852]_  = A167 & A168;
  assign \new_[33853]_  = A170 & \new_[33852]_ ;
  assign \new_[33856]_  = ~A232 & ~A166;
  assign \new_[33859]_  = ~A234 & A233;
  assign \new_[33860]_  = \new_[33859]_  & \new_[33856]_ ;
  assign \new_[33861]_  = \new_[33860]_  & \new_[33853]_ ;
  assign \new_[33864]_  = A236 & ~A235;
  assign \new_[33867]_  = ~A266 & ~A265;
  assign \new_[33868]_  = \new_[33867]_  & \new_[33864]_ ;
  assign \new_[33871]_  = A299 & ~A298;
  assign \new_[33874]_  = ~A302 & A300;
  assign \new_[33875]_  = \new_[33874]_  & \new_[33871]_ ;
  assign \new_[33876]_  = \new_[33875]_  & \new_[33868]_ ;
  assign \new_[33880]_  = A167 & A168;
  assign \new_[33881]_  = A170 & \new_[33880]_ ;
  assign \new_[33884]_  = A232 & ~A166;
  assign \new_[33887]_  = A234 & ~A233;
  assign \new_[33888]_  = \new_[33887]_  & \new_[33884]_ ;
  assign \new_[33889]_  = \new_[33888]_  & \new_[33881]_ ;
  assign \new_[33892]_  = A267 & A235;
  assign \new_[33895]_  = A269 & ~A268;
  assign \new_[33896]_  = \new_[33895]_  & \new_[33892]_ ;
  assign \new_[33899]_  = ~A299 & A298;
  assign \new_[33902]_  = A301 & A300;
  assign \new_[33903]_  = \new_[33902]_  & \new_[33899]_ ;
  assign \new_[33904]_  = \new_[33903]_  & \new_[33896]_ ;
  assign \new_[33908]_  = A167 & A168;
  assign \new_[33909]_  = A170 & \new_[33908]_ ;
  assign \new_[33912]_  = A232 & ~A166;
  assign \new_[33915]_  = A234 & ~A233;
  assign \new_[33916]_  = \new_[33915]_  & \new_[33912]_ ;
  assign \new_[33917]_  = \new_[33916]_  & \new_[33909]_ ;
  assign \new_[33920]_  = A267 & A235;
  assign \new_[33923]_  = A269 & ~A268;
  assign \new_[33924]_  = \new_[33923]_  & \new_[33920]_ ;
  assign \new_[33927]_  = ~A299 & A298;
  assign \new_[33930]_  = ~A302 & A300;
  assign \new_[33931]_  = \new_[33930]_  & \new_[33927]_ ;
  assign \new_[33932]_  = \new_[33931]_  & \new_[33924]_ ;
  assign \new_[33936]_  = A167 & A168;
  assign \new_[33937]_  = A170 & \new_[33936]_ ;
  assign \new_[33940]_  = A232 & ~A166;
  assign \new_[33943]_  = A234 & ~A233;
  assign \new_[33944]_  = \new_[33943]_  & \new_[33940]_ ;
  assign \new_[33945]_  = \new_[33944]_  & \new_[33937]_ ;
  assign \new_[33948]_  = A267 & A235;
  assign \new_[33951]_  = A269 & ~A268;
  assign \new_[33952]_  = \new_[33951]_  & \new_[33948]_ ;
  assign \new_[33955]_  = A299 & ~A298;
  assign \new_[33958]_  = A301 & A300;
  assign \new_[33959]_  = \new_[33958]_  & \new_[33955]_ ;
  assign \new_[33960]_  = \new_[33959]_  & \new_[33952]_ ;
  assign \new_[33964]_  = A167 & A168;
  assign \new_[33965]_  = A170 & \new_[33964]_ ;
  assign \new_[33968]_  = A232 & ~A166;
  assign \new_[33971]_  = A234 & ~A233;
  assign \new_[33972]_  = \new_[33971]_  & \new_[33968]_ ;
  assign \new_[33973]_  = \new_[33972]_  & \new_[33965]_ ;
  assign \new_[33976]_  = A267 & A235;
  assign \new_[33979]_  = A269 & ~A268;
  assign \new_[33980]_  = \new_[33979]_  & \new_[33976]_ ;
  assign \new_[33983]_  = A299 & ~A298;
  assign \new_[33986]_  = ~A302 & A300;
  assign \new_[33987]_  = \new_[33986]_  & \new_[33983]_ ;
  assign \new_[33988]_  = \new_[33987]_  & \new_[33980]_ ;
  assign \new_[33992]_  = A167 & A168;
  assign \new_[33993]_  = A170 & \new_[33992]_ ;
  assign \new_[33996]_  = A232 & ~A166;
  assign \new_[33999]_  = A234 & ~A233;
  assign \new_[34000]_  = \new_[33999]_  & \new_[33996]_ ;
  assign \new_[34001]_  = \new_[34000]_  & \new_[33993]_ ;
  assign \new_[34004]_  = ~A267 & A235;
  assign \new_[34007]_  = A298 & A268;
  assign \new_[34008]_  = \new_[34007]_  & \new_[34004]_ ;
  assign \new_[34011]_  = ~A300 & ~A299;
  assign \new_[34014]_  = A302 & ~A301;
  assign \new_[34015]_  = \new_[34014]_  & \new_[34011]_ ;
  assign \new_[34016]_  = \new_[34015]_  & \new_[34008]_ ;
  assign \new_[34020]_  = A167 & A168;
  assign \new_[34021]_  = A170 & \new_[34020]_ ;
  assign \new_[34024]_  = A232 & ~A166;
  assign \new_[34027]_  = A234 & ~A233;
  assign \new_[34028]_  = \new_[34027]_  & \new_[34024]_ ;
  assign \new_[34029]_  = \new_[34028]_  & \new_[34021]_ ;
  assign \new_[34032]_  = ~A267 & A235;
  assign \new_[34035]_  = ~A298 & A268;
  assign \new_[34036]_  = \new_[34035]_  & \new_[34032]_ ;
  assign \new_[34039]_  = ~A300 & A299;
  assign \new_[34042]_  = A302 & ~A301;
  assign \new_[34043]_  = \new_[34042]_  & \new_[34039]_ ;
  assign \new_[34044]_  = \new_[34043]_  & \new_[34036]_ ;
  assign \new_[34048]_  = A167 & A168;
  assign \new_[34049]_  = A170 & \new_[34048]_ ;
  assign \new_[34052]_  = A232 & ~A166;
  assign \new_[34055]_  = A234 & ~A233;
  assign \new_[34056]_  = \new_[34055]_  & \new_[34052]_ ;
  assign \new_[34057]_  = \new_[34056]_  & \new_[34049]_ ;
  assign \new_[34060]_  = ~A267 & A235;
  assign \new_[34063]_  = A298 & ~A269;
  assign \new_[34064]_  = \new_[34063]_  & \new_[34060]_ ;
  assign \new_[34067]_  = ~A300 & ~A299;
  assign \new_[34070]_  = A302 & ~A301;
  assign \new_[34071]_  = \new_[34070]_  & \new_[34067]_ ;
  assign \new_[34072]_  = \new_[34071]_  & \new_[34064]_ ;
  assign \new_[34076]_  = A167 & A168;
  assign \new_[34077]_  = A170 & \new_[34076]_ ;
  assign \new_[34080]_  = A232 & ~A166;
  assign \new_[34083]_  = A234 & ~A233;
  assign \new_[34084]_  = \new_[34083]_  & \new_[34080]_ ;
  assign \new_[34085]_  = \new_[34084]_  & \new_[34077]_ ;
  assign \new_[34088]_  = ~A267 & A235;
  assign \new_[34091]_  = ~A298 & ~A269;
  assign \new_[34092]_  = \new_[34091]_  & \new_[34088]_ ;
  assign \new_[34095]_  = ~A300 & A299;
  assign \new_[34098]_  = A302 & ~A301;
  assign \new_[34099]_  = \new_[34098]_  & \new_[34095]_ ;
  assign \new_[34100]_  = \new_[34099]_  & \new_[34092]_ ;
  assign \new_[34104]_  = A167 & A168;
  assign \new_[34105]_  = A170 & \new_[34104]_ ;
  assign \new_[34108]_  = A232 & ~A166;
  assign \new_[34111]_  = A234 & ~A233;
  assign \new_[34112]_  = \new_[34111]_  & \new_[34108]_ ;
  assign \new_[34113]_  = \new_[34112]_  & \new_[34105]_ ;
  assign \new_[34116]_  = A265 & A235;
  assign \new_[34119]_  = A298 & A266;
  assign \new_[34120]_  = \new_[34119]_  & \new_[34116]_ ;
  assign \new_[34123]_  = ~A300 & ~A299;
  assign \new_[34126]_  = A302 & ~A301;
  assign \new_[34127]_  = \new_[34126]_  & \new_[34123]_ ;
  assign \new_[34128]_  = \new_[34127]_  & \new_[34120]_ ;
  assign \new_[34132]_  = A167 & A168;
  assign \new_[34133]_  = A170 & \new_[34132]_ ;
  assign \new_[34136]_  = A232 & ~A166;
  assign \new_[34139]_  = A234 & ~A233;
  assign \new_[34140]_  = \new_[34139]_  & \new_[34136]_ ;
  assign \new_[34141]_  = \new_[34140]_  & \new_[34133]_ ;
  assign \new_[34144]_  = A265 & A235;
  assign \new_[34147]_  = ~A298 & A266;
  assign \new_[34148]_  = \new_[34147]_  & \new_[34144]_ ;
  assign \new_[34151]_  = ~A300 & A299;
  assign \new_[34154]_  = A302 & ~A301;
  assign \new_[34155]_  = \new_[34154]_  & \new_[34151]_ ;
  assign \new_[34156]_  = \new_[34155]_  & \new_[34148]_ ;
  assign \new_[34160]_  = A167 & A168;
  assign \new_[34161]_  = A170 & \new_[34160]_ ;
  assign \new_[34164]_  = A232 & ~A166;
  assign \new_[34167]_  = A234 & ~A233;
  assign \new_[34168]_  = \new_[34167]_  & \new_[34164]_ ;
  assign \new_[34169]_  = \new_[34168]_  & \new_[34161]_ ;
  assign \new_[34172]_  = ~A265 & A235;
  assign \new_[34175]_  = A298 & ~A266;
  assign \new_[34176]_  = \new_[34175]_  & \new_[34172]_ ;
  assign \new_[34179]_  = ~A300 & ~A299;
  assign \new_[34182]_  = A302 & ~A301;
  assign \new_[34183]_  = \new_[34182]_  & \new_[34179]_ ;
  assign \new_[34184]_  = \new_[34183]_  & \new_[34176]_ ;
  assign \new_[34188]_  = A167 & A168;
  assign \new_[34189]_  = A170 & \new_[34188]_ ;
  assign \new_[34192]_  = A232 & ~A166;
  assign \new_[34195]_  = A234 & ~A233;
  assign \new_[34196]_  = \new_[34195]_  & \new_[34192]_ ;
  assign \new_[34197]_  = \new_[34196]_  & \new_[34189]_ ;
  assign \new_[34200]_  = ~A265 & A235;
  assign \new_[34203]_  = ~A298 & ~A266;
  assign \new_[34204]_  = \new_[34203]_  & \new_[34200]_ ;
  assign \new_[34207]_  = ~A300 & A299;
  assign \new_[34210]_  = A302 & ~A301;
  assign \new_[34211]_  = \new_[34210]_  & \new_[34207]_ ;
  assign \new_[34212]_  = \new_[34211]_  & \new_[34204]_ ;
  assign \new_[34216]_  = A167 & A168;
  assign \new_[34217]_  = A170 & \new_[34216]_ ;
  assign \new_[34220]_  = A232 & ~A166;
  assign \new_[34223]_  = A234 & ~A233;
  assign \new_[34224]_  = \new_[34223]_  & \new_[34220]_ ;
  assign \new_[34225]_  = \new_[34224]_  & \new_[34217]_ ;
  assign \new_[34228]_  = A267 & ~A236;
  assign \new_[34231]_  = A269 & ~A268;
  assign \new_[34232]_  = \new_[34231]_  & \new_[34228]_ ;
  assign \new_[34235]_  = ~A299 & A298;
  assign \new_[34238]_  = A301 & A300;
  assign \new_[34239]_  = \new_[34238]_  & \new_[34235]_ ;
  assign \new_[34240]_  = \new_[34239]_  & \new_[34232]_ ;
  assign \new_[34244]_  = A167 & A168;
  assign \new_[34245]_  = A170 & \new_[34244]_ ;
  assign \new_[34248]_  = A232 & ~A166;
  assign \new_[34251]_  = A234 & ~A233;
  assign \new_[34252]_  = \new_[34251]_  & \new_[34248]_ ;
  assign \new_[34253]_  = \new_[34252]_  & \new_[34245]_ ;
  assign \new_[34256]_  = A267 & ~A236;
  assign \new_[34259]_  = A269 & ~A268;
  assign \new_[34260]_  = \new_[34259]_  & \new_[34256]_ ;
  assign \new_[34263]_  = ~A299 & A298;
  assign \new_[34266]_  = ~A302 & A300;
  assign \new_[34267]_  = \new_[34266]_  & \new_[34263]_ ;
  assign \new_[34268]_  = \new_[34267]_  & \new_[34260]_ ;
  assign \new_[34272]_  = A167 & A168;
  assign \new_[34273]_  = A170 & \new_[34272]_ ;
  assign \new_[34276]_  = A232 & ~A166;
  assign \new_[34279]_  = A234 & ~A233;
  assign \new_[34280]_  = \new_[34279]_  & \new_[34276]_ ;
  assign \new_[34281]_  = \new_[34280]_  & \new_[34273]_ ;
  assign \new_[34284]_  = A267 & ~A236;
  assign \new_[34287]_  = A269 & ~A268;
  assign \new_[34288]_  = \new_[34287]_  & \new_[34284]_ ;
  assign \new_[34291]_  = A299 & ~A298;
  assign \new_[34294]_  = A301 & A300;
  assign \new_[34295]_  = \new_[34294]_  & \new_[34291]_ ;
  assign \new_[34296]_  = \new_[34295]_  & \new_[34288]_ ;
  assign \new_[34300]_  = A167 & A168;
  assign \new_[34301]_  = A170 & \new_[34300]_ ;
  assign \new_[34304]_  = A232 & ~A166;
  assign \new_[34307]_  = A234 & ~A233;
  assign \new_[34308]_  = \new_[34307]_  & \new_[34304]_ ;
  assign \new_[34309]_  = \new_[34308]_  & \new_[34301]_ ;
  assign \new_[34312]_  = A267 & ~A236;
  assign \new_[34315]_  = A269 & ~A268;
  assign \new_[34316]_  = \new_[34315]_  & \new_[34312]_ ;
  assign \new_[34319]_  = A299 & ~A298;
  assign \new_[34322]_  = ~A302 & A300;
  assign \new_[34323]_  = \new_[34322]_  & \new_[34319]_ ;
  assign \new_[34324]_  = \new_[34323]_  & \new_[34316]_ ;
  assign \new_[34328]_  = A167 & A168;
  assign \new_[34329]_  = A170 & \new_[34328]_ ;
  assign \new_[34332]_  = A232 & ~A166;
  assign \new_[34335]_  = A234 & ~A233;
  assign \new_[34336]_  = \new_[34335]_  & \new_[34332]_ ;
  assign \new_[34337]_  = \new_[34336]_  & \new_[34329]_ ;
  assign \new_[34340]_  = ~A267 & ~A236;
  assign \new_[34343]_  = A298 & A268;
  assign \new_[34344]_  = \new_[34343]_  & \new_[34340]_ ;
  assign \new_[34347]_  = ~A300 & ~A299;
  assign \new_[34350]_  = A302 & ~A301;
  assign \new_[34351]_  = \new_[34350]_  & \new_[34347]_ ;
  assign \new_[34352]_  = \new_[34351]_  & \new_[34344]_ ;
  assign \new_[34356]_  = A167 & A168;
  assign \new_[34357]_  = A170 & \new_[34356]_ ;
  assign \new_[34360]_  = A232 & ~A166;
  assign \new_[34363]_  = A234 & ~A233;
  assign \new_[34364]_  = \new_[34363]_  & \new_[34360]_ ;
  assign \new_[34365]_  = \new_[34364]_  & \new_[34357]_ ;
  assign \new_[34368]_  = ~A267 & ~A236;
  assign \new_[34371]_  = ~A298 & A268;
  assign \new_[34372]_  = \new_[34371]_  & \new_[34368]_ ;
  assign \new_[34375]_  = ~A300 & A299;
  assign \new_[34378]_  = A302 & ~A301;
  assign \new_[34379]_  = \new_[34378]_  & \new_[34375]_ ;
  assign \new_[34380]_  = \new_[34379]_  & \new_[34372]_ ;
  assign \new_[34384]_  = A167 & A168;
  assign \new_[34385]_  = A170 & \new_[34384]_ ;
  assign \new_[34388]_  = A232 & ~A166;
  assign \new_[34391]_  = A234 & ~A233;
  assign \new_[34392]_  = \new_[34391]_  & \new_[34388]_ ;
  assign \new_[34393]_  = \new_[34392]_  & \new_[34385]_ ;
  assign \new_[34396]_  = ~A267 & ~A236;
  assign \new_[34399]_  = A298 & ~A269;
  assign \new_[34400]_  = \new_[34399]_  & \new_[34396]_ ;
  assign \new_[34403]_  = ~A300 & ~A299;
  assign \new_[34406]_  = A302 & ~A301;
  assign \new_[34407]_  = \new_[34406]_  & \new_[34403]_ ;
  assign \new_[34408]_  = \new_[34407]_  & \new_[34400]_ ;
  assign \new_[34412]_  = A167 & A168;
  assign \new_[34413]_  = A170 & \new_[34412]_ ;
  assign \new_[34416]_  = A232 & ~A166;
  assign \new_[34419]_  = A234 & ~A233;
  assign \new_[34420]_  = \new_[34419]_  & \new_[34416]_ ;
  assign \new_[34421]_  = \new_[34420]_  & \new_[34413]_ ;
  assign \new_[34424]_  = ~A267 & ~A236;
  assign \new_[34427]_  = ~A298 & ~A269;
  assign \new_[34428]_  = \new_[34427]_  & \new_[34424]_ ;
  assign \new_[34431]_  = ~A300 & A299;
  assign \new_[34434]_  = A302 & ~A301;
  assign \new_[34435]_  = \new_[34434]_  & \new_[34431]_ ;
  assign \new_[34436]_  = \new_[34435]_  & \new_[34428]_ ;
  assign \new_[34440]_  = A167 & A168;
  assign \new_[34441]_  = A170 & \new_[34440]_ ;
  assign \new_[34444]_  = A232 & ~A166;
  assign \new_[34447]_  = A234 & ~A233;
  assign \new_[34448]_  = \new_[34447]_  & \new_[34444]_ ;
  assign \new_[34449]_  = \new_[34448]_  & \new_[34441]_ ;
  assign \new_[34452]_  = A265 & ~A236;
  assign \new_[34455]_  = A298 & A266;
  assign \new_[34456]_  = \new_[34455]_  & \new_[34452]_ ;
  assign \new_[34459]_  = ~A300 & ~A299;
  assign \new_[34462]_  = A302 & ~A301;
  assign \new_[34463]_  = \new_[34462]_  & \new_[34459]_ ;
  assign \new_[34464]_  = \new_[34463]_  & \new_[34456]_ ;
  assign \new_[34468]_  = A167 & A168;
  assign \new_[34469]_  = A170 & \new_[34468]_ ;
  assign \new_[34472]_  = A232 & ~A166;
  assign \new_[34475]_  = A234 & ~A233;
  assign \new_[34476]_  = \new_[34475]_  & \new_[34472]_ ;
  assign \new_[34477]_  = \new_[34476]_  & \new_[34469]_ ;
  assign \new_[34480]_  = A265 & ~A236;
  assign \new_[34483]_  = ~A298 & A266;
  assign \new_[34484]_  = \new_[34483]_  & \new_[34480]_ ;
  assign \new_[34487]_  = ~A300 & A299;
  assign \new_[34490]_  = A302 & ~A301;
  assign \new_[34491]_  = \new_[34490]_  & \new_[34487]_ ;
  assign \new_[34492]_  = \new_[34491]_  & \new_[34484]_ ;
  assign \new_[34496]_  = A167 & A168;
  assign \new_[34497]_  = A170 & \new_[34496]_ ;
  assign \new_[34500]_  = A232 & ~A166;
  assign \new_[34503]_  = A234 & ~A233;
  assign \new_[34504]_  = \new_[34503]_  & \new_[34500]_ ;
  assign \new_[34505]_  = \new_[34504]_  & \new_[34497]_ ;
  assign \new_[34508]_  = ~A265 & ~A236;
  assign \new_[34511]_  = A298 & ~A266;
  assign \new_[34512]_  = \new_[34511]_  & \new_[34508]_ ;
  assign \new_[34515]_  = ~A300 & ~A299;
  assign \new_[34518]_  = A302 & ~A301;
  assign \new_[34519]_  = \new_[34518]_  & \new_[34515]_ ;
  assign \new_[34520]_  = \new_[34519]_  & \new_[34512]_ ;
  assign \new_[34524]_  = A167 & A168;
  assign \new_[34525]_  = A170 & \new_[34524]_ ;
  assign \new_[34528]_  = A232 & ~A166;
  assign \new_[34531]_  = A234 & ~A233;
  assign \new_[34532]_  = \new_[34531]_  & \new_[34528]_ ;
  assign \new_[34533]_  = \new_[34532]_  & \new_[34525]_ ;
  assign \new_[34536]_  = ~A265 & ~A236;
  assign \new_[34539]_  = ~A298 & ~A266;
  assign \new_[34540]_  = \new_[34539]_  & \new_[34536]_ ;
  assign \new_[34543]_  = ~A300 & A299;
  assign \new_[34546]_  = A302 & ~A301;
  assign \new_[34547]_  = \new_[34546]_  & \new_[34543]_ ;
  assign \new_[34548]_  = \new_[34547]_  & \new_[34540]_ ;
  assign \new_[34552]_  = A167 & A168;
  assign \new_[34553]_  = A170 & \new_[34552]_ ;
  assign \new_[34556]_  = A232 & ~A166;
  assign \new_[34559]_  = ~A234 & ~A233;
  assign \new_[34560]_  = \new_[34559]_  & \new_[34556]_ ;
  assign \new_[34561]_  = \new_[34560]_  & \new_[34553]_ ;
  assign \new_[34564]_  = A236 & ~A235;
  assign \new_[34567]_  = A268 & ~A267;
  assign \new_[34568]_  = \new_[34567]_  & \new_[34564]_ ;
  assign \new_[34571]_  = ~A299 & A298;
  assign \new_[34574]_  = A301 & A300;
  assign \new_[34575]_  = \new_[34574]_  & \new_[34571]_ ;
  assign \new_[34576]_  = \new_[34575]_  & \new_[34568]_ ;
  assign \new_[34580]_  = A167 & A168;
  assign \new_[34581]_  = A170 & \new_[34580]_ ;
  assign \new_[34584]_  = A232 & ~A166;
  assign \new_[34587]_  = ~A234 & ~A233;
  assign \new_[34588]_  = \new_[34587]_  & \new_[34584]_ ;
  assign \new_[34589]_  = \new_[34588]_  & \new_[34581]_ ;
  assign \new_[34592]_  = A236 & ~A235;
  assign \new_[34595]_  = A268 & ~A267;
  assign \new_[34596]_  = \new_[34595]_  & \new_[34592]_ ;
  assign \new_[34599]_  = ~A299 & A298;
  assign \new_[34602]_  = ~A302 & A300;
  assign \new_[34603]_  = \new_[34602]_  & \new_[34599]_ ;
  assign \new_[34604]_  = \new_[34603]_  & \new_[34596]_ ;
  assign \new_[34608]_  = A167 & A168;
  assign \new_[34609]_  = A170 & \new_[34608]_ ;
  assign \new_[34612]_  = A232 & ~A166;
  assign \new_[34615]_  = ~A234 & ~A233;
  assign \new_[34616]_  = \new_[34615]_  & \new_[34612]_ ;
  assign \new_[34617]_  = \new_[34616]_  & \new_[34609]_ ;
  assign \new_[34620]_  = A236 & ~A235;
  assign \new_[34623]_  = A268 & ~A267;
  assign \new_[34624]_  = \new_[34623]_  & \new_[34620]_ ;
  assign \new_[34627]_  = A299 & ~A298;
  assign \new_[34630]_  = A301 & A300;
  assign \new_[34631]_  = \new_[34630]_  & \new_[34627]_ ;
  assign \new_[34632]_  = \new_[34631]_  & \new_[34624]_ ;
  assign \new_[34636]_  = A167 & A168;
  assign \new_[34637]_  = A170 & \new_[34636]_ ;
  assign \new_[34640]_  = A232 & ~A166;
  assign \new_[34643]_  = ~A234 & ~A233;
  assign \new_[34644]_  = \new_[34643]_  & \new_[34640]_ ;
  assign \new_[34645]_  = \new_[34644]_  & \new_[34637]_ ;
  assign \new_[34648]_  = A236 & ~A235;
  assign \new_[34651]_  = A268 & ~A267;
  assign \new_[34652]_  = \new_[34651]_  & \new_[34648]_ ;
  assign \new_[34655]_  = A299 & ~A298;
  assign \new_[34658]_  = ~A302 & A300;
  assign \new_[34659]_  = \new_[34658]_  & \new_[34655]_ ;
  assign \new_[34660]_  = \new_[34659]_  & \new_[34652]_ ;
  assign \new_[34664]_  = A167 & A168;
  assign \new_[34665]_  = A170 & \new_[34664]_ ;
  assign \new_[34668]_  = A232 & ~A166;
  assign \new_[34671]_  = ~A234 & ~A233;
  assign \new_[34672]_  = \new_[34671]_  & \new_[34668]_ ;
  assign \new_[34673]_  = \new_[34672]_  & \new_[34665]_ ;
  assign \new_[34676]_  = A236 & ~A235;
  assign \new_[34679]_  = ~A269 & ~A267;
  assign \new_[34680]_  = \new_[34679]_  & \new_[34676]_ ;
  assign \new_[34683]_  = ~A299 & A298;
  assign \new_[34686]_  = A301 & A300;
  assign \new_[34687]_  = \new_[34686]_  & \new_[34683]_ ;
  assign \new_[34688]_  = \new_[34687]_  & \new_[34680]_ ;
  assign \new_[34692]_  = A167 & A168;
  assign \new_[34693]_  = A170 & \new_[34692]_ ;
  assign \new_[34696]_  = A232 & ~A166;
  assign \new_[34699]_  = ~A234 & ~A233;
  assign \new_[34700]_  = \new_[34699]_  & \new_[34696]_ ;
  assign \new_[34701]_  = \new_[34700]_  & \new_[34693]_ ;
  assign \new_[34704]_  = A236 & ~A235;
  assign \new_[34707]_  = ~A269 & ~A267;
  assign \new_[34708]_  = \new_[34707]_  & \new_[34704]_ ;
  assign \new_[34711]_  = ~A299 & A298;
  assign \new_[34714]_  = ~A302 & A300;
  assign \new_[34715]_  = \new_[34714]_  & \new_[34711]_ ;
  assign \new_[34716]_  = \new_[34715]_  & \new_[34708]_ ;
  assign \new_[34720]_  = A167 & A168;
  assign \new_[34721]_  = A170 & \new_[34720]_ ;
  assign \new_[34724]_  = A232 & ~A166;
  assign \new_[34727]_  = ~A234 & ~A233;
  assign \new_[34728]_  = \new_[34727]_  & \new_[34724]_ ;
  assign \new_[34729]_  = \new_[34728]_  & \new_[34721]_ ;
  assign \new_[34732]_  = A236 & ~A235;
  assign \new_[34735]_  = ~A269 & ~A267;
  assign \new_[34736]_  = \new_[34735]_  & \new_[34732]_ ;
  assign \new_[34739]_  = A299 & ~A298;
  assign \new_[34742]_  = A301 & A300;
  assign \new_[34743]_  = \new_[34742]_  & \new_[34739]_ ;
  assign \new_[34744]_  = \new_[34743]_  & \new_[34736]_ ;
  assign \new_[34748]_  = A167 & A168;
  assign \new_[34749]_  = A170 & \new_[34748]_ ;
  assign \new_[34752]_  = A232 & ~A166;
  assign \new_[34755]_  = ~A234 & ~A233;
  assign \new_[34756]_  = \new_[34755]_  & \new_[34752]_ ;
  assign \new_[34757]_  = \new_[34756]_  & \new_[34749]_ ;
  assign \new_[34760]_  = A236 & ~A235;
  assign \new_[34763]_  = ~A269 & ~A267;
  assign \new_[34764]_  = \new_[34763]_  & \new_[34760]_ ;
  assign \new_[34767]_  = A299 & ~A298;
  assign \new_[34770]_  = ~A302 & A300;
  assign \new_[34771]_  = \new_[34770]_  & \new_[34767]_ ;
  assign \new_[34772]_  = \new_[34771]_  & \new_[34764]_ ;
  assign \new_[34776]_  = A167 & A168;
  assign \new_[34777]_  = A170 & \new_[34776]_ ;
  assign \new_[34780]_  = A232 & ~A166;
  assign \new_[34783]_  = ~A234 & ~A233;
  assign \new_[34784]_  = \new_[34783]_  & \new_[34780]_ ;
  assign \new_[34785]_  = \new_[34784]_  & \new_[34777]_ ;
  assign \new_[34788]_  = A236 & ~A235;
  assign \new_[34791]_  = A266 & A265;
  assign \new_[34792]_  = \new_[34791]_  & \new_[34788]_ ;
  assign \new_[34795]_  = ~A299 & A298;
  assign \new_[34798]_  = A301 & A300;
  assign \new_[34799]_  = \new_[34798]_  & \new_[34795]_ ;
  assign \new_[34800]_  = \new_[34799]_  & \new_[34792]_ ;
  assign \new_[34804]_  = A167 & A168;
  assign \new_[34805]_  = A170 & \new_[34804]_ ;
  assign \new_[34808]_  = A232 & ~A166;
  assign \new_[34811]_  = ~A234 & ~A233;
  assign \new_[34812]_  = \new_[34811]_  & \new_[34808]_ ;
  assign \new_[34813]_  = \new_[34812]_  & \new_[34805]_ ;
  assign \new_[34816]_  = A236 & ~A235;
  assign \new_[34819]_  = A266 & A265;
  assign \new_[34820]_  = \new_[34819]_  & \new_[34816]_ ;
  assign \new_[34823]_  = ~A299 & A298;
  assign \new_[34826]_  = ~A302 & A300;
  assign \new_[34827]_  = \new_[34826]_  & \new_[34823]_ ;
  assign \new_[34828]_  = \new_[34827]_  & \new_[34820]_ ;
  assign \new_[34832]_  = A167 & A168;
  assign \new_[34833]_  = A170 & \new_[34832]_ ;
  assign \new_[34836]_  = A232 & ~A166;
  assign \new_[34839]_  = ~A234 & ~A233;
  assign \new_[34840]_  = \new_[34839]_  & \new_[34836]_ ;
  assign \new_[34841]_  = \new_[34840]_  & \new_[34833]_ ;
  assign \new_[34844]_  = A236 & ~A235;
  assign \new_[34847]_  = A266 & A265;
  assign \new_[34848]_  = \new_[34847]_  & \new_[34844]_ ;
  assign \new_[34851]_  = A299 & ~A298;
  assign \new_[34854]_  = A301 & A300;
  assign \new_[34855]_  = \new_[34854]_  & \new_[34851]_ ;
  assign \new_[34856]_  = \new_[34855]_  & \new_[34848]_ ;
  assign \new_[34860]_  = A167 & A168;
  assign \new_[34861]_  = A170 & \new_[34860]_ ;
  assign \new_[34864]_  = A232 & ~A166;
  assign \new_[34867]_  = ~A234 & ~A233;
  assign \new_[34868]_  = \new_[34867]_  & \new_[34864]_ ;
  assign \new_[34869]_  = \new_[34868]_  & \new_[34861]_ ;
  assign \new_[34872]_  = A236 & ~A235;
  assign \new_[34875]_  = A266 & A265;
  assign \new_[34876]_  = \new_[34875]_  & \new_[34872]_ ;
  assign \new_[34879]_  = A299 & ~A298;
  assign \new_[34882]_  = ~A302 & A300;
  assign \new_[34883]_  = \new_[34882]_  & \new_[34879]_ ;
  assign \new_[34884]_  = \new_[34883]_  & \new_[34876]_ ;
  assign \new_[34888]_  = A167 & A168;
  assign \new_[34889]_  = A170 & \new_[34888]_ ;
  assign \new_[34892]_  = A232 & ~A166;
  assign \new_[34895]_  = ~A234 & ~A233;
  assign \new_[34896]_  = \new_[34895]_  & \new_[34892]_ ;
  assign \new_[34897]_  = \new_[34896]_  & \new_[34889]_ ;
  assign \new_[34900]_  = A236 & ~A235;
  assign \new_[34903]_  = ~A266 & ~A265;
  assign \new_[34904]_  = \new_[34903]_  & \new_[34900]_ ;
  assign \new_[34907]_  = ~A299 & A298;
  assign \new_[34910]_  = A301 & A300;
  assign \new_[34911]_  = \new_[34910]_  & \new_[34907]_ ;
  assign \new_[34912]_  = \new_[34911]_  & \new_[34904]_ ;
  assign \new_[34916]_  = A167 & A168;
  assign \new_[34917]_  = A170 & \new_[34916]_ ;
  assign \new_[34920]_  = A232 & ~A166;
  assign \new_[34923]_  = ~A234 & ~A233;
  assign \new_[34924]_  = \new_[34923]_  & \new_[34920]_ ;
  assign \new_[34925]_  = \new_[34924]_  & \new_[34917]_ ;
  assign \new_[34928]_  = A236 & ~A235;
  assign \new_[34931]_  = ~A266 & ~A265;
  assign \new_[34932]_  = \new_[34931]_  & \new_[34928]_ ;
  assign \new_[34935]_  = ~A299 & A298;
  assign \new_[34938]_  = ~A302 & A300;
  assign \new_[34939]_  = \new_[34938]_  & \new_[34935]_ ;
  assign \new_[34940]_  = \new_[34939]_  & \new_[34932]_ ;
  assign \new_[34944]_  = A167 & A168;
  assign \new_[34945]_  = A170 & \new_[34944]_ ;
  assign \new_[34948]_  = A232 & ~A166;
  assign \new_[34951]_  = ~A234 & ~A233;
  assign \new_[34952]_  = \new_[34951]_  & \new_[34948]_ ;
  assign \new_[34953]_  = \new_[34952]_  & \new_[34945]_ ;
  assign \new_[34956]_  = A236 & ~A235;
  assign \new_[34959]_  = ~A266 & ~A265;
  assign \new_[34960]_  = \new_[34959]_  & \new_[34956]_ ;
  assign \new_[34963]_  = A299 & ~A298;
  assign \new_[34966]_  = A301 & A300;
  assign \new_[34967]_  = \new_[34966]_  & \new_[34963]_ ;
  assign \new_[34968]_  = \new_[34967]_  & \new_[34960]_ ;
  assign \new_[34972]_  = A167 & A168;
  assign \new_[34973]_  = A170 & \new_[34972]_ ;
  assign \new_[34976]_  = A232 & ~A166;
  assign \new_[34979]_  = ~A234 & ~A233;
  assign \new_[34980]_  = \new_[34979]_  & \new_[34976]_ ;
  assign \new_[34981]_  = \new_[34980]_  & \new_[34973]_ ;
  assign \new_[34984]_  = A236 & ~A235;
  assign \new_[34987]_  = ~A266 & ~A265;
  assign \new_[34988]_  = \new_[34987]_  & \new_[34984]_ ;
  assign \new_[34991]_  = A299 & ~A298;
  assign \new_[34994]_  = ~A302 & A300;
  assign \new_[34995]_  = \new_[34994]_  & \new_[34991]_ ;
  assign \new_[34996]_  = \new_[34995]_  & \new_[34988]_ ;
  assign \new_[35000]_  = ~A167 & A168;
  assign \new_[35001]_  = A170 & \new_[35000]_ ;
  assign \new_[35004]_  = ~A232 & A166;
  assign \new_[35007]_  = A234 & A233;
  assign \new_[35008]_  = \new_[35007]_  & \new_[35004]_ ;
  assign \new_[35009]_  = \new_[35008]_  & \new_[35001]_ ;
  assign \new_[35012]_  = A267 & A235;
  assign \new_[35015]_  = A269 & ~A268;
  assign \new_[35016]_  = \new_[35015]_  & \new_[35012]_ ;
  assign \new_[35019]_  = ~A299 & A298;
  assign \new_[35022]_  = A301 & A300;
  assign \new_[35023]_  = \new_[35022]_  & \new_[35019]_ ;
  assign \new_[35024]_  = \new_[35023]_  & \new_[35016]_ ;
  assign \new_[35028]_  = ~A167 & A168;
  assign \new_[35029]_  = A170 & \new_[35028]_ ;
  assign \new_[35032]_  = ~A232 & A166;
  assign \new_[35035]_  = A234 & A233;
  assign \new_[35036]_  = \new_[35035]_  & \new_[35032]_ ;
  assign \new_[35037]_  = \new_[35036]_  & \new_[35029]_ ;
  assign \new_[35040]_  = A267 & A235;
  assign \new_[35043]_  = A269 & ~A268;
  assign \new_[35044]_  = \new_[35043]_  & \new_[35040]_ ;
  assign \new_[35047]_  = ~A299 & A298;
  assign \new_[35050]_  = ~A302 & A300;
  assign \new_[35051]_  = \new_[35050]_  & \new_[35047]_ ;
  assign \new_[35052]_  = \new_[35051]_  & \new_[35044]_ ;
  assign \new_[35056]_  = ~A167 & A168;
  assign \new_[35057]_  = A170 & \new_[35056]_ ;
  assign \new_[35060]_  = ~A232 & A166;
  assign \new_[35063]_  = A234 & A233;
  assign \new_[35064]_  = \new_[35063]_  & \new_[35060]_ ;
  assign \new_[35065]_  = \new_[35064]_  & \new_[35057]_ ;
  assign \new_[35068]_  = A267 & A235;
  assign \new_[35071]_  = A269 & ~A268;
  assign \new_[35072]_  = \new_[35071]_  & \new_[35068]_ ;
  assign \new_[35075]_  = A299 & ~A298;
  assign \new_[35078]_  = A301 & A300;
  assign \new_[35079]_  = \new_[35078]_  & \new_[35075]_ ;
  assign \new_[35080]_  = \new_[35079]_  & \new_[35072]_ ;
  assign \new_[35084]_  = ~A167 & A168;
  assign \new_[35085]_  = A170 & \new_[35084]_ ;
  assign \new_[35088]_  = ~A232 & A166;
  assign \new_[35091]_  = A234 & A233;
  assign \new_[35092]_  = \new_[35091]_  & \new_[35088]_ ;
  assign \new_[35093]_  = \new_[35092]_  & \new_[35085]_ ;
  assign \new_[35096]_  = A267 & A235;
  assign \new_[35099]_  = A269 & ~A268;
  assign \new_[35100]_  = \new_[35099]_  & \new_[35096]_ ;
  assign \new_[35103]_  = A299 & ~A298;
  assign \new_[35106]_  = ~A302 & A300;
  assign \new_[35107]_  = \new_[35106]_  & \new_[35103]_ ;
  assign \new_[35108]_  = \new_[35107]_  & \new_[35100]_ ;
  assign \new_[35112]_  = ~A167 & A168;
  assign \new_[35113]_  = A170 & \new_[35112]_ ;
  assign \new_[35116]_  = ~A232 & A166;
  assign \new_[35119]_  = A234 & A233;
  assign \new_[35120]_  = \new_[35119]_  & \new_[35116]_ ;
  assign \new_[35121]_  = \new_[35120]_  & \new_[35113]_ ;
  assign \new_[35124]_  = ~A267 & A235;
  assign \new_[35127]_  = A298 & A268;
  assign \new_[35128]_  = \new_[35127]_  & \new_[35124]_ ;
  assign \new_[35131]_  = ~A300 & ~A299;
  assign \new_[35134]_  = A302 & ~A301;
  assign \new_[35135]_  = \new_[35134]_  & \new_[35131]_ ;
  assign \new_[35136]_  = \new_[35135]_  & \new_[35128]_ ;
  assign \new_[35140]_  = ~A167 & A168;
  assign \new_[35141]_  = A170 & \new_[35140]_ ;
  assign \new_[35144]_  = ~A232 & A166;
  assign \new_[35147]_  = A234 & A233;
  assign \new_[35148]_  = \new_[35147]_  & \new_[35144]_ ;
  assign \new_[35149]_  = \new_[35148]_  & \new_[35141]_ ;
  assign \new_[35152]_  = ~A267 & A235;
  assign \new_[35155]_  = ~A298 & A268;
  assign \new_[35156]_  = \new_[35155]_  & \new_[35152]_ ;
  assign \new_[35159]_  = ~A300 & A299;
  assign \new_[35162]_  = A302 & ~A301;
  assign \new_[35163]_  = \new_[35162]_  & \new_[35159]_ ;
  assign \new_[35164]_  = \new_[35163]_  & \new_[35156]_ ;
  assign \new_[35168]_  = ~A167 & A168;
  assign \new_[35169]_  = A170 & \new_[35168]_ ;
  assign \new_[35172]_  = ~A232 & A166;
  assign \new_[35175]_  = A234 & A233;
  assign \new_[35176]_  = \new_[35175]_  & \new_[35172]_ ;
  assign \new_[35177]_  = \new_[35176]_  & \new_[35169]_ ;
  assign \new_[35180]_  = ~A267 & A235;
  assign \new_[35183]_  = A298 & ~A269;
  assign \new_[35184]_  = \new_[35183]_  & \new_[35180]_ ;
  assign \new_[35187]_  = ~A300 & ~A299;
  assign \new_[35190]_  = A302 & ~A301;
  assign \new_[35191]_  = \new_[35190]_  & \new_[35187]_ ;
  assign \new_[35192]_  = \new_[35191]_  & \new_[35184]_ ;
  assign \new_[35196]_  = ~A167 & A168;
  assign \new_[35197]_  = A170 & \new_[35196]_ ;
  assign \new_[35200]_  = ~A232 & A166;
  assign \new_[35203]_  = A234 & A233;
  assign \new_[35204]_  = \new_[35203]_  & \new_[35200]_ ;
  assign \new_[35205]_  = \new_[35204]_  & \new_[35197]_ ;
  assign \new_[35208]_  = ~A267 & A235;
  assign \new_[35211]_  = ~A298 & ~A269;
  assign \new_[35212]_  = \new_[35211]_  & \new_[35208]_ ;
  assign \new_[35215]_  = ~A300 & A299;
  assign \new_[35218]_  = A302 & ~A301;
  assign \new_[35219]_  = \new_[35218]_  & \new_[35215]_ ;
  assign \new_[35220]_  = \new_[35219]_  & \new_[35212]_ ;
  assign \new_[35224]_  = ~A167 & A168;
  assign \new_[35225]_  = A170 & \new_[35224]_ ;
  assign \new_[35228]_  = ~A232 & A166;
  assign \new_[35231]_  = A234 & A233;
  assign \new_[35232]_  = \new_[35231]_  & \new_[35228]_ ;
  assign \new_[35233]_  = \new_[35232]_  & \new_[35225]_ ;
  assign \new_[35236]_  = A265 & A235;
  assign \new_[35239]_  = A298 & A266;
  assign \new_[35240]_  = \new_[35239]_  & \new_[35236]_ ;
  assign \new_[35243]_  = ~A300 & ~A299;
  assign \new_[35246]_  = A302 & ~A301;
  assign \new_[35247]_  = \new_[35246]_  & \new_[35243]_ ;
  assign \new_[35248]_  = \new_[35247]_  & \new_[35240]_ ;
  assign \new_[35252]_  = ~A167 & A168;
  assign \new_[35253]_  = A170 & \new_[35252]_ ;
  assign \new_[35256]_  = ~A232 & A166;
  assign \new_[35259]_  = A234 & A233;
  assign \new_[35260]_  = \new_[35259]_  & \new_[35256]_ ;
  assign \new_[35261]_  = \new_[35260]_  & \new_[35253]_ ;
  assign \new_[35264]_  = A265 & A235;
  assign \new_[35267]_  = ~A298 & A266;
  assign \new_[35268]_  = \new_[35267]_  & \new_[35264]_ ;
  assign \new_[35271]_  = ~A300 & A299;
  assign \new_[35274]_  = A302 & ~A301;
  assign \new_[35275]_  = \new_[35274]_  & \new_[35271]_ ;
  assign \new_[35276]_  = \new_[35275]_  & \new_[35268]_ ;
  assign \new_[35280]_  = ~A167 & A168;
  assign \new_[35281]_  = A170 & \new_[35280]_ ;
  assign \new_[35284]_  = ~A232 & A166;
  assign \new_[35287]_  = A234 & A233;
  assign \new_[35288]_  = \new_[35287]_  & \new_[35284]_ ;
  assign \new_[35289]_  = \new_[35288]_  & \new_[35281]_ ;
  assign \new_[35292]_  = ~A265 & A235;
  assign \new_[35295]_  = A298 & ~A266;
  assign \new_[35296]_  = \new_[35295]_  & \new_[35292]_ ;
  assign \new_[35299]_  = ~A300 & ~A299;
  assign \new_[35302]_  = A302 & ~A301;
  assign \new_[35303]_  = \new_[35302]_  & \new_[35299]_ ;
  assign \new_[35304]_  = \new_[35303]_  & \new_[35296]_ ;
  assign \new_[35308]_  = ~A167 & A168;
  assign \new_[35309]_  = A170 & \new_[35308]_ ;
  assign \new_[35312]_  = ~A232 & A166;
  assign \new_[35315]_  = A234 & A233;
  assign \new_[35316]_  = \new_[35315]_  & \new_[35312]_ ;
  assign \new_[35317]_  = \new_[35316]_  & \new_[35309]_ ;
  assign \new_[35320]_  = ~A265 & A235;
  assign \new_[35323]_  = ~A298 & ~A266;
  assign \new_[35324]_  = \new_[35323]_  & \new_[35320]_ ;
  assign \new_[35327]_  = ~A300 & A299;
  assign \new_[35330]_  = A302 & ~A301;
  assign \new_[35331]_  = \new_[35330]_  & \new_[35327]_ ;
  assign \new_[35332]_  = \new_[35331]_  & \new_[35324]_ ;
  assign \new_[35336]_  = ~A167 & A168;
  assign \new_[35337]_  = A170 & \new_[35336]_ ;
  assign \new_[35340]_  = ~A232 & A166;
  assign \new_[35343]_  = A234 & A233;
  assign \new_[35344]_  = \new_[35343]_  & \new_[35340]_ ;
  assign \new_[35345]_  = \new_[35344]_  & \new_[35337]_ ;
  assign \new_[35348]_  = A267 & ~A236;
  assign \new_[35351]_  = A269 & ~A268;
  assign \new_[35352]_  = \new_[35351]_  & \new_[35348]_ ;
  assign \new_[35355]_  = ~A299 & A298;
  assign \new_[35358]_  = A301 & A300;
  assign \new_[35359]_  = \new_[35358]_  & \new_[35355]_ ;
  assign \new_[35360]_  = \new_[35359]_  & \new_[35352]_ ;
  assign \new_[35364]_  = ~A167 & A168;
  assign \new_[35365]_  = A170 & \new_[35364]_ ;
  assign \new_[35368]_  = ~A232 & A166;
  assign \new_[35371]_  = A234 & A233;
  assign \new_[35372]_  = \new_[35371]_  & \new_[35368]_ ;
  assign \new_[35373]_  = \new_[35372]_  & \new_[35365]_ ;
  assign \new_[35376]_  = A267 & ~A236;
  assign \new_[35379]_  = A269 & ~A268;
  assign \new_[35380]_  = \new_[35379]_  & \new_[35376]_ ;
  assign \new_[35383]_  = ~A299 & A298;
  assign \new_[35386]_  = ~A302 & A300;
  assign \new_[35387]_  = \new_[35386]_  & \new_[35383]_ ;
  assign \new_[35388]_  = \new_[35387]_  & \new_[35380]_ ;
  assign \new_[35392]_  = ~A167 & A168;
  assign \new_[35393]_  = A170 & \new_[35392]_ ;
  assign \new_[35396]_  = ~A232 & A166;
  assign \new_[35399]_  = A234 & A233;
  assign \new_[35400]_  = \new_[35399]_  & \new_[35396]_ ;
  assign \new_[35401]_  = \new_[35400]_  & \new_[35393]_ ;
  assign \new_[35404]_  = A267 & ~A236;
  assign \new_[35407]_  = A269 & ~A268;
  assign \new_[35408]_  = \new_[35407]_  & \new_[35404]_ ;
  assign \new_[35411]_  = A299 & ~A298;
  assign \new_[35414]_  = A301 & A300;
  assign \new_[35415]_  = \new_[35414]_  & \new_[35411]_ ;
  assign \new_[35416]_  = \new_[35415]_  & \new_[35408]_ ;
  assign \new_[35420]_  = ~A167 & A168;
  assign \new_[35421]_  = A170 & \new_[35420]_ ;
  assign \new_[35424]_  = ~A232 & A166;
  assign \new_[35427]_  = A234 & A233;
  assign \new_[35428]_  = \new_[35427]_  & \new_[35424]_ ;
  assign \new_[35429]_  = \new_[35428]_  & \new_[35421]_ ;
  assign \new_[35432]_  = A267 & ~A236;
  assign \new_[35435]_  = A269 & ~A268;
  assign \new_[35436]_  = \new_[35435]_  & \new_[35432]_ ;
  assign \new_[35439]_  = A299 & ~A298;
  assign \new_[35442]_  = ~A302 & A300;
  assign \new_[35443]_  = \new_[35442]_  & \new_[35439]_ ;
  assign \new_[35444]_  = \new_[35443]_  & \new_[35436]_ ;
  assign \new_[35448]_  = ~A167 & A168;
  assign \new_[35449]_  = A170 & \new_[35448]_ ;
  assign \new_[35452]_  = ~A232 & A166;
  assign \new_[35455]_  = A234 & A233;
  assign \new_[35456]_  = \new_[35455]_  & \new_[35452]_ ;
  assign \new_[35457]_  = \new_[35456]_  & \new_[35449]_ ;
  assign \new_[35460]_  = ~A267 & ~A236;
  assign \new_[35463]_  = A298 & A268;
  assign \new_[35464]_  = \new_[35463]_  & \new_[35460]_ ;
  assign \new_[35467]_  = ~A300 & ~A299;
  assign \new_[35470]_  = A302 & ~A301;
  assign \new_[35471]_  = \new_[35470]_  & \new_[35467]_ ;
  assign \new_[35472]_  = \new_[35471]_  & \new_[35464]_ ;
  assign \new_[35476]_  = ~A167 & A168;
  assign \new_[35477]_  = A170 & \new_[35476]_ ;
  assign \new_[35480]_  = ~A232 & A166;
  assign \new_[35483]_  = A234 & A233;
  assign \new_[35484]_  = \new_[35483]_  & \new_[35480]_ ;
  assign \new_[35485]_  = \new_[35484]_  & \new_[35477]_ ;
  assign \new_[35488]_  = ~A267 & ~A236;
  assign \new_[35491]_  = ~A298 & A268;
  assign \new_[35492]_  = \new_[35491]_  & \new_[35488]_ ;
  assign \new_[35495]_  = ~A300 & A299;
  assign \new_[35498]_  = A302 & ~A301;
  assign \new_[35499]_  = \new_[35498]_  & \new_[35495]_ ;
  assign \new_[35500]_  = \new_[35499]_  & \new_[35492]_ ;
  assign \new_[35504]_  = ~A167 & A168;
  assign \new_[35505]_  = A170 & \new_[35504]_ ;
  assign \new_[35508]_  = ~A232 & A166;
  assign \new_[35511]_  = A234 & A233;
  assign \new_[35512]_  = \new_[35511]_  & \new_[35508]_ ;
  assign \new_[35513]_  = \new_[35512]_  & \new_[35505]_ ;
  assign \new_[35516]_  = ~A267 & ~A236;
  assign \new_[35519]_  = A298 & ~A269;
  assign \new_[35520]_  = \new_[35519]_  & \new_[35516]_ ;
  assign \new_[35523]_  = ~A300 & ~A299;
  assign \new_[35526]_  = A302 & ~A301;
  assign \new_[35527]_  = \new_[35526]_  & \new_[35523]_ ;
  assign \new_[35528]_  = \new_[35527]_  & \new_[35520]_ ;
  assign \new_[35532]_  = ~A167 & A168;
  assign \new_[35533]_  = A170 & \new_[35532]_ ;
  assign \new_[35536]_  = ~A232 & A166;
  assign \new_[35539]_  = A234 & A233;
  assign \new_[35540]_  = \new_[35539]_  & \new_[35536]_ ;
  assign \new_[35541]_  = \new_[35540]_  & \new_[35533]_ ;
  assign \new_[35544]_  = ~A267 & ~A236;
  assign \new_[35547]_  = ~A298 & ~A269;
  assign \new_[35548]_  = \new_[35547]_  & \new_[35544]_ ;
  assign \new_[35551]_  = ~A300 & A299;
  assign \new_[35554]_  = A302 & ~A301;
  assign \new_[35555]_  = \new_[35554]_  & \new_[35551]_ ;
  assign \new_[35556]_  = \new_[35555]_  & \new_[35548]_ ;
  assign \new_[35560]_  = ~A167 & A168;
  assign \new_[35561]_  = A170 & \new_[35560]_ ;
  assign \new_[35564]_  = ~A232 & A166;
  assign \new_[35567]_  = A234 & A233;
  assign \new_[35568]_  = \new_[35567]_  & \new_[35564]_ ;
  assign \new_[35569]_  = \new_[35568]_  & \new_[35561]_ ;
  assign \new_[35572]_  = A265 & ~A236;
  assign \new_[35575]_  = A298 & A266;
  assign \new_[35576]_  = \new_[35575]_  & \new_[35572]_ ;
  assign \new_[35579]_  = ~A300 & ~A299;
  assign \new_[35582]_  = A302 & ~A301;
  assign \new_[35583]_  = \new_[35582]_  & \new_[35579]_ ;
  assign \new_[35584]_  = \new_[35583]_  & \new_[35576]_ ;
  assign \new_[35588]_  = ~A167 & A168;
  assign \new_[35589]_  = A170 & \new_[35588]_ ;
  assign \new_[35592]_  = ~A232 & A166;
  assign \new_[35595]_  = A234 & A233;
  assign \new_[35596]_  = \new_[35595]_  & \new_[35592]_ ;
  assign \new_[35597]_  = \new_[35596]_  & \new_[35589]_ ;
  assign \new_[35600]_  = A265 & ~A236;
  assign \new_[35603]_  = ~A298 & A266;
  assign \new_[35604]_  = \new_[35603]_  & \new_[35600]_ ;
  assign \new_[35607]_  = ~A300 & A299;
  assign \new_[35610]_  = A302 & ~A301;
  assign \new_[35611]_  = \new_[35610]_  & \new_[35607]_ ;
  assign \new_[35612]_  = \new_[35611]_  & \new_[35604]_ ;
  assign \new_[35616]_  = ~A167 & A168;
  assign \new_[35617]_  = A170 & \new_[35616]_ ;
  assign \new_[35620]_  = ~A232 & A166;
  assign \new_[35623]_  = A234 & A233;
  assign \new_[35624]_  = \new_[35623]_  & \new_[35620]_ ;
  assign \new_[35625]_  = \new_[35624]_  & \new_[35617]_ ;
  assign \new_[35628]_  = ~A265 & ~A236;
  assign \new_[35631]_  = A298 & ~A266;
  assign \new_[35632]_  = \new_[35631]_  & \new_[35628]_ ;
  assign \new_[35635]_  = ~A300 & ~A299;
  assign \new_[35638]_  = A302 & ~A301;
  assign \new_[35639]_  = \new_[35638]_  & \new_[35635]_ ;
  assign \new_[35640]_  = \new_[35639]_  & \new_[35632]_ ;
  assign \new_[35644]_  = ~A167 & A168;
  assign \new_[35645]_  = A170 & \new_[35644]_ ;
  assign \new_[35648]_  = ~A232 & A166;
  assign \new_[35651]_  = A234 & A233;
  assign \new_[35652]_  = \new_[35651]_  & \new_[35648]_ ;
  assign \new_[35653]_  = \new_[35652]_  & \new_[35645]_ ;
  assign \new_[35656]_  = ~A265 & ~A236;
  assign \new_[35659]_  = ~A298 & ~A266;
  assign \new_[35660]_  = \new_[35659]_  & \new_[35656]_ ;
  assign \new_[35663]_  = ~A300 & A299;
  assign \new_[35666]_  = A302 & ~A301;
  assign \new_[35667]_  = \new_[35666]_  & \new_[35663]_ ;
  assign \new_[35668]_  = \new_[35667]_  & \new_[35660]_ ;
  assign \new_[35672]_  = ~A167 & A168;
  assign \new_[35673]_  = A170 & \new_[35672]_ ;
  assign \new_[35676]_  = ~A232 & A166;
  assign \new_[35679]_  = ~A234 & A233;
  assign \new_[35680]_  = \new_[35679]_  & \new_[35676]_ ;
  assign \new_[35681]_  = \new_[35680]_  & \new_[35673]_ ;
  assign \new_[35684]_  = A236 & ~A235;
  assign \new_[35687]_  = A268 & ~A267;
  assign \new_[35688]_  = \new_[35687]_  & \new_[35684]_ ;
  assign \new_[35691]_  = ~A299 & A298;
  assign \new_[35694]_  = A301 & A300;
  assign \new_[35695]_  = \new_[35694]_  & \new_[35691]_ ;
  assign \new_[35696]_  = \new_[35695]_  & \new_[35688]_ ;
  assign \new_[35700]_  = ~A167 & A168;
  assign \new_[35701]_  = A170 & \new_[35700]_ ;
  assign \new_[35704]_  = ~A232 & A166;
  assign \new_[35707]_  = ~A234 & A233;
  assign \new_[35708]_  = \new_[35707]_  & \new_[35704]_ ;
  assign \new_[35709]_  = \new_[35708]_  & \new_[35701]_ ;
  assign \new_[35712]_  = A236 & ~A235;
  assign \new_[35715]_  = A268 & ~A267;
  assign \new_[35716]_  = \new_[35715]_  & \new_[35712]_ ;
  assign \new_[35719]_  = ~A299 & A298;
  assign \new_[35722]_  = ~A302 & A300;
  assign \new_[35723]_  = \new_[35722]_  & \new_[35719]_ ;
  assign \new_[35724]_  = \new_[35723]_  & \new_[35716]_ ;
  assign \new_[35728]_  = ~A167 & A168;
  assign \new_[35729]_  = A170 & \new_[35728]_ ;
  assign \new_[35732]_  = ~A232 & A166;
  assign \new_[35735]_  = ~A234 & A233;
  assign \new_[35736]_  = \new_[35735]_  & \new_[35732]_ ;
  assign \new_[35737]_  = \new_[35736]_  & \new_[35729]_ ;
  assign \new_[35740]_  = A236 & ~A235;
  assign \new_[35743]_  = A268 & ~A267;
  assign \new_[35744]_  = \new_[35743]_  & \new_[35740]_ ;
  assign \new_[35747]_  = A299 & ~A298;
  assign \new_[35750]_  = A301 & A300;
  assign \new_[35751]_  = \new_[35750]_  & \new_[35747]_ ;
  assign \new_[35752]_  = \new_[35751]_  & \new_[35744]_ ;
  assign \new_[35756]_  = ~A167 & A168;
  assign \new_[35757]_  = A170 & \new_[35756]_ ;
  assign \new_[35760]_  = ~A232 & A166;
  assign \new_[35763]_  = ~A234 & A233;
  assign \new_[35764]_  = \new_[35763]_  & \new_[35760]_ ;
  assign \new_[35765]_  = \new_[35764]_  & \new_[35757]_ ;
  assign \new_[35768]_  = A236 & ~A235;
  assign \new_[35771]_  = A268 & ~A267;
  assign \new_[35772]_  = \new_[35771]_  & \new_[35768]_ ;
  assign \new_[35775]_  = A299 & ~A298;
  assign \new_[35778]_  = ~A302 & A300;
  assign \new_[35779]_  = \new_[35778]_  & \new_[35775]_ ;
  assign \new_[35780]_  = \new_[35779]_  & \new_[35772]_ ;
  assign \new_[35784]_  = ~A167 & A168;
  assign \new_[35785]_  = A170 & \new_[35784]_ ;
  assign \new_[35788]_  = ~A232 & A166;
  assign \new_[35791]_  = ~A234 & A233;
  assign \new_[35792]_  = \new_[35791]_  & \new_[35788]_ ;
  assign \new_[35793]_  = \new_[35792]_  & \new_[35785]_ ;
  assign \new_[35796]_  = A236 & ~A235;
  assign \new_[35799]_  = ~A269 & ~A267;
  assign \new_[35800]_  = \new_[35799]_  & \new_[35796]_ ;
  assign \new_[35803]_  = ~A299 & A298;
  assign \new_[35806]_  = A301 & A300;
  assign \new_[35807]_  = \new_[35806]_  & \new_[35803]_ ;
  assign \new_[35808]_  = \new_[35807]_  & \new_[35800]_ ;
  assign \new_[35812]_  = ~A167 & A168;
  assign \new_[35813]_  = A170 & \new_[35812]_ ;
  assign \new_[35816]_  = ~A232 & A166;
  assign \new_[35819]_  = ~A234 & A233;
  assign \new_[35820]_  = \new_[35819]_  & \new_[35816]_ ;
  assign \new_[35821]_  = \new_[35820]_  & \new_[35813]_ ;
  assign \new_[35824]_  = A236 & ~A235;
  assign \new_[35827]_  = ~A269 & ~A267;
  assign \new_[35828]_  = \new_[35827]_  & \new_[35824]_ ;
  assign \new_[35831]_  = ~A299 & A298;
  assign \new_[35834]_  = ~A302 & A300;
  assign \new_[35835]_  = \new_[35834]_  & \new_[35831]_ ;
  assign \new_[35836]_  = \new_[35835]_  & \new_[35828]_ ;
  assign \new_[35840]_  = ~A167 & A168;
  assign \new_[35841]_  = A170 & \new_[35840]_ ;
  assign \new_[35844]_  = ~A232 & A166;
  assign \new_[35847]_  = ~A234 & A233;
  assign \new_[35848]_  = \new_[35847]_  & \new_[35844]_ ;
  assign \new_[35849]_  = \new_[35848]_  & \new_[35841]_ ;
  assign \new_[35852]_  = A236 & ~A235;
  assign \new_[35855]_  = ~A269 & ~A267;
  assign \new_[35856]_  = \new_[35855]_  & \new_[35852]_ ;
  assign \new_[35859]_  = A299 & ~A298;
  assign \new_[35862]_  = A301 & A300;
  assign \new_[35863]_  = \new_[35862]_  & \new_[35859]_ ;
  assign \new_[35864]_  = \new_[35863]_  & \new_[35856]_ ;
  assign \new_[35868]_  = ~A167 & A168;
  assign \new_[35869]_  = A170 & \new_[35868]_ ;
  assign \new_[35872]_  = ~A232 & A166;
  assign \new_[35875]_  = ~A234 & A233;
  assign \new_[35876]_  = \new_[35875]_  & \new_[35872]_ ;
  assign \new_[35877]_  = \new_[35876]_  & \new_[35869]_ ;
  assign \new_[35880]_  = A236 & ~A235;
  assign \new_[35883]_  = ~A269 & ~A267;
  assign \new_[35884]_  = \new_[35883]_  & \new_[35880]_ ;
  assign \new_[35887]_  = A299 & ~A298;
  assign \new_[35890]_  = ~A302 & A300;
  assign \new_[35891]_  = \new_[35890]_  & \new_[35887]_ ;
  assign \new_[35892]_  = \new_[35891]_  & \new_[35884]_ ;
  assign \new_[35896]_  = ~A167 & A168;
  assign \new_[35897]_  = A170 & \new_[35896]_ ;
  assign \new_[35900]_  = ~A232 & A166;
  assign \new_[35903]_  = ~A234 & A233;
  assign \new_[35904]_  = \new_[35903]_  & \new_[35900]_ ;
  assign \new_[35905]_  = \new_[35904]_  & \new_[35897]_ ;
  assign \new_[35908]_  = A236 & ~A235;
  assign \new_[35911]_  = A266 & A265;
  assign \new_[35912]_  = \new_[35911]_  & \new_[35908]_ ;
  assign \new_[35915]_  = ~A299 & A298;
  assign \new_[35918]_  = A301 & A300;
  assign \new_[35919]_  = \new_[35918]_  & \new_[35915]_ ;
  assign \new_[35920]_  = \new_[35919]_  & \new_[35912]_ ;
  assign \new_[35924]_  = ~A167 & A168;
  assign \new_[35925]_  = A170 & \new_[35924]_ ;
  assign \new_[35928]_  = ~A232 & A166;
  assign \new_[35931]_  = ~A234 & A233;
  assign \new_[35932]_  = \new_[35931]_  & \new_[35928]_ ;
  assign \new_[35933]_  = \new_[35932]_  & \new_[35925]_ ;
  assign \new_[35936]_  = A236 & ~A235;
  assign \new_[35939]_  = A266 & A265;
  assign \new_[35940]_  = \new_[35939]_  & \new_[35936]_ ;
  assign \new_[35943]_  = ~A299 & A298;
  assign \new_[35946]_  = ~A302 & A300;
  assign \new_[35947]_  = \new_[35946]_  & \new_[35943]_ ;
  assign \new_[35948]_  = \new_[35947]_  & \new_[35940]_ ;
  assign \new_[35952]_  = ~A167 & A168;
  assign \new_[35953]_  = A170 & \new_[35952]_ ;
  assign \new_[35956]_  = ~A232 & A166;
  assign \new_[35959]_  = ~A234 & A233;
  assign \new_[35960]_  = \new_[35959]_  & \new_[35956]_ ;
  assign \new_[35961]_  = \new_[35960]_  & \new_[35953]_ ;
  assign \new_[35964]_  = A236 & ~A235;
  assign \new_[35967]_  = A266 & A265;
  assign \new_[35968]_  = \new_[35967]_  & \new_[35964]_ ;
  assign \new_[35971]_  = A299 & ~A298;
  assign \new_[35974]_  = A301 & A300;
  assign \new_[35975]_  = \new_[35974]_  & \new_[35971]_ ;
  assign \new_[35976]_  = \new_[35975]_  & \new_[35968]_ ;
  assign \new_[35980]_  = ~A167 & A168;
  assign \new_[35981]_  = A170 & \new_[35980]_ ;
  assign \new_[35984]_  = ~A232 & A166;
  assign \new_[35987]_  = ~A234 & A233;
  assign \new_[35988]_  = \new_[35987]_  & \new_[35984]_ ;
  assign \new_[35989]_  = \new_[35988]_  & \new_[35981]_ ;
  assign \new_[35992]_  = A236 & ~A235;
  assign \new_[35995]_  = A266 & A265;
  assign \new_[35996]_  = \new_[35995]_  & \new_[35992]_ ;
  assign \new_[35999]_  = A299 & ~A298;
  assign \new_[36002]_  = ~A302 & A300;
  assign \new_[36003]_  = \new_[36002]_  & \new_[35999]_ ;
  assign \new_[36004]_  = \new_[36003]_  & \new_[35996]_ ;
  assign \new_[36008]_  = ~A167 & A168;
  assign \new_[36009]_  = A170 & \new_[36008]_ ;
  assign \new_[36012]_  = ~A232 & A166;
  assign \new_[36015]_  = ~A234 & A233;
  assign \new_[36016]_  = \new_[36015]_  & \new_[36012]_ ;
  assign \new_[36017]_  = \new_[36016]_  & \new_[36009]_ ;
  assign \new_[36020]_  = A236 & ~A235;
  assign \new_[36023]_  = ~A266 & ~A265;
  assign \new_[36024]_  = \new_[36023]_  & \new_[36020]_ ;
  assign \new_[36027]_  = ~A299 & A298;
  assign \new_[36030]_  = A301 & A300;
  assign \new_[36031]_  = \new_[36030]_  & \new_[36027]_ ;
  assign \new_[36032]_  = \new_[36031]_  & \new_[36024]_ ;
  assign \new_[36036]_  = ~A167 & A168;
  assign \new_[36037]_  = A170 & \new_[36036]_ ;
  assign \new_[36040]_  = ~A232 & A166;
  assign \new_[36043]_  = ~A234 & A233;
  assign \new_[36044]_  = \new_[36043]_  & \new_[36040]_ ;
  assign \new_[36045]_  = \new_[36044]_  & \new_[36037]_ ;
  assign \new_[36048]_  = A236 & ~A235;
  assign \new_[36051]_  = ~A266 & ~A265;
  assign \new_[36052]_  = \new_[36051]_  & \new_[36048]_ ;
  assign \new_[36055]_  = ~A299 & A298;
  assign \new_[36058]_  = ~A302 & A300;
  assign \new_[36059]_  = \new_[36058]_  & \new_[36055]_ ;
  assign \new_[36060]_  = \new_[36059]_  & \new_[36052]_ ;
  assign \new_[36064]_  = ~A167 & A168;
  assign \new_[36065]_  = A170 & \new_[36064]_ ;
  assign \new_[36068]_  = ~A232 & A166;
  assign \new_[36071]_  = ~A234 & A233;
  assign \new_[36072]_  = \new_[36071]_  & \new_[36068]_ ;
  assign \new_[36073]_  = \new_[36072]_  & \new_[36065]_ ;
  assign \new_[36076]_  = A236 & ~A235;
  assign \new_[36079]_  = ~A266 & ~A265;
  assign \new_[36080]_  = \new_[36079]_  & \new_[36076]_ ;
  assign \new_[36083]_  = A299 & ~A298;
  assign \new_[36086]_  = A301 & A300;
  assign \new_[36087]_  = \new_[36086]_  & \new_[36083]_ ;
  assign \new_[36088]_  = \new_[36087]_  & \new_[36080]_ ;
  assign \new_[36092]_  = ~A167 & A168;
  assign \new_[36093]_  = A170 & \new_[36092]_ ;
  assign \new_[36096]_  = ~A232 & A166;
  assign \new_[36099]_  = ~A234 & A233;
  assign \new_[36100]_  = \new_[36099]_  & \new_[36096]_ ;
  assign \new_[36101]_  = \new_[36100]_  & \new_[36093]_ ;
  assign \new_[36104]_  = A236 & ~A235;
  assign \new_[36107]_  = ~A266 & ~A265;
  assign \new_[36108]_  = \new_[36107]_  & \new_[36104]_ ;
  assign \new_[36111]_  = A299 & ~A298;
  assign \new_[36114]_  = ~A302 & A300;
  assign \new_[36115]_  = \new_[36114]_  & \new_[36111]_ ;
  assign \new_[36116]_  = \new_[36115]_  & \new_[36108]_ ;
  assign \new_[36120]_  = ~A167 & A168;
  assign \new_[36121]_  = A170 & \new_[36120]_ ;
  assign \new_[36124]_  = A232 & A166;
  assign \new_[36127]_  = A234 & ~A233;
  assign \new_[36128]_  = \new_[36127]_  & \new_[36124]_ ;
  assign \new_[36129]_  = \new_[36128]_  & \new_[36121]_ ;
  assign \new_[36132]_  = A267 & A235;
  assign \new_[36135]_  = A269 & ~A268;
  assign \new_[36136]_  = \new_[36135]_  & \new_[36132]_ ;
  assign \new_[36139]_  = ~A299 & A298;
  assign \new_[36142]_  = A301 & A300;
  assign \new_[36143]_  = \new_[36142]_  & \new_[36139]_ ;
  assign \new_[36144]_  = \new_[36143]_  & \new_[36136]_ ;
  assign \new_[36148]_  = ~A167 & A168;
  assign \new_[36149]_  = A170 & \new_[36148]_ ;
  assign \new_[36152]_  = A232 & A166;
  assign \new_[36155]_  = A234 & ~A233;
  assign \new_[36156]_  = \new_[36155]_  & \new_[36152]_ ;
  assign \new_[36157]_  = \new_[36156]_  & \new_[36149]_ ;
  assign \new_[36160]_  = A267 & A235;
  assign \new_[36163]_  = A269 & ~A268;
  assign \new_[36164]_  = \new_[36163]_  & \new_[36160]_ ;
  assign \new_[36167]_  = ~A299 & A298;
  assign \new_[36170]_  = ~A302 & A300;
  assign \new_[36171]_  = \new_[36170]_  & \new_[36167]_ ;
  assign \new_[36172]_  = \new_[36171]_  & \new_[36164]_ ;
  assign \new_[36176]_  = ~A167 & A168;
  assign \new_[36177]_  = A170 & \new_[36176]_ ;
  assign \new_[36180]_  = A232 & A166;
  assign \new_[36183]_  = A234 & ~A233;
  assign \new_[36184]_  = \new_[36183]_  & \new_[36180]_ ;
  assign \new_[36185]_  = \new_[36184]_  & \new_[36177]_ ;
  assign \new_[36188]_  = A267 & A235;
  assign \new_[36191]_  = A269 & ~A268;
  assign \new_[36192]_  = \new_[36191]_  & \new_[36188]_ ;
  assign \new_[36195]_  = A299 & ~A298;
  assign \new_[36198]_  = A301 & A300;
  assign \new_[36199]_  = \new_[36198]_  & \new_[36195]_ ;
  assign \new_[36200]_  = \new_[36199]_  & \new_[36192]_ ;
  assign \new_[36204]_  = ~A167 & A168;
  assign \new_[36205]_  = A170 & \new_[36204]_ ;
  assign \new_[36208]_  = A232 & A166;
  assign \new_[36211]_  = A234 & ~A233;
  assign \new_[36212]_  = \new_[36211]_  & \new_[36208]_ ;
  assign \new_[36213]_  = \new_[36212]_  & \new_[36205]_ ;
  assign \new_[36216]_  = A267 & A235;
  assign \new_[36219]_  = A269 & ~A268;
  assign \new_[36220]_  = \new_[36219]_  & \new_[36216]_ ;
  assign \new_[36223]_  = A299 & ~A298;
  assign \new_[36226]_  = ~A302 & A300;
  assign \new_[36227]_  = \new_[36226]_  & \new_[36223]_ ;
  assign \new_[36228]_  = \new_[36227]_  & \new_[36220]_ ;
  assign \new_[36232]_  = ~A167 & A168;
  assign \new_[36233]_  = A170 & \new_[36232]_ ;
  assign \new_[36236]_  = A232 & A166;
  assign \new_[36239]_  = A234 & ~A233;
  assign \new_[36240]_  = \new_[36239]_  & \new_[36236]_ ;
  assign \new_[36241]_  = \new_[36240]_  & \new_[36233]_ ;
  assign \new_[36244]_  = ~A267 & A235;
  assign \new_[36247]_  = A298 & A268;
  assign \new_[36248]_  = \new_[36247]_  & \new_[36244]_ ;
  assign \new_[36251]_  = ~A300 & ~A299;
  assign \new_[36254]_  = A302 & ~A301;
  assign \new_[36255]_  = \new_[36254]_  & \new_[36251]_ ;
  assign \new_[36256]_  = \new_[36255]_  & \new_[36248]_ ;
  assign \new_[36260]_  = ~A167 & A168;
  assign \new_[36261]_  = A170 & \new_[36260]_ ;
  assign \new_[36264]_  = A232 & A166;
  assign \new_[36267]_  = A234 & ~A233;
  assign \new_[36268]_  = \new_[36267]_  & \new_[36264]_ ;
  assign \new_[36269]_  = \new_[36268]_  & \new_[36261]_ ;
  assign \new_[36272]_  = ~A267 & A235;
  assign \new_[36275]_  = ~A298 & A268;
  assign \new_[36276]_  = \new_[36275]_  & \new_[36272]_ ;
  assign \new_[36279]_  = ~A300 & A299;
  assign \new_[36282]_  = A302 & ~A301;
  assign \new_[36283]_  = \new_[36282]_  & \new_[36279]_ ;
  assign \new_[36284]_  = \new_[36283]_  & \new_[36276]_ ;
  assign \new_[36288]_  = ~A167 & A168;
  assign \new_[36289]_  = A170 & \new_[36288]_ ;
  assign \new_[36292]_  = A232 & A166;
  assign \new_[36295]_  = A234 & ~A233;
  assign \new_[36296]_  = \new_[36295]_  & \new_[36292]_ ;
  assign \new_[36297]_  = \new_[36296]_  & \new_[36289]_ ;
  assign \new_[36300]_  = ~A267 & A235;
  assign \new_[36303]_  = A298 & ~A269;
  assign \new_[36304]_  = \new_[36303]_  & \new_[36300]_ ;
  assign \new_[36307]_  = ~A300 & ~A299;
  assign \new_[36310]_  = A302 & ~A301;
  assign \new_[36311]_  = \new_[36310]_  & \new_[36307]_ ;
  assign \new_[36312]_  = \new_[36311]_  & \new_[36304]_ ;
  assign \new_[36316]_  = ~A167 & A168;
  assign \new_[36317]_  = A170 & \new_[36316]_ ;
  assign \new_[36320]_  = A232 & A166;
  assign \new_[36323]_  = A234 & ~A233;
  assign \new_[36324]_  = \new_[36323]_  & \new_[36320]_ ;
  assign \new_[36325]_  = \new_[36324]_  & \new_[36317]_ ;
  assign \new_[36328]_  = ~A267 & A235;
  assign \new_[36331]_  = ~A298 & ~A269;
  assign \new_[36332]_  = \new_[36331]_  & \new_[36328]_ ;
  assign \new_[36335]_  = ~A300 & A299;
  assign \new_[36338]_  = A302 & ~A301;
  assign \new_[36339]_  = \new_[36338]_  & \new_[36335]_ ;
  assign \new_[36340]_  = \new_[36339]_  & \new_[36332]_ ;
  assign \new_[36344]_  = ~A167 & A168;
  assign \new_[36345]_  = A170 & \new_[36344]_ ;
  assign \new_[36348]_  = A232 & A166;
  assign \new_[36351]_  = A234 & ~A233;
  assign \new_[36352]_  = \new_[36351]_  & \new_[36348]_ ;
  assign \new_[36353]_  = \new_[36352]_  & \new_[36345]_ ;
  assign \new_[36356]_  = A265 & A235;
  assign \new_[36359]_  = A298 & A266;
  assign \new_[36360]_  = \new_[36359]_  & \new_[36356]_ ;
  assign \new_[36363]_  = ~A300 & ~A299;
  assign \new_[36366]_  = A302 & ~A301;
  assign \new_[36367]_  = \new_[36366]_  & \new_[36363]_ ;
  assign \new_[36368]_  = \new_[36367]_  & \new_[36360]_ ;
  assign \new_[36372]_  = ~A167 & A168;
  assign \new_[36373]_  = A170 & \new_[36372]_ ;
  assign \new_[36376]_  = A232 & A166;
  assign \new_[36379]_  = A234 & ~A233;
  assign \new_[36380]_  = \new_[36379]_  & \new_[36376]_ ;
  assign \new_[36381]_  = \new_[36380]_  & \new_[36373]_ ;
  assign \new_[36384]_  = A265 & A235;
  assign \new_[36387]_  = ~A298 & A266;
  assign \new_[36388]_  = \new_[36387]_  & \new_[36384]_ ;
  assign \new_[36391]_  = ~A300 & A299;
  assign \new_[36394]_  = A302 & ~A301;
  assign \new_[36395]_  = \new_[36394]_  & \new_[36391]_ ;
  assign \new_[36396]_  = \new_[36395]_  & \new_[36388]_ ;
  assign \new_[36400]_  = ~A167 & A168;
  assign \new_[36401]_  = A170 & \new_[36400]_ ;
  assign \new_[36404]_  = A232 & A166;
  assign \new_[36407]_  = A234 & ~A233;
  assign \new_[36408]_  = \new_[36407]_  & \new_[36404]_ ;
  assign \new_[36409]_  = \new_[36408]_  & \new_[36401]_ ;
  assign \new_[36412]_  = ~A265 & A235;
  assign \new_[36415]_  = A298 & ~A266;
  assign \new_[36416]_  = \new_[36415]_  & \new_[36412]_ ;
  assign \new_[36419]_  = ~A300 & ~A299;
  assign \new_[36422]_  = A302 & ~A301;
  assign \new_[36423]_  = \new_[36422]_  & \new_[36419]_ ;
  assign \new_[36424]_  = \new_[36423]_  & \new_[36416]_ ;
  assign \new_[36428]_  = ~A167 & A168;
  assign \new_[36429]_  = A170 & \new_[36428]_ ;
  assign \new_[36432]_  = A232 & A166;
  assign \new_[36435]_  = A234 & ~A233;
  assign \new_[36436]_  = \new_[36435]_  & \new_[36432]_ ;
  assign \new_[36437]_  = \new_[36436]_  & \new_[36429]_ ;
  assign \new_[36440]_  = ~A265 & A235;
  assign \new_[36443]_  = ~A298 & ~A266;
  assign \new_[36444]_  = \new_[36443]_  & \new_[36440]_ ;
  assign \new_[36447]_  = ~A300 & A299;
  assign \new_[36450]_  = A302 & ~A301;
  assign \new_[36451]_  = \new_[36450]_  & \new_[36447]_ ;
  assign \new_[36452]_  = \new_[36451]_  & \new_[36444]_ ;
  assign \new_[36456]_  = ~A167 & A168;
  assign \new_[36457]_  = A170 & \new_[36456]_ ;
  assign \new_[36460]_  = A232 & A166;
  assign \new_[36463]_  = A234 & ~A233;
  assign \new_[36464]_  = \new_[36463]_  & \new_[36460]_ ;
  assign \new_[36465]_  = \new_[36464]_  & \new_[36457]_ ;
  assign \new_[36468]_  = A267 & ~A236;
  assign \new_[36471]_  = A269 & ~A268;
  assign \new_[36472]_  = \new_[36471]_  & \new_[36468]_ ;
  assign \new_[36475]_  = ~A299 & A298;
  assign \new_[36478]_  = A301 & A300;
  assign \new_[36479]_  = \new_[36478]_  & \new_[36475]_ ;
  assign \new_[36480]_  = \new_[36479]_  & \new_[36472]_ ;
  assign \new_[36484]_  = ~A167 & A168;
  assign \new_[36485]_  = A170 & \new_[36484]_ ;
  assign \new_[36488]_  = A232 & A166;
  assign \new_[36491]_  = A234 & ~A233;
  assign \new_[36492]_  = \new_[36491]_  & \new_[36488]_ ;
  assign \new_[36493]_  = \new_[36492]_  & \new_[36485]_ ;
  assign \new_[36496]_  = A267 & ~A236;
  assign \new_[36499]_  = A269 & ~A268;
  assign \new_[36500]_  = \new_[36499]_  & \new_[36496]_ ;
  assign \new_[36503]_  = ~A299 & A298;
  assign \new_[36506]_  = ~A302 & A300;
  assign \new_[36507]_  = \new_[36506]_  & \new_[36503]_ ;
  assign \new_[36508]_  = \new_[36507]_  & \new_[36500]_ ;
  assign \new_[36512]_  = ~A167 & A168;
  assign \new_[36513]_  = A170 & \new_[36512]_ ;
  assign \new_[36516]_  = A232 & A166;
  assign \new_[36519]_  = A234 & ~A233;
  assign \new_[36520]_  = \new_[36519]_  & \new_[36516]_ ;
  assign \new_[36521]_  = \new_[36520]_  & \new_[36513]_ ;
  assign \new_[36524]_  = A267 & ~A236;
  assign \new_[36527]_  = A269 & ~A268;
  assign \new_[36528]_  = \new_[36527]_  & \new_[36524]_ ;
  assign \new_[36531]_  = A299 & ~A298;
  assign \new_[36534]_  = A301 & A300;
  assign \new_[36535]_  = \new_[36534]_  & \new_[36531]_ ;
  assign \new_[36536]_  = \new_[36535]_  & \new_[36528]_ ;
  assign \new_[36540]_  = ~A167 & A168;
  assign \new_[36541]_  = A170 & \new_[36540]_ ;
  assign \new_[36544]_  = A232 & A166;
  assign \new_[36547]_  = A234 & ~A233;
  assign \new_[36548]_  = \new_[36547]_  & \new_[36544]_ ;
  assign \new_[36549]_  = \new_[36548]_  & \new_[36541]_ ;
  assign \new_[36552]_  = A267 & ~A236;
  assign \new_[36555]_  = A269 & ~A268;
  assign \new_[36556]_  = \new_[36555]_  & \new_[36552]_ ;
  assign \new_[36559]_  = A299 & ~A298;
  assign \new_[36562]_  = ~A302 & A300;
  assign \new_[36563]_  = \new_[36562]_  & \new_[36559]_ ;
  assign \new_[36564]_  = \new_[36563]_  & \new_[36556]_ ;
  assign \new_[36568]_  = ~A167 & A168;
  assign \new_[36569]_  = A170 & \new_[36568]_ ;
  assign \new_[36572]_  = A232 & A166;
  assign \new_[36575]_  = A234 & ~A233;
  assign \new_[36576]_  = \new_[36575]_  & \new_[36572]_ ;
  assign \new_[36577]_  = \new_[36576]_  & \new_[36569]_ ;
  assign \new_[36580]_  = ~A267 & ~A236;
  assign \new_[36583]_  = A298 & A268;
  assign \new_[36584]_  = \new_[36583]_  & \new_[36580]_ ;
  assign \new_[36587]_  = ~A300 & ~A299;
  assign \new_[36590]_  = A302 & ~A301;
  assign \new_[36591]_  = \new_[36590]_  & \new_[36587]_ ;
  assign \new_[36592]_  = \new_[36591]_  & \new_[36584]_ ;
  assign \new_[36596]_  = ~A167 & A168;
  assign \new_[36597]_  = A170 & \new_[36596]_ ;
  assign \new_[36600]_  = A232 & A166;
  assign \new_[36603]_  = A234 & ~A233;
  assign \new_[36604]_  = \new_[36603]_  & \new_[36600]_ ;
  assign \new_[36605]_  = \new_[36604]_  & \new_[36597]_ ;
  assign \new_[36608]_  = ~A267 & ~A236;
  assign \new_[36611]_  = ~A298 & A268;
  assign \new_[36612]_  = \new_[36611]_  & \new_[36608]_ ;
  assign \new_[36615]_  = ~A300 & A299;
  assign \new_[36618]_  = A302 & ~A301;
  assign \new_[36619]_  = \new_[36618]_  & \new_[36615]_ ;
  assign \new_[36620]_  = \new_[36619]_  & \new_[36612]_ ;
  assign \new_[36624]_  = ~A167 & A168;
  assign \new_[36625]_  = A170 & \new_[36624]_ ;
  assign \new_[36628]_  = A232 & A166;
  assign \new_[36631]_  = A234 & ~A233;
  assign \new_[36632]_  = \new_[36631]_  & \new_[36628]_ ;
  assign \new_[36633]_  = \new_[36632]_  & \new_[36625]_ ;
  assign \new_[36636]_  = ~A267 & ~A236;
  assign \new_[36639]_  = A298 & ~A269;
  assign \new_[36640]_  = \new_[36639]_  & \new_[36636]_ ;
  assign \new_[36643]_  = ~A300 & ~A299;
  assign \new_[36646]_  = A302 & ~A301;
  assign \new_[36647]_  = \new_[36646]_  & \new_[36643]_ ;
  assign \new_[36648]_  = \new_[36647]_  & \new_[36640]_ ;
  assign \new_[36652]_  = ~A167 & A168;
  assign \new_[36653]_  = A170 & \new_[36652]_ ;
  assign \new_[36656]_  = A232 & A166;
  assign \new_[36659]_  = A234 & ~A233;
  assign \new_[36660]_  = \new_[36659]_  & \new_[36656]_ ;
  assign \new_[36661]_  = \new_[36660]_  & \new_[36653]_ ;
  assign \new_[36664]_  = ~A267 & ~A236;
  assign \new_[36667]_  = ~A298 & ~A269;
  assign \new_[36668]_  = \new_[36667]_  & \new_[36664]_ ;
  assign \new_[36671]_  = ~A300 & A299;
  assign \new_[36674]_  = A302 & ~A301;
  assign \new_[36675]_  = \new_[36674]_  & \new_[36671]_ ;
  assign \new_[36676]_  = \new_[36675]_  & \new_[36668]_ ;
  assign \new_[36680]_  = ~A167 & A168;
  assign \new_[36681]_  = A170 & \new_[36680]_ ;
  assign \new_[36684]_  = A232 & A166;
  assign \new_[36687]_  = A234 & ~A233;
  assign \new_[36688]_  = \new_[36687]_  & \new_[36684]_ ;
  assign \new_[36689]_  = \new_[36688]_  & \new_[36681]_ ;
  assign \new_[36692]_  = A265 & ~A236;
  assign \new_[36695]_  = A298 & A266;
  assign \new_[36696]_  = \new_[36695]_  & \new_[36692]_ ;
  assign \new_[36699]_  = ~A300 & ~A299;
  assign \new_[36702]_  = A302 & ~A301;
  assign \new_[36703]_  = \new_[36702]_  & \new_[36699]_ ;
  assign \new_[36704]_  = \new_[36703]_  & \new_[36696]_ ;
  assign \new_[36708]_  = ~A167 & A168;
  assign \new_[36709]_  = A170 & \new_[36708]_ ;
  assign \new_[36712]_  = A232 & A166;
  assign \new_[36715]_  = A234 & ~A233;
  assign \new_[36716]_  = \new_[36715]_  & \new_[36712]_ ;
  assign \new_[36717]_  = \new_[36716]_  & \new_[36709]_ ;
  assign \new_[36720]_  = A265 & ~A236;
  assign \new_[36723]_  = ~A298 & A266;
  assign \new_[36724]_  = \new_[36723]_  & \new_[36720]_ ;
  assign \new_[36727]_  = ~A300 & A299;
  assign \new_[36730]_  = A302 & ~A301;
  assign \new_[36731]_  = \new_[36730]_  & \new_[36727]_ ;
  assign \new_[36732]_  = \new_[36731]_  & \new_[36724]_ ;
  assign \new_[36736]_  = ~A167 & A168;
  assign \new_[36737]_  = A170 & \new_[36736]_ ;
  assign \new_[36740]_  = A232 & A166;
  assign \new_[36743]_  = A234 & ~A233;
  assign \new_[36744]_  = \new_[36743]_  & \new_[36740]_ ;
  assign \new_[36745]_  = \new_[36744]_  & \new_[36737]_ ;
  assign \new_[36748]_  = ~A265 & ~A236;
  assign \new_[36751]_  = A298 & ~A266;
  assign \new_[36752]_  = \new_[36751]_  & \new_[36748]_ ;
  assign \new_[36755]_  = ~A300 & ~A299;
  assign \new_[36758]_  = A302 & ~A301;
  assign \new_[36759]_  = \new_[36758]_  & \new_[36755]_ ;
  assign \new_[36760]_  = \new_[36759]_  & \new_[36752]_ ;
  assign \new_[36764]_  = ~A167 & A168;
  assign \new_[36765]_  = A170 & \new_[36764]_ ;
  assign \new_[36768]_  = A232 & A166;
  assign \new_[36771]_  = A234 & ~A233;
  assign \new_[36772]_  = \new_[36771]_  & \new_[36768]_ ;
  assign \new_[36773]_  = \new_[36772]_  & \new_[36765]_ ;
  assign \new_[36776]_  = ~A265 & ~A236;
  assign \new_[36779]_  = ~A298 & ~A266;
  assign \new_[36780]_  = \new_[36779]_  & \new_[36776]_ ;
  assign \new_[36783]_  = ~A300 & A299;
  assign \new_[36786]_  = A302 & ~A301;
  assign \new_[36787]_  = \new_[36786]_  & \new_[36783]_ ;
  assign \new_[36788]_  = \new_[36787]_  & \new_[36780]_ ;
  assign \new_[36792]_  = ~A167 & A168;
  assign \new_[36793]_  = A170 & \new_[36792]_ ;
  assign \new_[36796]_  = A232 & A166;
  assign \new_[36799]_  = ~A234 & ~A233;
  assign \new_[36800]_  = \new_[36799]_  & \new_[36796]_ ;
  assign \new_[36801]_  = \new_[36800]_  & \new_[36793]_ ;
  assign \new_[36804]_  = A236 & ~A235;
  assign \new_[36807]_  = A268 & ~A267;
  assign \new_[36808]_  = \new_[36807]_  & \new_[36804]_ ;
  assign \new_[36811]_  = ~A299 & A298;
  assign \new_[36814]_  = A301 & A300;
  assign \new_[36815]_  = \new_[36814]_  & \new_[36811]_ ;
  assign \new_[36816]_  = \new_[36815]_  & \new_[36808]_ ;
  assign \new_[36820]_  = ~A167 & A168;
  assign \new_[36821]_  = A170 & \new_[36820]_ ;
  assign \new_[36824]_  = A232 & A166;
  assign \new_[36827]_  = ~A234 & ~A233;
  assign \new_[36828]_  = \new_[36827]_  & \new_[36824]_ ;
  assign \new_[36829]_  = \new_[36828]_  & \new_[36821]_ ;
  assign \new_[36832]_  = A236 & ~A235;
  assign \new_[36835]_  = A268 & ~A267;
  assign \new_[36836]_  = \new_[36835]_  & \new_[36832]_ ;
  assign \new_[36839]_  = ~A299 & A298;
  assign \new_[36842]_  = ~A302 & A300;
  assign \new_[36843]_  = \new_[36842]_  & \new_[36839]_ ;
  assign \new_[36844]_  = \new_[36843]_  & \new_[36836]_ ;
  assign \new_[36848]_  = ~A167 & A168;
  assign \new_[36849]_  = A170 & \new_[36848]_ ;
  assign \new_[36852]_  = A232 & A166;
  assign \new_[36855]_  = ~A234 & ~A233;
  assign \new_[36856]_  = \new_[36855]_  & \new_[36852]_ ;
  assign \new_[36857]_  = \new_[36856]_  & \new_[36849]_ ;
  assign \new_[36860]_  = A236 & ~A235;
  assign \new_[36863]_  = A268 & ~A267;
  assign \new_[36864]_  = \new_[36863]_  & \new_[36860]_ ;
  assign \new_[36867]_  = A299 & ~A298;
  assign \new_[36870]_  = A301 & A300;
  assign \new_[36871]_  = \new_[36870]_  & \new_[36867]_ ;
  assign \new_[36872]_  = \new_[36871]_  & \new_[36864]_ ;
  assign \new_[36876]_  = ~A167 & A168;
  assign \new_[36877]_  = A170 & \new_[36876]_ ;
  assign \new_[36880]_  = A232 & A166;
  assign \new_[36883]_  = ~A234 & ~A233;
  assign \new_[36884]_  = \new_[36883]_  & \new_[36880]_ ;
  assign \new_[36885]_  = \new_[36884]_  & \new_[36877]_ ;
  assign \new_[36888]_  = A236 & ~A235;
  assign \new_[36891]_  = A268 & ~A267;
  assign \new_[36892]_  = \new_[36891]_  & \new_[36888]_ ;
  assign \new_[36895]_  = A299 & ~A298;
  assign \new_[36898]_  = ~A302 & A300;
  assign \new_[36899]_  = \new_[36898]_  & \new_[36895]_ ;
  assign \new_[36900]_  = \new_[36899]_  & \new_[36892]_ ;
  assign \new_[36904]_  = ~A167 & A168;
  assign \new_[36905]_  = A170 & \new_[36904]_ ;
  assign \new_[36908]_  = A232 & A166;
  assign \new_[36911]_  = ~A234 & ~A233;
  assign \new_[36912]_  = \new_[36911]_  & \new_[36908]_ ;
  assign \new_[36913]_  = \new_[36912]_  & \new_[36905]_ ;
  assign \new_[36916]_  = A236 & ~A235;
  assign \new_[36919]_  = ~A269 & ~A267;
  assign \new_[36920]_  = \new_[36919]_  & \new_[36916]_ ;
  assign \new_[36923]_  = ~A299 & A298;
  assign \new_[36926]_  = A301 & A300;
  assign \new_[36927]_  = \new_[36926]_  & \new_[36923]_ ;
  assign \new_[36928]_  = \new_[36927]_  & \new_[36920]_ ;
  assign \new_[36932]_  = ~A167 & A168;
  assign \new_[36933]_  = A170 & \new_[36932]_ ;
  assign \new_[36936]_  = A232 & A166;
  assign \new_[36939]_  = ~A234 & ~A233;
  assign \new_[36940]_  = \new_[36939]_  & \new_[36936]_ ;
  assign \new_[36941]_  = \new_[36940]_  & \new_[36933]_ ;
  assign \new_[36944]_  = A236 & ~A235;
  assign \new_[36947]_  = ~A269 & ~A267;
  assign \new_[36948]_  = \new_[36947]_  & \new_[36944]_ ;
  assign \new_[36951]_  = ~A299 & A298;
  assign \new_[36954]_  = ~A302 & A300;
  assign \new_[36955]_  = \new_[36954]_  & \new_[36951]_ ;
  assign \new_[36956]_  = \new_[36955]_  & \new_[36948]_ ;
  assign \new_[36960]_  = ~A167 & A168;
  assign \new_[36961]_  = A170 & \new_[36960]_ ;
  assign \new_[36964]_  = A232 & A166;
  assign \new_[36967]_  = ~A234 & ~A233;
  assign \new_[36968]_  = \new_[36967]_  & \new_[36964]_ ;
  assign \new_[36969]_  = \new_[36968]_  & \new_[36961]_ ;
  assign \new_[36972]_  = A236 & ~A235;
  assign \new_[36975]_  = ~A269 & ~A267;
  assign \new_[36976]_  = \new_[36975]_  & \new_[36972]_ ;
  assign \new_[36979]_  = A299 & ~A298;
  assign \new_[36982]_  = A301 & A300;
  assign \new_[36983]_  = \new_[36982]_  & \new_[36979]_ ;
  assign \new_[36984]_  = \new_[36983]_  & \new_[36976]_ ;
  assign \new_[36988]_  = ~A167 & A168;
  assign \new_[36989]_  = A170 & \new_[36988]_ ;
  assign \new_[36992]_  = A232 & A166;
  assign \new_[36995]_  = ~A234 & ~A233;
  assign \new_[36996]_  = \new_[36995]_  & \new_[36992]_ ;
  assign \new_[36997]_  = \new_[36996]_  & \new_[36989]_ ;
  assign \new_[37000]_  = A236 & ~A235;
  assign \new_[37003]_  = ~A269 & ~A267;
  assign \new_[37004]_  = \new_[37003]_  & \new_[37000]_ ;
  assign \new_[37007]_  = A299 & ~A298;
  assign \new_[37010]_  = ~A302 & A300;
  assign \new_[37011]_  = \new_[37010]_  & \new_[37007]_ ;
  assign \new_[37012]_  = \new_[37011]_  & \new_[37004]_ ;
  assign \new_[37016]_  = ~A167 & A168;
  assign \new_[37017]_  = A170 & \new_[37016]_ ;
  assign \new_[37020]_  = A232 & A166;
  assign \new_[37023]_  = ~A234 & ~A233;
  assign \new_[37024]_  = \new_[37023]_  & \new_[37020]_ ;
  assign \new_[37025]_  = \new_[37024]_  & \new_[37017]_ ;
  assign \new_[37028]_  = A236 & ~A235;
  assign \new_[37031]_  = A266 & A265;
  assign \new_[37032]_  = \new_[37031]_  & \new_[37028]_ ;
  assign \new_[37035]_  = ~A299 & A298;
  assign \new_[37038]_  = A301 & A300;
  assign \new_[37039]_  = \new_[37038]_  & \new_[37035]_ ;
  assign \new_[37040]_  = \new_[37039]_  & \new_[37032]_ ;
  assign \new_[37044]_  = ~A167 & A168;
  assign \new_[37045]_  = A170 & \new_[37044]_ ;
  assign \new_[37048]_  = A232 & A166;
  assign \new_[37051]_  = ~A234 & ~A233;
  assign \new_[37052]_  = \new_[37051]_  & \new_[37048]_ ;
  assign \new_[37053]_  = \new_[37052]_  & \new_[37045]_ ;
  assign \new_[37056]_  = A236 & ~A235;
  assign \new_[37059]_  = A266 & A265;
  assign \new_[37060]_  = \new_[37059]_  & \new_[37056]_ ;
  assign \new_[37063]_  = ~A299 & A298;
  assign \new_[37066]_  = ~A302 & A300;
  assign \new_[37067]_  = \new_[37066]_  & \new_[37063]_ ;
  assign \new_[37068]_  = \new_[37067]_  & \new_[37060]_ ;
  assign \new_[37072]_  = ~A167 & A168;
  assign \new_[37073]_  = A170 & \new_[37072]_ ;
  assign \new_[37076]_  = A232 & A166;
  assign \new_[37079]_  = ~A234 & ~A233;
  assign \new_[37080]_  = \new_[37079]_  & \new_[37076]_ ;
  assign \new_[37081]_  = \new_[37080]_  & \new_[37073]_ ;
  assign \new_[37084]_  = A236 & ~A235;
  assign \new_[37087]_  = A266 & A265;
  assign \new_[37088]_  = \new_[37087]_  & \new_[37084]_ ;
  assign \new_[37091]_  = A299 & ~A298;
  assign \new_[37094]_  = A301 & A300;
  assign \new_[37095]_  = \new_[37094]_  & \new_[37091]_ ;
  assign \new_[37096]_  = \new_[37095]_  & \new_[37088]_ ;
  assign \new_[37100]_  = ~A167 & A168;
  assign \new_[37101]_  = A170 & \new_[37100]_ ;
  assign \new_[37104]_  = A232 & A166;
  assign \new_[37107]_  = ~A234 & ~A233;
  assign \new_[37108]_  = \new_[37107]_  & \new_[37104]_ ;
  assign \new_[37109]_  = \new_[37108]_  & \new_[37101]_ ;
  assign \new_[37112]_  = A236 & ~A235;
  assign \new_[37115]_  = A266 & A265;
  assign \new_[37116]_  = \new_[37115]_  & \new_[37112]_ ;
  assign \new_[37119]_  = A299 & ~A298;
  assign \new_[37122]_  = ~A302 & A300;
  assign \new_[37123]_  = \new_[37122]_  & \new_[37119]_ ;
  assign \new_[37124]_  = \new_[37123]_  & \new_[37116]_ ;
  assign \new_[37128]_  = ~A167 & A168;
  assign \new_[37129]_  = A170 & \new_[37128]_ ;
  assign \new_[37132]_  = A232 & A166;
  assign \new_[37135]_  = ~A234 & ~A233;
  assign \new_[37136]_  = \new_[37135]_  & \new_[37132]_ ;
  assign \new_[37137]_  = \new_[37136]_  & \new_[37129]_ ;
  assign \new_[37140]_  = A236 & ~A235;
  assign \new_[37143]_  = ~A266 & ~A265;
  assign \new_[37144]_  = \new_[37143]_  & \new_[37140]_ ;
  assign \new_[37147]_  = ~A299 & A298;
  assign \new_[37150]_  = A301 & A300;
  assign \new_[37151]_  = \new_[37150]_  & \new_[37147]_ ;
  assign \new_[37152]_  = \new_[37151]_  & \new_[37144]_ ;
  assign \new_[37156]_  = ~A167 & A168;
  assign \new_[37157]_  = A170 & \new_[37156]_ ;
  assign \new_[37160]_  = A232 & A166;
  assign \new_[37163]_  = ~A234 & ~A233;
  assign \new_[37164]_  = \new_[37163]_  & \new_[37160]_ ;
  assign \new_[37165]_  = \new_[37164]_  & \new_[37157]_ ;
  assign \new_[37168]_  = A236 & ~A235;
  assign \new_[37171]_  = ~A266 & ~A265;
  assign \new_[37172]_  = \new_[37171]_  & \new_[37168]_ ;
  assign \new_[37175]_  = ~A299 & A298;
  assign \new_[37178]_  = ~A302 & A300;
  assign \new_[37179]_  = \new_[37178]_  & \new_[37175]_ ;
  assign \new_[37180]_  = \new_[37179]_  & \new_[37172]_ ;
  assign \new_[37184]_  = ~A167 & A168;
  assign \new_[37185]_  = A170 & \new_[37184]_ ;
  assign \new_[37188]_  = A232 & A166;
  assign \new_[37191]_  = ~A234 & ~A233;
  assign \new_[37192]_  = \new_[37191]_  & \new_[37188]_ ;
  assign \new_[37193]_  = \new_[37192]_  & \new_[37185]_ ;
  assign \new_[37196]_  = A236 & ~A235;
  assign \new_[37199]_  = ~A266 & ~A265;
  assign \new_[37200]_  = \new_[37199]_  & \new_[37196]_ ;
  assign \new_[37203]_  = A299 & ~A298;
  assign \new_[37206]_  = A301 & A300;
  assign \new_[37207]_  = \new_[37206]_  & \new_[37203]_ ;
  assign \new_[37208]_  = \new_[37207]_  & \new_[37200]_ ;
  assign \new_[37212]_  = ~A167 & A168;
  assign \new_[37213]_  = A170 & \new_[37212]_ ;
  assign \new_[37216]_  = A232 & A166;
  assign \new_[37219]_  = ~A234 & ~A233;
  assign \new_[37220]_  = \new_[37219]_  & \new_[37216]_ ;
  assign \new_[37221]_  = \new_[37220]_  & \new_[37213]_ ;
  assign \new_[37224]_  = A236 & ~A235;
  assign \new_[37227]_  = ~A266 & ~A265;
  assign \new_[37228]_  = \new_[37227]_  & \new_[37224]_ ;
  assign \new_[37231]_  = A299 & ~A298;
  assign \new_[37234]_  = ~A302 & A300;
  assign \new_[37235]_  = \new_[37234]_  & \new_[37231]_ ;
  assign \new_[37236]_  = \new_[37235]_  & \new_[37228]_ ;
  assign \new_[37240]_  = A167 & A168;
  assign \new_[37241]_  = A169 & \new_[37240]_ ;
  assign \new_[37244]_  = ~A232 & ~A166;
  assign \new_[37247]_  = A234 & A233;
  assign \new_[37248]_  = \new_[37247]_  & \new_[37244]_ ;
  assign \new_[37249]_  = \new_[37248]_  & \new_[37241]_ ;
  assign \new_[37252]_  = A267 & A235;
  assign \new_[37255]_  = A269 & ~A268;
  assign \new_[37256]_  = \new_[37255]_  & \new_[37252]_ ;
  assign \new_[37259]_  = ~A299 & A298;
  assign \new_[37262]_  = A301 & A300;
  assign \new_[37263]_  = \new_[37262]_  & \new_[37259]_ ;
  assign \new_[37264]_  = \new_[37263]_  & \new_[37256]_ ;
  assign \new_[37268]_  = A167 & A168;
  assign \new_[37269]_  = A169 & \new_[37268]_ ;
  assign \new_[37272]_  = ~A232 & ~A166;
  assign \new_[37275]_  = A234 & A233;
  assign \new_[37276]_  = \new_[37275]_  & \new_[37272]_ ;
  assign \new_[37277]_  = \new_[37276]_  & \new_[37269]_ ;
  assign \new_[37280]_  = A267 & A235;
  assign \new_[37283]_  = A269 & ~A268;
  assign \new_[37284]_  = \new_[37283]_  & \new_[37280]_ ;
  assign \new_[37287]_  = ~A299 & A298;
  assign \new_[37290]_  = ~A302 & A300;
  assign \new_[37291]_  = \new_[37290]_  & \new_[37287]_ ;
  assign \new_[37292]_  = \new_[37291]_  & \new_[37284]_ ;
  assign \new_[37296]_  = A167 & A168;
  assign \new_[37297]_  = A169 & \new_[37296]_ ;
  assign \new_[37300]_  = ~A232 & ~A166;
  assign \new_[37303]_  = A234 & A233;
  assign \new_[37304]_  = \new_[37303]_  & \new_[37300]_ ;
  assign \new_[37305]_  = \new_[37304]_  & \new_[37297]_ ;
  assign \new_[37308]_  = A267 & A235;
  assign \new_[37311]_  = A269 & ~A268;
  assign \new_[37312]_  = \new_[37311]_  & \new_[37308]_ ;
  assign \new_[37315]_  = A299 & ~A298;
  assign \new_[37318]_  = A301 & A300;
  assign \new_[37319]_  = \new_[37318]_  & \new_[37315]_ ;
  assign \new_[37320]_  = \new_[37319]_  & \new_[37312]_ ;
  assign \new_[37324]_  = A167 & A168;
  assign \new_[37325]_  = A169 & \new_[37324]_ ;
  assign \new_[37328]_  = ~A232 & ~A166;
  assign \new_[37331]_  = A234 & A233;
  assign \new_[37332]_  = \new_[37331]_  & \new_[37328]_ ;
  assign \new_[37333]_  = \new_[37332]_  & \new_[37325]_ ;
  assign \new_[37336]_  = A267 & A235;
  assign \new_[37339]_  = A269 & ~A268;
  assign \new_[37340]_  = \new_[37339]_  & \new_[37336]_ ;
  assign \new_[37343]_  = A299 & ~A298;
  assign \new_[37346]_  = ~A302 & A300;
  assign \new_[37347]_  = \new_[37346]_  & \new_[37343]_ ;
  assign \new_[37348]_  = \new_[37347]_  & \new_[37340]_ ;
  assign \new_[37352]_  = A167 & A168;
  assign \new_[37353]_  = A169 & \new_[37352]_ ;
  assign \new_[37356]_  = ~A232 & ~A166;
  assign \new_[37359]_  = A234 & A233;
  assign \new_[37360]_  = \new_[37359]_  & \new_[37356]_ ;
  assign \new_[37361]_  = \new_[37360]_  & \new_[37353]_ ;
  assign \new_[37364]_  = ~A267 & A235;
  assign \new_[37367]_  = A298 & A268;
  assign \new_[37368]_  = \new_[37367]_  & \new_[37364]_ ;
  assign \new_[37371]_  = ~A300 & ~A299;
  assign \new_[37374]_  = A302 & ~A301;
  assign \new_[37375]_  = \new_[37374]_  & \new_[37371]_ ;
  assign \new_[37376]_  = \new_[37375]_  & \new_[37368]_ ;
  assign \new_[37380]_  = A167 & A168;
  assign \new_[37381]_  = A169 & \new_[37380]_ ;
  assign \new_[37384]_  = ~A232 & ~A166;
  assign \new_[37387]_  = A234 & A233;
  assign \new_[37388]_  = \new_[37387]_  & \new_[37384]_ ;
  assign \new_[37389]_  = \new_[37388]_  & \new_[37381]_ ;
  assign \new_[37392]_  = ~A267 & A235;
  assign \new_[37395]_  = ~A298 & A268;
  assign \new_[37396]_  = \new_[37395]_  & \new_[37392]_ ;
  assign \new_[37399]_  = ~A300 & A299;
  assign \new_[37402]_  = A302 & ~A301;
  assign \new_[37403]_  = \new_[37402]_  & \new_[37399]_ ;
  assign \new_[37404]_  = \new_[37403]_  & \new_[37396]_ ;
  assign \new_[37408]_  = A167 & A168;
  assign \new_[37409]_  = A169 & \new_[37408]_ ;
  assign \new_[37412]_  = ~A232 & ~A166;
  assign \new_[37415]_  = A234 & A233;
  assign \new_[37416]_  = \new_[37415]_  & \new_[37412]_ ;
  assign \new_[37417]_  = \new_[37416]_  & \new_[37409]_ ;
  assign \new_[37420]_  = ~A267 & A235;
  assign \new_[37423]_  = A298 & ~A269;
  assign \new_[37424]_  = \new_[37423]_  & \new_[37420]_ ;
  assign \new_[37427]_  = ~A300 & ~A299;
  assign \new_[37430]_  = A302 & ~A301;
  assign \new_[37431]_  = \new_[37430]_  & \new_[37427]_ ;
  assign \new_[37432]_  = \new_[37431]_  & \new_[37424]_ ;
  assign \new_[37436]_  = A167 & A168;
  assign \new_[37437]_  = A169 & \new_[37436]_ ;
  assign \new_[37440]_  = ~A232 & ~A166;
  assign \new_[37443]_  = A234 & A233;
  assign \new_[37444]_  = \new_[37443]_  & \new_[37440]_ ;
  assign \new_[37445]_  = \new_[37444]_  & \new_[37437]_ ;
  assign \new_[37448]_  = ~A267 & A235;
  assign \new_[37451]_  = ~A298 & ~A269;
  assign \new_[37452]_  = \new_[37451]_  & \new_[37448]_ ;
  assign \new_[37455]_  = ~A300 & A299;
  assign \new_[37458]_  = A302 & ~A301;
  assign \new_[37459]_  = \new_[37458]_  & \new_[37455]_ ;
  assign \new_[37460]_  = \new_[37459]_  & \new_[37452]_ ;
  assign \new_[37464]_  = A167 & A168;
  assign \new_[37465]_  = A169 & \new_[37464]_ ;
  assign \new_[37468]_  = ~A232 & ~A166;
  assign \new_[37471]_  = A234 & A233;
  assign \new_[37472]_  = \new_[37471]_  & \new_[37468]_ ;
  assign \new_[37473]_  = \new_[37472]_  & \new_[37465]_ ;
  assign \new_[37476]_  = A265 & A235;
  assign \new_[37479]_  = A298 & A266;
  assign \new_[37480]_  = \new_[37479]_  & \new_[37476]_ ;
  assign \new_[37483]_  = ~A300 & ~A299;
  assign \new_[37486]_  = A302 & ~A301;
  assign \new_[37487]_  = \new_[37486]_  & \new_[37483]_ ;
  assign \new_[37488]_  = \new_[37487]_  & \new_[37480]_ ;
  assign \new_[37492]_  = A167 & A168;
  assign \new_[37493]_  = A169 & \new_[37492]_ ;
  assign \new_[37496]_  = ~A232 & ~A166;
  assign \new_[37499]_  = A234 & A233;
  assign \new_[37500]_  = \new_[37499]_  & \new_[37496]_ ;
  assign \new_[37501]_  = \new_[37500]_  & \new_[37493]_ ;
  assign \new_[37504]_  = A265 & A235;
  assign \new_[37507]_  = ~A298 & A266;
  assign \new_[37508]_  = \new_[37507]_  & \new_[37504]_ ;
  assign \new_[37511]_  = ~A300 & A299;
  assign \new_[37514]_  = A302 & ~A301;
  assign \new_[37515]_  = \new_[37514]_  & \new_[37511]_ ;
  assign \new_[37516]_  = \new_[37515]_  & \new_[37508]_ ;
  assign \new_[37520]_  = A167 & A168;
  assign \new_[37521]_  = A169 & \new_[37520]_ ;
  assign \new_[37524]_  = ~A232 & ~A166;
  assign \new_[37527]_  = A234 & A233;
  assign \new_[37528]_  = \new_[37527]_  & \new_[37524]_ ;
  assign \new_[37529]_  = \new_[37528]_  & \new_[37521]_ ;
  assign \new_[37532]_  = ~A265 & A235;
  assign \new_[37535]_  = A298 & ~A266;
  assign \new_[37536]_  = \new_[37535]_  & \new_[37532]_ ;
  assign \new_[37539]_  = ~A300 & ~A299;
  assign \new_[37542]_  = A302 & ~A301;
  assign \new_[37543]_  = \new_[37542]_  & \new_[37539]_ ;
  assign \new_[37544]_  = \new_[37543]_  & \new_[37536]_ ;
  assign \new_[37548]_  = A167 & A168;
  assign \new_[37549]_  = A169 & \new_[37548]_ ;
  assign \new_[37552]_  = ~A232 & ~A166;
  assign \new_[37555]_  = A234 & A233;
  assign \new_[37556]_  = \new_[37555]_  & \new_[37552]_ ;
  assign \new_[37557]_  = \new_[37556]_  & \new_[37549]_ ;
  assign \new_[37560]_  = ~A265 & A235;
  assign \new_[37563]_  = ~A298 & ~A266;
  assign \new_[37564]_  = \new_[37563]_  & \new_[37560]_ ;
  assign \new_[37567]_  = ~A300 & A299;
  assign \new_[37570]_  = A302 & ~A301;
  assign \new_[37571]_  = \new_[37570]_  & \new_[37567]_ ;
  assign \new_[37572]_  = \new_[37571]_  & \new_[37564]_ ;
  assign \new_[37576]_  = A167 & A168;
  assign \new_[37577]_  = A169 & \new_[37576]_ ;
  assign \new_[37580]_  = ~A232 & ~A166;
  assign \new_[37583]_  = A234 & A233;
  assign \new_[37584]_  = \new_[37583]_  & \new_[37580]_ ;
  assign \new_[37585]_  = \new_[37584]_  & \new_[37577]_ ;
  assign \new_[37588]_  = A267 & ~A236;
  assign \new_[37591]_  = A269 & ~A268;
  assign \new_[37592]_  = \new_[37591]_  & \new_[37588]_ ;
  assign \new_[37595]_  = ~A299 & A298;
  assign \new_[37598]_  = A301 & A300;
  assign \new_[37599]_  = \new_[37598]_  & \new_[37595]_ ;
  assign \new_[37600]_  = \new_[37599]_  & \new_[37592]_ ;
  assign \new_[37604]_  = A167 & A168;
  assign \new_[37605]_  = A169 & \new_[37604]_ ;
  assign \new_[37608]_  = ~A232 & ~A166;
  assign \new_[37611]_  = A234 & A233;
  assign \new_[37612]_  = \new_[37611]_  & \new_[37608]_ ;
  assign \new_[37613]_  = \new_[37612]_  & \new_[37605]_ ;
  assign \new_[37616]_  = A267 & ~A236;
  assign \new_[37619]_  = A269 & ~A268;
  assign \new_[37620]_  = \new_[37619]_  & \new_[37616]_ ;
  assign \new_[37623]_  = ~A299 & A298;
  assign \new_[37626]_  = ~A302 & A300;
  assign \new_[37627]_  = \new_[37626]_  & \new_[37623]_ ;
  assign \new_[37628]_  = \new_[37627]_  & \new_[37620]_ ;
  assign \new_[37632]_  = A167 & A168;
  assign \new_[37633]_  = A169 & \new_[37632]_ ;
  assign \new_[37636]_  = ~A232 & ~A166;
  assign \new_[37639]_  = A234 & A233;
  assign \new_[37640]_  = \new_[37639]_  & \new_[37636]_ ;
  assign \new_[37641]_  = \new_[37640]_  & \new_[37633]_ ;
  assign \new_[37644]_  = A267 & ~A236;
  assign \new_[37647]_  = A269 & ~A268;
  assign \new_[37648]_  = \new_[37647]_  & \new_[37644]_ ;
  assign \new_[37651]_  = A299 & ~A298;
  assign \new_[37654]_  = A301 & A300;
  assign \new_[37655]_  = \new_[37654]_  & \new_[37651]_ ;
  assign \new_[37656]_  = \new_[37655]_  & \new_[37648]_ ;
  assign \new_[37660]_  = A167 & A168;
  assign \new_[37661]_  = A169 & \new_[37660]_ ;
  assign \new_[37664]_  = ~A232 & ~A166;
  assign \new_[37667]_  = A234 & A233;
  assign \new_[37668]_  = \new_[37667]_  & \new_[37664]_ ;
  assign \new_[37669]_  = \new_[37668]_  & \new_[37661]_ ;
  assign \new_[37672]_  = A267 & ~A236;
  assign \new_[37675]_  = A269 & ~A268;
  assign \new_[37676]_  = \new_[37675]_  & \new_[37672]_ ;
  assign \new_[37679]_  = A299 & ~A298;
  assign \new_[37682]_  = ~A302 & A300;
  assign \new_[37683]_  = \new_[37682]_  & \new_[37679]_ ;
  assign \new_[37684]_  = \new_[37683]_  & \new_[37676]_ ;
  assign \new_[37688]_  = A167 & A168;
  assign \new_[37689]_  = A169 & \new_[37688]_ ;
  assign \new_[37692]_  = ~A232 & ~A166;
  assign \new_[37695]_  = A234 & A233;
  assign \new_[37696]_  = \new_[37695]_  & \new_[37692]_ ;
  assign \new_[37697]_  = \new_[37696]_  & \new_[37689]_ ;
  assign \new_[37700]_  = ~A267 & ~A236;
  assign \new_[37703]_  = A298 & A268;
  assign \new_[37704]_  = \new_[37703]_  & \new_[37700]_ ;
  assign \new_[37707]_  = ~A300 & ~A299;
  assign \new_[37710]_  = A302 & ~A301;
  assign \new_[37711]_  = \new_[37710]_  & \new_[37707]_ ;
  assign \new_[37712]_  = \new_[37711]_  & \new_[37704]_ ;
  assign \new_[37716]_  = A167 & A168;
  assign \new_[37717]_  = A169 & \new_[37716]_ ;
  assign \new_[37720]_  = ~A232 & ~A166;
  assign \new_[37723]_  = A234 & A233;
  assign \new_[37724]_  = \new_[37723]_  & \new_[37720]_ ;
  assign \new_[37725]_  = \new_[37724]_  & \new_[37717]_ ;
  assign \new_[37728]_  = ~A267 & ~A236;
  assign \new_[37731]_  = ~A298 & A268;
  assign \new_[37732]_  = \new_[37731]_  & \new_[37728]_ ;
  assign \new_[37735]_  = ~A300 & A299;
  assign \new_[37738]_  = A302 & ~A301;
  assign \new_[37739]_  = \new_[37738]_  & \new_[37735]_ ;
  assign \new_[37740]_  = \new_[37739]_  & \new_[37732]_ ;
  assign \new_[37744]_  = A167 & A168;
  assign \new_[37745]_  = A169 & \new_[37744]_ ;
  assign \new_[37748]_  = ~A232 & ~A166;
  assign \new_[37751]_  = A234 & A233;
  assign \new_[37752]_  = \new_[37751]_  & \new_[37748]_ ;
  assign \new_[37753]_  = \new_[37752]_  & \new_[37745]_ ;
  assign \new_[37756]_  = ~A267 & ~A236;
  assign \new_[37759]_  = A298 & ~A269;
  assign \new_[37760]_  = \new_[37759]_  & \new_[37756]_ ;
  assign \new_[37763]_  = ~A300 & ~A299;
  assign \new_[37766]_  = A302 & ~A301;
  assign \new_[37767]_  = \new_[37766]_  & \new_[37763]_ ;
  assign \new_[37768]_  = \new_[37767]_  & \new_[37760]_ ;
  assign \new_[37772]_  = A167 & A168;
  assign \new_[37773]_  = A169 & \new_[37772]_ ;
  assign \new_[37776]_  = ~A232 & ~A166;
  assign \new_[37779]_  = A234 & A233;
  assign \new_[37780]_  = \new_[37779]_  & \new_[37776]_ ;
  assign \new_[37781]_  = \new_[37780]_  & \new_[37773]_ ;
  assign \new_[37784]_  = ~A267 & ~A236;
  assign \new_[37787]_  = ~A298 & ~A269;
  assign \new_[37788]_  = \new_[37787]_  & \new_[37784]_ ;
  assign \new_[37791]_  = ~A300 & A299;
  assign \new_[37794]_  = A302 & ~A301;
  assign \new_[37795]_  = \new_[37794]_  & \new_[37791]_ ;
  assign \new_[37796]_  = \new_[37795]_  & \new_[37788]_ ;
  assign \new_[37800]_  = A167 & A168;
  assign \new_[37801]_  = A169 & \new_[37800]_ ;
  assign \new_[37804]_  = ~A232 & ~A166;
  assign \new_[37807]_  = A234 & A233;
  assign \new_[37808]_  = \new_[37807]_  & \new_[37804]_ ;
  assign \new_[37809]_  = \new_[37808]_  & \new_[37801]_ ;
  assign \new_[37812]_  = A265 & ~A236;
  assign \new_[37815]_  = A298 & A266;
  assign \new_[37816]_  = \new_[37815]_  & \new_[37812]_ ;
  assign \new_[37819]_  = ~A300 & ~A299;
  assign \new_[37822]_  = A302 & ~A301;
  assign \new_[37823]_  = \new_[37822]_  & \new_[37819]_ ;
  assign \new_[37824]_  = \new_[37823]_  & \new_[37816]_ ;
  assign \new_[37828]_  = A167 & A168;
  assign \new_[37829]_  = A169 & \new_[37828]_ ;
  assign \new_[37832]_  = ~A232 & ~A166;
  assign \new_[37835]_  = A234 & A233;
  assign \new_[37836]_  = \new_[37835]_  & \new_[37832]_ ;
  assign \new_[37837]_  = \new_[37836]_  & \new_[37829]_ ;
  assign \new_[37840]_  = A265 & ~A236;
  assign \new_[37843]_  = ~A298 & A266;
  assign \new_[37844]_  = \new_[37843]_  & \new_[37840]_ ;
  assign \new_[37847]_  = ~A300 & A299;
  assign \new_[37850]_  = A302 & ~A301;
  assign \new_[37851]_  = \new_[37850]_  & \new_[37847]_ ;
  assign \new_[37852]_  = \new_[37851]_  & \new_[37844]_ ;
  assign \new_[37856]_  = A167 & A168;
  assign \new_[37857]_  = A169 & \new_[37856]_ ;
  assign \new_[37860]_  = ~A232 & ~A166;
  assign \new_[37863]_  = A234 & A233;
  assign \new_[37864]_  = \new_[37863]_  & \new_[37860]_ ;
  assign \new_[37865]_  = \new_[37864]_  & \new_[37857]_ ;
  assign \new_[37868]_  = ~A265 & ~A236;
  assign \new_[37871]_  = A298 & ~A266;
  assign \new_[37872]_  = \new_[37871]_  & \new_[37868]_ ;
  assign \new_[37875]_  = ~A300 & ~A299;
  assign \new_[37878]_  = A302 & ~A301;
  assign \new_[37879]_  = \new_[37878]_  & \new_[37875]_ ;
  assign \new_[37880]_  = \new_[37879]_  & \new_[37872]_ ;
  assign \new_[37884]_  = A167 & A168;
  assign \new_[37885]_  = A169 & \new_[37884]_ ;
  assign \new_[37888]_  = ~A232 & ~A166;
  assign \new_[37891]_  = A234 & A233;
  assign \new_[37892]_  = \new_[37891]_  & \new_[37888]_ ;
  assign \new_[37893]_  = \new_[37892]_  & \new_[37885]_ ;
  assign \new_[37896]_  = ~A265 & ~A236;
  assign \new_[37899]_  = ~A298 & ~A266;
  assign \new_[37900]_  = \new_[37899]_  & \new_[37896]_ ;
  assign \new_[37903]_  = ~A300 & A299;
  assign \new_[37906]_  = A302 & ~A301;
  assign \new_[37907]_  = \new_[37906]_  & \new_[37903]_ ;
  assign \new_[37908]_  = \new_[37907]_  & \new_[37900]_ ;
  assign \new_[37912]_  = A167 & A168;
  assign \new_[37913]_  = A169 & \new_[37912]_ ;
  assign \new_[37916]_  = ~A232 & ~A166;
  assign \new_[37919]_  = ~A234 & A233;
  assign \new_[37920]_  = \new_[37919]_  & \new_[37916]_ ;
  assign \new_[37921]_  = \new_[37920]_  & \new_[37913]_ ;
  assign \new_[37924]_  = A236 & ~A235;
  assign \new_[37927]_  = A268 & ~A267;
  assign \new_[37928]_  = \new_[37927]_  & \new_[37924]_ ;
  assign \new_[37931]_  = ~A299 & A298;
  assign \new_[37934]_  = A301 & A300;
  assign \new_[37935]_  = \new_[37934]_  & \new_[37931]_ ;
  assign \new_[37936]_  = \new_[37935]_  & \new_[37928]_ ;
  assign \new_[37940]_  = A167 & A168;
  assign \new_[37941]_  = A169 & \new_[37940]_ ;
  assign \new_[37944]_  = ~A232 & ~A166;
  assign \new_[37947]_  = ~A234 & A233;
  assign \new_[37948]_  = \new_[37947]_  & \new_[37944]_ ;
  assign \new_[37949]_  = \new_[37948]_  & \new_[37941]_ ;
  assign \new_[37952]_  = A236 & ~A235;
  assign \new_[37955]_  = A268 & ~A267;
  assign \new_[37956]_  = \new_[37955]_  & \new_[37952]_ ;
  assign \new_[37959]_  = ~A299 & A298;
  assign \new_[37962]_  = ~A302 & A300;
  assign \new_[37963]_  = \new_[37962]_  & \new_[37959]_ ;
  assign \new_[37964]_  = \new_[37963]_  & \new_[37956]_ ;
  assign \new_[37968]_  = A167 & A168;
  assign \new_[37969]_  = A169 & \new_[37968]_ ;
  assign \new_[37972]_  = ~A232 & ~A166;
  assign \new_[37975]_  = ~A234 & A233;
  assign \new_[37976]_  = \new_[37975]_  & \new_[37972]_ ;
  assign \new_[37977]_  = \new_[37976]_  & \new_[37969]_ ;
  assign \new_[37980]_  = A236 & ~A235;
  assign \new_[37983]_  = A268 & ~A267;
  assign \new_[37984]_  = \new_[37983]_  & \new_[37980]_ ;
  assign \new_[37987]_  = A299 & ~A298;
  assign \new_[37990]_  = A301 & A300;
  assign \new_[37991]_  = \new_[37990]_  & \new_[37987]_ ;
  assign \new_[37992]_  = \new_[37991]_  & \new_[37984]_ ;
  assign \new_[37996]_  = A167 & A168;
  assign \new_[37997]_  = A169 & \new_[37996]_ ;
  assign \new_[38000]_  = ~A232 & ~A166;
  assign \new_[38003]_  = ~A234 & A233;
  assign \new_[38004]_  = \new_[38003]_  & \new_[38000]_ ;
  assign \new_[38005]_  = \new_[38004]_  & \new_[37997]_ ;
  assign \new_[38008]_  = A236 & ~A235;
  assign \new_[38011]_  = A268 & ~A267;
  assign \new_[38012]_  = \new_[38011]_  & \new_[38008]_ ;
  assign \new_[38015]_  = A299 & ~A298;
  assign \new_[38018]_  = ~A302 & A300;
  assign \new_[38019]_  = \new_[38018]_  & \new_[38015]_ ;
  assign \new_[38020]_  = \new_[38019]_  & \new_[38012]_ ;
  assign \new_[38024]_  = A167 & A168;
  assign \new_[38025]_  = A169 & \new_[38024]_ ;
  assign \new_[38028]_  = ~A232 & ~A166;
  assign \new_[38031]_  = ~A234 & A233;
  assign \new_[38032]_  = \new_[38031]_  & \new_[38028]_ ;
  assign \new_[38033]_  = \new_[38032]_  & \new_[38025]_ ;
  assign \new_[38036]_  = A236 & ~A235;
  assign \new_[38039]_  = ~A269 & ~A267;
  assign \new_[38040]_  = \new_[38039]_  & \new_[38036]_ ;
  assign \new_[38043]_  = ~A299 & A298;
  assign \new_[38046]_  = A301 & A300;
  assign \new_[38047]_  = \new_[38046]_  & \new_[38043]_ ;
  assign \new_[38048]_  = \new_[38047]_  & \new_[38040]_ ;
  assign \new_[38052]_  = A167 & A168;
  assign \new_[38053]_  = A169 & \new_[38052]_ ;
  assign \new_[38056]_  = ~A232 & ~A166;
  assign \new_[38059]_  = ~A234 & A233;
  assign \new_[38060]_  = \new_[38059]_  & \new_[38056]_ ;
  assign \new_[38061]_  = \new_[38060]_  & \new_[38053]_ ;
  assign \new_[38064]_  = A236 & ~A235;
  assign \new_[38067]_  = ~A269 & ~A267;
  assign \new_[38068]_  = \new_[38067]_  & \new_[38064]_ ;
  assign \new_[38071]_  = ~A299 & A298;
  assign \new_[38074]_  = ~A302 & A300;
  assign \new_[38075]_  = \new_[38074]_  & \new_[38071]_ ;
  assign \new_[38076]_  = \new_[38075]_  & \new_[38068]_ ;
  assign \new_[38080]_  = A167 & A168;
  assign \new_[38081]_  = A169 & \new_[38080]_ ;
  assign \new_[38084]_  = ~A232 & ~A166;
  assign \new_[38087]_  = ~A234 & A233;
  assign \new_[38088]_  = \new_[38087]_  & \new_[38084]_ ;
  assign \new_[38089]_  = \new_[38088]_  & \new_[38081]_ ;
  assign \new_[38092]_  = A236 & ~A235;
  assign \new_[38095]_  = ~A269 & ~A267;
  assign \new_[38096]_  = \new_[38095]_  & \new_[38092]_ ;
  assign \new_[38099]_  = A299 & ~A298;
  assign \new_[38102]_  = A301 & A300;
  assign \new_[38103]_  = \new_[38102]_  & \new_[38099]_ ;
  assign \new_[38104]_  = \new_[38103]_  & \new_[38096]_ ;
  assign \new_[38108]_  = A167 & A168;
  assign \new_[38109]_  = A169 & \new_[38108]_ ;
  assign \new_[38112]_  = ~A232 & ~A166;
  assign \new_[38115]_  = ~A234 & A233;
  assign \new_[38116]_  = \new_[38115]_  & \new_[38112]_ ;
  assign \new_[38117]_  = \new_[38116]_  & \new_[38109]_ ;
  assign \new_[38120]_  = A236 & ~A235;
  assign \new_[38123]_  = ~A269 & ~A267;
  assign \new_[38124]_  = \new_[38123]_  & \new_[38120]_ ;
  assign \new_[38127]_  = A299 & ~A298;
  assign \new_[38130]_  = ~A302 & A300;
  assign \new_[38131]_  = \new_[38130]_  & \new_[38127]_ ;
  assign \new_[38132]_  = \new_[38131]_  & \new_[38124]_ ;
  assign \new_[38136]_  = A167 & A168;
  assign \new_[38137]_  = A169 & \new_[38136]_ ;
  assign \new_[38140]_  = ~A232 & ~A166;
  assign \new_[38143]_  = ~A234 & A233;
  assign \new_[38144]_  = \new_[38143]_  & \new_[38140]_ ;
  assign \new_[38145]_  = \new_[38144]_  & \new_[38137]_ ;
  assign \new_[38148]_  = A236 & ~A235;
  assign \new_[38151]_  = A266 & A265;
  assign \new_[38152]_  = \new_[38151]_  & \new_[38148]_ ;
  assign \new_[38155]_  = ~A299 & A298;
  assign \new_[38158]_  = A301 & A300;
  assign \new_[38159]_  = \new_[38158]_  & \new_[38155]_ ;
  assign \new_[38160]_  = \new_[38159]_  & \new_[38152]_ ;
  assign \new_[38164]_  = A167 & A168;
  assign \new_[38165]_  = A169 & \new_[38164]_ ;
  assign \new_[38168]_  = ~A232 & ~A166;
  assign \new_[38171]_  = ~A234 & A233;
  assign \new_[38172]_  = \new_[38171]_  & \new_[38168]_ ;
  assign \new_[38173]_  = \new_[38172]_  & \new_[38165]_ ;
  assign \new_[38176]_  = A236 & ~A235;
  assign \new_[38179]_  = A266 & A265;
  assign \new_[38180]_  = \new_[38179]_  & \new_[38176]_ ;
  assign \new_[38183]_  = ~A299 & A298;
  assign \new_[38186]_  = ~A302 & A300;
  assign \new_[38187]_  = \new_[38186]_  & \new_[38183]_ ;
  assign \new_[38188]_  = \new_[38187]_  & \new_[38180]_ ;
  assign \new_[38192]_  = A167 & A168;
  assign \new_[38193]_  = A169 & \new_[38192]_ ;
  assign \new_[38196]_  = ~A232 & ~A166;
  assign \new_[38199]_  = ~A234 & A233;
  assign \new_[38200]_  = \new_[38199]_  & \new_[38196]_ ;
  assign \new_[38201]_  = \new_[38200]_  & \new_[38193]_ ;
  assign \new_[38204]_  = A236 & ~A235;
  assign \new_[38207]_  = A266 & A265;
  assign \new_[38208]_  = \new_[38207]_  & \new_[38204]_ ;
  assign \new_[38211]_  = A299 & ~A298;
  assign \new_[38214]_  = A301 & A300;
  assign \new_[38215]_  = \new_[38214]_  & \new_[38211]_ ;
  assign \new_[38216]_  = \new_[38215]_  & \new_[38208]_ ;
  assign \new_[38220]_  = A167 & A168;
  assign \new_[38221]_  = A169 & \new_[38220]_ ;
  assign \new_[38224]_  = ~A232 & ~A166;
  assign \new_[38227]_  = ~A234 & A233;
  assign \new_[38228]_  = \new_[38227]_  & \new_[38224]_ ;
  assign \new_[38229]_  = \new_[38228]_  & \new_[38221]_ ;
  assign \new_[38232]_  = A236 & ~A235;
  assign \new_[38235]_  = A266 & A265;
  assign \new_[38236]_  = \new_[38235]_  & \new_[38232]_ ;
  assign \new_[38239]_  = A299 & ~A298;
  assign \new_[38242]_  = ~A302 & A300;
  assign \new_[38243]_  = \new_[38242]_  & \new_[38239]_ ;
  assign \new_[38244]_  = \new_[38243]_  & \new_[38236]_ ;
  assign \new_[38248]_  = A167 & A168;
  assign \new_[38249]_  = A169 & \new_[38248]_ ;
  assign \new_[38252]_  = ~A232 & ~A166;
  assign \new_[38255]_  = ~A234 & A233;
  assign \new_[38256]_  = \new_[38255]_  & \new_[38252]_ ;
  assign \new_[38257]_  = \new_[38256]_  & \new_[38249]_ ;
  assign \new_[38260]_  = A236 & ~A235;
  assign \new_[38263]_  = ~A266 & ~A265;
  assign \new_[38264]_  = \new_[38263]_  & \new_[38260]_ ;
  assign \new_[38267]_  = ~A299 & A298;
  assign \new_[38270]_  = A301 & A300;
  assign \new_[38271]_  = \new_[38270]_  & \new_[38267]_ ;
  assign \new_[38272]_  = \new_[38271]_  & \new_[38264]_ ;
  assign \new_[38276]_  = A167 & A168;
  assign \new_[38277]_  = A169 & \new_[38276]_ ;
  assign \new_[38280]_  = ~A232 & ~A166;
  assign \new_[38283]_  = ~A234 & A233;
  assign \new_[38284]_  = \new_[38283]_  & \new_[38280]_ ;
  assign \new_[38285]_  = \new_[38284]_  & \new_[38277]_ ;
  assign \new_[38288]_  = A236 & ~A235;
  assign \new_[38291]_  = ~A266 & ~A265;
  assign \new_[38292]_  = \new_[38291]_  & \new_[38288]_ ;
  assign \new_[38295]_  = ~A299 & A298;
  assign \new_[38298]_  = ~A302 & A300;
  assign \new_[38299]_  = \new_[38298]_  & \new_[38295]_ ;
  assign \new_[38300]_  = \new_[38299]_  & \new_[38292]_ ;
  assign \new_[38304]_  = A167 & A168;
  assign \new_[38305]_  = A169 & \new_[38304]_ ;
  assign \new_[38308]_  = ~A232 & ~A166;
  assign \new_[38311]_  = ~A234 & A233;
  assign \new_[38312]_  = \new_[38311]_  & \new_[38308]_ ;
  assign \new_[38313]_  = \new_[38312]_  & \new_[38305]_ ;
  assign \new_[38316]_  = A236 & ~A235;
  assign \new_[38319]_  = ~A266 & ~A265;
  assign \new_[38320]_  = \new_[38319]_  & \new_[38316]_ ;
  assign \new_[38323]_  = A299 & ~A298;
  assign \new_[38326]_  = A301 & A300;
  assign \new_[38327]_  = \new_[38326]_  & \new_[38323]_ ;
  assign \new_[38328]_  = \new_[38327]_  & \new_[38320]_ ;
  assign \new_[38332]_  = A167 & A168;
  assign \new_[38333]_  = A169 & \new_[38332]_ ;
  assign \new_[38336]_  = ~A232 & ~A166;
  assign \new_[38339]_  = ~A234 & A233;
  assign \new_[38340]_  = \new_[38339]_  & \new_[38336]_ ;
  assign \new_[38341]_  = \new_[38340]_  & \new_[38333]_ ;
  assign \new_[38344]_  = A236 & ~A235;
  assign \new_[38347]_  = ~A266 & ~A265;
  assign \new_[38348]_  = \new_[38347]_  & \new_[38344]_ ;
  assign \new_[38351]_  = A299 & ~A298;
  assign \new_[38354]_  = ~A302 & A300;
  assign \new_[38355]_  = \new_[38354]_  & \new_[38351]_ ;
  assign \new_[38356]_  = \new_[38355]_  & \new_[38348]_ ;
  assign \new_[38360]_  = A167 & A168;
  assign \new_[38361]_  = A169 & \new_[38360]_ ;
  assign \new_[38364]_  = A232 & ~A166;
  assign \new_[38367]_  = A234 & ~A233;
  assign \new_[38368]_  = \new_[38367]_  & \new_[38364]_ ;
  assign \new_[38369]_  = \new_[38368]_  & \new_[38361]_ ;
  assign \new_[38372]_  = A267 & A235;
  assign \new_[38375]_  = A269 & ~A268;
  assign \new_[38376]_  = \new_[38375]_  & \new_[38372]_ ;
  assign \new_[38379]_  = ~A299 & A298;
  assign \new_[38382]_  = A301 & A300;
  assign \new_[38383]_  = \new_[38382]_  & \new_[38379]_ ;
  assign \new_[38384]_  = \new_[38383]_  & \new_[38376]_ ;
  assign \new_[38388]_  = A167 & A168;
  assign \new_[38389]_  = A169 & \new_[38388]_ ;
  assign \new_[38392]_  = A232 & ~A166;
  assign \new_[38395]_  = A234 & ~A233;
  assign \new_[38396]_  = \new_[38395]_  & \new_[38392]_ ;
  assign \new_[38397]_  = \new_[38396]_  & \new_[38389]_ ;
  assign \new_[38400]_  = A267 & A235;
  assign \new_[38403]_  = A269 & ~A268;
  assign \new_[38404]_  = \new_[38403]_  & \new_[38400]_ ;
  assign \new_[38407]_  = ~A299 & A298;
  assign \new_[38410]_  = ~A302 & A300;
  assign \new_[38411]_  = \new_[38410]_  & \new_[38407]_ ;
  assign \new_[38412]_  = \new_[38411]_  & \new_[38404]_ ;
  assign \new_[38416]_  = A167 & A168;
  assign \new_[38417]_  = A169 & \new_[38416]_ ;
  assign \new_[38420]_  = A232 & ~A166;
  assign \new_[38423]_  = A234 & ~A233;
  assign \new_[38424]_  = \new_[38423]_  & \new_[38420]_ ;
  assign \new_[38425]_  = \new_[38424]_  & \new_[38417]_ ;
  assign \new_[38428]_  = A267 & A235;
  assign \new_[38431]_  = A269 & ~A268;
  assign \new_[38432]_  = \new_[38431]_  & \new_[38428]_ ;
  assign \new_[38435]_  = A299 & ~A298;
  assign \new_[38438]_  = A301 & A300;
  assign \new_[38439]_  = \new_[38438]_  & \new_[38435]_ ;
  assign \new_[38440]_  = \new_[38439]_  & \new_[38432]_ ;
  assign \new_[38444]_  = A167 & A168;
  assign \new_[38445]_  = A169 & \new_[38444]_ ;
  assign \new_[38448]_  = A232 & ~A166;
  assign \new_[38451]_  = A234 & ~A233;
  assign \new_[38452]_  = \new_[38451]_  & \new_[38448]_ ;
  assign \new_[38453]_  = \new_[38452]_  & \new_[38445]_ ;
  assign \new_[38456]_  = A267 & A235;
  assign \new_[38459]_  = A269 & ~A268;
  assign \new_[38460]_  = \new_[38459]_  & \new_[38456]_ ;
  assign \new_[38463]_  = A299 & ~A298;
  assign \new_[38466]_  = ~A302 & A300;
  assign \new_[38467]_  = \new_[38466]_  & \new_[38463]_ ;
  assign \new_[38468]_  = \new_[38467]_  & \new_[38460]_ ;
  assign \new_[38472]_  = A167 & A168;
  assign \new_[38473]_  = A169 & \new_[38472]_ ;
  assign \new_[38476]_  = A232 & ~A166;
  assign \new_[38479]_  = A234 & ~A233;
  assign \new_[38480]_  = \new_[38479]_  & \new_[38476]_ ;
  assign \new_[38481]_  = \new_[38480]_  & \new_[38473]_ ;
  assign \new_[38484]_  = ~A267 & A235;
  assign \new_[38487]_  = A298 & A268;
  assign \new_[38488]_  = \new_[38487]_  & \new_[38484]_ ;
  assign \new_[38491]_  = ~A300 & ~A299;
  assign \new_[38494]_  = A302 & ~A301;
  assign \new_[38495]_  = \new_[38494]_  & \new_[38491]_ ;
  assign \new_[38496]_  = \new_[38495]_  & \new_[38488]_ ;
  assign \new_[38500]_  = A167 & A168;
  assign \new_[38501]_  = A169 & \new_[38500]_ ;
  assign \new_[38504]_  = A232 & ~A166;
  assign \new_[38507]_  = A234 & ~A233;
  assign \new_[38508]_  = \new_[38507]_  & \new_[38504]_ ;
  assign \new_[38509]_  = \new_[38508]_  & \new_[38501]_ ;
  assign \new_[38512]_  = ~A267 & A235;
  assign \new_[38515]_  = ~A298 & A268;
  assign \new_[38516]_  = \new_[38515]_  & \new_[38512]_ ;
  assign \new_[38519]_  = ~A300 & A299;
  assign \new_[38522]_  = A302 & ~A301;
  assign \new_[38523]_  = \new_[38522]_  & \new_[38519]_ ;
  assign \new_[38524]_  = \new_[38523]_  & \new_[38516]_ ;
  assign \new_[38528]_  = A167 & A168;
  assign \new_[38529]_  = A169 & \new_[38528]_ ;
  assign \new_[38532]_  = A232 & ~A166;
  assign \new_[38535]_  = A234 & ~A233;
  assign \new_[38536]_  = \new_[38535]_  & \new_[38532]_ ;
  assign \new_[38537]_  = \new_[38536]_  & \new_[38529]_ ;
  assign \new_[38540]_  = ~A267 & A235;
  assign \new_[38543]_  = A298 & ~A269;
  assign \new_[38544]_  = \new_[38543]_  & \new_[38540]_ ;
  assign \new_[38547]_  = ~A300 & ~A299;
  assign \new_[38550]_  = A302 & ~A301;
  assign \new_[38551]_  = \new_[38550]_  & \new_[38547]_ ;
  assign \new_[38552]_  = \new_[38551]_  & \new_[38544]_ ;
  assign \new_[38556]_  = A167 & A168;
  assign \new_[38557]_  = A169 & \new_[38556]_ ;
  assign \new_[38560]_  = A232 & ~A166;
  assign \new_[38563]_  = A234 & ~A233;
  assign \new_[38564]_  = \new_[38563]_  & \new_[38560]_ ;
  assign \new_[38565]_  = \new_[38564]_  & \new_[38557]_ ;
  assign \new_[38568]_  = ~A267 & A235;
  assign \new_[38571]_  = ~A298 & ~A269;
  assign \new_[38572]_  = \new_[38571]_  & \new_[38568]_ ;
  assign \new_[38575]_  = ~A300 & A299;
  assign \new_[38578]_  = A302 & ~A301;
  assign \new_[38579]_  = \new_[38578]_  & \new_[38575]_ ;
  assign \new_[38580]_  = \new_[38579]_  & \new_[38572]_ ;
  assign \new_[38584]_  = A167 & A168;
  assign \new_[38585]_  = A169 & \new_[38584]_ ;
  assign \new_[38588]_  = A232 & ~A166;
  assign \new_[38591]_  = A234 & ~A233;
  assign \new_[38592]_  = \new_[38591]_  & \new_[38588]_ ;
  assign \new_[38593]_  = \new_[38592]_  & \new_[38585]_ ;
  assign \new_[38596]_  = A265 & A235;
  assign \new_[38599]_  = A298 & A266;
  assign \new_[38600]_  = \new_[38599]_  & \new_[38596]_ ;
  assign \new_[38603]_  = ~A300 & ~A299;
  assign \new_[38606]_  = A302 & ~A301;
  assign \new_[38607]_  = \new_[38606]_  & \new_[38603]_ ;
  assign \new_[38608]_  = \new_[38607]_  & \new_[38600]_ ;
  assign \new_[38612]_  = A167 & A168;
  assign \new_[38613]_  = A169 & \new_[38612]_ ;
  assign \new_[38616]_  = A232 & ~A166;
  assign \new_[38619]_  = A234 & ~A233;
  assign \new_[38620]_  = \new_[38619]_  & \new_[38616]_ ;
  assign \new_[38621]_  = \new_[38620]_  & \new_[38613]_ ;
  assign \new_[38624]_  = A265 & A235;
  assign \new_[38627]_  = ~A298 & A266;
  assign \new_[38628]_  = \new_[38627]_  & \new_[38624]_ ;
  assign \new_[38631]_  = ~A300 & A299;
  assign \new_[38634]_  = A302 & ~A301;
  assign \new_[38635]_  = \new_[38634]_  & \new_[38631]_ ;
  assign \new_[38636]_  = \new_[38635]_  & \new_[38628]_ ;
  assign \new_[38640]_  = A167 & A168;
  assign \new_[38641]_  = A169 & \new_[38640]_ ;
  assign \new_[38644]_  = A232 & ~A166;
  assign \new_[38647]_  = A234 & ~A233;
  assign \new_[38648]_  = \new_[38647]_  & \new_[38644]_ ;
  assign \new_[38649]_  = \new_[38648]_  & \new_[38641]_ ;
  assign \new_[38652]_  = ~A265 & A235;
  assign \new_[38655]_  = A298 & ~A266;
  assign \new_[38656]_  = \new_[38655]_  & \new_[38652]_ ;
  assign \new_[38659]_  = ~A300 & ~A299;
  assign \new_[38662]_  = A302 & ~A301;
  assign \new_[38663]_  = \new_[38662]_  & \new_[38659]_ ;
  assign \new_[38664]_  = \new_[38663]_  & \new_[38656]_ ;
  assign \new_[38668]_  = A167 & A168;
  assign \new_[38669]_  = A169 & \new_[38668]_ ;
  assign \new_[38672]_  = A232 & ~A166;
  assign \new_[38675]_  = A234 & ~A233;
  assign \new_[38676]_  = \new_[38675]_  & \new_[38672]_ ;
  assign \new_[38677]_  = \new_[38676]_  & \new_[38669]_ ;
  assign \new_[38680]_  = ~A265 & A235;
  assign \new_[38683]_  = ~A298 & ~A266;
  assign \new_[38684]_  = \new_[38683]_  & \new_[38680]_ ;
  assign \new_[38687]_  = ~A300 & A299;
  assign \new_[38690]_  = A302 & ~A301;
  assign \new_[38691]_  = \new_[38690]_  & \new_[38687]_ ;
  assign \new_[38692]_  = \new_[38691]_  & \new_[38684]_ ;
  assign \new_[38696]_  = A167 & A168;
  assign \new_[38697]_  = A169 & \new_[38696]_ ;
  assign \new_[38700]_  = A232 & ~A166;
  assign \new_[38703]_  = A234 & ~A233;
  assign \new_[38704]_  = \new_[38703]_  & \new_[38700]_ ;
  assign \new_[38705]_  = \new_[38704]_  & \new_[38697]_ ;
  assign \new_[38708]_  = A267 & ~A236;
  assign \new_[38711]_  = A269 & ~A268;
  assign \new_[38712]_  = \new_[38711]_  & \new_[38708]_ ;
  assign \new_[38715]_  = ~A299 & A298;
  assign \new_[38718]_  = A301 & A300;
  assign \new_[38719]_  = \new_[38718]_  & \new_[38715]_ ;
  assign \new_[38720]_  = \new_[38719]_  & \new_[38712]_ ;
  assign \new_[38724]_  = A167 & A168;
  assign \new_[38725]_  = A169 & \new_[38724]_ ;
  assign \new_[38728]_  = A232 & ~A166;
  assign \new_[38731]_  = A234 & ~A233;
  assign \new_[38732]_  = \new_[38731]_  & \new_[38728]_ ;
  assign \new_[38733]_  = \new_[38732]_  & \new_[38725]_ ;
  assign \new_[38736]_  = A267 & ~A236;
  assign \new_[38739]_  = A269 & ~A268;
  assign \new_[38740]_  = \new_[38739]_  & \new_[38736]_ ;
  assign \new_[38743]_  = ~A299 & A298;
  assign \new_[38746]_  = ~A302 & A300;
  assign \new_[38747]_  = \new_[38746]_  & \new_[38743]_ ;
  assign \new_[38748]_  = \new_[38747]_  & \new_[38740]_ ;
  assign \new_[38752]_  = A167 & A168;
  assign \new_[38753]_  = A169 & \new_[38752]_ ;
  assign \new_[38756]_  = A232 & ~A166;
  assign \new_[38759]_  = A234 & ~A233;
  assign \new_[38760]_  = \new_[38759]_  & \new_[38756]_ ;
  assign \new_[38761]_  = \new_[38760]_  & \new_[38753]_ ;
  assign \new_[38764]_  = A267 & ~A236;
  assign \new_[38767]_  = A269 & ~A268;
  assign \new_[38768]_  = \new_[38767]_  & \new_[38764]_ ;
  assign \new_[38771]_  = A299 & ~A298;
  assign \new_[38774]_  = A301 & A300;
  assign \new_[38775]_  = \new_[38774]_  & \new_[38771]_ ;
  assign \new_[38776]_  = \new_[38775]_  & \new_[38768]_ ;
  assign \new_[38780]_  = A167 & A168;
  assign \new_[38781]_  = A169 & \new_[38780]_ ;
  assign \new_[38784]_  = A232 & ~A166;
  assign \new_[38787]_  = A234 & ~A233;
  assign \new_[38788]_  = \new_[38787]_  & \new_[38784]_ ;
  assign \new_[38789]_  = \new_[38788]_  & \new_[38781]_ ;
  assign \new_[38792]_  = A267 & ~A236;
  assign \new_[38795]_  = A269 & ~A268;
  assign \new_[38796]_  = \new_[38795]_  & \new_[38792]_ ;
  assign \new_[38799]_  = A299 & ~A298;
  assign \new_[38802]_  = ~A302 & A300;
  assign \new_[38803]_  = \new_[38802]_  & \new_[38799]_ ;
  assign \new_[38804]_  = \new_[38803]_  & \new_[38796]_ ;
  assign \new_[38808]_  = A167 & A168;
  assign \new_[38809]_  = A169 & \new_[38808]_ ;
  assign \new_[38812]_  = A232 & ~A166;
  assign \new_[38815]_  = A234 & ~A233;
  assign \new_[38816]_  = \new_[38815]_  & \new_[38812]_ ;
  assign \new_[38817]_  = \new_[38816]_  & \new_[38809]_ ;
  assign \new_[38820]_  = ~A267 & ~A236;
  assign \new_[38823]_  = A298 & A268;
  assign \new_[38824]_  = \new_[38823]_  & \new_[38820]_ ;
  assign \new_[38827]_  = ~A300 & ~A299;
  assign \new_[38830]_  = A302 & ~A301;
  assign \new_[38831]_  = \new_[38830]_  & \new_[38827]_ ;
  assign \new_[38832]_  = \new_[38831]_  & \new_[38824]_ ;
  assign \new_[38836]_  = A167 & A168;
  assign \new_[38837]_  = A169 & \new_[38836]_ ;
  assign \new_[38840]_  = A232 & ~A166;
  assign \new_[38843]_  = A234 & ~A233;
  assign \new_[38844]_  = \new_[38843]_  & \new_[38840]_ ;
  assign \new_[38845]_  = \new_[38844]_  & \new_[38837]_ ;
  assign \new_[38848]_  = ~A267 & ~A236;
  assign \new_[38851]_  = ~A298 & A268;
  assign \new_[38852]_  = \new_[38851]_  & \new_[38848]_ ;
  assign \new_[38855]_  = ~A300 & A299;
  assign \new_[38858]_  = A302 & ~A301;
  assign \new_[38859]_  = \new_[38858]_  & \new_[38855]_ ;
  assign \new_[38860]_  = \new_[38859]_  & \new_[38852]_ ;
  assign \new_[38864]_  = A167 & A168;
  assign \new_[38865]_  = A169 & \new_[38864]_ ;
  assign \new_[38868]_  = A232 & ~A166;
  assign \new_[38871]_  = A234 & ~A233;
  assign \new_[38872]_  = \new_[38871]_  & \new_[38868]_ ;
  assign \new_[38873]_  = \new_[38872]_  & \new_[38865]_ ;
  assign \new_[38876]_  = ~A267 & ~A236;
  assign \new_[38879]_  = A298 & ~A269;
  assign \new_[38880]_  = \new_[38879]_  & \new_[38876]_ ;
  assign \new_[38883]_  = ~A300 & ~A299;
  assign \new_[38886]_  = A302 & ~A301;
  assign \new_[38887]_  = \new_[38886]_  & \new_[38883]_ ;
  assign \new_[38888]_  = \new_[38887]_  & \new_[38880]_ ;
  assign \new_[38892]_  = A167 & A168;
  assign \new_[38893]_  = A169 & \new_[38892]_ ;
  assign \new_[38896]_  = A232 & ~A166;
  assign \new_[38899]_  = A234 & ~A233;
  assign \new_[38900]_  = \new_[38899]_  & \new_[38896]_ ;
  assign \new_[38901]_  = \new_[38900]_  & \new_[38893]_ ;
  assign \new_[38904]_  = ~A267 & ~A236;
  assign \new_[38907]_  = ~A298 & ~A269;
  assign \new_[38908]_  = \new_[38907]_  & \new_[38904]_ ;
  assign \new_[38911]_  = ~A300 & A299;
  assign \new_[38914]_  = A302 & ~A301;
  assign \new_[38915]_  = \new_[38914]_  & \new_[38911]_ ;
  assign \new_[38916]_  = \new_[38915]_  & \new_[38908]_ ;
  assign \new_[38920]_  = A167 & A168;
  assign \new_[38921]_  = A169 & \new_[38920]_ ;
  assign \new_[38924]_  = A232 & ~A166;
  assign \new_[38927]_  = A234 & ~A233;
  assign \new_[38928]_  = \new_[38927]_  & \new_[38924]_ ;
  assign \new_[38929]_  = \new_[38928]_  & \new_[38921]_ ;
  assign \new_[38932]_  = A265 & ~A236;
  assign \new_[38935]_  = A298 & A266;
  assign \new_[38936]_  = \new_[38935]_  & \new_[38932]_ ;
  assign \new_[38939]_  = ~A300 & ~A299;
  assign \new_[38942]_  = A302 & ~A301;
  assign \new_[38943]_  = \new_[38942]_  & \new_[38939]_ ;
  assign \new_[38944]_  = \new_[38943]_  & \new_[38936]_ ;
  assign \new_[38948]_  = A167 & A168;
  assign \new_[38949]_  = A169 & \new_[38948]_ ;
  assign \new_[38952]_  = A232 & ~A166;
  assign \new_[38955]_  = A234 & ~A233;
  assign \new_[38956]_  = \new_[38955]_  & \new_[38952]_ ;
  assign \new_[38957]_  = \new_[38956]_  & \new_[38949]_ ;
  assign \new_[38960]_  = A265 & ~A236;
  assign \new_[38963]_  = ~A298 & A266;
  assign \new_[38964]_  = \new_[38963]_  & \new_[38960]_ ;
  assign \new_[38967]_  = ~A300 & A299;
  assign \new_[38970]_  = A302 & ~A301;
  assign \new_[38971]_  = \new_[38970]_  & \new_[38967]_ ;
  assign \new_[38972]_  = \new_[38971]_  & \new_[38964]_ ;
  assign \new_[38976]_  = A167 & A168;
  assign \new_[38977]_  = A169 & \new_[38976]_ ;
  assign \new_[38980]_  = A232 & ~A166;
  assign \new_[38983]_  = A234 & ~A233;
  assign \new_[38984]_  = \new_[38983]_  & \new_[38980]_ ;
  assign \new_[38985]_  = \new_[38984]_  & \new_[38977]_ ;
  assign \new_[38988]_  = ~A265 & ~A236;
  assign \new_[38991]_  = A298 & ~A266;
  assign \new_[38992]_  = \new_[38991]_  & \new_[38988]_ ;
  assign \new_[38995]_  = ~A300 & ~A299;
  assign \new_[38998]_  = A302 & ~A301;
  assign \new_[38999]_  = \new_[38998]_  & \new_[38995]_ ;
  assign \new_[39000]_  = \new_[38999]_  & \new_[38992]_ ;
  assign \new_[39004]_  = A167 & A168;
  assign \new_[39005]_  = A169 & \new_[39004]_ ;
  assign \new_[39008]_  = A232 & ~A166;
  assign \new_[39011]_  = A234 & ~A233;
  assign \new_[39012]_  = \new_[39011]_  & \new_[39008]_ ;
  assign \new_[39013]_  = \new_[39012]_  & \new_[39005]_ ;
  assign \new_[39016]_  = ~A265 & ~A236;
  assign \new_[39019]_  = ~A298 & ~A266;
  assign \new_[39020]_  = \new_[39019]_  & \new_[39016]_ ;
  assign \new_[39023]_  = ~A300 & A299;
  assign \new_[39026]_  = A302 & ~A301;
  assign \new_[39027]_  = \new_[39026]_  & \new_[39023]_ ;
  assign \new_[39028]_  = \new_[39027]_  & \new_[39020]_ ;
  assign \new_[39032]_  = A167 & A168;
  assign \new_[39033]_  = A169 & \new_[39032]_ ;
  assign \new_[39036]_  = A232 & ~A166;
  assign \new_[39039]_  = ~A234 & ~A233;
  assign \new_[39040]_  = \new_[39039]_  & \new_[39036]_ ;
  assign \new_[39041]_  = \new_[39040]_  & \new_[39033]_ ;
  assign \new_[39044]_  = A236 & ~A235;
  assign \new_[39047]_  = A268 & ~A267;
  assign \new_[39048]_  = \new_[39047]_  & \new_[39044]_ ;
  assign \new_[39051]_  = ~A299 & A298;
  assign \new_[39054]_  = A301 & A300;
  assign \new_[39055]_  = \new_[39054]_  & \new_[39051]_ ;
  assign \new_[39056]_  = \new_[39055]_  & \new_[39048]_ ;
  assign \new_[39060]_  = A167 & A168;
  assign \new_[39061]_  = A169 & \new_[39060]_ ;
  assign \new_[39064]_  = A232 & ~A166;
  assign \new_[39067]_  = ~A234 & ~A233;
  assign \new_[39068]_  = \new_[39067]_  & \new_[39064]_ ;
  assign \new_[39069]_  = \new_[39068]_  & \new_[39061]_ ;
  assign \new_[39072]_  = A236 & ~A235;
  assign \new_[39075]_  = A268 & ~A267;
  assign \new_[39076]_  = \new_[39075]_  & \new_[39072]_ ;
  assign \new_[39079]_  = ~A299 & A298;
  assign \new_[39082]_  = ~A302 & A300;
  assign \new_[39083]_  = \new_[39082]_  & \new_[39079]_ ;
  assign \new_[39084]_  = \new_[39083]_  & \new_[39076]_ ;
  assign \new_[39088]_  = A167 & A168;
  assign \new_[39089]_  = A169 & \new_[39088]_ ;
  assign \new_[39092]_  = A232 & ~A166;
  assign \new_[39095]_  = ~A234 & ~A233;
  assign \new_[39096]_  = \new_[39095]_  & \new_[39092]_ ;
  assign \new_[39097]_  = \new_[39096]_  & \new_[39089]_ ;
  assign \new_[39100]_  = A236 & ~A235;
  assign \new_[39103]_  = A268 & ~A267;
  assign \new_[39104]_  = \new_[39103]_  & \new_[39100]_ ;
  assign \new_[39107]_  = A299 & ~A298;
  assign \new_[39110]_  = A301 & A300;
  assign \new_[39111]_  = \new_[39110]_  & \new_[39107]_ ;
  assign \new_[39112]_  = \new_[39111]_  & \new_[39104]_ ;
  assign \new_[39116]_  = A167 & A168;
  assign \new_[39117]_  = A169 & \new_[39116]_ ;
  assign \new_[39120]_  = A232 & ~A166;
  assign \new_[39123]_  = ~A234 & ~A233;
  assign \new_[39124]_  = \new_[39123]_  & \new_[39120]_ ;
  assign \new_[39125]_  = \new_[39124]_  & \new_[39117]_ ;
  assign \new_[39128]_  = A236 & ~A235;
  assign \new_[39131]_  = A268 & ~A267;
  assign \new_[39132]_  = \new_[39131]_  & \new_[39128]_ ;
  assign \new_[39135]_  = A299 & ~A298;
  assign \new_[39138]_  = ~A302 & A300;
  assign \new_[39139]_  = \new_[39138]_  & \new_[39135]_ ;
  assign \new_[39140]_  = \new_[39139]_  & \new_[39132]_ ;
  assign \new_[39144]_  = A167 & A168;
  assign \new_[39145]_  = A169 & \new_[39144]_ ;
  assign \new_[39148]_  = A232 & ~A166;
  assign \new_[39151]_  = ~A234 & ~A233;
  assign \new_[39152]_  = \new_[39151]_  & \new_[39148]_ ;
  assign \new_[39153]_  = \new_[39152]_  & \new_[39145]_ ;
  assign \new_[39156]_  = A236 & ~A235;
  assign \new_[39159]_  = ~A269 & ~A267;
  assign \new_[39160]_  = \new_[39159]_  & \new_[39156]_ ;
  assign \new_[39163]_  = ~A299 & A298;
  assign \new_[39166]_  = A301 & A300;
  assign \new_[39167]_  = \new_[39166]_  & \new_[39163]_ ;
  assign \new_[39168]_  = \new_[39167]_  & \new_[39160]_ ;
  assign \new_[39172]_  = A167 & A168;
  assign \new_[39173]_  = A169 & \new_[39172]_ ;
  assign \new_[39176]_  = A232 & ~A166;
  assign \new_[39179]_  = ~A234 & ~A233;
  assign \new_[39180]_  = \new_[39179]_  & \new_[39176]_ ;
  assign \new_[39181]_  = \new_[39180]_  & \new_[39173]_ ;
  assign \new_[39184]_  = A236 & ~A235;
  assign \new_[39187]_  = ~A269 & ~A267;
  assign \new_[39188]_  = \new_[39187]_  & \new_[39184]_ ;
  assign \new_[39191]_  = ~A299 & A298;
  assign \new_[39194]_  = ~A302 & A300;
  assign \new_[39195]_  = \new_[39194]_  & \new_[39191]_ ;
  assign \new_[39196]_  = \new_[39195]_  & \new_[39188]_ ;
  assign \new_[39200]_  = A167 & A168;
  assign \new_[39201]_  = A169 & \new_[39200]_ ;
  assign \new_[39204]_  = A232 & ~A166;
  assign \new_[39207]_  = ~A234 & ~A233;
  assign \new_[39208]_  = \new_[39207]_  & \new_[39204]_ ;
  assign \new_[39209]_  = \new_[39208]_  & \new_[39201]_ ;
  assign \new_[39212]_  = A236 & ~A235;
  assign \new_[39215]_  = ~A269 & ~A267;
  assign \new_[39216]_  = \new_[39215]_  & \new_[39212]_ ;
  assign \new_[39219]_  = A299 & ~A298;
  assign \new_[39222]_  = A301 & A300;
  assign \new_[39223]_  = \new_[39222]_  & \new_[39219]_ ;
  assign \new_[39224]_  = \new_[39223]_  & \new_[39216]_ ;
  assign \new_[39228]_  = A167 & A168;
  assign \new_[39229]_  = A169 & \new_[39228]_ ;
  assign \new_[39232]_  = A232 & ~A166;
  assign \new_[39235]_  = ~A234 & ~A233;
  assign \new_[39236]_  = \new_[39235]_  & \new_[39232]_ ;
  assign \new_[39237]_  = \new_[39236]_  & \new_[39229]_ ;
  assign \new_[39240]_  = A236 & ~A235;
  assign \new_[39243]_  = ~A269 & ~A267;
  assign \new_[39244]_  = \new_[39243]_  & \new_[39240]_ ;
  assign \new_[39247]_  = A299 & ~A298;
  assign \new_[39250]_  = ~A302 & A300;
  assign \new_[39251]_  = \new_[39250]_  & \new_[39247]_ ;
  assign \new_[39252]_  = \new_[39251]_  & \new_[39244]_ ;
  assign \new_[39256]_  = A167 & A168;
  assign \new_[39257]_  = A169 & \new_[39256]_ ;
  assign \new_[39260]_  = A232 & ~A166;
  assign \new_[39263]_  = ~A234 & ~A233;
  assign \new_[39264]_  = \new_[39263]_  & \new_[39260]_ ;
  assign \new_[39265]_  = \new_[39264]_  & \new_[39257]_ ;
  assign \new_[39268]_  = A236 & ~A235;
  assign \new_[39271]_  = A266 & A265;
  assign \new_[39272]_  = \new_[39271]_  & \new_[39268]_ ;
  assign \new_[39275]_  = ~A299 & A298;
  assign \new_[39278]_  = A301 & A300;
  assign \new_[39279]_  = \new_[39278]_  & \new_[39275]_ ;
  assign \new_[39280]_  = \new_[39279]_  & \new_[39272]_ ;
  assign \new_[39284]_  = A167 & A168;
  assign \new_[39285]_  = A169 & \new_[39284]_ ;
  assign \new_[39288]_  = A232 & ~A166;
  assign \new_[39291]_  = ~A234 & ~A233;
  assign \new_[39292]_  = \new_[39291]_  & \new_[39288]_ ;
  assign \new_[39293]_  = \new_[39292]_  & \new_[39285]_ ;
  assign \new_[39296]_  = A236 & ~A235;
  assign \new_[39299]_  = A266 & A265;
  assign \new_[39300]_  = \new_[39299]_  & \new_[39296]_ ;
  assign \new_[39303]_  = ~A299 & A298;
  assign \new_[39306]_  = ~A302 & A300;
  assign \new_[39307]_  = \new_[39306]_  & \new_[39303]_ ;
  assign \new_[39308]_  = \new_[39307]_  & \new_[39300]_ ;
  assign \new_[39312]_  = A167 & A168;
  assign \new_[39313]_  = A169 & \new_[39312]_ ;
  assign \new_[39316]_  = A232 & ~A166;
  assign \new_[39319]_  = ~A234 & ~A233;
  assign \new_[39320]_  = \new_[39319]_  & \new_[39316]_ ;
  assign \new_[39321]_  = \new_[39320]_  & \new_[39313]_ ;
  assign \new_[39324]_  = A236 & ~A235;
  assign \new_[39327]_  = A266 & A265;
  assign \new_[39328]_  = \new_[39327]_  & \new_[39324]_ ;
  assign \new_[39331]_  = A299 & ~A298;
  assign \new_[39334]_  = A301 & A300;
  assign \new_[39335]_  = \new_[39334]_  & \new_[39331]_ ;
  assign \new_[39336]_  = \new_[39335]_  & \new_[39328]_ ;
  assign \new_[39340]_  = A167 & A168;
  assign \new_[39341]_  = A169 & \new_[39340]_ ;
  assign \new_[39344]_  = A232 & ~A166;
  assign \new_[39347]_  = ~A234 & ~A233;
  assign \new_[39348]_  = \new_[39347]_  & \new_[39344]_ ;
  assign \new_[39349]_  = \new_[39348]_  & \new_[39341]_ ;
  assign \new_[39352]_  = A236 & ~A235;
  assign \new_[39355]_  = A266 & A265;
  assign \new_[39356]_  = \new_[39355]_  & \new_[39352]_ ;
  assign \new_[39359]_  = A299 & ~A298;
  assign \new_[39362]_  = ~A302 & A300;
  assign \new_[39363]_  = \new_[39362]_  & \new_[39359]_ ;
  assign \new_[39364]_  = \new_[39363]_  & \new_[39356]_ ;
  assign \new_[39368]_  = A167 & A168;
  assign \new_[39369]_  = A169 & \new_[39368]_ ;
  assign \new_[39372]_  = A232 & ~A166;
  assign \new_[39375]_  = ~A234 & ~A233;
  assign \new_[39376]_  = \new_[39375]_  & \new_[39372]_ ;
  assign \new_[39377]_  = \new_[39376]_  & \new_[39369]_ ;
  assign \new_[39380]_  = A236 & ~A235;
  assign \new_[39383]_  = ~A266 & ~A265;
  assign \new_[39384]_  = \new_[39383]_  & \new_[39380]_ ;
  assign \new_[39387]_  = ~A299 & A298;
  assign \new_[39390]_  = A301 & A300;
  assign \new_[39391]_  = \new_[39390]_  & \new_[39387]_ ;
  assign \new_[39392]_  = \new_[39391]_  & \new_[39384]_ ;
  assign \new_[39396]_  = A167 & A168;
  assign \new_[39397]_  = A169 & \new_[39396]_ ;
  assign \new_[39400]_  = A232 & ~A166;
  assign \new_[39403]_  = ~A234 & ~A233;
  assign \new_[39404]_  = \new_[39403]_  & \new_[39400]_ ;
  assign \new_[39405]_  = \new_[39404]_  & \new_[39397]_ ;
  assign \new_[39408]_  = A236 & ~A235;
  assign \new_[39411]_  = ~A266 & ~A265;
  assign \new_[39412]_  = \new_[39411]_  & \new_[39408]_ ;
  assign \new_[39415]_  = ~A299 & A298;
  assign \new_[39418]_  = ~A302 & A300;
  assign \new_[39419]_  = \new_[39418]_  & \new_[39415]_ ;
  assign \new_[39420]_  = \new_[39419]_  & \new_[39412]_ ;
  assign \new_[39424]_  = A167 & A168;
  assign \new_[39425]_  = A169 & \new_[39424]_ ;
  assign \new_[39428]_  = A232 & ~A166;
  assign \new_[39431]_  = ~A234 & ~A233;
  assign \new_[39432]_  = \new_[39431]_  & \new_[39428]_ ;
  assign \new_[39433]_  = \new_[39432]_  & \new_[39425]_ ;
  assign \new_[39436]_  = A236 & ~A235;
  assign \new_[39439]_  = ~A266 & ~A265;
  assign \new_[39440]_  = \new_[39439]_  & \new_[39436]_ ;
  assign \new_[39443]_  = A299 & ~A298;
  assign \new_[39446]_  = A301 & A300;
  assign \new_[39447]_  = \new_[39446]_  & \new_[39443]_ ;
  assign \new_[39448]_  = \new_[39447]_  & \new_[39440]_ ;
  assign \new_[39452]_  = A167 & A168;
  assign \new_[39453]_  = A169 & \new_[39452]_ ;
  assign \new_[39456]_  = A232 & ~A166;
  assign \new_[39459]_  = ~A234 & ~A233;
  assign \new_[39460]_  = \new_[39459]_  & \new_[39456]_ ;
  assign \new_[39461]_  = \new_[39460]_  & \new_[39453]_ ;
  assign \new_[39464]_  = A236 & ~A235;
  assign \new_[39467]_  = ~A266 & ~A265;
  assign \new_[39468]_  = \new_[39467]_  & \new_[39464]_ ;
  assign \new_[39471]_  = A299 & ~A298;
  assign \new_[39474]_  = ~A302 & A300;
  assign \new_[39475]_  = \new_[39474]_  & \new_[39471]_ ;
  assign \new_[39476]_  = \new_[39475]_  & \new_[39468]_ ;
  assign \new_[39480]_  = ~A167 & A168;
  assign \new_[39481]_  = A169 & \new_[39480]_ ;
  assign \new_[39484]_  = ~A232 & A166;
  assign \new_[39487]_  = A234 & A233;
  assign \new_[39488]_  = \new_[39487]_  & \new_[39484]_ ;
  assign \new_[39489]_  = \new_[39488]_  & \new_[39481]_ ;
  assign \new_[39492]_  = A267 & A235;
  assign \new_[39495]_  = A269 & ~A268;
  assign \new_[39496]_  = \new_[39495]_  & \new_[39492]_ ;
  assign \new_[39499]_  = ~A299 & A298;
  assign \new_[39502]_  = A301 & A300;
  assign \new_[39503]_  = \new_[39502]_  & \new_[39499]_ ;
  assign \new_[39504]_  = \new_[39503]_  & \new_[39496]_ ;
  assign \new_[39508]_  = ~A167 & A168;
  assign \new_[39509]_  = A169 & \new_[39508]_ ;
  assign \new_[39512]_  = ~A232 & A166;
  assign \new_[39515]_  = A234 & A233;
  assign \new_[39516]_  = \new_[39515]_  & \new_[39512]_ ;
  assign \new_[39517]_  = \new_[39516]_  & \new_[39509]_ ;
  assign \new_[39520]_  = A267 & A235;
  assign \new_[39523]_  = A269 & ~A268;
  assign \new_[39524]_  = \new_[39523]_  & \new_[39520]_ ;
  assign \new_[39527]_  = ~A299 & A298;
  assign \new_[39530]_  = ~A302 & A300;
  assign \new_[39531]_  = \new_[39530]_  & \new_[39527]_ ;
  assign \new_[39532]_  = \new_[39531]_  & \new_[39524]_ ;
  assign \new_[39536]_  = ~A167 & A168;
  assign \new_[39537]_  = A169 & \new_[39536]_ ;
  assign \new_[39540]_  = ~A232 & A166;
  assign \new_[39543]_  = A234 & A233;
  assign \new_[39544]_  = \new_[39543]_  & \new_[39540]_ ;
  assign \new_[39545]_  = \new_[39544]_  & \new_[39537]_ ;
  assign \new_[39548]_  = A267 & A235;
  assign \new_[39551]_  = A269 & ~A268;
  assign \new_[39552]_  = \new_[39551]_  & \new_[39548]_ ;
  assign \new_[39555]_  = A299 & ~A298;
  assign \new_[39558]_  = A301 & A300;
  assign \new_[39559]_  = \new_[39558]_  & \new_[39555]_ ;
  assign \new_[39560]_  = \new_[39559]_  & \new_[39552]_ ;
  assign \new_[39564]_  = ~A167 & A168;
  assign \new_[39565]_  = A169 & \new_[39564]_ ;
  assign \new_[39568]_  = ~A232 & A166;
  assign \new_[39571]_  = A234 & A233;
  assign \new_[39572]_  = \new_[39571]_  & \new_[39568]_ ;
  assign \new_[39573]_  = \new_[39572]_  & \new_[39565]_ ;
  assign \new_[39576]_  = A267 & A235;
  assign \new_[39579]_  = A269 & ~A268;
  assign \new_[39580]_  = \new_[39579]_  & \new_[39576]_ ;
  assign \new_[39583]_  = A299 & ~A298;
  assign \new_[39586]_  = ~A302 & A300;
  assign \new_[39587]_  = \new_[39586]_  & \new_[39583]_ ;
  assign \new_[39588]_  = \new_[39587]_  & \new_[39580]_ ;
  assign \new_[39592]_  = ~A167 & A168;
  assign \new_[39593]_  = A169 & \new_[39592]_ ;
  assign \new_[39596]_  = ~A232 & A166;
  assign \new_[39599]_  = A234 & A233;
  assign \new_[39600]_  = \new_[39599]_  & \new_[39596]_ ;
  assign \new_[39601]_  = \new_[39600]_  & \new_[39593]_ ;
  assign \new_[39604]_  = ~A267 & A235;
  assign \new_[39607]_  = A298 & A268;
  assign \new_[39608]_  = \new_[39607]_  & \new_[39604]_ ;
  assign \new_[39611]_  = ~A300 & ~A299;
  assign \new_[39614]_  = A302 & ~A301;
  assign \new_[39615]_  = \new_[39614]_  & \new_[39611]_ ;
  assign \new_[39616]_  = \new_[39615]_  & \new_[39608]_ ;
  assign \new_[39620]_  = ~A167 & A168;
  assign \new_[39621]_  = A169 & \new_[39620]_ ;
  assign \new_[39624]_  = ~A232 & A166;
  assign \new_[39627]_  = A234 & A233;
  assign \new_[39628]_  = \new_[39627]_  & \new_[39624]_ ;
  assign \new_[39629]_  = \new_[39628]_  & \new_[39621]_ ;
  assign \new_[39632]_  = ~A267 & A235;
  assign \new_[39635]_  = ~A298 & A268;
  assign \new_[39636]_  = \new_[39635]_  & \new_[39632]_ ;
  assign \new_[39639]_  = ~A300 & A299;
  assign \new_[39642]_  = A302 & ~A301;
  assign \new_[39643]_  = \new_[39642]_  & \new_[39639]_ ;
  assign \new_[39644]_  = \new_[39643]_  & \new_[39636]_ ;
  assign \new_[39648]_  = ~A167 & A168;
  assign \new_[39649]_  = A169 & \new_[39648]_ ;
  assign \new_[39652]_  = ~A232 & A166;
  assign \new_[39655]_  = A234 & A233;
  assign \new_[39656]_  = \new_[39655]_  & \new_[39652]_ ;
  assign \new_[39657]_  = \new_[39656]_  & \new_[39649]_ ;
  assign \new_[39660]_  = ~A267 & A235;
  assign \new_[39663]_  = A298 & ~A269;
  assign \new_[39664]_  = \new_[39663]_  & \new_[39660]_ ;
  assign \new_[39667]_  = ~A300 & ~A299;
  assign \new_[39670]_  = A302 & ~A301;
  assign \new_[39671]_  = \new_[39670]_  & \new_[39667]_ ;
  assign \new_[39672]_  = \new_[39671]_  & \new_[39664]_ ;
  assign \new_[39676]_  = ~A167 & A168;
  assign \new_[39677]_  = A169 & \new_[39676]_ ;
  assign \new_[39680]_  = ~A232 & A166;
  assign \new_[39683]_  = A234 & A233;
  assign \new_[39684]_  = \new_[39683]_  & \new_[39680]_ ;
  assign \new_[39685]_  = \new_[39684]_  & \new_[39677]_ ;
  assign \new_[39688]_  = ~A267 & A235;
  assign \new_[39691]_  = ~A298 & ~A269;
  assign \new_[39692]_  = \new_[39691]_  & \new_[39688]_ ;
  assign \new_[39695]_  = ~A300 & A299;
  assign \new_[39698]_  = A302 & ~A301;
  assign \new_[39699]_  = \new_[39698]_  & \new_[39695]_ ;
  assign \new_[39700]_  = \new_[39699]_  & \new_[39692]_ ;
  assign \new_[39704]_  = ~A167 & A168;
  assign \new_[39705]_  = A169 & \new_[39704]_ ;
  assign \new_[39708]_  = ~A232 & A166;
  assign \new_[39711]_  = A234 & A233;
  assign \new_[39712]_  = \new_[39711]_  & \new_[39708]_ ;
  assign \new_[39713]_  = \new_[39712]_  & \new_[39705]_ ;
  assign \new_[39716]_  = A265 & A235;
  assign \new_[39719]_  = A298 & A266;
  assign \new_[39720]_  = \new_[39719]_  & \new_[39716]_ ;
  assign \new_[39723]_  = ~A300 & ~A299;
  assign \new_[39726]_  = A302 & ~A301;
  assign \new_[39727]_  = \new_[39726]_  & \new_[39723]_ ;
  assign \new_[39728]_  = \new_[39727]_  & \new_[39720]_ ;
  assign \new_[39732]_  = ~A167 & A168;
  assign \new_[39733]_  = A169 & \new_[39732]_ ;
  assign \new_[39736]_  = ~A232 & A166;
  assign \new_[39739]_  = A234 & A233;
  assign \new_[39740]_  = \new_[39739]_  & \new_[39736]_ ;
  assign \new_[39741]_  = \new_[39740]_  & \new_[39733]_ ;
  assign \new_[39744]_  = A265 & A235;
  assign \new_[39747]_  = ~A298 & A266;
  assign \new_[39748]_  = \new_[39747]_  & \new_[39744]_ ;
  assign \new_[39751]_  = ~A300 & A299;
  assign \new_[39754]_  = A302 & ~A301;
  assign \new_[39755]_  = \new_[39754]_  & \new_[39751]_ ;
  assign \new_[39756]_  = \new_[39755]_  & \new_[39748]_ ;
  assign \new_[39760]_  = ~A167 & A168;
  assign \new_[39761]_  = A169 & \new_[39760]_ ;
  assign \new_[39764]_  = ~A232 & A166;
  assign \new_[39767]_  = A234 & A233;
  assign \new_[39768]_  = \new_[39767]_  & \new_[39764]_ ;
  assign \new_[39769]_  = \new_[39768]_  & \new_[39761]_ ;
  assign \new_[39772]_  = ~A265 & A235;
  assign \new_[39775]_  = A298 & ~A266;
  assign \new_[39776]_  = \new_[39775]_  & \new_[39772]_ ;
  assign \new_[39779]_  = ~A300 & ~A299;
  assign \new_[39782]_  = A302 & ~A301;
  assign \new_[39783]_  = \new_[39782]_  & \new_[39779]_ ;
  assign \new_[39784]_  = \new_[39783]_  & \new_[39776]_ ;
  assign \new_[39788]_  = ~A167 & A168;
  assign \new_[39789]_  = A169 & \new_[39788]_ ;
  assign \new_[39792]_  = ~A232 & A166;
  assign \new_[39795]_  = A234 & A233;
  assign \new_[39796]_  = \new_[39795]_  & \new_[39792]_ ;
  assign \new_[39797]_  = \new_[39796]_  & \new_[39789]_ ;
  assign \new_[39800]_  = ~A265 & A235;
  assign \new_[39803]_  = ~A298 & ~A266;
  assign \new_[39804]_  = \new_[39803]_  & \new_[39800]_ ;
  assign \new_[39807]_  = ~A300 & A299;
  assign \new_[39810]_  = A302 & ~A301;
  assign \new_[39811]_  = \new_[39810]_  & \new_[39807]_ ;
  assign \new_[39812]_  = \new_[39811]_  & \new_[39804]_ ;
  assign \new_[39816]_  = ~A167 & A168;
  assign \new_[39817]_  = A169 & \new_[39816]_ ;
  assign \new_[39820]_  = ~A232 & A166;
  assign \new_[39823]_  = A234 & A233;
  assign \new_[39824]_  = \new_[39823]_  & \new_[39820]_ ;
  assign \new_[39825]_  = \new_[39824]_  & \new_[39817]_ ;
  assign \new_[39828]_  = A267 & ~A236;
  assign \new_[39831]_  = A269 & ~A268;
  assign \new_[39832]_  = \new_[39831]_  & \new_[39828]_ ;
  assign \new_[39835]_  = ~A299 & A298;
  assign \new_[39838]_  = A301 & A300;
  assign \new_[39839]_  = \new_[39838]_  & \new_[39835]_ ;
  assign \new_[39840]_  = \new_[39839]_  & \new_[39832]_ ;
  assign \new_[39844]_  = ~A167 & A168;
  assign \new_[39845]_  = A169 & \new_[39844]_ ;
  assign \new_[39848]_  = ~A232 & A166;
  assign \new_[39851]_  = A234 & A233;
  assign \new_[39852]_  = \new_[39851]_  & \new_[39848]_ ;
  assign \new_[39853]_  = \new_[39852]_  & \new_[39845]_ ;
  assign \new_[39856]_  = A267 & ~A236;
  assign \new_[39859]_  = A269 & ~A268;
  assign \new_[39860]_  = \new_[39859]_  & \new_[39856]_ ;
  assign \new_[39863]_  = ~A299 & A298;
  assign \new_[39866]_  = ~A302 & A300;
  assign \new_[39867]_  = \new_[39866]_  & \new_[39863]_ ;
  assign \new_[39868]_  = \new_[39867]_  & \new_[39860]_ ;
  assign \new_[39872]_  = ~A167 & A168;
  assign \new_[39873]_  = A169 & \new_[39872]_ ;
  assign \new_[39876]_  = ~A232 & A166;
  assign \new_[39879]_  = A234 & A233;
  assign \new_[39880]_  = \new_[39879]_  & \new_[39876]_ ;
  assign \new_[39881]_  = \new_[39880]_  & \new_[39873]_ ;
  assign \new_[39884]_  = A267 & ~A236;
  assign \new_[39887]_  = A269 & ~A268;
  assign \new_[39888]_  = \new_[39887]_  & \new_[39884]_ ;
  assign \new_[39891]_  = A299 & ~A298;
  assign \new_[39894]_  = A301 & A300;
  assign \new_[39895]_  = \new_[39894]_  & \new_[39891]_ ;
  assign \new_[39896]_  = \new_[39895]_  & \new_[39888]_ ;
  assign \new_[39900]_  = ~A167 & A168;
  assign \new_[39901]_  = A169 & \new_[39900]_ ;
  assign \new_[39904]_  = ~A232 & A166;
  assign \new_[39907]_  = A234 & A233;
  assign \new_[39908]_  = \new_[39907]_  & \new_[39904]_ ;
  assign \new_[39909]_  = \new_[39908]_  & \new_[39901]_ ;
  assign \new_[39912]_  = A267 & ~A236;
  assign \new_[39915]_  = A269 & ~A268;
  assign \new_[39916]_  = \new_[39915]_  & \new_[39912]_ ;
  assign \new_[39919]_  = A299 & ~A298;
  assign \new_[39922]_  = ~A302 & A300;
  assign \new_[39923]_  = \new_[39922]_  & \new_[39919]_ ;
  assign \new_[39924]_  = \new_[39923]_  & \new_[39916]_ ;
  assign \new_[39928]_  = ~A167 & A168;
  assign \new_[39929]_  = A169 & \new_[39928]_ ;
  assign \new_[39932]_  = ~A232 & A166;
  assign \new_[39935]_  = A234 & A233;
  assign \new_[39936]_  = \new_[39935]_  & \new_[39932]_ ;
  assign \new_[39937]_  = \new_[39936]_  & \new_[39929]_ ;
  assign \new_[39940]_  = ~A267 & ~A236;
  assign \new_[39943]_  = A298 & A268;
  assign \new_[39944]_  = \new_[39943]_  & \new_[39940]_ ;
  assign \new_[39947]_  = ~A300 & ~A299;
  assign \new_[39950]_  = A302 & ~A301;
  assign \new_[39951]_  = \new_[39950]_  & \new_[39947]_ ;
  assign \new_[39952]_  = \new_[39951]_  & \new_[39944]_ ;
  assign \new_[39956]_  = ~A167 & A168;
  assign \new_[39957]_  = A169 & \new_[39956]_ ;
  assign \new_[39960]_  = ~A232 & A166;
  assign \new_[39963]_  = A234 & A233;
  assign \new_[39964]_  = \new_[39963]_  & \new_[39960]_ ;
  assign \new_[39965]_  = \new_[39964]_  & \new_[39957]_ ;
  assign \new_[39968]_  = ~A267 & ~A236;
  assign \new_[39971]_  = ~A298 & A268;
  assign \new_[39972]_  = \new_[39971]_  & \new_[39968]_ ;
  assign \new_[39975]_  = ~A300 & A299;
  assign \new_[39978]_  = A302 & ~A301;
  assign \new_[39979]_  = \new_[39978]_  & \new_[39975]_ ;
  assign \new_[39980]_  = \new_[39979]_  & \new_[39972]_ ;
  assign \new_[39984]_  = ~A167 & A168;
  assign \new_[39985]_  = A169 & \new_[39984]_ ;
  assign \new_[39988]_  = ~A232 & A166;
  assign \new_[39991]_  = A234 & A233;
  assign \new_[39992]_  = \new_[39991]_  & \new_[39988]_ ;
  assign \new_[39993]_  = \new_[39992]_  & \new_[39985]_ ;
  assign \new_[39996]_  = ~A267 & ~A236;
  assign \new_[39999]_  = A298 & ~A269;
  assign \new_[40000]_  = \new_[39999]_  & \new_[39996]_ ;
  assign \new_[40003]_  = ~A300 & ~A299;
  assign \new_[40006]_  = A302 & ~A301;
  assign \new_[40007]_  = \new_[40006]_  & \new_[40003]_ ;
  assign \new_[40008]_  = \new_[40007]_  & \new_[40000]_ ;
  assign \new_[40012]_  = ~A167 & A168;
  assign \new_[40013]_  = A169 & \new_[40012]_ ;
  assign \new_[40016]_  = ~A232 & A166;
  assign \new_[40019]_  = A234 & A233;
  assign \new_[40020]_  = \new_[40019]_  & \new_[40016]_ ;
  assign \new_[40021]_  = \new_[40020]_  & \new_[40013]_ ;
  assign \new_[40024]_  = ~A267 & ~A236;
  assign \new_[40027]_  = ~A298 & ~A269;
  assign \new_[40028]_  = \new_[40027]_  & \new_[40024]_ ;
  assign \new_[40031]_  = ~A300 & A299;
  assign \new_[40034]_  = A302 & ~A301;
  assign \new_[40035]_  = \new_[40034]_  & \new_[40031]_ ;
  assign \new_[40036]_  = \new_[40035]_  & \new_[40028]_ ;
  assign \new_[40040]_  = ~A167 & A168;
  assign \new_[40041]_  = A169 & \new_[40040]_ ;
  assign \new_[40044]_  = ~A232 & A166;
  assign \new_[40047]_  = A234 & A233;
  assign \new_[40048]_  = \new_[40047]_  & \new_[40044]_ ;
  assign \new_[40049]_  = \new_[40048]_  & \new_[40041]_ ;
  assign \new_[40052]_  = A265 & ~A236;
  assign \new_[40055]_  = A298 & A266;
  assign \new_[40056]_  = \new_[40055]_  & \new_[40052]_ ;
  assign \new_[40059]_  = ~A300 & ~A299;
  assign \new_[40062]_  = A302 & ~A301;
  assign \new_[40063]_  = \new_[40062]_  & \new_[40059]_ ;
  assign \new_[40064]_  = \new_[40063]_  & \new_[40056]_ ;
  assign \new_[40068]_  = ~A167 & A168;
  assign \new_[40069]_  = A169 & \new_[40068]_ ;
  assign \new_[40072]_  = ~A232 & A166;
  assign \new_[40075]_  = A234 & A233;
  assign \new_[40076]_  = \new_[40075]_  & \new_[40072]_ ;
  assign \new_[40077]_  = \new_[40076]_  & \new_[40069]_ ;
  assign \new_[40080]_  = A265 & ~A236;
  assign \new_[40083]_  = ~A298 & A266;
  assign \new_[40084]_  = \new_[40083]_  & \new_[40080]_ ;
  assign \new_[40087]_  = ~A300 & A299;
  assign \new_[40090]_  = A302 & ~A301;
  assign \new_[40091]_  = \new_[40090]_  & \new_[40087]_ ;
  assign \new_[40092]_  = \new_[40091]_  & \new_[40084]_ ;
  assign \new_[40096]_  = ~A167 & A168;
  assign \new_[40097]_  = A169 & \new_[40096]_ ;
  assign \new_[40100]_  = ~A232 & A166;
  assign \new_[40103]_  = A234 & A233;
  assign \new_[40104]_  = \new_[40103]_  & \new_[40100]_ ;
  assign \new_[40105]_  = \new_[40104]_  & \new_[40097]_ ;
  assign \new_[40108]_  = ~A265 & ~A236;
  assign \new_[40111]_  = A298 & ~A266;
  assign \new_[40112]_  = \new_[40111]_  & \new_[40108]_ ;
  assign \new_[40115]_  = ~A300 & ~A299;
  assign \new_[40118]_  = A302 & ~A301;
  assign \new_[40119]_  = \new_[40118]_  & \new_[40115]_ ;
  assign \new_[40120]_  = \new_[40119]_  & \new_[40112]_ ;
  assign \new_[40124]_  = ~A167 & A168;
  assign \new_[40125]_  = A169 & \new_[40124]_ ;
  assign \new_[40128]_  = ~A232 & A166;
  assign \new_[40131]_  = A234 & A233;
  assign \new_[40132]_  = \new_[40131]_  & \new_[40128]_ ;
  assign \new_[40133]_  = \new_[40132]_  & \new_[40125]_ ;
  assign \new_[40136]_  = ~A265 & ~A236;
  assign \new_[40139]_  = ~A298 & ~A266;
  assign \new_[40140]_  = \new_[40139]_  & \new_[40136]_ ;
  assign \new_[40143]_  = ~A300 & A299;
  assign \new_[40146]_  = A302 & ~A301;
  assign \new_[40147]_  = \new_[40146]_  & \new_[40143]_ ;
  assign \new_[40148]_  = \new_[40147]_  & \new_[40140]_ ;
  assign \new_[40152]_  = ~A167 & A168;
  assign \new_[40153]_  = A169 & \new_[40152]_ ;
  assign \new_[40156]_  = ~A232 & A166;
  assign \new_[40159]_  = ~A234 & A233;
  assign \new_[40160]_  = \new_[40159]_  & \new_[40156]_ ;
  assign \new_[40161]_  = \new_[40160]_  & \new_[40153]_ ;
  assign \new_[40164]_  = A236 & ~A235;
  assign \new_[40167]_  = A268 & ~A267;
  assign \new_[40168]_  = \new_[40167]_  & \new_[40164]_ ;
  assign \new_[40171]_  = ~A299 & A298;
  assign \new_[40174]_  = A301 & A300;
  assign \new_[40175]_  = \new_[40174]_  & \new_[40171]_ ;
  assign \new_[40176]_  = \new_[40175]_  & \new_[40168]_ ;
  assign \new_[40180]_  = ~A167 & A168;
  assign \new_[40181]_  = A169 & \new_[40180]_ ;
  assign \new_[40184]_  = ~A232 & A166;
  assign \new_[40187]_  = ~A234 & A233;
  assign \new_[40188]_  = \new_[40187]_  & \new_[40184]_ ;
  assign \new_[40189]_  = \new_[40188]_  & \new_[40181]_ ;
  assign \new_[40192]_  = A236 & ~A235;
  assign \new_[40195]_  = A268 & ~A267;
  assign \new_[40196]_  = \new_[40195]_  & \new_[40192]_ ;
  assign \new_[40199]_  = ~A299 & A298;
  assign \new_[40202]_  = ~A302 & A300;
  assign \new_[40203]_  = \new_[40202]_  & \new_[40199]_ ;
  assign \new_[40204]_  = \new_[40203]_  & \new_[40196]_ ;
  assign \new_[40208]_  = ~A167 & A168;
  assign \new_[40209]_  = A169 & \new_[40208]_ ;
  assign \new_[40212]_  = ~A232 & A166;
  assign \new_[40215]_  = ~A234 & A233;
  assign \new_[40216]_  = \new_[40215]_  & \new_[40212]_ ;
  assign \new_[40217]_  = \new_[40216]_  & \new_[40209]_ ;
  assign \new_[40220]_  = A236 & ~A235;
  assign \new_[40223]_  = A268 & ~A267;
  assign \new_[40224]_  = \new_[40223]_  & \new_[40220]_ ;
  assign \new_[40227]_  = A299 & ~A298;
  assign \new_[40230]_  = A301 & A300;
  assign \new_[40231]_  = \new_[40230]_  & \new_[40227]_ ;
  assign \new_[40232]_  = \new_[40231]_  & \new_[40224]_ ;
  assign \new_[40236]_  = ~A167 & A168;
  assign \new_[40237]_  = A169 & \new_[40236]_ ;
  assign \new_[40240]_  = ~A232 & A166;
  assign \new_[40243]_  = ~A234 & A233;
  assign \new_[40244]_  = \new_[40243]_  & \new_[40240]_ ;
  assign \new_[40245]_  = \new_[40244]_  & \new_[40237]_ ;
  assign \new_[40248]_  = A236 & ~A235;
  assign \new_[40251]_  = A268 & ~A267;
  assign \new_[40252]_  = \new_[40251]_  & \new_[40248]_ ;
  assign \new_[40255]_  = A299 & ~A298;
  assign \new_[40258]_  = ~A302 & A300;
  assign \new_[40259]_  = \new_[40258]_  & \new_[40255]_ ;
  assign \new_[40260]_  = \new_[40259]_  & \new_[40252]_ ;
  assign \new_[40264]_  = ~A167 & A168;
  assign \new_[40265]_  = A169 & \new_[40264]_ ;
  assign \new_[40268]_  = ~A232 & A166;
  assign \new_[40271]_  = ~A234 & A233;
  assign \new_[40272]_  = \new_[40271]_  & \new_[40268]_ ;
  assign \new_[40273]_  = \new_[40272]_  & \new_[40265]_ ;
  assign \new_[40276]_  = A236 & ~A235;
  assign \new_[40279]_  = ~A269 & ~A267;
  assign \new_[40280]_  = \new_[40279]_  & \new_[40276]_ ;
  assign \new_[40283]_  = ~A299 & A298;
  assign \new_[40286]_  = A301 & A300;
  assign \new_[40287]_  = \new_[40286]_  & \new_[40283]_ ;
  assign \new_[40288]_  = \new_[40287]_  & \new_[40280]_ ;
  assign \new_[40292]_  = ~A167 & A168;
  assign \new_[40293]_  = A169 & \new_[40292]_ ;
  assign \new_[40296]_  = ~A232 & A166;
  assign \new_[40299]_  = ~A234 & A233;
  assign \new_[40300]_  = \new_[40299]_  & \new_[40296]_ ;
  assign \new_[40301]_  = \new_[40300]_  & \new_[40293]_ ;
  assign \new_[40304]_  = A236 & ~A235;
  assign \new_[40307]_  = ~A269 & ~A267;
  assign \new_[40308]_  = \new_[40307]_  & \new_[40304]_ ;
  assign \new_[40311]_  = ~A299 & A298;
  assign \new_[40314]_  = ~A302 & A300;
  assign \new_[40315]_  = \new_[40314]_  & \new_[40311]_ ;
  assign \new_[40316]_  = \new_[40315]_  & \new_[40308]_ ;
  assign \new_[40320]_  = ~A167 & A168;
  assign \new_[40321]_  = A169 & \new_[40320]_ ;
  assign \new_[40324]_  = ~A232 & A166;
  assign \new_[40327]_  = ~A234 & A233;
  assign \new_[40328]_  = \new_[40327]_  & \new_[40324]_ ;
  assign \new_[40329]_  = \new_[40328]_  & \new_[40321]_ ;
  assign \new_[40332]_  = A236 & ~A235;
  assign \new_[40335]_  = ~A269 & ~A267;
  assign \new_[40336]_  = \new_[40335]_  & \new_[40332]_ ;
  assign \new_[40339]_  = A299 & ~A298;
  assign \new_[40342]_  = A301 & A300;
  assign \new_[40343]_  = \new_[40342]_  & \new_[40339]_ ;
  assign \new_[40344]_  = \new_[40343]_  & \new_[40336]_ ;
  assign \new_[40348]_  = ~A167 & A168;
  assign \new_[40349]_  = A169 & \new_[40348]_ ;
  assign \new_[40352]_  = ~A232 & A166;
  assign \new_[40355]_  = ~A234 & A233;
  assign \new_[40356]_  = \new_[40355]_  & \new_[40352]_ ;
  assign \new_[40357]_  = \new_[40356]_  & \new_[40349]_ ;
  assign \new_[40360]_  = A236 & ~A235;
  assign \new_[40363]_  = ~A269 & ~A267;
  assign \new_[40364]_  = \new_[40363]_  & \new_[40360]_ ;
  assign \new_[40367]_  = A299 & ~A298;
  assign \new_[40370]_  = ~A302 & A300;
  assign \new_[40371]_  = \new_[40370]_  & \new_[40367]_ ;
  assign \new_[40372]_  = \new_[40371]_  & \new_[40364]_ ;
  assign \new_[40376]_  = ~A167 & A168;
  assign \new_[40377]_  = A169 & \new_[40376]_ ;
  assign \new_[40380]_  = ~A232 & A166;
  assign \new_[40383]_  = ~A234 & A233;
  assign \new_[40384]_  = \new_[40383]_  & \new_[40380]_ ;
  assign \new_[40385]_  = \new_[40384]_  & \new_[40377]_ ;
  assign \new_[40388]_  = A236 & ~A235;
  assign \new_[40391]_  = A266 & A265;
  assign \new_[40392]_  = \new_[40391]_  & \new_[40388]_ ;
  assign \new_[40395]_  = ~A299 & A298;
  assign \new_[40398]_  = A301 & A300;
  assign \new_[40399]_  = \new_[40398]_  & \new_[40395]_ ;
  assign \new_[40400]_  = \new_[40399]_  & \new_[40392]_ ;
  assign \new_[40404]_  = ~A167 & A168;
  assign \new_[40405]_  = A169 & \new_[40404]_ ;
  assign \new_[40408]_  = ~A232 & A166;
  assign \new_[40411]_  = ~A234 & A233;
  assign \new_[40412]_  = \new_[40411]_  & \new_[40408]_ ;
  assign \new_[40413]_  = \new_[40412]_  & \new_[40405]_ ;
  assign \new_[40416]_  = A236 & ~A235;
  assign \new_[40419]_  = A266 & A265;
  assign \new_[40420]_  = \new_[40419]_  & \new_[40416]_ ;
  assign \new_[40423]_  = ~A299 & A298;
  assign \new_[40426]_  = ~A302 & A300;
  assign \new_[40427]_  = \new_[40426]_  & \new_[40423]_ ;
  assign \new_[40428]_  = \new_[40427]_  & \new_[40420]_ ;
  assign \new_[40432]_  = ~A167 & A168;
  assign \new_[40433]_  = A169 & \new_[40432]_ ;
  assign \new_[40436]_  = ~A232 & A166;
  assign \new_[40439]_  = ~A234 & A233;
  assign \new_[40440]_  = \new_[40439]_  & \new_[40436]_ ;
  assign \new_[40441]_  = \new_[40440]_  & \new_[40433]_ ;
  assign \new_[40444]_  = A236 & ~A235;
  assign \new_[40447]_  = A266 & A265;
  assign \new_[40448]_  = \new_[40447]_  & \new_[40444]_ ;
  assign \new_[40451]_  = A299 & ~A298;
  assign \new_[40454]_  = A301 & A300;
  assign \new_[40455]_  = \new_[40454]_  & \new_[40451]_ ;
  assign \new_[40456]_  = \new_[40455]_  & \new_[40448]_ ;
  assign \new_[40460]_  = ~A167 & A168;
  assign \new_[40461]_  = A169 & \new_[40460]_ ;
  assign \new_[40464]_  = ~A232 & A166;
  assign \new_[40467]_  = ~A234 & A233;
  assign \new_[40468]_  = \new_[40467]_  & \new_[40464]_ ;
  assign \new_[40469]_  = \new_[40468]_  & \new_[40461]_ ;
  assign \new_[40472]_  = A236 & ~A235;
  assign \new_[40475]_  = A266 & A265;
  assign \new_[40476]_  = \new_[40475]_  & \new_[40472]_ ;
  assign \new_[40479]_  = A299 & ~A298;
  assign \new_[40482]_  = ~A302 & A300;
  assign \new_[40483]_  = \new_[40482]_  & \new_[40479]_ ;
  assign \new_[40484]_  = \new_[40483]_  & \new_[40476]_ ;
  assign \new_[40488]_  = ~A167 & A168;
  assign \new_[40489]_  = A169 & \new_[40488]_ ;
  assign \new_[40492]_  = ~A232 & A166;
  assign \new_[40495]_  = ~A234 & A233;
  assign \new_[40496]_  = \new_[40495]_  & \new_[40492]_ ;
  assign \new_[40497]_  = \new_[40496]_  & \new_[40489]_ ;
  assign \new_[40500]_  = A236 & ~A235;
  assign \new_[40503]_  = ~A266 & ~A265;
  assign \new_[40504]_  = \new_[40503]_  & \new_[40500]_ ;
  assign \new_[40507]_  = ~A299 & A298;
  assign \new_[40510]_  = A301 & A300;
  assign \new_[40511]_  = \new_[40510]_  & \new_[40507]_ ;
  assign \new_[40512]_  = \new_[40511]_  & \new_[40504]_ ;
  assign \new_[40516]_  = ~A167 & A168;
  assign \new_[40517]_  = A169 & \new_[40516]_ ;
  assign \new_[40520]_  = ~A232 & A166;
  assign \new_[40523]_  = ~A234 & A233;
  assign \new_[40524]_  = \new_[40523]_  & \new_[40520]_ ;
  assign \new_[40525]_  = \new_[40524]_  & \new_[40517]_ ;
  assign \new_[40528]_  = A236 & ~A235;
  assign \new_[40531]_  = ~A266 & ~A265;
  assign \new_[40532]_  = \new_[40531]_  & \new_[40528]_ ;
  assign \new_[40535]_  = ~A299 & A298;
  assign \new_[40538]_  = ~A302 & A300;
  assign \new_[40539]_  = \new_[40538]_  & \new_[40535]_ ;
  assign \new_[40540]_  = \new_[40539]_  & \new_[40532]_ ;
  assign \new_[40544]_  = ~A167 & A168;
  assign \new_[40545]_  = A169 & \new_[40544]_ ;
  assign \new_[40548]_  = ~A232 & A166;
  assign \new_[40551]_  = ~A234 & A233;
  assign \new_[40552]_  = \new_[40551]_  & \new_[40548]_ ;
  assign \new_[40553]_  = \new_[40552]_  & \new_[40545]_ ;
  assign \new_[40556]_  = A236 & ~A235;
  assign \new_[40559]_  = ~A266 & ~A265;
  assign \new_[40560]_  = \new_[40559]_  & \new_[40556]_ ;
  assign \new_[40563]_  = A299 & ~A298;
  assign \new_[40566]_  = A301 & A300;
  assign \new_[40567]_  = \new_[40566]_  & \new_[40563]_ ;
  assign \new_[40568]_  = \new_[40567]_  & \new_[40560]_ ;
  assign \new_[40572]_  = ~A167 & A168;
  assign \new_[40573]_  = A169 & \new_[40572]_ ;
  assign \new_[40576]_  = ~A232 & A166;
  assign \new_[40579]_  = ~A234 & A233;
  assign \new_[40580]_  = \new_[40579]_  & \new_[40576]_ ;
  assign \new_[40581]_  = \new_[40580]_  & \new_[40573]_ ;
  assign \new_[40584]_  = A236 & ~A235;
  assign \new_[40587]_  = ~A266 & ~A265;
  assign \new_[40588]_  = \new_[40587]_  & \new_[40584]_ ;
  assign \new_[40591]_  = A299 & ~A298;
  assign \new_[40594]_  = ~A302 & A300;
  assign \new_[40595]_  = \new_[40594]_  & \new_[40591]_ ;
  assign \new_[40596]_  = \new_[40595]_  & \new_[40588]_ ;
  assign \new_[40600]_  = ~A167 & A168;
  assign \new_[40601]_  = A169 & \new_[40600]_ ;
  assign \new_[40604]_  = A232 & A166;
  assign \new_[40607]_  = A234 & ~A233;
  assign \new_[40608]_  = \new_[40607]_  & \new_[40604]_ ;
  assign \new_[40609]_  = \new_[40608]_  & \new_[40601]_ ;
  assign \new_[40612]_  = A267 & A235;
  assign \new_[40615]_  = A269 & ~A268;
  assign \new_[40616]_  = \new_[40615]_  & \new_[40612]_ ;
  assign \new_[40619]_  = ~A299 & A298;
  assign \new_[40622]_  = A301 & A300;
  assign \new_[40623]_  = \new_[40622]_  & \new_[40619]_ ;
  assign \new_[40624]_  = \new_[40623]_  & \new_[40616]_ ;
  assign \new_[40628]_  = ~A167 & A168;
  assign \new_[40629]_  = A169 & \new_[40628]_ ;
  assign \new_[40632]_  = A232 & A166;
  assign \new_[40635]_  = A234 & ~A233;
  assign \new_[40636]_  = \new_[40635]_  & \new_[40632]_ ;
  assign \new_[40637]_  = \new_[40636]_  & \new_[40629]_ ;
  assign \new_[40640]_  = A267 & A235;
  assign \new_[40643]_  = A269 & ~A268;
  assign \new_[40644]_  = \new_[40643]_  & \new_[40640]_ ;
  assign \new_[40647]_  = ~A299 & A298;
  assign \new_[40650]_  = ~A302 & A300;
  assign \new_[40651]_  = \new_[40650]_  & \new_[40647]_ ;
  assign \new_[40652]_  = \new_[40651]_  & \new_[40644]_ ;
  assign \new_[40656]_  = ~A167 & A168;
  assign \new_[40657]_  = A169 & \new_[40656]_ ;
  assign \new_[40660]_  = A232 & A166;
  assign \new_[40663]_  = A234 & ~A233;
  assign \new_[40664]_  = \new_[40663]_  & \new_[40660]_ ;
  assign \new_[40665]_  = \new_[40664]_  & \new_[40657]_ ;
  assign \new_[40668]_  = A267 & A235;
  assign \new_[40671]_  = A269 & ~A268;
  assign \new_[40672]_  = \new_[40671]_  & \new_[40668]_ ;
  assign \new_[40675]_  = A299 & ~A298;
  assign \new_[40678]_  = A301 & A300;
  assign \new_[40679]_  = \new_[40678]_  & \new_[40675]_ ;
  assign \new_[40680]_  = \new_[40679]_  & \new_[40672]_ ;
  assign \new_[40684]_  = ~A167 & A168;
  assign \new_[40685]_  = A169 & \new_[40684]_ ;
  assign \new_[40688]_  = A232 & A166;
  assign \new_[40691]_  = A234 & ~A233;
  assign \new_[40692]_  = \new_[40691]_  & \new_[40688]_ ;
  assign \new_[40693]_  = \new_[40692]_  & \new_[40685]_ ;
  assign \new_[40696]_  = A267 & A235;
  assign \new_[40699]_  = A269 & ~A268;
  assign \new_[40700]_  = \new_[40699]_  & \new_[40696]_ ;
  assign \new_[40703]_  = A299 & ~A298;
  assign \new_[40706]_  = ~A302 & A300;
  assign \new_[40707]_  = \new_[40706]_  & \new_[40703]_ ;
  assign \new_[40708]_  = \new_[40707]_  & \new_[40700]_ ;
  assign \new_[40712]_  = ~A167 & A168;
  assign \new_[40713]_  = A169 & \new_[40712]_ ;
  assign \new_[40716]_  = A232 & A166;
  assign \new_[40719]_  = A234 & ~A233;
  assign \new_[40720]_  = \new_[40719]_  & \new_[40716]_ ;
  assign \new_[40721]_  = \new_[40720]_  & \new_[40713]_ ;
  assign \new_[40724]_  = ~A267 & A235;
  assign \new_[40727]_  = A298 & A268;
  assign \new_[40728]_  = \new_[40727]_  & \new_[40724]_ ;
  assign \new_[40731]_  = ~A300 & ~A299;
  assign \new_[40734]_  = A302 & ~A301;
  assign \new_[40735]_  = \new_[40734]_  & \new_[40731]_ ;
  assign \new_[40736]_  = \new_[40735]_  & \new_[40728]_ ;
  assign \new_[40740]_  = ~A167 & A168;
  assign \new_[40741]_  = A169 & \new_[40740]_ ;
  assign \new_[40744]_  = A232 & A166;
  assign \new_[40747]_  = A234 & ~A233;
  assign \new_[40748]_  = \new_[40747]_  & \new_[40744]_ ;
  assign \new_[40749]_  = \new_[40748]_  & \new_[40741]_ ;
  assign \new_[40752]_  = ~A267 & A235;
  assign \new_[40755]_  = ~A298 & A268;
  assign \new_[40756]_  = \new_[40755]_  & \new_[40752]_ ;
  assign \new_[40759]_  = ~A300 & A299;
  assign \new_[40762]_  = A302 & ~A301;
  assign \new_[40763]_  = \new_[40762]_  & \new_[40759]_ ;
  assign \new_[40764]_  = \new_[40763]_  & \new_[40756]_ ;
  assign \new_[40768]_  = ~A167 & A168;
  assign \new_[40769]_  = A169 & \new_[40768]_ ;
  assign \new_[40772]_  = A232 & A166;
  assign \new_[40775]_  = A234 & ~A233;
  assign \new_[40776]_  = \new_[40775]_  & \new_[40772]_ ;
  assign \new_[40777]_  = \new_[40776]_  & \new_[40769]_ ;
  assign \new_[40780]_  = ~A267 & A235;
  assign \new_[40783]_  = A298 & ~A269;
  assign \new_[40784]_  = \new_[40783]_  & \new_[40780]_ ;
  assign \new_[40787]_  = ~A300 & ~A299;
  assign \new_[40790]_  = A302 & ~A301;
  assign \new_[40791]_  = \new_[40790]_  & \new_[40787]_ ;
  assign \new_[40792]_  = \new_[40791]_  & \new_[40784]_ ;
  assign \new_[40796]_  = ~A167 & A168;
  assign \new_[40797]_  = A169 & \new_[40796]_ ;
  assign \new_[40800]_  = A232 & A166;
  assign \new_[40803]_  = A234 & ~A233;
  assign \new_[40804]_  = \new_[40803]_  & \new_[40800]_ ;
  assign \new_[40805]_  = \new_[40804]_  & \new_[40797]_ ;
  assign \new_[40808]_  = ~A267 & A235;
  assign \new_[40811]_  = ~A298 & ~A269;
  assign \new_[40812]_  = \new_[40811]_  & \new_[40808]_ ;
  assign \new_[40815]_  = ~A300 & A299;
  assign \new_[40818]_  = A302 & ~A301;
  assign \new_[40819]_  = \new_[40818]_  & \new_[40815]_ ;
  assign \new_[40820]_  = \new_[40819]_  & \new_[40812]_ ;
  assign \new_[40824]_  = ~A167 & A168;
  assign \new_[40825]_  = A169 & \new_[40824]_ ;
  assign \new_[40828]_  = A232 & A166;
  assign \new_[40831]_  = A234 & ~A233;
  assign \new_[40832]_  = \new_[40831]_  & \new_[40828]_ ;
  assign \new_[40833]_  = \new_[40832]_  & \new_[40825]_ ;
  assign \new_[40836]_  = A265 & A235;
  assign \new_[40839]_  = A298 & A266;
  assign \new_[40840]_  = \new_[40839]_  & \new_[40836]_ ;
  assign \new_[40843]_  = ~A300 & ~A299;
  assign \new_[40846]_  = A302 & ~A301;
  assign \new_[40847]_  = \new_[40846]_  & \new_[40843]_ ;
  assign \new_[40848]_  = \new_[40847]_  & \new_[40840]_ ;
  assign \new_[40852]_  = ~A167 & A168;
  assign \new_[40853]_  = A169 & \new_[40852]_ ;
  assign \new_[40856]_  = A232 & A166;
  assign \new_[40859]_  = A234 & ~A233;
  assign \new_[40860]_  = \new_[40859]_  & \new_[40856]_ ;
  assign \new_[40861]_  = \new_[40860]_  & \new_[40853]_ ;
  assign \new_[40864]_  = A265 & A235;
  assign \new_[40867]_  = ~A298 & A266;
  assign \new_[40868]_  = \new_[40867]_  & \new_[40864]_ ;
  assign \new_[40871]_  = ~A300 & A299;
  assign \new_[40874]_  = A302 & ~A301;
  assign \new_[40875]_  = \new_[40874]_  & \new_[40871]_ ;
  assign \new_[40876]_  = \new_[40875]_  & \new_[40868]_ ;
  assign \new_[40880]_  = ~A167 & A168;
  assign \new_[40881]_  = A169 & \new_[40880]_ ;
  assign \new_[40884]_  = A232 & A166;
  assign \new_[40887]_  = A234 & ~A233;
  assign \new_[40888]_  = \new_[40887]_  & \new_[40884]_ ;
  assign \new_[40889]_  = \new_[40888]_  & \new_[40881]_ ;
  assign \new_[40892]_  = ~A265 & A235;
  assign \new_[40895]_  = A298 & ~A266;
  assign \new_[40896]_  = \new_[40895]_  & \new_[40892]_ ;
  assign \new_[40899]_  = ~A300 & ~A299;
  assign \new_[40902]_  = A302 & ~A301;
  assign \new_[40903]_  = \new_[40902]_  & \new_[40899]_ ;
  assign \new_[40904]_  = \new_[40903]_  & \new_[40896]_ ;
  assign \new_[40908]_  = ~A167 & A168;
  assign \new_[40909]_  = A169 & \new_[40908]_ ;
  assign \new_[40912]_  = A232 & A166;
  assign \new_[40915]_  = A234 & ~A233;
  assign \new_[40916]_  = \new_[40915]_  & \new_[40912]_ ;
  assign \new_[40917]_  = \new_[40916]_  & \new_[40909]_ ;
  assign \new_[40920]_  = ~A265 & A235;
  assign \new_[40923]_  = ~A298 & ~A266;
  assign \new_[40924]_  = \new_[40923]_  & \new_[40920]_ ;
  assign \new_[40927]_  = ~A300 & A299;
  assign \new_[40930]_  = A302 & ~A301;
  assign \new_[40931]_  = \new_[40930]_  & \new_[40927]_ ;
  assign \new_[40932]_  = \new_[40931]_  & \new_[40924]_ ;
  assign \new_[40936]_  = ~A167 & A168;
  assign \new_[40937]_  = A169 & \new_[40936]_ ;
  assign \new_[40940]_  = A232 & A166;
  assign \new_[40943]_  = A234 & ~A233;
  assign \new_[40944]_  = \new_[40943]_  & \new_[40940]_ ;
  assign \new_[40945]_  = \new_[40944]_  & \new_[40937]_ ;
  assign \new_[40948]_  = A267 & ~A236;
  assign \new_[40951]_  = A269 & ~A268;
  assign \new_[40952]_  = \new_[40951]_  & \new_[40948]_ ;
  assign \new_[40955]_  = ~A299 & A298;
  assign \new_[40958]_  = A301 & A300;
  assign \new_[40959]_  = \new_[40958]_  & \new_[40955]_ ;
  assign \new_[40960]_  = \new_[40959]_  & \new_[40952]_ ;
  assign \new_[40964]_  = ~A167 & A168;
  assign \new_[40965]_  = A169 & \new_[40964]_ ;
  assign \new_[40968]_  = A232 & A166;
  assign \new_[40971]_  = A234 & ~A233;
  assign \new_[40972]_  = \new_[40971]_  & \new_[40968]_ ;
  assign \new_[40973]_  = \new_[40972]_  & \new_[40965]_ ;
  assign \new_[40976]_  = A267 & ~A236;
  assign \new_[40979]_  = A269 & ~A268;
  assign \new_[40980]_  = \new_[40979]_  & \new_[40976]_ ;
  assign \new_[40983]_  = ~A299 & A298;
  assign \new_[40986]_  = ~A302 & A300;
  assign \new_[40987]_  = \new_[40986]_  & \new_[40983]_ ;
  assign \new_[40988]_  = \new_[40987]_  & \new_[40980]_ ;
  assign \new_[40992]_  = ~A167 & A168;
  assign \new_[40993]_  = A169 & \new_[40992]_ ;
  assign \new_[40996]_  = A232 & A166;
  assign \new_[40999]_  = A234 & ~A233;
  assign \new_[41000]_  = \new_[40999]_  & \new_[40996]_ ;
  assign \new_[41001]_  = \new_[41000]_  & \new_[40993]_ ;
  assign \new_[41004]_  = A267 & ~A236;
  assign \new_[41007]_  = A269 & ~A268;
  assign \new_[41008]_  = \new_[41007]_  & \new_[41004]_ ;
  assign \new_[41011]_  = A299 & ~A298;
  assign \new_[41014]_  = A301 & A300;
  assign \new_[41015]_  = \new_[41014]_  & \new_[41011]_ ;
  assign \new_[41016]_  = \new_[41015]_  & \new_[41008]_ ;
  assign \new_[41020]_  = ~A167 & A168;
  assign \new_[41021]_  = A169 & \new_[41020]_ ;
  assign \new_[41024]_  = A232 & A166;
  assign \new_[41027]_  = A234 & ~A233;
  assign \new_[41028]_  = \new_[41027]_  & \new_[41024]_ ;
  assign \new_[41029]_  = \new_[41028]_  & \new_[41021]_ ;
  assign \new_[41032]_  = A267 & ~A236;
  assign \new_[41035]_  = A269 & ~A268;
  assign \new_[41036]_  = \new_[41035]_  & \new_[41032]_ ;
  assign \new_[41039]_  = A299 & ~A298;
  assign \new_[41042]_  = ~A302 & A300;
  assign \new_[41043]_  = \new_[41042]_  & \new_[41039]_ ;
  assign \new_[41044]_  = \new_[41043]_  & \new_[41036]_ ;
  assign \new_[41048]_  = ~A167 & A168;
  assign \new_[41049]_  = A169 & \new_[41048]_ ;
  assign \new_[41052]_  = A232 & A166;
  assign \new_[41055]_  = A234 & ~A233;
  assign \new_[41056]_  = \new_[41055]_  & \new_[41052]_ ;
  assign \new_[41057]_  = \new_[41056]_  & \new_[41049]_ ;
  assign \new_[41060]_  = ~A267 & ~A236;
  assign \new_[41063]_  = A298 & A268;
  assign \new_[41064]_  = \new_[41063]_  & \new_[41060]_ ;
  assign \new_[41067]_  = ~A300 & ~A299;
  assign \new_[41070]_  = A302 & ~A301;
  assign \new_[41071]_  = \new_[41070]_  & \new_[41067]_ ;
  assign \new_[41072]_  = \new_[41071]_  & \new_[41064]_ ;
  assign \new_[41076]_  = ~A167 & A168;
  assign \new_[41077]_  = A169 & \new_[41076]_ ;
  assign \new_[41080]_  = A232 & A166;
  assign \new_[41083]_  = A234 & ~A233;
  assign \new_[41084]_  = \new_[41083]_  & \new_[41080]_ ;
  assign \new_[41085]_  = \new_[41084]_  & \new_[41077]_ ;
  assign \new_[41088]_  = ~A267 & ~A236;
  assign \new_[41091]_  = ~A298 & A268;
  assign \new_[41092]_  = \new_[41091]_  & \new_[41088]_ ;
  assign \new_[41095]_  = ~A300 & A299;
  assign \new_[41098]_  = A302 & ~A301;
  assign \new_[41099]_  = \new_[41098]_  & \new_[41095]_ ;
  assign \new_[41100]_  = \new_[41099]_  & \new_[41092]_ ;
  assign \new_[41104]_  = ~A167 & A168;
  assign \new_[41105]_  = A169 & \new_[41104]_ ;
  assign \new_[41108]_  = A232 & A166;
  assign \new_[41111]_  = A234 & ~A233;
  assign \new_[41112]_  = \new_[41111]_  & \new_[41108]_ ;
  assign \new_[41113]_  = \new_[41112]_  & \new_[41105]_ ;
  assign \new_[41116]_  = ~A267 & ~A236;
  assign \new_[41119]_  = A298 & ~A269;
  assign \new_[41120]_  = \new_[41119]_  & \new_[41116]_ ;
  assign \new_[41123]_  = ~A300 & ~A299;
  assign \new_[41126]_  = A302 & ~A301;
  assign \new_[41127]_  = \new_[41126]_  & \new_[41123]_ ;
  assign \new_[41128]_  = \new_[41127]_  & \new_[41120]_ ;
  assign \new_[41132]_  = ~A167 & A168;
  assign \new_[41133]_  = A169 & \new_[41132]_ ;
  assign \new_[41136]_  = A232 & A166;
  assign \new_[41139]_  = A234 & ~A233;
  assign \new_[41140]_  = \new_[41139]_  & \new_[41136]_ ;
  assign \new_[41141]_  = \new_[41140]_  & \new_[41133]_ ;
  assign \new_[41144]_  = ~A267 & ~A236;
  assign \new_[41147]_  = ~A298 & ~A269;
  assign \new_[41148]_  = \new_[41147]_  & \new_[41144]_ ;
  assign \new_[41151]_  = ~A300 & A299;
  assign \new_[41154]_  = A302 & ~A301;
  assign \new_[41155]_  = \new_[41154]_  & \new_[41151]_ ;
  assign \new_[41156]_  = \new_[41155]_  & \new_[41148]_ ;
  assign \new_[41160]_  = ~A167 & A168;
  assign \new_[41161]_  = A169 & \new_[41160]_ ;
  assign \new_[41164]_  = A232 & A166;
  assign \new_[41167]_  = A234 & ~A233;
  assign \new_[41168]_  = \new_[41167]_  & \new_[41164]_ ;
  assign \new_[41169]_  = \new_[41168]_  & \new_[41161]_ ;
  assign \new_[41172]_  = A265 & ~A236;
  assign \new_[41175]_  = A298 & A266;
  assign \new_[41176]_  = \new_[41175]_  & \new_[41172]_ ;
  assign \new_[41179]_  = ~A300 & ~A299;
  assign \new_[41182]_  = A302 & ~A301;
  assign \new_[41183]_  = \new_[41182]_  & \new_[41179]_ ;
  assign \new_[41184]_  = \new_[41183]_  & \new_[41176]_ ;
  assign \new_[41188]_  = ~A167 & A168;
  assign \new_[41189]_  = A169 & \new_[41188]_ ;
  assign \new_[41192]_  = A232 & A166;
  assign \new_[41195]_  = A234 & ~A233;
  assign \new_[41196]_  = \new_[41195]_  & \new_[41192]_ ;
  assign \new_[41197]_  = \new_[41196]_  & \new_[41189]_ ;
  assign \new_[41200]_  = A265 & ~A236;
  assign \new_[41203]_  = ~A298 & A266;
  assign \new_[41204]_  = \new_[41203]_  & \new_[41200]_ ;
  assign \new_[41207]_  = ~A300 & A299;
  assign \new_[41210]_  = A302 & ~A301;
  assign \new_[41211]_  = \new_[41210]_  & \new_[41207]_ ;
  assign \new_[41212]_  = \new_[41211]_  & \new_[41204]_ ;
  assign \new_[41216]_  = ~A167 & A168;
  assign \new_[41217]_  = A169 & \new_[41216]_ ;
  assign \new_[41220]_  = A232 & A166;
  assign \new_[41223]_  = A234 & ~A233;
  assign \new_[41224]_  = \new_[41223]_  & \new_[41220]_ ;
  assign \new_[41225]_  = \new_[41224]_  & \new_[41217]_ ;
  assign \new_[41228]_  = ~A265 & ~A236;
  assign \new_[41231]_  = A298 & ~A266;
  assign \new_[41232]_  = \new_[41231]_  & \new_[41228]_ ;
  assign \new_[41235]_  = ~A300 & ~A299;
  assign \new_[41238]_  = A302 & ~A301;
  assign \new_[41239]_  = \new_[41238]_  & \new_[41235]_ ;
  assign \new_[41240]_  = \new_[41239]_  & \new_[41232]_ ;
  assign \new_[41244]_  = ~A167 & A168;
  assign \new_[41245]_  = A169 & \new_[41244]_ ;
  assign \new_[41248]_  = A232 & A166;
  assign \new_[41251]_  = A234 & ~A233;
  assign \new_[41252]_  = \new_[41251]_  & \new_[41248]_ ;
  assign \new_[41253]_  = \new_[41252]_  & \new_[41245]_ ;
  assign \new_[41256]_  = ~A265 & ~A236;
  assign \new_[41259]_  = ~A298 & ~A266;
  assign \new_[41260]_  = \new_[41259]_  & \new_[41256]_ ;
  assign \new_[41263]_  = ~A300 & A299;
  assign \new_[41266]_  = A302 & ~A301;
  assign \new_[41267]_  = \new_[41266]_  & \new_[41263]_ ;
  assign \new_[41268]_  = \new_[41267]_  & \new_[41260]_ ;
  assign \new_[41272]_  = ~A167 & A168;
  assign \new_[41273]_  = A169 & \new_[41272]_ ;
  assign \new_[41276]_  = A232 & A166;
  assign \new_[41279]_  = ~A234 & ~A233;
  assign \new_[41280]_  = \new_[41279]_  & \new_[41276]_ ;
  assign \new_[41281]_  = \new_[41280]_  & \new_[41273]_ ;
  assign \new_[41284]_  = A236 & ~A235;
  assign \new_[41287]_  = A268 & ~A267;
  assign \new_[41288]_  = \new_[41287]_  & \new_[41284]_ ;
  assign \new_[41291]_  = ~A299 & A298;
  assign \new_[41294]_  = A301 & A300;
  assign \new_[41295]_  = \new_[41294]_  & \new_[41291]_ ;
  assign \new_[41296]_  = \new_[41295]_  & \new_[41288]_ ;
  assign \new_[41300]_  = ~A167 & A168;
  assign \new_[41301]_  = A169 & \new_[41300]_ ;
  assign \new_[41304]_  = A232 & A166;
  assign \new_[41307]_  = ~A234 & ~A233;
  assign \new_[41308]_  = \new_[41307]_  & \new_[41304]_ ;
  assign \new_[41309]_  = \new_[41308]_  & \new_[41301]_ ;
  assign \new_[41312]_  = A236 & ~A235;
  assign \new_[41315]_  = A268 & ~A267;
  assign \new_[41316]_  = \new_[41315]_  & \new_[41312]_ ;
  assign \new_[41319]_  = ~A299 & A298;
  assign \new_[41322]_  = ~A302 & A300;
  assign \new_[41323]_  = \new_[41322]_  & \new_[41319]_ ;
  assign \new_[41324]_  = \new_[41323]_  & \new_[41316]_ ;
  assign \new_[41328]_  = ~A167 & A168;
  assign \new_[41329]_  = A169 & \new_[41328]_ ;
  assign \new_[41332]_  = A232 & A166;
  assign \new_[41335]_  = ~A234 & ~A233;
  assign \new_[41336]_  = \new_[41335]_  & \new_[41332]_ ;
  assign \new_[41337]_  = \new_[41336]_  & \new_[41329]_ ;
  assign \new_[41340]_  = A236 & ~A235;
  assign \new_[41343]_  = A268 & ~A267;
  assign \new_[41344]_  = \new_[41343]_  & \new_[41340]_ ;
  assign \new_[41347]_  = A299 & ~A298;
  assign \new_[41350]_  = A301 & A300;
  assign \new_[41351]_  = \new_[41350]_  & \new_[41347]_ ;
  assign \new_[41352]_  = \new_[41351]_  & \new_[41344]_ ;
  assign \new_[41356]_  = ~A167 & A168;
  assign \new_[41357]_  = A169 & \new_[41356]_ ;
  assign \new_[41360]_  = A232 & A166;
  assign \new_[41363]_  = ~A234 & ~A233;
  assign \new_[41364]_  = \new_[41363]_  & \new_[41360]_ ;
  assign \new_[41365]_  = \new_[41364]_  & \new_[41357]_ ;
  assign \new_[41368]_  = A236 & ~A235;
  assign \new_[41371]_  = A268 & ~A267;
  assign \new_[41372]_  = \new_[41371]_  & \new_[41368]_ ;
  assign \new_[41375]_  = A299 & ~A298;
  assign \new_[41378]_  = ~A302 & A300;
  assign \new_[41379]_  = \new_[41378]_  & \new_[41375]_ ;
  assign \new_[41380]_  = \new_[41379]_  & \new_[41372]_ ;
  assign \new_[41384]_  = ~A167 & A168;
  assign \new_[41385]_  = A169 & \new_[41384]_ ;
  assign \new_[41388]_  = A232 & A166;
  assign \new_[41391]_  = ~A234 & ~A233;
  assign \new_[41392]_  = \new_[41391]_  & \new_[41388]_ ;
  assign \new_[41393]_  = \new_[41392]_  & \new_[41385]_ ;
  assign \new_[41396]_  = A236 & ~A235;
  assign \new_[41399]_  = ~A269 & ~A267;
  assign \new_[41400]_  = \new_[41399]_  & \new_[41396]_ ;
  assign \new_[41403]_  = ~A299 & A298;
  assign \new_[41406]_  = A301 & A300;
  assign \new_[41407]_  = \new_[41406]_  & \new_[41403]_ ;
  assign \new_[41408]_  = \new_[41407]_  & \new_[41400]_ ;
  assign \new_[41412]_  = ~A167 & A168;
  assign \new_[41413]_  = A169 & \new_[41412]_ ;
  assign \new_[41416]_  = A232 & A166;
  assign \new_[41419]_  = ~A234 & ~A233;
  assign \new_[41420]_  = \new_[41419]_  & \new_[41416]_ ;
  assign \new_[41421]_  = \new_[41420]_  & \new_[41413]_ ;
  assign \new_[41424]_  = A236 & ~A235;
  assign \new_[41427]_  = ~A269 & ~A267;
  assign \new_[41428]_  = \new_[41427]_  & \new_[41424]_ ;
  assign \new_[41431]_  = ~A299 & A298;
  assign \new_[41434]_  = ~A302 & A300;
  assign \new_[41435]_  = \new_[41434]_  & \new_[41431]_ ;
  assign \new_[41436]_  = \new_[41435]_  & \new_[41428]_ ;
  assign \new_[41440]_  = ~A167 & A168;
  assign \new_[41441]_  = A169 & \new_[41440]_ ;
  assign \new_[41444]_  = A232 & A166;
  assign \new_[41447]_  = ~A234 & ~A233;
  assign \new_[41448]_  = \new_[41447]_  & \new_[41444]_ ;
  assign \new_[41449]_  = \new_[41448]_  & \new_[41441]_ ;
  assign \new_[41452]_  = A236 & ~A235;
  assign \new_[41455]_  = ~A269 & ~A267;
  assign \new_[41456]_  = \new_[41455]_  & \new_[41452]_ ;
  assign \new_[41459]_  = A299 & ~A298;
  assign \new_[41462]_  = A301 & A300;
  assign \new_[41463]_  = \new_[41462]_  & \new_[41459]_ ;
  assign \new_[41464]_  = \new_[41463]_  & \new_[41456]_ ;
  assign \new_[41468]_  = ~A167 & A168;
  assign \new_[41469]_  = A169 & \new_[41468]_ ;
  assign \new_[41472]_  = A232 & A166;
  assign \new_[41475]_  = ~A234 & ~A233;
  assign \new_[41476]_  = \new_[41475]_  & \new_[41472]_ ;
  assign \new_[41477]_  = \new_[41476]_  & \new_[41469]_ ;
  assign \new_[41480]_  = A236 & ~A235;
  assign \new_[41483]_  = ~A269 & ~A267;
  assign \new_[41484]_  = \new_[41483]_  & \new_[41480]_ ;
  assign \new_[41487]_  = A299 & ~A298;
  assign \new_[41490]_  = ~A302 & A300;
  assign \new_[41491]_  = \new_[41490]_  & \new_[41487]_ ;
  assign \new_[41492]_  = \new_[41491]_  & \new_[41484]_ ;
  assign \new_[41496]_  = ~A167 & A168;
  assign \new_[41497]_  = A169 & \new_[41496]_ ;
  assign \new_[41500]_  = A232 & A166;
  assign \new_[41503]_  = ~A234 & ~A233;
  assign \new_[41504]_  = \new_[41503]_  & \new_[41500]_ ;
  assign \new_[41505]_  = \new_[41504]_  & \new_[41497]_ ;
  assign \new_[41508]_  = A236 & ~A235;
  assign \new_[41511]_  = A266 & A265;
  assign \new_[41512]_  = \new_[41511]_  & \new_[41508]_ ;
  assign \new_[41515]_  = ~A299 & A298;
  assign \new_[41518]_  = A301 & A300;
  assign \new_[41519]_  = \new_[41518]_  & \new_[41515]_ ;
  assign \new_[41520]_  = \new_[41519]_  & \new_[41512]_ ;
  assign \new_[41524]_  = ~A167 & A168;
  assign \new_[41525]_  = A169 & \new_[41524]_ ;
  assign \new_[41528]_  = A232 & A166;
  assign \new_[41531]_  = ~A234 & ~A233;
  assign \new_[41532]_  = \new_[41531]_  & \new_[41528]_ ;
  assign \new_[41533]_  = \new_[41532]_  & \new_[41525]_ ;
  assign \new_[41536]_  = A236 & ~A235;
  assign \new_[41539]_  = A266 & A265;
  assign \new_[41540]_  = \new_[41539]_  & \new_[41536]_ ;
  assign \new_[41543]_  = ~A299 & A298;
  assign \new_[41546]_  = ~A302 & A300;
  assign \new_[41547]_  = \new_[41546]_  & \new_[41543]_ ;
  assign \new_[41548]_  = \new_[41547]_  & \new_[41540]_ ;
  assign \new_[41552]_  = ~A167 & A168;
  assign \new_[41553]_  = A169 & \new_[41552]_ ;
  assign \new_[41556]_  = A232 & A166;
  assign \new_[41559]_  = ~A234 & ~A233;
  assign \new_[41560]_  = \new_[41559]_  & \new_[41556]_ ;
  assign \new_[41561]_  = \new_[41560]_  & \new_[41553]_ ;
  assign \new_[41564]_  = A236 & ~A235;
  assign \new_[41567]_  = A266 & A265;
  assign \new_[41568]_  = \new_[41567]_  & \new_[41564]_ ;
  assign \new_[41571]_  = A299 & ~A298;
  assign \new_[41574]_  = A301 & A300;
  assign \new_[41575]_  = \new_[41574]_  & \new_[41571]_ ;
  assign \new_[41576]_  = \new_[41575]_  & \new_[41568]_ ;
  assign \new_[41580]_  = ~A167 & A168;
  assign \new_[41581]_  = A169 & \new_[41580]_ ;
  assign \new_[41584]_  = A232 & A166;
  assign \new_[41587]_  = ~A234 & ~A233;
  assign \new_[41588]_  = \new_[41587]_  & \new_[41584]_ ;
  assign \new_[41589]_  = \new_[41588]_  & \new_[41581]_ ;
  assign \new_[41592]_  = A236 & ~A235;
  assign \new_[41595]_  = A266 & A265;
  assign \new_[41596]_  = \new_[41595]_  & \new_[41592]_ ;
  assign \new_[41599]_  = A299 & ~A298;
  assign \new_[41602]_  = ~A302 & A300;
  assign \new_[41603]_  = \new_[41602]_  & \new_[41599]_ ;
  assign \new_[41604]_  = \new_[41603]_  & \new_[41596]_ ;
  assign \new_[41608]_  = ~A167 & A168;
  assign \new_[41609]_  = A169 & \new_[41608]_ ;
  assign \new_[41612]_  = A232 & A166;
  assign \new_[41615]_  = ~A234 & ~A233;
  assign \new_[41616]_  = \new_[41615]_  & \new_[41612]_ ;
  assign \new_[41617]_  = \new_[41616]_  & \new_[41609]_ ;
  assign \new_[41620]_  = A236 & ~A235;
  assign \new_[41623]_  = ~A266 & ~A265;
  assign \new_[41624]_  = \new_[41623]_  & \new_[41620]_ ;
  assign \new_[41627]_  = ~A299 & A298;
  assign \new_[41630]_  = A301 & A300;
  assign \new_[41631]_  = \new_[41630]_  & \new_[41627]_ ;
  assign \new_[41632]_  = \new_[41631]_  & \new_[41624]_ ;
  assign \new_[41636]_  = ~A167 & A168;
  assign \new_[41637]_  = A169 & \new_[41636]_ ;
  assign \new_[41640]_  = A232 & A166;
  assign \new_[41643]_  = ~A234 & ~A233;
  assign \new_[41644]_  = \new_[41643]_  & \new_[41640]_ ;
  assign \new_[41645]_  = \new_[41644]_  & \new_[41637]_ ;
  assign \new_[41648]_  = A236 & ~A235;
  assign \new_[41651]_  = ~A266 & ~A265;
  assign \new_[41652]_  = \new_[41651]_  & \new_[41648]_ ;
  assign \new_[41655]_  = ~A299 & A298;
  assign \new_[41658]_  = ~A302 & A300;
  assign \new_[41659]_  = \new_[41658]_  & \new_[41655]_ ;
  assign \new_[41660]_  = \new_[41659]_  & \new_[41652]_ ;
  assign \new_[41664]_  = ~A167 & A168;
  assign \new_[41665]_  = A169 & \new_[41664]_ ;
  assign \new_[41668]_  = A232 & A166;
  assign \new_[41671]_  = ~A234 & ~A233;
  assign \new_[41672]_  = \new_[41671]_  & \new_[41668]_ ;
  assign \new_[41673]_  = \new_[41672]_  & \new_[41665]_ ;
  assign \new_[41676]_  = A236 & ~A235;
  assign \new_[41679]_  = ~A266 & ~A265;
  assign \new_[41680]_  = \new_[41679]_  & \new_[41676]_ ;
  assign \new_[41683]_  = A299 & ~A298;
  assign \new_[41686]_  = A301 & A300;
  assign \new_[41687]_  = \new_[41686]_  & \new_[41683]_ ;
  assign \new_[41688]_  = \new_[41687]_  & \new_[41680]_ ;
  assign \new_[41692]_  = ~A167 & A168;
  assign \new_[41693]_  = A169 & \new_[41692]_ ;
  assign \new_[41696]_  = A232 & A166;
  assign \new_[41699]_  = ~A234 & ~A233;
  assign \new_[41700]_  = \new_[41699]_  & \new_[41696]_ ;
  assign \new_[41701]_  = \new_[41700]_  & \new_[41693]_ ;
  assign \new_[41704]_  = A236 & ~A235;
  assign \new_[41707]_  = ~A266 & ~A265;
  assign \new_[41708]_  = \new_[41707]_  & \new_[41704]_ ;
  assign \new_[41711]_  = A299 & ~A298;
  assign \new_[41714]_  = ~A302 & A300;
  assign \new_[41715]_  = \new_[41714]_  & \new_[41711]_ ;
  assign \new_[41716]_  = \new_[41715]_  & \new_[41708]_ ;
  assign \new_[41720]_  = ~A168 & ~A169;
  assign \new_[41721]_  = ~A170 & \new_[41720]_ ;
  assign \new_[41724]_  = ~A166 & A167;
  assign \new_[41727]_  = A233 & ~A232;
  assign \new_[41728]_  = \new_[41727]_  & \new_[41724]_ ;
  assign \new_[41729]_  = \new_[41728]_  & \new_[41721]_ ;
  assign \new_[41732]_  = A235 & A234;
  assign \new_[41735]_  = A268 & ~A267;
  assign \new_[41736]_  = \new_[41735]_  & \new_[41732]_ ;
  assign \new_[41739]_  = ~A299 & A298;
  assign \new_[41742]_  = A301 & A300;
  assign \new_[41743]_  = \new_[41742]_  & \new_[41739]_ ;
  assign \new_[41744]_  = \new_[41743]_  & \new_[41736]_ ;
  assign \new_[41748]_  = ~A168 & ~A169;
  assign \new_[41749]_  = ~A170 & \new_[41748]_ ;
  assign \new_[41752]_  = ~A166 & A167;
  assign \new_[41755]_  = A233 & ~A232;
  assign \new_[41756]_  = \new_[41755]_  & \new_[41752]_ ;
  assign \new_[41757]_  = \new_[41756]_  & \new_[41749]_ ;
  assign \new_[41760]_  = A235 & A234;
  assign \new_[41763]_  = A268 & ~A267;
  assign \new_[41764]_  = \new_[41763]_  & \new_[41760]_ ;
  assign \new_[41767]_  = ~A299 & A298;
  assign \new_[41770]_  = ~A302 & A300;
  assign \new_[41771]_  = \new_[41770]_  & \new_[41767]_ ;
  assign \new_[41772]_  = \new_[41771]_  & \new_[41764]_ ;
  assign \new_[41776]_  = ~A168 & ~A169;
  assign \new_[41777]_  = ~A170 & \new_[41776]_ ;
  assign \new_[41780]_  = ~A166 & A167;
  assign \new_[41783]_  = A233 & ~A232;
  assign \new_[41784]_  = \new_[41783]_  & \new_[41780]_ ;
  assign \new_[41785]_  = \new_[41784]_  & \new_[41777]_ ;
  assign \new_[41788]_  = A235 & A234;
  assign \new_[41791]_  = A268 & ~A267;
  assign \new_[41792]_  = \new_[41791]_  & \new_[41788]_ ;
  assign \new_[41795]_  = A299 & ~A298;
  assign \new_[41798]_  = A301 & A300;
  assign \new_[41799]_  = \new_[41798]_  & \new_[41795]_ ;
  assign \new_[41800]_  = \new_[41799]_  & \new_[41792]_ ;
  assign \new_[41804]_  = ~A168 & ~A169;
  assign \new_[41805]_  = ~A170 & \new_[41804]_ ;
  assign \new_[41808]_  = ~A166 & A167;
  assign \new_[41811]_  = A233 & ~A232;
  assign \new_[41812]_  = \new_[41811]_  & \new_[41808]_ ;
  assign \new_[41813]_  = \new_[41812]_  & \new_[41805]_ ;
  assign \new_[41816]_  = A235 & A234;
  assign \new_[41819]_  = A268 & ~A267;
  assign \new_[41820]_  = \new_[41819]_  & \new_[41816]_ ;
  assign \new_[41823]_  = A299 & ~A298;
  assign \new_[41826]_  = ~A302 & A300;
  assign \new_[41827]_  = \new_[41826]_  & \new_[41823]_ ;
  assign \new_[41828]_  = \new_[41827]_  & \new_[41820]_ ;
  assign \new_[41832]_  = ~A168 & ~A169;
  assign \new_[41833]_  = ~A170 & \new_[41832]_ ;
  assign \new_[41836]_  = ~A166 & A167;
  assign \new_[41839]_  = A233 & ~A232;
  assign \new_[41840]_  = \new_[41839]_  & \new_[41836]_ ;
  assign \new_[41841]_  = \new_[41840]_  & \new_[41833]_ ;
  assign \new_[41844]_  = A235 & A234;
  assign \new_[41847]_  = ~A269 & ~A267;
  assign \new_[41848]_  = \new_[41847]_  & \new_[41844]_ ;
  assign \new_[41851]_  = ~A299 & A298;
  assign \new_[41854]_  = A301 & A300;
  assign \new_[41855]_  = \new_[41854]_  & \new_[41851]_ ;
  assign \new_[41856]_  = \new_[41855]_  & \new_[41848]_ ;
  assign \new_[41860]_  = ~A168 & ~A169;
  assign \new_[41861]_  = ~A170 & \new_[41860]_ ;
  assign \new_[41864]_  = ~A166 & A167;
  assign \new_[41867]_  = A233 & ~A232;
  assign \new_[41868]_  = \new_[41867]_  & \new_[41864]_ ;
  assign \new_[41869]_  = \new_[41868]_  & \new_[41861]_ ;
  assign \new_[41872]_  = A235 & A234;
  assign \new_[41875]_  = ~A269 & ~A267;
  assign \new_[41876]_  = \new_[41875]_  & \new_[41872]_ ;
  assign \new_[41879]_  = ~A299 & A298;
  assign \new_[41882]_  = ~A302 & A300;
  assign \new_[41883]_  = \new_[41882]_  & \new_[41879]_ ;
  assign \new_[41884]_  = \new_[41883]_  & \new_[41876]_ ;
  assign \new_[41888]_  = ~A168 & ~A169;
  assign \new_[41889]_  = ~A170 & \new_[41888]_ ;
  assign \new_[41892]_  = ~A166 & A167;
  assign \new_[41895]_  = A233 & ~A232;
  assign \new_[41896]_  = \new_[41895]_  & \new_[41892]_ ;
  assign \new_[41897]_  = \new_[41896]_  & \new_[41889]_ ;
  assign \new_[41900]_  = A235 & A234;
  assign \new_[41903]_  = ~A269 & ~A267;
  assign \new_[41904]_  = \new_[41903]_  & \new_[41900]_ ;
  assign \new_[41907]_  = A299 & ~A298;
  assign \new_[41910]_  = A301 & A300;
  assign \new_[41911]_  = \new_[41910]_  & \new_[41907]_ ;
  assign \new_[41912]_  = \new_[41911]_  & \new_[41904]_ ;
  assign \new_[41916]_  = ~A168 & ~A169;
  assign \new_[41917]_  = ~A170 & \new_[41916]_ ;
  assign \new_[41920]_  = ~A166 & A167;
  assign \new_[41923]_  = A233 & ~A232;
  assign \new_[41924]_  = \new_[41923]_  & \new_[41920]_ ;
  assign \new_[41925]_  = \new_[41924]_  & \new_[41917]_ ;
  assign \new_[41928]_  = A235 & A234;
  assign \new_[41931]_  = ~A269 & ~A267;
  assign \new_[41932]_  = \new_[41931]_  & \new_[41928]_ ;
  assign \new_[41935]_  = A299 & ~A298;
  assign \new_[41938]_  = ~A302 & A300;
  assign \new_[41939]_  = \new_[41938]_  & \new_[41935]_ ;
  assign \new_[41940]_  = \new_[41939]_  & \new_[41932]_ ;
  assign \new_[41944]_  = ~A168 & ~A169;
  assign \new_[41945]_  = ~A170 & \new_[41944]_ ;
  assign \new_[41948]_  = ~A166 & A167;
  assign \new_[41951]_  = A233 & ~A232;
  assign \new_[41952]_  = \new_[41951]_  & \new_[41948]_ ;
  assign \new_[41953]_  = \new_[41952]_  & \new_[41945]_ ;
  assign \new_[41956]_  = A235 & A234;
  assign \new_[41959]_  = A266 & A265;
  assign \new_[41960]_  = \new_[41959]_  & \new_[41956]_ ;
  assign \new_[41963]_  = ~A299 & A298;
  assign \new_[41966]_  = A301 & A300;
  assign \new_[41967]_  = \new_[41966]_  & \new_[41963]_ ;
  assign \new_[41968]_  = \new_[41967]_  & \new_[41960]_ ;
  assign \new_[41972]_  = ~A168 & ~A169;
  assign \new_[41973]_  = ~A170 & \new_[41972]_ ;
  assign \new_[41976]_  = ~A166 & A167;
  assign \new_[41979]_  = A233 & ~A232;
  assign \new_[41980]_  = \new_[41979]_  & \new_[41976]_ ;
  assign \new_[41981]_  = \new_[41980]_  & \new_[41973]_ ;
  assign \new_[41984]_  = A235 & A234;
  assign \new_[41987]_  = A266 & A265;
  assign \new_[41988]_  = \new_[41987]_  & \new_[41984]_ ;
  assign \new_[41991]_  = ~A299 & A298;
  assign \new_[41994]_  = ~A302 & A300;
  assign \new_[41995]_  = \new_[41994]_  & \new_[41991]_ ;
  assign \new_[41996]_  = \new_[41995]_  & \new_[41988]_ ;
  assign \new_[42000]_  = ~A168 & ~A169;
  assign \new_[42001]_  = ~A170 & \new_[42000]_ ;
  assign \new_[42004]_  = ~A166 & A167;
  assign \new_[42007]_  = A233 & ~A232;
  assign \new_[42008]_  = \new_[42007]_  & \new_[42004]_ ;
  assign \new_[42009]_  = \new_[42008]_  & \new_[42001]_ ;
  assign \new_[42012]_  = A235 & A234;
  assign \new_[42015]_  = A266 & A265;
  assign \new_[42016]_  = \new_[42015]_  & \new_[42012]_ ;
  assign \new_[42019]_  = A299 & ~A298;
  assign \new_[42022]_  = A301 & A300;
  assign \new_[42023]_  = \new_[42022]_  & \new_[42019]_ ;
  assign \new_[42024]_  = \new_[42023]_  & \new_[42016]_ ;
  assign \new_[42028]_  = ~A168 & ~A169;
  assign \new_[42029]_  = ~A170 & \new_[42028]_ ;
  assign \new_[42032]_  = ~A166 & A167;
  assign \new_[42035]_  = A233 & ~A232;
  assign \new_[42036]_  = \new_[42035]_  & \new_[42032]_ ;
  assign \new_[42037]_  = \new_[42036]_  & \new_[42029]_ ;
  assign \new_[42040]_  = A235 & A234;
  assign \new_[42043]_  = A266 & A265;
  assign \new_[42044]_  = \new_[42043]_  & \new_[42040]_ ;
  assign \new_[42047]_  = A299 & ~A298;
  assign \new_[42050]_  = ~A302 & A300;
  assign \new_[42051]_  = \new_[42050]_  & \new_[42047]_ ;
  assign \new_[42052]_  = \new_[42051]_  & \new_[42044]_ ;
  assign \new_[42056]_  = ~A168 & ~A169;
  assign \new_[42057]_  = ~A170 & \new_[42056]_ ;
  assign \new_[42060]_  = ~A166 & A167;
  assign \new_[42063]_  = A233 & ~A232;
  assign \new_[42064]_  = \new_[42063]_  & \new_[42060]_ ;
  assign \new_[42065]_  = \new_[42064]_  & \new_[42057]_ ;
  assign \new_[42068]_  = A235 & A234;
  assign \new_[42071]_  = ~A266 & ~A265;
  assign \new_[42072]_  = \new_[42071]_  & \new_[42068]_ ;
  assign \new_[42075]_  = ~A299 & A298;
  assign \new_[42078]_  = A301 & A300;
  assign \new_[42079]_  = \new_[42078]_  & \new_[42075]_ ;
  assign \new_[42080]_  = \new_[42079]_  & \new_[42072]_ ;
  assign \new_[42084]_  = ~A168 & ~A169;
  assign \new_[42085]_  = ~A170 & \new_[42084]_ ;
  assign \new_[42088]_  = ~A166 & A167;
  assign \new_[42091]_  = A233 & ~A232;
  assign \new_[42092]_  = \new_[42091]_  & \new_[42088]_ ;
  assign \new_[42093]_  = \new_[42092]_  & \new_[42085]_ ;
  assign \new_[42096]_  = A235 & A234;
  assign \new_[42099]_  = ~A266 & ~A265;
  assign \new_[42100]_  = \new_[42099]_  & \new_[42096]_ ;
  assign \new_[42103]_  = ~A299 & A298;
  assign \new_[42106]_  = ~A302 & A300;
  assign \new_[42107]_  = \new_[42106]_  & \new_[42103]_ ;
  assign \new_[42108]_  = \new_[42107]_  & \new_[42100]_ ;
  assign \new_[42112]_  = ~A168 & ~A169;
  assign \new_[42113]_  = ~A170 & \new_[42112]_ ;
  assign \new_[42116]_  = ~A166 & A167;
  assign \new_[42119]_  = A233 & ~A232;
  assign \new_[42120]_  = \new_[42119]_  & \new_[42116]_ ;
  assign \new_[42121]_  = \new_[42120]_  & \new_[42113]_ ;
  assign \new_[42124]_  = A235 & A234;
  assign \new_[42127]_  = ~A266 & ~A265;
  assign \new_[42128]_  = \new_[42127]_  & \new_[42124]_ ;
  assign \new_[42131]_  = A299 & ~A298;
  assign \new_[42134]_  = A301 & A300;
  assign \new_[42135]_  = \new_[42134]_  & \new_[42131]_ ;
  assign \new_[42136]_  = \new_[42135]_  & \new_[42128]_ ;
  assign \new_[42140]_  = ~A168 & ~A169;
  assign \new_[42141]_  = ~A170 & \new_[42140]_ ;
  assign \new_[42144]_  = ~A166 & A167;
  assign \new_[42147]_  = A233 & ~A232;
  assign \new_[42148]_  = \new_[42147]_  & \new_[42144]_ ;
  assign \new_[42149]_  = \new_[42148]_  & \new_[42141]_ ;
  assign \new_[42152]_  = A235 & A234;
  assign \new_[42155]_  = ~A266 & ~A265;
  assign \new_[42156]_  = \new_[42155]_  & \new_[42152]_ ;
  assign \new_[42159]_  = A299 & ~A298;
  assign \new_[42162]_  = ~A302 & A300;
  assign \new_[42163]_  = \new_[42162]_  & \new_[42159]_ ;
  assign \new_[42164]_  = \new_[42163]_  & \new_[42156]_ ;
  assign \new_[42168]_  = ~A168 & ~A169;
  assign \new_[42169]_  = ~A170 & \new_[42168]_ ;
  assign \new_[42172]_  = ~A166 & A167;
  assign \new_[42175]_  = A233 & ~A232;
  assign \new_[42176]_  = \new_[42175]_  & \new_[42172]_ ;
  assign \new_[42177]_  = \new_[42176]_  & \new_[42169]_ ;
  assign \new_[42180]_  = ~A236 & A234;
  assign \new_[42183]_  = A268 & ~A267;
  assign \new_[42184]_  = \new_[42183]_  & \new_[42180]_ ;
  assign \new_[42187]_  = ~A299 & A298;
  assign \new_[42190]_  = A301 & A300;
  assign \new_[42191]_  = \new_[42190]_  & \new_[42187]_ ;
  assign \new_[42192]_  = \new_[42191]_  & \new_[42184]_ ;
  assign \new_[42196]_  = ~A168 & ~A169;
  assign \new_[42197]_  = ~A170 & \new_[42196]_ ;
  assign \new_[42200]_  = ~A166 & A167;
  assign \new_[42203]_  = A233 & ~A232;
  assign \new_[42204]_  = \new_[42203]_  & \new_[42200]_ ;
  assign \new_[42205]_  = \new_[42204]_  & \new_[42197]_ ;
  assign \new_[42208]_  = ~A236 & A234;
  assign \new_[42211]_  = A268 & ~A267;
  assign \new_[42212]_  = \new_[42211]_  & \new_[42208]_ ;
  assign \new_[42215]_  = ~A299 & A298;
  assign \new_[42218]_  = ~A302 & A300;
  assign \new_[42219]_  = \new_[42218]_  & \new_[42215]_ ;
  assign \new_[42220]_  = \new_[42219]_  & \new_[42212]_ ;
  assign \new_[42224]_  = ~A168 & ~A169;
  assign \new_[42225]_  = ~A170 & \new_[42224]_ ;
  assign \new_[42228]_  = ~A166 & A167;
  assign \new_[42231]_  = A233 & ~A232;
  assign \new_[42232]_  = \new_[42231]_  & \new_[42228]_ ;
  assign \new_[42233]_  = \new_[42232]_  & \new_[42225]_ ;
  assign \new_[42236]_  = ~A236 & A234;
  assign \new_[42239]_  = A268 & ~A267;
  assign \new_[42240]_  = \new_[42239]_  & \new_[42236]_ ;
  assign \new_[42243]_  = A299 & ~A298;
  assign \new_[42246]_  = A301 & A300;
  assign \new_[42247]_  = \new_[42246]_  & \new_[42243]_ ;
  assign \new_[42248]_  = \new_[42247]_  & \new_[42240]_ ;
  assign \new_[42252]_  = ~A168 & ~A169;
  assign \new_[42253]_  = ~A170 & \new_[42252]_ ;
  assign \new_[42256]_  = ~A166 & A167;
  assign \new_[42259]_  = A233 & ~A232;
  assign \new_[42260]_  = \new_[42259]_  & \new_[42256]_ ;
  assign \new_[42261]_  = \new_[42260]_  & \new_[42253]_ ;
  assign \new_[42264]_  = ~A236 & A234;
  assign \new_[42267]_  = A268 & ~A267;
  assign \new_[42268]_  = \new_[42267]_  & \new_[42264]_ ;
  assign \new_[42271]_  = A299 & ~A298;
  assign \new_[42274]_  = ~A302 & A300;
  assign \new_[42275]_  = \new_[42274]_  & \new_[42271]_ ;
  assign \new_[42276]_  = \new_[42275]_  & \new_[42268]_ ;
  assign \new_[42280]_  = ~A168 & ~A169;
  assign \new_[42281]_  = ~A170 & \new_[42280]_ ;
  assign \new_[42284]_  = ~A166 & A167;
  assign \new_[42287]_  = A233 & ~A232;
  assign \new_[42288]_  = \new_[42287]_  & \new_[42284]_ ;
  assign \new_[42289]_  = \new_[42288]_  & \new_[42281]_ ;
  assign \new_[42292]_  = ~A236 & A234;
  assign \new_[42295]_  = ~A269 & ~A267;
  assign \new_[42296]_  = \new_[42295]_  & \new_[42292]_ ;
  assign \new_[42299]_  = ~A299 & A298;
  assign \new_[42302]_  = A301 & A300;
  assign \new_[42303]_  = \new_[42302]_  & \new_[42299]_ ;
  assign \new_[42304]_  = \new_[42303]_  & \new_[42296]_ ;
  assign \new_[42308]_  = ~A168 & ~A169;
  assign \new_[42309]_  = ~A170 & \new_[42308]_ ;
  assign \new_[42312]_  = ~A166 & A167;
  assign \new_[42315]_  = A233 & ~A232;
  assign \new_[42316]_  = \new_[42315]_  & \new_[42312]_ ;
  assign \new_[42317]_  = \new_[42316]_  & \new_[42309]_ ;
  assign \new_[42320]_  = ~A236 & A234;
  assign \new_[42323]_  = ~A269 & ~A267;
  assign \new_[42324]_  = \new_[42323]_  & \new_[42320]_ ;
  assign \new_[42327]_  = ~A299 & A298;
  assign \new_[42330]_  = ~A302 & A300;
  assign \new_[42331]_  = \new_[42330]_  & \new_[42327]_ ;
  assign \new_[42332]_  = \new_[42331]_  & \new_[42324]_ ;
  assign \new_[42336]_  = ~A168 & ~A169;
  assign \new_[42337]_  = ~A170 & \new_[42336]_ ;
  assign \new_[42340]_  = ~A166 & A167;
  assign \new_[42343]_  = A233 & ~A232;
  assign \new_[42344]_  = \new_[42343]_  & \new_[42340]_ ;
  assign \new_[42345]_  = \new_[42344]_  & \new_[42337]_ ;
  assign \new_[42348]_  = ~A236 & A234;
  assign \new_[42351]_  = ~A269 & ~A267;
  assign \new_[42352]_  = \new_[42351]_  & \new_[42348]_ ;
  assign \new_[42355]_  = A299 & ~A298;
  assign \new_[42358]_  = A301 & A300;
  assign \new_[42359]_  = \new_[42358]_  & \new_[42355]_ ;
  assign \new_[42360]_  = \new_[42359]_  & \new_[42352]_ ;
  assign \new_[42364]_  = ~A168 & ~A169;
  assign \new_[42365]_  = ~A170 & \new_[42364]_ ;
  assign \new_[42368]_  = ~A166 & A167;
  assign \new_[42371]_  = A233 & ~A232;
  assign \new_[42372]_  = \new_[42371]_  & \new_[42368]_ ;
  assign \new_[42373]_  = \new_[42372]_  & \new_[42365]_ ;
  assign \new_[42376]_  = ~A236 & A234;
  assign \new_[42379]_  = ~A269 & ~A267;
  assign \new_[42380]_  = \new_[42379]_  & \new_[42376]_ ;
  assign \new_[42383]_  = A299 & ~A298;
  assign \new_[42386]_  = ~A302 & A300;
  assign \new_[42387]_  = \new_[42386]_  & \new_[42383]_ ;
  assign \new_[42388]_  = \new_[42387]_  & \new_[42380]_ ;
  assign \new_[42392]_  = ~A168 & ~A169;
  assign \new_[42393]_  = ~A170 & \new_[42392]_ ;
  assign \new_[42396]_  = ~A166 & A167;
  assign \new_[42399]_  = A233 & ~A232;
  assign \new_[42400]_  = \new_[42399]_  & \new_[42396]_ ;
  assign \new_[42401]_  = \new_[42400]_  & \new_[42393]_ ;
  assign \new_[42404]_  = ~A236 & A234;
  assign \new_[42407]_  = A266 & A265;
  assign \new_[42408]_  = \new_[42407]_  & \new_[42404]_ ;
  assign \new_[42411]_  = ~A299 & A298;
  assign \new_[42414]_  = A301 & A300;
  assign \new_[42415]_  = \new_[42414]_  & \new_[42411]_ ;
  assign \new_[42416]_  = \new_[42415]_  & \new_[42408]_ ;
  assign \new_[42420]_  = ~A168 & ~A169;
  assign \new_[42421]_  = ~A170 & \new_[42420]_ ;
  assign \new_[42424]_  = ~A166 & A167;
  assign \new_[42427]_  = A233 & ~A232;
  assign \new_[42428]_  = \new_[42427]_  & \new_[42424]_ ;
  assign \new_[42429]_  = \new_[42428]_  & \new_[42421]_ ;
  assign \new_[42432]_  = ~A236 & A234;
  assign \new_[42435]_  = A266 & A265;
  assign \new_[42436]_  = \new_[42435]_  & \new_[42432]_ ;
  assign \new_[42439]_  = ~A299 & A298;
  assign \new_[42442]_  = ~A302 & A300;
  assign \new_[42443]_  = \new_[42442]_  & \new_[42439]_ ;
  assign \new_[42444]_  = \new_[42443]_  & \new_[42436]_ ;
  assign \new_[42448]_  = ~A168 & ~A169;
  assign \new_[42449]_  = ~A170 & \new_[42448]_ ;
  assign \new_[42452]_  = ~A166 & A167;
  assign \new_[42455]_  = A233 & ~A232;
  assign \new_[42456]_  = \new_[42455]_  & \new_[42452]_ ;
  assign \new_[42457]_  = \new_[42456]_  & \new_[42449]_ ;
  assign \new_[42460]_  = ~A236 & A234;
  assign \new_[42463]_  = A266 & A265;
  assign \new_[42464]_  = \new_[42463]_  & \new_[42460]_ ;
  assign \new_[42467]_  = A299 & ~A298;
  assign \new_[42470]_  = A301 & A300;
  assign \new_[42471]_  = \new_[42470]_  & \new_[42467]_ ;
  assign \new_[42472]_  = \new_[42471]_  & \new_[42464]_ ;
  assign \new_[42476]_  = ~A168 & ~A169;
  assign \new_[42477]_  = ~A170 & \new_[42476]_ ;
  assign \new_[42480]_  = ~A166 & A167;
  assign \new_[42483]_  = A233 & ~A232;
  assign \new_[42484]_  = \new_[42483]_  & \new_[42480]_ ;
  assign \new_[42485]_  = \new_[42484]_  & \new_[42477]_ ;
  assign \new_[42488]_  = ~A236 & A234;
  assign \new_[42491]_  = A266 & A265;
  assign \new_[42492]_  = \new_[42491]_  & \new_[42488]_ ;
  assign \new_[42495]_  = A299 & ~A298;
  assign \new_[42498]_  = ~A302 & A300;
  assign \new_[42499]_  = \new_[42498]_  & \new_[42495]_ ;
  assign \new_[42500]_  = \new_[42499]_  & \new_[42492]_ ;
  assign \new_[42504]_  = ~A168 & ~A169;
  assign \new_[42505]_  = ~A170 & \new_[42504]_ ;
  assign \new_[42508]_  = ~A166 & A167;
  assign \new_[42511]_  = A233 & ~A232;
  assign \new_[42512]_  = \new_[42511]_  & \new_[42508]_ ;
  assign \new_[42513]_  = \new_[42512]_  & \new_[42505]_ ;
  assign \new_[42516]_  = ~A236 & A234;
  assign \new_[42519]_  = ~A266 & ~A265;
  assign \new_[42520]_  = \new_[42519]_  & \new_[42516]_ ;
  assign \new_[42523]_  = ~A299 & A298;
  assign \new_[42526]_  = A301 & A300;
  assign \new_[42527]_  = \new_[42526]_  & \new_[42523]_ ;
  assign \new_[42528]_  = \new_[42527]_  & \new_[42520]_ ;
  assign \new_[42532]_  = ~A168 & ~A169;
  assign \new_[42533]_  = ~A170 & \new_[42532]_ ;
  assign \new_[42536]_  = ~A166 & A167;
  assign \new_[42539]_  = A233 & ~A232;
  assign \new_[42540]_  = \new_[42539]_  & \new_[42536]_ ;
  assign \new_[42541]_  = \new_[42540]_  & \new_[42533]_ ;
  assign \new_[42544]_  = ~A236 & A234;
  assign \new_[42547]_  = ~A266 & ~A265;
  assign \new_[42548]_  = \new_[42547]_  & \new_[42544]_ ;
  assign \new_[42551]_  = ~A299 & A298;
  assign \new_[42554]_  = ~A302 & A300;
  assign \new_[42555]_  = \new_[42554]_  & \new_[42551]_ ;
  assign \new_[42556]_  = \new_[42555]_  & \new_[42548]_ ;
  assign \new_[42560]_  = ~A168 & ~A169;
  assign \new_[42561]_  = ~A170 & \new_[42560]_ ;
  assign \new_[42564]_  = ~A166 & A167;
  assign \new_[42567]_  = A233 & ~A232;
  assign \new_[42568]_  = \new_[42567]_  & \new_[42564]_ ;
  assign \new_[42569]_  = \new_[42568]_  & \new_[42561]_ ;
  assign \new_[42572]_  = ~A236 & A234;
  assign \new_[42575]_  = ~A266 & ~A265;
  assign \new_[42576]_  = \new_[42575]_  & \new_[42572]_ ;
  assign \new_[42579]_  = A299 & ~A298;
  assign \new_[42582]_  = A301 & A300;
  assign \new_[42583]_  = \new_[42582]_  & \new_[42579]_ ;
  assign \new_[42584]_  = \new_[42583]_  & \new_[42576]_ ;
  assign \new_[42588]_  = ~A168 & ~A169;
  assign \new_[42589]_  = ~A170 & \new_[42588]_ ;
  assign \new_[42592]_  = ~A166 & A167;
  assign \new_[42595]_  = A233 & ~A232;
  assign \new_[42596]_  = \new_[42595]_  & \new_[42592]_ ;
  assign \new_[42597]_  = \new_[42596]_  & \new_[42589]_ ;
  assign \new_[42600]_  = ~A236 & A234;
  assign \new_[42603]_  = ~A266 & ~A265;
  assign \new_[42604]_  = \new_[42603]_  & \new_[42600]_ ;
  assign \new_[42607]_  = A299 & ~A298;
  assign \new_[42610]_  = ~A302 & A300;
  assign \new_[42611]_  = \new_[42610]_  & \new_[42607]_ ;
  assign \new_[42612]_  = \new_[42611]_  & \new_[42604]_ ;
  assign \new_[42616]_  = ~A168 & ~A169;
  assign \new_[42617]_  = ~A170 & \new_[42616]_ ;
  assign \new_[42620]_  = ~A166 & A167;
  assign \new_[42623]_  = ~A233 & A232;
  assign \new_[42624]_  = \new_[42623]_  & \new_[42620]_ ;
  assign \new_[42625]_  = \new_[42624]_  & \new_[42617]_ ;
  assign \new_[42628]_  = A235 & A234;
  assign \new_[42631]_  = A268 & ~A267;
  assign \new_[42632]_  = \new_[42631]_  & \new_[42628]_ ;
  assign \new_[42635]_  = ~A299 & A298;
  assign \new_[42638]_  = A301 & A300;
  assign \new_[42639]_  = \new_[42638]_  & \new_[42635]_ ;
  assign \new_[42640]_  = \new_[42639]_  & \new_[42632]_ ;
  assign \new_[42644]_  = ~A168 & ~A169;
  assign \new_[42645]_  = ~A170 & \new_[42644]_ ;
  assign \new_[42648]_  = ~A166 & A167;
  assign \new_[42651]_  = ~A233 & A232;
  assign \new_[42652]_  = \new_[42651]_  & \new_[42648]_ ;
  assign \new_[42653]_  = \new_[42652]_  & \new_[42645]_ ;
  assign \new_[42656]_  = A235 & A234;
  assign \new_[42659]_  = A268 & ~A267;
  assign \new_[42660]_  = \new_[42659]_  & \new_[42656]_ ;
  assign \new_[42663]_  = ~A299 & A298;
  assign \new_[42666]_  = ~A302 & A300;
  assign \new_[42667]_  = \new_[42666]_  & \new_[42663]_ ;
  assign \new_[42668]_  = \new_[42667]_  & \new_[42660]_ ;
  assign \new_[42672]_  = ~A168 & ~A169;
  assign \new_[42673]_  = ~A170 & \new_[42672]_ ;
  assign \new_[42676]_  = ~A166 & A167;
  assign \new_[42679]_  = ~A233 & A232;
  assign \new_[42680]_  = \new_[42679]_  & \new_[42676]_ ;
  assign \new_[42681]_  = \new_[42680]_  & \new_[42673]_ ;
  assign \new_[42684]_  = A235 & A234;
  assign \new_[42687]_  = A268 & ~A267;
  assign \new_[42688]_  = \new_[42687]_  & \new_[42684]_ ;
  assign \new_[42691]_  = A299 & ~A298;
  assign \new_[42694]_  = A301 & A300;
  assign \new_[42695]_  = \new_[42694]_  & \new_[42691]_ ;
  assign \new_[42696]_  = \new_[42695]_  & \new_[42688]_ ;
  assign \new_[42700]_  = ~A168 & ~A169;
  assign \new_[42701]_  = ~A170 & \new_[42700]_ ;
  assign \new_[42704]_  = ~A166 & A167;
  assign \new_[42707]_  = ~A233 & A232;
  assign \new_[42708]_  = \new_[42707]_  & \new_[42704]_ ;
  assign \new_[42709]_  = \new_[42708]_  & \new_[42701]_ ;
  assign \new_[42712]_  = A235 & A234;
  assign \new_[42715]_  = A268 & ~A267;
  assign \new_[42716]_  = \new_[42715]_  & \new_[42712]_ ;
  assign \new_[42719]_  = A299 & ~A298;
  assign \new_[42722]_  = ~A302 & A300;
  assign \new_[42723]_  = \new_[42722]_  & \new_[42719]_ ;
  assign \new_[42724]_  = \new_[42723]_  & \new_[42716]_ ;
  assign \new_[42728]_  = ~A168 & ~A169;
  assign \new_[42729]_  = ~A170 & \new_[42728]_ ;
  assign \new_[42732]_  = ~A166 & A167;
  assign \new_[42735]_  = ~A233 & A232;
  assign \new_[42736]_  = \new_[42735]_  & \new_[42732]_ ;
  assign \new_[42737]_  = \new_[42736]_  & \new_[42729]_ ;
  assign \new_[42740]_  = A235 & A234;
  assign \new_[42743]_  = ~A269 & ~A267;
  assign \new_[42744]_  = \new_[42743]_  & \new_[42740]_ ;
  assign \new_[42747]_  = ~A299 & A298;
  assign \new_[42750]_  = A301 & A300;
  assign \new_[42751]_  = \new_[42750]_  & \new_[42747]_ ;
  assign \new_[42752]_  = \new_[42751]_  & \new_[42744]_ ;
  assign \new_[42756]_  = ~A168 & ~A169;
  assign \new_[42757]_  = ~A170 & \new_[42756]_ ;
  assign \new_[42760]_  = ~A166 & A167;
  assign \new_[42763]_  = ~A233 & A232;
  assign \new_[42764]_  = \new_[42763]_  & \new_[42760]_ ;
  assign \new_[42765]_  = \new_[42764]_  & \new_[42757]_ ;
  assign \new_[42768]_  = A235 & A234;
  assign \new_[42771]_  = ~A269 & ~A267;
  assign \new_[42772]_  = \new_[42771]_  & \new_[42768]_ ;
  assign \new_[42775]_  = ~A299 & A298;
  assign \new_[42778]_  = ~A302 & A300;
  assign \new_[42779]_  = \new_[42778]_  & \new_[42775]_ ;
  assign \new_[42780]_  = \new_[42779]_  & \new_[42772]_ ;
  assign \new_[42784]_  = ~A168 & ~A169;
  assign \new_[42785]_  = ~A170 & \new_[42784]_ ;
  assign \new_[42788]_  = ~A166 & A167;
  assign \new_[42791]_  = ~A233 & A232;
  assign \new_[42792]_  = \new_[42791]_  & \new_[42788]_ ;
  assign \new_[42793]_  = \new_[42792]_  & \new_[42785]_ ;
  assign \new_[42796]_  = A235 & A234;
  assign \new_[42799]_  = ~A269 & ~A267;
  assign \new_[42800]_  = \new_[42799]_  & \new_[42796]_ ;
  assign \new_[42803]_  = A299 & ~A298;
  assign \new_[42806]_  = A301 & A300;
  assign \new_[42807]_  = \new_[42806]_  & \new_[42803]_ ;
  assign \new_[42808]_  = \new_[42807]_  & \new_[42800]_ ;
  assign \new_[42812]_  = ~A168 & ~A169;
  assign \new_[42813]_  = ~A170 & \new_[42812]_ ;
  assign \new_[42816]_  = ~A166 & A167;
  assign \new_[42819]_  = ~A233 & A232;
  assign \new_[42820]_  = \new_[42819]_  & \new_[42816]_ ;
  assign \new_[42821]_  = \new_[42820]_  & \new_[42813]_ ;
  assign \new_[42824]_  = A235 & A234;
  assign \new_[42827]_  = ~A269 & ~A267;
  assign \new_[42828]_  = \new_[42827]_  & \new_[42824]_ ;
  assign \new_[42831]_  = A299 & ~A298;
  assign \new_[42834]_  = ~A302 & A300;
  assign \new_[42835]_  = \new_[42834]_  & \new_[42831]_ ;
  assign \new_[42836]_  = \new_[42835]_  & \new_[42828]_ ;
  assign \new_[42840]_  = ~A168 & ~A169;
  assign \new_[42841]_  = ~A170 & \new_[42840]_ ;
  assign \new_[42844]_  = ~A166 & A167;
  assign \new_[42847]_  = ~A233 & A232;
  assign \new_[42848]_  = \new_[42847]_  & \new_[42844]_ ;
  assign \new_[42849]_  = \new_[42848]_  & \new_[42841]_ ;
  assign \new_[42852]_  = A235 & A234;
  assign \new_[42855]_  = A266 & A265;
  assign \new_[42856]_  = \new_[42855]_  & \new_[42852]_ ;
  assign \new_[42859]_  = ~A299 & A298;
  assign \new_[42862]_  = A301 & A300;
  assign \new_[42863]_  = \new_[42862]_  & \new_[42859]_ ;
  assign \new_[42864]_  = \new_[42863]_  & \new_[42856]_ ;
  assign \new_[42868]_  = ~A168 & ~A169;
  assign \new_[42869]_  = ~A170 & \new_[42868]_ ;
  assign \new_[42872]_  = ~A166 & A167;
  assign \new_[42875]_  = ~A233 & A232;
  assign \new_[42876]_  = \new_[42875]_  & \new_[42872]_ ;
  assign \new_[42877]_  = \new_[42876]_  & \new_[42869]_ ;
  assign \new_[42880]_  = A235 & A234;
  assign \new_[42883]_  = A266 & A265;
  assign \new_[42884]_  = \new_[42883]_  & \new_[42880]_ ;
  assign \new_[42887]_  = ~A299 & A298;
  assign \new_[42890]_  = ~A302 & A300;
  assign \new_[42891]_  = \new_[42890]_  & \new_[42887]_ ;
  assign \new_[42892]_  = \new_[42891]_  & \new_[42884]_ ;
  assign \new_[42896]_  = ~A168 & ~A169;
  assign \new_[42897]_  = ~A170 & \new_[42896]_ ;
  assign \new_[42900]_  = ~A166 & A167;
  assign \new_[42903]_  = ~A233 & A232;
  assign \new_[42904]_  = \new_[42903]_  & \new_[42900]_ ;
  assign \new_[42905]_  = \new_[42904]_  & \new_[42897]_ ;
  assign \new_[42908]_  = A235 & A234;
  assign \new_[42911]_  = A266 & A265;
  assign \new_[42912]_  = \new_[42911]_  & \new_[42908]_ ;
  assign \new_[42915]_  = A299 & ~A298;
  assign \new_[42918]_  = A301 & A300;
  assign \new_[42919]_  = \new_[42918]_  & \new_[42915]_ ;
  assign \new_[42920]_  = \new_[42919]_  & \new_[42912]_ ;
  assign \new_[42924]_  = ~A168 & ~A169;
  assign \new_[42925]_  = ~A170 & \new_[42924]_ ;
  assign \new_[42928]_  = ~A166 & A167;
  assign \new_[42931]_  = ~A233 & A232;
  assign \new_[42932]_  = \new_[42931]_  & \new_[42928]_ ;
  assign \new_[42933]_  = \new_[42932]_  & \new_[42925]_ ;
  assign \new_[42936]_  = A235 & A234;
  assign \new_[42939]_  = A266 & A265;
  assign \new_[42940]_  = \new_[42939]_  & \new_[42936]_ ;
  assign \new_[42943]_  = A299 & ~A298;
  assign \new_[42946]_  = ~A302 & A300;
  assign \new_[42947]_  = \new_[42946]_  & \new_[42943]_ ;
  assign \new_[42948]_  = \new_[42947]_  & \new_[42940]_ ;
  assign \new_[42952]_  = ~A168 & ~A169;
  assign \new_[42953]_  = ~A170 & \new_[42952]_ ;
  assign \new_[42956]_  = ~A166 & A167;
  assign \new_[42959]_  = ~A233 & A232;
  assign \new_[42960]_  = \new_[42959]_  & \new_[42956]_ ;
  assign \new_[42961]_  = \new_[42960]_  & \new_[42953]_ ;
  assign \new_[42964]_  = A235 & A234;
  assign \new_[42967]_  = ~A266 & ~A265;
  assign \new_[42968]_  = \new_[42967]_  & \new_[42964]_ ;
  assign \new_[42971]_  = ~A299 & A298;
  assign \new_[42974]_  = A301 & A300;
  assign \new_[42975]_  = \new_[42974]_  & \new_[42971]_ ;
  assign \new_[42976]_  = \new_[42975]_  & \new_[42968]_ ;
  assign \new_[42980]_  = ~A168 & ~A169;
  assign \new_[42981]_  = ~A170 & \new_[42980]_ ;
  assign \new_[42984]_  = ~A166 & A167;
  assign \new_[42987]_  = ~A233 & A232;
  assign \new_[42988]_  = \new_[42987]_  & \new_[42984]_ ;
  assign \new_[42989]_  = \new_[42988]_  & \new_[42981]_ ;
  assign \new_[42992]_  = A235 & A234;
  assign \new_[42995]_  = ~A266 & ~A265;
  assign \new_[42996]_  = \new_[42995]_  & \new_[42992]_ ;
  assign \new_[42999]_  = ~A299 & A298;
  assign \new_[43002]_  = ~A302 & A300;
  assign \new_[43003]_  = \new_[43002]_  & \new_[42999]_ ;
  assign \new_[43004]_  = \new_[43003]_  & \new_[42996]_ ;
  assign \new_[43008]_  = ~A168 & ~A169;
  assign \new_[43009]_  = ~A170 & \new_[43008]_ ;
  assign \new_[43012]_  = ~A166 & A167;
  assign \new_[43015]_  = ~A233 & A232;
  assign \new_[43016]_  = \new_[43015]_  & \new_[43012]_ ;
  assign \new_[43017]_  = \new_[43016]_  & \new_[43009]_ ;
  assign \new_[43020]_  = A235 & A234;
  assign \new_[43023]_  = ~A266 & ~A265;
  assign \new_[43024]_  = \new_[43023]_  & \new_[43020]_ ;
  assign \new_[43027]_  = A299 & ~A298;
  assign \new_[43030]_  = A301 & A300;
  assign \new_[43031]_  = \new_[43030]_  & \new_[43027]_ ;
  assign \new_[43032]_  = \new_[43031]_  & \new_[43024]_ ;
  assign \new_[43036]_  = ~A168 & ~A169;
  assign \new_[43037]_  = ~A170 & \new_[43036]_ ;
  assign \new_[43040]_  = ~A166 & A167;
  assign \new_[43043]_  = ~A233 & A232;
  assign \new_[43044]_  = \new_[43043]_  & \new_[43040]_ ;
  assign \new_[43045]_  = \new_[43044]_  & \new_[43037]_ ;
  assign \new_[43048]_  = A235 & A234;
  assign \new_[43051]_  = ~A266 & ~A265;
  assign \new_[43052]_  = \new_[43051]_  & \new_[43048]_ ;
  assign \new_[43055]_  = A299 & ~A298;
  assign \new_[43058]_  = ~A302 & A300;
  assign \new_[43059]_  = \new_[43058]_  & \new_[43055]_ ;
  assign \new_[43060]_  = \new_[43059]_  & \new_[43052]_ ;
  assign \new_[43064]_  = ~A168 & ~A169;
  assign \new_[43065]_  = ~A170 & \new_[43064]_ ;
  assign \new_[43068]_  = ~A166 & A167;
  assign \new_[43071]_  = ~A233 & A232;
  assign \new_[43072]_  = \new_[43071]_  & \new_[43068]_ ;
  assign \new_[43073]_  = \new_[43072]_  & \new_[43065]_ ;
  assign \new_[43076]_  = ~A236 & A234;
  assign \new_[43079]_  = A268 & ~A267;
  assign \new_[43080]_  = \new_[43079]_  & \new_[43076]_ ;
  assign \new_[43083]_  = ~A299 & A298;
  assign \new_[43086]_  = A301 & A300;
  assign \new_[43087]_  = \new_[43086]_  & \new_[43083]_ ;
  assign \new_[43088]_  = \new_[43087]_  & \new_[43080]_ ;
  assign \new_[43092]_  = ~A168 & ~A169;
  assign \new_[43093]_  = ~A170 & \new_[43092]_ ;
  assign \new_[43096]_  = ~A166 & A167;
  assign \new_[43099]_  = ~A233 & A232;
  assign \new_[43100]_  = \new_[43099]_  & \new_[43096]_ ;
  assign \new_[43101]_  = \new_[43100]_  & \new_[43093]_ ;
  assign \new_[43104]_  = ~A236 & A234;
  assign \new_[43107]_  = A268 & ~A267;
  assign \new_[43108]_  = \new_[43107]_  & \new_[43104]_ ;
  assign \new_[43111]_  = ~A299 & A298;
  assign \new_[43114]_  = ~A302 & A300;
  assign \new_[43115]_  = \new_[43114]_  & \new_[43111]_ ;
  assign \new_[43116]_  = \new_[43115]_  & \new_[43108]_ ;
  assign \new_[43120]_  = ~A168 & ~A169;
  assign \new_[43121]_  = ~A170 & \new_[43120]_ ;
  assign \new_[43124]_  = ~A166 & A167;
  assign \new_[43127]_  = ~A233 & A232;
  assign \new_[43128]_  = \new_[43127]_  & \new_[43124]_ ;
  assign \new_[43129]_  = \new_[43128]_  & \new_[43121]_ ;
  assign \new_[43132]_  = ~A236 & A234;
  assign \new_[43135]_  = A268 & ~A267;
  assign \new_[43136]_  = \new_[43135]_  & \new_[43132]_ ;
  assign \new_[43139]_  = A299 & ~A298;
  assign \new_[43142]_  = A301 & A300;
  assign \new_[43143]_  = \new_[43142]_  & \new_[43139]_ ;
  assign \new_[43144]_  = \new_[43143]_  & \new_[43136]_ ;
  assign \new_[43148]_  = ~A168 & ~A169;
  assign \new_[43149]_  = ~A170 & \new_[43148]_ ;
  assign \new_[43152]_  = ~A166 & A167;
  assign \new_[43155]_  = ~A233 & A232;
  assign \new_[43156]_  = \new_[43155]_  & \new_[43152]_ ;
  assign \new_[43157]_  = \new_[43156]_  & \new_[43149]_ ;
  assign \new_[43160]_  = ~A236 & A234;
  assign \new_[43163]_  = A268 & ~A267;
  assign \new_[43164]_  = \new_[43163]_  & \new_[43160]_ ;
  assign \new_[43167]_  = A299 & ~A298;
  assign \new_[43170]_  = ~A302 & A300;
  assign \new_[43171]_  = \new_[43170]_  & \new_[43167]_ ;
  assign \new_[43172]_  = \new_[43171]_  & \new_[43164]_ ;
  assign \new_[43176]_  = ~A168 & ~A169;
  assign \new_[43177]_  = ~A170 & \new_[43176]_ ;
  assign \new_[43180]_  = ~A166 & A167;
  assign \new_[43183]_  = ~A233 & A232;
  assign \new_[43184]_  = \new_[43183]_  & \new_[43180]_ ;
  assign \new_[43185]_  = \new_[43184]_  & \new_[43177]_ ;
  assign \new_[43188]_  = ~A236 & A234;
  assign \new_[43191]_  = ~A269 & ~A267;
  assign \new_[43192]_  = \new_[43191]_  & \new_[43188]_ ;
  assign \new_[43195]_  = ~A299 & A298;
  assign \new_[43198]_  = A301 & A300;
  assign \new_[43199]_  = \new_[43198]_  & \new_[43195]_ ;
  assign \new_[43200]_  = \new_[43199]_  & \new_[43192]_ ;
  assign \new_[43204]_  = ~A168 & ~A169;
  assign \new_[43205]_  = ~A170 & \new_[43204]_ ;
  assign \new_[43208]_  = ~A166 & A167;
  assign \new_[43211]_  = ~A233 & A232;
  assign \new_[43212]_  = \new_[43211]_  & \new_[43208]_ ;
  assign \new_[43213]_  = \new_[43212]_  & \new_[43205]_ ;
  assign \new_[43216]_  = ~A236 & A234;
  assign \new_[43219]_  = ~A269 & ~A267;
  assign \new_[43220]_  = \new_[43219]_  & \new_[43216]_ ;
  assign \new_[43223]_  = ~A299 & A298;
  assign \new_[43226]_  = ~A302 & A300;
  assign \new_[43227]_  = \new_[43226]_  & \new_[43223]_ ;
  assign \new_[43228]_  = \new_[43227]_  & \new_[43220]_ ;
  assign \new_[43232]_  = ~A168 & ~A169;
  assign \new_[43233]_  = ~A170 & \new_[43232]_ ;
  assign \new_[43236]_  = ~A166 & A167;
  assign \new_[43239]_  = ~A233 & A232;
  assign \new_[43240]_  = \new_[43239]_  & \new_[43236]_ ;
  assign \new_[43241]_  = \new_[43240]_  & \new_[43233]_ ;
  assign \new_[43244]_  = ~A236 & A234;
  assign \new_[43247]_  = ~A269 & ~A267;
  assign \new_[43248]_  = \new_[43247]_  & \new_[43244]_ ;
  assign \new_[43251]_  = A299 & ~A298;
  assign \new_[43254]_  = A301 & A300;
  assign \new_[43255]_  = \new_[43254]_  & \new_[43251]_ ;
  assign \new_[43256]_  = \new_[43255]_  & \new_[43248]_ ;
  assign \new_[43260]_  = ~A168 & ~A169;
  assign \new_[43261]_  = ~A170 & \new_[43260]_ ;
  assign \new_[43264]_  = ~A166 & A167;
  assign \new_[43267]_  = ~A233 & A232;
  assign \new_[43268]_  = \new_[43267]_  & \new_[43264]_ ;
  assign \new_[43269]_  = \new_[43268]_  & \new_[43261]_ ;
  assign \new_[43272]_  = ~A236 & A234;
  assign \new_[43275]_  = ~A269 & ~A267;
  assign \new_[43276]_  = \new_[43275]_  & \new_[43272]_ ;
  assign \new_[43279]_  = A299 & ~A298;
  assign \new_[43282]_  = ~A302 & A300;
  assign \new_[43283]_  = \new_[43282]_  & \new_[43279]_ ;
  assign \new_[43284]_  = \new_[43283]_  & \new_[43276]_ ;
  assign \new_[43288]_  = ~A168 & ~A169;
  assign \new_[43289]_  = ~A170 & \new_[43288]_ ;
  assign \new_[43292]_  = ~A166 & A167;
  assign \new_[43295]_  = ~A233 & A232;
  assign \new_[43296]_  = \new_[43295]_  & \new_[43292]_ ;
  assign \new_[43297]_  = \new_[43296]_  & \new_[43289]_ ;
  assign \new_[43300]_  = ~A236 & A234;
  assign \new_[43303]_  = A266 & A265;
  assign \new_[43304]_  = \new_[43303]_  & \new_[43300]_ ;
  assign \new_[43307]_  = ~A299 & A298;
  assign \new_[43310]_  = A301 & A300;
  assign \new_[43311]_  = \new_[43310]_  & \new_[43307]_ ;
  assign \new_[43312]_  = \new_[43311]_  & \new_[43304]_ ;
  assign \new_[43316]_  = ~A168 & ~A169;
  assign \new_[43317]_  = ~A170 & \new_[43316]_ ;
  assign \new_[43320]_  = ~A166 & A167;
  assign \new_[43323]_  = ~A233 & A232;
  assign \new_[43324]_  = \new_[43323]_  & \new_[43320]_ ;
  assign \new_[43325]_  = \new_[43324]_  & \new_[43317]_ ;
  assign \new_[43328]_  = ~A236 & A234;
  assign \new_[43331]_  = A266 & A265;
  assign \new_[43332]_  = \new_[43331]_  & \new_[43328]_ ;
  assign \new_[43335]_  = ~A299 & A298;
  assign \new_[43338]_  = ~A302 & A300;
  assign \new_[43339]_  = \new_[43338]_  & \new_[43335]_ ;
  assign \new_[43340]_  = \new_[43339]_  & \new_[43332]_ ;
  assign \new_[43344]_  = ~A168 & ~A169;
  assign \new_[43345]_  = ~A170 & \new_[43344]_ ;
  assign \new_[43348]_  = ~A166 & A167;
  assign \new_[43351]_  = ~A233 & A232;
  assign \new_[43352]_  = \new_[43351]_  & \new_[43348]_ ;
  assign \new_[43353]_  = \new_[43352]_  & \new_[43345]_ ;
  assign \new_[43356]_  = ~A236 & A234;
  assign \new_[43359]_  = A266 & A265;
  assign \new_[43360]_  = \new_[43359]_  & \new_[43356]_ ;
  assign \new_[43363]_  = A299 & ~A298;
  assign \new_[43366]_  = A301 & A300;
  assign \new_[43367]_  = \new_[43366]_  & \new_[43363]_ ;
  assign \new_[43368]_  = \new_[43367]_  & \new_[43360]_ ;
  assign \new_[43372]_  = ~A168 & ~A169;
  assign \new_[43373]_  = ~A170 & \new_[43372]_ ;
  assign \new_[43376]_  = ~A166 & A167;
  assign \new_[43379]_  = ~A233 & A232;
  assign \new_[43380]_  = \new_[43379]_  & \new_[43376]_ ;
  assign \new_[43381]_  = \new_[43380]_  & \new_[43373]_ ;
  assign \new_[43384]_  = ~A236 & A234;
  assign \new_[43387]_  = A266 & A265;
  assign \new_[43388]_  = \new_[43387]_  & \new_[43384]_ ;
  assign \new_[43391]_  = A299 & ~A298;
  assign \new_[43394]_  = ~A302 & A300;
  assign \new_[43395]_  = \new_[43394]_  & \new_[43391]_ ;
  assign \new_[43396]_  = \new_[43395]_  & \new_[43388]_ ;
  assign \new_[43400]_  = ~A168 & ~A169;
  assign \new_[43401]_  = ~A170 & \new_[43400]_ ;
  assign \new_[43404]_  = ~A166 & A167;
  assign \new_[43407]_  = ~A233 & A232;
  assign \new_[43408]_  = \new_[43407]_  & \new_[43404]_ ;
  assign \new_[43409]_  = \new_[43408]_  & \new_[43401]_ ;
  assign \new_[43412]_  = ~A236 & A234;
  assign \new_[43415]_  = ~A266 & ~A265;
  assign \new_[43416]_  = \new_[43415]_  & \new_[43412]_ ;
  assign \new_[43419]_  = ~A299 & A298;
  assign \new_[43422]_  = A301 & A300;
  assign \new_[43423]_  = \new_[43422]_  & \new_[43419]_ ;
  assign \new_[43424]_  = \new_[43423]_  & \new_[43416]_ ;
  assign \new_[43428]_  = ~A168 & ~A169;
  assign \new_[43429]_  = ~A170 & \new_[43428]_ ;
  assign \new_[43432]_  = ~A166 & A167;
  assign \new_[43435]_  = ~A233 & A232;
  assign \new_[43436]_  = \new_[43435]_  & \new_[43432]_ ;
  assign \new_[43437]_  = \new_[43436]_  & \new_[43429]_ ;
  assign \new_[43440]_  = ~A236 & A234;
  assign \new_[43443]_  = ~A266 & ~A265;
  assign \new_[43444]_  = \new_[43443]_  & \new_[43440]_ ;
  assign \new_[43447]_  = ~A299 & A298;
  assign \new_[43450]_  = ~A302 & A300;
  assign \new_[43451]_  = \new_[43450]_  & \new_[43447]_ ;
  assign \new_[43452]_  = \new_[43451]_  & \new_[43444]_ ;
  assign \new_[43456]_  = ~A168 & ~A169;
  assign \new_[43457]_  = ~A170 & \new_[43456]_ ;
  assign \new_[43460]_  = ~A166 & A167;
  assign \new_[43463]_  = ~A233 & A232;
  assign \new_[43464]_  = \new_[43463]_  & \new_[43460]_ ;
  assign \new_[43465]_  = \new_[43464]_  & \new_[43457]_ ;
  assign \new_[43468]_  = ~A236 & A234;
  assign \new_[43471]_  = ~A266 & ~A265;
  assign \new_[43472]_  = \new_[43471]_  & \new_[43468]_ ;
  assign \new_[43475]_  = A299 & ~A298;
  assign \new_[43478]_  = A301 & A300;
  assign \new_[43479]_  = \new_[43478]_  & \new_[43475]_ ;
  assign \new_[43480]_  = \new_[43479]_  & \new_[43472]_ ;
  assign \new_[43484]_  = ~A168 & ~A169;
  assign \new_[43485]_  = ~A170 & \new_[43484]_ ;
  assign \new_[43488]_  = ~A166 & A167;
  assign \new_[43491]_  = ~A233 & A232;
  assign \new_[43492]_  = \new_[43491]_  & \new_[43488]_ ;
  assign \new_[43493]_  = \new_[43492]_  & \new_[43485]_ ;
  assign \new_[43496]_  = ~A236 & A234;
  assign \new_[43499]_  = ~A266 & ~A265;
  assign \new_[43500]_  = \new_[43499]_  & \new_[43496]_ ;
  assign \new_[43503]_  = A299 & ~A298;
  assign \new_[43506]_  = ~A302 & A300;
  assign \new_[43507]_  = \new_[43506]_  & \new_[43503]_ ;
  assign \new_[43508]_  = \new_[43507]_  & \new_[43500]_ ;
  assign \new_[43512]_  = ~A168 & ~A169;
  assign \new_[43513]_  = ~A170 & \new_[43512]_ ;
  assign \new_[43516]_  = A166 & ~A167;
  assign \new_[43519]_  = A233 & ~A232;
  assign \new_[43520]_  = \new_[43519]_  & \new_[43516]_ ;
  assign \new_[43521]_  = \new_[43520]_  & \new_[43513]_ ;
  assign \new_[43524]_  = A235 & A234;
  assign \new_[43527]_  = A268 & ~A267;
  assign \new_[43528]_  = \new_[43527]_  & \new_[43524]_ ;
  assign \new_[43531]_  = ~A299 & A298;
  assign \new_[43534]_  = A301 & A300;
  assign \new_[43535]_  = \new_[43534]_  & \new_[43531]_ ;
  assign \new_[43536]_  = \new_[43535]_  & \new_[43528]_ ;
  assign \new_[43540]_  = ~A168 & ~A169;
  assign \new_[43541]_  = ~A170 & \new_[43540]_ ;
  assign \new_[43544]_  = A166 & ~A167;
  assign \new_[43547]_  = A233 & ~A232;
  assign \new_[43548]_  = \new_[43547]_  & \new_[43544]_ ;
  assign \new_[43549]_  = \new_[43548]_  & \new_[43541]_ ;
  assign \new_[43552]_  = A235 & A234;
  assign \new_[43555]_  = A268 & ~A267;
  assign \new_[43556]_  = \new_[43555]_  & \new_[43552]_ ;
  assign \new_[43559]_  = ~A299 & A298;
  assign \new_[43562]_  = ~A302 & A300;
  assign \new_[43563]_  = \new_[43562]_  & \new_[43559]_ ;
  assign \new_[43564]_  = \new_[43563]_  & \new_[43556]_ ;
  assign \new_[43568]_  = ~A168 & ~A169;
  assign \new_[43569]_  = ~A170 & \new_[43568]_ ;
  assign \new_[43572]_  = A166 & ~A167;
  assign \new_[43575]_  = A233 & ~A232;
  assign \new_[43576]_  = \new_[43575]_  & \new_[43572]_ ;
  assign \new_[43577]_  = \new_[43576]_  & \new_[43569]_ ;
  assign \new_[43580]_  = A235 & A234;
  assign \new_[43583]_  = A268 & ~A267;
  assign \new_[43584]_  = \new_[43583]_  & \new_[43580]_ ;
  assign \new_[43587]_  = A299 & ~A298;
  assign \new_[43590]_  = A301 & A300;
  assign \new_[43591]_  = \new_[43590]_  & \new_[43587]_ ;
  assign \new_[43592]_  = \new_[43591]_  & \new_[43584]_ ;
  assign \new_[43596]_  = ~A168 & ~A169;
  assign \new_[43597]_  = ~A170 & \new_[43596]_ ;
  assign \new_[43600]_  = A166 & ~A167;
  assign \new_[43603]_  = A233 & ~A232;
  assign \new_[43604]_  = \new_[43603]_  & \new_[43600]_ ;
  assign \new_[43605]_  = \new_[43604]_  & \new_[43597]_ ;
  assign \new_[43608]_  = A235 & A234;
  assign \new_[43611]_  = A268 & ~A267;
  assign \new_[43612]_  = \new_[43611]_  & \new_[43608]_ ;
  assign \new_[43615]_  = A299 & ~A298;
  assign \new_[43618]_  = ~A302 & A300;
  assign \new_[43619]_  = \new_[43618]_  & \new_[43615]_ ;
  assign \new_[43620]_  = \new_[43619]_  & \new_[43612]_ ;
  assign \new_[43624]_  = ~A168 & ~A169;
  assign \new_[43625]_  = ~A170 & \new_[43624]_ ;
  assign \new_[43628]_  = A166 & ~A167;
  assign \new_[43631]_  = A233 & ~A232;
  assign \new_[43632]_  = \new_[43631]_  & \new_[43628]_ ;
  assign \new_[43633]_  = \new_[43632]_  & \new_[43625]_ ;
  assign \new_[43636]_  = A235 & A234;
  assign \new_[43639]_  = ~A269 & ~A267;
  assign \new_[43640]_  = \new_[43639]_  & \new_[43636]_ ;
  assign \new_[43643]_  = ~A299 & A298;
  assign \new_[43646]_  = A301 & A300;
  assign \new_[43647]_  = \new_[43646]_  & \new_[43643]_ ;
  assign \new_[43648]_  = \new_[43647]_  & \new_[43640]_ ;
  assign \new_[43652]_  = ~A168 & ~A169;
  assign \new_[43653]_  = ~A170 & \new_[43652]_ ;
  assign \new_[43656]_  = A166 & ~A167;
  assign \new_[43659]_  = A233 & ~A232;
  assign \new_[43660]_  = \new_[43659]_  & \new_[43656]_ ;
  assign \new_[43661]_  = \new_[43660]_  & \new_[43653]_ ;
  assign \new_[43664]_  = A235 & A234;
  assign \new_[43667]_  = ~A269 & ~A267;
  assign \new_[43668]_  = \new_[43667]_  & \new_[43664]_ ;
  assign \new_[43671]_  = ~A299 & A298;
  assign \new_[43674]_  = ~A302 & A300;
  assign \new_[43675]_  = \new_[43674]_  & \new_[43671]_ ;
  assign \new_[43676]_  = \new_[43675]_  & \new_[43668]_ ;
  assign \new_[43680]_  = ~A168 & ~A169;
  assign \new_[43681]_  = ~A170 & \new_[43680]_ ;
  assign \new_[43684]_  = A166 & ~A167;
  assign \new_[43687]_  = A233 & ~A232;
  assign \new_[43688]_  = \new_[43687]_  & \new_[43684]_ ;
  assign \new_[43689]_  = \new_[43688]_  & \new_[43681]_ ;
  assign \new_[43692]_  = A235 & A234;
  assign \new_[43695]_  = ~A269 & ~A267;
  assign \new_[43696]_  = \new_[43695]_  & \new_[43692]_ ;
  assign \new_[43699]_  = A299 & ~A298;
  assign \new_[43702]_  = A301 & A300;
  assign \new_[43703]_  = \new_[43702]_  & \new_[43699]_ ;
  assign \new_[43704]_  = \new_[43703]_  & \new_[43696]_ ;
  assign \new_[43708]_  = ~A168 & ~A169;
  assign \new_[43709]_  = ~A170 & \new_[43708]_ ;
  assign \new_[43712]_  = A166 & ~A167;
  assign \new_[43715]_  = A233 & ~A232;
  assign \new_[43716]_  = \new_[43715]_  & \new_[43712]_ ;
  assign \new_[43717]_  = \new_[43716]_  & \new_[43709]_ ;
  assign \new_[43720]_  = A235 & A234;
  assign \new_[43723]_  = ~A269 & ~A267;
  assign \new_[43724]_  = \new_[43723]_  & \new_[43720]_ ;
  assign \new_[43727]_  = A299 & ~A298;
  assign \new_[43730]_  = ~A302 & A300;
  assign \new_[43731]_  = \new_[43730]_  & \new_[43727]_ ;
  assign \new_[43732]_  = \new_[43731]_  & \new_[43724]_ ;
  assign \new_[43736]_  = ~A168 & ~A169;
  assign \new_[43737]_  = ~A170 & \new_[43736]_ ;
  assign \new_[43740]_  = A166 & ~A167;
  assign \new_[43743]_  = A233 & ~A232;
  assign \new_[43744]_  = \new_[43743]_  & \new_[43740]_ ;
  assign \new_[43745]_  = \new_[43744]_  & \new_[43737]_ ;
  assign \new_[43748]_  = A235 & A234;
  assign \new_[43751]_  = A266 & A265;
  assign \new_[43752]_  = \new_[43751]_  & \new_[43748]_ ;
  assign \new_[43755]_  = ~A299 & A298;
  assign \new_[43758]_  = A301 & A300;
  assign \new_[43759]_  = \new_[43758]_  & \new_[43755]_ ;
  assign \new_[43760]_  = \new_[43759]_  & \new_[43752]_ ;
  assign \new_[43764]_  = ~A168 & ~A169;
  assign \new_[43765]_  = ~A170 & \new_[43764]_ ;
  assign \new_[43768]_  = A166 & ~A167;
  assign \new_[43771]_  = A233 & ~A232;
  assign \new_[43772]_  = \new_[43771]_  & \new_[43768]_ ;
  assign \new_[43773]_  = \new_[43772]_  & \new_[43765]_ ;
  assign \new_[43776]_  = A235 & A234;
  assign \new_[43779]_  = A266 & A265;
  assign \new_[43780]_  = \new_[43779]_  & \new_[43776]_ ;
  assign \new_[43783]_  = ~A299 & A298;
  assign \new_[43786]_  = ~A302 & A300;
  assign \new_[43787]_  = \new_[43786]_  & \new_[43783]_ ;
  assign \new_[43788]_  = \new_[43787]_  & \new_[43780]_ ;
  assign \new_[43792]_  = ~A168 & ~A169;
  assign \new_[43793]_  = ~A170 & \new_[43792]_ ;
  assign \new_[43796]_  = A166 & ~A167;
  assign \new_[43799]_  = A233 & ~A232;
  assign \new_[43800]_  = \new_[43799]_  & \new_[43796]_ ;
  assign \new_[43801]_  = \new_[43800]_  & \new_[43793]_ ;
  assign \new_[43804]_  = A235 & A234;
  assign \new_[43807]_  = A266 & A265;
  assign \new_[43808]_  = \new_[43807]_  & \new_[43804]_ ;
  assign \new_[43811]_  = A299 & ~A298;
  assign \new_[43814]_  = A301 & A300;
  assign \new_[43815]_  = \new_[43814]_  & \new_[43811]_ ;
  assign \new_[43816]_  = \new_[43815]_  & \new_[43808]_ ;
  assign \new_[43820]_  = ~A168 & ~A169;
  assign \new_[43821]_  = ~A170 & \new_[43820]_ ;
  assign \new_[43824]_  = A166 & ~A167;
  assign \new_[43827]_  = A233 & ~A232;
  assign \new_[43828]_  = \new_[43827]_  & \new_[43824]_ ;
  assign \new_[43829]_  = \new_[43828]_  & \new_[43821]_ ;
  assign \new_[43832]_  = A235 & A234;
  assign \new_[43835]_  = A266 & A265;
  assign \new_[43836]_  = \new_[43835]_  & \new_[43832]_ ;
  assign \new_[43839]_  = A299 & ~A298;
  assign \new_[43842]_  = ~A302 & A300;
  assign \new_[43843]_  = \new_[43842]_  & \new_[43839]_ ;
  assign \new_[43844]_  = \new_[43843]_  & \new_[43836]_ ;
  assign \new_[43848]_  = ~A168 & ~A169;
  assign \new_[43849]_  = ~A170 & \new_[43848]_ ;
  assign \new_[43852]_  = A166 & ~A167;
  assign \new_[43855]_  = A233 & ~A232;
  assign \new_[43856]_  = \new_[43855]_  & \new_[43852]_ ;
  assign \new_[43857]_  = \new_[43856]_  & \new_[43849]_ ;
  assign \new_[43860]_  = A235 & A234;
  assign \new_[43863]_  = ~A266 & ~A265;
  assign \new_[43864]_  = \new_[43863]_  & \new_[43860]_ ;
  assign \new_[43867]_  = ~A299 & A298;
  assign \new_[43870]_  = A301 & A300;
  assign \new_[43871]_  = \new_[43870]_  & \new_[43867]_ ;
  assign \new_[43872]_  = \new_[43871]_  & \new_[43864]_ ;
  assign \new_[43876]_  = ~A168 & ~A169;
  assign \new_[43877]_  = ~A170 & \new_[43876]_ ;
  assign \new_[43880]_  = A166 & ~A167;
  assign \new_[43883]_  = A233 & ~A232;
  assign \new_[43884]_  = \new_[43883]_  & \new_[43880]_ ;
  assign \new_[43885]_  = \new_[43884]_  & \new_[43877]_ ;
  assign \new_[43888]_  = A235 & A234;
  assign \new_[43891]_  = ~A266 & ~A265;
  assign \new_[43892]_  = \new_[43891]_  & \new_[43888]_ ;
  assign \new_[43895]_  = ~A299 & A298;
  assign \new_[43898]_  = ~A302 & A300;
  assign \new_[43899]_  = \new_[43898]_  & \new_[43895]_ ;
  assign \new_[43900]_  = \new_[43899]_  & \new_[43892]_ ;
  assign \new_[43904]_  = ~A168 & ~A169;
  assign \new_[43905]_  = ~A170 & \new_[43904]_ ;
  assign \new_[43908]_  = A166 & ~A167;
  assign \new_[43911]_  = A233 & ~A232;
  assign \new_[43912]_  = \new_[43911]_  & \new_[43908]_ ;
  assign \new_[43913]_  = \new_[43912]_  & \new_[43905]_ ;
  assign \new_[43916]_  = A235 & A234;
  assign \new_[43919]_  = ~A266 & ~A265;
  assign \new_[43920]_  = \new_[43919]_  & \new_[43916]_ ;
  assign \new_[43923]_  = A299 & ~A298;
  assign \new_[43926]_  = A301 & A300;
  assign \new_[43927]_  = \new_[43926]_  & \new_[43923]_ ;
  assign \new_[43928]_  = \new_[43927]_  & \new_[43920]_ ;
  assign \new_[43932]_  = ~A168 & ~A169;
  assign \new_[43933]_  = ~A170 & \new_[43932]_ ;
  assign \new_[43936]_  = A166 & ~A167;
  assign \new_[43939]_  = A233 & ~A232;
  assign \new_[43940]_  = \new_[43939]_  & \new_[43936]_ ;
  assign \new_[43941]_  = \new_[43940]_  & \new_[43933]_ ;
  assign \new_[43944]_  = A235 & A234;
  assign \new_[43947]_  = ~A266 & ~A265;
  assign \new_[43948]_  = \new_[43947]_  & \new_[43944]_ ;
  assign \new_[43951]_  = A299 & ~A298;
  assign \new_[43954]_  = ~A302 & A300;
  assign \new_[43955]_  = \new_[43954]_  & \new_[43951]_ ;
  assign \new_[43956]_  = \new_[43955]_  & \new_[43948]_ ;
  assign \new_[43960]_  = ~A168 & ~A169;
  assign \new_[43961]_  = ~A170 & \new_[43960]_ ;
  assign \new_[43964]_  = A166 & ~A167;
  assign \new_[43967]_  = A233 & ~A232;
  assign \new_[43968]_  = \new_[43967]_  & \new_[43964]_ ;
  assign \new_[43969]_  = \new_[43968]_  & \new_[43961]_ ;
  assign \new_[43972]_  = ~A236 & A234;
  assign \new_[43975]_  = A268 & ~A267;
  assign \new_[43976]_  = \new_[43975]_  & \new_[43972]_ ;
  assign \new_[43979]_  = ~A299 & A298;
  assign \new_[43982]_  = A301 & A300;
  assign \new_[43983]_  = \new_[43982]_  & \new_[43979]_ ;
  assign \new_[43984]_  = \new_[43983]_  & \new_[43976]_ ;
  assign \new_[43988]_  = ~A168 & ~A169;
  assign \new_[43989]_  = ~A170 & \new_[43988]_ ;
  assign \new_[43992]_  = A166 & ~A167;
  assign \new_[43995]_  = A233 & ~A232;
  assign \new_[43996]_  = \new_[43995]_  & \new_[43992]_ ;
  assign \new_[43997]_  = \new_[43996]_  & \new_[43989]_ ;
  assign \new_[44000]_  = ~A236 & A234;
  assign \new_[44003]_  = A268 & ~A267;
  assign \new_[44004]_  = \new_[44003]_  & \new_[44000]_ ;
  assign \new_[44007]_  = ~A299 & A298;
  assign \new_[44010]_  = ~A302 & A300;
  assign \new_[44011]_  = \new_[44010]_  & \new_[44007]_ ;
  assign \new_[44012]_  = \new_[44011]_  & \new_[44004]_ ;
  assign \new_[44016]_  = ~A168 & ~A169;
  assign \new_[44017]_  = ~A170 & \new_[44016]_ ;
  assign \new_[44020]_  = A166 & ~A167;
  assign \new_[44023]_  = A233 & ~A232;
  assign \new_[44024]_  = \new_[44023]_  & \new_[44020]_ ;
  assign \new_[44025]_  = \new_[44024]_  & \new_[44017]_ ;
  assign \new_[44028]_  = ~A236 & A234;
  assign \new_[44031]_  = A268 & ~A267;
  assign \new_[44032]_  = \new_[44031]_  & \new_[44028]_ ;
  assign \new_[44035]_  = A299 & ~A298;
  assign \new_[44038]_  = A301 & A300;
  assign \new_[44039]_  = \new_[44038]_  & \new_[44035]_ ;
  assign \new_[44040]_  = \new_[44039]_  & \new_[44032]_ ;
  assign \new_[44044]_  = ~A168 & ~A169;
  assign \new_[44045]_  = ~A170 & \new_[44044]_ ;
  assign \new_[44048]_  = A166 & ~A167;
  assign \new_[44051]_  = A233 & ~A232;
  assign \new_[44052]_  = \new_[44051]_  & \new_[44048]_ ;
  assign \new_[44053]_  = \new_[44052]_  & \new_[44045]_ ;
  assign \new_[44056]_  = ~A236 & A234;
  assign \new_[44059]_  = A268 & ~A267;
  assign \new_[44060]_  = \new_[44059]_  & \new_[44056]_ ;
  assign \new_[44063]_  = A299 & ~A298;
  assign \new_[44066]_  = ~A302 & A300;
  assign \new_[44067]_  = \new_[44066]_  & \new_[44063]_ ;
  assign \new_[44068]_  = \new_[44067]_  & \new_[44060]_ ;
  assign \new_[44072]_  = ~A168 & ~A169;
  assign \new_[44073]_  = ~A170 & \new_[44072]_ ;
  assign \new_[44076]_  = A166 & ~A167;
  assign \new_[44079]_  = A233 & ~A232;
  assign \new_[44080]_  = \new_[44079]_  & \new_[44076]_ ;
  assign \new_[44081]_  = \new_[44080]_  & \new_[44073]_ ;
  assign \new_[44084]_  = ~A236 & A234;
  assign \new_[44087]_  = ~A269 & ~A267;
  assign \new_[44088]_  = \new_[44087]_  & \new_[44084]_ ;
  assign \new_[44091]_  = ~A299 & A298;
  assign \new_[44094]_  = A301 & A300;
  assign \new_[44095]_  = \new_[44094]_  & \new_[44091]_ ;
  assign \new_[44096]_  = \new_[44095]_  & \new_[44088]_ ;
  assign \new_[44100]_  = ~A168 & ~A169;
  assign \new_[44101]_  = ~A170 & \new_[44100]_ ;
  assign \new_[44104]_  = A166 & ~A167;
  assign \new_[44107]_  = A233 & ~A232;
  assign \new_[44108]_  = \new_[44107]_  & \new_[44104]_ ;
  assign \new_[44109]_  = \new_[44108]_  & \new_[44101]_ ;
  assign \new_[44112]_  = ~A236 & A234;
  assign \new_[44115]_  = ~A269 & ~A267;
  assign \new_[44116]_  = \new_[44115]_  & \new_[44112]_ ;
  assign \new_[44119]_  = ~A299 & A298;
  assign \new_[44122]_  = ~A302 & A300;
  assign \new_[44123]_  = \new_[44122]_  & \new_[44119]_ ;
  assign \new_[44124]_  = \new_[44123]_  & \new_[44116]_ ;
  assign \new_[44128]_  = ~A168 & ~A169;
  assign \new_[44129]_  = ~A170 & \new_[44128]_ ;
  assign \new_[44132]_  = A166 & ~A167;
  assign \new_[44135]_  = A233 & ~A232;
  assign \new_[44136]_  = \new_[44135]_  & \new_[44132]_ ;
  assign \new_[44137]_  = \new_[44136]_  & \new_[44129]_ ;
  assign \new_[44140]_  = ~A236 & A234;
  assign \new_[44143]_  = ~A269 & ~A267;
  assign \new_[44144]_  = \new_[44143]_  & \new_[44140]_ ;
  assign \new_[44147]_  = A299 & ~A298;
  assign \new_[44150]_  = A301 & A300;
  assign \new_[44151]_  = \new_[44150]_  & \new_[44147]_ ;
  assign \new_[44152]_  = \new_[44151]_  & \new_[44144]_ ;
  assign \new_[44156]_  = ~A168 & ~A169;
  assign \new_[44157]_  = ~A170 & \new_[44156]_ ;
  assign \new_[44160]_  = A166 & ~A167;
  assign \new_[44163]_  = A233 & ~A232;
  assign \new_[44164]_  = \new_[44163]_  & \new_[44160]_ ;
  assign \new_[44165]_  = \new_[44164]_  & \new_[44157]_ ;
  assign \new_[44168]_  = ~A236 & A234;
  assign \new_[44171]_  = ~A269 & ~A267;
  assign \new_[44172]_  = \new_[44171]_  & \new_[44168]_ ;
  assign \new_[44175]_  = A299 & ~A298;
  assign \new_[44178]_  = ~A302 & A300;
  assign \new_[44179]_  = \new_[44178]_  & \new_[44175]_ ;
  assign \new_[44180]_  = \new_[44179]_  & \new_[44172]_ ;
  assign \new_[44184]_  = ~A168 & ~A169;
  assign \new_[44185]_  = ~A170 & \new_[44184]_ ;
  assign \new_[44188]_  = A166 & ~A167;
  assign \new_[44191]_  = A233 & ~A232;
  assign \new_[44192]_  = \new_[44191]_  & \new_[44188]_ ;
  assign \new_[44193]_  = \new_[44192]_  & \new_[44185]_ ;
  assign \new_[44196]_  = ~A236 & A234;
  assign \new_[44199]_  = A266 & A265;
  assign \new_[44200]_  = \new_[44199]_  & \new_[44196]_ ;
  assign \new_[44203]_  = ~A299 & A298;
  assign \new_[44206]_  = A301 & A300;
  assign \new_[44207]_  = \new_[44206]_  & \new_[44203]_ ;
  assign \new_[44208]_  = \new_[44207]_  & \new_[44200]_ ;
  assign \new_[44212]_  = ~A168 & ~A169;
  assign \new_[44213]_  = ~A170 & \new_[44212]_ ;
  assign \new_[44216]_  = A166 & ~A167;
  assign \new_[44219]_  = A233 & ~A232;
  assign \new_[44220]_  = \new_[44219]_  & \new_[44216]_ ;
  assign \new_[44221]_  = \new_[44220]_  & \new_[44213]_ ;
  assign \new_[44224]_  = ~A236 & A234;
  assign \new_[44227]_  = A266 & A265;
  assign \new_[44228]_  = \new_[44227]_  & \new_[44224]_ ;
  assign \new_[44231]_  = ~A299 & A298;
  assign \new_[44234]_  = ~A302 & A300;
  assign \new_[44235]_  = \new_[44234]_  & \new_[44231]_ ;
  assign \new_[44236]_  = \new_[44235]_  & \new_[44228]_ ;
  assign \new_[44240]_  = ~A168 & ~A169;
  assign \new_[44241]_  = ~A170 & \new_[44240]_ ;
  assign \new_[44244]_  = A166 & ~A167;
  assign \new_[44247]_  = A233 & ~A232;
  assign \new_[44248]_  = \new_[44247]_  & \new_[44244]_ ;
  assign \new_[44249]_  = \new_[44248]_  & \new_[44241]_ ;
  assign \new_[44252]_  = ~A236 & A234;
  assign \new_[44255]_  = A266 & A265;
  assign \new_[44256]_  = \new_[44255]_  & \new_[44252]_ ;
  assign \new_[44259]_  = A299 & ~A298;
  assign \new_[44262]_  = A301 & A300;
  assign \new_[44263]_  = \new_[44262]_  & \new_[44259]_ ;
  assign \new_[44264]_  = \new_[44263]_  & \new_[44256]_ ;
  assign \new_[44268]_  = ~A168 & ~A169;
  assign \new_[44269]_  = ~A170 & \new_[44268]_ ;
  assign \new_[44272]_  = A166 & ~A167;
  assign \new_[44275]_  = A233 & ~A232;
  assign \new_[44276]_  = \new_[44275]_  & \new_[44272]_ ;
  assign \new_[44277]_  = \new_[44276]_  & \new_[44269]_ ;
  assign \new_[44280]_  = ~A236 & A234;
  assign \new_[44283]_  = A266 & A265;
  assign \new_[44284]_  = \new_[44283]_  & \new_[44280]_ ;
  assign \new_[44287]_  = A299 & ~A298;
  assign \new_[44290]_  = ~A302 & A300;
  assign \new_[44291]_  = \new_[44290]_  & \new_[44287]_ ;
  assign \new_[44292]_  = \new_[44291]_  & \new_[44284]_ ;
  assign \new_[44296]_  = ~A168 & ~A169;
  assign \new_[44297]_  = ~A170 & \new_[44296]_ ;
  assign \new_[44300]_  = A166 & ~A167;
  assign \new_[44303]_  = A233 & ~A232;
  assign \new_[44304]_  = \new_[44303]_  & \new_[44300]_ ;
  assign \new_[44305]_  = \new_[44304]_  & \new_[44297]_ ;
  assign \new_[44308]_  = ~A236 & A234;
  assign \new_[44311]_  = ~A266 & ~A265;
  assign \new_[44312]_  = \new_[44311]_  & \new_[44308]_ ;
  assign \new_[44315]_  = ~A299 & A298;
  assign \new_[44318]_  = A301 & A300;
  assign \new_[44319]_  = \new_[44318]_  & \new_[44315]_ ;
  assign \new_[44320]_  = \new_[44319]_  & \new_[44312]_ ;
  assign \new_[44324]_  = ~A168 & ~A169;
  assign \new_[44325]_  = ~A170 & \new_[44324]_ ;
  assign \new_[44328]_  = A166 & ~A167;
  assign \new_[44331]_  = A233 & ~A232;
  assign \new_[44332]_  = \new_[44331]_  & \new_[44328]_ ;
  assign \new_[44333]_  = \new_[44332]_  & \new_[44325]_ ;
  assign \new_[44336]_  = ~A236 & A234;
  assign \new_[44339]_  = ~A266 & ~A265;
  assign \new_[44340]_  = \new_[44339]_  & \new_[44336]_ ;
  assign \new_[44343]_  = ~A299 & A298;
  assign \new_[44346]_  = ~A302 & A300;
  assign \new_[44347]_  = \new_[44346]_  & \new_[44343]_ ;
  assign \new_[44348]_  = \new_[44347]_  & \new_[44340]_ ;
  assign \new_[44352]_  = ~A168 & ~A169;
  assign \new_[44353]_  = ~A170 & \new_[44352]_ ;
  assign \new_[44356]_  = A166 & ~A167;
  assign \new_[44359]_  = A233 & ~A232;
  assign \new_[44360]_  = \new_[44359]_  & \new_[44356]_ ;
  assign \new_[44361]_  = \new_[44360]_  & \new_[44353]_ ;
  assign \new_[44364]_  = ~A236 & A234;
  assign \new_[44367]_  = ~A266 & ~A265;
  assign \new_[44368]_  = \new_[44367]_  & \new_[44364]_ ;
  assign \new_[44371]_  = A299 & ~A298;
  assign \new_[44374]_  = A301 & A300;
  assign \new_[44375]_  = \new_[44374]_  & \new_[44371]_ ;
  assign \new_[44376]_  = \new_[44375]_  & \new_[44368]_ ;
  assign \new_[44380]_  = ~A168 & ~A169;
  assign \new_[44381]_  = ~A170 & \new_[44380]_ ;
  assign \new_[44384]_  = A166 & ~A167;
  assign \new_[44387]_  = A233 & ~A232;
  assign \new_[44388]_  = \new_[44387]_  & \new_[44384]_ ;
  assign \new_[44389]_  = \new_[44388]_  & \new_[44381]_ ;
  assign \new_[44392]_  = ~A236 & A234;
  assign \new_[44395]_  = ~A266 & ~A265;
  assign \new_[44396]_  = \new_[44395]_  & \new_[44392]_ ;
  assign \new_[44399]_  = A299 & ~A298;
  assign \new_[44402]_  = ~A302 & A300;
  assign \new_[44403]_  = \new_[44402]_  & \new_[44399]_ ;
  assign \new_[44404]_  = \new_[44403]_  & \new_[44396]_ ;
  assign \new_[44408]_  = ~A168 & ~A169;
  assign \new_[44409]_  = ~A170 & \new_[44408]_ ;
  assign \new_[44412]_  = A166 & ~A167;
  assign \new_[44415]_  = ~A233 & A232;
  assign \new_[44416]_  = \new_[44415]_  & \new_[44412]_ ;
  assign \new_[44417]_  = \new_[44416]_  & \new_[44409]_ ;
  assign \new_[44420]_  = A235 & A234;
  assign \new_[44423]_  = A268 & ~A267;
  assign \new_[44424]_  = \new_[44423]_  & \new_[44420]_ ;
  assign \new_[44427]_  = ~A299 & A298;
  assign \new_[44430]_  = A301 & A300;
  assign \new_[44431]_  = \new_[44430]_  & \new_[44427]_ ;
  assign \new_[44432]_  = \new_[44431]_  & \new_[44424]_ ;
  assign \new_[44436]_  = ~A168 & ~A169;
  assign \new_[44437]_  = ~A170 & \new_[44436]_ ;
  assign \new_[44440]_  = A166 & ~A167;
  assign \new_[44443]_  = ~A233 & A232;
  assign \new_[44444]_  = \new_[44443]_  & \new_[44440]_ ;
  assign \new_[44445]_  = \new_[44444]_  & \new_[44437]_ ;
  assign \new_[44448]_  = A235 & A234;
  assign \new_[44451]_  = A268 & ~A267;
  assign \new_[44452]_  = \new_[44451]_  & \new_[44448]_ ;
  assign \new_[44455]_  = ~A299 & A298;
  assign \new_[44458]_  = ~A302 & A300;
  assign \new_[44459]_  = \new_[44458]_  & \new_[44455]_ ;
  assign \new_[44460]_  = \new_[44459]_  & \new_[44452]_ ;
  assign \new_[44464]_  = ~A168 & ~A169;
  assign \new_[44465]_  = ~A170 & \new_[44464]_ ;
  assign \new_[44468]_  = A166 & ~A167;
  assign \new_[44471]_  = ~A233 & A232;
  assign \new_[44472]_  = \new_[44471]_  & \new_[44468]_ ;
  assign \new_[44473]_  = \new_[44472]_  & \new_[44465]_ ;
  assign \new_[44476]_  = A235 & A234;
  assign \new_[44479]_  = A268 & ~A267;
  assign \new_[44480]_  = \new_[44479]_  & \new_[44476]_ ;
  assign \new_[44483]_  = A299 & ~A298;
  assign \new_[44486]_  = A301 & A300;
  assign \new_[44487]_  = \new_[44486]_  & \new_[44483]_ ;
  assign \new_[44488]_  = \new_[44487]_  & \new_[44480]_ ;
  assign \new_[44492]_  = ~A168 & ~A169;
  assign \new_[44493]_  = ~A170 & \new_[44492]_ ;
  assign \new_[44496]_  = A166 & ~A167;
  assign \new_[44499]_  = ~A233 & A232;
  assign \new_[44500]_  = \new_[44499]_  & \new_[44496]_ ;
  assign \new_[44501]_  = \new_[44500]_  & \new_[44493]_ ;
  assign \new_[44504]_  = A235 & A234;
  assign \new_[44507]_  = A268 & ~A267;
  assign \new_[44508]_  = \new_[44507]_  & \new_[44504]_ ;
  assign \new_[44511]_  = A299 & ~A298;
  assign \new_[44514]_  = ~A302 & A300;
  assign \new_[44515]_  = \new_[44514]_  & \new_[44511]_ ;
  assign \new_[44516]_  = \new_[44515]_  & \new_[44508]_ ;
  assign \new_[44520]_  = ~A168 & ~A169;
  assign \new_[44521]_  = ~A170 & \new_[44520]_ ;
  assign \new_[44524]_  = A166 & ~A167;
  assign \new_[44527]_  = ~A233 & A232;
  assign \new_[44528]_  = \new_[44527]_  & \new_[44524]_ ;
  assign \new_[44529]_  = \new_[44528]_  & \new_[44521]_ ;
  assign \new_[44532]_  = A235 & A234;
  assign \new_[44535]_  = ~A269 & ~A267;
  assign \new_[44536]_  = \new_[44535]_  & \new_[44532]_ ;
  assign \new_[44539]_  = ~A299 & A298;
  assign \new_[44542]_  = A301 & A300;
  assign \new_[44543]_  = \new_[44542]_  & \new_[44539]_ ;
  assign \new_[44544]_  = \new_[44543]_  & \new_[44536]_ ;
  assign \new_[44548]_  = ~A168 & ~A169;
  assign \new_[44549]_  = ~A170 & \new_[44548]_ ;
  assign \new_[44552]_  = A166 & ~A167;
  assign \new_[44555]_  = ~A233 & A232;
  assign \new_[44556]_  = \new_[44555]_  & \new_[44552]_ ;
  assign \new_[44557]_  = \new_[44556]_  & \new_[44549]_ ;
  assign \new_[44560]_  = A235 & A234;
  assign \new_[44563]_  = ~A269 & ~A267;
  assign \new_[44564]_  = \new_[44563]_  & \new_[44560]_ ;
  assign \new_[44567]_  = ~A299 & A298;
  assign \new_[44570]_  = ~A302 & A300;
  assign \new_[44571]_  = \new_[44570]_  & \new_[44567]_ ;
  assign \new_[44572]_  = \new_[44571]_  & \new_[44564]_ ;
  assign \new_[44576]_  = ~A168 & ~A169;
  assign \new_[44577]_  = ~A170 & \new_[44576]_ ;
  assign \new_[44580]_  = A166 & ~A167;
  assign \new_[44583]_  = ~A233 & A232;
  assign \new_[44584]_  = \new_[44583]_  & \new_[44580]_ ;
  assign \new_[44585]_  = \new_[44584]_  & \new_[44577]_ ;
  assign \new_[44588]_  = A235 & A234;
  assign \new_[44591]_  = ~A269 & ~A267;
  assign \new_[44592]_  = \new_[44591]_  & \new_[44588]_ ;
  assign \new_[44595]_  = A299 & ~A298;
  assign \new_[44598]_  = A301 & A300;
  assign \new_[44599]_  = \new_[44598]_  & \new_[44595]_ ;
  assign \new_[44600]_  = \new_[44599]_  & \new_[44592]_ ;
  assign \new_[44604]_  = ~A168 & ~A169;
  assign \new_[44605]_  = ~A170 & \new_[44604]_ ;
  assign \new_[44608]_  = A166 & ~A167;
  assign \new_[44611]_  = ~A233 & A232;
  assign \new_[44612]_  = \new_[44611]_  & \new_[44608]_ ;
  assign \new_[44613]_  = \new_[44612]_  & \new_[44605]_ ;
  assign \new_[44616]_  = A235 & A234;
  assign \new_[44619]_  = ~A269 & ~A267;
  assign \new_[44620]_  = \new_[44619]_  & \new_[44616]_ ;
  assign \new_[44623]_  = A299 & ~A298;
  assign \new_[44626]_  = ~A302 & A300;
  assign \new_[44627]_  = \new_[44626]_  & \new_[44623]_ ;
  assign \new_[44628]_  = \new_[44627]_  & \new_[44620]_ ;
  assign \new_[44632]_  = ~A168 & ~A169;
  assign \new_[44633]_  = ~A170 & \new_[44632]_ ;
  assign \new_[44636]_  = A166 & ~A167;
  assign \new_[44639]_  = ~A233 & A232;
  assign \new_[44640]_  = \new_[44639]_  & \new_[44636]_ ;
  assign \new_[44641]_  = \new_[44640]_  & \new_[44633]_ ;
  assign \new_[44644]_  = A235 & A234;
  assign \new_[44647]_  = A266 & A265;
  assign \new_[44648]_  = \new_[44647]_  & \new_[44644]_ ;
  assign \new_[44651]_  = ~A299 & A298;
  assign \new_[44654]_  = A301 & A300;
  assign \new_[44655]_  = \new_[44654]_  & \new_[44651]_ ;
  assign \new_[44656]_  = \new_[44655]_  & \new_[44648]_ ;
  assign \new_[44660]_  = ~A168 & ~A169;
  assign \new_[44661]_  = ~A170 & \new_[44660]_ ;
  assign \new_[44664]_  = A166 & ~A167;
  assign \new_[44667]_  = ~A233 & A232;
  assign \new_[44668]_  = \new_[44667]_  & \new_[44664]_ ;
  assign \new_[44669]_  = \new_[44668]_  & \new_[44661]_ ;
  assign \new_[44672]_  = A235 & A234;
  assign \new_[44675]_  = A266 & A265;
  assign \new_[44676]_  = \new_[44675]_  & \new_[44672]_ ;
  assign \new_[44679]_  = ~A299 & A298;
  assign \new_[44682]_  = ~A302 & A300;
  assign \new_[44683]_  = \new_[44682]_  & \new_[44679]_ ;
  assign \new_[44684]_  = \new_[44683]_  & \new_[44676]_ ;
  assign \new_[44688]_  = ~A168 & ~A169;
  assign \new_[44689]_  = ~A170 & \new_[44688]_ ;
  assign \new_[44692]_  = A166 & ~A167;
  assign \new_[44695]_  = ~A233 & A232;
  assign \new_[44696]_  = \new_[44695]_  & \new_[44692]_ ;
  assign \new_[44697]_  = \new_[44696]_  & \new_[44689]_ ;
  assign \new_[44700]_  = A235 & A234;
  assign \new_[44703]_  = A266 & A265;
  assign \new_[44704]_  = \new_[44703]_  & \new_[44700]_ ;
  assign \new_[44707]_  = A299 & ~A298;
  assign \new_[44710]_  = A301 & A300;
  assign \new_[44711]_  = \new_[44710]_  & \new_[44707]_ ;
  assign \new_[44712]_  = \new_[44711]_  & \new_[44704]_ ;
  assign \new_[44716]_  = ~A168 & ~A169;
  assign \new_[44717]_  = ~A170 & \new_[44716]_ ;
  assign \new_[44720]_  = A166 & ~A167;
  assign \new_[44723]_  = ~A233 & A232;
  assign \new_[44724]_  = \new_[44723]_  & \new_[44720]_ ;
  assign \new_[44725]_  = \new_[44724]_  & \new_[44717]_ ;
  assign \new_[44728]_  = A235 & A234;
  assign \new_[44731]_  = A266 & A265;
  assign \new_[44732]_  = \new_[44731]_  & \new_[44728]_ ;
  assign \new_[44735]_  = A299 & ~A298;
  assign \new_[44738]_  = ~A302 & A300;
  assign \new_[44739]_  = \new_[44738]_  & \new_[44735]_ ;
  assign \new_[44740]_  = \new_[44739]_  & \new_[44732]_ ;
  assign \new_[44744]_  = ~A168 & ~A169;
  assign \new_[44745]_  = ~A170 & \new_[44744]_ ;
  assign \new_[44748]_  = A166 & ~A167;
  assign \new_[44751]_  = ~A233 & A232;
  assign \new_[44752]_  = \new_[44751]_  & \new_[44748]_ ;
  assign \new_[44753]_  = \new_[44752]_  & \new_[44745]_ ;
  assign \new_[44756]_  = A235 & A234;
  assign \new_[44759]_  = ~A266 & ~A265;
  assign \new_[44760]_  = \new_[44759]_  & \new_[44756]_ ;
  assign \new_[44763]_  = ~A299 & A298;
  assign \new_[44766]_  = A301 & A300;
  assign \new_[44767]_  = \new_[44766]_  & \new_[44763]_ ;
  assign \new_[44768]_  = \new_[44767]_  & \new_[44760]_ ;
  assign \new_[44772]_  = ~A168 & ~A169;
  assign \new_[44773]_  = ~A170 & \new_[44772]_ ;
  assign \new_[44776]_  = A166 & ~A167;
  assign \new_[44779]_  = ~A233 & A232;
  assign \new_[44780]_  = \new_[44779]_  & \new_[44776]_ ;
  assign \new_[44781]_  = \new_[44780]_  & \new_[44773]_ ;
  assign \new_[44784]_  = A235 & A234;
  assign \new_[44787]_  = ~A266 & ~A265;
  assign \new_[44788]_  = \new_[44787]_  & \new_[44784]_ ;
  assign \new_[44791]_  = ~A299 & A298;
  assign \new_[44794]_  = ~A302 & A300;
  assign \new_[44795]_  = \new_[44794]_  & \new_[44791]_ ;
  assign \new_[44796]_  = \new_[44795]_  & \new_[44788]_ ;
  assign \new_[44800]_  = ~A168 & ~A169;
  assign \new_[44801]_  = ~A170 & \new_[44800]_ ;
  assign \new_[44804]_  = A166 & ~A167;
  assign \new_[44807]_  = ~A233 & A232;
  assign \new_[44808]_  = \new_[44807]_  & \new_[44804]_ ;
  assign \new_[44809]_  = \new_[44808]_  & \new_[44801]_ ;
  assign \new_[44812]_  = A235 & A234;
  assign \new_[44815]_  = ~A266 & ~A265;
  assign \new_[44816]_  = \new_[44815]_  & \new_[44812]_ ;
  assign \new_[44819]_  = A299 & ~A298;
  assign \new_[44822]_  = A301 & A300;
  assign \new_[44823]_  = \new_[44822]_  & \new_[44819]_ ;
  assign \new_[44824]_  = \new_[44823]_  & \new_[44816]_ ;
  assign \new_[44828]_  = ~A168 & ~A169;
  assign \new_[44829]_  = ~A170 & \new_[44828]_ ;
  assign \new_[44832]_  = A166 & ~A167;
  assign \new_[44835]_  = ~A233 & A232;
  assign \new_[44836]_  = \new_[44835]_  & \new_[44832]_ ;
  assign \new_[44837]_  = \new_[44836]_  & \new_[44829]_ ;
  assign \new_[44840]_  = A235 & A234;
  assign \new_[44843]_  = ~A266 & ~A265;
  assign \new_[44844]_  = \new_[44843]_  & \new_[44840]_ ;
  assign \new_[44847]_  = A299 & ~A298;
  assign \new_[44850]_  = ~A302 & A300;
  assign \new_[44851]_  = \new_[44850]_  & \new_[44847]_ ;
  assign \new_[44852]_  = \new_[44851]_  & \new_[44844]_ ;
  assign \new_[44856]_  = ~A168 & ~A169;
  assign \new_[44857]_  = ~A170 & \new_[44856]_ ;
  assign \new_[44860]_  = A166 & ~A167;
  assign \new_[44863]_  = ~A233 & A232;
  assign \new_[44864]_  = \new_[44863]_  & \new_[44860]_ ;
  assign \new_[44865]_  = \new_[44864]_  & \new_[44857]_ ;
  assign \new_[44868]_  = ~A236 & A234;
  assign \new_[44871]_  = A268 & ~A267;
  assign \new_[44872]_  = \new_[44871]_  & \new_[44868]_ ;
  assign \new_[44875]_  = ~A299 & A298;
  assign \new_[44878]_  = A301 & A300;
  assign \new_[44879]_  = \new_[44878]_  & \new_[44875]_ ;
  assign \new_[44880]_  = \new_[44879]_  & \new_[44872]_ ;
  assign \new_[44884]_  = ~A168 & ~A169;
  assign \new_[44885]_  = ~A170 & \new_[44884]_ ;
  assign \new_[44888]_  = A166 & ~A167;
  assign \new_[44891]_  = ~A233 & A232;
  assign \new_[44892]_  = \new_[44891]_  & \new_[44888]_ ;
  assign \new_[44893]_  = \new_[44892]_  & \new_[44885]_ ;
  assign \new_[44896]_  = ~A236 & A234;
  assign \new_[44899]_  = A268 & ~A267;
  assign \new_[44900]_  = \new_[44899]_  & \new_[44896]_ ;
  assign \new_[44903]_  = ~A299 & A298;
  assign \new_[44906]_  = ~A302 & A300;
  assign \new_[44907]_  = \new_[44906]_  & \new_[44903]_ ;
  assign \new_[44908]_  = \new_[44907]_  & \new_[44900]_ ;
  assign \new_[44912]_  = ~A168 & ~A169;
  assign \new_[44913]_  = ~A170 & \new_[44912]_ ;
  assign \new_[44916]_  = A166 & ~A167;
  assign \new_[44919]_  = ~A233 & A232;
  assign \new_[44920]_  = \new_[44919]_  & \new_[44916]_ ;
  assign \new_[44921]_  = \new_[44920]_  & \new_[44913]_ ;
  assign \new_[44924]_  = ~A236 & A234;
  assign \new_[44927]_  = A268 & ~A267;
  assign \new_[44928]_  = \new_[44927]_  & \new_[44924]_ ;
  assign \new_[44931]_  = A299 & ~A298;
  assign \new_[44934]_  = A301 & A300;
  assign \new_[44935]_  = \new_[44934]_  & \new_[44931]_ ;
  assign \new_[44936]_  = \new_[44935]_  & \new_[44928]_ ;
  assign \new_[44940]_  = ~A168 & ~A169;
  assign \new_[44941]_  = ~A170 & \new_[44940]_ ;
  assign \new_[44944]_  = A166 & ~A167;
  assign \new_[44947]_  = ~A233 & A232;
  assign \new_[44948]_  = \new_[44947]_  & \new_[44944]_ ;
  assign \new_[44949]_  = \new_[44948]_  & \new_[44941]_ ;
  assign \new_[44952]_  = ~A236 & A234;
  assign \new_[44955]_  = A268 & ~A267;
  assign \new_[44956]_  = \new_[44955]_  & \new_[44952]_ ;
  assign \new_[44959]_  = A299 & ~A298;
  assign \new_[44962]_  = ~A302 & A300;
  assign \new_[44963]_  = \new_[44962]_  & \new_[44959]_ ;
  assign \new_[44964]_  = \new_[44963]_  & \new_[44956]_ ;
  assign \new_[44968]_  = ~A168 & ~A169;
  assign \new_[44969]_  = ~A170 & \new_[44968]_ ;
  assign \new_[44972]_  = A166 & ~A167;
  assign \new_[44975]_  = ~A233 & A232;
  assign \new_[44976]_  = \new_[44975]_  & \new_[44972]_ ;
  assign \new_[44977]_  = \new_[44976]_  & \new_[44969]_ ;
  assign \new_[44980]_  = ~A236 & A234;
  assign \new_[44983]_  = ~A269 & ~A267;
  assign \new_[44984]_  = \new_[44983]_  & \new_[44980]_ ;
  assign \new_[44987]_  = ~A299 & A298;
  assign \new_[44990]_  = A301 & A300;
  assign \new_[44991]_  = \new_[44990]_  & \new_[44987]_ ;
  assign \new_[44992]_  = \new_[44991]_  & \new_[44984]_ ;
  assign \new_[44996]_  = ~A168 & ~A169;
  assign \new_[44997]_  = ~A170 & \new_[44996]_ ;
  assign \new_[45000]_  = A166 & ~A167;
  assign \new_[45003]_  = ~A233 & A232;
  assign \new_[45004]_  = \new_[45003]_  & \new_[45000]_ ;
  assign \new_[45005]_  = \new_[45004]_  & \new_[44997]_ ;
  assign \new_[45008]_  = ~A236 & A234;
  assign \new_[45011]_  = ~A269 & ~A267;
  assign \new_[45012]_  = \new_[45011]_  & \new_[45008]_ ;
  assign \new_[45015]_  = ~A299 & A298;
  assign \new_[45018]_  = ~A302 & A300;
  assign \new_[45019]_  = \new_[45018]_  & \new_[45015]_ ;
  assign \new_[45020]_  = \new_[45019]_  & \new_[45012]_ ;
  assign \new_[45024]_  = ~A168 & ~A169;
  assign \new_[45025]_  = ~A170 & \new_[45024]_ ;
  assign \new_[45028]_  = A166 & ~A167;
  assign \new_[45031]_  = ~A233 & A232;
  assign \new_[45032]_  = \new_[45031]_  & \new_[45028]_ ;
  assign \new_[45033]_  = \new_[45032]_  & \new_[45025]_ ;
  assign \new_[45036]_  = ~A236 & A234;
  assign \new_[45039]_  = ~A269 & ~A267;
  assign \new_[45040]_  = \new_[45039]_  & \new_[45036]_ ;
  assign \new_[45043]_  = A299 & ~A298;
  assign \new_[45046]_  = A301 & A300;
  assign \new_[45047]_  = \new_[45046]_  & \new_[45043]_ ;
  assign \new_[45048]_  = \new_[45047]_  & \new_[45040]_ ;
  assign \new_[45052]_  = ~A168 & ~A169;
  assign \new_[45053]_  = ~A170 & \new_[45052]_ ;
  assign \new_[45056]_  = A166 & ~A167;
  assign \new_[45059]_  = ~A233 & A232;
  assign \new_[45060]_  = \new_[45059]_  & \new_[45056]_ ;
  assign \new_[45061]_  = \new_[45060]_  & \new_[45053]_ ;
  assign \new_[45064]_  = ~A236 & A234;
  assign \new_[45067]_  = ~A269 & ~A267;
  assign \new_[45068]_  = \new_[45067]_  & \new_[45064]_ ;
  assign \new_[45071]_  = A299 & ~A298;
  assign \new_[45074]_  = ~A302 & A300;
  assign \new_[45075]_  = \new_[45074]_  & \new_[45071]_ ;
  assign \new_[45076]_  = \new_[45075]_  & \new_[45068]_ ;
  assign \new_[45080]_  = ~A168 & ~A169;
  assign \new_[45081]_  = ~A170 & \new_[45080]_ ;
  assign \new_[45084]_  = A166 & ~A167;
  assign \new_[45087]_  = ~A233 & A232;
  assign \new_[45088]_  = \new_[45087]_  & \new_[45084]_ ;
  assign \new_[45089]_  = \new_[45088]_  & \new_[45081]_ ;
  assign \new_[45092]_  = ~A236 & A234;
  assign \new_[45095]_  = A266 & A265;
  assign \new_[45096]_  = \new_[45095]_  & \new_[45092]_ ;
  assign \new_[45099]_  = ~A299 & A298;
  assign \new_[45102]_  = A301 & A300;
  assign \new_[45103]_  = \new_[45102]_  & \new_[45099]_ ;
  assign \new_[45104]_  = \new_[45103]_  & \new_[45096]_ ;
  assign \new_[45108]_  = ~A168 & ~A169;
  assign \new_[45109]_  = ~A170 & \new_[45108]_ ;
  assign \new_[45112]_  = A166 & ~A167;
  assign \new_[45115]_  = ~A233 & A232;
  assign \new_[45116]_  = \new_[45115]_  & \new_[45112]_ ;
  assign \new_[45117]_  = \new_[45116]_  & \new_[45109]_ ;
  assign \new_[45120]_  = ~A236 & A234;
  assign \new_[45123]_  = A266 & A265;
  assign \new_[45124]_  = \new_[45123]_  & \new_[45120]_ ;
  assign \new_[45127]_  = ~A299 & A298;
  assign \new_[45130]_  = ~A302 & A300;
  assign \new_[45131]_  = \new_[45130]_  & \new_[45127]_ ;
  assign \new_[45132]_  = \new_[45131]_  & \new_[45124]_ ;
  assign \new_[45136]_  = ~A168 & ~A169;
  assign \new_[45137]_  = ~A170 & \new_[45136]_ ;
  assign \new_[45140]_  = A166 & ~A167;
  assign \new_[45143]_  = ~A233 & A232;
  assign \new_[45144]_  = \new_[45143]_  & \new_[45140]_ ;
  assign \new_[45145]_  = \new_[45144]_  & \new_[45137]_ ;
  assign \new_[45148]_  = ~A236 & A234;
  assign \new_[45151]_  = A266 & A265;
  assign \new_[45152]_  = \new_[45151]_  & \new_[45148]_ ;
  assign \new_[45155]_  = A299 & ~A298;
  assign \new_[45158]_  = A301 & A300;
  assign \new_[45159]_  = \new_[45158]_  & \new_[45155]_ ;
  assign \new_[45160]_  = \new_[45159]_  & \new_[45152]_ ;
  assign \new_[45164]_  = ~A168 & ~A169;
  assign \new_[45165]_  = ~A170 & \new_[45164]_ ;
  assign \new_[45168]_  = A166 & ~A167;
  assign \new_[45171]_  = ~A233 & A232;
  assign \new_[45172]_  = \new_[45171]_  & \new_[45168]_ ;
  assign \new_[45173]_  = \new_[45172]_  & \new_[45165]_ ;
  assign \new_[45176]_  = ~A236 & A234;
  assign \new_[45179]_  = A266 & A265;
  assign \new_[45180]_  = \new_[45179]_  & \new_[45176]_ ;
  assign \new_[45183]_  = A299 & ~A298;
  assign \new_[45186]_  = ~A302 & A300;
  assign \new_[45187]_  = \new_[45186]_  & \new_[45183]_ ;
  assign \new_[45188]_  = \new_[45187]_  & \new_[45180]_ ;
  assign \new_[45192]_  = ~A168 & ~A169;
  assign \new_[45193]_  = ~A170 & \new_[45192]_ ;
  assign \new_[45196]_  = A166 & ~A167;
  assign \new_[45199]_  = ~A233 & A232;
  assign \new_[45200]_  = \new_[45199]_  & \new_[45196]_ ;
  assign \new_[45201]_  = \new_[45200]_  & \new_[45193]_ ;
  assign \new_[45204]_  = ~A236 & A234;
  assign \new_[45207]_  = ~A266 & ~A265;
  assign \new_[45208]_  = \new_[45207]_  & \new_[45204]_ ;
  assign \new_[45211]_  = ~A299 & A298;
  assign \new_[45214]_  = A301 & A300;
  assign \new_[45215]_  = \new_[45214]_  & \new_[45211]_ ;
  assign \new_[45216]_  = \new_[45215]_  & \new_[45208]_ ;
  assign \new_[45220]_  = ~A168 & ~A169;
  assign \new_[45221]_  = ~A170 & \new_[45220]_ ;
  assign \new_[45224]_  = A166 & ~A167;
  assign \new_[45227]_  = ~A233 & A232;
  assign \new_[45228]_  = \new_[45227]_  & \new_[45224]_ ;
  assign \new_[45229]_  = \new_[45228]_  & \new_[45221]_ ;
  assign \new_[45232]_  = ~A236 & A234;
  assign \new_[45235]_  = ~A266 & ~A265;
  assign \new_[45236]_  = \new_[45235]_  & \new_[45232]_ ;
  assign \new_[45239]_  = ~A299 & A298;
  assign \new_[45242]_  = ~A302 & A300;
  assign \new_[45243]_  = \new_[45242]_  & \new_[45239]_ ;
  assign \new_[45244]_  = \new_[45243]_  & \new_[45236]_ ;
  assign \new_[45248]_  = ~A168 & ~A169;
  assign \new_[45249]_  = ~A170 & \new_[45248]_ ;
  assign \new_[45252]_  = A166 & ~A167;
  assign \new_[45255]_  = ~A233 & A232;
  assign \new_[45256]_  = \new_[45255]_  & \new_[45252]_ ;
  assign \new_[45257]_  = \new_[45256]_  & \new_[45249]_ ;
  assign \new_[45260]_  = ~A236 & A234;
  assign \new_[45263]_  = ~A266 & ~A265;
  assign \new_[45264]_  = \new_[45263]_  & \new_[45260]_ ;
  assign \new_[45267]_  = A299 & ~A298;
  assign \new_[45270]_  = A301 & A300;
  assign \new_[45271]_  = \new_[45270]_  & \new_[45267]_ ;
  assign \new_[45272]_  = \new_[45271]_  & \new_[45264]_ ;
  assign \new_[45276]_  = ~A168 & ~A169;
  assign \new_[45277]_  = ~A170 & \new_[45276]_ ;
  assign \new_[45280]_  = A166 & ~A167;
  assign \new_[45283]_  = ~A233 & A232;
  assign \new_[45284]_  = \new_[45283]_  & \new_[45280]_ ;
  assign \new_[45285]_  = \new_[45284]_  & \new_[45277]_ ;
  assign \new_[45288]_  = ~A236 & A234;
  assign \new_[45291]_  = ~A266 & ~A265;
  assign \new_[45292]_  = \new_[45291]_  & \new_[45288]_ ;
  assign \new_[45295]_  = A299 & ~A298;
  assign \new_[45298]_  = ~A302 & A300;
  assign \new_[45299]_  = \new_[45298]_  & \new_[45295]_ ;
  assign \new_[45300]_  = \new_[45299]_  & \new_[45292]_ ;
  assign \new_[45303]_  = A200 & ~A199;
  assign \new_[45306]_  = A202 & A201;
  assign \new_[45307]_  = \new_[45306]_  & \new_[45303]_ ;
  assign \new_[45310]_  = A233 & ~A232;
  assign \new_[45313]_  = A235 & A234;
  assign \new_[45314]_  = \new_[45313]_  & \new_[45310]_ ;
  assign \new_[45315]_  = \new_[45314]_  & \new_[45307]_ ;
  assign \new_[45318]_  = ~A268 & A267;
  assign \new_[45321]_  = A298 & A269;
  assign \new_[45322]_  = \new_[45321]_  & \new_[45318]_ ;
  assign \new_[45325]_  = ~A300 & ~A299;
  assign \new_[45328]_  = A302 & ~A301;
  assign \new_[45329]_  = \new_[45328]_  & \new_[45325]_ ;
  assign \new_[45330]_  = \new_[45329]_  & \new_[45322]_ ;
  assign \new_[45333]_  = A200 & ~A199;
  assign \new_[45336]_  = A202 & A201;
  assign \new_[45337]_  = \new_[45336]_  & \new_[45333]_ ;
  assign \new_[45340]_  = A233 & ~A232;
  assign \new_[45343]_  = A235 & A234;
  assign \new_[45344]_  = \new_[45343]_  & \new_[45340]_ ;
  assign \new_[45345]_  = \new_[45344]_  & \new_[45337]_ ;
  assign \new_[45348]_  = ~A268 & A267;
  assign \new_[45351]_  = ~A298 & A269;
  assign \new_[45352]_  = \new_[45351]_  & \new_[45348]_ ;
  assign \new_[45355]_  = ~A300 & A299;
  assign \new_[45358]_  = A302 & ~A301;
  assign \new_[45359]_  = \new_[45358]_  & \new_[45355]_ ;
  assign \new_[45360]_  = \new_[45359]_  & \new_[45352]_ ;
  assign \new_[45363]_  = A200 & ~A199;
  assign \new_[45366]_  = A202 & A201;
  assign \new_[45367]_  = \new_[45366]_  & \new_[45363]_ ;
  assign \new_[45370]_  = A233 & ~A232;
  assign \new_[45373]_  = ~A236 & A234;
  assign \new_[45374]_  = \new_[45373]_  & \new_[45370]_ ;
  assign \new_[45375]_  = \new_[45374]_  & \new_[45367]_ ;
  assign \new_[45378]_  = ~A268 & A267;
  assign \new_[45381]_  = A298 & A269;
  assign \new_[45382]_  = \new_[45381]_  & \new_[45378]_ ;
  assign \new_[45385]_  = ~A300 & ~A299;
  assign \new_[45388]_  = A302 & ~A301;
  assign \new_[45389]_  = \new_[45388]_  & \new_[45385]_ ;
  assign \new_[45390]_  = \new_[45389]_  & \new_[45382]_ ;
  assign \new_[45393]_  = A200 & ~A199;
  assign \new_[45396]_  = A202 & A201;
  assign \new_[45397]_  = \new_[45396]_  & \new_[45393]_ ;
  assign \new_[45400]_  = A233 & ~A232;
  assign \new_[45403]_  = ~A236 & A234;
  assign \new_[45404]_  = \new_[45403]_  & \new_[45400]_ ;
  assign \new_[45405]_  = \new_[45404]_  & \new_[45397]_ ;
  assign \new_[45408]_  = ~A268 & A267;
  assign \new_[45411]_  = ~A298 & A269;
  assign \new_[45412]_  = \new_[45411]_  & \new_[45408]_ ;
  assign \new_[45415]_  = ~A300 & A299;
  assign \new_[45418]_  = A302 & ~A301;
  assign \new_[45419]_  = \new_[45418]_  & \new_[45415]_ ;
  assign \new_[45420]_  = \new_[45419]_  & \new_[45412]_ ;
  assign \new_[45423]_  = A200 & ~A199;
  assign \new_[45426]_  = A202 & A201;
  assign \new_[45427]_  = \new_[45426]_  & \new_[45423]_ ;
  assign \new_[45430]_  = A233 & ~A232;
  assign \new_[45433]_  = ~A235 & ~A234;
  assign \new_[45434]_  = \new_[45433]_  & \new_[45430]_ ;
  assign \new_[45435]_  = \new_[45434]_  & \new_[45427]_ ;
  assign \new_[45438]_  = A267 & A236;
  assign \new_[45441]_  = A269 & ~A268;
  assign \new_[45442]_  = \new_[45441]_  & \new_[45438]_ ;
  assign \new_[45445]_  = ~A299 & A298;
  assign \new_[45448]_  = A301 & A300;
  assign \new_[45449]_  = \new_[45448]_  & \new_[45445]_ ;
  assign \new_[45450]_  = \new_[45449]_  & \new_[45442]_ ;
  assign \new_[45453]_  = A200 & ~A199;
  assign \new_[45456]_  = A202 & A201;
  assign \new_[45457]_  = \new_[45456]_  & \new_[45453]_ ;
  assign \new_[45460]_  = A233 & ~A232;
  assign \new_[45463]_  = ~A235 & ~A234;
  assign \new_[45464]_  = \new_[45463]_  & \new_[45460]_ ;
  assign \new_[45465]_  = \new_[45464]_  & \new_[45457]_ ;
  assign \new_[45468]_  = A267 & A236;
  assign \new_[45471]_  = A269 & ~A268;
  assign \new_[45472]_  = \new_[45471]_  & \new_[45468]_ ;
  assign \new_[45475]_  = ~A299 & A298;
  assign \new_[45478]_  = ~A302 & A300;
  assign \new_[45479]_  = \new_[45478]_  & \new_[45475]_ ;
  assign \new_[45480]_  = \new_[45479]_  & \new_[45472]_ ;
  assign \new_[45483]_  = A200 & ~A199;
  assign \new_[45486]_  = A202 & A201;
  assign \new_[45487]_  = \new_[45486]_  & \new_[45483]_ ;
  assign \new_[45490]_  = A233 & ~A232;
  assign \new_[45493]_  = ~A235 & ~A234;
  assign \new_[45494]_  = \new_[45493]_  & \new_[45490]_ ;
  assign \new_[45495]_  = \new_[45494]_  & \new_[45487]_ ;
  assign \new_[45498]_  = A267 & A236;
  assign \new_[45501]_  = A269 & ~A268;
  assign \new_[45502]_  = \new_[45501]_  & \new_[45498]_ ;
  assign \new_[45505]_  = A299 & ~A298;
  assign \new_[45508]_  = A301 & A300;
  assign \new_[45509]_  = \new_[45508]_  & \new_[45505]_ ;
  assign \new_[45510]_  = \new_[45509]_  & \new_[45502]_ ;
  assign \new_[45513]_  = A200 & ~A199;
  assign \new_[45516]_  = A202 & A201;
  assign \new_[45517]_  = \new_[45516]_  & \new_[45513]_ ;
  assign \new_[45520]_  = A233 & ~A232;
  assign \new_[45523]_  = ~A235 & ~A234;
  assign \new_[45524]_  = \new_[45523]_  & \new_[45520]_ ;
  assign \new_[45525]_  = \new_[45524]_  & \new_[45517]_ ;
  assign \new_[45528]_  = A267 & A236;
  assign \new_[45531]_  = A269 & ~A268;
  assign \new_[45532]_  = \new_[45531]_  & \new_[45528]_ ;
  assign \new_[45535]_  = A299 & ~A298;
  assign \new_[45538]_  = ~A302 & A300;
  assign \new_[45539]_  = \new_[45538]_  & \new_[45535]_ ;
  assign \new_[45540]_  = \new_[45539]_  & \new_[45532]_ ;
  assign \new_[45543]_  = A200 & ~A199;
  assign \new_[45546]_  = A202 & A201;
  assign \new_[45547]_  = \new_[45546]_  & \new_[45543]_ ;
  assign \new_[45550]_  = A233 & ~A232;
  assign \new_[45553]_  = ~A235 & ~A234;
  assign \new_[45554]_  = \new_[45553]_  & \new_[45550]_ ;
  assign \new_[45555]_  = \new_[45554]_  & \new_[45547]_ ;
  assign \new_[45558]_  = ~A267 & A236;
  assign \new_[45561]_  = A298 & A268;
  assign \new_[45562]_  = \new_[45561]_  & \new_[45558]_ ;
  assign \new_[45565]_  = ~A300 & ~A299;
  assign \new_[45568]_  = A302 & ~A301;
  assign \new_[45569]_  = \new_[45568]_  & \new_[45565]_ ;
  assign \new_[45570]_  = \new_[45569]_  & \new_[45562]_ ;
  assign \new_[45573]_  = A200 & ~A199;
  assign \new_[45576]_  = A202 & A201;
  assign \new_[45577]_  = \new_[45576]_  & \new_[45573]_ ;
  assign \new_[45580]_  = A233 & ~A232;
  assign \new_[45583]_  = ~A235 & ~A234;
  assign \new_[45584]_  = \new_[45583]_  & \new_[45580]_ ;
  assign \new_[45585]_  = \new_[45584]_  & \new_[45577]_ ;
  assign \new_[45588]_  = ~A267 & A236;
  assign \new_[45591]_  = ~A298 & A268;
  assign \new_[45592]_  = \new_[45591]_  & \new_[45588]_ ;
  assign \new_[45595]_  = ~A300 & A299;
  assign \new_[45598]_  = A302 & ~A301;
  assign \new_[45599]_  = \new_[45598]_  & \new_[45595]_ ;
  assign \new_[45600]_  = \new_[45599]_  & \new_[45592]_ ;
  assign \new_[45603]_  = A200 & ~A199;
  assign \new_[45606]_  = A202 & A201;
  assign \new_[45607]_  = \new_[45606]_  & \new_[45603]_ ;
  assign \new_[45610]_  = A233 & ~A232;
  assign \new_[45613]_  = ~A235 & ~A234;
  assign \new_[45614]_  = \new_[45613]_  & \new_[45610]_ ;
  assign \new_[45615]_  = \new_[45614]_  & \new_[45607]_ ;
  assign \new_[45618]_  = ~A267 & A236;
  assign \new_[45621]_  = A298 & ~A269;
  assign \new_[45622]_  = \new_[45621]_  & \new_[45618]_ ;
  assign \new_[45625]_  = ~A300 & ~A299;
  assign \new_[45628]_  = A302 & ~A301;
  assign \new_[45629]_  = \new_[45628]_  & \new_[45625]_ ;
  assign \new_[45630]_  = \new_[45629]_  & \new_[45622]_ ;
  assign \new_[45633]_  = A200 & ~A199;
  assign \new_[45636]_  = A202 & A201;
  assign \new_[45637]_  = \new_[45636]_  & \new_[45633]_ ;
  assign \new_[45640]_  = A233 & ~A232;
  assign \new_[45643]_  = ~A235 & ~A234;
  assign \new_[45644]_  = \new_[45643]_  & \new_[45640]_ ;
  assign \new_[45645]_  = \new_[45644]_  & \new_[45637]_ ;
  assign \new_[45648]_  = ~A267 & A236;
  assign \new_[45651]_  = ~A298 & ~A269;
  assign \new_[45652]_  = \new_[45651]_  & \new_[45648]_ ;
  assign \new_[45655]_  = ~A300 & A299;
  assign \new_[45658]_  = A302 & ~A301;
  assign \new_[45659]_  = \new_[45658]_  & \new_[45655]_ ;
  assign \new_[45660]_  = \new_[45659]_  & \new_[45652]_ ;
  assign \new_[45663]_  = A200 & ~A199;
  assign \new_[45666]_  = A202 & A201;
  assign \new_[45667]_  = \new_[45666]_  & \new_[45663]_ ;
  assign \new_[45670]_  = A233 & ~A232;
  assign \new_[45673]_  = ~A235 & ~A234;
  assign \new_[45674]_  = \new_[45673]_  & \new_[45670]_ ;
  assign \new_[45675]_  = \new_[45674]_  & \new_[45667]_ ;
  assign \new_[45678]_  = A265 & A236;
  assign \new_[45681]_  = A298 & A266;
  assign \new_[45682]_  = \new_[45681]_  & \new_[45678]_ ;
  assign \new_[45685]_  = ~A300 & ~A299;
  assign \new_[45688]_  = A302 & ~A301;
  assign \new_[45689]_  = \new_[45688]_  & \new_[45685]_ ;
  assign \new_[45690]_  = \new_[45689]_  & \new_[45682]_ ;
  assign \new_[45693]_  = A200 & ~A199;
  assign \new_[45696]_  = A202 & A201;
  assign \new_[45697]_  = \new_[45696]_  & \new_[45693]_ ;
  assign \new_[45700]_  = A233 & ~A232;
  assign \new_[45703]_  = ~A235 & ~A234;
  assign \new_[45704]_  = \new_[45703]_  & \new_[45700]_ ;
  assign \new_[45705]_  = \new_[45704]_  & \new_[45697]_ ;
  assign \new_[45708]_  = A265 & A236;
  assign \new_[45711]_  = ~A298 & A266;
  assign \new_[45712]_  = \new_[45711]_  & \new_[45708]_ ;
  assign \new_[45715]_  = ~A300 & A299;
  assign \new_[45718]_  = A302 & ~A301;
  assign \new_[45719]_  = \new_[45718]_  & \new_[45715]_ ;
  assign \new_[45720]_  = \new_[45719]_  & \new_[45712]_ ;
  assign \new_[45723]_  = A200 & ~A199;
  assign \new_[45726]_  = A202 & A201;
  assign \new_[45727]_  = \new_[45726]_  & \new_[45723]_ ;
  assign \new_[45730]_  = A233 & ~A232;
  assign \new_[45733]_  = ~A235 & ~A234;
  assign \new_[45734]_  = \new_[45733]_  & \new_[45730]_ ;
  assign \new_[45735]_  = \new_[45734]_  & \new_[45727]_ ;
  assign \new_[45738]_  = ~A265 & A236;
  assign \new_[45741]_  = A298 & ~A266;
  assign \new_[45742]_  = \new_[45741]_  & \new_[45738]_ ;
  assign \new_[45745]_  = ~A300 & ~A299;
  assign \new_[45748]_  = A302 & ~A301;
  assign \new_[45749]_  = \new_[45748]_  & \new_[45745]_ ;
  assign \new_[45750]_  = \new_[45749]_  & \new_[45742]_ ;
  assign \new_[45753]_  = A200 & ~A199;
  assign \new_[45756]_  = A202 & A201;
  assign \new_[45757]_  = \new_[45756]_  & \new_[45753]_ ;
  assign \new_[45760]_  = A233 & ~A232;
  assign \new_[45763]_  = ~A235 & ~A234;
  assign \new_[45764]_  = \new_[45763]_  & \new_[45760]_ ;
  assign \new_[45765]_  = \new_[45764]_  & \new_[45757]_ ;
  assign \new_[45768]_  = ~A265 & A236;
  assign \new_[45771]_  = ~A298 & ~A266;
  assign \new_[45772]_  = \new_[45771]_  & \new_[45768]_ ;
  assign \new_[45775]_  = ~A300 & A299;
  assign \new_[45778]_  = A302 & ~A301;
  assign \new_[45779]_  = \new_[45778]_  & \new_[45775]_ ;
  assign \new_[45780]_  = \new_[45779]_  & \new_[45772]_ ;
  assign \new_[45783]_  = A200 & ~A199;
  assign \new_[45786]_  = A202 & A201;
  assign \new_[45787]_  = \new_[45786]_  & \new_[45783]_ ;
  assign \new_[45790]_  = ~A233 & A232;
  assign \new_[45793]_  = A235 & A234;
  assign \new_[45794]_  = \new_[45793]_  & \new_[45790]_ ;
  assign \new_[45795]_  = \new_[45794]_  & \new_[45787]_ ;
  assign \new_[45798]_  = ~A268 & A267;
  assign \new_[45801]_  = A298 & A269;
  assign \new_[45802]_  = \new_[45801]_  & \new_[45798]_ ;
  assign \new_[45805]_  = ~A300 & ~A299;
  assign \new_[45808]_  = A302 & ~A301;
  assign \new_[45809]_  = \new_[45808]_  & \new_[45805]_ ;
  assign \new_[45810]_  = \new_[45809]_  & \new_[45802]_ ;
  assign \new_[45813]_  = A200 & ~A199;
  assign \new_[45816]_  = A202 & A201;
  assign \new_[45817]_  = \new_[45816]_  & \new_[45813]_ ;
  assign \new_[45820]_  = ~A233 & A232;
  assign \new_[45823]_  = A235 & A234;
  assign \new_[45824]_  = \new_[45823]_  & \new_[45820]_ ;
  assign \new_[45825]_  = \new_[45824]_  & \new_[45817]_ ;
  assign \new_[45828]_  = ~A268 & A267;
  assign \new_[45831]_  = ~A298 & A269;
  assign \new_[45832]_  = \new_[45831]_  & \new_[45828]_ ;
  assign \new_[45835]_  = ~A300 & A299;
  assign \new_[45838]_  = A302 & ~A301;
  assign \new_[45839]_  = \new_[45838]_  & \new_[45835]_ ;
  assign \new_[45840]_  = \new_[45839]_  & \new_[45832]_ ;
  assign \new_[45843]_  = A200 & ~A199;
  assign \new_[45846]_  = A202 & A201;
  assign \new_[45847]_  = \new_[45846]_  & \new_[45843]_ ;
  assign \new_[45850]_  = ~A233 & A232;
  assign \new_[45853]_  = ~A236 & A234;
  assign \new_[45854]_  = \new_[45853]_  & \new_[45850]_ ;
  assign \new_[45855]_  = \new_[45854]_  & \new_[45847]_ ;
  assign \new_[45858]_  = ~A268 & A267;
  assign \new_[45861]_  = A298 & A269;
  assign \new_[45862]_  = \new_[45861]_  & \new_[45858]_ ;
  assign \new_[45865]_  = ~A300 & ~A299;
  assign \new_[45868]_  = A302 & ~A301;
  assign \new_[45869]_  = \new_[45868]_  & \new_[45865]_ ;
  assign \new_[45870]_  = \new_[45869]_  & \new_[45862]_ ;
  assign \new_[45873]_  = A200 & ~A199;
  assign \new_[45876]_  = A202 & A201;
  assign \new_[45877]_  = \new_[45876]_  & \new_[45873]_ ;
  assign \new_[45880]_  = ~A233 & A232;
  assign \new_[45883]_  = ~A236 & A234;
  assign \new_[45884]_  = \new_[45883]_  & \new_[45880]_ ;
  assign \new_[45885]_  = \new_[45884]_  & \new_[45877]_ ;
  assign \new_[45888]_  = ~A268 & A267;
  assign \new_[45891]_  = ~A298 & A269;
  assign \new_[45892]_  = \new_[45891]_  & \new_[45888]_ ;
  assign \new_[45895]_  = ~A300 & A299;
  assign \new_[45898]_  = A302 & ~A301;
  assign \new_[45899]_  = \new_[45898]_  & \new_[45895]_ ;
  assign \new_[45900]_  = \new_[45899]_  & \new_[45892]_ ;
  assign \new_[45903]_  = A200 & ~A199;
  assign \new_[45906]_  = A202 & A201;
  assign \new_[45907]_  = \new_[45906]_  & \new_[45903]_ ;
  assign \new_[45910]_  = ~A233 & A232;
  assign \new_[45913]_  = ~A235 & ~A234;
  assign \new_[45914]_  = \new_[45913]_  & \new_[45910]_ ;
  assign \new_[45915]_  = \new_[45914]_  & \new_[45907]_ ;
  assign \new_[45918]_  = A267 & A236;
  assign \new_[45921]_  = A269 & ~A268;
  assign \new_[45922]_  = \new_[45921]_  & \new_[45918]_ ;
  assign \new_[45925]_  = ~A299 & A298;
  assign \new_[45928]_  = A301 & A300;
  assign \new_[45929]_  = \new_[45928]_  & \new_[45925]_ ;
  assign \new_[45930]_  = \new_[45929]_  & \new_[45922]_ ;
  assign \new_[45933]_  = A200 & ~A199;
  assign \new_[45936]_  = A202 & A201;
  assign \new_[45937]_  = \new_[45936]_  & \new_[45933]_ ;
  assign \new_[45940]_  = ~A233 & A232;
  assign \new_[45943]_  = ~A235 & ~A234;
  assign \new_[45944]_  = \new_[45943]_  & \new_[45940]_ ;
  assign \new_[45945]_  = \new_[45944]_  & \new_[45937]_ ;
  assign \new_[45948]_  = A267 & A236;
  assign \new_[45951]_  = A269 & ~A268;
  assign \new_[45952]_  = \new_[45951]_  & \new_[45948]_ ;
  assign \new_[45955]_  = ~A299 & A298;
  assign \new_[45958]_  = ~A302 & A300;
  assign \new_[45959]_  = \new_[45958]_  & \new_[45955]_ ;
  assign \new_[45960]_  = \new_[45959]_  & \new_[45952]_ ;
  assign \new_[45963]_  = A200 & ~A199;
  assign \new_[45966]_  = A202 & A201;
  assign \new_[45967]_  = \new_[45966]_  & \new_[45963]_ ;
  assign \new_[45970]_  = ~A233 & A232;
  assign \new_[45973]_  = ~A235 & ~A234;
  assign \new_[45974]_  = \new_[45973]_  & \new_[45970]_ ;
  assign \new_[45975]_  = \new_[45974]_  & \new_[45967]_ ;
  assign \new_[45978]_  = A267 & A236;
  assign \new_[45981]_  = A269 & ~A268;
  assign \new_[45982]_  = \new_[45981]_  & \new_[45978]_ ;
  assign \new_[45985]_  = A299 & ~A298;
  assign \new_[45988]_  = A301 & A300;
  assign \new_[45989]_  = \new_[45988]_  & \new_[45985]_ ;
  assign \new_[45990]_  = \new_[45989]_  & \new_[45982]_ ;
  assign \new_[45993]_  = A200 & ~A199;
  assign \new_[45996]_  = A202 & A201;
  assign \new_[45997]_  = \new_[45996]_  & \new_[45993]_ ;
  assign \new_[46000]_  = ~A233 & A232;
  assign \new_[46003]_  = ~A235 & ~A234;
  assign \new_[46004]_  = \new_[46003]_  & \new_[46000]_ ;
  assign \new_[46005]_  = \new_[46004]_  & \new_[45997]_ ;
  assign \new_[46008]_  = A267 & A236;
  assign \new_[46011]_  = A269 & ~A268;
  assign \new_[46012]_  = \new_[46011]_  & \new_[46008]_ ;
  assign \new_[46015]_  = A299 & ~A298;
  assign \new_[46018]_  = ~A302 & A300;
  assign \new_[46019]_  = \new_[46018]_  & \new_[46015]_ ;
  assign \new_[46020]_  = \new_[46019]_  & \new_[46012]_ ;
  assign \new_[46023]_  = A200 & ~A199;
  assign \new_[46026]_  = A202 & A201;
  assign \new_[46027]_  = \new_[46026]_  & \new_[46023]_ ;
  assign \new_[46030]_  = ~A233 & A232;
  assign \new_[46033]_  = ~A235 & ~A234;
  assign \new_[46034]_  = \new_[46033]_  & \new_[46030]_ ;
  assign \new_[46035]_  = \new_[46034]_  & \new_[46027]_ ;
  assign \new_[46038]_  = ~A267 & A236;
  assign \new_[46041]_  = A298 & A268;
  assign \new_[46042]_  = \new_[46041]_  & \new_[46038]_ ;
  assign \new_[46045]_  = ~A300 & ~A299;
  assign \new_[46048]_  = A302 & ~A301;
  assign \new_[46049]_  = \new_[46048]_  & \new_[46045]_ ;
  assign \new_[46050]_  = \new_[46049]_  & \new_[46042]_ ;
  assign \new_[46053]_  = A200 & ~A199;
  assign \new_[46056]_  = A202 & A201;
  assign \new_[46057]_  = \new_[46056]_  & \new_[46053]_ ;
  assign \new_[46060]_  = ~A233 & A232;
  assign \new_[46063]_  = ~A235 & ~A234;
  assign \new_[46064]_  = \new_[46063]_  & \new_[46060]_ ;
  assign \new_[46065]_  = \new_[46064]_  & \new_[46057]_ ;
  assign \new_[46068]_  = ~A267 & A236;
  assign \new_[46071]_  = ~A298 & A268;
  assign \new_[46072]_  = \new_[46071]_  & \new_[46068]_ ;
  assign \new_[46075]_  = ~A300 & A299;
  assign \new_[46078]_  = A302 & ~A301;
  assign \new_[46079]_  = \new_[46078]_  & \new_[46075]_ ;
  assign \new_[46080]_  = \new_[46079]_  & \new_[46072]_ ;
  assign \new_[46083]_  = A200 & ~A199;
  assign \new_[46086]_  = A202 & A201;
  assign \new_[46087]_  = \new_[46086]_  & \new_[46083]_ ;
  assign \new_[46090]_  = ~A233 & A232;
  assign \new_[46093]_  = ~A235 & ~A234;
  assign \new_[46094]_  = \new_[46093]_  & \new_[46090]_ ;
  assign \new_[46095]_  = \new_[46094]_  & \new_[46087]_ ;
  assign \new_[46098]_  = ~A267 & A236;
  assign \new_[46101]_  = A298 & ~A269;
  assign \new_[46102]_  = \new_[46101]_  & \new_[46098]_ ;
  assign \new_[46105]_  = ~A300 & ~A299;
  assign \new_[46108]_  = A302 & ~A301;
  assign \new_[46109]_  = \new_[46108]_  & \new_[46105]_ ;
  assign \new_[46110]_  = \new_[46109]_  & \new_[46102]_ ;
  assign \new_[46113]_  = A200 & ~A199;
  assign \new_[46116]_  = A202 & A201;
  assign \new_[46117]_  = \new_[46116]_  & \new_[46113]_ ;
  assign \new_[46120]_  = ~A233 & A232;
  assign \new_[46123]_  = ~A235 & ~A234;
  assign \new_[46124]_  = \new_[46123]_  & \new_[46120]_ ;
  assign \new_[46125]_  = \new_[46124]_  & \new_[46117]_ ;
  assign \new_[46128]_  = ~A267 & A236;
  assign \new_[46131]_  = ~A298 & ~A269;
  assign \new_[46132]_  = \new_[46131]_  & \new_[46128]_ ;
  assign \new_[46135]_  = ~A300 & A299;
  assign \new_[46138]_  = A302 & ~A301;
  assign \new_[46139]_  = \new_[46138]_  & \new_[46135]_ ;
  assign \new_[46140]_  = \new_[46139]_  & \new_[46132]_ ;
  assign \new_[46143]_  = A200 & ~A199;
  assign \new_[46146]_  = A202 & A201;
  assign \new_[46147]_  = \new_[46146]_  & \new_[46143]_ ;
  assign \new_[46150]_  = ~A233 & A232;
  assign \new_[46153]_  = ~A235 & ~A234;
  assign \new_[46154]_  = \new_[46153]_  & \new_[46150]_ ;
  assign \new_[46155]_  = \new_[46154]_  & \new_[46147]_ ;
  assign \new_[46158]_  = A265 & A236;
  assign \new_[46161]_  = A298 & A266;
  assign \new_[46162]_  = \new_[46161]_  & \new_[46158]_ ;
  assign \new_[46165]_  = ~A300 & ~A299;
  assign \new_[46168]_  = A302 & ~A301;
  assign \new_[46169]_  = \new_[46168]_  & \new_[46165]_ ;
  assign \new_[46170]_  = \new_[46169]_  & \new_[46162]_ ;
  assign \new_[46173]_  = A200 & ~A199;
  assign \new_[46176]_  = A202 & A201;
  assign \new_[46177]_  = \new_[46176]_  & \new_[46173]_ ;
  assign \new_[46180]_  = ~A233 & A232;
  assign \new_[46183]_  = ~A235 & ~A234;
  assign \new_[46184]_  = \new_[46183]_  & \new_[46180]_ ;
  assign \new_[46185]_  = \new_[46184]_  & \new_[46177]_ ;
  assign \new_[46188]_  = A265 & A236;
  assign \new_[46191]_  = ~A298 & A266;
  assign \new_[46192]_  = \new_[46191]_  & \new_[46188]_ ;
  assign \new_[46195]_  = ~A300 & A299;
  assign \new_[46198]_  = A302 & ~A301;
  assign \new_[46199]_  = \new_[46198]_  & \new_[46195]_ ;
  assign \new_[46200]_  = \new_[46199]_  & \new_[46192]_ ;
  assign \new_[46203]_  = A200 & ~A199;
  assign \new_[46206]_  = A202 & A201;
  assign \new_[46207]_  = \new_[46206]_  & \new_[46203]_ ;
  assign \new_[46210]_  = ~A233 & A232;
  assign \new_[46213]_  = ~A235 & ~A234;
  assign \new_[46214]_  = \new_[46213]_  & \new_[46210]_ ;
  assign \new_[46215]_  = \new_[46214]_  & \new_[46207]_ ;
  assign \new_[46218]_  = ~A265 & A236;
  assign \new_[46221]_  = A298 & ~A266;
  assign \new_[46222]_  = \new_[46221]_  & \new_[46218]_ ;
  assign \new_[46225]_  = ~A300 & ~A299;
  assign \new_[46228]_  = A302 & ~A301;
  assign \new_[46229]_  = \new_[46228]_  & \new_[46225]_ ;
  assign \new_[46230]_  = \new_[46229]_  & \new_[46222]_ ;
  assign \new_[46233]_  = A200 & ~A199;
  assign \new_[46236]_  = A202 & A201;
  assign \new_[46237]_  = \new_[46236]_  & \new_[46233]_ ;
  assign \new_[46240]_  = ~A233 & A232;
  assign \new_[46243]_  = ~A235 & ~A234;
  assign \new_[46244]_  = \new_[46243]_  & \new_[46240]_ ;
  assign \new_[46245]_  = \new_[46244]_  & \new_[46237]_ ;
  assign \new_[46248]_  = ~A265 & A236;
  assign \new_[46251]_  = ~A298 & ~A266;
  assign \new_[46252]_  = \new_[46251]_  & \new_[46248]_ ;
  assign \new_[46255]_  = ~A300 & A299;
  assign \new_[46258]_  = A302 & ~A301;
  assign \new_[46259]_  = \new_[46258]_  & \new_[46255]_ ;
  assign \new_[46260]_  = \new_[46259]_  & \new_[46252]_ ;
  assign \new_[46263]_  = A200 & ~A199;
  assign \new_[46266]_  = ~A203 & A201;
  assign \new_[46267]_  = \new_[46266]_  & \new_[46263]_ ;
  assign \new_[46270]_  = A233 & ~A232;
  assign \new_[46273]_  = A235 & A234;
  assign \new_[46274]_  = \new_[46273]_  & \new_[46270]_ ;
  assign \new_[46275]_  = \new_[46274]_  & \new_[46267]_ ;
  assign \new_[46278]_  = ~A268 & A267;
  assign \new_[46281]_  = A298 & A269;
  assign \new_[46282]_  = \new_[46281]_  & \new_[46278]_ ;
  assign \new_[46285]_  = ~A300 & ~A299;
  assign \new_[46288]_  = A302 & ~A301;
  assign \new_[46289]_  = \new_[46288]_  & \new_[46285]_ ;
  assign \new_[46290]_  = \new_[46289]_  & \new_[46282]_ ;
  assign \new_[46293]_  = A200 & ~A199;
  assign \new_[46296]_  = ~A203 & A201;
  assign \new_[46297]_  = \new_[46296]_  & \new_[46293]_ ;
  assign \new_[46300]_  = A233 & ~A232;
  assign \new_[46303]_  = A235 & A234;
  assign \new_[46304]_  = \new_[46303]_  & \new_[46300]_ ;
  assign \new_[46305]_  = \new_[46304]_  & \new_[46297]_ ;
  assign \new_[46308]_  = ~A268 & A267;
  assign \new_[46311]_  = ~A298 & A269;
  assign \new_[46312]_  = \new_[46311]_  & \new_[46308]_ ;
  assign \new_[46315]_  = ~A300 & A299;
  assign \new_[46318]_  = A302 & ~A301;
  assign \new_[46319]_  = \new_[46318]_  & \new_[46315]_ ;
  assign \new_[46320]_  = \new_[46319]_  & \new_[46312]_ ;
  assign \new_[46323]_  = A200 & ~A199;
  assign \new_[46326]_  = ~A203 & A201;
  assign \new_[46327]_  = \new_[46326]_  & \new_[46323]_ ;
  assign \new_[46330]_  = A233 & ~A232;
  assign \new_[46333]_  = ~A236 & A234;
  assign \new_[46334]_  = \new_[46333]_  & \new_[46330]_ ;
  assign \new_[46335]_  = \new_[46334]_  & \new_[46327]_ ;
  assign \new_[46338]_  = ~A268 & A267;
  assign \new_[46341]_  = A298 & A269;
  assign \new_[46342]_  = \new_[46341]_  & \new_[46338]_ ;
  assign \new_[46345]_  = ~A300 & ~A299;
  assign \new_[46348]_  = A302 & ~A301;
  assign \new_[46349]_  = \new_[46348]_  & \new_[46345]_ ;
  assign \new_[46350]_  = \new_[46349]_  & \new_[46342]_ ;
  assign \new_[46353]_  = A200 & ~A199;
  assign \new_[46356]_  = ~A203 & A201;
  assign \new_[46357]_  = \new_[46356]_  & \new_[46353]_ ;
  assign \new_[46360]_  = A233 & ~A232;
  assign \new_[46363]_  = ~A236 & A234;
  assign \new_[46364]_  = \new_[46363]_  & \new_[46360]_ ;
  assign \new_[46365]_  = \new_[46364]_  & \new_[46357]_ ;
  assign \new_[46368]_  = ~A268 & A267;
  assign \new_[46371]_  = ~A298 & A269;
  assign \new_[46372]_  = \new_[46371]_  & \new_[46368]_ ;
  assign \new_[46375]_  = ~A300 & A299;
  assign \new_[46378]_  = A302 & ~A301;
  assign \new_[46379]_  = \new_[46378]_  & \new_[46375]_ ;
  assign \new_[46380]_  = \new_[46379]_  & \new_[46372]_ ;
  assign \new_[46383]_  = A200 & ~A199;
  assign \new_[46386]_  = ~A203 & A201;
  assign \new_[46387]_  = \new_[46386]_  & \new_[46383]_ ;
  assign \new_[46390]_  = A233 & ~A232;
  assign \new_[46393]_  = ~A235 & ~A234;
  assign \new_[46394]_  = \new_[46393]_  & \new_[46390]_ ;
  assign \new_[46395]_  = \new_[46394]_  & \new_[46387]_ ;
  assign \new_[46398]_  = A267 & A236;
  assign \new_[46401]_  = A269 & ~A268;
  assign \new_[46402]_  = \new_[46401]_  & \new_[46398]_ ;
  assign \new_[46405]_  = ~A299 & A298;
  assign \new_[46408]_  = A301 & A300;
  assign \new_[46409]_  = \new_[46408]_  & \new_[46405]_ ;
  assign \new_[46410]_  = \new_[46409]_  & \new_[46402]_ ;
  assign \new_[46413]_  = A200 & ~A199;
  assign \new_[46416]_  = ~A203 & A201;
  assign \new_[46417]_  = \new_[46416]_  & \new_[46413]_ ;
  assign \new_[46420]_  = A233 & ~A232;
  assign \new_[46423]_  = ~A235 & ~A234;
  assign \new_[46424]_  = \new_[46423]_  & \new_[46420]_ ;
  assign \new_[46425]_  = \new_[46424]_  & \new_[46417]_ ;
  assign \new_[46428]_  = A267 & A236;
  assign \new_[46431]_  = A269 & ~A268;
  assign \new_[46432]_  = \new_[46431]_  & \new_[46428]_ ;
  assign \new_[46435]_  = ~A299 & A298;
  assign \new_[46438]_  = ~A302 & A300;
  assign \new_[46439]_  = \new_[46438]_  & \new_[46435]_ ;
  assign \new_[46440]_  = \new_[46439]_  & \new_[46432]_ ;
  assign \new_[46443]_  = A200 & ~A199;
  assign \new_[46446]_  = ~A203 & A201;
  assign \new_[46447]_  = \new_[46446]_  & \new_[46443]_ ;
  assign \new_[46450]_  = A233 & ~A232;
  assign \new_[46453]_  = ~A235 & ~A234;
  assign \new_[46454]_  = \new_[46453]_  & \new_[46450]_ ;
  assign \new_[46455]_  = \new_[46454]_  & \new_[46447]_ ;
  assign \new_[46458]_  = A267 & A236;
  assign \new_[46461]_  = A269 & ~A268;
  assign \new_[46462]_  = \new_[46461]_  & \new_[46458]_ ;
  assign \new_[46465]_  = A299 & ~A298;
  assign \new_[46468]_  = A301 & A300;
  assign \new_[46469]_  = \new_[46468]_  & \new_[46465]_ ;
  assign \new_[46470]_  = \new_[46469]_  & \new_[46462]_ ;
  assign \new_[46473]_  = A200 & ~A199;
  assign \new_[46476]_  = ~A203 & A201;
  assign \new_[46477]_  = \new_[46476]_  & \new_[46473]_ ;
  assign \new_[46480]_  = A233 & ~A232;
  assign \new_[46483]_  = ~A235 & ~A234;
  assign \new_[46484]_  = \new_[46483]_  & \new_[46480]_ ;
  assign \new_[46485]_  = \new_[46484]_  & \new_[46477]_ ;
  assign \new_[46488]_  = A267 & A236;
  assign \new_[46491]_  = A269 & ~A268;
  assign \new_[46492]_  = \new_[46491]_  & \new_[46488]_ ;
  assign \new_[46495]_  = A299 & ~A298;
  assign \new_[46498]_  = ~A302 & A300;
  assign \new_[46499]_  = \new_[46498]_  & \new_[46495]_ ;
  assign \new_[46500]_  = \new_[46499]_  & \new_[46492]_ ;
  assign \new_[46503]_  = A200 & ~A199;
  assign \new_[46506]_  = ~A203 & A201;
  assign \new_[46507]_  = \new_[46506]_  & \new_[46503]_ ;
  assign \new_[46510]_  = A233 & ~A232;
  assign \new_[46513]_  = ~A235 & ~A234;
  assign \new_[46514]_  = \new_[46513]_  & \new_[46510]_ ;
  assign \new_[46515]_  = \new_[46514]_  & \new_[46507]_ ;
  assign \new_[46518]_  = ~A267 & A236;
  assign \new_[46521]_  = A298 & A268;
  assign \new_[46522]_  = \new_[46521]_  & \new_[46518]_ ;
  assign \new_[46525]_  = ~A300 & ~A299;
  assign \new_[46528]_  = A302 & ~A301;
  assign \new_[46529]_  = \new_[46528]_  & \new_[46525]_ ;
  assign \new_[46530]_  = \new_[46529]_  & \new_[46522]_ ;
  assign \new_[46533]_  = A200 & ~A199;
  assign \new_[46536]_  = ~A203 & A201;
  assign \new_[46537]_  = \new_[46536]_  & \new_[46533]_ ;
  assign \new_[46540]_  = A233 & ~A232;
  assign \new_[46543]_  = ~A235 & ~A234;
  assign \new_[46544]_  = \new_[46543]_  & \new_[46540]_ ;
  assign \new_[46545]_  = \new_[46544]_  & \new_[46537]_ ;
  assign \new_[46548]_  = ~A267 & A236;
  assign \new_[46551]_  = ~A298 & A268;
  assign \new_[46552]_  = \new_[46551]_  & \new_[46548]_ ;
  assign \new_[46555]_  = ~A300 & A299;
  assign \new_[46558]_  = A302 & ~A301;
  assign \new_[46559]_  = \new_[46558]_  & \new_[46555]_ ;
  assign \new_[46560]_  = \new_[46559]_  & \new_[46552]_ ;
  assign \new_[46563]_  = A200 & ~A199;
  assign \new_[46566]_  = ~A203 & A201;
  assign \new_[46567]_  = \new_[46566]_  & \new_[46563]_ ;
  assign \new_[46570]_  = A233 & ~A232;
  assign \new_[46573]_  = ~A235 & ~A234;
  assign \new_[46574]_  = \new_[46573]_  & \new_[46570]_ ;
  assign \new_[46575]_  = \new_[46574]_  & \new_[46567]_ ;
  assign \new_[46578]_  = ~A267 & A236;
  assign \new_[46581]_  = A298 & ~A269;
  assign \new_[46582]_  = \new_[46581]_  & \new_[46578]_ ;
  assign \new_[46585]_  = ~A300 & ~A299;
  assign \new_[46588]_  = A302 & ~A301;
  assign \new_[46589]_  = \new_[46588]_  & \new_[46585]_ ;
  assign \new_[46590]_  = \new_[46589]_  & \new_[46582]_ ;
  assign \new_[46593]_  = A200 & ~A199;
  assign \new_[46596]_  = ~A203 & A201;
  assign \new_[46597]_  = \new_[46596]_  & \new_[46593]_ ;
  assign \new_[46600]_  = A233 & ~A232;
  assign \new_[46603]_  = ~A235 & ~A234;
  assign \new_[46604]_  = \new_[46603]_  & \new_[46600]_ ;
  assign \new_[46605]_  = \new_[46604]_  & \new_[46597]_ ;
  assign \new_[46608]_  = ~A267 & A236;
  assign \new_[46611]_  = ~A298 & ~A269;
  assign \new_[46612]_  = \new_[46611]_  & \new_[46608]_ ;
  assign \new_[46615]_  = ~A300 & A299;
  assign \new_[46618]_  = A302 & ~A301;
  assign \new_[46619]_  = \new_[46618]_  & \new_[46615]_ ;
  assign \new_[46620]_  = \new_[46619]_  & \new_[46612]_ ;
  assign \new_[46623]_  = A200 & ~A199;
  assign \new_[46626]_  = ~A203 & A201;
  assign \new_[46627]_  = \new_[46626]_  & \new_[46623]_ ;
  assign \new_[46630]_  = A233 & ~A232;
  assign \new_[46633]_  = ~A235 & ~A234;
  assign \new_[46634]_  = \new_[46633]_  & \new_[46630]_ ;
  assign \new_[46635]_  = \new_[46634]_  & \new_[46627]_ ;
  assign \new_[46638]_  = A265 & A236;
  assign \new_[46641]_  = A298 & A266;
  assign \new_[46642]_  = \new_[46641]_  & \new_[46638]_ ;
  assign \new_[46645]_  = ~A300 & ~A299;
  assign \new_[46648]_  = A302 & ~A301;
  assign \new_[46649]_  = \new_[46648]_  & \new_[46645]_ ;
  assign \new_[46650]_  = \new_[46649]_  & \new_[46642]_ ;
  assign \new_[46653]_  = A200 & ~A199;
  assign \new_[46656]_  = ~A203 & A201;
  assign \new_[46657]_  = \new_[46656]_  & \new_[46653]_ ;
  assign \new_[46660]_  = A233 & ~A232;
  assign \new_[46663]_  = ~A235 & ~A234;
  assign \new_[46664]_  = \new_[46663]_  & \new_[46660]_ ;
  assign \new_[46665]_  = \new_[46664]_  & \new_[46657]_ ;
  assign \new_[46668]_  = A265 & A236;
  assign \new_[46671]_  = ~A298 & A266;
  assign \new_[46672]_  = \new_[46671]_  & \new_[46668]_ ;
  assign \new_[46675]_  = ~A300 & A299;
  assign \new_[46678]_  = A302 & ~A301;
  assign \new_[46679]_  = \new_[46678]_  & \new_[46675]_ ;
  assign \new_[46680]_  = \new_[46679]_  & \new_[46672]_ ;
  assign \new_[46683]_  = A200 & ~A199;
  assign \new_[46686]_  = ~A203 & A201;
  assign \new_[46687]_  = \new_[46686]_  & \new_[46683]_ ;
  assign \new_[46690]_  = A233 & ~A232;
  assign \new_[46693]_  = ~A235 & ~A234;
  assign \new_[46694]_  = \new_[46693]_  & \new_[46690]_ ;
  assign \new_[46695]_  = \new_[46694]_  & \new_[46687]_ ;
  assign \new_[46698]_  = ~A265 & A236;
  assign \new_[46701]_  = A298 & ~A266;
  assign \new_[46702]_  = \new_[46701]_  & \new_[46698]_ ;
  assign \new_[46705]_  = ~A300 & ~A299;
  assign \new_[46708]_  = A302 & ~A301;
  assign \new_[46709]_  = \new_[46708]_  & \new_[46705]_ ;
  assign \new_[46710]_  = \new_[46709]_  & \new_[46702]_ ;
  assign \new_[46713]_  = A200 & ~A199;
  assign \new_[46716]_  = ~A203 & A201;
  assign \new_[46717]_  = \new_[46716]_  & \new_[46713]_ ;
  assign \new_[46720]_  = A233 & ~A232;
  assign \new_[46723]_  = ~A235 & ~A234;
  assign \new_[46724]_  = \new_[46723]_  & \new_[46720]_ ;
  assign \new_[46725]_  = \new_[46724]_  & \new_[46717]_ ;
  assign \new_[46728]_  = ~A265 & A236;
  assign \new_[46731]_  = ~A298 & ~A266;
  assign \new_[46732]_  = \new_[46731]_  & \new_[46728]_ ;
  assign \new_[46735]_  = ~A300 & A299;
  assign \new_[46738]_  = A302 & ~A301;
  assign \new_[46739]_  = \new_[46738]_  & \new_[46735]_ ;
  assign \new_[46740]_  = \new_[46739]_  & \new_[46732]_ ;
  assign \new_[46743]_  = A200 & ~A199;
  assign \new_[46746]_  = ~A203 & A201;
  assign \new_[46747]_  = \new_[46746]_  & \new_[46743]_ ;
  assign \new_[46750]_  = ~A233 & A232;
  assign \new_[46753]_  = A235 & A234;
  assign \new_[46754]_  = \new_[46753]_  & \new_[46750]_ ;
  assign \new_[46755]_  = \new_[46754]_  & \new_[46747]_ ;
  assign \new_[46758]_  = ~A268 & A267;
  assign \new_[46761]_  = A298 & A269;
  assign \new_[46762]_  = \new_[46761]_  & \new_[46758]_ ;
  assign \new_[46765]_  = ~A300 & ~A299;
  assign \new_[46768]_  = A302 & ~A301;
  assign \new_[46769]_  = \new_[46768]_  & \new_[46765]_ ;
  assign \new_[46770]_  = \new_[46769]_  & \new_[46762]_ ;
  assign \new_[46773]_  = A200 & ~A199;
  assign \new_[46776]_  = ~A203 & A201;
  assign \new_[46777]_  = \new_[46776]_  & \new_[46773]_ ;
  assign \new_[46780]_  = ~A233 & A232;
  assign \new_[46783]_  = A235 & A234;
  assign \new_[46784]_  = \new_[46783]_  & \new_[46780]_ ;
  assign \new_[46785]_  = \new_[46784]_  & \new_[46777]_ ;
  assign \new_[46788]_  = ~A268 & A267;
  assign \new_[46791]_  = ~A298 & A269;
  assign \new_[46792]_  = \new_[46791]_  & \new_[46788]_ ;
  assign \new_[46795]_  = ~A300 & A299;
  assign \new_[46798]_  = A302 & ~A301;
  assign \new_[46799]_  = \new_[46798]_  & \new_[46795]_ ;
  assign \new_[46800]_  = \new_[46799]_  & \new_[46792]_ ;
  assign \new_[46803]_  = A200 & ~A199;
  assign \new_[46806]_  = ~A203 & A201;
  assign \new_[46807]_  = \new_[46806]_  & \new_[46803]_ ;
  assign \new_[46810]_  = ~A233 & A232;
  assign \new_[46813]_  = ~A236 & A234;
  assign \new_[46814]_  = \new_[46813]_  & \new_[46810]_ ;
  assign \new_[46815]_  = \new_[46814]_  & \new_[46807]_ ;
  assign \new_[46818]_  = ~A268 & A267;
  assign \new_[46821]_  = A298 & A269;
  assign \new_[46822]_  = \new_[46821]_  & \new_[46818]_ ;
  assign \new_[46825]_  = ~A300 & ~A299;
  assign \new_[46828]_  = A302 & ~A301;
  assign \new_[46829]_  = \new_[46828]_  & \new_[46825]_ ;
  assign \new_[46830]_  = \new_[46829]_  & \new_[46822]_ ;
  assign \new_[46833]_  = A200 & ~A199;
  assign \new_[46836]_  = ~A203 & A201;
  assign \new_[46837]_  = \new_[46836]_  & \new_[46833]_ ;
  assign \new_[46840]_  = ~A233 & A232;
  assign \new_[46843]_  = ~A236 & A234;
  assign \new_[46844]_  = \new_[46843]_  & \new_[46840]_ ;
  assign \new_[46845]_  = \new_[46844]_  & \new_[46837]_ ;
  assign \new_[46848]_  = ~A268 & A267;
  assign \new_[46851]_  = ~A298 & A269;
  assign \new_[46852]_  = \new_[46851]_  & \new_[46848]_ ;
  assign \new_[46855]_  = ~A300 & A299;
  assign \new_[46858]_  = A302 & ~A301;
  assign \new_[46859]_  = \new_[46858]_  & \new_[46855]_ ;
  assign \new_[46860]_  = \new_[46859]_  & \new_[46852]_ ;
  assign \new_[46863]_  = A200 & ~A199;
  assign \new_[46866]_  = ~A203 & A201;
  assign \new_[46867]_  = \new_[46866]_  & \new_[46863]_ ;
  assign \new_[46870]_  = ~A233 & A232;
  assign \new_[46873]_  = ~A235 & ~A234;
  assign \new_[46874]_  = \new_[46873]_  & \new_[46870]_ ;
  assign \new_[46875]_  = \new_[46874]_  & \new_[46867]_ ;
  assign \new_[46878]_  = A267 & A236;
  assign \new_[46881]_  = A269 & ~A268;
  assign \new_[46882]_  = \new_[46881]_  & \new_[46878]_ ;
  assign \new_[46885]_  = ~A299 & A298;
  assign \new_[46888]_  = A301 & A300;
  assign \new_[46889]_  = \new_[46888]_  & \new_[46885]_ ;
  assign \new_[46890]_  = \new_[46889]_  & \new_[46882]_ ;
  assign \new_[46893]_  = A200 & ~A199;
  assign \new_[46896]_  = ~A203 & A201;
  assign \new_[46897]_  = \new_[46896]_  & \new_[46893]_ ;
  assign \new_[46900]_  = ~A233 & A232;
  assign \new_[46903]_  = ~A235 & ~A234;
  assign \new_[46904]_  = \new_[46903]_  & \new_[46900]_ ;
  assign \new_[46905]_  = \new_[46904]_  & \new_[46897]_ ;
  assign \new_[46908]_  = A267 & A236;
  assign \new_[46911]_  = A269 & ~A268;
  assign \new_[46912]_  = \new_[46911]_  & \new_[46908]_ ;
  assign \new_[46915]_  = ~A299 & A298;
  assign \new_[46918]_  = ~A302 & A300;
  assign \new_[46919]_  = \new_[46918]_  & \new_[46915]_ ;
  assign \new_[46920]_  = \new_[46919]_  & \new_[46912]_ ;
  assign \new_[46923]_  = A200 & ~A199;
  assign \new_[46926]_  = ~A203 & A201;
  assign \new_[46927]_  = \new_[46926]_  & \new_[46923]_ ;
  assign \new_[46930]_  = ~A233 & A232;
  assign \new_[46933]_  = ~A235 & ~A234;
  assign \new_[46934]_  = \new_[46933]_  & \new_[46930]_ ;
  assign \new_[46935]_  = \new_[46934]_  & \new_[46927]_ ;
  assign \new_[46938]_  = A267 & A236;
  assign \new_[46941]_  = A269 & ~A268;
  assign \new_[46942]_  = \new_[46941]_  & \new_[46938]_ ;
  assign \new_[46945]_  = A299 & ~A298;
  assign \new_[46948]_  = A301 & A300;
  assign \new_[46949]_  = \new_[46948]_  & \new_[46945]_ ;
  assign \new_[46950]_  = \new_[46949]_  & \new_[46942]_ ;
  assign \new_[46953]_  = A200 & ~A199;
  assign \new_[46956]_  = ~A203 & A201;
  assign \new_[46957]_  = \new_[46956]_  & \new_[46953]_ ;
  assign \new_[46960]_  = ~A233 & A232;
  assign \new_[46963]_  = ~A235 & ~A234;
  assign \new_[46964]_  = \new_[46963]_  & \new_[46960]_ ;
  assign \new_[46965]_  = \new_[46964]_  & \new_[46957]_ ;
  assign \new_[46968]_  = A267 & A236;
  assign \new_[46971]_  = A269 & ~A268;
  assign \new_[46972]_  = \new_[46971]_  & \new_[46968]_ ;
  assign \new_[46975]_  = A299 & ~A298;
  assign \new_[46978]_  = ~A302 & A300;
  assign \new_[46979]_  = \new_[46978]_  & \new_[46975]_ ;
  assign \new_[46980]_  = \new_[46979]_  & \new_[46972]_ ;
  assign \new_[46983]_  = A200 & ~A199;
  assign \new_[46986]_  = ~A203 & A201;
  assign \new_[46987]_  = \new_[46986]_  & \new_[46983]_ ;
  assign \new_[46990]_  = ~A233 & A232;
  assign \new_[46993]_  = ~A235 & ~A234;
  assign \new_[46994]_  = \new_[46993]_  & \new_[46990]_ ;
  assign \new_[46995]_  = \new_[46994]_  & \new_[46987]_ ;
  assign \new_[46998]_  = ~A267 & A236;
  assign \new_[47001]_  = A298 & A268;
  assign \new_[47002]_  = \new_[47001]_  & \new_[46998]_ ;
  assign \new_[47005]_  = ~A300 & ~A299;
  assign \new_[47008]_  = A302 & ~A301;
  assign \new_[47009]_  = \new_[47008]_  & \new_[47005]_ ;
  assign \new_[47010]_  = \new_[47009]_  & \new_[47002]_ ;
  assign \new_[47013]_  = A200 & ~A199;
  assign \new_[47016]_  = ~A203 & A201;
  assign \new_[47017]_  = \new_[47016]_  & \new_[47013]_ ;
  assign \new_[47020]_  = ~A233 & A232;
  assign \new_[47023]_  = ~A235 & ~A234;
  assign \new_[47024]_  = \new_[47023]_  & \new_[47020]_ ;
  assign \new_[47025]_  = \new_[47024]_  & \new_[47017]_ ;
  assign \new_[47028]_  = ~A267 & A236;
  assign \new_[47031]_  = ~A298 & A268;
  assign \new_[47032]_  = \new_[47031]_  & \new_[47028]_ ;
  assign \new_[47035]_  = ~A300 & A299;
  assign \new_[47038]_  = A302 & ~A301;
  assign \new_[47039]_  = \new_[47038]_  & \new_[47035]_ ;
  assign \new_[47040]_  = \new_[47039]_  & \new_[47032]_ ;
  assign \new_[47043]_  = A200 & ~A199;
  assign \new_[47046]_  = ~A203 & A201;
  assign \new_[47047]_  = \new_[47046]_  & \new_[47043]_ ;
  assign \new_[47050]_  = ~A233 & A232;
  assign \new_[47053]_  = ~A235 & ~A234;
  assign \new_[47054]_  = \new_[47053]_  & \new_[47050]_ ;
  assign \new_[47055]_  = \new_[47054]_  & \new_[47047]_ ;
  assign \new_[47058]_  = ~A267 & A236;
  assign \new_[47061]_  = A298 & ~A269;
  assign \new_[47062]_  = \new_[47061]_  & \new_[47058]_ ;
  assign \new_[47065]_  = ~A300 & ~A299;
  assign \new_[47068]_  = A302 & ~A301;
  assign \new_[47069]_  = \new_[47068]_  & \new_[47065]_ ;
  assign \new_[47070]_  = \new_[47069]_  & \new_[47062]_ ;
  assign \new_[47073]_  = A200 & ~A199;
  assign \new_[47076]_  = ~A203 & A201;
  assign \new_[47077]_  = \new_[47076]_  & \new_[47073]_ ;
  assign \new_[47080]_  = ~A233 & A232;
  assign \new_[47083]_  = ~A235 & ~A234;
  assign \new_[47084]_  = \new_[47083]_  & \new_[47080]_ ;
  assign \new_[47085]_  = \new_[47084]_  & \new_[47077]_ ;
  assign \new_[47088]_  = ~A267 & A236;
  assign \new_[47091]_  = ~A298 & ~A269;
  assign \new_[47092]_  = \new_[47091]_  & \new_[47088]_ ;
  assign \new_[47095]_  = ~A300 & A299;
  assign \new_[47098]_  = A302 & ~A301;
  assign \new_[47099]_  = \new_[47098]_  & \new_[47095]_ ;
  assign \new_[47100]_  = \new_[47099]_  & \new_[47092]_ ;
  assign \new_[47103]_  = A200 & ~A199;
  assign \new_[47106]_  = ~A203 & A201;
  assign \new_[47107]_  = \new_[47106]_  & \new_[47103]_ ;
  assign \new_[47110]_  = ~A233 & A232;
  assign \new_[47113]_  = ~A235 & ~A234;
  assign \new_[47114]_  = \new_[47113]_  & \new_[47110]_ ;
  assign \new_[47115]_  = \new_[47114]_  & \new_[47107]_ ;
  assign \new_[47118]_  = A265 & A236;
  assign \new_[47121]_  = A298 & A266;
  assign \new_[47122]_  = \new_[47121]_  & \new_[47118]_ ;
  assign \new_[47125]_  = ~A300 & ~A299;
  assign \new_[47128]_  = A302 & ~A301;
  assign \new_[47129]_  = \new_[47128]_  & \new_[47125]_ ;
  assign \new_[47130]_  = \new_[47129]_  & \new_[47122]_ ;
  assign \new_[47133]_  = A200 & ~A199;
  assign \new_[47136]_  = ~A203 & A201;
  assign \new_[47137]_  = \new_[47136]_  & \new_[47133]_ ;
  assign \new_[47140]_  = ~A233 & A232;
  assign \new_[47143]_  = ~A235 & ~A234;
  assign \new_[47144]_  = \new_[47143]_  & \new_[47140]_ ;
  assign \new_[47145]_  = \new_[47144]_  & \new_[47137]_ ;
  assign \new_[47148]_  = A265 & A236;
  assign \new_[47151]_  = ~A298 & A266;
  assign \new_[47152]_  = \new_[47151]_  & \new_[47148]_ ;
  assign \new_[47155]_  = ~A300 & A299;
  assign \new_[47158]_  = A302 & ~A301;
  assign \new_[47159]_  = \new_[47158]_  & \new_[47155]_ ;
  assign \new_[47160]_  = \new_[47159]_  & \new_[47152]_ ;
  assign \new_[47163]_  = A200 & ~A199;
  assign \new_[47166]_  = ~A203 & A201;
  assign \new_[47167]_  = \new_[47166]_  & \new_[47163]_ ;
  assign \new_[47170]_  = ~A233 & A232;
  assign \new_[47173]_  = ~A235 & ~A234;
  assign \new_[47174]_  = \new_[47173]_  & \new_[47170]_ ;
  assign \new_[47175]_  = \new_[47174]_  & \new_[47167]_ ;
  assign \new_[47178]_  = ~A265 & A236;
  assign \new_[47181]_  = A298 & ~A266;
  assign \new_[47182]_  = \new_[47181]_  & \new_[47178]_ ;
  assign \new_[47185]_  = ~A300 & ~A299;
  assign \new_[47188]_  = A302 & ~A301;
  assign \new_[47189]_  = \new_[47188]_  & \new_[47185]_ ;
  assign \new_[47190]_  = \new_[47189]_  & \new_[47182]_ ;
  assign \new_[47193]_  = A200 & ~A199;
  assign \new_[47196]_  = ~A203 & A201;
  assign \new_[47197]_  = \new_[47196]_  & \new_[47193]_ ;
  assign \new_[47200]_  = ~A233 & A232;
  assign \new_[47203]_  = ~A235 & ~A234;
  assign \new_[47204]_  = \new_[47203]_  & \new_[47200]_ ;
  assign \new_[47205]_  = \new_[47204]_  & \new_[47197]_ ;
  assign \new_[47208]_  = ~A265 & A236;
  assign \new_[47211]_  = ~A298 & ~A266;
  assign \new_[47212]_  = \new_[47211]_  & \new_[47208]_ ;
  assign \new_[47215]_  = ~A300 & A299;
  assign \new_[47218]_  = A302 & ~A301;
  assign \new_[47219]_  = \new_[47218]_  & \new_[47215]_ ;
  assign \new_[47220]_  = \new_[47219]_  & \new_[47212]_ ;
  assign \new_[47223]_  = A200 & ~A199;
  assign \new_[47226]_  = ~A202 & ~A201;
  assign \new_[47227]_  = \new_[47226]_  & \new_[47223]_ ;
  assign \new_[47230]_  = ~A232 & A203;
  assign \new_[47233]_  = A234 & A233;
  assign \new_[47234]_  = \new_[47233]_  & \new_[47230]_ ;
  assign \new_[47235]_  = \new_[47234]_  & \new_[47227]_ ;
  assign \new_[47238]_  = A267 & A235;
  assign \new_[47241]_  = A269 & ~A268;
  assign \new_[47242]_  = \new_[47241]_  & \new_[47238]_ ;
  assign \new_[47245]_  = ~A299 & A298;
  assign \new_[47248]_  = A301 & A300;
  assign \new_[47249]_  = \new_[47248]_  & \new_[47245]_ ;
  assign \new_[47250]_  = \new_[47249]_  & \new_[47242]_ ;
  assign \new_[47253]_  = A200 & ~A199;
  assign \new_[47256]_  = ~A202 & ~A201;
  assign \new_[47257]_  = \new_[47256]_  & \new_[47253]_ ;
  assign \new_[47260]_  = ~A232 & A203;
  assign \new_[47263]_  = A234 & A233;
  assign \new_[47264]_  = \new_[47263]_  & \new_[47260]_ ;
  assign \new_[47265]_  = \new_[47264]_  & \new_[47257]_ ;
  assign \new_[47268]_  = A267 & A235;
  assign \new_[47271]_  = A269 & ~A268;
  assign \new_[47272]_  = \new_[47271]_  & \new_[47268]_ ;
  assign \new_[47275]_  = ~A299 & A298;
  assign \new_[47278]_  = ~A302 & A300;
  assign \new_[47279]_  = \new_[47278]_  & \new_[47275]_ ;
  assign \new_[47280]_  = \new_[47279]_  & \new_[47272]_ ;
  assign \new_[47283]_  = A200 & ~A199;
  assign \new_[47286]_  = ~A202 & ~A201;
  assign \new_[47287]_  = \new_[47286]_  & \new_[47283]_ ;
  assign \new_[47290]_  = ~A232 & A203;
  assign \new_[47293]_  = A234 & A233;
  assign \new_[47294]_  = \new_[47293]_  & \new_[47290]_ ;
  assign \new_[47295]_  = \new_[47294]_  & \new_[47287]_ ;
  assign \new_[47298]_  = A267 & A235;
  assign \new_[47301]_  = A269 & ~A268;
  assign \new_[47302]_  = \new_[47301]_  & \new_[47298]_ ;
  assign \new_[47305]_  = A299 & ~A298;
  assign \new_[47308]_  = A301 & A300;
  assign \new_[47309]_  = \new_[47308]_  & \new_[47305]_ ;
  assign \new_[47310]_  = \new_[47309]_  & \new_[47302]_ ;
  assign \new_[47313]_  = A200 & ~A199;
  assign \new_[47316]_  = ~A202 & ~A201;
  assign \new_[47317]_  = \new_[47316]_  & \new_[47313]_ ;
  assign \new_[47320]_  = ~A232 & A203;
  assign \new_[47323]_  = A234 & A233;
  assign \new_[47324]_  = \new_[47323]_  & \new_[47320]_ ;
  assign \new_[47325]_  = \new_[47324]_  & \new_[47317]_ ;
  assign \new_[47328]_  = A267 & A235;
  assign \new_[47331]_  = A269 & ~A268;
  assign \new_[47332]_  = \new_[47331]_  & \new_[47328]_ ;
  assign \new_[47335]_  = A299 & ~A298;
  assign \new_[47338]_  = ~A302 & A300;
  assign \new_[47339]_  = \new_[47338]_  & \new_[47335]_ ;
  assign \new_[47340]_  = \new_[47339]_  & \new_[47332]_ ;
  assign \new_[47343]_  = A200 & ~A199;
  assign \new_[47346]_  = ~A202 & ~A201;
  assign \new_[47347]_  = \new_[47346]_  & \new_[47343]_ ;
  assign \new_[47350]_  = ~A232 & A203;
  assign \new_[47353]_  = A234 & A233;
  assign \new_[47354]_  = \new_[47353]_  & \new_[47350]_ ;
  assign \new_[47355]_  = \new_[47354]_  & \new_[47347]_ ;
  assign \new_[47358]_  = ~A267 & A235;
  assign \new_[47361]_  = A298 & A268;
  assign \new_[47362]_  = \new_[47361]_  & \new_[47358]_ ;
  assign \new_[47365]_  = ~A300 & ~A299;
  assign \new_[47368]_  = A302 & ~A301;
  assign \new_[47369]_  = \new_[47368]_  & \new_[47365]_ ;
  assign \new_[47370]_  = \new_[47369]_  & \new_[47362]_ ;
  assign \new_[47373]_  = A200 & ~A199;
  assign \new_[47376]_  = ~A202 & ~A201;
  assign \new_[47377]_  = \new_[47376]_  & \new_[47373]_ ;
  assign \new_[47380]_  = ~A232 & A203;
  assign \new_[47383]_  = A234 & A233;
  assign \new_[47384]_  = \new_[47383]_  & \new_[47380]_ ;
  assign \new_[47385]_  = \new_[47384]_  & \new_[47377]_ ;
  assign \new_[47388]_  = ~A267 & A235;
  assign \new_[47391]_  = ~A298 & A268;
  assign \new_[47392]_  = \new_[47391]_  & \new_[47388]_ ;
  assign \new_[47395]_  = ~A300 & A299;
  assign \new_[47398]_  = A302 & ~A301;
  assign \new_[47399]_  = \new_[47398]_  & \new_[47395]_ ;
  assign \new_[47400]_  = \new_[47399]_  & \new_[47392]_ ;
  assign \new_[47403]_  = A200 & ~A199;
  assign \new_[47406]_  = ~A202 & ~A201;
  assign \new_[47407]_  = \new_[47406]_  & \new_[47403]_ ;
  assign \new_[47410]_  = ~A232 & A203;
  assign \new_[47413]_  = A234 & A233;
  assign \new_[47414]_  = \new_[47413]_  & \new_[47410]_ ;
  assign \new_[47415]_  = \new_[47414]_  & \new_[47407]_ ;
  assign \new_[47418]_  = ~A267 & A235;
  assign \new_[47421]_  = A298 & ~A269;
  assign \new_[47422]_  = \new_[47421]_  & \new_[47418]_ ;
  assign \new_[47425]_  = ~A300 & ~A299;
  assign \new_[47428]_  = A302 & ~A301;
  assign \new_[47429]_  = \new_[47428]_  & \new_[47425]_ ;
  assign \new_[47430]_  = \new_[47429]_  & \new_[47422]_ ;
  assign \new_[47433]_  = A200 & ~A199;
  assign \new_[47436]_  = ~A202 & ~A201;
  assign \new_[47437]_  = \new_[47436]_  & \new_[47433]_ ;
  assign \new_[47440]_  = ~A232 & A203;
  assign \new_[47443]_  = A234 & A233;
  assign \new_[47444]_  = \new_[47443]_  & \new_[47440]_ ;
  assign \new_[47445]_  = \new_[47444]_  & \new_[47437]_ ;
  assign \new_[47448]_  = ~A267 & A235;
  assign \new_[47451]_  = ~A298 & ~A269;
  assign \new_[47452]_  = \new_[47451]_  & \new_[47448]_ ;
  assign \new_[47455]_  = ~A300 & A299;
  assign \new_[47458]_  = A302 & ~A301;
  assign \new_[47459]_  = \new_[47458]_  & \new_[47455]_ ;
  assign \new_[47460]_  = \new_[47459]_  & \new_[47452]_ ;
  assign \new_[47463]_  = A200 & ~A199;
  assign \new_[47466]_  = ~A202 & ~A201;
  assign \new_[47467]_  = \new_[47466]_  & \new_[47463]_ ;
  assign \new_[47470]_  = ~A232 & A203;
  assign \new_[47473]_  = A234 & A233;
  assign \new_[47474]_  = \new_[47473]_  & \new_[47470]_ ;
  assign \new_[47475]_  = \new_[47474]_  & \new_[47467]_ ;
  assign \new_[47478]_  = A265 & A235;
  assign \new_[47481]_  = A298 & A266;
  assign \new_[47482]_  = \new_[47481]_  & \new_[47478]_ ;
  assign \new_[47485]_  = ~A300 & ~A299;
  assign \new_[47488]_  = A302 & ~A301;
  assign \new_[47489]_  = \new_[47488]_  & \new_[47485]_ ;
  assign \new_[47490]_  = \new_[47489]_  & \new_[47482]_ ;
  assign \new_[47493]_  = A200 & ~A199;
  assign \new_[47496]_  = ~A202 & ~A201;
  assign \new_[47497]_  = \new_[47496]_  & \new_[47493]_ ;
  assign \new_[47500]_  = ~A232 & A203;
  assign \new_[47503]_  = A234 & A233;
  assign \new_[47504]_  = \new_[47503]_  & \new_[47500]_ ;
  assign \new_[47505]_  = \new_[47504]_  & \new_[47497]_ ;
  assign \new_[47508]_  = A265 & A235;
  assign \new_[47511]_  = ~A298 & A266;
  assign \new_[47512]_  = \new_[47511]_  & \new_[47508]_ ;
  assign \new_[47515]_  = ~A300 & A299;
  assign \new_[47518]_  = A302 & ~A301;
  assign \new_[47519]_  = \new_[47518]_  & \new_[47515]_ ;
  assign \new_[47520]_  = \new_[47519]_  & \new_[47512]_ ;
  assign \new_[47523]_  = A200 & ~A199;
  assign \new_[47526]_  = ~A202 & ~A201;
  assign \new_[47527]_  = \new_[47526]_  & \new_[47523]_ ;
  assign \new_[47530]_  = ~A232 & A203;
  assign \new_[47533]_  = A234 & A233;
  assign \new_[47534]_  = \new_[47533]_  & \new_[47530]_ ;
  assign \new_[47535]_  = \new_[47534]_  & \new_[47527]_ ;
  assign \new_[47538]_  = ~A265 & A235;
  assign \new_[47541]_  = A298 & ~A266;
  assign \new_[47542]_  = \new_[47541]_  & \new_[47538]_ ;
  assign \new_[47545]_  = ~A300 & ~A299;
  assign \new_[47548]_  = A302 & ~A301;
  assign \new_[47549]_  = \new_[47548]_  & \new_[47545]_ ;
  assign \new_[47550]_  = \new_[47549]_  & \new_[47542]_ ;
  assign \new_[47553]_  = A200 & ~A199;
  assign \new_[47556]_  = ~A202 & ~A201;
  assign \new_[47557]_  = \new_[47556]_  & \new_[47553]_ ;
  assign \new_[47560]_  = ~A232 & A203;
  assign \new_[47563]_  = A234 & A233;
  assign \new_[47564]_  = \new_[47563]_  & \new_[47560]_ ;
  assign \new_[47565]_  = \new_[47564]_  & \new_[47557]_ ;
  assign \new_[47568]_  = ~A265 & A235;
  assign \new_[47571]_  = ~A298 & ~A266;
  assign \new_[47572]_  = \new_[47571]_  & \new_[47568]_ ;
  assign \new_[47575]_  = ~A300 & A299;
  assign \new_[47578]_  = A302 & ~A301;
  assign \new_[47579]_  = \new_[47578]_  & \new_[47575]_ ;
  assign \new_[47580]_  = \new_[47579]_  & \new_[47572]_ ;
  assign \new_[47583]_  = A200 & ~A199;
  assign \new_[47586]_  = ~A202 & ~A201;
  assign \new_[47587]_  = \new_[47586]_  & \new_[47583]_ ;
  assign \new_[47590]_  = ~A232 & A203;
  assign \new_[47593]_  = A234 & A233;
  assign \new_[47594]_  = \new_[47593]_  & \new_[47590]_ ;
  assign \new_[47595]_  = \new_[47594]_  & \new_[47587]_ ;
  assign \new_[47598]_  = A267 & ~A236;
  assign \new_[47601]_  = A269 & ~A268;
  assign \new_[47602]_  = \new_[47601]_  & \new_[47598]_ ;
  assign \new_[47605]_  = ~A299 & A298;
  assign \new_[47608]_  = A301 & A300;
  assign \new_[47609]_  = \new_[47608]_  & \new_[47605]_ ;
  assign \new_[47610]_  = \new_[47609]_  & \new_[47602]_ ;
  assign \new_[47613]_  = A200 & ~A199;
  assign \new_[47616]_  = ~A202 & ~A201;
  assign \new_[47617]_  = \new_[47616]_  & \new_[47613]_ ;
  assign \new_[47620]_  = ~A232 & A203;
  assign \new_[47623]_  = A234 & A233;
  assign \new_[47624]_  = \new_[47623]_  & \new_[47620]_ ;
  assign \new_[47625]_  = \new_[47624]_  & \new_[47617]_ ;
  assign \new_[47628]_  = A267 & ~A236;
  assign \new_[47631]_  = A269 & ~A268;
  assign \new_[47632]_  = \new_[47631]_  & \new_[47628]_ ;
  assign \new_[47635]_  = ~A299 & A298;
  assign \new_[47638]_  = ~A302 & A300;
  assign \new_[47639]_  = \new_[47638]_  & \new_[47635]_ ;
  assign \new_[47640]_  = \new_[47639]_  & \new_[47632]_ ;
  assign \new_[47643]_  = A200 & ~A199;
  assign \new_[47646]_  = ~A202 & ~A201;
  assign \new_[47647]_  = \new_[47646]_  & \new_[47643]_ ;
  assign \new_[47650]_  = ~A232 & A203;
  assign \new_[47653]_  = A234 & A233;
  assign \new_[47654]_  = \new_[47653]_  & \new_[47650]_ ;
  assign \new_[47655]_  = \new_[47654]_  & \new_[47647]_ ;
  assign \new_[47658]_  = A267 & ~A236;
  assign \new_[47661]_  = A269 & ~A268;
  assign \new_[47662]_  = \new_[47661]_  & \new_[47658]_ ;
  assign \new_[47665]_  = A299 & ~A298;
  assign \new_[47668]_  = A301 & A300;
  assign \new_[47669]_  = \new_[47668]_  & \new_[47665]_ ;
  assign \new_[47670]_  = \new_[47669]_  & \new_[47662]_ ;
  assign \new_[47673]_  = A200 & ~A199;
  assign \new_[47676]_  = ~A202 & ~A201;
  assign \new_[47677]_  = \new_[47676]_  & \new_[47673]_ ;
  assign \new_[47680]_  = ~A232 & A203;
  assign \new_[47683]_  = A234 & A233;
  assign \new_[47684]_  = \new_[47683]_  & \new_[47680]_ ;
  assign \new_[47685]_  = \new_[47684]_  & \new_[47677]_ ;
  assign \new_[47688]_  = A267 & ~A236;
  assign \new_[47691]_  = A269 & ~A268;
  assign \new_[47692]_  = \new_[47691]_  & \new_[47688]_ ;
  assign \new_[47695]_  = A299 & ~A298;
  assign \new_[47698]_  = ~A302 & A300;
  assign \new_[47699]_  = \new_[47698]_  & \new_[47695]_ ;
  assign \new_[47700]_  = \new_[47699]_  & \new_[47692]_ ;
  assign \new_[47703]_  = A200 & ~A199;
  assign \new_[47706]_  = ~A202 & ~A201;
  assign \new_[47707]_  = \new_[47706]_  & \new_[47703]_ ;
  assign \new_[47710]_  = ~A232 & A203;
  assign \new_[47713]_  = A234 & A233;
  assign \new_[47714]_  = \new_[47713]_  & \new_[47710]_ ;
  assign \new_[47715]_  = \new_[47714]_  & \new_[47707]_ ;
  assign \new_[47718]_  = ~A267 & ~A236;
  assign \new_[47721]_  = A298 & A268;
  assign \new_[47722]_  = \new_[47721]_  & \new_[47718]_ ;
  assign \new_[47725]_  = ~A300 & ~A299;
  assign \new_[47728]_  = A302 & ~A301;
  assign \new_[47729]_  = \new_[47728]_  & \new_[47725]_ ;
  assign \new_[47730]_  = \new_[47729]_  & \new_[47722]_ ;
  assign \new_[47733]_  = A200 & ~A199;
  assign \new_[47736]_  = ~A202 & ~A201;
  assign \new_[47737]_  = \new_[47736]_  & \new_[47733]_ ;
  assign \new_[47740]_  = ~A232 & A203;
  assign \new_[47743]_  = A234 & A233;
  assign \new_[47744]_  = \new_[47743]_  & \new_[47740]_ ;
  assign \new_[47745]_  = \new_[47744]_  & \new_[47737]_ ;
  assign \new_[47748]_  = ~A267 & ~A236;
  assign \new_[47751]_  = ~A298 & A268;
  assign \new_[47752]_  = \new_[47751]_  & \new_[47748]_ ;
  assign \new_[47755]_  = ~A300 & A299;
  assign \new_[47758]_  = A302 & ~A301;
  assign \new_[47759]_  = \new_[47758]_  & \new_[47755]_ ;
  assign \new_[47760]_  = \new_[47759]_  & \new_[47752]_ ;
  assign \new_[47763]_  = A200 & ~A199;
  assign \new_[47766]_  = ~A202 & ~A201;
  assign \new_[47767]_  = \new_[47766]_  & \new_[47763]_ ;
  assign \new_[47770]_  = ~A232 & A203;
  assign \new_[47773]_  = A234 & A233;
  assign \new_[47774]_  = \new_[47773]_  & \new_[47770]_ ;
  assign \new_[47775]_  = \new_[47774]_  & \new_[47767]_ ;
  assign \new_[47778]_  = ~A267 & ~A236;
  assign \new_[47781]_  = A298 & ~A269;
  assign \new_[47782]_  = \new_[47781]_  & \new_[47778]_ ;
  assign \new_[47785]_  = ~A300 & ~A299;
  assign \new_[47788]_  = A302 & ~A301;
  assign \new_[47789]_  = \new_[47788]_  & \new_[47785]_ ;
  assign \new_[47790]_  = \new_[47789]_  & \new_[47782]_ ;
  assign \new_[47793]_  = A200 & ~A199;
  assign \new_[47796]_  = ~A202 & ~A201;
  assign \new_[47797]_  = \new_[47796]_  & \new_[47793]_ ;
  assign \new_[47800]_  = ~A232 & A203;
  assign \new_[47803]_  = A234 & A233;
  assign \new_[47804]_  = \new_[47803]_  & \new_[47800]_ ;
  assign \new_[47805]_  = \new_[47804]_  & \new_[47797]_ ;
  assign \new_[47808]_  = ~A267 & ~A236;
  assign \new_[47811]_  = ~A298 & ~A269;
  assign \new_[47812]_  = \new_[47811]_  & \new_[47808]_ ;
  assign \new_[47815]_  = ~A300 & A299;
  assign \new_[47818]_  = A302 & ~A301;
  assign \new_[47819]_  = \new_[47818]_  & \new_[47815]_ ;
  assign \new_[47820]_  = \new_[47819]_  & \new_[47812]_ ;
  assign \new_[47823]_  = A200 & ~A199;
  assign \new_[47826]_  = ~A202 & ~A201;
  assign \new_[47827]_  = \new_[47826]_  & \new_[47823]_ ;
  assign \new_[47830]_  = ~A232 & A203;
  assign \new_[47833]_  = A234 & A233;
  assign \new_[47834]_  = \new_[47833]_  & \new_[47830]_ ;
  assign \new_[47835]_  = \new_[47834]_  & \new_[47827]_ ;
  assign \new_[47838]_  = A265 & ~A236;
  assign \new_[47841]_  = A298 & A266;
  assign \new_[47842]_  = \new_[47841]_  & \new_[47838]_ ;
  assign \new_[47845]_  = ~A300 & ~A299;
  assign \new_[47848]_  = A302 & ~A301;
  assign \new_[47849]_  = \new_[47848]_  & \new_[47845]_ ;
  assign \new_[47850]_  = \new_[47849]_  & \new_[47842]_ ;
  assign \new_[47853]_  = A200 & ~A199;
  assign \new_[47856]_  = ~A202 & ~A201;
  assign \new_[47857]_  = \new_[47856]_  & \new_[47853]_ ;
  assign \new_[47860]_  = ~A232 & A203;
  assign \new_[47863]_  = A234 & A233;
  assign \new_[47864]_  = \new_[47863]_  & \new_[47860]_ ;
  assign \new_[47865]_  = \new_[47864]_  & \new_[47857]_ ;
  assign \new_[47868]_  = A265 & ~A236;
  assign \new_[47871]_  = ~A298 & A266;
  assign \new_[47872]_  = \new_[47871]_  & \new_[47868]_ ;
  assign \new_[47875]_  = ~A300 & A299;
  assign \new_[47878]_  = A302 & ~A301;
  assign \new_[47879]_  = \new_[47878]_  & \new_[47875]_ ;
  assign \new_[47880]_  = \new_[47879]_  & \new_[47872]_ ;
  assign \new_[47883]_  = A200 & ~A199;
  assign \new_[47886]_  = ~A202 & ~A201;
  assign \new_[47887]_  = \new_[47886]_  & \new_[47883]_ ;
  assign \new_[47890]_  = ~A232 & A203;
  assign \new_[47893]_  = A234 & A233;
  assign \new_[47894]_  = \new_[47893]_  & \new_[47890]_ ;
  assign \new_[47895]_  = \new_[47894]_  & \new_[47887]_ ;
  assign \new_[47898]_  = ~A265 & ~A236;
  assign \new_[47901]_  = A298 & ~A266;
  assign \new_[47902]_  = \new_[47901]_  & \new_[47898]_ ;
  assign \new_[47905]_  = ~A300 & ~A299;
  assign \new_[47908]_  = A302 & ~A301;
  assign \new_[47909]_  = \new_[47908]_  & \new_[47905]_ ;
  assign \new_[47910]_  = \new_[47909]_  & \new_[47902]_ ;
  assign \new_[47913]_  = A200 & ~A199;
  assign \new_[47916]_  = ~A202 & ~A201;
  assign \new_[47917]_  = \new_[47916]_  & \new_[47913]_ ;
  assign \new_[47920]_  = ~A232 & A203;
  assign \new_[47923]_  = A234 & A233;
  assign \new_[47924]_  = \new_[47923]_  & \new_[47920]_ ;
  assign \new_[47925]_  = \new_[47924]_  & \new_[47917]_ ;
  assign \new_[47928]_  = ~A265 & ~A236;
  assign \new_[47931]_  = ~A298 & ~A266;
  assign \new_[47932]_  = \new_[47931]_  & \new_[47928]_ ;
  assign \new_[47935]_  = ~A300 & A299;
  assign \new_[47938]_  = A302 & ~A301;
  assign \new_[47939]_  = \new_[47938]_  & \new_[47935]_ ;
  assign \new_[47940]_  = \new_[47939]_  & \new_[47932]_ ;
  assign \new_[47943]_  = A200 & ~A199;
  assign \new_[47946]_  = ~A202 & ~A201;
  assign \new_[47947]_  = \new_[47946]_  & \new_[47943]_ ;
  assign \new_[47950]_  = ~A232 & A203;
  assign \new_[47953]_  = ~A234 & A233;
  assign \new_[47954]_  = \new_[47953]_  & \new_[47950]_ ;
  assign \new_[47955]_  = \new_[47954]_  & \new_[47947]_ ;
  assign \new_[47958]_  = A236 & ~A235;
  assign \new_[47961]_  = A268 & ~A267;
  assign \new_[47962]_  = \new_[47961]_  & \new_[47958]_ ;
  assign \new_[47965]_  = ~A299 & A298;
  assign \new_[47968]_  = A301 & A300;
  assign \new_[47969]_  = \new_[47968]_  & \new_[47965]_ ;
  assign \new_[47970]_  = \new_[47969]_  & \new_[47962]_ ;
  assign \new_[47973]_  = A200 & ~A199;
  assign \new_[47976]_  = ~A202 & ~A201;
  assign \new_[47977]_  = \new_[47976]_  & \new_[47973]_ ;
  assign \new_[47980]_  = ~A232 & A203;
  assign \new_[47983]_  = ~A234 & A233;
  assign \new_[47984]_  = \new_[47983]_  & \new_[47980]_ ;
  assign \new_[47985]_  = \new_[47984]_  & \new_[47977]_ ;
  assign \new_[47988]_  = A236 & ~A235;
  assign \new_[47991]_  = A268 & ~A267;
  assign \new_[47992]_  = \new_[47991]_  & \new_[47988]_ ;
  assign \new_[47995]_  = ~A299 & A298;
  assign \new_[47998]_  = ~A302 & A300;
  assign \new_[47999]_  = \new_[47998]_  & \new_[47995]_ ;
  assign \new_[48000]_  = \new_[47999]_  & \new_[47992]_ ;
  assign \new_[48003]_  = A200 & ~A199;
  assign \new_[48006]_  = ~A202 & ~A201;
  assign \new_[48007]_  = \new_[48006]_  & \new_[48003]_ ;
  assign \new_[48010]_  = ~A232 & A203;
  assign \new_[48013]_  = ~A234 & A233;
  assign \new_[48014]_  = \new_[48013]_  & \new_[48010]_ ;
  assign \new_[48015]_  = \new_[48014]_  & \new_[48007]_ ;
  assign \new_[48018]_  = A236 & ~A235;
  assign \new_[48021]_  = A268 & ~A267;
  assign \new_[48022]_  = \new_[48021]_  & \new_[48018]_ ;
  assign \new_[48025]_  = A299 & ~A298;
  assign \new_[48028]_  = A301 & A300;
  assign \new_[48029]_  = \new_[48028]_  & \new_[48025]_ ;
  assign \new_[48030]_  = \new_[48029]_  & \new_[48022]_ ;
  assign \new_[48033]_  = A200 & ~A199;
  assign \new_[48036]_  = ~A202 & ~A201;
  assign \new_[48037]_  = \new_[48036]_  & \new_[48033]_ ;
  assign \new_[48040]_  = ~A232 & A203;
  assign \new_[48043]_  = ~A234 & A233;
  assign \new_[48044]_  = \new_[48043]_  & \new_[48040]_ ;
  assign \new_[48045]_  = \new_[48044]_  & \new_[48037]_ ;
  assign \new_[48048]_  = A236 & ~A235;
  assign \new_[48051]_  = A268 & ~A267;
  assign \new_[48052]_  = \new_[48051]_  & \new_[48048]_ ;
  assign \new_[48055]_  = A299 & ~A298;
  assign \new_[48058]_  = ~A302 & A300;
  assign \new_[48059]_  = \new_[48058]_  & \new_[48055]_ ;
  assign \new_[48060]_  = \new_[48059]_  & \new_[48052]_ ;
  assign \new_[48063]_  = A200 & ~A199;
  assign \new_[48066]_  = ~A202 & ~A201;
  assign \new_[48067]_  = \new_[48066]_  & \new_[48063]_ ;
  assign \new_[48070]_  = ~A232 & A203;
  assign \new_[48073]_  = ~A234 & A233;
  assign \new_[48074]_  = \new_[48073]_  & \new_[48070]_ ;
  assign \new_[48075]_  = \new_[48074]_  & \new_[48067]_ ;
  assign \new_[48078]_  = A236 & ~A235;
  assign \new_[48081]_  = ~A269 & ~A267;
  assign \new_[48082]_  = \new_[48081]_  & \new_[48078]_ ;
  assign \new_[48085]_  = ~A299 & A298;
  assign \new_[48088]_  = A301 & A300;
  assign \new_[48089]_  = \new_[48088]_  & \new_[48085]_ ;
  assign \new_[48090]_  = \new_[48089]_  & \new_[48082]_ ;
  assign \new_[48093]_  = A200 & ~A199;
  assign \new_[48096]_  = ~A202 & ~A201;
  assign \new_[48097]_  = \new_[48096]_  & \new_[48093]_ ;
  assign \new_[48100]_  = ~A232 & A203;
  assign \new_[48103]_  = ~A234 & A233;
  assign \new_[48104]_  = \new_[48103]_  & \new_[48100]_ ;
  assign \new_[48105]_  = \new_[48104]_  & \new_[48097]_ ;
  assign \new_[48108]_  = A236 & ~A235;
  assign \new_[48111]_  = ~A269 & ~A267;
  assign \new_[48112]_  = \new_[48111]_  & \new_[48108]_ ;
  assign \new_[48115]_  = ~A299 & A298;
  assign \new_[48118]_  = ~A302 & A300;
  assign \new_[48119]_  = \new_[48118]_  & \new_[48115]_ ;
  assign \new_[48120]_  = \new_[48119]_  & \new_[48112]_ ;
  assign \new_[48123]_  = A200 & ~A199;
  assign \new_[48126]_  = ~A202 & ~A201;
  assign \new_[48127]_  = \new_[48126]_  & \new_[48123]_ ;
  assign \new_[48130]_  = ~A232 & A203;
  assign \new_[48133]_  = ~A234 & A233;
  assign \new_[48134]_  = \new_[48133]_  & \new_[48130]_ ;
  assign \new_[48135]_  = \new_[48134]_  & \new_[48127]_ ;
  assign \new_[48138]_  = A236 & ~A235;
  assign \new_[48141]_  = ~A269 & ~A267;
  assign \new_[48142]_  = \new_[48141]_  & \new_[48138]_ ;
  assign \new_[48145]_  = A299 & ~A298;
  assign \new_[48148]_  = A301 & A300;
  assign \new_[48149]_  = \new_[48148]_  & \new_[48145]_ ;
  assign \new_[48150]_  = \new_[48149]_  & \new_[48142]_ ;
  assign \new_[48153]_  = A200 & ~A199;
  assign \new_[48156]_  = ~A202 & ~A201;
  assign \new_[48157]_  = \new_[48156]_  & \new_[48153]_ ;
  assign \new_[48160]_  = ~A232 & A203;
  assign \new_[48163]_  = ~A234 & A233;
  assign \new_[48164]_  = \new_[48163]_  & \new_[48160]_ ;
  assign \new_[48165]_  = \new_[48164]_  & \new_[48157]_ ;
  assign \new_[48168]_  = A236 & ~A235;
  assign \new_[48171]_  = ~A269 & ~A267;
  assign \new_[48172]_  = \new_[48171]_  & \new_[48168]_ ;
  assign \new_[48175]_  = A299 & ~A298;
  assign \new_[48178]_  = ~A302 & A300;
  assign \new_[48179]_  = \new_[48178]_  & \new_[48175]_ ;
  assign \new_[48180]_  = \new_[48179]_  & \new_[48172]_ ;
  assign \new_[48183]_  = A200 & ~A199;
  assign \new_[48186]_  = ~A202 & ~A201;
  assign \new_[48187]_  = \new_[48186]_  & \new_[48183]_ ;
  assign \new_[48190]_  = ~A232 & A203;
  assign \new_[48193]_  = ~A234 & A233;
  assign \new_[48194]_  = \new_[48193]_  & \new_[48190]_ ;
  assign \new_[48195]_  = \new_[48194]_  & \new_[48187]_ ;
  assign \new_[48198]_  = A236 & ~A235;
  assign \new_[48201]_  = A266 & A265;
  assign \new_[48202]_  = \new_[48201]_  & \new_[48198]_ ;
  assign \new_[48205]_  = ~A299 & A298;
  assign \new_[48208]_  = A301 & A300;
  assign \new_[48209]_  = \new_[48208]_  & \new_[48205]_ ;
  assign \new_[48210]_  = \new_[48209]_  & \new_[48202]_ ;
  assign \new_[48213]_  = A200 & ~A199;
  assign \new_[48216]_  = ~A202 & ~A201;
  assign \new_[48217]_  = \new_[48216]_  & \new_[48213]_ ;
  assign \new_[48220]_  = ~A232 & A203;
  assign \new_[48223]_  = ~A234 & A233;
  assign \new_[48224]_  = \new_[48223]_  & \new_[48220]_ ;
  assign \new_[48225]_  = \new_[48224]_  & \new_[48217]_ ;
  assign \new_[48228]_  = A236 & ~A235;
  assign \new_[48231]_  = A266 & A265;
  assign \new_[48232]_  = \new_[48231]_  & \new_[48228]_ ;
  assign \new_[48235]_  = ~A299 & A298;
  assign \new_[48238]_  = ~A302 & A300;
  assign \new_[48239]_  = \new_[48238]_  & \new_[48235]_ ;
  assign \new_[48240]_  = \new_[48239]_  & \new_[48232]_ ;
  assign \new_[48243]_  = A200 & ~A199;
  assign \new_[48246]_  = ~A202 & ~A201;
  assign \new_[48247]_  = \new_[48246]_  & \new_[48243]_ ;
  assign \new_[48250]_  = ~A232 & A203;
  assign \new_[48253]_  = ~A234 & A233;
  assign \new_[48254]_  = \new_[48253]_  & \new_[48250]_ ;
  assign \new_[48255]_  = \new_[48254]_  & \new_[48247]_ ;
  assign \new_[48258]_  = A236 & ~A235;
  assign \new_[48261]_  = A266 & A265;
  assign \new_[48262]_  = \new_[48261]_  & \new_[48258]_ ;
  assign \new_[48265]_  = A299 & ~A298;
  assign \new_[48268]_  = A301 & A300;
  assign \new_[48269]_  = \new_[48268]_  & \new_[48265]_ ;
  assign \new_[48270]_  = \new_[48269]_  & \new_[48262]_ ;
  assign \new_[48273]_  = A200 & ~A199;
  assign \new_[48276]_  = ~A202 & ~A201;
  assign \new_[48277]_  = \new_[48276]_  & \new_[48273]_ ;
  assign \new_[48280]_  = ~A232 & A203;
  assign \new_[48283]_  = ~A234 & A233;
  assign \new_[48284]_  = \new_[48283]_  & \new_[48280]_ ;
  assign \new_[48285]_  = \new_[48284]_  & \new_[48277]_ ;
  assign \new_[48288]_  = A236 & ~A235;
  assign \new_[48291]_  = A266 & A265;
  assign \new_[48292]_  = \new_[48291]_  & \new_[48288]_ ;
  assign \new_[48295]_  = A299 & ~A298;
  assign \new_[48298]_  = ~A302 & A300;
  assign \new_[48299]_  = \new_[48298]_  & \new_[48295]_ ;
  assign \new_[48300]_  = \new_[48299]_  & \new_[48292]_ ;
  assign \new_[48303]_  = A200 & ~A199;
  assign \new_[48306]_  = ~A202 & ~A201;
  assign \new_[48307]_  = \new_[48306]_  & \new_[48303]_ ;
  assign \new_[48310]_  = ~A232 & A203;
  assign \new_[48313]_  = ~A234 & A233;
  assign \new_[48314]_  = \new_[48313]_  & \new_[48310]_ ;
  assign \new_[48315]_  = \new_[48314]_  & \new_[48307]_ ;
  assign \new_[48318]_  = A236 & ~A235;
  assign \new_[48321]_  = ~A266 & ~A265;
  assign \new_[48322]_  = \new_[48321]_  & \new_[48318]_ ;
  assign \new_[48325]_  = ~A299 & A298;
  assign \new_[48328]_  = A301 & A300;
  assign \new_[48329]_  = \new_[48328]_  & \new_[48325]_ ;
  assign \new_[48330]_  = \new_[48329]_  & \new_[48322]_ ;
  assign \new_[48333]_  = A200 & ~A199;
  assign \new_[48336]_  = ~A202 & ~A201;
  assign \new_[48337]_  = \new_[48336]_  & \new_[48333]_ ;
  assign \new_[48340]_  = ~A232 & A203;
  assign \new_[48343]_  = ~A234 & A233;
  assign \new_[48344]_  = \new_[48343]_  & \new_[48340]_ ;
  assign \new_[48345]_  = \new_[48344]_  & \new_[48337]_ ;
  assign \new_[48348]_  = A236 & ~A235;
  assign \new_[48351]_  = ~A266 & ~A265;
  assign \new_[48352]_  = \new_[48351]_  & \new_[48348]_ ;
  assign \new_[48355]_  = ~A299 & A298;
  assign \new_[48358]_  = ~A302 & A300;
  assign \new_[48359]_  = \new_[48358]_  & \new_[48355]_ ;
  assign \new_[48360]_  = \new_[48359]_  & \new_[48352]_ ;
  assign \new_[48363]_  = A200 & ~A199;
  assign \new_[48366]_  = ~A202 & ~A201;
  assign \new_[48367]_  = \new_[48366]_  & \new_[48363]_ ;
  assign \new_[48370]_  = ~A232 & A203;
  assign \new_[48373]_  = ~A234 & A233;
  assign \new_[48374]_  = \new_[48373]_  & \new_[48370]_ ;
  assign \new_[48375]_  = \new_[48374]_  & \new_[48367]_ ;
  assign \new_[48378]_  = A236 & ~A235;
  assign \new_[48381]_  = ~A266 & ~A265;
  assign \new_[48382]_  = \new_[48381]_  & \new_[48378]_ ;
  assign \new_[48385]_  = A299 & ~A298;
  assign \new_[48388]_  = A301 & A300;
  assign \new_[48389]_  = \new_[48388]_  & \new_[48385]_ ;
  assign \new_[48390]_  = \new_[48389]_  & \new_[48382]_ ;
  assign \new_[48393]_  = A200 & ~A199;
  assign \new_[48396]_  = ~A202 & ~A201;
  assign \new_[48397]_  = \new_[48396]_  & \new_[48393]_ ;
  assign \new_[48400]_  = ~A232 & A203;
  assign \new_[48403]_  = ~A234 & A233;
  assign \new_[48404]_  = \new_[48403]_  & \new_[48400]_ ;
  assign \new_[48405]_  = \new_[48404]_  & \new_[48397]_ ;
  assign \new_[48408]_  = A236 & ~A235;
  assign \new_[48411]_  = ~A266 & ~A265;
  assign \new_[48412]_  = \new_[48411]_  & \new_[48408]_ ;
  assign \new_[48415]_  = A299 & ~A298;
  assign \new_[48418]_  = ~A302 & A300;
  assign \new_[48419]_  = \new_[48418]_  & \new_[48415]_ ;
  assign \new_[48420]_  = \new_[48419]_  & \new_[48412]_ ;
  assign \new_[48423]_  = A200 & ~A199;
  assign \new_[48426]_  = ~A202 & ~A201;
  assign \new_[48427]_  = \new_[48426]_  & \new_[48423]_ ;
  assign \new_[48430]_  = A232 & A203;
  assign \new_[48433]_  = A234 & ~A233;
  assign \new_[48434]_  = \new_[48433]_  & \new_[48430]_ ;
  assign \new_[48435]_  = \new_[48434]_  & \new_[48427]_ ;
  assign \new_[48438]_  = A267 & A235;
  assign \new_[48441]_  = A269 & ~A268;
  assign \new_[48442]_  = \new_[48441]_  & \new_[48438]_ ;
  assign \new_[48445]_  = ~A299 & A298;
  assign \new_[48448]_  = A301 & A300;
  assign \new_[48449]_  = \new_[48448]_  & \new_[48445]_ ;
  assign \new_[48450]_  = \new_[48449]_  & \new_[48442]_ ;
  assign \new_[48453]_  = A200 & ~A199;
  assign \new_[48456]_  = ~A202 & ~A201;
  assign \new_[48457]_  = \new_[48456]_  & \new_[48453]_ ;
  assign \new_[48460]_  = A232 & A203;
  assign \new_[48463]_  = A234 & ~A233;
  assign \new_[48464]_  = \new_[48463]_  & \new_[48460]_ ;
  assign \new_[48465]_  = \new_[48464]_  & \new_[48457]_ ;
  assign \new_[48468]_  = A267 & A235;
  assign \new_[48471]_  = A269 & ~A268;
  assign \new_[48472]_  = \new_[48471]_  & \new_[48468]_ ;
  assign \new_[48475]_  = ~A299 & A298;
  assign \new_[48478]_  = ~A302 & A300;
  assign \new_[48479]_  = \new_[48478]_  & \new_[48475]_ ;
  assign \new_[48480]_  = \new_[48479]_  & \new_[48472]_ ;
  assign \new_[48483]_  = A200 & ~A199;
  assign \new_[48486]_  = ~A202 & ~A201;
  assign \new_[48487]_  = \new_[48486]_  & \new_[48483]_ ;
  assign \new_[48490]_  = A232 & A203;
  assign \new_[48493]_  = A234 & ~A233;
  assign \new_[48494]_  = \new_[48493]_  & \new_[48490]_ ;
  assign \new_[48495]_  = \new_[48494]_  & \new_[48487]_ ;
  assign \new_[48498]_  = A267 & A235;
  assign \new_[48501]_  = A269 & ~A268;
  assign \new_[48502]_  = \new_[48501]_  & \new_[48498]_ ;
  assign \new_[48505]_  = A299 & ~A298;
  assign \new_[48508]_  = A301 & A300;
  assign \new_[48509]_  = \new_[48508]_  & \new_[48505]_ ;
  assign \new_[48510]_  = \new_[48509]_  & \new_[48502]_ ;
  assign \new_[48513]_  = A200 & ~A199;
  assign \new_[48516]_  = ~A202 & ~A201;
  assign \new_[48517]_  = \new_[48516]_  & \new_[48513]_ ;
  assign \new_[48520]_  = A232 & A203;
  assign \new_[48523]_  = A234 & ~A233;
  assign \new_[48524]_  = \new_[48523]_  & \new_[48520]_ ;
  assign \new_[48525]_  = \new_[48524]_  & \new_[48517]_ ;
  assign \new_[48528]_  = A267 & A235;
  assign \new_[48531]_  = A269 & ~A268;
  assign \new_[48532]_  = \new_[48531]_  & \new_[48528]_ ;
  assign \new_[48535]_  = A299 & ~A298;
  assign \new_[48538]_  = ~A302 & A300;
  assign \new_[48539]_  = \new_[48538]_  & \new_[48535]_ ;
  assign \new_[48540]_  = \new_[48539]_  & \new_[48532]_ ;
  assign \new_[48543]_  = A200 & ~A199;
  assign \new_[48546]_  = ~A202 & ~A201;
  assign \new_[48547]_  = \new_[48546]_  & \new_[48543]_ ;
  assign \new_[48550]_  = A232 & A203;
  assign \new_[48553]_  = A234 & ~A233;
  assign \new_[48554]_  = \new_[48553]_  & \new_[48550]_ ;
  assign \new_[48555]_  = \new_[48554]_  & \new_[48547]_ ;
  assign \new_[48558]_  = ~A267 & A235;
  assign \new_[48561]_  = A298 & A268;
  assign \new_[48562]_  = \new_[48561]_  & \new_[48558]_ ;
  assign \new_[48565]_  = ~A300 & ~A299;
  assign \new_[48568]_  = A302 & ~A301;
  assign \new_[48569]_  = \new_[48568]_  & \new_[48565]_ ;
  assign \new_[48570]_  = \new_[48569]_  & \new_[48562]_ ;
  assign \new_[48573]_  = A200 & ~A199;
  assign \new_[48576]_  = ~A202 & ~A201;
  assign \new_[48577]_  = \new_[48576]_  & \new_[48573]_ ;
  assign \new_[48580]_  = A232 & A203;
  assign \new_[48583]_  = A234 & ~A233;
  assign \new_[48584]_  = \new_[48583]_  & \new_[48580]_ ;
  assign \new_[48585]_  = \new_[48584]_  & \new_[48577]_ ;
  assign \new_[48588]_  = ~A267 & A235;
  assign \new_[48591]_  = ~A298 & A268;
  assign \new_[48592]_  = \new_[48591]_  & \new_[48588]_ ;
  assign \new_[48595]_  = ~A300 & A299;
  assign \new_[48598]_  = A302 & ~A301;
  assign \new_[48599]_  = \new_[48598]_  & \new_[48595]_ ;
  assign \new_[48600]_  = \new_[48599]_  & \new_[48592]_ ;
  assign \new_[48603]_  = A200 & ~A199;
  assign \new_[48606]_  = ~A202 & ~A201;
  assign \new_[48607]_  = \new_[48606]_  & \new_[48603]_ ;
  assign \new_[48610]_  = A232 & A203;
  assign \new_[48613]_  = A234 & ~A233;
  assign \new_[48614]_  = \new_[48613]_  & \new_[48610]_ ;
  assign \new_[48615]_  = \new_[48614]_  & \new_[48607]_ ;
  assign \new_[48618]_  = ~A267 & A235;
  assign \new_[48621]_  = A298 & ~A269;
  assign \new_[48622]_  = \new_[48621]_  & \new_[48618]_ ;
  assign \new_[48625]_  = ~A300 & ~A299;
  assign \new_[48628]_  = A302 & ~A301;
  assign \new_[48629]_  = \new_[48628]_  & \new_[48625]_ ;
  assign \new_[48630]_  = \new_[48629]_  & \new_[48622]_ ;
  assign \new_[48633]_  = A200 & ~A199;
  assign \new_[48636]_  = ~A202 & ~A201;
  assign \new_[48637]_  = \new_[48636]_  & \new_[48633]_ ;
  assign \new_[48640]_  = A232 & A203;
  assign \new_[48643]_  = A234 & ~A233;
  assign \new_[48644]_  = \new_[48643]_  & \new_[48640]_ ;
  assign \new_[48645]_  = \new_[48644]_  & \new_[48637]_ ;
  assign \new_[48648]_  = ~A267 & A235;
  assign \new_[48651]_  = ~A298 & ~A269;
  assign \new_[48652]_  = \new_[48651]_  & \new_[48648]_ ;
  assign \new_[48655]_  = ~A300 & A299;
  assign \new_[48658]_  = A302 & ~A301;
  assign \new_[48659]_  = \new_[48658]_  & \new_[48655]_ ;
  assign \new_[48660]_  = \new_[48659]_  & \new_[48652]_ ;
  assign \new_[48663]_  = A200 & ~A199;
  assign \new_[48666]_  = ~A202 & ~A201;
  assign \new_[48667]_  = \new_[48666]_  & \new_[48663]_ ;
  assign \new_[48670]_  = A232 & A203;
  assign \new_[48673]_  = A234 & ~A233;
  assign \new_[48674]_  = \new_[48673]_  & \new_[48670]_ ;
  assign \new_[48675]_  = \new_[48674]_  & \new_[48667]_ ;
  assign \new_[48678]_  = A265 & A235;
  assign \new_[48681]_  = A298 & A266;
  assign \new_[48682]_  = \new_[48681]_  & \new_[48678]_ ;
  assign \new_[48685]_  = ~A300 & ~A299;
  assign \new_[48688]_  = A302 & ~A301;
  assign \new_[48689]_  = \new_[48688]_  & \new_[48685]_ ;
  assign \new_[48690]_  = \new_[48689]_  & \new_[48682]_ ;
  assign \new_[48693]_  = A200 & ~A199;
  assign \new_[48696]_  = ~A202 & ~A201;
  assign \new_[48697]_  = \new_[48696]_  & \new_[48693]_ ;
  assign \new_[48700]_  = A232 & A203;
  assign \new_[48703]_  = A234 & ~A233;
  assign \new_[48704]_  = \new_[48703]_  & \new_[48700]_ ;
  assign \new_[48705]_  = \new_[48704]_  & \new_[48697]_ ;
  assign \new_[48708]_  = A265 & A235;
  assign \new_[48711]_  = ~A298 & A266;
  assign \new_[48712]_  = \new_[48711]_  & \new_[48708]_ ;
  assign \new_[48715]_  = ~A300 & A299;
  assign \new_[48718]_  = A302 & ~A301;
  assign \new_[48719]_  = \new_[48718]_  & \new_[48715]_ ;
  assign \new_[48720]_  = \new_[48719]_  & \new_[48712]_ ;
  assign \new_[48723]_  = A200 & ~A199;
  assign \new_[48726]_  = ~A202 & ~A201;
  assign \new_[48727]_  = \new_[48726]_  & \new_[48723]_ ;
  assign \new_[48730]_  = A232 & A203;
  assign \new_[48733]_  = A234 & ~A233;
  assign \new_[48734]_  = \new_[48733]_  & \new_[48730]_ ;
  assign \new_[48735]_  = \new_[48734]_  & \new_[48727]_ ;
  assign \new_[48738]_  = ~A265 & A235;
  assign \new_[48741]_  = A298 & ~A266;
  assign \new_[48742]_  = \new_[48741]_  & \new_[48738]_ ;
  assign \new_[48745]_  = ~A300 & ~A299;
  assign \new_[48748]_  = A302 & ~A301;
  assign \new_[48749]_  = \new_[48748]_  & \new_[48745]_ ;
  assign \new_[48750]_  = \new_[48749]_  & \new_[48742]_ ;
  assign \new_[48753]_  = A200 & ~A199;
  assign \new_[48756]_  = ~A202 & ~A201;
  assign \new_[48757]_  = \new_[48756]_  & \new_[48753]_ ;
  assign \new_[48760]_  = A232 & A203;
  assign \new_[48763]_  = A234 & ~A233;
  assign \new_[48764]_  = \new_[48763]_  & \new_[48760]_ ;
  assign \new_[48765]_  = \new_[48764]_  & \new_[48757]_ ;
  assign \new_[48768]_  = ~A265 & A235;
  assign \new_[48771]_  = ~A298 & ~A266;
  assign \new_[48772]_  = \new_[48771]_  & \new_[48768]_ ;
  assign \new_[48775]_  = ~A300 & A299;
  assign \new_[48778]_  = A302 & ~A301;
  assign \new_[48779]_  = \new_[48778]_  & \new_[48775]_ ;
  assign \new_[48780]_  = \new_[48779]_  & \new_[48772]_ ;
  assign \new_[48783]_  = A200 & ~A199;
  assign \new_[48786]_  = ~A202 & ~A201;
  assign \new_[48787]_  = \new_[48786]_  & \new_[48783]_ ;
  assign \new_[48790]_  = A232 & A203;
  assign \new_[48793]_  = A234 & ~A233;
  assign \new_[48794]_  = \new_[48793]_  & \new_[48790]_ ;
  assign \new_[48795]_  = \new_[48794]_  & \new_[48787]_ ;
  assign \new_[48798]_  = A267 & ~A236;
  assign \new_[48801]_  = A269 & ~A268;
  assign \new_[48802]_  = \new_[48801]_  & \new_[48798]_ ;
  assign \new_[48805]_  = ~A299 & A298;
  assign \new_[48808]_  = A301 & A300;
  assign \new_[48809]_  = \new_[48808]_  & \new_[48805]_ ;
  assign \new_[48810]_  = \new_[48809]_  & \new_[48802]_ ;
  assign \new_[48813]_  = A200 & ~A199;
  assign \new_[48816]_  = ~A202 & ~A201;
  assign \new_[48817]_  = \new_[48816]_  & \new_[48813]_ ;
  assign \new_[48820]_  = A232 & A203;
  assign \new_[48823]_  = A234 & ~A233;
  assign \new_[48824]_  = \new_[48823]_  & \new_[48820]_ ;
  assign \new_[48825]_  = \new_[48824]_  & \new_[48817]_ ;
  assign \new_[48828]_  = A267 & ~A236;
  assign \new_[48831]_  = A269 & ~A268;
  assign \new_[48832]_  = \new_[48831]_  & \new_[48828]_ ;
  assign \new_[48835]_  = ~A299 & A298;
  assign \new_[48838]_  = ~A302 & A300;
  assign \new_[48839]_  = \new_[48838]_  & \new_[48835]_ ;
  assign \new_[48840]_  = \new_[48839]_  & \new_[48832]_ ;
  assign \new_[48843]_  = A200 & ~A199;
  assign \new_[48846]_  = ~A202 & ~A201;
  assign \new_[48847]_  = \new_[48846]_  & \new_[48843]_ ;
  assign \new_[48850]_  = A232 & A203;
  assign \new_[48853]_  = A234 & ~A233;
  assign \new_[48854]_  = \new_[48853]_  & \new_[48850]_ ;
  assign \new_[48855]_  = \new_[48854]_  & \new_[48847]_ ;
  assign \new_[48858]_  = A267 & ~A236;
  assign \new_[48861]_  = A269 & ~A268;
  assign \new_[48862]_  = \new_[48861]_  & \new_[48858]_ ;
  assign \new_[48865]_  = A299 & ~A298;
  assign \new_[48868]_  = A301 & A300;
  assign \new_[48869]_  = \new_[48868]_  & \new_[48865]_ ;
  assign \new_[48870]_  = \new_[48869]_  & \new_[48862]_ ;
  assign \new_[48873]_  = A200 & ~A199;
  assign \new_[48876]_  = ~A202 & ~A201;
  assign \new_[48877]_  = \new_[48876]_  & \new_[48873]_ ;
  assign \new_[48880]_  = A232 & A203;
  assign \new_[48883]_  = A234 & ~A233;
  assign \new_[48884]_  = \new_[48883]_  & \new_[48880]_ ;
  assign \new_[48885]_  = \new_[48884]_  & \new_[48877]_ ;
  assign \new_[48888]_  = A267 & ~A236;
  assign \new_[48891]_  = A269 & ~A268;
  assign \new_[48892]_  = \new_[48891]_  & \new_[48888]_ ;
  assign \new_[48895]_  = A299 & ~A298;
  assign \new_[48898]_  = ~A302 & A300;
  assign \new_[48899]_  = \new_[48898]_  & \new_[48895]_ ;
  assign \new_[48900]_  = \new_[48899]_  & \new_[48892]_ ;
  assign \new_[48903]_  = A200 & ~A199;
  assign \new_[48906]_  = ~A202 & ~A201;
  assign \new_[48907]_  = \new_[48906]_  & \new_[48903]_ ;
  assign \new_[48910]_  = A232 & A203;
  assign \new_[48913]_  = A234 & ~A233;
  assign \new_[48914]_  = \new_[48913]_  & \new_[48910]_ ;
  assign \new_[48915]_  = \new_[48914]_  & \new_[48907]_ ;
  assign \new_[48918]_  = ~A267 & ~A236;
  assign \new_[48921]_  = A298 & A268;
  assign \new_[48922]_  = \new_[48921]_  & \new_[48918]_ ;
  assign \new_[48925]_  = ~A300 & ~A299;
  assign \new_[48928]_  = A302 & ~A301;
  assign \new_[48929]_  = \new_[48928]_  & \new_[48925]_ ;
  assign \new_[48930]_  = \new_[48929]_  & \new_[48922]_ ;
  assign \new_[48933]_  = A200 & ~A199;
  assign \new_[48936]_  = ~A202 & ~A201;
  assign \new_[48937]_  = \new_[48936]_  & \new_[48933]_ ;
  assign \new_[48940]_  = A232 & A203;
  assign \new_[48943]_  = A234 & ~A233;
  assign \new_[48944]_  = \new_[48943]_  & \new_[48940]_ ;
  assign \new_[48945]_  = \new_[48944]_  & \new_[48937]_ ;
  assign \new_[48948]_  = ~A267 & ~A236;
  assign \new_[48951]_  = ~A298 & A268;
  assign \new_[48952]_  = \new_[48951]_  & \new_[48948]_ ;
  assign \new_[48955]_  = ~A300 & A299;
  assign \new_[48958]_  = A302 & ~A301;
  assign \new_[48959]_  = \new_[48958]_  & \new_[48955]_ ;
  assign \new_[48960]_  = \new_[48959]_  & \new_[48952]_ ;
  assign \new_[48963]_  = A200 & ~A199;
  assign \new_[48966]_  = ~A202 & ~A201;
  assign \new_[48967]_  = \new_[48966]_  & \new_[48963]_ ;
  assign \new_[48970]_  = A232 & A203;
  assign \new_[48973]_  = A234 & ~A233;
  assign \new_[48974]_  = \new_[48973]_  & \new_[48970]_ ;
  assign \new_[48975]_  = \new_[48974]_  & \new_[48967]_ ;
  assign \new_[48978]_  = ~A267 & ~A236;
  assign \new_[48981]_  = A298 & ~A269;
  assign \new_[48982]_  = \new_[48981]_  & \new_[48978]_ ;
  assign \new_[48985]_  = ~A300 & ~A299;
  assign \new_[48988]_  = A302 & ~A301;
  assign \new_[48989]_  = \new_[48988]_  & \new_[48985]_ ;
  assign \new_[48990]_  = \new_[48989]_  & \new_[48982]_ ;
  assign \new_[48993]_  = A200 & ~A199;
  assign \new_[48996]_  = ~A202 & ~A201;
  assign \new_[48997]_  = \new_[48996]_  & \new_[48993]_ ;
  assign \new_[49000]_  = A232 & A203;
  assign \new_[49003]_  = A234 & ~A233;
  assign \new_[49004]_  = \new_[49003]_  & \new_[49000]_ ;
  assign \new_[49005]_  = \new_[49004]_  & \new_[48997]_ ;
  assign \new_[49008]_  = ~A267 & ~A236;
  assign \new_[49011]_  = ~A298 & ~A269;
  assign \new_[49012]_  = \new_[49011]_  & \new_[49008]_ ;
  assign \new_[49015]_  = ~A300 & A299;
  assign \new_[49018]_  = A302 & ~A301;
  assign \new_[49019]_  = \new_[49018]_  & \new_[49015]_ ;
  assign \new_[49020]_  = \new_[49019]_  & \new_[49012]_ ;
  assign \new_[49023]_  = A200 & ~A199;
  assign \new_[49026]_  = ~A202 & ~A201;
  assign \new_[49027]_  = \new_[49026]_  & \new_[49023]_ ;
  assign \new_[49030]_  = A232 & A203;
  assign \new_[49033]_  = A234 & ~A233;
  assign \new_[49034]_  = \new_[49033]_  & \new_[49030]_ ;
  assign \new_[49035]_  = \new_[49034]_  & \new_[49027]_ ;
  assign \new_[49038]_  = A265 & ~A236;
  assign \new_[49041]_  = A298 & A266;
  assign \new_[49042]_  = \new_[49041]_  & \new_[49038]_ ;
  assign \new_[49045]_  = ~A300 & ~A299;
  assign \new_[49048]_  = A302 & ~A301;
  assign \new_[49049]_  = \new_[49048]_  & \new_[49045]_ ;
  assign \new_[49050]_  = \new_[49049]_  & \new_[49042]_ ;
  assign \new_[49053]_  = A200 & ~A199;
  assign \new_[49056]_  = ~A202 & ~A201;
  assign \new_[49057]_  = \new_[49056]_  & \new_[49053]_ ;
  assign \new_[49060]_  = A232 & A203;
  assign \new_[49063]_  = A234 & ~A233;
  assign \new_[49064]_  = \new_[49063]_  & \new_[49060]_ ;
  assign \new_[49065]_  = \new_[49064]_  & \new_[49057]_ ;
  assign \new_[49068]_  = A265 & ~A236;
  assign \new_[49071]_  = ~A298 & A266;
  assign \new_[49072]_  = \new_[49071]_  & \new_[49068]_ ;
  assign \new_[49075]_  = ~A300 & A299;
  assign \new_[49078]_  = A302 & ~A301;
  assign \new_[49079]_  = \new_[49078]_  & \new_[49075]_ ;
  assign \new_[49080]_  = \new_[49079]_  & \new_[49072]_ ;
  assign \new_[49083]_  = A200 & ~A199;
  assign \new_[49086]_  = ~A202 & ~A201;
  assign \new_[49087]_  = \new_[49086]_  & \new_[49083]_ ;
  assign \new_[49090]_  = A232 & A203;
  assign \new_[49093]_  = A234 & ~A233;
  assign \new_[49094]_  = \new_[49093]_  & \new_[49090]_ ;
  assign \new_[49095]_  = \new_[49094]_  & \new_[49087]_ ;
  assign \new_[49098]_  = ~A265 & ~A236;
  assign \new_[49101]_  = A298 & ~A266;
  assign \new_[49102]_  = \new_[49101]_  & \new_[49098]_ ;
  assign \new_[49105]_  = ~A300 & ~A299;
  assign \new_[49108]_  = A302 & ~A301;
  assign \new_[49109]_  = \new_[49108]_  & \new_[49105]_ ;
  assign \new_[49110]_  = \new_[49109]_  & \new_[49102]_ ;
  assign \new_[49113]_  = A200 & ~A199;
  assign \new_[49116]_  = ~A202 & ~A201;
  assign \new_[49117]_  = \new_[49116]_  & \new_[49113]_ ;
  assign \new_[49120]_  = A232 & A203;
  assign \new_[49123]_  = A234 & ~A233;
  assign \new_[49124]_  = \new_[49123]_  & \new_[49120]_ ;
  assign \new_[49125]_  = \new_[49124]_  & \new_[49117]_ ;
  assign \new_[49128]_  = ~A265 & ~A236;
  assign \new_[49131]_  = ~A298 & ~A266;
  assign \new_[49132]_  = \new_[49131]_  & \new_[49128]_ ;
  assign \new_[49135]_  = ~A300 & A299;
  assign \new_[49138]_  = A302 & ~A301;
  assign \new_[49139]_  = \new_[49138]_  & \new_[49135]_ ;
  assign \new_[49140]_  = \new_[49139]_  & \new_[49132]_ ;
  assign \new_[49143]_  = A200 & ~A199;
  assign \new_[49146]_  = ~A202 & ~A201;
  assign \new_[49147]_  = \new_[49146]_  & \new_[49143]_ ;
  assign \new_[49150]_  = A232 & A203;
  assign \new_[49153]_  = ~A234 & ~A233;
  assign \new_[49154]_  = \new_[49153]_  & \new_[49150]_ ;
  assign \new_[49155]_  = \new_[49154]_  & \new_[49147]_ ;
  assign \new_[49158]_  = A236 & ~A235;
  assign \new_[49161]_  = A268 & ~A267;
  assign \new_[49162]_  = \new_[49161]_  & \new_[49158]_ ;
  assign \new_[49165]_  = ~A299 & A298;
  assign \new_[49168]_  = A301 & A300;
  assign \new_[49169]_  = \new_[49168]_  & \new_[49165]_ ;
  assign \new_[49170]_  = \new_[49169]_  & \new_[49162]_ ;
  assign \new_[49173]_  = A200 & ~A199;
  assign \new_[49176]_  = ~A202 & ~A201;
  assign \new_[49177]_  = \new_[49176]_  & \new_[49173]_ ;
  assign \new_[49180]_  = A232 & A203;
  assign \new_[49183]_  = ~A234 & ~A233;
  assign \new_[49184]_  = \new_[49183]_  & \new_[49180]_ ;
  assign \new_[49185]_  = \new_[49184]_  & \new_[49177]_ ;
  assign \new_[49188]_  = A236 & ~A235;
  assign \new_[49191]_  = A268 & ~A267;
  assign \new_[49192]_  = \new_[49191]_  & \new_[49188]_ ;
  assign \new_[49195]_  = ~A299 & A298;
  assign \new_[49198]_  = ~A302 & A300;
  assign \new_[49199]_  = \new_[49198]_  & \new_[49195]_ ;
  assign \new_[49200]_  = \new_[49199]_  & \new_[49192]_ ;
  assign \new_[49203]_  = A200 & ~A199;
  assign \new_[49206]_  = ~A202 & ~A201;
  assign \new_[49207]_  = \new_[49206]_  & \new_[49203]_ ;
  assign \new_[49210]_  = A232 & A203;
  assign \new_[49213]_  = ~A234 & ~A233;
  assign \new_[49214]_  = \new_[49213]_  & \new_[49210]_ ;
  assign \new_[49215]_  = \new_[49214]_  & \new_[49207]_ ;
  assign \new_[49218]_  = A236 & ~A235;
  assign \new_[49221]_  = A268 & ~A267;
  assign \new_[49222]_  = \new_[49221]_  & \new_[49218]_ ;
  assign \new_[49225]_  = A299 & ~A298;
  assign \new_[49228]_  = A301 & A300;
  assign \new_[49229]_  = \new_[49228]_  & \new_[49225]_ ;
  assign \new_[49230]_  = \new_[49229]_  & \new_[49222]_ ;
  assign \new_[49233]_  = A200 & ~A199;
  assign \new_[49236]_  = ~A202 & ~A201;
  assign \new_[49237]_  = \new_[49236]_  & \new_[49233]_ ;
  assign \new_[49240]_  = A232 & A203;
  assign \new_[49243]_  = ~A234 & ~A233;
  assign \new_[49244]_  = \new_[49243]_  & \new_[49240]_ ;
  assign \new_[49245]_  = \new_[49244]_  & \new_[49237]_ ;
  assign \new_[49248]_  = A236 & ~A235;
  assign \new_[49251]_  = A268 & ~A267;
  assign \new_[49252]_  = \new_[49251]_  & \new_[49248]_ ;
  assign \new_[49255]_  = A299 & ~A298;
  assign \new_[49258]_  = ~A302 & A300;
  assign \new_[49259]_  = \new_[49258]_  & \new_[49255]_ ;
  assign \new_[49260]_  = \new_[49259]_  & \new_[49252]_ ;
  assign \new_[49263]_  = A200 & ~A199;
  assign \new_[49266]_  = ~A202 & ~A201;
  assign \new_[49267]_  = \new_[49266]_  & \new_[49263]_ ;
  assign \new_[49270]_  = A232 & A203;
  assign \new_[49273]_  = ~A234 & ~A233;
  assign \new_[49274]_  = \new_[49273]_  & \new_[49270]_ ;
  assign \new_[49275]_  = \new_[49274]_  & \new_[49267]_ ;
  assign \new_[49278]_  = A236 & ~A235;
  assign \new_[49281]_  = ~A269 & ~A267;
  assign \new_[49282]_  = \new_[49281]_  & \new_[49278]_ ;
  assign \new_[49285]_  = ~A299 & A298;
  assign \new_[49288]_  = A301 & A300;
  assign \new_[49289]_  = \new_[49288]_  & \new_[49285]_ ;
  assign \new_[49290]_  = \new_[49289]_  & \new_[49282]_ ;
  assign \new_[49293]_  = A200 & ~A199;
  assign \new_[49296]_  = ~A202 & ~A201;
  assign \new_[49297]_  = \new_[49296]_  & \new_[49293]_ ;
  assign \new_[49300]_  = A232 & A203;
  assign \new_[49303]_  = ~A234 & ~A233;
  assign \new_[49304]_  = \new_[49303]_  & \new_[49300]_ ;
  assign \new_[49305]_  = \new_[49304]_  & \new_[49297]_ ;
  assign \new_[49308]_  = A236 & ~A235;
  assign \new_[49311]_  = ~A269 & ~A267;
  assign \new_[49312]_  = \new_[49311]_  & \new_[49308]_ ;
  assign \new_[49315]_  = ~A299 & A298;
  assign \new_[49318]_  = ~A302 & A300;
  assign \new_[49319]_  = \new_[49318]_  & \new_[49315]_ ;
  assign \new_[49320]_  = \new_[49319]_  & \new_[49312]_ ;
  assign \new_[49323]_  = A200 & ~A199;
  assign \new_[49326]_  = ~A202 & ~A201;
  assign \new_[49327]_  = \new_[49326]_  & \new_[49323]_ ;
  assign \new_[49330]_  = A232 & A203;
  assign \new_[49333]_  = ~A234 & ~A233;
  assign \new_[49334]_  = \new_[49333]_  & \new_[49330]_ ;
  assign \new_[49335]_  = \new_[49334]_  & \new_[49327]_ ;
  assign \new_[49338]_  = A236 & ~A235;
  assign \new_[49341]_  = ~A269 & ~A267;
  assign \new_[49342]_  = \new_[49341]_  & \new_[49338]_ ;
  assign \new_[49345]_  = A299 & ~A298;
  assign \new_[49348]_  = A301 & A300;
  assign \new_[49349]_  = \new_[49348]_  & \new_[49345]_ ;
  assign \new_[49350]_  = \new_[49349]_  & \new_[49342]_ ;
  assign \new_[49353]_  = A200 & ~A199;
  assign \new_[49356]_  = ~A202 & ~A201;
  assign \new_[49357]_  = \new_[49356]_  & \new_[49353]_ ;
  assign \new_[49360]_  = A232 & A203;
  assign \new_[49363]_  = ~A234 & ~A233;
  assign \new_[49364]_  = \new_[49363]_  & \new_[49360]_ ;
  assign \new_[49365]_  = \new_[49364]_  & \new_[49357]_ ;
  assign \new_[49368]_  = A236 & ~A235;
  assign \new_[49371]_  = ~A269 & ~A267;
  assign \new_[49372]_  = \new_[49371]_  & \new_[49368]_ ;
  assign \new_[49375]_  = A299 & ~A298;
  assign \new_[49378]_  = ~A302 & A300;
  assign \new_[49379]_  = \new_[49378]_  & \new_[49375]_ ;
  assign \new_[49380]_  = \new_[49379]_  & \new_[49372]_ ;
  assign \new_[49383]_  = A200 & ~A199;
  assign \new_[49386]_  = ~A202 & ~A201;
  assign \new_[49387]_  = \new_[49386]_  & \new_[49383]_ ;
  assign \new_[49390]_  = A232 & A203;
  assign \new_[49393]_  = ~A234 & ~A233;
  assign \new_[49394]_  = \new_[49393]_  & \new_[49390]_ ;
  assign \new_[49395]_  = \new_[49394]_  & \new_[49387]_ ;
  assign \new_[49398]_  = A236 & ~A235;
  assign \new_[49401]_  = A266 & A265;
  assign \new_[49402]_  = \new_[49401]_  & \new_[49398]_ ;
  assign \new_[49405]_  = ~A299 & A298;
  assign \new_[49408]_  = A301 & A300;
  assign \new_[49409]_  = \new_[49408]_  & \new_[49405]_ ;
  assign \new_[49410]_  = \new_[49409]_  & \new_[49402]_ ;
  assign \new_[49413]_  = A200 & ~A199;
  assign \new_[49416]_  = ~A202 & ~A201;
  assign \new_[49417]_  = \new_[49416]_  & \new_[49413]_ ;
  assign \new_[49420]_  = A232 & A203;
  assign \new_[49423]_  = ~A234 & ~A233;
  assign \new_[49424]_  = \new_[49423]_  & \new_[49420]_ ;
  assign \new_[49425]_  = \new_[49424]_  & \new_[49417]_ ;
  assign \new_[49428]_  = A236 & ~A235;
  assign \new_[49431]_  = A266 & A265;
  assign \new_[49432]_  = \new_[49431]_  & \new_[49428]_ ;
  assign \new_[49435]_  = ~A299 & A298;
  assign \new_[49438]_  = ~A302 & A300;
  assign \new_[49439]_  = \new_[49438]_  & \new_[49435]_ ;
  assign \new_[49440]_  = \new_[49439]_  & \new_[49432]_ ;
  assign \new_[49443]_  = A200 & ~A199;
  assign \new_[49446]_  = ~A202 & ~A201;
  assign \new_[49447]_  = \new_[49446]_  & \new_[49443]_ ;
  assign \new_[49450]_  = A232 & A203;
  assign \new_[49453]_  = ~A234 & ~A233;
  assign \new_[49454]_  = \new_[49453]_  & \new_[49450]_ ;
  assign \new_[49455]_  = \new_[49454]_  & \new_[49447]_ ;
  assign \new_[49458]_  = A236 & ~A235;
  assign \new_[49461]_  = A266 & A265;
  assign \new_[49462]_  = \new_[49461]_  & \new_[49458]_ ;
  assign \new_[49465]_  = A299 & ~A298;
  assign \new_[49468]_  = A301 & A300;
  assign \new_[49469]_  = \new_[49468]_  & \new_[49465]_ ;
  assign \new_[49470]_  = \new_[49469]_  & \new_[49462]_ ;
  assign \new_[49473]_  = A200 & ~A199;
  assign \new_[49476]_  = ~A202 & ~A201;
  assign \new_[49477]_  = \new_[49476]_  & \new_[49473]_ ;
  assign \new_[49480]_  = A232 & A203;
  assign \new_[49483]_  = ~A234 & ~A233;
  assign \new_[49484]_  = \new_[49483]_  & \new_[49480]_ ;
  assign \new_[49485]_  = \new_[49484]_  & \new_[49477]_ ;
  assign \new_[49488]_  = A236 & ~A235;
  assign \new_[49491]_  = A266 & A265;
  assign \new_[49492]_  = \new_[49491]_  & \new_[49488]_ ;
  assign \new_[49495]_  = A299 & ~A298;
  assign \new_[49498]_  = ~A302 & A300;
  assign \new_[49499]_  = \new_[49498]_  & \new_[49495]_ ;
  assign \new_[49500]_  = \new_[49499]_  & \new_[49492]_ ;
  assign \new_[49503]_  = A200 & ~A199;
  assign \new_[49506]_  = ~A202 & ~A201;
  assign \new_[49507]_  = \new_[49506]_  & \new_[49503]_ ;
  assign \new_[49510]_  = A232 & A203;
  assign \new_[49513]_  = ~A234 & ~A233;
  assign \new_[49514]_  = \new_[49513]_  & \new_[49510]_ ;
  assign \new_[49515]_  = \new_[49514]_  & \new_[49507]_ ;
  assign \new_[49518]_  = A236 & ~A235;
  assign \new_[49521]_  = ~A266 & ~A265;
  assign \new_[49522]_  = \new_[49521]_  & \new_[49518]_ ;
  assign \new_[49525]_  = ~A299 & A298;
  assign \new_[49528]_  = A301 & A300;
  assign \new_[49529]_  = \new_[49528]_  & \new_[49525]_ ;
  assign \new_[49530]_  = \new_[49529]_  & \new_[49522]_ ;
  assign \new_[49533]_  = A200 & ~A199;
  assign \new_[49536]_  = ~A202 & ~A201;
  assign \new_[49537]_  = \new_[49536]_  & \new_[49533]_ ;
  assign \new_[49540]_  = A232 & A203;
  assign \new_[49543]_  = ~A234 & ~A233;
  assign \new_[49544]_  = \new_[49543]_  & \new_[49540]_ ;
  assign \new_[49545]_  = \new_[49544]_  & \new_[49537]_ ;
  assign \new_[49548]_  = A236 & ~A235;
  assign \new_[49551]_  = ~A266 & ~A265;
  assign \new_[49552]_  = \new_[49551]_  & \new_[49548]_ ;
  assign \new_[49555]_  = ~A299 & A298;
  assign \new_[49558]_  = ~A302 & A300;
  assign \new_[49559]_  = \new_[49558]_  & \new_[49555]_ ;
  assign \new_[49560]_  = \new_[49559]_  & \new_[49552]_ ;
  assign \new_[49563]_  = A200 & ~A199;
  assign \new_[49566]_  = ~A202 & ~A201;
  assign \new_[49567]_  = \new_[49566]_  & \new_[49563]_ ;
  assign \new_[49570]_  = A232 & A203;
  assign \new_[49573]_  = ~A234 & ~A233;
  assign \new_[49574]_  = \new_[49573]_  & \new_[49570]_ ;
  assign \new_[49575]_  = \new_[49574]_  & \new_[49567]_ ;
  assign \new_[49578]_  = A236 & ~A235;
  assign \new_[49581]_  = ~A266 & ~A265;
  assign \new_[49582]_  = \new_[49581]_  & \new_[49578]_ ;
  assign \new_[49585]_  = A299 & ~A298;
  assign \new_[49588]_  = A301 & A300;
  assign \new_[49589]_  = \new_[49588]_  & \new_[49585]_ ;
  assign \new_[49590]_  = \new_[49589]_  & \new_[49582]_ ;
  assign \new_[49593]_  = A200 & ~A199;
  assign \new_[49596]_  = ~A202 & ~A201;
  assign \new_[49597]_  = \new_[49596]_  & \new_[49593]_ ;
  assign \new_[49600]_  = A232 & A203;
  assign \new_[49603]_  = ~A234 & ~A233;
  assign \new_[49604]_  = \new_[49603]_  & \new_[49600]_ ;
  assign \new_[49605]_  = \new_[49604]_  & \new_[49597]_ ;
  assign \new_[49608]_  = A236 & ~A235;
  assign \new_[49611]_  = ~A266 & ~A265;
  assign \new_[49612]_  = \new_[49611]_  & \new_[49608]_ ;
  assign \new_[49615]_  = A299 & ~A298;
  assign \new_[49618]_  = ~A302 & A300;
  assign \new_[49619]_  = \new_[49618]_  & \new_[49615]_ ;
  assign \new_[49620]_  = \new_[49619]_  & \new_[49612]_ ;
  assign \new_[49623]_  = ~A200 & A199;
  assign \new_[49626]_  = A202 & A201;
  assign \new_[49627]_  = \new_[49626]_  & \new_[49623]_ ;
  assign \new_[49630]_  = A233 & ~A232;
  assign \new_[49633]_  = A235 & A234;
  assign \new_[49634]_  = \new_[49633]_  & \new_[49630]_ ;
  assign \new_[49635]_  = \new_[49634]_  & \new_[49627]_ ;
  assign \new_[49638]_  = ~A268 & A267;
  assign \new_[49641]_  = A298 & A269;
  assign \new_[49642]_  = \new_[49641]_  & \new_[49638]_ ;
  assign \new_[49645]_  = ~A300 & ~A299;
  assign \new_[49648]_  = A302 & ~A301;
  assign \new_[49649]_  = \new_[49648]_  & \new_[49645]_ ;
  assign \new_[49650]_  = \new_[49649]_  & \new_[49642]_ ;
  assign \new_[49653]_  = ~A200 & A199;
  assign \new_[49656]_  = A202 & A201;
  assign \new_[49657]_  = \new_[49656]_  & \new_[49653]_ ;
  assign \new_[49660]_  = A233 & ~A232;
  assign \new_[49663]_  = A235 & A234;
  assign \new_[49664]_  = \new_[49663]_  & \new_[49660]_ ;
  assign \new_[49665]_  = \new_[49664]_  & \new_[49657]_ ;
  assign \new_[49668]_  = ~A268 & A267;
  assign \new_[49671]_  = ~A298 & A269;
  assign \new_[49672]_  = \new_[49671]_  & \new_[49668]_ ;
  assign \new_[49675]_  = ~A300 & A299;
  assign \new_[49678]_  = A302 & ~A301;
  assign \new_[49679]_  = \new_[49678]_  & \new_[49675]_ ;
  assign \new_[49680]_  = \new_[49679]_  & \new_[49672]_ ;
  assign \new_[49683]_  = ~A200 & A199;
  assign \new_[49686]_  = A202 & A201;
  assign \new_[49687]_  = \new_[49686]_  & \new_[49683]_ ;
  assign \new_[49690]_  = A233 & ~A232;
  assign \new_[49693]_  = ~A236 & A234;
  assign \new_[49694]_  = \new_[49693]_  & \new_[49690]_ ;
  assign \new_[49695]_  = \new_[49694]_  & \new_[49687]_ ;
  assign \new_[49698]_  = ~A268 & A267;
  assign \new_[49701]_  = A298 & A269;
  assign \new_[49702]_  = \new_[49701]_  & \new_[49698]_ ;
  assign \new_[49705]_  = ~A300 & ~A299;
  assign \new_[49708]_  = A302 & ~A301;
  assign \new_[49709]_  = \new_[49708]_  & \new_[49705]_ ;
  assign \new_[49710]_  = \new_[49709]_  & \new_[49702]_ ;
  assign \new_[49713]_  = ~A200 & A199;
  assign \new_[49716]_  = A202 & A201;
  assign \new_[49717]_  = \new_[49716]_  & \new_[49713]_ ;
  assign \new_[49720]_  = A233 & ~A232;
  assign \new_[49723]_  = ~A236 & A234;
  assign \new_[49724]_  = \new_[49723]_  & \new_[49720]_ ;
  assign \new_[49725]_  = \new_[49724]_  & \new_[49717]_ ;
  assign \new_[49728]_  = ~A268 & A267;
  assign \new_[49731]_  = ~A298 & A269;
  assign \new_[49732]_  = \new_[49731]_  & \new_[49728]_ ;
  assign \new_[49735]_  = ~A300 & A299;
  assign \new_[49738]_  = A302 & ~A301;
  assign \new_[49739]_  = \new_[49738]_  & \new_[49735]_ ;
  assign \new_[49740]_  = \new_[49739]_  & \new_[49732]_ ;
  assign \new_[49743]_  = ~A200 & A199;
  assign \new_[49746]_  = A202 & A201;
  assign \new_[49747]_  = \new_[49746]_  & \new_[49743]_ ;
  assign \new_[49750]_  = A233 & ~A232;
  assign \new_[49753]_  = ~A235 & ~A234;
  assign \new_[49754]_  = \new_[49753]_  & \new_[49750]_ ;
  assign \new_[49755]_  = \new_[49754]_  & \new_[49747]_ ;
  assign \new_[49758]_  = A267 & A236;
  assign \new_[49761]_  = A269 & ~A268;
  assign \new_[49762]_  = \new_[49761]_  & \new_[49758]_ ;
  assign \new_[49765]_  = ~A299 & A298;
  assign \new_[49768]_  = A301 & A300;
  assign \new_[49769]_  = \new_[49768]_  & \new_[49765]_ ;
  assign \new_[49770]_  = \new_[49769]_  & \new_[49762]_ ;
  assign \new_[49773]_  = ~A200 & A199;
  assign \new_[49776]_  = A202 & A201;
  assign \new_[49777]_  = \new_[49776]_  & \new_[49773]_ ;
  assign \new_[49780]_  = A233 & ~A232;
  assign \new_[49783]_  = ~A235 & ~A234;
  assign \new_[49784]_  = \new_[49783]_  & \new_[49780]_ ;
  assign \new_[49785]_  = \new_[49784]_  & \new_[49777]_ ;
  assign \new_[49788]_  = A267 & A236;
  assign \new_[49791]_  = A269 & ~A268;
  assign \new_[49792]_  = \new_[49791]_  & \new_[49788]_ ;
  assign \new_[49795]_  = ~A299 & A298;
  assign \new_[49798]_  = ~A302 & A300;
  assign \new_[49799]_  = \new_[49798]_  & \new_[49795]_ ;
  assign \new_[49800]_  = \new_[49799]_  & \new_[49792]_ ;
  assign \new_[49803]_  = ~A200 & A199;
  assign \new_[49806]_  = A202 & A201;
  assign \new_[49807]_  = \new_[49806]_  & \new_[49803]_ ;
  assign \new_[49810]_  = A233 & ~A232;
  assign \new_[49813]_  = ~A235 & ~A234;
  assign \new_[49814]_  = \new_[49813]_  & \new_[49810]_ ;
  assign \new_[49815]_  = \new_[49814]_  & \new_[49807]_ ;
  assign \new_[49818]_  = A267 & A236;
  assign \new_[49821]_  = A269 & ~A268;
  assign \new_[49822]_  = \new_[49821]_  & \new_[49818]_ ;
  assign \new_[49825]_  = A299 & ~A298;
  assign \new_[49828]_  = A301 & A300;
  assign \new_[49829]_  = \new_[49828]_  & \new_[49825]_ ;
  assign \new_[49830]_  = \new_[49829]_  & \new_[49822]_ ;
  assign \new_[49833]_  = ~A200 & A199;
  assign \new_[49836]_  = A202 & A201;
  assign \new_[49837]_  = \new_[49836]_  & \new_[49833]_ ;
  assign \new_[49840]_  = A233 & ~A232;
  assign \new_[49843]_  = ~A235 & ~A234;
  assign \new_[49844]_  = \new_[49843]_  & \new_[49840]_ ;
  assign \new_[49845]_  = \new_[49844]_  & \new_[49837]_ ;
  assign \new_[49848]_  = A267 & A236;
  assign \new_[49851]_  = A269 & ~A268;
  assign \new_[49852]_  = \new_[49851]_  & \new_[49848]_ ;
  assign \new_[49855]_  = A299 & ~A298;
  assign \new_[49858]_  = ~A302 & A300;
  assign \new_[49859]_  = \new_[49858]_  & \new_[49855]_ ;
  assign \new_[49860]_  = \new_[49859]_  & \new_[49852]_ ;
  assign \new_[49863]_  = ~A200 & A199;
  assign \new_[49866]_  = A202 & A201;
  assign \new_[49867]_  = \new_[49866]_  & \new_[49863]_ ;
  assign \new_[49870]_  = A233 & ~A232;
  assign \new_[49873]_  = ~A235 & ~A234;
  assign \new_[49874]_  = \new_[49873]_  & \new_[49870]_ ;
  assign \new_[49875]_  = \new_[49874]_  & \new_[49867]_ ;
  assign \new_[49878]_  = ~A267 & A236;
  assign \new_[49881]_  = A298 & A268;
  assign \new_[49882]_  = \new_[49881]_  & \new_[49878]_ ;
  assign \new_[49885]_  = ~A300 & ~A299;
  assign \new_[49888]_  = A302 & ~A301;
  assign \new_[49889]_  = \new_[49888]_  & \new_[49885]_ ;
  assign \new_[49890]_  = \new_[49889]_  & \new_[49882]_ ;
  assign \new_[49893]_  = ~A200 & A199;
  assign \new_[49896]_  = A202 & A201;
  assign \new_[49897]_  = \new_[49896]_  & \new_[49893]_ ;
  assign \new_[49900]_  = A233 & ~A232;
  assign \new_[49903]_  = ~A235 & ~A234;
  assign \new_[49904]_  = \new_[49903]_  & \new_[49900]_ ;
  assign \new_[49905]_  = \new_[49904]_  & \new_[49897]_ ;
  assign \new_[49908]_  = ~A267 & A236;
  assign \new_[49911]_  = ~A298 & A268;
  assign \new_[49912]_  = \new_[49911]_  & \new_[49908]_ ;
  assign \new_[49915]_  = ~A300 & A299;
  assign \new_[49918]_  = A302 & ~A301;
  assign \new_[49919]_  = \new_[49918]_  & \new_[49915]_ ;
  assign \new_[49920]_  = \new_[49919]_  & \new_[49912]_ ;
  assign \new_[49923]_  = ~A200 & A199;
  assign \new_[49926]_  = A202 & A201;
  assign \new_[49927]_  = \new_[49926]_  & \new_[49923]_ ;
  assign \new_[49930]_  = A233 & ~A232;
  assign \new_[49933]_  = ~A235 & ~A234;
  assign \new_[49934]_  = \new_[49933]_  & \new_[49930]_ ;
  assign \new_[49935]_  = \new_[49934]_  & \new_[49927]_ ;
  assign \new_[49938]_  = ~A267 & A236;
  assign \new_[49941]_  = A298 & ~A269;
  assign \new_[49942]_  = \new_[49941]_  & \new_[49938]_ ;
  assign \new_[49945]_  = ~A300 & ~A299;
  assign \new_[49948]_  = A302 & ~A301;
  assign \new_[49949]_  = \new_[49948]_  & \new_[49945]_ ;
  assign \new_[49950]_  = \new_[49949]_  & \new_[49942]_ ;
  assign \new_[49953]_  = ~A200 & A199;
  assign \new_[49956]_  = A202 & A201;
  assign \new_[49957]_  = \new_[49956]_  & \new_[49953]_ ;
  assign \new_[49960]_  = A233 & ~A232;
  assign \new_[49963]_  = ~A235 & ~A234;
  assign \new_[49964]_  = \new_[49963]_  & \new_[49960]_ ;
  assign \new_[49965]_  = \new_[49964]_  & \new_[49957]_ ;
  assign \new_[49968]_  = ~A267 & A236;
  assign \new_[49971]_  = ~A298 & ~A269;
  assign \new_[49972]_  = \new_[49971]_  & \new_[49968]_ ;
  assign \new_[49975]_  = ~A300 & A299;
  assign \new_[49978]_  = A302 & ~A301;
  assign \new_[49979]_  = \new_[49978]_  & \new_[49975]_ ;
  assign \new_[49980]_  = \new_[49979]_  & \new_[49972]_ ;
  assign \new_[49983]_  = ~A200 & A199;
  assign \new_[49986]_  = A202 & A201;
  assign \new_[49987]_  = \new_[49986]_  & \new_[49983]_ ;
  assign \new_[49990]_  = A233 & ~A232;
  assign \new_[49993]_  = ~A235 & ~A234;
  assign \new_[49994]_  = \new_[49993]_  & \new_[49990]_ ;
  assign \new_[49995]_  = \new_[49994]_  & \new_[49987]_ ;
  assign \new_[49998]_  = A265 & A236;
  assign \new_[50001]_  = A298 & A266;
  assign \new_[50002]_  = \new_[50001]_  & \new_[49998]_ ;
  assign \new_[50005]_  = ~A300 & ~A299;
  assign \new_[50008]_  = A302 & ~A301;
  assign \new_[50009]_  = \new_[50008]_  & \new_[50005]_ ;
  assign \new_[50010]_  = \new_[50009]_  & \new_[50002]_ ;
  assign \new_[50013]_  = ~A200 & A199;
  assign \new_[50016]_  = A202 & A201;
  assign \new_[50017]_  = \new_[50016]_  & \new_[50013]_ ;
  assign \new_[50020]_  = A233 & ~A232;
  assign \new_[50023]_  = ~A235 & ~A234;
  assign \new_[50024]_  = \new_[50023]_  & \new_[50020]_ ;
  assign \new_[50025]_  = \new_[50024]_  & \new_[50017]_ ;
  assign \new_[50028]_  = A265 & A236;
  assign \new_[50031]_  = ~A298 & A266;
  assign \new_[50032]_  = \new_[50031]_  & \new_[50028]_ ;
  assign \new_[50035]_  = ~A300 & A299;
  assign \new_[50038]_  = A302 & ~A301;
  assign \new_[50039]_  = \new_[50038]_  & \new_[50035]_ ;
  assign \new_[50040]_  = \new_[50039]_  & \new_[50032]_ ;
  assign \new_[50043]_  = ~A200 & A199;
  assign \new_[50046]_  = A202 & A201;
  assign \new_[50047]_  = \new_[50046]_  & \new_[50043]_ ;
  assign \new_[50050]_  = A233 & ~A232;
  assign \new_[50053]_  = ~A235 & ~A234;
  assign \new_[50054]_  = \new_[50053]_  & \new_[50050]_ ;
  assign \new_[50055]_  = \new_[50054]_  & \new_[50047]_ ;
  assign \new_[50058]_  = ~A265 & A236;
  assign \new_[50061]_  = A298 & ~A266;
  assign \new_[50062]_  = \new_[50061]_  & \new_[50058]_ ;
  assign \new_[50065]_  = ~A300 & ~A299;
  assign \new_[50068]_  = A302 & ~A301;
  assign \new_[50069]_  = \new_[50068]_  & \new_[50065]_ ;
  assign \new_[50070]_  = \new_[50069]_  & \new_[50062]_ ;
  assign \new_[50073]_  = ~A200 & A199;
  assign \new_[50076]_  = A202 & A201;
  assign \new_[50077]_  = \new_[50076]_  & \new_[50073]_ ;
  assign \new_[50080]_  = A233 & ~A232;
  assign \new_[50083]_  = ~A235 & ~A234;
  assign \new_[50084]_  = \new_[50083]_  & \new_[50080]_ ;
  assign \new_[50085]_  = \new_[50084]_  & \new_[50077]_ ;
  assign \new_[50088]_  = ~A265 & A236;
  assign \new_[50091]_  = ~A298 & ~A266;
  assign \new_[50092]_  = \new_[50091]_  & \new_[50088]_ ;
  assign \new_[50095]_  = ~A300 & A299;
  assign \new_[50098]_  = A302 & ~A301;
  assign \new_[50099]_  = \new_[50098]_  & \new_[50095]_ ;
  assign \new_[50100]_  = \new_[50099]_  & \new_[50092]_ ;
  assign \new_[50103]_  = ~A200 & A199;
  assign \new_[50106]_  = A202 & A201;
  assign \new_[50107]_  = \new_[50106]_  & \new_[50103]_ ;
  assign \new_[50110]_  = ~A233 & A232;
  assign \new_[50113]_  = A235 & A234;
  assign \new_[50114]_  = \new_[50113]_  & \new_[50110]_ ;
  assign \new_[50115]_  = \new_[50114]_  & \new_[50107]_ ;
  assign \new_[50118]_  = ~A268 & A267;
  assign \new_[50121]_  = A298 & A269;
  assign \new_[50122]_  = \new_[50121]_  & \new_[50118]_ ;
  assign \new_[50125]_  = ~A300 & ~A299;
  assign \new_[50128]_  = A302 & ~A301;
  assign \new_[50129]_  = \new_[50128]_  & \new_[50125]_ ;
  assign \new_[50130]_  = \new_[50129]_  & \new_[50122]_ ;
  assign \new_[50133]_  = ~A200 & A199;
  assign \new_[50136]_  = A202 & A201;
  assign \new_[50137]_  = \new_[50136]_  & \new_[50133]_ ;
  assign \new_[50140]_  = ~A233 & A232;
  assign \new_[50143]_  = A235 & A234;
  assign \new_[50144]_  = \new_[50143]_  & \new_[50140]_ ;
  assign \new_[50145]_  = \new_[50144]_  & \new_[50137]_ ;
  assign \new_[50148]_  = ~A268 & A267;
  assign \new_[50151]_  = ~A298 & A269;
  assign \new_[50152]_  = \new_[50151]_  & \new_[50148]_ ;
  assign \new_[50155]_  = ~A300 & A299;
  assign \new_[50158]_  = A302 & ~A301;
  assign \new_[50159]_  = \new_[50158]_  & \new_[50155]_ ;
  assign \new_[50160]_  = \new_[50159]_  & \new_[50152]_ ;
  assign \new_[50163]_  = ~A200 & A199;
  assign \new_[50166]_  = A202 & A201;
  assign \new_[50167]_  = \new_[50166]_  & \new_[50163]_ ;
  assign \new_[50170]_  = ~A233 & A232;
  assign \new_[50173]_  = ~A236 & A234;
  assign \new_[50174]_  = \new_[50173]_  & \new_[50170]_ ;
  assign \new_[50175]_  = \new_[50174]_  & \new_[50167]_ ;
  assign \new_[50178]_  = ~A268 & A267;
  assign \new_[50181]_  = A298 & A269;
  assign \new_[50182]_  = \new_[50181]_  & \new_[50178]_ ;
  assign \new_[50185]_  = ~A300 & ~A299;
  assign \new_[50188]_  = A302 & ~A301;
  assign \new_[50189]_  = \new_[50188]_  & \new_[50185]_ ;
  assign \new_[50190]_  = \new_[50189]_  & \new_[50182]_ ;
  assign \new_[50193]_  = ~A200 & A199;
  assign \new_[50196]_  = A202 & A201;
  assign \new_[50197]_  = \new_[50196]_  & \new_[50193]_ ;
  assign \new_[50200]_  = ~A233 & A232;
  assign \new_[50203]_  = ~A236 & A234;
  assign \new_[50204]_  = \new_[50203]_  & \new_[50200]_ ;
  assign \new_[50205]_  = \new_[50204]_  & \new_[50197]_ ;
  assign \new_[50208]_  = ~A268 & A267;
  assign \new_[50211]_  = ~A298 & A269;
  assign \new_[50212]_  = \new_[50211]_  & \new_[50208]_ ;
  assign \new_[50215]_  = ~A300 & A299;
  assign \new_[50218]_  = A302 & ~A301;
  assign \new_[50219]_  = \new_[50218]_  & \new_[50215]_ ;
  assign \new_[50220]_  = \new_[50219]_  & \new_[50212]_ ;
  assign \new_[50223]_  = ~A200 & A199;
  assign \new_[50226]_  = A202 & A201;
  assign \new_[50227]_  = \new_[50226]_  & \new_[50223]_ ;
  assign \new_[50230]_  = ~A233 & A232;
  assign \new_[50233]_  = ~A235 & ~A234;
  assign \new_[50234]_  = \new_[50233]_  & \new_[50230]_ ;
  assign \new_[50235]_  = \new_[50234]_  & \new_[50227]_ ;
  assign \new_[50238]_  = A267 & A236;
  assign \new_[50241]_  = A269 & ~A268;
  assign \new_[50242]_  = \new_[50241]_  & \new_[50238]_ ;
  assign \new_[50245]_  = ~A299 & A298;
  assign \new_[50248]_  = A301 & A300;
  assign \new_[50249]_  = \new_[50248]_  & \new_[50245]_ ;
  assign \new_[50250]_  = \new_[50249]_  & \new_[50242]_ ;
  assign \new_[50253]_  = ~A200 & A199;
  assign \new_[50256]_  = A202 & A201;
  assign \new_[50257]_  = \new_[50256]_  & \new_[50253]_ ;
  assign \new_[50260]_  = ~A233 & A232;
  assign \new_[50263]_  = ~A235 & ~A234;
  assign \new_[50264]_  = \new_[50263]_  & \new_[50260]_ ;
  assign \new_[50265]_  = \new_[50264]_  & \new_[50257]_ ;
  assign \new_[50268]_  = A267 & A236;
  assign \new_[50271]_  = A269 & ~A268;
  assign \new_[50272]_  = \new_[50271]_  & \new_[50268]_ ;
  assign \new_[50275]_  = ~A299 & A298;
  assign \new_[50278]_  = ~A302 & A300;
  assign \new_[50279]_  = \new_[50278]_  & \new_[50275]_ ;
  assign \new_[50280]_  = \new_[50279]_  & \new_[50272]_ ;
  assign \new_[50283]_  = ~A200 & A199;
  assign \new_[50286]_  = A202 & A201;
  assign \new_[50287]_  = \new_[50286]_  & \new_[50283]_ ;
  assign \new_[50290]_  = ~A233 & A232;
  assign \new_[50293]_  = ~A235 & ~A234;
  assign \new_[50294]_  = \new_[50293]_  & \new_[50290]_ ;
  assign \new_[50295]_  = \new_[50294]_  & \new_[50287]_ ;
  assign \new_[50298]_  = A267 & A236;
  assign \new_[50301]_  = A269 & ~A268;
  assign \new_[50302]_  = \new_[50301]_  & \new_[50298]_ ;
  assign \new_[50305]_  = A299 & ~A298;
  assign \new_[50308]_  = A301 & A300;
  assign \new_[50309]_  = \new_[50308]_  & \new_[50305]_ ;
  assign \new_[50310]_  = \new_[50309]_  & \new_[50302]_ ;
  assign \new_[50313]_  = ~A200 & A199;
  assign \new_[50316]_  = A202 & A201;
  assign \new_[50317]_  = \new_[50316]_  & \new_[50313]_ ;
  assign \new_[50320]_  = ~A233 & A232;
  assign \new_[50323]_  = ~A235 & ~A234;
  assign \new_[50324]_  = \new_[50323]_  & \new_[50320]_ ;
  assign \new_[50325]_  = \new_[50324]_  & \new_[50317]_ ;
  assign \new_[50328]_  = A267 & A236;
  assign \new_[50331]_  = A269 & ~A268;
  assign \new_[50332]_  = \new_[50331]_  & \new_[50328]_ ;
  assign \new_[50335]_  = A299 & ~A298;
  assign \new_[50338]_  = ~A302 & A300;
  assign \new_[50339]_  = \new_[50338]_  & \new_[50335]_ ;
  assign \new_[50340]_  = \new_[50339]_  & \new_[50332]_ ;
  assign \new_[50343]_  = ~A200 & A199;
  assign \new_[50346]_  = A202 & A201;
  assign \new_[50347]_  = \new_[50346]_  & \new_[50343]_ ;
  assign \new_[50350]_  = ~A233 & A232;
  assign \new_[50353]_  = ~A235 & ~A234;
  assign \new_[50354]_  = \new_[50353]_  & \new_[50350]_ ;
  assign \new_[50355]_  = \new_[50354]_  & \new_[50347]_ ;
  assign \new_[50358]_  = ~A267 & A236;
  assign \new_[50361]_  = A298 & A268;
  assign \new_[50362]_  = \new_[50361]_  & \new_[50358]_ ;
  assign \new_[50365]_  = ~A300 & ~A299;
  assign \new_[50368]_  = A302 & ~A301;
  assign \new_[50369]_  = \new_[50368]_  & \new_[50365]_ ;
  assign \new_[50370]_  = \new_[50369]_  & \new_[50362]_ ;
  assign \new_[50373]_  = ~A200 & A199;
  assign \new_[50376]_  = A202 & A201;
  assign \new_[50377]_  = \new_[50376]_  & \new_[50373]_ ;
  assign \new_[50380]_  = ~A233 & A232;
  assign \new_[50383]_  = ~A235 & ~A234;
  assign \new_[50384]_  = \new_[50383]_  & \new_[50380]_ ;
  assign \new_[50385]_  = \new_[50384]_  & \new_[50377]_ ;
  assign \new_[50388]_  = ~A267 & A236;
  assign \new_[50391]_  = ~A298 & A268;
  assign \new_[50392]_  = \new_[50391]_  & \new_[50388]_ ;
  assign \new_[50395]_  = ~A300 & A299;
  assign \new_[50398]_  = A302 & ~A301;
  assign \new_[50399]_  = \new_[50398]_  & \new_[50395]_ ;
  assign \new_[50400]_  = \new_[50399]_  & \new_[50392]_ ;
  assign \new_[50403]_  = ~A200 & A199;
  assign \new_[50406]_  = A202 & A201;
  assign \new_[50407]_  = \new_[50406]_  & \new_[50403]_ ;
  assign \new_[50410]_  = ~A233 & A232;
  assign \new_[50413]_  = ~A235 & ~A234;
  assign \new_[50414]_  = \new_[50413]_  & \new_[50410]_ ;
  assign \new_[50415]_  = \new_[50414]_  & \new_[50407]_ ;
  assign \new_[50418]_  = ~A267 & A236;
  assign \new_[50421]_  = A298 & ~A269;
  assign \new_[50422]_  = \new_[50421]_  & \new_[50418]_ ;
  assign \new_[50425]_  = ~A300 & ~A299;
  assign \new_[50428]_  = A302 & ~A301;
  assign \new_[50429]_  = \new_[50428]_  & \new_[50425]_ ;
  assign \new_[50430]_  = \new_[50429]_  & \new_[50422]_ ;
  assign \new_[50433]_  = ~A200 & A199;
  assign \new_[50436]_  = A202 & A201;
  assign \new_[50437]_  = \new_[50436]_  & \new_[50433]_ ;
  assign \new_[50440]_  = ~A233 & A232;
  assign \new_[50443]_  = ~A235 & ~A234;
  assign \new_[50444]_  = \new_[50443]_  & \new_[50440]_ ;
  assign \new_[50445]_  = \new_[50444]_  & \new_[50437]_ ;
  assign \new_[50448]_  = ~A267 & A236;
  assign \new_[50451]_  = ~A298 & ~A269;
  assign \new_[50452]_  = \new_[50451]_  & \new_[50448]_ ;
  assign \new_[50455]_  = ~A300 & A299;
  assign \new_[50458]_  = A302 & ~A301;
  assign \new_[50459]_  = \new_[50458]_  & \new_[50455]_ ;
  assign \new_[50460]_  = \new_[50459]_  & \new_[50452]_ ;
  assign \new_[50463]_  = ~A200 & A199;
  assign \new_[50466]_  = A202 & A201;
  assign \new_[50467]_  = \new_[50466]_  & \new_[50463]_ ;
  assign \new_[50470]_  = ~A233 & A232;
  assign \new_[50473]_  = ~A235 & ~A234;
  assign \new_[50474]_  = \new_[50473]_  & \new_[50470]_ ;
  assign \new_[50475]_  = \new_[50474]_  & \new_[50467]_ ;
  assign \new_[50478]_  = A265 & A236;
  assign \new_[50481]_  = A298 & A266;
  assign \new_[50482]_  = \new_[50481]_  & \new_[50478]_ ;
  assign \new_[50485]_  = ~A300 & ~A299;
  assign \new_[50488]_  = A302 & ~A301;
  assign \new_[50489]_  = \new_[50488]_  & \new_[50485]_ ;
  assign \new_[50490]_  = \new_[50489]_  & \new_[50482]_ ;
  assign \new_[50493]_  = ~A200 & A199;
  assign \new_[50496]_  = A202 & A201;
  assign \new_[50497]_  = \new_[50496]_  & \new_[50493]_ ;
  assign \new_[50500]_  = ~A233 & A232;
  assign \new_[50503]_  = ~A235 & ~A234;
  assign \new_[50504]_  = \new_[50503]_  & \new_[50500]_ ;
  assign \new_[50505]_  = \new_[50504]_  & \new_[50497]_ ;
  assign \new_[50508]_  = A265 & A236;
  assign \new_[50511]_  = ~A298 & A266;
  assign \new_[50512]_  = \new_[50511]_  & \new_[50508]_ ;
  assign \new_[50515]_  = ~A300 & A299;
  assign \new_[50518]_  = A302 & ~A301;
  assign \new_[50519]_  = \new_[50518]_  & \new_[50515]_ ;
  assign \new_[50520]_  = \new_[50519]_  & \new_[50512]_ ;
  assign \new_[50523]_  = ~A200 & A199;
  assign \new_[50526]_  = A202 & A201;
  assign \new_[50527]_  = \new_[50526]_  & \new_[50523]_ ;
  assign \new_[50530]_  = ~A233 & A232;
  assign \new_[50533]_  = ~A235 & ~A234;
  assign \new_[50534]_  = \new_[50533]_  & \new_[50530]_ ;
  assign \new_[50535]_  = \new_[50534]_  & \new_[50527]_ ;
  assign \new_[50538]_  = ~A265 & A236;
  assign \new_[50541]_  = A298 & ~A266;
  assign \new_[50542]_  = \new_[50541]_  & \new_[50538]_ ;
  assign \new_[50545]_  = ~A300 & ~A299;
  assign \new_[50548]_  = A302 & ~A301;
  assign \new_[50549]_  = \new_[50548]_  & \new_[50545]_ ;
  assign \new_[50550]_  = \new_[50549]_  & \new_[50542]_ ;
  assign \new_[50553]_  = ~A200 & A199;
  assign \new_[50556]_  = A202 & A201;
  assign \new_[50557]_  = \new_[50556]_  & \new_[50553]_ ;
  assign \new_[50560]_  = ~A233 & A232;
  assign \new_[50563]_  = ~A235 & ~A234;
  assign \new_[50564]_  = \new_[50563]_  & \new_[50560]_ ;
  assign \new_[50565]_  = \new_[50564]_  & \new_[50557]_ ;
  assign \new_[50568]_  = ~A265 & A236;
  assign \new_[50571]_  = ~A298 & ~A266;
  assign \new_[50572]_  = \new_[50571]_  & \new_[50568]_ ;
  assign \new_[50575]_  = ~A300 & A299;
  assign \new_[50578]_  = A302 & ~A301;
  assign \new_[50579]_  = \new_[50578]_  & \new_[50575]_ ;
  assign \new_[50580]_  = \new_[50579]_  & \new_[50572]_ ;
  assign \new_[50583]_  = ~A200 & A199;
  assign \new_[50586]_  = ~A203 & A201;
  assign \new_[50587]_  = \new_[50586]_  & \new_[50583]_ ;
  assign \new_[50590]_  = A233 & ~A232;
  assign \new_[50593]_  = A235 & A234;
  assign \new_[50594]_  = \new_[50593]_  & \new_[50590]_ ;
  assign \new_[50595]_  = \new_[50594]_  & \new_[50587]_ ;
  assign \new_[50598]_  = ~A268 & A267;
  assign \new_[50601]_  = A298 & A269;
  assign \new_[50602]_  = \new_[50601]_  & \new_[50598]_ ;
  assign \new_[50605]_  = ~A300 & ~A299;
  assign \new_[50608]_  = A302 & ~A301;
  assign \new_[50609]_  = \new_[50608]_  & \new_[50605]_ ;
  assign \new_[50610]_  = \new_[50609]_  & \new_[50602]_ ;
  assign \new_[50613]_  = ~A200 & A199;
  assign \new_[50616]_  = ~A203 & A201;
  assign \new_[50617]_  = \new_[50616]_  & \new_[50613]_ ;
  assign \new_[50620]_  = A233 & ~A232;
  assign \new_[50623]_  = A235 & A234;
  assign \new_[50624]_  = \new_[50623]_  & \new_[50620]_ ;
  assign \new_[50625]_  = \new_[50624]_  & \new_[50617]_ ;
  assign \new_[50628]_  = ~A268 & A267;
  assign \new_[50631]_  = ~A298 & A269;
  assign \new_[50632]_  = \new_[50631]_  & \new_[50628]_ ;
  assign \new_[50635]_  = ~A300 & A299;
  assign \new_[50638]_  = A302 & ~A301;
  assign \new_[50639]_  = \new_[50638]_  & \new_[50635]_ ;
  assign \new_[50640]_  = \new_[50639]_  & \new_[50632]_ ;
  assign \new_[50643]_  = ~A200 & A199;
  assign \new_[50646]_  = ~A203 & A201;
  assign \new_[50647]_  = \new_[50646]_  & \new_[50643]_ ;
  assign \new_[50650]_  = A233 & ~A232;
  assign \new_[50653]_  = ~A236 & A234;
  assign \new_[50654]_  = \new_[50653]_  & \new_[50650]_ ;
  assign \new_[50655]_  = \new_[50654]_  & \new_[50647]_ ;
  assign \new_[50658]_  = ~A268 & A267;
  assign \new_[50661]_  = A298 & A269;
  assign \new_[50662]_  = \new_[50661]_  & \new_[50658]_ ;
  assign \new_[50665]_  = ~A300 & ~A299;
  assign \new_[50668]_  = A302 & ~A301;
  assign \new_[50669]_  = \new_[50668]_  & \new_[50665]_ ;
  assign \new_[50670]_  = \new_[50669]_  & \new_[50662]_ ;
  assign \new_[50673]_  = ~A200 & A199;
  assign \new_[50676]_  = ~A203 & A201;
  assign \new_[50677]_  = \new_[50676]_  & \new_[50673]_ ;
  assign \new_[50680]_  = A233 & ~A232;
  assign \new_[50683]_  = ~A236 & A234;
  assign \new_[50684]_  = \new_[50683]_  & \new_[50680]_ ;
  assign \new_[50685]_  = \new_[50684]_  & \new_[50677]_ ;
  assign \new_[50688]_  = ~A268 & A267;
  assign \new_[50691]_  = ~A298 & A269;
  assign \new_[50692]_  = \new_[50691]_  & \new_[50688]_ ;
  assign \new_[50695]_  = ~A300 & A299;
  assign \new_[50698]_  = A302 & ~A301;
  assign \new_[50699]_  = \new_[50698]_  & \new_[50695]_ ;
  assign \new_[50700]_  = \new_[50699]_  & \new_[50692]_ ;
  assign \new_[50703]_  = ~A200 & A199;
  assign \new_[50706]_  = ~A203 & A201;
  assign \new_[50707]_  = \new_[50706]_  & \new_[50703]_ ;
  assign \new_[50710]_  = A233 & ~A232;
  assign \new_[50713]_  = ~A235 & ~A234;
  assign \new_[50714]_  = \new_[50713]_  & \new_[50710]_ ;
  assign \new_[50715]_  = \new_[50714]_  & \new_[50707]_ ;
  assign \new_[50718]_  = A267 & A236;
  assign \new_[50721]_  = A269 & ~A268;
  assign \new_[50722]_  = \new_[50721]_  & \new_[50718]_ ;
  assign \new_[50725]_  = ~A299 & A298;
  assign \new_[50728]_  = A301 & A300;
  assign \new_[50729]_  = \new_[50728]_  & \new_[50725]_ ;
  assign \new_[50730]_  = \new_[50729]_  & \new_[50722]_ ;
  assign \new_[50733]_  = ~A200 & A199;
  assign \new_[50736]_  = ~A203 & A201;
  assign \new_[50737]_  = \new_[50736]_  & \new_[50733]_ ;
  assign \new_[50740]_  = A233 & ~A232;
  assign \new_[50743]_  = ~A235 & ~A234;
  assign \new_[50744]_  = \new_[50743]_  & \new_[50740]_ ;
  assign \new_[50745]_  = \new_[50744]_  & \new_[50737]_ ;
  assign \new_[50748]_  = A267 & A236;
  assign \new_[50751]_  = A269 & ~A268;
  assign \new_[50752]_  = \new_[50751]_  & \new_[50748]_ ;
  assign \new_[50755]_  = ~A299 & A298;
  assign \new_[50758]_  = ~A302 & A300;
  assign \new_[50759]_  = \new_[50758]_  & \new_[50755]_ ;
  assign \new_[50760]_  = \new_[50759]_  & \new_[50752]_ ;
  assign \new_[50763]_  = ~A200 & A199;
  assign \new_[50766]_  = ~A203 & A201;
  assign \new_[50767]_  = \new_[50766]_  & \new_[50763]_ ;
  assign \new_[50770]_  = A233 & ~A232;
  assign \new_[50773]_  = ~A235 & ~A234;
  assign \new_[50774]_  = \new_[50773]_  & \new_[50770]_ ;
  assign \new_[50775]_  = \new_[50774]_  & \new_[50767]_ ;
  assign \new_[50778]_  = A267 & A236;
  assign \new_[50781]_  = A269 & ~A268;
  assign \new_[50782]_  = \new_[50781]_  & \new_[50778]_ ;
  assign \new_[50785]_  = A299 & ~A298;
  assign \new_[50788]_  = A301 & A300;
  assign \new_[50789]_  = \new_[50788]_  & \new_[50785]_ ;
  assign \new_[50790]_  = \new_[50789]_  & \new_[50782]_ ;
  assign \new_[50793]_  = ~A200 & A199;
  assign \new_[50796]_  = ~A203 & A201;
  assign \new_[50797]_  = \new_[50796]_  & \new_[50793]_ ;
  assign \new_[50800]_  = A233 & ~A232;
  assign \new_[50803]_  = ~A235 & ~A234;
  assign \new_[50804]_  = \new_[50803]_  & \new_[50800]_ ;
  assign \new_[50805]_  = \new_[50804]_  & \new_[50797]_ ;
  assign \new_[50808]_  = A267 & A236;
  assign \new_[50811]_  = A269 & ~A268;
  assign \new_[50812]_  = \new_[50811]_  & \new_[50808]_ ;
  assign \new_[50815]_  = A299 & ~A298;
  assign \new_[50818]_  = ~A302 & A300;
  assign \new_[50819]_  = \new_[50818]_  & \new_[50815]_ ;
  assign \new_[50820]_  = \new_[50819]_  & \new_[50812]_ ;
  assign \new_[50823]_  = ~A200 & A199;
  assign \new_[50826]_  = ~A203 & A201;
  assign \new_[50827]_  = \new_[50826]_  & \new_[50823]_ ;
  assign \new_[50830]_  = A233 & ~A232;
  assign \new_[50833]_  = ~A235 & ~A234;
  assign \new_[50834]_  = \new_[50833]_  & \new_[50830]_ ;
  assign \new_[50835]_  = \new_[50834]_  & \new_[50827]_ ;
  assign \new_[50838]_  = ~A267 & A236;
  assign \new_[50841]_  = A298 & A268;
  assign \new_[50842]_  = \new_[50841]_  & \new_[50838]_ ;
  assign \new_[50845]_  = ~A300 & ~A299;
  assign \new_[50848]_  = A302 & ~A301;
  assign \new_[50849]_  = \new_[50848]_  & \new_[50845]_ ;
  assign \new_[50850]_  = \new_[50849]_  & \new_[50842]_ ;
  assign \new_[50853]_  = ~A200 & A199;
  assign \new_[50856]_  = ~A203 & A201;
  assign \new_[50857]_  = \new_[50856]_  & \new_[50853]_ ;
  assign \new_[50860]_  = A233 & ~A232;
  assign \new_[50863]_  = ~A235 & ~A234;
  assign \new_[50864]_  = \new_[50863]_  & \new_[50860]_ ;
  assign \new_[50865]_  = \new_[50864]_  & \new_[50857]_ ;
  assign \new_[50868]_  = ~A267 & A236;
  assign \new_[50871]_  = ~A298 & A268;
  assign \new_[50872]_  = \new_[50871]_  & \new_[50868]_ ;
  assign \new_[50875]_  = ~A300 & A299;
  assign \new_[50878]_  = A302 & ~A301;
  assign \new_[50879]_  = \new_[50878]_  & \new_[50875]_ ;
  assign \new_[50880]_  = \new_[50879]_  & \new_[50872]_ ;
  assign \new_[50883]_  = ~A200 & A199;
  assign \new_[50886]_  = ~A203 & A201;
  assign \new_[50887]_  = \new_[50886]_  & \new_[50883]_ ;
  assign \new_[50890]_  = A233 & ~A232;
  assign \new_[50893]_  = ~A235 & ~A234;
  assign \new_[50894]_  = \new_[50893]_  & \new_[50890]_ ;
  assign \new_[50895]_  = \new_[50894]_  & \new_[50887]_ ;
  assign \new_[50898]_  = ~A267 & A236;
  assign \new_[50901]_  = A298 & ~A269;
  assign \new_[50902]_  = \new_[50901]_  & \new_[50898]_ ;
  assign \new_[50905]_  = ~A300 & ~A299;
  assign \new_[50908]_  = A302 & ~A301;
  assign \new_[50909]_  = \new_[50908]_  & \new_[50905]_ ;
  assign \new_[50910]_  = \new_[50909]_  & \new_[50902]_ ;
  assign \new_[50913]_  = ~A200 & A199;
  assign \new_[50916]_  = ~A203 & A201;
  assign \new_[50917]_  = \new_[50916]_  & \new_[50913]_ ;
  assign \new_[50920]_  = A233 & ~A232;
  assign \new_[50923]_  = ~A235 & ~A234;
  assign \new_[50924]_  = \new_[50923]_  & \new_[50920]_ ;
  assign \new_[50925]_  = \new_[50924]_  & \new_[50917]_ ;
  assign \new_[50928]_  = ~A267 & A236;
  assign \new_[50931]_  = ~A298 & ~A269;
  assign \new_[50932]_  = \new_[50931]_  & \new_[50928]_ ;
  assign \new_[50935]_  = ~A300 & A299;
  assign \new_[50938]_  = A302 & ~A301;
  assign \new_[50939]_  = \new_[50938]_  & \new_[50935]_ ;
  assign \new_[50940]_  = \new_[50939]_  & \new_[50932]_ ;
  assign \new_[50943]_  = ~A200 & A199;
  assign \new_[50946]_  = ~A203 & A201;
  assign \new_[50947]_  = \new_[50946]_  & \new_[50943]_ ;
  assign \new_[50950]_  = A233 & ~A232;
  assign \new_[50953]_  = ~A235 & ~A234;
  assign \new_[50954]_  = \new_[50953]_  & \new_[50950]_ ;
  assign \new_[50955]_  = \new_[50954]_  & \new_[50947]_ ;
  assign \new_[50958]_  = A265 & A236;
  assign \new_[50961]_  = A298 & A266;
  assign \new_[50962]_  = \new_[50961]_  & \new_[50958]_ ;
  assign \new_[50965]_  = ~A300 & ~A299;
  assign \new_[50968]_  = A302 & ~A301;
  assign \new_[50969]_  = \new_[50968]_  & \new_[50965]_ ;
  assign \new_[50970]_  = \new_[50969]_  & \new_[50962]_ ;
  assign \new_[50973]_  = ~A200 & A199;
  assign \new_[50976]_  = ~A203 & A201;
  assign \new_[50977]_  = \new_[50976]_  & \new_[50973]_ ;
  assign \new_[50980]_  = A233 & ~A232;
  assign \new_[50983]_  = ~A235 & ~A234;
  assign \new_[50984]_  = \new_[50983]_  & \new_[50980]_ ;
  assign \new_[50985]_  = \new_[50984]_  & \new_[50977]_ ;
  assign \new_[50988]_  = A265 & A236;
  assign \new_[50991]_  = ~A298 & A266;
  assign \new_[50992]_  = \new_[50991]_  & \new_[50988]_ ;
  assign \new_[50995]_  = ~A300 & A299;
  assign \new_[50998]_  = A302 & ~A301;
  assign \new_[50999]_  = \new_[50998]_  & \new_[50995]_ ;
  assign \new_[51000]_  = \new_[50999]_  & \new_[50992]_ ;
  assign \new_[51003]_  = ~A200 & A199;
  assign \new_[51006]_  = ~A203 & A201;
  assign \new_[51007]_  = \new_[51006]_  & \new_[51003]_ ;
  assign \new_[51010]_  = A233 & ~A232;
  assign \new_[51013]_  = ~A235 & ~A234;
  assign \new_[51014]_  = \new_[51013]_  & \new_[51010]_ ;
  assign \new_[51015]_  = \new_[51014]_  & \new_[51007]_ ;
  assign \new_[51018]_  = ~A265 & A236;
  assign \new_[51021]_  = A298 & ~A266;
  assign \new_[51022]_  = \new_[51021]_  & \new_[51018]_ ;
  assign \new_[51025]_  = ~A300 & ~A299;
  assign \new_[51028]_  = A302 & ~A301;
  assign \new_[51029]_  = \new_[51028]_  & \new_[51025]_ ;
  assign \new_[51030]_  = \new_[51029]_  & \new_[51022]_ ;
  assign \new_[51033]_  = ~A200 & A199;
  assign \new_[51036]_  = ~A203 & A201;
  assign \new_[51037]_  = \new_[51036]_  & \new_[51033]_ ;
  assign \new_[51040]_  = A233 & ~A232;
  assign \new_[51043]_  = ~A235 & ~A234;
  assign \new_[51044]_  = \new_[51043]_  & \new_[51040]_ ;
  assign \new_[51045]_  = \new_[51044]_  & \new_[51037]_ ;
  assign \new_[51048]_  = ~A265 & A236;
  assign \new_[51051]_  = ~A298 & ~A266;
  assign \new_[51052]_  = \new_[51051]_  & \new_[51048]_ ;
  assign \new_[51055]_  = ~A300 & A299;
  assign \new_[51058]_  = A302 & ~A301;
  assign \new_[51059]_  = \new_[51058]_  & \new_[51055]_ ;
  assign \new_[51060]_  = \new_[51059]_  & \new_[51052]_ ;
  assign \new_[51063]_  = ~A200 & A199;
  assign \new_[51066]_  = ~A203 & A201;
  assign \new_[51067]_  = \new_[51066]_  & \new_[51063]_ ;
  assign \new_[51070]_  = ~A233 & A232;
  assign \new_[51073]_  = A235 & A234;
  assign \new_[51074]_  = \new_[51073]_  & \new_[51070]_ ;
  assign \new_[51075]_  = \new_[51074]_  & \new_[51067]_ ;
  assign \new_[51078]_  = ~A268 & A267;
  assign \new_[51081]_  = A298 & A269;
  assign \new_[51082]_  = \new_[51081]_  & \new_[51078]_ ;
  assign \new_[51085]_  = ~A300 & ~A299;
  assign \new_[51088]_  = A302 & ~A301;
  assign \new_[51089]_  = \new_[51088]_  & \new_[51085]_ ;
  assign \new_[51090]_  = \new_[51089]_  & \new_[51082]_ ;
  assign \new_[51093]_  = ~A200 & A199;
  assign \new_[51096]_  = ~A203 & A201;
  assign \new_[51097]_  = \new_[51096]_  & \new_[51093]_ ;
  assign \new_[51100]_  = ~A233 & A232;
  assign \new_[51103]_  = A235 & A234;
  assign \new_[51104]_  = \new_[51103]_  & \new_[51100]_ ;
  assign \new_[51105]_  = \new_[51104]_  & \new_[51097]_ ;
  assign \new_[51108]_  = ~A268 & A267;
  assign \new_[51111]_  = ~A298 & A269;
  assign \new_[51112]_  = \new_[51111]_  & \new_[51108]_ ;
  assign \new_[51115]_  = ~A300 & A299;
  assign \new_[51118]_  = A302 & ~A301;
  assign \new_[51119]_  = \new_[51118]_  & \new_[51115]_ ;
  assign \new_[51120]_  = \new_[51119]_  & \new_[51112]_ ;
  assign \new_[51123]_  = ~A200 & A199;
  assign \new_[51126]_  = ~A203 & A201;
  assign \new_[51127]_  = \new_[51126]_  & \new_[51123]_ ;
  assign \new_[51130]_  = ~A233 & A232;
  assign \new_[51133]_  = ~A236 & A234;
  assign \new_[51134]_  = \new_[51133]_  & \new_[51130]_ ;
  assign \new_[51135]_  = \new_[51134]_  & \new_[51127]_ ;
  assign \new_[51138]_  = ~A268 & A267;
  assign \new_[51141]_  = A298 & A269;
  assign \new_[51142]_  = \new_[51141]_  & \new_[51138]_ ;
  assign \new_[51145]_  = ~A300 & ~A299;
  assign \new_[51148]_  = A302 & ~A301;
  assign \new_[51149]_  = \new_[51148]_  & \new_[51145]_ ;
  assign \new_[51150]_  = \new_[51149]_  & \new_[51142]_ ;
  assign \new_[51153]_  = ~A200 & A199;
  assign \new_[51156]_  = ~A203 & A201;
  assign \new_[51157]_  = \new_[51156]_  & \new_[51153]_ ;
  assign \new_[51160]_  = ~A233 & A232;
  assign \new_[51163]_  = ~A236 & A234;
  assign \new_[51164]_  = \new_[51163]_  & \new_[51160]_ ;
  assign \new_[51165]_  = \new_[51164]_  & \new_[51157]_ ;
  assign \new_[51168]_  = ~A268 & A267;
  assign \new_[51171]_  = ~A298 & A269;
  assign \new_[51172]_  = \new_[51171]_  & \new_[51168]_ ;
  assign \new_[51175]_  = ~A300 & A299;
  assign \new_[51178]_  = A302 & ~A301;
  assign \new_[51179]_  = \new_[51178]_  & \new_[51175]_ ;
  assign \new_[51180]_  = \new_[51179]_  & \new_[51172]_ ;
  assign \new_[51183]_  = ~A200 & A199;
  assign \new_[51186]_  = ~A203 & A201;
  assign \new_[51187]_  = \new_[51186]_  & \new_[51183]_ ;
  assign \new_[51190]_  = ~A233 & A232;
  assign \new_[51193]_  = ~A235 & ~A234;
  assign \new_[51194]_  = \new_[51193]_  & \new_[51190]_ ;
  assign \new_[51195]_  = \new_[51194]_  & \new_[51187]_ ;
  assign \new_[51198]_  = A267 & A236;
  assign \new_[51201]_  = A269 & ~A268;
  assign \new_[51202]_  = \new_[51201]_  & \new_[51198]_ ;
  assign \new_[51205]_  = ~A299 & A298;
  assign \new_[51208]_  = A301 & A300;
  assign \new_[51209]_  = \new_[51208]_  & \new_[51205]_ ;
  assign \new_[51210]_  = \new_[51209]_  & \new_[51202]_ ;
  assign \new_[51213]_  = ~A200 & A199;
  assign \new_[51216]_  = ~A203 & A201;
  assign \new_[51217]_  = \new_[51216]_  & \new_[51213]_ ;
  assign \new_[51220]_  = ~A233 & A232;
  assign \new_[51223]_  = ~A235 & ~A234;
  assign \new_[51224]_  = \new_[51223]_  & \new_[51220]_ ;
  assign \new_[51225]_  = \new_[51224]_  & \new_[51217]_ ;
  assign \new_[51228]_  = A267 & A236;
  assign \new_[51231]_  = A269 & ~A268;
  assign \new_[51232]_  = \new_[51231]_  & \new_[51228]_ ;
  assign \new_[51235]_  = ~A299 & A298;
  assign \new_[51238]_  = ~A302 & A300;
  assign \new_[51239]_  = \new_[51238]_  & \new_[51235]_ ;
  assign \new_[51240]_  = \new_[51239]_  & \new_[51232]_ ;
  assign \new_[51243]_  = ~A200 & A199;
  assign \new_[51246]_  = ~A203 & A201;
  assign \new_[51247]_  = \new_[51246]_  & \new_[51243]_ ;
  assign \new_[51250]_  = ~A233 & A232;
  assign \new_[51253]_  = ~A235 & ~A234;
  assign \new_[51254]_  = \new_[51253]_  & \new_[51250]_ ;
  assign \new_[51255]_  = \new_[51254]_  & \new_[51247]_ ;
  assign \new_[51258]_  = A267 & A236;
  assign \new_[51261]_  = A269 & ~A268;
  assign \new_[51262]_  = \new_[51261]_  & \new_[51258]_ ;
  assign \new_[51265]_  = A299 & ~A298;
  assign \new_[51268]_  = A301 & A300;
  assign \new_[51269]_  = \new_[51268]_  & \new_[51265]_ ;
  assign \new_[51270]_  = \new_[51269]_  & \new_[51262]_ ;
  assign \new_[51273]_  = ~A200 & A199;
  assign \new_[51276]_  = ~A203 & A201;
  assign \new_[51277]_  = \new_[51276]_  & \new_[51273]_ ;
  assign \new_[51280]_  = ~A233 & A232;
  assign \new_[51283]_  = ~A235 & ~A234;
  assign \new_[51284]_  = \new_[51283]_  & \new_[51280]_ ;
  assign \new_[51285]_  = \new_[51284]_  & \new_[51277]_ ;
  assign \new_[51288]_  = A267 & A236;
  assign \new_[51291]_  = A269 & ~A268;
  assign \new_[51292]_  = \new_[51291]_  & \new_[51288]_ ;
  assign \new_[51295]_  = A299 & ~A298;
  assign \new_[51298]_  = ~A302 & A300;
  assign \new_[51299]_  = \new_[51298]_  & \new_[51295]_ ;
  assign \new_[51300]_  = \new_[51299]_  & \new_[51292]_ ;
  assign \new_[51303]_  = ~A200 & A199;
  assign \new_[51306]_  = ~A203 & A201;
  assign \new_[51307]_  = \new_[51306]_  & \new_[51303]_ ;
  assign \new_[51310]_  = ~A233 & A232;
  assign \new_[51313]_  = ~A235 & ~A234;
  assign \new_[51314]_  = \new_[51313]_  & \new_[51310]_ ;
  assign \new_[51315]_  = \new_[51314]_  & \new_[51307]_ ;
  assign \new_[51318]_  = ~A267 & A236;
  assign \new_[51321]_  = A298 & A268;
  assign \new_[51322]_  = \new_[51321]_  & \new_[51318]_ ;
  assign \new_[51325]_  = ~A300 & ~A299;
  assign \new_[51328]_  = A302 & ~A301;
  assign \new_[51329]_  = \new_[51328]_  & \new_[51325]_ ;
  assign \new_[51330]_  = \new_[51329]_  & \new_[51322]_ ;
  assign \new_[51333]_  = ~A200 & A199;
  assign \new_[51336]_  = ~A203 & A201;
  assign \new_[51337]_  = \new_[51336]_  & \new_[51333]_ ;
  assign \new_[51340]_  = ~A233 & A232;
  assign \new_[51343]_  = ~A235 & ~A234;
  assign \new_[51344]_  = \new_[51343]_  & \new_[51340]_ ;
  assign \new_[51345]_  = \new_[51344]_  & \new_[51337]_ ;
  assign \new_[51348]_  = ~A267 & A236;
  assign \new_[51351]_  = ~A298 & A268;
  assign \new_[51352]_  = \new_[51351]_  & \new_[51348]_ ;
  assign \new_[51355]_  = ~A300 & A299;
  assign \new_[51358]_  = A302 & ~A301;
  assign \new_[51359]_  = \new_[51358]_  & \new_[51355]_ ;
  assign \new_[51360]_  = \new_[51359]_  & \new_[51352]_ ;
  assign \new_[51363]_  = ~A200 & A199;
  assign \new_[51366]_  = ~A203 & A201;
  assign \new_[51367]_  = \new_[51366]_  & \new_[51363]_ ;
  assign \new_[51370]_  = ~A233 & A232;
  assign \new_[51373]_  = ~A235 & ~A234;
  assign \new_[51374]_  = \new_[51373]_  & \new_[51370]_ ;
  assign \new_[51375]_  = \new_[51374]_  & \new_[51367]_ ;
  assign \new_[51378]_  = ~A267 & A236;
  assign \new_[51381]_  = A298 & ~A269;
  assign \new_[51382]_  = \new_[51381]_  & \new_[51378]_ ;
  assign \new_[51385]_  = ~A300 & ~A299;
  assign \new_[51388]_  = A302 & ~A301;
  assign \new_[51389]_  = \new_[51388]_  & \new_[51385]_ ;
  assign \new_[51390]_  = \new_[51389]_  & \new_[51382]_ ;
  assign \new_[51393]_  = ~A200 & A199;
  assign \new_[51396]_  = ~A203 & A201;
  assign \new_[51397]_  = \new_[51396]_  & \new_[51393]_ ;
  assign \new_[51400]_  = ~A233 & A232;
  assign \new_[51403]_  = ~A235 & ~A234;
  assign \new_[51404]_  = \new_[51403]_  & \new_[51400]_ ;
  assign \new_[51405]_  = \new_[51404]_  & \new_[51397]_ ;
  assign \new_[51408]_  = ~A267 & A236;
  assign \new_[51411]_  = ~A298 & ~A269;
  assign \new_[51412]_  = \new_[51411]_  & \new_[51408]_ ;
  assign \new_[51415]_  = ~A300 & A299;
  assign \new_[51418]_  = A302 & ~A301;
  assign \new_[51419]_  = \new_[51418]_  & \new_[51415]_ ;
  assign \new_[51420]_  = \new_[51419]_  & \new_[51412]_ ;
  assign \new_[51423]_  = ~A200 & A199;
  assign \new_[51426]_  = ~A203 & A201;
  assign \new_[51427]_  = \new_[51426]_  & \new_[51423]_ ;
  assign \new_[51430]_  = ~A233 & A232;
  assign \new_[51433]_  = ~A235 & ~A234;
  assign \new_[51434]_  = \new_[51433]_  & \new_[51430]_ ;
  assign \new_[51435]_  = \new_[51434]_  & \new_[51427]_ ;
  assign \new_[51438]_  = A265 & A236;
  assign \new_[51441]_  = A298 & A266;
  assign \new_[51442]_  = \new_[51441]_  & \new_[51438]_ ;
  assign \new_[51445]_  = ~A300 & ~A299;
  assign \new_[51448]_  = A302 & ~A301;
  assign \new_[51449]_  = \new_[51448]_  & \new_[51445]_ ;
  assign \new_[51450]_  = \new_[51449]_  & \new_[51442]_ ;
  assign \new_[51453]_  = ~A200 & A199;
  assign \new_[51456]_  = ~A203 & A201;
  assign \new_[51457]_  = \new_[51456]_  & \new_[51453]_ ;
  assign \new_[51460]_  = ~A233 & A232;
  assign \new_[51463]_  = ~A235 & ~A234;
  assign \new_[51464]_  = \new_[51463]_  & \new_[51460]_ ;
  assign \new_[51465]_  = \new_[51464]_  & \new_[51457]_ ;
  assign \new_[51468]_  = A265 & A236;
  assign \new_[51471]_  = ~A298 & A266;
  assign \new_[51472]_  = \new_[51471]_  & \new_[51468]_ ;
  assign \new_[51475]_  = ~A300 & A299;
  assign \new_[51478]_  = A302 & ~A301;
  assign \new_[51479]_  = \new_[51478]_  & \new_[51475]_ ;
  assign \new_[51480]_  = \new_[51479]_  & \new_[51472]_ ;
  assign \new_[51483]_  = ~A200 & A199;
  assign \new_[51486]_  = ~A203 & A201;
  assign \new_[51487]_  = \new_[51486]_  & \new_[51483]_ ;
  assign \new_[51490]_  = ~A233 & A232;
  assign \new_[51493]_  = ~A235 & ~A234;
  assign \new_[51494]_  = \new_[51493]_  & \new_[51490]_ ;
  assign \new_[51495]_  = \new_[51494]_  & \new_[51487]_ ;
  assign \new_[51498]_  = ~A265 & A236;
  assign \new_[51501]_  = A298 & ~A266;
  assign \new_[51502]_  = \new_[51501]_  & \new_[51498]_ ;
  assign \new_[51505]_  = ~A300 & ~A299;
  assign \new_[51508]_  = A302 & ~A301;
  assign \new_[51509]_  = \new_[51508]_  & \new_[51505]_ ;
  assign \new_[51510]_  = \new_[51509]_  & \new_[51502]_ ;
  assign \new_[51513]_  = ~A200 & A199;
  assign \new_[51516]_  = ~A203 & A201;
  assign \new_[51517]_  = \new_[51516]_  & \new_[51513]_ ;
  assign \new_[51520]_  = ~A233 & A232;
  assign \new_[51523]_  = ~A235 & ~A234;
  assign \new_[51524]_  = \new_[51523]_  & \new_[51520]_ ;
  assign \new_[51525]_  = \new_[51524]_  & \new_[51517]_ ;
  assign \new_[51528]_  = ~A265 & A236;
  assign \new_[51531]_  = ~A298 & ~A266;
  assign \new_[51532]_  = \new_[51531]_  & \new_[51528]_ ;
  assign \new_[51535]_  = ~A300 & A299;
  assign \new_[51538]_  = A302 & ~A301;
  assign \new_[51539]_  = \new_[51538]_  & \new_[51535]_ ;
  assign \new_[51540]_  = \new_[51539]_  & \new_[51532]_ ;
  assign \new_[51543]_  = ~A200 & A199;
  assign \new_[51546]_  = ~A202 & ~A201;
  assign \new_[51547]_  = \new_[51546]_  & \new_[51543]_ ;
  assign \new_[51550]_  = ~A232 & A203;
  assign \new_[51553]_  = A234 & A233;
  assign \new_[51554]_  = \new_[51553]_  & \new_[51550]_ ;
  assign \new_[51555]_  = \new_[51554]_  & \new_[51547]_ ;
  assign \new_[51558]_  = A267 & A235;
  assign \new_[51561]_  = A269 & ~A268;
  assign \new_[51562]_  = \new_[51561]_  & \new_[51558]_ ;
  assign \new_[51565]_  = ~A299 & A298;
  assign \new_[51568]_  = A301 & A300;
  assign \new_[51569]_  = \new_[51568]_  & \new_[51565]_ ;
  assign \new_[51570]_  = \new_[51569]_  & \new_[51562]_ ;
  assign \new_[51573]_  = ~A200 & A199;
  assign \new_[51576]_  = ~A202 & ~A201;
  assign \new_[51577]_  = \new_[51576]_  & \new_[51573]_ ;
  assign \new_[51580]_  = ~A232 & A203;
  assign \new_[51583]_  = A234 & A233;
  assign \new_[51584]_  = \new_[51583]_  & \new_[51580]_ ;
  assign \new_[51585]_  = \new_[51584]_  & \new_[51577]_ ;
  assign \new_[51588]_  = A267 & A235;
  assign \new_[51591]_  = A269 & ~A268;
  assign \new_[51592]_  = \new_[51591]_  & \new_[51588]_ ;
  assign \new_[51595]_  = ~A299 & A298;
  assign \new_[51598]_  = ~A302 & A300;
  assign \new_[51599]_  = \new_[51598]_  & \new_[51595]_ ;
  assign \new_[51600]_  = \new_[51599]_  & \new_[51592]_ ;
  assign \new_[51603]_  = ~A200 & A199;
  assign \new_[51606]_  = ~A202 & ~A201;
  assign \new_[51607]_  = \new_[51606]_  & \new_[51603]_ ;
  assign \new_[51610]_  = ~A232 & A203;
  assign \new_[51613]_  = A234 & A233;
  assign \new_[51614]_  = \new_[51613]_  & \new_[51610]_ ;
  assign \new_[51615]_  = \new_[51614]_  & \new_[51607]_ ;
  assign \new_[51618]_  = A267 & A235;
  assign \new_[51621]_  = A269 & ~A268;
  assign \new_[51622]_  = \new_[51621]_  & \new_[51618]_ ;
  assign \new_[51625]_  = A299 & ~A298;
  assign \new_[51628]_  = A301 & A300;
  assign \new_[51629]_  = \new_[51628]_  & \new_[51625]_ ;
  assign \new_[51630]_  = \new_[51629]_  & \new_[51622]_ ;
  assign \new_[51633]_  = ~A200 & A199;
  assign \new_[51636]_  = ~A202 & ~A201;
  assign \new_[51637]_  = \new_[51636]_  & \new_[51633]_ ;
  assign \new_[51640]_  = ~A232 & A203;
  assign \new_[51643]_  = A234 & A233;
  assign \new_[51644]_  = \new_[51643]_  & \new_[51640]_ ;
  assign \new_[51645]_  = \new_[51644]_  & \new_[51637]_ ;
  assign \new_[51648]_  = A267 & A235;
  assign \new_[51651]_  = A269 & ~A268;
  assign \new_[51652]_  = \new_[51651]_  & \new_[51648]_ ;
  assign \new_[51655]_  = A299 & ~A298;
  assign \new_[51658]_  = ~A302 & A300;
  assign \new_[51659]_  = \new_[51658]_  & \new_[51655]_ ;
  assign \new_[51660]_  = \new_[51659]_  & \new_[51652]_ ;
  assign \new_[51663]_  = ~A200 & A199;
  assign \new_[51666]_  = ~A202 & ~A201;
  assign \new_[51667]_  = \new_[51666]_  & \new_[51663]_ ;
  assign \new_[51670]_  = ~A232 & A203;
  assign \new_[51673]_  = A234 & A233;
  assign \new_[51674]_  = \new_[51673]_  & \new_[51670]_ ;
  assign \new_[51675]_  = \new_[51674]_  & \new_[51667]_ ;
  assign \new_[51678]_  = ~A267 & A235;
  assign \new_[51681]_  = A298 & A268;
  assign \new_[51682]_  = \new_[51681]_  & \new_[51678]_ ;
  assign \new_[51685]_  = ~A300 & ~A299;
  assign \new_[51688]_  = A302 & ~A301;
  assign \new_[51689]_  = \new_[51688]_  & \new_[51685]_ ;
  assign \new_[51690]_  = \new_[51689]_  & \new_[51682]_ ;
  assign \new_[51693]_  = ~A200 & A199;
  assign \new_[51696]_  = ~A202 & ~A201;
  assign \new_[51697]_  = \new_[51696]_  & \new_[51693]_ ;
  assign \new_[51700]_  = ~A232 & A203;
  assign \new_[51703]_  = A234 & A233;
  assign \new_[51704]_  = \new_[51703]_  & \new_[51700]_ ;
  assign \new_[51705]_  = \new_[51704]_  & \new_[51697]_ ;
  assign \new_[51708]_  = ~A267 & A235;
  assign \new_[51711]_  = ~A298 & A268;
  assign \new_[51712]_  = \new_[51711]_  & \new_[51708]_ ;
  assign \new_[51715]_  = ~A300 & A299;
  assign \new_[51718]_  = A302 & ~A301;
  assign \new_[51719]_  = \new_[51718]_  & \new_[51715]_ ;
  assign \new_[51720]_  = \new_[51719]_  & \new_[51712]_ ;
  assign \new_[51723]_  = ~A200 & A199;
  assign \new_[51726]_  = ~A202 & ~A201;
  assign \new_[51727]_  = \new_[51726]_  & \new_[51723]_ ;
  assign \new_[51730]_  = ~A232 & A203;
  assign \new_[51733]_  = A234 & A233;
  assign \new_[51734]_  = \new_[51733]_  & \new_[51730]_ ;
  assign \new_[51735]_  = \new_[51734]_  & \new_[51727]_ ;
  assign \new_[51738]_  = ~A267 & A235;
  assign \new_[51741]_  = A298 & ~A269;
  assign \new_[51742]_  = \new_[51741]_  & \new_[51738]_ ;
  assign \new_[51745]_  = ~A300 & ~A299;
  assign \new_[51748]_  = A302 & ~A301;
  assign \new_[51749]_  = \new_[51748]_  & \new_[51745]_ ;
  assign \new_[51750]_  = \new_[51749]_  & \new_[51742]_ ;
  assign \new_[51753]_  = ~A200 & A199;
  assign \new_[51756]_  = ~A202 & ~A201;
  assign \new_[51757]_  = \new_[51756]_  & \new_[51753]_ ;
  assign \new_[51760]_  = ~A232 & A203;
  assign \new_[51763]_  = A234 & A233;
  assign \new_[51764]_  = \new_[51763]_  & \new_[51760]_ ;
  assign \new_[51765]_  = \new_[51764]_  & \new_[51757]_ ;
  assign \new_[51768]_  = ~A267 & A235;
  assign \new_[51771]_  = ~A298 & ~A269;
  assign \new_[51772]_  = \new_[51771]_  & \new_[51768]_ ;
  assign \new_[51775]_  = ~A300 & A299;
  assign \new_[51778]_  = A302 & ~A301;
  assign \new_[51779]_  = \new_[51778]_  & \new_[51775]_ ;
  assign \new_[51780]_  = \new_[51779]_  & \new_[51772]_ ;
  assign \new_[51783]_  = ~A200 & A199;
  assign \new_[51786]_  = ~A202 & ~A201;
  assign \new_[51787]_  = \new_[51786]_  & \new_[51783]_ ;
  assign \new_[51790]_  = ~A232 & A203;
  assign \new_[51793]_  = A234 & A233;
  assign \new_[51794]_  = \new_[51793]_  & \new_[51790]_ ;
  assign \new_[51795]_  = \new_[51794]_  & \new_[51787]_ ;
  assign \new_[51798]_  = A265 & A235;
  assign \new_[51801]_  = A298 & A266;
  assign \new_[51802]_  = \new_[51801]_  & \new_[51798]_ ;
  assign \new_[51805]_  = ~A300 & ~A299;
  assign \new_[51808]_  = A302 & ~A301;
  assign \new_[51809]_  = \new_[51808]_  & \new_[51805]_ ;
  assign \new_[51810]_  = \new_[51809]_  & \new_[51802]_ ;
  assign \new_[51813]_  = ~A200 & A199;
  assign \new_[51816]_  = ~A202 & ~A201;
  assign \new_[51817]_  = \new_[51816]_  & \new_[51813]_ ;
  assign \new_[51820]_  = ~A232 & A203;
  assign \new_[51823]_  = A234 & A233;
  assign \new_[51824]_  = \new_[51823]_  & \new_[51820]_ ;
  assign \new_[51825]_  = \new_[51824]_  & \new_[51817]_ ;
  assign \new_[51828]_  = A265 & A235;
  assign \new_[51831]_  = ~A298 & A266;
  assign \new_[51832]_  = \new_[51831]_  & \new_[51828]_ ;
  assign \new_[51835]_  = ~A300 & A299;
  assign \new_[51838]_  = A302 & ~A301;
  assign \new_[51839]_  = \new_[51838]_  & \new_[51835]_ ;
  assign \new_[51840]_  = \new_[51839]_  & \new_[51832]_ ;
  assign \new_[51843]_  = ~A200 & A199;
  assign \new_[51846]_  = ~A202 & ~A201;
  assign \new_[51847]_  = \new_[51846]_  & \new_[51843]_ ;
  assign \new_[51850]_  = ~A232 & A203;
  assign \new_[51853]_  = A234 & A233;
  assign \new_[51854]_  = \new_[51853]_  & \new_[51850]_ ;
  assign \new_[51855]_  = \new_[51854]_  & \new_[51847]_ ;
  assign \new_[51858]_  = ~A265 & A235;
  assign \new_[51861]_  = A298 & ~A266;
  assign \new_[51862]_  = \new_[51861]_  & \new_[51858]_ ;
  assign \new_[51865]_  = ~A300 & ~A299;
  assign \new_[51868]_  = A302 & ~A301;
  assign \new_[51869]_  = \new_[51868]_  & \new_[51865]_ ;
  assign \new_[51870]_  = \new_[51869]_  & \new_[51862]_ ;
  assign \new_[51873]_  = ~A200 & A199;
  assign \new_[51876]_  = ~A202 & ~A201;
  assign \new_[51877]_  = \new_[51876]_  & \new_[51873]_ ;
  assign \new_[51880]_  = ~A232 & A203;
  assign \new_[51883]_  = A234 & A233;
  assign \new_[51884]_  = \new_[51883]_  & \new_[51880]_ ;
  assign \new_[51885]_  = \new_[51884]_  & \new_[51877]_ ;
  assign \new_[51888]_  = ~A265 & A235;
  assign \new_[51891]_  = ~A298 & ~A266;
  assign \new_[51892]_  = \new_[51891]_  & \new_[51888]_ ;
  assign \new_[51895]_  = ~A300 & A299;
  assign \new_[51898]_  = A302 & ~A301;
  assign \new_[51899]_  = \new_[51898]_  & \new_[51895]_ ;
  assign \new_[51900]_  = \new_[51899]_  & \new_[51892]_ ;
  assign \new_[51903]_  = ~A200 & A199;
  assign \new_[51906]_  = ~A202 & ~A201;
  assign \new_[51907]_  = \new_[51906]_  & \new_[51903]_ ;
  assign \new_[51910]_  = ~A232 & A203;
  assign \new_[51913]_  = A234 & A233;
  assign \new_[51914]_  = \new_[51913]_  & \new_[51910]_ ;
  assign \new_[51915]_  = \new_[51914]_  & \new_[51907]_ ;
  assign \new_[51918]_  = A267 & ~A236;
  assign \new_[51921]_  = A269 & ~A268;
  assign \new_[51922]_  = \new_[51921]_  & \new_[51918]_ ;
  assign \new_[51925]_  = ~A299 & A298;
  assign \new_[51928]_  = A301 & A300;
  assign \new_[51929]_  = \new_[51928]_  & \new_[51925]_ ;
  assign \new_[51930]_  = \new_[51929]_  & \new_[51922]_ ;
  assign \new_[51933]_  = ~A200 & A199;
  assign \new_[51936]_  = ~A202 & ~A201;
  assign \new_[51937]_  = \new_[51936]_  & \new_[51933]_ ;
  assign \new_[51940]_  = ~A232 & A203;
  assign \new_[51943]_  = A234 & A233;
  assign \new_[51944]_  = \new_[51943]_  & \new_[51940]_ ;
  assign \new_[51945]_  = \new_[51944]_  & \new_[51937]_ ;
  assign \new_[51948]_  = A267 & ~A236;
  assign \new_[51951]_  = A269 & ~A268;
  assign \new_[51952]_  = \new_[51951]_  & \new_[51948]_ ;
  assign \new_[51955]_  = ~A299 & A298;
  assign \new_[51958]_  = ~A302 & A300;
  assign \new_[51959]_  = \new_[51958]_  & \new_[51955]_ ;
  assign \new_[51960]_  = \new_[51959]_  & \new_[51952]_ ;
  assign \new_[51963]_  = ~A200 & A199;
  assign \new_[51966]_  = ~A202 & ~A201;
  assign \new_[51967]_  = \new_[51966]_  & \new_[51963]_ ;
  assign \new_[51970]_  = ~A232 & A203;
  assign \new_[51973]_  = A234 & A233;
  assign \new_[51974]_  = \new_[51973]_  & \new_[51970]_ ;
  assign \new_[51975]_  = \new_[51974]_  & \new_[51967]_ ;
  assign \new_[51978]_  = A267 & ~A236;
  assign \new_[51981]_  = A269 & ~A268;
  assign \new_[51982]_  = \new_[51981]_  & \new_[51978]_ ;
  assign \new_[51985]_  = A299 & ~A298;
  assign \new_[51988]_  = A301 & A300;
  assign \new_[51989]_  = \new_[51988]_  & \new_[51985]_ ;
  assign \new_[51990]_  = \new_[51989]_  & \new_[51982]_ ;
  assign \new_[51993]_  = ~A200 & A199;
  assign \new_[51996]_  = ~A202 & ~A201;
  assign \new_[51997]_  = \new_[51996]_  & \new_[51993]_ ;
  assign \new_[52000]_  = ~A232 & A203;
  assign \new_[52003]_  = A234 & A233;
  assign \new_[52004]_  = \new_[52003]_  & \new_[52000]_ ;
  assign \new_[52005]_  = \new_[52004]_  & \new_[51997]_ ;
  assign \new_[52008]_  = A267 & ~A236;
  assign \new_[52011]_  = A269 & ~A268;
  assign \new_[52012]_  = \new_[52011]_  & \new_[52008]_ ;
  assign \new_[52015]_  = A299 & ~A298;
  assign \new_[52018]_  = ~A302 & A300;
  assign \new_[52019]_  = \new_[52018]_  & \new_[52015]_ ;
  assign \new_[52020]_  = \new_[52019]_  & \new_[52012]_ ;
  assign \new_[52023]_  = ~A200 & A199;
  assign \new_[52026]_  = ~A202 & ~A201;
  assign \new_[52027]_  = \new_[52026]_  & \new_[52023]_ ;
  assign \new_[52030]_  = ~A232 & A203;
  assign \new_[52033]_  = A234 & A233;
  assign \new_[52034]_  = \new_[52033]_  & \new_[52030]_ ;
  assign \new_[52035]_  = \new_[52034]_  & \new_[52027]_ ;
  assign \new_[52038]_  = ~A267 & ~A236;
  assign \new_[52041]_  = A298 & A268;
  assign \new_[52042]_  = \new_[52041]_  & \new_[52038]_ ;
  assign \new_[52045]_  = ~A300 & ~A299;
  assign \new_[52048]_  = A302 & ~A301;
  assign \new_[52049]_  = \new_[52048]_  & \new_[52045]_ ;
  assign \new_[52050]_  = \new_[52049]_  & \new_[52042]_ ;
  assign \new_[52053]_  = ~A200 & A199;
  assign \new_[52056]_  = ~A202 & ~A201;
  assign \new_[52057]_  = \new_[52056]_  & \new_[52053]_ ;
  assign \new_[52060]_  = ~A232 & A203;
  assign \new_[52063]_  = A234 & A233;
  assign \new_[52064]_  = \new_[52063]_  & \new_[52060]_ ;
  assign \new_[52065]_  = \new_[52064]_  & \new_[52057]_ ;
  assign \new_[52068]_  = ~A267 & ~A236;
  assign \new_[52071]_  = ~A298 & A268;
  assign \new_[52072]_  = \new_[52071]_  & \new_[52068]_ ;
  assign \new_[52075]_  = ~A300 & A299;
  assign \new_[52078]_  = A302 & ~A301;
  assign \new_[52079]_  = \new_[52078]_  & \new_[52075]_ ;
  assign \new_[52080]_  = \new_[52079]_  & \new_[52072]_ ;
  assign \new_[52083]_  = ~A200 & A199;
  assign \new_[52086]_  = ~A202 & ~A201;
  assign \new_[52087]_  = \new_[52086]_  & \new_[52083]_ ;
  assign \new_[52090]_  = ~A232 & A203;
  assign \new_[52093]_  = A234 & A233;
  assign \new_[52094]_  = \new_[52093]_  & \new_[52090]_ ;
  assign \new_[52095]_  = \new_[52094]_  & \new_[52087]_ ;
  assign \new_[52098]_  = ~A267 & ~A236;
  assign \new_[52101]_  = A298 & ~A269;
  assign \new_[52102]_  = \new_[52101]_  & \new_[52098]_ ;
  assign \new_[52105]_  = ~A300 & ~A299;
  assign \new_[52108]_  = A302 & ~A301;
  assign \new_[52109]_  = \new_[52108]_  & \new_[52105]_ ;
  assign \new_[52110]_  = \new_[52109]_  & \new_[52102]_ ;
  assign \new_[52113]_  = ~A200 & A199;
  assign \new_[52116]_  = ~A202 & ~A201;
  assign \new_[52117]_  = \new_[52116]_  & \new_[52113]_ ;
  assign \new_[52120]_  = ~A232 & A203;
  assign \new_[52123]_  = A234 & A233;
  assign \new_[52124]_  = \new_[52123]_  & \new_[52120]_ ;
  assign \new_[52125]_  = \new_[52124]_  & \new_[52117]_ ;
  assign \new_[52128]_  = ~A267 & ~A236;
  assign \new_[52131]_  = ~A298 & ~A269;
  assign \new_[52132]_  = \new_[52131]_  & \new_[52128]_ ;
  assign \new_[52135]_  = ~A300 & A299;
  assign \new_[52138]_  = A302 & ~A301;
  assign \new_[52139]_  = \new_[52138]_  & \new_[52135]_ ;
  assign \new_[52140]_  = \new_[52139]_  & \new_[52132]_ ;
  assign \new_[52143]_  = ~A200 & A199;
  assign \new_[52146]_  = ~A202 & ~A201;
  assign \new_[52147]_  = \new_[52146]_  & \new_[52143]_ ;
  assign \new_[52150]_  = ~A232 & A203;
  assign \new_[52153]_  = A234 & A233;
  assign \new_[52154]_  = \new_[52153]_  & \new_[52150]_ ;
  assign \new_[52155]_  = \new_[52154]_  & \new_[52147]_ ;
  assign \new_[52158]_  = A265 & ~A236;
  assign \new_[52161]_  = A298 & A266;
  assign \new_[52162]_  = \new_[52161]_  & \new_[52158]_ ;
  assign \new_[52165]_  = ~A300 & ~A299;
  assign \new_[52168]_  = A302 & ~A301;
  assign \new_[52169]_  = \new_[52168]_  & \new_[52165]_ ;
  assign \new_[52170]_  = \new_[52169]_  & \new_[52162]_ ;
  assign \new_[52173]_  = ~A200 & A199;
  assign \new_[52176]_  = ~A202 & ~A201;
  assign \new_[52177]_  = \new_[52176]_  & \new_[52173]_ ;
  assign \new_[52180]_  = ~A232 & A203;
  assign \new_[52183]_  = A234 & A233;
  assign \new_[52184]_  = \new_[52183]_  & \new_[52180]_ ;
  assign \new_[52185]_  = \new_[52184]_  & \new_[52177]_ ;
  assign \new_[52188]_  = A265 & ~A236;
  assign \new_[52191]_  = ~A298 & A266;
  assign \new_[52192]_  = \new_[52191]_  & \new_[52188]_ ;
  assign \new_[52195]_  = ~A300 & A299;
  assign \new_[52198]_  = A302 & ~A301;
  assign \new_[52199]_  = \new_[52198]_  & \new_[52195]_ ;
  assign \new_[52200]_  = \new_[52199]_  & \new_[52192]_ ;
  assign \new_[52203]_  = ~A200 & A199;
  assign \new_[52206]_  = ~A202 & ~A201;
  assign \new_[52207]_  = \new_[52206]_  & \new_[52203]_ ;
  assign \new_[52210]_  = ~A232 & A203;
  assign \new_[52213]_  = A234 & A233;
  assign \new_[52214]_  = \new_[52213]_  & \new_[52210]_ ;
  assign \new_[52215]_  = \new_[52214]_  & \new_[52207]_ ;
  assign \new_[52218]_  = ~A265 & ~A236;
  assign \new_[52221]_  = A298 & ~A266;
  assign \new_[52222]_  = \new_[52221]_  & \new_[52218]_ ;
  assign \new_[52225]_  = ~A300 & ~A299;
  assign \new_[52228]_  = A302 & ~A301;
  assign \new_[52229]_  = \new_[52228]_  & \new_[52225]_ ;
  assign \new_[52230]_  = \new_[52229]_  & \new_[52222]_ ;
  assign \new_[52233]_  = ~A200 & A199;
  assign \new_[52236]_  = ~A202 & ~A201;
  assign \new_[52237]_  = \new_[52236]_  & \new_[52233]_ ;
  assign \new_[52240]_  = ~A232 & A203;
  assign \new_[52243]_  = A234 & A233;
  assign \new_[52244]_  = \new_[52243]_  & \new_[52240]_ ;
  assign \new_[52245]_  = \new_[52244]_  & \new_[52237]_ ;
  assign \new_[52248]_  = ~A265 & ~A236;
  assign \new_[52251]_  = ~A298 & ~A266;
  assign \new_[52252]_  = \new_[52251]_  & \new_[52248]_ ;
  assign \new_[52255]_  = ~A300 & A299;
  assign \new_[52258]_  = A302 & ~A301;
  assign \new_[52259]_  = \new_[52258]_  & \new_[52255]_ ;
  assign \new_[52260]_  = \new_[52259]_  & \new_[52252]_ ;
  assign \new_[52263]_  = ~A200 & A199;
  assign \new_[52266]_  = ~A202 & ~A201;
  assign \new_[52267]_  = \new_[52266]_  & \new_[52263]_ ;
  assign \new_[52270]_  = ~A232 & A203;
  assign \new_[52273]_  = ~A234 & A233;
  assign \new_[52274]_  = \new_[52273]_  & \new_[52270]_ ;
  assign \new_[52275]_  = \new_[52274]_  & \new_[52267]_ ;
  assign \new_[52278]_  = A236 & ~A235;
  assign \new_[52281]_  = A268 & ~A267;
  assign \new_[52282]_  = \new_[52281]_  & \new_[52278]_ ;
  assign \new_[52285]_  = ~A299 & A298;
  assign \new_[52288]_  = A301 & A300;
  assign \new_[52289]_  = \new_[52288]_  & \new_[52285]_ ;
  assign \new_[52290]_  = \new_[52289]_  & \new_[52282]_ ;
  assign \new_[52293]_  = ~A200 & A199;
  assign \new_[52296]_  = ~A202 & ~A201;
  assign \new_[52297]_  = \new_[52296]_  & \new_[52293]_ ;
  assign \new_[52300]_  = ~A232 & A203;
  assign \new_[52303]_  = ~A234 & A233;
  assign \new_[52304]_  = \new_[52303]_  & \new_[52300]_ ;
  assign \new_[52305]_  = \new_[52304]_  & \new_[52297]_ ;
  assign \new_[52308]_  = A236 & ~A235;
  assign \new_[52311]_  = A268 & ~A267;
  assign \new_[52312]_  = \new_[52311]_  & \new_[52308]_ ;
  assign \new_[52315]_  = ~A299 & A298;
  assign \new_[52318]_  = ~A302 & A300;
  assign \new_[52319]_  = \new_[52318]_  & \new_[52315]_ ;
  assign \new_[52320]_  = \new_[52319]_  & \new_[52312]_ ;
  assign \new_[52323]_  = ~A200 & A199;
  assign \new_[52326]_  = ~A202 & ~A201;
  assign \new_[52327]_  = \new_[52326]_  & \new_[52323]_ ;
  assign \new_[52330]_  = ~A232 & A203;
  assign \new_[52333]_  = ~A234 & A233;
  assign \new_[52334]_  = \new_[52333]_  & \new_[52330]_ ;
  assign \new_[52335]_  = \new_[52334]_  & \new_[52327]_ ;
  assign \new_[52338]_  = A236 & ~A235;
  assign \new_[52341]_  = A268 & ~A267;
  assign \new_[52342]_  = \new_[52341]_  & \new_[52338]_ ;
  assign \new_[52345]_  = A299 & ~A298;
  assign \new_[52348]_  = A301 & A300;
  assign \new_[52349]_  = \new_[52348]_  & \new_[52345]_ ;
  assign \new_[52350]_  = \new_[52349]_  & \new_[52342]_ ;
  assign \new_[52353]_  = ~A200 & A199;
  assign \new_[52356]_  = ~A202 & ~A201;
  assign \new_[52357]_  = \new_[52356]_  & \new_[52353]_ ;
  assign \new_[52360]_  = ~A232 & A203;
  assign \new_[52363]_  = ~A234 & A233;
  assign \new_[52364]_  = \new_[52363]_  & \new_[52360]_ ;
  assign \new_[52365]_  = \new_[52364]_  & \new_[52357]_ ;
  assign \new_[52368]_  = A236 & ~A235;
  assign \new_[52371]_  = A268 & ~A267;
  assign \new_[52372]_  = \new_[52371]_  & \new_[52368]_ ;
  assign \new_[52375]_  = A299 & ~A298;
  assign \new_[52378]_  = ~A302 & A300;
  assign \new_[52379]_  = \new_[52378]_  & \new_[52375]_ ;
  assign \new_[52380]_  = \new_[52379]_  & \new_[52372]_ ;
  assign \new_[52383]_  = ~A200 & A199;
  assign \new_[52386]_  = ~A202 & ~A201;
  assign \new_[52387]_  = \new_[52386]_  & \new_[52383]_ ;
  assign \new_[52390]_  = ~A232 & A203;
  assign \new_[52393]_  = ~A234 & A233;
  assign \new_[52394]_  = \new_[52393]_  & \new_[52390]_ ;
  assign \new_[52395]_  = \new_[52394]_  & \new_[52387]_ ;
  assign \new_[52398]_  = A236 & ~A235;
  assign \new_[52401]_  = ~A269 & ~A267;
  assign \new_[52402]_  = \new_[52401]_  & \new_[52398]_ ;
  assign \new_[52405]_  = ~A299 & A298;
  assign \new_[52408]_  = A301 & A300;
  assign \new_[52409]_  = \new_[52408]_  & \new_[52405]_ ;
  assign \new_[52410]_  = \new_[52409]_  & \new_[52402]_ ;
  assign \new_[52413]_  = ~A200 & A199;
  assign \new_[52416]_  = ~A202 & ~A201;
  assign \new_[52417]_  = \new_[52416]_  & \new_[52413]_ ;
  assign \new_[52420]_  = ~A232 & A203;
  assign \new_[52423]_  = ~A234 & A233;
  assign \new_[52424]_  = \new_[52423]_  & \new_[52420]_ ;
  assign \new_[52425]_  = \new_[52424]_  & \new_[52417]_ ;
  assign \new_[52428]_  = A236 & ~A235;
  assign \new_[52431]_  = ~A269 & ~A267;
  assign \new_[52432]_  = \new_[52431]_  & \new_[52428]_ ;
  assign \new_[52435]_  = ~A299 & A298;
  assign \new_[52438]_  = ~A302 & A300;
  assign \new_[52439]_  = \new_[52438]_  & \new_[52435]_ ;
  assign \new_[52440]_  = \new_[52439]_  & \new_[52432]_ ;
  assign \new_[52443]_  = ~A200 & A199;
  assign \new_[52446]_  = ~A202 & ~A201;
  assign \new_[52447]_  = \new_[52446]_  & \new_[52443]_ ;
  assign \new_[52450]_  = ~A232 & A203;
  assign \new_[52453]_  = ~A234 & A233;
  assign \new_[52454]_  = \new_[52453]_  & \new_[52450]_ ;
  assign \new_[52455]_  = \new_[52454]_  & \new_[52447]_ ;
  assign \new_[52458]_  = A236 & ~A235;
  assign \new_[52461]_  = ~A269 & ~A267;
  assign \new_[52462]_  = \new_[52461]_  & \new_[52458]_ ;
  assign \new_[52465]_  = A299 & ~A298;
  assign \new_[52468]_  = A301 & A300;
  assign \new_[52469]_  = \new_[52468]_  & \new_[52465]_ ;
  assign \new_[52470]_  = \new_[52469]_  & \new_[52462]_ ;
  assign \new_[52473]_  = ~A200 & A199;
  assign \new_[52476]_  = ~A202 & ~A201;
  assign \new_[52477]_  = \new_[52476]_  & \new_[52473]_ ;
  assign \new_[52480]_  = ~A232 & A203;
  assign \new_[52483]_  = ~A234 & A233;
  assign \new_[52484]_  = \new_[52483]_  & \new_[52480]_ ;
  assign \new_[52485]_  = \new_[52484]_  & \new_[52477]_ ;
  assign \new_[52488]_  = A236 & ~A235;
  assign \new_[52491]_  = ~A269 & ~A267;
  assign \new_[52492]_  = \new_[52491]_  & \new_[52488]_ ;
  assign \new_[52495]_  = A299 & ~A298;
  assign \new_[52498]_  = ~A302 & A300;
  assign \new_[52499]_  = \new_[52498]_  & \new_[52495]_ ;
  assign \new_[52500]_  = \new_[52499]_  & \new_[52492]_ ;
  assign \new_[52503]_  = ~A200 & A199;
  assign \new_[52506]_  = ~A202 & ~A201;
  assign \new_[52507]_  = \new_[52506]_  & \new_[52503]_ ;
  assign \new_[52510]_  = ~A232 & A203;
  assign \new_[52513]_  = ~A234 & A233;
  assign \new_[52514]_  = \new_[52513]_  & \new_[52510]_ ;
  assign \new_[52515]_  = \new_[52514]_  & \new_[52507]_ ;
  assign \new_[52518]_  = A236 & ~A235;
  assign \new_[52521]_  = A266 & A265;
  assign \new_[52522]_  = \new_[52521]_  & \new_[52518]_ ;
  assign \new_[52525]_  = ~A299 & A298;
  assign \new_[52528]_  = A301 & A300;
  assign \new_[52529]_  = \new_[52528]_  & \new_[52525]_ ;
  assign \new_[52530]_  = \new_[52529]_  & \new_[52522]_ ;
  assign \new_[52533]_  = ~A200 & A199;
  assign \new_[52536]_  = ~A202 & ~A201;
  assign \new_[52537]_  = \new_[52536]_  & \new_[52533]_ ;
  assign \new_[52540]_  = ~A232 & A203;
  assign \new_[52543]_  = ~A234 & A233;
  assign \new_[52544]_  = \new_[52543]_  & \new_[52540]_ ;
  assign \new_[52545]_  = \new_[52544]_  & \new_[52537]_ ;
  assign \new_[52548]_  = A236 & ~A235;
  assign \new_[52551]_  = A266 & A265;
  assign \new_[52552]_  = \new_[52551]_  & \new_[52548]_ ;
  assign \new_[52555]_  = ~A299 & A298;
  assign \new_[52558]_  = ~A302 & A300;
  assign \new_[52559]_  = \new_[52558]_  & \new_[52555]_ ;
  assign \new_[52560]_  = \new_[52559]_  & \new_[52552]_ ;
  assign \new_[52563]_  = ~A200 & A199;
  assign \new_[52566]_  = ~A202 & ~A201;
  assign \new_[52567]_  = \new_[52566]_  & \new_[52563]_ ;
  assign \new_[52570]_  = ~A232 & A203;
  assign \new_[52573]_  = ~A234 & A233;
  assign \new_[52574]_  = \new_[52573]_  & \new_[52570]_ ;
  assign \new_[52575]_  = \new_[52574]_  & \new_[52567]_ ;
  assign \new_[52578]_  = A236 & ~A235;
  assign \new_[52581]_  = A266 & A265;
  assign \new_[52582]_  = \new_[52581]_  & \new_[52578]_ ;
  assign \new_[52585]_  = A299 & ~A298;
  assign \new_[52588]_  = A301 & A300;
  assign \new_[52589]_  = \new_[52588]_  & \new_[52585]_ ;
  assign \new_[52590]_  = \new_[52589]_  & \new_[52582]_ ;
  assign \new_[52593]_  = ~A200 & A199;
  assign \new_[52596]_  = ~A202 & ~A201;
  assign \new_[52597]_  = \new_[52596]_  & \new_[52593]_ ;
  assign \new_[52600]_  = ~A232 & A203;
  assign \new_[52603]_  = ~A234 & A233;
  assign \new_[52604]_  = \new_[52603]_  & \new_[52600]_ ;
  assign \new_[52605]_  = \new_[52604]_  & \new_[52597]_ ;
  assign \new_[52608]_  = A236 & ~A235;
  assign \new_[52611]_  = A266 & A265;
  assign \new_[52612]_  = \new_[52611]_  & \new_[52608]_ ;
  assign \new_[52615]_  = A299 & ~A298;
  assign \new_[52618]_  = ~A302 & A300;
  assign \new_[52619]_  = \new_[52618]_  & \new_[52615]_ ;
  assign \new_[52620]_  = \new_[52619]_  & \new_[52612]_ ;
  assign \new_[52623]_  = ~A200 & A199;
  assign \new_[52626]_  = ~A202 & ~A201;
  assign \new_[52627]_  = \new_[52626]_  & \new_[52623]_ ;
  assign \new_[52630]_  = ~A232 & A203;
  assign \new_[52633]_  = ~A234 & A233;
  assign \new_[52634]_  = \new_[52633]_  & \new_[52630]_ ;
  assign \new_[52635]_  = \new_[52634]_  & \new_[52627]_ ;
  assign \new_[52638]_  = A236 & ~A235;
  assign \new_[52641]_  = ~A266 & ~A265;
  assign \new_[52642]_  = \new_[52641]_  & \new_[52638]_ ;
  assign \new_[52645]_  = ~A299 & A298;
  assign \new_[52648]_  = A301 & A300;
  assign \new_[52649]_  = \new_[52648]_  & \new_[52645]_ ;
  assign \new_[52650]_  = \new_[52649]_  & \new_[52642]_ ;
  assign \new_[52653]_  = ~A200 & A199;
  assign \new_[52656]_  = ~A202 & ~A201;
  assign \new_[52657]_  = \new_[52656]_  & \new_[52653]_ ;
  assign \new_[52660]_  = ~A232 & A203;
  assign \new_[52663]_  = ~A234 & A233;
  assign \new_[52664]_  = \new_[52663]_  & \new_[52660]_ ;
  assign \new_[52665]_  = \new_[52664]_  & \new_[52657]_ ;
  assign \new_[52668]_  = A236 & ~A235;
  assign \new_[52671]_  = ~A266 & ~A265;
  assign \new_[52672]_  = \new_[52671]_  & \new_[52668]_ ;
  assign \new_[52675]_  = ~A299 & A298;
  assign \new_[52678]_  = ~A302 & A300;
  assign \new_[52679]_  = \new_[52678]_  & \new_[52675]_ ;
  assign \new_[52680]_  = \new_[52679]_  & \new_[52672]_ ;
  assign \new_[52683]_  = ~A200 & A199;
  assign \new_[52686]_  = ~A202 & ~A201;
  assign \new_[52687]_  = \new_[52686]_  & \new_[52683]_ ;
  assign \new_[52690]_  = ~A232 & A203;
  assign \new_[52693]_  = ~A234 & A233;
  assign \new_[52694]_  = \new_[52693]_  & \new_[52690]_ ;
  assign \new_[52695]_  = \new_[52694]_  & \new_[52687]_ ;
  assign \new_[52698]_  = A236 & ~A235;
  assign \new_[52701]_  = ~A266 & ~A265;
  assign \new_[52702]_  = \new_[52701]_  & \new_[52698]_ ;
  assign \new_[52705]_  = A299 & ~A298;
  assign \new_[52708]_  = A301 & A300;
  assign \new_[52709]_  = \new_[52708]_  & \new_[52705]_ ;
  assign \new_[52710]_  = \new_[52709]_  & \new_[52702]_ ;
  assign \new_[52713]_  = ~A200 & A199;
  assign \new_[52716]_  = ~A202 & ~A201;
  assign \new_[52717]_  = \new_[52716]_  & \new_[52713]_ ;
  assign \new_[52720]_  = ~A232 & A203;
  assign \new_[52723]_  = ~A234 & A233;
  assign \new_[52724]_  = \new_[52723]_  & \new_[52720]_ ;
  assign \new_[52725]_  = \new_[52724]_  & \new_[52717]_ ;
  assign \new_[52728]_  = A236 & ~A235;
  assign \new_[52731]_  = ~A266 & ~A265;
  assign \new_[52732]_  = \new_[52731]_  & \new_[52728]_ ;
  assign \new_[52735]_  = A299 & ~A298;
  assign \new_[52738]_  = ~A302 & A300;
  assign \new_[52739]_  = \new_[52738]_  & \new_[52735]_ ;
  assign \new_[52740]_  = \new_[52739]_  & \new_[52732]_ ;
  assign \new_[52743]_  = ~A200 & A199;
  assign \new_[52746]_  = ~A202 & ~A201;
  assign \new_[52747]_  = \new_[52746]_  & \new_[52743]_ ;
  assign \new_[52750]_  = A232 & A203;
  assign \new_[52753]_  = A234 & ~A233;
  assign \new_[52754]_  = \new_[52753]_  & \new_[52750]_ ;
  assign \new_[52755]_  = \new_[52754]_  & \new_[52747]_ ;
  assign \new_[52758]_  = A267 & A235;
  assign \new_[52761]_  = A269 & ~A268;
  assign \new_[52762]_  = \new_[52761]_  & \new_[52758]_ ;
  assign \new_[52765]_  = ~A299 & A298;
  assign \new_[52768]_  = A301 & A300;
  assign \new_[52769]_  = \new_[52768]_  & \new_[52765]_ ;
  assign \new_[52770]_  = \new_[52769]_  & \new_[52762]_ ;
  assign \new_[52773]_  = ~A200 & A199;
  assign \new_[52776]_  = ~A202 & ~A201;
  assign \new_[52777]_  = \new_[52776]_  & \new_[52773]_ ;
  assign \new_[52780]_  = A232 & A203;
  assign \new_[52783]_  = A234 & ~A233;
  assign \new_[52784]_  = \new_[52783]_  & \new_[52780]_ ;
  assign \new_[52785]_  = \new_[52784]_  & \new_[52777]_ ;
  assign \new_[52788]_  = A267 & A235;
  assign \new_[52791]_  = A269 & ~A268;
  assign \new_[52792]_  = \new_[52791]_  & \new_[52788]_ ;
  assign \new_[52795]_  = ~A299 & A298;
  assign \new_[52798]_  = ~A302 & A300;
  assign \new_[52799]_  = \new_[52798]_  & \new_[52795]_ ;
  assign \new_[52800]_  = \new_[52799]_  & \new_[52792]_ ;
  assign \new_[52803]_  = ~A200 & A199;
  assign \new_[52806]_  = ~A202 & ~A201;
  assign \new_[52807]_  = \new_[52806]_  & \new_[52803]_ ;
  assign \new_[52810]_  = A232 & A203;
  assign \new_[52813]_  = A234 & ~A233;
  assign \new_[52814]_  = \new_[52813]_  & \new_[52810]_ ;
  assign \new_[52815]_  = \new_[52814]_  & \new_[52807]_ ;
  assign \new_[52818]_  = A267 & A235;
  assign \new_[52821]_  = A269 & ~A268;
  assign \new_[52822]_  = \new_[52821]_  & \new_[52818]_ ;
  assign \new_[52825]_  = A299 & ~A298;
  assign \new_[52828]_  = A301 & A300;
  assign \new_[52829]_  = \new_[52828]_  & \new_[52825]_ ;
  assign \new_[52830]_  = \new_[52829]_  & \new_[52822]_ ;
  assign \new_[52833]_  = ~A200 & A199;
  assign \new_[52836]_  = ~A202 & ~A201;
  assign \new_[52837]_  = \new_[52836]_  & \new_[52833]_ ;
  assign \new_[52840]_  = A232 & A203;
  assign \new_[52843]_  = A234 & ~A233;
  assign \new_[52844]_  = \new_[52843]_  & \new_[52840]_ ;
  assign \new_[52845]_  = \new_[52844]_  & \new_[52837]_ ;
  assign \new_[52848]_  = A267 & A235;
  assign \new_[52851]_  = A269 & ~A268;
  assign \new_[52852]_  = \new_[52851]_  & \new_[52848]_ ;
  assign \new_[52855]_  = A299 & ~A298;
  assign \new_[52858]_  = ~A302 & A300;
  assign \new_[52859]_  = \new_[52858]_  & \new_[52855]_ ;
  assign \new_[52860]_  = \new_[52859]_  & \new_[52852]_ ;
  assign \new_[52863]_  = ~A200 & A199;
  assign \new_[52866]_  = ~A202 & ~A201;
  assign \new_[52867]_  = \new_[52866]_  & \new_[52863]_ ;
  assign \new_[52870]_  = A232 & A203;
  assign \new_[52873]_  = A234 & ~A233;
  assign \new_[52874]_  = \new_[52873]_  & \new_[52870]_ ;
  assign \new_[52875]_  = \new_[52874]_  & \new_[52867]_ ;
  assign \new_[52878]_  = ~A267 & A235;
  assign \new_[52881]_  = A298 & A268;
  assign \new_[52882]_  = \new_[52881]_  & \new_[52878]_ ;
  assign \new_[52885]_  = ~A300 & ~A299;
  assign \new_[52888]_  = A302 & ~A301;
  assign \new_[52889]_  = \new_[52888]_  & \new_[52885]_ ;
  assign \new_[52890]_  = \new_[52889]_  & \new_[52882]_ ;
  assign \new_[52893]_  = ~A200 & A199;
  assign \new_[52896]_  = ~A202 & ~A201;
  assign \new_[52897]_  = \new_[52896]_  & \new_[52893]_ ;
  assign \new_[52900]_  = A232 & A203;
  assign \new_[52903]_  = A234 & ~A233;
  assign \new_[52904]_  = \new_[52903]_  & \new_[52900]_ ;
  assign \new_[52905]_  = \new_[52904]_  & \new_[52897]_ ;
  assign \new_[52908]_  = ~A267 & A235;
  assign \new_[52911]_  = ~A298 & A268;
  assign \new_[52912]_  = \new_[52911]_  & \new_[52908]_ ;
  assign \new_[52915]_  = ~A300 & A299;
  assign \new_[52918]_  = A302 & ~A301;
  assign \new_[52919]_  = \new_[52918]_  & \new_[52915]_ ;
  assign \new_[52920]_  = \new_[52919]_  & \new_[52912]_ ;
  assign \new_[52923]_  = ~A200 & A199;
  assign \new_[52926]_  = ~A202 & ~A201;
  assign \new_[52927]_  = \new_[52926]_  & \new_[52923]_ ;
  assign \new_[52930]_  = A232 & A203;
  assign \new_[52933]_  = A234 & ~A233;
  assign \new_[52934]_  = \new_[52933]_  & \new_[52930]_ ;
  assign \new_[52935]_  = \new_[52934]_  & \new_[52927]_ ;
  assign \new_[52938]_  = ~A267 & A235;
  assign \new_[52941]_  = A298 & ~A269;
  assign \new_[52942]_  = \new_[52941]_  & \new_[52938]_ ;
  assign \new_[52945]_  = ~A300 & ~A299;
  assign \new_[52948]_  = A302 & ~A301;
  assign \new_[52949]_  = \new_[52948]_  & \new_[52945]_ ;
  assign \new_[52950]_  = \new_[52949]_  & \new_[52942]_ ;
  assign \new_[52953]_  = ~A200 & A199;
  assign \new_[52956]_  = ~A202 & ~A201;
  assign \new_[52957]_  = \new_[52956]_  & \new_[52953]_ ;
  assign \new_[52960]_  = A232 & A203;
  assign \new_[52963]_  = A234 & ~A233;
  assign \new_[52964]_  = \new_[52963]_  & \new_[52960]_ ;
  assign \new_[52965]_  = \new_[52964]_  & \new_[52957]_ ;
  assign \new_[52968]_  = ~A267 & A235;
  assign \new_[52971]_  = ~A298 & ~A269;
  assign \new_[52972]_  = \new_[52971]_  & \new_[52968]_ ;
  assign \new_[52975]_  = ~A300 & A299;
  assign \new_[52978]_  = A302 & ~A301;
  assign \new_[52979]_  = \new_[52978]_  & \new_[52975]_ ;
  assign \new_[52980]_  = \new_[52979]_  & \new_[52972]_ ;
  assign \new_[52983]_  = ~A200 & A199;
  assign \new_[52986]_  = ~A202 & ~A201;
  assign \new_[52987]_  = \new_[52986]_  & \new_[52983]_ ;
  assign \new_[52990]_  = A232 & A203;
  assign \new_[52993]_  = A234 & ~A233;
  assign \new_[52994]_  = \new_[52993]_  & \new_[52990]_ ;
  assign \new_[52995]_  = \new_[52994]_  & \new_[52987]_ ;
  assign \new_[52998]_  = A265 & A235;
  assign \new_[53001]_  = A298 & A266;
  assign \new_[53002]_  = \new_[53001]_  & \new_[52998]_ ;
  assign \new_[53005]_  = ~A300 & ~A299;
  assign \new_[53008]_  = A302 & ~A301;
  assign \new_[53009]_  = \new_[53008]_  & \new_[53005]_ ;
  assign \new_[53010]_  = \new_[53009]_  & \new_[53002]_ ;
  assign \new_[53013]_  = ~A200 & A199;
  assign \new_[53016]_  = ~A202 & ~A201;
  assign \new_[53017]_  = \new_[53016]_  & \new_[53013]_ ;
  assign \new_[53020]_  = A232 & A203;
  assign \new_[53023]_  = A234 & ~A233;
  assign \new_[53024]_  = \new_[53023]_  & \new_[53020]_ ;
  assign \new_[53025]_  = \new_[53024]_  & \new_[53017]_ ;
  assign \new_[53028]_  = A265 & A235;
  assign \new_[53031]_  = ~A298 & A266;
  assign \new_[53032]_  = \new_[53031]_  & \new_[53028]_ ;
  assign \new_[53035]_  = ~A300 & A299;
  assign \new_[53038]_  = A302 & ~A301;
  assign \new_[53039]_  = \new_[53038]_  & \new_[53035]_ ;
  assign \new_[53040]_  = \new_[53039]_  & \new_[53032]_ ;
  assign \new_[53043]_  = ~A200 & A199;
  assign \new_[53046]_  = ~A202 & ~A201;
  assign \new_[53047]_  = \new_[53046]_  & \new_[53043]_ ;
  assign \new_[53050]_  = A232 & A203;
  assign \new_[53053]_  = A234 & ~A233;
  assign \new_[53054]_  = \new_[53053]_  & \new_[53050]_ ;
  assign \new_[53055]_  = \new_[53054]_  & \new_[53047]_ ;
  assign \new_[53058]_  = ~A265 & A235;
  assign \new_[53061]_  = A298 & ~A266;
  assign \new_[53062]_  = \new_[53061]_  & \new_[53058]_ ;
  assign \new_[53065]_  = ~A300 & ~A299;
  assign \new_[53068]_  = A302 & ~A301;
  assign \new_[53069]_  = \new_[53068]_  & \new_[53065]_ ;
  assign \new_[53070]_  = \new_[53069]_  & \new_[53062]_ ;
  assign \new_[53073]_  = ~A200 & A199;
  assign \new_[53076]_  = ~A202 & ~A201;
  assign \new_[53077]_  = \new_[53076]_  & \new_[53073]_ ;
  assign \new_[53080]_  = A232 & A203;
  assign \new_[53083]_  = A234 & ~A233;
  assign \new_[53084]_  = \new_[53083]_  & \new_[53080]_ ;
  assign \new_[53085]_  = \new_[53084]_  & \new_[53077]_ ;
  assign \new_[53088]_  = ~A265 & A235;
  assign \new_[53091]_  = ~A298 & ~A266;
  assign \new_[53092]_  = \new_[53091]_  & \new_[53088]_ ;
  assign \new_[53095]_  = ~A300 & A299;
  assign \new_[53098]_  = A302 & ~A301;
  assign \new_[53099]_  = \new_[53098]_  & \new_[53095]_ ;
  assign \new_[53100]_  = \new_[53099]_  & \new_[53092]_ ;
  assign \new_[53103]_  = ~A200 & A199;
  assign \new_[53106]_  = ~A202 & ~A201;
  assign \new_[53107]_  = \new_[53106]_  & \new_[53103]_ ;
  assign \new_[53110]_  = A232 & A203;
  assign \new_[53113]_  = A234 & ~A233;
  assign \new_[53114]_  = \new_[53113]_  & \new_[53110]_ ;
  assign \new_[53115]_  = \new_[53114]_  & \new_[53107]_ ;
  assign \new_[53118]_  = A267 & ~A236;
  assign \new_[53121]_  = A269 & ~A268;
  assign \new_[53122]_  = \new_[53121]_  & \new_[53118]_ ;
  assign \new_[53125]_  = ~A299 & A298;
  assign \new_[53128]_  = A301 & A300;
  assign \new_[53129]_  = \new_[53128]_  & \new_[53125]_ ;
  assign \new_[53130]_  = \new_[53129]_  & \new_[53122]_ ;
  assign \new_[53133]_  = ~A200 & A199;
  assign \new_[53136]_  = ~A202 & ~A201;
  assign \new_[53137]_  = \new_[53136]_  & \new_[53133]_ ;
  assign \new_[53140]_  = A232 & A203;
  assign \new_[53143]_  = A234 & ~A233;
  assign \new_[53144]_  = \new_[53143]_  & \new_[53140]_ ;
  assign \new_[53145]_  = \new_[53144]_  & \new_[53137]_ ;
  assign \new_[53148]_  = A267 & ~A236;
  assign \new_[53151]_  = A269 & ~A268;
  assign \new_[53152]_  = \new_[53151]_  & \new_[53148]_ ;
  assign \new_[53155]_  = ~A299 & A298;
  assign \new_[53158]_  = ~A302 & A300;
  assign \new_[53159]_  = \new_[53158]_  & \new_[53155]_ ;
  assign \new_[53160]_  = \new_[53159]_  & \new_[53152]_ ;
  assign \new_[53163]_  = ~A200 & A199;
  assign \new_[53166]_  = ~A202 & ~A201;
  assign \new_[53167]_  = \new_[53166]_  & \new_[53163]_ ;
  assign \new_[53170]_  = A232 & A203;
  assign \new_[53173]_  = A234 & ~A233;
  assign \new_[53174]_  = \new_[53173]_  & \new_[53170]_ ;
  assign \new_[53175]_  = \new_[53174]_  & \new_[53167]_ ;
  assign \new_[53178]_  = A267 & ~A236;
  assign \new_[53181]_  = A269 & ~A268;
  assign \new_[53182]_  = \new_[53181]_  & \new_[53178]_ ;
  assign \new_[53185]_  = A299 & ~A298;
  assign \new_[53188]_  = A301 & A300;
  assign \new_[53189]_  = \new_[53188]_  & \new_[53185]_ ;
  assign \new_[53190]_  = \new_[53189]_  & \new_[53182]_ ;
  assign \new_[53193]_  = ~A200 & A199;
  assign \new_[53196]_  = ~A202 & ~A201;
  assign \new_[53197]_  = \new_[53196]_  & \new_[53193]_ ;
  assign \new_[53200]_  = A232 & A203;
  assign \new_[53203]_  = A234 & ~A233;
  assign \new_[53204]_  = \new_[53203]_  & \new_[53200]_ ;
  assign \new_[53205]_  = \new_[53204]_  & \new_[53197]_ ;
  assign \new_[53208]_  = A267 & ~A236;
  assign \new_[53211]_  = A269 & ~A268;
  assign \new_[53212]_  = \new_[53211]_  & \new_[53208]_ ;
  assign \new_[53215]_  = A299 & ~A298;
  assign \new_[53218]_  = ~A302 & A300;
  assign \new_[53219]_  = \new_[53218]_  & \new_[53215]_ ;
  assign \new_[53220]_  = \new_[53219]_  & \new_[53212]_ ;
  assign \new_[53223]_  = ~A200 & A199;
  assign \new_[53226]_  = ~A202 & ~A201;
  assign \new_[53227]_  = \new_[53226]_  & \new_[53223]_ ;
  assign \new_[53230]_  = A232 & A203;
  assign \new_[53233]_  = A234 & ~A233;
  assign \new_[53234]_  = \new_[53233]_  & \new_[53230]_ ;
  assign \new_[53235]_  = \new_[53234]_  & \new_[53227]_ ;
  assign \new_[53238]_  = ~A267 & ~A236;
  assign \new_[53241]_  = A298 & A268;
  assign \new_[53242]_  = \new_[53241]_  & \new_[53238]_ ;
  assign \new_[53245]_  = ~A300 & ~A299;
  assign \new_[53248]_  = A302 & ~A301;
  assign \new_[53249]_  = \new_[53248]_  & \new_[53245]_ ;
  assign \new_[53250]_  = \new_[53249]_  & \new_[53242]_ ;
  assign \new_[53253]_  = ~A200 & A199;
  assign \new_[53256]_  = ~A202 & ~A201;
  assign \new_[53257]_  = \new_[53256]_  & \new_[53253]_ ;
  assign \new_[53260]_  = A232 & A203;
  assign \new_[53263]_  = A234 & ~A233;
  assign \new_[53264]_  = \new_[53263]_  & \new_[53260]_ ;
  assign \new_[53265]_  = \new_[53264]_  & \new_[53257]_ ;
  assign \new_[53268]_  = ~A267 & ~A236;
  assign \new_[53271]_  = ~A298 & A268;
  assign \new_[53272]_  = \new_[53271]_  & \new_[53268]_ ;
  assign \new_[53275]_  = ~A300 & A299;
  assign \new_[53278]_  = A302 & ~A301;
  assign \new_[53279]_  = \new_[53278]_  & \new_[53275]_ ;
  assign \new_[53280]_  = \new_[53279]_  & \new_[53272]_ ;
  assign \new_[53283]_  = ~A200 & A199;
  assign \new_[53286]_  = ~A202 & ~A201;
  assign \new_[53287]_  = \new_[53286]_  & \new_[53283]_ ;
  assign \new_[53290]_  = A232 & A203;
  assign \new_[53293]_  = A234 & ~A233;
  assign \new_[53294]_  = \new_[53293]_  & \new_[53290]_ ;
  assign \new_[53295]_  = \new_[53294]_  & \new_[53287]_ ;
  assign \new_[53298]_  = ~A267 & ~A236;
  assign \new_[53301]_  = A298 & ~A269;
  assign \new_[53302]_  = \new_[53301]_  & \new_[53298]_ ;
  assign \new_[53305]_  = ~A300 & ~A299;
  assign \new_[53308]_  = A302 & ~A301;
  assign \new_[53309]_  = \new_[53308]_  & \new_[53305]_ ;
  assign \new_[53310]_  = \new_[53309]_  & \new_[53302]_ ;
  assign \new_[53313]_  = ~A200 & A199;
  assign \new_[53316]_  = ~A202 & ~A201;
  assign \new_[53317]_  = \new_[53316]_  & \new_[53313]_ ;
  assign \new_[53320]_  = A232 & A203;
  assign \new_[53323]_  = A234 & ~A233;
  assign \new_[53324]_  = \new_[53323]_  & \new_[53320]_ ;
  assign \new_[53325]_  = \new_[53324]_  & \new_[53317]_ ;
  assign \new_[53328]_  = ~A267 & ~A236;
  assign \new_[53331]_  = ~A298 & ~A269;
  assign \new_[53332]_  = \new_[53331]_  & \new_[53328]_ ;
  assign \new_[53335]_  = ~A300 & A299;
  assign \new_[53338]_  = A302 & ~A301;
  assign \new_[53339]_  = \new_[53338]_  & \new_[53335]_ ;
  assign \new_[53340]_  = \new_[53339]_  & \new_[53332]_ ;
  assign \new_[53343]_  = ~A200 & A199;
  assign \new_[53346]_  = ~A202 & ~A201;
  assign \new_[53347]_  = \new_[53346]_  & \new_[53343]_ ;
  assign \new_[53350]_  = A232 & A203;
  assign \new_[53353]_  = A234 & ~A233;
  assign \new_[53354]_  = \new_[53353]_  & \new_[53350]_ ;
  assign \new_[53355]_  = \new_[53354]_  & \new_[53347]_ ;
  assign \new_[53358]_  = A265 & ~A236;
  assign \new_[53361]_  = A298 & A266;
  assign \new_[53362]_  = \new_[53361]_  & \new_[53358]_ ;
  assign \new_[53365]_  = ~A300 & ~A299;
  assign \new_[53368]_  = A302 & ~A301;
  assign \new_[53369]_  = \new_[53368]_  & \new_[53365]_ ;
  assign \new_[53370]_  = \new_[53369]_  & \new_[53362]_ ;
  assign \new_[53373]_  = ~A200 & A199;
  assign \new_[53376]_  = ~A202 & ~A201;
  assign \new_[53377]_  = \new_[53376]_  & \new_[53373]_ ;
  assign \new_[53380]_  = A232 & A203;
  assign \new_[53383]_  = A234 & ~A233;
  assign \new_[53384]_  = \new_[53383]_  & \new_[53380]_ ;
  assign \new_[53385]_  = \new_[53384]_  & \new_[53377]_ ;
  assign \new_[53388]_  = A265 & ~A236;
  assign \new_[53391]_  = ~A298 & A266;
  assign \new_[53392]_  = \new_[53391]_  & \new_[53388]_ ;
  assign \new_[53395]_  = ~A300 & A299;
  assign \new_[53398]_  = A302 & ~A301;
  assign \new_[53399]_  = \new_[53398]_  & \new_[53395]_ ;
  assign \new_[53400]_  = \new_[53399]_  & \new_[53392]_ ;
  assign \new_[53403]_  = ~A200 & A199;
  assign \new_[53406]_  = ~A202 & ~A201;
  assign \new_[53407]_  = \new_[53406]_  & \new_[53403]_ ;
  assign \new_[53410]_  = A232 & A203;
  assign \new_[53413]_  = A234 & ~A233;
  assign \new_[53414]_  = \new_[53413]_  & \new_[53410]_ ;
  assign \new_[53415]_  = \new_[53414]_  & \new_[53407]_ ;
  assign \new_[53418]_  = ~A265 & ~A236;
  assign \new_[53421]_  = A298 & ~A266;
  assign \new_[53422]_  = \new_[53421]_  & \new_[53418]_ ;
  assign \new_[53425]_  = ~A300 & ~A299;
  assign \new_[53428]_  = A302 & ~A301;
  assign \new_[53429]_  = \new_[53428]_  & \new_[53425]_ ;
  assign \new_[53430]_  = \new_[53429]_  & \new_[53422]_ ;
  assign \new_[53433]_  = ~A200 & A199;
  assign \new_[53436]_  = ~A202 & ~A201;
  assign \new_[53437]_  = \new_[53436]_  & \new_[53433]_ ;
  assign \new_[53440]_  = A232 & A203;
  assign \new_[53443]_  = A234 & ~A233;
  assign \new_[53444]_  = \new_[53443]_  & \new_[53440]_ ;
  assign \new_[53445]_  = \new_[53444]_  & \new_[53437]_ ;
  assign \new_[53448]_  = ~A265 & ~A236;
  assign \new_[53451]_  = ~A298 & ~A266;
  assign \new_[53452]_  = \new_[53451]_  & \new_[53448]_ ;
  assign \new_[53455]_  = ~A300 & A299;
  assign \new_[53458]_  = A302 & ~A301;
  assign \new_[53459]_  = \new_[53458]_  & \new_[53455]_ ;
  assign \new_[53460]_  = \new_[53459]_  & \new_[53452]_ ;
  assign \new_[53463]_  = ~A200 & A199;
  assign \new_[53466]_  = ~A202 & ~A201;
  assign \new_[53467]_  = \new_[53466]_  & \new_[53463]_ ;
  assign \new_[53470]_  = A232 & A203;
  assign \new_[53473]_  = ~A234 & ~A233;
  assign \new_[53474]_  = \new_[53473]_  & \new_[53470]_ ;
  assign \new_[53475]_  = \new_[53474]_  & \new_[53467]_ ;
  assign \new_[53478]_  = A236 & ~A235;
  assign \new_[53481]_  = A268 & ~A267;
  assign \new_[53482]_  = \new_[53481]_  & \new_[53478]_ ;
  assign \new_[53485]_  = ~A299 & A298;
  assign \new_[53488]_  = A301 & A300;
  assign \new_[53489]_  = \new_[53488]_  & \new_[53485]_ ;
  assign \new_[53490]_  = \new_[53489]_  & \new_[53482]_ ;
  assign \new_[53493]_  = ~A200 & A199;
  assign \new_[53496]_  = ~A202 & ~A201;
  assign \new_[53497]_  = \new_[53496]_  & \new_[53493]_ ;
  assign \new_[53500]_  = A232 & A203;
  assign \new_[53503]_  = ~A234 & ~A233;
  assign \new_[53504]_  = \new_[53503]_  & \new_[53500]_ ;
  assign \new_[53505]_  = \new_[53504]_  & \new_[53497]_ ;
  assign \new_[53508]_  = A236 & ~A235;
  assign \new_[53511]_  = A268 & ~A267;
  assign \new_[53512]_  = \new_[53511]_  & \new_[53508]_ ;
  assign \new_[53515]_  = ~A299 & A298;
  assign \new_[53518]_  = ~A302 & A300;
  assign \new_[53519]_  = \new_[53518]_  & \new_[53515]_ ;
  assign \new_[53520]_  = \new_[53519]_  & \new_[53512]_ ;
  assign \new_[53523]_  = ~A200 & A199;
  assign \new_[53526]_  = ~A202 & ~A201;
  assign \new_[53527]_  = \new_[53526]_  & \new_[53523]_ ;
  assign \new_[53530]_  = A232 & A203;
  assign \new_[53533]_  = ~A234 & ~A233;
  assign \new_[53534]_  = \new_[53533]_  & \new_[53530]_ ;
  assign \new_[53535]_  = \new_[53534]_  & \new_[53527]_ ;
  assign \new_[53538]_  = A236 & ~A235;
  assign \new_[53541]_  = A268 & ~A267;
  assign \new_[53542]_  = \new_[53541]_  & \new_[53538]_ ;
  assign \new_[53545]_  = A299 & ~A298;
  assign \new_[53548]_  = A301 & A300;
  assign \new_[53549]_  = \new_[53548]_  & \new_[53545]_ ;
  assign \new_[53550]_  = \new_[53549]_  & \new_[53542]_ ;
  assign \new_[53553]_  = ~A200 & A199;
  assign \new_[53556]_  = ~A202 & ~A201;
  assign \new_[53557]_  = \new_[53556]_  & \new_[53553]_ ;
  assign \new_[53560]_  = A232 & A203;
  assign \new_[53563]_  = ~A234 & ~A233;
  assign \new_[53564]_  = \new_[53563]_  & \new_[53560]_ ;
  assign \new_[53565]_  = \new_[53564]_  & \new_[53557]_ ;
  assign \new_[53568]_  = A236 & ~A235;
  assign \new_[53571]_  = A268 & ~A267;
  assign \new_[53572]_  = \new_[53571]_  & \new_[53568]_ ;
  assign \new_[53575]_  = A299 & ~A298;
  assign \new_[53578]_  = ~A302 & A300;
  assign \new_[53579]_  = \new_[53578]_  & \new_[53575]_ ;
  assign \new_[53580]_  = \new_[53579]_  & \new_[53572]_ ;
  assign \new_[53583]_  = ~A200 & A199;
  assign \new_[53586]_  = ~A202 & ~A201;
  assign \new_[53587]_  = \new_[53586]_  & \new_[53583]_ ;
  assign \new_[53590]_  = A232 & A203;
  assign \new_[53593]_  = ~A234 & ~A233;
  assign \new_[53594]_  = \new_[53593]_  & \new_[53590]_ ;
  assign \new_[53595]_  = \new_[53594]_  & \new_[53587]_ ;
  assign \new_[53598]_  = A236 & ~A235;
  assign \new_[53601]_  = ~A269 & ~A267;
  assign \new_[53602]_  = \new_[53601]_  & \new_[53598]_ ;
  assign \new_[53605]_  = ~A299 & A298;
  assign \new_[53608]_  = A301 & A300;
  assign \new_[53609]_  = \new_[53608]_  & \new_[53605]_ ;
  assign \new_[53610]_  = \new_[53609]_  & \new_[53602]_ ;
  assign \new_[53613]_  = ~A200 & A199;
  assign \new_[53616]_  = ~A202 & ~A201;
  assign \new_[53617]_  = \new_[53616]_  & \new_[53613]_ ;
  assign \new_[53620]_  = A232 & A203;
  assign \new_[53623]_  = ~A234 & ~A233;
  assign \new_[53624]_  = \new_[53623]_  & \new_[53620]_ ;
  assign \new_[53625]_  = \new_[53624]_  & \new_[53617]_ ;
  assign \new_[53628]_  = A236 & ~A235;
  assign \new_[53631]_  = ~A269 & ~A267;
  assign \new_[53632]_  = \new_[53631]_  & \new_[53628]_ ;
  assign \new_[53635]_  = ~A299 & A298;
  assign \new_[53638]_  = ~A302 & A300;
  assign \new_[53639]_  = \new_[53638]_  & \new_[53635]_ ;
  assign \new_[53640]_  = \new_[53639]_  & \new_[53632]_ ;
  assign \new_[53643]_  = ~A200 & A199;
  assign \new_[53646]_  = ~A202 & ~A201;
  assign \new_[53647]_  = \new_[53646]_  & \new_[53643]_ ;
  assign \new_[53650]_  = A232 & A203;
  assign \new_[53653]_  = ~A234 & ~A233;
  assign \new_[53654]_  = \new_[53653]_  & \new_[53650]_ ;
  assign \new_[53655]_  = \new_[53654]_  & \new_[53647]_ ;
  assign \new_[53658]_  = A236 & ~A235;
  assign \new_[53661]_  = ~A269 & ~A267;
  assign \new_[53662]_  = \new_[53661]_  & \new_[53658]_ ;
  assign \new_[53665]_  = A299 & ~A298;
  assign \new_[53668]_  = A301 & A300;
  assign \new_[53669]_  = \new_[53668]_  & \new_[53665]_ ;
  assign \new_[53670]_  = \new_[53669]_  & \new_[53662]_ ;
  assign \new_[53673]_  = ~A200 & A199;
  assign \new_[53676]_  = ~A202 & ~A201;
  assign \new_[53677]_  = \new_[53676]_  & \new_[53673]_ ;
  assign \new_[53680]_  = A232 & A203;
  assign \new_[53683]_  = ~A234 & ~A233;
  assign \new_[53684]_  = \new_[53683]_  & \new_[53680]_ ;
  assign \new_[53685]_  = \new_[53684]_  & \new_[53677]_ ;
  assign \new_[53688]_  = A236 & ~A235;
  assign \new_[53691]_  = ~A269 & ~A267;
  assign \new_[53692]_  = \new_[53691]_  & \new_[53688]_ ;
  assign \new_[53695]_  = A299 & ~A298;
  assign \new_[53698]_  = ~A302 & A300;
  assign \new_[53699]_  = \new_[53698]_  & \new_[53695]_ ;
  assign \new_[53700]_  = \new_[53699]_  & \new_[53692]_ ;
  assign \new_[53703]_  = ~A200 & A199;
  assign \new_[53706]_  = ~A202 & ~A201;
  assign \new_[53707]_  = \new_[53706]_  & \new_[53703]_ ;
  assign \new_[53710]_  = A232 & A203;
  assign \new_[53713]_  = ~A234 & ~A233;
  assign \new_[53714]_  = \new_[53713]_  & \new_[53710]_ ;
  assign \new_[53715]_  = \new_[53714]_  & \new_[53707]_ ;
  assign \new_[53718]_  = A236 & ~A235;
  assign \new_[53721]_  = A266 & A265;
  assign \new_[53722]_  = \new_[53721]_  & \new_[53718]_ ;
  assign \new_[53725]_  = ~A299 & A298;
  assign \new_[53728]_  = A301 & A300;
  assign \new_[53729]_  = \new_[53728]_  & \new_[53725]_ ;
  assign \new_[53730]_  = \new_[53729]_  & \new_[53722]_ ;
  assign \new_[53733]_  = ~A200 & A199;
  assign \new_[53736]_  = ~A202 & ~A201;
  assign \new_[53737]_  = \new_[53736]_  & \new_[53733]_ ;
  assign \new_[53740]_  = A232 & A203;
  assign \new_[53743]_  = ~A234 & ~A233;
  assign \new_[53744]_  = \new_[53743]_  & \new_[53740]_ ;
  assign \new_[53745]_  = \new_[53744]_  & \new_[53737]_ ;
  assign \new_[53748]_  = A236 & ~A235;
  assign \new_[53751]_  = A266 & A265;
  assign \new_[53752]_  = \new_[53751]_  & \new_[53748]_ ;
  assign \new_[53755]_  = ~A299 & A298;
  assign \new_[53758]_  = ~A302 & A300;
  assign \new_[53759]_  = \new_[53758]_  & \new_[53755]_ ;
  assign \new_[53760]_  = \new_[53759]_  & \new_[53752]_ ;
  assign \new_[53763]_  = ~A200 & A199;
  assign \new_[53766]_  = ~A202 & ~A201;
  assign \new_[53767]_  = \new_[53766]_  & \new_[53763]_ ;
  assign \new_[53770]_  = A232 & A203;
  assign \new_[53773]_  = ~A234 & ~A233;
  assign \new_[53774]_  = \new_[53773]_  & \new_[53770]_ ;
  assign \new_[53775]_  = \new_[53774]_  & \new_[53767]_ ;
  assign \new_[53778]_  = A236 & ~A235;
  assign \new_[53781]_  = A266 & A265;
  assign \new_[53782]_  = \new_[53781]_  & \new_[53778]_ ;
  assign \new_[53785]_  = A299 & ~A298;
  assign \new_[53788]_  = A301 & A300;
  assign \new_[53789]_  = \new_[53788]_  & \new_[53785]_ ;
  assign \new_[53790]_  = \new_[53789]_  & \new_[53782]_ ;
  assign \new_[53793]_  = ~A200 & A199;
  assign \new_[53796]_  = ~A202 & ~A201;
  assign \new_[53797]_  = \new_[53796]_  & \new_[53793]_ ;
  assign \new_[53800]_  = A232 & A203;
  assign \new_[53803]_  = ~A234 & ~A233;
  assign \new_[53804]_  = \new_[53803]_  & \new_[53800]_ ;
  assign \new_[53805]_  = \new_[53804]_  & \new_[53797]_ ;
  assign \new_[53808]_  = A236 & ~A235;
  assign \new_[53811]_  = A266 & A265;
  assign \new_[53812]_  = \new_[53811]_  & \new_[53808]_ ;
  assign \new_[53815]_  = A299 & ~A298;
  assign \new_[53818]_  = ~A302 & A300;
  assign \new_[53819]_  = \new_[53818]_  & \new_[53815]_ ;
  assign \new_[53820]_  = \new_[53819]_  & \new_[53812]_ ;
  assign \new_[53823]_  = ~A200 & A199;
  assign \new_[53826]_  = ~A202 & ~A201;
  assign \new_[53827]_  = \new_[53826]_  & \new_[53823]_ ;
  assign \new_[53830]_  = A232 & A203;
  assign \new_[53833]_  = ~A234 & ~A233;
  assign \new_[53834]_  = \new_[53833]_  & \new_[53830]_ ;
  assign \new_[53835]_  = \new_[53834]_  & \new_[53827]_ ;
  assign \new_[53838]_  = A236 & ~A235;
  assign \new_[53841]_  = ~A266 & ~A265;
  assign \new_[53842]_  = \new_[53841]_  & \new_[53838]_ ;
  assign \new_[53845]_  = ~A299 & A298;
  assign \new_[53848]_  = A301 & A300;
  assign \new_[53849]_  = \new_[53848]_  & \new_[53845]_ ;
  assign \new_[53850]_  = \new_[53849]_  & \new_[53842]_ ;
  assign \new_[53853]_  = ~A200 & A199;
  assign \new_[53856]_  = ~A202 & ~A201;
  assign \new_[53857]_  = \new_[53856]_  & \new_[53853]_ ;
  assign \new_[53860]_  = A232 & A203;
  assign \new_[53863]_  = ~A234 & ~A233;
  assign \new_[53864]_  = \new_[53863]_  & \new_[53860]_ ;
  assign \new_[53865]_  = \new_[53864]_  & \new_[53857]_ ;
  assign \new_[53868]_  = A236 & ~A235;
  assign \new_[53871]_  = ~A266 & ~A265;
  assign \new_[53872]_  = \new_[53871]_  & \new_[53868]_ ;
  assign \new_[53875]_  = ~A299 & A298;
  assign \new_[53878]_  = ~A302 & A300;
  assign \new_[53879]_  = \new_[53878]_  & \new_[53875]_ ;
  assign \new_[53880]_  = \new_[53879]_  & \new_[53872]_ ;
  assign \new_[53883]_  = ~A200 & A199;
  assign \new_[53886]_  = ~A202 & ~A201;
  assign \new_[53887]_  = \new_[53886]_  & \new_[53883]_ ;
  assign \new_[53890]_  = A232 & A203;
  assign \new_[53893]_  = ~A234 & ~A233;
  assign \new_[53894]_  = \new_[53893]_  & \new_[53890]_ ;
  assign \new_[53895]_  = \new_[53894]_  & \new_[53887]_ ;
  assign \new_[53898]_  = A236 & ~A235;
  assign \new_[53901]_  = ~A266 & ~A265;
  assign \new_[53902]_  = \new_[53901]_  & \new_[53898]_ ;
  assign \new_[53905]_  = A299 & ~A298;
  assign \new_[53908]_  = A301 & A300;
  assign \new_[53909]_  = \new_[53908]_  & \new_[53905]_ ;
  assign \new_[53910]_  = \new_[53909]_  & \new_[53902]_ ;
  assign \new_[53913]_  = ~A200 & A199;
  assign \new_[53916]_  = ~A202 & ~A201;
  assign \new_[53917]_  = \new_[53916]_  & \new_[53913]_ ;
  assign \new_[53920]_  = A232 & A203;
  assign \new_[53923]_  = ~A234 & ~A233;
  assign \new_[53924]_  = \new_[53923]_  & \new_[53920]_ ;
  assign \new_[53925]_  = \new_[53924]_  & \new_[53917]_ ;
  assign \new_[53928]_  = A236 & ~A235;
  assign \new_[53931]_  = ~A266 & ~A265;
  assign \new_[53932]_  = \new_[53931]_  & \new_[53928]_ ;
  assign \new_[53935]_  = A299 & ~A298;
  assign \new_[53938]_  = ~A302 & A300;
  assign \new_[53939]_  = \new_[53938]_  & \new_[53935]_ ;
  assign \new_[53940]_  = \new_[53939]_  & \new_[53932]_ ;
  assign \new_[53943]_  = A168 & A170;
  assign \new_[53946]_  = ~A166 & A167;
  assign \new_[53947]_  = \new_[53946]_  & \new_[53943]_ ;
  assign \new_[53950]_  = A233 & ~A232;
  assign \new_[53953]_  = A235 & A234;
  assign \new_[53954]_  = \new_[53953]_  & \new_[53950]_ ;
  assign \new_[53955]_  = \new_[53954]_  & \new_[53947]_ ;
  assign \new_[53958]_  = ~A268 & A267;
  assign \new_[53961]_  = A298 & A269;
  assign \new_[53962]_  = \new_[53961]_  & \new_[53958]_ ;
  assign \new_[53965]_  = ~A300 & ~A299;
  assign \new_[53968]_  = A302 & ~A301;
  assign \new_[53969]_  = \new_[53968]_  & \new_[53965]_ ;
  assign \new_[53970]_  = \new_[53969]_  & \new_[53962]_ ;
  assign \new_[53973]_  = A168 & A170;
  assign \new_[53976]_  = ~A166 & A167;
  assign \new_[53977]_  = \new_[53976]_  & \new_[53973]_ ;
  assign \new_[53980]_  = A233 & ~A232;
  assign \new_[53983]_  = A235 & A234;
  assign \new_[53984]_  = \new_[53983]_  & \new_[53980]_ ;
  assign \new_[53985]_  = \new_[53984]_  & \new_[53977]_ ;
  assign \new_[53988]_  = ~A268 & A267;
  assign \new_[53991]_  = ~A298 & A269;
  assign \new_[53992]_  = \new_[53991]_  & \new_[53988]_ ;
  assign \new_[53995]_  = ~A300 & A299;
  assign \new_[53998]_  = A302 & ~A301;
  assign \new_[53999]_  = \new_[53998]_  & \new_[53995]_ ;
  assign \new_[54000]_  = \new_[53999]_  & \new_[53992]_ ;
  assign \new_[54003]_  = A168 & A170;
  assign \new_[54006]_  = ~A166 & A167;
  assign \new_[54007]_  = \new_[54006]_  & \new_[54003]_ ;
  assign \new_[54010]_  = A233 & ~A232;
  assign \new_[54013]_  = ~A236 & A234;
  assign \new_[54014]_  = \new_[54013]_  & \new_[54010]_ ;
  assign \new_[54015]_  = \new_[54014]_  & \new_[54007]_ ;
  assign \new_[54018]_  = ~A268 & A267;
  assign \new_[54021]_  = A298 & A269;
  assign \new_[54022]_  = \new_[54021]_  & \new_[54018]_ ;
  assign \new_[54025]_  = ~A300 & ~A299;
  assign \new_[54028]_  = A302 & ~A301;
  assign \new_[54029]_  = \new_[54028]_  & \new_[54025]_ ;
  assign \new_[54030]_  = \new_[54029]_  & \new_[54022]_ ;
  assign \new_[54033]_  = A168 & A170;
  assign \new_[54036]_  = ~A166 & A167;
  assign \new_[54037]_  = \new_[54036]_  & \new_[54033]_ ;
  assign \new_[54040]_  = A233 & ~A232;
  assign \new_[54043]_  = ~A236 & A234;
  assign \new_[54044]_  = \new_[54043]_  & \new_[54040]_ ;
  assign \new_[54045]_  = \new_[54044]_  & \new_[54037]_ ;
  assign \new_[54048]_  = ~A268 & A267;
  assign \new_[54051]_  = ~A298 & A269;
  assign \new_[54052]_  = \new_[54051]_  & \new_[54048]_ ;
  assign \new_[54055]_  = ~A300 & A299;
  assign \new_[54058]_  = A302 & ~A301;
  assign \new_[54059]_  = \new_[54058]_  & \new_[54055]_ ;
  assign \new_[54060]_  = \new_[54059]_  & \new_[54052]_ ;
  assign \new_[54063]_  = A168 & A170;
  assign \new_[54066]_  = ~A166 & A167;
  assign \new_[54067]_  = \new_[54066]_  & \new_[54063]_ ;
  assign \new_[54070]_  = A233 & ~A232;
  assign \new_[54073]_  = ~A235 & ~A234;
  assign \new_[54074]_  = \new_[54073]_  & \new_[54070]_ ;
  assign \new_[54075]_  = \new_[54074]_  & \new_[54067]_ ;
  assign \new_[54078]_  = A267 & A236;
  assign \new_[54081]_  = A269 & ~A268;
  assign \new_[54082]_  = \new_[54081]_  & \new_[54078]_ ;
  assign \new_[54085]_  = ~A299 & A298;
  assign \new_[54088]_  = A301 & A300;
  assign \new_[54089]_  = \new_[54088]_  & \new_[54085]_ ;
  assign \new_[54090]_  = \new_[54089]_  & \new_[54082]_ ;
  assign \new_[54093]_  = A168 & A170;
  assign \new_[54096]_  = ~A166 & A167;
  assign \new_[54097]_  = \new_[54096]_  & \new_[54093]_ ;
  assign \new_[54100]_  = A233 & ~A232;
  assign \new_[54103]_  = ~A235 & ~A234;
  assign \new_[54104]_  = \new_[54103]_  & \new_[54100]_ ;
  assign \new_[54105]_  = \new_[54104]_  & \new_[54097]_ ;
  assign \new_[54108]_  = A267 & A236;
  assign \new_[54111]_  = A269 & ~A268;
  assign \new_[54112]_  = \new_[54111]_  & \new_[54108]_ ;
  assign \new_[54115]_  = ~A299 & A298;
  assign \new_[54118]_  = ~A302 & A300;
  assign \new_[54119]_  = \new_[54118]_  & \new_[54115]_ ;
  assign \new_[54120]_  = \new_[54119]_  & \new_[54112]_ ;
  assign \new_[54123]_  = A168 & A170;
  assign \new_[54126]_  = ~A166 & A167;
  assign \new_[54127]_  = \new_[54126]_  & \new_[54123]_ ;
  assign \new_[54130]_  = A233 & ~A232;
  assign \new_[54133]_  = ~A235 & ~A234;
  assign \new_[54134]_  = \new_[54133]_  & \new_[54130]_ ;
  assign \new_[54135]_  = \new_[54134]_  & \new_[54127]_ ;
  assign \new_[54138]_  = A267 & A236;
  assign \new_[54141]_  = A269 & ~A268;
  assign \new_[54142]_  = \new_[54141]_  & \new_[54138]_ ;
  assign \new_[54145]_  = A299 & ~A298;
  assign \new_[54148]_  = A301 & A300;
  assign \new_[54149]_  = \new_[54148]_  & \new_[54145]_ ;
  assign \new_[54150]_  = \new_[54149]_  & \new_[54142]_ ;
  assign \new_[54153]_  = A168 & A170;
  assign \new_[54156]_  = ~A166 & A167;
  assign \new_[54157]_  = \new_[54156]_  & \new_[54153]_ ;
  assign \new_[54160]_  = A233 & ~A232;
  assign \new_[54163]_  = ~A235 & ~A234;
  assign \new_[54164]_  = \new_[54163]_  & \new_[54160]_ ;
  assign \new_[54165]_  = \new_[54164]_  & \new_[54157]_ ;
  assign \new_[54168]_  = A267 & A236;
  assign \new_[54171]_  = A269 & ~A268;
  assign \new_[54172]_  = \new_[54171]_  & \new_[54168]_ ;
  assign \new_[54175]_  = A299 & ~A298;
  assign \new_[54178]_  = ~A302 & A300;
  assign \new_[54179]_  = \new_[54178]_  & \new_[54175]_ ;
  assign \new_[54180]_  = \new_[54179]_  & \new_[54172]_ ;
  assign \new_[54183]_  = A168 & A170;
  assign \new_[54186]_  = ~A166 & A167;
  assign \new_[54187]_  = \new_[54186]_  & \new_[54183]_ ;
  assign \new_[54190]_  = A233 & ~A232;
  assign \new_[54193]_  = ~A235 & ~A234;
  assign \new_[54194]_  = \new_[54193]_  & \new_[54190]_ ;
  assign \new_[54195]_  = \new_[54194]_  & \new_[54187]_ ;
  assign \new_[54198]_  = ~A267 & A236;
  assign \new_[54201]_  = A298 & A268;
  assign \new_[54202]_  = \new_[54201]_  & \new_[54198]_ ;
  assign \new_[54205]_  = ~A300 & ~A299;
  assign \new_[54208]_  = A302 & ~A301;
  assign \new_[54209]_  = \new_[54208]_  & \new_[54205]_ ;
  assign \new_[54210]_  = \new_[54209]_  & \new_[54202]_ ;
  assign \new_[54213]_  = A168 & A170;
  assign \new_[54216]_  = ~A166 & A167;
  assign \new_[54217]_  = \new_[54216]_  & \new_[54213]_ ;
  assign \new_[54220]_  = A233 & ~A232;
  assign \new_[54223]_  = ~A235 & ~A234;
  assign \new_[54224]_  = \new_[54223]_  & \new_[54220]_ ;
  assign \new_[54225]_  = \new_[54224]_  & \new_[54217]_ ;
  assign \new_[54228]_  = ~A267 & A236;
  assign \new_[54231]_  = ~A298 & A268;
  assign \new_[54232]_  = \new_[54231]_  & \new_[54228]_ ;
  assign \new_[54235]_  = ~A300 & A299;
  assign \new_[54238]_  = A302 & ~A301;
  assign \new_[54239]_  = \new_[54238]_  & \new_[54235]_ ;
  assign \new_[54240]_  = \new_[54239]_  & \new_[54232]_ ;
  assign \new_[54243]_  = A168 & A170;
  assign \new_[54246]_  = ~A166 & A167;
  assign \new_[54247]_  = \new_[54246]_  & \new_[54243]_ ;
  assign \new_[54250]_  = A233 & ~A232;
  assign \new_[54253]_  = ~A235 & ~A234;
  assign \new_[54254]_  = \new_[54253]_  & \new_[54250]_ ;
  assign \new_[54255]_  = \new_[54254]_  & \new_[54247]_ ;
  assign \new_[54258]_  = ~A267 & A236;
  assign \new_[54261]_  = A298 & ~A269;
  assign \new_[54262]_  = \new_[54261]_  & \new_[54258]_ ;
  assign \new_[54265]_  = ~A300 & ~A299;
  assign \new_[54268]_  = A302 & ~A301;
  assign \new_[54269]_  = \new_[54268]_  & \new_[54265]_ ;
  assign \new_[54270]_  = \new_[54269]_  & \new_[54262]_ ;
  assign \new_[54273]_  = A168 & A170;
  assign \new_[54276]_  = ~A166 & A167;
  assign \new_[54277]_  = \new_[54276]_  & \new_[54273]_ ;
  assign \new_[54280]_  = A233 & ~A232;
  assign \new_[54283]_  = ~A235 & ~A234;
  assign \new_[54284]_  = \new_[54283]_  & \new_[54280]_ ;
  assign \new_[54285]_  = \new_[54284]_  & \new_[54277]_ ;
  assign \new_[54288]_  = ~A267 & A236;
  assign \new_[54291]_  = ~A298 & ~A269;
  assign \new_[54292]_  = \new_[54291]_  & \new_[54288]_ ;
  assign \new_[54295]_  = ~A300 & A299;
  assign \new_[54298]_  = A302 & ~A301;
  assign \new_[54299]_  = \new_[54298]_  & \new_[54295]_ ;
  assign \new_[54300]_  = \new_[54299]_  & \new_[54292]_ ;
  assign \new_[54303]_  = A168 & A170;
  assign \new_[54306]_  = ~A166 & A167;
  assign \new_[54307]_  = \new_[54306]_  & \new_[54303]_ ;
  assign \new_[54310]_  = A233 & ~A232;
  assign \new_[54313]_  = ~A235 & ~A234;
  assign \new_[54314]_  = \new_[54313]_  & \new_[54310]_ ;
  assign \new_[54315]_  = \new_[54314]_  & \new_[54307]_ ;
  assign \new_[54318]_  = A265 & A236;
  assign \new_[54321]_  = A298 & A266;
  assign \new_[54322]_  = \new_[54321]_  & \new_[54318]_ ;
  assign \new_[54325]_  = ~A300 & ~A299;
  assign \new_[54328]_  = A302 & ~A301;
  assign \new_[54329]_  = \new_[54328]_  & \new_[54325]_ ;
  assign \new_[54330]_  = \new_[54329]_  & \new_[54322]_ ;
  assign \new_[54333]_  = A168 & A170;
  assign \new_[54336]_  = ~A166 & A167;
  assign \new_[54337]_  = \new_[54336]_  & \new_[54333]_ ;
  assign \new_[54340]_  = A233 & ~A232;
  assign \new_[54343]_  = ~A235 & ~A234;
  assign \new_[54344]_  = \new_[54343]_  & \new_[54340]_ ;
  assign \new_[54345]_  = \new_[54344]_  & \new_[54337]_ ;
  assign \new_[54348]_  = A265 & A236;
  assign \new_[54351]_  = ~A298 & A266;
  assign \new_[54352]_  = \new_[54351]_  & \new_[54348]_ ;
  assign \new_[54355]_  = ~A300 & A299;
  assign \new_[54358]_  = A302 & ~A301;
  assign \new_[54359]_  = \new_[54358]_  & \new_[54355]_ ;
  assign \new_[54360]_  = \new_[54359]_  & \new_[54352]_ ;
  assign \new_[54363]_  = A168 & A170;
  assign \new_[54366]_  = ~A166 & A167;
  assign \new_[54367]_  = \new_[54366]_  & \new_[54363]_ ;
  assign \new_[54370]_  = A233 & ~A232;
  assign \new_[54373]_  = ~A235 & ~A234;
  assign \new_[54374]_  = \new_[54373]_  & \new_[54370]_ ;
  assign \new_[54375]_  = \new_[54374]_  & \new_[54367]_ ;
  assign \new_[54378]_  = ~A265 & A236;
  assign \new_[54381]_  = A298 & ~A266;
  assign \new_[54382]_  = \new_[54381]_  & \new_[54378]_ ;
  assign \new_[54385]_  = ~A300 & ~A299;
  assign \new_[54388]_  = A302 & ~A301;
  assign \new_[54389]_  = \new_[54388]_  & \new_[54385]_ ;
  assign \new_[54390]_  = \new_[54389]_  & \new_[54382]_ ;
  assign \new_[54393]_  = A168 & A170;
  assign \new_[54396]_  = ~A166 & A167;
  assign \new_[54397]_  = \new_[54396]_  & \new_[54393]_ ;
  assign \new_[54400]_  = A233 & ~A232;
  assign \new_[54403]_  = ~A235 & ~A234;
  assign \new_[54404]_  = \new_[54403]_  & \new_[54400]_ ;
  assign \new_[54405]_  = \new_[54404]_  & \new_[54397]_ ;
  assign \new_[54408]_  = ~A265 & A236;
  assign \new_[54411]_  = ~A298 & ~A266;
  assign \new_[54412]_  = \new_[54411]_  & \new_[54408]_ ;
  assign \new_[54415]_  = ~A300 & A299;
  assign \new_[54418]_  = A302 & ~A301;
  assign \new_[54419]_  = \new_[54418]_  & \new_[54415]_ ;
  assign \new_[54420]_  = \new_[54419]_  & \new_[54412]_ ;
  assign \new_[54423]_  = A168 & A170;
  assign \new_[54426]_  = ~A166 & A167;
  assign \new_[54427]_  = \new_[54426]_  & \new_[54423]_ ;
  assign \new_[54430]_  = ~A233 & A232;
  assign \new_[54433]_  = A235 & A234;
  assign \new_[54434]_  = \new_[54433]_  & \new_[54430]_ ;
  assign \new_[54435]_  = \new_[54434]_  & \new_[54427]_ ;
  assign \new_[54438]_  = ~A268 & A267;
  assign \new_[54441]_  = A298 & A269;
  assign \new_[54442]_  = \new_[54441]_  & \new_[54438]_ ;
  assign \new_[54445]_  = ~A300 & ~A299;
  assign \new_[54448]_  = A302 & ~A301;
  assign \new_[54449]_  = \new_[54448]_  & \new_[54445]_ ;
  assign \new_[54450]_  = \new_[54449]_  & \new_[54442]_ ;
  assign \new_[54453]_  = A168 & A170;
  assign \new_[54456]_  = ~A166 & A167;
  assign \new_[54457]_  = \new_[54456]_  & \new_[54453]_ ;
  assign \new_[54460]_  = ~A233 & A232;
  assign \new_[54463]_  = A235 & A234;
  assign \new_[54464]_  = \new_[54463]_  & \new_[54460]_ ;
  assign \new_[54465]_  = \new_[54464]_  & \new_[54457]_ ;
  assign \new_[54468]_  = ~A268 & A267;
  assign \new_[54471]_  = ~A298 & A269;
  assign \new_[54472]_  = \new_[54471]_  & \new_[54468]_ ;
  assign \new_[54475]_  = ~A300 & A299;
  assign \new_[54478]_  = A302 & ~A301;
  assign \new_[54479]_  = \new_[54478]_  & \new_[54475]_ ;
  assign \new_[54480]_  = \new_[54479]_  & \new_[54472]_ ;
  assign \new_[54483]_  = A168 & A170;
  assign \new_[54486]_  = ~A166 & A167;
  assign \new_[54487]_  = \new_[54486]_  & \new_[54483]_ ;
  assign \new_[54490]_  = ~A233 & A232;
  assign \new_[54493]_  = ~A236 & A234;
  assign \new_[54494]_  = \new_[54493]_  & \new_[54490]_ ;
  assign \new_[54495]_  = \new_[54494]_  & \new_[54487]_ ;
  assign \new_[54498]_  = ~A268 & A267;
  assign \new_[54501]_  = A298 & A269;
  assign \new_[54502]_  = \new_[54501]_  & \new_[54498]_ ;
  assign \new_[54505]_  = ~A300 & ~A299;
  assign \new_[54508]_  = A302 & ~A301;
  assign \new_[54509]_  = \new_[54508]_  & \new_[54505]_ ;
  assign \new_[54510]_  = \new_[54509]_  & \new_[54502]_ ;
  assign \new_[54513]_  = A168 & A170;
  assign \new_[54516]_  = ~A166 & A167;
  assign \new_[54517]_  = \new_[54516]_  & \new_[54513]_ ;
  assign \new_[54520]_  = ~A233 & A232;
  assign \new_[54523]_  = ~A236 & A234;
  assign \new_[54524]_  = \new_[54523]_  & \new_[54520]_ ;
  assign \new_[54525]_  = \new_[54524]_  & \new_[54517]_ ;
  assign \new_[54528]_  = ~A268 & A267;
  assign \new_[54531]_  = ~A298 & A269;
  assign \new_[54532]_  = \new_[54531]_  & \new_[54528]_ ;
  assign \new_[54535]_  = ~A300 & A299;
  assign \new_[54538]_  = A302 & ~A301;
  assign \new_[54539]_  = \new_[54538]_  & \new_[54535]_ ;
  assign \new_[54540]_  = \new_[54539]_  & \new_[54532]_ ;
  assign \new_[54543]_  = A168 & A170;
  assign \new_[54546]_  = ~A166 & A167;
  assign \new_[54547]_  = \new_[54546]_  & \new_[54543]_ ;
  assign \new_[54550]_  = ~A233 & A232;
  assign \new_[54553]_  = ~A235 & ~A234;
  assign \new_[54554]_  = \new_[54553]_  & \new_[54550]_ ;
  assign \new_[54555]_  = \new_[54554]_  & \new_[54547]_ ;
  assign \new_[54558]_  = A267 & A236;
  assign \new_[54561]_  = A269 & ~A268;
  assign \new_[54562]_  = \new_[54561]_  & \new_[54558]_ ;
  assign \new_[54565]_  = ~A299 & A298;
  assign \new_[54568]_  = A301 & A300;
  assign \new_[54569]_  = \new_[54568]_  & \new_[54565]_ ;
  assign \new_[54570]_  = \new_[54569]_  & \new_[54562]_ ;
  assign \new_[54573]_  = A168 & A170;
  assign \new_[54576]_  = ~A166 & A167;
  assign \new_[54577]_  = \new_[54576]_  & \new_[54573]_ ;
  assign \new_[54580]_  = ~A233 & A232;
  assign \new_[54583]_  = ~A235 & ~A234;
  assign \new_[54584]_  = \new_[54583]_  & \new_[54580]_ ;
  assign \new_[54585]_  = \new_[54584]_  & \new_[54577]_ ;
  assign \new_[54588]_  = A267 & A236;
  assign \new_[54591]_  = A269 & ~A268;
  assign \new_[54592]_  = \new_[54591]_  & \new_[54588]_ ;
  assign \new_[54595]_  = ~A299 & A298;
  assign \new_[54598]_  = ~A302 & A300;
  assign \new_[54599]_  = \new_[54598]_  & \new_[54595]_ ;
  assign \new_[54600]_  = \new_[54599]_  & \new_[54592]_ ;
  assign \new_[54603]_  = A168 & A170;
  assign \new_[54606]_  = ~A166 & A167;
  assign \new_[54607]_  = \new_[54606]_  & \new_[54603]_ ;
  assign \new_[54610]_  = ~A233 & A232;
  assign \new_[54613]_  = ~A235 & ~A234;
  assign \new_[54614]_  = \new_[54613]_  & \new_[54610]_ ;
  assign \new_[54615]_  = \new_[54614]_  & \new_[54607]_ ;
  assign \new_[54618]_  = A267 & A236;
  assign \new_[54621]_  = A269 & ~A268;
  assign \new_[54622]_  = \new_[54621]_  & \new_[54618]_ ;
  assign \new_[54625]_  = A299 & ~A298;
  assign \new_[54628]_  = A301 & A300;
  assign \new_[54629]_  = \new_[54628]_  & \new_[54625]_ ;
  assign \new_[54630]_  = \new_[54629]_  & \new_[54622]_ ;
  assign \new_[54633]_  = A168 & A170;
  assign \new_[54636]_  = ~A166 & A167;
  assign \new_[54637]_  = \new_[54636]_  & \new_[54633]_ ;
  assign \new_[54640]_  = ~A233 & A232;
  assign \new_[54643]_  = ~A235 & ~A234;
  assign \new_[54644]_  = \new_[54643]_  & \new_[54640]_ ;
  assign \new_[54645]_  = \new_[54644]_  & \new_[54637]_ ;
  assign \new_[54648]_  = A267 & A236;
  assign \new_[54651]_  = A269 & ~A268;
  assign \new_[54652]_  = \new_[54651]_  & \new_[54648]_ ;
  assign \new_[54655]_  = A299 & ~A298;
  assign \new_[54658]_  = ~A302 & A300;
  assign \new_[54659]_  = \new_[54658]_  & \new_[54655]_ ;
  assign \new_[54660]_  = \new_[54659]_  & \new_[54652]_ ;
  assign \new_[54663]_  = A168 & A170;
  assign \new_[54666]_  = ~A166 & A167;
  assign \new_[54667]_  = \new_[54666]_  & \new_[54663]_ ;
  assign \new_[54670]_  = ~A233 & A232;
  assign \new_[54673]_  = ~A235 & ~A234;
  assign \new_[54674]_  = \new_[54673]_  & \new_[54670]_ ;
  assign \new_[54675]_  = \new_[54674]_  & \new_[54667]_ ;
  assign \new_[54678]_  = ~A267 & A236;
  assign \new_[54681]_  = A298 & A268;
  assign \new_[54682]_  = \new_[54681]_  & \new_[54678]_ ;
  assign \new_[54685]_  = ~A300 & ~A299;
  assign \new_[54688]_  = A302 & ~A301;
  assign \new_[54689]_  = \new_[54688]_  & \new_[54685]_ ;
  assign \new_[54690]_  = \new_[54689]_  & \new_[54682]_ ;
  assign \new_[54693]_  = A168 & A170;
  assign \new_[54696]_  = ~A166 & A167;
  assign \new_[54697]_  = \new_[54696]_  & \new_[54693]_ ;
  assign \new_[54700]_  = ~A233 & A232;
  assign \new_[54703]_  = ~A235 & ~A234;
  assign \new_[54704]_  = \new_[54703]_  & \new_[54700]_ ;
  assign \new_[54705]_  = \new_[54704]_  & \new_[54697]_ ;
  assign \new_[54708]_  = ~A267 & A236;
  assign \new_[54711]_  = ~A298 & A268;
  assign \new_[54712]_  = \new_[54711]_  & \new_[54708]_ ;
  assign \new_[54715]_  = ~A300 & A299;
  assign \new_[54718]_  = A302 & ~A301;
  assign \new_[54719]_  = \new_[54718]_  & \new_[54715]_ ;
  assign \new_[54720]_  = \new_[54719]_  & \new_[54712]_ ;
  assign \new_[54723]_  = A168 & A170;
  assign \new_[54726]_  = ~A166 & A167;
  assign \new_[54727]_  = \new_[54726]_  & \new_[54723]_ ;
  assign \new_[54730]_  = ~A233 & A232;
  assign \new_[54733]_  = ~A235 & ~A234;
  assign \new_[54734]_  = \new_[54733]_  & \new_[54730]_ ;
  assign \new_[54735]_  = \new_[54734]_  & \new_[54727]_ ;
  assign \new_[54738]_  = ~A267 & A236;
  assign \new_[54741]_  = A298 & ~A269;
  assign \new_[54742]_  = \new_[54741]_  & \new_[54738]_ ;
  assign \new_[54745]_  = ~A300 & ~A299;
  assign \new_[54748]_  = A302 & ~A301;
  assign \new_[54749]_  = \new_[54748]_  & \new_[54745]_ ;
  assign \new_[54750]_  = \new_[54749]_  & \new_[54742]_ ;
  assign \new_[54753]_  = A168 & A170;
  assign \new_[54756]_  = ~A166 & A167;
  assign \new_[54757]_  = \new_[54756]_  & \new_[54753]_ ;
  assign \new_[54760]_  = ~A233 & A232;
  assign \new_[54763]_  = ~A235 & ~A234;
  assign \new_[54764]_  = \new_[54763]_  & \new_[54760]_ ;
  assign \new_[54765]_  = \new_[54764]_  & \new_[54757]_ ;
  assign \new_[54768]_  = ~A267 & A236;
  assign \new_[54771]_  = ~A298 & ~A269;
  assign \new_[54772]_  = \new_[54771]_  & \new_[54768]_ ;
  assign \new_[54775]_  = ~A300 & A299;
  assign \new_[54778]_  = A302 & ~A301;
  assign \new_[54779]_  = \new_[54778]_  & \new_[54775]_ ;
  assign \new_[54780]_  = \new_[54779]_  & \new_[54772]_ ;
  assign \new_[54783]_  = A168 & A170;
  assign \new_[54786]_  = ~A166 & A167;
  assign \new_[54787]_  = \new_[54786]_  & \new_[54783]_ ;
  assign \new_[54790]_  = ~A233 & A232;
  assign \new_[54793]_  = ~A235 & ~A234;
  assign \new_[54794]_  = \new_[54793]_  & \new_[54790]_ ;
  assign \new_[54795]_  = \new_[54794]_  & \new_[54787]_ ;
  assign \new_[54798]_  = A265 & A236;
  assign \new_[54801]_  = A298 & A266;
  assign \new_[54802]_  = \new_[54801]_  & \new_[54798]_ ;
  assign \new_[54805]_  = ~A300 & ~A299;
  assign \new_[54808]_  = A302 & ~A301;
  assign \new_[54809]_  = \new_[54808]_  & \new_[54805]_ ;
  assign \new_[54810]_  = \new_[54809]_  & \new_[54802]_ ;
  assign \new_[54813]_  = A168 & A170;
  assign \new_[54816]_  = ~A166 & A167;
  assign \new_[54817]_  = \new_[54816]_  & \new_[54813]_ ;
  assign \new_[54820]_  = ~A233 & A232;
  assign \new_[54823]_  = ~A235 & ~A234;
  assign \new_[54824]_  = \new_[54823]_  & \new_[54820]_ ;
  assign \new_[54825]_  = \new_[54824]_  & \new_[54817]_ ;
  assign \new_[54828]_  = A265 & A236;
  assign \new_[54831]_  = ~A298 & A266;
  assign \new_[54832]_  = \new_[54831]_  & \new_[54828]_ ;
  assign \new_[54835]_  = ~A300 & A299;
  assign \new_[54838]_  = A302 & ~A301;
  assign \new_[54839]_  = \new_[54838]_  & \new_[54835]_ ;
  assign \new_[54840]_  = \new_[54839]_  & \new_[54832]_ ;
  assign \new_[54843]_  = A168 & A170;
  assign \new_[54846]_  = ~A166 & A167;
  assign \new_[54847]_  = \new_[54846]_  & \new_[54843]_ ;
  assign \new_[54850]_  = ~A233 & A232;
  assign \new_[54853]_  = ~A235 & ~A234;
  assign \new_[54854]_  = \new_[54853]_  & \new_[54850]_ ;
  assign \new_[54855]_  = \new_[54854]_  & \new_[54847]_ ;
  assign \new_[54858]_  = ~A265 & A236;
  assign \new_[54861]_  = A298 & ~A266;
  assign \new_[54862]_  = \new_[54861]_  & \new_[54858]_ ;
  assign \new_[54865]_  = ~A300 & ~A299;
  assign \new_[54868]_  = A302 & ~A301;
  assign \new_[54869]_  = \new_[54868]_  & \new_[54865]_ ;
  assign \new_[54870]_  = \new_[54869]_  & \new_[54862]_ ;
  assign \new_[54873]_  = A168 & A170;
  assign \new_[54876]_  = ~A166 & A167;
  assign \new_[54877]_  = \new_[54876]_  & \new_[54873]_ ;
  assign \new_[54880]_  = ~A233 & A232;
  assign \new_[54883]_  = ~A235 & ~A234;
  assign \new_[54884]_  = \new_[54883]_  & \new_[54880]_ ;
  assign \new_[54885]_  = \new_[54884]_  & \new_[54877]_ ;
  assign \new_[54888]_  = ~A265 & A236;
  assign \new_[54891]_  = ~A298 & ~A266;
  assign \new_[54892]_  = \new_[54891]_  & \new_[54888]_ ;
  assign \new_[54895]_  = ~A300 & A299;
  assign \new_[54898]_  = A302 & ~A301;
  assign \new_[54899]_  = \new_[54898]_  & \new_[54895]_ ;
  assign \new_[54900]_  = \new_[54899]_  & \new_[54892]_ ;
  assign \new_[54903]_  = A168 & A170;
  assign \new_[54906]_  = A166 & ~A167;
  assign \new_[54907]_  = \new_[54906]_  & \new_[54903]_ ;
  assign \new_[54910]_  = A233 & ~A232;
  assign \new_[54913]_  = A235 & A234;
  assign \new_[54914]_  = \new_[54913]_  & \new_[54910]_ ;
  assign \new_[54915]_  = \new_[54914]_  & \new_[54907]_ ;
  assign \new_[54918]_  = ~A268 & A267;
  assign \new_[54921]_  = A298 & A269;
  assign \new_[54922]_  = \new_[54921]_  & \new_[54918]_ ;
  assign \new_[54925]_  = ~A300 & ~A299;
  assign \new_[54928]_  = A302 & ~A301;
  assign \new_[54929]_  = \new_[54928]_  & \new_[54925]_ ;
  assign \new_[54930]_  = \new_[54929]_  & \new_[54922]_ ;
  assign \new_[54933]_  = A168 & A170;
  assign \new_[54936]_  = A166 & ~A167;
  assign \new_[54937]_  = \new_[54936]_  & \new_[54933]_ ;
  assign \new_[54940]_  = A233 & ~A232;
  assign \new_[54943]_  = A235 & A234;
  assign \new_[54944]_  = \new_[54943]_  & \new_[54940]_ ;
  assign \new_[54945]_  = \new_[54944]_  & \new_[54937]_ ;
  assign \new_[54948]_  = ~A268 & A267;
  assign \new_[54951]_  = ~A298 & A269;
  assign \new_[54952]_  = \new_[54951]_  & \new_[54948]_ ;
  assign \new_[54955]_  = ~A300 & A299;
  assign \new_[54958]_  = A302 & ~A301;
  assign \new_[54959]_  = \new_[54958]_  & \new_[54955]_ ;
  assign \new_[54960]_  = \new_[54959]_  & \new_[54952]_ ;
  assign \new_[54963]_  = A168 & A170;
  assign \new_[54966]_  = A166 & ~A167;
  assign \new_[54967]_  = \new_[54966]_  & \new_[54963]_ ;
  assign \new_[54970]_  = A233 & ~A232;
  assign \new_[54973]_  = ~A236 & A234;
  assign \new_[54974]_  = \new_[54973]_  & \new_[54970]_ ;
  assign \new_[54975]_  = \new_[54974]_  & \new_[54967]_ ;
  assign \new_[54978]_  = ~A268 & A267;
  assign \new_[54981]_  = A298 & A269;
  assign \new_[54982]_  = \new_[54981]_  & \new_[54978]_ ;
  assign \new_[54985]_  = ~A300 & ~A299;
  assign \new_[54988]_  = A302 & ~A301;
  assign \new_[54989]_  = \new_[54988]_  & \new_[54985]_ ;
  assign \new_[54990]_  = \new_[54989]_  & \new_[54982]_ ;
  assign \new_[54993]_  = A168 & A170;
  assign \new_[54996]_  = A166 & ~A167;
  assign \new_[54997]_  = \new_[54996]_  & \new_[54993]_ ;
  assign \new_[55000]_  = A233 & ~A232;
  assign \new_[55003]_  = ~A236 & A234;
  assign \new_[55004]_  = \new_[55003]_  & \new_[55000]_ ;
  assign \new_[55005]_  = \new_[55004]_  & \new_[54997]_ ;
  assign \new_[55008]_  = ~A268 & A267;
  assign \new_[55011]_  = ~A298 & A269;
  assign \new_[55012]_  = \new_[55011]_  & \new_[55008]_ ;
  assign \new_[55015]_  = ~A300 & A299;
  assign \new_[55018]_  = A302 & ~A301;
  assign \new_[55019]_  = \new_[55018]_  & \new_[55015]_ ;
  assign \new_[55020]_  = \new_[55019]_  & \new_[55012]_ ;
  assign \new_[55023]_  = A168 & A170;
  assign \new_[55026]_  = A166 & ~A167;
  assign \new_[55027]_  = \new_[55026]_  & \new_[55023]_ ;
  assign \new_[55030]_  = A233 & ~A232;
  assign \new_[55033]_  = ~A235 & ~A234;
  assign \new_[55034]_  = \new_[55033]_  & \new_[55030]_ ;
  assign \new_[55035]_  = \new_[55034]_  & \new_[55027]_ ;
  assign \new_[55038]_  = A267 & A236;
  assign \new_[55041]_  = A269 & ~A268;
  assign \new_[55042]_  = \new_[55041]_  & \new_[55038]_ ;
  assign \new_[55045]_  = ~A299 & A298;
  assign \new_[55048]_  = A301 & A300;
  assign \new_[55049]_  = \new_[55048]_  & \new_[55045]_ ;
  assign \new_[55050]_  = \new_[55049]_  & \new_[55042]_ ;
  assign \new_[55053]_  = A168 & A170;
  assign \new_[55056]_  = A166 & ~A167;
  assign \new_[55057]_  = \new_[55056]_  & \new_[55053]_ ;
  assign \new_[55060]_  = A233 & ~A232;
  assign \new_[55063]_  = ~A235 & ~A234;
  assign \new_[55064]_  = \new_[55063]_  & \new_[55060]_ ;
  assign \new_[55065]_  = \new_[55064]_  & \new_[55057]_ ;
  assign \new_[55068]_  = A267 & A236;
  assign \new_[55071]_  = A269 & ~A268;
  assign \new_[55072]_  = \new_[55071]_  & \new_[55068]_ ;
  assign \new_[55075]_  = ~A299 & A298;
  assign \new_[55078]_  = ~A302 & A300;
  assign \new_[55079]_  = \new_[55078]_  & \new_[55075]_ ;
  assign \new_[55080]_  = \new_[55079]_  & \new_[55072]_ ;
  assign \new_[55083]_  = A168 & A170;
  assign \new_[55086]_  = A166 & ~A167;
  assign \new_[55087]_  = \new_[55086]_  & \new_[55083]_ ;
  assign \new_[55090]_  = A233 & ~A232;
  assign \new_[55093]_  = ~A235 & ~A234;
  assign \new_[55094]_  = \new_[55093]_  & \new_[55090]_ ;
  assign \new_[55095]_  = \new_[55094]_  & \new_[55087]_ ;
  assign \new_[55098]_  = A267 & A236;
  assign \new_[55101]_  = A269 & ~A268;
  assign \new_[55102]_  = \new_[55101]_  & \new_[55098]_ ;
  assign \new_[55105]_  = A299 & ~A298;
  assign \new_[55108]_  = A301 & A300;
  assign \new_[55109]_  = \new_[55108]_  & \new_[55105]_ ;
  assign \new_[55110]_  = \new_[55109]_  & \new_[55102]_ ;
  assign \new_[55113]_  = A168 & A170;
  assign \new_[55116]_  = A166 & ~A167;
  assign \new_[55117]_  = \new_[55116]_  & \new_[55113]_ ;
  assign \new_[55120]_  = A233 & ~A232;
  assign \new_[55123]_  = ~A235 & ~A234;
  assign \new_[55124]_  = \new_[55123]_  & \new_[55120]_ ;
  assign \new_[55125]_  = \new_[55124]_  & \new_[55117]_ ;
  assign \new_[55128]_  = A267 & A236;
  assign \new_[55131]_  = A269 & ~A268;
  assign \new_[55132]_  = \new_[55131]_  & \new_[55128]_ ;
  assign \new_[55135]_  = A299 & ~A298;
  assign \new_[55138]_  = ~A302 & A300;
  assign \new_[55139]_  = \new_[55138]_  & \new_[55135]_ ;
  assign \new_[55140]_  = \new_[55139]_  & \new_[55132]_ ;
  assign \new_[55143]_  = A168 & A170;
  assign \new_[55146]_  = A166 & ~A167;
  assign \new_[55147]_  = \new_[55146]_  & \new_[55143]_ ;
  assign \new_[55150]_  = A233 & ~A232;
  assign \new_[55153]_  = ~A235 & ~A234;
  assign \new_[55154]_  = \new_[55153]_  & \new_[55150]_ ;
  assign \new_[55155]_  = \new_[55154]_  & \new_[55147]_ ;
  assign \new_[55158]_  = ~A267 & A236;
  assign \new_[55161]_  = A298 & A268;
  assign \new_[55162]_  = \new_[55161]_  & \new_[55158]_ ;
  assign \new_[55165]_  = ~A300 & ~A299;
  assign \new_[55168]_  = A302 & ~A301;
  assign \new_[55169]_  = \new_[55168]_  & \new_[55165]_ ;
  assign \new_[55170]_  = \new_[55169]_  & \new_[55162]_ ;
  assign \new_[55173]_  = A168 & A170;
  assign \new_[55176]_  = A166 & ~A167;
  assign \new_[55177]_  = \new_[55176]_  & \new_[55173]_ ;
  assign \new_[55180]_  = A233 & ~A232;
  assign \new_[55183]_  = ~A235 & ~A234;
  assign \new_[55184]_  = \new_[55183]_  & \new_[55180]_ ;
  assign \new_[55185]_  = \new_[55184]_  & \new_[55177]_ ;
  assign \new_[55188]_  = ~A267 & A236;
  assign \new_[55191]_  = ~A298 & A268;
  assign \new_[55192]_  = \new_[55191]_  & \new_[55188]_ ;
  assign \new_[55195]_  = ~A300 & A299;
  assign \new_[55198]_  = A302 & ~A301;
  assign \new_[55199]_  = \new_[55198]_  & \new_[55195]_ ;
  assign \new_[55200]_  = \new_[55199]_  & \new_[55192]_ ;
  assign \new_[55203]_  = A168 & A170;
  assign \new_[55206]_  = A166 & ~A167;
  assign \new_[55207]_  = \new_[55206]_  & \new_[55203]_ ;
  assign \new_[55210]_  = A233 & ~A232;
  assign \new_[55213]_  = ~A235 & ~A234;
  assign \new_[55214]_  = \new_[55213]_  & \new_[55210]_ ;
  assign \new_[55215]_  = \new_[55214]_  & \new_[55207]_ ;
  assign \new_[55218]_  = ~A267 & A236;
  assign \new_[55221]_  = A298 & ~A269;
  assign \new_[55222]_  = \new_[55221]_  & \new_[55218]_ ;
  assign \new_[55225]_  = ~A300 & ~A299;
  assign \new_[55228]_  = A302 & ~A301;
  assign \new_[55229]_  = \new_[55228]_  & \new_[55225]_ ;
  assign \new_[55230]_  = \new_[55229]_  & \new_[55222]_ ;
  assign \new_[55233]_  = A168 & A170;
  assign \new_[55236]_  = A166 & ~A167;
  assign \new_[55237]_  = \new_[55236]_  & \new_[55233]_ ;
  assign \new_[55240]_  = A233 & ~A232;
  assign \new_[55243]_  = ~A235 & ~A234;
  assign \new_[55244]_  = \new_[55243]_  & \new_[55240]_ ;
  assign \new_[55245]_  = \new_[55244]_  & \new_[55237]_ ;
  assign \new_[55248]_  = ~A267 & A236;
  assign \new_[55251]_  = ~A298 & ~A269;
  assign \new_[55252]_  = \new_[55251]_  & \new_[55248]_ ;
  assign \new_[55255]_  = ~A300 & A299;
  assign \new_[55258]_  = A302 & ~A301;
  assign \new_[55259]_  = \new_[55258]_  & \new_[55255]_ ;
  assign \new_[55260]_  = \new_[55259]_  & \new_[55252]_ ;
  assign \new_[55263]_  = A168 & A170;
  assign \new_[55266]_  = A166 & ~A167;
  assign \new_[55267]_  = \new_[55266]_  & \new_[55263]_ ;
  assign \new_[55270]_  = A233 & ~A232;
  assign \new_[55273]_  = ~A235 & ~A234;
  assign \new_[55274]_  = \new_[55273]_  & \new_[55270]_ ;
  assign \new_[55275]_  = \new_[55274]_  & \new_[55267]_ ;
  assign \new_[55278]_  = A265 & A236;
  assign \new_[55281]_  = A298 & A266;
  assign \new_[55282]_  = \new_[55281]_  & \new_[55278]_ ;
  assign \new_[55285]_  = ~A300 & ~A299;
  assign \new_[55288]_  = A302 & ~A301;
  assign \new_[55289]_  = \new_[55288]_  & \new_[55285]_ ;
  assign \new_[55290]_  = \new_[55289]_  & \new_[55282]_ ;
  assign \new_[55293]_  = A168 & A170;
  assign \new_[55296]_  = A166 & ~A167;
  assign \new_[55297]_  = \new_[55296]_  & \new_[55293]_ ;
  assign \new_[55300]_  = A233 & ~A232;
  assign \new_[55303]_  = ~A235 & ~A234;
  assign \new_[55304]_  = \new_[55303]_  & \new_[55300]_ ;
  assign \new_[55305]_  = \new_[55304]_  & \new_[55297]_ ;
  assign \new_[55308]_  = A265 & A236;
  assign \new_[55311]_  = ~A298 & A266;
  assign \new_[55312]_  = \new_[55311]_  & \new_[55308]_ ;
  assign \new_[55315]_  = ~A300 & A299;
  assign \new_[55318]_  = A302 & ~A301;
  assign \new_[55319]_  = \new_[55318]_  & \new_[55315]_ ;
  assign \new_[55320]_  = \new_[55319]_  & \new_[55312]_ ;
  assign \new_[55323]_  = A168 & A170;
  assign \new_[55326]_  = A166 & ~A167;
  assign \new_[55327]_  = \new_[55326]_  & \new_[55323]_ ;
  assign \new_[55330]_  = A233 & ~A232;
  assign \new_[55333]_  = ~A235 & ~A234;
  assign \new_[55334]_  = \new_[55333]_  & \new_[55330]_ ;
  assign \new_[55335]_  = \new_[55334]_  & \new_[55327]_ ;
  assign \new_[55338]_  = ~A265 & A236;
  assign \new_[55341]_  = A298 & ~A266;
  assign \new_[55342]_  = \new_[55341]_  & \new_[55338]_ ;
  assign \new_[55345]_  = ~A300 & ~A299;
  assign \new_[55348]_  = A302 & ~A301;
  assign \new_[55349]_  = \new_[55348]_  & \new_[55345]_ ;
  assign \new_[55350]_  = \new_[55349]_  & \new_[55342]_ ;
  assign \new_[55353]_  = A168 & A170;
  assign \new_[55356]_  = A166 & ~A167;
  assign \new_[55357]_  = \new_[55356]_  & \new_[55353]_ ;
  assign \new_[55360]_  = A233 & ~A232;
  assign \new_[55363]_  = ~A235 & ~A234;
  assign \new_[55364]_  = \new_[55363]_  & \new_[55360]_ ;
  assign \new_[55365]_  = \new_[55364]_  & \new_[55357]_ ;
  assign \new_[55368]_  = ~A265 & A236;
  assign \new_[55371]_  = ~A298 & ~A266;
  assign \new_[55372]_  = \new_[55371]_  & \new_[55368]_ ;
  assign \new_[55375]_  = ~A300 & A299;
  assign \new_[55378]_  = A302 & ~A301;
  assign \new_[55379]_  = \new_[55378]_  & \new_[55375]_ ;
  assign \new_[55380]_  = \new_[55379]_  & \new_[55372]_ ;
  assign \new_[55383]_  = A168 & A170;
  assign \new_[55386]_  = A166 & ~A167;
  assign \new_[55387]_  = \new_[55386]_  & \new_[55383]_ ;
  assign \new_[55390]_  = ~A233 & A232;
  assign \new_[55393]_  = A235 & A234;
  assign \new_[55394]_  = \new_[55393]_  & \new_[55390]_ ;
  assign \new_[55395]_  = \new_[55394]_  & \new_[55387]_ ;
  assign \new_[55398]_  = ~A268 & A267;
  assign \new_[55401]_  = A298 & A269;
  assign \new_[55402]_  = \new_[55401]_  & \new_[55398]_ ;
  assign \new_[55405]_  = ~A300 & ~A299;
  assign \new_[55408]_  = A302 & ~A301;
  assign \new_[55409]_  = \new_[55408]_  & \new_[55405]_ ;
  assign \new_[55410]_  = \new_[55409]_  & \new_[55402]_ ;
  assign \new_[55413]_  = A168 & A170;
  assign \new_[55416]_  = A166 & ~A167;
  assign \new_[55417]_  = \new_[55416]_  & \new_[55413]_ ;
  assign \new_[55420]_  = ~A233 & A232;
  assign \new_[55423]_  = A235 & A234;
  assign \new_[55424]_  = \new_[55423]_  & \new_[55420]_ ;
  assign \new_[55425]_  = \new_[55424]_  & \new_[55417]_ ;
  assign \new_[55428]_  = ~A268 & A267;
  assign \new_[55431]_  = ~A298 & A269;
  assign \new_[55432]_  = \new_[55431]_  & \new_[55428]_ ;
  assign \new_[55435]_  = ~A300 & A299;
  assign \new_[55438]_  = A302 & ~A301;
  assign \new_[55439]_  = \new_[55438]_  & \new_[55435]_ ;
  assign \new_[55440]_  = \new_[55439]_  & \new_[55432]_ ;
  assign \new_[55443]_  = A168 & A170;
  assign \new_[55446]_  = A166 & ~A167;
  assign \new_[55447]_  = \new_[55446]_  & \new_[55443]_ ;
  assign \new_[55450]_  = ~A233 & A232;
  assign \new_[55453]_  = ~A236 & A234;
  assign \new_[55454]_  = \new_[55453]_  & \new_[55450]_ ;
  assign \new_[55455]_  = \new_[55454]_  & \new_[55447]_ ;
  assign \new_[55458]_  = ~A268 & A267;
  assign \new_[55461]_  = A298 & A269;
  assign \new_[55462]_  = \new_[55461]_  & \new_[55458]_ ;
  assign \new_[55465]_  = ~A300 & ~A299;
  assign \new_[55468]_  = A302 & ~A301;
  assign \new_[55469]_  = \new_[55468]_  & \new_[55465]_ ;
  assign \new_[55470]_  = \new_[55469]_  & \new_[55462]_ ;
  assign \new_[55473]_  = A168 & A170;
  assign \new_[55476]_  = A166 & ~A167;
  assign \new_[55477]_  = \new_[55476]_  & \new_[55473]_ ;
  assign \new_[55480]_  = ~A233 & A232;
  assign \new_[55483]_  = ~A236 & A234;
  assign \new_[55484]_  = \new_[55483]_  & \new_[55480]_ ;
  assign \new_[55485]_  = \new_[55484]_  & \new_[55477]_ ;
  assign \new_[55488]_  = ~A268 & A267;
  assign \new_[55491]_  = ~A298 & A269;
  assign \new_[55492]_  = \new_[55491]_  & \new_[55488]_ ;
  assign \new_[55495]_  = ~A300 & A299;
  assign \new_[55498]_  = A302 & ~A301;
  assign \new_[55499]_  = \new_[55498]_  & \new_[55495]_ ;
  assign \new_[55500]_  = \new_[55499]_  & \new_[55492]_ ;
  assign \new_[55503]_  = A168 & A170;
  assign \new_[55506]_  = A166 & ~A167;
  assign \new_[55507]_  = \new_[55506]_  & \new_[55503]_ ;
  assign \new_[55510]_  = ~A233 & A232;
  assign \new_[55513]_  = ~A235 & ~A234;
  assign \new_[55514]_  = \new_[55513]_  & \new_[55510]_ ;
  assign \new_[55515]_  = \new_[55514]_  & \new_[55507]_ ;
  assign \new_[55518]_  = A267 & A236;
  assign \new_[55521]_  = A269 & ~A268;
  assign \new_[55522]_  = \new_[55521]_  & \new_[55518]_ ;
  assign \new_[55525]_  = ~A299 & A298;
  assign \new_[55528]_  = A301 & A300;
  assign \new_[55529]_  = \new_[55528]_  & \new_[55525]_ ;
  assign \new_[55530]_  = \new_[55529]_  & \new_[55522]_ ;
  assign \new_[55533]_  = A168 & A170;
  assign \new_[55536]_  = A166 & ~A167;
  assign \new_[55537]_  = \new_[55536]_  & \new_[55533]_ ;
  assign \new_[55540]_  = ~A233 & A232;
  assign \new_[55543]_  = ~A235 & ~A234;
  assign \new_[55544]_  = \new_[55543]_  & \new_[55540]_ ;
  assign \new_[55545]_  = \new_[55544]_  & \new_[55537]_ ;
  assign \new_[55548]_  = A267 & A236;
  assign \new_[55551]_  = A269 & ~A268;
  assign \new_[55552]_  = \new_[55551]_  & \new_[55548]_ ;
  assign \new_[55555]_  = ~A299 & A298;
  assign \new_[55558]_  = ~A302 & A300;
  assign \new_[55559]_  = \new_[55558]_  & \new_[55555]_ ;
  assign \new_[55560]_  = \new_[55559]_  & \new_[55552]_ ;
  assign \new_[55563]_  = A168 & A170;
  assign \new_[55566]_  = A166 & ~A167;
  assign \new_[55567]_  = \new_[55566]_  & \new_[55563]_ ;
  assign \new_[55570]_  = ~A233 & A232;
  assign \new_[55573]_  = ~A235 & ~A234;
  assign \new_[55574]_  = \new_[55573]_  & \new_[55570]_ ;
  assign \new_[55575]_  = \new_[55574]_  & \new_[55567]_ ;
  assign \new_[55578]_  = A267 & A236;
  assign \new_[55581]_  = A269 & ~A268;
  assign \new_[55582]_  = \new_[55581]_  & \new_[55578]_ ;
  assign \new_[55585]_  = A299 & ~A298;
  assign \new_[55588]_  = A301 & A300;
  assign \new_[55589]_  = \new_[55588]_  & \new_[55585]_ ;
  assign \new_[55590]_  = \new_[55589]_  & \new_[55582]_ ;
  assign \new_[55593]_  = A168 & A170;
  assign \new_[55596]_  = A166 & ~A167;
  assign \new_[55597]_  = \new_[55596]_  & \new_[55593]_ ;
  assign \new_[55600]_  = ~A233 & A232;
  assign \new_[55603]_  = ~A235 & ~A234;
  assign \new_[55604]_  = \new_[55603]_  & \new_[55600]_ ;
  assign \new_[55605]_  = \new_[55604]_  & \new_[55597]_ ;
  assign \new_[55608]_  = A267 & A236;
  assign \new_[55611]_  = A269 & ~A268;
  assign \new_[55612]_  = \new_[55611]_  & \new_[55608]_ ;
  assign \new_[55615]_  = A299 & ~A298;
  assign \new_[55618]_  = ~A302 & A300;
  assign \new_[55619]_  = \new_[55618]_  & \new_[55615]_ ;
  assign \new_[55620]_  = \new_[55619]_  & \new_[55612]_ ;
  assign \new_[55623]_  = A168 & A170;
  assign \new_[55626]_  = A166 & ~A167;
  assign \new_[55627]_  = \new_[55626]_  & \new_[55623]_ ;
  assign \new_[55630]_  = ~A233 & A232;
  assign \new_[55633]_  = ~A235 & ~A234;
  assign \new_[55634]_  = \new_[55633]_  & \new_[55630]_ ;
  assign \new_[55635]_  = \new_[55634]_  & \new_[55627]_ ;
  assign \new_[55638]_  = ~A267 & A236;
  assign \new_[55641]_  = A298 & A268;
  assign \new_[55642]_  = \new_[55641]_  & \new_[55638]_ ;
  assign \new_[55645]_  = ~A300 & ~A299;
  assign \new_[55648]_  = A302 & ~A301;
  assign \new_[55649]_  = \new_[55648]_  & \new_[55645]_ ;
  assign \new_[55650]_  = \new_[55649]_  & \new_[55642]_ ;
  assign \new_[55653]_  = A168 & A170;
  assign \new_[55656]_  = A166 & ~A167;
  assign \new_[55657]_  = \new_[55656]_  & \new_[55653]_ ;
  assign \new_[55660]_  = ~A233 & A232;
  assign \new_[55663]_  = ~A235 & ~A234;
  assign \new_[55664]_  = \new_[55663]_  & \new_[55660]_ ;
  assign \new_[55665]_  = \new_[55664]_  & \new_[55657]_ ;
  assign \new_[55668]_  = ~A267 & A236;
  assign \new_[55671]_  = ~A298 & A268;
  assign \new_[55672]_  = \new_[55671]_  & \new_[55668]_ ;
  assign \new_[55675]_  = ~A300 & A299;
  assign \new_[55678]_  = A302 & ~A301;
  assign \new_[55679]_  = \new_[55678]_  & \new_[55675]_ ;
  assign \new_[55680]_  = \new_[55679]_  & \new_[55672]_ ;
  assign \new_[55683]_  = A168 & A170;
  assign \new_[55686]_  = A166 & ~A167;
  assign \new_[55687]_  = \new_[55686]_  & \new_[55683]_ ;
  assign \new_[55690]_  = ~A233 & A232;
  assign \new_[55693]_  = ~A235 & ~A234;
  assign \new_[55694]_  = \new_[55693]_  & \new_[55690]_ ;
  assign \new_[55695]_  = \new_[55694]_  & \new_[55687]_ ;
  assign \new_[55698]_  = ~A267 & A236;
  assign \new_[55701]_  = A298 & ~A269;
  assign \new_[55702]_  = \new_[55701]_  & \new_[55698]_ ;
  assign \new_[55705]_  = ~A300 & ~A299;
  assign \new_[55708]_  = A302 & ~A301;
  assign \new_[55709]_  = \new_[55708]_  & \new_[55705]_ ;
  assign \new_[55710]_  = \new_[55709]_  & \new_[55702]_ ;
  assign \new_[55713]_  = A168 & A170;
  assign \new_[55716]_  = A166 & ~A167;
  assign \new_[55717]_  = \new_[55716]_  & \new_[55713]_ ;
  assign \new_[55720]_  = ~A233 & A232;
  assign \new_[55723]_  = ~A235 & ~A234;
  assign \new_[55724]_  = \new_[55723]_  & \new_[55720]_ ;
  assign \new_[55725]_  = \new_[55724]_  & \new_[55717]_ ;
  assign \new_[55728]_  = ~A267 & A236;
  assign \new_[55731]_  = ~A298 & ~A269;
  assign \new_[55732]_  = \new_[55731]_  & \new_[55728]_ ;
  assign \new_[55735]_  = ~A300 & A299;
  assign \new_[55738]_  = A302 & ~A301;
  assign \new_[55739]_  = \new_[55738]_  & \new_[55735]_ ;
  assign \new_[55740]_  = \new_[55739]_  & \new_[55732]_ ;
  assign \new_[55743]_  = A168 & A170;
  assign \new_[55746]_  = A166 & ~A167;
  assign \new_[55747]_  = \new_[55746]_  & \new_[55743]_ ;
  assign \new_[55750]_  = ~A233 & A232;
  assign \new_[55753]_  = ~A235 & ~A234;
  assign \new_[55754]_  = \new_[55753]_  & \new_[55750]_ ;
  assign \new_[55755]_  = \new_[55754]_  & \new_[55747]_ ;
  assign \new_[55758]_  = A265 & A236;
  assign \new_[55761]_  = A298 & A266;
  assign \new_[55762]_  = \new_[55761]_  & \new_[55758]_ ;
  assign \new_[55765]_  = ~A300 & ~A299;
  assign \new_[55768]_  = A302 & ~A301;
  assign \new_[55769]_  = \new_[55768]_  & \new_[55765]_ ;
  assign \new_[55770]_  = \new_[55769]_  & \new_[55762]_ ;
  assign \new_[55773]_  = A168 & A170;
  assign \new_[55776]_  = A166 & ~A167;
  assign \new_[55777]_  = \new_[55776]_  & \new_[55773]_ ;
  assign \new_[55780]_  = ~A233 & A232;
  assign \new_[55783]_  = ~A235 & ~A234;
  assign \new_[55784]_  = \new_[55783]_  & \new_[55780]_ ;
  assign \new_[55785]_  = \new_[55784]_  & \new_[55777]_ ;
  assign \new_[55788]_  = A265 & A236;
  assign \new_[55791]_  = ~A298 & A266;
  assign \new_[55792]_  = \new_[55791]_  & \new_[55788]_ ;
  assign \new_[55795]_  = ~A300 & A299;
  assign \new_[55798]_  = A302 & ~A301;
  assign \new_[55799]_  = \new_[55798]_  & \new_[55795]_ ;
  assign \new_[55800]_  = \new_[55799]_  & \new_[55792]_ ;
  assign \new_[55803]_  = A168 & A170;
  assign \new_[55806]_  = A166 & ~A167;
  assign \new_[55807]_  = \new_[55806]_  & \new_[55803]_ ;
  assign \new_[55810]_  = ~A233 & A232;
  assign \new_[55813]_  = ~A235 & ~A234;
  assign \new_[55814]_  = \new_[55813]_  & \new_[55810]_ ;
  assign \new_[55815]_  = \new_[55814]_  & \new_[55807]_ ;
  assign \new_[55818]_  = ~A265 & A236;
  assign \new_[55821]_  = A298 & ~A266;
  assign \new_[55822]_  = \new_[55821]_  & \new_[55818]_ ;
  assign \new_[55825]_  = ~A300 & ~A299;
  assign \new_[55828]_  = A302 & ~A301;
  assign \new_[55829]_  = \new_[55828]_  & \new_[55825]_ ;
  assign \new_[55830]_  = \new_[55829]_  & \new_[55822]_ ;
  assign \new_[55833]_  = A168 & A170;
  assign \new_[55836]_  = A166 & ~A167;
  assign \new_[55837]_  = \new_[55836]_  & \new_[55833]_ ;
  assign \new_[55840]_  = ~A233 & A232;
  assign \new_[55843]_  = ~A235 & ~A234;
  assign \new_[55844]_  = \new_[55843]_  & \new_[55840]_ ;
  assign \new_[55845]_  = \new_[55844]_  & \new_[55837]_ ;
  assign \new_[55848]_  = ~A265 & A236;
  assign \new_[55851]_  = ~A298 & ~A266;
  assign \new_[55852]_  = \new_[55851]_  & \new_[55848]_ ;
  assign \new_[55855]_  = ~A300 & A299;
  assign \new_[55858]_  = A302 & ~A301;
  assign \new_[55859]_  = \new_[55858]_  & \new_[55855]_ ;
  assign \new_[55860]_  = \new_[55859]_  & \new_[55852]_ ;
  assign \new_[55863]_  = A168 & A169;
  assign \new_[55866]_  = ~A166 & A167;
  assign \new_[55867]_  = \new_[55866]_  & \new_[55863]_ ;
  assign \new_[55870]_  = A233 & ~A232;
  assign \new_[55873]_  = A235 & A234;
  assign \new_[55874]_  = \new_[55873]_  & \new_[55870]_ ;
  assign \new_[55875]_  = \new_[55874]_  & \new_[55867]_ ;
  assign \new_[55878]_  = ~A268 & A267;
  assign \new_[55881]_  = A298 & A269;
  assign \new_[55882]_  = \new_[55881]_  & \new_[55878]_ ;
  assign \new_[55885]_  = ~A300 & ~A299;
  assign \new_[55888]_  = A302 & ~A301;
  assign \new_[55889]_  = \new_[55888]_  & \new_[55885]_ ;
  assign \new_[55890]_  = \new_[55889]_  & \new_[55882]_ ;
  assign \new_[55893]_  = A168 & A169;
  assign \new_[55896]_  = ~A166 & A167;
  assign \new_[55897]_  = \new_[55896]_  & \new_[55893]_ ;
  assign \new_[55900]_  = A233 & ~A232;
  assign \new_[55903]_  = A235 & A234;
  assign \new_[55904]_  = \new_[55903]_  & \new_[55900]_ ;
  assign \new_[55905]_  = \new_[55904]_  & \new_[55897]_ ;
  assign \new_[55908]_  = ~A268 & A267;
  assign \new_[55911]_  = ~A298 & A269;
  assign \new_[55912]_  = \new_[55911]_  & \new_[55908]_ ;
  assign \new_[55915]_  = ~A300 & A299;
  assign \new_[55918]_  = A302 & ~A301;
  assign \new_[55919]_  = \new_[55918]_  & \new_[55915]_ ;
  assign \new_[55920]_  = \new_[55919]_  & \new_[55912]_ ;
  assign \new_[55923]_  = A168 & A169;
  assign \new_[55926]_  = ~A166 & A167;
  assign \new_[55927]_  = \new_[55926]_  & \new_[55923]_ ;
  assign \new_[55930]_  = A233 & ~A232;
  assign \new_[55933]_  = ~A236 & A234;
  assign \new_[55934]_  = \new_[55933]_  & \new_[55930]_ ;
  assign \new_[55935]_  = \new_[55934]_  & \new_[55927]_ ;
  assign \new_[55938]_  = ~A268 & A267;
  assign \new_[55941]_  = A298 & A269;
  assign \new_[55942]_  = \new_[55941]_  & \new_[55938]_ ;
  assign \new_[55945]_  = ~A300 & ~A299;
  assign \new_[55948]_  = A302 & ~A301;
  assign \new_[55949]_  = \new_[55948]_  & \new_[55945]_ ;
  assign \new_[55950]_  = \new_[55949]_  & \new_[55942]_ ;
  assign \new_[55953]_  = A168 & A169;
  assign \new_[55956]_  = ~A166 & A167;
  assign \new_[55957]_  = \new_[55956]_  & \new_[55953]_ ;
  assign \new_[55960]_  = A233 & ~A232;
  assign \new_[55963]_  = ~A236 & A234;
  assign \new_[55964]_  = \new_[55963]_  & \new_[55960]_ ;
  assign \new_[55965]_  = \new_[55964]_  & \new_[55957]_ ;
  assign \new_[55968]_  = ~A268 & A267;
  assign \new_[55971]_  = ~A298 & A269;
  assign \new_[55972]_  = \new_[55971]_  & \new_[55968]_ ;
  assign \new_[55975]_  = ~A300 & A299;
  assign \new_[55978]_  = A302 & ~A301;
  assign \new_[55979]_  = \new_[55978]_  & \new_[55975]_ ;
  assign \new_[55980]_  = \new_[55979]_  & \new_[55972]_ ;
  assign \new_[55983]_  = A168 & A169;
  assign \new_[55986]_  = ~A166 & A167;
  assign \new_[55987]_  = \new_[55986]_  & \new_[55983]_ ;
  assign \new_[55990]_  = A233 & ~A232;
  assign \new_[55993]_  = ~A235 & ~A234;
  assign \new_[55994]_  = \new_[55993]_  & \new_[55990]_ ;
  assign \new_[55995]_  = \new_[55994]_  & \new_[55987]_ ;
  assign \new_[55998]_  = A267 & A236;
  assign \new_[56001]_  = A269 & ~A268;
  assign \new_[56002]_  = \new_[56001]_  & \new_[55998]_ ;
  assign \new_[56005]_  = ~A299 & A298;
  assign \new_[56008]_  = A301 & A300;
  assign \new_[56009]_  = \new_[56008]_  & \new_[56005]_ ;
  assign \new_[56010]_  = \new_[56009]_  & \new_[56002]_ ;
  assign \new_[56013]_  = A168 & A169;
  assign \new_[56016]_  = ~A166 & A167;
  assign \new_[56017]_  = \new_[56016]_  & \new_[56013]_ ;
  assign \new_[56020]_  = A233 & ~A232;
  assign \new_[56023]_  = ~A235 & ~A234;
  assign \new_[56024]_  = \new_[56023]_  & \new_[56020]_ ;
  assign \new_[56025]_  = \new_[56024]_  & \new_[56017]_ ;
  assign \new_[56028]_  = A267 & A236;
  assign \new_[56031]_  = A269 & ~A268;
  assign \new_[56032]_  = \new_[56031]_  & \new_[56028]_ ;
  assign \new_[56035]_  = ~A299 & A298;
  assign \new_[56038]_  = ~A302 & A300;
  assign \new_[56039]_  = \new_[56038]_  & \new_[56035]_ ;
  assign \new_[56040]_  = \new_[56039]_  & \new_[56032]_ ;
  assign \new_[56043]_  = A168 & A169;
  assign \new_[56046]_  = ~A166 & A167;
  assign \new_[56047]_  = \new_[56046]_  & \new_[56043]_ ;
  assign \new_[56050]_  = A233 & ~A232;
  assign \new_[56053]_  = ~A235 & ~A234;
  assign \new_[56054]_  = \new_[56053]_  & \new_[56050]_ ;
  assign \new_[56055]_  = \new_[56054]_  & \new_[56047]_ ;
  assign \new_[56058]_  = A267 & A236;
  assign \new_[56061]_  = A269 & ~A268;
  assign \new_[56062]_  = \new_[56061]_  & \new_[56058]_ ;
  assign \new_[56065]_  = A299 & ~A298;
  assign \new_[56068]_  = A301 & A300;
  assign \new_[56069]_  = \new_[56068]_  & \new_[56065]_ ;
  assign \new_[56070]_  = \new_[56069]_  & \new_[56062]_ ;
  assign \new_[56073]_  = A168 & A169;
  assign \new_[56076]_  = ~A166 & A167;
  assign \new_[56077]_  = \new_[56076]_  & \new_[56073]_ ;
  assign \new_[56080]_  = A233 & ~A232;
  assign \new_[56083]_  = ~A235 & ~A234;
  assign \new_[56084]_  = \new_[56083]_  & \new_[56080]_ ;
  assign \new_[56085]_  = \new_[56084]_  & \new_[56077]_ ;
  assign \new_[56088]_  = A267 & A236;
  assign \new_[56091]_  = A269 & ~A268;
  assign \new_[56092]_  = \new_[56091]_  & \new_[56088]_ ;
  assign \new_[56095]_  = A299 & ~A298;
  assign \new_[56098]_  = ~A302 & A300;
  assign \new_[56099]_  = \new_[56098]_  & \new_[56095]_ ;
  assign \new_[56100]_  = \new_[56099]_  & \new_[56092]_ ;
  assign \new_[56103]_  = A168 & A169;
  assign \new_[56106]_  = ~A166 & A167;
  assign \new_[56107]_  = \new_[56106]_  & \new_[56103]_ ;
  assign \new_[56110]_  = A233 & ~A232;
  assign \new_[56113]_  = ~A235 & ~A234;
  assign \new_[56114]_  = \new_[56113]_  & \new_[56110]_ ;
  assign \new_[56115]_  = \new_[56114]_  & \new_[56107]_ ;
  assign \new_[56118]_  = ~A267 & A236;
  assign \new_[56121]_  = A298 & A268;
  assign \new_[56122]_  = \new_[56121]_  & \new_[56118]_ ;
  assign \new_[56125]_  = ~A300 & ~A299;
  assign \new_[56128]_  = A302 & ~A301;
  assign \new_[56129]_  = \new_[56128]_  & \new_[56125]_ ;
  assign \new_[56130]_  = \new_[56129]_  & \new_[56122]_ ;
  assign \new_[56133]_  = A168 & A169;
  assign \new_[56136]_  = ~A166 & A167;
  assign \new_[56137]_  = \new_[56136]_  & \new_[56133]_ ;
  assign \new_[56140]_  = A233 & ~A232;
  assign \new_[56143]_  = ~A235 & ~A234;
  assign \new_[56144]_  = \new_[56143]_  & \new_[56140]_ ;
  assign \new_[56145]_  = \new_[56144]_  & \new_[56137]_ ;
  assign \new_[56148]_  = ~A267 & A236;
  assign \new_[56151]_  = ~A298 & A268;
  assign \new_[56152]_  = \new_[56151]_  & \new_[56148]_ ;
  assign \new_[56155]_  = ~A300 & A299;
  assign \new_[56158]_  = A302 & ~A301;
  assign \new_[56159]_  = \new_[56158]_  & \new_[56155]_ ;
  assign \new_[56160]_  = \new_[56159]_  & \new_[56152]_ ;
  assign \new_[56163]_  = A168 & A169;
  assign \new_[56166]_  = ~A166 & A167;
  assign \new_[56167]_  = \new_[56166]_  & \new_[56163]_ ;
  assign \new_[56170]_  = A233 & ~A232;
  assign \new_[56173]_  = ~A235 & ~A234;
  assign \new_[56174]_  = \new_[56173]_  & \new_[56170]_ ;
  assign \new_[56175]_  = \new_[56174]_  & \new_[56167]_ ;
  assign \new_[56178]_  = ~A267 & A236;
  assign \new_[56181]_  = A298 & ~A269;
  assign \new_[56182]_  = \new_[56181]_  & \new_[56178]_ ;
  assign \new_[56185]_  = ~A300 & ~A299;
  assign \new_[56188]_  = A302 & ~A301;
  assign \new_[56189]_  = \new_[56188]_  & \new_[56185]_ ;
  assign \new_[56190]_  = \new_[56189]_  & \new_[56182]_ ;
  assign \new_[56193]_  = A168 & A169;
  assign \new_[56196]_  = ~A166 & A167;
  assign \new_[56197]_  = \new_[56196]_  & \new_[56193]_ ;
  assign \new_[56200]_  = A233 & ~A232;
  assign \new_[56203]_  = ~A235 & ~A234;
  assign \new_[56204]_  = \new_[56203]_  & \new_[56200]_ ;
  assign \new_[56205]_  = \new_[56204]_  & \new_[56197]_ ;
  assign \new_[56208]_  = ~A267 & A236;
  assign \new_[56211]_  = ~A298 & ~A269;
  assign \new_[56212]_  = \new_[56211]_  & \new_[56208]_ ;
  assign \new_[56215]_  = ~A300 & A299;
  assign \new_[56218]_  = A302 & ~A301;
  assign \new_[56219]_  = \new_[56218]_  & \new_[56215]_ ;
  assign \new_[56220]_  = \new_[56219]_  & \new_[56212]_ ;
  assign \new_[56223]_  = A168 & A169;
  assign \new_[56226]_  = ~A166 & A167;
  assign \new_[56227]_  = \new_[56226]_  & \new_[56223]_ ;
  assign \new_[56230]_  = A233 & ~A232;
  assign \new_[56233]_  = ~A235 & ~A234;
  assign \new_[56234]_  = \new_[56233]_  & \new_[56230]_ ;
  assign \new_[56235]_  = \new_[56234]_  & \new_[56227]_ ;
  assign \new_[56238]_  = A265 & A236;
  assign \new_[56241]_  = A298 & A266;
  assign \new_[56242]_  = \new_[56241]_  & \new_[56238]_ ;
  assign \new_[56245]_  = ~A300 & ~A299;
  assign \new_[56248]_  = A302 & ~A301;
  assign \new_[56249]_  = \new_[56248]_  & \new_[56245]_ ;
  assign \new_[56250]_  = \new_[56249]_  & \new_[56242]_ ;
  assign \new_[56253]_  = A168 & A169;
  assign \new_[56256]_  = ~A166 & A167;
  assign \new_[56257]_  = \new_[56256]_  & \new_[56253]_ ;
  assign \new_[56260]_  = A233 & ~A232;
  assign \new_[56263]_  = ~A235 & ~A234;
  assign \new_[56264]_  = \new_[56263]_  & \new_[56260]_ ;
  assign \new_[56265]_  = \new_[56264]_  & \new_[56257]_ ;
  assign \new_[56268]_  = A265 & A236;
  assign \new_[56271]_  = ~A298 & A266;
  assign \new_[56272]_  = \new_[56271]_  & \new_[56268]_ ;
  assign \new_[56275]_  = ~A300 & A299;
  assign \new_[56278]_  = A302 & ~A301;
  assign \new_[56279]_  = \new_[56278]_  & \new_[56275]_ ;
  assign \new_[56280]_  = \new_[56279]_  & \new_[56272]_ ;
  assign \new_[56283]_  = A168 & A169;
  assign \new_[56286]_  = ~A166 & A167;
  assign \new_[56287]_  = \new_[56286]_  & \new_[56283]_ ;
  assign \new_[56290]_  = A233 & ~A232;
  assign \new_[56293]_  = ~A235 & ~A234;
  assign \new_[56294]_  = \new_[56293]_  & \new_[56290]_ ;
  assign \new_[56295]_  = \new_[56294]_  & \new_[56287]_ ;
  assign \new_[56298]_  = ~A265 & A236;
  assign \new_[56301]_  = A298 & ~A266;
  assign \new_[56302]_  = \new_[56301]_  & \new_[56298]_ ;
  assign \new_[56305]_  = ~A300 & ~A299;
  assign \new_[56308]_  = A302 & ~A301;
  assign \new_[56309]_  = \new_[56308]_  & \new_[56305]_ ;
  assign \new_[56310]_  = \new_[56309]_  & \new_[56302]_ ;
  assign \new_[56313]_  = A168 & A169;
  assign \new_[56316]_  = ~A166 & A167;
  assign \new_[56317]_  = \new_[56316]_  & \new_[56313]_ ;
  assign \new_[56320]_  = A233 & ~A232;
  assign \new_[56323]_  = ~A235 & ~A234;
  assign \new_[56324]_  = \new_[56323]_  & \new_[56320]_ ;
  assign \new_[56325]_  = \new_[56324]_  & \new_[56317]_ ;
  assign \new_[56328]_  = ~A265 & A236;
  assign \new_[56331]_  = ~A298 & ~A266;
  assign \new_[56332]_  = \new_[56331]_  & \new_[56328]_ ;
  assign \new_[56335]_  = ~A300 & A299;
  assign \new_[56338]_  = A302 & ~A301;
  assign \new_[56339]_  = \new_[56338]_  & \new_[56335]_ ;
  assign \new_[56340]_  = \new_[56339]_  & \new_[56332]_ ;
  assign \new_[56343]_  = A168 & A169;
  assign \new_[56346]_  = ~A166 & A167;
  assign \new_[56347]_  = \new_[56346]_  & \new_[56343]_ ;
  assign \new_[56350]_  = ~A233 & A232;
  assign \new_[56353]_  = A235 & A234;
  assign \new_[56354]_  = \new_[56353]_  & \new_[56350]_ ;
  assign \new_[56355]_  = \new_[56354]_  & \new_[56347]_ ;
  assign \new_[56358]_  = ~A268 & A267;
  assign \new_[56361]_  = A298 & A269;
  assign \new_[56362]_  = \new_[56361]_  & \new_[56358]_ ;
  assign \new_[56365]_  = ~A300 & ~A299;
  assign \new_[56368]_  = A302 & ~A301;
  assign \new_[56369]_  = \new_[56368]_  & \new_[56365]_ ;
  assign \new_[56370]_  = \new_[56369]_  & \new_[56362]_ ;
  assign \new_[56373]_  = A168 & A169;
  assign \new_[56376]_  = ~A166 & A167;
  assign \new_[56377]_  = \new_[56376]_  & \new_[56373]_ ;
  assign \new_[56380]_  = ~A233 & A232;
  assign \new_[56383]_  = A235 & A234;
  assign \new_[56384]_  = \new_[56383]_  & \new_[56380]_ ;
  assign \new_[56385]_  = \new_[56384]_  & \new_[56377]_ ;
  assign \new_[56388]_  = ~A268 & A267;
  assign \new_[56391]_  = ~A298 & A269;
  assign \new_[56392]_  = \new_[56391]_  & \new_[56388]_ ;
  assign \new_[56395]_  = ~A300 & A299;
  assign \new_[56398]_  = A302 & ~A301;
  assign \new_[56399]_  = \new_[56398]_  & \new_[56395]_ ;
  assign \new_[56400]_  = \new_[56399]_  & \new_[56392]_ ;
  assign \new_[56403]_  = A168 & A169;
  assign \new_[56406]_  = ~A166 & A167;
  assign \new_[56407]_  = \new_[56406]_  & \new_[56403]_ ;
  assign \new_[56410]_  = ~A233 & A232;
  assign \new_[56413]_  = ~A236 & A234;
  assign \new_[56414]_  = \new_[56413]_  & \new_[56410]_ ;
  assign \new_[56415]_  = \new_[56414]_  & \new_[56407]_ ;
  assign \new_[56418]_  = ~A268 & A267;
  assign \new_[56421]_  = A298 & A269;
  assign \new_[56422]_  = \new_[56421]_  & \new_[56418]_ ;
  assign \new_[56425]_  = ~A300 & ~A299;
  assign \new_[56428]_  = A302 & ~A301;
  assign \new_[56429]_  = \new_[56428]_  & \new_[56425]_ ;
  assign \new_[56430]_  = \new_[56429]_  & \new_[56422]_ ;
  assign \new_[56433]_  = A168 & A169;
  assign \new_[56436]_  = ~A166 & A167;
  assign \new_[56437]_  = \new_[56436]_  & \new_[56433]_ ;
  assign \new_[56440]_  = ~A233 & A232;
  assign \new_[56443]_  = ~A236 & A234;
  assign \new_[56444]_  = \new_[56443]_  & \new_[56440]_ ;
  assign \new_[56445]_  = \new_[56444]_  & \new_[56437]_ ;
  assign \new_[56448]_  = ~A268 & A267;
  assign \new_[56451]_  = ~A298 & A269;
  assign \new_[56452]_  = \new_[56451]_  & \new_[56448]_ ;
  assign \new_[56455]_  = ~A300 & A299;
  assign \new_[56458]_  = A302 & ~A301;
  assign \new_[56459]_  = \new_[56458]_  & \new_[56455]_ ;
  assign \new_[56460]_  = \new_[56459]_  & \new_[56452]_ ;
  assign \new_[56463]_  = A168 & A169;
  assign \new_[56466]_  = ~A166 & A167;
  assign \new_[56467]_  = \new_[56466]_  & \new_[56463]_ ;
  assign \new_[56470]_  = ~A233 & A232;
  assign \new_[56473]_  = ~A235 & ~A234;
  assign \new_[56474]_  = \new_[56473]_  & \new_[56470]_ ;
  assign \new_[56475]_  = \new_[56474]_  & \new_[56467]_ ;
  assign \new_[56478]_  = A267 & A236;
  assign \new_[56481]_  = A269 & ~A268;
  assign \new_[56482]_  = \new_[56481]_  & \new_[56478]_ ;
  assign \new_[56485]_  = ~A299 & A298;
  assign \new_[56488]_  = A301 & A300;
  assign \new_[56489]_  = \new_[56488]_  & \new_[56485]_ ;
  assign \new_[56490]_  = \new_[56489]_  & \new_[56482]_ ;
  assign \new_[56493]_  = A168 & A169;
  assign \new_[56496]_  = ~A166 & A167;
  assign \new_[56497]_  = \new_[56496]_  & \new_[56493]_ ;
  assign \new_[56500]_  = ~A233 & A232;
  assign \new_[56503]_  = ~A235 & ~A234;
  assign \new_[56504]_  = \new_[56503]_  & \new_[56500]_ ;
  assign \new_[56505]_  = \new_[56504]_  & \new_[56497]_ ;
  assign \new_[56508]_  = A267 & A236;
  assign \new_[56511]_  = A269 & ~A268;
  assign \new_[56512]_  = \new_[56511]_  & \new_[56508]_ ;
  assign \new_[56515]_  = ~A299 & A298;
  assign \new_[56518]_  = ~A302 & A300;
  assign \new_[56519]_  = \new_[56518]_  & \new_[56515]_ ;
  assign \new_[56520]_  = \new_[56519]_  & \new_[56512]_ ;
  assign \new_[56523]_  = A168 & A169;
  assign \new_[56526]_  = ~A166 & A167;
  assign \new_[56527]_  = \new_[56526]_  & \new_[56523]_ ;
  assign \new_[56530]_  = ~A233 & A232;
  assign \new_[56533]_  = ~A235 & ~A234;
  assign \new_[56534]_  = \new_[56533]_  & \new_[56530]_ ;
  assign \new_[56535]_  = \new_[56534]_  & \new_[56527]_ ;
  assign \new_[56538]_  = A267 & A236;
  assign \new_[56541]_  = A269 & ~A268;
  assign \new_[56542]_  = \new_[56541]_  & \new_[56538]_ ;
  assign \new_[56545]_  = A299 & ~A298;
  assign \new_[56548]_  = A301 & A300;
  assign \new_[56549]_  = \new_[56548]_  & \new_[56545]_ ;
  assign \new_[56550]_  = \new_[56549]_  & \new_[56542]_ ;
  assign \new_[56553]_  = A168 & A169;
  assign \new_[56556]_  = ~A166 & A167;
  assign \new_[56557]_  = \new_[56556]_  & \new_[56553]_ ;
  assign \new_[56560]_  = ~A233 & A232;
  assign \new_[56563]_  = ~A235 & ~A234;
  assign \new_[56564]_  = \new_[56563]_  & \new_[56560]_ ;
  assign \new_[56565]_  = \new_[56564]_  & \new_[56557]_ ;
  assign \new_[56568]_  = A267 & A236;
  assign \new_[56571]_  = A269 & ~A268;
  assign \new_[56572]_  = \new_[56571]_  & \new_[56568]_ ;
  assign \new_[56575]_  = A299 & ~A298;
  assign \new_[56578]_  = ~A302 & A300;
  assign \new_[56579]_  = \new_[56578]_  & \new_[56575]_ ;
  assign \new_[56580]_  = \new_[56579]_  & \new_[56572]_ ;
  assign \new_[56583]_  = A168 & A169;
  assign \new_[56586]_  = ~A166 & A167;
  assign \new_[56587]_  = \new_[56586]_  & \new_[56583]_ ;
  assign \new_[56590]_  = ~A233 & A232;
  assign \new_[56593]_  = ~A235 & ~A234;
  assign \new_[56594]_  = \new_[56593]_  & \new_[56590]_ ;
  assign \new_[56595]_  = \new_[56594]_  & \new_[56587]_ ;
  assign \new_[56598]_  = ~A267 & A236;
  assign \new_[56601]_  = A298 & A268;
  assign \new_[56602]_  = \new_[56601]_  & \new_[56598]_ ;
  assign \new_[56605]_  = ~A300 & ~A299;
  assign \new_[56608]_  = A302 & ~A301;
  assign \new_[56609]_  = \new_[56608]_  & \new_[56605]_ ;
  assign \new_[56610]_  = \new_[56609]_  & \new_[56602]_ ;
  assign \new_[56613]_  = A168 & A169;
  assign \new_[56616]_  = ~A166 & A167;
  assign \new_[56617]_  = \new_[56616]_  & \new_[56613]_ ;
  assign \new_[56620]_  = ~A233 & A232;
  assign \new_[56623]_  = ~A235 & ~A234;
  assign \new_[56624]_  = \new_[56623]_  & \new_[56620]_ ;
  assign \new_[56625]_  = \new_[56624]_  & \new_[56617]_ ;
  assign \new_[56628]_  = ~A267 & A236;
  assign \new_[56631]_  = ~A298 & A268;
  assign \new_[56632]_  = \new_[56631]_  & \new_[56628]_ ;
  assign \new_[56635]_  = ~A300 & A299;
  assign \new_[56638]_  = A302 & ~A301;
  assign \new_[56639]_  = \new_[56638]_  & \new_[56635]_ ;
  assign \new_[56640]_  = \new_[56639]_  & \new_[56632]_ ;
  assign \new_[56643]_  = A168 & A169;
  assign \new_[56646]_  = ~A166 & A167;
  assign \new_[56647]_  = \new_[56646]_  & \new_[56643]_ ;
  assign \new_[56650]_  = ~A233 & A232;
  assign \new_[56653]_  = ~A235 & ~A234;
  assign \new_[56654]_  = \new_[56653]_  & \new_[56650]_ ;
  assign \new_[56655]_  = \new_[56654]_  & \new_[56647]_ ;
  assign \new_[56658]_  = ~A267 & A236;
  assign \new_[56661]_  = A298 & ~A269;
  assign \new_[56662]_  = \new_[56661]_  & \new_[56658]_ ;
  assign \new_[56665]_  = ~A300 & ~A299;
  assign \new_[56668]_  = A302 & ~A301;
  assign \new_[56669]_  = \new_[56668]_  & \new_[56665]_ ;
  assign \new_[56670]_  = \new_[56669]_  & \new_[56662]_ ;
  assign \new_[56673]_  = A168 & A169;
  assign \new_[56676]_  = ~A166 & A167;
  assign \new_[56677]_  = \new_[56676]_  & \new_[56673]_ ;
  assign \new_[56680]_  = ~A233 & A232;
  assign \new_[56683]_  = ~A235 & ~A234;
  assign \new_[56684]_  = \new_[56683]_  & \new_[56680]_ ;
  assign \new_[56685]_  = \new_[56684]_  & \new_[56677]_ ;
  assign \new_[56688]_  = ~A267 & A236;
  assign \new_[56691]_  = ~A298 & ~A269;
  assign \new_[56692]_  = \new_[56691]_  & \new_[56688]_ ;
  assign \new_[56695]_  = ~A300 & A299;
  assign \new_[56698]_  = A302 & ~A301;
  assign \new_[56699]_  = \new_[56698]_  & \new_[56695]_ ;
  assign \new_[56700]_  = \new_[56699]_  & \new_[56692]_ ;
  assign \new_[56703]_  = A168 & A169;
  assign \new_[56706]_  = ~A166 & A167;
  assign \new_[56707]_  = \new_[56706]_  & \new_[56703]_ ;
  assign \new_[56710]_  = ~A233 & A232;
  assign \new_[56713]_  = ~A235 & ~A234;
  assign \new_[56714]_  = \new_[56713]_  & \new_[56710]_ ;
  assign \new_[56715]_  = \new_[56714]_  & \new_[56707]_ ;
  assign \new_[56718]_  = A265 & A236;
  assign \new_[56721]_  = A298 & A266;
  assign \new_[56722]_  = \new_[56721]_  & \new_[56718]_ ;
  assign \new_[56725]_  = ~A300 & ~A299;
  assign \new_[56728]_  = A302 & ~A301;
  assign \new_[56729]_  = \new_[56728]_  & \new_[56725]_ ;
  assign \new_[56730]_  = \new_[56729]_  & \new_[56722]_ ;
  assign \new_[56733]_  = A168 & A169;
  assign \new_[56736]_  = ~A166 & A167;
  assign \new_[56737]_  = \new_[56736]_  & \new_[56733]_ ;
  assign \new_[56740]_  = ~A233 & A232;
  assign \new_[56743]_  = ~A235 & ~A234;
  assign \new_[56744]_  = \new_[56743]_  & \new_[56740]_ ;
  assign \new_[56745]_  = \new_[56744]_  & \new_[56737]_ ;
  assign \new_[56748]_  = A265 & A236;
  assign \new_[56751]_  = ~A298 & A266;
  assign \new_[56752]_  = \new_[56751]_  & \new_[56748]_ ;
  assign \new_[56755]_  = ~A300 & A299;
  assign \new_[56758]_  = A302 & ~A301;
  assign \new_[56759]_  = \new_[56758]_  & \new_[56755]_ ;
  assign \new_[56760]_  = \new_[56759]_  & \new_[56752]_ ;
  assign \new_[56763]_  = A168 & A169;
  assign \new_[56766]_  = ~A166 & A167;
  assign \new_[56767]_  = \new_[56766]_  & \new_[56763]_ ;
  assign \new_[56770]_  = ~A233 & A232;
  assign \new_[56773]_  = ~A235 & ~A234;
  assign \new_[56774]_  = \new_[56773]_  & \new_[56770]_ ;
  assign \new_[56775]_  = \new_[56774]_  & \new_[56767]_ ;
  assign \new_[56778]_  = ~A265 & A236;
  assign \new_[56781]_  = A298 & ~A266;
  assign \new_[56782]_  = \new_[56781]_  & \new_[56778]_ ;
  assign \new_[56785]_  = ~A300 & ~A299;
  assign \new_[56788]_  = A302 & ~A301;
  assign \new_[56789]_  = \new_[56788]_  & \new_[56785]_ ;
  assign \new_[56790]_  = \new_[56789]_  & \new_[56782]_ ;
  assign \new_[56793]_  = A168 & A169;
  assign \new_[56796]_  = ~A166 & A167;
  assign \new_[56797]_  = \new_[56796]_  & \new_[56793]_ ;
  assign \new_[56800]_  = ~A233 & A232;
  assign \new_[56803]_  = ~A235 & ~A234;
  assign \new_[56804]_  = \new_[56803]_  & \new_[56800]_ ;
  assign \new_[56805]_  = \new_[56804]_  & \new_[56797]_ ;
  assign \new_[56808]_  = ~A265 & A236;
  assign \new_[56811]_  = ~A298 & ~A266;
  assign \new_[56812]_  = \new_[56811]_  & \new_[56808]_ ;
  assign \new_[56815]_  = ~A300 & A299;
  assign \new_[56818]_  = A302 & ~A301;
  assign \new_[56819]_  = \new_[56818]_  & \new_[56815]_ ;
  assign \new_[56820]_  = \new_[56819]_  & \new_[56812]_ ;
  assign \new_[56823]_  = A168 & A169;
  assign \new_[56826]_  = A166 & ~A167;
  assign \new_[56827]_  = \new_[56826]_  & \new_[56823]_ ;
  assign \new_[56830]_  = A233 & ~A232;
  assign \new_[56833]_  = A235 & A234;
  assign \new_[56834]_  = \new_[56833]_  & \new_[56830]_ ;
  assign \new_[56835]_  = \new_[56834]_  & \new_[56827]_ ;
  assign \new_[56838]_  = ~A268 & A267;
  assign \new_[56841]_  = A298 & A269;
  assign \new_[56842]_  = \new_[56841]_  & \new_[56838]_ ;
  assign \new_[56845]_  = ~A300 & ~A299;
  assign \new_[56848]_  = A302 & ~A301;
  assign \new_[56849]_  = \new_[56848]_  & \new_[56845]_ ;
  assign \new_[56850]_  = \new_[56849]_  & \new_[56842]_ ;
  assign \new_[56853]_  = A168 & A169;
  assign \new_[56856]_  = A166 & ~A167;
  assign \new_[56857]_  = \new_[56856]_  & \new_[56853]_ ;
  assign \new_[56860]_  = A233 & ~A232;
  assign \new_[56863]_  = A235 & A234;
  assign \new_[56864]_  = \new_[56863]_  & \new_[56860]_ ;
  assign \new_[56865]_  = \new_[56864]_  & \new_[56857]_ ;
  assign \new_[56868]_  = ~A268 & A267;
  assign \new_[56871]_  = ~A298 & A269;
  assign \new_[56872]_  = \new_[56871]_  & \new_[56868]_ ;
  assign \new_[56875]_  = ~A300 & A299;
  assign \new_[56878]_  = A302 & ~A301;
  assign \new_[56879]_  = \new_[56878]_  & \new_[56875]_ ;
  assign \new_[56880]_  = \new_[56879]_  & \new_[56872]_ ;
  assign \new_[56883]_  = A168 & A169;
  assign \new_[56886]_  = A166 & ~A167;
  assign \new_[56887]_  = \new_[56886]_  & \new_[56883]_ ;
  assign \new_[56890]_  = A233 & ~A232;
  assign \new_[56893]_  = ~A236 & A234;
  assign \new_[56894]_  = \new_[56893]_  & \new_[56890]_ ;
  assign \new_[56895]_  = \new_[56894]_  & \new_[56887]_ ;
  assign \new_[56898]_  = ~A268 & A267;
  assign \new_[56901]_  = A298 & A269;
  assign \new_[56902]_  = \new_[56901]_  & \new_[56898]_ ;
  assign \new_[56905]_  = ~A300 & ~A299;
  assign \new_[56908]_  = A302 & ~A301;
  assign \new_[56909]_  = \new_[56908]_  & \new_[56905]_ ;
  assign \new_[56910]_  = \new_[56909]_  & \new_[56902]_ ;
  assign \new_[56913]_  = A168 & A169;
  assign \new_[56916]_  = A166 & ~A167;
  assign \new_[56917]_  = \new_[56916]_  & \new_[56913]_ ;
  assign \new_[56920]_  = A233 & ~A232;
  assign \new_[56923]_  = ~A236 & A234;
  assign \new_[56924]_  = \new_[56923]_  & \new_[56920]_ ;
  assign \new_[56925]_  = \new_[56924]_  & \new_[56917]_ ;
  assign \new_[56928]_  = ~A268 & A267;
  assign \new_[56931]_  = ~A298 & A269;
  assign \new_[56932]_  = \new_[56931]_  & \new_[56928]_ ;
  assign \new_[56935]_  = ~A300 & A299;
  assign \new_[56938]_  = A302 & ~A301;
  assign \new_[56939]_  = \new_[56938]_  & \new_[56935]_ ;
  assign \new_[56940]_  = \new_[56939]_  & \new_[56932]_ ;
  assign \new_[56943]_  = A168 & A169;
  assign \new_[56946]_  = A166 & ~A167;
  assign \new_[56947]_  = \new_[56946]_  & \new_[56943]_ ;
  assign \new_[56950]_  = A233 & ~A232;
  assign \new_[56953]_  = ~A235 & ~A234;
  assign \new_[56954]_  = \new_[56953]_  & \new_[56950]_ ;
  assign \new_[56955]_  = \new_[56954]_  & \new_[56947]_ ;
  assign \new_[56958]_  = A267 & A236;
  assign \new_[56961]_  = A269 & ~A268;
  assign \new_[56962]_  = \new_[56961]_  & \new_[56958]_ ;
  assign \new_[56965]_  = ~A299 & A298;
  assign \new_[56968]_  = A301 & A300;
  assign \new_[56969]_  = \new_[56968]_  & \new_[56965]_ ;
  assign \new_[56970]_  = \new_[56969]_  & \new_[56962]_ ;
  assign \new_[56973]_  = A168 & A169;
  assign \new_[56976]_  = A166 & ~A167;
  assign \new_[56977]_  = \new_[56976]_  & \new_[56973]_ ;
  assign \new_[56980]_  = A233 & ~A232;
  assign \new_[56983]_  = ~A235 & ~A234;
  assign \new_[56984]_  = \new_[56983]_  & \new_[56980]_ ;
  assign \new_[56985]_  = \new_[56984]_  & \new_[56977]_ ;
  assign \new_[56988]_  = A267 & A236;
  assign \new_[56991]_  = A269 & ~A268;
  assign \new_[56992]_  = \new_[56991]_  & \new_[56988]_ ;
  assign \new_[56995]_  = ~A299 & A298;
  assign \new_[56998]_  = ~A302 & A300;
  assign \new_[56999]_  = \new_[56998]_  & \new_[56995]_ ;
  assign \new_[57000]_  = \new_[56999]_  & \new_[56992]_ ;
  assign \new_[57003]_  = A168 & A169;
  assign \new_[57006]_  = A166 & ~A167;
  assign \new_[57007]_  = \new_[57006]_  & \new_[57003]_ ;
  assign \new_[57010]_  = A233 & ~A232;
  assign \new_[57013]_  = ~A235 & ~A234;
  assign \new_[57014]_  = \new_[57013]_  & \new_[57010]_ ;
  assign \new_[57015]_  = \new_[57014]_  & \new_[57007]_ ;
  assign \new_[57018]_  = A267 & A236;
  assign \new_[57021]_  = A269 & ~A268;
  assign \new_[57022]_  = \new_[57021]_  & \new_[57018]_ ;
  assign \new_[57025]_  = A299 & ~A298;
  assign \new_[57028]_  = A301 & A300;
  assign \new_[57029]_  = \new_[57028]_  & \new_[57025]_ ;
  assign \new_[57030]_  = \new_[57029]_  & \new_[57022]_ ;
  assign \new_[57033]_  = A168 & A169;
  assign \new_[57036]_  = A166 & ~A167;
  assign \new_[57037]_  = \new_[57036]_  & \new_[57033]_ ;
  assign \new_[57040]_  = A233 & ~A232;
  assign \new_[57043]_  = ~A235 & ~A234;
  assign \new_[57044]_  = \new_[57043]_  & \new_[57040]_ ;
  assign \new_[57045]_  = \new_[57044]_  & \new_[57037]_ ;
  assign \new_[57048]_  = A267 & A236;
  assign \new_[57051]_  = A269 & ~A268;
  assign \new_[57052]_  = \new_[57051]_  & \new_[57048]_ ;
  assign \new_[57055]_  = A299 & ~A298;
  assign \new_[57058]_  = ~A302 & A300;
  assign \new_[57059]_  = \new_[57058]_  & \new_[57055]_ ;
  assign \new_[57060]_  = \new_[57059]_  & \new_[57052]_ ;
  assign \new_[57063]_  = A168 & A169;
  assign \new_[57066]_  = A166 & ~A167;
  assign \new_[57067]_  = \new_[57066]_  & \new_[57063]_ ;
  assign \new_[57070]_  = A233 & ~A232;
  assign \new_[57073]_  = ~A235 & ~A234;
  assign \new_[57074]_  = \new_[57073]_  & \new_[57070]_ ;
  assign \new_[57075]_  = \new_[57074]_  & \new_[57067]_ ;
  assign \new_[57078]_  = ~A267 & A236;
  assign \new_[57081]_  = A298 & A268;
  assign \new_[57082]_  = \new_[57081]_  & \new_[57078]_ ;
  assign \new_[57085]_  = ~A300 & ~A299;
  assign \new_[57088]_  = A302 & ~A301;
  assign \new_[57089]_  = \new_[57088]_  & \new_[57085]_ ;
  assign \new_[57090]_  = \new_[57089]_  & \new_[57082]_ ;
  assign \new_[57093]_  = A168 & A169;
  assign \new_[57096]_  = A166 & ~A167;
  assign \new_[57097]_  = \new_[57096]_  & \new_[57093]_ ;
  assign \new_[57100]_  = A233 & ~A232;
  assign \new_[57103]_  = ~A235 & ~A234;
  assign \new_[57104]_  = \new_[57103]_  & \new_[57100]_ ;
  assign \new_[57105]_  = \new_[57104]_  & \new_[57097]_ ;
  assign \new_[57108]_  = ~A267 & A236;
  assign \new_[57111]_  = ~A298 & A268;
  assign \new_[57112]_  = \new_[57111]_  & \new_[57108]_ ;
  assign \new_[57115]_  = ~A300 & A299;
  assign \new_[57118]_  = A302 & ~A301;
  assign \new_[57119]_  = \new_[57118]_  & \new_[57115]_ ;
  assign \new_[57120]_  = \new_[57119]_  & \new_[57112]_ ;
  assign \new_[57123]_  = A168 & A169;
  assign \new_[57126]_  = A166 & ~A167;
  assign \new_[57127]_  = \new_[57126]_  & \new_[57123]_ ;
  assign \new_[57130]_  = A233 & ~A232;
  assign \new_[57133]_  = ~A235 & ~A234;
  assign \new_[57134]_  = \new_[57133]_  & \new_[57130]_ ;
  assign \new_[57135]_  = \new_[57134]_  & \new_[57127]_ ;
  assign \new_[57138]_  = ~A267 & A236;
  assign \new_[57141]_  = A298 & ~A269;
  assign \new_[57142]_  = \new_[57141]_  & \new_[57138]_ ;
  assign \new_[57145]_  = ~A300 & ~A299;
  assign \new_[57148]_  = A302 & ~A301;
  assign \new_[57149]_  = \new_[57148]_  & \new_[57145]_ ;
  assign \new_[57150]_  = \new_[57149]_  & \new_[57142]_ ;
  assign \new_[57153]_  = A168 & A169;
  assign \new_[57156]_  = A166 & ~A167;
  assign \new_[57157]_  = \new_[57156]_  & \new_[57153]_ ;
  assign \new_[57160]_  = A233 & ~A232;
  assign \new_[57163]_  = ~A235 & ~A234;
  assign \new_[57164]_  = \new_[57163]_  & \new_[57160]_ ;
  assign \new_[57165]_  = \new_[57164]_  & \new_[57157]_ ;
  assign \new_[57168]_  = ~A267 & A236;
  assign \new_[57171]_  = ~A298 & ~A269;
  assign \new_[57172]_  = \new_[57171]_  & \new_[57168]_ ;
  assign \new_[57175]_  = ~A300 & A299;
  assign \new_[57178]_  = A302 & ~A301;
  assign \new_[57179]_  = \new_[57178]_  & \new_[57175]_ ;
  assign \new_[57180]_  = \new_[57179]_  & \new_[57172]_ ;
  assign \new_[57183]_  = A168 & A169;
  assign \new_[57186]_  = A166 & ~A167;
  assign \new_[57187]_  = \new_[57186]_  & \new_[57183]_ ;
  assign \new_[57190]_  = A233 & ~A232;
  assign \new_[57193]_  = ~A235 & ~A234;
  assign \new_[57194]_  = \new_[57193]_  & \new_[57190]_ ;
  assign \new_[57195]_  = \new_[57194]_  & \new_[57187]_ ;
  assign \new_[57198]_  = A265 & A236;
  assign \new_[57201]_  = A298 & A266;
  assign \new_[57202]_  = \new_[57201]_  & \new_[57198]_ ;
  assign \new_[57205]_  = ~A300 & ~A299;
  assign \new_[57208]_  = A302 & ~A301;
  assign \new_[57209]_  = \new_[57208]_  & \new_[57205]_ ;
  assign \new_[57210]_  = \new_[57209]_  & \new_[57202]_ ;
  assign \new_[57213]_  = A168 & A169;
  assign \new_[57216]_  = A166 & ~A167;
  assign \new_[57217]_  = \new_[57216]_  & \new_[57213]_ ;
  assign \new_[57220]_  = A233 & ~A232;
  assign \new_[57223]_  = ~A235 & ~A234;
  assign \new_[57224]_  = \new_[57223]_  & \new_[57220]_ ;
  assign \new_[57225]_  = \new_[57224]_  & \new_[57217]_ ;
  assign \new_[57228]_  = A265 & A236;
  assign \new_[57231]_  = ~A298 & A266;
  assign \new_[57232]_  = \new_[57231]_  & \new_[57228]_ ;
  assign \new_[57235]_  = ~A300 & A299;
  assign \new_[57238]_  = A302 & ~A301;
  assign \new_[57239]_  = \new_[57238]_  & \new_[57235]_ ;
  assign \new_[57240]_  = \new_[57239]_  & \new_[57232]_ ;
  assign \new_[57243]_  = A168 & A169;
  assign \new_[57246]_  = A166 & ~A167;
  assign \new_[57247]_  = \new_[57246]_  & \new_[57243]_ ;
  assign \new_[57250]_  = A233 & ~A232;
  assign \new_[57253]_  = ~A235 & ~A234;
  assign \new_[57254]_  = \new_[57253]_  & \new_[57250]_ ;
  assign \new_[57255]_  = \new_[57254]_  & \new_[57247]_ ;
  assign \new_[57258]_  = ~A265 & A236;
  assign \new_[57261]_  = A298 & ~A266;
  assign \new_[57262]_  = \new_[57261]_  & \new_[57258]_ ;
  assign \new_[57265]_  = ~A300 & ~A299;
  assign \new_[57268]_  = A302 & ~A301;
  assign \new_[57269]_  = \new_[57268]_  & \new_[57265]_ ;
  assign \new_[57270]_  = \new_[57269]_  & \new_[57262]_ ;
  assign \new_[57273]_  = A168 & A169;
  assign \new_[57276]_  = A166 & ~A167;
  assign \new_[57277]_  = \new_[57276]_  & \new_[57273]_ ;
  assign \new_[57280]_  = A233 & ~A232;
  assign \new_[57283]_  = ~A235 & ~A234;
  assign \new_[57284]_  = \new_[57283]_  & \new_[57280]_ ;
  assign \new_[57285]_  = \new_[57284]_  & \new_[57277]_ ;
  assign \new_[57288]_  = ~A265 & A236;
  assign \new_[57291]_  = ~A298 & ~A266;
  assign \new_[57292]_  = \new_[57291]_  & \new_[57288]_ ;
  assign \new_[57295]_  = ~A300 & A299;
  assign \new_[57298]_  = A302 & ~A301;
  assign \new_[57299]_  = \new_[57298]_  & \new_[57295]_ ;
  assign \new_[57300]_  = \new_[57299]_  & \new_[57292]_ ;
  assign \new_[57303]_  = A168 & A169;
  assign \new_[57306]_  = A166 & ~A167;
  assign \new_[57307]_  = \new_[57306]_  & \new_[57303]_ ;
  assign \new_[57310]_  = ~A233 & A232;
  assign \new_[57313]_  = A235 & A234;
  assign \new_[57314]_  = \new_[57313]_  & \new_[57310]_ ;
  assign \new_[57315]_  = \new_[57314]_  & \new_[57307]_ ;
  assign \new_[57318]_  = ~A268 & A267;
  assign \new_[57321]_  = A298 & A269;
  assign \new_[57322]_  = \new_[57321]_  & \new_[57318]_ ;
  assign \new_[57325]_  = ~A300 & ~A299;
  assign \new_[57328]_  = A302 & ~A301;
  assign \new_[57329]_  = \new_[57328]_  & \new_[57325]_ ;
  assign \new_[57330]_  = \new_[57329]_  & \new_[57322]_ ;
  assign \new_[57333]_  = A168 & A169;
  assign \new_[57336]_  = A166 & ~A167;
  assign \new_[57337]_  = \new_[57336]_  & \new_[57333]_ ;
  assign \new_[57340]_  = ~A233 & A232;
  assign \new_[57343]_  = A235 & A234;
  assign \new_[57344]_  = \new_[57343]_  & \new_[57340]_ ;
  assign \new_[57345]_  = \new_[57344]_  & \new_[57337]_ ;
  assign \new_[57348]_  = ~A268 & A267;
  assign \new_[57351]_  = ~A298 & A269;
  assign \new_[57352]_  = \new_[57351]_  & \new_[57348]_ ;
  assign \new_[57355]_  = ~A300 & A299;
  assign \new_[57358]_  = A302 & ~A301;
  assign \new_[57359]_  = \new_[57358]_  & \new_[57355]_ ;
  assign \new_[57360]_  = \new_[57359]_  & \new_[57352]_ ;
  assign \new_[57363]_  = A168 & A169;
  assign \new_[57366]_  = A166 & ~A167;
  assign \new_[57367]_  = \new_[57366]_  & \new_[57363]_ ;
  assign \new_[57370]_  = ~A233 & A232;
  assign \new_[57373]_  = ~A236 & A234;
  assign \new_[57374]_  = \new_[57373]_  & \new_[57370]_ ;
  assign \new_[57375]_  = \new_[57374]_  & \new_[57367]_ ;
  assign \new_[57378]_  = ~A268 & A267;
  assign \new_[57381]_  = A298 & A269;
  assign \new_[57382]_  = \new_[57381]_  & \new_[57378]_ ;
  assign \new_[57385]_  = ~A300 & ~A299;
  assign \new_[57388]_  = A302 & ~A301;
  assign \new_[57389]_  = \new_[57388]_  & \new_[57385]_ ;
  assign \new_[57390]_  = \new_[57389]_  & \new_[57382]_ ;
  assign \new_[57393]_  = A168 & A169;
  assign \new_[57396]_  = A166 & ~A167;
  assign \new_[57397]_  = \new_[57396]_  & \new_[57393]_ ;
  assign \new_[57400]_  = ~A233 & A232;
  assign \new_[57403]_  = ~A236 & A234;
  assign \new_[57404]_  = \new_[57403]_  & \new_[57400]_ ;
  assign \new_[57405]_  = \new_[57404]_  & \new_[57397]_ ;
  assign \new_[57408]_  = ~A268 & A267;
  assign \new_[57411]_  = ~A298 & A269;
  assign \new_[57412]_  = \new_[57411]_  & \new_[57408]_ ;
  assign \new_[57415]_  = ~A300 & A299;
  assign \new_[57418]_  = A302 & ~A301;
  assign \new_[57419]_  = \new_[57418]_  & \new_[57415]_ ;
  assign \new_[57420]_  = \new_[57419]_  & \new_[57412]_ ;
  assign \new_[57423]_  = A168 & A169;
  assign \new_[57426]_  = A166 & ~A167;
  assign \new_[57427]_  = \new_[57426]_  & \new_[57423]_ ;
  assign \new_[57430]_  = ~A233 & A232;
  assign \new_[57433]_  = ~A235 & ~A234;
  assign \new_[57434]_  = \new_[57433]_  & \new_[57430]_ ;
  assign \new_[57435]_  = \new_[57434]_  & \new_[57427]_ ;
  assign \new_[57438]_  = A267 & A236;
  assign \new_[57441]_  = A269 & ~A268;
  assign \new_[57442]_  = \new_[57441]_  & \new_[57438]_ ;
  assign \new_[57445]_  = ~A299 & A298;
  assign \new_[57448]_  = A301 & A300;
  assign \new_[57449]_  = \new_[57448]_  & \new_[57445]_ ;
  assign \new_[57450]_  = \new_[57449]_  & \new_[57442]_ ;
  assign \new_[57453]_  = A168 & A169;
  assign \new_[57456]_  = A166 & ~A167;
  assign \new_[57457]_  = \new_[57456]_  & \new_[57453]_ ;
  assign \new_[57460]_  = ~A233 & A232;
  assign \new_[57463]_  = ~A235 & ~A234;
  assign \new_[57464]_  = \new_[57463]_  & \new_[57460]_ ;
  assign \new_[57465]_  = \new_[57464]_  & \new_[57457]_ ;
  assign \new_[57468]_  = A267 & A236;
  assign \new_[57471]_  = A269 & ~A268;
  assign \new_[57472]_  = \new_[57471]_  & \new_[57468]_ ;
  assign \new_[57475]_  = ~A299 & A298;
  assign \new_[57478]_  = ~A302 & A300;
  assign \new_[57479]_  = \new_[57478]_  & \new_[57475]_ ;
  assign \new_[57480]_  = \new_[57479]_  & \new_[57472]_ ;
  assign \new_[57483]_  = A168 & A169;
  assign \new_[57486]_  = A166 & ~A167;
  assign \new_[57487]_  = \new_[57486]_  & \new_[57483]_ ;
  assign \new_[57490]_  = ~A233 & A232;
  assign \new_[57493]_  = ~A235 & ~A234;
  assign \new_[57494]_  = \new_[57493]_  & \new_[57490]_ ;
  assign \new_[57495]_  = \new_[57494]_  & \new_[57487]_ ;
  assign \new_[57498]_  = A267 & A236;
  assign \new_[57501]_  = A269 & ~A268;
  assign \new_[57502]_  = \new_[57501]_  & \new_[57498]_ ;
  assign \new_[57505]_  = A299 & ~A298;
  assign \new_[57508]_  = A301 & A300;
  assign \new_[57509]_  = \new_[57508]_  & \new_[57505]_ ;
  assign \new_[57510]_  = \new_[57509]_  & \new_[57502]_ ;
  assign \new_[57513]_  = A168 & A169;
  assign \new_[57516]_  = A166 & ~A167;
  assign \new_[57517]_  = \new_[57516]_  & \new_[57513]_ ;
  assign \new_[57520]_  = ~A233 & A232;
  assign \new_[57523]_  = ~A235 & ~A234;
  assign \new_[57524]_  = \new_[57523]_  & \new_[57520]_ ;
  assign \new_[57525]_  = \new_[57524]_  & \new_[57517]_ ;
  assign \new_[57528]_  = A267 & A236;
  assign \new_[57531]_  = A269 & ~A268;
  assign \new_[57532]_  = \new_[57531]_  & \new_[57528]_ ;
  assign \new_[57535]_  = A299 & ~A298;
  assign \new_[57538]_  = ~A302 & A300;
  assign \new_[57539]_  = \new_[57538]_  & \new_[57535]_ ;
  assign \new_[57540]_  = \new_[57539]_  & \new_[57532]_ ;
  assign \new_[57543]_  = A168 & A169;
  assign \new_[57546]_  = A166 & ~A167;
  assign \new_[57547]_  = \new_[57546]_  & \new_[57543]_ ;
  assign \new_[57550]_  = ~A233 & A232;
  assign \new_[57553]_  = ~A235 & ~A234;
  assign \new_[57554]_  = \new_[57553]_  & \new_[57550]_ ;
  assign \new_[57555]_  = \new_[57554]_  & \new_[57547]_ ;
  assign \new_[57558]_  = ~A267 & A236;
  assign \new_[57561]_  = A298 & A268;
  assign \new_[57562]_  = \new_[57561]_  & \new_[57558]_ ;
  assign \new_[57565]_  = ~A300 & ~A299;
  assign \new_[57568]_  = A302 & ~A301;
  assign \new_[57569]_  = \new_[57568]_  & \new_[57565]_ ;
  assign \new_[57570]_  = \new_[57569]_  & \new_[57562]_ ;
  assign \new_[57573]_  = A168 & A169;
  assign \new_[57576]_  = A166 & ~A167;
  assign \new_[57577]_  = \new_[57576]_  & \new_[57573]_ ;
  assign \new_[57580]_  = ~A233 & A232;
  assign \new_[57583]_  = ~A235 & ~A234;
  assign \new_[57584]_  = \new_[57583]_  & \new_[57580]_ ;
  assign \new_[57585]_  = \new_[57584]_  & \new_[57577]_ ;
  assign \new_[57588]_  = ~A267 & A236;
  assign \new_[57591]_  = ~A298 & A268;
  assign \new_[57592]_  = \new_[57591]_  & \new_[57588]_ ;
  assign \new_[57595]_  = ~A300 & A299;
  assign \new_[57598]_  = A302 & ~A301;
  assign \new_[57599]_  = \new_[57598]_  & \new_[57595]_ ;
  assign \new_[57600]_  = \new_[57599]_  & \new_[57592]_ ;
  assign \new_[57603]_  = A168 & A169;
  assign \new_[57606]_  = A166 & ~A167;
  assign \new_[57607]_  = \new_[57606]_  & \new_[57603]_ ;
  assign \new_[57610]_  = ~A233 & A232;
  assign \new_[57613]_  = ~A235 & ~A234;
  assign \new_[57614]_  = \new_[57613]_  & \new_[57610]_ ;
  assign \new_[57615]_  = \new_[57614]_  & \new_[57607]_ ;
  assign \new_[57618]_  = ~A267 & A236;
  assign \new_[57621]_  = A298 & ~A269;
  assign \new_[57622]_  = \new_[57621]_  & \new_[57618]_ ;
  assign \new_[57625]_  = ~A300 & ~A299;
  assign \new_[57628]_  = A302 & ~A301;
  assign \new_[57629]_  = \new_[57628]_  & \new_[57625]_ ;
  assign \new_[57630]_  = \new_[57629]_  & \new_[57622]_ ;
  assign \new_[57633]_  = A168 & A169;
  assign \new_[57636]_  = A166 & ~A167;
  assign \new_[57637]_  = \new_[57636]_  & \new_[57633]_ ;
  assign \new_[57640]_  = ~A233 & A232;
  assign \new_[57643]_  = ~A235 & ~A234;
  assign \new_[57644]_  = \new_[57643]_  & \new_[57640]_ ;
  assign \new_[57645]_  = \new_[57644]_  & \new_[57637]_ ;
  assign \new_[57648]_  = ~A267 & A236;
  assign \new_[57651]_  = ~A298 & ~A269;
  assign \new_[57652]_  = \new_[57651]_  & \new_[57648]_ ;
  assign \new_[57655]_  = ~A300 & A299;
  assign \new_[57658]_  = A302 & ~A301;
  assign \new_[57659]_  = \new_[57658]_  & \new_[57655]_ ;
  assign \new_[57660]_  = \new_[57659]_  & \new_[57652]_ ;
  assign \new_[57663]_  = A168 & A169;
  assign \new_[57666]_  = A166 & ~A167;
  assign \new_[57667]_  = \new_[57666]_  & \new_[57663]_ ;
  assign \new_[57670]_  = ~A233 & A232;
  assign \new_[57673]_  = ~A235 & ~A234;
  assign \new_[57674]_  = \new_[57673]_  & \new_[57670]_ ;
  assign \new_[57675]_  = \new_[57674]_  & \new_[57667]_ ;
  assign \new_[57678]_  = A265 & A236;
  assign \new_[57681]_  = A298 & A266;
  assign \new_[57682]_  = \new_[57681]_  & \new_[57678]_ ;
  assign \new_[57685]_  = ~A300 & ~A299;
  assign \new_[57688]_  = A302 & ~A301;
  assign \new_[57689]_  = \new_[57688]_  & \new_[57685]_ ;
  assign \new_[57690]_  = \new_[57689]_  & \new_[57682]_ ;
  assign \new_[57693]_  = A168 & A169;
  assign \new_[57696]_  = A166 & ~A167;
  assign \new_[57697]_  = \new_[57696]_  & \new_[57693]_ ;
  assign \new_[57700]_  = ~A233 & A232;
  assign \new_[57703]_  = ~A235 & ~A234;
  assign \new_[57704]_  = \new_[57703]_  & \new_[57700]_ ;
  assign \new_[57705]_  = \new_[57704]_  & \new_[57697]_ ;
  assign \new_[57708]_  = A265 & A236;
  assign \new_[57711]_  = ~A298 & A266;
  assign \new_[57712]_  = \new_[57711]_  & \new_[57708]_ ;
  assign \new_[57715]_  = ~A300 & A299;
  assign \new_[57718]_  = A302 & ~A301;
  assign \new_[57719]_  = \new_[57718]_  & \new_[57715]_ ;
  assign \new_[57720]_  = \new_[57719]_  & \new_[57712]_ ;
  assign \new_[57723]_  = A168 & A169;
  assign \new_[57726]_  = A166 & ~A167;
  assign \new_[57727]_  = \new_[57726]_  & \new_[57723]_ ;
  assign \new_[57730]_  = ~A233 & A232;
  assign \new_[57733]_  = ~A235 & ~A234;
  assign \new_[57734]_  = \new_[57733]_  & \new_[57730]_ ;
  assign \new_[57735]_  = \new_[57734]_  & \new_[57727]_ ;
  assign \new_[57738]_  = ~A265 & A236;
  assign \new_[57741]_  = A298 & ~A266;
  assign \new_[57742]_  = \new_[57741]_  & \new_[57738]_ ;
  assign \new_[57745]_  = ~A300 & ~A299;
  assign \new_[57748]_  = A302 & ~A301;
  assign \new_[57749]_  = \new_[57748]_  & \new_[57745]_ ;
  assign \new_[57750]_  = \new_[57749]_  & \new_[57742]_ ;
  assign \new_[57753]_  = A168 & A169;
  assign \new_[57756]_  = A166 & ~A167;
  assign \new_[57757]_  = \new_[57756]_  & \new_[57753]_ ;
  assign \new_[57760]_  = ~A233 & A232;
  assign \new_[57763]_  = ~A235 & ~A234;
  assign \new_[57764]_  = \new_[57763]_  & \new_[57760]_ ;
  assign \new_[57765]_  = \new_[57764]_  & \new_[57757]_ ;
  assign \new_[57768]_  = ~A265 & A236;
  assign \new_[57771]_  = ~A298 & ~A266;
  assign \new_[57772]_  = \new_[57771]_  & \new_[57768]_ ;
  assign \new_[57775]_  = ~A300 & A299;
  assign \new_[57778]_  = A302 & ~A301;
  assign \new_[57779]_  = \new_[57778]_  & \new_[57775]_ ;
  assign \new_[57780]_  = \new_[57779]_  & \new_[57772]_ ;
  assign \new_[57783]_  = ~A169 & ~A170;
  assign \new_[57786]_  = A167 & ~A168;
  assign \new_[57787]_  = \new_[57786]_  & \new_[57783]_ ;
  assign \new_[57790]_  = ~A232 & ~A166;
  assign \new_[57793]_  = A234 & A233;
  assign \new_[57794]_  = \new_[57793]_  & \new_[57790]_ ;
  assign \new_[57795]_  = \new_[57794]_  & \new_[57787]_ ;
  assign \new_[57798]_  = A267 & A235;
  assign \new_[57801]_  = A269 & ~A268;
  assign \new_[57802]_  = \new_[57801]_  & \new_[57798]_ ;
  assign \new_[57805]_  = ~A299 & A298;
  assign \new_[57808]_  = A301 & A300;
  assign \new_[57809]_  = \new_[57808]_  & \new_[57805]_ ;
  assign \new_[57810]_  = \new_[57809]_  & \new_[57802]_ ;
  assign \new_[57813]_  = ~A169 & ~A170;
  assign \new_[57816]_  = A167 & ~A168;
  assign \new_[57817]_  = \new_[57816]_  & \new_[57813]_ ;
  assign \new_[57820]_  = ~A232 & ~A166;
  assign \new_[57823]_  = A234 & A233;
  assign \new_[57824]_  = \new_[57823]_  & \new_[57820]_ ;
  assign \new_[57825]_  = \new_[57824]_  & \new_[57817]_ ;
  assign \new_[57828]_  = A267 & A235;
  assign \new_[57831]_  = A269 & ~A268;
  assign \new_[57832]_  = \new_[57831]_  & \new_[57828]_ ;
  assign \new_[57835]_  = ~A299 & A298;
  assign \new_[57838]_  = ~A302 & A300;
  assign \new_[57839]_  = \new_[57838]_  & \new_[57835]_ ;
  assign \new_[57840]_  = \new_[57839]_  & \new_[57832]_ ;
  assign \new_[57843]_  = ~A169 & ~A170;
  assign \new_[57846]_  = A167 & ~A168;
  assign \new_[57847]_  = \new_[57846]_  & \new_[57843]_ ;
  assign \new_[57850]_  = ~A232 & ~A166;
  assign \new_[57853]_  = A234 & A233;
  assign \new_[57854]_  = \new_[57853]_  & \new_[57850]_ ;
  assign \new_[57855]_  = \new_[57854]_  & \new_[57847]_ ;
  assign \new_[57858]_  = A267 & A235;
  assign \new_[57861]_  = A269 & ~A268;
  assign \new_[57862]_  = \new_[57861]_  & \new_[57858]_ ;
  assign \new_[57865]_  = A299 & ~A298;
  assign \new_[57868]_  = A301 & A300;
  assign \new_[57869]_  = \new_[57868]_  & \new_[57865]_ ;
  assign \new_[57870]_  = \new_[57869]_  & \new_[57862]_ ;
  assign \new_[57873]_  = ~A169 & ~A170;
  assign \new_[57876]_  = A167 & ~A168;
  assign \new_[57877]_  = \new_[57876]_  & \new_[57873]_ ;
  assign \new_[57880]_  = ~A232 & ~A166;
  assign \new_[57883]_  = A234 & A233;
  assign \new_[57884]_  = \new_[57883]_  & \new_[57880]_ ;
  assign \new_[57885]_  = \new_[57884]_  & \new_[57877]_ ;
  assign \new_[57888]_  = A267 & A235;
  assign \new_[57891]_  = A269 & ~A268;
  assign \new_[57892]_  = \new_[57891]_  & \new_[57888]_ ;
  assign \new_[57895]_  = A299 & ~A298;
  assign \new_[57898]_  = ~A302 & A300;
  assign \new_[57899]_  = \new_[57898]_  & \new_[57895]_ ;
  assign \new_[57900]_  = \new_[57899]_  & \new_[57892]_ ;
  assign \new_[57903]_  = ~A169 & ~A170;
  assign \new_[57906]_  = A167 & ~A168;
  assign \new_[57907]_  = \new_[57906]_  & \new_[57903]_ ;
  assign \new_[57910]_  = ~A232 & ~A166;
  assign \new_[57913]_  = A234 & A233;
  assign \new_[57914]_  = \new_[57913]_  & \new_[57910]_ ;
  assign \new_[57915]_  = \new_[57914]_  & \new_[57907]_ ;
  assign \new_[57918]_  = ~A267 & A235;
  assign \new_[57921]_  = A298 & A268;
  assign \new_[57922]_  = \new_[57921]_  & \new_[57918]_ ;
  assign \new_[57925]_  = ~A300 & ~A299;
  assign \new_[57928]_  = A302 & ~A301;
  assign \new_[57929]_  = \new_[57928]_  & \new_[57925]_ ;
  assign \new_[57930]_  = \new_[57929]_  & \new_[57922]_ ;
  assign \new_[57933]_  = ~A169 & ~A170;
  assign \new_[57936]_  = A167 & ~A168;
  assign \new_[57937]_  = \new_[57936]_  & \new_[57933]_ ;
  assign \new_[57940]_  = ~A232 & ~A166;
  assign \new_[57943]_  = A234 & A233;
  assign \new_[57944]_  = \new_[57943]_  & \new_[57940]_ ;
  assign \new_[57945]_  = \new_[57944]_  & \new_[57937]_ ;
  assign \new_[57948]_  = ~A267 & A235;
  assign \new_[57951]_  = ~A298 & A268;
  assign \new_[57952]_  = \new_[57951]_  & \new_[57948]_ ;
  assign \new_[57955]_  = ~A300 & A299;
  assign \new_[57958]_  = A302 & ~A301;
  assign \new_[57959]_  = \new_[57958]_  & \new_[57955]_ ;
  assign \new_[57960]_  = \new_[57959]_  & \new_[57952]_ ;
  assign \new_[57963]_  = ~A169 & ~A170;
  assign \new_[57966]_  = A167 & ~A168;
  assign \new_[57967]_  = \new_[57966]_  & \new_[57963]_ ;
  assign \new_[57970]_  = ~A232 & ~A166;
  assign \new_[57973]_  = A234 & A233;
  assign \new_[57974]_  = \new_[57973]_  & \new_[57970]_ ;
  assign \new_[57975]_  = \new_[57974]_  & \new_[57967]_ ;
  assign \new_[57978]_  = ~A267 & A235;
  assign \new_[57981]_  = A298 & ~A269;
  assign \new_[57982]_  = \new_[57981]_  & \new_[57978]_ ;
  assign \new_[57985]_  = ~A300 & ~A299;
  assign \new_[57988]_  = A302 & ~A301;
  assign \new_[57989]_  = \new_[57988]_  & \new_[57985]_ ;
  assign \new_[57990]_  = \new_[57989]_  & \new_[57982]_ ;
  assign \new_[57993]_  = ~A169 & ~A170;
  assign \new_[57996]_  = A167 & ~A168;
  assign \new_[57997]_  = \new_[57996]_  & \new_[57993]_ ;
  assign \new_[58000]_  = ~A232 & ~A166;
  assign \new_[58003]_  = A234 & A233;
  assign \new_[58004]_  = \new_[58003]_  & \new_[58000]_ ;
  assign \new_[58005]_  = \new_[58004]_  & \new_[57997]_ ;
  assign \new_[58008]_  = ~A267 & A235;
  assign \new_[58011]_  = ~A298 & ~A269;
  assign \new_[58012]_  = \new_[58011]_  & \new_[58008]_ ;
  assign \new_[58015]_  = ~A300 & A299;
  assign \new_[58018]_  = A302 & ~A301;
  assign \new_[58019]_  = \new_[58018]_  & \new_[58015]_ ;
  assign \new_[58020]_  = \new_[58019]_  & \new_[58012]_ ;
  assign \new_[58023]_  = ~A169 & ~A170;
  assign \new_[58026]_  = A167 & ~A168;
  assign \new_[58027]_  = \new_[58026]_  & \new_[58023]_ ;
  assign \new_[58030]_  = ~A232 & ~A166;
  assign \new_[58033]_  = A234 & A233;
  assign \new_[58034]_  = \new_[58033]_  & \new_[58030]_ ;
  assign \new_[58035]_  = \new_[58034]_  & \new_[58027]_ ;
  assign \new_[58038]_  = A265 & A235;
  assign \new_[58041]_  = A298 & A266;
  assign \new_[58042]_  = \new_[58041]_  & \new_[58038]_ ;
  assign \new_[58045]_  = ~A300 & ~A299;
  assign \new_[58048]_  = A302 & ~A301;
  assign \new_[58049]_  = \new_[58048]_  & \new_[58045]_ ;
  assign \new_[58050]_  = \new_[58049]_  & \new_[58042]_ ;
  assign \new_[58053]_  = ~A169 & ~A170;
  assign \new_[58056]_  = A167 & ~A168;
  assign \new_[58057]_  = \new_[58056]_  & \new_[58053]_ ;
  assign \new_[58060]_  = ~A232 & ~A166;
  assign \new_[58063]_  = A234 & A233;
  assign \new_[58064]_  = \new_[58063]_  & \new_[58060]_ ;
  assign \new_[58065]_  = \new_[58064]_  & \new_[58057]_ ;
  assign \new_[58068]_  = A265 & A235;
  assign \new_[58071]_  = ~A298 & A266;
  assign \new_[58072]_  = \new_[58071]_  & \new_[58068]_ ;
  assign \new_[58075]_  = ~A300 & A299;
  assign \new_[58078]_  = A302 & ~A301;
  assign \new_[58079]_  = \new_[58078]_  & \new_[58075]_ ;
  assign \new_[58080]_  = \new_[58079]_  & \new_[58072]_ ;
  assign \new_[58083]_  = ~A169 & ~A170;
  assign \new_[58086]_  = A167 & ~A168;
  assign \new_[58087]_  = \new_[58086]_  & \new_[58083]_ ;
  assign \new_[58090]_  = ~A232 & ~A166;
  assign \new_[58093]_  = A234 & A233;
  assign \new_[58094]_  = \new_[58093]_  & \new_[58090]_ ;
  assign \new_[58095]_  = \new_[58094]_  & \new_[58087]_ ;
  assign \new_[58098]_  = ~A265 & A235;
  assign \new_[58101]_  = A298 & ~A266;
  assign \new_[58102]_  = \new_[58101]_  & \new_[58098]_ ;
  assign \new_[58105]_  = ~A300 & ~A299;
  assign \new_[58108]_  = A302 & ~A301;
  assign \new_[58109]_  = \new_[58108]_  & \new_[58105]_ ;
  assign \new_[58110]_  = \new_[58109]_  & \new_[58102]_ ;
  assign \new_[58113]_  = ~A169 & ~A170;
  assign \new_[58116]_  = A167 & ~A168;
  assign \new_[58117]_  = \new_[58116]_  & \new_[58113]_ ;
  assign \new_[58120]_  = ~A232 & ~A166;
  assign \new_[58123]_  = A234 & A233;
  assign \new_[58124]_  = \new_[58123]_  & \new_[58120]_ ;
  assign \new_[58125]_  = \new_[58124]_  & \new_[58117]_ ;
  assign \new_[58128]_  = ~A265 & A235;
  assign \new_[58131]_  = ~A298 & ~A266;
  assign \new_[58132]_  = \new_[58131]_  & \new_[58128]_ ;
  assign \new_[58135]_  = ~A300 & A299;
  assign \new_[58138]_  = A302 & ~A301;
  assign \new_[58139]_  = \new_[58138]_  & \new_[58135]_ ;
  assign \new_[58140]_  = \new_[58139]_  & \new_[58132]_ ;
  assign \new_[58143]_  = ~A169 & ~A170;
  assign \new_[58146]_  = A167 & ~A168;
  assign \new_[58147]_  = \new_[58146]_  & \new_[58143]_ ;
  assign \new_[58150]_  = ~A232 & ~A166;
  assign \new_[58153]_  = A234 & A233;
  assign \new_[58154]_  = \new_[58153]_  & \new_[58150]_ ;
  assign \new_[58155]_  = \new_[58154]_  & \new_[58147]_ ;
  assign \new_[58158]_  = A267 & ~A236;
  assign \new_[58161]_  = A269 & ~A268;
  assign \new_[58162]_  = \new_[58161]_  & \new_[58158]_ ;
  assign \new_[58165]_  = ~A299 & A298;
  assign \new_[58168]_  = A301 & A300;
  assign \new_[58169]_  = \new_[58168]_  & \new_[58165]_ ;
  assign \new_[58170]_  = \new_[58169]_  & \new_[58162]_ ;
  assign \new_[58173]_  = ~A169 & ~A170;
  assign \new_[58176]_  = A167 & ~A168;
  assign \new_[58177]_  = \new_[58176]_  & \new_[58173]_ ;
  assign \new_[58180]_  = ~A232 & ~A166;
  assign \new_[58183]_  = A234 & A233;
  assign \new_[58184]_  = \new_[58183]_  & \new_[58180]_ ;
  assign \new_[58185]_  = \new_[58184]_  & \new_[58177]_ ;
  assign \new_[58188]_  = A267 & ~A236;
  assign \new_[58191]_  = A269 & ~A268;
  assign \new_[58192]_  = \new_[58191]_  & \new_[58188]_ ;
  assign \new_[58195]_  = ~A299 & A298;
  assign \new_[58198]_  = ~A302 & A300;
  assign \new_[58199]_  = \new_[58198]_  & \new_[58195]_ ;
  assign \new_[58200]_  = \new_[58199]_  & \new_[58192]_ ;
  assign \new_[58203]_  = ~A169 & ~A170;
  assign \new_[58206]_  = A167 & ~A168;
  assign \new_[58207]_  = \new_[58206]_  & \new_[58203]_ ;
  assign \new_[58210]_  = ~A232 & ~A166;
  assign \new_[58213]_  = A234 & A233;
  assign \new_[58214]_  = \new_[58213]_  & \new_[58210]_ ;
  assign \new_[58215]_  = \new_[58214]_  & \new_[58207]_ ;
  assign \new_[58218]_  = A267 & ~A236;
  assign \new_[58221]_  = A269 & ~A268;
  assign \new_[58222]_  = \new_[58221]_  & \new_[58218]_ ;
  assign \new_[58225]_  = A299 & ~A298;
  assign \new_[58228]_  = A301 & A300;
  assign \new_[58229]_  = \new_[58228]_  & \new_[58225]_ ;
  assign \new_[58230]_  = \new_[58229]_  & \new_[58222]_ ;
  assign \new_[58233]_  = ~A169 & ~A170;
  assign \new_[58236]_  = A167 & ~A168;
  assign \new_[58237]_  = \new_[58236]_  & \new_[58233]_ ;
  assign \new_[58240]_  = ~A232 & ~A166;
  assign \new_[58243]_  = A234 & A233;
  assign \new_[58244]_  = \new_[58243]_  & \new_[58240]_ ;
  assign \new_[58245]_  = \new_[58244]_  & \new_[58237]_ ;
  assign \new_[58248]_  = A267 & ~A236;
  assign \new_[58251]_  = A269 & ~A268;
  assign \new_[58252]_  = \new_[58251]_  & \new_[58248]_ ;
  assign \new_[58255]_  = A299 & ~A298;
  assign \new_[58258]_  = ~A302 & A300;
  assign \new_[58259]_  = \new_[58258]_  & \new_[58255]_ ;
  assign \new_[58260]_  = \new_[58259]_  & \new_[58252]_ ;
  assign \new_[58263]_  = ~A169 & ~A170;
  assign \new_[58266]_  = A167 & ~A168;
  assign \new_[58267]_  = \new_[58266]_  & \new_[58263]_ ;
  assign \new_[58270]_  = ~A232 & ~A166;
  assign \new_[58273]_  = A234 & A233;
  assign \new_[58274]_  = \new_[58273]_  & \new_[58270]_ ;
  assign \new_[58275]_  = \new_[58274]_  & \new_[58267]_ ;
  assign \new_[58278]_  = ~A267 & ~A236;
  assign \new_[58281]_  = A298 & A268;
  assign \new_[58282]_  = \new_[58281]_  & \new_[58278]_ ;
  assign \new_[58285]_  = ~A300 & ~A299;
  assign \new_[58288]_  = A302 & ~A301;
  assign \new_[58289]_  = \new_[58288]_  & \new_[58285]_ ;
  assign \new_[58290]_  = \new_[58289]_  & \new_[58282]_ ;
  assign \new_[58293]_  = ~A169 & ~A170;
  assign \new_[58296]_  = A167 & ~A168;
  assign \new_[58297]_  = \new_[58296]_  & \new_[58293]_ ;
  assign \new_[58300]_  = ~A232 & ~A166;
  assign \new_[58303]_  = A234 & A233;
  assign \new_[58304]_  = \new_[58303]_  & \new_[58300]_ ;
  assign \new_[58305]_  = \new_[58304]_  & \new_[58297]_ ;
  assign \new_[58308]_  = ~A267 & ~A236;
  assign \new_[58311]_  = ~A298 & A268;
  assign \new_[58312]_  = \new_[58311]_  & \new_[58308]_ ;
  assign \new_[58315]_  = ~A300 & A299;
  assign \new_[58318]_  = A302 & ~A301;
  assign \new_[58319]_  = \new_[58318]_  & \new_[58315]_ ;
  assign \new_[58320]_  = \new_[58319]_  & \new_[58312]_ ;
  assign \new_[58323]_  = ~A169 & ~A170;
  assign \new_[58326]_  = A167 & ~A168;
  assign \new_[58327]_  = \new_[58326]_  & \new_[58323]_ ;
  assign \new_[58330]_  = ~A232 & ~A166;
  assign \new_[58333]_  = A234 & A233;
  assign \new_[58334]_  = \new_[58333]_  & \new_[58330]_ ;
  assign \new_[58335]_  = \new_[58334]_  & \new_[58327]_ ;
  assign \new_[58338]_  = ~A267 & ~A236;
  assign \new_[58341]_  = A298 & ~A269;
  assign \new_[58342]_  = \new_[58341]_  & \new_[58338]_ ;
  assign \new_[58345]_  = ~A300 & ~A299;
  assign \new_[58348]_  = A302 & ~A301;
  assign \new_[58349]_  = \new_[58348]_  & \new_[58345]_ ;
  assign \new_[58350]_  = \new_[58349]_  & \new_[58342]_ ;
  assign \new_[58353]_  = ~A169 & ~A170;
  assign \new_[58356]_  = A167 & ~A168;
  assign \new_[58357]_  = \new_[58356]_  & \new_[58353]_ ;
  assign \new_[58360]_  = ~A232 & ~A166;
  assign \new_[58363]_  = A234 & A233;
  assign \new_[58364]_  = \new_[58363]_  & \new_[58360]_ ;
  assign \new_[58365]_  = \new_[58364]_  & \new_[58357]_ ;
  assign \new_[58368]_  = ~A267 & ~A236;
  assign \new_[58371]_  = ~A298 & ~A269;
  assign \new_[58372]_  = \new_[58371]_  & \new_[58368]_ ;
  assign \new_[58375]_  = ~A300 & A299;
  assign \new_[58378]_  = A302 & ~A301;
  assign \new_[58379]_  = \new_[58378]_  & \new_[58375]_ ;
  assign \new_[58380]_  = \new_[58379]_  & \new_[58372]_ ;
  assign \new_[58383]_  = ~A169 & ~A170;
  assign \new_[58386]_  = A167 & ~A168;
  assign \new_[58387]_  = \new_[58386]_  & \new_[58383]_ ;
  assign \new_[58390]_  = ~A232 & ~A166;
  assign \new_[58393]_  = A234 & A233;
  assign \new_[58394]_  = \new_[58393]_  & \new_[58390]_ ;
  assign \new_[58395]_  = \new_[58394]_  & \new_[58387]_ ;
  assign \new_[58398]_  = A265 & ~A236;
  assign \new_[58401]_  = A298 & A266;
  assign \new_[58402]_  = \new_[58401]_  & \new_[58398]_ ;
  assign \new_[58405]_  = ~A300 & ~A299;
  assign \new_[58408]_  = A302 & ~A301;
  assign \new_[58409]_  = \new_[58408]_  & \new_[58405]_ ;
  assign \new_[58410]_  = \new_[58409]_  & \new_[58402]_ ;
  assign \new_[58413]_  = ~A169 & ~A170;
  assign \new_[58416]_  = A167 & ~A168;
  assign \new_[58417]_  = \new_[58416]_  & \new_[58413]_ ;
  assign \new_[58420]_  = ~A232 & ~A166;
  assign \new_[58423]_  = A234 & A233;
  assign \new_[58424]_  = \new_[58423]_  & \new_[58420]_ ;
  assign \new_[58425]_  = \new_[58424]_  & \new_[58417]_ ;
  assign \new_[58428]_  = A265 & ~A236;
  assign \new_[58431]_  = ~A298 & A266;
  assign \new_[58432]_  = \new_[58431]_  & \new_[58428]_ ;
  assign \new_[58435]_  = ~A300 & A299;
  assign \new_[58438]_  = A302 & ~A301;
  assign \new_[58439]_  = \new_[58438]_  & \new_[58435]_ ;
  assign \new_[58440]_  = \new_[58439]_  & \new_[58432]_ ;
  assign \new_[58443]_  = ~A169 & ~A170;
  assign \new_[58446]_  = A167 & ~A168;
  assign \new_[58447]_  = \new_[58446]_  & \new_[58443]_ ;
  assign \new_[58450]_  = ~A232 & ~A166;
  assign \new_[58453]_  = A234 & A233;
  assign \new_[58454]_  = \new_[58453]_  & \new_[58450]_ ;
  assign \new_[58455]_  = \new_[58454]_  & \new_[58447]_ ;
  assign \new_[58458]_  = ~A265 & ~A236;
  assign \new_[58461]_  = A298 & ~A266;
  assign \new_[58462]_  = \new_[58461]_  & \new_[58458]_ ;
  assign \new_[58465]_  = ~A300 & ~A299;
  assign \new_[58468]_  = A302 & ~A301;
  assign \new_[58469]_  = \new_[58468]_  & \new_[58465]_ ;
  assign \new_[58470]_  = \new_[58469]_  & \new_[58462]_ ;
  assign \new_[58473]_  = ~A169 & ~A170;
  assign \new_[58476]_  = A167 & ~A168;
  assign \new_[58477]_  = \new_[58476]_  & \new_[58473]_ ;
  assign \new_[58480]_  = ~A232 & ~A166;
  assign \new_[58483]_  = A234 & A233;
  assign \new_[58484]_  = \new_[58483]_  & \new_[58480]_ ;
  assign \new_[58485]_  = \new_[58484]_  & \new_[58477]_ ;
  assign \new_[58488]_  = ~A265 & ~A236;
  assign \new_[58491]_  = ~A298 & ~A266;
  assign \new_[58492]_  = \new_[58491]_  & \new_[58488]_ ;
  assign \new_[58495]_  = ~A300 & A299;
  assign \new_[58498]_  = A302 & ~A301;
  assign \new_[58499]_  = \new_[58498]_  & \new_[58495]_ ;
  assign \new_[58500]_  = \new_[58499]_  & \new_[58492]_ ;
  assign \new_[58503]_  = ~A169 & ~A170;
  assign \new_[58506]_  = A167 & ~A168;
  assign \new_[58507]_  = \new_[58506]_  & \new_[58503]_ ;
  assign \new_[58510]_  = ~A232 & ~A166;
  assign \new_[58513]_  = ~A234 & A233;
  assign \new_[58514]_  = \new_[58513]_  & \new_[58510]_ ;
  assign \new_[58515]_  = \new_[58514]_  & \new_[58507]_ ;
  assign \new_[58518]_  = A236 & ~A235;
  assign \new_[58521]_  = A268 & ~A267;
  assign \new_[58522]_  = \new_[58521]_  & \new_[58518]_ ;
  assign \new_[58525]_  = ~A299 & A298;
  assign \new_[58528]_  = A301 & A300;
  assign \new_[58529]_  = \new_[58528]_  & \new_[58525]_ ;
  assign \new_[58530]_  = \new_[58529]_  & \new_[58522]_ ;
  assign \new_[58533]_  = ~A169 & ~A170;
  assign \new_[58536]_  = A167 & ~A168;
  assign \new_[58537]_  = \new_[58536]_  & \new_[58533]_ ;
  assign \new_[58540]_  = ~A232 & ~A166;
  assign \new_[58543]_  = ~A234 & A233;
  assign \new_[58544]_  = \new_[58543]_  & \new_[58540]_ ;
  assign \new_[58545]_  = \new_[58544]_  & \new_[58537]_ ;
  assign \new_[58548]_  = A236 & ~A235;
  assign \new_[58551]_  = A268 & ~A267;
  assign \new_[58552]_  = \new_[58551]_  & \new_[58548]_ ;
  assign \new_[58555]_  = ~A299 & A298;
  assign \new_[58558]_  = ~A302 & A300;
  assign \new_[58559]_  = \new_[58558]_  & \new_[58555]_ ;
  assign \new_[58560]_  = \new_[58559]_  & \new_[58552]_ ;
  assign \new_[58563]_  = ~A169 & ~A170;
  assign \new_[58566]_  = A167 & ~A168;
  assign \new_[58567]_  = \new_[58566]_  & \new_[58563]_ ;
  assign \new_[58570]_  = ~A232 & ~A166;
  assign \new_[58573]_  = ~A234 & A233;
  assign \new_[58574]_  = \new_[58573]_  & \new_[58570]_ ;
  assign \new_[58575]_  = \new_[58574]_  & \new_[58567]_ ;
  assign \new_[58578]_  = A236 & ~A235;
  assign \new_[58581]_  = A268 & ~A267;
  assign \new_[58582]_  = \new_[58581]_  & \new_[58578]_ ;
  assign \new_[58585]_  = A299 & ~A298;
  assign \new_[58588]_  = A301 & A300;
  assign \new_[58589]_  = \new_[58588]_  & \new_[58585]_ ;
  assign \new_[58590]_  = \new_[58589]_  & \new_[58582]_ ;
  assign \new_[58593]_  = ~A169 & ~A170;
  assign \new_[58596]_  = A167 & ~A168;
  assign \new_[58597]_  = \new_[58596]_  & \new_[58593]_ ;
  assign \new_[58600]_  = ~A232 & ~A166;
  assign \new_[58603]_  = ~A234 & A233;
  assign \new_[58604]_  = \new_[58603]_  & \new_[58600]_ ;
  assign \new_[58605]_  = \new_[58604]_  & \new_[58597]_ ;
  assign \new_[58608]_  = A236 & ~A235;
  assign \new_[58611]_  = A268 & ~A267;
  assign \new_[58612]_  = \new_[58611]_  & \new_[58608]_ ;
  assign \new_[58615]_  = A299 & ~A298;
  assign \new_[58618]_  = ~A302 & A300;
  assign \new_[58619]_  = \new_[58618]_  & \new_[58615]_ ;
  assign \new_[58620]_  = \new_[58619]_  & \new_[58612]_ ;
  assign \new_[58623]_  = ~A169 & ~A170;
  assign \new_[58626]_  = A167 & ~A168;
  assign \new_[58627]_  = \new_[58626]_  & \new_[58623]_ ;
  assign \new_[58630]_  = ~A232 & ~A166;
  assign \new_[58633]_  = ~A234 & A233;
  assign \new_[58634]_  = \new_[58633]_  & \new_[58630]_ ;
  assign \new_[58635]_  = \new_[58634]_  & \new_[58627]_ ;
  assign \new_[58638]_  = A236 & ~A235;
  assign \new_[58641]_  = ~A269 & ~A267;
  assign \new_[58642]_  = \new_[58641]_  & \new_[58638]_ ;
  assign \new_[58645]_  = ~A299 & A298;
  assign \new_[58648]_  = A301 & A300;
  assign \new_[58649]_  = \new_[58648]_  & \new_[58645]_ ;
  assign \new_[58650]_  = \new_[58649]_  & \new_[58642]_ ;
  assign \new_[58653]_  = ~A169 & ~A170;
  assign \new_[58656]_  = A167 & ~A168;
  assign \new_[58657]_  = \new_[58656]_  & \new_[58653]_ ;
  assign \new_[58660]_  = ~A232 & ~A166;
  assign \new_[58663]_  = ~A234 & A233;
  assign \new_[58664]_  = \new_[58663]_  & \new_[58660]_ ;
  assign \new_[58665]_  = \new_[58664]_  & \new_[58657]_ ;
  assign \new_[58668]_  = A236 & ~A235;
  assign \new_[58671]_  = ~A269 & ~A267;
  assign \new_[58672]_  = \new_[58671]_  & \new_[58668]_ ;
  assign \new_[58675]_  = ~A299 & A298;
  assign \new_[58678]_  = ~A302 & A300;
  assign \new_[58679]_  = \new_[58678]_  & \new_[58675]_ ;
  assign \new_[58680]_  = \new_[58679]_  & \new_[58672]_ ;
  assign \new_[58683]_  = ~A169 & ~A170;
  assign \new_[58686]_  = A167 & ~A168;
  assign \new_[58687]_  = \new_[58686]_  & \new_[58683]_ ;
  assign \new_[58690]_  = ~A232 & ~A166;
  assign \new_[58693]_  = ~A234 & A233;
  assign \new_[58694]_  = \new_[58693]_  & \new_[58690]_ ;
  assign \new_[58695]_  = \new_[58694]_  & \new_[58687]_ ;
  assign \new_[58698]_  = A236 & ~A235;
  assign \new_[58701]_  = ~A269 & ~A267;
  assign \new_[58702]_  = \new_[58701]_  & \new_[58698]_ ;
  assign \new_[58705]_  = A299 & ~A298;
  assign \new_[58708]_  = A301 & A300;
  assign \new_[58709]_  = \new_[58708]_  & \new_[58705]_ ;
  assign \new_[58710]_  = \new_[58709]_  & \new_[58702]_ ;
  assign \new_[58713]_  = ~A169 & ~A170;
  assign \new_[58716]_  = A167 & ~A168;
  assign \new_[58717]_  = \new_[58716]_  & \new_[58713]_ ;
  assign \new_[58720]_  = ~A232 & ~A166;
  assign \new_[58723]_  = ~A234 & A233;
  assign \new_[58724]_  = \new_[58723]_  & \new_[58720]_ ;
  assign \new_[58725]_  = \new_[58724]_  & \new_[58717]_ ;
  assign \new_[58728]_  = A236 & ~A235;
  assign \new_[58731]_  = ~A269 & ~A267;
  assign \new_[58732]_  = \new_[58731]_  & \new_[58728]_ ;
  assign \new_[58735]_  = A299 & ~A298;
  assign \new_[58738]_  = ~A302 & A300;
  assign \new_[58739]_  = \new_[58738]_  & \new_[58735]_ ;
  assign \new_[58740]_  = \new_[58739]_  & \new_[58732]_ ;
  assign \new_[58743]_  = ~A169 & ~A170;
  assign \new_[58746]_  = A167 & ~A168;
  assign \new_[58747]_  = \new_[58746]_  & \new_[58743]_ ;
  assign \new_[58750]_  = ~A232 & ~A166;
  assign \new_[58753]_  = ~A234 & A233;
  assign \new_[58754]_  = \new_[58753]_  & \new_[58750]_ ;
  assign \new_[58755]_  = \new_[58754]_  & \new_[58747]_ ;
  assign \new_[58758]_  = A236 & ~A235;
  assign \new_[58761]_  = A266 & A265;
  assign \new_[58762]_  = \new_[58761]_  & \new_[58758]_ ;
  assign \new_[58765]_  = ~A299 & A298;
  assign \new_[58768]_  = A301 & A300;
  assign \new_[58769]_  = \new_[58768]_  & \new_[58765]_ ;
  assign \new_[58770]_  = \new_[58769]_  & \new_[58762]_ ;
  assign \new_[58773]_  = ~A169 & ~A170;
  assign \new_[58776]_  = A167 & ~A168;
  assign \new_[58777]_  = \new_[58776]_  & \new_[58773]_ ;
  assign \new_[58780]_  = ~A232 & ~A166;
  assign \new_[58783]_  = ~A234 & A233;
  assign \new_[58784]_  = \new_[58783]_  & \new_[58780]_ ;
  assign \new_[58785]_  = \new_[58784]_  & \new_[58777]_ ;
  assign \new_[58788]_  = A236 & ~A235;
  assign \new_[58791]_  = A266 & A265;
  assign \new_[58792]_  = \new_[58791]_  & \new_[58788]_ ;
  assign \new_[58795]_  = ~A299 & A298;
  assign \new_[58798]_  = ~A302 & A300;
  assign \new_[58799]_  = \new_[58798]_  & \new_[58795]_ ;
  assign \new_[58800]_  = \new_[58799]_  & \new_[58792]_ ;
  assign \new_[58803]_  = ~A169 & ~A170;
  assign \new_[58806]_  = A167 & ~A168;
  assign \new_[58807]_  = \new_[58806]_  & \new_[58803]_ ;
  assign \new_[58810]_  = ~A232 & ~A166;
  assign \new_[58813]_  = ~A234 & A233;
  assign \new_[58814]_  = \new_[58813]_  & \new_[58810]_ ;
  assign \new_[58815]_  = \new_[58814]_  & \new_[58807]_ ;
  assign \new_[58818]_  = A236 & ~A235;
  assign \new_[58821]_  = A266 & A265;
  assign \new_[58822]_  = \new_[58821]_  & \new_[58818]_ ;
  assign \new_[58825]_  = A299 & ~A298;
  assign \new_[58828]_  = A301 & A300;
  assign \new_[58829]_  = \new_[58828]_  & \new_[58825]_ ;
  assign \new_[58830]_  = \new_[58829]_  & \new_[58822]_ ;
  assign \new_[58833]_  = ~A169 & ~A170;
  assign \new_[58836]_  = A167 & ~A168;
  assign \new_[58837]_  = \new_[58836]_  & \new_[58833]_ ;
  assign \new_[58840]_  = ~A232 & ~A166;
  assign \new_[58843]_  = ~A234 & A233;
  assign \new_[58844]_  = \new_[58843]_  & \new_[58840]_ ;
  assign \new_[58845]_  = \new_[58844]_  & \new_[58837]_ ;
  assign \new_[58848]_  = A236 & ~A235;
  assign \new_[58851]_  = A266 & A265;
  assign \new_[58852]_  = \new_[58851]_  & \new_[58848]_ ;
  assign \new_[58855]_  = A299 & ~A298;
  assign \new_[58858]_  = ~A302 & A300;
  assign \new_[58859]_  = \new_[58858]_  & \new_[58855]_ ;
  assign \new_[58860]_  = \new_[58859]_  & \new_[58852]_ ;
  assign \new_[58863]_  = ~A169 & ~A170;
  assign \new_[58866]_  = A167 & ~A168;
  assign \new_[58867]_  = \new_[58866]_  & \new_[58863]_ ;
  assign \new_[58870]_  = ~A232 & ~A166;
  assign \new_[58873]_  = ~A234 & A233;
  assign \new_[58874]_  = \new_[58873]_  & \new_[58870]_ ;
  assign \new_[58875]_  = \new_[58874]_  & \new_[58867]_ ;
  assign \new_[58878]_  = A236 & ~A235;
  assign \new_[58881]_  = ~A266 & ~A265;
  assign \new_[58882]_  = \new_[58881]_  & \new_[58878]_ ;
  assign \new_[58885]_  = ~A299 & A298;
  assign \new_[58888]_  = A301 & A300;
  assign \new_[58889]_  = \new_[58888]_  & \new_[58885]_ ;
  assign \new_[58890]_  = \new_[58889]_  & \new_[58882]_ ;
  assign \new_[58893]_  = ~A169 & ~A170;
  assign \new_[58896]_  = A167 & ~A168;
  assign \new_[58897]_  = \new_[58896]_  & \new_[58893]_ ;
  assign \new_[58900]_  = ~A232 & ~A166;
  assign \new_[58903]_  = ~A234 & A233;
  assign \new_[58904]_  = \new_[58903]_  & \new_[58900]_ ;
  assign \new_[58905]_  = \new_[58904]_  & \new_[58897]_ ;
  assign \new_[58908]_  = A236 & ~A235;
  assign \new_[58911]_  = ~A266 & ~A265;
  assign \new_[58912]_  = \new_[58911]_  & \new_[58908]_ ;
  assign \new_[58915]_  = ~A299 & A298;
  assign \new_[58918]_  = ~A302 & A300;
  assign \new_[58919]_  = \new_[58918]_  & \new_[58915]_ ;
  assign \new_[58920]_  = \new_[58919]_  & \new_[58912]_ ;
  assign \new_[58923]_  = ~A169 & ~A170;
  assign \new_[58926]_  = A167 & ~A168;
  assign \new_[58927]_  = \new_[58926]_  & \new_[58923]_ ;
  assign \new_[58930]_  = ~A232 & ~A166;
  assign \new_[58933]_  = ~A234 & A233;
  assign \new_[58934]_  = \new_[58933]_  & \new_[58930]_ ;
  assign \new_[58935]_  = \new_[58934]_  & \new_[58927]_ ;
  assign \new_[58938]_  = A236 & ~A235;
  assign \new_[58941]_  = ~A266 & ~A265;
  assign \new_[58942]_  = \new_[58941]_  & \new_[58938]_ ;
  assign \new_[58945]_  = A299 & ~A298;
  assign \new_[58948]_  = A301 & A300;
  assign \new_[58949]_  = \new_[58948]_  & \new_[58945]_ ;
  assign \new_[58950]_  = \new_[58949]_  & \new_[58942]_ ;
  assign \new_[58953]_  = ~A169 & ~A170;
  assign \new_[58956]_  = A167 & ~A168;
  assign \new_[58957]_  = \new_[58956]_  & \new_[58953]_ ;
  assign \new_[58960]_  = ~A232 & ~A166;
  assign \new_[58963]_  = ~A234 & A233;
  assign \new_[58964]_  = \new_[58963]_  & \new_[58960]_ ;
  assign \new_[58965]_  = \new_[58964]_  & \new_[58957]_ ;
  assign \new_[58968]_  = A236 & ~A235;
  assign \new_[58971]_  = ~A266 & ~A265;
  assign \new_[58972]_  = \new_[58971]_  & \new_[58968]_ ;
  assign \new_[58975]_  = A299 & ~A298;
  assign \new_[58978]_  = ~A302 & A300;
  assign \new_[58979]_  = \new_[58978]_  & \new_[58975]_ ;
  assign \new_[58980]_  = \new_[58979]_  & \new_[58972]_ ;
  assign \new_[58983]_  = ~A169 & ~A170;
  assign \new_[58986]_  = A167 & ~A168;
  assign \new_[58987]_  = \new_[58986]_  & \new_[58983]_ ;
  assign \new_[58990]_  = A232 & ~A166;
  assign \new_[58993]_  = A234 & ~A233;
  assign \new_[58994]_  = \new_[58993]_  & \new_[58990]_ ;
  assign \new_[58995]_  = \new_[58994]_  & \new_[58987]_ ;
  assign \new_[58998]_  = A267 & A235;
  assign \new_[59001]_  = A269 & ~A268;
  assign \new_[59002]_  = \new_[59001]_  & \new_[58998]_ ;
  assign \new_[59005]_  = ~A299 & A298;
  assign \new_[59008]_  = A301 & A300;
  assign \new_[59009]_  = \new_[59008]_  & \new_[59005]_ ;
  assign \new_[59010]_  = \new_[59009]_  & \new_[59002]_ ;
  assign \new_[59013]_  = ~A169 & ~A170;
  assign \new_[59016]_  = A167 & ~A168;
  assign \new_[59017]_  = \new_[59016]_  & \new_[59013]_ ;
  assign \new_[59020]_  = A232 & ~A166;
  assign \new_[59023]_  = A234 & ~A233;
  assign \new_[59024]_  = \new_[59023]_  & \new_[59020]_ ;
  assign \new_[59025]_  = \new_[59024]_  & \new_[59017]_ ;
  assign \new_[59028]_  = A267 & A235;
  assign \new_[59031]_  = A269 & ~A268;
  assign \new_[59032]_  = \new_[59031]_  & \new_[59028]_ ;
  assign \new_[59035]_  = ~A299 & A298;
  assign \new_[59038]_  = ~A302 & A300;
  assign \new_[59039]_  = \new_[59038]_  & \new_[59035]_ ;
  assign \new_[59040]_  = \new_[59039]_  & \new_[59032]_ ;
  assign \new_[59043]_  = ~A169 & ~A170;
  assign \new_[59046]_  = A167 & ~A168;
  assign \new_[59047]_  = \new_[59046]_  & \new_[59043]_ ;
  assign \new_[59050]_  = A232 & ~A166;
  assign \new_[59053]_  = A234 & ~A233;
  assign \new_[59054]_  = \new_[59053]_  & \new_[59050]_ ;
  assign \new_[59055]_  = \new_[59054]_  & \new_[59047]_ ;
  assign \new_[59058]_  = A267 & A235;
  assign \new_[59061]_  = A269 & ~A268;
  assign \new_[59062]_  = \new_[59061]_  & \new_[59058]_ ;
  assign \new_[59065]_  = A299 & ~A298;
  assign \new_[59068]_  = A301 & A300;
  assign \new_[59069]_  = \new_[59068]_  & \new_[59065]_ ;
  assign \new_[59070]_  = \new_[59069]_  & \new_[59062]_ ;
  assign \new_[59073]_  = ~A169 & ~A170;
  assign \new_[59076]_  = A167 & ~A168;
  assign \new_[59077]_  = \new_[59076]_  & \new_[59073]_ ;
  assign \new_[59080]_  = A232 & ~A166;
  assign \new_[59083]_  = A234 & ~A233;
  assign \new_[59084]_  = \new_[59083]_  & \new_[59080]_ ;
  assign \new_[59085]_  = \new_[59084]_  & \new_[59077]_ ;
  assign \new_[59088]_  = A267 & A235;
  assign \new_[59091]_  = A269 & ~A268;
  assign \new_[59092]_  = \new_[59091]_  & \new_[59088]_ ;
  assign \new_[59095]_  = A299 & ~A298;
  assign \new_[59098]_  = ~A302 & A300;
  assign \new_[59099]_  = \new_[59098]_  & \new_[59095]_ ;
  assign \new_[59100]_  = \new_[59099]_  & \new_[59092]_ ;
  assign \new_[59103]_  = ~A169 & ~A170;
  assign \new_[59106]_  = A167 & ~A168;
  assign \new_[59107]_  = \new_[59106]_  & \new_[59103]_ ;
  assign \new_[59110]_  = A232 & ~A166;
  assign \new_[59113]_  = A234 & ~A233;
  assign \new_[59114]_  = \new_[59113]_  & \new_[59110]_ ;
  assign \new_[59115]_  = \new_[59114]_  & \new_[59107]_ ;
  assign \new_[59118]_  = ~A267 & A235;
  assign \new_[59121]_  = A298 & A268;
  assign \new_[59122]_  = \new_[59121]_  & \new_[59118]_ ;
  assign \new_[59125]_  = ~A300 & ~A299;
  assign \new_[59128]_  = A302 & ~A301;
  assign \new_[59129]_  = \new_[59128]_  & \new_[59125]_ ;
  assign \new_[59130]_  = \new_[59129]_  & \new_[59122]_ ;
  assign \new_[59133]_  = ~A169 & ~A170;
  assign \new_[59136]_  = A167 & ~A168;
  assign \new_[59137]_  = \new_[59136]_  & \new_[59133]_ ;
  assign \new_[59140]_  = A232 & ~A166;
  assign \new_[59143]_  = A234 & ~A233;
  assign \new_[59144]_  = \new_[59143]_  & \new_[59140]_ ;
  assign \new_[59145]_  = \new_[59144]_  & \new_[59137]_ ;
  assign \new_[59148]_  = ~A267 & A235;
  assign \new_[59151]_  = ~A298 & A268;
  assign \new_[59152]_  = \new_[59151]_  & \new_[59148]_ ;
  assign \new_[59155]_  = ~A300 & A299;
  assign \new_[59158]_  = A302 & ~A301;
  assign \new_[59159]_  = \new_[59158]_  & \new_[59155]_ ;
  assign \new_[59160]_  = \new_[59159]_  & \new_[59152]_ ;
  assign \new_[59163]_  = ~A169 & ~A170;
  assign \new_[59166]_  = A167 & ~A168;
  assign \new_[59167]_  = \new_[59166]_  & \new_[59163]_ ;
  assign \new_[59170]_  = A232 & ~A166;
  assign \new_[59173]_  = A234 & ~A233;
  assign \new_[59174]_  = \new_[59173]_  & \new_[59170]_ ;
  assign \new_[59175]_  = \new_[59174]_  & \new_[59167]_ ;
  assign \new_[59178]_  = ~A267 & A235;
  assign \new_[59181]_  = A298 & ~A269;
  assign \new_[59182]_  = \new_[59181]_  & \new_[59178]_ ;
  assign \new_[59185]_  = ~A300 & ~A299;
  assign \new_[59188]_  = A302 & ~A301;
  assign \new_[59189]_  = \new_[59188]_  & \new_[59185]_ ;
  assign \new_[59190]_  = \new_[59189]_  & \new_[59182]_ ;
  assign \new_[59193]_  = ~A169 & ~A170;
  assign \new_[59196]_  = A167 & ~A168;
  assign \new_[59197]_  = \new_[59196]_  & \new_[59193]_ ;
  assign \new_[59200]_  = A232 & ~A166;
  assign \new_[59203]_  = A234 & ~A233;
  assign \new_[59204]_  = \new_[59203]_  & \new_[59200]_ ;
  assign \new_[59205]_  = \new_[59204]_  & \new_[59197]_ ;
  assign \new_[59208]_  = ~A267 & A235;
  assign \new_[59211]_  = ~A298 & ~A269;
  assign \new_[59212]_  = \new_[59211]_  & \new_[59208]_ ;
  assign \new_[59215]_  = ~A300 & A299;
  assign \new_[59218]_  = A302 & ~A301;
  assign \new_[59219]_  = \new_[59218]_  & \new_[59215]_ ;
  assign \new_[59220]_  = \new_[59219]_  & \new_[59212]_ ;
  assign \new_[59223]_  = ~A169 & ~A170;
  assign \new_[59226]_  = A167 & ~A168;
  assign \new_[59227]_  = \new_[59226]_  & \new_[59223]_ ;
  assign \new_[59230]_  = A232 & ~A166;
  assign \new_[59233]_  = A234 & ~A233;
  assign \new_[59234]_  = \new_[59233]_  & \new_[59230]_ ;
  assign \new_[59235]_  = \new_[59234]_  & \new_[59227]_ ;
  assign \new_[59238]_  = A265 & A235;
  assign \new_[59241]_  = A298 & A266;
  assign \new_[59242]_  = \new_[59241]_  & \new_[59238]_ ;
  assign \new_[59245]_  = ~A300 & ~A299;
  assign \new_[59248]_  = A302 & ~A301;
  assign \new_[59249]_  = \new_[59248]_  & \new_[59245]_ ;
  assign \new_[59250]_  = \new_[59249]_  & \new_[59242]_ ;
  assign \new_[59253]_  = ~A169 & ~A170;
  assign \new_[59256]_  = A167 & ~A168;
  assign \new_[59257]_  = \new_[59256]_  & \new_[59253]_ ;
  assign \new_[59260]_  = A232 & ~A166;
  assign \new_[59263]_  = A234 & ~A233;
  assign \new_[59264]_  = \new_[59263]_  & \new_[59260]_ ;
  assign \new_[59265]_  = \new_[59264]_  & \new_[59257]_ ;
  assign \new_[59268]_  = A265 & A235;
  assign \new_[59271]_  = ~A298 & A266;
  assign \new_[59272]_  = \new_[59271]_  & \new_[59268]_ ;
  assign \new_[59275]_  = ~A300 & A299;
  assign \new_[59278]_  = A302 & ~A301;
  assign \new_[59279]_  = \new_[59278]_  & \new_[59275]_ ;
  assign \new_[59280]_  = \new_[59279]_  & \new_[59272]_ ;
  assign \new_[59283]_  = ~A169 & ~A170;
  assign \new_[59286]_  = A167 & ~A168;
  assign \new_[59287]_  = \new_[59286]_  & \new_[59283]_ ;
  assign \new_[59290]_  = A232 & ~A166;
  assign \new_[59293]_  = A234 & ~A233;
  assign \new_[59294]_  = \new_[59293]_  & \new_[59290]_ ;
  assign \new_[59295]_  = \new_[59294]_  & \new_[59287]_ ;
  assign \new_[59298]_  = ~A265 & A235;
  assign \new_[59301]_  = A298 & ~A266;
  assign \new_[59302]_  = \new_[59301]_  & \new_[59298]_ ;
  assign \new_[59305]_  = ~A300 & ~A299;
  assign \new_[59308]_  = A302 & ~A301;
  assign \new_[59309]_  = \new_[59308]_  & \new_[59305]_ ;
  assign \new_[59310]_  = \new_[59309]_  & \new_[59302]_ ;
  assign \new_[59313]_  = ~A169 & ~A170;
  assign \new_[59316]_  = A167 & ~A168;
  assign \new_[59317]_  = \new_[59316]_  & \new_[59313]_ ;
  assign \new_[59320]_  = A232 & ~A166;
  assign \new_[59323]_  = A234 & ~A233;
  assign \new_[59324]_  = \new_[59323]_  & \new_[59320]_ ;
  assign \new_[59325]_  = \new_[59324]_  & \new_[59317]_ ;
  assign \new_[59328]_  = ~A265 & A235;
  assign \new_[59331]_  = ~A298 & ~A266;
  assign \new_[59332]_  = \new_[59331]_  & \new_[59328]_ ;
  assign \new_[59335]_  = ~A300 & A299;
  assign \new_[59338]_  = A302 & ~A301;
  assign \new_[59339]_  = \new_[59338]_  & \new_[59335]_ ;
  assign \new_[59340]_  = \new_[59339]_  & \new_[59332]_ ;
  assign \new_[59343]_  = ~A169 & ~A170;
  assign \new_[59346]_  = A167 & ~A168;
  assign \new_[59347]_  = \new_[59346]_  & \new_[59343]_ ;
  assign \new_[59350]_  = A232 & ~A166;
  assign \new_[59353]_  = A234 & ~A233;
  assign \new_[59354]_  = \new_[59353]_  & \new_[59350]_ ;
  assign \new_[59355]_  = \new_[59354]_  & \new_[59347]_ ;
  assign \new_[59358]_  = A267 & ~A236;
  assign \new_[59361]_  = A269 & ~A268;
  assign \new_[59362]_  = \new_[59361]_  & \new_[59358]_ ;
  assign \new_[59365]_  = ~A299 & A298;
  assign \new_[59368]_  = A301 & A300;
  assign \new_[59369]_  = \new_[59368]_  & \new_[59365]_ ;
  assign \new_[59370]_  = \new_[59369]_  & \new_[59362]_ ;
  assign \new_[59373]_  = ~A169 & ~A170;
  assign \new_[59376]_  = A167 & ~A168;
  assign \new_[59377]_  = \new_[59376]_  & \new_[59373]_ ;
  assign \new_[59380]_  = A232 & ~A166;
  assign \new_[59383]_  = A234 & ~A233;
  assign \new_[59384]_  = \new_[59383]_  & \new_[59380]_ ;
  assign \new_[59385]_  = \new_[59384]_  & \new_[59377]_ ;
  assign \new_[59388]_  = A267 & ~A236;
  assign \new_[59391]_  = A269 & ~A268;
  assign \new_[59392]_  = \new_[59391]_  & \new_[59388]_ ;
  assign \new_[59395]_  = ~A299 & A298;
  assign \new_[59398]_  = ~A302 & A300;
  assign \new_[59399]_  = \new_[59398]_  & \new_[59395]_ ;
  assign \new_[59400]_  = \new_[59399]_  & \new_[59392]_ ;
  assign \new_[59403]_  = ~A169 & ~A170;
  assign \new_[59406]_  = A167 & ~A168;
  assign \new_[59407]_  = \new_[59406]_  & \new_[59403]_ ;
  assign \new_[59410]_  = A232 & ~A166;
  assign \new_[59413]_  = A234 & ~A233;
  assign \new_[59414]_  = \new_[59413]_  & \new_[59410]_ ;
  assign \new_[59415]_  = \new_[59414]_  & \new_[59407]_ ;
  assign \new_[59418]_  = A267 & ~A236;
  assign \new_[59421]_  = A269 & ~A268;
  assign \new_[59422]_  = \new_[59421]_  & \new_[59418]_ ;
  assign \new_[59425]_  = A299 & ~A298;
  assign \new_[59428]_  = A301 & A300;
  assign \new_[59429]_  = \new_[59428]_  & \new_[59425]_ ;
  assign \new_[59430]_  = \new_[59429]_  & \new_[59422]_ ;
  assign \new_[59433]_  = ~A169 & ~A170;
  assign \new_[59436]_  = A167 & ~A168;
  assign \new_[59437]_  = \new_[59436]_  & \new_[59433]_ ;
  assign \new_[59440]_  = A232 & ~A166;
  assign \new_[59443]_  = A234 & ~A233;
  assign \new_[59444]_  = \new_[59443]_  & \new_[59440]_ ;
  assign \new_[59445]_  = \new_[59444]_  & \new_[59437]_ ;
  assign \new_[59448]_  = A267 & ~A236;
  assign \new_[59451]_  = A269 & ~A268;
  assign \new_[59452]_  = \new_[59451]_  & \new_[59448]_ ;
  assign \new_[59455]_  = A299 & ~A298;
  assign \new_[59458]_  = ~A302 & A300;
  assign \new_[59459]_  = \new_[59458]_  & \new_[59455]_ ;
  assign \new_[59460]_  = \new_[59459]_  & \new_[59452]_ ;
  assign \new_[59463]_  = ~A169 & ~A170;
  assign \new_[59466]_  = A167 & ~A168;
  assign \new_[59467]_  = \new_[59466]_  & \new_[59463]_ ;
  assign \new_[59470]_  = A232 & ~A166;
  assign \new_[59473]_  = A234 & ~A233;
  assign \new_[59474]_  = \new_[59473]_  & \new_[59470]_ ;
  assign \new_[59475]_  = \new_[59474]_  & \new_[59467]_ ;
  assign \new_[59478]_  = ~A267 & ~A236;
  assign \new_[59481]_  = A298 & A268;
  assign \new_[59482]_  = \new_[59481]_  & \new_[59478]_ ;
  assign \new_[59485]_  = ~A300 & ~A299;
  assign \new_[59488]_  = A302 & ~A301;
  assign \new_[59489]_  = \new_[59488]_  & \new_[59485]_ ;
  assign \new_[59490]_  = \new_[59489]_  & \new_[59482]_ ;
  assign \new_[59493]_  = ~A169 & ~A170;
  assign \new_[59496]_  = A167 & ~A168;
  assign \new_[59497]_  = \new_[59496]_  & \new_[59493]_ ;
  assign \new_[59500]_  = A232 & ~A166;
  assign \new_[59503]_  = A234 & ~A233;
  assign \new_[59504]_  = \new_[59503]_  & \new_[59500]_ ;
  assign \new_[59505]_  = \new_[59504]_  & \new_[59497]_ ;
  assign \new_[59508]_  = ~A267 & ~A236;
  assign \new_[59511]_  = ~A298 & A268;
  assign \new_[59512]_  = \new_[59511]_  & \new_[59508]_ ;
  assign \new_[59515]_  = ~A300 & A299;
  assign \new_[59518]_  = A302 & ~A301;
  assign \new_[59519]_  = \new_[59518]_  & \new_[59515]_ ;
  assign \new_[59520]_  = \new_[59519]_  & \new_[59512]_ ;
  assign \new_[59523]_  = ~A169 & ~A170;
  assign \new_[59526]_  = A167 & ~A168;
  assign \new_[59527]_  = \new_[59526]_  & \new_[59523]_ ;
  assign \new_[59530]_  = A232 & ~A166;
  assign \new_[59533]_  = A234 & ~A233;
  assign \new_[59534]_  = \new_[59533]_  & \new_[59530]_ ;
  assign \new_[59535]_  = \new_[59534]_  & \new_[59527]_ ;
  assign \new_[59538]_  = ~A267 & ~A236;
  assign \new_[59541]_  = A298 & ~A269;
  assign \new_[59542]_  = \new_[59541]_  & \new_[59538]_ ;
  assign \new_[59545]_  = ~A300 & ~A299;
  assign \new_[59548]_  = A302 & ~A301;
  assign \new_[59549]_  = \new_[59548]_  & \new_[59545]_ ;
  assign \new_[59550]_  = \new_[59549]_  & \new_[59542]_ ;
  assign \new_[59553]_  = ~A169 & ~A170;
  assign \new_[59556]_  = A167 & ~A168;
  assign \new_[59557]_  = \new_[59556]_  & \new_[59553]_ ;
  assign \new_[59560]_  = A232 & ~A166;
  assign \new_[59563]_  = A234 & ~A233;
  assign \new_[59564]_  = \new_[59563]_  & \new_[59560]_ ;
  assign \new_[59565]_  = \new_[59564]_  & \new_[59557]_ ;
  assign \new_[59568]_  = ~A267 & ~A236;
  assign \new_[59571]_  = ~A298 & ~A269;
  assign \new_[59572]_  = \new_[59571]_  & \new_[59568]_ ;
  assign \new_[59575]_  = ~A300 & A299;
  assign \new_[59578]_  = A302 & ~A301;
  assign \new_[59579]_  = \new_[59578]_  & \new_[59575]_ ;
  assign \new_[59580]_  = \new_[59579]_  & \new_[59572]_ ;
  assign \new_[59583]_  = ~A169 & ~A170;
  assign \new_[59586]_  = A167 & ~A168;
  assign \new_[59587]_  = \new_[59586]_  & \new_[59583]_ ;
  assign \new_[59590]_  = A232 & ~A166;
  assign \new_[59593]_  = A234 & ~A233;
  assign \new_[59594]_  = \new_[59593]_  & \new_[59590]_ ;
  assign \new_[59595]_  = \new_[59594]_  & \new_[59587]_ ;
  assign \new_[59598]_  = A265 & ~A236;
  assign \new_[59601]_  = A298 & A266;
  assign \new_[59602]_  = \new_[59601]_  & \new_[59598]_ ;
  assign \new_[59605]_  = ~A300 & ~A299;
  assign \new_[59608]_  = A302 & ~A301;
  assign \new_[59609]_  = \new_[59608]_  & \new_[59605]_ ;
  assign \new_[59610]_  = \new_[59609]_  & \new_[59602]_ ;
  assign \new_[59613]_  = ~A169 & ~A170;
  assign \new_[59616]_  = A167 & ~A168;
  assign \new_[59617]_  = \new_[59616]_  & \new_[59613]_ ;
  assign \new_[59620]_  = A232 & ~A166;
  assign \new_[59623]_  = A234 & ~A233;
  assign \new_[59624]_  = \new_[59623]_  & \new_[59620]_ ;
  assign \new_[59625]_  = \new_[59624]_  & \new_[59617]_ ;
  assign \new_[59628]_  = A265 & ~A236;
  assign \new_[59631]_  = ~A298 & A266;
  assign \new_[59632]_  = \new_[59631]_  & \new_[59628]_ ;
  assign \new_[59635]_  = ~A300 & A299;
  assign \new_[59638]_  = A302 & ~A301;
  assign \new_[59639]_  = \new_[59638]_  & \new_[59635]_ ;
  assign \new_[59640]_  = \new_[59639]_  & \new_[59632]_ ;
  assign \new_[59643]_  = ~A169 & ~A170;
  assign \new_[59646]_  = A167 & ~A168;
  assign \new_[59647]_  = \new_[59646]_  & \new_[59643]_ ;
  assign \new_[59650]_  = A232 & ~A166;
  assign \new_[59653]_  = A234 & ~A233;
  assign \new_[59654]_  = \new_[59653]_  & \new_[59650]_ ;
  assign \new_[59655]_  = \new_[59654]_  & \new_[59647]_ ;
  assign \new_[59658]_  = ~A265 & ~A236;
  assign \new_[59661]_  = A298 & ~A266;
  assign \new_[59662]_  = \new_[59661]_  & \new_[59658]_ ;
  assign \new_[59665]_  = ~A300 & ~A299;
  assign \new_[59668]_  = A302 & ~A301;
  assign \new_[59669]_  = \new_[59668]_  & \new_[59665]_ ;
  assign \new_[59670]_  = \new_[59669]_  & \new_[59662]_ ;
  assign \new_[59673]_  = ~A169 & ~A170;
  assign \new_[59676]_  = A167 & ~A168;
  assign \new_[59677]_  = \new_[59676]_  & \new_[59673]_ ;
  assign \new_[59680]_  = A232 & ~A166;
  assign \new_[59683]_  = A234 & ~A233;
  assign \new_[59684]_  = \new_[59683]_  & \new_[59680]_ ;
  assign \new_[59685]_  = \new_[59684]_  & \new_[59677]_ ;
  assign \new_[59688]_  = ~A265 & ~A236;
  assign \new_[59691]_  = ~A298 & ~A266;
  assign \new_[59692]_  = \new_[59691]_  & \new_[59688]_ ;
  assign \new_[59695]_  = ~A300 & A299;
  assign \new_[59698]_  = A302 & ~A301;
  assign \new_[59699]_  = \new_[59698]_  & \new_[59695]_ ;
  assign \new_[59700]_  = \new_[59699]_  & \new_[59692]_ ;
  assign \new_[59703]_  = ~A169 & ~A170;
  assign \new_[59706]_  = A167 & ~A168;
  assign \new_[59707]_  = \new_[59706]_  & \new_[59703]_ ;
  assign \new_[59710]_  = A232 & ~A166;
  assign \new_[59713]_  = ~A234 & ~A233;
  assign \new_[59714]_  = \new_[59713]_  & \new_[59710]_ ;
  assign \new_[59715]_  = \new_[59714]_  & \new_[59707]_ ;
  assign \new_[59718]_  = A236 & ~A235;
  assign \new_[59721]_  = A268 & ~A267;
  assign \new_[59722]_  = \new_[59721]_  & \new_[59718]_ ;
  assign \new_[59725]_  = ~A299 & A298;
  assign \new_[59728]_  = A301 & A300;
  assign \new_[59729]_  = \new_[59728]_  & \new_[59725]_ ;
  assign \new_[59730]_  = \new_[59729]_  & \new_[59722]_ ;
  assign \new_[59733]_  = ~A169 & ~A170;
  assign \new_[59736]_  = A167 & ~A168;
  assign \new_[59737]_  = \new_[59736]_  & \new_[59733]_ ;
  assign \new_[59740]_  = A232 & ~A166;
  assign \new_[59743]_  = ~A234 & ~A233;
  assign \new_[59744]_  = \new_[59743]_  & \new_[59740]_ ;
  assign \new_[59745]_  = \new_[59744]_  & \new_[59737]_ ;
  assign \new_[59748]_  = A236 & ~A235;
  assign \new_[59751]_  = A268 & ~A267;
  assign \new_[59752]_  = \new_[59751]_  & \new_[59748]_ ;
  assign \new_[59755]_  = ~A299 & A298;
  assign \new_[59758]_  = ~A302 & A300;
  assign \new_[59759]_  = \new_[59758]_  & \new_[59755]_ ;
  assign \new_[59760]_  = \new_[59759]_  & \new_[59752]_ ;
  assign \new_[59763]_  = ~A169 & ~A170;
  assign \new_[59766]_  = A167 & ~A168;
  assign \new_[59767]_  = \new_[59766]_  & \new_[59763]_ ;
  assign \new_[59770]_  = A232 & ~A166;
  assign \new_[59773]_  = ~A234 & ~A233;
  assign \new_[59774]_  = \new_[59773]_  & \new_[59770]_ ;
  assign \new_[59775]_  = \new_[59774]_  & \new_[59767]_ ;
  assign \new_[59778]_  = A236 & ~A235;
  assign \new_[59781]_  = A268 & ~A267;
  assign \new_[59782]_  = \new_[59781]_  & \new_[59778]_ ;
  assign \new_[59785]_  = A299 & ~A298;
  assign \new_[59788]_  = A301 & A300;
  assign \new_[59789]_  = \new_[59788]_  & \new_[59785]_ ;
  assign \new_[59790]_  = \new_[59789]_  & \new_[59782]_ ;
  assign \new_[59793]_  = ~A169 & ~A170;
  assign \new_[59796]_  = A167 & ~A168;
  assign \new_[59797]_  = \new_[59796]_  & \new_[59793]_ ;
  assign \new_[59800]_  = A232 & ~A166;
  assign \new_[59803]_  = ~A234 & ~A233;
  assign \new_[59804]_  = \new_[59803]_  & \new_[59800]_ ;
  assign \new_[59805]_  = \new_[59804]_  & \new_[59797]_ ;
  assign \new_[59808]_  = A236 & ~A235;
  assign \new_[59811]_  = A268 & ~A267;
  assign \new_[59812]_  = \new_[59811]_  & \new_[59808]_ ;
  assign \new_[59815]_  = A299 & ~A298;
  assign \new_[59818]_  = ~A302 & A300;
  assign \new_[59819]_  = \new_[59818]_  & \new_[59815]_ ;
  assign \new_[59820]_  = \new_[59819]_  & \new_[59812]_ ;
  assign \new_[59823]_  = ~A169 & ~A170;
  assign \new_[59826]_  = A167 & ~A168;
  assign \new_[59827]_  = \new_[59826]_  & \new_[59823]_ ;
  assign \new_[59830]_  = A232 & ~A166;
  assign \new_[59833]_  = ~A234 & ~A233;
  assign \new_[59834]_  = \new_[59833]_  & \new_[59830]_ ;
  assign \new_[59835]_  = \new_[59834]_  & \new_[59827]_ ;
  assign \new_[59838]_  = A236 & ~A235;
  assign \new_[59841]_  = ~A269 & ~A267;
  assign \new_[59842]_  = \new_[59841]_  & \new_[59838]_ ;
  assign \new_[59845]_  = ~A299 & A298;
  assign \new_[59848]_  = A301 & A300;
  assign \new_[59849]_  = \new_[59848]_  & \new_[59845]_ ;
  assign \new_[59850]_  = \new_[59849]_  & \new_[59842]_ ;
  assign \new_[59853]_  = ~A169 & ~A170;
  assign \new_[59856]_  = A167 & ~A168;
  assign \new_[59857]_  = \new_[59856]_  & \new_[59853]_ ;
  assign \new_[59860]_  = A232 & ~A166;
  assign \new_[59863]_  = ~A234 & ~A233;
  assign \new_[59864]_  = \new_[59863]_  & \new_[59860]_ ;
  assign \new_[59865]_  = \new_[59864]_  & \new_[59857]_ ;
  assign \new_[59868]_  = A236 & ~A235;
  assign \new_[59871]_  = ~A269 & ~A267;
  assign \new_[59872]_  = \new_[59871]_  & \new_[59868]_ ;
  assign \new_[59875]_  = ~A299 & A298;
  assign \new_[59878]_  = ~A302 & A300;
  assign \new_[59879]_  = \new_[59878]_  & \new_[59875]_ ;
  assign \new_[59880]_  = \new_[59879]_  & \new_[59872]_ ;
  assign \new_[59883]_  = ~A169 & ~A170;
  assign \new_[59886]_  = A167 & ~A168;
  assign \new_[59887]_  = \new_[59886]_  & \new_[59883]_ ;
  assign \new_[59890]_  = A232 & ~A166;
  assign \new_[59893]_  = ~A234 & ~A233;
  assign \new_[59894]_  = \new_[59893]_  & \new_[59890]_ ;
  assign \new_[59895]_  = \new_[59894]_  & \new_[59887]_ ;
  assign \new_[59898]_  = A236 & ~A235;
  assign \new_[59901]_  = ~A269 & ~A267;
  assign \new_[59902]_  = \new_[59901]_  & \new_[59898]_ ;
  assign \new_[59905]_  = A299 & ~A298;
  assign \new_[59908]_  = A301 & A300;
  assign \new_[59909]_  = \new_[59908]_  & \new_[59905]_ ;
  assign \new_[59910]_  = \new_[59909]_  & \new_[59902]_ ;
  assign \new_[59913]_  = ~A169 & ~A170;
  assign \new_[59916]_  = A167 & ~A168;
  assign \new_[59917]_  = \new_[59916]_  & \new_[59913]_ ;
  assign \new_[59920]_  = A232 & ~A166;
  assign \new_[59923]_  = ~A234 & ~A233;
  assign \new_[59924]_  = \new_[59923]_  & \new_[59920]_ ;
  assign \new_[59925]_  = \new_[59924]_  & \new_[59917]_ ;
  assign \new_[59928]_  = A236 & ~A235;
  assign \new_[59931]_  = ~A269 & ~A267;
  assign \new_[59932]_  = \new_[59931]_  & \new_[59928]_ ;
  assign \new_[59935]_  = A299 & ~A298;
  assign \new_[59938]_  = ~A302 & A300;
  assign \new_[59939]_  = \new_[59938]_  & \new_[59935]_ ;
  assign \new_[59940]_  = \new_[59939]_  & \new_[59932]_ ;
  assign \new_[59943]_  = ~A169 & ~A170;
  assign \new_[59946]_  = A167 & ~A168;
  assign \new_[59947]_  = \new_[59946]_  & \new_[59943]_ ;
  assign \new_[59950]_  = A232 & ~A166;
  assign \new_[59953]_  = ~A234 & ~A233;
  assign \new_[59954]_  = \new_[59953]_  & \new_[59950]_ ;
  assign \new_[59955]_  = \new_[59954]_  & \new_[59947]_ ;
  assign \new_[59958]_  = A236 & ~A235;
  assign \new_[59961]_  = A266 & A265;
  assign \new_[59962]_  = \new_[59961]_  & \new_[59958]_ ;
  assign \new_[59965]_  = ~A299 & A298;
  assign \new_[59968]_  = A301 & A300;
  assign \new_[59969]_  = \new_[59968]_  & \new_[59965]_ ;
  assign \new_[59970]_  = \new_[59969]_  & \new_[59962]_ ;
  assign \new_[59973]_  = ~A169 & ~A170;
  assign \new_[59976]_  = A167 & ~A168;
  assign \new_[59977]_  = \new_[59976]_  & \new_[59973]_ ;
  assign \new_[59980]_  = A232 & ~A166;
  assign \new_[59983]_  = ~A234 & ~A233;
  assign \new_[59984]_  = \new_[59983]_  & \new_[59980]_ ;
  assign \new_[59985]_  = \new_[59984]_  & \new_[59977]_ ;
  assign \new_[59988]_  = A236 & ~A235;
  assign \new_[59991]_  = A266 & A265;
  assign \new_[59992]_  = \new_[59991]_  & \new_[59988]_ ;
  assign \new_[59995]_  = ~A299 & A298;
  assign \new_[59998]_  = ~A302 & A300;
  assign \new_[59999]_  = \new_[59998]_  & \new_[59995]_ ;
  assign \new_[60000]_  = \new_[59999]_  & \new_[59992]_ ;
  assign \new_[60003]_  = ~A169 & ~A170;
  assign \new_[60006]_  = A167 & ~A168;
  assign \new_[60007]_  = \new_[60006]_  & \new_[60003]_ ;
  assign \new_[60010]_  = A232 & ~A166;
  assign \new_[60013]_  = ~A234 & ~A233;
  assign \new_[60014]_  = \new_[60013]_  & \new_[60010]_ ;
  assign \new_[60015]_  = \new_[60014]_  & \new_[60007]_ ;
  assign \new_[60018]_  = A236 & ~A235;
  assign \new_[60021]_  = A266 & A265;
  assign \new_[60022]_  = \new_[60021]_  & \new_[60018]_ ;
  assign \new_[60025]_  = A299 & ~A298;
  assign \new_[60028]_  = A301 & A300;
  assign \new_[60029]_  = \new_[60028]_  & \new_[60025]_ ;
  assign \new_[60030]_  = \new_[60029]_  & \new_[60022]_ ;
  assign \new_[60033]_  = ~A169 & ~A170;
  assign \new_[60036]_  = A167 & ~A168;
  assign \new_[60037]_  = \new_[60036]_  & \new_[60033]_ ;
  assign \new_[60040]_  = A232 & ~A166;
  assign \new_[60043]_  = ~A234 & ~A233;
  assign \new_[60044]_  = \new_[60043]_  & \new_[60040]_ ;
  assign \new_[60045]_  = \new_[60044]_  & \new_[60037]_ ;
  assign \new_[60048]_  = A236 & ~A235;
  assign \new_[60051]_  = A266 & A265;
  assign \new_[60052]_  = \new_[60051]_  & \new_[60048]_ ;
  assign \new_[60055]_  = A299 & ~A298;
  assign \new_[60058]_  = ~A302 & A300;
  assign \new_[60059]_  = \new_[60058]_  & \new_[60055]_ ;
  assign \new_[60060]_  = \new_[60059]_  & \new_[60052]_ ;
  assign \new_[60063]_  = ~A169 & ~A170;
  assign \new_[60066]_  = A167 & ~A168;
  assign \new_[60067]_  = \new_[60066]_  & \new_[60063]_ ;
  assign \new_[60070]_  = A232 & ~A166;
  assign \new_[60073]_  = ~A234 & ~A233;
  assign \new_[60074]_  = \new_[60073]_  & \new_[60070]_ ;
  assign \new_[60075]_  = \new_[60074]_  & \new_[60067]_ ;
  assign \new_[60078]_  = A236 & ~A235;
  assign \new_[60081]_  = ~A266 & ~A265;
  assign \new_[60082]_  = \new_[60081]_  & \new_[60078]_ ;
  assign \new_[60085]_  = ~A299 & A298;
  assign \new_[60088]_  = A301 & A300;
  assign \new_[60089]_  = \new_[60088]_  & \new_[60085]_ ;
  assign \new_[60090]_  = \new_[60089]_  & \new_[60082]_ ;
  assign \new_[60093]_  = ~A169 & ~A170;
  assign \new_[60096]_  = A167 & ~A168;
  assign \new_[60097]_  = \new_[60096]_  & \new_[60093]_ ;
  assign \new_[60100]_  = A232 & ~A166;
  assign \new_[60103]_  = ~A234 & ~A233;
  assign \new_[60104]_  = \new_[60103]_  & \new_[60100]_ ;
  assign \new_[60105]_  = \new_[60104]_  & \new_[60097]_ ;
  assign \new_[60108]_  = A236 & ~A235;
  assign \new_[60111]_  = ~A266 & ~A265;
  assign \new_[60112]_  = \new_[60111]_  & \new_[60108]_ ;
  assign \new_[60115]_  = ~A299 & A298;
  assign \new_[60118]_  = ~A302 & A300;
  assign \new_[60119]_  = \new_[60118]_  & \new_[60115]_ ;
  assign \new_[60120]_  = \new_[60119]_  & \new_[60112]_ ;
  assign \new_[60123]_  = ~A169 & ~A170;
  assign \new_[60126]_  = A167 & ~A168;
  assign \new_[60127]_  = \new_[60126]_  & \new_[60123]_ ;
  assign \new_[60130]_  = A232 & ~A166;
  assign \new_[60133]_  = ~A234 & ~A233;
  assign \new_[60134]_  = \new_[60133]_  & \new_[60130]_ ;
  assign \new_[60135]_  = \new_[60134]_  & \new_[60127]_ ;
  assign \new_[60138]_  = A236 & ~A235;
  assign \new_[60141]_  = ~A266 & ~A265;
  assign \new_[60142]_  = \new_[60141]_  & \new_[60138]_ ;
  assign \new_[60145]_  = A299 & ~A298;
  assign \new_[60148]_  = A301 & A300;
  assign \new_[60149]_  = \new_[60148]_  & \new_[60145]_ ;
  assign \new_[60150]_  = \new_[60149]_  & \new_[60142]_ ;
  assign \new_[60153]_  = ~A169 & ~A170;
  assign \new_[60156]_  = A167 & ~A168;
  assign \new_[60157]_  = \new_[60156]_  & \new_[60153]_ ;
  assign \new_[60160]_  = A232 & ~A166;
  assign \new_[60163]_  = ~A234 & ~A233;
  assign \new_[60164]_  = \new_[60163]_  & \new_[60160]_ ;
  assign \new_[60165]_  = \new_[60164]_  & \new_[60157]_ ;
  assign \new_[60168]_  = A236 & ~A235;
  assign \new_[60171]_  = ~A266 & ~A265;
  assign \new_[60172]_  = \new_[60171]_  & \new_[60168]_ ;
  assign \new_[60175]_  = A299 & ~A298;
  assign \new_[60178]_  = ~A302 & A300;
  assign \new_[60179]_  = \new_[60178]_  & \new_[60175]_ ;
  assign \new_[60180]_  = \new_[60179]_  & \new_[60172]_ ;
  assign \new_[60183]_  = ~A169 & ~A170;
  assign \new_[60186]_  = ~A167 & ~A168;
  assign \new_[60187]_  = \new_[60186]_  & \new_[60183]_ ;
  assign \new_[60190]_  = ~A232 & A166;
  assign \new_[60193]_  = A234 & A233;
  assign \new_[60194]_  = \new_[60193]_  & \new_[60190]_ ;
  assign \new_[60195]_  = \new_[60194]_  & \new_[60187]_ ;
  assign \new_[60198]_  = A267 & A235;
  assign \new_[60201]_  = A269 & ~A268;
  assign \new_[60202]_  = \new_[60201]_  & \new_[60198]_ ;
  assign \new_[60205]_  = ~A299 & A298;
  assign \new_[60208]_  = A301 & A300;
  assign \new_[60209]_  = \new_[60208]_  & \new_[60205]_ ;
  assign \new_[60210]_  = \new_[60209]_  & \new_[60202]_ ;
  assign \new_[60213]_  = ~A169 & ~A170;
  assign \new_[60216]_  = ~A167 & ~A168;
  assign \new_[60217]_  = \new_[60216]_  & \new_[60213]_ ;
  assign \new_[60220]_  = ~A232 & A166;
  assign \new_[60223]_  = A234 & A233;
  assign \new_[60224]_  = \new_[60223]_  & \new_[60220]_ ;
  assign \new_[60225]_  = \new_[60224]_  & \new_[60217]_ ;
  assign \new_[60228]_  = A267 & A235;
  assign \new_[60231]_  = A269 & ~A268;
  assign \new_[60232]_  = \new_[60231]_  & \new_[60228]_ ;
  assign \new_[60235]_  = ~A299 & A298;
  assign \new_[60238]_  = ~A302 & A300;
  assign \new_[60239]_  = \new_[60238]_  & \new_[60235]_ ;
  assign \new_[60240]_  = \new_[60239]_  & \new_[60232]_ ;
  assign \new_[60243]_  = ~A169 & ~A170;
  assign \new_[60246]_  = ~A167 & ~A168;
  assign \new_[60247]_  = \new_[60246]_  & \new_[60243]_ ;
  assign \new_[60250]_  = ~A232 & A166;
  assign \new_[60253]_  = A234 & A233;
  assign \new_[60254]_  = \new_[60253]_  & \new_[60250]_ ;
  assign \new_[60255]_  = \new_[60254]_  & \new_[60247]_ ;
  assign \new_[60258]_  = A267 & A235;
  assign \new_[60261]_  = A269 & ~A268;
  assign \new_[60262]_  = \new_[60261]_  & \new_[60258]_ ;
  assign \new_[60265]_  = A299 & ~A298;
  assign \new_[60268]_  = A301 & A300;
  assign \new_[60269]_  = \new_[60268]_  & \new_[60265]_ ;
  assign \new_[60270]_  = \new_[60269]_  & \new_[60262]_ ;
  assign \new_[60273]_  = ~A169 & ~A170;
  assign \new_[60276]_  = ~A167 & ~A168;
  assign \new_[60277]_  = \new_[60276]_  & \new_[60273]_ ;
  assign \new_[60280]_  = ~A232 & A166;
  assign \new_[60283]_  = A234 & A233;
  assign \new_[60284]_  = \new_[60283]_  & \new_[60280]_ ;
  assign \new_[60285]_  = \new_[60284]_  & \new_[60277]_ ;
  assign \new_[60288]_  = A267 & A235;
  assign \new_[60291]_  = A269 & ~A268;
  assign \new_[60292]_  = \new_[60291]_  & \new_[60288]_ ;
  assign \new_[60295]_  = A299 & ~A298;
  assign \new_[60298]_  = ~A302 & A300;
  assign \new_[60299]_  = \new_[60298]_  & \new_[60295]_ ;
  assign \new_[60300]_  = \new_[60299]_  & \new_[60292]_ ;
  assign \new_[60303]_  = ~A169 & ~A170;
  assign \new_[60306]_  = ~A167 & ~A168;
  assign \new_[60307]_  = \new_[60306]_  & \new_[60303]_ ;
  assign \new_[60310]_  = ~A232 & A166;
  assign \new_[60313]_  = A234 & A233;
  assign \new_[60314]_  = \new_[60313]_  & \new_[60310]_ ;
  assign \new_[60315]_  = \new_[60314]_  & \new_[60307]_ ;
  assign \new_[60318]_  = ~A267 & A235;
  assign \new_[60321]_  = A298 & A268;
  assign \new_[60322]_  = \new_[60321]_  & \new_[60318]_ ;
  assign \new_[60325]_  = ~A300 & ~A299;
  assign \new_[60328]_  = A302 & ~A301;
  assign \new_[60329]_  = \new_[60328]_  & \new_[60325]_ ;
  assign \new_[60330]_  = \new_[60329]_  & \new_[60322]_ ;
  assign \new_[60333]_  = ~A169 & ~A170;
  assign \new_[60336]_  = ~A167 & ~A168;
  assign \new_[60337]_  = \new_[60336]_  & \new_[60333]_ ;
  assign \new_[60340]_  = ~A232 & A166;
  assign \new_[60343]_  = A234 & A233;
  assign \new_[60344]_  = \new_[60343]_  & \new_[60340]_ ;
  assign \new_[60345]_  = \new_[60344]_  & \new_[60337]_ ;
  assign \new_[60348]_  = ~A267 & A235;
  assign \new_[60351]_  = ~A298 & A268;
  assign \new_[60352]_  = \new_[60351]_  & \new_[60348]_ ;
  assign \new_[60355]_  = ~A300 & A299;
  assign \new_[60358]_  = A302 & ~A301;
  assign \new_[60359]_  = \new_[60358]_  & \new_[60355]_ ;
  assign \new_[60360]_  = \new_[60359]_  & \new_[60352]_ ;
  assign \new_[60363]_  = ~A169 & ~A170;
  assign \new_[60366]_  = ~A167 & ~A168;
  assign \new_[60367]_  = \new_[60366]_  & \new_[60363]_ ;
  assign \new_[60370]_  = ~A232 & A166;
  assign \new_[60373]_  = A234 & A233;
  assign \new_[60374]_  = \new_[60373]_  & \new_[60370]_ ;
  assign \new_[60375]_  = \new_[60374]_  & \new_[60367]_ ;
  assign \new_[60378]_  = ~A267 & A235;
  assign \new_[60381]_  = A298 & ~A269;
  assign \new_[60382]_  = \new_[60381]_  & \new_[60378]_ ;
  assign \new_[60385]_  = ~A300 & ~A299;
  assign \new_[60388]_  = A302 & ~A301;
  assign \new_[60389]_  = \new_[60388]_  & \new_[60385]_ ;
  assign \new_[60390]_  = \new_[60389]_  & \new_[60382]_ ;
  assign \new_[60393]_  = ~A169 & ~A170;
  assign \new_[60396]_  = ~A167 & ~A168;
  assign \new_[60397]_  = \new_[60396]_  & \new_[60393]_ ;
  assign \new_[60400]_  = ~A232 & A166;
  assign \new_[60403]_  = A234 & A233;
  assign \new_[60404]_  = \new_[60403]_  & \new_[60400]_ ;
  assign \new_[60405]_  = \new_[60404]_  & \new_[60397]_ ;
  assign \new_[60408]_  = ~A267 & A235;
  assign \new_[60411]_  = ~A298 & ~A269;
  assign \new_[60412]_  = \new_[60411]_  & \new_[60408]_ ;
  assign \new_[60415]_  = ~A300 & A299;
  assign \new_[60418]_  = A302 & ~A301;
  assign \new_[60419]_  = \new_[60418]_  & \new_[60415]_ ;
  assign \new_[60420]_  = \new_[60419]_  & \new_[60412]_ ;
  assign \new_[60423]_  = ~A169 & ~A170;
  assign \new_[60426]_  = ~A167 & ~A168;
  assign \new_[60427]_  = \new_[60426]_  & \new_[60423]_ ;
  assign \new_[60430]_  = ~A232 & A166;
  assign \new_[60433]_  = A234 & A233;
  assign \new_[60434]_  = \new_[60433]_  & \new_[60430]_ ;
  assign \new_[60435]_  = \new_[60434]_  & \new_[60427]_ ;
  assign \new_[60438]_  = A265 & A235;
  assign \new_[60441]_  = A298 & A266;
  assign \new_[60442]_  = \new_[60441]_  & \new_[60438]_ ;
  assign \new_[60445]_  = ~A300 & ~A299;
  assign \new_[60448]_  = A302 & ~A301;
  assign \new_[60449]_  = \new_[60448]_  & \new_[60445]_ ;
  assign \new_[60450]_  = \new_[60449]_  & \new_[60442]_ ;
  assign \new_[60453]_  = ~A169 & ~A170;
  assign \new_[60456]_  = ~A167 & ~A168;
  assign \new_[60457]_  = \new_[60456]_  & \new_[60453]_ ;
  assign \new_[60460]_  = ~A232 & A166;
  assign \new_[60463]_  = A234 & A233;
  assign \new_[60464]_  = \new_[60463]_  & \new_[60460]_ ;
  assign \new_[60465]_  = \new_[60464]_  & \new_[60457]_ ;
  assign \new_[60468]_  = A265 & A235;
  assign \new_[60471]_  = ~A298 & A266;
  assign \new_[60472]_  = \new_[60471]_  & \new_[60468]_ ;
  assign \new_[60475]_  = ~A300 & A299;
  assign \new_[60478]_  = A302 & ~A301;
  assign \new_[60479]_  = \new_[60478]_  & \new_[60475]_ ;
  assign \new_[60480]_  = \new_[60479]_  & \new_[60472]_ ;
  assign \new_[60483]_  = ~A169 & ~A170;
  assign \new_[60486]_  = ~A167 & ~A168;
  assign \new_[60487]_  = \new_[60486]_  & \new_[60483]_ ;
  assign \new_[60490]_  = ~A232 & A166;
  assign \new_[60493]_  = A234 & A233;
  assign \new_[60494]_  = \new_[60493]_  & \new_[60490]_ ;
  assign \new_[60495]_  = \new_[60494]_  & \new_[60487]_ ;
  assign \new_[60498]_  = ~A265 & A235;
  assign \new_[60501]_  = A298 & ~A266;
  assign \new_[60502]_  = \new_[60501]_  & \new_[60498]_ ;
  assign \new_[60505]_  = ~A300 & ~A299;
  assign \new_[60508]_  = A302 & ~A301;
  assign \new_[60509]_  = \new_[60508]_  & \new_[60505]_ ;
  assign \new_[60510]_  = \new_[60509]_  & \new_[60502]_ ;
  assign \new_[60513]_  = ~A169 & ~A170;
  assign \new_[60516]_  = ~A167 & ~A168;
  assign \new_[60517]_  = \new_[60516]_  & \new_[60513]_ ;
  assign \new_[60520]_  = ~A232 & A166;
  assign \new_[60523]_  = A234 & A233;
  assign \new_[60524]_  = \new_[60523]_  & \new_[60520]_ ;
  assign \new_[60525]_  = \new_[60524]_  & \new_[60517]_ ;
  assign \new_[60528]_  = ~A265 & A235;
  assign \new_[60531]_  = ~A298 & ~A266;
  assign \new_[60532]_  = \new_[60531]_  & \new_[60528]_ ;
  assign \new_[60535]_  = ~A300 & A299;
  assign \new_[60538]_  = A302 & ~A301;
  assign \new_[60539]_  = \new_[60538]_  & \new_[60535]_ ;
  assign \new_[60540]_  = \new_[60539]_  & \new_[60532]_ ;
  assign \new_[60543]_  = ~A169 & ~A170;
  assign \new_[60546]_  = ~A167 & ~A168;
  assign \new_[60547]_  = \new_[60546]_  & \new_[60543]_ ;
  assign \new_[60550]_  = ~A232 & A166;
  assign \new_[60553]_  = A234 & A233;
  assign \new_[60554]_  = \new_[60553]_  & \new_[60550]_ ;
  assign \new_[60555]_  = \new_[60554]_  & \new_[60547]_ ;
  assign \new_[60558]_  = A267 & ~A236;
  assign \new_[60561]_  = A269 & ~A268;
  assign \new_[60562]_  = \new_[60561]_  & \new_[60558]_ ;
  assign \new_[60565]_  = ~A299 & A298;
  assign \new_[60568]_  = A301 & A300;
  assign \new_[60569]_  = \new_[60568]_  & \new_[60565]_ ;
  assign \new_[60570]_  = \new_[60569]_  & \new_[60562]_ ;
  assign \new_[60573]_  = ~A169 & ~A170;
  assign \new_[60576]_  = ~A167 & ~A168;
  assign \new_[60577]_  = \new_[60576]_  & \new_[60573]_ ;
  assign \new_[60580]_  = ~A232 & A166;
  assign \new_[60583]_  = A234 & A233;
  assign \new_[60584]_  = \new_[60583]_  & \new_[60580]_ ;
  assign \new_[60585]_  = \new_[60584]_  & \new_[60577]_ ;
  assign \new_[60588]_  = A267 & ~A236;
  assign \new_[60591]_  = A269 & ~A268;
  assign \new_[60592]_  = \new_[60591]_  & \new_[60588]_ ;
  assign \new_[60595]_  = ~A299 & A298;
  assign \new_[60598]_  = ~A302 & A300;
  assign \new_[60599]_  = \new_[60598]_  & \new_[60595]_ ;
  assign \new_[60600]_  = \new_[60599]_  & \new_[60592]_ ;
  assign \new_[60603]_  = ~A169 & ~A170;
  assign \new_[60606]_  = ~A167 & ~A168;
  assign \new_[60607]_  = \new_[60606]_  & \new_[60603]_ ;
  assign \new_[60610]_  = ~A232 & A166;
  assign \new_[60613]_  = A234 & A233;
  assign \new_[60614]_  = \new_[60613]_  & \new_[60610]_ ;
  assign \new_[60615]_  = \new_[60614]_  & \new_[60607]_ ;
  assign \new_[60618]_  = A267 & ~A236;
  assign \new_[60621]_  = A269 & ~A268;
  assign \new_[60622]_  = \new_[60621]_  & \new_[60618]_ ;
  assign \new_[60625]_  = A299 & ~A298;
  assign \new_[60628]_  = A301 & A300;
  assign \new_[60629]_  = \new_[60628]_  & \new_[60625]_ ;
  assign \new_[60630]_  = \new_[60629]_  & \new_[60622]_ ;
  assign \new_[60633]_  = ~A169 & ~A170;
  assign \new_[60636]_  = ~A167 & ~A168;
  assign \new_[60637]_  = \new_[60636]_  & \new_[60633]_ ;
  assign \new_[60640]_  = ~A232 & A166;
  assign \new_[60643]_  = A234 & A233;
  assign \new_[60644]_  = \new_[60643]_  & \new_[60640]_ ;
  assign \new_[60645]_  = \new_[60644]_  & \new_[60637]_ ;
  assign \new_[60648]_  = A267 & ~A236;
  assign \new_[60651]_  = A269 & ~A268;
  assign \new_[60652]_  = \new_[60651]_  & \new_[60648]_ ;
  assign \new_[60655]_  = A299 & ~A298;
  assign \new_[60658]_  = ~A302 & A300;
  assign \new_[60659]_  = \new_[60658]_  & \new_[60655]_ ;
  assign \new_[60660]_  = \new_[60659]_  & \new_[60652]_ ;
  assign \new_[60663]_  = ~A169 & ~A170;
  assign \new_[60666]_  = ~A167 & ~A168;
  assign \new_[60667]_  = \new_[60666]_  & \new_[60663]_ ;
  assign \new_[60670]_  = ~A232 & A166;
  assign \new_[60673]_  = A234 & A233;
  assign \new_[60674]_  = \new_[60673]_  & \new_[60670]_ ;
  assign \new_[60675]_  = \new_[60674]_  & \new_[60667]_ ;
  assign \new_[60678]_  = ~A267 & ~A236;
  assign \new_[60681]_  = A298 & A268;
  assign \new_[60682]_  = \new_[60681]_  & \new_[60678]_ ;
  assign \new_[60685]_  = ~A300 & ~A299;
  assign \new_[60688]_  = A302 & ~A301;
  assign \new_[60689]_  = \new_[60688]_  & \new_[60685]_ ;
  assign \new_[60690]_  = \new_[60689]_  & \new_[60682]_ ;
  assign \new_[60693]_  = ~A169 & ~A170;
  assign \new_[60696]_  = ~A167 & ~A168;
  assign \new_[60697]_  = \new_[60696]_  & \new_[60693]_ ;
  assign \new_[60700]_  = ~A232 & A166;
  assign \new_[60703]_  = A234 & A233;
  assign \new_[60704]_  = \new_[60703]_  & \new_[60700]_ ;
  assign \new_[60705]_  = \new_[60704]_  & \new_[60697]_ ;
  assign \new_[60708]_  = ~A267 & ~A236;
  assign \new_[60711]_  = ~A298 & A268;
  assign \new_[60712]_  = \new_[60711]_  & \new_[60708]_ ;
  assign \new_[60715]_  = ~A300 & A299;
  assign \new_[60718]_  = A302 & ~A301;
  assign \new_[60719]_  = \new_[60718]_  & \new_[60715]_ ;
  assign \new_[60720]_  = \new_[60719]_  & \new_[60712]_ ;
  assign \new_[60723]_  = ~A169 & ~A170;
  assign \new_[60726]_  = ~A167 & ~A168;
  assign \new_[60727]_  = \new_[60726]_  & \new_[60723]_ ;
  assign \new_[60730]_  = ~A232 & A166;
  assign \new_[60733]_  = A234 & A233;
  assign \new_[60734]_  = \new_[60733]_  & \new_[60730]_ ;
  assign \new_[60735]_  = \new_[60734]_  & \new_[60727]_ ;
  assign \new_[60738]_  = ~A267 & ~A236;
  assign \new_[60741]_  = A298 & ~A269;
  assign \new_[60742]_  = \new_[60741]_  & \new_[60738]_ ;
  assign \new_[60745]_  = ~A300 & ~A299;
  assign \new_[60748]_  = A302 & ~A301;
  assign \new_[60749]_  = \new_[60748]_  & \new_[60745]_ ;
  assign \new_[60750]_  = \new_[60749]_  & \new_[60742]_ ;
  assign \new_[60753]_  = ~A169 & ~A170;
  assign \new_[60756]_  = ~A167 & ~A168;
  assign \new_[60757]_  = \new_[60756]_  & \new_[60753]_ ;
  assign \new_[60760]_  = ~A232 & A166;
  assign \new_[60763]_  = A234 & A233;
  assign \new_[60764]_  = \new_[60763]_  & \new_[60760]_ ;
  assign \new_[60765]_  = \new_[60764]_  & \new_[60757]_ ;
  assign \new_[60768]_  = ~A267 & ~A236;
  assign \new_[60771]_  = ~A298 & ~A269;
  assign \new_[60772]_  = \new_[60771]_  & \new_[60768]_ ;
  assign \new_[60775]_  = ~A300 & A299;
  assign \new_[60778]_  = A302 & ~A301;
  assign \new_[60779]_  = \new_[60778]_  & \new_[60775]_ ;
  assign \new_[60780]_  = \new_[60779]_  & \new_[60772]_ ;
  assign \new_[60783]_  = ~A169 & ~A170;
  assign \new_[60786]_  = ~A167 & ~A168;
  assign \new_[60787]_  = \new_[60786]_  & \new_[60783]_ ;
  assign \new_[60790]_  = ~A232 & A166;
  assign \new_[60793]_  = A234 & A233;
  assign \new_[60794]_  = \new_[60793]_  & \new_[60790]_ ;
  assign \new_[60795]_  = \new_[60794]_  & \new_[60787]_ ;
  assign \new_[60798]_  = A265 & ~A236;
  assign \new_[60801]_  = A298 & A266;
  assign \new_[60802]_  = \new_[60801]_  & \new_[60798]_ ;
  assign \new_[60805]_  = ~A300 & ~A299;
  assign \new_[60808]_  = A302 & ~A301;
  assign \new_[60809]_  = \new_[60808]_  & \new_[60805]_ ;
  assign \new_[60810]_  = \new_[60809]_  & \new_[60802]_ ;
  assign \new_[60813]_  = ~A169 & ~A170;
  assign \new_[60816]_  = ~A167 & ~A168;
  assign \new_[60817]_  = \new_[60816]_  & \new_[60813]_ ;
  assign \new_[60820]_  = ~A232 & A166;
  assign \new_[60823]_  = A234 & A233;
  assign \new_[60824]_  = \new_[60823]_  & \new_[60820]_ ;
  assign \new_[60825]_  = \new_[60824]_  & \new_[60817]_ ;
  assign \new_[60828]_  = A265 & ~A236;
  assign \new_[60831]_  = ~A298 & A266;
  assign \new_[60832]_  = \new_[60831]_  & \new_[60828]_ ;
  assign \new_[60835]_  = ~A300 & A299;
  assign \new_[60838]_  = A302 & ~A301;
  assign \new_[60839]_  = \new_[60838]_  & \new_[60835]_ ;
  assign \new_[60840]_  = \new_[60839]_  & \new_[60832]_ ;
  assign \new_[60843]_  = ~A169 & ~A170;
  assign \new_[60846]_  = ~A167 & ~A168;
  assign \new_[60847]_  = \new_[60846]_  & \new_[60843]_ ;
  assign \new_[60850]_  = ~A232 & A166;
  assign \new_[60853]_  = A234 & A233;
  assign \new_[60854]_  = \new_[60853]_  & \new_[60850]_ ;
  assign \new_[60855]_  = \new_[60854]_  & \new_[60847]_ ;
  assign \new_[60858]_  = ~A265 & ~A236;
  assign \new_[60861]_  = A298 & ~A266;
  assign \new_[60862]_  = \new_[60861]_  & \new_[60858]_ ;
  assign \new_[60865]_  = ~A300 & ~A299;
  assign \new_[60868]_  = A302 & ~A301;
  assign \new_[60869]_  = \new_[60868]_  & \new_[60865]_ ;
  assign \new_[60870]_  = \new_[60869]_  & \new_[60862]_ ;
  assign \new_[60873]_  = ~A169 & ~A170;
  assign \new_[60876]_  = ~A167 & ~A168;
  assign \new_[60877]_  = \new_[60876]_  & \new_[60873]_ ;
  assign \new_[60880]_  = ~A232 & A166;
  assign \new_[60883]_  = A234 & A233;
  assign \new_[60884]_  = \new_[60883]_  & \new_[60880]_ ;
  assign \new_[60885]_  = \new_[60884]_  & \new_[60877]_ ;
  assign \new_[60888]_  = ~A265 & ~A236;
  assign \new_[60891]_  = ~A298 & ~A266;
  assign \new_[60892]_  = \new_[60891]_  & \new_[60888]_ ;
  assign \new_[60895]_  = ~A300 & A299;
  assign \new_[60898]_  = A302 & ~A301;
  assign \new_[60899]_  = \new_[60898]_  & \new_[60895]_ ;
  assign \new_[60900]_  = \new_[60899]_  & \new_[60892]_ ;
  assign \new_[60903]_  = ~A169 & ~A170;
  assign \new_[60906]_  = ~A167 & ~A168;
  assign \new_[60907]_  = \new_[60906]_  & \new_[60903]_ ;
  assign \new_[60910]_  = ~A232 & A166;
  assign \new_[60913]_  = ~A234 & A233;
  assign \new_[60914]_  = \new_[60913]_  & \new_[60910]_ ;
  assign \new_[60915]_  = \new_[60914]_  & \new_[60907]_ ;
  assign \new_[60918]_  = A236 & ~A235;
  assign \new_[60921]_  = A268 & ~A267;
  assign \new_[60922]_  = \new_[60921]_  & \new_[60918]_ ;
  assign \new_[60925]_  = ~A299 & A298;
  assign \new_[60928]_  = A301 & A300;
  assign \new_[60929]_  = \new_[60928]_  & \new_[60925]_ ;
  assign \new_[60930]_  = \new_[60929]_  & \new_[60922]_ ;
  assign \new_[60933]_  = ~A169 & ~A170;
  assign \new_[60936]_  = ~A167 & ~A168;
  assign \new_[60937]_  = \new_[60936]_  & \new_[60933]_ ;
  assign \new_[60940]_  = ~A232 & A166;
  assign \new_[60943]_  = ~A234 & A233;
  assign \new_[60944]_  = \new_[60943]_  & \new_[60940]_ ;
  assign \new_[60945]_  = \new_[60944]_  & \new_[60937]_ ;
  assign \new_[60948]_  = A236 & ~A235;
  assign \new_[60951]_  = A268 & ~A267;
  assign \new_[60952]_  = \new_[60951]_  & \new_[60948]_ ;
  assign \new_[60955]_  = ~A299 & A298;
  assign \new_[60958]_  = ~A302 & A300;
  assign \new_[60959]_  = \new_[60958]_  & \new_[60955]_ ;
  assign \new_[60960]_  = \new_[60959]_  & \new_[60952]_ ;
  assign \new_[60963]_  = ~A169 & ~A170;
  assign \new_[60966]_  = ~A167 & ~A168;
  assign \new_[60967]_  = \new_[60966]_  & \new_[60963]_ ;
  assign \new_[60970]_  = ~A232 & A166;
  assign \new_[60973]_  = ~A234 & A233;
  assign \new_[60974]_  = \new_[60973]_  & \new_[60970]_ ;
  assign \new_[60975]_  = \new_[60974]_  & \new_[60967]_ ;
  assign \new_[60978]_  = A236 & ~A235;
  assign \new_[60981]_  = A268 & ~A267;
  assign \new_[60982]_  = \new_[60981]_  & \new_[60978]_ ;
  assign \new_[60985]_  = A299 & ~A298;
  assign \new_[60988]_  = A301 & A300;
  assign \new_[60989]_  = \new_[60988]_  & \new_[60985]_ ;
  assign \new_[60990]_  = \new_[60989]_  & \new_[60982]_ ;
  assign \new_[60993]_  = ~A169 & ~A170;
  assign \new_[60996]_  = ~A167 & ~A168;
  assign \new_[60997]_  = \new_[60996]_  & \new_[60993]_ ;
  assign \new_[61000]_  = ~A232 & A166;
  assign \new_[61003]_  = ~A234 & A233;
  assign \new_[61004]_  = \new_[61003]_  & \new_[61000]_ ;
  assign \new_[61005]_  = \new_[61004]_  & \new_[60997]_ ;
  assign \new_[61008]_  = A236 & ~A235;
  assign \new_[61011]_  = A268 & ~A267;
  assign \new_[61012]_  = \new_[61011]_  & \new_[61008]_ ;
  assign \new_[61015]_  = A299 & ~A298;
  assign \new_[61018]_  = ~A302 & A300;
  assign \new_[61019]_  = \new_[61018]_  & \new_[61015]_ ;
  assign \new_[61020]_  = \new_[61019]_  & \new_[61012]_ ;
  assign \new_[61023]_  = ~A169 & ~A170;
  assign \new_[61026]_  = ~A167 & ~A168;
  assign \new_[61027]_  = \new_[61026]_  & \new_[61023]_ ;
  assign \new_[61030]_  = ~A232 & A166;
  assign \new_[61033]_  = ~A234 & A233;
  assign \new_[61034]_  = \new_[61033]_  & \new_[61030]_ ;
  assign \new_[61035]_  = \new_[61034]_  & \new_[61027]_ ;
  assign \new_[61038]_  = A236 & ~A235;
  assign \new_[61041]_  = ~A269 & ~A267;
  assign \new_[61042]_  = \new_[61041]_  & \new_[61038]_ ;
  assign \new_[61045]_  = ~A299 & A298;
  assign \new_[61048]_  = A301 & A300;
  assign \new_[61049]_  = \new_[61048]_  & \new_[61045]_ ;
  assign \new_[61050]_  = \new_[61049]_  & \new_[61042]_ ;
  assign \new_[61053]_  = ~A169 & ~A170;
  assign \new_[61056]_  = ~A167 & ~A168;
  assign \new_[61057]_  = \new_[61056]_  & \new_[61053]_ ;
  assign \new_[61060]_  = ~A232 & A166;
  assign \new_[61063]_  = ~A234 & A233;
  assign \new_[61064]_  = \new_[61063]_  & \new_[61060]_ ;
  assign \new_[61065]_  = \new_[61064]_  & \new_[61057]_ ;
  assign \new_[61068]_  = A236 & ~A235;
  assign \new_[61071]_  = ~A269 & ~A267;
  assign \new_[61072]_  = \new_[61071]_  & \new_[61068]_ ;
  assign \new_[61075]_  = ~A299 & A298;
  assign \new_[61078]_  = ~A302 & A300;
  assign \new_[61079]_  = \new_[61078]_  & \new_[61075]_ ;
  assign \new_[61080]_  = \new_[61079]_  & \new_[61072]_ ;
  assign \new_[61083]_  = ~A169 & ~A170;
  assign \new_[61086]_  = ~A167 & ~A168;
  assign \new_[61087]_  = \new_[61086]_  & \new_[61083]_ ;
  assign \new_[61090]_  = ~A232 & A166;
  assign \new_[61093]_  = ~A234 & A233;
  assign \new_[61094]_  = \new_[61093]_  & \new_[61090]_ ;
  assign \new_[61095]_  = \new_[61094]_  & \new_[61087]_ ;
  assign \new_[61098]_  = A236 & ~A235;
  assign \new_[61101]_  = ~A269 & ~A267;
  assign \new_[61102]_  = \new_[61101]_  & \new_[61098]_ ;
  assign \new_[61105]_  = A299 & ~A298;
  assign \new_[61108]_  = A301 & A300;
  assign \new_[61109]_  = \new_[61108]_  & \new_[61105]_ ;
  assign \new_[61110]_  = \new_[61109]_  & \new_[61102]_ ;
  assign \new_[61113]_  = ~A169 & ~A170;
  assign \new_[61116]_  = ~A167 & ~A168;
  assign \new_[61117]_  = \new_[61116]_  & \new_[61113]_ ;
  assign \new_[61120]_  = ~A232 & A166;
  assign \new_[61123]_  = ~A234 & A233;
  assign \new_[61124]_  = \new_[61123]_  & \new_[61120]_ ;
  assign \new_[61125]_  = \new_[61124]_  & \new_[61117]_ ;
  assign \new_[61128]_  = A236 & ~A235;
  assign \new_[61131]_  = ~A269 & ~A267;
  assign \new_[61132]_  = \new_[61131]_  & \new_[61128]_ ;
  assign \new_[61135]_  = A299 & ~A298;
  assign \new_[61138]_  = ~A302 & A300;
  assign \new_[61139]_  = \new_[61138]_  & \new_[61135]_ ;
  assign \new_[61140]_  = \new_[61139]_  & \new_[61132]_ ;
  assign \new_[61143]_  = ~A169 & ~A170;
  assign \new_[61146]_  = ~A167 & ~A168;
  assign \new_[61147]_  = \new_[61146]_  & \new_[61143]_ ;
  assign \new_[61150]_  = ~A232 & A166;
  assign \new_[61153]_  = ~A234 & A233;
  assign \new_[61154]_  = \new_[61153]_  & \new_[61150]_ ;
  assign \new_[61155]_  = \new_[61154]_  & \new_[61147]_ ;
  assign \new_[61158]_  = A236 & ~A235;
  assign \new_[61161]_  = A266 & A265;
  assign \new_[61162]_  = \new_[61161]_  & \new_[61158]_ ;
  assign \new_[61165]_  = ~A299 & A298;
  assign \new_[61168]_  = A301 & A300;
  assign \new_[61169]_  = \new_[61168]_  & \new_[61165]_ ;
  assign \new_[61170]_  = \new_[61169]_  & \new_[61162]_ ;
  assign \new_[61173]_  = ~A169 & ~A170;
  assign \new_[61176]_  = ~A167 & ~A168;
  assign \new_[61177]_  = \new_[61176]_  & \new_[61173]_ ;
  assign \new_[61180]_  = ~A232 & A166;
  assign \new_[61183]_  = ~A234 & A233;
  assign \new_[61184]_  = \new_[61183]_  & \new_[61180]_ ;
  assign \new_[61185]_  = \new_[61184]_  & \new_[61177]_ ;
  assign \new_[61188]_  = A236 & ~A235;
  assign \new_[61191]_  = A266 & A265;
  assign \new_[61192]_  = \new_[61191]_  & \new_[61188]_ ;
  assign \new_[61195]_  = ~A299 & A298;
  assign \new_[61198]_  = ~A302 & A300;
  assign \new_[61199]_  = \new_[61198]_  & \new_[61195]_ ;
  assign \new_[61200]_  = \new_[61199]_  & \new_[61192]_ ;
  assign \new_[61203]_  = ~A169 & ~A170;
  assign \new_[61206]_  = ~A167 & ~A168;
  assign \new_[61207]_  = \new_[61206]_  & \new_[61203]_ ;
  assign \new_[61210]_  = ~A232 & A166;
  assign \new_[61213]_  = ~A234 & A233;
  assign \new_[61214]_  = \new_[61213]_  & \new_[61210]_ ;
  assign \new_[61215]_  = \new_[61214]_  & \new_[61207]_ ;
  assign \new_[61218]_  = A236 & ~A235;
  assign \new_[61221]_  = A266 & A265;
  assign \new_[61222]_  = \new_[61221]_  & \new_[61218]_ ;
  assign \new_[61225]_  = A299 & ~A298;
  assign \new_[61228]_  = A301 & A300;
  assign \new_[61229]_  = \new_[61228]_  & \new_[61225]_ ;
  assign \new_[61230]_  = \new_[61229]_  & \new_[61222]_ ;
  assign \new_[61233]_  = ~A169 & ~A170;
  assign \new_[61236]_  = ~A167 & ~A168;
  assign \new_[61237]_  = \new_[61236]_  & \new_[61233]_ ;
  assign \new_[61240]_  = ~A232 & A166;
  assign \new_[61243]_  = ~A234 & A233;
  assign \new_[61244]_  = \new_[61243]_  & \new_[61240]_ ;
  assign \new_[61245]_  = \new_[61244]_  & \new_[61237]_ ;
  assign \new_[61248]_  = A236 & ~A235;
  assign \new_[61251]_  = A266 & A265;
  assign \new_[61252]_  = \new_[61251]_  & \new_[61248]_ ;
  assign \new_[61255]_  = A299 & ~A298;
  assign \new_[61258]_  = ~A302 & A300;
  assign \new_[61259]_  = \new_[61258]_  & \new_[61255]_ ;
  assign \new_[61260]_  = \new_[61259]_  & \new_[61252]_ ;
  assign \new_[61263]_  = ~A169 & ~A170;
  assign \new_[61266]_  = ~A167 & ~A168;
  assign \new_[61267]_  = \new_[61266]_  & \new_[61263]_ ;
  assign \new_[61270]_  = ~A232 & A166;
  assign \new_[61273]_  = ~A234 & A233;
  assign \new_[61274]_  = \new_[61273]_  & \new_[61270]_ ;
  assign \new_[61275]_  = \new_[61274]_  & \new_[61267]_ ;
  assign \new_[61278]_  = A236 & ~A235;
  assign \new_[61281]_  = ~A266 & ~A265;
  assign \new_[61282]_  = \new_[61281]_  & \new_[61278]_ ;
  assign \new_[61285]_  = ~A299 & A298;
  assign \new_[61288]_  = A301 & A300;
  assign \new_[61289]_  = \new_[61288]_  & \new_[61285]_ ;
  assign \new_[61290]_  = \new_[61289]_  & \new_[61282]_ ;
  assign \new_[61293]_  = ~A169 & ~A170;
  assign \new_[61296]_  = ~A167 & ~A168;
  assign \new_[61297]_  = \new_[61296]_  & \new_[61293]_ ;
  assign \new_[61300]_  = ~A232 & A166;
  assign \new_[61303]_  = ~A234 & A233;
  assign \new_[61304]_  = \new_[61303]_  & \new_[61300]_ ;
  assign \new_[61305]_  = \new_[61304]_  & \new_[61297]_ ;
  assign \new_[61308]_  = A236 & ~A235;
  assign \new_[61311]_  = ~A266 & ~A265;
  assign \new_[61312]_  = \new_[61311]_  & \new_[61308]_ ;
  assign \new_[61315]_  = ~A299 & A298;
  assign \new_[61318]_  = ~A302 & A300;
  assign \new_[61319]_  = \new_[61318]_  & \new_[61315]_ ;
  assign \new_[61320]_  = \new_[61319]_  & \new_[61312]_ ;
  assign \new_[61323]_  = ~A169 & ~A170;
  assign \new_[61326]_  = ~A167 & ~A168;
  assign \new_[61327]_  = \new_[61326]_  & \new_[61323]_ ;
  assign \new_[61330]_  = ~A232 & A166;
  assign \new_[61333]_  = ~A234 & A233;
  assign \new_[61334]_  = \new_[61333]_  & \new_[61330]_ ;
  assign \new_[61335]_  = \new_[61334]_  & \new_[61327]_ ;
  assign \new_[61338]_  = A236 & ~A235;
  assign \new_[61341]_  = ~A266 & ~A265;
  assign \new_[61342]_  = \new_[61341]_  & \new_[61338]_ ;
  assign \new_[61345]_  = A299 & ~A298;
  assign \new_[61348]_  = A301 & A300;
  assign \new_[61349]_  = \new_[61348]_  & \new_[61345]_ ;
  assign \new_[61350]_  = \new_[61349]_  & \new_[61342]_ ;
  assign \new_[61353]_  = ~A169 & ~A170;
  assign \new_[61356]_  = ~A167 & ~A168;
  assign \new_[61357]_  = \new_[61356]_  & \new_[61353]_ ;
  assign \new_[61360]_  = ~A232 & A166;
  assign \new_[61363]_  = ~A234 & A233;
  assign \new_[61364]_  = \new_[61363]_  & \new_[61360]_ ;
  assign \new_[61365]_  = \new_[61364]_  & \new_[61357]_ ;
  assign \new_[61368]_  = A236 & ~A235;
  assign \new_[61371]_  = ~A266 & ~A265;
  assign \new_[61372]_  = \new_[61371]_  & \new_[61368]_ ;
  assign \new_[61375]_  = A299 & ~A298;
  assign \new_[61378]_  = ~A302 & A300;
  assign \new_[61379]_  = \new_[61378]_  & \new_[61375]_ ;
  assign \new_[61380]_  = \new_[61379]_  & \new_[61372]_ ;
  assign \new_[61383]_  = ~A169 & ~A170;
  assign \new_[61386]_  = ~A167 & ~A168;
  assign \new_[61387]_  = \new_[61386]_  & \new_[61383]_ ;
  assign \new_[61390]_  = A232 & A166;
  assign \new_[61393]_  = A234 & ~A233;
  assign \new_[61394]_  = \new_[61393]_  & \new_[61390]_ ;
  assign \new_[61395]_  = \new_[61394]_  & \new_[61387]_ ;
  assign \new_[61398]_  = A267 & A235;
  assign \new_[61401]_  = A269 & ~A268;
  assign \new_[61402]_  = \new_[61401]_  & \new_[61398]_ ;
  assign \new_[61405]_  = ~A299 & A298;
  assign \new_[61408]_  = A301 & A300;
  assign \new_[61409]_  = \new_[61408]_  & \new_[61405]_ ;
  assign \new_[61410]_  = \new_[61409]_  & \new_[61402]_ ;
  assign \new_[61413]_  = ~A169 & ~A170;
  assign \new_[61416]_  = ~A167 & ~A168;
  assign \new_[61417]_  = \new_[61416]_  & \new_[61413]_ ;
  assign \new_[61420]_  = A232 & A166;
  assign \new_[61423]_  = A234 & ~A233;
  assign \new_[61424]_  = \new_[61423]_  & \new_[61420]_ ;
  assign \new_[61425]_  = \new_[61424]_  & \new_[61417]_ ;
  assign \new_[61428]_  = A267 & A235;
  assign \new_[61431]_  = A269 & ~A268;
  assign \new_[61432]_  = \new_[61431]_  & \new_[61428]_ ;
  assign \new_[61435]_  = ~A299 & A298;
  assign \new_[61438]_  = ~A302 & A300;
  assign \new_[61439]_  = \new_[61438]_  & \new_[61435]_ ;
  assign \new_[61440]_  = \new_[61439]_  & \new_[61432]_ ;
  assign \new_[61443]_  = ~A169 & ~A170;
  assign \new_[61446]_  = ~A167 & ~A168;
  assign \new_[61447]_  = \new_[61446]_  & \new_[61443]_ ;
  assign \new_[61450]_  = A232 & A166;
  assign \new_[61453]_  = A234 & ~A233;
  assign \new_[61454]_  = \new_[61453]_  & \new_[61450]_ ;
  assign \new_[61455]_  = \new_[61454]_  & \new_[61447]_ ;
  assign \new_[61458]_  = A267 & A235;
  assign \new_[61461]_  = A269 & ~A268;
  assign \new_[61462]_  = \new_[61461]_  & \new_[61458]_ ;
  assign \new_[61465]_  = A299 & ~A298;
  assign \new_[61468]_  = A301 & A300;
  assign \new_[61469]_  = \new_[61468]_  & \new_[61465]_ ;
  assign \new_[61470]_  = \new_[61469]_  & \new_[61462]_ ;
  assign \new_[61473]_  = ~A169 & ~A170;
  assign \new_[61476]_  = ~A167 & ~A168;
  assign \new_[61477]_  = \new_[61476]_  & \new_[61473]_ ;
  assign \new_[61480]_  = A232 & A166;
  assign \new_[61483]_  = A234 & ~A233;
  assign \new_[61484]_  = \new_[61483]_  & \new_[61480]_ ;
  assign \new_[61485]_  = \new_[61484]_  & \new_[61477]_ ;
  assign \new_[61488]_  = A267 & A235;
  assign \new_[61491]_  = A269 & ~A268;
  assign \new_[61492]_  = \new_[61491]_  & \new_[61488]_ ;
  assign \new_[61495]_  = A299 & ~A298;
  assign \new_[61498]_  = ~A302 & A300;
  assign \new_[61499]_  = \new_[61498]_  & \new_[61495]_ ;
  assign \new_[61500]_  = \new_[61499]_  & \new_[61492]_ ;
  assign \new_[61503]_  = ~A169 & ~A170;
  assign \new_[61506]_  = ~A167 & ~A168;
  assign \new_[61507]_  = \new_[61506]_  & \new_[61503]_ ;
  assign \new_[61510]_  = A232 & A166;
  assign \new_[61513]_  = A234 & ~A233;
  assign \new_[61514]_  = \new_[61513]_  & \new_[61510]_ ;
  assign \new_[61515]_  = \new_[61514]_  & \new_[61507]_ ;
  assign \new_[61518]_  = ~A267 & A235;
  assign \new_[61521]_  = A298 & A268;
  assign \new_[61522]_  = \new_[61521]_  & \new_[61518]_ ;
  assign \new_[61525]_  = ~A300 & ~A299;
  assign \new_[61528]_  = A302 & ~A301;
  assign \new_[61529]_  = \new_[61528]_  & \new_[61525]_ ;
  assign \new_[61530]_  = \new_[61529]_  & \new_[61522]_ ;
  assign \new_[61533]_  = ~A169 & ~A170;
  assign \new_[61536]_  = ~A167 & ~A168;
  assign \new_[61537]_  = \new_[61536]_  & \new_[61533]_ ;
  assign \new_[61540]_  = A232 & A166;
  assign \new_[61543]_  = A234 & ~A233;
  assign \new_[61544]_  = \new_[61543]_  & \new_[61540]_ ;
  assign \new_[61545]_  = \new_[61544]_  & \new_[61537]_ ;
  assign \new_[61548]_  = ~A267 & A235;
  assign \new_[61551]_  = ~A298 & A268;
  assign \new_[61552]_  = \new_[61551]_  & \new_[61548]_ ;
  assign \new_[61555]_  = ~A300 & A299;
  assign \new_[61558]_  = A302 & ~A301;
  assign \new_[61559]_  = \new_[61558]_  & \new_[61555]_ ;
  assign \new_[61560]_  = \new_[61559]_  & \new_[61552]_ ;
  assign \new_[61563]_  = ~A169 & ~A170;
  assign \new_[61566]_  = ~A167 & ~A168;
  assign \new_[61567]_  = \new_[61566]_  & \new_[61563]_ ;
  assign \new_[61570]_  = A232 & A166;
  assign \new_[61573]_  = A234 & ~A233;
  assign \new_[61574]_  = \new_[61573]_  & \new_[61570]_ ;
  assign \new_[61575]_  = \new_[61574]_  & \new_[61567]_ ;
  assign \new_[61578]_  = ~A267 & A235;
  assign \new_[61581]_  = A298 & ~A269;
  assign \new_[61582]_  = \new_[61581]_  & \new_[61578]_ ;
  assign \new_[61585]_  = ~A300 & ~A299;
  assign \new_[61588]_  = A302 & ~A301;
  assign \new_[61589]_  = \new_[61588]_  & \new_[61585]_ ;
  assign \new_[61590]_  = \new_[61589]_  & \new_[61582]_ ;
  assign \new_[61593]_  = ~A169 & ~A170;
  assign \new_[61596]_  = ~A167 & ~A168;
  assign \new_[61597]_  = \new_[61596]_  & \new_[61593]_ ;
  assign \new_[61600]_  = A232 & A166;
  assign \new_[61603]_  = A234 & ~A233;
  assign \new_[61604]_  = \new_[61603]_  & \new_[61600]_ ;
  assign \new_[61605]_  = \new_[61604]_  & \new_[61597]_ ;
  assign \new_[61608]_  = ~A267 & A235;
  assign \new_[61611]_  = ~A298 & ~A269;
  assign \new_[61612]_  = \new_[61611]_  & \new_[61608]_ ;
  assign \new_[61615]_  = ~A300 & A299;
  assign \new_[61618]_  = A302 & ~A301;
  assign \new_[61619]_  = \new_[61618]_  & \new_[61615]_ ;
  assign \new_[61620]_  = \new_[61619]_  & \new_[61612]_ ;
  assign \new_[61623]_  = ~A169 & ~A170;
  assign \new_[61626]_  = ~A167 & ~A168;
  assign \new_[61627]_  = \new_[61626]_  & \new_[61623]_ ;
  assign \new_[61630]_  = A232 & A166;
  assign \new_[61633]_  = A234 & ~A233;
  assign \new_[61634]_  = \new_[61633]_  & \new_[61630]_ ;
  assign \new_[61635]_  = \new_[61634]_  & \new_[61627]_ ;
  assign \new_[61638]_  = A265 & A235;
  assign \new_[61641]_  = A298 & A266;
  assign \new_[61642]_  = \new_[61641]_  & \new_[61638]_ ;
  assign \new_[61645]_  = ~A300 & ~A299;
  assign \new_[61648]_  = A302 & ~A301;
  assign \new_[61649]_  = \new_[61648]_  & \new_[61645]_ ;
  assign \new_[61650]_  = \new_[61649]_  & \new_[61642]_ ;
  assign \new_[61653]_  = ~A169 & ~A170;
  assign \new_[61656]_  = ~A167 & ~A168;
  assign \new_[61657]_  = \new_[61656]_  & \new_[61653]_ ;
  assign \new_[61660]_  = A232 & A166;
  assign \new_[61663]_  = A234 & ~A233;
  assign \new_[61664]_  = \new_[61663]_  & \new_[61660]_ ;
  assign \new_[61665]_  = \new_[61664]_  & \new_[61657]_ ;
  assign \new_[61668]_  = A265 & A235;
  assign \new_[61671]_  = ~A298 & A266;
  assign \new_[61672]_  = \new_[61671]_  & \new_[61668]_ ;
  assign \new_[61675]_  = ~A300 & A299;
  assign \new_[61678]_  = A302 & ~A301;
  assign \new_[61679]_  = \new_[61678]_  & \new_[61675]_ ;
  assign \new_[61680]_  = \new_[61679]_  & \new_[61672]_ ;
  assign \new_[61683]_  = ~A169 & ~A170;
  assign \new_[61686]_  = ~A167 & ~A168;
  assign \new_[61687]_  = \new_[61686]_  & \new_[61683]_ ;
  assign \new_[61690]_  = A232 & A166;
  assign \new_[61693]_  = A234 & ~A233;
  assign \new_[61694]_  = \new_[61693]_  & \new_[61690]_ ;
  assign \new_[61695]_  = \new_[61694]_  & \new_[61687]_ ;
  assign \new_[61698]_  = ~A265 & A235;
  assign \new_[61701]_  = A298 & ~A266;
  assign \new_[61702]_  = \new_[61701]_  & \new_[61698]_ ;
  assign \new_[61705]_  = ~A300 & ~A299;
  assign \new_[61708]_  = A302 & ~A301;
  assign \new_[61709]_  = \new_[61708]_  & \new_[61705]_ ;
  assign \new_[61710]_  = \new_[61709]_  & \new_[61702]_ ;
  assign \new_[61713]_  = ~A169 & ~A170;
  assign \new_[61716]_  = ~A167 & ~A168;
  assign \new_[61717]_  = \new_[61716]_  & \new_[61713]_ ;
  assign \new_[61720]_  = A232 & A166;
  assign \new_[61723]_  = A234 & ~A233;
  assign \new_[61724]_  = \new_[61723]_  & \new_[61720]_ ;
  assign \new_[61725]_  = \new_[61724]_  & \new_[61717]_ ;
  assign \new_[61728]_  = ~A265 & A235;
  assign \new_[61731]_  = ~A298 & ~A266;
  assign \new_[61732]_  = \new_[61731]_  & \new_[61728]_ ;
  assign \new_[61735]_  = ~A300 & A299;
  assign \new_[61738]_  = A302 & ~A301;
  assign \new_[61739]_  = \new_[61738]_  & \new_[61735]_ ;
  assign \new_[61740]_  = \new_[61739]_  & \new_[61732]_ ;
  assign \new_[61743]_  = ~A169 & ~A170;
  assign \new_[61746]_  = ~A167 & ~A168;
  assign \new_[61747]_  = \new_[61746]_  & \new_[61743]_ ;
  assign \new_[61750]_  = A232 & A166;
  assign \new_[61753]_  = A234 & ~A233;
  assign \new_[61754]_  = \new_[61753]_  & \new_[61750]_ ;
  assign \new_[61755]_  = \new_[61754]_  & \new_[61747]_ ;
  assign \new_[61758]_  = A267 & ~A236;
  assign \new_[61761]_  = A269 & ~A268;
  assign \new_[61762]_  = \new_[61761]_  & \new_[61758]_ ;
  assign \new_[61765]_  = ~A299 & A298;
  assign \new_[61768]_  = A301 & A300;
  assign \new_[61769]_  = \new_[61768]_  & \new_[61765]_ ;
  assign \new_[61770]_  = \new_[61769]_  & \new_[61762]_ ;
  assign \new_[61773]_  = ~A169 & ~A170;
  assign \new_[61776]_  = ~A167 & ~A168;
  assign \new_[61777]_  = \new_[61776]_  & \new_[61773]_ ;
  assign \new_[61780]_  = A232 & A166;
  assign \new_[61783]_  = A234 & ~A233;
  assign \new_[61784]_  = \new_[61783]_  & \new_[61780]_ ;
  assign \new_[61785]_  = \new_[61784]_  & \new_[61777]_ ;
  assign \new_[61788]_  = A267 & ~A236;
  assign \new_[61791]_  = A269 & ~A268;
  assign \new_[61792]_  = \new_[61791]_  & \new_[61788]_ ;
  assign \new_[61795]_  = ~A299 & A298;
  assign \new_[61798]_  = ~A302 & A300;
  assign \new_[61799]_  = \new_[61798]_  & \new_[61795]_ ;
  assign \new_[61800]_  = \new_[61799]_  & \new_[61792]_ ;
  assign \new_[61803]_  = ~A169 & ~A170;
  assign \new_[61806]_  = ~A167 & ~A168;
  assign \new_[61807]_  = \new_[61806]_  & \new_[61803]_ ;
  assign \new_[61810]_  = A232 & A166;
  assign \new_[61813]_  = A234 & ~A233;
  assign \new_[61814]_  = \new_[61813]_  & \new_[61810]_ ;
  assign \new_[61815]_  = \new_[61814]_  & \new_[61807]_ ;
  assign \new_[61818]_  = A267 & ~A236;
  assign \new_[61821]_  = A269 & ~A268;
  assign \new_[61822]_  = \new_[61821]_  & \new_[61818]_ ;
  assign \new_[61825]_  = A299 & ~A298;
  assign \new_[61828]_  = A301 & A300;
  assign \new_[61829]_  = \new_[61828]_  & \new_[61825]_ ;
  assign \new_[61830]_  = \new_[61829]_  & \new_[61822]_ ;
  assign \new_[61833]_  = ~A169 & ~A170;
  assign \new_[61836]_  = ~A167 & ~A168;
  assign \new_[61837]_  = \new_[61836]_  & \new_[61833]_ ;
  assign \new_[61840]_  = A232 & A166;
  assign \new_[61843]_  = A234 & ~A233;
  assign \new_[61844]_  = \new_[61843]_  & \new_[61840]_ ;
  assign \new_[61845]_  = \new_[61844]_  & \new_[61837]_ ;
  assign \new_[61848]_  = A267 & ~A236;
  assign \new_[61851]_  = A269 & ~A268;
  assign \new_[61852]_  = \new_[61851]_  & \new_[61848]_ ;
  assign \new_[61855]_  = A299 & ~A298;
  assign \new_[61858]_  = ~A302 & A300;
  assign \new_[61859]_  = \new_[61858]_  & \new_[61855]_ ;
  assign \new_[61860]_  = \new_[61859]_  & \new_[61852]_ ;
  assign \new_[61863]_  = ~A169 & ~A170;
  assign \new_[61866]_  = ~A167 & ~A168;
  assign \new_[61867]_  = \new_[61866]_  & \new_[61863]_ ;
  assign \new_[61870]_  = A232 & A166;
  assign \new_[61873]_  = A234 & ~A233;
  assign \new_[61874]_  = \new_[61873]_  & \new_[61870]_ ;
  assign \new_[61875]_  = \new_[61874]_  & \new_[61867]_ ;
  assign \new_[61878]_  = ~A267 & ~A236;
  assign \new_[61881]_  = A298 & A268;
  assign \new_[61882]_  = \new_[61881]_  & \new_[61878]_ ;
  assign \new_[61885]_  = ~A300 & ~A299;
  assign \new_[61888]_  = A302 & ~A301;
  assign \new_[61889]_  = \new_[61888]_  & \new_[61885]_ ;
  assign \new_[61890]_  = \new_[61889]_  & \new_[61882]_ ;
  assign \new_[61893]_  = ~A169 & ~A170;
  assign \new_[61896]_  = ~A167 & ~A168;
  assign \new_[61897]_  = \new_[61896]_  & \new_[61893]_ ;
  assign \new_[61900]_  = A232 & A166;
  assign \new_[61903]_  = A234 & ~A233;
  assign \new_[61904]_  = \new_[61903]_  & \new_[61900]_ ;
  assign \new_[61905]_  = \new_[61904]_  & \new_[61897]_ ;
  assign \new_[61908]_  = ~A267 & ~A236;
  assign \new_[61911]_  = ~A298 & A268;
  assign \new_[61912]_  = \new_[61911]_  & \new_[61908]_ ;
  assign \new_[61915]_  = ~A300 & A299;
  assign \new_[61918]_  = A302 & ~A301;
  assign \new_[61919]_  = \new_[61918]_  & \new_[61915]_ ;
  assign \new_[61920]_  = \new_[61919]_  & \new_[61912]_ ;
  assign \new_[61923]_  = ~A169 & ~A170;
  assign \new_[61926]_  = ~A167 & ~A168;
  assign \new_[61927]_  = \new_[61926]_  & \new_[61923]_ ;
  assign \new_[61930]_  = A232 & A166;
  assign \new_[61933]_  = A234 & ~A233;
  assign \new_[61934]_  = \new_[61933]_  & \new_[61930]_ ;
  assign \new_[61935]_  = \new_[61934]_  & \new_[61927]_ ;
  assign \new_[61938]_  = ~A267 & ~A236;
  assign \new_[61941]_  = A298 & ~A269;
  assign \new_[61942]_  = \new_[61941]_  & \new_[61938]_ ;
  assign \new_[61945]_  = ~A300 & ~A299;
  assign \new_[61948]_  = A302 & ~A301;
  assign \new_[61949]_  = \new_[61948]_  & \new_[61945]_ ;
  assign \new_[61950]_  = \new_[61949]_  & \new_[61942]_ ;
  assign \new_[61953]_  = ~A169 & ~A170;
  assign \new_[61956]_  = ~A167 & ~A168;
  assign \new_[61957]_  = \new_[61956]_  & \new_[61953]_ ;
  assign \new_[61960]_  = A232 & A166;
  assign \new_[61963]_  = A234 & ~A233;
  assign \new_[61964]_  = \new_[61963]_  & \new_[61960]_ ;
  assign \new_[61965]_  = \new_[61964]_  & \new_[61957]_ ;
  assign \new_[61968]_  = ~A267 & ~A236;
  assign \new_[61971]_  = ~A298 & ~A269;
  assign \new_[61972]_  = \new_[61971]_  & \new_[61968]_ ;
  assign \new_[61975]_  = ~A300 & A299;
  assign \new_[61978]_  = A302 & ~A301;
  assign \new_[61979]_  = \new_[61978]_  & \new_[61975]_ ;
  assign \new_[61980]_  = \new_[61979]_  & \new_[61972]_ ;
  assign \new_[61983]_  = ~A169 & ~A170;
  assign \new_[61986]_  = ~A167 & ~A168;
  assign \new_[61987]_  = \new_[61986]_  & \new_[61983]_ ;
  assign \new_[61990]_  = A232 & A166;
  assign \new_[61993]_  = A234 & ~A233;
  assign \new_[61994]_  = \new_[61993]_  & \new_[61990]_ ;
  assign \new_[61995]_  = \new_[61994]_  & \new_[61987]_ ;
  assign \new_[61998]_  = A265 & ~A236;
  assign \new_[62001]_  = A298 & A266;
  assign \new_[62002]_  = \new_[62001]_  & \new_[61998]_ ;
  assign \new_[62005]_  = ~A300 & ~A299;
  assign \new_[62008]_  = A302 & ~A301;
  assign \new_[62009]_  = \new_[62008]_  & \new_[62005]_ ;
  assign \new_[62010]_  = \new_[62009]_  & \new_[62002]_ ;
  assign \new_[62013]_  = ~A169 & ~A170;
  assign \new_[62016]_  = ~A167 & ~A168;
  assign \new_[62017]_  = \new_[62016]_  & \new_[62013]_ ;
  assign \new_[62020]_  = A232 & A166;
  assign \new_[62023]_  = A234 & ~A233;
  assign \new_[62024]_  = \new_[62023]_  & \new_[62020]_ ;
  assign \new_[62025]_  = \new_[62024]_  & \new_[62017]_ ;
  assign \new_[62028]_  = A265 & ~A236;
  assign \new_[62031]_  = ~A298 & A266;
  assign \new_[62032]_  = \new_[62031]_  & \new_[62028]_ ;
  assign \new_[62035]_  = ~A300 & A299;
  assign \new_[62038]_  = A302 & ~A301;
  assign \new_[62039]_  = \new_[62038]_  & \new_[62035]_ ;
  assign \new_[62040]_  = \new_[62039]_  & \new_[62032]_ ;
  assign \new_[62043]_  = ~A169 & ~A170;
  assign \new_[62046]_  = ~A167 & ~A168;
  assign \new_[62047]_  = \new_[62046]_  & \new_[62043]_ ;
  assign \new_[62050]_  = A232 & A166;
  assign \new_[62053]_  = A234 & ~A233;
  assign \new_[62054]_  = \new_[62053]_  & \new_[62050]_ ;
  assign \new_[62055]_  = \new_[62054]_  & \new_[62047]_ ;
  assign \new_[62058]_  = ~A265 & ~A236;
  assign \new_[62061]_  = A298 & ~A266;
  assign \new_[62062]_  = \new_[62061]_  & \new_[62058]_ ;
  assign \new_[62065]_  = ~A300 & ~A299;
  assign \new_[62068]_  = A302 & ~A301;
  assign \new_[62069]_  = \new_[62068]_  & \new_[62065]_ ;
  assign \new_[62070]_  = \new_[62069]_  & \new_[62062]_ ;
  assign \new_[62073]_  = ~A169 & ~A170;
  assign \new_[62076]_  = ~A167 & ~A168;
  assign \new_[62077]_  = \new_[62076]_  & \new_[62073]_ ;
  assign \new_[62080]_  = A232 & A166;
  assign \new_[62083]_  = A234 & ~A233;
  assign \new_[62084]_  = \new_[62083]_  & \new_[62080]_ ;
  assign \new_[62085]_  = \new_[62084]_  & \new_[62077]_ ;
  assign \new_[62088]_  = ~A265 & ~A236;
  assign \new_[62091]_  = ~A298 & ~A266;
  assign \new_[62092]_  = \new_[62091]_  & \new_[62088]_ ;
  assign \new_[62095]_  = ~A300 & A299;
  assign \new_[62098]_  = A302 & ~A301;
  assign \new_[62099]_  = \new_[62098]_  & \new_[62095]_ ;
  assign \new_[62100]_  = \new_[62099]_  & \new_[62092]_ ;
  assign \new_[62103]_  = ~A169 & ~A170;
  assign \new_[62106]_  = ~A167 & ~A168;
  assign \new_[62107]_  = \new_[62106]_  & \new_[62103]_ ;
  assign \new_[62110]_  = A232 & A166;
  assign \new_[62113]_  = ~A234 & ~A233;
  assign \new_[62114]_  = \new_[62113]_  & \new_[62110]_ ;
  assign \new_[62115]_  = \new_[62114]_  & \new_[62107]_ ;
  assign \new_[62118]_  = A236 & ~A235;
  assign \new_[62121]_  = A268 & ~A267;
  assign \new_[62122]_  = \new_[62121]_  & \new_[62118]_ ;
  assign \new_[62125]_  = ~A299 & A298;
  assign \new_[62128]_  = A301 & A300;
  assign \new_[62129]_  = \new_[62128]_  & \new_[62125]_ ;
  assign \new_[62130]_  = \new_[62129]_  & \new_[62122]_ ;
  assign \new_[62133]_  = ~A169 & ~A170;
  assign \new_[62136]_  = ~A167 & ~A168;
  assign \new_[62137]_  = \new_[62136]_  & \new_[62133]_ ;
  assign \new_[62140]_  = A232 & A166;
  assign \new_[62143]_  = ~A234 & ~A233;
  assign \new_[62144]_  = \new_[62143]_  & \new_[62140]_ ;
  assign \new_[62145]_  = \new_[62144]_  & \new_[62137]_ ;
  assign \new_[62148]_  = A236 & ~A235;
  assign \new_[62151]_  = A268 & ~A267;
  assign \new_[62152]_  = \new_[62151]_  & \new_[62148]_ ;
  assign \new_[62155]_  = ~A299 & A298;
  assign \new_[62158]_  = ~A302 & A300;
  assign \new_[62159]_  = \new_[62158]_  & \new_[62155]_ ;
  assign \new_[62160]_  = \new_[62159]_  & \new_[62152]_ ;
  assign \new_[62163]_  = ~A169 & ~A170;
  assign \new_[62166]_  = ~A167 & ~A168;
  assign \new_[62167]_  = \new_[62166]_  & \new_[62163]_ ;
  assign \new_[62170]_  = A232 & A166;
  assign \new_[62173]_  = ~A234 & ~A233;
  assign \new_[62174]_  = \new_[62173]_  & \new_[62170]_ ;
  assign \new_[62175]_  = \new_[62174]_  & \new_[62167]_ ;
  assign \new_[62178]_  = A236 & ~A235;
  assign \new_[62181]_  = A268 & ~A267;
  assign \new_[62182]_  = \new_[62181]_  & \new_[62178]_ ;
  assign \new_[62185]_  = A299 & ~A298;
  assign \new_[62188]_  = A301 & A300;
  assign \new_[62189]_  = \new_[62188]_  & \new_[62185]_ ;
  assign \new_[62190]_  = \new_[62189]_  & \new_[62182]_ ;
  assign \new_[62193]_  = ~A169 & ~A170;
  assign \new_[62196]_  = ~A167 & ~A168;
  assign \new_[62197]_  = \new_[62196]_  & \new_[62193]_ ;
  assign \new_[62200]_  = A232 & A166;
  assign \new_[62203]_  = ~A234 & ~A233;
  assign \new_[62204]_  = \new_[62203]_  & \new_[62200]_ ;
  assign \new_[62205]_  = \new_[62204]_  & \new_[62197]_ ;
  assign \new_[62208]_  = A236 & ~A235;
  assign \new_[62211]_  = A268 & ~A267;
  assign \new_[62212]_  = \new_[62211]_  & \new_[62208]_ ;
  assign \new_[62215]_  = A299 & ~A298;
  assign \new_[62218]_  = ~A302 & A300;
  assign \new_[62219]_  = \new_[62218]_  & \new_[62215]_ ;
  assign \new_[62220]_  = \new_[62219]_  & \new_[62212]_ ;
  assign \new_[62223]_  = ~A169 & ~A170;
  assign \new_[62226]_  = ~A167 & ~A168;
  assign \new_[62227]_  = \new_[62226]_  & \new_[62223]_ ;
  assign \new_[62230]_  = A232 & A166;
  assign \new_[62233]_  = ~A234 & ~A233;
  assign \new_[62234]_  = \new_[62233]_  & \new_[62230]_ ;
  assign \new_[62235]_  = \new_[62234]_  & \new_[62227]_ ;
  assign \new_[62238]_  = A236 & ~A235;
  assign \new_[62241]_  = ~A269 & ~A267;
  assign \new_[62242]_  = \new_[62241]_  & \new_[62238]_ ;
  assign \new_[62245]_  = ~A299 & A298;
  assign \new_[62248]_  = A301 & A300;
  assign \new_[62249]_  = \new_[62248]_  & \new_[62245]_ ;
  assign \new_[62250]_  = \new_[62249]_  & \new_[62242]_ ;
  assign \new_[62253]_  = ~A169 & ~A170;
  assign \new_[62256]_  = ~A167 & ~A168;
  assign \new_[62257]_  = \new_[62256]_  & \new_[62253]_ ;
  assign \new_[62260]_  = A232 & A166;
  assign \new_[62263]_  = ~A234 & ~A233;
  assign \new_[62264]_  = \new_[62263]_  & \new_[62260]_ ;
  assign \new_[62265]_  = \new_[62264]_  & \new_[62257]_ ;
  assign \new_[62268]_  = A236 & ~A235;
  assign \new_[62271]_  = ~A269 & ~A267;
  assign \new_[62272]_  = \new_[62271]_  & \new_[62268]_ ;
  assign \new_[62275]_  = ~A299 & A298;
  assign \new_[62278]_  = ~A302 & A300;
  assign \new_[62279]_  = \new_[62278]_  & \new_[62275]_ ;
  assign \new_[62280]_  = \new_[62279]_  & \new_[62272]_ ;
  assign \new_[62283]_  = ~A169 & ~A170;
  assign \new_[62286]_  = ~A167 & ~A168;
  assign \new_[62287]_  = \new_[62286]_  & \new_[62283]_ ;
  assign \new_[62290]_  = A232 & A166;
  assign \new_[62293]_  = ~A234 & ~A233;
  assign \new_[62294]_  = \new_[62293]_  & \new_[62290]_ ;
  assign \new_[62295]_  = \new_[62294]_  & \new_[62287]_ ;
  assign \new_[62298]_  = A236 & ~A235;
  assign \new_[62301]_  = ~A269 & ~A267;
  assign \new_[62302]_  = \new_[62301]_  & \new_[62298]_ ;
  assign \new_[62305]_  = A299 & ~A298;
  assign \new_[62308]_  = A301 & A300;
  assign \new_[62309]_  = \new_[62308]_  & \new_[62305]_ ;
  assign \new_[62310]_  = \new_[62309]_  & \new_[62302]_ ;
  assign \new_[62313]_  = ~A169 & ~A170;
  assign \new_[62316]_  = ~A167 & ~A168;
  assign \new_[62317]_  = \new_[62316]_  & \new_[62313]_ ;
  assign \new_[62320]_  = A232 & A166;
  assign \new_[62323]_  = ~A234 & ~A233;
  assign \new_[62324]_  = \new_[62323]_  & \new_[62320]_ ;
  assign \new_[62325]_  = \new_[62324]_  & \new_[62317]_ ;
  assign \new_[62328]_  = A236 & ~A235;
  assign \new_[62331]_  = ~A269 & ~A267;
  assign \new_[62332]_  = \new_[62331]_  & \new_[62328]_ ;
  assign \new_[62335]_  = A299 & ~A298;
  assign \new_[62338]_  = ~A302 & A300;
  assign \new_[62339]_  = \new_[62338]_  & \new_[62335]_ ;
  assign \new_[62340]_  = \new_[62339]_  & \new_[62332]_ ;
  assign \new_[62343]_  = ~A169 & ~A170;
  assign \new_[62346]_  = ~A167 & ~A168;
  assign \new_[62347]_  = \new_[62346]_  & \new_[62343]_ ;
  assign \new_[62350]_  = A232 & A166;
  assign \new_[62353]_  = ~A234 & ~A233;
  assign \new_[62354]_  = \new_[62353]_  & \new_[62350]_ ;
  assign \new_[62355]_  = \new_[62354]_  & \new_[62347]_ ;
  assign \new_[62358]_  = A236 & ~A235;
  assign \new_[62361]_  = A266 & A265;
  assign \new_[62362]_  = \new_[62361]_  & \new_[62358]_ ;
  assign \new_[62365]_  = ~A299 & A298;
  assign \new_[62368]_  = A301 & A300;
  assign \new_[62369]_  = \new_[62368]_  & \new_[62365]_ ;
  assign \new_[62370]_  = \new_[62369]_  & \new_[62362]_ ;
  assign \new_[62373]_  = ~A169 & ~A170;
  assign \new_[62376]_  = ~A167 & ~A168;
  assign \new_[62377]_  = \new_[62376]_  & \new_[62373]_ ;
  assign \new_[62380]_  = A232 & A166;
  assign \new_[62383]_  = ~A234 & ~A233;
  assign \new_[62384]_  = \new_[62383]_  & \new_[62380]_ ;
  assign \new_[62385]_  = \new_[62384]_  & \new_[62377]_ ;
  assign \new_[62388]_  = A236 & ~A235;
  assign \new_[62391]_  = A266 & A265;
  assign \new_[62392]_  = \new_[62391]_  & \new_[62388]_ ;
  assign \new_[62395]_  = ~A299 & A298;
  assign \new_[62398]_  = ~A302 & A300;
  assign \new_[62399]_  = \new_[62398]_  & \new_[62395]_ ;
  assign \new_[62400]_  = \new_[62399]_  & \new_[62392]_ ;
  assign \new_[62403]_  = ~A169 & ~A170;
  assign \new_[62406]_  = ~A167 & ~A168;
  assign \new_[62407]_  = \new_[62406]_  & \new_[62403]_ ;
  assign \new_[62410]_  = A232 & A166;
  assign \new_[62413]_  = ~A234 & ~A233;
  assign \new_[62414]_  = \new_[62413]_  & \new_[62410]_ ;
  assign \new_[62415]_  = \new_[62414]_  & \new_[62407]_ ;
  assign \new_[62418]_  = A236 & ~A235;
  assign \new_[62421]_  = A266 & A265;
  assign \new_[62422]_  = \new_[62421]_  & \new_[62418]_ ;
  assign \new_[62425]_  = A299 & ~A298;
  assign \new_[62428]_  = A301 & A300;
  assign \new_[62429]_  = \new_[62428]_  & \new_[62425]_ ;
  assign \new_[62430]_  = \new_[62429]_  & \new_[62422]_ ;
  assign \new_[62433]_  = ~A169 & ~A170;
  assign \new_[62436]_  = ~A167 & ~A168;
  assign \new_[62437]_  = \new_[62436]_  & \new_[62433]_ ;
  assign \new_[62440]_  = A232 & A166;
  assign \new_[62443]_  = ~A234 & ~A233;
  assign \new_[62444]_  = \new_[62443]_  & \new_[62440]_ ;
  assign \new_[62445]_  = \new_[62444]_  & \new_[62437]_ ;
  assign \new_[62448]_  = A236 & ~A235;
  assign \new_[62451]_  = A266 & A265;
  assign \new_[62452]_  = \new_[62451]_  & \new_[62448]_ ;
  assign \new_[62455]_  = A299 & ~A298;
  assign \new_[62458]_  = ~A302 & A300;
  assign \new_[62459]_  = \new_[62458]_  & \new_[62455]_ ;
  assign \new_[62460]_  = \new_[62459]_  & \new_[62452]_ ;
  assign \new_[62463]_  = ~A169 & ~A170;
  assign \new_[62466]_  = ~A167 & ~A168;
  assign \new_[62467]_  = \new_[62466]_  & \new_[62463]_ ;
  assign \new_[62470]_  = A232 & A166;
  assign \new_[62473]_  = ~A234 & ~A233;
  assign \new_[62474]_  = \new_[62473]_  & \new_[62470]_ ;
  assign \new_[62475]_  = \new_[62474]_  & \new_[62467]_ ;
  assign \new_[62478]_  = A236 & ~A235;
  assign \new_[62481]_  = ~A266 & ~A265;
  assign \new_[62482]_  = \new_[62481]_  & \new_[62478]_ ;
  assign \new_[62485]_  = ~A299 & A298;
  assign \new_[62488]_  = A301 & A300;
  assign \new_[62489]_  = \new_[62488]_  & \new_[62485]_ ;
  assign \new_[62490]_  = \new_[62489]_  & \new_[62482]_ ;
  assign \new_[62493]_  = ~A169 & ~A170;
  assign \new_[62496]_  = ~A167 & ~A168;
  assign \new_[62497]_  = \new_[62496]_  & \new_[62493]_ ;
  assign \new_[62500]_  = A232 & A166;
  assign \new_[62503]_  = ~A234 & ~A233;
  assign \new_[62504]_  = \new_[62503]_  & \new_[62500]_ ;
  assign \new_[62505]_  = \new_[62504]_  & \new_[62497]_ ;
  assign \new_[62508]_  = A236 & ~A235;
  assign \new_[62511]_  = ~A266 & ~A265;
  assign \new_[62512]_  = \new_[62511]_  & \new_[62508]_ ;
  assign \new_[62515]_  = ~A299 & A298;
  assign \new_[62518]_  = ~A302 & A300;
  assign \new_[62519]_  = \new_[62518]_  & \new_[62515]_ ;
  assign \new_[62520]_  = \new_[62519]_  & \new_[62512]_ ;
  assign \new_[62523]_  = ~A169 & ~A170;
  assign \new_[62526]_  = ~A167 & ~A168;
  assign \new_[62527]_  = \new_[62526]_  & \new_[62523]_ ;
  assign \new_[62530]_  = A232 & A166;
  assign \new_[62533]_  = ~A234 & ~A233;
  assign \new_[62534]_  = \new_[62533]_  & \new_[62530]_ ;
  assign \new_[62535]_  = \new_[62534]_  & \new_[62527]_ ;
  assign \new_[62538]_  = A236 & ~A235;
  assign \new_[62541]_  = ~A266 & ~A265;
  assign \new_[62542]_  = \new_[62541]_  & \new_[62538]_ ;
  assign \new_[62545]_  = A299 & ~A298;
  assign \new_[62548]_  = A301 & A300;
  assign \new_[62549]_  = \new_[62548]_  & \new_[62545]_ ;
  assign \new_[62550]_  = \new_[62549]_  & \new_[62542]_ ;
  assign \new_[62553]_  = ~A169 & ~A170;
  assign \new_[62556]_  = ~A167 & ~A168;
  assign \new_[62557]_  = \new_[62556]_  & \new_[62553]_ ;
  assign \new_[62560]_  = A232 & A166;
  assign \new_[62563]_  = ~A234 & ~A233;
  assign \new_[62564]_  = \new_[62563]_  & \new_[62560]_ ;
  assign \new_[62565]_  = \new_[62564]_  & \new_[62557]_ ;
  assign \new_[62568]_  = A236 & ~A235;
  assign \new_[62571]_  = ~A266 & ~A265;
  assign \new_[62572]_  = \new_[62571]_  & \new_[62568]_ ;
  assign \new_[62575]_  = A299 & ~A298;
  assign \new_[62578]_  = ~A302 & A300;
  assign \new_[62579]_  = \new_[62578]_  & \new_[62575]_ ;
  assign \new_[62580]_  = \new_[62579]_  & \new_[62572]_ ;
  assign \new_[62583]_  = A200 & ~A199;
  assign \new_[62586]_  = A202 & A201;
  assign \new_[62587]_  = \new_[62586]_  & \new_[62583]_ ;
  assign \new_[62590]_  = A233 & ~A232;
  assign \new_[62593]_  = ~A235 & ~A234;
  assign \new_[62594]_  = \new_[62593]_  & \new_[62590]_ ;
  assign \new_[62595]_  = \new_[62594]_  & \new_[62587]_ ;
  assign \new_[62598]_  = A267 & A236;
  assign \new_[62601]_  = A269 & ~A268;
  assign \new_[62602]_  = \new_[62601]_  & \new_[62598]_ ;
  assign \new_[62605]_  = ~A299 & A298;
  assign \new_[62609]_  = A302 & ~A301;
  assign \new_[62610]_  = ~A300 & \new_[62609]_ ;
  assign \new_[62611]_  = \new_[62610]_  & \new_[62605]_ ;
  assign \new_[62612]_  = \new_[62611]_  & \new_[62602]_ ;
  assign \new_[62615]_  = A200 & ~A199;
  assign \new_[62618]_  = A202 & A201;
  assign \new_[62619]_  = \new_[62618]_  & \new_[62615]_ ;
  assign \new_[62622]_  = A233 & ~A232;
  assign \new_[62625]_  = ~A235 & ~A234;
  assign \new_[62626]_  = \new_[62625]_  & \new_[62622]_ ;
  assign \new_[62627]_  = \new_[62626]_  & \new_[62619]_ ;
  assign \new_[62630]_  = A267 & A236;
  assign \new_[62633]_  = A269 & ~A268;
  assign \new_[62634]_  = \new_[62633]_  & \new_[62630]_ ;
  assign \new_[62637]_  = A299 & ~A298;
  assign \new_[62641]_  = A302 & ~A301;
  assign \new_[62642]_  = ~A300 & \new_[62641]_ ;
  assign \new_[62643]_  = \new_[62642]_  & \new_[62637]_ ;
  assign \new_[62644]_  = \new_[62643]_  & \new_[62634]_ ;
  assign \new_[62647]_  = A200 & ~A199;
  assign \new_[62650]_  = A202 & A201;
  assign \new_[62651]_  = \new_[62650]_  & \new_[62647]_ ;
  assign \new_[62654]_  = ~A233 & A232;
  assign \new_[62657]_  = ~A235 & ~A234;
  assign \new_[62658]_  = \new_[62657]_  & \new_[62654]_ ;
  assign \new_[62659]_  = \new_[62658]_  & \new_[62651]_ ;
  assign \new_[62662]_  = A267 & A236;
  assign \new_[62665]_  = A269 & ~A268;
  assign \new_[62666]_  = \new_[62665]_  & \new_[62662]_ ;
  assign \new_[62669]_  = ~A299 & A298;
  assign \new_[62673]_  = A302 & ~A301;
  assign \new_[62674]_  = ~A300 & \new_[62673]_ ;
  assign \new_[62675]_  = \new_[62674]_  & \new_[62669]_ ;
  assign \new_[62676]_  = \new_[62675]_  & \new_[62666]_ ;
  assign \new_[62679]_  = A200 & ~A199;
  assign \new_[62682]_  = A202 & A201;
  assign \new_[62683]_  = \new_[62682]_  & \new_[62679]_ ;
  assign \new_[62686]_  = ~A233 & A232;
  assign \new_[62689]_  = ~A235 & ~A234;
  assign \new_[62690]_  = \new_[62689]_  & \new_[62686]_ ;
  assign \new_[62691]_  = \new_[62690]_  & \new_[62683]_ ;
  assign \new_[62694]_  = A267 & A236;
  assign \new_[62697]_  = A269 & ~A268;
  assign \new_[62698]_  = \new_[62697]_  & \new_[62694]_ ;
  assign \new_[62701]_  = A299 & ~A298;
  assign \new_[62705]_  = A302 & ~A301;
  assign \new_[62706]_  = ~A300 & \new_[62705]_ ;
  assign \new_[62707]_  = \new_[62706]_  & \new_[62701]_ ;
  assign \new_[62708]_  = \new_[62707]_  & \new_[62698]_ ;
  assign \new_[62711]_  = A200 & ~A199;
  assign \new_[62714]_  = ~A203 & A201;
  assign \new_[62715]_  = \new_[62714]_  & \new_[62711]_ ;
  assign \new_[62718]_  = A233 & ~A232;
  assign \new_[62721]_  = ~A235 & ~A234;
  assign \new_[62722]_  = \new_[62721]_  & \new_[62718]_ ;
  assign \new_[62723]_  = \new_[62722]_  & \new_[62715]_ ;
  assign \new_[62726]_  = A267 & A236;
  assign \new_[62729]_  = A269 & ~A268;
  assign \new_[62730]_  = \new_[62729]_  & \new_[62726]_ ;
  assign \new_[62733]_  = ~A299 & A298;
  assign \new_[62737]_  = A302 & ~A301;
  assign \new_[62738]_  = ~A300 & \new_[62737]_ ;
  assign \new_[62739]_  = \new_[62738]_  & \new_[62733]_ ;
  assign \new_[62740]_  = \new_[62739]_  & \new_[62730]_ ;
  assign \new_[62743]_  = A200 & ~A199;
  assign \new_[62746]_  = ~A203 & A201;
  assign \new_[62747]_  = \new_[62746]_  & \new_[62743]_ ;
  assign \new_[62750]_  = A233 & ~A232;
  assign \new_[62753]_  = ~A235 & ~A234;
  assign \new_[62754]_  = \new_[62753]_  & \new_[62750]_ ;
  assign \new_[62755]_  = \new_[62754]_  & \new_[62747]_ ;
  assign \new_[62758]_  = A267 & A236;
  assign \new_[62761]_  = A269 & ~A268;
  assign \new_[62762]_  = \new_[62761]_  & \new_[62758]_ ;
  assign \new_[62765]_  = A299 & ~A298;
  assign \new_[62769]_  = A302 & ~A301;
  assign \new_[62770]_  = ~A300 & \new_[62769]_ ;
  assign \new_[62771]_  = \new_[62770]_  & \new_[62765]_ ;
  assign \new_[62772]_  = \new_[62771]_  & \new_[62762]_ ;
  assign \new_[62775]_  = A200 & ~A199;
  assign \new_[62778]_  = ~A203 & A201;
  assign \new_[62779]_  = \new_[62778]_  & \new_[62775]_ ;
  assign \new_[62782]_  = ~A233 & A232;
  assign \new_[62785]_  = ~A235 & ~A234;
  assign \new_[62786]_  = \new_[62785]_  & \new_[62782]_ ;
  assign \new_[62787]_  = \new_[62786]_  & \new_[62779]_ ;
  assign \new_[62790]_  = A267 & A236;
  assign \new_[62793]_  = A269 & ~A268;
  assign \new_[62794]_  = \new_[62793]_  & \new_[62790]_ ;
  assign \new_[62797]_  = ~A299 & A298;
  assign \new_[62801]_  = A302 & ~A301;
  assign \new_[62802]_  = ~A300 & \new_[62801]_ ;
  assign \new_[62803]_  = \new_[62802]_  & \new_[62797]_ ;
  assign \new_[62804]_  = \new_[62803]_  & \new_[62794]_ ;
  assign \new_[62807]_  = A200 & ~A199;
  assign \new_[62810]_  = ~A203 & A201;
  assign \new_[62811]_  = \new_[62810]_  & \new_[62807]_ ;
  assign \new_[62814]_  = ~A233 & A232;
  assign \new_[62817]_  = ~A235 & ~A234;
  assign \new_[62818]_  = \new_[62817]_  & \new_[62814]_ ;
  assign \new_[62819]_  = \new_[62818]_  & \new_[62811]_ ;
  assign \new_[62822]_  = A267 & A236;
  assign \new_[62825]_  = A269 & ~A268;
  assign \new_[62826]_  = \new_[62825]_  & \new_[62822]_ ;
  assign \new_[62829]_  = A299 & ~A298;
  assign \new_[62833]_  = A302 & ~A301;
  assign \new_[62834]_  = ~A300 & \new_[62833]_ ;
  assign \new_[62835]_  = \new_[62834]_  & \new_[62829]_ ;
  assign \new_[62836]_  = \new_[62835]_  & \new_[62826]_ ;
  assign \new_[62839]_  = A200 & ~A199;
  assign \new_[62842]_  = ~A202 & ~A201;
  assign \new_[62843]_  = \new_[62842]_  & \new_[62839]_ ;
  assign \new_[62846]_  = ~A232 & A203;
  assign \new_[62849]_  = A234 & A233;
  assign \new_[62850]_  = \new_[62849]_  & \new_[62846]_ ;
  assign \new_[62851]_  = \new_[62850]_  & \new_[62843]_ ;
  assign \new_[62854]_  = A267 & A235;
  assign \new_[62857]_  = A269 & ~A268;
  assign \new_[62858]_  = \new_[62857]_  & \new_[62854]_ ;
  assign \new_[62861]_  = ~A299 & A298;
  assign \new_[62865]_  = A302 & ~A301;
  assign \new_[62866]_  = ~A300 & \new_[62865]_ ;
  assign \new_[62867]_  = \new_[62866]_  & \new_[62861]_ ;
  assign \new_[62868]_  = \new_[62867]_  & \new_[62858]_ ;
  assign \new_[62871]_  = A200 & ~A199;
  assign \new_[62874]_  = ~A202 & ~A201;
  assign \new_[62875]_  = \new_[62874]_  & \new_[62871]_ ;
  assign \new_[62878]_  = ~A232 & A203;
  assign \new_[62881]_  = A234 & A233;
  assign \new_[62882]_  = \new_[62881]_  & \new_[62878]_ ;
  assign \new_[62883]_  = \new_[62882]_  & \new_[62875]_ ;
  assign \new_[62886]_  = A267 & A235;
  assign \new_[62889]_  = A269 & ~A268;
  assign \new_[62890]_  = \new_[62889]_  & \new_[62886]_ ;
  assign \new_[62893]_  = A299 & ~A298;
  assign \new_[62897]_  = A302 & ~A301;
  assign \new_[62898]_  = ~A300 & \new_[62897]_ ;
  assign \new_[62899]_  = \new_[62898]_  & \new_[62893]_ ;
  assign \new_[62900]_  = \new_[62899]_  & \new_[62890]_ ;
  assign \new_[62903]_  = A200 & ~A199;
  assign \new_[62906]_  = ~A202 & ~A201;
  assign \new_[62907]_  = \new_[62906]_  & \new_[62903]_ ;
  assign \new_[62910]_  = ~A232 & A203;
  assign \new_[62913]_  = A234 & A233;
  assign \new_[62914]_  = \new_[62913]_  & \new_[62910]_ ;
  assign \new_[62915]_  = \new_[62914]_  & \new_[62907]_ ;
  assign \new_[62918]_  = A267 & ~A236;
  assign \new_[62921]_  = A269 & ~A268;
  assign \new_[62922]_  = \new_[62921]_  & \new_[62918]_ ;
  assign \new_[62925]_  = ~A299 & A298;
  assign \new_[62929]_  = A302 & ~A301;
  assign \new_[62930]_  = ~A300 & \new_[62929]_ ;
  assign \new_[62931]_  = \new_[62930]_  & \new_[62925]_ ;
  assign \new_[62932]_  = \new_[62931]_  & \new_[62922]_ ;
  assign \new_[62935]_  = A200 & ~A199;
  assign \new_[62938]_  = ~A202 & ~A201;
  assign \new_[62939]_  = \new_[62938]_  & \new_[62935]_ ;
  assign \new_[62942]_  = ~A232 & A203;
  assign \new_[62945]_  = A234 & A233;
  assign \new_[62946]_  = \new_[62945]_  & \new_[62942]_ ;
  assign \new_[62947]_  = \new_[62946]_  & \new_[62939]_ ;
  assign \new_[62950]_  = A267 & ~A236;
  assign \new_[62953]_  = A269 & ~A268;
  assign \new_[62954]_  = \new_[62953]_  & \new_[62950]_ ;
  assign \new_[62957]_  = A299 & ~A298;
  assign \new_[62961]_  = A302 & ~A301;
  assign \new_[62962]_  = ~A300 & \new_[62961]_ ;
  assign \new_[62963]_  = \new_[62962]_  & \new_[62957]_ ;
  assign \new_[62964]_  = \new_[62963]_  & \new_[62954]_ ;
  assign \new_[62967]_  = A200 & ~A199;
  assign \new_[62970]_  = ~A202 & ~A201;
  assign \new_[62971]_  = \new_[62970]_  & \new_[62967]_ ;
  assign \new_[62974]_  = ~A232 & A203;
  assign \new_[62977]_  = ~A234 & A233;
  assign \new_[62978]_  = \new_[62977]_  & \new_[62974]_ ;
  assign \new_[62979]_  = \new_[62978]_  & \new_[62971]_ ;
  assign \new_[62982]_  = A236 & ~A235;
  assign \new_[62985]_  = ~A268 & A267;
  assign \new_[62986]_  = \new_[62985]_  & \new_[62982]_ ;
  assign \new_[62989]_  = A298 & A269;
  assign \new_[62993]_  = A301 & A300;
  assign \new_[62994]_  = ~A299 & \new_[62993]_ ;
  assign \new_[62995]_  = \new_[62994]_  & \new_[62989]_ ;
  assign \new_[62996]_  = \new_[62995]_  & \new_[62986]_ ;
  assign \new_[62999]_  = A200 & ~A199;
  assign \new_[63002]_  = ~A202 & ~A201;
  assign \new_[63003]_  = \new_[63002]_  & \new_[62999]_ ;
  assign \new_[63006]_  = ~A232 & A203;
  assign \new_[63009]_  = ~A234 & A233;
  assign \new_[63010]_  = \new_[63009]_  & \new_[63006]_ ;
  assign \new_[63011]_  = \new_[63010]_  & \new_[63003]_ ;
  assign \new_[63014]_  = A236 & ~A235;
  assign \new_[63017]_  = ~A268 & A267;
  assign \new_[63018]_  = \new_[63017]_  & \new_[63014]_ ;
  assign \new_[63021]_  = A298 & A269;
  assign \new_[63025]_  = ~A302 & A300;
  assign \new_[63026]_  = ~A299 & \new_[63025]_ ;
  assign \new_[63027]_  = \new_[63026]_  & \new_[63021]_ ;
  assign \new_[63028]_  = \new_[63027]_  & \new_[63018]_ ;
  assign \new_[63031]_  = A200 & ~A199;
  assign \new_[63034]_  = ~A202 & ~A201;
  assign \new_[63035]_  = \new_[63034]_  & \new_[63031]_ ;
  assign \new_[63038]_  = ~A232 & A203;
  assign \new_[63041]_  = ~A234 & A233;
  assign \new_[63042]_  = \new_[63041]_  & \new_[63038]_ ;
  assign \new_[63043]_  = \new_[63042]_  & \new_[63035]_ ;
  assign \new_[63046]_  = A236 & ~A235;
  assign \new_[63049]_  = ~A268 & A267;
  assign \new_[63050]_  = \new_[63049]_  & \new_[63046]_ ;
  assign \new_[63053]_  = ~A298 & A269;
  assign \new_[63057]_  = A301 & A300;
  assign \new_[63058]_  = A299 & \new_[63057]_ ;
  assign \new_[63059]_  = \new_[63058]_  & \new_[63053]_ ;
  assign \new_[63060]_  = \new_[63059]_  & \new_[63050]_ ;
  assign \new_[63063]_  = A200 & ~A199;
  assign \new_[63066]_  = ~A202 & ~A201;
  assign \new_[63067]_  = \new_[63066]_  & \new_[63063]_ ;
  assign \new_[63070]_  = ~A232 & A203;
  assign \new_[63073]_  = ~A234 & A233;
  assign \new_[63074]_  = \new_[63073]_  & \new_[63070]_ ;
  assign \new_[63075]_  = \new_[63074]_  & \new_[63067]_ ;
  assign \new_[63078]_  = A236 & ~A235;
  assign \new_[63081]_  = ~A268 & A267;
  assign \new_[63082]_  = \new_[63081]_  & \new_[63078]_ ;
  assign \new_[63085]_  = ~A298 & A269;
  assign \new_[63089]_  = ~A302 & A300;
  assign \new_[63090]_  = A299 & \new_[63089]_ ;
  assign \new_[63091]_  = \new_[63090]_  & \new_[63085]_ ;
  assign \new_[63092]_  = \new_[63091]_  & \new_[63082]_ ;
  assign \new_[63095]_  = A200 & ~A199;
  assign \new_[63098]_  = ~A202 & ~A201;
  assign \new_[63099]_  = \new_[63098]_  & \new_[63095]_ ;
  assign \new_[63102]_  = ~A232 & A203;
  assign \new_[63105]_  = ~A234 & A233;
  assign \new_[63106]_  = \new_[63105]_  & \new_[63102]_ ;
  assign \new_[63107]_  = \new_[63106]_  & \new_[63099]_ ;
  assign \new_[63110]_  = A236 & ~A235;
  assign \new_[63113]_  = A268 & ~A267;
  assign \new_[63114]_  = \new_[63113]_  & \new_[63110]_ ;
  assign \new_[63117]_  = ~A299 & A298;
  assign \new_[63121]_  = A302 & ~A301;
  assign \new_[63122]_  = ~A300 & \new_[63121]_ ;
  assign \new_[63123]_  = \new_[63122]_  & \new_[63117]_ ;
  assign \new_[63124]_  = \new_[63123]_  & \new_[63114]_ ;
  assign \new_[63127]_  = A200 & ~A199;
  assign \new_[63130]_  = ~A202 & ~A201;
  assign \new_[63131]_  = \new_[63130]_  & \new_[63127]_ ;
  assign \new_[63134]_  = ~A232 & A203;
  assign \new_[63137]_  = ~A234 & A233;
  assign \new_[63138]_  = \new_[63137]_  & \new_[63134]_ ;
  assign \new_[63139]_  = \new_[63138]_  & \new_[63131]_ ;
  assign \new_[63142]_  = A236 & ~A235;
  assign \new_[63145]_  = A268 & ~A267;
  assign \new_[63146]_  = \new_[63145]_  & \new_[63142]_ ;
  assign \new_[63149]_  = A299 & ~A298;
  assign \new_[63153]_  = A302 & ~A301;
  assign \new_[63154]_  = ~A300 & \new_[63153]_ ;
  assign \new_[63155]_  = \new_[63154]_  & \new_[63149]_ ;
  assign \new_[63156]_  = \new_[63155]_  & \new_[63146]_ ;
  assign \new_[63159]_  = A200 & ~A199;
  assign \new_[63162]_  = ~A202 & ~A201;
  assign \new_[63163]_  = \new_[63162]_  & \new_[63159]_ ;
  assign \new_[63166]_  = ~A232 & A203;
  assign \new_[63169]_  = ~A234 & A233;
  assign \new_[63170]_  = \new_[63169]_  & \new_[63166]_ ;
  assign \new_[63171]_  = \new_[63170]_  & \new_[63163]_ ;
  assign \new_[63174]_  = A236 & ~A235;
  assign \new_[63177]_  = ~A269 & ~A267;
  assign \new_[63178]_  = \new_[63177]_  & \new_[63174]_ ;
  assign \new_[63181]_  = ~A299 & A298;
  assign \new_[63185]_  = A302 & ~A301;
  assign \new_[63186]_  = ~A300 & \new_[63185]_ ;
  assign \new_[63187]_  = \new_[63186]_  & \new_[63181]_ ;
  assign \new_[63188]_  = \new_[63187]_  & \new_[63178]_ ;
  assign \new_[63191]_  = A200 & ~A199;
  assign \new_[63194]_  = ~A202 & ~A201;
  assign \new_[63195]_  = \new_[63194]_  & \new_[63191]_ ;
  assign \new_[63198]_  = ~A232 & A203;
  assign \new_[63201]_  = ~A234 & A233;
  assign \new_[63202]_  = \new_[63201]_  & \new_[63198]_ ;
  assign \new_[63203]_  = \new_[63202]_  & \new_[63195]_ ;
  assign \new_[63206]_  = A236 & ~A235;
  assign \new_[63209]_  = ~A269 & ~A267;
  assign \new_[63210]_  = \new_[63209]_  & \new_[63206]_ ;
  assign \new_[63213]_  = A299 & ~A298;
  assign \new_[63217]_  = A302 & ~A301;
  assign \new_[63218]_  = ~A300 & \new_[63217]_ ;
  assign \new_[63219]_  = \new_[63218]_  & \new_[63213]_ ;
  assign \new_[63220]_  = \new_[63219]_  & \new_[63210]_ ;
  assign \new_[63223]_  = A200 & ~A199;
  assign \new_[63226]_  = ~A202 & ~A201;
  assign \new_[63227]_  = \new_[63226]_  & \new_[63223]_ ;
  assign \new_[63230]_  = ~A232 & A203;
  assign \new_[63233]_  = ~A234 & A233;
  assign \new_[63234]_  = \new_[63233]_  & \new_[63230]_ ;
  assign \new_[63235]_  = \new_[63234]_  & \new_[63227]_ ;
  assign \new_[63238]_  = A236 & ~A235;
  assign \new_[63241]_  = A266 & A265;
  assign \new_[63242]_  = \new_[63241]_  & \new_[63238]_ ;
  assign \new_[63245]_  = ~A299 & A298;
  assign \new_[63249]_  = A302 & ~A301;
  assign \new_[63250]_  = ~A300 & \new_[63249]_ ;
  assign \new_[63251]_  = \new_[63250]_  & \new_[63245]_ ;
  assign \new_[63252]_  = \new_[63251]_  & \new_[63242]_ ;
  assign \new_[63255]_  = A200 & ~A199;
  assign \new_[63258]_  = ~A202 & ~A201;
  assign \new_[63259]_  = \new_[63258]_  & \new_[63255]_ ;
  assign \new_[63262]_  = ~A232 & A203;
  assign \new_[63265]_  = ~A234 & A233;
  assign \new_[63266]_  = \new_[63265]_  & \new_[63262]_ ;
  assign \new_[63267]_  = \new_[63266]_  & \new_[63259]_ ;
  assign \new_[63270]_  = A236 & ~A235;
  assign \new_[63273]_  = A266 & A265;
  assign \new_[63274]_  = \new_[63273]_  & \new_[63270]_ ;
  assign \new_[63277]_  = A299 & ~A298;
  assign \new_[63281]_  = A302 & ~A301;
  assign \new_[63282]_  = ~A300 & \new_[63281]_ ;
  assign \new_[63283]_  = \new_[63282]_  & \new_[63277]_ ;
  assign \new_[63284]_  = \new_[63283]_  & \new_[63274]_ ;
  assign \new_[63287]_  = A200 & ~A199;
  assign \new_[63290]_  = ~A202 & ~A201;
  assign \new_[63291]_  = \new_[63290]_  & \new_[63287]_ ;
  assign \new_[63294]_  = ~A232 & A203;
  assign \new_[63297]_  = ~A234 & A233;
  assign \new_[63298]_  = \new_[63297]_  & \new_[63294]_ ;
  assign \new_[63299]_  = \new_[63298]_  & \new_[63291]_ ;
  assign \new_[63302]_  = A236 & ~A235;
  assign \new_[63305]_  = ~A266 & ~A265;
  assign \new_[63306]_  = \new_[63305]_  & \new_[63302]_ ;
  assign \new_[63309]_  = ~A299 & A298;
  assign \new_[63313]_  = A302 & ~A301;
  assign \new_[63314]_  = ~A300 & \new_[63313]_ ;
  assign \new_[63315]_  = \new_[63314]_  & \new_[63309]_ ;
  assign \new_[63316]_  = \new_[63315]_  & \new_[63306]_ ;
  assign \new_[63319]_  = A200 & ~A199;
  assign \new_[63322]_  = ~A202 & ~A201;
  assign \new_[63323]_  = \new_[63322]_  & \new_[63319]_ ;
  assign \new_[63326]_  = ~A232 & A203;
  assign \new_[63329]_  = ~A234 & A233;
  assign \new_[63330]_  = \new_[63329]_  & \new_[63326]_ ;
  assign \new_[63331]_  = \new_[63330]_  & \new_[63323]_ ;
  assign \new_[63334]_  = A236 & ~A235;
  assign \new_[63337]_  = ~A266 & ~A265;
  assign \new_[63338]_  = \new_[63337]_  & \new_[63334]_ ;
  assign \new_[63341]_  = A299 & ~A298;
  assign \new_[63345]_  = A302 & ~A301;
  assign \new_[63346]_  = ~A300 & \new_[63345]_ ;
  assign \new_[63347]_  = \new_[63346]_  & \new_[63341]_ ;
  assign \new_[63348]_  = \new_[63347]_  & \new_[63338]_ ;
  assign \new_[63351]_  = A200 & ~A199;
  assign \new_[63354]_  = ~A202 & ~A201;
  assign \new_[63355]_  = \new_[63354]_  & \new_[63351]_ ;
  assign \new_[63358]_  = A232 & A203;
  assign \new_[63361]_  = A234 & ~A233;
  assign \new_[63362]_  = \new_[63361]_  & \new_[63358]_ ;
  assign \new_[63363]_  = \new_[63362]_  & \new_[63355]_ ;
  assign \new_[63366]_  = A267 & A235;
  assign \new_[63369]_  = A269 & ~A268;
  assign \new_[63370]_  = \new_[63369]_  & \new_[63366]_ ;
  assign \new_[63373]_  = ~A299 & A298;
  assign \new_[63377]_  = A302 & ~A301;
  assign \new_[63378]_  = ~A300 & \new_[63377]_ ;
  assign \new_[63379]_  = \new_[63378]_  & \new_[63373]_ ;
  assign \new_[63380]_  = \new_[63379]_  & \new_[63370]_ ;
  assign \new_[63383]_  = A200 & ~A199;
  assign \new_[63386]_  = ~A202 & ~A201;
  assign \new_[63387]_  = \new_[63386]_  & \new_[63383]_ ;
  assign \new_[63390]_  = A232 & A203;
  assign \new_[63393]_  = A234 & ~A233;
  assign \new_[63394]_  = \new_[63393]_  & \new_[63390]_ ;
  assign \new_[63395]_  = \new_[63394]_  & \new_[63387]_ ;
  assign \new_[63398]_  = A267 & A235;
  assign \new_[63401]_  = A269 & ~A268;
  assign \new_[63402]_  = \new_[63401]_  & \new_[63398]_ ;
  assign \new_[63405]_  = A299 & ~A298;
  assign \new_[63409]_  = A302 & ~A301;
  assign \new_[63410]_  = ~A300 & \new_[63409]_ ;
  assign \new_[63411]_  = \new_[63410]_  & \new_[63405]_ ;
  assign \new_[63412]_  = \new_[63411]_  & \new_[63402]_ ;
  assign \new_[63415]_  = A200 & ~A199;
  assign \new_[63418]_  = ~A202 & ~A201;
  assign \new_[63419]_  = \new_[63418]_  & \new_[63415]_ ;
  assign \new_[63422]_  = A232 & A203;
  assign \new_[63425]_  = A234 & ~A233;
  assign \new_[63426]_  = \new_[63425]_  & \new_[63422]_ ;
  assign \new_[63427]_  = \new_[63426]_  & \new_[63419]_ ;
  assign \new_[63430]_  = A267 & ~A236;
  assign \new_[63433]_  = A269 & ~A268;
  assign \new_[63434]_  = \new_[63433]_  & \new_[63430]_ ;
  assign \new_[63437]_  = ~A299 & A298;
  assign \new_[63441]_  = A302 & ~A301;
  assign \new_[63442]_  = ~A300 & \new_[63441]_ ;
  assign \new_[63443]_  = \new_[63442]_  & \new_[63437]_ ;
  assign \new_[63444]_  = \new_[63443]_  & \new_[63434]_ ;
  assign \new_[63447]_  = A200 & ~A199;
  assign \new_[63450]_  = ~A202 & ~A201;
  assign \new_[63451]_  = \new_[63450]_  & \new_[63447]_ ;
  assign \new_[63454]_  = A232 & A203;
  assign \new_[63457]_  = A234 & ~A233;
  assign \new_[63458]_  = \new_[63457]_  & \new_[63454]_ ;
  assign \new_[63459]_  = \new_[63458]_  & \new_[63451]_ ;
  assign \new_[63462]_  = A267 & ~A236;
  assign \new_[63465]_  = A269 & ~A268;
  assign \new_[63466]_  = \new_[63465]_  & \new_[63462]_ ;
  assign \new_[63469]_  = A299 & ~A298;
  assign \new_[63473]_  = A302 & ~A301;
  assign \new_[63474]_  = ~A300 & \new_[63473]_ ;
  assign \new_[63475]_  = \new_[63474]_  & \new_[63469]_ ;
  assign \new_[63476]_  = \new_[63475]_  & \new_[63466]_ ;
  assign \new_[63479]_  = A200 & ~A199;
  assign \new_[63482]_  = ~A202 & ~A201;
  assign \new_[63483]_  = \new_[63482]_  & \new_[63479]_ ;
  assign \new_[63486]_  = A232 & A203;
  assign \new_[63489]_  = ~A234 & ~A233;
  assign \new_[63490]_  = \new_[63489]_  & \new_[63486]_ ;
  assign \new_[63491]_  = \new_[63490]_  & \new_[63483]_ ;
  assign \new_[63494]_  = A236 & ~A235;
  assign \new_[63497]_  = ~A268 & A267;
  assign \new_[63498]_  = \new_[63497]_  & \new_[63494]_ ;
  assign \new_[63501]_  = A298 & A269;
  assign \new_[63505]_  = A301 & A300;
  assign \new_[63506]_  = ~A299 & \new_[63505]_ ;
  assign \new_[63507]_  = \new_[63506]_  & \new_[63501]_ ;
  assign \new_[63508]_  = \new_[63507]_  & \new_[63498]_ ;
  assign \new_[63511]_  = A200 & ~A199;
  assign \new_[63514]_  = ~A202 & ~A201;
  assign \new_[63515]_  = \new_[63514]_  & \new_[63511]_ ;
  assign \new_[63518]_  = A232 & A203;
  assign \new_[63521]_  = ~A234 & ~A233;
  assign \new_[63522]_  = \new_[63521]_  & \new_[63518]_ ;
  assign \new_[63523]_  = \new_[63522]_  & \new_[63515]_ ;
  assign \new_[63526]_  = A236 & ~A235;
  assign \new_[63529]_  = ~A268 & A267;
  assign \new_[63530]_  = \new_[63529]_  & \new_[63526]_ ;
  assign \new_[63533]_  = A298 & A269;
  assign \new_[63537]_  = ~A302 & A300;
  assign \new_[63538]_  = ~A299 & \new_[63537]_ ;
  assign \new_[63539]_  = \new_[63538]_  & \new_[63533]_ ;
  assign \new_[63540]_  = \new_[63539]_  & \new_[63530]_ ;
  assign \new_[63543]_  = A200 & ~A199;
  assign \new_[63546]_  = ~A202 & ~A201;
  assign \new_[63547]_  = \new_[63546]_  & \new_[63543]_ ;
  assign \new_[63550]_  = A232 & A203;
  assign \new_[63553]_  = ~A234 & ~A233;
  assign \new_[63554]_  = \new_[63553]_  & \new_[63550]_ ;
  assign \new_[63555]_  = \new_[63554]_  & \new_[63547]_ ;
  assign \new_[63558]_  = A236 & ~A235;
  assign \new_[63561]_  = ~A268 & A267;
  assign \new_[63562]_  = \new_[63561]_  & \new_[63558]_ ;
  assign \new_[63565]_  = ~A298 & A269;
  assign \new_[63569]_  = A301 & A300;
  assign \new_[63570]_  = A299 & \new_[63569]_ ;
  assign \new_[63571]_  = \new_[63570]_  & \new_[63565]_ ;
  assign \new_[63572]_  = \new_[63571]_  & \new_[63562]_ ;
  assign \new_[63575]_  = A200 & ~A199;
  assign \new_[63578]_  = ~A202 & ~A201;
  assign \new_[63579]_  = \new_[63578]_  & \new_[63575]_ ;
  assign \new_[63582]_  = A232 & A203;
  assign \new_[63585]_  = ~A234 & ~A233;
  assign \new_[63586]_  = \new_[63585]_  & \new_[63582]_ ;
  assign \new_[63587]_  = \new_[63586]_  & \new_[63579]_ ;
  assign \new_[63590]_  = A236 & ~A235;
  assign \new_[63593]_  = ~A268 & A267;
  assign \new_[63594]_  = \new_[63593]_  & \new_[63590]_ ;
  assign \new_[63597]_  = ~A298 & A269;
  assign \new_[63601]_  = ~A302 & A300;
  assign \new_[63602]_  = A299 & \new_[63601]_ ;
  assign \new_[63603]_  = \new_[63602]_  & \new_[63597]_ ;
  assign \new_[63604]_  = \new_[63603]_  & \new_[63594]_ ;
  assign \new_[63607]_  = A200 & ~A199;
  assign \new_[63610]_  = ~A202 & ~A201;
  assign \new_[63611]_  = \new_[63610]_  & \new_[63607]_ ;
  assign \new_[63614]_  = A232 & A203;
  assign \new_[63617]_  = ~A234 & ~A233;
  assign \new_[63618]_  = \new_[63617]_  & \new_[63614]_ ;
  assign \new_[63619]_  = \new_[63618]_  & \new_[63611]_ ;
  assign \new_[63622]_  = A236 & ~A235;
  assign \new_[63625]_  = A268 & ~A267;
  assign \new_[63626]_  = \new_[63625]_  & \new_[63622]_ ;
  assign \new_[63629]_  = ~A299 & A298;
  assign \new_[63633]_  = A302 & ~A301;
  assign \new_[63634]_  = ~A300 & \new_[63633]_ ;
  assign \new_[63635]_  = \new_[63634]_  & \new_[63629]_ ;
  assign \new_[63636]_  = \new_[63635]_  & \new_[63626]_ ;
  assign \new_[63639]_  = A200 & ~A199;
  assign \new_[63642]_  = ~A202 & ~A201;
  assign \new_[63643]_  = \new_[63642]_  & \new_[63639]_ ;
  assign \new_[63646]_  = A232 & A203;
  assign \new_[63649]_  = ~A234 & ~A233;
  assign \new_[63650]_  = \new_[63649]_  & \new_[63646]_ ;
  assign \new_[63651]_  = \new_[63650]_  & \new_[63643]_ ;
  assign \new_[63654]_  = A236 & ~A235;
  assign \new_[63657]_  = A268 & ~A267;
  assign \new_[63658]_  = \new_[63657]_  & \new_[63654]_ ;
  assign \new_[63661]_  = A299 & ~A298;
  assign \new_[63665]_  = A302 & ~A301;
  assign \new_[63666]_  = ~A300 & \new_[63665]_ ;
  assign \new_[63667]_  = \new_[63666]_  & \new_[63661]_ ;
  assign \new_[63668]_  = \new_[63667]_  & \new_[63658]_ ;
  assign \new_[63671]_  = A200 & ~A199;
  assign \new_[63674]_  = ~A202 & ~A201;
  assign \new_[63675]_  = \new_[63674]_  & \new_[63671]_ ;
  assign \new_[63678]_  = A232 & A203;
  assign \new_[63681]_  = ~A234 & ~A233;
  assign \new_[63682]_  = \new_[63681]_  & \new_[63678]_ ;
  assign \new_[63683]_  = \new_[63682]_  & \new_[63675]_ ;
  assign \new_[63686]_  = A236 & ~A235;
  assign \new_[63689]_  = ~A269 & ~A267;
  assign \new_[63690]_  = \new_[63689]_  & \new_[63686]_ ;
  assign \new_[63693]_  = ~A299 & A298;
  assign \new_[63697]_  = A302 & ~A301;
  assign \new_[63698]_  = ~A300 & \new_[63697]_ ;
  assign \new_[63699]_  = \new_[63698]_  & \new_[63693]_ ;
  assign \new_[63700]_  = \new_[63699]_  & \new_[63690]_ ;
  assign \new_[63703]_  = A200 & ~A199;
  assign \new_[63706]_  = ~A202 & ~A201;
  assign \new_[63707]_  = \new_[63706]_  & \new_[63703]_ ;
  assign \new_[63710]_  = A232 & A203;
  assign \new_[63713]_  = ~A234 & ~A233;
  assign \new_[63714]_  = \new_[63713]_  & \new_[63710]_ ;
  assign \new_[63715]_  = \new_[63714]_  & \new_[63707]_ ;
  assign \new_[63718]_  = A236 & ~A235;
  assign \new_[63721]_  = ~A269 & ~A267;
  assign \new_[63722]_  = \new_[63721]_  & \new_[63718]_ ;
  assign \new_[63725]_  = A299 & ~A298;
  assign \new_[63729]_  = A302 & ~A301;
  assign \new_[63730]_  = ~A300 & \new_[63729]_ ;
  assign \new_[63731]_  = \new_[63730]_  & \new_[63725]_ ;
  assign \new_[63732]_  = \new_[63731]_  & \new_[63722]_ ;
  assign \new_[63735]_  = A200 & ~A199;
  assign \new_[63738]_  = ~A202 & ~A201;
  assign \new_[63739]_  = \new_[63738]_  & \new_[63735]_ ;
  assign \new_[63742]_  = A232 & A203;
  assign \new_[63745]_  = ~A234 & ~A233;
  assign \new_[63746]_  = \new_[63745]_  & \new_[63742]_ ;
  assign \new_[63747]_  = \new_[63746]_  & \new_[63739]_ ;
  assign \new_[63750]_  = A236 & ~A235;
  assign \new_[63753]_  = A266 & A265;
  assign \new_[63754]_  = \new_[63753]_  & \new_[63750]_ ;
  assign \new_[63757]_  = ~A299 & A298;
  assign \new_[63761]_  = A302 & ~A301;
  assign \new_[63762]_  = ~A300 & \new_[63761]_ ;
  assign \new_[63763]_  = \new_[63762]_  & \new_[63757]_ ;
  assign \new_[63764]_  = \new_[63763]_  & \new_[63754]_ ;
  assign \new_[63767]_  = A200 & ~A199;
  assign \new_[63770]_  = ~A202 & ~A201;
  assign \new_[63771]_  = \new_[63770]_  & \new_[63767]_ ;
  assign \new_[63774]_  = A232 & A203;
  assign \new_[63777]_  = ~A234 & ~A233;
  assign \new_[63778]_  = \new_[63777]_  & \new_[63774]_ ;
  assign \new_[63779]_  = \new_[63778]_  & \new_[63771]_ ;
  assign \new_[63782]_  = A236 & ~A235;
  assign \new_[63785]_  = A266 & A265;
  assign \new_[63786]_  = \new_[63785]_  & \new_[63782]_ ;
  assign \new_[63789]_  = A299 & ~A298;
  assign \new_[63793]_  = A302 & ~A301;
  assign \new_[63794]_  = ~A300 & \new_[63793]_ ;
  assign \new_[63795]_  = \new_[63794]_  & \new_[63789]_ ;
  assign \new_[63796]_  = \new_[63795]_  & \new_[63786]_ ;
  assign \new_[63799]_  = A200 & ~A199;
  assign \new_[63802]_  = ~A202 & ~A201;
  assign \new_[63803]_  = \new_[63802]_  & \new_[63799]_ ;
  assign \new_[63806]_  = A232 & A203;
  assign \new_[63809]_  = ~A234 & ~A233;
  assign \new_[63810]_  = \new_[63809]_  & \new_[63806]_ ;
  assign \new_[63811]_  = \new_[63810]_  & \new_[63803]_ ;
  assign \new_[63814]_  = A236 & ~A235;
  assign \new_[63817]_  = ~A266 & ~A265;
  assign \new_[63818]_  = \new_[63817]_  & \new_[63814]_ ;
  assign \new_[63821]_  = ~A299 & A298;
  assign \new_[63825]_  = A302 & ~A301;
  assign \new_[63826]_  = ~A300 & \new_[63825]_ ;
  assign \new_[63827]_  = \new_[63826]_  & \new_[63821]_ ;
  assign \new_[63828]_  = \new_[63827]_  & \new_[63818]_ ;
  assign \new_[63831]_  = A200 & ~A199;
  assign \new_[63834]_  = ~A202 & ~A201;
  assign \new_[63835]_  = \new_[63834]_  & \new_[63831]_ ;
  assign \new_[63838]_  = A232 & A203;
  assign \new_[63841]_  = ~A234 & ~A233;
  assign \new_[63842]_  = \new_[63841]_  & \new_[63838]_ ;
  assign \new_[63843]_  = \new_[63842]_  & \new_[63835]_ ;
  assign \new_[63846]_  = A236 & ~A235;
  assign \new_[63849]_  = ~A266 & ~A265;
  assign \new_[63850]_  = \new_[63849]_  & \new_[63846]_ ;
  assign \new_[63853]_  = A299 & ~A298;
  assign \new_[63857]_  = A302 & ~A301;
  assign \new_[63858]_  = ~A300 & \new_[63857]_ ;
  assign \new_[63859]_  = \new_[63858]_  & \new_[63853]_ ;
  assign \new_[63860]_  = \new_[63859]_  & \new_[63850]_ ;
  assign \new_[63863]_  = ~A200 & A199;
  assign \new_[63866]_  = A202 & A201;
  assign \new_[63867]_  = \new_[63866]_  & \new_[63863]_ ;
  assign \new_[63870]_  = A233 & ~A232;
  assign \new_[63873]_  = ~A235 & ~A234;
  assign \new_[63874]_  = \new_[63873]_  & \new_[63870]_ ;
  assign \new_[63875]_  = \new_[63874]_  & \new_[63867]_ ;
  assign \new_[63878]_  = A267 & A236;
  assign \new_[63881]_  = A269 & ~A268;
  assign \new_[63882]_  = \new_[63881]_  & \new_[63878]_ ;
  assign \new_[63885]_  = ~A299 & A298;
  assign \new_[63889]_  = A302 & ~A301;
  assign \new_[63890]_  = ~A300 & \new_[63889]_ ;
  assign \new_[63891]_  = \new_[63890]_  & \new_[63885]_ ;
  assign \new_[63892]_  = \new_[63891]_  & \new_[63882]_ ;
  assign \new_[63895]_  = ~A200 & A199;
  assign \new_[63898]_  = A202 & A201;
  assign \new_[63899]_  = \new_[63898]_  & \new_[63895]_ ;
  assign \new_[63902]_  = A233 & ~A232;
  assign \new_[63905]_  = ~A235 & ~A234;
  assign \new_[63906]_  = \new_[63905]_  & \new_[63902]_ ;
  assign \new_[63907]_  = \new_[63906]_  & \new_[63899]_ ;
  assign \new_[63910]_  = A267 & A236;
  assign \new_[63913]_  = A269 & ~A268;
  assign \new_[63914]_  = \new_[63913]_  & \new_[63910]_ ;
  assign \new_[63917]_  = A299 & ~A298;
  assign \new_[63921]_  = A302 & ~A301;
  assign \new_[63922]_  = ~A300 & \new_[63921]_ ;
  assign \new_[63923]_  = \new_[63922]_  & \new_[63917]_ ;
  assign \new_[63924]_  = \new_[63923]_  & \new_[63914]_ ;
  assign \new_[63927]_  = ~A200 & A199;
  assign \new_[63930]_  = A202 & A201;
  assign \new_[63931]_  = \new_[63930]_  & \new_[63927]_ ;
  assign \new_[63934]_  = ~A233 & A232;
  assign \new_[63937]_  = ~A235 & ~A234;
  assign \new_[63938]_  = \new_[63937]_  & \new_[63934]_ ;
  assign \new_[63939]_  = \new_[63938]_  & \new_[63931]_ ;
  assign \new_[63942]_  = A267 & A236;
  assign \new_[63945]_  = A269 & ~A268;
  assign \new_[63946]_  = \new_[63945]_  & \new_[63942]_ ;
  assign \new_[63949]_  = ~A299 & A298;
  assign \new_[63953]_  = A302 & ~A301;
  assign \new_[63954]_  = ~A300 & \new_[63953]_ ;
  assign \new_[63955]_  = \new_[63954]_  & \new_[63949]_ ;
  assign \new_[63956]_  = \new_[63955]_  & \new_[63946]_ ;
  assign \new_[63959]_  = ~A200 & A199;
  assign \new_[63962]_  = A202 & A201;
  assign \new_[63963]_  = \new_[63962]_  & \new_[63959]_ ;
  assign \new_[63966]_  = ~A233 & A232;
  assign \new_[63969]_  = ~A235 & ~A234;
  assign \new_[63970]_  = \new_[63969]_  & \new_[63966]_ ;
  assign \new_[63971]_  = \new_[63970]_  & \new_[63963]_ ;
  assign \new_[63974]_  = A267 & A236;
  assign \new_[63977]_  = A269 & ~A268;
  assign \new_[63978]_  = \new_[63977]_  & \new_[63974]_ ;
  assign \new_[63981]_  = A299 & ~A298;
  assign \new_[63985]_  = A302 & ~A301;
  assign \new_[63986]_  = ~A300 & \new_[63985]_ ;
  assign \new_[63987]_  = \new_[63986]_  & \new_[63981]_ ;
  assign \new_[63988]_  = \new_[63987]_  & \new_[63978]_ ;
  assign \new_[63991]_  = ~A200 & A199;
  assign \new_[63994]_  = ~A203 & A201;
  assign \new_[63995]_  = \new_[63994]_  & \new_[63991]_ ;
  assign \new_[63998]_  = A233 & ~A232;
  assign \new_[64001]_  = ~A235 & ~A234;
  assign \new_[64002]_  = \new_[64001]_  & \new_[63998]_ ;
  assign \new_[64003]_  = \new_[64002]_  & \new_[63995]_ ;
  assign \new_[64006]_  = A267 & A236;
  assign \new_[64009]_  = A269 & ~A268;
  assign \new_[64010]_  = \new_[64009]_  & \new_[64006]_ ;
  assign \new_[64013]_  = ~A299 & A298;
  assign \new_[64017]_  = A302 & ~A301;
  assign \new_[64018]_  = ~A300 & \new_[64017]_ ;
  assign \new_[64019]_  = \new_[64018]_  & \new_[64013]_ ;
  assign \new_[64020]_  = \new_[64019]_  & \new_[64010]_ ;
  assign \new_[64023]_  = ~A200 & A199;
  assign \new_[64026]_  = ~A203 & A201;
  assign \new_[64027]_  = \new_[64026]_  & \new_[64023]_ ;
  assign \new_[64030]_  = A233 & ~A232;
  assign \new_[64033]_  = ~A235 & ~A234;
  assign \new_[64034]_  = \new_[64033]_  & \new_[64030]_ ;
  assign \new_[64035]_  = \new_[64034]_  & \new_[64027]_ ;
  assign \new_[64038]_  = A267 & A236;
  assign \new_[64041]_  = A269 & ~A268;
  assign \new_[64042]_  = \new_[64041]_  & \new_[64038]_ ;
  assign \new_[64045]_  = A299 & ~A298;
  assign \new_[64049]_  = A302 & ~A301;
  assign \new_[64050]_  = ~A300 & \new_[64049]_ ;
  assign \new_[64051]_  = \new_[64050]_  & \new_[64045]_ ;
  assign \new_[64052]_  = \new_[64051]_  & \new_[64042]_ ;
  assign \new_[64055]_  = ~A200 & A199;
  assign \new_[64058]_  = ~A203 & A201;
  assign \new_[64059]_  = \new_[64058]_  & \new_[64055]_ ;
  assign \new_[64062]_  = ~A233 & A232;
  assign \new_[64065]_  = ~A235 & ~A234;
  assign \new_[64066]_  = \new_[64065]_  & \new_[64062]_ ;
  assign \new_[64067]_  = \new_[64066]_  & \new_[64059]_ ;
  assign \new_[64070]_  = A267 & A236;
  assign \new_[64073]_  = A269 & ~A268;
  assign \new_[64074]_  = \new_[64073]_  & \new_[64070]_ ;
  assign \new_[64077]_  = ~A299 & A298;
  assign \new_[64081]_  = A302 & ~A301;
  assign \new_[64082]_  = ~A300 & \new_[64081]_ ;
  assign \new_[64083]_  = \new_[64082]_  & \new_[64077]_ ;
  assign \new_[64084]_  = \new_[64083]_  & \new_[64074]_ ;
  assign \new_[64087]_  = ~A200 & A199;
  assign \new_[64090]_  = ~A203 & A201;
  assign \new_[64091]_  = \new_[64090]_  & \new_[64087]_ ;
  assign \new_[64094]_  = ~A233 & A232;
  assign \new_[64097]_  = ~A235 & ~A234;
  assign \new_[64098]_  = \new_[64097]_  & \new_[64094]_ ;
  assign \new_[64099]_  = \new_[64098]_  & \new_[64091]_ ;
  assign \new_[64102]_  = A267 & A236;
  assign \new_[64105]_  = A269 & ~A268;
  assign \new_[64106]_  = \new_[64105]_  & \new_[64102]_ ;
  assign \new_[64109]_  = A299 & ~A298;
  assign \new_[64113]_  = A302 & ~A301;
  assign \new_[64114]_  = ~A300 & \new_[64113]_ ;
  assign \new_[64115]_  = \new_[64114]_  & \new_[64109]_ ;
  assign \new_[64116]_  = \new_[64115]_  & \new_[64106]_ ;
  assign \new_[64119]_  = ~A200 & A199;
  assign \new_[64122]_  = ~A202 & ~A201;
  assign \new_[64123]_  = \new_[64122]_  & \new_[64119]_ ;
  assign \new_[64126]_  = ~A232 & A203;
  assign \new_[64129]_  = A234 & A233;
  assign \new_[64130]_  = \new_[64129]_  & \new_[64126]_ ;
  assign \new_[64131]_  = \new_[64130]_  & \new_[64123]_ ;
  assign \new_[64134]_  = A267 & A235;
  assign \new_[64137]_  = A269 & ~A268;
  assign \new_[64138]_  = \new_[64137]_  & \new_[64134]_ ;
  assign \new_[64141]_  = ~A299 & A298;
  assign \new_[64145]_  = A302 & ~A301;
  assign \new_[64146]_  = ~A300 & \new_[64145]_ ;
  assign \new_[64147]_  = \new_[64146]_  & \new_[64141]_ ;
  assign \new_[64148]_  = \new_[64147]_  & \new_[64138]_ ;
  assign \new_[64151]_  = ~A200 & A199;
  assign \new_[64154]_  = ~A202 & ~A201;
  assign \new_[64155]_  = \new_[64154]_  & \new_[64151]_ ;
  assign \new_[64158]_  = ~A232 & A203;
  assign \new_[64161]_  = A234 & A233;
  assign \new_[64162]_  = \new_[64161]_  & \new_[64158]_ ;
  assign \new_[64163]_  = \new_[64162]_  & \new_[64155]_ ;
  assign \new_[64166]_  = A267 & A235;
  assign \new_[64169]_  = A269 & ~A268;
  assign \new_[64170]_  = \new_[64169]_  & \new_[64166]_ ;
  assign \new_[64173]_  = A299 & ~A298;
  assign \new_[64177]_  = A302 & ~A301;
  assign \new_[64178]_  = ~A300 & \new_[64177]_ ;
  assign \new_[64179]_  = \new_[64178]_  & \new_[64173]_ ;
  assign \new_[64180]_  = \new_[64179]_  & \new_[64170]_ ;
  assign \new_[64183]_  = ~A200 & A199;
  assign \new_[64186]_  = ~A202 & ~A201;
  assign \new_[64187]_  = \new_[64186]_  & \new_[64183]_ ;
  assign \new_[64190]_  = ~A232 & A203;
  assign \new_[64193]_  = A234 & A233;
  assign \new_[64194]_  = \new_[64193]_  & \new_[64190]_ ;
  assign \new_[64195]_  = \new_[64194]_  & \new_[64187]_ ;
  assign \new_[64198]_  = A267 & ~A236;
  assign \new_[64201]_  = A269 & ~A268;
  assign \new_[64202]_  = \new_[64201]_  & \new_[64198]_ ;
  assign \new_[64205]_  = ~A299 & A298;
  assign \new_[64209]_  = A302 & ~A301;
  assign \new_[64210]_  = ~A300 & \new_[64209]_ ;
  assign \new_[64211]_  = \new_[64210]_  & \new_[64205]_ ;
  assign \new_[64212]_  = \new_[64211]_  & \new_[64202]_ ;
  assign \new_[64215]_  = ~A200 & A199;
  assign \new_[64218]_  = ~A202 & ~A201;
  assign \new_[64219]_  = \new_[64218]_  & \new_[64215]_ ;
  assign \new_[64222]_  = ~A232 & A203;
  assign \new_[64225]_  = A234 & A233;
  assign \new_[64226]_  = \new_[64225]_  & \new_[64222]_ ;
  assign \new_[64227]_  = \new_[64226]_  & \new_[64219]_ ;
  assign \new_[64230]_  = A267 & ~A236;
  assign \new_[64233]_  = A269 & ~A268;
  assign \new_[64234]_  = \new_[64233]_  & \new_[64230]_ ;
  assign \new_[64237]_  = A299 & ~A298;
  assign \new_[64241]_  = A302 & ~A301;
  assign \new_[64242]_  = ~A300 & \new_[64241]_ ;
  assign \new_[64243]_  = \new_[64242]_  & \new_[64237]_ ;
  assign \new_[64244]_  = \new_[64243]_  & \new_[64234]_ ;
  assign \new_[64247]_  = ~A200 & A199;
  assign \new_[64250]_  = ~A202 & ~A201;
  assign \new_[64251]_  = \new_[64250]_  & \new_[64247]_ ;
  assign \new_[64254]_  = ~A232 & A203;
  assign \new_[64257]_  = ~A234 & A233;
  assign \new_[64258]_  = \new_[64257]_  & \new_[64254]_ ;
  assign \new_[64259]_  = \new_[64258]_  & \new_[64251]_ ;
  assign \new_[64262]_  = A236 & ~A235;
  assign \new_[64265]_  = ~A268 & A267;
  assign \new_[64266]_  = \new_[64265]_  & \new_[64262]_ ;
  assign \new_[64269]_  = A298 & A269;
  assign \new_[64273]_  = A301 & A300;
  assign \new_[64274]_  = ~A299 & \new_[64273]_ ;
  assign \new_[64275]_  = \new_[64274]_  & \new_[64269]_ ;
  assign \new_[64276]_  = \new_[64275]_  & \new_[64266]_ ;
  assign \new_[64279]_  = ~A200 & A199;
  assign \new_[64282]_  = ~A202 & ~A201;
  assign \new_[64283]_  = \new_[64282]_  & \new_[64279]_ ;
  assign \new_[64286]_  = ~A232 & A203;
  assign \new_[64289]_  = ~A234 & A233;
  assign \new_[64290]_  = \new_[64289]_  & \new_[64286]_ ;
  assign \new_[64291]_  = \new_[64290]_  & \new_[64283]_ ;
  assign \new_[64294]_  = A236 & ~A235;
  assign \new_[64297]_  = ~A268 & A267;
  assign \new_[64298]_  = \new_[64297]_  & \new_[64294]_ ;
  assign \new_[64301]_  = A298 & A269;
  assign \new_[64305]_  = ~A302 & A300;
  assign \new_[64306]_  = ~A299 & \new_[64305]_ ;
  assign \new_[64307]_  = \new_[64306]_  & \new_[64301]_ ;
  assign \new_[64308]_  = \new_[64307]_  & \new_[64298]_ ;
  assign \new_[64311]_  = ~A200 & A199;
  assign \new_[64314]_  = ~A202 & ~A201;
  assign \new_[64315]_  = \new_[64314]_  & \new_[64311]_ ;
  assign \new_[64318]_  = ~A232 & A203;
  assign \new_[64321]_  = ~A234 & A233;
  assign \new_[64322]_  = \new_[64321]_  & \new_[64318]_ ;
  assign \new_[64323]_  = \new_[64322]_  & \new_[64315]_ ;
  assign \new_[64326]_  = A236 & ~A235;
  assign \new_[64329]_  = ~A268 & A267;
  assign \new_[64330]_  = \new_[64329]_  & \new_[64326]_ ;
  assign \new_[64333]_  = ~A298 & A269;
  assign \new_[64337]_  = A301 & A300;
  assign \new_[64338]_  = A299 & \new_[64337]_ ;
  assign \new_[64339]_  = \new_[64338]_  & \new_[64333]_ ;
  assign \new_[64340]_  = \new_[64339]_  & \new_[64330]_ ;
  assign \new_[64343]_  = ~A200 & A199;
  assign \new_[64346]_  = ~A202 & ~A201;
  assign \new_[64347]_  = \new_[64346]_  & \new_[64343]_ ;
  assign \new_[64350]_  = ~A232 & A203;
  assign \new_[64353]_  = ~A234 & A233;
  assign \new_[64354]_  = \new_[64353]_  & \new_[64350]_ ;
  assign \new_[64355]_  = \new_[64354]_  & \new_[64347]_ ;
  assign \new_[64358]_  = A236 & ~A235;
  assign \new_[64361]_  = ~A268 & A267;
  assign \new_[64362]_  = \new_[64361]_  & \new_[64358]_ ;
  assign \new_[64365]_  = ~A298 & A269;
  assign \new_[64369]_  = ~A302 & A300;
  assign \new_[64370]_  = A299 & \new_[64369]_ ;
  assign \new_[64371]_  = \new_[64370]_  & \new_[64365]_ ;
  assign \new_[64372]_  = \new_[64371]_  & \new_[64362]_ ;
  assign \new_[64375]_  = ~A200 & A199;
  assign \new_[64378]_  = ~A202 & ~A201;
  assign \new_[64379]_  = \new_[64378]_  & \new_[64375]_ ;
  assign \new_[64382]_  = ~A232 & A203;
  assign \new_[64385]_  = ~A234 & A233;
  assign \new_[64386]_  = \new_[64385]_  & \new_[64382]_ ;
  assign \new_[64387]_  = \new_[64386]_  & \new_[64379]_ ;
  assign \new_[64390]_  = A236 & ~A235;
  assign \new_[64393]_  = A268 & ~A267;
  assign \new_[64394]_  = \new_[64393]_  & \new_[64390]_ ;
  assign \new_[64397]_  = ~A299 & A298;
  assign \new_[64401]_  = A302 & ~A301;
  assign \new_[64402]_  = ~A300 & \new_[64401]_ ;
  assign \new_[64403]_  = \new_[64402]_  & \new_[64397]_ ;
  assign \new_[64404]_  = \new_[64403]_  & \new_[64394]_ ;
  assign \new_[64407]_  = ~A200 & A199;
  assign \new_[64410]_  = ~A202 & ~A201;
  assign \new_[64411]_  = \new_[64410]_  & \new_[64407]_ ;
  assign \new_[64414]_  = ~A232 & A203;
  assign \new_[64417]_  = ~A234 & A233;
  assign \new_[64418]_  = \new_[64417]_  & \new_[64414]_ ;
  assign \new_[64419]_  = \new_[64418]_  & \new_[64411]_ ;
  assign \new_[64422]_  = A236 & ~A235;
  assign \new_[64425]_  = A268 & ~A267;
  assign \new_[64426]_  = \new_[64425]_  & \new_[64422]_ ;
  assign \new_[64429]_  = A299 & ~A298;
  assign \new_[64433]_  = A302 & ~A301;
  assign \new_[64434]_  = ~A300 & \new_[64433]_ ;
  assign \new_[64435]_  = \new_[64434]_  & \new_[64429]_ ;
  assign \new_[64436]_  = \new_[64435]_  & \new_[64426]_ ;
  assign \new_[64439]_  = ~A200 & A199;
  assign \new_[64442]_  = ~A202 & ~A201;
  assign \new_[64443]_  = \new_[64442]_  & \new_[64439]_ ;
  assign \new_[64446]_  = ~A232 & A203;
  assign \new_[64449]_  = ~A234 & A233;
  assign \new_[64450]_  = \new_[64449]_  & \new_[64446]_ ;
  assign \new_[64451]_  = \new_[64450]_  & \new_[64443]_ ;
  assign \new_[64454]_  = A236 & ~A235;
  assign \new_[64457]_  = ~A269 & ~A267;
  assign \new_[64458]_  = \new_[64457]_  & \new_[64454]_ ;
  assign \new_[64461]_  = ~A299 & A298;
  assign \new_[64465]_  = A302 & ~A301;
  assign \new_[64466]_  = ~A300 & \new_[64465]_ ;
  assign \new_[64467]_  = \new_[64466]_  & \new_[64461]_ ;
  assign \new_[64468]_  = \new_[64467]_  & \new_[64458]_ ;
  assign \new_[64471]_  = ~A200 & A199;
  assign \new_[64474]_  = ~A202 & ~A201;
  assign \new_[64475]_  = \new_[64474]_  & \new_[64471]_ ;
  assign \new_[64478]_  = ~A232 & A203;
  assign \new_[64481]_  = ~A234 & A233;
  assign \new_[64482]_  = \new_[64481]_  & \new_[64478]_ ;
  assign \new_[64483]_  = \new_[64482]_  & \new_[64475]_ ;
  assign \new_[64486]_  = A236 & ~A235;
  assign \new_[64489]_  = ~A269 & ~A267;
  assign \new_[64490]_  = \new_[64489]_  & \new_[64486]_ ;
  assign \new_[64493]_  = A299 & ~A298;
  assign \new_[64497]_  = A302 & ~A301;
  assign \new_[64498]_  = ~A300 & \new_[64497]_ ;
  assign \new_[64499]_  = \new_[64498]_  & \new_[64493]_ ;
  assign \new_[64500]_  = \new_[64499]_  & \new_[64490]_ ;
  assign \new_[64503]_  = ~A200 & A199;
  assign \new_[64506]_  = ~A202 & ~A201;
  assign \new_[64507]_  = \new_[64506]_  & \new_[64503]_ ;
  assign \new_[64510]_  = ~A232 & A203;
  assign \new_[64513]_  = ~A234 & A233;
  assign \new_[64514]_  = \new_[64513]_  & \new_[64510]_ ;
  assign \new_[64515]_  = \new_[64514]_  & \new_[64507]_ ;
  assign \new_[64518]_  = A236 & ~A235;
  assign \new_[64521]_  = A266 & A265;
  assign \new_[64522]_  = \new_[64521]_  & \new_[64518]_ ;
  assign \new_[64525]_  = ~A299 & A298;
  assign \new_[64529]_  = A302 & ~A301;
  assign \new_[64530]_  = ~A300 & \new_[64529]_ ;
  assign \new_[64531]_  = \new_[64530]_  & \new_[64525]_ ;
  assign \new_[64532]_  = \new_[64531]_  & \new_[64522]_ ;
  assign \new_[64535]_  = ~A200 & A199;
  assign \new_[64538]_  = ~A202 & ~A201;
  assign \new_[64539]_  = \new_[64538]_  & \new_[64535]_ ;
  assign \new_[64542]_  = ~A232 & A203;
  assign \new_[64545]_  = ~A234 & A233;
  assign \new_[64546]_  = \new_[64545]_  & \new_[64542]_ ;
  assign \new_[64547]_  = \new_[64546]_  & \new_[64539]_ ;
  assign \new_[64550]_  = A236 & ~A235;
  assign \new_[64553]_  = A266 & A265;
  assign \new_[64554]_  = \new_[64553]_  & \new_[64550]_ ;
  assign \new_[64557]_  = A299 & ~A298;
  assign \new_[64561]_  = A302 & ~A301;
  assign \new_[64562]_  = ~A300 & \new_[64561]_ ;
  assign \new_[64563]_  = \new_[64562]_  & \new_[64557]_ ;
  assign \new_[64564]_  = \new_[64563]_  & \new_[64554]_ ;
  assign \new_[64567]_  = ~A200 & A199;
  assign \new_[64570]_  = ~A202 & ~A201;
  assign \new_[64571]_  = \new_[64570]_  & \new_[64567]_ ;
  assign \new_[64574]_  = ~A232 & A203;
  assign \new_[64577]_  = ~A234 & A233;
  assign \new_[64578]_  = \new_[64577]_  & \new_[64574]_ ;
  assign \new_[64579]_  = \new_[64578]_  & \new_[64571]_ ;
  assign \new_[64582]_  = A236 & ~A235;
  assign \new_[64585]_  = ~A266 & ~A265;
  assign \new_[64586]_  = \new_[64585]_  & \new_[64582]_ ;
  assign \new_[64589]_  = ~A299 & A298;
  assign \new_[64593]_  = A302 & ~A301;
  assign \new_[64594]_  = ~A300 & \new_[64593]_ ;
  assign \new_[64595]_  = \new_[64594]_  & \new_[64589]_ ;
  assign \new_[64596]_  = \new_[64595]_  & \new_[64586]_ ;
  assign \new_[64599]_  = ~A200 & A199;
  assign \new_[64602]_  = ~A202 & ~A201;
  assign \new_[64603]_  = \new_[64602]_  & \new_[64599]_ ;
  assign \new_[64606]_  = ~A232 & A203;
  assign \new_[64609]_  = ~A234 & A233;
  assign \new_[64610]_  = \new_[64609]_  & \new_[64606]_ ;
  assign \new_[64611]_  = \new_[64610]_  & \new_[64603]_ ;
  assign \new_[64614]_  = A236 & ~A235;
  assign \new_[64617]_  = ~A266 & ~A265;
  assign \new_[64618]_  = \new_[64617]_  & \new_[64614]_ ;
  assign \new_[64621]_  = A299 & ~A298;
  assign \new_[64625]_  = A302 & ~A301;
  assign \new_[64626]_  = ~A300 & \new_[64625]_ ;
  assign \new_[64627]_  = \new_[64626]_  & \new_[64621]_ ;
  assign \new_[64628]_  = \new_[64627]_  & \new_[64618]_ ;
  assign \new_[64631]_  = ~A200 & A199;
  assign \new_[64634]_  = ~A202 & ~A201;
  assign \new_[64635]_  = \new_[64634]_  & \new_[64631]_ ;
  assign \new_[64638]_  = A232 & A203;
  assign \new_[64641]_  = A234 & ~A233;
  assign \new_[64642]_  = \new_[64641]_  & \new_[64638]_ ;
  assign \new_[64643]_  = \new_[64642]_  & \new_[64635]_ ;
  assign \new_[64646]_  = A267 & A235;
  assign \new_[64649]_  = A269 & ~A268;
  assign \new_[64650]_  = \new_[64649]_  & \new_[64646]_ ;
  assign \new_[64653]_  = ~A299 & A298;
  assign \new_[64657]_  = A302 & ~A301;
  assign \new_[64658]_  = ~A300 & \new_[64657]_ ;
  assign \new_[64659]_  = \new_[64658]_  & \new_[64653]_ ;
  assign \new_[64660]_  = \new_[64659]_  & \new_[64650]_ ;
  assign \new_[64663]_  = ~A200 & A199;
  assign \new_[64666]_  = ~A202 & ~A201;
  assign \new_[64667]_  = \new_[64666]_  & \new_[64663]_ ;
  assign \new_[64670]_  = A232 & A203;
  assign \new_[64673]_  = A234 & ~A233;
  assign \new_[64674]_  = \new_[64673]_  & \new_[64670]_ ;
  assign \new_[64675]_  = \new_[64674]_  & \new_[64667]_ ;
  assign \new_[64678]_  = A267 & A235;
  assign \new_[64681]_  = A269 & ~A268;
  assign \new_[64682]_  = \new_[64681]_  & \new_[64678]_ ;
  assign \new_[64685]_  = A299 & ~A298;
  assign \new_[64689]_  = A302 & ~A301;
  assign \new_[64690]_  = ~A300 & \new_[64689]_ ;
  assign \new_[64691]_  = \new_[64690]_  & \new_[64685]_ ;
  assign \new_[64692]_  = \new_[64691]_  & \new_[64682]_ ;
  assign \new_[64695]_  = ~A200 & A199;
  assign \new_[64698]_  = ~A202 & ~A201;
  assign \new_[64699]_  = \new_[64698]_  & \new_[64695]_ ;
  assign \new_[64702]_  = A232 & A203;
  assign \new_[64705]_  = A234 & ~A233;
  assign \new_[64706]_  = \new_[64705]_  & \new_[64702]_ ;
  assign \new_[64707]_  = \new_[64706]_  & \new_[64699]_ ;
  assign \new_[64710]_  = A267 & ~A236;
  assign \new_[64713]_  = A269 & ~A268;
  assign \new_[64714]_  = \new_[64713]_  & \new_[64710]_ ;
  assign \new_[64717]_  = ~A299 & A298;
  assign \new_[64721]_  = A302 & ~A301;
  assign \new_[64722]_  = ~A300 & \new_[64721]_ ;
  assign \new_[64723]_  = \new_[64722]_  & \new_[64717]_ ;
  assign \new_[64724]_  = \new_[64723]_  & \new_[64714]_ ;
  assign \new_[64727]_  = ~A200 & A199;
  assign \new_[64730]_  = ~A202 & ~A201;
  assign \new_[64731]_  = \new_[64730]_  & \new_[64727]_ ;
  assign \new_[64734]_  = A232 & A203;
  assign \new_[64737]_  = A234 & ~A233;
  assign \new_[64738]_  = \new_[64737]_  & \new_[64734]_ ;
  assign \new_[64739]_  = \new_[64738]_  & \new_[64731]_ ;
  assign \new_[64742]_  = A267 & ~A236;
  assign \new_[64745]_  = A269 & ~A268;
  assign \new_[64746]_  = \new_[64745]_  & \new_[64742]_ ;
  assign \new_[64749]_  = A299 & ~A298;
  assign \new_[64753]_  = A302 & ~A301;
  assign \new_[64754]_  = ~A300 & \new_[64753]_ ;
  assign \new_[64755]_  = \new_[64754]_  & \new_[64749]_ ;
  assign \new_[64756]_  = \new_[64755]_  & \new_[64746]_ ;
  assign \new_[64759]_  = ~A200 & A199;
  assign \new_[64762]_  = ~A202 & ~A201;
  assign \new_[64763]_  = \new_[64762]_  & \new_[64759]_ ;
  assign \new_[64766]_  = A232 & A203;
  assign \new_[64769]_  = ~A234 & ~A233;
  assign \new_[64770]_  = \new_[64769]_  & \new_[64766]_ ;
  assign \new_[64771]_  = \new_[64770]_  & \new_[64763]_ ;
  assign \new_[64774]_  = A236 & ~A235;
  assign \new_[64777]_  = ~A268 & A267;
  assign \new_[64778]_  = \new_[64777]_  & \new_[64774]_ ;
  assign \new_[64781]_  = A298 & A269;
  assign \new_[64785]_  = A301 & A300;
  assign \new_[64786]_  = ~A299 & \new_[64785]_ ;
  assign \new_[64787]_  = \new_[64786]_  & \new_[64781]_ ;
  assign \new_[64788]_  = \new_[64787]_  & \new_[64778]_ ;
  assign \new_[64791]_  = ~A200 & A199;
  assign \new_[64794]_  = ~A202 & ~A201;
  assign \new_[64795]_  = \new_[64794]_  & \new_[64791]_ ;
  assign \new_[64798]_  = A232 & A203;
  assign \new_[64801]_  = ~A234 & ~A233;
  assign \new_[64802]_  = \new_[64801]_  & \new_[64798]_ ;
  assign \new_[64803]_  = \new_[64802]_  & \new_[64795]_ ;
  assign \new_[64806]_  = A236 & ~A235;
  assign \new_[64809]_  = ~A268 & A267;
  assign \new_[64810]_  = \new_[64809]_  & \new_[64806]_ ;
  assign \new_[64813]_  = A298 & A269;
  assign \new_[64817]_  = ~A302 & A300;
  assign \new_[64818]_  = ~A299 & \new_[64817]_ ;
  assign \new_[64819]_  = \new_[64818]_  & \new_[64813]_ ;
  assign \new_[64820]_  = \new_[64819]_  & \new_[64810]_ ;
  assign \new_[64823]_  = ~A200 & A199;
  assign \new_[64826]_  = ~A202 & ~A201;
  assign \new_[64827]_  = \new_[64826]_  & \new_[64823]_ ;
  assign \new_[64830]_  = A232 & A203;
  assign \new_[64833]_  = ~A234 & ~A233;
  assign \new_[64834]_  = \new_[64833]_  & \new_[64830]_ ;
  assign \new_[64835]_  = \new_[64834]_  & \new_[64827]_ ;
  assign \new_[64838]_  = A236 & ~A235;
  assign \new_[64841]_  = ~A268 & A267;
  assign \new_[64842]_  = \new_[64841]_  & \new_[64838]_ ;
  assign \new_[64845]_  = ~A298 & A269;
  assign \new_[64849]_  = A301 & A300;
  assign \new_[64850]_  = A299 & \new_[64849]_ ;
  assign \new_[64851]_  = \new_[64850]_  & \new_[64845]_ ;
  assign \new_[64852]_  = \new_[64851]_  & \new_[64842]_ ;
  assign \new_[64855]_  = ~A200 & A199;
  assign \new_[64858]_  = ~A202 & ~A201;
  assign \new_[64859]_  = \new_[64858]_  & \new_[64855]_ ;
  assign \new_[64862]_  = A232 & A203;
  assign \new_[64865]_  = ~A234 & ~A233;
  assign \new_[64866]_  = \new_[64865]_  & \new_[64862]_ ;
  assign \new_[64867]_  = \new_[64866]_  & \new_[64859]_ ;
  assign \new_[64870]_  = A236 & ~A235;
  assign \new_[64873]_  = ~A268 & A267;
  assign \new_[64874]_  = \new_[64873]_  & \new_[64870]_ ;
  assign \new_[64877]_  = ~A298 & A269;
  assign \new_[64881]_  = ~A302 & A300;
  assign \new_[64882]_  = A299 & \new_[64881]_ ;
  assign \new_[64883]_  = \new_[64882]_  & \new_[64877]_ ;
  assign \new_[64884]_  = \new_[64883]_  & \new_[64874]_ ;
  assign \new_[64887]_  = ~A200 & A199;
  assign \new_[64890]_  = ~A202 & ~A201;
  assign \new_[64891]_  = \new_[64890]_  & \new_[64887]_ ;
  assign \new_[64894]_  = A232 & A203;
  assign \new_[64897]_  = ~A234 & ~A233;
  assign \new_[64898]_  = \new_[64897]_  & \new_[64894]_ ;
  assign \new_[64899]_  = \new_[64898]_  & \new_[64891]_ ;
  assign \new_[64902]_  = A236 & ~A235;
  assign \new_[64905]_  = A268 & ~A267;
  assign \new_[64906]_  = \new_[64905]_  & \new_[64902]_ ;
  assign \new_[64909]_  = ~A299 & A298;
  assign \new_[64913]_  = A302 & ~A301;
  assign \new_[64914]_  = ~A300 & \new_[64913]_ ;
  assign \new_[64915]_  = \new_[64914]_  & \new_[64909]_ ;
  assign \new_[64916]_  = \new_[64915]_  & \new_[64906]_ ;
  assign \new_[64919]_  = ~A200 & A199;
  assign \new_[64922]_  = ~A202 & ~A201;
  assign \new_[64923]_  = \new_[64922]_  & \new_[64919]_ ;
  assign \new_[64926]_  = A232 & A203;
  assign \new_[64929]_  = ~A234 & ~A233;
  assign \new_[64930]_  = \new_[64929]_  & \new_[64926]_ ;
  assign \new_[64931]_  = \new_[64930]_  & \new_[64923]_ ;
  assign \new_[64934]_  = A236 & ~A235;
  assign \new_[64937]_  = A268 & ~A267;
  assign \new_[64938]_  = \new_[64937]_  & \new_[64934]_ ;
  assign \new_[64941]_  = A299 & ~A298;
  assign \new_[64945]_  = A302 & ~A301;
  assign \new_[64946]_  = ~A300 & \new_[64945]_ ;
  assign \new_[64947]_  = \new_[64946]_  & \new_[64941]_ ;
  assign \new_[64948]_  = \new_[64947]_  & \new_[64938]_ ;
  assign \new_[64951]_  = ~A200 & A199;
  assign \new_[64954]_  = ~A202 & ~A201;
  assign \new_[64955]_  = \new_[64954]_  & \new_[64951]_ ;
  assign \new_[64958]_  = A232 & A203;
  assign \new_[64961]_  = ~A234 & ~A233;
  assign \new_[64962]_  = \new_[64961]_  & \new_[64958]_ ;
  assign \new_[64963]_  = \new_[64962]_  & \new_[64955]_ ;
  assign \new_[64966]_  = A236 & ~A235;
  assign \new_[64969]_  = ~A269 & ~A267;
  assign \new_[64970]_  = \new_[64969]_  & \new_[64966]_ ;
  assign \new_[64973]_  = ~A299 & A298;
  assign \new_[64977]_  = A302 & ~A301;
  assign \new_[64978]_  = ~A300 & \new_[64977]_ ;
  assign \new_[64979]_  = \new_[64978]_  & \new_[64973]_ ;
  assign \new_[64980]_  = \new_[64979]_  & \new_[64970]_ ;
  assign \new_[64983]_  = ~A200 & A199;
  assign \new_[64986]_  = ~A202 & ~A201;
  assign \new_[64987]_  = \new_[64986]_  & \new_[64983]_ ;
  assign \new_[64990]_  = A232 & A203;
  assign \new_[64993]_  = ~A234 & ~A233;
  assign \new_[64994]_  = \new_[64993]_  & \new_[64990]_ ;
  assign \new_[64995]_  = \new_[64994]_  & \new_[64987]_ ;
  assign \new_[64998]_  = A236 & ~A235;
  assign \new_[65001]_  = ~A269 & ~A267;
  assign \new_[65002]_  = \new_[65001]_  & \new_[64998]_ ;
  assign \new_[65005]_  = A299 & ~A298;
  assign \new_[65009]_  = A302 & ~A301;
  assign \new_[65010]_  = ~A300 & \new_[65009]_ ;
  assign \new_[65011]_  = \new_[65010]_  & \new_[65005]_ ;
  assign \new_[65012]_  = \new_[65011]_  & \new_[65002]_ ;
  assign \new_[65015]_  = ~A200 & A199;
  assign \new_[65018]_  = ~A202 & ~A201;
  assign \new_[65019]_  = \new_[65018]_  & \new_[65015]_ ;
  assign \new_[65022]_  = A232 & A203;
  assign \new_[65025]_  = ~A234 & ~A233;
  assign \new_[65026]_  = \new_[65025]_  & \new_[65022]_ ;
  assign \new_[65027]_  = \new_[65026]_  & \new_[65019]_ ;
  assign \new_[65030]_  = A236 & ~A235;
  assign \new_[65033]_  = A266 & A265;
  assign \new_[65034]_  = \new_[65033]_  & \new_[65030]_ ;
  assign \new_[65037]_  = ~A299 & A298;
  assign \new_[65041]_  = A302 & ~A301;
  assign \new_[65042]_  = ~A300 & \new_[65041]_ ;
  assign \new_[65043]_  = \new_[65042]_  & \new_[65037]_ ;
  assign \new_[65044]_  = \new_[65043]_  & \new_[65034]_ ;
  assign \new_[65047]_  = ~A200 & A199;
  assign \new_[65050]_  = ~A202 & ~A201;
  assign \new_[65051]_  = \new_[65050]_  & \new_[65047]_ ;
  assign \new_[65054]_  = A232 & A203;
  assign \new_[65057]_  = ~A234 & ~A233;
  assign \new_[65058]_  = \new_[65057]_  & \new_[65054]_ ;
  assign \new_[65059]_  = \new_[65058]_  & \new_[65051]_ ;
  assign \new_[65062]_  = A236 & ~A235;
  assign \new_[65065]_  = A266 & A265;
  assign \new_[65066]_  = \new_[65065]_  & \new_[65062]_ ;
  assign \new_[65069]_  = A299 & ~A298;
  assign \new_[65073]_  = A302 & ~A301;
  assign \new_[65074]_  = ~A300 & \new_[65073]_ ;
  assign \new_[65075]_  = \new_[65074]_  & \new_[65069]_ ;
  assign \new_[65076]_  = \new_[65075]_  & \new_[65066]_ ;
  assign \new_[65079]_  = ~A200 & A199;
  assign \new_[65082]_  = ~A202 & ~A201;
  assign \new_[65083]_  = \new_[65082]_  & \new_[65079]_ ;
  assign \new_[65086]_  = A232 & A203;
  assign \new_[65089]_  = ~A234 & ~A233;
  assign \new_[65090]_  = \new_[65089]_  & \new_[65086]_ ;
  assign \new_[65091]_  = \new_[65090]_  & \new_[65083]_ ;
  assign \new_[65094]_  = A236 & ~A235;
  assign \new_[65097]_  = ~A266 & ~A265;
  assign \new_[65098]_  = \new_[65097]_  & \new_[65094]_ ;
  assign \new_[65101]_  = ~A299 & A298;
  assign \new_[65105]_  = A302 & ~A301;
  assign \new_[65106]_  = ~A300 & \new_[65105]_ ;
  assign \new_[65107]_  = \new_[65106]_  & \new_[65101]_ ;
  assign \new_[65108]_  = \new_[65107]_  & \new_[65098]_ ;
  assign \new_[65111]_  = ~A200 & A199;
  assign \new_[65114]_  = ~A202 & ~A201;
  assign \new_[65115]_  = \new_[65114]_  & \new_[65111]_ ;
  assign \new_[65118]_  = A232 & A203;
  assign \new_[65121]_  = ~A234 & ~A233;
  assign \new_[65122]_  = \new_[65121]_  & \new_[65118]_ ;
  assign \new_[65123]_  = \new_[65122]_  & \new_[65115]_ ;
  assign \new_[65126]_  = A236 & ~A235;
  assign \new_[65129]_  = ~A266 & ~A265;
  assign \new_[65130]_  = \new_[65129]_  & \new_[65126]_ ;
  assign \new_[65133]_  = A299 & ~A298;
  assign \new_[65137]_  = A302 & ~A301;
  assign \new_[65138]_  = ~A300 & \new_[65137]_ ;
  assign \new_[65139]_  = \new_[65138]_  & \new_[65133]_ ;
  assign \new_[65140]_  = \new_[65139]_  & \new_[65130]_ ;
  assign \new_[65143]_  = A168 & A170;
  assign \new_[65146]_  = ~A166 & A167;
  assign \new_[65147]_  = \new_[65146]_  & \new_[65143]_ ;
  assign \new_[65150]_  = A233 & ~A232;
  assign \new_[65153]_  = ~A235 & ~A234;
  assign \new_[65154]_  = \new_[65153]_  & \new_[65150]_ ;
  assign \new_[65155]_  = \new_[65154]_  & \new_[65147]_ ;
  assign \new_[65158]_  = A267 & A236;
  assign \new_[65161]_  = A269 & ~A268;
  assign \new_[65162]_  = \new_[65161]_  & \new_[65158]_ ;
  assign \new_[65165]_  = ~A299 & A298;
  assign \new_[65169]_  = A302 & ~A301;
  assign \new_[65170]_  = ~A300 & \new_[65169]_ ;
  assign \new_[65171]_  = \new_[65170]_  & \new_[65165]_ ;
  assign \new_[65172]_  = \new_[65171]_  & \new_[65162]_ ;
  assign \new_[65175]_  = A168 & A170;
  assign \new_[65178]_  = ~A166 & A167;
  assign \new_[65179]_  = \new_[65178]_  & \new_[65175]_ ;
  assign \new_[65182]_  = A233 & ~A232;
  assign \new_[65185]_  = ~A235 & ~A234;
  assign \new_[65186]_  = \new_[65185]_  & \new_[65182]_ ;
  assign \new_[65187]_  = \new_[65186]_  & \new_[65179]_ ;
  assign \new_[65190]_  = A267 & A236;
  assign \new_[65193]_  = A269 & ~A268;
  assign \new_[65194]_  = \new_[65193]_  & \new_[65190]_ ;
  assign \new_[65197]_  = A299 & ~A298;
  assign \new_[65201]_  = A302 & ~A301;
  assign \new_[65202]_  = ~A300 & \new_[65201]_ ;
  assign \new_[65203]_  = \new_[65202]_  & \new_[65197]_ ;
  assign \new_[65204]_  = \new_[65203]_  & \new_[65194]_ ;
  assign \new_[65207]_  = A168 & A170;
  assign \new_[65210]_  = ~A166 & A167;
  assign \new_[65211]_  = \new_[65210]_  & \new_[65207]_ ;
  assign \new_[65214]_  = ~A233 & A232;
  assign \new_[65217]_  = ~A235 & ~A234;
  assign \new_[65218]_  = \new_[65217]_  & \new_[65214]_ ;
  assign \new_[65219]_  = \new_[65218]_  & \new_[65211]_ ;
  assign \new_[65222]_  = A267 & A236;
  assign \new_[65225]_  = A269 & ~A268;
  assign \new_[65226]_  = \new_[65225]_  & \new_[65222]_ ;
  assign \new_[65229]_  = ~A299 & A298;
  assign \new_[65233]_  = A302 & ~A301;
  assign \new_[65234]_  = ~A300 & \new_[65233]_ ;
  assign \new_[65235]_  = \new_[65234]_  & \new_[65229]_ ;
  assign \new_[65236]_  = \new_[65235]_  & \new_[65226]_ ;
  assign \new_[65239]_  = A168 & A170;
  assign \new_[65242]_  = ~A166 & A167;
  assign \new_[65243]_  = \new_[65242]_  & \new_[65239]_ ;
  assign \new_[65246]_  = ~A233 & A232;
  assign \new_[65249]_  = ~A235 & ~A234;
  assign \new_[65250]_  = \new_[65249]_  & \new_[65246]_ ;
  assign \new_[65251]_  = \new_[65250]_  & \new_[65243]_ ;
  assign \new_[65254]_  = A267 & A236;
  assign \new_[65257]_  = A269 & ~A268;
  assign \new_[65258]_  = \new_[65257]_  & \new_[65254]_ ;
  assign \new_[65261]_  = A299 & ~A298;
  assign \new_[65265]_  = A302 & ~A301;
  assign \new_[65266]_  = ~A300 & \new_[65265]_ ;
  assign \new_[65267]_  = \new_[65266]_  & \new_[65261]_ ;
  assign \new_[65268]_  = \new_[65267]_  & \new_[65258]_ ;
  assign \new_[65271]_  = A168 & A170;
  assign \new_[65274]_  = A166 & ~A167;
  assign \new_[65275]_  = \new_[65274]_  & \new_[65271]_ ;
  assign \new_[65278]_  = A233 & ~A232;
  assign \new_[65281]_  = ~A235 & ~A234;
  assign \new_[65282]_  = \new_[65281]_  & \new_[65278]_ ;
  assign \new_[65283]_  = \new_[65282]_  & \new_[65275]_ ;
  assign \new_[65286]_  = A267 & A236;
  assign \new_[65289]_  = A269 & ~A268;
  assign \new_[65290]_  = \new_[65289]_  & \new_[65286]_ ;
  assign \new_[65293]_  = ~A299 & A298;
  assign \new_[65297]_  = A302 & ~A301;
  assign \new_[65298]_  = ~A300 & \new_[65297]_ ;
  assign \new_[65299]_  = \new_[65298]_  & \new_[65293]_ ;
  assign \new_[65300]_  = \new_[65299]_  & \new_[65290]_ ;
  assign \new_[65303]_  = A168 & A170;
  assign \new_[65306]_  = A166 & ~A167;
  assign \new_[65307]_  = \new_[65306]_  & \new_[65303]_ ;
  assign \new_[65310]_  = A233 & ~A232;
  assign \new_[65313]_  = ~A235 & ~A234;
  assign \new_[65314]_  = \new_[65313]_  & \new_[65310]_ ;
  assign \new_[65315]_  = \new_[65314]_  & \new_[65307]_ ;
  assign \new_[65318]_  = A267 & A236;
  assign \new_[65321]_  = A269 & ~A268;
  assign \new_[65322]_  = \new_[65321]_  & \new_[65318]_ ;
  assign \new_[65325]_  = A299 & ~A298;
  assign \new_[65329]_  = A302 & ~A301;
  assign \new_[65330]_  = ~A300 & \new_[65329]_ ;
  assign \new_[65331]_  = \new_[65330]_  & \new_[65325]_ ;
  assign \new_[65332]_  = \new_[65331]_  & \new_[65322]_ ;
  assign \new_[65335]_  = A168 & A170;
  assign \new_[65338]_  = A166 & ~A167;
  assign \new_[65339]_  = \new_[65338]_  & \new_[65335]_ ;
  assign \new_[65342]_  = ~A233 & A232;
  assign \new_[65345]_  = ~A235 & ~A234;
  assign \new_[65346]_  = \new_[65345]_  & \new_[65342]_ ;
  assign \new_[65347]_  = \new_[65346]_  & \new_[65339]_ ;
  assign \new_[65350]_  = A267 & A236;
  assign \new_[65353]_  = A269 & ~A268;
  assign \new_[65354]_  = \new_[65353]_  & \new_[65350]_ ;
  assign \new_[65357]_  = ~A299 & A298;
  assign \new_[65361]_  = A302 & ~A301;
  assign \new_[65362]_  = ~A300 & \new_[65361]_ ;
  assign \new_[65363]_  = \new_[65362]_  & \new_[65357]_ ;
  assign \new_[65364]_  = \new_[65363]_  & \new_[65354]_ ;
  assign \new_[65367]_  = A168 & A170;
  assign \new_[65370]_  = A166 & ~A167;
  assign \new_[65371]_  = \new_[65370]_  & \new_[65367]_ ;
  assign \new_[65374]_  = ~A233 & A232;
  assign \new_[65377]_  = ~A235 & ~A234;
  assign \new_[65378]_  = \new_[65377]_  & \new_[65374]_ ;
  assign \new_[65379]_  = \new_[65378]_  & \new_[65371]_ ;
  assign \new_[65382]_  = A267 & A236;
  assign \new_[65385]_  = A269 & ~A268;
  assign \new_[65386]_  = \new_[65385]_  & \new_[65382]_ ;
  assign \new_[65389]_  = A299 & ~A298;
  assign \new_[65393]_  = A302 & ~A301;
  assign \new_[65394]_  = ~A300 & \new_[65393]_ ;
  assign \new_[65395]_  = \new_[65394]_  & \new_[65389]_ ;
  assign \new_[65396]_  = \new_[65395]_  & \new_[65386]_ ;
  assign \new_[65399]_  = A168 & A169;
  assign \new_[65402]_  = ~A166 & A167;
  assign \new_[65403]_  = \new_[65402]_  & \new_[65399]_ ;
  assign \new_[65406]_  = A233 & ~A232;
  assign \new_[65409]_  = ~A235 & ~A234;
  assign \new_[65410]_  = \new_[65409]_  & \new_[65406]_ ;
  assign \new_[65411]_  = \new_[65410]_  & \new_[65403]_ ;
  assign \new_[65414]_  = A267 & A236;
  assign \new_[65417]_  = A269 & ~A268;
  assign \new_[65418]_  = \new_[65417]_  & \new_[65414]_ ;
  assign \new_[65421]_  = ~A299 & A298;
  assign \new_[65425]_  = A302 & ~A301;
  assign \new_[65426]_  = ~A300 & \new_[65425]_ ;
  assign \new_[65427]_  = \new_[65426]_  & \new_[65421]_ ;
  assign \new_[65428]_  = \new_[65427]_  & \new_[65418]_ ;
  assign \new_[65431]_  = A168 & A169;
  assign \new_[65434]_  = ~A166 & A167;
  assign \new_[65435]_  = \new_[65434]_  & \new_[65431]_ ;
  assign \new_[65438]_  = A233 & ~A232;
  assign \new_[65441]_  = ~A235 & ~A234;
  assign \new_[65442]_  = \new_[65441]_  & \new_[65438]_ ;
  assign \new_[65443]_  = \new_[65442]_  & \new_[65435]_ ;
  assign \new_[65446]_  = A267 & A236;
  assign \new_[65449]_  = A269 & ~A268;
  assign \new_[65450]_  = \new_[65449]_  & \new_[65446]_ ;
  assign \new_[65453]_  = A299 & ~A298;
  assign \new_[65457]_  = A302 & ~A301;
  assign \new_[65458]_  = ~A300 & \new_[65457]_ ;
  assign \new_[65459]_  = \new_[65458]_  & \new_[65453]_ ;
  assign \new_[65460]_  = \new_[65459]_  & \new_[65450]_ ;
  assign \new_[65463]_  = A168 & A169;
  assign \new_[65466]_  = ~A166 & A167;
  assign \new_[65467]_  = \new_[65466]_  & \new_[65463]_ ;
  assign \new_[65470]_  = ~A233 & A232;
  assign \new_[65473]_  = ~A235 & ~A234;
  assign \new_[65474]_  = \new_[65473]_  & \new_[65470]_ ;
  assign \new_[65475]_  = \new_[65474]_  & \new_[65467]_ ;
  assign \new_[65478]_  = A267 & A236;
  assign \new_[65481]_  = A269 & ~A268;
  assign \new_[65482]_  = \new_[65481]_  & \new_[65478]_ ;
  assign \new_[65485]_  = ~A299 & A298;
  assign \new_[65489]_  = A302 & ~A301;
  assign \new_[65490]_  = ~A300 & \new_[65489]_ ;
  assign \new_[65491]_  = \new_[65490]_  & \new_[65485]_ ;
  assign \new_[65492]_  = \new_[65491]_  & \new_[65482]_ ;
  assign \new_[65495]_  = A168 & A169;
  assign \new_[65498]_  = ~A166 & A167;
  assign \new_[65499]_  = \new_[65498]_  & \new_[65495]_ ;
  assign \new_[65502]_  = ~A233 & A232;
  assign \new_[65505]_  = ~A235 & ~A234;
  assign \new_[65506]_  = \new_[65505]_  & \new_[65502]_ ;
  assign \new_[65507]_  = \new_[65506]_  & \new_[65499]_ ;
  assign \new_[65510]_  = A267 & A236;
  assign \new_[65513]_  = A269 & ~A268;
  assign \new_[65514]_  = \new_[65513]_  & \new_[65510]_ ;
  assign \new_[65517]_  = A299 & ~A298;
  assign \new_[65521]_  = A302 & ~A301;
  assign \new_[65522]_  = ~A300 & \new_[65521]_ ;
  assign \new_[65523]_  = \new_[65522]_  & \new_[65517]_ ;
  assign \new_[65524]_  = \new_[65523]_  & \new_[65514]_ ;
  assign \new_[65527]_  = A168 & A169;
  assign \new_[65530]_  = A166 & ~A167;
  assign \new_[65531]_  = \new_[65530]_  & \new_[65527]_ ;
  assign \new_[65534]_  = A233 & ~A232;
  assign \new_[65537]_  = ~A235 & ~A234;
  assign \new_[65538]_  = \new_[65537]_  & \new_[65534]_ ;
  assign \new_[65539]_  = \new_[65538]_  & \new_[65531]_ ;
  assign \new_[65542]_  = A267 & A236;
  assign \new_[65545]_  = A269 & ~A268;
  assign \new_[65546]_  = \new_[65545]_  & \new_[65542]_ ;
  assign \new_[65549]_  = ~A299 & A298;
  assign \new_[65553]_  = A302 & ~A301;
  assign \new_[65554]_  = ~A300 & \new_[65553]_ ;
  assign \new_[65555]_  = \new_[65554]_  & \new_[65549]_ ;
  assign \new_[65556]_  = \new_[65555]_  & \new_[65546]_ ;
  assign \new_[65559]_  = A168 & A169;
  assign \new_[65562]_  = A166 & ~A167;
  assign \new_[65563]_  = \new_[65562]_  & \new_[65559]_ ;
  assign \new_[65566]_  = A233 & ~A232;
  assign \new_[65569]_  = ~A235 & ~A234;
  assign \new_[65570]_  = \new_[65569]_  & \new_[65566]_ ;
  assign \new_[65571]_  = \new_[65570]_  & \new_[65563]_ ;
  assign \new_[65574]_  = A267 & A236;
  assign \new_[65577]_  = A269 & ~A268;
  assign \new_[65578]_  = \new_[65577]_  & \new_[65574]_ ;
  assign \new_[65581]_  = A299 & ~A298;
  assign \new_[65585]_  = A302 & ~A301;
  assign \new_[65586]_  = ~A300 & \new_[65585]_ ;
  assign \new_[65587]_  = \new_[65586]_  & \new_[65581]_ ;
  assign \new_[65588]_  = \new_[65587]_  & \new_[65578]_ ;
  assign \new_[65591]_  = A168 & A169;
  assign \new_[65594]_  = A166 & ~A167;
  assign \new_[65595]_  = \new_[65594]_  & \new_[65591]_ ;
  assign \new_[65598]_  = ~A233 & A232;
  assign \new_[65601]_  = ~A235 & ~A234;
  assign \new_[65602]_  = \new_[65601]_  & \new_[65598]_ ;
  assign \new_[65603]_  = \new_[65602]_  & \new_[65595]_ ;
  assign \new_[65606]_  = A267 & A236;
  assign \new_[65609]_  = A269 & ~A268;
  assign \new_[65610]_  = \new_[65609]_  & \new_[65606]_ ;
  assign \new_[65613]_  = ~A299 & A298;
  assign \new_[65617]_  = A302 & ~A301;
  assign \new_[65618]_  = ~A300 & \new_[65617]_ ;
  assign \new_[65619]_  = \new_[65618]_  & \new_[65613]_ ;
  assign \new_[65620]_  = \new_[65619]_  & \new_[65610]_ ;
  assign \new_[65623]_  = A168 & A169;
  assign \new_[65626]_  = A166 & ~A167;
  assign \new_[65627]_  = \new_[65626]_  & \new_[65623]_ ;
  assign \new_[65630]_  = ~A233 & A232;
  assign \new_[65633]_  = ~A235 & ~A234;
  assign \new_[65634]_  = \new_[65633]_  & \new_[65630]_ ;
  assign \new_[65635]_  = \new_[65634]_  & \new_[65627]_ ;
  assign \new_[65638]_  = A267 & A236;
  assign \new_[65641]_  = A269 & ~A268;
  assign \new_[65642]_  = \new_[65641]_  & \new_[65638]_ ;
  assign \new_[65645]_  = A299 & ~A298;
  assign \new_[65649]_  = A302 & ~A301;
  assign \new_[65650]_  = ~A300 & \new_[65649]_ ;
  assign \new_[65651]_  = \new_[65650]_  & \new_[65645]_ ;
  assign \new_[65652]_  = \new_[65651]_  & \new_[65642]_ ;
  assign \new_[65655]_  = ~A169 & ~A170;
  assign \new_[65658]_  = A167 & ~A168;
  assign \new_[65659]_  = \new_[65658]_  & \new_[65655]_ ;
  assign \new_[65662]_  = ~A232 & ~A166;
  assign \new_[65665]_  = A234 & A233;
  assign \new_[65666]_  = \new_[65665]_  & \new_[65662]_ ;
  assign \new_[65667]_  = \new_[65666]_  & \new_[65659]_ ;
  assign \new_[65670]_  = A267 & A235;
  assign \new_[65673]_  = A269 & ~A268;
  assign \new_[65674]_  = \new_[65673]_  & \new_[65670]_ ;
  assign \new_[65677]_  = ~A299 & A298;
  assign \new_[65681]_  = A302 & ~A301;
  assign \new_[65682]_  = ~A300 & \new_[65681]_ ;
  assign \new_[65683]_  = \new_[65682]_  & \new_[65677]_ ;
  assign \new_[65684]_  = \new_[65683]_  & \new_[65674]_ ;
  assign \new_[65687]_  = ~A169 & ~A170;
  assign \new_[65690]_  = A167 & ~A168;
  assign \new_[65691]_  = \new_[65690]_  & \new_[65687]_ ;
  assign \new_[65694]_  = ~A232 & ~A166;
  assign \new_[65697]_  = A234 & A233;
  assign \new_[65698]_  = \new_[65697]_  & \new_[65694]_ ;
  assign \new_[65699]_  = \new_[65698]_  & \new_[65691]_ ;
  assign \new_[65702]_  = A267 & A235;
  assign \new_[65705]_  = A269 & ~A268;
  assign \new_[65706]_  = \new_[65705]_  & \new_[65702]_ ;
  assign \new_[65709]_  = A299 & ~A298;
  assign \new_[65713]_  = A302 & ~A301;
  assign \new_[65714]_  = ~A300 & \new_[65713]_ ;
  assign \new_[65715]_  = \new_[65714]_  & \new_[65709]_ ;
  assign \new_[65716]_  = \new_[65715]_  & \new_[65706]_ ;
  assign \new_[65719]_  = ~A169 & ~A170;
  assign \new_[65722]_  = A167 & ~A168;
  assign \new_[65723]_  = \new_[65722]_  & \new_[65719]_ ;
  assign \new_[65726]_  = ~A232 & ~A166;
  assign \new_[65729]_  = A234 & A233;
  assign \new_[65730]_  = \new_[65729]_  & \new_[65726]_ ;
  assign \new_[65731]_  = \new_[65730]_  & \new_[65723]_ ;
  assign \new_[65734]_  = A267 & ~A236;
  assign \new_[65737]_  = A269 & ~A268;
  assign \new_[65738]_  = \new_[65737]_  & \new_[65734]_ ;
  assign \new_[65741]_  = ~A299 & A298;
  assign \new_[65745]_  = A302 & ~A301;
  assign \new_[65746]_  = ~A300 & \new_[65745]_ ;
  assign \new_[65747]_  = \new_[65746]_  & \new_[65741]_ ;
  assign \new_[65748]_  = \new_[65747]_  & \new_[65738]_ ;
  assign \new_[65751]_  = ~A169 & ~A170;
  assign \new_[65754]_  = A167 & ~A168;
  assign \new_[65755]_  = \new_[65754]_  & \new_[65751]_ ;
  assign \new_[65758]_  = ~A232 & ~A166;
  assign \new_[65761]_  = A234 & A233;
  assign \new_[65762]_  = \new_[65761]_  & \new_[65758]_ ;
  assign \new_[65763]_  = \new_[65762]_  & \new_[65755]_ ;
  assign \new_[65766]_  = A267 & ~A236;
  assign \new_[65769]_  = A269 & ~A268;
  assign \new_[65770]_  = \new_[65769]_  & \new_[65766]_ ;
  assign \new_[65773]_  = A299 & ~A298;
  assign \new_[65777]_  = A302 & ~A301;
  assign \new_[65778]_  = ~A300 & \new_[65777]_ ;
  assign \new_[65779]_  = \new_[65778]_  & \new_[65773]_ ;
  assign \new_[65780]_  = \new_[65779]_  & \new_[65770]_ ;
  assign \new_[65783]_  = ~A169 & ~A170;
  assign \new_[65786]_  = A167 & ~A168;
  assign \new_[65787]_  = \new_[65786]_  & \new_[65783]_ ;
  assign \new_[65790]_  = ~A232 & ~A166;
  assign \new_[65793]_  = ~A234 & A233;
  assign \new_[65794]_  = \new_[65793]_  & \new_[65790]_ ;
  assign \new_[65795]_  = \new_[65794]_  & \new_[65787]_ ;
  assign \new_[65798]_  = A236 & ~A235;
  assign \new_[65801]_  = ~A268 & A267;
  assign \new_[65802]_  = \new_[65801]_  & \new_[65798]_ ;
  assign \new_[65805]_  = A298 & A269;
  assign \new_[65809]_  = A301 & A300;
  assign \new_[65810]_  = ~A299 & \new_[65809]_ ;
  assign \new_[65811]_  = \new_[65810]_  & \new_[65805]_ ;
  assign \new_[65812]_  = \new_[65811]_  & \new_[65802]_ ;
  assign \new_[65815]_  = ~A169 & ~A170;
  assign \new_[65818]_  = A167 & ~A168;
  assign \new_[65819]_  = \new_[65818]_  & \new_[65815]_ ;
  assign \new_[65822]_  = ~A232 & ~A166;
  assign \new_[65825]_  = ~A234 & A233;
  assign \new_[65826]_  = \new_[65825]_  & \new_[65822]_ ;
  assign \new_[65827]_  = \new_[65826]_  & \new_[65819]_ ;
  assign \new_[65830]_  = A236 & ~A235;
  assign \new_[65833]_  = ~A268 & A267;
  assign \new_[65834]_  = \new_[65833]_  & \new_[65830]_ ;
  assign \new_[65837]_  = A298 & A269;
  assign \new_[65841]_  = ~A302 & A300;
  assign \new_[65842]_  = ~A299 & \new_[65841]_ ;
  assign \new_[65843]_  = \new_[65842]_  & \new_[65837]_ ;
  assign \new_[65844]_  = \new_[65843]_  & \new_[65834]_ ;
  assign \new_[65847]_  = ~A169 & ~A170;
  assign \new_[65850]_  = A167 & ~A168;
  assign \new_[65851]_  = \new_[65850]_  & \new_[65847]_ ;
  assign \new_[65854]_  = ~A232 & ~A166;
  assign \new_[65857]_  = ~A234 & A233;
  assign \new_[65858]_  = \new_[65857]_  & \new_[65854]_ ;
  assign \new_[65859]_  = \new_[65858]_  & \new_[65851]_ ;
  assign \new_[65862]_  = A236 & ~A235;
  assign \new_[65865]_  = ~A268 & A267;
  assign \new_[65866]_  = \new_[65865]_  & \new_[65862]_ ;
  assign \new_[65869]_  = ~A298 & A269;
  assign \new_[65873]_  = A301 & A300;
  assign \new_[65874]_  = A299 & \new_[65873]_ ;
  assign \new_[65875]_  = \new_[65874]_  & \new_[65869]_ ;
  assign \new_[65876]_  = \new_[65875]_  & \new_[65866]_ ;
  assign \new_[65879]_  = ~A169 & ~A170;
  assign \new_[65882]_  = A167 & ~A168;
  assign \new_[65883]_  = \new_[65882]_  & \new_[65879]_ ;
  assign \new_[65886]_  = ~A232 & ~A166;
  assign \new_[65889]_  = ~A234 & A233;
  assign \new_[65890]_  = \new_[65889]_  & \new_[65886]_ ;
  assign \new_[65891]_  = \new_[65890]_  & \new_[65883]_ ;
  assign \new_[65894]_  = A236 & ~A235;
  assign \new_[65897]_  = ~A268 & A267;
  assign \new_[65898]_  = \new_[65897]_  & \new_[65894]_ ;
  assign \new_[65901]_  = ~A298 & A269;
  assign \new_[65905]_  = ~A302 & A300;
  assign \new_[65906]_  = A299 & \new_[65905]_ ;
  assign \new_[65907]_  = \new_[65906]_  & \new_[65901]_ ;
  assign \new_[65908]_  = \new_[65907]_  & \new_[65898]_ ;
  assign \new_[65911]_  = ~A169 & ~A170;
  assign \new_[65914]_  = A167 & ~A168;
  assign \new_[65915]_  = \new_[65914]_  & \new_[65911]_ ;
  assign \new_[65918]_  = ~A232 & ~A166;
  assign \new_[65921]_  = ~A234 & A233;
  assign \new_[65922]_  = \new_[65921]_  & \new_[65918]_ ;
  assign \new_[65923]_  = \new_[65922]_  & \new_[65915]_ ;
  assign \new_[65926]_  = A236 & ~A235;
  assign \new_[65929]_  = A268 & ~A267;
  assign \new_[65930]_  = \new_[65929]_  & \new_[65926]_ ;
  assign \new_[65933]_  = ~A299 & A298;
  assign \new_[65937]_  = A302 & ~A301;
  assign \new_[65938]_  = ~A300 & \new_[65937]_ ;
  assign \new_[65939]_  = \new_[65938]_  & \new_[65933]_ ;
  assign \new_[65940]_  = \new_[65939]_  & \new_[65930]_ ;
  assign \new_[65943]_  = ~A169 & ~A170;
  assign \new_[65946]_  = A167 & ~A168;
  assign \new_[65947]_  = \new_[65946]_  & \new_[65943]_ ;
  assign \new_[65950]_  = ~A232 & ~A166;
  assign \new_[65953]_  = ~A234 & A233;
  assign \new_[65954]_  = \new_[65953]_  & \new_[65950]_ ;
  assign \new_[65955]_  = \new_[65954]_  & \new_[65947]_ ;
  assign \new_[65958]_  = A236 & ~A235;
  assign \new_[65961]_  = A268 & ~A267;
  assign \new_[65962]_  = \new_[65961]_  & \new_[65958]_ ;
  assign \new_[65965]_  = A299 & ~A298;
  assign \new_[65969]_  = A302 & ~A301;
  assign \new_[65970]_  = ~A300 & \new_[65969]_ ;
  assign \new_[65971]_  = \new_[65970]_  & \new_[65965]_ ;
  assign \new_[65972]_  = \new_[65971]_  & \new_[65962]_ ;
  assign \new_[65975]_  = ~A169 & ~A170;
  assign \new_[65978]_  = A167 & ~A168;
  assign \new_[65979]_  = \new_[65978]_  & \new_[65975]_ ;
  assign \new_[65982]_  = ~A232 & ~A166;
  assign \new_[65985]_  = ~A234 & A233;
  assign \new_[65986]_  = \new_[65985]_  & \new_[65982]_ ;
  assign \new_[65987]_  = \new_[65986]_  & \new_[65979]_ ;
  assign \new_[65990]_  = A236 & ~A235;
  assign \new_[65993]_  = ~A269 & ~A267;
  assign \new_[65994]_  = \new_[65993]_  & \new_[65990]_ ;
  assign \new_[65997]_  = ~A299 & A298;
  assign \new_[66001]_  = A302 & ~A301;
  assign \new_[66002]_  = ~A300 & \new_[66001]_ ;
  assign \new_[66003]_  = \new_[66002]_  & \new_[65997]_ ;
  assign \new_[66004]_  = \new_[66003]_  & \new_[65994]_ ;
  assign \new_[66007]_  = ~A169 & ~A170;
  assign \new_[66010]_  = A167 & ~A168;
  assign \new_[66011]_  = \new_[66010]_  & \new_[66007]_ ;
  assign \new_[66014]_  = ~A232 & ~A166;
  assign \new_[66017]_  = ~A234 & A233;
  assign \new_[66018]_  = \new_[66017]_  & \new_[66014]_ ;
  assign \new_[66019]_  = \new_[66018]_  & \new_[66011]_ ;
  assign \new_[66022]_  = A236 & ~A235;
  assign \new_[66025]_  = ~A269 & ~A267;
  assign \new_[66026]_  = \new_[66025]_  & \new_[66022]_ ;
  assign \new_[66029]_  = A299 & ~A298;
  assign \new_[66033]_  = A302 & ~A301;
  assign \new_[66034]_  = ~A300 & \new_[66033]_ ;
  assign \new_[66035]_  = \new_[66034]_  & \new_[66029]_ ;
  assign \new_[66036]_  = \new_[66035]_  & \new_[66026]_ ;
  assign \new_[66039]_  = ~A169 & ~A170;
  assign \new_[66042]_  = A167 & ~A168;
  assign \new_[66043]_  = \new_[66042]_  & \new_[66039]_ ;
  assign \new_[66046]_  = ~A232 & ~A166;
  assign \new_[66049]_  = ~A234 & A233;
  assign \new_[66050]_  = \new_[66049]_  & \new_[66046]_ ;
  assign \new_[66051]_  = \new_[66050]_  & \new_[66043]_ ;
  assign \new_[66054]_  = A236 & ~A235;
  assign \new_[66057]_  = A266 & A265;
  assign \new_[66058]_  = \new_[66057]_  & \new_[66054]_ ;
  assign \new_[66061]_  = ~A299 & A298;
  assign \new_[66065]_  = A302 & ~A301;
  assign \new_[66066]_  = ~A300 & \new_[66065]_ ;
  assign \new_[66067]_  = \new_[66066]_  & \new_[66061]_ ;
  assign \new_[66068]_  = \new_[66067]_  & \new_[66058]_ ;
  assign \new_[66071]_  = ~A169 & ~A170;
  assign \new_[66074]_  = A167 & ~A168;
  assign \new_[66075]_  = \new_[66074]_  & \new_[66071]_ ;
  assign \new_[66078]_  = ~A232 & ~A166;
  assign \new_[66081]_  = ~A234 & A233;
  assign \new_[66082]_  = \new_[66081]_  & \new_[66078]_ ;
  assign \new_[66083]_  = \new_[66082]_  & \new_[66075]_ ;
  assign \new_[66086]_  = A236 & ~A235;
  assign \new_[66089]_  = A266 & A265;
  assign \new_[66090]_  = \new_[66089]_  & \new_[66086]_ ;
  assign \new_[66093]_  = A299 & ~A298;
  assign \new_[66097]_  = A302 & ~A301;
  assign \new_[66098]_  = ~A300 & \new_[66097]_ ;
  assign \new_[66099]_  = \new_[66098]_  & \new_[66093]_ ;
  assign \new_[66100]_  = \new_[66099]_  & \new_[66090]_ ;
  assign \new_[66103]_  = ~A169 & ~A170;
  assign \new_[66106]_  = A167 & ~A168;
  assign \new_[66107]_  = \new_[66106]_  & \new_[66103]_ ;
  assign \new_[66110]_  = ~A232 & ~A166;
  assign \new_[66113]_  = ~A234 & A233;
  assign \new_[66114]_  = \new_[66113]_  & \new_[66110]_ ;
  assign \new_[66115]_  = \new_[66114]_  & \new_[66107]_ ;
  assign \new_[66118]_  = A236 & ~A235;
  assign \new_[66121]_  = ~A266 & ~A265;
  assign \new_[66122]_  = \new_[66121]_  & \new_[66118]_ ;
  assign \new_[66125]_  = ~A299 & A298;
  assign \new_[66129]_  = A302 & ~A301;
  assign \new_[66130]_  = ~A300 & \new_[66129]_ ;
  assign \new_[66131]_  = \new_[66130]_  & \new_[66125]_ ;
  assign \new_[66132]_  = \new_[66131]_  & \new_[66122]_ ;
  assign \new_[66135]_  = ~A169 & ~A170;
  assign \new_[66138]_  = A167 & ~A168;
  assign \new_[66139]_  = \new_[66138]_  & \new_[66135]_ ;
  assign \new_[66142]_  = ~A232 & ~A166;
  assign \new_[66145]_  = ~A234 & A233;
  assign \new_[66146]_  = \new_[66145]_  & \new_[66142]_ ;
  assign \new_[66147]_  = \new_[66146]_  & \new_[66139]_ ;
  assign \new_[66150]_  = A236 & ~A235;
  assign \new_[66153]_  = ~A266 & ~A265;
  assign \new_[66154]_  = \new_[66153]_  & \new_[66150]_ ;
  assign \new_[66157]_  = A299 & ~A298;
  assign \new_[66161]_  = A302 & ~A301;
  assign \new_[66162]_  = ~A300 & \new_[66161]_ ;
  assign \new_[66163]_  = \new_[66162]_  & \new_[66157]_ ;
  assign \new_[66164]_  = \new_[66163]_  & \new_[66154]_ ;
  assign \new_[66167]_  = ~A169 & ~A170;
  assign \new_[66170]_  = A167 & ~A168;
  assign \new_[66171]_  = \new_[66170]_  & \new_[66167]_ ;
  assign \new_[66174]_  = A232 & ~A166;
  assign \new_[66177]_  = A234 & ~A233;
  assign \new_[66178]_  = \new_[66177]_  & \new_[66174]_ ;
  assign \new_[66179]_  = \new_[66178]_  & \new_[66171]_ ;
  assign \new_[66182]_  = A267 & A235;
  assign \new_[66185]_  = A269 & ~A268;
  assign \new_[66186]_  = \new_[66185]_  & \new_[66182]_ ;
  assign \new_[66189]_  = ~A299 & A298;
  assign \new_[66193]_  = A302 & ~A301;
  assign \new_[66194]_  = ~A300 & \new_[66193]_ ;
  assign \new_[66195]_  = \new_[66194]_  & \new_[66189]_ ;
  assign \new_[66196]_  = \new_[66195]_  & \new_[66186]_ ;
  assign \new_[66199]_  = ~A169 & ~A170;
  assign \new_[66202]_  = A167 & ~A168;
  assign \new_[66203]_  = \new_[66202]_  & \new_[66199]_ ;
  assign \new_[66206]_  = A232 & ~A166;
  assign \new_[66209]_  = A234 & ~A233;
  assign \new_[66210]_  = \new_[66209]_  & \new_[66206]_ ;
  assign \new_[66211]_  = \new_[66210]_  & \new_[66203]_ ;
  assign \new_[66214]_  = A267 & A235;
  assign \new_[66217]_  = A269 & ~A268;
  assign \new_[66218]_  = \new_[66217]_  & \new_[66214]_ ;
  assign \new_[66221]_  = A299 & ~A298;
  assign \new_[66225]_  = A302 & ~A301;
  assign \new_[66226]_  = ~A300 & \new_[66225]_ ;
  assign \new_[66227]_  = \new_[66226]_  & \new_[66221]_ ;
  assign \new_[66228]_  = \new_[66227]_  & \new_[66218]_ ;
  assign \new_[66231]_  = ~A169 & ~A170;
  assign \new_[66234]_  = A167 & ~A168;
  assign \new_[66235]_  = \new_[66234]_  & \new_[66231]_ ;
  assign \new_[66238]_  = A232 & ~A166;
  assign \new_[66241]_  = A234 & ~A233;
  assign \new_[66242]_  = \new_[66241]_  & \new_[66238]_ ;
  assign \new_[66243]_  = \new_[66242]_  & \new_[66235]_ ;
  assign \new_[66246]_  = A267 & ~A236;
  assign \new_[66249]_  = A269 & ~A268;
  assign \new_[66250]_  = \new_[66249]_  & \new_[66246]_ ;
  assign \new_[66253]_  = ~A299 & A298;
  assign \new_[66257]_  = A302 & ~A301;
  assign \new_[66258]_  = ~A300 & \new_[66257]_ ;
  assign \new_[66259]_  = \new_[66258]_  & \new_[66253]_ ;
  assign \new_[66260]_  = \new_[66259]_  & \new_[66250]_ ;
  assign \new_[66263]_  = ~A169 & ~A170;
  assign \new_[66266]_  = A167 & ~A168;
  assign \new_[66267]_  = \new_[66266]_  & \new_[66263]_ ;
  assign \new_[66270]_  = A232 & ~A166;
  assign \new_[66273]_  = A234 & ~A233;
  assign \new_[66274]_  = \new_[66273]_  & \new_[66270]_ ;
  assign \new_[66275]_  = \new_[66274]_  & \new_[66267]_ ;
  assign \new_[66278]_  = A267 & ~A236;
  assign \new_[66281]_  = A269 & ~A268;
  assign \new_[66282]_  = \new_[66281]_  & \new_[66278]_ ;
  assign \new_[66285]_  = A299 & ~A298;
  assign \new_[66289]_  = A302 & ~A301;
  assign \new_[66290]_  = ~A300 & \new_[66289]_ ;
  assign \new_[66291]_  = \new_[66290]_  & \new_[66285]_ ;
  assign \new_[66292]_  = \new_[66291]_  & \new_[66282]_ ;
  assign \new_[66295]_  = ~A169 & ~A170;
  assign \new_[66298]_  = A167 & ~A168;
  assign \new_[66299]_  = \new_[66298]_  & \new_[66295]_ ;
  assign \new_[66302]_  = A232 & ~A166;
  assign \new_[66305]_  = ~A234 & ~A233;
  assign \new_[66306]_  = \new_[66305]_  & \new_[66302]_ ;
  assign \new_[66307]_  = \new_[66306]_  & \new_[66299]_ ;
  assign \new_[66310]_  = A236 & ~A235;
  assign \new_[66313]_  = ~A268 & A267;
  assign \new_[66314]_  = \new_[66313]_  & \new_[66310]_ ;
  assign \new_[66317]_  = A298 & A269;
  assign \new_[66321]_  = A301 & A300;
  assign \new_[66322]_  = ~A299 & \new_[66321]_ ;
  assign \new_[66323]_  = \new_[66322]_  & \new_[66317]_ ;
  assign \new_[66324]_  = \new_[66323]_  & \new_[66314]_ ;
  assign \new_[66327]_  = ~A169 & ~A170;
  assign \new_[66330]_  = A167 & ~A168;
  assign \new_[66331]_  = \new_[66330]_  & \new_[66327]_ ;
  assign \new_[66334]_  = A232 & ~A166;
  assign \new_[66337]_  = ~A234 & ~A233;
  assign \new_[66338]_  = \new_[66337]_  & \new_[66334]_ ;
  assign \new_[66339]_  = \new_[66338]_  & \new_[66331]_ ;
  assign \new_[66342]_  = A236 & ~A235;
  assign \new_[66345]_  = ~A268 & A267;
  assign \new_[66346]_  = \new_[66345]_  & \new_[66342]_ ;
  assign \new_[66349]_  = A298 & A269;
  assign \new_[66353]_  = ~A302 & A300;
  assign \new_[66354]_  = ~A299 & \new_[66353]_ ;
  assign \new_[66355]_  = \new_[66354]_  & \new_[66349]_ ;
  assign \new_[66356]_  = \new_[66355]_  & \new_[66346]_ ;
  assign \new_[66359]_  = ~A169 & ~A170;
  assign \new_[66362]_  = A167 & ~A168;
  assign \new_[66363]_  = \new_[66362]_  & \new_[66359]_ ;
  assign \new_[66366]_  = A232 & ~A166;
  assign \new_[66369]_  = ~A234 & ~A233;
  assign \new_[66370]_  = \new_[66369]_  & \new_[66366]_ ;
  assign \new_[66371]_  = \new_[66370]_  & \new_[66363]_ ;
  assign \new_[66374]_  = A236 & ~A235;
  assign \new_[66377]_  = ~A268 & A267;
  assign \new_[66378]_  = \new_[66377]_  & \new_[66374]_ ;
  assign \new_[66381]_  = ~A298 & A269;
  assign \new_[66385]_  = A301 & A300;
  assign \new_[66386]_  = A299 & \new_[66385]_ ;
  assign \new_[66387]_  = \new_[66386]_  & \new_[66381]_ ;
  assign \new_[66388]_  = \new_[66387]_  & \new_[66378]_ ;
  assign \new_[66391]_  = ~A169 & ~A170;
  assign \new_[66394]_  = A167 & ~A168;
  assign \new_[66395]_  = \new_[66394]_  & \new_[66391]_ ;
  assign \new_[66398]_  = A232 & ~A166;
  assign \new_[66401]_  = ~A234 & ~A233;
  assign \new_[66402]_  = \new_[66401]_  & \new_[66398]_ ;
  assign \new_[66403]_  = \new_[66402]_  & \new_[66395]_ ;
  assign \new_[66406]_  = A236 & ~A235;
  assign \new_[66409]_  = ~A268 & A267;
  assign \new_[66410]_  = \new_[66409]_  & \new_[66406]_ ;
  assign \new_[66413]_  = ~A298 & A269;
  assign \new_[66417]_  = ~A302 & A300;
  assign \new_[66418]_  = A299 & \new_[66417]_ ;
  assign \new_[66419]_  = \new_[66418]_  & \new_[66413]_ ;
  assign \new_[66420]_  = \new_[66419]_  & \new_[66410]_ ;
  assign \new_[66423]_  = ~A169 & ~A170;
  assign \new_[66426]_  = A167 & ~A168;
  assign \new_[66427]_  = \new_[66426]_  & \new_[66423]_ ;
  assign \new_[66430]_  = A232 & ~A166;
  assign \new_[66433]_  = ~A234 & ~A233;
  assign \new_[66434]_  = \new_[66433]_  & \new_[66430]_ ;
  assign \new_[66435]_  = \new_[66434]_  & \new_[66427]_ ;
  assign \new_[66438]_  = A236 & ~A235;
  assign \new_[66441]_  = A268 & ~A267;
  assign \new_[66442]_  = \new_[66441]_  & \new_[66438]_ ;
  assign \new_[66445]_  = ~A299 & A298;
  assign \new_[66449]_  = A302 & ~A301;
  assign \new_[66450]_  = ~A300 & \new_[66449]_ ;
  assign \new_[66451]_  = \new_[66450]_  & \new_[66445]_ ;
  assign \new_[66452]_  = \new_[66451]_  & \new_[66442]_ ;
  assign \new_[66455]_  = ~A169 & ~A170;
  assign \new_[66458]_  = A167 & ~A168;
  assign \new_[66459]_  = \new_[66458]_  & \new_[66455]_ ;
  assign \new_[66462]_  = A232 & ~A166;
  assign \new_[66465]_  = ~A234 & ~A233;
  assign \new_[66466]_  = \new_[66465]_  & \new_[66462]_ ;
  assign \new_[66467]_  = \new_[66466]_  & \new_[66459]_ ;
  assign \new_[66470]_  = A236 & ~A235;
  assign \new_[66473]_  = A268 & ~A267;
  assign \new_[66474]_  = \new_[66473]_  & \new_[66470]_ ;
  assign \new_[66477]_  = A299 & ~A298;
  assign \new_[66481]_  = A302 & ~A301;
  assign \new_[66482]_  = ~A300 & \new_[66481]_ ;
  assign \new_[66483]_  = \new_[66482]_  & \new_[66477]_ ;
  assign \new_[66484]_  = \new_[66483]_  & \new_[66474]_ ;
  assign \new_[66487]_  = ~A169 & ~A170;
  assign \new_[66490]_  = A167 & ~A168;
  assign \new_[66491]_  = \new_[66490]_  & \new_[66487]_ ;
  assign \new_[66494]_  = A232 & ~A166;
  assign \new_[66497]_  = ~A234 & ~A233;
  assign \new_[66498]_  = \new_[66497]_  & \new_[66494]_ ;
  assign \new_[66499]_  = \new_[66498]_  & \new_[66491]_ ;
  assign \new_[66502]_  = A236 & ~A235;
  assign \new_[66505]_  = ~A269 & ~A267;
  assign \new_[66506]_  = \new_[66505]_  & \new_[66502]_ ;
  assign \new_[66509]_  = ~A299 & A298;
  assign \new_[66513]_  = A302 & ~A301;
  assign \new_[66514]_  = ~A300 & \new_[66513]_ ;
  assign \new_[66515]_  = \new_[66514]_  & \new_[66509]_ ;
  assign \new_[66516]_  = \new_[66515]_  & \new_[66506]_ ;
  assign \new_[66519]_  = ~A169 & ~A170;
  assign \new_[66522]_  = A167 & ~A168;
  assign \new_[66523]_  = \new_[66522]_  & \new_[66519]_ ;
  assign \new_[66526]_  = A232 & ~A166;
  assign \new_[66529]_  = ~A234 & ~A233;
  assign \new_[66530]_  = \new_[66529]_  & \new_[66526]_ ;
  assign \new_[66531]_  = \new_[66530]_  & \new_[66523]_ ;
  assign \new_[66534]_  = A236 & ~A235;
  assign \new_[66537]_  = ~A269 & ~A267;
  assign \new_[66538]_  = \new_[66537]_  & \new_[66534]_ ;
  assign \new_[66541]_  = A299 & ~A298;
  assign \new_[66545]_  = A302 & ~A301;
  assign \new_[66546]_  = ~A300 & \new_[66545]_ ;
  assign \new_[66547]_  = \new_[66546]_  & \new_[66541]_ ;
  assign \new_[66548]_  = \new_[66547]_  & \new_[66538]_ ;
  assign \new_[66551]_  = ~A169 & ~A170;
  assign \new_[66554]_  = A167 & ~A168;
  assign \new_[66555]_  = \new_[66554]_  & \new_[66551]_ ;
  assign \new_[66558]_  = A232 & ~A166;
  assign \new_[66561]_  = ~A234 & ~A233;
  assign \new_[66562]_  = \new_[66561]_  & \new_[66558]_ ;
  assign \new_[66563]_  = \new_[66562]_  & \new_[66555]_ ;
  assign \new_[66566]_  = A236 & ~A235;
  assign \new_[66569]_  = A266 & A265;
  assign \new_[66570]_  = \new_[66569]_  & \new_[66566]_ ;
  assign \new_[66573]_  = ~A299 & A298;
  assign \new_[66577]_  = A302 & ~A301;
  assign \new_[66578]_  = ~A300 & \new_[66577]_ ;
  assign \new_[66579]_  = \new_[66578]_  & \new_[66573]_ ;
  assign \new_[66580]_  = \new_[66579]_  & \new_[66570]_ ;
  assign \new_[66583]_  = ~A169 & ~A170;
  assign \new_[66586]_  = A167 & ~A168;
  assign \new_[66587]_  = \new_[66586]_  & \new_[66583]_ ;
  assign \new_[66590]_  = A232 & ~A166;
  assign \new_[66593]_  = ~A234 & ~A233;
  assign \new_[66594]_  = \new_[66593]_  & \new_[66590]_ ;
  assign \new_[66595]_  = \new_[66594]_  & \new_[66587]_ ;
  assign \new_[66598]_  = A236 & ~A235;
  assign \new_[66601]_  = A266 & A265;
  assign \new_[66602]_  = \new_[66601]_  & \new_[66598]_ ;
  assign \new_[66605]_  = A299 & ~A298;
  assign \new_[66609]_  = A302 & ~A301;
  assign \new_[66610]_  = ~A300 & \new_[66609]_ ;
  assign \new_[66611]_  = \new_[66610]_  & \new_[66605]_ ;
  assign \new_[66612]_  = \new_[66611]_  & \new_[66602]_ ;
  assign \new_[66615]_  = ~A169 & ~A170;
  assign \new_[66618]_  = A167 & ~A168;
  assign \new_[66619]_  = \new_[66618]_  & \new_[66615]_ ;
  assign \new_[66622]_  = A232 & ~A166;
  assign \new_[66625]_  = ~A234 & ~A233;
  assign \new_[66626]_  = \new_[66625]_  & \new_[66622]_ ;
  assign \new_[66627]_  = \new_[66626]_  & \new_[66619]_ ;
  assign \new_[66630]_  = A236 & ~A235;
  assign \new_[66633]_  = ~A266 & ~A265;
  assign \new_[66634]_  = \new_[66633]_  & \new_[66630]_ ;
  assign \new_[66637]_  = ~A299 & A298;
  assign \new_[66641]_  = A302 & ~A301;
  assign \new_[66642]_  = ~A300 & \new_[66641]_ ;
  assign \new_[66643]_  = \new_[66642]_  & \new_[66637]_ ;
  assign \new_[66644]_  = \new_[66643]_  & \new_[66634]_ ;
  assign \new_[66647]_  = ~A169 & ~A170;
  assign \new_[66650]_  = A167 & ~A168;
  assign \new_[66651]_  = \new_[66650]_  & \new_[66647]_ ;
  assign \new_[66654]_  = A232 & ~A166;
  assign \new_[66657]_  = ~A234 & ~A233;
  assign \new_[66658]_  = \new_[66657]_  & \new_[66654]_ ;
  assign \new_[66659]_  = \new_[66658]_  & \new_[66651]_ ;
  assign \new_[66662]_  = A236 & ~A235;
  assign \new_[66665]_  = ~A266 & ~A265;
  assign \new_[66666]_  = \new_[66665]_  & \new_[66662]_ ;
  assign \new_[66669]_  = A299 & ~A298;
  assign \new_[66673]_  = A302 & ~A301;
  assign \new_[66674]_  = ~A300 & \new_[66673]_ ;
  assign \new_[66675]_  = \new_[66674]_  & \new_[66669]_ ;
  assign \new_[66676]_  = \new_[66675]_  & \new_[66666]_ ;
  assign \new_[66679]_  = ~A169 & ~A170;
  assign \new_[66682]_  = ~A167 & ~A168;
  assign \new_[66683]_  = \new_[66682]_  & \new_[66679]_ ;
  assign \new_[66686]_  = ~A232 & A166;
  assign \new_[66689]_  = A234 & A233;
  assign \new_[66690]_  = \new_[66689]_  & \new_[66686]_ ;
  assign \new_[66691]_  = \new_[66690]_  & \new_[66683]_ ;
  assign \new_[66694]_  = A267 & A235;
  assign \new_[66697]_  = A269 & ~A268;
  assign \new_[66698]_  = \new_[66697]_  & \new_[66694]_ ;
  assign \new_[66701]_  = ~A299 & A298;
  assign \new_[66705]_  = A302 & ~A301;
  assign \new_[66706]_  = ~A300 & \new_[66705]_ ;
  assign \new_[66707]_  = \new_[66706]_  & \new_[66701]_ ;
  assign \new_[66708]_  = \new_[66707]_  & \new_[66698]_ ;
  assign \new_[66711]_  = ~A169 & ~A170;
  assign \new_[66714]_  = ~A167 & ~A168;
  assign \new_[66715]_  = \new_[66714]_  & \new_[66711]_ ;
  assign \new_[66718]_  = ~A232 & A166;
  assign \new_[66721]_  = A234 & A233;
  assign \new_[66722]_  = \new_[66721]_  & \new_[66718]_ ;
  assign \new_[66723]_  = \new_[66722]_  & \new_[66715]_ ;
  assign \new_[66726]_  = A267 & A235;
  assign \new_[66729]_  = A269 & ~A268;
  assign \new_[66730]_  = \new_[66729]_  & \new_[66726]_ ;
  assign \new_[66733]_  = A299 & ~A298;
  assign \new_[66737]_  = A302 & ~A301;
  assign \new_[66738]_  = ~A300 & \new_[66737]_ ;
  assign \new_[66739]_  = \new_[66738]_  & \new_[66733]_ ;
  assign \new_[66740]_  = \new_[66739]_  & \new_[66730]_ ;
  assign \new_[66743]_  = ~A169 & ~A170;
  assign \new_[66746]_  = ~A167 & ~A168;
  assign \new_[66747]_  = \new_[66746]_  & \new_[66743]_ ;
  assign \new_[66750]_  = ~A232 & A166;
  assign \new_[66753]_  = A234 & A233;
  assign \new_[66754]_  = \new_[66753]_  & \new_[66750]_ ;
  assign \new_[66755]_  = \new_[66754]_  & \new_[66747]_ ;
  assign \new_[66758]_  = A267 & ~A236;
  assign \new_[66761]_  = A269 & ~A268;
  assign \new_[66762]_  = \new_[66761]_  & \new_[66758]_ ;
  assign \new_[66765]_  = ~A299 & A298;
  assign \new_[66769]_  = A302 & ~A301;
  assign \new_[66770]_  = ~A300 & \new_[66769]_ ;
  assign \new_[66771]_  = \new_[66770]_  & \new_[66765]_ ;
  assign \new_[66772]_  = \new_[66771]_  & \new_[66762]_ ;
  assign \new_[66775]_  = ~A169 & ~A170;
  assign \new_[66778]_  = ~A167 & ~A168;
  assign \new_[66779]_  = \new_[66778]_  & \new_[66775]_ ;
  assign \new_[66782]_  = ~A232 & A166;
  assign \new_[66785]_  = A234 & A233;
  assign \new_[66786]_  = \new_[66785]_  & \new_[66782]_ ;
  assign \new_[66787]_  = \new_[66786]_  & \new_[66779]_ ;
  assign \new_[66790]_  = A267 & ~A236;
  assign \new_[66793]_  = A269 & ~A268;
  assign \new_[66794]_  = \new_[66793]_  & \new_[66790]_ ;
  assign \new_[66797]_  = A299 & ~A298;
  assign \new_[66801]_  = A302 & ~A301;
  assign \new_[66802]_  = ~A300 & \new_[66801]_ ;
  assign \new_[66803]_  = \new_[66802]_  & \new_[66797]_ ;
  assign \new_[66804]_  = \new_[66803]_  & \new_[66794]_ ;
  assign \new_[66807]_  = ~A169 & ~A170;
  assign \new_[66810]_  = ~A167 & ~A168;
  assign \new_[66811]_  = \new_[66810]_  & \new_[66807]_ ;
  assign \new_[66814]_  = ~A232 & A166;
  assign \new_[66817]_  = ~A234 & A233;
  assign \new_[66818]_  = \new_[66817]_  & \new_[66814]_ ;
  assign \new_[66819]_  = \new_[66818]_  & \new_[66811]_ ;
  assign \new_[66822]_  = A236 & ~A235;
  assign \new_[66825]_  = ~A268 & A267;
  assign \new_[66826]_  = \new_[66825]_  & \new_[66822]_ ;
  assign \new_[66829]_  = A298 & A269;
  assign \new_[66833]_  = A301 & A300;
  assign \new_[66834]_  = ~A299 & \new_[66833]_ ;
  assign \new_[66835]_  = \new_[66834]_  & \new_[66829]_ ;
  assign \new_[66836]_  = \new_[66835]_  & \new_[66826]_ ;
  assign \new_[66839]_  = ~A169 & ~A170;
  assign \new_[66842]_  = ~A167 & ~A168;
  assign \new_[66843]_  = \new_[66842]_  & \new_[66839]_ ;
  assign \new_[66846]_  = ~A232 & A166;
  assign \new_[66849]_  = ~A234 & A233;
  assign \new_[66850]_  = \new_[66849]_  & \new_[66846]_ ;
  assign \new_[66851]_  = \new_[66850]_  & \new_[66843]_ ;
  assign \new_[66854]_  = A236 & ~A235;
  assign \new_[66857]_  = ~A268 & A267;
  assign \new_[66858]_  = \new_[66857]_  & \new_[66854]_ ;
  assign \new_[66861]_  = A298 & A269;
  assign \new_[66865]_  = ~A302 & A300;
  assign \new_[66866]_  = ~A299 & \new_[66865]_ ;
  assign \new_[66867]_  = \new_[66866]_  & \new_[66861]_ ;
  assign \new_[66868]_  = \new_[66867]_  & \new_[66858]_ ;
  assign \new_[66871]_  = ~A169 & ~A170;
  assign \new_[66874]_  = ~A167 & ~A168;
  assign \new_[66875]_  = \new_[66874]_  & \new_[66871]_ ;
  assign \new_[66878]_  = ~A232 & A166;
  assign \new_[66881]_  = ~A234 & A233;
  assign \new_[66882]_  = \new_[66881]_  & \new_[66878]_ ;
  assign \new_[66883]_  = \new_[66882]_  & \new_[66875]_ ;
  assign \new_[66886]_  = A236 & ~A235;
  assign \new_[66889]_  = ~A268 & A267;
  assign \new_[66890]_  = \new_[66889]_  & \new_[66886]_ ;
  assign \new_[66893]_  = ~A298 & A269;
  assign \new_[66897]_  = A301 & A300;
  assign \new_[66898]_  = A299 & \new_[66897]_ ;
  assign \new_[66899]_  = \new_[66898]_  & \new_[66893]_ ;
  assign \new_[66900]_  = \new_[66899]_  & \new_[66890]_ ;
  assign \new_[66903]_  = ~A169 & ~A170;
  assign \new_[66906]_  = ~A167 & ~A168;
  assign \new_[66907]_  = \new_[66906]_  & \new_[66903]_ ;
  assign \new_[66910]_  = ~A232 & A166;
  assign \new_[66913]_  = ~A234 & A233;
  assign \new_[66914]_  = \new_[66913]_  & \new_[66910]_ ;
  assign \new_[66915]_  = \new_[66914]_  & \new_[66907]_ ;
  assign \new_[66918]_  = A236 & ~A235;
  assign \new_[66921]_  = ~A268 & A267;
  assign \new_[66922]_  = \new_[66921]_  & \new_[66918]_ ;
  assign \new_[66925]_  = ~A298 & A269;
  assign \new_[66929]_  = ~A302 & A300;
  assign \new_[66930]_  = A299 & \new_[66929]_ ;
  assign \new_[66931]_  = \new_[66930]_  & \new_[66925]_ ;
  assign \new_[66932]_  = \new_[66931]_  & \new_[66922]_ ;
  assign \new_[66935]_  = ~A169 & ~A170;
  assign \new_[66938]_  = ~A167 & ~A168;
  assign \new_[66939]_  = \new_[66938]_  & \new_[66935]_ ;
  assign \new_[66942]_  = ~A232 & A166;
  assign \new_[66945]_  = ~A234 & A233;
  assign \new_[66946]_  = \new_[66945]_  & \new_[66942]_ ;
  assign \new_[66947]_  = \new_[66946]_  & \new_[66939]_ ;
  assign \new_[66950]_  = A236 & ~A235;
  assign \new_[66953]_  = A268 & ~A267;
  assign \new_[66954]_  = \new_[66953]_  & \new_[66950]_ ;
  assign \new_[66957]_  = ~A299 & A298;
  assign \new_[66961]_  = A302 & ~A301;
  assign \new_[66962]_  = ~A300 & \new_[66961]_ ;
  assign \new_[66963]_  = \new_[66962]_  & \new_[66957]_ ;
  assign \new_[66964]_  = \new_[66963]_  & \new_[66954]_ ;
  assign \new_[66967]_  = ~A169 & ~A170;
  assign \new_[66970]_  = ~A167 & ~A168;
  assign \new_[66971]_  = \new_[66970]_  & \new_[66967]_ ;
  assign \new_[66974]_  = ~A232 & A166;
  assign \new_[66977]_  = ~A234 & A233;
  assign \new_[66978]_  = \new_[66977]_  & \new_[66974]_ ;
  assign \new_[66979]_  = \new_[66978]_  & \new_[66971]_ ;
  assign \new_[66982]_  = A236 & ~A235;
  assign \new_[66985]_  = A268 & ~A267;
  assign \new_[66986]_  = \new_[66985]_  & \new_[66982]_ ;
  assign \new_[66989]_  = A299 & ~A298;
  assign \new_[66993]_  = A302 & ~A301;
  assign \new_[66994]_  = ~A300 & \new_[66993]_ ;
  assign \new_[66995]_  = \new_[66994]_  & \new_[66989]_ ;
  assign \new_[66996]_  = \new_[66995]_  & \new_[66986]_ ;
  assign \new_[66999]_  = ~A169 & ~A170;
  assign \new_[67002]_  = ~A167 & ~A168;
  assign \new_[67003]_  = \new_[67002]_  & \new_[66999]_ ;
  assign \new_[67006]_  = ~A232 & A166;
  assign \new_[67009]_  = ~A234 & A233;
  assign \new_[67010]_  = \new_[67009]_  & \new_[67006]_ ;
  assign \new_[67011]_  = \new_[67010]_  & \new_[67003]_ ;
  assign \new_[67014]_  = A236 & ~A235;
  assign \new_[67017]_  = ~A269 & ~A267;
  assign \new_[67018]_  = \new_[67017]_  & \new_[67014]_ ;
  assign \new_[67021]_  = ~A299 & A298;
  assign \new_[67025]_  = A302 & ~A301;
  assign \new_[67026]_  = ~A300 & \new_[67025]_ ;
  assign \new_[67027]_  = \new_[67026]_  & \new_[67021]_ ;
  assign \new_[67028]_  = \new_[67027]_  & \new_[67018]_ ;
  assign \new_[67031]_  = ~A169 & ~A170;
  assign \new_[67034]_  = ~A167 & ~A168;
  assign \new_[67035]_  = \new_[67034]_  & \new_[67031]_ ;
  assign \new_[67038]_  = ~A232 & A166;
  assign \new_[67041]_  = ~A234 & A233;
  assign \new_[67042]_  = \new_[67041]_  & \new_[67038]_ ;
  assign \new_[67043]_  = \new_[67042]_  & \new_[67035]_ ;
  assign \new_[67046]_  = A236 & ~A235;
  assign \new_[67049]_  = ~A269 & ~A267;
  assign \new_[67050]_  = \new_[67049]_  & \new_[67046]_ ;
  assign \new_[67053]_  = A299 & ~A298;
  assign \new_[67057]_  = A302 & ~A301;
  assign \new_[67058]_  = ~A300 & \new_[67057]_ ;
  assign \new_[67059]_  = \new_[67058]_  & \new_[67053]_ ;
  assign \new_[67060]_  = \new_[67059]_  & \new_[67050]_ ;
  assign \new_[67063]_  = ~A169 & ~A170;
  assign \new_[67066]_  = ~A167 & ~A168;
  assign \new_[67067]_  = \new_[67066]_  & \new_[67063]_ ;
  assign \new_[67070]_  = ~A232 & A166;
  assign \new_[67073]_  = ~A234 & A233;
  assign \new_[67074]_  = \new_[67073]_  & \new_[67070]_ ;
  assign \new_[67075]_  = \new_[67074]_  & \new_[67067]_ ;
  assign \new_[67078]_  = A236 & ~A235;
  assign \new_[67081]_  = A266 & A265;
  assign \new_[67082]_  = \new_[67081]_  & \new_[67078]_ ;
  assign \new_[67085]_  = ~A299 & A298;
  assign \new_[67089]_  = A302 & ~A301;
  assign \new_[67090]_  = ~A300 & \new_[67089]_ ;
  assign \new_[67091]_  = \new_[67090]_  & \new_[67085]_ ;
  assign \new_[67092]_  = \new_[67091]_  & \new_[67082]_ ;
  assign \new_[67095]_  = ~A169 & ~A170;
  assign \new_[67098]_  = ~A167 & ~A168;
  assign \new_[67099]_  = \new_[67098]_  & \new_[67095]_ ;
  assign \new_[67102]_  = ~A232 & A166;
  assign \new_[67105]_  = ~A234 & A233;
  assign \new_[67106]_  = \new_[67105]_  & \new_[67102]_ ;
  assign \new_[67107]_  = \new_[67106]_  & \new_[67099]_ ;
  assign \new_[67110]_  = A236 & ~A235;
  assign \new_[67113]_  = A266 & A265;
  assign \new_[67114]_  = \new_[67113]_  & \new_[67110]_ ;
  assign \new_[67117]_  = A299 & ~A298;
  assign \new_[67121]_  = A302 & ~A301;
  assign \new_[67122]_  = ~A300 & \new_[67121]_ ;
  assign \new_[67123]_  = \new_[67122]_  & \new_[67117]_ ;
  assign \new_[67124]_  = \new_[67123]_  & \new_[67114]_ ;
  assign \new_[67127]_  = ~A169 & ~A170;
  assign \new_[67130]_  = ~A167 & ~A168;
  assign \new_[67131]_  = \new_[67130]_  & \new_[67127]_ ;
  assign \new_[67134]_  = ~A232 & A166;
  assign \new_[67137]_  = ~A234 & A233;
  assign \new_[67138]_  = \new_[67137]_  & \new_[67134]_ ;
  assign \new_[67139]_  = \new_[67138]_  & \new_[67131]_ ;
  assign \new_[67142]_  = A236 & ~A235;
  assign \new_[67145]_  = ~A266 & ~A265;
  assign \new_[67146]_  = \new_[67145]_  & \new_[67142]_ ;
  assign \new_[67149]_  = ~A299 & A298;
  assign \new_[67153]_  = A302 & ~A301;
  assign \new_[67154]_  = ~A300 & \new_[67153]_ ;
  assign \new_[67155]_  = \new_[67154]_  & \new_[67149]_ ;
  assign \new_[67156]_  = \new_[67155]_  & \new_[67146]_ ;
  assign \new_[67159]_  = ~A169 & ~A170;
  assign \new_[67162]_  = ~A167 & ~A168;
  assign \new_[67163]_  = \new_[67162]_  & \new_[67159]_ ;
  assign \new_[67166]_  = ~A232 & A166;
  assign \new_[67169]_  = ~A234 & A233;
  assign \new_[67170]_  = \new_[67169]_  & \new_[67166]_ ;
  assign \new_[67171]_  = \new_[67170]_  & \new_[67163]_ ;
  assign \new_[67174]_  = A236 & ~A235;
  assign \new_[67177]_  = ~A266 & ~A265;
  assign \new_[67178]_  = \new_[67177]_  & \new_[67174]_ ;
  assign \new_[67181]_  = A299 & ~A298;
  assign \new_[67185]_  = A302 & ~A301;
  assign \new_[67186]_  = ~A300 & \new_[67185]_ ;
  assign \new_[67187]_  = \new_[67186]_  & \new_[67181]_ ;
  assign \new_[67188]_  = \new_[67187]_  & \new_[67178]_ ;
  assign \new_[67191]_  = ~A169 & ~A170;
  assign \new_[67194]_  = ~A167 & ~A168;
  assign \new_[67195]_  = \new_[67194]_  & \new_[67191]_ ;
  assign \new_[67198]_  = A232 & A166;
  assign \new_[67201]_  = A234 & ~A233;
  assign \new_[67202]_  = \new_[67201]_  & \new_[67198]_ ;
  assign \new_[67203]_  = \new_[67202]_  & \new_[67195]_ ;
  assign \new_[67206]_  = A267 & A235;
  assign \new_[67209]_  = A269 & ~A268;
  assign \new_[67210]_  = \new_[67209]_  & \new_[67206]_ ;
  assign \new_[67213]_  = ~A299 & A298;
  assign \new_[67217]_  = A302 & ~A301;
  assign \new_[67218]_  = ~A300 & \new_[67217]_ ;
  assign \new_[67219]_  = \new_[67218]_  & \new_[67213]_ ;
  assign \new_[67220]_  = \new_[67219]_  & \new_[67210]_ ;
  assign \new_[67223]_  = ~A169 & ~A170;
  assign \new_[67226]_  = ~A167 & ~A168;
  assign \new_[67227]_  = \new_[67226]_  & \new_[67223]_ ;
  assign \new_[67230]_  = A232 & A166;
  assign \new_[67233]_  = A234 & ~A233;
  assign \new_[67234]_  = \new_[67233]_  & \new_[67230]_ ;
  assign \new_[67235]_  = \new_[67234]_  & \new_[67227]_ ;
  assign \new_[67238]_  = A267 & A235;
  assign \new_[67241]_  = A269 & ~A268;
  assign \new_[67242]_  = \new_[67241]_  & \new_[67238]_ ;
  assign \new_[67245]_  = A299 & ~A298;
  assign \new_[67249]_  = A302 & ~A301;
  assign \new_[67250]_  = ~A300 & \new_[67249]_ ;
  assign \new_[67251]_  = \new_[67250]_  & \new_[67245]_ ;
  assign \new_[67252]_  = \new_[67251]_  & \new_[67242]_ ;
  assign \new_[67255]_  = ~A169 & ~A170;
  assign \new_[67258]_  = ~A167 & ~A168;
  assign \new_[67259]_  = \new_[67258]_  & \new_[67255]_ ;
  assign \new_[67262]_  = A232 & A166;
  assign \new_[67265]_  = A234 & ~A233;
  assign \new_[67266]_  = \new_[67265]_  & \new_[67262]_ ;
  assign \new_[67267]_  = \new_[67266]_  & \new_[67259]_ ;
  assign \new_[67270]_  = A267 & ~A236;
  assign \new_[67273]_  = A269 & ~A268;
  assign \new_[67274]_  = \new_[67273]_  & \new_[67270]_ ;
  assign \new_[67277]_  = ~A299 & A298;
  assign \new_[67281]_  = A302 & ~A301;
  assign \new_[67282]_  = ~A300 & \new_[67281]_ ;
  assign \new_[67283]_  = \new_[67282]_  & \new_[67277]_ ;
  assign \new_[67284]_  = \new_[67283]_  & \new_[67274]_ ;
  assign \new_[67287]_  = ~A169 & ~A170;
  assign \new_[67290]_  = ~A167 & ~A168;
  assign \new_[67291]_  = \new_[67290]_  & \new_[67287]_ ;
  assign \new_[67294]_  = A232 & A166;
  assign \new_[67297]_  = A234 & ~A233;
  assign \new_[67298]_  = \new_[67297]_  & \new_[67294]_ ;
  assign \new_[67299]_  = \new_[67298]_  & \new_[67291]_ ;
  assign \new_[67302]_  = A267 & ~A236;
  assign \new_[67305]_  = A269 & ~A268;
  assign \new_[67306]_  = \new_[67305]_  & \new_[67302]_ ;
  assign \new_[67309]_  = A299 & ~A298;
  assign \new_[67313]_  = A302 & ~A301;
  assign \new_[67314]_  = ~A300 & \new_[67313]_ ;
  assign \new_[67315]_  = \new_[67314]_  & \new_[67309]_ ;
  assign \new_[67316]_  = \new_[67315]_  & \new_[67306]_ ;
  assign \new_[67319]_  = ~A169 & ~A170;
  assign \new_[67322]_  = ~A167 & ~A168;
  assign \new_[67323]_  = \new_[67322]_  & \new_[67319]_ ;
  assign \new_[67326]_  = A232 & A166;
  assign \new_[67329]_  = ~A234 & ~A233;
  assign \new_[67330]_  = \new_[67329]_  & \new_[67326]_ ;
  assign \new_[67331]_  = \new_[67330]_  & \new_[67323]_ ;
  assign \new_[67334]_  = A236 & ~A235;
  assign \new_[67337]_  = ~A268 & A267;
  assign \new_[67338]_  = \new_[67337]_  & \new_[67334]_ ;
  assign \new_[67341]_  = A298 & A269;
  assign \new_[67345]_  = A301 & A300;
  assign \new_[67346]_  = ~A299 & \new_[67345]_ ;
  assign \new_[67347]_  = \new_[67346]_  & \new_[67341]_ ;
  assign \new_[67348]_  = \new_[67347]_  & \new_[67338]_ ;
  assign \new_[67351]_  = ~A169 & ~A170;
  assign \new_[67354]_  = ~A167 & ~A168;
  assign \new_[67355]_  = \new_[67354]_  & \new_[67351]_ ;
  assign \new_[67358]_  = A232 & A166;
  assign \new_[67361]_  = ~A234 & ~A233;
  assign \new_[67362]_  = \new_[67361]_  & \new_[67358]_ ;
  assign \new_[67363]_  = \new_[67362]_  & \new_[67355]_ ;
  assign \new_[67366]_  = A236 & ~A235;
  assign \new_[67369]_  = ~A268 & A267;
  assign \new_[67370]_  = \new_[67369]_  & \new_[67366]_ ;
  assign \new_[67373]_  = A298 & A269;
  assign \new_[67377]_  = ~A302 & A300;
  assign \new_[67378]_  = ~A299 & \new_[67377]_ ;
  assign \new_[67379]_  = \new_[67378]_  & \new_[67373]_ ;
  assign \new_[67380]_  = \new_[67379]_  & \new_[67370]_ ;
  assign \new_[67383]_  = ~A169 & ~A170;
  assign \new_[67386]_  = ~A167 & ~A168;
  assign \new_[67387]_  = \new_[67386]_  & \new_[67383]_ ;
  assign \new_[67390]_  = A232 & A166;
  assign \new_[67393]_  = ~A234 & ~A233;
  assign \new_[67394]_  = \new_[67393]_  & \new_[67390]_ ;
  assign \new_[67395]_  = \new_[67394]_  & \new_[67387]_ ;
  assign \new_[67398]_  = A236 & ~A235;
  assign \new_[67401]_  = ~A268 & A267;
  assign \new_[67402]_  = \new_[67401]_  & \new_[67398]_ ;
  assign \new_[67405]_  = ~A298 & A269;
  assign \new_[67409]_  = A301 & A300;
  assign \new_[67410]_  = A299 & \new_[67409]_ ;
  assign \new_[67411]_  = \new_[67410]_  & \new_[67405]_ ;
  assign \new_[67412]_  = \new_[67411]_  & \new_[67402]_ ;
  assign \new_[67415]_  = ~A169 & ~A170;
  assign \new_[67418]_  = ~A167 & ~A168;
  assign \new_[67419]_  = \new_[67418]_  & \new_[67415]_ ;
  assign \new_[67422]_  = A232 & A166;
  assign \new_[67425]_  = ~A234 & ~A233;
  assign \new_[67426]_  = \new_[67425]_  & \new_[67422]_ ;
  assign \new_[67427]_  = \new_[67426]_  & \new_[67419]_ ;
  assign \new_[67430]_  = A236 & ~A235;
  assign \new_[67433]_  = ~A268 & A267;
  assign \new_[67434]_  = \new_[67433]_  & \new_[67430]_ ;
  assign \new_[67437]_  = ~A298 & A269;
  assign \new_[67441]_  = ~A302 & A300;
  assign \new_[67442]_  = A299 & \new_[67441]_ ;
  assign \new_[67443]_  = \new_[67442]_  & \new_[67437]_ ;
  assign \new_[67444]_  = \new_[67443]_  & \new_[67434]_ ;
  assign \new_[67447]_  = ~A169 & ~A170;
  assign \new_[67450]_  = ~A167 & ~A168;
  assign \new_[67451]_  = \new_[67450]_  & \new_[67447]_ ;
  assign \new_[67454]_  = A232 & A166;
  assign \new_[67457]_  = ~A234 & ~A233;
  assign \new_[67458]_  = \new_[67457]_  & \new_[67454]_ ;
  assign \new_[67459]_  = \new_[67458]_  & \new_[67451]_ ;
  assign \new_[67462]_  = A236 & ~A235;
  assign \new_[67465]_  = A268 & ~A267;
  assign \new_[67466]_  = \new_[67465]_  & \new_[67462]_ ;
  assign \new_[67469]_  = ~A299 & A298;
  assign \new_[67473]_  = A302 & ~A301;
  assign \new_[67474]_  = ~A300 & \new_[67473]_ ;
  assign \new_[67475]_  = \new_[67474]_  & \new_[67469]_ ;
  assign \new_[67476]_  = \new_[67475]_  & \new_[67466]_ ;
  assign \new_[67479]_  = ~A169 & ~A170;
  assign \new_[67482]_  = ~A167 & ~A168;
  assign \new_[67483]_  = \new_[67482]_  & \new_[67479]_ ;
  assign \new_[67486]_  = A232 & A166;
  assign \new_[67489]_  = ~A234 & ~A233;
  assign \new_[67490]_  = \new_[67489]_  & \new_[67486]_ ;
  assign \new_[67491]_  = \new_[67490]_  & \new_[67483]_ ;
  assign \new_[67494]_  = A236 & ~A235;
  assign \new_[67497]_  = A268 & ~A267;
  assign \new_[67498]_  = \new_[67497]_  & \new_[67494]_ ;
  assign \new_[67501]_  = A299 & ~A298;
  assign \new_[67505]_  = A302 & ~A301;
  assign \new_[67506]_  = ~A300 & \new_[67505]_ ;
  assign \new_[67507]_  = \new_[67506]_  & \new_[67501]_ ;
  assign \new_[67508]_  = \new_[67507]_  & \new_[67498]_ ;
  assign \new_[67511]_  = ~A169 & ~A170;
  assign \new_[67514]_  = ~A167 & ~A168;
  assign \new_[67515]_  = \new_[67514]_  & \new_[67511]_ ;
  assign \new_[67518]_  = A232 & A166;
  assign \new_[67521]_  = ~A234 & ~A233;
  assign \new_[67522]_  = \new_[67521]_  & \new_[67518]_ ;
  assign \new_[67523]_  = \new_[67522]_  & \new_[67515]_ ;
  assign \new_[67526]_  = A236 & ~A235;
  assign \new_[67529]_  = ~A269 & ~A267;
  assign \new_[67530]_  = \new_[67529]_  & \new_[67526]_ ;
  assign \new_[67533]_  = ~A299 & A298;
  assign \new_[67537]_  = A302 & ~A301;
  assign \new_[67538]_  = ~A300 & \new_[67537]_ ;
  assign \new_[67539]_  = \new_[67538]_  & \new_[67533]_ ;
  assign \new_[67540]_  = \new_[67539]_  & \new_[67530]_ ;
  assign \new_[67543]_  = ~A169 & ~A170;
  assign \new_[67546]_  = ~A167 & ~A168;
  assign \new_[67547]_  = \new_[67546]_  & \new_[67543]_ ;
  assign \new_[67550]_  = A232 & A166;
  assign \new_[67553]_  = ~A234 & ~A233;
  assign \new_[67554]_  = \new_[67553]_  & \new_[67550]_ ;
  assign \new_[67555]_  = \new_[67554]_  & \new_[67547]_ ;
  assign \new_[67558]_  = A236 & ~A235;
  assign \new_[67561]_  = ~A269 & ~A267;
  assign \new_[67562]_  = \new_[67561]_  & \new_[67558]_ ;
  assign \new_[67565]_  = A299 & ~A298;
  assign \new_[67569]_  = A302 & ~A301;
  assign \new_[67570]_  = ~A300 & \new_[67569]_ ;
  assign \new_[67571]_  = \new_[67570]_  & \new_[67565]_ ;
  assign \new_[67572]_  = \new_[67571]_  & \new_[67562]_ ;
  assign \new_[67575]_  = ~A169 & ~A170;
  assign \new_[67578]_  = ~A167 & ~A168;
  assign \new_[67579]_  = \new_[67578]_  & \new_[67575]_ ;
  assign \new_[67582]_  = A232 & A166;
  assign \new_[67585]_  = ~A234 & ~A233;
  assign \new_[67586]_  = \new_[67585]_  & \new_[67582]_ ;
  assign \new_[67587]_  = \new_[67586]_  & \new_[67579]_ ;
  assign \new_[67590]_  = A236 & ~A235;
  assign \new_[67593]_  = A266 & A265;
  assign \new_[67594]_  = \new_[67593]_  & \new_[67590]_ ;
  assign \new_[67597]_  = ~A299 & A298;
  assign \new_[67601]_  = A302 & ~A301;
  assign \new_[67602]_  = ~A300 & \new_[67601]_ ;
  assign \new_[67603]_  = \new_[67602]_  & \new_[67597]_ ;
  assign \new_[67604]_  = \new_[67603]_  & \new_[67594]_ ;
  assign \new_[67607]_  = ~A169 & ~A170;
  assign \new_[67610]_  = ~A167 & ~A168;
  assign \new_[67611]_  = \new_[67610]_  & \new_[67607]_ ;
  assign \new_[67614]_  = A232 & A166;
  assign \new_[67617]_  = ~A234 & ~A233;
  assign \new_[67618]_  = \new_[67617]_  & \new_[67614]_ ;
  assign \new_[67619]_  = \new_[67618]_  & \new_[67611]_ ;
  assign \new_[67622]_  = A236 & ~A235;
  assign \new_[67625]_  = A266 & A265;
  assign \new_[67626]_  = \new_[67625]_  & \new_[67622]_ ;
  assign \new_[67629]_  = A299 & ~A298;
  assign \new_[67633]_  = A302 & ~A301;
  assign \new_[67634]_  = ~A300 & \new_[67633]_ ;
  assign \new_[67635]_  = \new_[67634]_  & \new_[67629]_ ;
  assign \new_[67636]_  = \new_[67635]_  & \new_[67626]_ ;
  assign \new_[67639]_  = ~A169 & ~A170;
  assign \new_[67642]_  = ~A167 & ~A168;
  assign \new_[67643]_  = \new_[67642]_  & \new_[67639]_ ;
  assign \new_[67646]_  = A232 & A166;
  assign \new_[67649]_  = ~A234 & ~A233;
  assign \new_[67650]_  = \new_[67649]_  & \new_[67646]_ ;
  assign \new_[67651]_  = \new_[67650]_  & \new_[67643]_ ;
  assign \new_[67654]_  = A236 & ~A235;
  assign \new_[67657]_  = ~A266 & ~A265;
  assign \new_[67658]_  = \new_[67657]_  & \new_[67654]_ ;
  assign \new_[67661]_  = ~A299 & A298;
  assign \new_[67665]_  = A302 & ~A301;
  assign \new_[67666]_  = ~A300 & \new_[67665]_ ;
  assign \new_[67667]_  = \new_[67666]_  & \new_[67661]_ ;
  assign \new_[67668]_  = \new_[67667]_  & \new_[67658]_ ;
  assign \new_[67671]_  = ~A169 & ~A170;
  assign \new_[67674]_  = ~A167 & ~A168;
  assign \new_[67675]_  = \new_[67674]_  & \new_[67671]_ ;
  assign \new_[67678]_  = A232 & A166;
  assign \new_[67681]_  = ~A234 & ~A233;
  assign \new_[67682]_  = \new_[67681]_  & \new_[67678]_ ;
  assign \new_[67683]_  = \new_[67682]_  & \new_[67675]_ ;
  assign \new_[67686]_  = A236 & ~A235;
  assign \new_[67689]_  = ~A266 & ~A265;
  assign \new_[67690]_  = \new_[67689]_  & \new_[67686]_ ;
  assign \new_[67693]_  = A299 & ~A298;
  assign \new_[67697]_  = A302 & ~A301;
  assign \new_[67698]_  = ~A300 & \new_[67697]_ ;
  assign \new_[67699]_  = \new_[67698]_  & \new_[67693]_ ;
  assign \new_[67700]_  = \new_[67699]_  & \new_[67690]_ ;
  assign \new_[67703]_  = A200 & ~A199;
  assign \new_[67706]_  = ~A202 & ~A201;
  assign \new_[67707]_  = \new_[67706]_  & \new_[67703]_ ;
  assign \new_[67710]_  = ~A232 & A203;
  assign \new_[67714]_  = ~A235 & ~A234;
  assign \new_[67715]_  = A233 & \new_[67714]_ ;
  assign \new_[67716]_  = \new_[67715]_  & \new_[67710]_ ;
  assign \new_[67717]_  = \new_[67716]_  & \new_[67707]_ ;
  assign \new_[67720]_  = A267 & A236;
  assign \new_[67723]_  = A269 & ~A268;
  assign \new_[67724]_  = \new_[67723]_  & \new_[67720]_ ;
  assign \new_[67727]_  = ~A299 & A298;
  assign \new_[67731]_  = A302 & ~A301;
  assign \new_[67732]_  = ~A300 & \new_[67731]_ ;
  assign \new_[67733]_  = \new_[67732]_  & \new_[67727]_ ;
  assign \new_[67734]_  = \new_[67733]_  & \new_[67724]_ ;
  assign \new_[67737]_  = A200 & ~A199;
  assign \new_[67740]_  = ~A202 & ~A201;
  assign \new_[67741]_  = \new_[67740]_  & \new_[67737]_ ;
  assign \new_[67744]_  = ~A232 & A203;
  assign \new_[67748]_  = ~A235 & ~A234;
  assign \new_[67749]_  = A233 & \new_[67748]_ ;
  assign \new_[67750]_  = \new_[67749]_  & \new_[67744]_ ;
  assign \new_[67751]_  = \new_[67750]_  & \new_[67741]_ ;
  assign \new_[67754]_  = A267 & A236;
  assign \new_[67757]_  = A269 & ~A268;
  assign \new_[67758]_  = \new_[67757]_  & \new_[67754]_ ;
  assign \new_[67761]_  = A299 & ~A298;
  assign \new_[67765]_  = A302 & ~A301;
  assign \new_[67766]_  = ~A300 & \new_[67765]_ ;
  assign \new_[67767]_  = \new_[67766]_  & \new_[67761]_ ;
  assign \new_[67768]_  = \new_[67767]_  & \new_[67758]_ ;
  assign \new_[67771]_  = A200 & ~A199;
  assign \new_[67774]_  = ~A202 & ~A201;
  assign \new_[67775]_  = \new_[67774]_  & \new_[67771]_ ;
  assign \new_[67778]_  = A232 & A203;
  assign \new_[67782]_  = ~A235 & ~A234;
  assign \new_[67783]_  = ~A233 & \new_[67782]_ ;
  assign \new_[67784]_  = \new_[67783]_  & \new_[67778]_ ;
  assign \new_[67785]_  = \new_[67784]_  & \new_[67775]_ ;
  assign \new_[67788]_  = A267 & A236;
  assign \new_[67791]_  = A269 & ~A268;
  assign \new_[67792]_  = \new_[67791]_  & \new_[67788]_ ;
  assign \new_[67795]_  = ~A299 & A298;
  assign \new_[67799]_  = A302 & ~A301;
  assign \new_[67800]_  = ~A300 & \new_[67799]_ ;
  assign \new_[67801]_  = \new_[67800]_  & \new_[67795]_ ;
  assign \new_[67802]_  = \new_[67801]_  & \new_[67792]_ ;
  assign \new_[67805]_  = A200 & ~A199;
  assign \new_[67808]_  = ~A202 & ~A201;
  assign \new_[67809]_  = \new_[67808]_  & \new_[67805]_ ;
  assign \new_[67812]_  = A232 & A203;
  assign \new_[67816]_  = ~A235 & ~A234;
  assign \new_[67817]_  = ~A233 & \new_[67816]_ ;
  assign \new_[67818]_  = \new_[67817]_  & \new_[67812]_ ;
  assign \new_[67819]_  = \new_[67818]_  & \new_[67809]_ ;
  assign \new_[67822]_  = A267 & A236;
  assign \new_[67825]_  = A269 & ~A268;
  assign \new_[67826]_  = \new_[67825]_  & \new_[67822]_ ;
  assign \new_[67829]_  = A299 & ~A298;
  assign \new_[67833]_  = A302 & ~A301;
  assign \new_[67834]_  = ~A300 & \new_[67833]_ ;
  assign \new_[67835]_  = \new_[67834]_  & \new_[67829]_ ;
  assign \new_[67836]_  = \new_[67835]_  & \new_[67826]_ ;
  assign \new_[67839]_  = ~A200 & A199;
  assign \new_[67842]_  = ~A202 & ~A201;
  assign \new_[67843]_  = \new_[67842]_  & \new_[67839]_ ;
  assign \new_[67846]_  = ~A232 & A203;
  assign \new_[67850]_  = ~A235 & ~A234;
  assign \new_[67851]_  = A233 & \new_[67850]_ ;
  assign \new_[67852]_  = \new_[67851]_  & \new_[67846]_ ;
  assign \new_[67853]_  = \new_[67852]_  & \new_[67843]_ ;
  assign \new_[67856]_  = A267 & A236;
  assign \new_[67859]_  = A269 & ~A268;
  assign \new_[67860]_  = \new_[67859]_  & \new_[67856]_ ;
  assign \new_[67863]_  = ~A299 & A298;
  assign \new_[67867]_  = A302 & ~A301;
  assign \new_[67868]_  = ~A300 & \new_[67867]_ ;
  assign \new_[67869]_  = \new_[67868]_  & \new_[67863]_ ;
  assign \new_[67870]_  = \new_[67869]_  & \new_[67860]_ ;
  assign \new_[67873]_  = ~A200 & A199;
  assign \new_[67876]_  = ~A202 & ~A201;
  assign \new_[67877]_  = \new_[67876]_  & \new_[67873]_ ;
  assign \new_[67880]_  = ~A232 & A203;
  assign \new_[67884]_  = ~A235 & ~A234;
  assign \new_[67885]_  = A233 & \new_[67884]_ ;
  assign \new_[67886]_  = \new_[67885]_  & \new_[67880]_ ;
  assign \new_[67887]_  = \new_[67886]_  & \new_[67877]_ ;
  assign \new_[67890]_  = A267 & A236;
  assign \new_[67893]_  = A269 & ~A268;
  assign \new_[67894]_  = \new_[67893]_  & \new_[67890]_ ;
  assign \new_[67897]_  = A299 & ~A298;
  assign \new_[67901]_  = A302 & ~A301;
  assign \new_[67902]_  = ~A300 & \new_[67901]_ ;
  assign \new_[67903]_  = \new_[67902]_  & \new_[67897]_ ;
  assign \new_[67904]_  = \new_[67903]_  & \new_[67894]_ ;
  assign \new_[67907]_  = ~A200 & A199;
  assign \new_[67910]_  = ~A202 & ~A201;
  assign \new_[67911]_  = \new_[67910]_  & \new_[67907]_ ;
  assign \new_[67914]_  = A232 & A203;
  assign \new_[67918]_  = ~A235 & ~A234;
  assign \new_[67919]_  = ~A233 & \new_[67918]_ ;
  assign \new_[67920]_  = \new_[67919]_  & \new_[67914]_ ;
  assign \new_[67921]_  = \new_[67920]_  & \new_[67911]_ ;
  assign \new_[67924]_  = A267 & A236;
  assign \new_[67927]_  = A269 & ~A268;
  assign \new_[67928]_  = \new_[67927]_  & \new_[67924]_ ;
  assign \new_[67931]_  = ~A299 & A298;
  assign \new_[67935]_  = A302 & ~A301;
  assign \new_[67936]_  = ~A300 & \new_[67935]_ ;
  assign \new_[67937]_  = \new_[67936]_  & \new_[67931]_ ;
  assign \new_[67938]_  = \new_[67937]_  & \new_[67928]_ ;
  assign \new_[67941]_  = ~A200 & A199;
  assign \new_[67944]_  = ~A202 & ~A201;
  assign \new_[67945]_  = \new_[67944]_  & \new_[67941]_ ;
  assign \new_[67948]_  = A232 & A203;
  assign \new_[67952]_  = ~A235 & ~A234;
  assign \new_[67953]_  = ~A233 & \new_[67952]_ ;
  assign \new_[67954]_  = \new_[67953]_  & \new_[67948]_ ;
  assign \new_[67955]_  = \new_[67954]_  & \new_[67945]_ ;
  assign \new_[67958]_  = A267 & A236;
  assign \new_[67961]_  = A269 & ~A268;
  assign \new_[67962]_  = \new_[67961]_  & \new_[67958]_ ;
  assign \new_[67965]_  = A299 & ~A298;
  assign \new_[67969]_  = A302 & ~A301;
  assign \new_[67970]_  = ~A300 & \new_[67969]_ ;
  assign \new_[67971]_  = \new_[67970]_  & \new_[67965]_ ;
  assign \new_[67972]_  = \new_[67971]_  & \new_[67962]_ ;
  assign \new_[67975]_  = ~A169 & ~A170;
  assign \new_[67978]_  = A167 & ~A168;
  assign \new_[67979]_  = \new_[67978]_  & \new_[67975]_ ;
  assign \new_[67982]_  = ~A232 & ~A166;
  assign \new_[67986]_  = ~A235 & ~A234;
  assign \new_[67987]_  = A233 & \new_[67986]_ ;
  assign \new_[67988]_  = \new_[67987]_  & \new_[67982]_ ;
  assign \new_[67989]_  = \new_[67988]_  & \new_[67979]_ ;
  assign \new_[67992]_  = A267 & A236;
  assign \new_[67995]_  = A269 & ~A268;
  assign \new_[67996]_  = \new_[67995]_  & \new_[67992]_ ;
  assign \new_[67999]_  = ~A299 & A298;
  assign \new_[68003]_  = A302 & ~A301;
  assign \new_[68004]_  = ~A300 & \new_[68003]_ ;
  assign \new_[68005]_  = \new_[68004]_  & \new_[67999]_ ;
  assign \new_[68006]_  = \new_[68005]_  & \new_[67996]_ ;
  assign \new_[68009]_  = ~A169 & ~A170;
  assign \new_[68012]_  = A167 & ~A168;
  assign \new_[68013]_  = \new_[68012]_  & \new_[68009]_ ;
  assign \new_[68016]_  = ~A232 & ~A166;
  assign \new_[68020]_  = ~A235 & ~A234;
  assign \new_[68021]_  = A233 & \new_[68020]_ ;
  assign \new_[68022]_  = \new_[68021]_  & \new_[68016]_ ;
  assign \new_[68023]_  = \new_[68022]_  & \new_[68013]_ ;
  assign \new_[68026]_  = A267 & A236;
  assign \new_[68029]_  = A269 & ~A268;
  assign \new_[68030]_  = \new_[68029]_  & \new_[68026]_ ;
  assign \new_[68033]_  = A299 & ~A298;
  assign \new_[68037]_  = A302 & ~A301;
  assign \new_[68038]_  = ~A300 & \new_[68037]_ ;
  assign \new_[68039]_  = \new_[68038]_  & \new_[68033]_ ;
  assign \new_[68040]_  = \new_[68039]_  & \new_[68030]_ ;
  assign \new_[68043]_  = ~A169 & ~A170;
  assign \new_[68046]_  = A167 & ~A168;
  assign \new_[68047]_  = \new_[68046]_  & \new_[68043]_ ;
  assign \new_[68050]_  = A232 & ~A166;
  assign \new_[68054]_  = ~A235 & ~A234;
  assign \new_[68055]_  = ~A233 & \new_[68054]_ ;
  assign \new_[68056]_  = \new_[68055]_  & \new_[68050]_ ;
  assign \new_[68057]_  = \new_[68056]_  & \new_[68047]_ ;
  assign \new_[68060]_  = A267 & A236;
  assign \new_[68063]_  = A269 & ~A268;
  assign \new_[68064]_  = \new_[68063]_  & \new_[68060]_ ;
  assign \new_[68067]_  = ~A299 & A298;
  assign \new_[68071]_  = A302 & ~A301;
  assign \new_[68072]_  = ~A300 & \new_[68071]_ ;
  assign \new_[68073]_  = \new_[68072]_  & \new_[68067]_ ;
  assign \new_[68074]_  = \new_[68073]_  & \new_[68064]_ ;
  assign \new_[68077]_  = ~A169 & ~A170;
  assign \new_[68080]_  = A167 & ~A168;
  assign \new_[68081]_  = \new_[68080]_  & \new_[68077]_ ;
  assign \new_[68084]_  = A232 & ~A166;
  assign \new_[68088]_  = ~A235 & ~A234;
  assign \new_[68089]_  = ~A233 & \new_[68088]_ ;
  assign \new_[68090]_  = \new_[68089]_  & \new_[68084]_ ;
  assign \new_[68091]_  = \new_[68090]_  & \new_[68081]_ ;
  assign \new_[68094]_  = A267 & A236;
  assign \new_[68097]_  = A269 & ~A268;
  assign \new_[68098]_  = \new_[68097]_  & \new_[68094]_ ;
  assign \new_[68101]_  = A299 & ~A298;
  assign \new_[68105]_  = A302 & ~A301;
  assign \new_[68106]_  = ~A300 & \new_[68105]_ ;
  assign \new_[68107]_  = \new_[68106]_  & \new_[68101]_ ;
  assign \new_[68108]_  = \new_[68107]_  & \new_[68098]_ ;
  assign \new_[68111]_  = ~A169 & ~A170;
  assign \new_[68114]_  = ~A167 & ~A168;
  assign \new_[68115]_  = \new_[68114]_  & \new_[68111]_ ;
  assign \new_[68118]_  = ~A232 & A166;
  assign \new_[68122]_  = ~A235 & ~A234;
  assign \new_[68123]_  = A233 & \new_[68122]_ ;
  assign \new_[68124]_  = \new_[68123]_  & \new_[68118]_ ;
  assign \new_[68125]_  = \new_[68124]_  & \new_[68115]_ ;
  assign \new_[68128]_  = A267 & A236;
  assign \new_[68131]_  = A269 & ~A268;
  assign \new_[68132]_  = \new_[68131]_  & \new_[68128]_ ;
  assign \new_[68135]_  = ~A299 & A298;
  assign \new_[68139]_  = A302 & ~A301;
  assign \new_[68140]_  = ~A300 & \new_[68139]_ ;
  assign \new_[68141]_  = \new_[68140]_  & \new_[68135]_ ;
  assign \new_[68142]_  = \new_[68141]_  & \new_[68132]_ ;
  assign \new_[68145]_  = ~A169 & ~A170;
  assign \new_[68148]_  = ~A167 & ~A168;
  assign \new_[68149]_  = \new_[68148]_  & \new_[68145]_ ;
  assign \new_[68152]_  = ~A232 & A166;
  assign \new_[68156]_  = ~A235 & ~A234;
  assign \new_[68157]_  = A233 & \new_[68156]_ ;
  assign \new_[68158]_  = \new_[68157]_  & \new_[68152]_ ;
  assign \new_[68159]_  = \new_[68158]_  & \new_[68149]_ ;
  assign \new_[68162]_  = A267 & A236;
  assign \new_[68165]_  = A269 & ~A268;
  assign \new_[68166]_  = \new_[68165]_  & \new_[68162]_ ;
  assign \new_[68169]_  = A299 & ~A298;
  assign \new_[68173]_  = A302 & ~A301;
  assign \new_[68174]_  = ~A300 & \new_[68173]_ ;
  assign \new_[68175]_  = \new_[68174]_  & \new_[68169]_ ;
  assign \new_[68176]_  = \new_[68175]_  & \new_[68166]_ ;
  assign \new_[68179]_  = ~A169 & ~A170;
  assign \new_[68182]_  = ~A167 & ~A168;
  assign \new_[68183]_  = \new_[68182]_  & \new_[68179]_ ;
  assign \new_[68186]_  = A232 & A166;
  assign \new_[68190]_  = ~A235 & ~A234;
  assign \new_[68191]_  = ~A233 & \new_[68190]_ ;
  assign \new_[68192]_  = \new_[68191]_  & \new_[68186]_ ;
  assign \new_[68193]_  = \new_[68192]_  & \new_[68183]_ ;
  assign \new_[68196]_  = A267 & A236;
  assign \new_[68199]_  = A269 & ~A268;
  assign \new_[68200]_  = \new_[68199]_  & \new_[68196]_ ;
  assign \new_[68203]_  = ~A299 & A298;
  assign \new_[68207]_  = A302 & ~A301;
  assign \new_[68208]_  = ~A300 & \new_[68207]_ ;
  assign \new_[68209]_  = \new_[68208]_  & \new_[68203]_ ;
  assign \new_[68210]_  = \new_[68209]_  & \new_[68200]_ ;
  assign \new_[68213]_  = ~A169 & ~A170;
  assign \new_[68216]_  = ~A167 & ~A168;
  assign \new_[68217]_  = \new_[68216]_  & \new_[68213]_ ;
  assign \new_[68220]_  = A232 & A166;
  assign \new_[68224]_  = ~A235 & ~A234;
  assign \new_[68225]_  = ~A233 & \new_[68224]_ ;
  assign \new_[68226]_  = \new_[68225]_  & \new_[68220]_ ;
  assign \new_[68227]_  = \new_[68226]_  & \new_[68217]_ ;
  assign \new_[68230]_  = A267 & A236;
  assign \new_[68233]_  = A269 & ~A268;
  assign \new_[68234]_  = \new_[68233]_  & \new_[68230]_ ;
  assign \new_[68237]_  = A299 & ~A298;
  assign \new_[68241]_  = A302 & ~A301;
  assign \new_[68242]_  = ~A300 & \new_[68241]_ ;
  assign \new_[68243]_  = \new_[68242]_  & \new_[68237]_ ;
  assign \new_[68244]_  = \new_[68243]_  & \new_[68234]_ ;
endmodule


