// Benchmark "testing" written by ABC on Thu Oct  8 22:16:32 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A43  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A43;
  wire new_n_32_, new_n_33_, new_n_37_, new_n_38_, new_n_39_, new_n_40_,
    new_n_46_, new_n_47_, new_n_48_, new_n_49_, new_n_55_, new_n_56_,
    new_n_57_, new_n_58_, new_n_59_, new_n_60_, new_n_66_, new_n_67_,
    new_n_68_, new_n_69_, new_n_72_, new_n_73_, new_n_74_, new_n_81_,
    new_n_82_, new_n_83_, new_n_84_, new_n_87_, new_n_88_, new_n_91_,
    new_n_94_, new_n_97_, new_n_98_, new_n_99_, new_n_104_, new_n_105_,
    new_n_106_, new_n_107_, new_n_108_, new_n_109_, new_n_114_, new_n_120_,
    new_n_121_, new_n_122_, new_n_123_, new_n_126_, new_n_127_, new_n_128_,
    new_n_129_, new_n_130_, new_n_135_, new_n_136_, new_n_140_, new_n_141_,
    new_n_142_, new_n_143_, new_n_149_, new_n_150_, new_n_151_, new_n_152_,
    new_n_158_, new_n_159_, new_n_160_, new_n_161_, new_n_166_, new_n_167_,
    new_n_171_, new_n_172_, new_n_173_, new_n_174_, new_n_180_, new_n_181_,
    new_n_182_, new_n_183_, new_n_189_, new_n_190_, new_n_191_, new_n_192_,
    new_n_193_, new_n_194_, new_n_195_, new_n_196_, new_n_197_, new_n_201_,
    new_n_204_, new_n_207_, new_n_208_, new_n_209_, new_n_214_, new_n_215_,
    new_n_216_, new_n_217_, new_n_218_, new_n_223_, new_n_224_, new_n_225_,
    new_n_226_, new_n_227_, new_n_234_, new_n_235_, new_n_239_, new_n_240_,
    new_n_241_, new_n_242_, new_n_248_, new_n_249_, new_n_250_, new_n_251_,
    new_n_257_, new_n_258_, new_n_259_, new_n_260_, new_n_261_, new_n_262_,
    new_n_265_, new_n_268_, new_n_271_, new_n_272_, new_n_275_, new_n_278_,
    new_n_281_, new_n_282_, new_n_283_, new_n_288_, new_n_289_, new_n_290_,
    new_n_291_, new_n_292_, new_n_293_, new_n_298_, new_n_301_, new_n_304_,
    new_n_307_, new_n_308_, new_n_309_, new_n_314_, new_n_315_, new_n_316_,
    new_n_317_, new_n_318_, new_n_319_, new_n_320_, new_n_321_, new_n_322_,
    new_n_323_, new_n_328_, new_n_333_, new_n_334_, new_n_338_, new_n_339_,
    new_n_340_, new_n_341_, new_n_347_, new_n_348_, new_n_349_, new_n_350_,
    new_n_356_, new_n_357_, new_n_358_, new_n_359_, new_n_360_, new_n_361_,
    new_n_364_, new_n_367_, new_n_370_, new_n_371_, new_n_372_, new_n_377_,
    new_n_378_, new_n_379_, new_n_380_, new_n_381_, new_n_382_, new_n_383_,
    new_n_384_, new_n_385_, new_n_386_, new_n_391_, new_n_397_, new_n_398_,
    new_n_402_, new_n_403_, new_n_404_, new_n_405_, new_n_411_, new_n_412_,
    new_n_413_, new_n_414_, new_n_420_, new_n_421_, new_n_422_, new_n_423_,
    new_n_424_, new_n_425_, new_n_428_, new_n_431_, new_n_434_, new_n_435_,
    new_n_436_, new_n_441_, new_n_442_, new_n_443_, new_n_444_, new_n_445_,
    new_n_446_, new_n_451_, new_n_456_, new_n_457_, new_n_461_, new_n_462_,
    new_n_463_, new_n_464_, new_n_470_, new_n_471_, new_n_472_, new_n_473_,
    new_n_479_, new_n_480_, new_n_481_, new_n_482_, new_n_483_, new_n_484_,
    new_n_485_, new_n_486_, new_n_487_, new_n_488_, new_n_489_, new_n_490_,
    new_n_491_, new_n_492_, new_n_493_, new_n_494_, new_n_495_, new_n_496_;
  assign A43 = ~new_n_496_;
  assign new_n_32_ = ~A202 & A203;
  assign new_n_33_ = A200 & new_n_32_;
  assign new_n_37_ = A202 & ~A203;
  assign new_n_38_ = ~A200 & new_n_37_;
  assign new_n_39_ = new_n_33_ | new_n_38_;
  assign new_n_40_ = ~A199 & new_n_39_;
  assign new_n_46_ = A202 & ~A203;
  assign new_n_47_ = A199 & new_n_46_;
  assign new_n_48_ = A201 | new_n_47_;
  assign new_n_49_ = A200 & new_n_48_;
  assign new_n_55_ = ~A202 & A203;
  assign new_n_56_ = ~A200 & new_n_55_;
  assign new_n_57_ = A201 | new_n_56_;
  assign new_n_58_ = A199 & new_n_57_;
  assign new_n_59_ = new_n_49_ | new_n_58_;
  assign new_n_60_ = new_n_40_ | new_n_59_;
  assign new_n_66_ = A169 | A170;
  assign new_n_67_ = A168 & new_n_66_;
  assign new_n_68_ = ~A167 & new_n_67_;
  assign new_n_69_ = A166 & new_n_68_;
  assign new_n_72_ = ~A166 & A167;
  assign new_n_73_ = new_n_69_ | new_n_72_;
  assign new_n_74_ = new_n_60_ & new_n_73_;
  assign new_n_81_ = ~A169 & ~A170;
  assign new_n_82_ = ~A168 | new_n_81_;
  assign new_n_83_ = ~A166 | new_n_82_;
  assign new_n_84_ = ~A167 & new_n_83_;
  assign new_n_87_ = A166 & A167;
  assign new_n_88_ = new_n_84_ | new_n_87_;
  assign new_n_91_ = A202 | ~A203;
  assign new_n_94_ = ~A199 & A200;
  assign new_n_97_ = A199 & ~A200;
  assign new_n_98_ = new_n_94_ | new_n_97_;
  assign new_n_99_ = new_n_91_ & new_n_98_;
  assign new_n_104_ = ~A202 | A203;
  assign new_n_105_ = A200 & new_n_104_;
  assign new_n_106_ = A199 & new_n_105_;
  assign new_n_107_ = new_n_99_ | new_n_106_;
  assign new_n_108_ = new_n_88_ & new_n_107_;
  assign new_n_109_ = ~A201 & new_n_108_;
  assign new_n_114_ = ~A202 | A203;
  assign new_n_120_ = ~A169 & ~A170;
  assign new_n_121_ = ~A168 | new_n_120_;
  assign new_n_122_ = ~A166 | new_n_121_;
  assign new_n_123_ = ~A167 & new_n_122_;
  assign new_n_126_ = A166 & A167;
  assign new_n_127_ = new_n_123_ | new_n_126_;
  assign new_n_128_ = new_n_114_ & new_n_127_;
  assign new_n_129_ = ~A200 & new_n_128_;
  assign new_n_130_ = ~A199 & new_n_129_;
  assign new_n_135_ = ~A268 & A269;
  assign new_n_136_ = A266 & new_n_135_;
  assign new_n_140_ = A268 & ~A269;
  assign new_n_141_ = ~A266 & new_n_140_;
  assign new_n_142_ = new_n_136_ | new_n_141_;
  assign new_n_143_ = ~A265 & new_n_142_;
  assign new_n_149_ = A268 & ~A269;
  assign new_n_150_ = A265 & new_n_149_;
  assign new_n_151_ = A267 | new_n_150_;
  assign new_n_152_ = A266 & new_n_151_;
  assign new_n_158_ = ~A268 & A269;
  assign new_n_159_ = ~A266 & new_n_158_;
  assign new_n_160_ = A267 | new_n_159_;
  assign new_n_161_ = A265 & new_n_160_;
  assign new_n_166_ = ~A301 & A302;
  assign new_n_167_ = A299 & new_n_166_;
  assign new_n_171_ = A301 & ~A302;
  assign new_n_172_ = ~A299 & new_n_171_;
  assign new_n_173_ = new_n_167_ | new_n_172_;
  assign new_n_174_ = ~A298 & new_n_173_;
  assign new_n_180_ = A301 & ~A302;
  assign new_n_181_ = A298 & new_n_180_;
  assign new_n_182_ = A300 | new_n_181_;
  assign new_n_183_ = A299 & new_n_182_;
  assign new_n_189_ = ~A301 & A302;
  assign new_n_190_ = ~A299 & new_n_189_;
  assign new_n_191_ = A300 | new_n_190_;
  assign new_n_192_ = A298 & new_n_191_;
  assign new_n_193_ = new_n_183_ | new_n_192_;
  assign new_n_194_ = new_n_174_ | new_n_193_;
  assign new_n_195_ = new_n_161_ | new_n_194_;
  assign new_n_196_ = new_n_152_ | new_n_195_;
  assign new_n_197_ = new_n_143_ | new_n_196_;
  assign new_n_201_ = A235 | ~A236;
  assign new_n_204_ = ~A232 & A233;
  assign new_n_207_ = A232 & ~A233;
  assign new_n_208_ = new_n_204_ | new_n_207_;
  assign new_n_209_ = new_n_201_ & new_n_208_;
  assign new_n_214_ = ~A235 | A236;
  assign new_n_215_ = A233 & new_n_214_;
  assign new_n_216_ = A232 & new_n_215_;
  assign new_n_217_ = new_n_209_ | new_n_216_;
  assign new_n_218_ = ~A234 & new_n_217_;
  assign new_n_223_ = ~A235 | A236;
  assign new_n_224_ = ~A233 & new_n_223_;
  assign new_n_225_ = ~A232 & new_n_224_;
  assign new_n_226_ = new_n_218_ | new_n_225_;
  assign new_n_227_ = new_n_197_ & new_n_226_;
  assign new_n_234_ = ~A235 & A236;
  assign new_n_235_ = A233 & new_n_234_;
  assign new_n_239_ = A235 & ~A236;
  assign new_n_240_ = ~A233 & new_n_239_;
  assign new_n_241_ = new_n_235_ | new_n_240_;
  assign new_n_242_ = ~A232 & new_n_241_;
  assign new_n_248_ = A235 & ~A236;
  assign new_n_249_ = A232 & new_n_248_;
  assign new_n_250_ = A234 | new_n_249_;
  assign new_n_251_ = A233 & new_n_250_;
  assign new_n_257_ = ~A235 & A236;
  assign new_n_258_ = ~A233 & new_n_257_;
  assign new_n_259_ = A234 | new_n_258_;
  assign new_n_260_ = A232 & new_n_259_;
  assign new_n_261_ = new_n_251_ | new_n_260_;
  assign new_n_262_ = new_n_242_ | new_n_261_;
  assign new_n_265_ = A301 | ~A302;
  assign new_n_268_ = ~A298 & A299;
  assign new_n_271_ = A298 & ~A299;
  assign new_n_272_ = new_n_268_ | new_n_271_;
  assign new_n_275_ = A268 | ~A269;
  assign new_n_278_ = ~A265 & A266;
  assign new_n_281_ = A265 & ~A266;
  assign new_n_282_ = new_n_278_ | new_n_281_;
  assign new_n_283_ = new_n_275_ & new_n_282_;
  assign new_n_288_ = ~A268 | A269;
  assign new_n_289_ = A266 & new_n_288_;
  assign new_n_290_ = A265 & new_n_289_;
  assign new_n_291_ = new_n_283_ | new_n_290_;
  assign new_n_292_ = new_n_272_ & new_n_291_;
  assign new_n_293_ = new_n_265_ & new_n_292_;
  assign new_n_298_ = ~A301 | A302;
  assign new_n_301_ = A268 | ~A269;
  assign new_n_304_ = ~A265 & A266;
  assign new_n_307_ = A265 & ~A266;
  assign new_n_308_ = new_n_304_ | new_n_307_;
  assign new_n_309_ = new_n_301_ & new_n_308_;
  assign new_n_314_ = ~A268 | A269;
  assign new_n_315_ = A266 & new_n_314_;
  assign new_n_316_ = A265 & new_n_315_;
  assign new_n_317_ = new_n_309_ | new_n_316_;
  assign new_n_318_ = new_n_298_ & new_n_317_;
  assign new_n_319_ = A299 & new_n_318_;
  assign new_n_320_ = A298 & new_n_319_;
  assign new_n_321_ = new_n_293_ | new_n_320_;
  assign new_n_322_ = new_n_262_ & new_n_321_;
  assign new_n_323_ = ~A267 & new_n_322_;
  assign new_n_328_ = ~A268 | A269;
  assign new_n_333_ = ~A235 & A236;
  assign new_n_334_ = A233 & new_n_333_;
  assign new_n_338_ = A235 & ~A236;
  assign new_n_339_ = ~A233 & new_n_338_;
  assign new_n_340_ = new_n_334_ | new_n_339_;
  assign new_n_341_ = ~A232 & new_n_340_;
  assign new_n_347_ = A235 & ~A236;
  assign new_n_348_ = A232 & new_n_347_;
  assign new_n_349_ = A234 | new_n_348_;
  assign new_n_350_ = A233 & new_n_349_;
  assign new_n_356_ = ~A235 & A236;
  assign new_n_357_ = ~A233 & new_n_356_;
  assign new_n_358_ = A234 | new_n_357_;
  assign new_n_359_ = A232 & new_n_358_;
  assign new_n_360_ = new_n_350_ | new_n_359_;
  assign new_n_361_ = new_n_341_ | new_n_360_;
  assign new_n_364_ = A301 | ~A302;
  assign new_n_367_ = ~A298 & A299;
  assign new_n_370_ = A298 & ~A299;
  assign new_n_371_ = new_n_367_ | new_n_370_;
  assign new_n_372_ = new_n_364_ & new_n_371_;
  assign new_n_377_ = ~A301 | A302;
  assign new_n_378_ = A299 & new_n_377_;
  assign new_n_379_ = A298 & new_n_378_;
  assign new_n_380_ = new_n_372_ | new_n_379_;
  assign new_n_381_ = new_n_361_ & new_n_380_;
  assign new_n_382_ = new_n_328_ & new_n_381_;
  assign new_n_383_ = ~A266 & new_n_382_;
  assign new_n_384_ = ~A265 & new_n_383_;
  assign new_n_385_ = new_n_323_ | new_n_384_;
  assign new_n_386_ = ~A300 & new_n_385_;
  assign new_n_391_ = ~A301 | A302;
  assign new_n_397_ = ~A235 & A236;
  assign new_n_398_ = A233 & new_n_397_;
  assign new_n_402_ = A235 & ~A236;
  assign new_n_403_ = ~A233 & new_n_402_;
  assign new_n_404_ = new_n_398_ | new_n_403_;
  assign new_n_405_ = ~A232 & new_n_404_;
  assign new_n_411_ = A235 & ~A236;
  assign new_n_412_ = A232 & new_n_411_;
  assign new_n_413_ = A234 | new_n_412_;
  assign new_n_414_ = A233 & new_n_413_;
  assign new_n_420_ = ~A235 & A236;
  assign new_n_421_ = ~A233 & new_n_420_;
  assign new_n_422_ = A234 | new_n_421_;
  assign new_n_423_ = A232 & new_n_422_;
  assign new_n_424_ = new_n_414_ | new_n_423_;
  assign new_n_425_ = new_n_405_ | new_n_424_;
  assign new_n_428_ = A268 | ~A269;
  assign new_n_431_ = ~A265 & A266;
  assign new_n_434_ = A265 & ~A266;
  assign new_n_435_ = new_n_431_ | new_n_434_;
  assign new_n_436_ = new_n_428_ & new_n_435_;
  assign new_n_441_ = ~A268 | A269;
  assign new_n_442_ = A266 & new_n_441_;
  assign new_n_443_ = A265 & new_n_442_;
  assign new_n_444_ = new_n_436_ | new_n_443_;
  assign new_n_445_ = new_n_425_ & new_n_444_;
  assign new_n_446_ = ~A267 & new_n_445_;
  assign new_n_451_ = ~A268 | A269;
  assign new_n_456_ = ~A235 & A236;
  assign new_n_457_ = A233 & new_n_456_;
  assign new_n_461_ = A235 & ~A236;
  assign new_n_462_ = ~A233 & new_n_461_;
  assign new_n_463_ = new_n_457_ | new_n_462_;
  assign new_n_464_ = ~A232 & new_n_463_;
  assign new_n_470_ = A235 & ~A236;
  assign new_n_471_ = A232 & new_n_470_;
  assign new_n_472_ = A234 | new_n_471_;
  assign new_n_473_ = A233 & new_n_472_;
  assign new_n_479_ = ~A235 & A236;
  assign new_n_480_ = ~A233 & new_n_479_;
  assign new_n_481_ = A234 | new_n_480_;
  assign new_n_482_ = A232 & new_n_481_;
  assign new_n_483_ = new_n_473_ | new_n_482_;
  assign new_n_484_ = new_n_464_ | new_n_483_;
  assign new_n_485_ = new_n_451_ & new_n_484_;
  assign new_n_486_ = ~A266 & new_n_485_;
  assign new_n_487_ = ~A265 & new_n_486_;
  assign new_n_488_ = new_n_446_ | new_n_487_;
  assign new_n_489_ = new_n_391_ & new_n_488_;
  assign new_n_490_ = ~A299 & new_n_489_;
  assign new_n_491_ = ~A298 & new_n_490_;
  assign new_n_492_ = new_n_386_ | new_n_491_;
  assign new_n_493_ = new_n_227_ | new_n_492_;
  assign new_n_494_ = new_n_130_ | new_n_493_;
  assign new_n_495_ = new_n_109_ | new_n_494_;
  assign new_n_496_ = new_n_74_ | new_n_495_;
endmodule


