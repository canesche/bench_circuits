module top ( 
    txwrd3, a, qpr4, txwrd2, b, i1zzz0, txwrd5, c, p1zzz0, txwrd4, xzfs,
    i1zzz2, i2zzz1, p1zzz1, p2zzz0, qpr1, i1zzz1, i2zzz0, p1zzz2, p2zzz1,
    qpr0, i1zzz4, i2zzz3, infin, p1zzz3, p2zzz2, qpr3, txwrd1, vybb1,
    i1zzz3, i2zzz2, p1zzz4, p2zzz3, qpr2, txwrd0, vybb0, comppar, psrw,
    xz323, cbt2, mmerr, ryz, xz324, esrsum, v1zzz7, v2zzz6, xz161, pfin,
    stw_n, v2zzz7, vzzze, xz162, xz320, cbt1, slad0, v1zzz5, v2zzz4, xz163,
    xz321, cbt0, slad1, v1zzz6, v2zzz5, xz322, pybb5, slad2, txwrd14,
    v1zzz3, v2zzz2, xz160_n, pybb4, slad3, txwrd13, v1zzz4, v2zzz3, iclr,
    pybb3, rptwin, txwrd12, v1zzz1, v2zzz0, pybb2, txwrd11, v1zzz2, v2zzz1,
    axz1, inzzze, axz0, pybb8, v1zzz0, inybb8, pybb7, xzfr0, enwin, ofs1,
    pybb6, pzzze, txmess_n, txwrd15, xzfr1, i1zzz6, i2zzz5, inybb6, ofs2,
    p1zzz5, p2zzz4, rxz0, i1zzz5, i2zzz4, inybb7, p1zzz6, p2zzz5, rpten,
    rxz1, i2zzz7, inybb4, p1zzz7, p2zzz6, i1zzz7, i2zzz6, inybb5, p2zzz7,
    inybb2, pybb1, txwrd7, txwrd10, inybb3, pybb0, txwrd6, inybb0, txwrd9,
    inybb1, psync, txwrd8, vfin,
    i1zzz0_p, v1zzz0_p, i1zzz3_p, i2zzz2_p, txwrd8_p, v1zzz2_p, v2zzz1_p,
    i1zzz4_p, i2zzz3_p, stw_f, txwrd9_p, v1zzz1_p, v2zzz0_p, xz163_p, c_p,
    enwin_p, i1zzz1_p, i2zzz0_p, txwrd6_p, v1zzz4_p, v2zzz3_p, i1zzz2_p,
    i2zzz1_p, txwrd7_p, v1zzz3_p, v2zzz2_p, p1zzz4_p, p2zzz3_p, xz162_p,
    b_p, p1zzz3_p, p2zzz2_p, p1zzz2_p, p2zzz1_p, xzfr1_p, p1zzz1_p,
    p2zzz0_p, txwrd14_p, xz161_p, a_p, p1zzz0_p, axz0_p, txwrd15_p, axz1_p,
    td_p, fsesr_p, rptwin_p, txwrd12_p, txwrd11_p, xz322_p, p2zzz7_p,
    txwrd13_p, xz324_p, xzfs_p, p1zzz7_p, p2zzz6_p, xzfr0_p, p1zzz6_p,
    p2zzz5_p, rxz1_p, comppar_p, ofs2_p, p1zzz5_p, p2zzz4_p, rxz0_p,
    xz323_p, i1zzz7_p, i2zzz6_p, ofs1_p, ryz_p, sbuff, txwrd4_p, v1zzz6_p,
    v2zzz5_p, xz160_f, xz320_p, i2zzz7_p, txwrd5_p, v1zzz5_p, v2zzz4_p,
    i1zzz5_p, i2zzz4_p, qpr4_p, txwrd2_p, v2zzz7_p, i1zzz6_p, i2zzz5_p,
    txwrd3_p, v1zzz7_p, v2zzz6_p, qpr2_p, txwrd0_p, qpr3_p, txwrd1_p,
    xz321_p, qpr0_p, qpr1_p, txmess_f, txwrd10_p  );
  input  txwrd3, a, qpr4, txwrd2, b, i1zzz0, txwrd5, c, p1zzz0, txwrd4,
    xzfs, i1zzz2, i2zzz1, p1zzz1, p2zzz0, qpr1, i1zzz1, i2zzz0, p1zzz2,
    p2zzz1, qpr0, i1zzz4, i2zzz3, infin, p1zzz3, p2zzz2, qpr3, txwrd1,
    vybb1, i1zzz3, i2zzz2, p1zzz4, p2zzz3, qpr2, txwrd0, vybb0, comppar,
    psrw, xz323, cbt2, mmerr, ryz, xz324, esrsum, v1zzz7, v2zzz6, xz161,
    pfin, stw_n, v2zzz7, vzzze, xz162, xz320, cbt1, slad0, v1zzz5, v2zzz4,
    xz163, xz321, cbt0, slad1, v1zzz6, v2zzz5, xz322, pybb5, slad2,
    txwrd14, v1zzz3, v2zzz2, xz160_n, pybb4, slad3, txwrd13, v1zzz4,
    v2zzz3, iclr, pybb3, rptwin, txwrd12, v1zzz1, v2zzz0, pybb2, txwrd11,
    v1zzz2, v2zzz1, axz1, inzzze, axz0, pybb8, v1zzz0, inybb8, pybb7,
    xzfr0, enwin, ofs1, pybb6, pzzze, txmess_n, txwrd15, xzfr1, i1zzz6,
    i2zzz5, inybb6, ofs2, p1zzz5, p2zzz4, rxz0, i1zzz5, i2zzz4, inybb7,
    p1zzz6, p2zzz5, rpten, rxz1, i2zzz7, inybb4, p1zzz7, p2zzz6, i1zzz7,
    i2zzz6, inybb5, p2zzz7, inybb2, pybb1, txwrd7, txwrd10, inybb3, pybb0,
    txwrd6, inybb0, txwrd9, inybb1, psync, txwrd8, vfin;
  output i1zzz0_p, v1zzz0_p, i1zzz3_p, i2zzz2_p, txwrd8_p, v1zzz2_p, v2zzz1_p,
    i1zzz4_p, i2zzz3_p, stw_f, txwrd9_p, v1zzz1_p, v2zzz0_p, xz163_p, c_p,
    enwin_p, i1zzz1_p, i2zzz0_p, txwrd6_p, v1zzz4_p, v2zzz3_p, i1zzz2_p,
    i2zzz1_p, txwrd7_p, v1zzz3_p, v2zzz2_p, p1zzz4_p, p2zzz3_p, xz162_p,
    b_p, p1zzz3_p, p2zzz2_p, p1zzz2_p, p2zzz1_p, xzfr1_p, p1zzz1_p,
    p2zzz0_p, txwrd14_p, xz161_p, a_p, p1zzz0_p, axz0_p, txwrd15_p, axz1_p,
    td_p, fsesr_p, rptwin_p, txwrd12_p, txwrd11_p, xz322_p, p2zzz7_p,
    txwrd13_p, xz324_p, xzfs_p, p1zzz7_p, p2zzz6_p, xzfr0_p, p1zzz6_p,
    p2zzz5_p, rxz1_p, comppar_p, ofs2_p, p1zzz5_p, p2zzz4_p, rxz0_p,
    xz323_p, i1zzz7_p, i2zzz6_p, ofs1_p, ryz_p, sbuff, txwrd4_p, v1zzz6_p,
    v2zzz5_p, xz160_f, xz320_p, i2zzz7_p, txwrd5_p, v1zzz5_p, v2zzz4_p,
    i1zzz5_p, i2zzz4_p, qpr4_p, txwrd2_p, v2zzz7_p, i1zzz6_p, i2zzz5_p,
    txwrd3_p, v1zzz7_p, v2zzz6_p, qpr2_p, txwrd0_p, qpr3_p, txwrd1_p,
    xz321_p, qpr0_p, qpr1_p, txmess_f, txwrd10_p;
  wire new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n241_,
    new_n242_, new_n243_, new_n244_, new_n245_, new_n247_, new_n248_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n274_, new_n275_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n283_,
    new_n284_, new_n286_, new_n287_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n310_, new_n311_,
    new_n313_, new_n314_, new_n316_, new_n317_, new_n318_, new_n319_,
    new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n330_, new_n331_, new_n332_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n353_, new_n354_,
    new_n356_, new_n357_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n369_,
    new_n370_, new_n372_, new_n373_, new_n375_, new_n376_, new_n378_,
    new_n379_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n393_, new_n394_, new_n396_, new_n397_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n431_, new_n432_, new_n434_, new_n435_,
    new_n437_, new_n438_, new_n440_, new_n441_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n457_,
    new_n458_, new_n460_, new_n461_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n473_, new_n474_, new_n475_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n486_,
    new_n487_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_,
    new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n547_, new_n548_, new_n549_, new_n552_, new_n553_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n746_, new_n747_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n842_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n878_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_;
  assign new_n235_ = ~inzzze & inybb0;
  assign new_n236_ = ~ryz & new_n235_;
  assign new_n237_ = inybb1 & new_n236_;
  assign new_n238_ = ~ryz & ~new_n235_;
  assign new_n239_ = i1zzz0 & new_n238_;
  assign i1zzz0_p = new_n237_ | new_n239_;
  assign new_n241_ = vybb0 & ~vzzze;
  assign new_n242_ = ~ryz & new_n241_;
  assign new_n243_ = v1zzz1 & new_n242_;
  assign new_n244_ = ~ryz & ~new_n241_;
  assign new_n245_ = v1zzz0 & new_n244_;
  assign v1zzz0_p = new_n243_ | new_n245_;
  assign new_n247_ = inybb4 & new_n236_;
  assign new_n248_ = i1zzz3 & new_n238_;
  assign i1zzz3_p = new_n247_ | new_n248_;
  assign new_n250_ = inzzze & inybb0;
  assign new_n251_ = ~ryz & new_n250_;
  assign new_n252_ = inybb3 & new_n251_;
  assign new_n253_ = ~ryz & ~new_n250_;
  assign new_n254_ = i2zzz2 & new_n253_;
  assign i2zzz2_p = new_n252_ | new_n254_;
  assign new_n256_ = ~infin & ~ryz;
  assign new_n257_ = pfin & new_n256_;
  assign new_n258_ = p2zzz0 & new_n257_;
  assign new_n259_ = ~pfin & new_n256_;
  assign new_n260_ = ~b & ~c;
  assign new_n261_ = ~txmess_n & ~new_n260_;
  assign new_n262_ = ~vfin & ~new_n261_;
  assign new_n263_ = txwrd8 & new_n262_;
  assign new_n264_ = ~vfin & new_n261_;
  assign new_n265_ = txwrd9 & new_n264_;
  assign new_n266_ = v2zzz0 & vfin;
  assign new_n267_ = ~new_n263_ & ~new_n265_;
  assign new_n268_ = ~new_n266_ & new_n267_;
  assign new_n269_ = new_n259_ & ~new_n268_;
  assign new_n270_ = infin & ~ryz;
  assign new_n271_ = i2zzz0 & new_n270_;
  assign new_n272_ = ~new_n258_ & ~new_n269_;
  assign txwrd8_p = new_n271_ | ~new_n272_;
  assign new_n274_ = v1zzz3 & new_n242_;
  assign new_n275_ = v1zzz2 & new_n244_;
  assign v1zzz2_p = new_n274_ | new_n275_;
  assign new_n277_ = vybb0 & vzzze;
  assign new_n278_ = ~ryz & new_n277_;
  assign new_n279_ = v2zzz2 & new_n278_;
  assign new_n280_ = ~ryz & ~new_n277_;
  assign new_n281_ = v2zzz1 & new_n280_;
  assign v2zzz1_p = new_n279_ | new_n281_;
  assign new_n283_ = inybb5 & new_n236_;
  assign new_n284_ = i1zzz4 & new_n238_;
  assign i1zzz4_p = new_n283_ | new_n284_;
  assign new_n286_ = inybb4 & new_n251_;
  assign new_n287_ = i2zzz3 & new_n253_;
  assign i2zzz3_p = new_n286_ | new_n287_;
  assign new_n289_ = ~infin & ~pfin;
  assign new_n290_ = axz1 & axz0;
  assign new_n291_ = ~txmess_n & new_n290_;
  assign new_n292_ = a & new_n291_;
  assign new_n293_ = ~stw_n & ~new_n292_;
  assign new_n294_ = new_n289_ & ~new_n293_;
  assign new_n295_ = ~vfin & new_n294_;
  assign stw_f = ryz | new_n295_;
  assign new_n297_ = ~pfin & vfin;
  assign new_n298_ = v2zzz1 & new_n297_;
  assign new_n299_ = ~pfin & new_n262_;
  assign new_n300_ = txwrd9 & new_n299_;
  assign new_n301_ = ~pfin & new_n264_;
  assign new_n302_ = txwrd10 & new_n301_;
  assign new_n303_ = p2zzz1 & pfin;
  assign new_n304_ = ~new_n298_ & ~new_n300_;
  assign new_n305_ = ~new_n302_ & ~new_n303_;
  assign new_n306_ = new_n304_ & new_n305_;
  assign new_n307_ = new_n256_ & ~new_n306_;
  assign new_n308_ = i2zzz1 & new_n270_;
  assign txwrd9_p = new_n307_ | new_n308_;
  assign new_n310_ = v1zzz2 & new_n242_;
  assign new_n311_ = v1zzz1 & new_n244_;
  assign v1zzz1_p = new_n310_ | new_n311_;
  assign new_n313_ = v2zzz1 & new_n278_;
  assign new_n314_ = v2zzz0 & new_n280_;
  assign v2zzz0_p = new_n313_ | new_n314_;
  assign new_n316_ = ~iclr & ~psync;
  assign new_n317_ = xz321 & xz322;
  assign new_n318_ = xz324 & new_n317_;
  assign new_n319_ = xz323 & new_n318_;
  assign new_n320_ = ~xz160_n & new_n319_;
  assign new_n321_ = xz161 & new_n320_;
  assign new_n322_ = xz320 & new_n321_;
  assign new_n323_ = xz162 & new_n316_;
  assign new_n324_ = ~xz163 & new_n323_;
  assign new_n325_ = new_n322_ & new_n324_;
  assign new_n326_ = xz161 & xz162;
  assign new_n327_ = new_n316_ & ~new_n326_;
  assign new_n328_ = new_n316_ & ~new_n320_;
  assign xz320_p = ~xz320 & new_n316_;
  assign new_n330_ = ~new_n328_ & ~xz320_p;
  assign new_n331_ = ~new_n327_ & new_n330_;
  assign new_n332_ = xz163 & ~new_n331_;
  assign xz163_p = new_n325_ | new_n332_;
  assign new_n334_ = cbt2 & ~cbt1;
  assign new_n335_ = ~cbt0 & new_n334_;
  assign new_n336_ = ~qpr4 & ~new_n335_;
  assign new_n337_ = ~qpr1 & qpr2;
  assign new_n338_ = qpr0 & new_n337_;
  assign new_n339_ = ~qpr3 & ~new_n336_;
  assign new_n340_ = ~txmess_n & new_n338_;
  assign new_n341_ = new_n339_ & new_n340_;
  assign new_n342_ = ~c & new_n341_;
  assign new_n343_ = c & ~new_n341_;
  assign new_n344_ = ~new_n342_ & ~new_n343_;
  assign c_p = ~ryz & ~new_n344_;
  assign ofs1_p = ~iclr & psync;
  assign new_n347_ = xzfs & ofs1_p;
  assign new_n348_ = ~iclr & enwin;
  assign new_n349_ = ~new_n347_ & ~new_n348_;
  assign new_n350_ = ofs1 & ofs2;
  assign new_n351_ = ~new_n349_ & ~new_n350_;
  assign enwin_p = psrw & new_n351_;
  assign new_n353_ = inybb2 & new_n236_;
  assign new_n354_ = i1zzz1 & new_n238_;
  assign i1zzz1_p = new_n353_ | new_n354_;
  assign new_n356_ = inybb1 & new_n251_;
  assign new_n357_ = i2zzz0 & new_n253_;
  assign i2zzz0_p = new_n356_ | new_n357_;
  assign new_n359_ = p1zzz6 & new_n257_;
  assign new_n360_ = txwrd6 & new_n262_;
  assign new_n361_ = txwrd7 & new_n264_;
  assign new_n362_ = v1zzz6 & vfin;
  assign new_n363_ = ~new_n360_ & ~new_n361_;
  assign new_n364_ = ~new_n362_ & new_n363_;
  assign new_n365_ = new_n259_ & ~new_n364_;
  assign new_n366_ = i1zzz6 & new_n270_;
  assign new_n367_ = ~new_n359_ & ~new_n365_;
  assign txwrd6_p = new_n366_ | ~new_n367_;
  assign new_n369_ = v1zzz5 & new_n242_;
  assign new_n370_ = v1zzz4 & new_n244_;
  assign v1zzz4_p = new_n369_ | new_n370_;
  assign new_n372_ = v2zzz4 & new_n278_;
  assign new_n373_ = v2zzz3 & new_n280_;
  assign v2zzz3_p = new_n372_ | new_n373_;
  assign new_n375_ = inybb3 & new_n236_;
  assign new_n376_ = i1zzz2 & new_n238_;
  assign i1zzz2_p = new_n375_ | new_n376_;
  assign new_n378_ = inybb2 & new_n251_;
  assign new_n379_ = i2zzz1 & new_n253_;
  assign i2zzz1_p = new_n378_ | new_n379_;
  assign new_n381_ = infin & i1zzz7;
  assign new_n382_ = ~infin & pfin;
  assign new_n383_ = p1zzz7 & new_n382_;
  assign new_n384_ = txwrd7 & new_n262_;
  assign new_n385_ = txwrd8 & new_n264_;
  assign new_n386_ = v1zzz7 & vfin;
  assign new_n387_ = ~new_n384_ & ~new_n385_;
  assign new_n388_ = ~new_n386_ & new_n387_;
  assign new_n389_ = new_n289_ & ~new_n388_;
  assign new_n390_ = ~new_n381_ & ~new_n383_;
  assign new_n391_ = ~new_n389_ & new_n390_;
  assign txwrd7_p = ~ryz & ~new_n391_;
  assign new_n393_ = v1zzz4 & new_n242_;
  assign new_n394_ = v1zzz3 & new_n244_;
  assign v1zzz3_p = new_n393_ | new_n394_;
  assign new_n396_ = v2zzz3 & new_n278_;
  assign new_n397_ = v2zzz2 & new_n280_;
  assign v2zzz2_p = new_n396_ | new_n397_;
  assign new_n399_ = ~pzzze & pybb0;
  assign new_n400_ = ~ryz & new_n399_;
  assign new_n401_ = pybb5 & new_n400_;
  assign new_n402_ = ~ryz & ~new_n399_;
  assign new_n403_ = p1zzz4 & new_n402_;
  assign p1zzz4_p = new_n401_ | new_n403_;
  assign new_n405_ = pzzze & pybb0;
  assign new_n406_ = ~ryz & new_n405_;
  assign new_n407_ = pybb4 & new_n406_;
  assign new_n408_ = ~ryz & ~new_n405_;
  assign new_n409_ = p2zzz3 & new_n408_;
  assign p2zzz3_p = new_n407_ | new_n409_;
  assign new_n411_ = ~xz162 & new_n316_;
  assign new_n412_ = new_n322_ & new_n411_;
  assign new_n413_ = ~xz161 & new_n316_;
  assign new_n414_ = new_n330_ & ~new_n413_;
  assign new_n415_ = xz162 & ~new_n414_;
  assign xz162_p = new_n412_ | new_n415_;
  assign new_n417_ = ~cbt1 & ~cbt0;
  assign new_n418_ = cbt2 & ~new_n417_;
  assign new_n419_ = ~qpr4 & ~qpr3;
  assign new_n420_ = new_n338_ & new_n419_;
  assign new_n421_ = ~b & new_n420_;
  assign new_n422_ = new_n418_ & new_n421_;
  assign new_n423_ = ~txmess_n & new_n422_;
  assign new_n424_ = ~qpr3 & ~new_n418_;
  assign new_n425_ = new_n338_ & ~new_n424_;
  assign new_n426_ = ~qpr4 & ~txmess_n;
  assign new_n427_ = new_n425_ & new_n426_;
  assign new_n428_ = b & ~new_n427_;
  assign new_n429_ = ~new_n423_ & ~new_n428_;
  assign b_p = ~ryz & ~new_n429_;
  assign new_n431_ = pybb4 & new_n400_;
  assign new_n432_ = p1zzz3 & new_n402_;
  assign p1zzz3_p = new_n431_ | new_n432_;
  assign new_n434_ = pybb3 & new_n406_;
  assign new_n435_ = p2zzz2 & new_n408_;
  assign p2zzz2_p = new_n434_ | new_n435_;
  assign new_n437_ = pybb3 & new_n400_;
  assign new_n438_ = p1zzz2 & new_n402_;
  assign p1zzz2_p = new_n437_ | new_n438_;
  assign new_n440_ = pybb2 & new_n406_;
  assign new_n441_ = p2zzz1 & new_n408_;
  assign p2zzz1_p = new_n440_ | new_n441_;
  assign new_n443_ = ~xz163 & new_n319_;
  assign new_n444_ = ~xz161 & new_n443_;
  assign new_n445_ = ~xz162 & xz160_n;
  assign new_n446_ = new_n444_ & new_n445_;
  assign new_n447_ = xz320 & new_n316_;
  assign new_n448_ = ~xzfr1 & new_n446_;
  assign new_n449_ = new_n447_ & new_n448_;
  assign new_n450_ = xzfr0 & new_n449_;
  assign new_n451_ = ~xzfr0 & new_n316_;
  assign new_n452_ = new_n316_ & ~new_n446_;
  assign new_n453_ = ~xz320_p & ~new_n452_;
  assign new_n454_ = ~new_n451_ & new_n453_;
  assign new_n455_ = xzfr1 & ~new_n454_;
  assign xzfr1_p = new_n450_ | new_n455_;
  assign new_n457_ = pybb2 & new_n400_;
  assign new_n458_ = p1zzz1 & new_n402_;
  assign p1zzz1_p = new_n457_ | new_n458_;
  assign new_n460_ = pybb1 & new_n406_;
  assign new_n461_ = p2zzz0 & new_n408_;
  assign p2zzz0_p = new_n460_ | new_n461_;
  assign new_n463_ = i2zzz6 & new_n270_;
  assign new_n464_ = txwrd14 & new_n262_;
  assign new_n465_ = txwrd15 & new_n264_;
  assign new_n466_ = v2zzz6 & vfin;
  assign new_n467_ = ~new_n464_ & ~new_n465_;
  assign new_n468_ = ~new_n466_ & new_n467_;
  assign new_n469_ = new_n259_ & ~new_n468_;
  assign new_n470_ = p2zzz6 & new_n257_;
  assign new_n471_ = ~new_n463_ & ~new_n469_;
  assign txwrd14_p = new_n470_ | ~new_n471_;
  assign new_n473_ = new_n320_ & new_n447_;
  assign new_n474_ = ~xz161 & new_n473_;
  assign new_n475_ = xz161 & ~new_n330_;
  assign xz161_p = new_n474_ | new_n475_;
  assign new_n477_ = ~qpr4 & b;
  assign new_n478_ = qpr3 & new_n477_;
  assign new_n479_ = ~qpr4 & cbt2;
  assign new_n480_ = ~qpr3 & ~new_n479_;
  assign new_n481_ = ~new_n478_ & ~new_n480_;
  assign new_n482_ = new_n338_ & ~new_n481_;
  assign new_n483_ = ~txmess_n & new_n482_;
  assign new_n484_ = ~a & ~new_n483_;
  assign a_p = ~ryz & ~new_n484_;
  assign new_n486_ = pybb1 & new_n400_;
  assign new_n487_ = p1zzz0 & new_n402_;
  assign p1zzz0_p = new_n486_ | new_n487_;
  assign new_n489_ = ~a & ~new_n482_;
  assign new_n490_ = ~txmess_n & ~new_n489_;
  assign new_n491_ = ~axz0 & new_n490_;
  assign new_n492_ = axz0 & ~new_n490_;
  assign new_n493_ = ~new_n491_ & ~new_n492_;
  assign axz0_p = ~ryz & ~new_n493_;
  assign new_n495_ = txwrd15 & new_n299_;
  assign new_n496_ = v2zzz7 & new_n297_;
  assign new_n497_ = pfin & p2zzz7;
  assign new_n498_ = ~new_n495_ & ~new_n496_;
  assign new_n499_ = ~new_n497_ & new_n498_;
  assign new_n500_ = new_n256_ & ~new_n499_;
  assign new_n501_ = i2zzz7 & new_n270_;
  assign txwrd15_p = new_n500_ | new_n501_;
  assign new_n503_ = ~axz1 & axz0;
  assign new_n504_ = new_n490_ & new_n503_;
  assign new_n505_ = axz0 & new_n490_;
  assign new_n506_ = axz1 & ~new_n505_;
  assign new_n507_ = ~new_n504_ & ~new_n506_;
  assign axz1_p = ~ryz & ~new_n507_;
  assign new_n509_ = rxz0 & ~rxz1;
  assign new_n510_ = ~esrsum & new_n509_;
  assign new_n511_ = ~rxz0 & rxz1;
  assign new_n512_ = esrsum & new_n511_;
  assign new_n513_ = ~new_n510_ & ~new_n512_;
  assign new_n514_ = rpten & ~new_n513_;
  assign new_n515_ = rptwin & new_n514_;
  assign new_n516_ = ~axz1 & ~axz0;
  assign new_n517_ = a & ~new_n516_;
  assign new_n518_ = new_n260_ & ~new_n517_;
  assign new_n519_ = ~rptwin & new_n518_;
  assign sbuff = rptwin | ~txmess_n;
  assign new_n521_ = ~new_n519_ & sbuff;
  assign new_n522_ = ~qpr0 & slad1;
  assign new_n523_ = qpr0 & slad0;
  assign new_n524_ = ~new_n522_ & ~new_n523_;
  assign new_n525_ = qpr2 & ~new_n524_;
  assign new_n526_ = ~qpr1 & new_n525_;
  assign new_n527_ = ~qpr0 & slad3;
  assign new_n528_ = qpr0 & slad2;
  assign new_n529_ = ~new_n527_ & ~new_n528_;
  assign new_n530_ = ~qpr2 & ~new_n529_;
  assign new_n531_ = qpr1 & new_n530_;
  assign new_n532_ = ~new_n526_ & ~new_n531_;
  assign new_n533_ = ~qpr3 & ~new_n521_;
  assign new_n534_ = ~qpr4 & new_n533_;
  assign new_n535_ = ~new_n532_ & new_n534_;
  assign new_n536_ = txwrd0 & ~new_n517_;
  assign new_n537_ = ~new_n260_ & new_n536_;
  assign new_n538_ = ~mmerr & new_n503_;
  assign new_n539_ = ~comppar & axz0;
  assign new_n540_ = esrsum & ~axz0;
  assign new_n541_ = ~new_n539_ & ~new_n540_;
  assign new_n542_ = axz1 & ~new_n541_;
  assign new_n543_ = ~new_n538_ & ~new_n542_;
  assign new_n544_ = a & ~new_n543_;
  assign new_n545_ = ~new_n537_ & ~new_n544_;
  assign new_n546_ = ~txmess_n & ~new_n545_;
  assign new_n547_ = ~rptwin & new_n546_;
  assign new_n548_ = ~new_n515_ & ~new_n535_;
  assign new_n549_ = ~new_n547_ & new_n548_;
  assign td_p = ~ryz & ~new_n549_;
  assign ofs2_p = ~iclr & ofs1;
  assign new_n552_ = ofs2 & ofs2_p;
  assign new_n553_ = ~iclr & xzfr1;
  assign fsesr_p = new_n552_ | new_n553_;
  assign new_n555_ = rxz0 & rxz1;
  assign new_n556_ = rptwin & ~new_n555_;
  assign new_n557_ = xzfs & ~slad3;
  assign new_n558_ = ~slad2 & psync;
  assign new_n559_ = new_n557_ & new_n558_;
  assign new_n560_ = ~slad1 & new_n559_;
  assign new_n561_ = ~slad0 & new_n560_;
  assign new_n562_ = ~xz162 & ~slad2;
  assign new_n563_ = xz162 & slad2;
  assign new_n564_ = ~new_n562_ & ~new_n563_;
  assign new_n565_ = ~xz163 & ~slad3;
  assign new_n566_ = xz163 & slad3;
  assign new_n567_ = ~new_n565_ & ~new_n566_;
  assign new_n568_ = ~new_n564_ & ~new_n567_;
  assign new_n569_ = ~xz161 & ~slad1;
  assign new_n570_ = xz161 & slad1;
  assign new_n571_ = ~new_n569_ & ~new_n570_;
  assign new_n572_ = xz323 & new_n317_;
  assign new_n573_ = xz320 & new_n572_;
  assign new_n574_ = ~slad0 & xz160_n;
  assign new_n575_ = slad0 & ~xz160_n;
  assign new_n576_ = ~new_n574_ & ~new_n575_;
  assign new_n577_ = new_n568_ & ~new_n571_;
  assign new_n578_ = enwin & new_n577_;
  assign new_n579_ = new_n573_ & new_n578_;
  assign new_n580_ = xz324 & new_n579_;
  assign new_n581_ = ~new_n576_ & new_n580_;
  assign new_n582_ = ~new_n556_ & ~new_n561_;
  assign new_n583_ = ~new_n581_ & new_n582_;
  assign rptwin_p = ~ryz & ~new_n583_;
  assign new_n585_ = txwrd12 & new_n262_;
  assign new_n586_ = txwrd13 & new_n264_;
  assign new_n587_ = v2zzz4 & vfin;
  assign new_n588_ = ~new_n585_ & ~new_n586_;
  assign new_n589_ = ~new_n587_ & new_n588_;
  assign new_n590_ = new_n289_ & ~new_n589_;
  assign new_n591_ = infin & i2zzz4;
  assign new_n592_ = p2zzz4 & new_n382_;
  assign new_n593_ = ~new_n590_ & ~new_n591_;
  assign new_n594_ = ~new_n592_ & new_n593_;
  assign txwrd12_p = ~ryz & ~new_n594_;
  assign new_n596_ = txwrd11 & new_n262_;
  assign new_n597_ = txwrd12 & new_n264_;
  assign new_n598_ = v2zzz3 & vfin;
  assign new_n599_ = ~new_n596_ & ~new_n597_;
  assign new_n600_ = ~new_n598_ & new_n599_;
  assign new_n601_ = new_n289_ & ~new_n600_;
  assign new_n602_ = i2zzz3 & infin;
  assign new_n603_ = p2zzz3 & new_n382_;
  assign new_n604_ = ~new_n601_ & ~new_n602_;
  assign new_n605_ = ~new_n603_ & new_n604_;
  assign txwrd11_p = ~ryz & ~new_n605_;
  assign new_n607_ = ~xz322 & new_n447_;
  assign new_n608_ = xz321 & new_n607_;
  assign new_n609_ = ~xz321 & new_n316_;
  assign new_n610_ = ~xz320_p & ~new_n609_;
  assign new_n611_ = xz322 & ~new_n610_;
  assign xz322_p = new_n608_ | new_n611_;
  assign new_n613_ = pybb8 & new_n406_;
  assign new_n614_ = p2zzz7 & new_n408_;
  assign p2zzz7_p = new_n613_ | new_n614_;
  assign new_n616_ = i2zzz5 & new_n270_;
  assign new_n617_ = txwrd13 & new_n262_;
  assign new_n618_ = txwrd14 & new_n264_;
  assign new_n619_ = v2zzz5 & vfin;
  assign new_n620_ = ~new_n617_ & ~new_n618_;
  assign new_n621_ = ~new_n619_ & new_n620_;
  assign new_n622_ = new_n259_ & ~new_n621_;
  assign new_n623_ = p2zzz5 & new_n257_;
  assign new_n624_ = ~new_n616_ & ~new_n622_;
  assign txwrd13_p = new_n623_ | ~new_n624_;
  assign new_n626_ = new_n316_ & new_n573_;
  assign new_n627_ = ~xz324 & new_n626_;
  assign new_n628_ = xz323 & xz322;
  assign new_n629_ = new_n316_ & ~new_n628_;
  assign new_n630_ = new_n610_ & ~new_n629_;
  assign new_n631_ = xz324 & ~new_n630_;
  assign xz324_p = new_n627_ | new_n631_;
  assign new_n633_ = xzfs & ~iclr;
  assign new_n634_ = ~ofs1_p & ~new_n633_;
  assign new_n635_ = ~new_n350_ & ~new_n634_;
  assign xzfs_p = psrw & new_n635_;
  assign new_n637_ = pybb8 & new_n400_;
  assign new_n638_ = p1zzz7 & new_n402_;
  assign p1zzz7_p = new_n637_ | new_n638_;
  assign new_n640_ = pybb7 & new_n406_;
  assign new_n641_ = p2zzz6 & new_n408_;
  assign p2zzz6_p = new_n640_ | new_n641_;
  assign new_n643_ = new_n446_ & new_n447_;
  assign new_n644_ = ~xzfr0 & new_n643_;
  assign new_n645_ = xzfr0 & ~new_n453_;
  assign xzfr0_p = new_n644_ | new_n645_;
  assign new_n647_ = pybb7 & new_n400_;
  assign new_n648_ = p1zzz6 & new_n402_;
  assign p1zzz6_p = new_n647_ | new_n648_;
  assign new_n650_ = pybb6 & new_n406_;
  assign new_n651_ = p2zzz5 & new_n408_;
  assign p2zzz5_p = new_n650_ | new_n651_;
  assign new_n653_ = ~slad1 & ~slad2;
  assign new_n654_ = xzfs & new_n653_;
  assign new_n655_ = ~slad0 & new_n654_;
  assign new_n656_ = ofs1_p & new_n655_;
  assign new_n657_ = ~slad3 & new_n656_;
  assign new_n658_ = ~rptwin & ~new_n581_;
  assign new_n659_ = ~iclr & ~new_n658_;
  assign new_n660_ = ~new_n657_ & ~new_n659_;
  assign new_n661_ = ~rxz1 & ~new_n660_;
  assign new_n662_ = rxz0 & new_n661_;
  assign new_n663_ = ~iclr & ~rxz0;
  assign new_n664_ = xz162 & ~slad2;
  assign new_n665_ = xz163 & ~slad3;
  assign new_n666_ = ~new_n664_ & ~new_n665_;
  assign new_n667_ = ~psync & ~new_n666_;
  assign new_n668_ = xz161 & ~slad1;
  assign new_n669_ = enwin & ~new_n668_;
  assign new_n670_ = ~slad0 & ~xz160_n;
  assign new_n671_ = new_n319_ & ~new_n670_;
  assign new_n672_ = new_n669_ & new_n671_;
  assign new_n673_ = ~new_n559_ & ~new_n672_;
  assign new_n674_ = xz320 & new_n666_;
  assign new_n675_ = enwin & new_n674_;
  assign new_n676_ = xz161 & new_n671_;
  assign new_n677_ = new_n675_ & new_n676_;
  assign new_n678_ = slad1 & ~new_n677_;
  assign new_n679_ = xz320 & ~new_n664_;
  assign new_n680_ = xz163 & new_n679_;
  assign new_n681_ = slad3 & ~new_n680_;
  assign new_n682_ = xz320 & ~new_n665_;
  assign new_n683_ = xz162 & new_n682_;
  assign new_n684_ = slad2 & ~new_n683_;
  assign new_n685_ = new_n669_ & new_n674_;
  assign new_n686_ = new_n320_ & new_n685_;
  assign new_n687_ = slad0 & ~new_n686_;
  assign new_n688_ = ~xzfs & ~new_n674_;
  assign new_n689_ = ~new_n667_ & ~new_n673_;
  assign new_n690_ = ~new_n678_ & ~new_n681_;
  assign new_n691_ = new_n689_ & new_n690_;
  assign new_n692_ = ~new_n684_ & ~new_n687_;
  assign new_n693_ = ~new_n688_ & new_n692_;
  assign new_n694_ = new_n691_ & new_n693_;
  assign new_n695_ = ~iclr & ~new_n694_;
  assign new_n696_ = ~xz320_p & ~new_n695_;
  assign new_n697_ = ~rptwin & ~new_n696_;
  assign new_n698_ = ~new_n663_ & ~new_n697_;
  assign new_n699_ = rxz1 & ~new_n698_;
  assign rxz1_p = new_n662_ | new_n699_;
  assign new_n701_ = ~qpr3 & ~new_n532_;
  assign new_n702_ = ~qpr4 & new_n701_;
  assign new_n703_ = new_n260_ & new_n702_;
  assign new_n704_ = txwrd0 & ~new_n260_;
  assign new_n705_ = ~new_n703_ & ~new_n704_;
  assign new_n706_ = ~new_n517_ & new_n705_;
  assign new_n707_ = ~txmess_n & ~new_n706_;
  assign new_n708_ = comppar & ~new_n707_;
  assign new_n709_ = ~comppar & ~new_n517_;
  assign new_n710_ = ~txmess_n & new_n709_;
  assign new_n711_ = ~new_n705_ & new_n710_;
  assign new_n712_ = ~esrsum & axz1;
  assign new_n713_ = mmerr & axz0;
  assign new_n714_ = ~new_n712_ & ~new_n713_;
  assign new_n715_ = comppar & ~new_n714_;
  assign new_n716_ = esrsum & axz1;
  assign new_n717_ = ~mmerr & axz0;
  assign new_n718_ = ~new_n716_ & ~new_n717_;
  assign new_n719_ = ~comppar & ~txmess_n;
  assign new_n720_ = ~new_n718_ & new_n719_;
  assign new_n721_ = ~new_n715_ & ~new_n720_;
  assign new_n722_ = ~new_n291_ & new_n721_;
  assign new_n723_ = a & ~new_n722_;
  assign new_n724_ = ~new_n708_ & ~new_n711_;
  assign new_n725_ = ~new_n723_ & new_n724_;
  assign comppar_p = ~ryz & ~new_n725_;
  assign new_n727_ = pybb6 & new_n400_;
  assign new_n728_ = p1zzz5 & new_n402_;
  assign p1zzz5_p = new_n727_ | new_n728_;
  assign new_n730_ = pybb5 & new_n406_;
  assign new_n731_ = p2zzz4 & new_n408_;
  assign p2zzz4_p = new_n730_ | new_n731_;
  assign new_n733_ = rxz0 & ~new_n696_;
  assign new_n734_ = ~rptwin & new_n733_;
  assign new_n735_ = ~rxz0 & ~new_n660_;
  assign rxz0_p = new_n734_ | new_n735_;
  assign new_n737_ = new_n317_ & new_n447_;
  assign new_n738_ = ~xz323 & new_n737_;
  assign new_n739_ = ~xz322 & new_n316_;
  assign new_n740_ = new_n610_ & ~new_n739_;
  assign new_n741_ = xz323 & ~new_n740_;
  assign xz323_p = new_n738_ | new_n741_;
  assign new_n743_ = inybb8 & new_n236_;
  assign new_n744_ = i1zzz7 & new_n238_;
  assign i1zzz7_p = new_n743_ | new_n744_;
  assign new_n746_ = inybb7 & new_n251_;
  assign new_n747_ = i2zzz6 & new_n253_;
  assign i2zzz6_p = new_n746_ | new_n747_;
  assign ryz_p = iclr | new_n292_;
  assign new_n750_ = p1zzz4 & new_n257_;
  assign new_n751_ = txwrd4 & new_n262_;
  assign new_n752_ = txwrd5 & new_n264_;
  assign new_n753_ = v1zzz4 & vfin;
  assign new_n754_ = ~new_n751_ & ~new_n752_;
  assign new_n755_ = ~new_n753_ & new_n754_;
  assign new_n756_ = new_n259_ & ~new_n755_;
  assign new_n757_ = i1zzz4 & new_n270_;
  assign new_n758_ = ~new_n750_ & ~new_n756_;
  assign txwrd4_p = new_n757_ | ~new_n758_;
  assign new_n760_ = v1zzz7 & new_n242_;
  assign new_n761_ = v1zzz6 & new_n244_;
  assign v1zzz6_p = new_n760_ | new_n761_;
  assign new_n763_ = v2zzz6 & new_n278_;
  assign new_n764_ = v2zzz5 & new_n280_;
  assign v2zzz5_p = new_n763_ | new_n764_;
  assign new_n766_ = new_n316_ & ~new_n319_;
  assign new_n767_ = ~xz320_p & ~new_n766_;
  assign new_n768_ = xz160_n & ~new_n767_;
  assign xz160_f = new_n473_ | new_n768_;
  assign new_n770_ = inybb8 & new_n251_;
  assign new_n771_ = i2zzz7 & new_n253_;
  assign i2zzz7_p = new_n770_ | new_n771_;
  assign new_n773_ = p1zzz5 & new_n257_;
  assign new_n774_ = txwrd5 & new_n262_;
  assign new_n775_ = txwrd6 & new_n264_;
  assign new_n776_ = v1zzz5 & vfin;
  assign new_n777_ = ~new_n774_ & ~new_n775_;
  assign new_n778_ = ~new_n776_ & new_n777_;
  assign new_n779_ = new_n259_ & ~new_n778_;
  assign new_n780_ = i1zzz5 & new_n270_;
  assign new_n781_ = ~new_n773_ & ~new_n779_;
  assign txwrd5_p = new_n780_ | ~new_n781_;
  assign new_n783_ = v1zzz6 & new_n242_;
  assign new_n784_ = v1zzz5 & new_n244_;
  assign v1zzz5_p = new_n783_ | new_n784_;
  assign new_n786_ = v2zzz5 & new_n278_;
  assign new_n787_ = v2zzz4 & new_n280_;
  assign v2zzz4_p = new_n786_ | new_n787_;
  assign new_n789_ = inybb6 & new_n236_;
  assign new_n790_ = i1zzz5 & new_n238_;
  assign i1zzz5_p = new_n789_ | new_n790_;
  assign new_n792_ = inybb5 & new_n251_;
  assign new_n793_ = i2zzz4 & new_n253_;
  assign i2zzz4_p = new_n792_ | new_n793_;
  assign new_n795_ = ~vfin & new_n289_;
  assign new_n796_ = txmess_n & new_n795_;
  assign txmess_f = ryz | new_n796_;
  assign new_n798_ = qpr0 & ~txmess_f;
  assign new_n799_ = qpr1 & new_n798_;
  assign new_n800_ = qpr3 & new_n799_;
  assign new_n801_ = ~qpr4 & new_n800_;
  assign new_n802_ = qpr2 & new_n801_;
  assign new_n803_ = qpr0 & ~new_n796_;
  assign new_n804_ = qpr1 & new_n803_;
  assign new_n805_ = qpr2 & new_n804_;
  assign new_n806_ = qpr3 & new_n805_;
  assign new_n807_ = qpr4 & ~ryz;
  assign new_n808_ = ~new_n806_ & new_n807_;
  assign qpr4_p = new_n802_ | new_n808_;
  assign new_n810_ = i1zzz2 & new_n270_;
  assign new_n811_ = v1zzz2 & new_n297_;
  assign new_n812_ = txwrd2 & new_n299_;
  assign new_n813_ = txwrd3 & new_n301_;
  assign new_n814_ = p1zzz2 & pfin;
  assign new_n815_ = ~new_n811_ & ~new_n812_;
  assign new_n816_ = ~new_n813_ & ~new_n814_;
  assign new_n817_ = new_n815_ & new_n816_;
  assign new_n818_ = new_n256_ & ~new_n817_;
  assign txwrd2_p = new_n810_ | new_n818_;
  assign new_n820_ = vybb1 & new_n278_;
  assign new_n821_ = v2zzz7 & new_n280_;
  assign v2zzz7_p = new_n820_ | new_n821_;
  assign new_n823_ = inybb7 & new_n236_;
  assign new_n824_ = i1zzz6 & new_n238_;
  assign i1zzz6_p = new_n823_ | new_n824_;
  assign new_n826_ = inybb6 & new_n251_;
  assign new_n827_ = i2zzz5 & new_n253_;
  assign i2zzz5_p = new_n826_ | new_n827_;
  assign new_n829_ = p1zzz3 & new_n257_;
  assign new_n830_ = txwrd3 & new_n262_;
  assign new_n831_ = txwrd4 & new_n264_;
  assign new_n832_ = v1zzz3 & vfin;
  assign new_n833_ = ~new_n830_ & ~new_n831_;
  assign new_n834_ = ~new_n832_ & new_n833_;
  assign new_n835_ = new_n259_ & ~new_n834_;
  assign new_n836_ = i1zzz3 & new_n270_;
  assign new_n837_ = ~new_n829_ & ~new_n835_;
  assign txwrd3_p = new_n836_ | ~new_n837_;
  assign new_n839_ = vybb1 & new_n242_;
  assign new_n840_ = v1zzz7 & new_n244_;
  assign v1zzz7_p = new_n839_ | new_n840_;
  assign new_n842_ = v2zzz7 & new_n278_;
  assign new_n843_ = v2zzz6 & new_n280_;
  assign v2zzz6_p = new_n842_ | new_n843_;
  assign new_n845_ = ~ryz & ~new_n804_;
  assign new_n846_ = qpr2 & new_n845_;
  assign new_n847_ = ~qpr2 & new_n799_;
  assign qpr2_p = new_n846_ | new_n847_;
  assign new_n849_ = txwrd0 & new_n262_;
  assign new_n850_ = txwrd1 & new_n264_;
  assign new_n851_ = v1zzz0 & vfin;
  assign new_n852_ = ~new_n849_ & ~new_n850_;
  assign new_n853_ = ~new_n851_ & new_n852_;
  assign new_n854_ = new_n289_ & ~new_n853_;
  assign new_n855_ = p1zzz0 & new_n382_;
  assign new_n856_ = i1zzz0 & infin;
  assign new_n857_ = ~new_n854_ & ~new_n855_;
  assign new_n858_ = ~new_n856_ & new_n857_;
  assign txwrd0_p = ~ryz & ~new_n858_;
  assign new_n860_ = ~ryz & ~new_n805_;
  assign new_n861_ = qpr3 & new_n860_;
  assign new_n862_ = ~qpr3 & new_n799_;
  assign new_n863_ = qpr2 & new_n862_;
  assign qpr3_p = new_n861_ | new_n863_;
  assign new_n865_ = v1zzz1 & new_n297_;
  assign new_n866_ = txwrd1 & new_n299_;
  assign new_n867_ = txwrd2 & new_n301_;
  assign new_n868_ = p1zzz1 & pfin;
  assign new_n869_ = ~new_n865_ & ~new_n866_;
  assign new_n870_ = ~new_n867_ & ~new_n868_;
  assign new_n871_ = new_n869_ & new_n870_;
  assign new_n872_ = new_n256_ & ~new_n871_;
  assign new_n873_ = i1zzz1 & new_n270_;
  assign txwrd1_p = new_n872_ | new_n873_;
  assign new_n875_ = xz321 & xz320_p;
  assign new_n876_ = ~xz321 & new_n447_;
  assign xz321_p = new_n875_ | new_n876_;
  assign new_n878_ = qpr0 & new_n796_;
  assign new_n879_ = ~ryz & new_n878_;
  assign new_n880_ = ~qpr0 & ~txmess_f;
  assign qpr0_p = new_n879_ | new_n880_;
  assign new_n882_ = ~ryz & ~new_n803_;
  assign new_n883_ = qpr1 & new_n882_;
  assign new_n884_ = ~qpr1 & ~txmess_f;
  assign new_n885_ = qpr0 & new_n884_;
  assign qpr1_p = new_n883_ | new_n885_;
  assign new_n887_ = txwrd10 & new_n262_;
  assign new_n888_ = txwrd11 & new_n264_;
  assign new_n889_ = v2zzz2 & vfin;
  assign new_n890_ = ~new_n887_ & ~new_n888_;
  assign new_n891_ = ~new_n889_ & new_n890_;
  assign new_n892_ = new_n289_ & ~new_n891_;
  assign new_n893_ = infin & i2zzz2;
  assign new_n894_ = p2zzz2 & new_n382_;
  assign new_n895_ = ~new_n892_ & ~new_n893_;
  assign new_n896_ = ~new_n894_ & new_n895_;
  assign txwrd10_p = ~ryz & ~new_n896_;
endmodule

