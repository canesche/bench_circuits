module lal ( 
    a, b, c, d, e, f, g, h, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x, y,
    z, a0,
    b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0,
    t0  );
  input  a, b, c, d, e, f, g, h, j, k, l, m, n, o, p, q, r, s, t, u, v,
    w, x, y, z, a0;
  output b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0,
    s0, t0;
  wire new_n47_, new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_,
    new_n54_, new_n55_, new_n56_, new_n57_, new_n59_, new_n60_, new_n61_,
    new_n62_, new_n63_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_,
    new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_,
    new_n77_, new_n78_, new_n79_, new_n84_, new_n85_, new_n87_, new_n88_,
    new_n90_, new_n91_, new_n92_, new_n94_, new_n95_, new_n96_, new_n97_,
    new_n98_, new_n99_, new_n101_, new_n102_, new_n103_, new_n104_,
    new_n105_, new_n106_, new_n107_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_, new_n114_, new_n115_, new_n116_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_,
    new_n152_, new_n153_;
  assign b0 = j & ~r;
  assign new_n47_ = ~t & ~u;
  assign new_n48_ = ~s & new_n47_;
  assign new_n49_ = ~v & ~new_n48_;
  assign new_n50_ = w & x;
  assign new_n51_ = ~new_n49_ & new_n50_;
  assign new_n52_ = ~z & ~a0;
  assign new_n53_ = e & f;
  assign new_n54_ = ~new_n52_ & ~new_n53_;
  assign new_n55_ = ~h & new_n54_;
  assign new_n56_ = ~y & ~new_n51_;
  assign new_n57_ = ~a0 & new_n56_;
  assign c0 = ~new_n55_ | new_n57_;
  assign new_n59_ = x & z;
  assign new_n60_ = y & z;
  assign new_n61_ = ~a0 & ~new_n60_;
  assign new_n62_ = ~new_n49_ & new_n59_;
  assign new_n63_ = w & new_n62_;
  assign e0 = new_n61_ & ~new_n63_;
  assign new_n65_ = ~b & l;
  assign new_n66_ = ~c & m;
  assign new_n67_ = ~new_n65_ & ~new_n66_;
  assign new_n68_ = ~d & n;
  assign new_n69_ = new_n67_ & ~new_n68_;
  assign new_n70_ = ~a & k;
  assign new_n71_ = new_n69_ & ~new_n70_;
  assign new_n72_ = c & ~m;
  assign new_n73_ = d & ~n;
  assign new_n74_ = ~new_n72_ & ~new_n73_;
  assign new_n75_ = new_n71_ & new_n74_;
  assign new_n76_ = a & ~k;
  assign new_n77_ = b & ~l;
  assign new_n78_ = ~new_n76_ & ~new_n77_;
  assign new_n79_ = new_n75_ & new_n78_;
  assign f0 = ~j & ~new_n79_;
  assign g0 = ~j & ~o;
  assign h0 = ~j & p;
  assign i0 = ~g | j;
  assign new_n84_ = f & ~h;
  assign new_n85_ = e & new_n84_;
  assign k0 = ~q & new_n85_;
  assign new_n87_ = ~h & ~new_n53_;
  assign new_n88_ = ~q & new_n87_;
  assign l0 = ~s & new_n88_;
  assign new_n90_ = ~s & t;
  assign new_n91_ = s & ~t;
  assign new_n92_ = ~new_n90_ & ~new_n91_;
  assign m0 = new_n88_ & ~new_n92_;
  assign new_n94_ = ~q & ~new_n53_;
  assign new_n95_ = ~h & new_n94_;
  assign new_n96_ = s & t;
  assign new_n97_ = u & new_n96_;
  assign new_n98_ = new_n95_ & ~new_n97_;
  assign new_n99_ = ~u & ~new_n96_;
  assign n0 = new_n98_ & ~new_n99_;
  assign new_n101_ = t & u;
  assign new_n102_ = s & new_n101_;
  assign new_n103_ = ~v & new_n102_;
  assign new_n104_ = ~new_n53_ & ~new_n103_;
  assign new_n105_ = ~q & new_n104_;
  assign new_n106_ = v & ~new_n102_;
  assign new_n107_ = ~h & ~new_n106_;
  assign o0 = ~new_n105_ | ~new_n107_;
  assign new_n109_ = u & ~v;
  assign new_n110_ = new_n96_ & new_n109_;
  assign new_n111_ = ~v & ~w;
  assign new_n112_ = new_n102_ & new_n111_;
  assign new_n113_ = ~new_n53_ & ~new_n112_;
  assign new_n114_ = ~q & new_n113_;
  assign new_n115_ = w & ~new_n110_;
  assign new_n116_ = ~h & ~new_n115_;
  assign p0 = ~new_n114_ | ~new_n116_;
  assign new_n118_ = u & new_n111_;
  assign new_n119_ = new_n96_ & new_n118_;
  assign new_n120_ = ~w & ~x;
  assign new_n121_ = new_n110_ & new_n120_;
  assign new_n122_ = ~new_n53_ & ~new_n121_;
  assign new_n123_ = ~q & new_n122_;
  assign new_n124_ = x & ~new_n119_;
  assign new_n125_ = ~h & ~new_n124_;
  assign q0 = ~new_n123_ | ~new_n125_;
  assign new_n127_ = ~v & new_n120_;
  assign new_n128_ = new_n102_ & new_n127_;
  assign new_n129_ = ~x & ~y;
  assign new_n130_ = new_n119_ & new_n129_;
  assign new_n131_ = ~new_n53_ & ~new_n130_;
  assign new_n132_ = ~q & new_n131_;
  assign new_n133_ = y & ~new_n128_;
  assign new_n134_ = ~h & ~new_n133_;
  assign r0 = ~new_n132_ | ~new_n134_;
  assign new_n136_ = t & new_n109_;
  assign new_n137_ = ~w & new_n129_;
  assign new_n138_ = s & new_n136_;
  assign new_n139_ = new_n137_ & new_n138_;
  assign new_n140_ = ~y & ~z;
  assign new_n141_ = new_n128_ & new_n140_;
  assign new_n142_ = ~new_n53_ & ~new_n141_;
  assign new_n143_ = ~q & new_n142_;
  assign new_n144_ = z & ~new_n139_;
  assign new_n145_ = ~h & ~new_n144_;
  assign s0 = ~new_n143_ | ~new_n145_;
  assign new_n147_ = ~x & new_n140_;
  assign new_n148_ = new_n119_ & new_n147_;
  assign new_n149_ = new_n52_ & new_n139_;
  assign new_n150_ = ~new_n53_ & ~new_n149_;
  assign new_n151_ = ~q & new_n150_;
  assign new_n152_ = a0 & ~new_n148_;
  assign new_n153_ = ~h & ~new_n152_;
  assign t0 = ~new_n151_ | ~new_n153_;
  assign j0 = ~e0;
  assign d0 = r;
endmodule

