module top ( 
    pa, pb, pc, pd, pe, pf, pg, ph, pi,
    pp, pa0, pq, pb0, pr, ps, pt, pu, pv, pw, px, py, pz, pj, pk, pl, pm,
    pn, po  );
  input  pa, pb, pc, pd, pe, pf, pg, ph, pi;
  output pp, pa0, pq, pb0, pr, ps, pt, pu, pv, pw, px, py, pz, pj, pk, pl, pm,
    pn, po;
  wire new_n29_, new_n30_, new_n31_, new_n32_, new_n34_, new_n35_, new_n37_,
    new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_,
    new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n55_, new_n56_, new_n58_, new_n59_, new_n60_,
    new_n61_, new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_,
    new_n68_, new_n69_, new_n70_, new_n71_, new_n72_, new_n74_, new_n76_,
    new_n78_, new_n79_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n95_, new_n96_, new_n98_, new_n99_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n111_, new_n112_, new_n113_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n127_, new_n128_, new_n129_,
    new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n136_,
    new_n137_, new_n138_;
  assign new_n29_ = ~pa & pc;
  assign new_n30_ = ~pb & new_n29_;
  assign new_n31_ = pi & new_n30_;
  assign new_n32_ = ~pi & new_n30_;
  assign pp = new_n31_ | new_n32_;
  assign new_n34_ = pa & pc;
  assign new_n35_ = ~pb & new_n34_;
  assign pu = pi & new_n35_;
  assign new_n37_ = ~pb & ~pc;
  assign new_n38_ = ~pe & new_n37_;
  assign new_n39_ = ~pd & new_n38_;
  assign new_n40_ = pf & new_n39_;
  assign new_n41_ = ~pa & new_n40_;
  assign new_n42_ = ~pa & ~pb;
  assign new_n43_ = ~pd & new_n42_;
  assign new_n44_ = ~pc & new_n43_;
  assign new_n45_ = pe & new_n44_;
  assign new_n46_ = ~pc & ~pd;
  assign new_n47_ = ~pf & new_n46_;
  assign new_n48_ = ~pe & new_n47_;
  assign new_n49_ = pg & new_n48_;
  assign new_n50_ = ~pb & new_n49_;
  assign new_n51_ = ~pa & new_n50_;
  assign new_n52_ = ~pu & ~new_n41_;
  assign new_n53_ = ~new_n45_ & ~new_n51_;
  assign pa0 = ~new_n52_ | ~new_n53_;
  assign new_n55_ = ~pa & ~pc;
  assign new_n56_ = ~pb & new_n55_;
  assign pb0 = pd & new_n56_;
  assign new_n58_ = ~pd & ~pe;
  assign new_n59_ = ~pg & new_n58_;
  assign new_n60_ = ~pf & new_n59_;
  assign new_n61_ = ph & new_n60_;
  assign new_n62_ = ~pa & new_n61_;
  assign new_n63_ = ~pc & new_n62_;
  assign new_n64_ = ~pb & new_n63_;
  assign new_n65_ = ~ph & new_n60_;
  assign new_n66_ = ~pa & new_n65_;
  assign new_n67_ = ~pc & new_n66_;
  assign new_n68_ = ~pb & new_n67_;
  assign new_n69_ = ~new_n64_ & ~new_n68_;
  assign new_n70_ = ~new_n41_ & new_n69_;
  assign new_n71_ = ~new_n45_ & ~pb0;
  assign new_n72_ = ~new_n51_ & new_n71_;
  assign pq = ~new_n70_ | ~new_n72_;
  assign new_n74_ = pb & new_n55_;
  assign pr = pi & new_n74_;
  assign new_n76_ = pb & new_n29_;
  assign ps = pi & new_n76_;
  assign new_n78_ = pa & ~pc;
  assign new_n79_ = ~pb & new_n78_;
  assign pt = pi & new_n79_;
  assign new_n81_ = ~pi & new_n35_;
  assign new_n82_ = ~ps & ~pt;
  assign new_n83_ = ~pu & ~new_n81_;
  assign new_n84_ = new_n82_ & new_n83_;
  assign new_n85_ = ~new_n41_ & ~new_n64_;
  assign new_n86_ = ~new_n45_ & ~pr;
  assign new_n87_ = ~new_n51_ & new_n86_;
  assign new_n88_ = new_n85_ & new_n87_;
  assign pv = ~new_n84_ | ~new_n88_;
  assign new_n90_ = ~pu & ~new_n64_;
  assign new_n91_ = new_n82_ & new_n90_;
  assign new_n92_ = ~new_n41_ & ~new_n51_;
  assign new_n93_ = new_n86_ & new_n92_;
  assign pw = ~new_n91_ | ~new_n93_;
  assign new_n95_ = ~new_n45_ & ~pt;
  assign new_n96_ = ~new_n51_ & ~pr;
  assign py = ~new_n95_ | ~new_n96_;
  assign new_n98_ = ~pu & ~new_n45_;
  assign new_n99_ = ~new_n64_ & ~pr;
  assign pz = ~new_n98_ | ~new_n99_;
  assign new_n101_ = pb & new_n78_;
  assign new_n102_ = pi & new_n101_;
  assign new_n103_ = ~pi & new_n101_;
  assign new_n104_ = ~pi & new_n79_;
  assign new_n105_ = ~new_n31_ & ~new_n64_;
  assign new_n106_ = ~new_n102_ & new_n105_;
  assign new_n107_ = ~pr & ~ps;
  assign new_n108_ = ~new_n51_ & new_n107_;
  assign new_n109_ = new_n106_ & new_n108_;
  assign pn = pt | new_n104_;
  assign new_n111_ = ~new_n81_ & ~new_n103_;
  assign new_n112_ = ~pu & new_n111_;
  assign new_n113_ = ~pn & new_n112_;
  assign pj = ~new_n109_ | ~new_n113_;
  assign new_n115_ = ~pi & new_n74_;
  assign new_n116_ = ~pi & new_n76_;
  assign new_n117_ = ~new_n31_ & ~new_n41_;
  assign new_n118_ = ~new_n102_ & new_n117_;
  assign new_n119_ = ~pr & ~new_n115_;
  assign new_n120_ = ~new_n45_ & new_n119_;
  assign new_n121_ = new_n118_ & new_n120_;
  assign new_n122_ = ~ps & ~new_n116_;
  assign new_n123_ = ~pt & ~new_n103_;
  assign new_n124_ = ~pu & new_n123_;
  assign new_n125_ = new_n122_ & new_n124_;
  assign pk = ~new_n121_ | ~new_n125_;
  assign new_n127_ = ~pb0 & ~new_n64_;
  assign new_n128_ = ~new_n102_ & new_n127_;
  assign new_n129_ = ~pp & ~new_n41_;
  assign new_n130_ = new_n128_ & new_n129_;
  assign new_n131_ = ~pr & ~new_n116_;
  assign new_n132_ = ~ps & ~new_n81_;
  assign new_n133_ = ~pt & new_n132_;
  assign new_n134_ = new_n131_ & new_n133_;
  assign pl = ~new_n130_ | ~new_n134_;
  assign new_n136_ = ~new_n115_ & ~new_n116_;
  assign new_n137_ = ~pu & new_n136_;
  assign new_n138_ = ~pr & new_n132_;
  assign pm = ~new_n137_ | ~new_n138_;
  assign po = new_n102_ | new_n103_;
  assign px = pw;
endmodule

