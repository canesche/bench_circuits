module top ( 
    i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, i_13_, i_4_,
    i_12_, i_1_, i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_, i_21_,
    i_16_, i_22_, i_15_, i_19_,
    o_1_, o_2_, o_0_, o_7_, o_5_, o_6_, o_3_, o_4_  );
  input  i_20_, i_9_, i_10_, i_7_, i_8_, i_5_, i_6_, i_14_, i_3_, i_13_,
    i_4_, i_12_, i_1_, i_11_, i_2_, i_23_, i_18_, i_24_, i_17_, i_0_,
    i_21_, i_16_, i_22_, i_15_, i_19_;
  output o_1_, o_2_, o_0_, o_7_, o_5_, o_6_, o_3_, o_4_;
  wire new_n34_, new_n35_, new_n36_, new_n37_, new_n38_, new_n39_, new_n40_,
    new_n41_, new_n42_, new_n43_, new_n44_, new_n45_, new_n46_, new_n47_,
    new_n48_, new_n49_, new_n50_, new_n51_, new_n52_, new_n53_, new_n54_,
    new_n55_, new_n56_, new_n57_, new_n58_, new_n59_, new_n60_, new_n61_,
    new_n62_, new_n63_, new_n64_, new_n65_, new_n66_, new_n67_, new_n68_,
    new_n69_, new_n70_, new_n71_, new_n72_, new_n73_, new_n74_, new_n75_,
    new_n76_, new_n77_, new_n78_, new_n79_, new_n80_, new_n81_, new_n82_,
    new_n83_, new_n84_, new_n85_, new_n86_, new_n87_, new_n88_, new_n89_,
    new_n90_, new_n91_, new_n92_, new_n93_, new_n94_, new_n95_, new_n96_,
    new_n97_, new_n98_, new_n99_, new_n100_, new_n101_, new_n102_,
    new_n103_, new_n104_, new_n105_, new_n106_, new_n107_, new_n108_,
    new_n109_, new_n110_, new_n111_, new_n112_, new_n113_, new_n114_,
    new_n115_, new_n116_, new_n117_, new_n118_, new_n119_, new_n120_,
    new_n121_, new_n122_, new_n123_, new_n124_, new_n125_, new_n126_,
    new_n127_, new_n128_, new_n129_, new_n130_, new_n131_, new_n132_,
    new_n133_, new_n134_, new_n135_, new_n136_, new_n137_, new_n138_,
    new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_,
    new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_,
    new_n151_, new_n152_, new_n153_, new_n154_, new_n156_, new_n157_,
    new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_,
    new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_,
    new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_,
    new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_,
    new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_,
    new_n188_, new_n189_, new_n190_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_;
  assign new_n34_ = i_20_ & i_22_;
  assign new_n35_ = i_18_ & new_n34_;
  assign new_n36_ = i_23_ & i_24_;
  assign new_n37_ = i_17_ & i_16_;
  assign new_n38_ = i_14_ & new_n37_;
  assign new_n39_ = new_n35_ & new_n36_;
  assign new_n40_ = new_n38_ & new_n39_;
  assign new_n41_ = i_9_ & i_8_;
  assign new_n42_ = i_6_ & new_n41_;
  assign new_n43_ = i_13_ & i_12_;
  assign new_n44_ = i_11_ & new_n43_;
  assign new_n45_ = i_3_ & i_4_;
  assign new_n46_ = i_1_ & new_n45_;
  assign new_n47_ = new_n42_ & new_n44_;
  assign new_n48_ = new_n46_ & new_n47_;
  assign new_n49_ = new_n40_ & new_n48_;
  assign new_n50_ = i_8_ & i_6_;
  assign new_n51_ = i_5_ & new_n50_;
  assign new_n52_ = i_12_ & i_11_;
  assign new_n53_ = i_9_ & new_n52_;
  assign new_n54_ = new_n51_ & new_n53_;
  assign new_n55_ = new_n46_ & new_n54_;
  assign new_n56_ = new_n40_ & new_n55_;
  assign new_n57_ = i_20_ & i_21_;
  assign new_n58_ = i_17_ & new_n57_;
  assign new_n59_ = i_23_ & ~i_24_;
  assign new_n60_ = i_22_ & new_n59_;
  assign new_n61_ = i_14_ & i_16_;
  assign new_n62_ = i_12_ & new_n61_;
  assign new_n63_ = new_n58_ & new_n60_;
  assign new_n64_ = new_n62_ & new_n63_;
  assign new_n65_ = i_4_ & new_n50_;
  assign new_n66_ = ~i_10_ & i_11_;
  assign new_n67_ = i_9_ & new_n66_;
  assign new_n68_ = i_3_ & ~i_2_;
  assign new_n69_ = i_1_ & new_n68_;
  assign new_n70_ = new_n65_ & new_n67_;
  assign new_n71_ = new_n69_ & new_n70_;
  assign new_n72_ = new_n64_ & new_n71_;
  assign new_n73_ = i_20_ & i_17_;
  assign new_n74_ = i_16_ & new_n73_;
  assign new_n75_ = i_14_ & i_15_;
  assign new_n76_ = i_13_ & new_n75_;
  assign new_n77_ = new_n60_ & new_n74_;
  assign new_n78_ = new_n76_ & new_n77_;
  assign new_n79_ = new_n55_ & new_n78_;
  assign new_n80_ = ~new_n56_ & ~new_n72_;
  assign new_n81_ = ~new_n79_ & new_n80_;
  assign new_n82_ = ~i_20_ & ~i_22_;
  assign new_n83_ = ~i_17_ & new_n82_;
  assign new_n84_ = ~i_23_ & i_24_;
  assign new_n85_ = ~i_14_ & ~i_16_;
  assign new_n86_ = ~i_12_ & new_n85_;
  assign new_n87_ = new_n83_ & new_n84_;
  assign new_n88_ = new_n86_ & new_n87_;
  assign new_n89_ = i_7_ & ~i_6_;
  assign new_n90_ = i_5_ & new_n89_;
  assign new_n91_ = ~i_9_ & ~i_11_;
  assign new_n92_ = ~i_8_ & new_n91_;
  assign new_n93_ = ~i_3_ & ~i_4_;
  assign new_n94_ = ~i_1_ & new_n93_;
  assign new_n95_ = new_n90_ & new_n92_;
  assign new_n96_ = new_n94_ & new_n95_;
  assign new_n97_ = new_n88_ & new_n96_;
  assign new_n98_ = ~i_20_ & ~i_17_;
  assign new_n99_ = ~i_16_ & new_n98_;
  assign new_n100_ = ~i_23_ & ~i_24_;
  assign new_n101_ = ~i_22_ & new_n100_;
  assign new_n102_ = ~i_14_ & ~i_12_;
  assign new_n103_ = ~i_11_ & new_n102_;
  assign new_n104_ = new_n99_ & new_n101_;
  assign new_n105_ = new_n103_ & new_n104_;
  assign new_n106_ = ~i_6_ & ~i_4_;
  assign new_n107_ = ~i_3_ & new_n106_;
  assign new_n108_ = ~i_9_ & ~i_10_;
  assign new_n109_ = ~i_8_ & new_n108_;
  assign new_n110_ = ~i_1_ & ~i_2_;
  assign new_n111_ = i_0_ & new_n110_;
  assign new_n112_ = new_n107_ & new_n109_;
  assign new_n113_ = new_n111_ & new_n112_;
  assign new_n114_ = new_n105_ & new_n113_;
  assign new_n115_ = ~i_20_ & i_19_;
  assign new_n116_ = ~i_17_ & new_n115_;
  assign new_n117_ = i_13_ & new_n85_;
  assign new_n118_ = new_n101_ & new_n116_;
  assign new_n119_ = new_n117_ & new_n118_;
  assign new_n120_ = ~i_8_ & ~i_6_;
  assign new_n121_ = i_5_ & new_n120_;
  assign new_n122_ = ~i_12_ & ~i_11_;
  assign new_n123_ = ~i_9_ & new_n122_;
  assign new_n124_ = new_n121_ & new_n123_;
  assign new_n125_ = new_n94_ & new_n124_;
  assign new_n126_ = new_n119_ & new_n125_;
  assign new_n127_ = ~new_n97_ & ~new_n114_;
  assign new_n128_ = ~new_n126_ & new_n127_;
  assign new_n129_ = ~i_23_ & ~i_22_;
  assign new_n130_ = ~i_13_ & new_n85_;
  assign new_n131_ = new_n116_ & new_n129_;
  assign new_n132_ = new_n130_ & new_n131_;
  assign new_n133_ = ~i_5_ & new_n120_;
  assign new_n134_ = new_n123_ & new_n133_;
  assign new_n135_ = new_n94_ & new_n134_;
  assign new_n136_ = new_n132_ & new_n135_;
  assign new_n137_ = new_n87_ & new_n117_;
  assign new_n138_ = i_7_ & ~i_8_;
  assign new_n139_ = ~i_6_ & new_n138_;
  assign new_n140_ = new_n123_ & new_n139_;
  assign new_n141_ = new_n94_ & new_n140_;
  assign new_n142_ = new_n137_ & new_n141_;
  assign new_n143_ = i_23_ & i_22_;
  assign new_n144_ = ~i_13_ & new_n75_;
  assign new_n145_ = new_n74_ & new_n143_;
  assign new_n146_ = new_n144_ & new_n145_;
  assign new_n147_ = ~i_5_ & new_n50_;
  assign new_n148_ = new_n53_ & new_n147_;
  assign new_n149_ = new_n46_ & new_n148_;
  assign new_n150_ = new_n146_ & new_n149_;
  assign new_n151_ = ~new_n136_ & ~new_n142_;
  assign new_n152_ = ~new_n150_ & new_n151_;
  assign new_n153_ = new_n81_ & new_n128_;
  assign new_n154_ = new_n152_ & new_n153_;
  assign o_1_ = new_n49_ | ~new_n154_;
  assign new_n156_ = i_14_ & i_13_;
  assign new_n157_ = i_11_ & new_n156_;
  assign new_n158_ = i_20_ & i_24_;
  assign new_n159_ = i_18_ & new_n158_;
  assign new_n160_ = i_6_ & i_3_;
  assign new_n161_ = i_1_ & new_n160_;
  assign new_n162_ = new_n157_ & new_n159_;
  assign new_n163_ = new_n161_ & new_n162_;
  assign new_n164_ = i_6_ & new_n66_;
  assign new_n165_ = i_14_ & new_n57_;
  assign new_n166_ = new_n164_ & new_n165_;
  assign new_n167_ = new_n69_ & new_n166_;
  assign new_n168_ = ~i_24_ & new_n167_;
  assign new_n169_ = ~new_n163_ & ~new_n168_;
  assign new_n170_ = i_13_ & i_11_;
  assign new_n171_ = i_6_ & new_n170_;
  assign new_n172_ = i_20_ & i_15_;
  assign new_n173_ = i_14_ & new_n172_;
  assign new_n174_ = i_5_ & i_3_;
  assign new_n175_ = i_1_ & new_n174_;
  assign new_n176_ = new_n171_ & new_n173_;
  assign new_n177_ = new_n175_ & new_n176_;
  assign new_n178_ = ~i_24_ & new_n177_;
  assign new_n179_ = i_14_ & i_11_;
  assign new_n180_ = i_6_ & new_n179_;
  assign new_n181_ = new_n159_ & new_n180_;
  assign new_n182_ = new_n175_ & new_n181_;
  assign new_n183_ = ~i_13_ & i_11_;
  assign new_n184_ = i_6_ & new_n183_;
  assign new_n185_ = ~i_5_ & i_3_;
  assign new_n186_ = i_1_ & new_n185_;
  assign new_n187_ = new_n173_ & new_n184_;
  assign new_n188_ = new_n186_ & new_n187_;
  assign new_n189_ = ~new_n178_ & ~new_n182_;
  assign new_n190_ = ~new_n188_ & new_n189_;
  assign o_2_ = ~new_n169_ | ~new_n190_;
  assign new_n192_ = i_13_ & ~i_11_;
  assign new_n193_ = i_7_ & new_n192_;
  assign new_n194_ = ~i_20_ & i_24_;
  assign new_n195_ = ~i_14_ & new_n194_;
  assign new_n196_ = ~i_6_ & ~i_3_;
  assign new_n197_ = ~i_1_ & new_n196_;
  assign new_n198_ = new_n193_ & new_n195_;
  assign new_n199_ = new_n197_ & new_n198_;
  assign new_n200_ = ~i_10_ & ~i_6_;
  assign new_n201_ = ~i_3_ & new_n200_;
  assign new_n202_ = ~i_20_ & ~i_14_;
  assign new_n203_ = ~i_11_ & new_n202_;
  assign new_n204_ = new_n201_ & new_n203_;
  assign new_n205_ = new_n111_ & new_n204_;
  assign new_n206_ = ~i_24_ & new_n205_;
  assign new_n207_ = ~new_n199_ & ~new_n206_;
  assign new_n208_ = ~i_6_ & new_n192_;
  assign new_n209_ = ~i_14_ & new_n115_;
  assign new_n210_ = i_5_ & ~i_3_;
  assign new_n211_ = ~i_1_ & new_n210_;
  assign new_n212_ = new_n208_ & new_n209_;
  assign new_n213_ = new_n211_ & new_n212_;
  assign new_n214_ = ~i_24_ & new_n213_;
  assign new_n215_ = i_7_ & ~i_11_;
  assign new_n216_ = ~i_6_ & new_n215_;
  assign new_n217_ = new_n195_ & new_n216_;
  assign new_n218_ = new_n211_ & new_n217_;
  assign new_n219_ = ~i_13_ & ~i_11_;
  assign new_n220_ = ~i_6_ & new_n219_;
  assign new_n221_ = ~i_5_ & ~i_3_;
  assign new_n222_ = ~i_1_ & new_n221_;
  assign new_n223_ = new_n209_ & new_n220_;
  assign new_n224_ = new_n222_ & new_n223_;
  assign new_n225_ = ~new_n214_ & ~new_n218_;
  assign new_n226_ = ~new_n224_ & new_n225_;
  assign o_0_ = ~new_n207_ | ~new_n226_;
  assign new_n228_ = i_18_ & i_24_;
  assign new_n229_ = i_5_ & new_n228_;
  assign new_n230_ = ~i_10_ & i_21_;
  assign new_n231_ = ~i_2_ & new_n230_;
  assign new_n232_ = ~i_24_ & new_n231_;
  assign new_n233_ = ~new_n229_ & ~new_n232_;
  assign new_n234_ = i_13_ & new_n228_;
  assign new_n235_ = i_13_ & i_15_;
  assign new_n236_ = i_5_ & new_n235_;
  assign new_n237_ = ~i_24_ & new_n236_;
  assign new_n238_ = ~i_13_ & i_15_;
  assign new_n239_ = ~i_5_ & new_n238_;
  assign new_n240_ = ~new_n234_ & ~new_n237_;
  assign new_n241_ = ~new_n239_ & new_n240_;
  assign o_7_ = ~new_n233_ | ~new_n241_;
  assign new_n243_ = i_13_ & i_24_;
  assign new_n244_ = i_7_ & new_n243_;
  assign new_n245_ = ~i_10_ & ~i_2_;
  assign new_n246_ = i_0_ & new_n245_;
  assign new_n247_ = ~i_24_ & new_n246_;
  assign new_n248_ = ~new_n244_ & ~new_n247_;
  assign new_n249_ = i_13_ & i_19_;
  assign new_n250_ = i_5_ & new_n249_;
  assign new_n251_ = ~i_24_ & new_n250_;
  assign new_n252_ = i_7_ & i_24_;
  assign new_n253_ = i_5_ & new_n252_;
  assign new_n254_ = ~i_13_ & i_19_;
  assign new_n255_ = ~i_5_ & new_n254_;
  assign new_n256_ = ~new_n251_ & ~new_n253_;
  assign new_n257_ = ~new_n255_ & new_n256_;
  assign o_5_ = ~new_n248_ | ~new_n257_;
  assign new_n259_ = ~i_20_ & i_21_;
  assign new_n260_ = i_14_ & new_n259_;
  assign new_n261_ = ~i_2_ & new_n66_;
  assign new_n262_ = ~i_24_ & new_n260_;
  assign new_n263_ = new_n261_ & new_n262_;
  assign new_n264_ = i_7_ & i_13_;
  assign new_n265_ = i_3_ & new_n264_;
  assign new_n266_ = i_24_ & new_n265_;
  assign new_n267_ = i_20_ & ~i_14_;
  assign new_n268_ = ~i_11_ & new_n267_;
  assign new_n269_ = ~i_24_ & new_n268_;
  assign new_n270_ = new_n246_ & new_n269_;
  assign new_n271_ = ~new_n263_ & ~new_n266_;
  assign new_n272_ = ~new_n270_ & new_n271_;
  assign new_n273_ = i_6_ & ~i_11_;
  assign new_n274_ = ~i_5_ & new_n273_;
  assign new_n275_ = new_n254_ & new_n274_;
  assign new_n276_ = ~i_24_ & i_19_;
  assign new_n277_ = i_13_ & new_n276_;
  assign new_n278_ = i_5_ & new_n273_;
  assign new_n279_ = new_n277_ & new_n278_;
  assign new_n280_ = i_6_ & new_n215_;
  assign new_n281_ = new_n243_ & new_n280_;
  assign new_n282_ = ~new_n275_ & ~new_n279_;
  assign new_n283_ = ~new_n281_ & new_n282_;
  assign new_n284_ = ~i_24_ & i_15_;
  assign new_n285_ = i_13_ & new_n284_;
  assign new_n286_ = ~i_6_ & i_11_;
  assign new_n287_ = i_5_ & new_n286_;
  assign new_n288_ = new_n285_ & new_n287_;
  assign new_n289_ = ~i_11_ & ~i_24_;
  assign new_n290_ = ~i_10_ & new_n289_;
  assign new_n291_ = i_6_ & ~i_2_;
  assign new_n292_ = i_0_ & new_n291_;
  assign new_n293_ = new_n290_ & new_n292_;
  assign new_n294_ = ~i_24_ & i_21_;
  assign new_n295_ = i_11_ & new_n294_;
  assign new_n296_ = ~i_2_ & new_n200_;
  assign new_n297_ = new_n295_ & new_n296_;
  assign new_n298_ = ~new_n288_ & ~new_n293_;
  assign new_n299_ = ~new_n297_ & new_n298_;
  assign new_n300_ = ~i_5_ & new_n286_;
  assign new_n301_ = new_n238_ & new_n300_;
  assign new_n302_ = ~i_6_ & new_n170_;
  assign new_n303_ = new_n228_ & new_n302_;
  assign new_n304_ = ~i_11_ & i_24_;
  assign new_n305_ = i_7_ & i_6_;
  assign new_n306_ = i_5_ & new_n305_;
  assign new_n307_ = new_n304_ & new_n306_;
  assign new_n308_ = ~new_n301_ & ~new_n303_;
  assign new_n309_ = ~new_n307_ & new_n308_;
  assign new_n310_ = new_n283_ & new_n299_;
  assign new_n311_ = new_n309_ & new_n310_;
  assign new_n312_ = i_20_ & i_19_;
  assign new_n313_ = ~i_14_ & new_n312_;
  assign new_n314_ = ~i_5_ & new_n219_;
  assign new_n315_ = new_n313_ & new_n314_;
  assign new_n316_ = ~i_20_ & i_15_;
  assign new_n317_ = i_14_ & new_n316_;
  assign new_n318_ = ~i_5_ & new_n183_;
  assign new_n319_ = new_n317_ & new_n318_;
  assign new_n320_ = ~i_14_ & new_n158_;
  assign new_n321_ = new_n193_ & new_n320_;
  assign new_n322_ = ~new_n315_ & ~new_n319_;
  assign new_n323_ = ~new_n321_ & new_n322_;
  assign new_n324_ = i_5_ & new_n170_;
  assign new_n325_ = ~i_24_ & new_n317_;
  assign new_n326_ = new_n324_ & new_n325_;
  assign new_n327_ = i_18_ & new_n194_;
  assign new_n328_ = i_5_ & new_n179_;
  assign new_n329_ = new_n327_ & new_n328_;
  assign new_n330_ = i_5_ & new_n192_;
  assign new_n331_ = ~i_24_ & new_n313_;
  assign new_n332_ = new_n330_ & new_n331_;
  assign new_n333_ = ~new_n326_ & ~new_n329_;
  assign new_n334_ = ~new_n332_ & new_n333_;
  assign new_n335_ = i_5_ & new_n215_;
  assign new_n336_ = new_n320_ & new_n335_;
  assign new_n337_ = new_n157_ & new_n327_;
  assign new_n338_ = new_n228_ & new_n287_;
  assign new_n339_ = ~new_n336_ & ~new_n337_;
  assign new_n340_ = ~new_n338_ & new_n339_;
  assign new_n341_ = new_n323_ & new_n334_;
  assign new_n342_ = new_n340_ & new_n341_;
  assign new_n343_ = i_7_ & i_5_;
  assign new_n344_ = i_3_ & new_n343_;
  assign new_n345_ = i_24_ & new_n344_;
  assign new_n346_ = ~i_10_ & ~i_24_;
  assign new_n347_ = i_0_ & new_n68_;
  assign new_n348_ = new_n346_ & new_n347_;
  assign new_n349_ = ~i_10_ & ~i_3_;
  assign new_n350_ = ~i_2_ & new_n349_;
  assign new_n351_ = new_n294_ & new_n350_;
  assign new_n352_ = ~new_n345_ & ~new_n348_;
  assign new_n353_ = ~new_n351_ & new_n352_;
  assign new_n354_ = i_5_ & i_13_;
  assign new_n355_ = i_3_ & new_n354_;
  assign new_n356_ = new_n276_ & new_n355_;
  assign new_n357_ = ~i_3_ & new_n354_;
  assign new_n358_ = new_n284_ & new_n357_;
  assign new_n359_ = i_5_ & i_18_;
  assign new_n360_ = ~i_3_ & new_n359_;
  assign new_n361_ = i_24_ & new_n360_;
  assign new_n362_ = ~new_n356_ & ~new_n358_;
  assign new_n363_ = ~new_n361_ & new_n362_;
  assign new_n364_ = i_13_ & i_18_;
  assign new_n365_ = ~i_3_ & new_n364_;
  assign new_n366_ = i_24_ & new_n365_;
  assign new_n367_ = ~i_5_ & ~i_13_;
  assign new_n368_ = ~i_3_ & new_n367_;
  assign new_n369_ = i_15_ & new_n368_;
  assign new_n370_ = i_3_ & new_n367_;
  assign new_n371_ = i_19_ & new_n370_;
  assign new_n372_ = ~new_n366_ & ~new_n369_;
  assign new_n373_ = ~new_n371_ & new_n372_;
  assign new_n374_ = new_n353_ & new_n363_;
  assign new_n375_ = new_n373_ & new_n374_;
  assign new_n376_ = new_n311_ & new_n342_;
  assign new_n377_ = new_n375_ & new_n376_;
  assign o_6_ = ~new_n272_ | ~new_n377_;
  assign new_n379_ = i_8_ & new_n170_;
  assign new_n380_ = i_20_ & i_18_;
  assign new_n381_ = i_14_ & new_n380_;
  assign new_n382_ = new_n379_ & new_n381_;
  assign new_n383_ = new_n161_ & new_n382_;
  assign new_n384_ = i_24_ & new_n383_;
  assign new_n385_ = i_8_ & i_11_;
  assign new_n386_ = i_6_ & new_n385_;
  assign new_n387_ = new_n381_ & new_n386_;
  assign new_n388_ = new_n175_ & new_n387_;
  assign new_n389_ = i_24_ & new_n388_;
  assign new_n390_ = ~i_10_ & i_8_;
  assign new_n391_ = i_6_ & new_n390_;
  assign new_n392_ = i_20_ & i_14_;
  assign new_n393_ = i_11_ & new_n392_;
  assign new_n394_ = new_n391_ & new_n393_;
  assign new_n395_ = new_n69_ & new_n394_;
  assign new_n396_ = new_n294_ & new_n395_;
  assign new_n397_ = i_20_ & ~i_24_;
  assign new_n398_ = new_n76_ & new_n386_;
  assign new_n399_ = new_n175_ & new_n398_;
  assign new_n400_ = new_n397_ & new_n399_;
  assign new_n401_ = ~new_n389_ & ~new_n396_;
  assign new_n402_ = ~new_n400_ & new_n401_;
  assign new_n403_ = ~i_20_ & ~i_24_;
  assign new_n404_ = ~i_8_ & ~i_11_;
  assign new_n405_ = ~i_6_ & new_n404_;
  assign new_n406_ = ~i_14_ & i_19_;
  assign new_n407_ = i_13_ & new_n406_;
  assign new_n408_ = new_n405_ & new_n407_;
  assign new_n409_ = new_n211_ & new_n408_;
  assign new_n410_ = new_n403_ & new_n409_;
  assign new_n411_ = ~i_3_ & new_n120_;
  assign new_n412_ = ~i_14_ & ~i_11_;
  assign new_n413_ = ~i_10_ & new_n412_;
  assign new_n414_ = new_n411_ & new_n413_;
  assign new_n415_ = new_n111_ & new_n414_;
  assign new_n416_ = new_n403_ & new_n415_;
  assign new_n417_ = new_n139_ & new_n203_;
  assign new_n418_ = new_n211_ & new_n417_;
  assign new_n419_ = i_24_ & new_n418_;
  assign new_n420_ = ~new_n410_ & ~new_n416_;
  assign new_n421_ = ~new_n419_ & new_n420_;
  assign new_n422_ = ~i_13_ & new_n406_;
  assign new_n423_ = new_n405_ & new_n422_;
  assign new_n424_ = new_n222_ & new_n423_;
  assign new_n425_ = ~i_20_ & new_n424_;
  assign new_n426_ = i_7_ & new_n404_;
  assign new_n427_ = i_13_ & new_n202_;
  assign new_n428_ = new_n426_ & new_n427_;
  assign new_n429_ = new_n197_ & new_n428_;
  assign new_n430_ = i_24_ & new_n429_;
  assign new_n431_ = new_n144_ & new_n386_;
  assign new_n432_ = new_n186_ & new_n431_;
  assign new_n433_ = i_20_ & new_n432_;
  assign new_n434_ = ~new_n425_ & ~new_n430_;
  assign new_n435_ = ~new_n433_ & new_n434_;
  assign new_n436_ = new_n402_ & new_n421_;
  assign new_n437_ = new_n435_ & new_n436_;
  assign o_3_ = new_n384_ | ~new_n437_;
  assign new_n439_ = i_8_ & i_13_;
  assign new_n440_ = i_7_ & new_n439_;
  assign new_n441_ = i_24_ & new_n440_;
  assign new_n442_ = i_21_ & i_22_;
  assign new_n443_ = i_16_ & new_n442_;
  assign new_n444_ = ~i_10_ & ~i_4_;
  assign new_n445_ = ~i_2_ & new_n444_;
  assign new_n446_ = new_n59_ & new_n443_;
  assign new_n447_ = new_n445_ & new_n446_;
  assign new_n448_ = ~i_16_ & ~i_22_;
  assign new_n449_ = ~i_10_ & new_n448_;
  assign new_n450_ = i_4_ & ~i_2_;
  assign new_n451_ = i_0_ & new_n450_;
  assign new_n452_ = new_n100_ & new_n449_;
  assign new_n453_ = new_n451_ & new_n452_;
  assign new_n454_ = i_16_ & i_22_;
  assign new_n455_ = i_15_ & new_n454_;
  assign new_n456_ = ~i_4_ & new_n354_;
  assign new_n457_ = new_n59_ & new_n455_;
  assign new_n458_ = new_n456_ & new_n457_;
  assign new_n459_ = ~new_n447_ & ~new_n453_;
  assign new_n460_ = ~new_n458_ & new_n459_;
  assign new_n461_ = ~new_n441_ & new_n460_;
  assign new_n462_ = ~i_22_ & i_19_;
  assign new_n463_ = ~i_16_ & new_n462_;
  assign new_n464_ = i_4_ & new_n367_;
  assign new_n465_ = ~i_23_ & new_n463_;
  assign new_n466_ = new_n464_ & new_n465_;
  assign new_n467_ = ~i_16_ & new_n129_;
  assign new_n468_ = i_4_ & new_n264_;
  assign new_n469_ = i_24_ & new_n467_;
  assign new_n470_ = new_n468_ & new_n469_;
  assign new_n471_ = ~i_4_ & new_n367_;
  assign new_n472_ = i_23_ & new_n455_;
  assign new_n473_ = new_n471_ & new_n472_;
  assign new_n474_ = ~new_n466_ & ~new_n470_;
  assign new_n475_ = ~new_n473_ & new_n474_;
  assign new_n476_ = i_4_ & new_n354_;
  assign new_n477_ = new_n100_ & new_n463_;
  assign new_n478_ = new_n476_ & new_n477_;
  assign new_n479_ = i_4_ & new_n343_;
  assign new_n480_ = new_n469_ & new_n479_;
  assign new_n481_ = i_18_ & new_n143_;
  assign new_n482_ = i_5_ & i_16_;
  assign new_n483_ = ~i_4_ & new_n482_;
  assign new_n484_ = i_24_ & new_n481_;
  assign new_n485_ = new_n483_ & new_n484_;
  assign new_n486_ = ~new_n478_ & ~new_n480_;
  assign new_n487_ = ~new_n485_ & new_n486_;
  assign new_n488_ = i_17_ & ~i_22_;
  assign new_n489_ = ~i_16_ & new_n488_;
  assign new_n490_ = ~i_24_ & new_n489_;
  assign new_n491_ = new_n246_ & new_n490_;
  assign new_n492_ = i_13_ & i_16_;
  assign new_n493_ = ~i_4_ & new_n492_;
  assign new_n494_ = new_n484_ & new_n493_;
  assign new_n495_ = ~i_17_ & i_22_;
  assign new_n496_ = i_16_ & new_n495_;
  assign new_n497_ = ~i_24_ & new_n496_;
  assign new_n498_ = new_n236_ & new_n497_;
  assign new_n499_ = ~new_n491_ & ~new_n494_;
  assign new_n500_ = ~new_n498_ & new_n499_;
  assign new_n501_ = new_n475_ & new_n487_;
  assign new_n502_ = new_n500_ & new_n501_;
  assign new_n503_ = new_n461_ & new_n502_;
  assign new_n504_ = ~i_9_ & i_16_;
  assign new_n505_ = i_5_ & new_n504_;
  assign new_n506_ = new_n228_ & new_n505_;
  assign new_n507_ = i_24_ & ~i_16_;
  assign new_n508_ = i_9_ & i_7_;
  assign new_n509_ = i_5_ & new_n508_;
  assign new_n510_ = new_n507_ & new_n509_;
  assign new_n511_ = i_16_ & i_15_;
  assign new_n512_ = ~i_9_ & ~i_13_;
  assign new_n513_ = ~i_5_ & new_n512_;
  assign new_n514_ = new_n511_ & new_n513_;
  assign new_n515_ = ~new_n506_ & ~new_n510_;
  assign new_n516_ = ~new_n514_ & new_n515_;
  assign new_n517_ = ~i_16_ & new_n276_;
  assign new_n518_ = i_9_ & i_13_;
  assign new_n519_ = i_5_ & new_n518_;
  assign new_n520_ = new_n517_ & new_n519_;
  assign new_n521_ = i_16_ & new_n294_;
  assign new_n522_ = ~i_2_ & new_n108_;
  assign new_n523_ = new_n521_ & new_n522_;
  assign new_n524_ = ~i_24_ & i_16_;
  assign new_n525_ = i_15_ & new_n524_;
  assign new_n526_ = ~i_9_ & i_13_;
  assign new_n527_ = i_5_ & new_n526_;
  assign new_n528_ = new_n525_ & new_n527_;
  assign new_n529_ = ~new_n520_ & ~new_n523_;
  assign new_n530_ = ~new_n528_ & new_n529_;
  assign new_n531_ = i_7_ & new_n518_;
  assign new_n532_ = new_n507_ & new_n531_;
  assign new_n533_ = ~i_16_ & i_19_;
  assign new_n534_ = i_9_ & ~i_13_;
  assign new_n535_ = ~i_5_ & new_n534_;
  assign new_n536_ = new_n533_ & new_n535_;
  assign new_n537_ = ~i_9_ & new_n492_;
  assign new_n538_ = new_n228_ & new_n537_;
  assign new_n539_ = ~new_n532_ & ~new_n536_;
  assign new_n540_ = ~new_n538_ & new_n539_;
  assign new_n541_ = new_n516_ & new_n530_;
  assign new_n542_ = new_n540_ & new_n541_;
  assign new_n543_ = i_24_ & ~i_22_;
  assign new_n544_ = i_17_ & new_n543_;
  assign new_n545_ = i_13_ & ~i_16_;
  assign new_n546_ = i_7_ & new_n545_;
  assign new_n547_ = new_n544_ & new_n546_;
  assign new_n548_ = i_7_ & ~i_16_;
  assign new_n549_ = i_5_ & new_n548_;
  assign new_n550_ = new_n544_ & new_n549_;
  assign new_n551_ = new_n239_ & new_n496_;
  assign new_n552_ = ~new_n547_ & ~new_n550_;
  assign new_n553_ = ~new_n551_ & new_n552_;
  assign new_n554_ = i_24_ & i_22_;
  assign new_n555_ = i_18_ & new_n554_;
  assign new_n556_ = ~i_17_ & i_16_;
  assign new_n557_ = i_5_ & new_n556_;
  assign new_n558_ = new_n555_ & new_n557_;
  assign new_n559_ = ~i_17_ & new_n442_;
  assign new_n560_ = ~i_10_ & i_16_;
  assign new_n561_ = ~i_2_ & new_n560_;
  assign new_n562_ = ~i_24_ & new_n559_;
  assign new_n563_ = new_n561_ & new_n562_;
  assign new_n564_ = i_17_ & new_n462_;
  assign new_n565_ = i_5_ & new_n545_;
  assign new_n566_ = ~i_24_ & new_n564_;
  assign new_n567_ = new_n565_ & new_n566_;
  assign new_n568_ = ~new_n558_ & ~new_n563_;
  assign new_n569_ = ~new_n567_ & new_n568_;
  assign new_n570_ = ~i_13_ & ~i_16_;
  assign new_n571_ = ~i_5_ & new_n570_;
  assign new_n572_ = new_n564_ & new_n571_;
  assign new_n573_ = i_13_ & new_n556_;
  assign new_n574_ = new_n555_ & new_n573_;
  assign new_n575_ = ~i_24_ & ~i_16_;
  assign new_n576_ = ~i_10_ & new_n575_;
  assign new_n577_ = i_9_ & ~i_2_;
  assign new_n578_ = i_0_ & new_n577_;
  assign new_n579_ = new_n576_ & new_n578_;
  assign new_n580_ = ~new_n572_ & ~new_n574_;
  assign new_n581_ = ~new_n579_ & new_n580_;
  assign new_n582_ = new_n553_ & new_n569_;
  assign new_n583_ = new_n581_ & new_n582_;
  assign new_n584_ = i_5_ & new_n439_;
  assign new_n585_ = new_n276_ & new_n584_;
  assign new_n586_ = ~i_8_ & i_18_;
  assign new_n587_ = i_5_ & new_n586_;
  assign new_n588_ = i_24_ & new_n587_;
  assign new_n589_ = i_7_ & i_8_;
  assign new_n590_ = i_5_ & new_n589_;
  assign new_n591_ = i_24_ & new_n590_;
  assign new_n592_ = ~new_n585_ & ~new_n588_;
  assign new_n593_ = ~new_n591_ & new_n592_;
  assign new_n594_ = ~i_10_ & ~i_8_;
  assign new_n595_ = ~i_2_ & new_n594_;
  assign new_n596_ = new_n294_ & new_n595_;
  assign new_n597_ = ~i_8_ & i_13_;
  assign new_n598_ = i_5_ & new_n597_;
  assign new_n599_ = new_n284_ & new_n598_;
  assign new_n600_ = i_8_ & ~i_2_;
  assign new_n601_ = i_0_ & new_n600_;
  assign new_n602_ = new_n346_ & new_n601_;
  assign new_n603_ = ~new_n596_ & ~new_n599_;
  assign new_n604_ = ~new_n602_ & new_n603_;
  assign new_n605_ = ~i_8_ & new_n364_;
  assign new_n606_ = i_24_ & new_n605_;
  assign new_n607_ = ~i_8_ & ~i_13_;
  assign new_n608_ = ~i_5_ & new_n607_;
  assign new_n609_ = i_15_ & new_n608_;
  assign new_n610_ = i_8_ & ~i_13_;
  assign new_n611_ = ~i_5_ & new_n610_;
  assign new_n612_ = i_19_ & new_n611_;
  assign new_n613_ = ~new_n606_ & ~new_n609_;
  assign new_n614_ = ~new_n612_ & new_n613_;
  assign new_n615_ = new_n593_ & new_n604_;
  assign new_n616_ = new_n614_ & new_n615_;
  assign new_n617_ = new_n542_ & new_n583_;
  assign new_n618_ = new_n616_ & new_n617_;
  assign o_4_ = ~new_n503_ | ~new_n618_;
endmodule

