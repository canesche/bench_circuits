// Benchmark "ac97_ctrl" written by ABC on Thu Oct  8 22:03:22 2020

module ac97_ctrl ( clock, 
    clk_i, rst_i, wb_we_i, wb_cyc_i, wb_stb_i, bit_clk_pad_i, sdata_pad_i,
    \wb_data_i[0] , \wb_data_i[1] , \wb_data_i[2] , \wb_data_i[3] ,
    \wb_data_i[4] , \wb_data_i[5] , \wb_data_i[6] , \wb_data_i[7] ,
    \wb_data_i[8] , \wb_data_i[9] , \wb_data_i[10] , \wb_data_i[11] ,
    \wb_data_i[12] , \wb_data_i[13] , \wb_data_i[14] , \wb_data_i[15] ,
    \wb_data_i[16] , \wb_data_i[17] , \wb_data_i[18] , \wb_data_i[19] ,
    \wb_data_i[20] , \wb_data_i[21] , \wb_data_i[22] , \wb_data_i[23] ,
    \wb_data_i[24] , \wb_data_i[25] , \wb_data_i[26] , \wb_data_i[27] ,
    \wb_data_i[28] , \wb_data_i[29] , \wb_data_i[30] , \wb_data_i[31] ,
    \wb_addr_i[0] , \wb_addr_i[1] , \wb_addr_i[2] , \wb_addr_i[3] ,
    \wb_addr_i[4] , \wb_addr_i[5] , \wb_addr_i[6] , \wb_addr_i[7] ,
    \wb_addr_i[8] , \wb_addr_i[9] , \wb_addr_i[10] , \wb_addr_i[11] ,
    \wb_addr_i[12] , \wb_addr_i[13] , \wb_addr_i[14] , \wb_addr_i[15] ,
    \wb_addr_i[16] , \wb_addr_i[17] , \wb_addr_i[18] , \wb_addr_i[19] ,
    \wb_addr_i[20] , \wb_addr_i[21] , \wb_addr_i[22] , \wb_addr_i[23] ,
    \wb_addr_i[24] , \wb_addr_i[25] , \wb_addr_i[26] , \wb_addr_i[27] ,
    \wb_addr_i[28] , \wb_addr_i[29] , \wb_addr_i[30] , \wb_addr_i[31] ,
    \wb_sel_i[0] , \wb_sel_i[1] , \wb_sel_i[2] , \wb_sel_i[3] ,
    \dma_ack_i[0] , \dma_ack_i[1] , \dma_ack_i[2] , \dma_ack_i[3] ,
    \dma_ack_i[4] , \dma_ack_i[5] , \dma_ack_i[6] , \dma_ack_i[7] ,
    \dma_ack_i[8] ,
    \wb_data_o[0] , \wb_data_o[1] , \wb_data_o[2] , \wb_data_o[3] ,
    \wb_data_o[4] , \wb_data_o[5] , \wb_data_o[6] , \wb_data_o[7] ,
    \wb_data_o[8] , \wb_data_o[9] , \wb_data_o[10] , \wb_data_o[11] ,
    \wb_data_o[12] , \wb_data_o[13] , \wb_data_o[14] , \wb_data_o[15] ,
    \wb_data_o[16] , \wb_data_o[17] , \wb_data_o[18] , \wb_data_o[19] ,
    \wb_data_o[20] , \wb_data_o[21] , \wb_data_o[22] , \wb_data_o[23] ,
    \wb_data_o[24] , \wb_data_o[25] , \wb_data_o[26] , \wb_data_o[27] ,
    \wb_data_o[28] , \wb_data_o[29] , \wb_data_o[30] , \wb_data_o[31] ,
    wb_ack_o, wb_err_o, int_o, suspended_o, sync_pad_o, sdata_pad_o,
    ac97_reset_pad_o_, \dma_req_o[0] , \dma_req_o[1] , \dma_req_o[2] ,
    \dma_req_o[3] , \dma_req_o[4] , \dma_req_o[5] , \dma_req_o[6] ,
    \dma_req_o[7] , \dma_req_o[8]   );
  input  clock;
  input  clk_i, rst_i, wb_we_i, wb_cyc_i, wb_stb_i, bit_clk_pad_i,
    sdata_pad_i, \wb_data_i[0] , \wb_data_i[1] , \wb_data_i[2] ,
    \wb_data_i[3] , \wb_data_i[4] , \wb_data_i[5] , \wb_data_i[6] ,
    \wb_data_i[7] , \wb_data_i[8] , \wb_data_i[9] , \wb_data_i[10] ,
    \wb_data_i[11] , \wb_data_i[12] , \wb_data_i[13] , \wb_data_i[14] ,
    \wb_data_i[15] , \wb_data_i[16] , \wb_data_i[17] , \wb_data_i[18] ,
    \wb_data_i[19] , \wb_data_i[20] , \wb_data_i[21] , \wb_data_i[22] ,
    \wb_data_i[23] , \wb_data_i[24] , \wb_data_i[25] , \wb_data_i[26] ,
    \wb_data_i[27] , \wb_data_i[28] , \wb_data_i[29] , \wb_data_i[30] ,
    \wb_data_i[31] , \wb_addr_i[0] , \wb_addr_i[1] , \wb_addr_i[2] ,
    \wb_addr_i[3] , \wb_addr_i[4] , \wb_addr_i[5] , \wb_addr_i[6] ,
    \wb_addr_i[7] , \wb_addr_i[8] , \wb_addr_i[9] , \wb_addr_i[10] ,
    \wb_addr_i[11] , \wb_addr_i[12] , \wb_addr_i[13] , \wb_addr_i[14] ,
    \wb_addr_i[15] , \wb_addr_i[16] , \wb_addr_i[17] , \wb_addr_i[18] ,
    \wb_addr_i[19] , \wb_addr_i[20] , \wb_addr_i[21] , \wb_addr_i[22] ,
    \wb_addr_i[23] , \wb_addr_i[24] , \wb_addr_i[25] , \wb_addr_i[26] ,
    \wb_addr_i[27] , \wb_addr_i[28] , \wb_addr_i[29] , \wb_addr_i[30] ,
    \wb_addr_i[31] , \wb_sel_i[0] , \wb_sel_i[1] , \wb_sel_i[2] ,
    \wb_sel_i[3] , \dma_ack_i[0] , \dma_ack_i[1] , \dma_ack_i[2] ,
    \dma_ack_i[3] , \dma_ack_i[4] , \dma_ack_i[5] , \dma_ack_i[6] ,
    \dma_ack_i[7] , \dma_ack_i[8] ;
  output \wb_data_o[0] , \wb_data_o[1] , \wb_data_o[2] , \wb_data_o[3] ,
    \wb_data_o[4] , \wb_data_o[5] , \wb_data_o[6] , \wb_data_o[7] ,
    \wb_data_o[8] , \wb_data_o[9] , \wb_data_o[10] , \wb_data_o[11] ,
    \wb_data_o[12] , \wb_data_o[13] , \wb_data_o[14] , \wb_data_o[15] ,
    \wb_data_o[16] , \wb_data_o[17] , \wb_data_o[18] , \wb_data_o[19] ,
    \wb_data_o[20] , \wb_data_o[21] , \wb_data_o[22] , \wb_data_o[23] ,
    \wb_data_o[24] , \wb_data_o[25] , \wb_data_o[26] , \wb_data_o[27] ,
    \wb_data_o[28] , \wb_data_o[29] , \wb_data_o[30] , \wb_data_o[31] ,
    wb_ack_o, wb_err_o, int_o, suspended_o, sync_pad_o, sdata_pad_o,
    ac97_reset_pad_o_, \dma_req_o[0] , \dma_req_o[1] , \dma_req_o[2] ,
    \dma_req_o[3] , \dma_req_o[4] , \dma_req_o[5] , \dma_req_o[6] ,
    \dma_req_o[7] , \dma_req_o[8] ;
  reg \\u0_slt0_r_reg[15] , \\u0_slt0_r_reg[14] , \\u0_slt0_r_reg[13] ,
    \\u0_slt0_r_reg[12] , \\u0_slt0_r_reg[11] , \\u0_slt0_r_reg[10] ,
    \\u0_slt0_r_reg[9] , \\u0_slt0_r_reg[8] , \\u0_slt0_r_reg[7] ,
    \\u0_slt0_r_reg[6] , \\u0_slt0_r_reg[5] , \\u0_slt0_r_reg[4] ,
    \\u0_slt0_r_reg[3] , \\u0_slt0_r_reg[2] , \\u0_slt0_r_reg[1] ,
    \\u0_slt0_r_reg[0] , \\u0_slt1_r_reg[19] , \\u0_slt1_r_reg[18] ,
    \\u0_slt1_r_reg[17] , \\u0_slt1_r_reg[16] , \\u0_slt1_r_reg[15] ,
    \\u0_slt1_r_reg[14] , \\u0_slt1_r_reg[13] , \\u0_slt1_r_reg[12] ,
    \\u0_slt1_r_reg[11] , \\u0_slt1_r_reg[10] , \\u0_slt1_r_reg[9] ,
    \\u0_slt1_r_reg[8] , \\u0_slt1_r_reg[7] , \\u0_slt1_r_reg[6] ,
    \\u0_slt1_r_reg[5] , \\u0_slt1_r_reg[4] , \\u0_slt1_r_reg[3] ,
    \\u0_slt1_r_reg[2] , \\u0_slt1_r_reg[1] , \\u0_slt1_r_reg[0] ,
    \\u0_slt2_r_reg[19] , \\u0_slt2_r_reg[18] , \\u0_slt2_r_reg[17] ,
    \\u0_slt2_r_reg[16] , \\u0_slt2_r_reg[15] , \\u0_slt2_r_reg[14] ,
    \\u0_slt2_r_reg[13] , \\u0_slt2_r_reg[12] , \\u0_slt2_r_reg[11] ,
    \\u0_slt2_r_reg[10] , \\u0_slt2_r_reg[9] , \\u0_slt2_r_reg[8] ,
    \\u0_slt2_r_reg[7] , \\u0_slt2_r_reg[6] , \\u0_slt2_r_reg[5] ,
    \\u0_slt2_r_reg[4] , \\u0_slt2_r_reg[3] , \\u0_slt2_r_reg[2] ,
    \\u0_slt2_r_reg[1] , \\u0_slt2_r_reg[0] , \\u0_slt3_r_reg[19] ,
    \\u0_slt3_r_reg[18] , \\u0_slt3_r_reg[17] , \\u0_slt3_r_reg[16] ,
    \\u0_slt3_r_reg[15] , \\u0_slt3_r_reg[14] , \\u0_slt3_r_reg[13] ,
    \\u0_slt3_r_reg[12] , \\u0_slt3_r_reg[11] , \\u0_slt3_r_reg[10] ,
    \\u0_slt3_r_reg[9] , \\u0_slt3_r_reg[8] , \\u0_slt3_r_reg[7] ,
    \\u0_slt3_r_reg[6] , \\u0_slt3_r_reg[5] , \\u0_slt3_r_reg[4] ,
    \\u0_slt3_r_reg[3] , \\u0_slt3_r_reg[2] , \\u0_slt3_r_reg[1] ,
    \\u0_slt3_r_reg[0] , \\u0_slt4_r_reg[19] , \\u0_slt4_r_reg[18] ,
    \\u0_slt4_r_reg[17] , \\u0_slt4_r_reg[16] , \\u0_slt4_r_reg[15] ,
    \\u0_slt4_r_reg[14] , \\u0_slt4_r_reg[13] , \\u0_slt4_r_reg[12] ,
    \\u0_slt4_r_reg[11] , \\u0_slt4_r_reg[10] , \\u0_slt4_r_reg[9] ,
    \\u0_slt4_r_reg[8] , \\u0_slt4_r_reg[7] , \\u0_slt4_r_reg[6] ,
    \\u0_slt4_r_reg[5] , \\u0_slt4_r_reg[4] , \\u0_slt4_r_reg[3] ,
    \\u0_slt4_r_reg[2] , \\u0_slt4_r_reg[1] , \\u0_slt4_r_reg[0] ,
    \\u0_slt5_r_reg[19] , \\u0_slt5_r_reg[18] , \\u0_slt5_r_reg[17] ,
    \\u0_slt5_r_reg[16] , \\u0_slt5_r_reg[15] , \\u0_slt5_r_reg[14] ,
    \\u0_slt5_r_reg[13] , \\u0_slt5_r_reg[12] , \\u0_slt5_r_reg[11] ,
    \\u0_slt5_r_reg[10] , \\u0_slt5_r_reg[9] , \\u0_slt5_r_reg[8] ,
    \\u0_slt5_r_reg[7] , \\u0_slt5_r_reg[6] , \\u0_slt5_r_reg[5] ,
    \\u0_slt5_r_reg[4] , \\u0_slt5_r_reg[3] , \\u0_slt5_r_reg[2] ,
    \\u0_slt5_r_reg[1] , \\u0_slt5_r_reg[0] , \\u0_slt6_r_reg[19] ,
    \\u0_slt6_r_reg[18] , \\u0_slt6_r_reg[17] , \\u0_slt6_r_reg[16] ,
    \\u0_slt6_r_reg[15] , \\u0_slt6_r_reg[14] , \\u0_slt6_r_reg[13] ,
    \\u0_slt6_r_reg[12] , \\u0_slt6_r_reg[11] , \\u0_slt6_r_reg[10] ,
    \\u0_slt6_r_reg[9] , \\u0_slt6_r_reg[8] , \\u0_slt6_r_reg[7] ,
    \\u0_slt6_r_reg[6] , \\u0_slt6_r_reg[5] , \\u0_slt6_r_reg[4] ,
    \\u0_slt6_r_reg[3] , \\u0_slt6_r_reg[2] , \\u0_slt6_r_reg[1] ,
    \\u0_slt6_r_reg[0] , \\u0_slt7_r_reg[19] , \\u0_slt7_r_reg[18] ,
    \\u0_slt7_r_reg[17] , \\u0_slt7_r_reg[16] , \\u0_slt7_r_reg[15] ,
    \\u0_slt7_r_reg[14] , \\u0_slt7_r_reg[13] , \\u0_slt7_r_reg[12] ,
    \\u0_slt7_r_reg[11] , \\u0_slt7_r_reg[10] , \\u0_slt7_r_reg[9] ,
    \\u0_slt7_r_reg[8] , \\u0_slt7_r_reg[7] , \\u0_slt7_r_reg[6] ,
    \\u0_slt7_r_reg[5] , \\u0_slt7_r_reg[4] , \\u0_slt7_r_reg[3] ,
    \\u0_slt7_r_reg[2] , \\u0_slt7_r_reg[1] , \\u0_slt7_r_reg[0] ,
    \\u0_slt8_r_reg[19] , \\u0_slt8_r_reg[18] , \\u0_slt8_r_reg[17] ,
    \\u0_slt8_r_reg[16] , \\u0_slt8_r_reg[15] , \\u0_slt8_r_reg[14] ,
    \\u0_slt8_r_reg[13] , \\u0_slt8_r_reg[12] , \\u0_slt8_r_reg[11] ,
    \\u0_slt8_r_reg[10] , \\u0_slt8_r_reg[9] , \\u0_slt8_r_reg[8] ,
    \\u0_slt8_r_reg[7] , \\u0_slt8_r_reg[6] , \\u0_slt8_r_reg[5] ,
    \\u0_slt8_r_reg[4] , \\u0_slt8_r_reg[3] , \\u0_slt8_r_reg[2] ,
    \\u0_slt8_r_reg[1] , \\u0_slt8_r_reg[0] , \\u0_slt9_r_reg[19] ,
    \\u0_slt9_r_reg[18] , \\u0_slt9_r_reg[17] , \\u0_slt9_r_reg[16] ,
    \\u0_slt9_r_reg[15] , \\u0_slt9_r_reg[14] , \\u0_slt9_r_reg[13] ,
    \\u0_slt9_r_reg[12] , \\u0_slt9_r_reg[11] , \\u0_slt9_r_reg[10] ,
    \\u0_slt9_r_reg[9] , \\u0_slt9_r_reg[8] , \\u0_slt9_r_reg[7] ,
    \\u0_slt9_r_reg[6] , \\u1_slt2_reg[19] , \\u1_slt3_reg[19] ,
    \\u1_slt4_reg[19] , \\u1_slt6_reg[19] , \\u1_slt2_reg[18] ,
    \\u1_slt3_reg[18] , \\u1_slt4_reg[18] , \\u1_slt6_reg[18] ,
    u16_u1_dma_req_reg, u16_u3_dma_req_reg, \\u0_slt9_r_reg[5] ,
    u16_u0_dma_req_reg, u16_u2_dma_req_reg, u16_u4_dma_req_reg,
    u16_u5_dma_req_reg, \\u1_slt2_reg[17] , \\u1_slt3_reg[17] ,
    \\u1_slt4_reg[17] , \\u1_slt6_reg[17] , \\u1_sr_reg[19] ,
    \\u1_slt2_reg[16] , \\u1_slt3_reg[16] , \\u1_slt4_reg[16] ,
    \\u1_slt6_reg[16] , \\u4_rp_reg[2] , \\u5_rp_reg[2] , \\u8_rp_reg[2] ,
    \\u3_rp_reg[2] , \\u6_rp_reg[2] , \\u7_rp_reg[2] , \\u8_rp_reg[3] ,
    \\u3_rp_reg[3] , \\u6_rp_reg[3] , \\u7_rp_reg[3] , \\u8_rp_reg[1] ,
    \\u3_rp_reg[1] , \\u7_rp_reg[1] , \\u6_rp_reg[1] , \\u1_sr_reg[18] ,
    \\u13_ints_r_reg[11] , \\u13_ints_r_reg[5] , \\u1_slt3_reg[15] ,
    \\u1_slt0_reg[15] , \\u1_slt6_reg[15] , \\u1_slt2_reg[15] ,
    \\u1_slt4_reg[15] , \\u4_rp_reg[1] , \\u4_rp_reg[3] , \\u5_rp_reg[1] ,
    \\u5_rp_reg[3] , \\u6_dout_reg[2] , \\u6_dout_reg[3] ,
    \\u7_dout_reg[2] , \\u7_dout_reg[3] , \\u3_dout_reg[2] ,
    \\u3_dout_reg[3] , \\u8_dout_reg[2] , \\u8_dout_reg[3] ,
    \\u13_ints_r_reg[14] , \\u13_ints_r_reg[17] , \\u13_ints_r_reg[2] ,
    \\u13_ints_r_reg[8] , \\u6_dout_reg[0] , \\u6_dout_reg[1] ,
    \\u7_dout_reg[0] , \\u7_dout_reg[1] , \\u3_dout_reg[0] ,
    \\u8_dout_reg[0] , \\u3_dout_reg[1] , \\u8_dout_reg[1] ,
    \\u8_rp_reg[0] , \\u3_rp_reg[0] , \\u6_rp_reg[0] , \\u7_rp_reg[0] ,
    \\u6_dout_reg[12] , \\u6_dout_reg[13] , \\u6_dout_reg[14] ,
    \\u6_dout_reg[15] , \\u6_dout_reg[10] , \\u6_dout_reg[11] ,
    \\u6_dout_reg[18] , \\u6_dout_reg[19] , \\u6_dout_reg[16] ,
    \\u6_dout_reg[17] , \\u6_dout_reg[4] , \\u6_dout_reg[5] ,
    \\u6_dout_reg[6] , \\u6_dout_reg[7] , \\u6_dout_reg[8] ,
    \\u6_dout_reg[9] , \\u7_dout_reg[10] , \\u7_dout_reg[11] ,
    \\u7_dout_reg[12] , \\u7_dout_reg[13] , \\u7_dout_reg[14] ,
    \\u7_dout_reg[17] , \\u7_dout_reg[15] , \\u7_dout_reg[19] ,
    \\u7_dout_reg[16] , \\u7_dout_reg[18] , \\u7_dout_reg[4] ,
    \\u7_dout_reg[5] , \\u7_dout_reg[6] , \\u7_dout_reg[7] ,
    \\u7_dout_reg[8] , \\u7_dout_reg[9] , \\u3_dout_reg[10] ,
    \\u3_dout_reg[11] , \\u3_dout_reg[13] , \\u3_dout_reg[14] ,
    \\u3_dout_reg[15] , \\u3_dout_reg[16] , \\u3_dout_reg[17] ,
    \\u3_dout_reg[18] , \\u8_dout_reg[10] , \\u3_dout_reg[19] ,
    \\u8_dout_reg[11] , \\u8_dout_reg[12] , \\u3_dout_reg[12] ,
    \\u8_dout_reg[13] , \\u8_dout_reg[14] , \\u3_dout_reg[4] ,
    \\u8_dout_reg[16] , \\u3_dout_reg[6] , \\u8_dout_reg[17] ,
    \\u3_dout_reg[7] , \\u8_dout_reg[18] , \\u3_dout_reg[8] ,
    \\u8_dout_reg[15] , \\u3_dout_reg[5] , \\u8_dout_reg[19] ,
    \\u3_dout_reg[9] , \\u8_dout_reg[4] , \\u8_dout_reg[5] ,
    \\u8_dout_reg[6] , \\u8_dout_reg[7] , \\u8_dout_reg[8] ,
    \\u8_dout_reg[9] , \\u0_slt9_r_reg[4] , u16_u1_dma_req_r1_reg,
    u16_u3_dma_req_r1_reg, \\u1_sr_reg[17] , u16_u8_dma_req_reg,
    \\u1_slt3_reg[14] , \\u1_slt4_reg[14] , \\u1_slt6_reg[14] ,
    \\u1_slt2_reg[14] , \\u4_dout_reg[3] , \\u5_dout_reg[3] ,
    \\u5_dout_reg[2] , \\u4_dout_reg[2] , u16_u0_dma_req_r1_reg,
    u16_u2_dma_req_r1_reg, u16_u4_dma_req_r1_reg, u16_u5_dma_req_r1_reg,
    \\u4_dout_reg[4] , \\u11_wp_reg[3] , u16_u6_dma_req_reg,
    u16_u7_dma_req_reg, \\u5_dout_reg[0] , \\u5_dout_reg[1] ,
    \\u4_dout_reg[1] , \\u4_dout_reg[0] , \\u4_rp_reg[0] , \\u5_rp_reg[0] ,
    \\u11_mem_reg[0][18] , \\u11_mem_reg[0][19] , \\u11_mem_reg[1][18] ,
    \\u11_mem_reg[1][19] , \\u11_mem_reg[1][20] , \\u11_mem_reg[1][21] ,
    \\u11_mem_reg[1][22] , \\u11_mem_reg[1][23] , \\u11_mem_reg[1][24] ,
    \\u11_mem_reg[1][25] , \\u11_mem_reg[1][26] , \\u11_mem_reg[1][27] ,
    \\u11_mem_reg[1][28] , \\u11_mem_reg[1][29] , \\u11_mem_reg[1][30] ,
    \\u11_mem_reg[1][31] , \\u11_mem_reg[2][18] , \\u11_mem_reg[2][19] ,
    \\u11_mem_reg[2][20] , \\u11_mem_reg[2][21] , \\u11_mem_reg[2][22] ,
    \\u11_mem_reg[2][23] , \\u11_mem_reg[2][24] , \\u11_mem_reg[2][25] ,
    \\u11_mem_reg[2][26] , \\u11_mem_reg[2][27] , \\u11_mem_reg[2][28] ,
    \\u11_mem_reg[2][29] , \\u11_mem_reg[2][30] , \\u11_mem_reg[2][31] ,
    \\u11_mem_reg[3][18] , \\u11_mem_reg[3][19] , \\u11_mem_reg[3][20] ,
    \\u11_mem_reg[3][21] , \\u11_mem_reg[3][22] , \\u11_mem_reg[3][23] ,
    \\u11_mem_reg[3][24] , \\u11_mem_reg[3][25] , \\u11_mem_reg[3][26] ,
    \\u11_mem_reg[3][27] , \\u11_mem_reg[3][28] , \\u11_mem_reg[3][29] ,
    \\u11_mem_reg[3][30] , \\u11_mem_reg[3][31] , \\u11_mem_reg[3][7] ,
    \\u11_mem_reg[1][12] , \\u11_mem_reg[1][13] , \\u11_mem_reg[1][16] ,
    \\u11_mem_reg[2][17] , \\u11_mem_reg[2][1] , \\u11_mem_reg[2][7] ,
    \\u11_mem_reg[2][8] , \\u11_mem_reg[3][16] , \\u11_mem_reg[3][17] ,
    \\u11_mem_reg[3][5] , \\u11_mem_reg[3][6] , \\u11_wp_reg[1] ,
    \\u11_wp_reg[2] , \\u4_dout_reg[10] , \\u4_dout_reg[13] ,
    \\u4_dout_reg[14] , \\u4_dout_reg[15] , \\u4_dout_reg[16] ,
    \\u4_dout_reg[11] , \\u4_dout_reg[18] , \\u4_dout_reg[12] ,
    \\u4_dout_reg[19] , \\u4_dout_reg[17] , \\u4_dout_reg[5] ,
    \\u4_dout_reg[6] , \\u4_dout_reg[7] , \\u4_dout_reg[8] ,
    \\u4_dout_reg[9] , \\u5_dout_reg[10] , \\u5_dout_reg[11] ,
    \\u5_dout_reg[12] , \\u5_dout_reg[14] , \\u5_dout_reg[15] ,
    \\u5_dout_reg[16] , \\u5_dout_reg[18] , \\u5_dout_reg[19] ,
    \\u5_dout_reg[4] , \\u5_dout_reg[5] , \\u5_dout_reg[6] ,
    \\u5_dout_reg[8] , \\u5_dout_reg[9] , \\u11_mem_reg[0][0] ,
    \\u11_mem_reg[0][10] , \\u11_mem_reg[0][11] , \\u11_mem_reg[0][12] ,
    \\u11_mem_reg[0][13] , \\u11_mem_reg[0][14] , \\u11_mem_reg[0][15] ,
    \\u11_mem_reg[0][1] , u15_crac_rd_reg, \\u17_int_set_reg[1] ,
    \\u20_int_set_reg[1] , \\u21_int_set_reg[1] , \\u22_int_set_reg[1] ,
    \\u5_dout_reg[7] , \\u5_dout_reg[17] , \\u1_sr_reg[16] ,
    \\u5_dout_reg[13] , \\u10_mem_reg[0][18] , \\u10_mem_reg[3][28] ,
    \\u10_mem_reg[3][24] , \\u9_mem_reg[3][30] , \\u9_mem_reg[3][26] ,
    \\u10_wp_reg[3] , \\u9_mem_reg[3][22] , \\u9_mem_reg[2][28] ,
    \\u9_mem_reg[2][24] , \\u9_mem_reg[2][20] , \\u9_mem_reg[1][28] ,
    \\u9_mem_reg[1][25] , \\u9_mem_reg[1][22] , \\u10_mem_reg[2][24] ,
    \\u11_mem_reg[3][14] , \\u11_mem_reg[3][0] , \\u11_mem_reg[3][13] ,
    \\u10_mem_reg[1][0] , \\u11_mem_reg[1][15] , \\u11_mem_reg[1][6] ,
    \\u1_slt2_reg[13] , \\u1_slt4_reg[13] , \\u1_slt6_reg[13] ,
    \\u1_slt3_reg[13] , \\u10_mem_reg[2][18] , \\u10_mem_reg[2][19] ,
    \\u10_mem_reg[2][20] , \\u10_mem_reg[2][21] , \\u10_mem_reg[2][22] ,
    \\u9_mem_reg[0][18] , \\u9_mem_reg[0][19] , \\u10_mem_reg[2][23] ,
    \\u10_mem_reg[2][25] , \\u10_mem_reg[2][26] , \\u10_mem_reg[2][27] ,
    \\u9_mem_reg[1][18] , \\u9_mem_reg[1][19] , \\u9_mem_reg[1][20] ,
    \\u9_mem_reg[1][21] , \\u10_mem_reg[2][28] , \\u9_mem_reg[1][23] ,
    \\u9_mem_reg[1][24] , \\u9_mem_reg[1][26] , \\u10_mem_reg[2][29] ,
    \\u9_mem_reg[1][27] , \\u9_mem_reg[1][29] , \\u9_mem_reg[1][30] ,
    \\u9_mem_reg[1][31] , \\u10_mem_reg[2][30] , \\u9_mem_reg[2][18] ,
    \\u9_mem_reg[2][19] , \\u10_mem_reg[2][31] , \\u9_mem_reg[2][21] ,
    \\u9_mem_reg[2][22] , \\u9_mem_reg[2][23] , \\u9_mem_reg[2][25] ,
    \\u9_mem_reg[2][26] , \\u9_mem_reg[2][27] , \\u9_mem_reg[2][29] ,
    \\u9_mem_reg[2][30] , \\u9_mem_reg[2][31] , \\u9_mem_reg[3][18] ,
    \\u9_mem_reg[3][19] , \\u9_mem_reg[3][20] , \\u9_mem_reg[3][21] ,
    \\u9_mem_reg[3][23] , \\u9_mem_reg[3][24] , \\u9_mem_reg[3][25] ,
    \\u9_mem_reg[3][27] , \\u9_mem_reg[3][28] , \\u9_mem_reg[3][29] ,
    \\u9_mem_reg[3][31] , \\u10_mem_reg[3][18] , \\u10_mem_reg[3][19] ,
    \\u10_mem_reg[3][20] , \\u10_mem_reg[3][21] , \\u10_mem_reg[3][22] ,
    \\u10_mem_reg[3][23] , \\u10_mem_reg[3][25] , \\u10_mem_reg[3][26] ,
    \\u10_mem_reg[3][27] , \\u10_mem_reg[3][29] , \\u10_mem_reg[3][30] ,
    \\u10_mem_reg[3][31] , \\u10_mem_reg[0][19] , \\u10_mem_reg[1][18] ,
    \\u10_mem_reg[1][19] , \\u10_mem_reg[1][21] , \\u10_mem_reg[1][22] ,
    \\u10_mem_reg[1][23] , \\u10_mem_reg[1][24] , \\u10_mem_reg[1][25] ,
    \\u10_mem_reg[1][26] , \\u10_mem_reg[1][27] , \\u10_mem_reg[1][28] ,
    \\u10_mem_reg[1][29] , \\u10_mem_reg[1][20] , \\u10_mem_reg[1][30] ,
    \\u10_mem_reg[1][31] , \\u11_mem_reg[3][8] , \\u11_mem_reg[3][9] ,
    \\u10_mem_reg[2][1] , \\u10_mem_reg[2][5] , \\u10_mem_reg[2][6] ,
    \\u10_mem_reg[3][3] , \\u10_mem_reg[2][9] , \\u11_mem_reg[1][0] ,
    \\u11_mem_reg[1][10] , \\u11_mem_reg[1][11] , \\u10_mem_reg[3][2] ,
    \\u10_mem_reg[3][9] , \\u11_mem_reg[1][14] , \\u11_mem_reg[1][1] ,
    \\u11_mem_reg[1][2] , \\u11_mem_reg[1][3] , \\u11_mem_reg[1][4] ,
    \\u11_mem_reg[1][5] , \\u11_mem_reg[1][7] , \\u11_mem_reg[1][8] ,
    \\u11_mem_reg[1][9] , \\u11_mem_reg[2][0] , \\u11_mem_reg[2][10] ,
    \\u11_mem_reg[2][11] , \\u11_mem_reg[2][13] , \\u11_mem_reg[2][14] ,
    \\u11_mem_reg[2][15] , \\u11_mem_reg[2][16] , \\u11_mem_reg[1][17] ,
    \\u11_mem_reg[2][12] , \\u11_mem_reg[2][2] , \\u11_mem_reg[2][3] ,
    \\u11_mem_reg[2][6] , \\u11_mem_reg[2][4] , \\u11_mem_reg[2][5] ,
    \\u11_mem_reg[2][9] , \\u11_mem_reg[3][11] , \\u11_mem_reg[3][12] ,
    \\u11_mem_reg[3][15] , \\u11_mem_reg[3][10] , \\u11_mem_reg[3][2] ,
    \\u11_mem_reg[3][3] , \\u11_mem_reg[3][4] , \\u11_mem_reg[3][1] ,
    \\u10_wp_reg[1] , \\u10_wp_reg[2] , \\u10_mem_reg[0][2] ,
    \\u11_mem_reg[0][5] , \\u10_mem_reg[0][13] , \\u10_mem_reg[0][12] ,
    \\u11_mem_reg[0][16] , \\u11_mem_reg[0][20] , \\u11_mem_reg[0][21] ,
    \\u11_mem_reg[0][22] , \\u11_mem_reg[0][23] , \\u11_mem_reg[0][24] ,
    \\u11_mem_reg[0][25] , \\u10_mem_reg[0][21] , \\u11_mem_reg[0][26] ,
    \\u11_mem_reg[0][27] , \\u10_mem_reg[0][22] , \\u11_mem_reg[0][28] ,
    \\u11_mem_reg[0][29] , \\u11_mem_reg[0][2] , \\u11_mem_reg[0][30] ,
    \\u11_mem_reg[0][31] , \\u11_mem_reg[0][3] , \\u10_mem_reg[0][25] ,
    \\u11_mem_reg[0][4] , \\u10_mem_reg[0][26] , \\u10_mem_reg[0][27] ,
    \\u11_mem_reg[0][6] , \\u10_mem_reg[0][28] , \\u11_mem_reg[0][7] ,
    \\u11_mem_reg[0][8] , \\u10_mem_reg[0][29] , \\u11_mem_reg[0][9] ,
    \\u10_mem_reg[0][5] , \\u11_wp_reg[0] , \\u25_int_set_reg[2] ,
    \\u10_mem_reg[0][1] , \\u11_mem_reg[0][17] , \\u10_mem_reg[3][17] ,
    \\u1_sr_reg[15] , \\u10_mem_reg[0][11] , \\u9_mem_reg[0][4] ,
    \\u9_wp_reg[3] , \\u9_mem_reg[0][8] , \\u10_mem_reg[1][8] ,
    \\u9_mem_reg[0][2] , \\u9_mem_reg[0][26] , \\u10_mem_reg[1][6] ,
    \\u9_mem_reg[0][17] , \\u9_mem_reg[0][13] , \\u10_mem_reg[1][1] ,
    \\u10_mem_reg[1][15] , \\u10_mem_reg[1][13] , \\u10_mem_reg[1][10] ,
    \\u10_mem_reg[3][8] , \\u10_mem_reg[0][23] , \\u11_din_tmp1_reg[8] ,
    \\u9_mem_reg[2][12] , \\u10_mem_reg[3][13] , \\u10_mem_reg[3][0] ,
    \\u9_mem_reg[3][4] , \\u9_mem_reg[3][1] , \\u9_mem_reg[3][15] ,
    \\u9_mem_reg[2][5] , \\u9_mem_reg[2][2] , \\u10_mem_reg[1][9] ,
    \\u10_mem_reg[2][0] , \\u10_mem_reg[2][11] , \\u10_mem_reg[2][12] ,
    \\u10_mem_reg[2][13] , \\u10_mem_reg[2][14] , \\u10_mem_reg[2][15] ,
    \\u10_mem_reg[2][16] , \\u10_mem_reg[2][10] , \\u9_mem_reg[1][0] ,
    \\u9_mem_reg[1][10] , \\u9_mem_reg[1][12] , \\u9_mem_reg[1][13] ,
    \\u9_mem_reg[1][14] , \\u9_mem_reg[1][16] , \\u9_mem_reg[1][17] ,
    \\u9_mem_reg[1][1] , \\u9_mem_reg[1][2] , \\u9_mem_reg[1][3] ,
    \\u9_mem_reg[1][4] , \\u9_mem_reg[1][5] , \\u9_mem_reg[1][6] ,
    \\u9_mem_reg[1][7] , \\u9_mem_reg[1][8] , \\u9_mem_reg[2][0] ,
    \\u9_mem_reg[2][10] , \\u9_mem_reg[2][11] , \\u9_mem_reg[2][14] ,
    \\u9_mem_reg[2][15] , \\u9_mem_reg[2][16] , \\u9_mem_reg[2][17] ,
    \\u9_mem_reg[2][1] , \\u10_mem_reg[2][3] , \\u9_mem_reg[2][3] ,
    \\u10_mem_reg[2][4] , \\u9_mem_reg[2][4] , \\u9_mem_reg[2][6] ,
    \\u9_mem_reg[2][7] , \\u9_mem_reg[2][8] , \\u9_mem_reg[3][0] ,
    \\u9_mem_reg[3][10] , \\u9_mem_reg[3][11] , \\u9_mem_reg[3][12] ,
    \\u9_mem_reg[3][13] , \\u9_mem_reg[3][14] , \\u9_mem_reg[2][13] ,
    \\u9_mem_reg[3][16] , \\u9_mem_reg[3][17] , \\u10_mem_reg[2][7] ,
    \\u9_mem_reg[3][2] , \\u9_mem_reg[3][3] , \\u9_mem_reg[3][5] ,
    \\u9_mem_reg[3][6] , \\u9_mem_reg[3][7] , \\u10_mem_reg[2][8] ,
    \\u9_mem_reg[3][9] , \\u9_mem_reg[3][8] , \\u10_mem_reg[3][10] ,
    \\u10_mem_reg[3][11] , \\u10_mem_reg[3][12] , \\u10_mem_reg[3][14] ,
    \\u10_mem_reg[3][15] , \\u10_mem_reg[3][16] , \\u10_mem_reg[3][1] ,
    \\u10_mem_reg[3][4] , \\u10_mem_reg[3][5] , \\u10_mem_reg[3][6] ,
    \\u10_mem_reg[3][7] , \\u10_mem_reg[1][11] , \\u10_mem_reg[1][12] ,
    \\u10_mem_reg[1][14] , \\u10_mem_reg[1][17] , \\u10_mem_reg[1][16] ,
    \\u9_mem_reg[1][9] , \\u10_mem_reg[1][3] , \\u10_mem_reg[1][4] ,
    \\u10_mem_reg[1][5] , \\u10_mem_reg[1][2] , \\u10_mem_reg[2][2] ,
    \\u10_mem_reg[1][7] , \\u9_wp_reg[2] , \\u9_mem_reg[1][15] ,
    \\u9_mem_reg[1][11] , \\u10_mem_reg[2][17] , \\u10_mem_reg[0][24] ,
    \\u11_din_tmp1_reg[4] , \\u10_mem_reg[0][8] , \\u10_mem_reg[0][4] ,
    \\u9_mem_reg[0][0] , \\u9_mem_reg[0][10] , \\u9_mem_reg[0][11] ,
    \\u9_mem_reg[0][12] , \\u9_mem_reg[0][14] , \\u9_mem_reg[0][15] ,
    \\u9_mem_reg[0][16] , \\u9_mem_reg[0][1] , \\u9_mem_reg[0][20] ,
    \\u9_mem_reg[0][21] , \\u9_mem_reg[0][22] , \\u9_mem_reg[0][23] ,
    \\u9_mem_reg[0][24] , \\u9_mem_reg[0][25] , \\u9_mem_reg[0][27] ,
    \\u9_mem_reg[0][28] , \\u9_mem_reg[0][29] , \\u9_mem_reg[0][30] ,
    \\u9_mem_reg[0][31] , \\u9_mem_reg[0][3] , \\u9_mem_reg[0][5] ,
    \\u9_mem_reg[0][6] , \\u9_mem_reg[0][7] , \\u9_mem_reg[0][9] ,
    \\u10_mem_reg[0][0] , \\u10_mem_reg[0][10] , \\u10_mem_reg[0][14] ,
    \\u10_mem_reg[0][15] , \\u10_mem_reg[0][16] , \\u10_mem_reg[0][17] ,
    \\u10_mem_reg[0][31] , \\u10_mem_reg[0][3] , \\u10_mem_reg[0][30] ,
    \\u10_mem_reg[0][6] , \\u10_mem_reg[0][7] , \\u10_mem_reg[0][9] ,
    \\u10_wp_reg[0] , \\u11_din_tmp1_reg[0] , \\u11_din_tmp1_reg[10] ,
    \\u11_din_tmp1_reg[11] , \\u11_din_tmp1_reg[12] ,
    \\u11_din_tmp1_reg[13] , \\u11_din_tmp1_reg[14] ,
    \\u11_din_tmp1_reg[15] , \\u11_din_tmp1_reg[1] ,
    \\u11_din_tmp1_reg[2] , \\u11_din_tmp1_reg[3] , \\u11_din_tmp1_reg[5] ,
    \\u11_din_tmp1_reg[6] , \\u11_din_tmp1_reg[7] , \\u11_din_tmp1_reg[9] ,
    \\u9_mem_reg[2][9] , \\u18_int_set_reg[1] , \\u19_int_set_reg[1] ,
    \\u24_int_set_reg[2] , u15_crac_wr_reg, \\u13_ints_r_reg[1] ,
    \\u10_mem_reg[0][20] , \\u0_slt9_r_reg[3] , \\u10_din_tmp1_reg[13] ,
    \\u1_slt6_reg[12] , \\u13_ints_r_reg[26] , \\u1_slt0_reg[12] ,
    \\u1_slt2_reg[12] , \\u1_slt3_reg[12] , \\u1_slt4_reg[12] ,
    \\u10_din_tmp1_reg[11] , \\u9_wp_reg[0] , \\u10_din_tmp1_reg[5] ,
    \\u10_din_tmp1_reg[3] , \\u10_din_tmp1_reg[1] , \\u10_din_tmp1_reg[2] ,
    \\u10_din_tmp1_reg[4] , \\u10_din_tmp1_reg[6] , \\u10_din_tmp1_reg[8] ,
    \\u10_din_tmp1_reg[9] , \\u10_din_tmp1_reg[7] , \\u10_din_tmp1_reg[0] ,
    \\u10_din_tmp1_reg[10] , \\u10_din_tmp1_reg[15] ,
    \\u10_din_tmp1_reg[14] , \\u10_din_tmp1_reg[12] , u15_rdd1_reg,
    u15_rdd2_reg, \\u20_int_set_reg[0] , \\u18_int_set_reg[0] ,
    \\u1_sr_reg[14] , \\u13_ints_r_reg[23] , \\u13_ints_r_reg[20] ,
    \\u9_wp_reg[1] , \\u9_din_tmp1_reg[9] , \\u9_din_tmp1_reg[3] ,
    \\u9_din_tmp1_reg[10] , \\u9_din_tmp1_reg[14] , \\u9_din_tmp1_reg[0] ,
    \\u9_din_tmp1_reg[11] , \\u9_din_tmp1_reg[12] , \\u9_din_tmp1_reg[13] ,
    \\u9_din_tmp1_reg[15] , \\u9_din_tmp1_reg[1] , \\u9_din_tmp1_reg[2] ,
    \\u9_din_tmp1_reg[5] , \\u9_din_tmp1_reg[6] , \\u9_din_tmp1_reg[4] ,
    \\u9_din_tmp1_reg[8] , \\u9_din_tmp1_reg[7] , u15_rdd3_reg,
    \\u21_int_set_reg[0] , \\u22_int_set_reg[0] , \\u17_int_set_reg[0] ,
    \\u19_int_set_reg[0] , u16_u8_dma_req_r1_reg, \\u1_slt4_reg[11] ,
    \\u1_slt0_reg[11] , \\u1_slt1_reg[11] , \\u1_slt2_reg[11] ,
    \\u1_slt3_reg[11] , \\u1_slt6_reg[11] , \\u23_int_set_reg[2] ,
    u15_crac_rd_done_reg, u16_u6_dma_req_r1_reg, u16_u7_dma_req_r1_reg,
    \\u1_sr_reg[13] , \\u1_slt6_reg[10] , \\u1_slt2_reg[10] ,
    u14_u4_en_out_l_reg, u2_sync_resume_reg, \\u1_slt1_reg[10] ,
    \\u1_slt4_reg[10] , \\u1_slt3_reg[10] , u14_u0_en_out_l_reg,
    u14_u1_en_out_l_reg, u14_u2_en_out_l_reg, u14_u3_en_out_l_reg,
    u14_u5_en_out_l_reg, u14_crac_valid_r_reg, \\u0_slt9_r_reg[2] ,
    \\u1_sr_reg[12] , \\u26_ps_cnt_reg[5] , \\u26_ps_cnt_reg[2] ,
    \\u26_ps_cnt_reg[0] , \\u26_ps_cnt_reg[1] , \\u26_ps_cnt_reg[4] ,
    \\u26_ps_cnt_reg[3] , \\u12_wb_data_o_reg[1] , \\u17_int_set_reg[2] ,
    \\u18_int_set_reg[2] , \\u21_int_set_reg[2] , \\u20_int_set_reg[2] ,
    u14_crac_wr_r_reg, \\u22_int_set_reg[2] , \\u19_int_set_reg[2] ,
    \\u1_slt2_reg[9] , u14_u3_full_empty_r_reg, \\u25_int_set_reg[0] ,
    u14_u0_full_empty_r_reg, u14_u1_full_empty_r_reg,
    u14_u2_full_empty_r_reg, u14_u5_full_empty_r_reg, \\u1_slt0_reg[9] ,
    u14_u4_full_empty_r_reg, \\u1_slt4_reg[9] , \\u1_slt3_reg[9] ,
    \\u8_wp_reg[0] , \\u3_wp_reg[0] , \\u4_wp_reg[0] , \\u5_wp_reg[0] ,
    \\u6_wp_reg[0] , \\u7_wp_reg[0] , \\u1_slt6_reg[9] , u26_ac97_rst__reg,
    \\u1_sr_reg[11] , \\u26_cnt_reg[2] , \\u23_int_set_reg[0] ,
    \\u24_int_set_reg[0] , u14_u8_en_out_l_reg, \\u5_wp_reg[1] ,
    \\u6_wp_reg[2] , \\u26_cnt_reg[0] , \\u26_cnt_reg[1] , \\u8_wp_reg[2] ,
    \\u3_wp_reg[2] , \\u5_wp_reg[2] , \\u7_wp_reg[2] , u14_u6_en_out_l_reg,
    u14_u7_en_out_l_reg, \\u8_wp_reg[1] , \\u3_wp_reg[1] , \\u4_wp_reg[1] ,
    \\u6_wp_reg[1] , \\u7_wp_reg[1] , \\u4_wp_reg[2] , u15_valid_r_reg,
    \\u1_slt6_reg[8] , \\u1_slt2_reg[8] , \\u1_slt1_reg[8] ,
    \\u1_slt4_reg[8] , \\u1_slt3_reg[8] , \\u4_mem_reg[0][13] ,
    \\u4_mem_reg[0][14] , \\u4_mem_reg[0][16] , \\u4_mem_reg[0][19] ,
    \\u4_mem_reg[0][22] , \\u4_mem_reg[0][24] , \\u4_mem_reg[0][31] ,
    \\u4_mem_reg[0][4] , \\u4_mem_reg[0][7] , \\u4_mem_reg[0][9] ,
    \\u5_mem_reg[0][13] , \\u5_mem_reg[0][14] , \\u5_mem_reg[0][16] ,
    \\u5_mem_reg[0][19] , \\u5_mem_reg[0][22] , \\u5_mem_reg[0][24] ,
    \\u5_mem_reg[0][31] , \\u5_mem_reg[0][4] , \\u5_mem_reg[0][7] ,
    \\u5_mem_reg[0][9] , \\u6_mem_reg[0][13] , \\u6_mem_reg[0][14] ,
    \\u6_mem_reg[0][16] , \\u6_mem_reg[0][19] , \\u6_mem_reg[0][22] ,
    \\u6_mem_reg[0][24] , \\u6_mem_reg[0][31] , \\u6_mem_reg[0][4] ,
    \\u6_mem_reg[0][7] , \\u6_mem_reg[0][9] , \\u7_mem_reg[0][13] ,
    \\u7_mem_reg[0][14] , \\u7_mem_reg[0][16] , \\u7_mem_reg[0][19] ,
    \\u7_mem_reg[0][22] , \\u7_mem_reg[0][24] , \\u7_mem_reg[0][31] ,
    \\u7_mem_reg[0][4] , \\u7_mem_reg[0][7] , \\u7_mem_reg[0][9] ,
    \\u3_mem_reg[0][11] , \\u3_mem_reg[0][12] , \\u3_mem_reg[0][15] ,
    \\u8_mem_reg[0][0] , \\u8_mem_reg[0][11] , \\u8_mem_reg[0][12] ,
    \\u8_mem_reg[0][17] , \\u3_mem_reg[0][1] , \\u3_mem_reg[0][21] ,
    \\u8_mem_reg[0][26] , \\u8_mem_reg[0][28] , \\u8_mem_reg[0][29] ,
    \\u8_mem_reg[0][30] , \\u3_mem_reg[0][27] , \\u8_mem_reg[0][4] ,
    \\u8_mem_reg[0][5] , \\u3_mem_reg[0][2] , \\u3_mem_reg[0][29] ,
    \\u3_mem_reg[0][6] , \\u3_mem_reg[0][5] , \\u13_crac_r_reg[6] ,
    \\u3_mem_reg[0][17] , \\u8_mem_reg[2][18] , \\u7_mem_reg[0][20] ,
    \\u8_mem_reg[2][25] , \\u8_mem_reg[2][28] , \\u4_mem_reg[2][16] ,
    \\u5_mem_reg[1][26] , \\u13_occ0_r_reg[11] , \\u5_mem_reg[1][22] ,
    \\u5_mem_reg[1][15] , \\u5_mem_reg[1][19] , \\u5_mem_reg[1][11] ,
    \\u3_mem_reg[1][22] , \\u8_mem_reg[2][20] , \\u4_mem_reg[3][9] ,
    \\u4_mem_reg[3][5] , \\u4_mem_reg[3][30] , \\u8_mem_reg[0][15] ,
    \\u3_mem_reg[0][16] , \\u4_mem_reg[3][23] , \\u4_mem_reg[3][27] ,
    \\u8_mem_reg[1][6] , \\u13_occ0_r_reg[8] , \\u13_icc_r_reg[8] ,
    \\u8_mem_reg[2][13] , \\u3_mem_reg[1][19] , \\u4_mem_reg[2][9] ,
    \\u4_mem_reg[3][16] , \\u4_mem_reg[3][12] , \\u4_mem_reg[2][5] ,
    \\u3_mem_reg[1][15] , \\u4_mem_reg[2][30] , \\u4_mem_reg[2][27] ,
    \\u4_mem_reg[2][23] , \\u7_mem_reg[0][30] , \\u3_mem_reg[2][2] ,
    \\u8_mem_reg[1][21] , \\u3_mem_reg[1][11] , \\u8_mem_reg[1][3] ,
    \\u4_mem_reg[2][12] , \\u4_mem_reg[1][30] , \\u4_mem_reg[1][9] ,
    \\u4_mem_reg[1][5] , \\u4_mem_reg[1][27] , \\u8_mem_reg[1][28] ,
    \\u3_mem_reg[0][13] , \\u8_mem_reg[1][25] , \\u4_mem_reg[1][23] ,
    \\u4_mem_reg[1][16] , \\u7_mem_reg[0][6] , \\u7_mem_reg[1][25] ,
    \\u3_mem_reg[3][3] , \\u4_mem_reg[1][12] , \\u7_mem_reg[3][3] ,
    \\u8_mem_reg[1][14] , \\u8_mem_reg[1][18] , \\u3_mem_reg[3][6] ,
    \\u3_mem_reg[3][22] , \\u3_mem_reg[3][30] , \\u3_mem_reg[3][27] ,
    \\u7_mem_reg[0][23] , \\u3_mem_reg[3][19] , u14_u0_en_out_l2_reg,
    u14_u1_en_out_l2_reg, u14_u2_en_out_l2_reg, u14_u3_en_out_l2_reg,
    u14_u4_en_out_l2_reg, u14_u5_en_out_l2_reg, \\u6_mem_reg[0][12] ,
    \\u8_mem_reg[1][10] , \\u7_mem_reg[3][7] , \\u3_mem_reg[3][15] ,
    \\u3_mem_reg[3][11] , \\u3_mem_reg[2][8] , \\u7_mem_reg[0][12] ,
    \\u7_mem_reg[3][14] , \\u7_mem_reg[3][25] , \\u7_mem_reg[3][29] ,
    \\u3_mem_reg[2][26] , \\u3_mem_reg[2][22] , \\u3_mem_reg[2][18] ,
    \\u8_mem_reg[3][8] , \\u8_mem_reg[3][6] , \\u7_mem_reg[3][21] ,
    \\u7_mem_reg[3][18] , \\u8_mem_reg[3][3] , \\u3_mem_reg[2][11] ,
    \\u8_mem_reg[3][28] , \\u7_mem_reg[0][17] , \\u7_mem_reg[0][0] ,
    \\u8_mem_reg[3][22] , \\u8_mem_reg[3][25] , \\u7_mem_reg[2][25] ,
    \\u7_mem_reg[2][7] , \\u7_mem_reg[3][10] , \\u8_mem_reg[3][18] ,
    \\u3_mem_reg[1][3] , \\u8_mem_reg[3][15] , \\u8_mem_reg[3][10] ,
    \\u7_mem_reg[2][3] , \\u7_mem_reg[2][29] , \\u3_mem_reg[1][2] ,
    \\u7_mem_reg[2][21] , \\u7_mem_reg[2][18] , \\u6_mem_reg[0][30] ,
    \\u6_mem_reg[0][6] , \\u7_mem_reg[2][14] , \\u7_mem_reg[2][10] ,
    \\u8_mem_reg[2][6] , \\u6_mem_reg[0][28] , \\u7_mem_reg[1][7] ,
    \\u6_mem_reg[3][8] , \\u13_crac_dout_r_reg[3] ,
    \\u13_crac_dout_r_reg[9] , \\u7_mem_reg[1][3] , \\u13_icc_r_reg[22] ,
    \\u13_crac_dout_r_reg[14] , \\u13_occ0_r_reg[2] , \\u13_occ0_r_reg[4] ,
    \\u13_intm_r_reg[7] , \\u13_intm_r_reg[22] , \\u13_icc_r_reg[11] ,
    \\u7_mem_reg[1][29] , \\u6_mem_reg[0][23] , \\u13_icc_r_reg[15] ,
    \\u13_icc_r_reg[19] , \\u13_crac_r_reg[0] , \\u13_crac_r_reg[1] ,
    \\u13_crac_r_reg[3] , \\u13_crac_r_reg[4] , \\u13_crac_r_reg[5] ,
    \\u13_crac_r_reg[7] , \\u13_icc_r_reg[0] , \\u13_icc_r_reg[10] ,
    \\u13_icc_r_reg[12] , \\u13_icc_r_reg[13] , \\u13_icc_r_reg[14] ,
    \\u13_icc_r_reg[16] , \\u13_icc_r_reg[17] , \\u13_icc_r_reg[18] ,
    \\u13_icc_r_reg[1] , \\u13_icc_r_reg[20] , \\u13_icc_r_reg[21] ,
    \\u13_icc_r_reg[23] , \\u13_icc_r_reg[2] , \\u13_icc_r_reg[3] ,
    \\u13_icc_r_reg[4] , \\u13_icc_r_reg[5] , \\u13_icc_r_reg[6] ,
    \\u13_icc_r_reg[7] , \\u13_icc_r_reg[9] , \\u13_occ0_r_reg[0] ,
    \\u13_occ0_r_reg[10] , \\u13_occ0_r_reg[12] , \\u13_occ0_r_reg[13] ,
    \\u13_occ0_r_reg[14] , \\u13_occ0_r_reg[16] , \\u13_occ0_r_reg[17] ,
    \\u13_occ0_r_reg[18] , \\u13_occ0_r_reg[1] , \\u13_occ0_r_reg[20] ,
    \\u13_occ0_r_reg[21] , \\u13_occ0_r_reg[23] , \\u13_occ0_r_reg[24] ,
    \\u13_occ0_r_reg[25] , \\u13_occ0_r_reg[27] , \\u13_occ0_r_reg[28] ,
    \\u13_occ0_r_reg[29] , \\u13_occ0_r_reg[30] , \\u13_occ0_r_reg[31] ,
    \\u13_occ0_r_reg[3] , \\u13_occ0_r_reg[5] , \\u13_occ0_r_reg[6] ,
    \\u13_occ0_r_reg[7] , \\u13_occ0_r_reg[9] , \\u13_intm_r_reg[0] ,
    \\u13_intm_r_reg[10] , \\u13_intm_r_reg[11] , \\u13_intm_r_reg[12] ,
    \\u13_intm_r_reg[13] , \\u13_intm_r_reg[14] , \\u13_intm_r_reg[16] ,
    \\u13_intm_r_reg[17] , \\u13_intm_r_reg[18] , \\u13_intm_r_reg[19] ,
    \\u13_intm_r_reg[1] , \\u13_intm_r_reg[20] , \\u13_intm_r_reg[21] ,
    \\u13_intm_r_reg[23] , \\u13_intm_r_reg[24] , \\u13_intm_r_reg[25] ,
    \\u13_intm_r_reg[27] , \\u13_intm_r_reg[28] , \\u13_intm_r_reg[2] ,
    \\u13_intm_r_reg[5] , \\u13_intm_r_reg[6] , \\u13_intm_r_reg[9] ,
    \\u13_intm_r_reg[4] , \\u13_intm_r_reg[15] , \\u13_crac_dout_r_reg[0] ,
    \\u13_crac_dout_r_reg[10] , \\u13_crac_dout_r_reg[11] ,
    \\u13_crac_dout_r_reg[12] , \\u13_crac_dout_r_reg[13] ,
    \\u13_crac_dout_r_reg[15] , \\u13_crac_dout_r_reg[1] ,
    \\u13_crac_dout_r_reg[2] , \\u13_crac_dout_r_reg[4] ,
    \\u13_crac_dout_r_reg[5] , \\u13_crac_dout_r_reg[6] ,
    \\u13_crac_dout_r_reg[8] , \\u8_mem_reg[2][4] , \\u3_mem_reg[1][28] ,
    \\u8_mem_reg[2][5] , \\u3_mem_reg[1][29] , \\u8_mem_reg[2][7] ,
    \\u8_mem_reg[2][8] , \\u8_mem_reg[2][9] , \\u8_mem_reg[3][0] ,
    \\u3_mem_reg[1][30] , \\u8_mem_reg[3][11] , \\u3_mem_reg[1][31] ,
    \\u8_mem_reg[3][12] , \\u8_mem_reg[3][13] , \\u3_mem_reg[1][4] ,
    \\u8_mem_reg[3][14] , \\u8_mem_reg[3][16] , \\u8_mem_reg[3][17] ,
    \\u3_mem_reg[1][5] , \\u8_mem_reg[3][19] , \\u3_mem_reg[1][6] ,
    \\u8_mem_reg[3][1] , \\u3_mem_reg[1][7] , \\u8_mem_reg[3][20] ,
    \\u8_mem_reg[3][21] , \\u3_mem_reg[1][8] , \\u8_mem_reg[3][23] ,
    \\u8_mem_reg[3][24] , \\u3_mem_reg[1][9] , \\u8_mem_reg[3][26] ,
    \\u3_mem_reg[2][0] , \\u8_mem_reg[3][27] , \\u3_mem_reg[2][10] ,
    \\u8_mem_reg[3][29] , \\u8_mem_reg[3][2] , \\u8_mem_reg[3][30] ,
    \\u8_mem_reg[3][31] , \\u3_mem_reg[2][12] , \\u8_mem_reg[3][4] ,
    \\u3_mem_reg[2][13] , \\u8_mem_reg[3][5] , \\u3_mem_reg[2][14] ,
    \\u8_mem_reg[3][7] , \\u3_mem_reg[2][15] , \\u8_mem_reg[3][9] ,
    \\u3_mem_reg[2][16] , \\u3_mem_reg[2][17] , \\u3_mem_reg[2][19] ,
    \\u3_mem_reg[2][1] , \\u3_mem_reg[2][21] , \\u3_mem_reg[2][23] ,
    \\u3_mem_reg[2][24] , \\u3_mem_reg[2][25] , \\u3_mem_reg[2][27] ,
    \\u3_mem_reg[2][28] , \\u3_mem_reg[2][29] , \\u3_mem_reg[2][30] ,
    \\u3_mem_reg[2][31] , \\u3_mem_reg[2][3] , \\u3_mem_reg[2][4] ,
    \\u3_mem_reg[2][5] , \\u3_mem_reg[2][6] , \\u3_mem_reg[2][7] ,
    \\u3_mem_reg[2][9] , \\u3_mem_reg[3][0] , \\u3_mem_reg[3][10] ,
    \\u3_mem_reg[3][12] , \\u3_mem_reg[3][13] , \\u3_mem_reg[3][14] ,
    \\u3_mem_reg[3][16] , \\u3_mem_reg[3][17] , \\u3_mem_reg[3][18] ,
    \\u3_mem_reg[3][1] , \\u3_mem_reg[3][20] , \\u3_mem_reg[3][21] ,
    \\u3_mem_reg[3][23] , \\u3_mem_reg[3][24] , \\u3_mem_reg[3][26] ,
    \\u3_mem_reg[3][28] , \\u3_mem_reg[3][29] , \\u3_mem_reg[3][2] ,
    \\u3_mem_reg[3][31] , \\u3_mem_reg[3][4] , \\u3_mem_reg[3][5] ,
    \\u3_mem_reg[3][7] , \\u3_mem_reg[3][9] , \\u3_mem_reg[3][25] ,
    \\u4_mem_reg[1][0] , \\u4_mem_reg[1][10] , \\u4_mem_reg[1][11] ,
    \\u4_mem_reg[1][13] , \\u4_mem_reg[1][14] , \\u4_mem_reg[1][15] ,
    \\u4_mem_reg[1][17] , \\u4_mem_reg[1][18] , \\u4_mem_reg[1][19] ,
    \\u4_mem_reg[1][1] , \\u4_mem_reg[1][20] , \\u4_mem_reg[1][21] ,
    \\u4_mem_reg[1][22] , \\u4_mem_reg[1][24] , \\u4_mem_reg[1][25] ,
    \\u4_mem_reg[1][26] , \\u4_mem_reg[1][28] , \\u4_mem_reg[1][29] ,
    \\u4_mem_reg[1][2] , \\u4_mem_reg[1][31] , \\u4_mem_reg[1][3] ,
    \\u4_mem_reg[1][4] , \\u4_mem_reg[1][6] , \\u4_mem_reg[1][7] ,
    \\u4_mem_reg[1][8] , \\u4_mem_reg[2][0] , \\u4_mem_reg[2][10] ,
    \\u4_mem_reg[2][11] , \\u4_mem_reg[2][13] , \\u4_mem_reg[2][14] ,
    \\u4_mem_reg[2][15] , \\u4_mem_reg[2][17] , \\u4_mem_reg[2][18] ,
    \\u4_mem_reg[2][19] , \\u4_mem_reg[2][1] , \\u4_mem_reg[2][20] ,
    \\u4_mem_reg[2][21] , \\u4_mem_reg[2][22] , \\u4_mem_reg[2][24] ,
    \\u4_mem_reg[2][25] , \\u4_mem_reg[2][26] , \\u4_mem_reg[2][28] ,
    \\u4_mem_reg[2][29] , \\u4_mem_reg[2][2] , \\u4_mem_reg[2][31] ,
    \\u4_mem_reg[2][3] , \\u4_mem_reg[2][4] , \\u4_mem_reg[2][6] ,
    \\u4_mem_reg[2][7] , \\u4_mem_reg[2][8] , \\u4_mem_reg[3][0] ,
    \\u4_mem_reg[3][10] , \\u4_mem_reg[3][11] , \\u4_mem_reg[3][13] ,
    \\u4_mem_reg[3][14] , \\u4_mem_reg[3][15] , \\u4_mem_reg[3][17] ,
    \\u4_mem_reg[3][18] , \\u4_mem_reg[3][19] , \\u4_mem_reg[3][1] ,
    \\u4_mem_reg[3][20] , \\u4_mem_reg[3][21] , \\u4_mem_reg[3][22] ,
    \\u4_mem_reg[3][24] , \\u4_mem_reg[3][25] , \\u4_mem_reg[3][26] ,
    \\u4_mem_reg[3][28] , \\u4_mem_reg[3][29] , \\u4_mem_reg[3][2] ,
    \\u4_mem_reg[3][31] , \\u4_mem_reg[3][3] , \\u4_mem_reg[3][4] ,
    \\u4_mem_reg[3][6] , \\u4_mem_reg[3][7] , \\u4_mem_reg[3][8] ,
    \\u3_mem_reg[2][20] , \\u5_mem_reg[1][0] , \\u5_mem_reg[1][10] ,
    \\u5_mem_reg[1][12] , \\u5_mem_reg[1][13] , \\u5_mem_reg[1][14] ,
    \\u7_mem_reg[1][14] , \\u5_mem_reg[1][16] , \\u5_mem_reg[1][17] ,
    \\u5_mem_reg[1][18] , \\u5_mem_reg[1][1] , \\u5_mem_reg[1][20] ,
    \\u5_mem_reg[1][21] , \\u5_mem_reg[1][23] , \\u5_mem_reg[1][24] ,
    \\u5_mem_reg[1][25] , \\u5_mem_reg[1][27] , \\u5_mem_reg[1][28] ,
    \\u5_mem_reg[1][29] , \\u5_mem_reg[1][30] , \\u5_mem_reg[1][31] ,
    \\u5_mem_reg[1][3] , \\u5_mem_reg[1][5] , \\u5_mem_reg[1][6] ,
    \\u5_mem_reg[1][7] , \\u5_mem_reg[1][9] , \\u5_mem_reg[2][0] ,
    \\u5_mem_reg[2][10] , \\u5_mem_reg[2][12] , \\u5_mem_reg[2][13] ,
    \\u5_mem_reg[2][14] , \\u5_mem_reg[2][16] , \\u5_mem_reg[2][17] ,
    \\u5_mem_reg[2][18] , \\u5_mem_reg[2][1] , \\u5_mem_reg[2][20] ,
    \\u5_mem_reg[2][21] , \\u5_mem_reg[2][23] , \\u5_mem_reg[2][24] ,
    \\u5_mem_reg[2][25] , \\u5_mem_reg[2][27] , \\u5_mem_reg[2][28] ,
    \\u5_mem_reg[2][29] , \\u5_mem_reg[2][30] , \\u5_mem_reg[2][31] ,
    \\u5_mem_reg[2][3] , \\u5_mem_reg[2][4] , \\u5_mem_reg[2][5] ,
    \\u5_mem_reg[2][6] , \\u5_mem_reg[2][7] , \\u5_mem_reg[2][9] ,
    \\u5_mem_reg[3][0] , \\u5_mem_reg[3][10] , \\u5_mem_reg[3][12] ,
    \\u5_mem_reg[3][13] , \\u5_mem_reg[3][14] , \\u5_mem_reg[3][16] ,
    \\u5_mem_reg[3][17] , \\u5_mem_reg[3][18] , \\u5_mem_reg[3][1] ,
    \\u5_mem_reg[3][20] , \\u5_mem_reg[3][21] , \\u6_mem_reg[0][17] ,
    \\u5_mem_reg[3][23] , \\u5_mem_reg[3][24] , \\u5_mem_reg[3][25] ,
    \\u5_mem_reg[3][27] , \\u5_mem_reg[3][28] , \\u5_mem_reg[3][29] ,
    \\u5_mem_reg[3][30] , \\u5_mem_reg[3][31] , \\u5_mem_reg[3][3] ,
    \\u5_mem_reg[3][5] , \\u5_mem_reg[3][6] , \\u5_mem_reg[3][7] ,
    \\u5_mem_reg[3][9] , \\u6_mem_reg[1][0] , \\u6_mem_reg[1][10] ,
    \\u6_mem_reg[1][12] , \\u6_mem_reg[1][13] , \\u6_mem_reg[1][14] ,
    \\u6_mem_reg[1][16] , \\u6_mem_reg[1][17] , \\u6_mem_reg[1][18] ,
    \\u6_mem_reg[1][19] , \\u6_mem_reg[1][1] , \\u6_mem_reg[1][20] ,
    \\u6_mem_reg[1][21] , \\u6_mem_reg[1][23] , \\u6_mem_reg[1][24] ,
    \\u6_mem_reg[1][25] , \\u6_mem_reg[1][27] , \\u6_mem_reg[1][28] ,
    \\u6_mem_reg[1][29] , \\u6_mem_reg[1][30] , \\u6_mem_reg[1][31] ,
    \\u6_mem_reg[1][3] , \\u6_mem_reg[1][5] , \\u6_mem_reg[1][6] ,
    \\u6_mem_reg[1][7] , \\u6_mem_reg[1][9] , \\u6_mem_reg[2][0] ,
    \\u6_mem_reg[2][10] , \\u6_mem_reg[2][12] , \\u6_mem_reg[2][13] ,
    \\u6_mem_reg[2][14] , \\u6_mem_reg[2][16] , \\u6_mem_reg[2][17] ,
    \\u6_mem_reg[2][18] , \\u6_mem_reg[2][1] , \\u6_mem_reg[2][20] ,
    \\u6_mem_reg[2][21] , \\u6_mem_reg[2][23] , \\u6_mem_reg[2][24] ,
    \\u6_mem_reg[2][25] , \\u6_mem_reg[2][27] , \\u6_mem_reg[2][28] ,
    \\u6_mem_reg[2][29] , \\u6_mem_reg[2][30] , \\u6_mem_reg[2][31] ,
    \\u6_mem_reg[2][3] , \\u6_mem_reg[2][5] , \\u6_mem_reg[2][6] ,
    \\u6_mem_reg[2][7] , \\u6_mem_reg[2][9] , \\u6_mem_reg[3][0] ,
    \\u6_mem_reg[3][10] , \\u6_mem_reg[3][12] , \\u6_mem_reg[3][13] ,
    \\u6_mem_reg[3][14] , \\u6_mem_reg[3][16] , \\u6_mem_reg[3][17] ,
    \\u6_mem_reg[3][18] , \\u6_mem_reg[3][1] , \\u6_mem_reg[3][20] ,
    \\u6_mem_reg[3][21] , \\u6_mem_reg[3][23] , \\u6_mem_reg[3][24] ,
    \\u6_mem_reg[3][25] , \\u6_mem_reg[3][27] , \\u6_mem_reg[3][28] ,
    \\u6_mem_reg[3][29] , \\u6_mem_reg[3][30] , \\u6_mem_reg[3][31] ,
    \\u6_mem_reg[3][3] , \\u6_mem_reg[3][5] , \\u6_mem_reg[3][6] ,
    \\u6_mem_reg[3][7] , \\u6_mem_reg[3][9] , \\u3_mem_reg[3][8] ,
    \\u7_mem_reg[1][0] , \\u7_mem_reg[1][11] , \\u7_mem_reg[1][12] ,
    \\u7_mem_reg[1][13] , \\u7_mem_reg[1][15] , \\u7_mem_reg[1][16] ,
    \\u7_mem_reg[1][17] , \\u7_mem_reg[1][18] , \\u7_mem_reg[1][19] ,
    \\u7_mem_reg[1][1] , \\u7_mem_reg[1][20] , \\u7_mem_reg[1][22] ,
    \\u7_mem_reg[1][23] , \\u7_mem_reg[1][24] , \\u7_mem_reg[1][26] ,
    \\u7_mem_reg[1][27] , \\u7_mem_reg[1][28] , \\u7_mem_reg[1][2] ,
    \\u7_mem_reg[1][30] , \\u7_mem_reg[1][31] , \\u7_mem_reg[1][4] ,
    \\u7_mem_reg[1][5] , \\u7_mem_reg[1][6] , \\u7_mem_reg[1][8] ,
    \\u7_mem_reg[1][9] , \\u7_mem_reg[2][0] , \\u7_mem_reg[2][11] ,
    \\u7_mem_reg[2][12] , \\u7_mem_reg[2][13] , \\u7_mem_reg[2][15] ,
    \\u7_mem_reg[2][16] , \\u7_mem_reg[2][17] , \\u7_mem_reg[2][19] ,
    \\u7_mem_reg[2][1] , \\u7_mem_reg[2][20] , \\u7_mem_reg[2][22] ,
    \\u7_mem_reg[2][23] , \\u7_mem_reg[2][24] , \\u7_mem_reg[2][26] ,
    \\u7_mem_reg[2][27] , \\u7_mem_reg[2][28] , \\u7_mem_reg[2][2] ,
    \\u7_mem_reg[2][30] , \\u7_mem_reg[2][31] , \\u7_mem_reg[2][4] ,
    \\u7_mem_reg[2][5] , \\u7_mem_reg[2][6] , \\u7_mem_reg[2][8] ,
    \\u7_mem_reg[2][9] , \\u7_mem_reg[3][0] , \\u7_mem_reg[3][11] ,
    \\u7_mem_reg[3][12] , \\u7_mem_reg[3][13] , \\u7_mem_reg[3][15] ,
    \\u7_mem_reg[3][16] , \\u7_mem_reg[3][17] , \\u7_mem_reg[3][19] ,
    \\u7_mem_reg[3][1] , \\u7_mem_reg[3][20] , \\u6_mem_reg[0][20] ,
    \\u7_mem_reg[3][22] , \\u7_mem_reg[3][23] , \\u7_mem_reg[3][24] ,
    \\u7_mem_reg[3][26] , \\u7_mem_reg[3][27] , \\u7_mem_reg[3][28] ,
    \\u7_mem_reg[3][2] , \\u7_mem_reg[3][30] , \\u7_mem_reg[3][31] ,
    \\u7_mem_reg[3][4] , \\u7_mem_reg[3][5] , \\u7_mem_reg[3][6] ,
    \\u7_mem_reg[3][8] , \\u7_mem_reg[3][9] , \\u8_mem_reg[1][0] ,
    \\u8_mem_reg[1][11] , \\u8_mem_reg[1][12] , \\u8_mem_reg[1][13] ,
    \\u8_mem_reg[1][15] , \\u8_mem_reg[1][16] , \\u8_mem_reg[1][17] ,
    \\u8_mem_reg[1][19] , \\u8_mem_reg[1][1] , \\u8_mem_reg[1][20] ,
    \\u8_mem_reg[1][22] , \\u8_mem_reg[1][23] , \\u8_mem_reg[1][24] ,
    \\u8_mem_reg[1][26] , \\u3_mem_reg[1][0] , \\u8_mem_reg[1][27] ,
    \\u3_mem_reg[1][10] , \\u8_mem_reg[1][29] , \\u8_mem_reg[1][2] ,
    \\u8_mem_reg[1][30] , \\u8_mem_reg[1][31] , \\u3_mem_reg[1][12] ,
    \\u8_mem_reg[1][4] , \\u3_mem_reg[1][13] , \\u8_mem_reg[1][5] ,
    \\u3_mem_reg[1][14] , \\u8_mem_reg[1][7] , \\u8_mem_reg[1][8] ,
    \\u8_mem_reg[1][9] , \\u8_mem_reg[2][0] , \\u3_mem_reg[1][16] ,
    \\u8_mem_reg[2][10] , \\u8_mem_reg[2][11] , \\u3_mem_reg[1][17] ,
    \\u8_mem_reg[2][12] , \\u3_mem_reg[1][18] , \\u8_mem_reg[2][14] ,
    \\u8_mem_reg[2][15] , \\u8_mem_reg[2][16] , \\u8_mem_reg[2][17] ,
    \\u3_mem_reg[1][1] , \\u8_mem_reg[2][19] , \\u3_mem_reg[1][20] ,
    \\u8_mem_reg[2][1] , \\u3_mem_reg[1][21] , \\u8_mem_reg[2][21] ,
    \\u8_mem_reg[2][22] , \\u8_mem_reg[2][23] , \\u8_mem_reg[2][24] ,
    \\u3_mem_reg[1][23] , \\u8_mem_reg[2][26] , \\u3_mem_reg[1][24] ,
    \\u8_mem_reg[2][27] , \\u3_mem_reg[1][25] , \\u8_mem_reg[2][29] ,
    \\u8_mem_reg[2][2] , \\u8_mem_reg[2][30] , \\u8_mem_reg[2][31] ,
    \\u3_mem_reg[1][27] , \\u4_mem_reg[0][0] , \\u4_mem_reg[0][10] ,
    \\u4_mem_reg[0][11] , \\u4_mem_reg[0][15] , \\u4_mem_reg[0][18] ,
    \\u4_mem_reg[0][1] , \\u4_mem_reg[0][21] , \\u4_mem_reg[0][25] ,
    \\u4_mem_reg[0][27] , \\u4_mem_reg[0][28] , \\u4_mem_reg[0][26] ,
    \\u4_mem_reg[0][2] , \\u4_mem_reg[0][29] , \\u4_mem_reg[0][3] ,
    \\u4_mem_reg[0][5] , \\u4_mem_reg[0][8] , \\u5_mem_reg[0][10] ,
    \\u5_mem_reg[0][11] , \\u5_mem_reg[0][15] , \\u5_mem_reg[0][18] ,
    \\u5_mem_reg[0][1] , \\u5_mem_reg[0][21] , \\u13_intm_r_reg[8] ,
    \\u5_mem_reg[0][26] , \\u5_mem_reg[0][27] , \\u5_mem_reg[0][25] ,
    \\u5_mem_reg[0][2] , \\u5_mem_reg[0][29] , \\u5_mem_reg[0][3] ,
    \\u5_mem_reg[0][5] , \\u5_mem_reg[0][8] , \\u6_mem_reg[0][10] ,
    \\u6_mem_reg[0][11] , \\u6_mem_reg[0][15] , \\u7_mem_reg[1][21] ,
    \\u6_mem_reg[0][18] , \\u6_mem_reg[0][1] , \\u6_mem_reg[0][21] ,
    \\u6_mem_reg[0][26] , \\u6_mem_reg[0][27] , \\u6_mem_reg[0][25] ,
    \\u6_mem_reg[0][2] , \\u6_mem_reg[0][29] , \\u6_mem_reg[0][3] ,
    \\u6_mem_reg[0][5] , \\u6_mem_reg[0][8] , \\u7_mem_reg[0][10] ,
    \\u7_mem_reg[0][11] , \\u7_mem_reg[0][15] , \\u7_mem_reg[0][18] ,
    \\u7_mem_reg[0][1] , \\u7_mem_reg[0][21] , \\u7_mem_reg[0][25] ,
    \\u7_mem_reg[0][27] , \\u7_mem_reg[0][28] , \\u7_mem_reg[0][26] ,
    \\u7_mem_reg[0][2] , \\u7_mem_reg[0][29] , \\u7_mem_reg[0][3] ,
    \\u7_mem_reg[0][5] , \\u7_mem_reg[0][8] , \\u3_mem_reg[0][10] ,
    \\u8_mem_reg[0][10] , \\u8_mem_reg[0][13] , \\u3_mem_reg[0][18] ,
    \\u8_mem_reg[0][14] , \\u3_mem_reg[0][19] , \\u8_mem_reg[0][18] ,
    \\u8_mem_reg[0][19] , \\u3_mem_reg[0][20] , \\u8_mem_reg[0][20] ,
    \\u8_mem_reg[0][21] , \\u3_mem_reg[0][22] , \\u8_mem_reg[0][23] ,
    \\u8_mem_reg[0][24] , \\u8_mem_reg[0][25] , \\u3_mem_reg[0][24] ,
    \\u3_mem_reg[0][25] , \\u3_mem_reg[0][26] , \\u3_mem_reg[0][28] ,
    \\u8_mem_reg[0][7] , \\u8_mem_reg[0][8] , \\u8_mem_reg[0][6] ,
    \\u8_mem_reg[0][9] , \\u3_mem_reg[0][30] , \\u3_mem_reg[0][3] ,
    \\u3_mem_reg[0][8] , \\u7_mem_reg[1][10] , \\u13_crac_dout_r_reg[7] ,
    \\u6_mem_reg[2][22] , \\u6_mem_reg[0][0] , \\u6_mem_reg[3][4] ,
    \\u13_intm_r_reg[26] , \\u6_mem_reg[3][2] , \\u13_occ0_r_reg[22] ,
    \\u6_mem_reg[3][26] , \\u6_mem_reg[3][22] , \\u6_mem_reg[3][15] ,
    \\u5_mem_reg[0][6] , \\u6_mem_reg[3][19] , \\u1_sr_reg[10] ,
    \\u5_mem_reg[0][30] , \\u5_mem_reg[0][23] , \\u13_crac_r_reg[2] ,
    \\u6_mem_reg[2][4] , \\u6_mem_reg[3][11] , \\u6_mem_reg[2][8] ,
    \\u6_mem_reg[2][2] , \\u3_mem_reg[0][9] , \\u13_occ0_r_reg[26] ,
    \\u5_mem_reg[0][28] , \\u13_intm_r_reg[3] , \\u6_mem_reg[2][26] ,
    \\u3_mem_reg[0][4] , \\u5_mem_reg[0][20] , \\u8_mem_reg[0][31] ,
    \\u6_mem_reg[2][15] , \\u6_mem_reg[1][15] , \\u6_mem_reg[2][19] ,
    \\u6_mem_reg[2][11] , \\u5_mem_reg[0][17] , \\u13_occ0_r_reg[19] ,
    \\u5_mem_reg[0][12] , \\u6_mem_reg[1][26] , \\u4_mem_reg[0][6] ,
    \\u6_mem_reg[1][4] , \\u6_mem_reg[1][8] , \\u6_mem_reg[1][2] ,
    \\u5_mem_reg[0][0] , \\u6_mem_reg[1][22] , \\u8_mem_reg[0][3] ,
    \\u4_mem_reg[0][30] , \\u8_mem_reg[0][16] , \\u5_mem_reg[3][8] ,
    \\u6_mem_reg[1][11] , \\u5_mem_reg[3][4] , \\u8_mem_reg[0][2] ,
    \\u5_mem_reg[2][8] , \\u4_mem_reg[0][23] , \\u3_mem_reg[0][23] ,
    \\u4_mem_reg[0][17] , \\u5_mem_reg[3][19] , \\u5_mem_reg[3][26] ,
    \\u5_mem_reg[3][2] , \\u5_mem_reg[3][22] , \\u5_mem_reg[3][15] ,
    \\u8_mem_reg[0][27] , \\u4_mem_reg[0][20] , \\u5_mem_reg[3][11] ,
    \\u5_mem_reg[2][2] , \\u4_mem_reg[0][12] , \\u5_mem_reg[2][26] ,
    \\u8_mem_reg[0][22] , \\u13_occ0_r_reg[15] , \\u5_mem_reg[1][2] ,
    \\u5_mem_reg[2][11] , \\u3_mem_reg[1][26] , \\u5_mem_reg[2][19] ,
    \\u5_mem_reg[2][22] , \\u5_mem_reg[2][15] , \\u8_mem_reg[2][3] ,
    \\u5_mem_reg[1][8] , \\u5_mem_reg[1][4] , \\u8_mem_reg[0][1] ,
    \\u13_occ1_r_reg[11] , \\u3_mem_reg[0][0] , u14_u8_en_out_l2_reg,
    \\u12_wb_data_o_reg[4] , \\u12_wb_data_o_reg[6] ,
    \\u12_wb_data_o_reg[10] , \\u13_occ1_r_reg[8] , \\u13_occ1_r_reg[0] ,
    \\u13_occ1_r_reg[10] , \\u13_occ1_r_reg[12] , \\u13_occ1_r_reg[13] ,
    \\u13_occ1_r_reg[14] , \\u13_occ1_r_reg[1] , \\u13_occ1_r_reg[2] ,
    \\u13_occ1_r_reg[3] , \\u13_occ1_r_reg[5] , \\u13_occ1_r_reg[6] ,
    \\u13_occ1_r_reg[7] , \\u1_slt1_reg[7] , \\u1_slt2_reg[7] ,
    \\u1_slt4_reg[7] , \\u1_slt3_reg[7] , \\u3_mem_reg[0][14] ,
    \\u3_mem_reg[0][7] , u14_u6_full_empty_r_reg, u14_u8_full_empty_r_reg,
    \\u12_wb_data_o_reg[0] , \\u12_wb_data_o_reg[14] ,
    \\u12_wb_data_o_reg[13] , \\u12_wb_data_o_reg[12] ,
    \\u12_wb_data_o_reg[11] , \\u12_wb_data_o_reg[9] ,
    \\u12_wb_data_o_reg[7] , \\u12_wb_data_o_reg[15] ,
    \\u12_wb_data_o_reg[5] , \\u12_wb_data_o_reg[3] ,
    \\u12_wb_data_o_reg[8] , \\u12_wb_data_o_reg[2] , \\u13_occ1_r_reg[9] ,
    \\u13_occ1_r_reg[15] , \\u3_mem_reg[0][31] , \\u13_occ1_r_reg[4] ,
    \\u0_slt9_r_reg[1] , \\u1_slt6_reg[7] , u14_u7_en_out_l2_reg,
    u14_u7_full_empty_r_reg, u13_ac97_rst_force_reg, u13_resume_req_reg,
    \\u1_sr_reg[9] , u14_u6_en_out_l2_reg, \\u12_wb_data_o_reg[31] ,
    \\u1_slt3_reg[6] , \\u1_slt1_reg[6] , \\u1_slt2_reg[6] ,
    \\u1_slt4_reg[6] , \\u12_wb_data_o_reg[23] , \\u12_wb_data_o_reg[22] ,
    \\u12_wb_data_o_reg[21] , \\u12_wb_data_o_reg[16] ,
    \\u12_wb_data_o_reg[20] , \\u12_wb_data_o_reg[19] ,
    \\u12_wb_data_o_reg[17] , \\u12_wb_data_o_reg[24] ,
    \\u12_wb_data_o_reg[30] , \\u12_wb_data_o_reg[28] ,
    \\u12_wb_data_o_reg[27] , \\u12_wb_data_o_reg[26] ,
    \\u12_wb_data_o_reg[29] , \\u12_wb_data_o_reg[25] , \\u1_slt6_reg[6] ,
    \\u12_wb_data_o_reg[18] , u4_empty_reg, u6_empty_reg,
    u15_crac_we_r_reg, \\u1_sr_reg[8] , u3_empty_reg, u5_empty_reg,
    u7_empty_reg, u8_empty_reg, \\u10_rp_reg[2] , \\u11_rp_reg[2] ,
    \\u23_int_set_reg[1] , \\u24_int_set_reg[1] , \\u11_rp_reg[1] ,
    \\u9_rp_reg[1] , \\u10_rp_reg[1] , \\u11_rp_reg[0] , \\u9_rp_reg[0] ,
    \\u9_rp_reg[2] , \\u10_rp_reg[0] , \\u1_slt1_reg[5] ,
    \\u1_slt2_reg[5] , \\u1_slt4_reg[5] , \\u1_slt3_reg[5] ,
    \\u1_slt6_reg[5] , \\u25_int_set_reg[1] , \\u1_sr_reg[7] ,
    \\u0_slt9_r_reg[0] , valid_s_reg, \\in_valid_s_reg[0] ,
    \\u1_slt2_reg[4] , \\u1_slt3_reg[4] , \\u1_slt4_reg[4] ,
    \\u1_slt6_reg[4] , u12_o7_we_reg, u12_o3_we_reg, u12_o4_we_reg,
    u12_o6_we_reg, u12_o8_we_reg, u12_o9_we_reg, \\u1_sr_reg[6] ,
    \\in_valid_s_reg[2] , \\u2_to_cnt_reg[5] , u13_int_reg,
    \\u13_ints_r_reg[21] , \\u1_slt3_reg[0] , \\u13_ints_r_reg[0] ,
    \\u13_ints_r_reg[27] , \\u13_ints_r_reg[15] , \\u2_cnt_reg[7] ,
    \\in_valid_s_reg[1] , valid_s1_reg, \\in_valid_s1_reg[0] ,
    \\u2_to_cnt_reg[3] , \\u2_res_cnt_reg[3] , \\u2_to_cnt_reg[4] ,
    \\u1_slt3_reg[2] , \\u1_slt3_reg[1] , \\u1_slt4_reg[1] ,
    \\u1_slt6_reg[1] , \\u1_slt6_reg[2] , u12_wb_ack_o_reg,
    \\u13_ints_r_reg[10] , \\u13_ints_r_reg[12] , \\u13_ints_r_reg[13] ,
    \\u13_ints_r_reg[16] , \\u13_ints_r_reg[18] , \\u13_ints_r_reg[19] ,
    \\u13_ints_r_reg[22] , \\u13_ints_r_reg[24] , \\u13_ints_r_reg[25] ,
    \\u13_ints_r_reg[28] , \\u13_ints_r_reg[3] , \\u13_ints_r_reg[4] ,
    \\u13_ints_r_reg[7] , \\u13_ints_r_reg[6] , \\u1_slt6_reg[3] ,
    \\u1_slt6_reg[0] , \\u1_slt4_reg[3] , \\u1_slt3_reg[3] ,
    \\u13_ints_r_reg[9] , \\u1_slt4_reg[2] , \\u1_slt4_reg[0] ,
    \\u2_cnt_reg[1] , \\u2_to_cnt_reg[2] , \\u4_status_reg[1] ,
    \\u5_status_reg[1] , u12_rf_we_reg, \\u2_res_cnt_reg[0] ,
    \\in_valid_s1_reg[2] , \\u1_sr_reg[5] , \\u2_cnt_reg[4] ,
    \\u2_cnt_reg[3] , \\u2_to_cnt_reg[0] , \\u2_to_cnt_reg[1] ,
    \\u2_cnt_reg[5] , \\u2_cnt_reg[6] , \\u2_cnt_reg[0] , \\u2_cnt_reg[2] ,
    \\u2_res_cnt_reg[2] , u2_valid_reg, \\u2_res_cnt_reg[1] ,
    \\u3_status_reg[1] , \\u6_status_reg[1] , \\u7_status_reg[1] ,
    \\u8_status_reg[1] , \\u11_status_reg[1] , u10_empty_reg, u9_empty_reg,
    \\in_valid_s1_reg[1] , \\u2_in_valid_reg[0] , u12_we1_reg,
    \\u1_sr_reg[4] , \\u2_in_valid_reg[2] , \\u10_status_reg[1] ,
    \\u9_status_reg[1] , u11_empty_reg, u2_sync_beat_reg, u11_full_reg,
    \\u10_dout_reg[14] , \\u10_dout_reg[15] , \\u10_dout_reg[17] ,
    \\u10_dout_reg[18] , \\u10_dout_reg[19] , \\u10_dout_reg[1] ,
    \\u10_dout_reg[20] , \\u10_dout_reg[21] , \\u10_dout_reg[22] ,
    \\u10_dout_reg[23] , u12_i4_re_reg, u2_ld_reg, u9_full_reg,
    u12_i6_re_reg, \\u2_out_le_reg[1] , u12_i3_re_reg,
    \\u2_in_valid_reg[1] , \\u10_dout_reg[11] , \\u10_dout_reg[0] ,
    \\u10_dout_reg[10] , \\u10_dout_reg[12] , \\u10_dout_reg[13] ,
    \\u10_dout_reg[25] , \\u10_dout_reg[27] , \\u10_dout_reg[28] ,
    \\u10_dout_reg[29] , \\u10_dout_reg[2] , \\u10_dout_reg[30] ,
    \\u10_dout_reg[3] , \\u10_dout_reg[4] , \\u10_dout_reg[6] ,
    \\u10_dout_reg[7] , \\u10_dout_reg[8] , \\u10_dout_reg[9] ,
    u10_full_reg, \\u2_out_le_reg[2] , \\u2_out_le_reg[4] ,
    \\u2_out_le_reg[5] , \\u2_out_le_reg[3] , \\u2_out_le_reg[0] ,
    \\u9_dout_reg[11] , \\u9_dout_reg[14] , \\u9_dout_reg[18] ,
    \\u9_dout_reg[19] , \\u9_dout_reg[20] , \\u9_dout_reg[21] ,
    \\u9_dout_reg[22] , \\u9_dout_reg[23] , \\u9_dout_reg[24] ,
    \\u9_dout_reg[25] , \\u9_dout_reg[16] , \\u10_dout_reg[16] ,
    \\u9_dout_reg[26] , \\u9_dout_reg[27] , \\u9_dout_reg[28] ,
    \\u9_dout_reg[29] , \\u9_dout_reg[2] , \\u9_dout_reg[30] ,
    \\u9_dout_reg[31] , \\u9_dout_reg[3] , \\u1_sr_reg[3] ,
    \\u9_dout_reg[4] , \\u9_dout_reg[5] , \\u9_dout_reg[6] ,
    \\u9_dout_reg[7] , \\u9_dout_reg[8] , \\u9_dout_reg[9] ,
    \\u10_dout_reg[24] , \\u10_dout_reg[26] , \\u9_dout_reg[13] ,
    \\u11_dout_reg[0] , \\u11_dout_reg[10] , \\u11_dout_reg[11] ,
    \\u11_dout_reg[12] , \\u11_dout_reg[13] , \\u10_dout_reg[31] ,
    \\u11_dout_reg[14] , \\u11_dout_reg[15] , \\u11_dout_reg[16] ,
    \\u11_dout_reg[17] , \\u11_dout_reg[18] , \\u11_dout_reg[19] ,
    \\u10_dout_reg[5] , \\u11_dout_reg[1] , \\u11_dout_reg[20] ,
    \\u11_dout_reg[21] , \\u11_dout_reg[22] , \\u11_dout_reg[23] ,
    \\u11_dout_reg[24] , \\u11_dout_reg[25] , \\u11_dout_reg[26] ,
    \\u11_dout_reg[27] , \\u11_dout_reg[28] , \\u11_dout_reg[29] ,
    \\u11_dout_reg[2] , \\u11_dout_reg[30] , \\u11_dout_reg[31] ,
    \\u11_dout_reg[3] , \\u11_dout_reg[4] , \\u11_dout_reg[5] ,
    \\u11_dout_reg[6] , \\u11_dout_reg[7] , \\u11_dout_reg[8] ,
    \\u11_dout_reg[9] , \\u9_dout_reg[15] , \\u9_dout_reg[17] ,
    \\u9_dout_reg[0] , \\u9_dout_reg[12] , \\u9_dout_reg[10] ,
    \\u9_dout_reg[1] , u12_re2_reg, u12_re1_reg, u2_bit_clk_e_reg,
    u2_suspended_reg, \\u10_status_reg[0] , \\u9_status_reg[0] ,
    \\u11_status_reg[0] , \\u6_status_reg[0] , \\u3_status_reg[0] ,
    \\u4_status_reg[0] , \\u7_status_reg[0] , \\u1_sr_reg[2] ,
    \\u15_crac_din_reg[6] , \\u15_crac_din_reg[9] ,
    \\u15_crac_din_reg[12] , \\u15_crac_din_reg[1] ,
    \\u15_crac_din_reg[7] , \\u15_crac_din_reg[14] ,
    \\u15_crac_din_reg[10] , \\u15_crac_din_reg[15] ,
    \\u15_crac_din_reg[4] , \\u15_crac_din_reg[8] ,
    \\u15_crac_din_reg[11] , \\u15_crac_din_reg[13] ,
    \\u15_crac_din_reg[2] , \\u15_crac_din_reg[0] , \\u15_crac_din_reg[5] ,
    \\u5_status_reg[0] , \\u8_status_reg[0] , \\u15_crac_din_reg[3] ,
    \\u1_sr_reg[1] , u12_we2_reg, u2_bit_clk_r1_reg, \\u1_sr_reg[0] ,
    u1_sdata_in_r_reg, \\u12_dout_reg[7] , \\u12_dout_reg[4] ,
    \\u12_dout_reg[12] , \\u12_dout_reg[24] , \\u12_dout_reg[26] ,
    \\u12_dout_reg[23] , \\u12_dout_reg[11] , \\u12_dout_reg[31] ,
    \\u12_dout_reg[13] , \\u12_dout_reg[29] , \\u12_dout_reg[22] ,
    \\u12_dout_reg[30] , \\u12_dout_reg[15] , \\u12_dout_reg[19] ,
    u2_bit_clk_r_reg, \\u12_dout_reg[27] , \\u12_dout_reg[28] ,
    \\u12_dout_reg[10] , \\u12_dout_reg[6] , \\u12_dout_reg[20] ,
    \\u12_dout_reg[0] , \\u12_dout_reg[21] , \\u12_dout_reg[5] ,
    \\u12_dout_reg[18] , \\u12_dout_reg[25] , \\u12_dout_reg[2] ,
    \\u12_dout_reg[9] , \\u12_dout_reg[17] , \\u12_dout_reg[3] ,
    \\u12_dout_reg[8] , \\u12_dout_reg[16] , \\u12_dout_reg[14] ,
    \\u12_dout_reg[1] ;
  wire \new_[2331]_ , \new_[2336]_ , \new_[2337]_ , \new_[2339]_ ,
    \new_[2341]_ , \new_[2343]_ , \new_[2345]_ , \new_[2347]_ ,
    \new_[2349]_ , \new_[2351]_ , \new_[2353]_ , \new_[2355]_ ,
    \new_[2356]_ , \new_[2358]_ , \new_[2360]_ , \new_[2362]_ ,
    \new_[2364]_ , \new_[2366]_ , \new_[2368]_ , \new_[2370]_ ,
    \new_[2372]_ , \new_[2374]_ , \new_[2376]_ , \new_[2378]_ ,
    \new_[2380]_ , \new_[2382]_ , \new_[2384]_ , \new_[2386]_ ,
    \new_[2388]_ , \new_[2390]_ , \new_[2392]_ , \new_[2394]_ ,
    \new_[2396]_ , \new_[2398]_ , \new_[2400]_ , \new_[2402]_ ,
    \new_[2404]_ , \new_[2406]_ , \new_[2408]_ , \new_[2410]_ ,
    \new_[2412]_ , \new_[2414]_ , \new_[2416]_ , \new_[2418]_ ,
    \new_[2420]_ , \new_[2422]_ , \new_[2424]_ , \new_[2426]_ ,
    \new_[2428]_ , \new_[2430]_ , \new_[2432]_ , \new_[2434]_ ,
    \new_[2436]_ , \new_[2438]_ , \new_[2440]_ , \new_[2442]_ ,
    \new_[2444]_ , \new_[2446]_ , \new_[2448]_ , \new_[2450]_ ,
    \new_[2452]_ , \new_[2454]_ , \new_[2456]_ , \new_[2458]_ ,
    \new_[2460]_ , \new_[2462]_ , \new_[2464]_ , \new_[2466]_ ,
    \new_[2468]_ , \new_[2470]_ , \new_[2472]_ , \new_[2474]_ ,
    \new_[2476]_ , \new_[2478]_ , \new_[2480]_ , \new_[2482]_ ,
    \new_[2484]_ , \new_[2486]_ , \new_[2488]_ , \new_[2490]_ ,
    \new_[2492]_ , \new_[2494]_ , \new_[2496]_ , \new_[2498]_ ,
    \new_[2500]_ , \new_[2502]_ , \new_[2504]_ , \new_[2506]_ ,
    \new_[2508]_ , \new_[2510]_ , \new_[2512]_ , \new_[2514]_ ,
    \new_[2516]_ , \new_[2518]_ , \new_[2520]_ , \new_[2522]_ ,
    \new_[2524]_ , \new_[2526]_ , \new_[2528]_ , \new_[2530]_ ,
    \new_[2532]_ , \new_[2534]_ , \new_[2536]_ , \new_[2538]_ ,
    \new_[2540]_ , \new_[2542]_ , \new_[2544]_ , \new_[2546]_ ,
    \new_[2548]_ , \new_[2550]_ , \new_[2552]_ , \new_[2554]_ ,
    \new_[2556]_ , \new_[2558]_ , \new_[2560]_ , \new_[2562]_ ,
    \new_[2564]_ , \new_[2566]_ , \new_[2568]_ , \new_[2570]_ ,
    \new_[2572]_ , \new_[2574]_ , \new_[2576]_ , \new_[2578]_ ,
    \new_[2580]_ , \new_[2582]_ , \new_[2584]_ , \new_[2586]_ ,
    \new_[2588]_ , \new_[2590]_ , \new_[2592]_ , \new_[2594]_ ,
    \new_[2596]_ , \new_[2598]_ , \new_[2600]_ , \new_[2602]_ ,
    \new_[2604]_ , \new_[2606]_ , \new_[2608]_ , \new_[2610]_ ,
    \new_[2612]_ , \new_[2614]_ , \new_[2616]_ , \new_[2618]_ ,
    \new_[2620]_ , \new_[2622]_ , \new_[2624]_ , \new_[2626]_ ,
    \new_[2628]_ , \new_[2630]_ , \new_[2632]_ , \new_[2634]_ ,
    \new_[2636]_ , \new_[2638]_ , \new_[2640]_ , \new_[2642]_ ,
    \new_[2644]_ , \new_[2646]_ , \new_[2648]_ , \new_[2650]_ ,
    \new_[2652]_ , \new_[2654]_ , \new_[2656]_ , \new_[2658]_ ,
    \new_[2660]_ , \new_[2662]_ , \new_[2664]_ , \new_[2666]_ ,
    \new_[2668]_ , \new_[2670]_ , \new_[2672]_ , \new_[2674]_ ,
    \new_[2676]_ , \new_[2678]_ , \new_[2680]_ , \new_[2682]_ ,
    \new_[2684]_ , \new_[2686]_ , \new_[2688]_ , \new_[2690]_ ,
    \new_[2692]_ , \new_[2694]_ , \new_[2696]_ , \new_[2698]_ ,
    \new_[2700]_ , \new_[2702]_ , \new_[2704]_ , \new_[2706]_ ,
    \new_[2708]_ , \new_[2710]_ , \new_[2712]_ , \new_[2714]_ ,
    \new_[2715]_ , \new_[2716]_ , \new_[2717]_ , \new_[2718]_ ,
    \new_[2724]_ , \new_[2725]_ , \new_[2726]_ , \new_[2727]_ ,
    \new_[2730]_ , \new_[2735]_ , \new_[2736]_ , \new_[2737]_ ,
    \new_[2738]_ , \new_[2745]_ , \new_[2746]_ , \new_[2747]_ ,
    \new_[2748]_ , \new_[2749]_ , \new_[2750]_ , \new_[2751]_ ,
    \new_[2752]_ , \new_[2753]_ , \new_[2754]_ , \new_[2755]_ ,
    \new_[2756]_ , \new_[2757]_ , \new_[2758]_ , \new_[2759]_ ,
    \new_[2769]_ , \new_[2770]_ , \new_[2771]_ , \new_[2772]_ ,
    \new_[2773]_ , \new_[2774]_ , \new_[2783]_ , \new_[2784]_ ,
    \new_[2785]_ , \new_[2786]_ , \new_[2787]_ , \new_[2788]_ ,
    \new_[2789]_ , \new_[2790]_ , \new_[2791]_ , \new_[2792]_ ,
    \new_[2793]_ , \new_[2794]_ , \new_[2795]_ , \new_[2796]_ ,
    \new_[2797]_ , \new_[2798]_ , \new_[2799]_ , \new_[2800]_ ,
    \new_[2801]_ , \new_[2802]_ , \new_[2803]_ , \new_[2804]_ ,
    \new_[2805]_ , \new_[2816]_ , \new_[2817]_ , \new_[2818]_ ,
    \new_[2819]_ , \new_[2820]_ , \new_[2821]_ , \new_[2822]_ ,
    \new_[2823]_ , \new_[2824]_ , \new_[2825]_ , \new_[2826]_ ,
    \new_[2827]_ , \new_[2828]_ , \new_[2829]_ , \new_[2830]_ ,
    \new_[2831]_ , \new_[2832]_ , \new_[2833]_ , \new_[2834]_ ,
    \new_[2835]_ , \new_[2836]_ , \new_[2837]_ , \new_[2838]_ ,
    \new_[2839]_ , \new_[2840]_ , \new_[2841]_ , \new_[2842]_ ,
    \new_[2843]_ , \new_[2844]_ , \new_[2845]_ , \new_[2846]_ ,
    \new_[2847]_ , \new_[2848]_ , \new_[2849]_ , \new_[2850]_ ,
    \new_[2851]_ , \new_[2852]_ , \new_[2853]_ , \new_[2854]_ ,
    \new_[2855]_ , \new_[2856]_ , \new_[2857]_ , \new_[2858]_ ,
    \new_[2859]_ , \new_[2860]_ , \new_[2861]_ , \new_[2862]_ ,
    \new_[2863]_ , \new_[2864]_ , \new_[2865]_ , \new_[2866]_ ,
    \new_[2867]_ , \new_[2868]_ , \new_[2869]_ , \new_[2870]_ ,
    \new_[2871]_ , \new_[2872]_ , \new_[2873]_ , \new_[2874]_ ,
    \new_[2875]_ , \new_[2876]_ , \new_[2877]_ , \new_[2878]_ ,
    \new_[2879]_ , \new_[2880]_ , \new_[2881]_ , \new_[2882]_ ,
    \new_[2883]_ , \new_[2884]_ , \new_[2885]_ , \new_[2886]_ ,
    \new_[2887]_ , \new_[2888]_ , \new_[2889]_ , \new_[2890]_ ,
    \new_[2891]_ , \new_[2892]_ , \new_[2893]_ , \new_[2894]_ ,
    \new_[2895]_ , \new_[2896]_ , \new_[2897]_ , \new_[2898]_ ,
    \new_[2904]_ , \new_[2905]_ , \new_[2910]_ , \new_[2911]_ ,
    \new_[2912]_ , \new_[2913]_ , \new_[2914]_ , \new_[2917]_ ,
    \new_[2920]_ , \new_[2922]_ , \new_[2923]_ , \new_[2924]_ ,
    \new_[2925]_ , \new_[2926]_ , \new_[2927]_ , \new_[2928]_ ,
    \new_[2929]_ , \new_[2930]_ , \new_[2931]_ , \new_[2932]_ ,
    \new_[2933]_ , \new_[2949]_ , \new_[2952]_ , \new_[3019]_ ,
    \new_[3020]_ , \new_[3021]_ , \new_[3022]_ , \new_[3023]_ ,
    \new_[3024]_ , \new_[3025]_ , \new_[3026]_ , \new_[3027]_ ,
    \new_[3028]_ , \new_[3029]_ , \new_[3030]_ , \new_[3031]_ ,
    \new_[3032]_ , \new_[3033]_ , \new_[3034]_ , \new_[3035]_ ,
    \new_[3036]_ , \new_[3037]_ , \new_[3038]_ , \new_[3039]_ ,
    \new_[3040]_ , \new_[3041]_ , \new_[3042]_ , \new_[3043]_ ,
    \new_[3044]_ , \new_[3045]_ , \new_[3046]_ , \new_[3047]_ ,
    \new_[3048]_ , \new_[3049]_ , \new_[3050]_ , \new_[3051]_ ,
    \new_[3052]_ , \new_[3053]_ , \new_[3054]_ , \new_[3055]_ ,
    \new_[3056]_ , \new_[3057]_ , \new_[3058]_ , \new_[3059]_ ,
    \new_[3060]_ , \new_[3061]_ , \new_[3062]_ , \new_[3063]_ ,
    \new_[3064]_ , \new_[3065]_ , \new_[3066]_ , \new_[3067]_ ,
    \new_[3068]_ , \new_[3069]_ , \new_[3070]_ , \new_[3071]_ ,
    \new_[3072]_ , \new_[3073]_ , \new_[3074]_ , \new_[3075]_ ,
    \new_[3076]_ , \new_[3077]_ , \new_[3078]_ , \new_[3079]_ ,
    \new_[3080]_ , \new_[3081]_ , \new_[3082]_ , \new_[3083]_ ,
    \new_[3084]_ , \new_[3085]_ , \new_[3086]_ , \new_[3087]_ ,
    \new_[3088]_ , \new_[3089]_ , \new_[3090]_ , \new_[3091]_ ,
    \new_[3092]_ , \new_[3093]_ , \new_[3094]_ , \new_[3095]_ ,
    \new_[3096]_ , \new_[3097]_ , \new_[3098]_ , \new_[3099]_ ,
    \new_[3100]_ , \new_[3101]_ , \new_[3102]_ , \new_[3103]_ ,
    \new_[3104]_ , \new_[3105]_ , \new_[3106]_ , \new_[3107]_ ,
    \new_[3108]_ , \new_[3109]_ , \new_[3110]_ , \new_[3111]_ ,
    \new_[3112]_ , \new_[3113]_ , \new_[3114]_ , \new_[3115]_ ,
    \new_[3116]_ , \new_[3117]_ , \new_[3118]_ , \new_[3119]_ ,
    \new_[3120]_ , \new_[3121]_ , \new_[3122]_ , \new_[3123]_ ,
    \new_[3128]_ , \new_[3130]_ , \new_[3134]_ , \new_[3137]_ ,
    \new_[3138]_ , \new_[3139]_ , \new_[3140]_ , \new_[3141]_ ,
    \new_[3142]_ , \new_[3143]_ , \new_[3144]_ , \new_[3145]_ ,
    \new_[3146]_ , \new_[3147]_ , \new_[3148]_ , \new_[3149]_ ,
    \new_[3150]_ , \new_[3151]_ , \new_[3152]_ , \new_[3153]_ ,
    \new_[3154]_ , \new_[3157]_ , \new_[3158]_ , \new_[3159]_ ,
    \new_[3161]_ , \new_[3163]_ , \new_[3164]_ , \new_[3165]_ ,
    \new_[3166]_ , \new_[3167]_ , \new_[3168]_ , \new_[3169]_ ,
    \new_[3170]_ , \new_[3171]_ , \new_[3172]_ , \new_[3173]_ ,
    \new_[3174]_ , \new_[3175]_ , \new_[3176]_ , \new_[3177]_ ,
    \new_[3178]_ , \new_[3179]_ , \new_[3180]_ , \new_[3181]_ ,
    \new_[3182]_ , \new_[3183]_ , \new_[3184]_ , \new_[3185]_ ,
    \new_[3186]_ , \new_[3187]_ , \new_[3188]_ , \new_[3189]_ ,
    \new_[3190]_ , \new_[3191]_ , \new_[3192]_ , \new_[3193]_ ,
    \new_[3194]_ , \new_[3195]_ , \new_[3196]_ , \new_[3197]_ ,
    \new_[3198]_ , \new_[3199]_ , \new_[3200]_ , \new_[3201]_ ,
    \new_[3202]_ , \new_[3203]_ , \new_[3204]_ , \new_[3205]_ ,
    \new_[3206]_ , \new_[3207]_ , \new_[3208]_ , \new_[3209]_ ,
    \new_[3210]_ , \new_[3211]_ , \new_[3212]_ , \new_[3213]_ ,
    \new_[3214]_ , \new_[3215]_ , \new_[3216]_ , \new_[3217]_ ,
    \new_[3218]_ , \new_[3219]_ , \new_[3220]_ , \new_[3221]_ ,
    \new_[3222]_ , \new_[3223]_ , \new_[3224]_ , \new_[3225]_ ,
    \new_[3226]_ , \new_[3227]_ , \new_[3228]_ , \new_[3229]_ ,
    \new_[3230]_ , \new_[3231]_ , \new_[3232]_ , \new_[3233]_ ,
    \new_[3234]_ , \new_[3235]_ , \new_[3236]_ , \new_[3237]_ ,
    \new_[3238]_ , \new_[3239]_ , \new_[3240]_ , \new_[3241]_ ,
    \new_[3242]_ , \new_[3243]_ , \new_[3244]_ , \new_[3245]_ ,
    \new_[3246]_ , \new_[3247]_ , \new_[3248]_ , \new_[3249]_ ,
    \new_[3250]_ , \new_[3251]_ , \new_[3252]_ , \new_[3253]_ ,
    \new_[3254]_ , \new_[3255]_ , \new_[3256]_ , \new_[3257]_ ,
    \new_[3258]_ , \new_[3259]_ , \new_[3260]_ , \new_[3261]_ ,
    \new_[3262]_ , \new_[3263]_ , \new_[3264]_ , \new_[3265]_ ,
    \new_[3266]_ , \new_[3267]_ , \new_[3268]_ , \new_[3269]_ ,
    \new_[3270]_ , \new_[3271]_ , \new_[3272]_ , \new_[3273]_ ,
    \new_[3274]_ , \new_[3275]_ , \new_[3276]_ , \new_[3277]_ ,
    \new_[3278]_ , \new_[3279]_ , \new_[3280]_ , \new_[3281]_ ,
    \new_[3282]_ , \new_[3283]_ , \new_[3284]_ , \new_[3285]_ ,
    \new_[3286]_ , \new_[3287]_ , \new_[3288]_ , \new_[3289]_ ,
    \new_[3290]_ , \new_[3291]_ , \new_[3292]_ , \new_[3293]_ ,
    \new_[3294]_ , \new_[3295]_ , \new_[3296]_ , \new_[3297]_ ,
    \new_[3298]_ , \new_[3299]_ , \new_[3300]_ , \new_[3301]_ ,
    \new_[3302]_ , \new_[3303]_ , \new_[3304]_ , \new_[3305]_ ,
    \new_[3306]_ , \new_[3307]_ , \new_[3308]_ , \new_[3309]_ ,
    \new_[3310]_ , \new_[3311]_ , \new_[3312]_ , \new_[3313]_ ,
    \new_[3314]_ , \new_[3315]_ , \new_[3316]_ , \new_[3317]_ ,
    \new_[3318]_ , \new_[3319]_ , \new_[3320]_ , \new_[3321]_ ,
    \new_[3322]_ , \new_[3323]_ , \new_[3324]_ , \new_[3325]_ ,
    \new_[3326]_ , \new_[3327]_ , \new_[3328]_ , \new_[3329]_ ,
    \new_[3330]_ , \new_[3331]_ , \new_[3332]_ , \new_[3333]_ ,
    \new_[3334]_ , \new_[3335]_ , \new_[3336]_ , \new_[3337]_ ,
    \new_[3338]_ , \new_[3339]_ , \new_[3340]_ , \new_[3341]_ ,
    \new_[3342]_ , \new_[3343]_ , \new_[3344]_ , \new_[3349]_ ,
    \new_[3351]_ , \new_[3353]_ , \new_[3354]_ , \new_[3357]_ ,
    \new_[3363]_ , \new_[3364]_ , \new_[3374]_ , \new_[3377]_ ,
    \new_[3404]_ , \new_[3405]_ , \new_[3406]_ , \new_[3407]_ ,
    \new_[3408]_ , \new_[3409]_ , \new_[3411]_ , \new_[3412]_ ,
    \new_[3413]_ , \new_[3414]_ , \new_[3415]_ , \new_[3448]_ ,
    \new_[3449]_ , \new_[3450]_ , \new_[3451]_ , \new_[3452]_ ,
    \new_[3453]_ , \new_[3454]_ , \new_[3455]_ , \new_[3456]_ ,
    \new_[3457]_ , \new_[3458]_ , \new_[3459]_ , \new_[3460]_ ,
    \new_[3461]_ , \new_[3462]_ , \new_[3463]_ , \new_[3464]_ ,
    \new_[3465]_ , \new_[3466]_ , \new_[3467]_ , \new_[3468]_ ,
    \new_[3469]_ , \new_[3470]_ , \new_[3471]_ , \new_[3472]_ ,
    \new_[3473]_ , \new_[3474]_ , \new_[3475]_ , \new_[3476]_ ,
    \new_[3477]_ , \new_[3478]_ , \new_[3479]_ , \new_[3480]_ ,
    \new_[3481]_ , \new_[3482]_ , \new_[3483]_ , \new_[3484]_ ,
    \new_[3485]_ , \new_[3486]_ , \new_[3487]_ , \new_[3488]_ ,
    \new_[3489]_ , \new_[3490]_ , \new_[3491]_ , \new_[3492]_ ,
    \new_[3493]_ , \new_[3494]_ , \new_[3495]_ , \new_[3496]_ ,
    \new_[3497]_ , \new_[3498]_ , \new_[3499]_ , \new_[3500]_ ,
    \new_[3501]_ , \new_[3502]_ , \new_[3503]_ , \new_[3504]_ ,
    \new_[3505]_ , \new_[3506]_ , \new_[3507]_ , \new_[3508]_ ,
    \new_[3509]_ , \new_[3510]_ , \new_[3511]_ , \new_[3512]_ ,
    \new_[3513]_ , \new_[3514]_ , \new_[3515]_ , \new_[3516]_ ,
    \new_[3517]_ , \new_[3518]_ , \new_[3519]_ , \new_[3520]_ ,
    \new_[3521]_ , \new_[3522]_ , \new_[3523]_ , \new_[3524]_ ,
    \new_[3525]_ , \new_[3527]_ , \new_[3528]_ , \new_[3529]_ ,
    \new_[3530]_ , \new_[3531]_ , \new_[3532]_ , \new_[3533]_ ,
    \new_[3534]_ , \new_[3535]_ , \new_[3536]_ , \new_[3537]_ ,
    \new_[3538]_ , \new_[3540]_ , \new_[3541]_ , \new_[3542]_ ,
    \new_[3543]_ , \new_[3544]_ , \new_[3546]_ , \new_[3547]_ ,
    \new_[3548]_ , \new_[3549]_ , \new_[3550]_ , \new_[3551]_ ,
    \new_[3552]_ , \new_[3553]_ , \new_[3554]_ , \new_[3555]_ ,
    \new_[3556]_ , \new_[3557]_ , \new_[3558]_ , \new_[3559]_ ,
    \new_[3560]_ , \new_[3561]_ , \new_[3562]_ , \new_[3563]_ ,
    \new_[3564]_ , \new_[3565]_ , \new_[3566]_ , \new_[3567]_ ,
    \new_[3568]_ , \new_[3569]_ , \new_[3570]_ , \new_[3571]_ ,
    \new_[3572]_ , \new_[3573]_ , \new_[3574]_ , \new_[3576]_ ,
    \new_[3577]_ , \new_[3578]_ , \new_[3579]_ , \new_[3581]_ ,
    \new_[3582]_ , \new_[3583]_ , \new_[3584]_ , \new_[3585]_ ,
    \new_[3586]_ , \new_[3587]_ , \new_[3588]_ , \new_[3589]_ ,
    \new_[3590]_ , \new_[3591]_ , \new_[3592]_ , \new_[3593]_ ,
    \new_[3594]_ , \new_[3595]_ , \new_[3596]_ , \new_[3597]_ ,
    \new_[3598]_ , \new_[3599]_ , \new_[3600]_ , \new_[3601]_ ,
    \new_[3602]_ , \new_[3603]_ , \new_[3604]_ , \new_[3605]_ ,
    \new_[3606]_ , \new_[3607]_ , \new_[3620]_ , \new_[3627]_ ,
    \new_[3628]_ , \new_[3629]_ , \new_[3630]_ , \new_[3634]_ ,
    \new_[3635]_ , \new_[3644]_ , \new_[3645]_ , \new_[3646]_ ,
    \new_[3647]_ , \new_[3650]_ , \new_[3657]_ , \new_[3658]_ ,
    \new_[3659]_ , \new_[3660]_ , \new_[3661]_ , \new_[3662]_ ,
    \new_[3663]_ , \new_[3665]_ , \new_[3666]_ , \new_[3667]_ ,
    \new_[3668]_ , \new_[3669]_ , \new_[3670]_ , \new_[3671]_ ,
    \new_[3672]_ , \new_[3676]_ , \new_[3677]_ , \new_[3678]_ ,
    \new_[3679]_ , \new_[3760]_ , \new_[3761]_ , \new_[3762]_ ,
    \new_[3763]_ , \new_[3764]_ , \new_[3766]_ , \new_[3771]_ ,
    \new_[3773]_ , \new_[3774]_ , \new_[3776]_ , \new_[3777]_ ,
    \new_[3778]_ , \new_[3779]_ , \new_[3780]_ , \new_[3781]_ ,
    \new_[3782]_ , \new_[3783]_ , \new_[3784]_ , \new_[3785]_ ,
    \new_[3786]_ , \new_[3787]_ , \new_[3788]_ , \new_[3789]_ ,
    \new_[3790]_ , \new_[3791]_ , \new_[3792]_ , \new_[3793]_ ,
    \new_[3798]_ , \new_[3800]_ , \new_[3801]_ , \new_[3802]_ ,
    \new_[3803]_ , \new_[3804]_ , \new_[3805]_ , \new_[3806]_ ,
    \new_[3807]_ , \new_[3808]_ , \new_[3809]_ , \new_[3810]_ ,
    \new_[3811]_ , \new_[3812]_ , \new_[3813]_ , \new_[3814]_ ,
    \new_[3815]_ , \new_[3816]_ , \new_[3817]_ , \new_[3818]_ ,
    \new_[3819]_ , \new_[3820]_ , \new_[3821]_ , \new_[3822]_ ,
    \new_[3823]_ , \new_[3824]_ , \new_[3825]_ , \new_[3826]_ ,
    \new_[3827]_ , \new_[3828]_ , \new_[3829]_ , \new_[3830]_ ,
    \new_[3831]_ , \new_[3832]_ , \new_[3833]_ , \new_[3834]_ ,
    \new_[3835]_ , \new_[3836]_ , \new_[3837]_ , \new_[3838]_ ,
    \new_[3839]_ , \new_[3840]_ , \new_[3841]_ , \new_[3843]_ ,
    \new_[3844]_ , \new_[3845]_ , \new_[3846]_ , \new_[3847]_ ,
    \new_[3848]_ , \new_[3849]_ , \new_[3850]_ , \new_[3851]_ ,
    \new_[3852]_ , \new_[3853]_ , \new_[3854]_ , \new_[3855]_ ,
    \new_[3856]_ , \new_[3857]_ , \new_[3858]_ , \new_[3859]_ ,
    \new_[3860]_ , \new_[3861]_ , \new_[3862]_ , \new_[3863]_ ,
    \new_[3864]_ , \new_[3865]_ , \new_[3866]_ , \new_[3867]_ ,
    \new_[3868]_ , \new_[3869]_ , \new_[3870]_ , \new_[3871]_ ,
    \new_[3895]_ , \new_[3897]_ , \new_[3898]_ , \new_[3899]_ ,
    \new_[3901]_ , \new_[3902]_ , \new_[3903]_ , \new_[3904]_ ,
    \new_[3905]_ , \new_[3906]_ , \new_[3908]_ , \new_[3909]_ ,
    \new_[3910]_ , \new_[3911]_ , \new_[3912]_ , \new_[3914]_ ,
    \new_[3915]_ , \new_[3917]_ , \new_[3918]_ , \new_[3921]_ ,
    \new_[3922]_ , \new_[3924]_ , \new_[3925]_ , \new_[3926]_ ,
    \new_[3928]_ , \new_[3929]_ , \new_[3930]_ , \new_[3931]_ ,
    \new_[3932]_ , \new_[3933]_ , \new_[3934]_ , \new_[3935]_ ,
    \new_[3936]_ , \new_[3938]_ , \new_[3939]_ , \new_[3940]_ ,
    \new_[3942]_ , \new_[3943]_ , \new_[3944]_ , \new_[3946]_ ,
    \new_[3947]_ , \new_[3948]_ , \new_[3950]_ , \new_[3961]_ ,
    \new_[3962]_ , \new_[3995]_ , \new_[3996]_ , \new_[3997]_ ,
    \new_[3998]_ , \new_[3999]_ , \new_[4000]_ , \new_[4001]_ ,
    \new_[4002]_ , \new_[4003]_ , \new_[4004]_ , \new_[4006]_ ,
    \new_[4007]_ , \new_[4008]_ , \new_[4009]_ , \new_[4011]_ ,
    \new_[4012]_ , \new_[4013]_ , \new_[4014]_ , \new_[4015]_ ,
    \new_[4016]_ , \new_[4017]_ , \new_[4018]_ , \new_[4019]_ ,
    \new_[4020]_ , \new_[4021]_ , \new_[4022]_ , \new_[4023]_ ,
    \new_[4024]_ , \new_[4025]_ , \new_[4026]_ , \new_[4027]_ ,
    \new_[4028]_ , \new_[4029]_ , \new_[4030]_ , \new_[4031]_ ,
    \new_[4032]_ , \new_[4033]_ , \new_[4034]_ , \new_[4035]_ ,
    \new_[4036]_ , \new_[4037]_ , \new_[4038]_ , \new_[4039]_ ,
    \new_[4040]_ , \new_[4041]_ , \new_[4042]_ , \new_[4043]_ ,
    \new_[4044]_ , \new_[4045]_ , \new_[4046]_ , \new_[4047]_ ,
    \new_[4048]_ , \new_[4049]_ , \new_[4050]_ , \new_[4051]_ ,
    \new_[4052]_ , \new_[4053]_ , \new_[4054]_ , \new_[4058]_ ,
    \new_[4059]_ , \new_[4062]_ , \new_[4063]_ , \new_[4066]_ ,
    \new_[4067]_ , \new_[4068]_ , \new_[4069]_ , \new_[4070]_ ,
    \new_[4071]_ , \new_[4072]_ , \new_[4073]_ , \new_[4074]_ ,
    \new_[4075]_ , \new_[4076]_ , \new_[4077]_ , \new_[4078]_ ,
    \new_[4079]_ , \new_[4080]_ , \new_[4081]_ , \new_[4082]_ ,
    \new_[4083]_ , \new_[4084]_ , \new_[4085]_ , \new_[4086]_ ,
    \new_[4087]_ , \new_[4088]_ , \new_[4089]_ , \new_[4144]_ ,
    \new_[4151]_ , \new_[4157]_ , \new_[4160]_ , \new_[4181]_ ,
    \new_[4182]_ , \new_[4183]_ , \new_[4185]_ , \new_[4186]_ ,
    \new_[4187]_ , \new_[4188]_ , \new_[4189]_ , \new_[4190]_ ,
    \new_[4192]_ , \new_[4194]_ , \new_[4196]_ , \new_[4197]_ ,
    \new_[4237]_ , \new_[4238]_ , \new_[4245]_ , \new_[4246]_ ,
    \new_[4247]_ , \new_[4249]_ , \new_[4277]_ , \new_[4278]_ ,
    \new_[4279]_ , \new_[4282]_ , \new_[4283]_ , \new_[4284]_ ,
    \new_[4285]_ , \new_[4286]_ , \new_[4287]_ , \new_[4288]_ ,
    \new_[4290]_ , \new_[4291]_ , \new_[4292]_ , \new_[4293]_ ,
    \new_[4294]_ , \new_[4295]_ , \new_[4296]_ , \new_[4297]_ ,
    \new_[4298]_ , \new_[4299]_ , \new_[4300]_ , \new_[4301]_ ,
    \new_[4302]_ , \new_[4303]_ , \new_[4304]_ , \new_[4305]_ ,
    \new_[4306]_ , \new_[4307]_ , \new_[4308]_ , \new_[4309]_ ,
    \new_[4310]_ , \new_[4311]_ , \new_[4312]_ , \new_[4313]_ ,
    \new_[4314]_ , \new_[4315]_ , \new_[4316]_ , \new_[4317]_ ,
    \new_[4318]_ , \new_[4319]_ , \new_[4320]_ , \new_[4321]_ ,
    \new_[4322]_ , \new_[4323]_ , \new_[4324]_ , \new_[4325]_ ,
    \new_[4326]_ , \new_[4327]_ , \new_[4328]_ , \new_[4329]_ ,
    \new_[4330]_ , \new_[4331]_ , \new_[4332]_ , \new_[4333]_ ,
    \new_[4334]_ , \new_[4335]_ , \new_[4336]_ , \new_[4337]_ ,
    \new_[4338]_ , \new_[4339]_ , \new_[4340]_ , \new_[4341]_ ,
    \new_[4342]_ , \new_[4343]_ , \new_[4344]_ , \new_[4345]_ ,
    \new_[4346]_ , \new_[4347]_ , \new_[4348]_ , \new_[4349]_ ,
    \new_[4350]_ , \new_[4351]_ , \new_[4352]_ , \new_[4353]_ ,
    \new_[4354]_ , \new_[4355]_ , \new_[4356]_ , \new_[4357]_ ,
    \new_[4358]_ , \new_[4359]_ , \new_[4360]_ , \new_[4361]_ ,
    \new_[4362]_ , \new_[4363]_ , \new_[4364]_ , \new_[4365]_ ,
    \new_[4366]_ , \new_[4367]_ , \new_[4368]_ , \new_[4369]_ ,
    \new_[4370]_ , \new_[4371]_ , \new_[4372]_ , \new_[4373]_ ,
    \new_[4374]_ , \new_[4375]_ , \new_[4376]_ , \new_[4377]_ ,
    \new_[4378]_ , \new_[4379]_ , \new_[4380]_ , \new_[4381]_ ,
    \new_[4382]_ , \new_[4383]_ , \new_[4384]_ , \new_[4385]_ ,
    \new_[4386]_ , \new_[4387]_ , \new_[4388]_ , \new_[4389]_ ,
    \new_[4390]_ , \new_[4391]_ , \new_[4392]_ , \new_[4393]_ ,
    \new_[4394]_ , \new_[4395]_ , \new_[4396]_ , \new_[4397]_ ,
    \new_[4398]_ , \new_[4406]_ , \new_[4407]_ , \new_[4408]_ ,
    \new_[4409]_ , \new_[4410]_ , \new_[4411]_ , \new_[4412]_ ,
    \new_[4413]_ , \new_[4414]_ , \new_[4415]_ , \new_[4416]_ ,
    \new_[4417]_ , \new_[4418]_ , \new_[4419]_ , \new_[4420]_ ,
    \new_[4421]_ , \new_[4422]_ , \new_[4423]_ , \new_[4424]_ ,
    \new_[4425]_ , \new_[4426]_ , \new_[4427]_ , \new_[4428]_ ,
    \new_[4429]_ , \new_[4430]_ , \new_[4431]_ , \new_[4432]_ ,
    \new_[4433]_ , \new_[4434]_ , \new_[4435]_ , \new_[4436]_ ,
    \new_[4437]_ , \new_[4438]_ , \new_[4439]_ , \new_[4440]_ ,
    \new_[4441]_ , \new_[4442]_ , \new_[4443]_ , \new_[4444]_ ,
    \new_[4445]_ , \new_[4446]_ , \new_[4447]_ , \new_[4448]_ ,
    \new_[4449]_ , \new_[4450]_ , \new_[4451]_ , \new_[4452]_ ,
    \new_[4453]_ , \new_[4454]_ , \new_[4455]_ , \new_[4456]_ ,
    \new_[4457]_ , \new_[4458]_ , \new_[4459]_ , \new_[4460]_ ,
    \new_[4461]_ , \new_[4462]_ , \new_[4463]_ , \new_[4464]_ ,
    \new_[4465]_ , \new_[4468]_ , \new_[4469]_ , \new_[4470]_ ,
    \new_[4471]_ , \new_[4472]_ , \new_[4473]_ , \new_[4474]_ ,
    \new_[4475]_ , \new_[4476]_ , \new_[4477]_ , \new_[4478]_ ,
    \new_[4495]_ , \new_[4496]_ , \new_[4503]_ , \new_[4504]_ ,
    \new_[4505]_ , \new_[4506]_ , \new_[4507]_ , \new_[4508]_ ,
    \new_[4509]_ , \new_[4511]_ , \new_[4512]_ , \new_[4513]_ ,
    \new_[4514]_ , \new_[4515]_ , \new_[4516]_ , \new_[4517]_ ,
    \new_[4518]_ , \new_[4519]_ , \new_[4520]_ , \new_[4521]_ ,
    \new_[4522]_ , \new_[4523]_ , \new_[4524]_ , \new_[4525]_ ,
    \new_[4526]_ , \new_[4527]_ , \new_[4528]_ , \new_[4529]_ ,
    \new_[4530]_ , \new_[4531]_ , \new_[4532]_ , \new_[4533]_ ,
    \new_[4534]_ , \new_[4535]_ , \new_[4536]_ , \new_[4537]_ ,
    \new_[4538]_ , \new_[4539]_ , \new_[4540]_ , \new_[4541]_ ,
    \new_[4542]_ , \new_[4543]_ , \new_[4545]_ , \new_[4546]_ ,
    \new_[4564]_ , \new_[4565]_ , \new_[4572]_ , \new_[4574]_ ,
    \new_[4575]_ , \new_[4576]_ , \new_[4577]_ , \new_[4578]_ ,
    \new_[4579]_ , \new_[4580]_ , \new_[4581]_ , \new_[4582]_ ,
    \new_[4583]_ , \new_[4584]_ , \new_[4585]_ , \new_[4586]_ ,
    \new_[4587]_ , \new_[4588]_ , \new_[4589]_ , \new_[4590]_ ,
    \new_[4591]_ , \new_[4592]_ , \new_[4593]_ , \new_[4594]_ ,
    \new_[4595]_ , \new_[4596]_ , \new_[4597]_ , \new_[4598]_ ,
    \new_[4599]_ , \new_[4600]_ , \new_[4601]_ , \new_[4602]_ ,
    \new_[4603]_ , \new_[4604]_ , \new_[4605]_ , \new_[4606]_ ,
    \new_[4607]_ , \new_[4608]_ , \new_[4609]_ , \new_[4610]_ ,
    \new_[4611]_ , \new_[4612]_ , \new_[4613]_ , \new_[4614]_ ,
    \new_[4615]_ , \new_[4616]_ , \new_[4618]_ , \new_[4619]_ ,
    \new_[4620]_ , \new_[4621]_ , \new_[4622]_ , \new_[4623]_ ,
    \new_[4624]_ , \new_[4625]_ , \new_[4626]_ , \new_[4627]_ ,
    \new_[4628]_ , \new_[4629]_ , \new_[4631]_ , \new_[4632]_ ,
    \new_[4633]_ , \new_[4634]_ , \new_[4635]_ , \new_[4636]_ ,
    \new_[4637]_ , \new_[4638]_ , \new_[4639]_ , \new_[4640]_ ,
    \new_[4641]_ , \new_[4642]_ , \new_[4644]_ , \new_[4645]_ ,
    \new_[4646]_ , \new_[4647]_ , \new_[4648]_ , \new_[4649]_ ,
    \new_[4650]_ , \new_[4651]_ , \new_[4652]_ , \new_[4653]_ ,
    \new_[4654]_ , \new_[4655]_ , \new_[4656]_ , \new_[4657]_ ,
    \new_[4658]_ , \new_[4659]_ , \new_[4660]_ , \new_[4661]_ ,
    \new_[4662]_ , \new_[4663]_ , \new_[4664]_ , \new_[4665]_ ,
    \new_[4666]_ , \new_[4667]_ , \new_[4668]_ , \new_[4669]_ ,
    \new_[4670]_ , \new_[4671]_ , \new_[4672]_ , \new_[4673]_ ,
    \new_[4674]_ , \new_[4675]_ , \new_[4676]_ , \new_[4677]_ ,
    \new_[4678]_ , \new_[4679]_ , \new_[4680]_ , \new_[4681]_ ,
    \new_[4682]_ , \new_[4683]_ , \new_[4684]_ , \new_[4685]_ ,
    \new_[4686]_ , \new_[4687]_ , \new_[4688]_ , \new_[4689]_ ,
    \new_[4690]_ , \new_[4691]_ , \new_[4692]_ , \new_[4693]_ ,
    \new_[4694]_ , \new_[4695]_ , \new_[4696]_ , \new_[4703]_ ,
    \new_[4704]_ , \new_[4705]_ , \new_[4706]_ , \new_[4707]_ ,
    \new_[4708]_ , \new_[4709]_ , \new_[4713]_ , \new_[4715]_ ,
    \new_[4716]_ , \new_[4717]_ , \new_[4720]_ , \new_[4722]_ ,
    \new_[4723]_ , \new_[4724]_ , \new_[4725]_ , \new_[4728]_ ,
    \new_[4730]_ , \new_[4731]_ , \new_[4733]_ , \new_[4734]_ ,
    \new_[4735]_ , \new_[4736]_ , \new_[4743]_ , \new_[4744]_ ,
    \new_[4745]_ , \new_[4746]_ , \new_[4747]_ , \new_[4748]_ ,
    \new_[4749]_ , \new_[4750]_ , \new_[4752]_ , \new_[4753]_ ,
    \new_[4754]_ , \new_[4755]_ , \new_[4756]_ , \new_[4757]_ ,
    \new_[4758]_ , \new_[4759]_ , \new_[4760]_ , \new_[4761]_ ,
    \new_[4762]_ , \new_[4763]_ , \new_[4764]_ , \new_[4765]_ ,
    \new_[4766]_ , \new_[4767]_ , \new_[4768]_ , \new_[4775]_ ,
    \new_[4776]_ , \new_[4777]_ , \new_[4778]_ , \new_[4779]_ ,
    \new_[4780]_ , \new_[4781]_ , \new_[4782]_ , \new_[4783]_ ,
    \new_[4784]_ , \new_[4785]_ , \new_[4786]_ , \new_[4787]_ ,
    \new_[4788]_ , \new_[4789]_ , \new_[4790]_ , \new_[4791]_ ,
    \new_[4792]_ , \new_[4793]_ , \new_[4806]_ , \new_[4807]_ ,
    \new_[4808]_ , \new_[4809]_ , \new_[4810]_ , \new_[4811]_ ,
    \new_[4812]_ , \new_[4813]_ , \new_[4814]_ , \new_[4815]_ ,
    \new_[4816]_ , \new_[4817]_ , \new_[4818]_ , \new_[4819]_ ,
    \new_[4820]_ , \new_[4821]_ , \new_[4822]_ , \new_[4823]_ ,
    \new_[4824]_ , \new_[4825]_ , \new_[4826]_ , \new_[4827]_ ,
    \new_[4828]_ , \new_[4829]_ , \new_[4830]_ , \new_[4831]_ ,
    \new_[4832]_ , \new_[4833]_ , \new_[4834]_ , \new_[4835]_ ,
    \new_[4836]_ , \new_[4837]_ , \new_[4838]_ , \new_[4839]_ ,
    \new_[4840]_ , \new_[4841]_ , \new_[4842]_ , \new_[4843]_ ,
    \new_[4844]_ , \new_[4845]_ , \new_[4846]_ , \new_[4847]_ ,
    \new_[4848]_ , \new_[4849]_ , \new_[4850]_ , \new_[4851]_ ,
    \new_[4852]_ , \new_[4853]_ , \new_[4854]_ , \new_[4855]_ ,
    \new_[4856]_ , \new_[4857]_ , \new_[4858]_ , \new_[4859]_ ,
    \new_[4860]_ , \new_[4861]_ , \new_[4862]_ , \new_[4863]_ ,
    \new_[4864]_ , \new_[4865]_ , \new_[4866]_ , \new_[4867]_ ,
    \new_[4868]_ , \new_[4869]_ , \new_[4870]_ , \new_[4871]_ ,
    \new_[4872]_ , \new_[4873]_ , \new_[4874]_ , \new_[4875]_ ,
    \new_[4876]_ , \new_[4877]_ , \new_[4879]_ , \new_[4885]_ ,
    \new_[4886]_ , \new_[4887]_ , \new_[4888]_ , \new_[4889]_ ,
    \new_[4890]_ , \new_[4891]_ , \new_[4892]_ , \new_[4893]_ ,
    \new_[4894]_ , \new_[4895]_ , \new_[4896]_ , \new_[4897]_ ,
    \new_[4898]_ , \new_[4899]_ , \new_[4900]_ , \new_[4901]_ ,
    \new_[4902]_ , \new_[4903]_ , \new_[4904]_ , \new_[4905]_ ,
    \new_[4906]_ , \new_[4907]_ , \new_[4908]_ , \new_[4909]_ ,
    \new_[4910]_ , \new_[4911]_ , \new_[4912]_ , \new_[4913]_ ,
    \new_[4914]_ , \new_[4915]_ , \new_[4916]_ , \new_[4917]_ ,
    \new_[4918]_ , \new_[4919]_ , \new_[4920]_ , \new_[4921]_ ,
    \new_[4922]_ , \new_[4923]_ , \new_[4924]_ , \new_[4925]_ ,
    \new_[4926]_ , \new_[4927]_ , \new_[4928]_ , \new_[4929]_ ,
    \new_[4930]_ , \new_[4931]_ , \new_[4932]_ , \new_[4934]_ ,
    \new_[4935]_ , \new_[4936]_ , \new_[4937]_ , \new_[4938]_ ,
    \new_[4941]_ , \new_[4942]_ , \new_[4943]_ , \new_[4945]_ ,
    \new_[4946]_ , \new_[4947]_ , \new_[4948]_ , \new_[4949]_ ,
    \new_[4950]_ , \new_[4951]_ , \new_[4952]_ , \new_[4953]_ ,
    \new_[4954]_ , \new_[4956]_ , \new_[4957]_ , \new_[4959]_ ,
    \new_[4960]_ , \new_[4961]_ , \new_[4962]_ , \new_[4963]_ ,
    \new_[4964]_ , \new_[4965]_ , \new_[4966]_ , \new_[4967]_ ,
    \new_[4968]_ , \new_[4969]_ , \new_[4970]_ , \new_[4971]_ ,
    \new_[4972]_ , \new_[4973]_ , \new_[4974]_ , \new_[4975]_ ,
    \new_[4976]_ , \new_[4977]_ , \new_[4978]_ , \new_[4979]_ ,
    \new_[4980]_ , \new_[4981]_ , \new_[4982]_ , \new_[4983]_ ,
    \new_[4984]_ , \new_[4985]_ , \new_[4986]_ , \new_[4987]_ ,
    \new_[4988]_ , \new_[4989]_ , \new_[4990]_ , \new_[4991]_ ,
    \new_[4992]_ , \new_[4993]_ , \new_[4994]_ , \new_[4995]_ ,
    \new_[4996]_ , \new_[4997]_ , \new_[4998]_ , \new_[4999]_ ,
    \new_[5000]_ , \new_[5001]_ , \new_[5002]_ , \new_[5003]_ ,
    \new_[5004]_ , \new_[5005]_ , \new_[5006]_ , \new_[5007]_ ,
    \new_[5008]_ , \new_[5009]_ , \new_[5010]_ , \new_[5011]_ ,
    \new_[5012]_ , \new_[5013]_ , \new_[5014]_ , \new_[5015]_ ,
    \new_[5016]_ , \new_[5017]_ , \new_[5018]_ , \new_[5019]_ ,
    \new_[5020]_ , \new_[5021]_ , \new_[5022]_ , \new_[5023]_ ,
    \new_[5024]_ , \new_[5025]_ , \new_[5026]_ , \new_[5027]_ ,
    \new_[5028]_ , \new_[5029]_ , \new_[5030]_ , \new_[5031]_ ,
    \new_[5032]_ , \new_[5033]_ , \new_[5034]_ , \new_[5035]_ ,
    \new_[5036]_ , \new_[5037]_ , \new_[5038]_ , \new_[5039]_ ,
    \new_[5040]_ , \new_[5041]_ , \new_[5042]_ , \new_[5043]_ ,
    \new_[5044]_ , \new_[5045]_ , \new_[5046]_ , \new_[5047]_ ,
    \new_[5048]_ , \new_[5049]_ , \new_[5050]_ , \new_[5051]_ ,
    \new_[5052]_ , \new_[5053]_ , \new_[5054]_ , \new_[5055]_ ,
    \new_[5056]_ , \new_[5057]_ , \new_[5058]_ , \new_[5059]_ ,
    \new_[5060]_ , \new_[5061]_ , \new_[5062]_ , \new_[5063]_ ,
    \new_[5064]_ , \new_[5065]_ , \new_[5066]_ , \new_[5067]_ ,
    \new_[5068]_ , \new_[5069]_ , \new_[5070]_ , \new_[5071]_ ,
    \new_[5072]_ , \new_[5073]_ , \new_[5074]_ , \new_[5075]_ ,
    \new_[5076]_ , \new_[5077]_ , \new_[5078]_ , \new_[5079]_ ,
    \new_[5080]_ , \new_[5081]_ , \new_[5082]_ , \new_[5083]_ ,
    \new_[5084]_ , \new_[5085]_ , \new_[5086]_ , \new_[5087]_ ,
    \new_[5088]_ , \new_[5089]_ , \new_[5090]_ , \new_[5091]_ ,
    \new_[5092]_ , \new_[5093]_ , \new_[5094]_ , \new_[5095]_ ,
    \new_[5096]_ , \new_[5097]_ , \new_[5098]_ , \new_[5099]_ ,
    \new_[5100]_ , \new_[5101]_ , \new_[5102]_ , \new_[5103]_ ,
    \new_[5104]_ , \new_[5105]_ , \new_[5106]_ , \new_[5107]_ ,
    \new_[5108]_ , \new_[5109]_ , \new_[5110]_ , \new_[5111]_ ,
    \new_[5112]_ , \new_[5113]_ , \new_[5114]_ , \new_[5115]_ ,
    \new_[5116]_ , \new_[5117]_ , \new_[5118]_ , \new_[5119]_ ,
    \new_[5120]_ , \new_[5121]_ , \new_[5122]_ , \new_[5123]_ ,
    \new_[5124]_ , \new_[5125]_ , \new_[5126]_ , \new_[5127]_ ,
    \new_[5128]_ , \new_[5129]_ , \new_[5130]_ , \new_[5131]_ ,
    \new_[5132]_ , \new_[5133]_ , \new_[5134]_ , \new_[5135]_ ,
    \new_[5136]_ , \new_[5137]_ , \new_[5138]_ , \new_[5139]_ ,
    \new_[5140]_ , \new_[5141]_ , \new_[5142]_ , \new_[5143]_ ,
    \new_[5144]_ , \new_[5145]_ , \new_[5146]_ , \new_[5147]_ ,
    \new_[5148]_ , \new_[5149]_ , \new_[5150]_ , \new_[5151]_ ,
    \new_[5152]_ , \new_[5153]_ , \new_[5154]_ , \new_[5155]_ ,
    \new_[5156]_ , \new_[5157]_ , \new_[5158]_ , \new_[5159]_ ,
    \new_[5160]_ , \new_[5161]_ , \new_[5162]_ , \new_[5163]_ ,
    \new_[5164]_ , \new_[5165]_ , \new_[5166]_ , \new_[5167]_ ,
    \new_[5168]_ , \new_[5169]_ , \new_[5170]_ , \new_[5171]_ ,
    \new_[5172]_ , \new_[5173]_ , \new_[5174]_ , \new_[5175]_ ,
    \new_[5176]_ , \new_[5177]_ , \new_[5178]_ , \new_[5179]_ ,
    \new_[5180]_ , \new_[5181]_ , \new_[5182]_ , \new_[5183]_ ,
    \new_[5184]_ , \new_[5185]_ , \new_[5186]_ , \new_[5187]_ ,
    \new_[5188]_ , \new_[5189]_ , \new_[5190]_ , \new_[5191]_ ,
    \new_[5192]_ , \new_[5193]_ , \new_[5194]_ , \new_[5195]_ ,
    \new_[5196]_ , \new_[5197]_ , \new_[5198]_ , \new_[5199]_ ,
    \new_[5200]_ , \new_[5201]_ , \new_[5202]_ , \new_[5203]_ ,
    \new_[5204]_ , \new_[5205]_ , \new_[5206]_ , \new_[5207]_ ,
    \new_[5208]_ , \new_[5209]_ , \new_[5210]_ , \new_[5211]_ ,
    \new_[5212]_ , \new_[5213]_ , \new_[5214]_ , \new_[5215]_ ,
    \new_[5216]_ , \new_[5217]_ , \new_[5218]_ , \new_[5219]_ ,
    \new_[5220]_ , \new_[5221]_ , \new_[5222]_ , \new_[5223]_ ,
    \new_[5224]_ , \new_[5225]_ , \new_[5226]_ , \new_[5227]_ ,
    \new_[5228]_ , \new_[5229]_ , \new_[5230]_ , \new_[5231]_ ,
    \new_[5232]_ , \new_[5233]_ , \new_[5234]_ , \new_[5235]_ ,
    \new_[5236]_ , \new_[5237]_ , \new_[5238]_ , \new_[5239]_ ,
    \new_[5240]_ , \new_[5241]_ , \new_[5242]_ , \new_[5243]_ ,
    \new_[5244]_ , \new_[5245]_ , \new_[5246]_ , \new_[5247]_ ,
    \new_[5248]_ , \new_[5249]_ , \new_[5250]_ , \new_[5251]_ ,
    \new_[5252]_ , \new_[5253]_ , \new_[5254]_ , \new_[5255]_ ,
    \new_[5256]_ , \new_[5257]_ , \new_[5258]_ , \new_[5259]_ ,
    \new_[5260]_ , \new_[5261]_ , \new_[5262]_ , \new_[5263]_ ,
    \new_[5264]_ , \new_[5265]_ , \new_[5266]_ , \new_[5267]_ ,
    \new_[5268]_ , \new_[5269]_ , \new_[5270]_ , \new_[5271]_ ,
    \new_[5272]_ , \new_[5273]_ , \new_[5274]_ , \new_[5275]_ ,
    \new_[5276]_ , \new_[5277]_ , \new_[5278]_ , \new_[5279]_ ,
    \new_[5280]_ , \new_[5281]_ , \new_[5282]_ , \new_[5283]_ ,
    \new_[5284]_ , \new_[5285]_ , \new_[5286]_ , \new_[5287]_ ,
    \new_[5288]_ , \new_[5289]_ , \new_[5290]_ , \new_[5291]_ ,
    \new_[5292]_ , \new_[5293]_ , \new_[5294]_ , \new_[5295]_ ,
    \new_[5296]_ , \new_[5297]_ , \new_[5298]_ , \new_[5299]_ ,
    \new_[5300]_ , \new_[5301]_ , \new_[5302]_ , \new_[5303]_ ,
    \new_[5304]_ , \new_[5305]_ , \new_[5306]_ , \new_[5307]_ ,
    \new_[5308]_ , \new_[5309]_ , \new_[5310]_ , \new_[5311]_ ,
    \new_[5312]_ , \new_[5313]_ , \new_[5314]_ , \new_[5315]_ ,
    \new_[5316]_ , \new_[5317]_ , \new_[5318]_ , \new_[5319]_ ,
    \new_[5320]_ , \new_[5321]_ , \new_[5322]_ , \new_[5323]_ ,
    \new_[5324]_ , \new_[5325]_ , \new_[5326]_ , \new_[5327]_ ,
    \new_[5328]_ , \new_[5329]_ , \new_[5330]_ , \new_[5331]_ ,
    \new_[5332]_ , \new_[5333]_ , \new_[5334]_ , \new_[5335]_ ,
    \new_[5336]_ , \new_[5337]_ , \new_[5338]_ , \new_[5339]_ ,
    \new_[5340]_ , \new_[5341]_ , \new_[5342]_ , \new_[5343]_ ,
    \new_[5344]_ , \new_[5345]_ , \new_[5346]_ , \new_[5347]_ ,
    \new_[5348]_ , \new_[5349]_ , \new_[5350]_ , \new_[5351]_ ,
    \new_[5352]_ , \new_[5353]_ , \new_[5354]_ , \new_[5355]_ ,
    \new_[5356]_ , \new_[5357]_ , \new_[5358]_ , \new_[5359]_ ,
    \new_[5360]_ , \new_[5361]_ , \new_[5362]_ , \new_[5363]_ ,
    \new_[5364]_ , \new_[5365]_ , \new_[5366]_ , \new_[5367]_ ,
    \new_[5368]_ , \new_[5369]_ , \new_[5370]_ , \new_[5371]_ ,
    \new_[5372]_ , \new_[5373]_ , \new_[5374]_ , \new_[5375]_ ,
    \new_[5376]_ , \new_[5377]_ , \new_[5378]_ , \new_[5379]_ ,
    \new_[5380]_ , \new_[5381]_ , \new_[5382]_ , \new_[5383]_ ,
    \new_[5384]_ , \new_[5385]_ , \new_[5386]_ , \new_[5387]_ ,
    \new_[5388]_ , \new_[5389]_ , \new_[5390]_ , \new_[5391]_ ,
    \new_[5392]_ , \new_[5393]_ , \new_[5394]_ , \new_[5395]_ ,
    \new_[5396]_ , \new_[5397]_ , \new_[5398]_ , \new_[5399]_ ,
    \new_[5400]_ , \new_[5401]_ , \new_[5402]_ , \new_[5403]_ ,
    \new_[5404]_ , \new_[5405]_ , \new_[5406]_ , \new_[5407]_ ,
    \new_[5408]_ , \new_[5409]_ , \new_[5410]_ , \new_[5411]_ ,
    \new_[5412]_ , \new_[5413]_ , \new_[5414]_ , \new_[5415]_ ,
    \new_[5416]_ , \new_[5417]_ , \new_[5418]_ , \new_[5419]_ ,
    \new_[5420]_ , \new_[5421]_ , \new_[5422]_ , \new_[5423]_ ,
    \new_[5424]_ , \new_[5425]_ , \new_[5426]_ , \new_[5427]_ ,
    \new_[5428]_ , \new_[5429]_ , \new_[5430]_ , \new_[5431]_ ,
    \new_[5432]_ , \new_[5433]_ , \new_[5434]_ , \new_[5435]_ ,
    \new_[5436]_ , \new_[5437]_ , \new_[5438]_ , \new_[5439]_ ,
    \new_[5440]_ , \new_[5441]_ , \new_[5442]_ , \new_[5443]_ ,
    \new_[5444]_ , \new_[5445]_ , \new_[5446]_ , \new_[5447]_ ,
    \new_[5448]_ , \new_[5449]_ , \new_[5450]_ , \new_[5451]_ ,
    \new_[5452]_ , \new_[5453]_ , \new_[5454]_ , \new_[5455]_ ,
    \new_[5456]_ , \new_[5457]_ , \new_[5458]_ , \new_[5459]_ ,
    \new_[5460]_ , \new_[5461]_ , \new_[5462]_ , \new_[5463]_ ,
    \new_[5464]_ , \new_[5465]_ , \new_[5466]_ , \new_[5467]_ ,
    \new_[5468]_ , \new_[5469]_ , \new_[5470]_ , \new_[5471]_ ,
    \new_[5472]_ , \new_[5473]_ , \new_[5474]_ , \new_[5475]_ ,
    \new_[5476]_ , \new_[5477]_ , \new_[5478]_ , \new_[5479]_ ,
    \new_[5480]_ , \new_[5481]_ , \new_[5482]_ , \new_[5483]_ ,
    \new_[5484]_ , \new_[5485]_ , \new_[5486]_ , \new_[5487]_ ,
    \new_[5488]_ , \new_[5489]_ , \new_[5490]_ , \new_[5491]_ ,
    \new_[5492]_ , \new_[5493]_ , \new_[5494]_ , \new_[5495]_ ,
    \new_[5496]_ , \new_[5497]_ , \new_[5498]_ , \new_[5499]_ ,
    \new_[5500]_ , \new_[5501]_ , \new_[5502]_ , \new_[5503]_ ,
    \new_[5504]_ , \new_[5505]_ , \new_[5506]_ , \new_[5507]_ ,
    \new_[5508]_ , \new_[5509]_ , \new_[5510]_ , \new_[5511]_ ,
    \new_[5512]_ , \new_[5513]_ , \new_[5514]_ , \new_[5515]_ ,
    \new_[5516]_ , \new_[5517]_ , \new_[5518]_ , \new_[5519]_ ,
    \new_[5520]_ , \new_[5521]_ , \new_[5522]_ , \new_[5523]_ ,
    \new_[5524]_ , \new_[5525]_ , \new_[5526]_ , \new_[5527]_ ,
    \new_[5528]_ , \new_[5529]_ , \new_[5530]_ , \new_[5531]_ ,
    \new_[5532]_ , \new_[5533]_ , \new_[5534]_ , \new_[5535]_ ,
    \new_[5536]_ , \new_[5537]_ , \new_[5538]_ , \new_[5539]_ ,
    \new_[5540]_ , \new_[5541]_ , \new_[5542]_ , \new_[5543]_ ,
    \new_[5544]_ , \new_[5545]_ , \new_[5546]_ , \new_[5547]_ ,
    \new_[5548]_ , \new_[5549]_ , \new_[5550]_ , \new_[5551]_ ,
    \new_[5552]_ , \new_[5553]_ , \new_[5554]_ , \new_[5555]_ ,
    \new_[5556]_ , \new_[5557]_ , \new_[5558]_ , \new_[5559]_ ,
    \new_[5560]_ , \new_[5561]_ , \new_[5562]_ , \new_[5563]_ ,
    \new_[5564]_ , \new_[5565]_ , \new_[5566]_ , \new_[5567]_ ,
    \new_[5568]_ , \new_[5569]_ , \new_[5570]_ , \new_[5571]_ ,
    \new_[5572]_ , \new_[5573]_ , \new_[5574]_ , \new_[5575]_ ,
    \new_[5576]_ , \new_[5577]_ , \new_[5578]_ , \new_[5579]_ ,
    \new_[5580]_ , \new_[5581]_ , \new_[5582]_ , \new_[5583]_ ,
    \new_[5584]_ , \new_[5585]_ , \new_[5586]_ , \new_[5587]_ ,
    \new_[5588]_ , \new_[5589]_ , \new_[5590]_ , \new_[5591]_ ,
    \new_[5592]_ , \new_[5593]_ , \new_[5594]_ , \new_[5595]_ ,
    \new_[5596]_ , \new_[5597]_ , \new_[5598]_ , \new_[5599]_ ,
    \new_[5600]_ , \new_[5601]_ , \new_[5602]_ , \new_[5603]_ ,
    \new_[5604]_ , \new_[5605]_ , \new_[5606]_ , \new_[5607]_ ,
    \new_[5608]_ , \new_[5609]_ , \new_[5610]_ , \new_[5611]_ ,
    \new_[5612]_ , \new_[5613]_ , \new_[5614]_ , \new_[5615]_ ,
    \new_[5616]_ , \new_[5617]_ , \new_[5618]_ , \new_[5619]_ ,
    \new_[5620]_ , \new_[5621]_ , \new_[5622]_ , \new_[5623]_ ,
    \new_[5624]_ , \new_[5625]_ , \new_[5626]_ , \new_[5627]_ ,
    \new_[5628]_ , \new_[5629]_ , \new_[5630]_ , \new_[5631]_ ,
    \new_[5632]_ , \new_[5633]_ , \new_[5634]_ , \new_[5635]_ ,
    \new_[5636]_ , \new_[5637]_ , \new_[5638]_ , \new_[5639]_ ,
    \new_[5640]_ , \new_[5641]_ , \new_[5642]_ , \new_[5643]_ ,
    \new_[5644]_ , \new_[5645]_ , \new_[5646]_ , \new_[5647]_ ,
    \new_[5648]_ , \new_[5649]_ , \new_[5650]_ , \new_[5651]_ ,
    \new_[5652]_ , \new_[5653]_ , \new_[5654]_ , \new_[5655]_ ,
    \new_[5656]_ , \new_[5657]_ , \new_[5658]_ , \new_[5659]_ ,
    \new_[5660]_ , \new_[5661]_ , \new_[5662]_ , \new_[5663]_ ,
    \new_[5664]_ , \new_[5665]_ , \new_[5666]_ , \new_[5667]_ ,
    \new_[5668]_ , \new_[5669]_ , \new_[5670]_ , \new_[5671]_ ,
    \new_[5672]_ , \new_[5673]_ , \new_[5674]_ , \new_[5675]_ ,
    \new_[5676]_ , \new_[5677]_ , \new_[5678]_ , \new_[5686]_ ,
    \new_[5687]_ , \new_[5688]_ , \new_[5689]_ , \new_[5690]_ ,
    \new_[5691]_ , \new_[5692]_ , \new_[5693]_ , \new_[5694]_ ,
    \new_[5695]_ , \new_[5696]_ , \new_[5697]_ , \new_[5701]_ ,
    \new_[5702]_ , \new_[5703]_ , \new_[5704]_ , \new_[5705]_ ,
    \new_[5708]_ , \new_[5713]_ , \new_[5714]_ , \new_[5715]_ ,
    \new_[5716]_ , \new_[5717]_ , \new_[5718]_ , \new_[5719]_ ,
    \new_[5720]_ , \new_[5721]_ , \new_[5722]_ , \new_[5723]_ ,
    \new_[5724]_ , \new_[5725]_ , \new_[5726]_ , \new_[5727]_ ,
    \new_[5728]_ , \new_[5729]_ , \new_[5730]_ , \new_[5731]_ ,
    \new_[5732]_ , \new_[5733]_ , \new_[5734]_ , \new_[5735]_ ,
    \new_[5736]_ , \new_[5737]_ , \new_[5738]_ , \new_[5739]_ ,
    \new_[5740]_ , \new_[5741]_ , \new_[5742]_ , \new_[5743]_ ,
    \new_[5744]_ , \new_[5745]_ , \new_[5746]_ , \new_[5747]_ ,
    \new_[5748]_ , \new_[5749]_ , \new_[5750]_ , \new_[5751]_ ,
    \new_[5752]_ , \new_[5753]_ , \new_[5754]_ , \new_[5755]_ ,
    \new_[5756]_ , \new_[5757]_ , \new_[5758]_ , \new_[5759]_ ,
    \new_[5760]_ , \new_[5761]_ , \new_[5762]_ , \new_[5763]_ ,
    \new_[5764]_ , \new_[5765]_ , \new_[5766]_ , \new_[5767]_ ,
    \new_[5768]_ , \new_[5769]_ , \new_[5777]_ , \new_[5831]_ ,
    \new_[5832]_ , \new_[5833]_ , \new_[5834]_ , \new_[5835]_ ,
    \new_[5836]_ , \new_[5837]_ , \new_[5841]_ , \new_[5842]_ ,
    \new_[5843]_ , \new_[5844]_ , \new_[5845]_ , \new_[5846]_ ,
    \new_[5847]_ , \new_[5848]_ , \new_[5849]_ , \new_[5850]_ ,
    \new_[5851]_ , \new_[5852]_ , \new_[5853]_ , \new_[5854]_ ,
    \new_[5855]_ , \new_[5856]_ , \new_[5857]_ , \new_[5858]_ ,
    \new_[5859]_ , \new_[5860]_ , \new_[5873]_ , \new_[5874]_ ,
    \new_[5875]_ , \new_[5876]_ , \new_[5877]_ , \new_[5878]_ ,
    \new_[5879]_ , \new_[5880]_ , \new_[5886]_ , \new_[5887]_ ,
    \new_[5888]_ , \new_[6237]_ , \new_[6241]_ , \new_[6289]_ ,
    \new_[6292]_ , \new_[6421]_ , \new_[6422]_ , \new_[6423]_ ,
    \new_[6424]_ , \new_[6425]_ , \new_[6426]_ , \new_[6427]_ ,
    \new_[6429]_ , \new_[6431]_ , \new_[6433]_ , \new_[6435]_ ,
    \new_[6437]_ , \new_[6439]_ , \new_[6440]_ , \new_[6441]_ ,
    \new_[6442]_ , \new_[6443]_ , \new_[6444]_ , \new_[6445]_ ,
    \new_[6446]_ , \new_[6447]_ , \new_[6448]_ , \new_[6449]_ ,
    \new_[6450]_ , \new_[6560]_ , \new_[6561]_ , \new_[6562]_ ,
    \new_[6564]_ , \new_[6565]_ , \new_[6566]_ , \new_[6567]_ ,
    \new_[6568]_ , \new_[6569]_ , \new_[6570]_ , \new_[6571]_ ,
    \new_[6572]_ , \new_[6573]_ , \new_[6759]_ , \new_[6760]_ ,
    \new_[6765]_ , \new_[6777]_ , \new_[6778]_ , \new_[6779]_ ,
    \new_[6780]_ , \new_[6785]_ , \new_[6786]_ , \new_[6787]_ ,
    \new_[6788]_ , \new_[6789]_ , \new_[6791]_ , \new_[6792]_ ,
    \new_[6793]_ , \new_[6794]_ , \new_[6809]_ , \new_[6810]_ ,
    \new_[6812]_ , \new_[6829]_ , \new_[6830]_ , \new_[6831]_ ,
    \new_[6832]_ , \new_[6833]_ , \new_[6834]_ , \new_[6835]_ ,
    \new_[6836]_ , \new_[6837]_ , \new_[6838]_ , \new_[6839]_ ,
    \new_[6840]_ , \new_[6841]_ , \new_[6843]_ , \new_[6844]_ ,
    \new_[6845]_ , \new_[6846]_ , \new_[6847]_ , \new_[6848]_ ,
    \new_[6849]_ , \new_[6850]_ , \new_[6851]_ , \new_[6852]_ ,
    \new_[6853]_ , \new_[6854]_ , \new_[6855]_ , \new_[6856]_ ,
    \new_[6857]_ , \new_[6858]_ , \new_[6859]_ , \new_[6860]_ ,
    \new_[6861]_ , \new_[6862]_ , \new_[6863]_ , \new_[6864]_ ,
    \new_[6865]_ , \new_[6866]_ , \new_[6867]_ , \new_[6868]_ ,
    \new_[6869]_ , \new_[6870]_ , \new_[6871]_ , \new_[6872]_ ,
    \new_[6873]_ , \new_[6874]_ , \new_[6875]_ , \new_[6876]_ ,
    \new_[6877]_ , \new_[6878]_ , \new_[6879]_ , \new_[6880]_ ,
    \new_[6881]_ , \new_[6882]_ , \new_[6883]_ , \new_[6884]_ ,
    \new_[6885]_ , \new_[6886]_ , \new_[6887]_ , \new_[6888]_ ,
    \new_[6889]_ , \new_[6890]_ , \new_[6891]_ , \new_[6892]_ ,
    \new_[6893]_ , \new_[6894]_ , \new_[6895]_ , \new_[6896]_ ,
    \new_[6897]_ , \new_[6898]_ , \new_[6899]_ , \new_[6900]_ ,
    \new_[6901]_ , \new_[6902]_ , \new_[6903]_ , \new_[6904]_ ,
    \new_[6905]_ , \new_[6906]_ , \new_[6907]_ , \new_[6908]_ ,
    \new_[6909]_ , \new_[6910]_ , \new_[6911]_ , \new_[6912]_ ,
    \new_[6913]_ , \new_[6914]_ , \new_[6915]_ , \new_[6916]_ ,
    \new_[6917]_ , \new_[6918]_ , \new_[6919]_ , \new_[6920]_ ,
    \new_[6921]_ , \new_[6922]_ , \new_[6923]_ , \new_[6924]_ ,
    \new_[6925]_ , \new_[6926]_ , \new_[6927]_ , \new_[6928]_ ,
    \new_[6929]_ , \new_[6930]_ , \new_[6931]_ , \new_[6932]_ ,
    \new_[6933]_ , \new_[6934]_ , \new_[6935]_ , \new_[6936]_ ,
    \new_[6937]_ , \new_[6938]_ , \new_[6939]_ , \new_[6940]_ ,
    \new_[6941]_ , \new_[6942]_ , \new_[6943]_ , \new_[6944]_ ,
    \new_[6945]_ , \new_[6946]_ , \new_[6947]_ , \new_[6948]_ ,
    \new_[6949]_ , \new_[6950]_ , \new_[6951]_ , \new_[6952]_ ,
    \new_[6953]_ , \new_[6954]_ , \new_[6955]_ , \new_[6956]_ ,
    \new_[6957]_ , \new_[6958]_ , \new_[6959]_ , \new_[6960]_ ,
    \new_[6961]_ , \new_[6962]_ , \new_[6963]_ , \new_[6964]_ ,
    \new_[6965]_ , \new_[6966]_ , \new_[6967]_ , \new_[6968]_ ,
    \new_[6969]_ , \new_[6970]_ , \new_[6971]_ , \new_[6972]_ ,
    \new_[6973]_ , \new_[6974]_ , \new_[6975]_ , \new_[6976]_ ,
    \new_[6977]_ , \new_[6978]_ , \new_[6979]_ , \new_[6980]_ ,
    \new_[6981]_ , \new_[6982]_ , \new_[6983]_ , \new_[6984]_ ,
    \new_[6985]_ , \new_[6986]_ , \new_[6987]_ , \new_[6988]_ ,
    \new_[6989]_ , \new_[6990]_ , \new_[6991]_ , \new_[6992]_ ,
    \new_[6993]_ , \new_[6994]_ , \new_[6995]_ , \new_[6996]_ ,
    \new_[6997]_ , \new_[6998]_ , \new_[6999]_ , \new_[7000]_ ,
    \new_[7001]_ , \new_[7002]_ , \new_[7003]_ , \new_[7004]_ ,
    \new_[7005]_ , \new_[7006]_ , \new_[7007]_ , \new_[7008]_ ,
    \new_[7009]_ , \new_[7010]_ , \new_[7011]_ , \new_[7012]_ ,
    \new_[7013]_ , \new_[7014]_ , \new_[7015]_ , \new_[7016]_ ,
    \new_[7017]_ , \new_[7018]_ , \new_[7019]_ , \new_[7020]_ ,
    \new_[7021]_ , \new_[7022]_ , \new_[7023]_ , \new_[7024]_ ,
    \new_[7025]_ , \new_[7026]_ , \new_[7027]_ , \new_[7028]_ ,
    \new_[7029]_ , \new_[7030]_ , \new_[7031]_ , \new_[7032]_ ,
    \new_[7033]_ , \new_[7034]_ , \new_[7035]_ , \new_[7036]_ ,
    \new_[7037]_ , \new_[7038]_ , \new_[7039]_ , \new_[7040]_ ,
    \new_[7041]_ , \new_[7042]_ , \new_[7043]_ , \new_[7044]_ ,
    \new_[7045]_ , \new_[7046]_ , \new_[7047]_ , \new_[7048]_ ,
    \new_[7049]_ , \new_[7050]_ , \new_[7051]_ , \new_[7052]_ ,
    \new_[7053]_ , \new_[7054]_ , \new_[7055]_ , \new_[7056]_ ,
    \new_[7057]_ , \new_[7058]_ , \new_[7059]_ , \new_[7060]_ ,
    \new_[7061]_ , \new_[7062]_ , \new_[7063]_ , \new_[7064]_ ,
    \new_[7065]_ , \new_[7066]_ , \new_[7067]_ , \new_[7068]_ ,
    \new_[7069]_ , \new_[7070]_ , \new_[7071]_ , \new_[7072]_ ,
    \new_[7073]_ , \new_[7074]_ , \new_[7075]_ , \new_[7076]_ ,
    \new_[7077]_ , \new_[7078]_ , \new_[7079]_ , \new_[7080]_ ,
    \new_[7081]_ , \new_[7082]_ , \new_[7083]_ , \new_[7084]_ ,
    \new_[7085]_ , \new_[7086]_ , \new_[7087]_ , \new_[7088]_ ,
    \new_[7089]_ , \new_[7090]_ , \new_[7091]_ , \new_[7092]_ ,
    \new_[7093]_ , \new_[7094]_ , \new_[7095]_ , \new_[7096]_ ,
    \new_[7097]_ , \new_[7098]_ , \new_[7099]_ , \new_[7100]_ ,
    \new_[7101]_ , \new_[7102]_ , \new_[7103]_ , \new_[7104]_ ,
    \new_[7105]_ , \new_[7106]_ , \new_[7107]_ , \new_[7108]_ ,
    \new_[7109]_ , \new_[7110]_ , \new_[7111]_ , \new_[7112]_ ,
    \new_[7113]_ , \new_[7114]_ , \new_[7115]_ , \new_[7116]_ ,
    \new_[7117]_ , \new_[7118]_ , \new_[7119]_ , \new_[7120]_ ,
    \new_[7121]_ , \new_[7122]_ , \new_[7123]_ , \new_[7124]_ ,
    \new_[7125]_ , \new_[7126]_ , \new_[7127]_ , \new_[7128]_ ,
    \new_[7129]_ , \new_[7130]_ , \new_[7131]_ , \new_[7132]_ ,
    \new_[7133]_ , \new_[7134]_ , \new_[7135]_ , \new_[7136]_ ,
    \new_[7137]_ , \new_[7138]_ , \new_[7139]_ , \new_[7140]_ ,
    \new_[7141]_ , \new_[7142]_ , \new_[7143]_ , \new_[7144]_ ,
    \new_[7145]_ , \new_[7146]_ , \new_[7147]_ , \new_[7148]_ ,
    \new_[7149]_ , \new_[7150]_ , \new_[7151]_ , \new_[7152]_ ,
    \new_[7153]_ , \new_[7154]_ , \new_[7155]_ , \new_[7156]_ ,
    \new_[7157]_ , \new_[7158]_ , \new_[7159]_ , \new_[7160]_ ,
    \new_[7161]_ , \new_[7162]_ , \new_[7163]_ , \new_[7164]_ ,
    \new_[7165]_ , \new_[7166]_ , \new_[7167]_ , \new_[7168]_ ,
    \new_[7169]_ , \new_[7170]_ , \new_[7171]_ , \new_[7172]_ ,
    \new_[7173]_ , \new_[7174]_ , \new_[7175]_ , \new_[7176]_ ,
    \new_[7177]_ , \new_[7178]_ , \new_[7179]_ , \new_[7180]_ ,
    \new_[7181]_ , \new_[7182]_ , \new_[7183]_ , \new_[7184]_ ,
    \new_[7185]_ , \new_[7186]_ , \new_[7187]_ , \new_[7188]_ ,
    \new_[7189]_ , \new_[7190]_ , \new_[7191]_ , \new_[7192]_ ,
    \new_[7193]_ , \new_[7194]_ , \new_[7195]_ , \new_[7196]_ ,
    \new_[7197]_ , \new_[7198]_ , \new_[7199]_ , \new_[7200]_ ,
    \new_[7201]_ , \new_[7202]_ , \new_[7203]_ , \new_[7204]_ ,
    \new_[7205]_ , \new_[7206]_ , \new_[7207]_ , \new_[7208]_ ,
    \new_[7209]_ , \new_[7210]_ , \new_[7211]_ , \new_[7212]_ ,
    \new_[7213]_ , \new_[7214]_ , \new_[7215]_ , \new_[7216]_ ,
    \new_[7217]_ , \new_[7218]_ , \new_[7219]_ , \new_[7220]_ ,
    \new_[7221]_ , \new_[7222]_ , \new_[7223]_ , \new_[7224]_ ,
    \new_[7225]_ , \new_[7226]_ , \new_[7227]_ , \new_[7228]_ ,
    \new_[7229]_ , \new_[7230]_ , \new_[7231]_ , \new_[7232]_ ,
    \new_[7233]_ , \new_[7234]_ , \new_[7235]_ , \new_[7236]_ ,
    \new_[7237]_ , \new_[7238]_ , \new_[7239]_ , \new_[7240]_ ,
    \new_[7241]_ , \new_[7242]_ , \new_[7243]_ , \new_[7244]_ ,
    \new_[7245]_ , \new_[7246]_ , \new_[7247]_ , \new_[7248]_ ,
    \new_[7249]_ , \new_[7250]_ , \new_[7251]_ , \new_[7252]_ ,
    \new_[7253]_ , \new_[7254]_ , \new_[7255]_ , \new_[7256]_ ,
    \new_[7257]_ , \new_[7258]_ , \new_[7259]_ , \new_[7260]_ ,
    \new_[7261]_ , \new_[7262]_ , \new_[7263]_ , \new_[7264]_ ,
    \new_[7265]_ , \new_[7266]_ , \new_[7267]_ , \new_[7268]_ ,
    \new_[7269]_ , \new_[7270]_ , \new_[7271]_ , \new_[7272]_ ,
    \new_[7273]_ , \new_[7274]_ , \new_[7275]_ , \new_[7276]_ ,
    \new_[7277]_ , \new_[7278]_ , \new_[7279]_ , \new_[7280]_ ,
    \new_[7281]_ , \new_[7282]_ , \new_[7283]_ , \new_[7284]_ ,
    \new_[7285]_ , \new_[7286]_ , \new_[7287]_ , \new_[7288]_ ,
    \new_[7289]_ , \new_[7290]_ , \new_[7291]_ , \new_[7292]_ ,
    \new_[7293]_ , \new_[7294]_ , \new_[7295]_ , \new_[7296]_ ,
    \new_[7297]_ , \new_[7298]_ , \new_[7299]_ , \new_[7300]_ ,
    \new_[7301]_ , \new_[7302]_ , \new_[7303]_ , \new_[7304]_ ,
    \new_[7305]_ , \new_[7306]_ , \new_[7307]_ , \new_[7308]_ ,
    \new_[7309]_ , \new_[7310]_ , \new_[7311]_ , \new_[7312]_ ,
    \new_[7313]_ , \new_[7314]_ , \new_[7315]_ , \new_[7316]_ ,
    \new_[7317]_ , \new_[7318]_ , \new_[7319]_ , \new_[7320]_ ,
    \new_[7321]_ , \new_[7322]_ , \new_[7323]_ , \new_[7324]_ ,
    \new_[7325]_ , \new_[7326]_ , \new_[7327]_ , \new_[7328]_ ,
    \new_[7329]_ , \new_[7330]_ , \new_[7331]_ , \new_[7332]_ ,
    \new_[7333]_ , \new_[7334]_ , \new_[7335]_ , \new_[7336]_ ,
    \new_[7337]_ , \new_[7338]_ , \new_[7339]_ , \new_[7340]_ ,
    \new_[7341]_ , \new_[7342]_ , \new_[7343]_ , \new_[7344]_ ,
    \new_[7345]_ , \new_[7346]_ , \new_[7347]_ , \new_[7348]_ ,
    \new_[7349]_ , \new_[7350]_ , \new_[7351]_ , \new_[7352]_ ,
    \new_[7353]_ , \new_[7354]_ , \new_[7355]_ , \new_[7356]_ ,
    \new_[7357]_ , \new_[7358]_ , \new_[7359]_ , \new_[7360]_ ,
    \new_[7361]_ , \new_[7362]_ , \new_[7363]_ , \new_[7364]_ ,
    \new_[7365]_ , \new_[7366]_ , \new_[7367]_ , \new_[7368]_ ,
    \new_[7369]_ , \new_[7370]_ , \new_[7371]_ , \new_[7372]_ ,
    \new_[7373]_ , \new_[7374]_ , \new_[7375]_ , \new_[7376]_ ,
    \new_[7377]_ , \new_[7378]_ , \new_[7379]_ , \new_[7380]_ ,
    \new_[7381]_ , \new_[7382]_ , \new_[7383]_ , \new_[7384]_ ,
    \new_[7385]_ , \new_[7386]_ , \new_[7387]_ , \new_[7388]_ ,
    \new_[7389]_ , \new_[7390]_ , \new_[7391]_ , \new_[7392]_ ,
    \new_[7393]_ , \new_[7394]_ , \new_[7395]_ , \new_[7396]_ ,
    \new_[7397]_ , \new_[7398]_ , \new_[7399]_ , \new_[7400]_ ,
    \new_[7401]_ , \new_[7402]_ , \new_[7403]_ , \new_[7404]_ ,
    \new_[7405]_ , \new_[7406]_ , \new_[7407]_ , \new_[7408]_ ,
    \new_[7409]_ , \new_[7410]_ , \new_[7411]_ , \new_[7412]_ ,
    \new_[7413]_ , \new_[7414]_ , \new_[7415]_ , \new_[7416]_ ,
    \new_[7417]_ , \new_[7418]_ , \new_[7420]_ , \new_[7421]_ ,
    \new_[7422]_ , \new_[7423]_ , \new_[7424]_ , \new_[7425]_ ,
    \new_[7427]_ , \new_[7428]_ , \new_[7429]_ , \new_[7430]_ ,
    \new_[7431]_ , \new_[7432]_ , \new_[7433]_ , \new_[7434]_ ,
    \new_[7437]_ , \new_[7438]_ , \new_[7439]_ , \new_[7441]_ ,
    \new_[7442]_ , \new_[7443]_ , \new_[7451]_ , \new_[7459]_ ,
    \new_[7461]_ , \new_[7462]_ , \new_[7463]_ , \new_[7465]_ ,
    \new_[7466]_ , \new_[7467]_ , \new_[7468]_ , \new_[7469]_ ,
    \new_[7470]_ , \new_[7471]_ , \new_[7472]_ , \new_[7473]_ ,
    \new_[7474]_ , \new_[7475]_ , \new_[7476]_ , \new_[7477]_ ,
    \new_[7478]_ , \new_[7479]_ , \new_[7480]_ , \new_[7481]_ ,
    \new_[7490]_ , \new_[7491]_ , \new_[7492]_ , \new_[7493]_ ,
    \new_[7494]_ , \new_[7495]_ , \new_[7496]_ , \new_[7497]_ ,
    \new_[7498]_ , \new_[7499]_ , \new_[7500]_ , \new_[7501]_ ,
    \new_[7502]_ , \new_[7503]_ , \new_[7504]_ , \new_[7505]_ ,
    \new_[7506]_ , \new_[7507]_ , \new_[7508]_ , \new_[7509]_ ,
    \new_[7510]_ , \new_[7511]_ , \new_[7512]_ , \new_[7513]_ ,
    \new_[7514]_ , \new_[7519]_ , \new_[7520]_ , \new_[7521]_ ,
    \new_[7522]_ , \new_[7523]_ , \new_[7524]_ , \new_[7525]_ ,
    \new_[7526]_ , \new_[7527]_ , \new_[7528]_ , \new_[7529]_ ,
    \new_[7530]_ , \new_[7531]_ , \new_[7532]_ , \new_[7533]_ ,
    \new_[7534]_ , \new_[7535]_ , \new_[7536]_ , \new_[7537]_ ,
    \new_[7538]_ , \new_[7539]_ , \new_[7540]_ , \new_[7541]_ ,
    \new_[7542]_ , \new_[7543]_ , \new_[7544]_ , \new_[7545]_ ,
    \new_[7546]_ , \new_[7547]_ , \new_[7548]_ , \new_[7549]_ ,
    \new_[7550]_ , \new_[7551]_ , \new_[7552]_ , \new_[7553]_ ,
    \new_[7554]_ , \new_[7555]_ , \new_[7556]_ , \new_[7557]_ ,
    \new_[7558]_ , \new_[7559]_ , \new_[7560]_ , \new_[7561]_ ,
    \new_[7562]_ , \new_[7563]_ , \new_[7564]_ , \new_[7565]_ ,
    \new_[7566]_ , \new_[7567]_ , \new_[7568]_ , \new_[7569]_ ,
    \new_[7570]_ , \new_[7571]_ , \new_[7572]_ , \new_[7573]_ ,
    \new_[7574]_ , \new_[7575]_ , \new_[7576]_ , \new_[7577]_ ,
    \new_[7578]_ , \new_[7579]_ , \new_[7580]_ , \new_[7581]_ ,
    \new_[7582]_ , \new_[7583]_ , \new_[7584]_ , \new_[7585]_ ,
    \new_[7586]_ , \new_[7587]_ , \new_[7588]_ , \new_[7589]_ ,
    \new_[7590]_ , \new_[7591]_ , \new_[7593]_ , \new_[7594]_ ,
    \new_[7595]_ , \new_[7596]_ , \new_[7597]_ , \new_[7598]_ ,
    \new_[7599]_ , \new_[7600]_ , \new_[7601]_ , \new_[7602]_ ,
    \new_[7603]_ , \new_[7604]_ , \new_[7605]_ , \new_[7606]_ ,
    \new_[7607]_ , \new_[7608]_ , \new_[7609]_ , \new_[7610]_ ,
    \new_[7611]_ , \new_[7612]_ , \new_[7613]_ , \new_[7614]_ ,
    \new_[7615]_ , \new_[7616]_ , \new_[7617]_ , \new_[7626]_ ,
    \new_[7628]_ , \new_[7636]_ , \new_[7637]_ , \new_[7638]_ ,
    \new_[7639]_ , \new_[7640]_ , \new_[7641]_ , \new_[7642]_ ,
    \new_[7643]_ , \new_[7644]_ , \new_[7645]_ , \new_[7646]_ ,
    \new_[7647]_ , \new_[7648]_ , \new_[7649]_ , \new_[7650]_ ,
    \new_[7651]_ , \new_[7652]_ , \new_[7653]_ , \new_[7654]_ ,
    \new_[7655]_ , \new_[7656]_ , \new_[7657]_ , \new_[7658]_ ,
    \new_[7659]_ , \new_[7660]_ , \new_[7661]_ , \new_[7662]_ ,
    \new_[7663]_ , \new_[7664]_ , \new_[7665]_ , \new_[7666]_ ,
    \new_[7667]_ , \new_[7668]_ , \new_[7669]_ , \new_[7670]_ ,
    \new_[7671]_ , \new_[7672]_ , \new_[7673]_ , \new_[7674]_ ,
    \new_[7675]_ , \new_[7676]_ , \new_[7677]_ , \new_[7678]_ ,
    \new_[7679]_ , \new_[7680]_ , \new_[7681]_ , \new_[7682]_ ,
    \new_[7683]_ , \new_[7684]_ , \new_[7685]_ , \new_[7686]_ ,
    \new_[7687]_ , \new_[7688]_ , \new_[7689]_ , \new_[7690]_ ,
    \new_[7691]_ , \new_[7692]_ , \new_[7693]_ , \new_[7694]_ ,
    \new_[7695]_ , \new_[7696]_ , \new_[7697]_ , \new_[7698]_ ,
    \new_[7699]_ , \new_[7700]_ , \new_[7701]_ , \new_[7702]_ ,
    \new_[7703]_ , \new_[7704]_ , \new_[7705]_ , \new_[7706]_ ,
    \new_[7707]_ , \new_[7708]_ , \new_[7709]_ , \new_[7710]_ ,
    \new_[7711]_ , \new_[7714]_ , \new_[7715]_ , \new_[7716]_ ,
    \new_[7717]_ , \new_[7718]_ , \new_[7719]_ , \new_[7720]_ ,
    \new_[7721]_ , \new_[7722]_ , \new_[7723]_ , \new_[7724]_ ,
    \new_[7725]_ , \new_[7726]_ , \new_[7727]_ , \new_[7728]_ ,
    \new_[7729]_ , \new_[7730]_ , \new_[7731]_ , \new_[7732]_ ,
    \new_[7733]_ , \new_[7734]_ , \new_[7735]_ , \new_[7736]_ ,
    \new_[7737]_ , \new_[7738]_ , \new_[7739]_ , \new_[7740]_ ,
    \new_[7741]_ , \new_[7742]_ , \new_[7743]_ , \new_[7744]_ ,
    \new_[7745]_ , \new_[7746]_ , \new_[7747]_ , \new_[7748]_ ,
    \new_[7749]_ , \new_[7751]_ , \new_[7752]_ , \new_[7753]_ ,
    \new_[7754]_ , \new_[7755]_ , \new_[7756]_ , \new_[7757]_ ,
    \new_[7758]_ , \new_[7759]_ , \new_[7760]_ , \new_[7761]_ ,
    \new_[7762]_ , \new_[7763]_ , \new_[7764]_ , \new_[7765]_ ,
    \new_[7766]_ , \new_[7767]_ , \new_[7768]_ , \new_[7769]_ ,
    \new_[7770]_ , \new_[7771]_ , \new_[7772]_ , \new_[7773]_ ,
    \new_[7774]_ , \new_[7775]_ , \new_[7776]_ , \new_[7777]_ ,
    \new_[7779]_ , \new_[7780]_ , \new_[7781]_ , \new_[7782]_ ,
    \new_[7783]_ , \new_[7784]_ , \new_[7785]_ , \new_[7786]_ ,
    \new_[7787]_ , \new_[7788]_ , \new_[7789]_ , \new_[7790]_ ,
    \new_[7791]_ , \new_[7792]_ , \new_[7793]_ , \new_[7794]_ ,
    \new_[7795]_ , \new_[7796]_ , \new_[7797]_ , \new_[7798]_ ,
    \new_[7799]_ , \new_[7800]_ , \new_[7801]_ , \new_[7802]_ ,
    \new_[7803]_ , \new_[7804]_ , \new_[7805]_ , \new_[7806]_ ,
    \new_[7807]_ , \new_[7808]_ , \new_[7809]_ , \new_[7810]_ ,
    \new_[7811]_ , \new_[7812]_ , \new_[7816]_ , \new_[7817]_ ,
    \new_[7818]_ , \new_[7819]_ , \new_[7820]_ , \new_[7821]_ ,
    \new_[7822]_ , \new_[7823]_ , \new_[7824]_ , \new_[7825]_ ,
    \new_[7827]_ , \new_[7828]_ , \new_[7829]_ , \new_[7832]_ ,
    \new_[7833]_ , \new_[7834]_ , \new_[7835]_ , \new_[7836]_ ,
    \new_[7837]_ , \new_[7838]_ , \new_[7839]_ , \new_[7840]_ ,
    \new_[7841]_ , \new_[7842]_ , \new_[7843]_ , \new_[7844]_ ,
    \new_[7845]_ , \new_[7846]_ , \new_[7847]_ , \new_[7848]_ ,
    \new_[7849]_ , \new_[7850]_ , \new_[7851]_ , \new_[7852]_ ,
    \new_[7853]_ , \new_[7854]_ , \new_[7855]_ , \new_[7856]_ ,
    \new_[7857]_ , \new_[7858]_ , \new_[7859]_ , \new_[7860]_ ,
    \new_[7861]_ , \new_[7862]_ , \new_[7863]_ , \new_[7864]_ ,
    \new_[7865]_ , \new_[7866]_ , \new_[7867]_ , \new_[7868]_ ,
    \new_[7869]_ , \new_[7870]_ , \new_[7871]_ , \new_[7872]_ ,
    \new_[7873]_ , \new_[7874]_ , \new_[7875]_ , \new_[7876]_ ,
    \new_[7877]_ , \new_[7878]_ , \new_[7879]_ , \new_[7881]_ ,
    \new_[7882]_ , \new_[7883]_ , \new_[7884]_ , \new_[7885]_ ,
    \new_[7886]_ , \new_[7887]_ , \new_[7888]_ , \new_[7889]_ ,
    \new_[7890]_ , \new_[7891]_ , \new_[7892]_ , \new_[7893]_ ,
    \new_[7894]_ , \new_[7895]_ , \new_[7896]_ , \new_[7897]_ ,
    \new_[7898]_ , \new_[7899]_ , \new_[7900]_ , \new_[7901]_ ,
    \new_[7902]_ , \new_[7903]_ , \new_[7904]_ , \new_[7905]_ ,
    \new_[7906]_ , \new_[7907]_ , \new_[7908]_ , \new_[7909]_ ,
    \new_[7910]_ , \new_[7911]_ , \new_[7912]_ , \new_[7913]_ ,
    \new_[7914]_ , \new_[7915]_ , \new_[7916]_ , \new_[7917]_ ,
    \new_[7918]_ , \new_[7919]_ , \new_[7920]_ , \new_[7921]_ ,
    \new_[7922]_ , \new_[7923]_ , \new_[7924]_ , \new_[7925]_ ,
    \new_[7926]_ , \new_[7927]_ , \new_[7928]_ , \new_[7929]_ ,
    \new_[7930]_ , \new_[7931]_ , \new_[7932]_ , \new_[7933]_ ,
    \new_[7934]_ , \new_[7935]_ , \new_[7936]_ , \new_[7937]_ ,
    \new_[7938]_ , \new_[7939]_ , \new_[7940]_ , \new_[7941]_ ,
    \new_[7942]_ , \new_[7943]_ , \new_[7945]_ , \new_[7946]_ ,
    \new_[7947]_ , \new_[7948]_ , \new_[7956]_ , \new_[7957]_ ,
    \new_[7960]_ , \new_[7961]_ , \new_[7962]_ , \new_[7963]_ ,
    \new_[7964]_ , \new_[7965]_ , \new_[7966]_ , \new_[7967]_ ,
    \new_[7968]_ , \new_[7969]_ , \new_[7970]_ , \new_[7971]_ ,
    \new_[7972]_ , \new_[7973]_ , \new_[7974]_ , \new_[7975]_ ,
    \new_[7976]_ , \new_[7977]_ , \new_[7978]_ , \new_[7979]_ ,
    \new_[7981]_ , \new_[7982]_ , \new_[7983]_ , \new_[7984]_ ,
    \new_[7985]_ , \new_[7986]_ , \new_[7987]_ , \new_[7988]_ ,
    \new_[7989]_ , \new_[7990]_ , \new_[7991]_ , \new_[7992]_ ,
    \new_[7993]_ , \new_[7994]_ , \new_[7995]_ , \new_[7996]_ ,
    \new_[7997]_ , \new_[7998]_ , \new_[7999]_ , \new_[8000]_ ,
    \new_[8001]_ , \new_[8002]_ , \new_[8003]_ , \new_[8004]_ ,
    \new_[8005]_ , \new_[8006]_ , \new_[8007]_ , \new_[8008]_ ,
    \new_[8009]_ , \new_[8010]_ , \new_[8011]_ , \new_[8012]_ ,
    \new_[8013]_ , \new_[8014]_ , \new_[8015]_ , \new_[8016]_ ,
    \new_[8017]_ , \new_[8018]_ , \new_[8019]_ , \new_[8020]_ ,
    \new_[8021]_ , \new_[8022]_ , \new_[8023]_ , \new_[8024]_ ,
    \new_[8025]_ , \new_[8026]_ , \new_[8027]_ , \new_[8028]_ ,
    \new_[8029]_ , \new_[8030]_ , \new_[8031]_ , \new_[8032]_ ,
    \new_[8033]_ , \new_[8034]_ , \new_[8035]_ , \new_[8036]_ ,
    \new_[8037]_ , \new_[8038]_ , \new_[8039]_ , \new_[8040]_ ,
    \new_[8041]_ , \new_[8042]_ , \new_[8043]_ , \new_[8044]_ ,
    \new_[8045]_ , \new_[8046]_ , \new_[8047]_ , \new_[8048]_ ,
    \new_[8049]_ , \new_[8050]_ , \new_[8051]_ , \new_[8052]_ ,
    \new_[8053]_ , \new_[8054]_ , \new_[8055]_ , \new_[8056]_ ,
    \new_[8057]_ , \new_[8058]_ , \new_[8059]_ , \new_[8060]_ ,
    \new_[8061]_ , \new_[8062]_ , \new_[8063]_ , \new_[8064]_ ,
    \new_[8065]_ , \new_[8066]_ , \new_[8067]_ , \new_[8068]_ ,
    \new_[8069]_ , \new_[8070]_ , \new_[8071]_ , \new_[8072]_ ,
    \new_[8073]_ , \new_[8074]_ , \new_[8075]_ , \new_[8076]_ ,
    \new_[8077]_ , \new_[8078]_ , \new_[8079]_ , \new_[8080]_ ,
    \new_[8081]_ , \new_[8082]_ , \new_[8083]_ , \new_[8084]_ ,
    \new_[8085]_ , \new_[8086]_ , \new_[8087]_ , \new_[8088]_ ,
    \new_[8089]_ , \new_[8090]_ , \new_[8091]_ , \new_[8094]_ ,
    \new_[8099]_ , \new_[8100]_ , \new_[8104]_ , \new_[8106]_ ,
    \new_[8112]_ , \new_[8113]_ , \new_[8114]_ , \new_[8115]_ ,
    \new_[8116]_ , \new_[8117]_ , \new_[8118]_ , \new_[8119]_ ,
    \new_[8120]_ , \new_[8134]_ , \new_[8135]_ , \new_[8136]_ ,
    \new_[8138]_ , \new_[8139]_ , \new_[8141]_ , \new_[8142]_ ,
    \new_[8143]_ , \new_[8144]_ , \new_[8145]_ , \new_[8146]_ ,
    \new_[8147]_ , \new_[8148]_ , \new_[8149]_ , \new_[8150]_ ,
    \new_[8151]_ , \new_[8152]_ , \new_[8153]_ , \new_[8154]_ ,
    \new_[8155]_ , \new_[8156]_ , \new_[8157]_ , \new_[8158]_ ,
    \new_[8159]_ , \new_[8160]_ , \new_[8161]_ , \new_[8162]_ ,
    \new_[8163]_ , \new_[8164]_ , \new_[8165]_ , \new_[8166]_ ,
    \new_[8167]_ , \new_[8168]_ , \new_[8169]_ , \new_[8170]_ ,
    \new_[8171]_ , \new_[8172]_ , \new_[8173]_ , \new_[8174]_ ,
    \new_[8178]_ , \new_[8179]_ , \new_[8180]_ , \new_[8181]_ ,
    \new_[8182]_ , \new_[8183]_ , \new_[8184]_ , \new_[8185]_ ,
    \new_[8186]_ , \new_[8187]_ , \new_[8188]_ , \new_[8189]_ ,
    \new_[8190]_ , \new_[8191]_ , \new_[8192]_ , \new_[8193]_ ,
    \new_[8194]_ , \new_[8195]_ , \new_[8196]_ , \new_[8197]_ ,
    \new_[8198]_ , \new_[8199]_ , \new_[8200]_ , \new_[8201]_ ,
    \new_[8202]_ , \new_[8203]_ , \new_[8204]_ , \new_[8205]_ ,
    \new_[8206]_ , \new_[8207]_ , \new_[8208]_ , \new_[8209]_ ,
    \new_[8210]_ , \new_[8211]_ , \new_[8212]_ , \new_[8213]_ ,
    \new_[8214]_ , \new_[8215]_ , \new_[8216]_ , \new_[8217]_ ,
    \new_[8218]_ , \new_[8219]_ , \new_[8220]_ , \new_[8221]_ ,
    \new_[8222]_ , \new_[8223]_ , \new_[8224]_ , \new_[8225]_ ,
    \new_[8226]_ , \new_[8227]_ , \new_[8228]_ , \new_[8229]_ ,
    \new_[8230]_ , \new_[8231]_ , \new_[8232]_ , \new_[8233]_ ,
    \new_[8234]_ , \new_[8235]_ , \new_[8236]_ , \new_[8237]_ ,
    \new_[8238]_ , \new_[8239]_ , \new_[8240]_ , \new_[8241]_ ,
    \new_[8242]_ , \new_[8243]_ , \new_[8244]_ , \new_[8245]_ ,
    \new_[8246]_ , \new_[8247]_ , \new_[8248]_ , \new_[8249]_ ,
    \new_[8250]_ , \new_[8251]_ , \new_[8252]_ , \new_[8253]_ ,
    \new_[8254]_ , \new_[8255]_ , \new_[8256]_ , \new_[8257]_ ,
    \new_[8258]_ , \new_[8259]_ , \new_[8260]_ , \new_[8261]_ ,
    \new_[8262]_ , \new_[8263]_ , \new_[8264]_ , \new_[8265]_ ,
    \new_[8266]_ , \new_[8267]_ , \new_[8268]_ , \new_[8269]_ ,
    \new_[8270]_ , \new_[8271]_ , \new_[8272]_ , \new_[8273]_ ,
    \new_[8274]_ , \new_[8275]_ , \new_[8276]_ , \new_[8277]_ ,
    \new_[8278]_ , \new_[8279]_ , \new_[8280]_ , \new_[8281]_ ,
    \new_[8282]_ , \new_[8283]_ , \new_[8284]_ , \new_[8285]_ ,
    \new_[8286]_ , \new_[8287]_ , \new_[8288]_ , \new_[8289]_ ,
    \new_[8290]_ , \new_[8291]_ , \new_[8292]_ , \new_[8293]_ ,
    \new_[8294]_ , \new_[8295]_ , \new_[8296]_ , \new_[8297]_ ,
    \new_[8298]_ , \new_[8299]_ , \new_[8300]_ , \new_[8301]_ ,
    \new_[8302]_ , \new_[8303]_ , \new_[8304]_ , \new_[8305]_ ,
    \new_[8306]_ , \new_[8307]_ , \new_[8308]_ , \new_[8309]_ ,
    \new_[8310]_ , \new_[8311]_ , \new_[8312]_ , \new_[8313]_ ,
    \new_[8314]_ , \new_[8315]_ , \new_[8316]_ , \new_[8317]_ ,
    \new_[8318]_ , \new_[8319]_ , \new_[8320]_ , \new_[8321]_ ,
    \new_[8322]_ , \new_[8323]_ , \new_[8324]_ , \new_[8325]_ ,
    \new_[8326]_ , \new_[8327]_ , \new_[8328]_ , \new_[8329]_ ,
    \new_[8330]_ , \new_[8331]_ , \new_[8332]_ , \new_[8333]_ ,
    \new_[8334]_ , \new_[8335]_ , \new_[8336]_ , \new_[8337]_ ,
    \new_[8338]_ , \new_[8339]_ , \new_[8340]_ , \new_[8341]_ ,
    \new_[8342]_ , \new_[8343]_ , \new_[8344]_ , \new_[8345]_ ,
    \new_[8346]_ , \new_[8347]_ , \new_[8348]_ , \new_[8349]_ ,
    \new_[8350]_ , \new_[8351]_ , \new_[8352]_ , \new_[8353]_ ,
    \new_[8354]_ , \new_[8355]_ , \new_[8356]_ , \new_[8357]_ ,
    \new_[8358]_ , \new_[8359]_ , \new_[8360]_ , \new_[8361]_ ,
    \new_[8362]_ , \new_[8363]_ , \new_[8364]_ , \new_[8365]_ ,
    \new_[8366]_ , \new_[8367]_ , \new_[8368]_ , \new_[8369]_ ,
    \new_[8370]_ , \new_[8371]_ , \new_[8372]_ , \new_[8373]_ ,
    \new_[8374]_ , \new_[8375]_ , \new_[8376]_ , \new_[8377]_ ,
    \new_[8378]_ , \new_[8379]_ , \new_[8380]_ , \new_[8381]_ ,
    \new_[8382]_ , \new_[8383]_ , \new_[8384]_ , \new_[8385]_ ,
    \new_[8386]_ , \new_[8387]_ , \new_[8388]_ , \new_[8389]_ ,
    \new_[8390]_ , \new_[8391]_ , \new_[8392]_ , \new_[8393]_ ,
    \new_[8394]_ , \new_[8395]_ , \new_[8396]_ , \new_[8397]_ ,
    \new_[8398]_ , \new_[8399]_ , \new_[8400]_ , \new_[8401]_ ,
    \new_[8402]_ , \new_[8403]_ , \new_[8404]_ , \new_[8405]_ ,
    \new_[8406]_ , \new_[8407]_ , \new_[8408]_ , \new_[8409]_ ,
    \new_[8410]_ , \new_[8411]_ , \new_[8412]_ , \new_[8413]_ ,
    \new_[8414]_ , \new_[8415]_ , \new_[8416]_ , \new_[8417]_ ,
    \new_[8418]_ , \new_[8419]_ , \new_[8420]_ , \new_[8421]_ ,
    \new_[8422]_ , \new_[8423]_ , \new_[8424]_ , \new_[8425]_ ,
    \new_[8426]_ , \new_[8427]_ , \new_[8428]_ , \new_[8429]_ ,
    \new_[8430]_ , \new_[8431]_ , \new_[8432]_ , \new_[8433]_ ,
    \new_[8434]_ , \new_[8435]_ , \new_[8436]_ , \new_[8437]_ ,
    \new_[8438]_ , \new_[8439]_ , \new_[8440]_ , \new_[8441]_ ,
    \new_[8442]_ , \new_[8443]_ , \new_[8444]_ , \new_[8445]_ ,
    \new_[8446]_ , \new_[8447]_ , \new_[8448]_ , \new_[8449]_ ,
    \new_[8450]_ , \new_[8451]_ , \new_[8452]_ , \new_[8453]_ ,
    \new_[8454]_ , \new_[8455]_ , \new_[8456]_ , \new_[8457]_ ,
    \new_[8458]_ , \new_[8459]_ , \new_[8460]_ , \new_[8461]_ ,
    \new_[8462]_ , \new_[8463]_ , \new_[8464]_ , \new_[8465]_ ,
    \new_[8466]_ , \new_[8467]_ , \new_[8468]_ , \new_[8469]_ ,
    \new_[8470]_ , \new_[8477]_ , \new_[8478]_ , \new_[8479]_ ,
    \new_[8483]_ , \new_[8484]_ , \new_[8485]_ , \new_[8487]_ ,
    \new_[8488]_ , \new_[8491]_ , \new_[8494]_ , \new_[8495]_ ,
    \new_[8496]_ , \new_[8497]_ , \new_[8498]_ , \new_[8499]_ ,
    \new_[8501]_ , \new_[8502]_ , \new_[8503]_ , \new_[8504]_ ,
    \new_[8505]_ , \new_[8506]_ , \new_[8507]_ , \new_[8508]_ ,
    \new_[8509]_ , \new_[8511]_ , \new_[8512]_ , \new_[8513]_ ,
    \new_[8514]_ , \new_[8515]_ , \new_[8516]_ , \new_[8517]_ ,
    \new_[8518]_ , \new_[8519]_ , \new_[8520]_ , \new_[8521]_ ,
    \new_[8522]_ , \new_[8523]_ , \new_[8524]_ , \new_[8525]_ ,
    \new_[8526]_ , \new_[8528]_ , \new_[8529]_ , \new_[8530]_ ,
    \new_[8531]_ , \new_[8532]_ , \new_[8533]_ , \new_[8534]_ ,
    \new_[8535]_ , \new_[8536]_ , \new_[8537]_ , \new_[8538]_ ,
    \new_[8539]_ , \new_[8540]_ , \new_[8541]_ , \new_[8542]_ ,
    \new_[8543]_ , \new_[8544]_ , \new_[8545]_ , \new_[8546]_ ,
    \new_[8547]_ , \new_[8548]_ , \new_[8549]_ , \new_[8550]_ ,
    \new_[8551]_ , \new_[8552]_ , \new_[8553]_ , \new_[8554]_ ,
    \new_[8555]_ , \new_[8556]_ , \new_[8557]_ , \new_[8558]_ ,
    \new_[8559]_ , \new_[8560]_ , \new_[8561]_ , \new_[8562]_ ,
    \new_[8563]_ , \new_[8564]_ , \new_[8565]_ , \new_[8566]_ ,
    \new_[8567]_ , \new_[8568]_ , \new_[8569]_ , \new_[8570]_ ,
    \new_[8571]_ , \new_[8572]_ , \new_[8573]_ , \new_[8574]_ ,
    \new_[8575]_ , \new_[8576]_ , \new_[8577]_ , \new_[8578]_ ,
    \new_[8579]_ , \new_[8580]_ , \new_[8581]_ , \new_[8582]_ ,
    \new_[8583]_ , \new_[8584]_ , \new_[8585]_ , \new_[8586]_ ,
    \new_[8587]_ , \new_[8588]_ , \new_[8589]_ , \new_[8590]_ ,
    \new_[8591]_ , \new_[8592]_ , \new_[8593]_ , \new_[8594]_ ,
    \new_[8596]_ , \new_[8597]_ , \new_[8598]_ , \new_[8599]_ ,
    \new_[8600]_ , \new_[8601]_ , \new_[8602]_ , \new_[8603]_ ,
    \new_[8604]_ , \new_[8605]_ , \new_[8606]_ , \new_[8607]_ ,
    \new_[8608]_ , \new_[8609]_ , \new_[8610]_ , \new_[8611]_ ,
    \new_[8612]_ , \new_[8613]_ , \new_[8614]_ , \new_[8615]_ ,
    \new_[8616]_ , \new_[8617]_ , \new_[8618]_ , \new_[8619]_ ,
    \new_[8620]_ , \new_[8621]_ , \new_[8622]_ , \new_[8623]_ ,
    \new_[8624]_ , \new_[8625]_ , \new_[8626]_ , \new_[8627]_ ,
    \new_[8628]_ , \new_[8629]_ , \new_[8630]_ , \new_[8634]_ ,
    \new_[8635]_ , \new_[8636]_ , \new_[8637]_ , \new_[8638]_ ,
    \new_[8639]_ , \new_[8640]_ , \new_[8641]_ , \new_[8642]_ ,
    \new_[8643]_ , \new_[8644]_ , \new_[8645]_ , \new_[8646]_ ,
    \new_[8647]_ , \new_[8648]_ , \new_[8649]_ , \new_[8650]_ ,
    \new_[8651]_ , \new_[8652]_ , \new_[8653]_ , \new_[8654]_ ,
    \new_[8655]_ , \new_[8656]_ , \new_[8657]_ , \new_[8658]_ ,
    \new_[8659]_ , \new_[8660]_ , \new_[8661]_ , \new_[8662]_ ,
    \new_[8663]_ , \new_[8664]_ , \new_[8665]_ , \new_[8666]_ ,
    \new_[8667]_ , \new_[8668]_ , \new_[8669]_ , \new_[8670]_ ,
    \new_[8671]_ , \new_[8672]_ , \new_[8673]_ , \new_[8674]_ ,
    \new_[8675]_ , \new_[8676]_ , \new_[8677]_ , \new_[8678]_ ,
    \new_[8679]_ , \new_[8680]_ , \new_[8681]_ , \new_[8682]_ ,
    \new_[8683]_ , \new_[8684]_ , \new_[8685]_ , \new_[8686]_ ,
    \new_[8687]_ , \new_[8688]_ , \new_[8689]_ , \new_[8690]_ ,
    \new_[8692]_ , \new_[8693]_ , \new_[8694]_ , \new_[8695]_ ,
    \new_[8696]_ , \new_[8697]_ , \new_[8698]_ , \new_[8699]_ ,
    \new_[8700]_ , \new_[8701]_ , \new_[8702]_ , \new_[8703]_ ,
    \new_[8704]_ , \new_[8705]_ , \new_[8706]_ , \new_[8707]_ ,
    \new_[8708]_ , \new_[8709]_ , \new_[8710]_ , \new_[8711]_ ,
    \new_[8712]_ , \new_[8713]_ , \new_[8714]_ , \new_[8715]_ ,
    \new_[8716]_ , \new_[8717]_ , \new_[8718]_ , \new_[8719]_ ,
    \new_[8720]_ , \new_[8721]_ , \new_[8722]_ , \new_[8723]_ ,
    \new_[8724]_ , \new_[8725]_ , \new_[8726]_ , \new_[8727]_ ,
    \new_[8728]_ , \new_[8729]_ , \new_[8730]_ , \new_[8731]_ ,
    \new_[8732]_ , \new_[8733]_ , \new_[8734]_ , \new_[8735]_ ,
    \new_[8736]_ , \new_[8737]_ , \new_[8738]_ , \new_[8739]_ ,
    \new_[8740]_ , \new_[8741]_ , \new_[8742]_ , \new_[8743]_ ,
    \new_[8744]_ , \new_[8745]_ , \new_[8746]_ , \new_[8747]_ ,
    \new_[8748]_ , \new_[8749]_ , \new_[8750]_ , \new_[8751]_ ,
    \new_[8752]_ , \new_[8753]_ , \new_[8754]_ , \new_[8755]_ ,
    \new_[8756]_ , \new_[8757]_ , \new_[8758]_ , \new_[8759]_ ,
    \new_[8760]_ , \new_[8761]_ , \new_[8762]_ , \new_[8763]_ ,
    \new_[8764]_ , \new_[8765]_ , \new_[8766]_ , \new_[8767]_ ,
    \new_[8768]_ , \new_[8769]_ , \new_[8770]_ , \new_[8771]_ ,
    \new_[8772]_ , \new_[8773]_ , \new_[8774]_ , \new_[8775]_ ,
    \new_[8776]_ , \new_[8777]_ , \new_[8778]_ , \new_[8779]_ ,
    \new_[8780]_ , \new_[8781]_ , \new_[8782]_ , \new_[8783]_ ,
    \new_[8784]_ , \new_[8786]_ , \new_[8787]_ , \new_[8788]_ ,
    \new_[8789]_ , \new_[8790]_ , \new_[8791]_ , \new_[8792]_ ,
    \new_[8795]_ , \new_[8796]_ , \new_[8801]_ , \new_[8802]_ ,
    \new_[8803]_ , \new_[8804]_ , \new_[8805]_ , \new_[8806]_ ,
    \new_[8810]_ , \new_[8811]_ , \new_[8812]_ , \new_[8813]_ ,
    \new_[8814]_ , \new_[8815]_ , \new_[8816]_ , \new_[8817]_ ,
    \new_[8818]_ , \new_[8819]_ , \new_[8820]_ , \new_[8821]_ ,
    \new_[8822]_ , \new_[8823]_ , \new_[8824]_ , \new_[8825]_ ,
    \new_[8826]_ , \new_[8827]_ , \new_[8829]_ , \new_[8830]_ ,
    \new_[8831]_ , \new_[8832]_ , \new_[8833]_ , \new_[8835]_ ,
    \new_[8836]_ , \new_[8837]_ , \new_[8838]_ , \new_[8839]_ ,
    \new_[8840]_ , \new_[8841]_ , \new_[8842]_ , \new_[8843]_ ,
    \new_[8844]_ , \new_[8845]_ , \new_[8846]_ , \new_[8847]_ ,
    \new_[8848]_ , \new_[8849]_ , \new_[8850]_ , \new_[8851]_ ,
    \new_[8852]_ , \new_[8853]_ , \new_[8854]_ , \new_[8855]_ ,
    \new_[8856]_ , \new_[8857]_ , \new_[8858]_ , \new_[8859]_ ,
    \new_[8860]_ , \new_[8861]_ , \new_[8862]_ , \new_[8863]_ ,
    \new_[8864]_ , \new_[8865]_ , \new_[8866]_ , \new_[8867]_ ,
    \new_[8868]_ , \new_[8869]_ , \new_[8870]_ , \new_[8871]_ ,
    \new_[8872]_ , \new_[8873]_ , \new_[8874]_ , \new_[8875]_ ,
    \new_[8876]_ , \new_[8877]_ , \new_[8878]_ , \new_[8879]_ ,
    \new_[8880]_ , \new_[8881]_ , \new_[8882]_ , \new_[8883]_ ,
    \new_[8884]_ , \new_[8885]_ , \new_[8886]_ , \new_[8887]_ ,
    \new_[8888]_ , \new_[8889]_ , \new_[8890]_ , \new_[8891]_ ,
    \new_[8892]_ , \new_[8893]_ , \new_[8894]_ , \new_[8895]_ ,
    \new_[8896]_ , \new_[8897]_ , \new_[8898]_ , \new_[8899]_ ,
    \new_[8900]_ , \new_[8901]_ , \new_[8902]_ , \new_[8903]_ ,
    \new_[8904]_ , \new_[8905]_ , \new_[8906]_ , \new_[8907]_ ,
    \new_[8908]_ , \new_[8909]_ , \new_[8910]_ , \new_[8911]_ ,
    \new_[8912]_ , \new_[8913]_ , \new_[8914]_ , \new_[8915]_ ,
    \new_[8916]_ , \new_[8917]_ , \new_[8918]_ , \new_[8919]_ ,
    \new_[8920]_ , \new_[8921]_ , \new_[8922]_ , \new_[8923]_ ,
    \new_[8924]_ , \new_[8925]_ , \new_[8926]_ , \new_[8927]_ ,
    \new_[8928]_ , \new_[8929]_ , \new_[8930]_ , \new_[8931]_ ,
    \new_[8932]_ , \new_[8933]_ , \new_[8934]_ , \new_[8935]_ ,
    \new_[8936]_ , \new_[8937]_ , \new_[8938]_ , \new_[8939]_ ,
    \new_[8940]_ , \new_[8941]_ , \new_[8942]_ , \new_[8943]_ ,
    \new_[8944]_ , \new_[8945]_ , \new_[8946]_ , \new_[8947]_ ,
    \new_[8948]_ , \new_[8949]_ , \new_[8950]_ , \new_[8951]_ ,
    \new_[8952]_ , \new_[8953]_ , \new_[8954]_ , \new_[8955]_ ,
    \new_[8956]_ , \new_[8957]_ , \new_[8958]_ , \new_[8959]_ ,
    \new_[8960]_ , \new_[8961]_ , \new_[8962]_ , \new_[8963]_ ,
    \new_[8964]_ , \new_[8965]_ , \new_[8966]_ , \new_[8967]_ ,
    \new_[8968]_ , \new_[8969]_ , \new_[8970]_ , \new_[8971]_ ,
    \new_[8972]_ , \new_[8973]_ , \new_[8974]_ , \new_[8975]_ ,
    \new_[8976]_ , \new_[8977]_ , \new_[8978]_ , \new_[8979]_ ,
    \new_[8980]_ , \new_[8981]_ , \new_[8982]_ , \new_[8983]_ ,
    \new_[8984]_ , \new_[8985]_ , \new_[8986]_ , \new_[8987]_ ,
    \new_[8988]_ , \new_[8989]_ , \new_[8990]_ , \new_[8991]_ ,
    \new_[8992]_ , \new_[8993]_ , \new_[8995]_ , \new_[8996]_ ,
    \new_[8997]_ , \new_[8998]_ , \new_[8999]_ , \new_[9000]_ ,
    \new_[9001]_ , \new_[9002]_ , \new_[9003]_ , \new_[9006]_ ,
    \new_[9007]_ , \new_[9008]_ , \new_[9009]_ , \new_[9010]_ ,
    \new_[9011]_ , \new_[9012]_ , \new_[9013]_ , \new_[9014]_ ,
    \new_[9015]_ , \new_[9016]_ , \new_[9017]_ , \new_[9018]_ ,
    \new_[9019]_ , \new_[9020]_ , \new_[9021]_ , \new_[9022]_ ,
    \new_[9023]_ , \new_[9024]_ , \new_[9025]_ , \new_[9026]_ ,
    \new_[9028]_ , \new_[9029]_ , \new_[9030]_ , \new_[9031]_ ,
    \new_[9032]_ , \new_[9033]_ , \new_[9034]_ , \new_[9035]_ ,
    \new_[9036]_ , \new_[9037]_ , \new_[9038]_ , \new_[9039]_ ,
    \new_[9040]_ , \new_[9041]_ , \new_[9042]_ , \new_[9043]_ ,
    \new_[9044]_ , \new_[9045]_ , \new_[9046]_ , \new_[9047]_ ,
    \new_[9048]_ , \new_[9049]_ , \new_[9050]_ , \new_[9051]_ ,
    \new_[9052]_ , \new_[9053]_ , \new_[9054]_ , \new_[9055]_ ,
    \new_[9056]_ , \new_[9057]_ , \new_[9058]_ , \new_[9059]_ ,
    \new_[9060]_ , \new_[9061]_ , \new_[9062]_ , \new_[9063]_ ,
    \new_[9064]_ , \new_[9065]_ , \new_[9066]_ , \new_[9067]_ ,
    \new_[9068]_ , \new_[9069]_ , \new_[9070]_ , \new_[9071]_ ,
    \new_[9072]_ , \new_[9073]_ , \new_[9074]_ , \new_[9075]_ ,
    \new_[9076]_ , \new_[9077]_ , \new_[9078]_ , \new_[9079]_ ,
    \new_[9080]_ , \new_[9081]_ , \new_[9082]_ , \new_[9085]_ ,
    \new_[9086]_ , \new_[9087]_ , \new_[9088]_ , \new_[9089]_ ,
    \new_[9090]_ , \new_[9091]_ , \new_[9092]_ , \new_[9093]_ ,
    \new_[9094]_ , \new_[9095]_ , \new_[9096]_ , \new_[9097]_ ,
    \new_[9098]_ , \new_[9099]_ , \new_[9100]_ , \new_[9101]_ ,
    \new_[9102]_ , \new_[9103]_ , \new_[9113]_ , \new_[9114]_ ,
    \new_[9115]_ , \new_[9116]_ , \new_[9117]_ , \new_[9118]_ ,
    \new_[9119]_ , \new_[9120]_ , \new_[9121]_ , \new_[9122]_ ,
    \new_[9123]_ , \new_[9124]_ , \new_[9125]_ , \new_[9128]_ ,
    \new_[9129]_ , \new_[9130]_ , \new_[9131]_ , \new_[9132]_ ,
    \new_[9133]_ , \new_[9134]_ , \new_[9135]_ , \new_[9136]_ ,
    \new_[9137]_ , \new_[9138]_ , \new_[9139]_ , \new_[9140]_ ,
    \new_[9141]_ , \new_[9142]_ , \new_[9143]_ , \new_[9144]_ ,
    \new_[9145]_ , \new_[9146]_ , \new_[9147]_ , \new_[9148]_ ,
    \new_[9149]_ , \new_[9150]_ , \new_[9151]_ , \new_[9152]_ ,
    \new_[9153]_ , \new_[9154]_ , \new_[9155]_ , \new_[9156]_ ,
    \new_[9157]_ , \new_[9158]_ , \new_[9159]_ , \new_[9160]_ ,
    \new_[9161]_ , \new_[9162]_ , \new_[9163]_ , \new_[9164]_ ,
    \new_[9165]_ , \new_[9166]_ , \new_[9167]_ , \new_[9168]_ ,
    \new_[9169]_ , \new_[9170]_ , \new_[9171]_ , \new_[9172]_ ,
    \new_[9173]_ , \new_[9174]_ , \new_[9175]_ , \new_[9176]_ ,
    \new_[9177]_ , \new_[9178]_ , \new_[9179]_ , \new_[9180]_ ,
    \new_[9181]_ , \new_[9182]_ , \new_[9183]_ , \new_[9184]_ ,
    \new_[9185]_ , \new_[9186]_ , \new_[9187]_ , \new_[9188]_ ,
    \new_[9189]_ , \new_[9190]_ , \new_[9191]_ , \new_[9192]_ ,
    \new_[9193]_ , \new_[9194]_ , \new_[9195]_ , \new_[9196]_ ,
    \new_[9197]_ , \new_[9198]_ , \new_[9199]_ , \new_[9200]_ ,
    \new_[9201]_ , \new_[9202]_ , \new_[9204]_ , \new_[9205]_ ,
    \new_[9206]_ , \new_[9207]_ , \new_[9208]_ , \new_[9209]_ ,
    \new_[9210]_ , \new_[9211]_ , \new_[9212]_ , \new_[9213]_ ,
    \new_[9214]_ , \new_[9215]_ , \new_[9216]_ , \new_[9217]_ ,
    \new_[9218]_ , \new_[9219]_ , \new_[9220]_ , \new_[9221]_ ,
    \new_[9222]_ , \new_[9223]_ , \new_[9224]_ , \new_[9225]_ ,
    \new_[9226]_ , \new_[9227]_ , \new_[9228]_ , \new_[9229]_ ,
    \new_[9230]_ , \new_[9231]_ , \new_[9232]_ , \new_[9233]_ ,
    \new_[9234]_ , \new_[9235]_ , \new_[9236]_ , \new_[9237]_ ,
    \new_[9238]_ , \new_[9239]_ , \new_[9240]_ , \new_[9241]_ ,
    \new_[9242]_ , \new_[9243]_ , \new_[9244]_ , \new_[9245]_ ,
    \new_[9246]_ , \new_[9247]_ , \new_[9248]_ , \new_[9249]_ ,
    \new_[9250]_ , \new_[9251]_ , \new_[9252]_ , \new_[9253]_ ,
    \new_[9254]_ , \new_[9255]_ , \new_[9256]_ , \new_[9257]_ ,
    \new_[9258]_ , \new_[9259]_ , \new_[9260]_ , \new_[9261]_ ,
    \new_[9262]_ , \new_[9263]_ , \new_[9264]_ , \new_[9265]_ ,
    \new_[9266]_ , \new_[9267]_ , \new_[9268]_ , \new_[9269]_ ,
    \new_[9270]_ , \new_[9271]_ , \new_[9272]_ , \new_[9273]_ ,
    \new_[9274]_ , \new_[9275]_ , \new_[9276]_ , \new_[9277]_ ,
    \new_[9278]_ , \new_[9279]_ , \new_[9280]_ , \new_[9281]_ ,
    \new_[9282]_ , \new_[9283]_ , \new_[9284]_ , \new_[9285]_ ,
    \new_[9286]_ , \new_[9287]_ , \new_[9288]_ , \new_[9289]_ ,
    \new_[9290]_ , \new_[9291]_ , \new_[9292]_ , \new_[9293]_ ,
    \new_[9294]_ , \new_[9295]_ , \new_[9296]_ , \new_[9297]_ ,
    \new_[9298]_ , \new_[9299]_ , \new_[9300]_ , \new_[9301]_ ,
    \new_[9302]_ , \new_[9303]_ , \new_[9304]_ , \new_[9305]_ ,
    \new_[9306]_ , \new_[9307]_ , \new_[9308]_ , \new_[9309]_ ,
    \new_[9310]_ , \new_[9311]_ , \new_[9312]_ , \new_[9313]_ ,
    \new_[9314]_ , \new_[9315]_ , \new_[9316]_ , \new_[9317]_ ,
    \new_[9318]_ , \new_[9319]_ , \new_[9320]_ , \new_[9321]_ ,
    \new_[9322]_ , \new_[9323]_ , \new_[9324]_ , \new_[9325]_ ,
    \new_[9326]_ , \new_[9327]_ , \new_[9328]_ , \new_[9329]_ ,
    \new_[9330]_ , \new_[9331]_ , \new_[9332]_ , \new_[9333]_ ,
    \new_[9334]_ , \new_[9335]_ , \new_[9336]_ , \new_[9337]_ ,
    \new_[9338]_ , \new_[9339]_ , \new_[9340]_ , \new_[9341]_ ,
    \new_[9342]_ , \new_[9343]_ , \new_[9344]_ , \new_[9345]_ ,
    \new_[9346]_ , \new_[9347]_ , \new_[9348]_ , \new_[9349]_ ,
    \new_[9350]_ , \new_[9351]_ , \new_[9352]_ , \new_[9353]_ ,
    \new_[9354]_ , \new_[9355]_ , \new_[9356]_ , \new_[9357]_ ,
    \new_[9358]_ , \new_[9359]_ , \new_[9360]_ , \new_[9361]_ ,
    \new_[9362]_ , \new_[9363]_ , \new_[9364]_ , \new_[9365]_ ,
    \new_[9366]_ , \new_[9367]_ , \new_[9368]_ , \new_[9369]_ ,
    \new_[9370]_ , \new_[9371]_ , \new_[9372]_ , \new_[9373]_ ,
    \new_[9374]_ , \new_[9375]_ , \new_[9376]_ , \new_[9377]_ ,
    \new_[9378]_ , \new_[9379]_ , \new_[9380]_ , \new_[9381]_ ,
    \new_[9382]_ , \new_[9383]_ , \new_[9384]_ , \new_[9385]_ ,
    \new_[9386]_ , \new_[9387]_ , \new_[9388]_ , \new_[9389]_ ,
    \new_[9390]_ , \new_[9391]_ , \new_[9392]_ , \new_[9393]_ ,
    \new_[9394]_ , \new_[9395]_ , \new_[9396]_ , \new_[9397]_ ,
    \new_[9398]_ , \new_[9399]_ , \new_[9400]_ , \new_[9401]_ ,
    \new_[9402]_ , \new_[9403]_ , \new_[9404]_ , \new_[9405]_ ,
    \new_[9406]_ , \new_[9407]_ , \new_[9408]_ , \new_[9409]_ ,
    \new_[9410]_ , \new_[9411]_ , \new_[9412]_ , \new_[9413]_ ,
    \new_[9414]_ , \new_[9415]_ , \new_[9416]_ , \new_[9417]_ ,
    \new_[9418]_ , \new_[9419]_ , \new_[9420]_ , \new_[9421]_ ,
    \new_[9422]_ , \new_[9423]_ , \new_[9424]_ , \new_[9425]_ ,
    \new_[9426]_ , \new_[9427]_ , \new_[9428]_ , \new_[9429]_ ,
    \new_[9430]_ , \new_[9431]_ , \new_[9432]_ , \new_[9433]_ ,
    \new_[9434]_ , \new_[9435]_ , \new_[9436]_ , \new_[9437]_ ,
    \new_[9438]_ , \new_[9439]_ , \new_[9440]_ , \new_[9441]_ ,
    \new_[9442]_ , \new_[9443]_ , \new_[9444]_ , \new_[9445]_ ,
    \new_[9446]_ , \new_[9447]_ , \new_[9448]_ , \new_[9449]_ ,
    \new_[9450]_ , \new_[9451]_ , \new_[9452]_ , \new_[9453]_ ,
    \new_[9454]_ , \new_[9455]_ , \new_[9456]_ , \new_[9457]_ ,
    \new_[9458]_ , \new_[9459]_ , \new_[9460]_ , \new_[9461]_ ,
    \new_[9462]_ , \new_[9463]_ , \new_[9464]_ , \new_[9465]_ ,
    \new_[9466]_ , \new_[9467]_ , \new_[9468]_ , \new_[9469]_ ,
    \new_[9470]_ , \new_[9471]_ , \new_[9472]_ , \new_[9473]_ ,
    \new_[9474]_ , \new_[9475]_ , \new_[9476]_ , \new_[9477]_ ,
    \new_[9478]_ , \new_[9479]_ , \new_[9480]_ , \new_[9481]_ ,
    \new_[9482]_ , \new_[9483]_ , \new_[9484]_ , \new_[9485]_ ,
    \new_[9486]_ , \new_[9487]_ , \new_[9488]_ , \new_[9489]_ ,
    \new_[9490]_ , \new_[9491]_ , \new_[9492]_ , \new_[9493]_ ,
    \new_[9494]_ , \new_[9495]_ , \new_[9496]_ , \new_[9497]_ ,
    \new_[9498]_ , \new_[9499]_ , \new_[9500]_ , \new_[9501]_ ,
    \new_[9502]_ , \new_[9503]_ , \new_[9504]_ , \new_[9505]_ ,
    \new_[9506]_ , \new_[9507]_ , \new_[9508]_ , \new_[9509]_ ,
    \new_[9510]_ , \new_[9511]_ , \new_[9512]_ , \new_[9513]_ ,
    \new_[9514]_ , \new_[9515]_ , \new_[9516]_ , \new_[9517]_ ,
    \new_[9518]_ , \new_[9519]_ , \new_[9520]_ , \new_[9521]_ ,
    \new_[9522]_ , \new_[9523]_ , \new_[9524]_ , \new_[9525]_ ,
    \new_[9526]_ , \new_[9527]_ , \new_[9528]_ , \new_[9529]_ ,
    \new_[9530]_ , \new_[9531]_ , \new_[9532]_ , \new_[9533]_ ,
    \new_[9534]_ , \new_[9535]_ , \new_[9536]_ , \new_[9537]_ ,
    \new_[9538]_ , \new_[9539]_ , \new_[9540]_ , \new_[9541]_ ,
    \new_[9542]_ , \new_[9543]_ , \new_[9544]_ , \new_[9545]_ ,
    \new_[9546]_ , \new_[9547]_ , \new_[9548]_ , \new_[9549]_ ,
    \new_[9550]_ , \new_[9551]_ , \new_[9552]_ , \new_[9553]_ ,
    \new_[9554]_ , \new_[9555]_ , \new_[9556]_ , \new_[9557]_ ,
    \new_[9558]_ , \new_[9559]_ , \new_[9560]_ , \new_[9561]_ ,
    \new_[9562]_ , \new_[9563]_ , \new_[9564]_ , \new_[9565]_ ,
    \new_[9566]_ , \new_[9567]_ , \new_[9568]_ , \new_[9569]_ ,
    \new_[9570]_ , \new_[9571]_ , \new_[9572]_ , \new_[9573]_ ,
    \new_[9574]_ , \new_[9575]_ , \new_[9576]_ , \new_[9577]_ ,
    \new_[9578]_ , \new_[9579]_ , \new_[9580]_ , \new_[9581]_ ,
    \new_[9582]_ , \new_[9583]_ , \new_[9584]_ , \new_[9585]_ ,
    \new_[9586]_ , \new_[9587]_ , \new_[9588]_ , \new_[9589]_ ,
    \new_[9590]_ , \new_[9591]_ , \new_[9592]_ , \new_[9593]_ ,
    \new_[9594]_ , \new_[9595]_ , \new_[9596]_ , \new_[9597]_ ,
    \new_[9598]_ , \new_[9599]_ , \new_[9600]_ , \new_[9601]_ ,
    \new_[9602]_ , \new_[9603]_ , \new_[9604]_ , \new_[9605]_ ,
    \new_[9606]_ , \new_[9607]_ , \new_[9608]_ , \new_[9609]_ ,
    \new_[9610]_ , \new_[9611]_ , \new_[9612]_ , \new_[9613]_ ,
    \new_[9614]_ , \new_[9615]_ , \new_[9616]_ , \new_[9617]_ ,
    \new_[9618]_ , \new_[9619]_ , \new_[9620]_ , \new_[9621]_ ,
    \new_[9622]_ , \new_[9623]_ , \new_[9624]_ , \new_[9625]_ ,
    \new_[9626]_ , \new_[9627]_ , \new_[9628]_ , \new_[9629]_ ,
    \new_[9630]_ , \new_[9631]_ , \new_[9632]_ , \new_[9633]_ ,
    \new_[9634]_ , \new_[9635]_ , \new_[9636]_ , \new_[9637]_ ,
    \new_[9638]_ , \new_[9639]_ , \new_[9640]_ , \new_[9641]_ ,
    \new_[9642]_ , \new_[9643]_ , \new_[9644]_ , \new_[9645]_ ,
    \new_[9647]_ , \new_[9648]_ , \new_[9649]_ , \new_[9650]_ ,
    \new_[9651]_ , \new_[9652]_ , \new_[9653]_ , \new_[9654]_ ,
    \new_[9655]_ , \new_[9656]_ , \new_[9660]_ , \new_[9661]_ ,
    \new_[9662]_ , \new_[9663]_ , \new_[9666]_ , \new_[9668]_ ,
    \new_[9669]_ , \new_[9670]_ , \new_[9672]_ , \new_[9673]_ ,
    \new_[9674]_ , \new_[9675]_ , \new_[9676]_ , \new_[9677]_ ,
    \new_[9682]_ , \new_[9683]_ , \new_[9697]_ , \new_[9698]_ ,
    \new_[9699]_ , \new_[9700]_ , \new_[9701]_ , \new_[9702]_ ,
    \new_[9703]_ , \new_[9704]_ , \new_[9705]_ , \new_[9706]_ ,
    \new_[9707]_ , \new_[9708]_ , \new_[9709]_ , \new_[9710]_ ,
    \new_[9711]_ , \new_[9712]_ , \new_[9713]_ , \new_[9714]_ ,
    \new_[9715]_ , \new_[9716]_ , \new_[9717]_ , \new_[9718]_ ,
    \new_[9719]_ , \new_[9720]_ , \new_[9721]_ , \new_[9722]_ ,
    \new_[9723]_ , \new_[9724]_ , \new_[9725]_ , \new_[9726]_ ,
    \new_[9727]_ , \new_[9728]_ , \new_[9729]_ , \new_[9730]_ ,
    \new_[9731]_ , \new_[9732]_ , \new_[9733]_ , \new_[9734]_ ,
    \new_[9735]_ , \new_[9736]_ , \new_[9737]_ , \new_[9738]_ ,
    \new_[9739]_ , \new_[9740]_ , \new_[9741]_ , \new_[9742]_ ,
    \new_[9743]_ , \new_[9744]_ , \new_[9745]_ , \new_[9746]_ ,
    \new_[9747]_ , \new_[9748]_ , \new_[9749]_ , \new_[9750]_ ,
    \new_[9751]_ , \new_[9752]_ , \new_[9753]_ , \new_[9754]_ ,
    \new_[9755]_ , \new_[9756]_ , \new_[9757]_ , \new_[9758]_ ,
    \new_[9759]_ , \new_[9760]_ , \new_[9761]_ , \new_[9762]_ ,
    \new_[9763]_ , \new_[9764]_ , \new_[9765]_ , \new_[9766]_ ,
    \new_[9767]_ , \new_[9768]_ , \new_[9769]_ , \new_[9770]_ ,
    \new_[9771]_ , \new_[9772]_ , \new_[9773]_ , \new_[9774]_ ,
    \new_[9775]_ , \new_[9776]_ , \new_[9777]_ , \new_[9778]_ ,
    \new_[9779]_ , \new_[9780]_ , \new_[9781]_ , \new_[9782]_ ,
    \new_[9783]_ , \new_[9784]_ , \new_[9785]_ , \new_[9786]_ ,
    \new_[9787]_ , \new_[9788]_ , \new_[9789]_ , \new_[9790]_ ,
    \new_[9791]_ , \new_[9792]_ , \new_[9793]_ , \new_[9794]_ ,
    \new_[9795]_ , \new_[9796]_ , \new_[9797]_ , \new_[9798]_ ,
    \new_[9799]_ , \new_[9800]_ , \new_[9801]_ , \new_[9802]_ ,
    \new_[9803]_ , \new_[9804]_ , \new_[9805]_ , \new_[9806]_ ,
    \new_[9807]_ , \new_[9808]_ , \new_[9809]_ , \new_[9810]_ ,
    \new_[9811]_ , \new_[9812]_ , \new_[9813]_ , \new_[9814]_ ,
    \new_[9815]_ , \new_[9816]_ , \new_[9817]_ , \new_[9818]_ ,
    \new_[9819]_ , \new_[9820]_ , \new_[9821]_ , \new_[9822]_ ,
    \new_[9823]_ , \new_[9824]_ , \new_[9825]_ , \new_[9826]_ ,
    \new_[9827]_ , \new_[9828]_ , \new_[9829]_ , \new_[9830]_ ,
    \new_[9831]_ , \new_[9832]_ , \new_[9833]_ , \new_[9834]_ ,
    \new_[9835]_ , \new_[9836]_ , \new_[9837]_ , \new_[9838]_ ,
    \new_[9839]_ , \new_[9840]_ , \new_[9841]_ , \new_[9842]_ ,
    \new_[9843]_ , \new_[9844]_ , \new_[9845]_ , \new_[9846]_ ,
    \new_[9847]_ , \new_[9848]_ , \new_[9849]_ , \new_[9850]_ ,
    \new_[9851]_ , \new_[9852]_ , \new_[9853]_ , \new_[9854]_ ,
    \new_[9855]_ , \new_[9856]_ , \new_[9857]_ , \new_[9858]_ ,
    \new_[9859]_ , \new_[9860]_ , \new_[9861]_ , \new_[9862]_ ,
    \new_[9863]_ , \new_[9864]_ , \new_[9865]_ , \new_[9866]_ ,
    \new_[9867]_ , \new_[9868]_ , \new_[9869]_ , \new_[9870]_ ,
    \new_[9871]_ , \new_[9872]_ , \new_[9873]_ , \new_[9874]_ ,
    \new_[9875]_ , \new_[9876]_ , \new_[9877]_ , \new_[9878]_ ,
    \new_[9879]_ , \new_[9880]_ , \new_[9881]_ , \new_[9882]_ ,
    \new_[9883]_ , \new_[9884]_ , \new_[9885]_ , \new_[9886]_ ,
    \new_[9887]_ , \new_[9888]_ , \new_[9889]_ , \new_[9890]_ ,
    \new_[9891]_ , \new_[9892]_ , \new_[9893]_ , \new_[9894]_ ,
    \new_[9895]_ , \new_[9896]_ , \new_[9897]_ , \new_[9898]_ ,
    \new_[9899]_ , \new_[9900]_ , \new_[9901]_ , \new_[9902]_ ,
    \new_[9903]_ , \new_[9904]_ , \new_[9905]_ , \new_[9906]_ ,
    \new_[9907]_ , \new_[9908]_ , \new_[9909]_ , \new_[9910]_ ,
    \new_[9911]_ , \new_[9912]_ , \new_[9913]_ , \new_[9914]_ ,
    \new_[9915]_ , \new_[9916]_ , \new_[9917]_ , \new_[9918]_ ,
    \new_[9919]_ , \new_[9920]_ , \new_[9921]_ , \new_[9922]_ ,
    \new_[9923]_ , \new_[9924]_ , \new_[9925]_ , \new_[9926]_ ,
    \new_[9927]_ , \new_[9928]_ , \new_[9929]_ , \new_[9930]_ ,
    \new_[9931]_ , \new_[9932]_ , \new_[9933]_ , \new_[9934]_ ,
    \new_[9935]_ , \new_[9936]_ , \new_[9937]_ , \new_[9938]_ ,
    \new_[9939]_ , \new_[9940]_ , \new_[9941]_ , \new_[9942]_ ,
    \new_[9943]_ , \new_[9944]_ , \new_[9945]_ , \new_[9946]_ ,
    \new_[9947]_ , \new_[9948]_ , \new_[9949]_ , \new_[9950]_ ,
    \new_[9951]_ , \new_[9952]_ , \new_[9953]_ , \new_[9954]_ ,
    \new_[9955]_ , \new_[9956]_ , \new_[9957]_ , \new_[9958]_ ,
    \new_[9959]_ , \new_[9960]_ , \new_[9961]_ , \new_[9962]_ ,
    \new_[9963]_ , \new_[9964]_ , \new_[9965]_ , \new_[9966]_ ,
    \new_[9967]_ , \new_[9968]_ , \new_[9969]_ , \new_[9970]_ ,
    \new_[9971]_ , \new_[9972]_ , \new_[9973]_ , \new_[9974]_ ,
    \new_[9975]_ , \new_[9976]_ , \new_[9977]_ , \new_[9978]_ ,
    \new_[9979]_ , \new_[9980]_ , \new_[9981]_ , \new_[9982]_ ,
    \new_[9983]_ , \new_[9984]_ , \new_[9985]_ , \new_[9986]_ ,
    \new_[9987]_ , \new_[9988]_ , \new_[9989]_ , \new_[9990]_ ,
    \new_[9991]_ , \new_[9992]_ , \new_[9993]_ , \new_[9994]_ ,
    \new_[9995]_ , \new_[9996]_ , \new_[9997]_ , \new_[9998]_ ,
    \new_[9999]_ , \new_[10000]_ , \new_[10001]_ , \new_[10002]_ ,
    \new_[10003]_ , \new_[10004]_ , \new_[10005]_ , \new_[10006]_ ,
    \new_[10007]_ , \new_[10008]_ , \new_[10009]_ , \new_[10010]_ ,
    \new_[10011]_ , \new_[10012]_ , \new_[10013]_ , \new_[10014]_ ,
    \new_[10015]_ , \new_[10016]_ , \new_[10017]_ , \new_[10018]_ ,
    \new_[10019]_ , \new_[10020]_ , \new_[10021]_ , \new_[10022]_ ,
    \new_[10023]_ , \new_[10024]_ , \new_[10025]_ , \new_[10026]_ ,
    \new_[10027]_ , \new_[10028]_ , \new_[10029]_ , \new_[10030]_ ,
    \new_[10031]_ , \new_[10032]_ , \new_[10033]_ , \new_[10034]_ ,
    \new_[10035]_ , \new_[10036]_ , \new_[10037]_ , \new_[10038]_ ,
    \new_[10039]_ , \new_[10040]_ , \new_[10041]_ , \new_[10042]_ ,
    \new_[10043]_ , \new_[10044]_ , \new_[10045]_ , \new_[10046]_ ,
    \new_[10047]_ , \new_[10048]_ , \new_[10049]_ , \new_[10050]_ ,
    \new_[10051]_ , \new_[10052]_ , \new_[10053]_ , \new_[10054]_ ,
    \new_[10055]_ , \new_[10056]_ , \new_[10057]_ , \new_[10058]_ ,
    \new_[10059]_ , \new_[10060]_ , \new_[10061]_ , \new_[10062]_ ,
    \new_[10063]_ , \new_[10064]_ , \new_[10065]_ , \new_[10066]_ ,
    \new_[10067]_ , \new_[10068]_ , \new_[10069]_ , \new_[10070]_ ,
    \new_[10071]_ , \new_[10072]_ , \new_[10073]_ , \new_[10074]_ ,
    \new_[10075]_ , \new_[10076]_ , \new_[10077]_ , \new_[10078]_ ,
    \new_[10079]_ , \new_[10080]_ , \new_[10081]_ , \new_[10082]_ ,
    \new_[10083]_ , \new_[10084]_ , \new_[10086]_ , \new_[10087]_ ,
    \new_[10088]_ , \new_[10089]_ , \new_[10090]_ , \new_[10091]_ ,
    \new_[10092]_ , \new_[10093]_ , \new_[10094]_ , \new_[10095]_ ,
    \new_[10096]_ , \new_[10097]_ , \new_[10098]_ , \new_[10099]_ ,
    \new_[10100]_ , \new_[10101]_ , \new_[10102]_ , \new_[10103]_ ,
    \new_[10104]_ , \new_[10105]_ , \new_[10106]_ , \new_[10107]_ ,
    \new_[10108]_ , \new_[10109]_ , \new_[10110]_ , \new_[10111]_ ,
    \new_[10112]_ , \new_[10113]_ , \new_[10114]_ , \new_[10115]_ ,
    \new_[10116]_ , \new_[10117]_ , \new_[10118]_ , \new_[10119]_ ,
    \new_[10120]_ , \new_[10121]_ , \new_[10122]_ , \new_[10123]_ ,
    \new_[10124]_ , \new_[10125]_ , \new_[10126]_ , \new_[10127]_ ,
    \new_[10128]_ , \new_[10129]_ , \new_[10130]_ , \new_[10131]_ ,
    \new_[10132]_ , \new_[10133]_ , \new_[10134]_ , \new_[10135]_ ,
    \new_[10136]_ , \new_[10137]_ , \new_[10138]_ , \new_[10139]_ ,
    \new_[10140]_ , \new_[10141]_ , \new_[10142]_ , \new_[10143]_ ,
    \new_[10144]_ , \new_[10145]_ , \new_[10146]_ , \new_[10147]_ ,
    \new_[10148]_ , \new_[10149]_ , \new_[10150]_ , \new_[10151]_ ,
    \new_[10152]_ , \new_[10153]_ , \new_[10154]_ , \new_[10155]_ ,
    \new_[10156]_ , \new_[10157]_ , \new_[10158]_ , \new_[10159]_ ,
    \new_[10160]_ , \new_[10161]_ , \new_[10162]_ , \new_[10163]_ ,
    \new_[10164]_ , \new_[10165]_ , \new_[10166]_ , \new_[10167]_ ,
    \new_[10168]_ , \new_[10169]_ , \new_[10170]_ , \new_[10171]_ ,
    \new_[10172]_ , \new_[10173]_ , \new_[10174]_ , \new_[10175]_ ,
    \new_[10176]_ , \new_[10177]_ , \new_[10178]_ , \new_[10179]_ ,
    \new_[10180]_ , \new_[10181]_ , \new_[10182]_ , \new_[10183]_ ,
    \new_[10184]_ , \new_[10185]_ , \new_[10186]_ , \new_[10187]_ ,
    \new_[10188]_ , \new_[10189]_ , \new_[10190]_ , \new_[10191]_ ,
    \new_[10192]_ , \new_[10193]_ , \new_[10194]_ , \new_[10195]_ ,
    \new_[10196]_ , \new_[10197]_ , \new_[10198]_ , \new_[10199]_ ,
    \new_[10200]_ , \new_[10201]_ , \new_[10202]_ , \new_[10203]_ ,
    \new_[10204]_ , \new_[10205]_ , \new_[10206]_ , \new_[10207]_ ,
    \new_[10208]_ , \new_[10209]_ , \new_[10210]_ , \new_[10211]_ ,
    \new_[10212]_ , \new_[10213]_ , \new_[10214]_ , \new_[10215]_ ,
    \new_[10216]_ , \new_[10217]_ , \new_[10218]_ , \new_[10219]_ ,
    \new_[10220]_ , \new_[10221]_ , \new_[10222]_ , \new_[10223]_ ,
    \new_[10224]_ , \new_[10225]_ , \new_[10226]_ , \new_[10227]_ ,
    \new_[10228]_ , \new_[10229]_ , \new_[10230]_ , \new_[10231]_ ,
    \new_[10232]_ , \new_[10233]_ , \new_[10234]_ , \new_[10235]_ ,
    \new_[10236]_ , \new_[10237]_ , \new_[10238]_ , \new_[10239]_ ,
    \new_[10240]_ , \new_[10241]_ , \new_[10242]_ , \new_[10243]_ ,
    \new_[10244]_ , \new_[10245]_ , \new_[10246]_ , \new_[10247]_ ,
    \new_[10248]_ , \new_[10249]_ , \new_[10250]_ , \new_[10251]_ ,
    \new_[10252]_ , \new_[10253]_ , \new_[10254]_ , \new_[10255]_ ,
    \new_[10256]_ , \new_[10257]_ , \new_[10258]_ , \new_[10259]_ ,
    \new_[10260]_ , \new_[10261]_ , \new_[10262]_ , \new_[10263]_ ,
    \new_[10264]_ , \new_[10265]_ , \new_[10266]_ , \new_[10267]_ ,
    \new_[10268]_ , \new_[10269]_ , \new_[10270]_ , \new_[10271]_ ,
    \new_[10272]_ , \new_[10273]_ , \new_[10274]_ , \new_[10275]_ ,
    \new_[10276]_ , \new_[10277]_ , \new_[10278]_ , \new_[10279]_ ,
    \new_[10280]_ , \new_[10281]_ , \new_[10282]_ , \new_[10283]_ ,
    \new_[10284]_ , \new_[10285]_ , \new_[10286]_ , \new_[10288]_ ,
    \new_[10290]_ , \new_[10291]_ , \new_[10292]_ , \new_[10293]_ ,
    \new_[10294]_ , \new_[10297]_ , \new_[10298]_ , \new_[10299]_ ,
    \new_[10300]_ , \new_[10301]_ , \new_[10302]_ , \new_[10303]_ ,
    \new_[10305]_ , \new_[10306]_ , \new_[10307]_ , \new_[10308]_ ,
    \new_[10309]_ , \new_[10310]_ , \new_[10311]_ , \new_[10313]_ ,
    \new_[10314]_ , \new_[10315]_ , \new_[10316]_ , \new_[10317]_ ,
    \new_[10318]_ , \new_[10319]_ , \new_[10320]_ , \new_[10321]_ ,
    \new_[10354]_ , \new_[10355]_ , \new_[10390]_ , \new_[10394]_ ,
    \new_[10395]_ , \new_[10396]_ , \new_[10397]_ , \new_[10398]_ ,
    \new_[10399]_ , \new_[10401]_ , \new_[10402]_ , \new_[10403]_ ,
    \new_[10404]_ , \new_[10405]_ , \new_[10406]_ , \new_[10407]_ ,
    \new_[10408]_ , \new_[10409]_ , \new_[10410]_ , \new_[10411]_ ,
    \new_[10412]_ , \new_[10413]_ , \new_[10414]_ , \new_[10415]_ ,
    \new_[10416]_ , \new_[10417]_ , \new_[10418]_ , \new_[10419]_ ,
    \new_[10420]_ , \new_[10421]_ , \new_[10422]_ , \new_[10423]_ ,
    \new_[10424]_ , \new_[10425]_ , \new_[10426]_ , \new_[10427]_ ,
    \new_[10428]_ , \new_[10429]_ , \new_[10430]_ , \new_[10431]_ ,
    \new_[10432]_ , \new_[10433]_ , \new_[10434]_ , \new_[10435]_ ,
    \new_[10436]_ , \new_[10437]_ , \new_[10438]_ , \new_[10439]_ ,
    \new_[10440]_ , \new_[10441]_ , \new_[10442]_ , \new_[10443]_ ,
    \new_[10444]_ , \new_[10445]_ , \new_[10446]_ , \new_[10447]_ ,
    \new_[10448]_ , \new_[10449]_ , \new_[10450]_ , \new_[10451]_ ,
    \new_[10452]_ , \new_[10453]_ , \new_[10454]_ , \new_[10455]_ ,
    \new_[10456]_ , \new_[10457]_ , \new_[10458]_ , \new_[10459]_ ,
    \new_[10460]_ , \new_[10461]_ , \new_[10462]_ , \new_[10463]_ ,
    \new_[10464]_ , \new_[10465]_ , \new_[10466]_ , \new_[10467]_ ,
    \new_[10468]_ , \new_[10469]_ , \new_[10470]_ , \new_[10471]_ ,
    \new_[10472]_ , \new_[10473]_ , \new_[10474]_ , \new_[10475]_ ,
    \new_[10476]_ , \new_[10477]_ , \new_[10478]_ , \new_[10479]_ ,
    \new_[10480]_ , \new_[10481]_ , \new_[10482]_ , \new_[10483]_ ,
    \new_[10484]_ , \new_[10485]_ , \new_[10486]_ , \new_[10487]_ ,
    \new_[10488]_ , \new_[10489]_ , \new_[10490]_ , \new_[10491]_ ,
    \new_[10492]_ , \new_[10493]_ , \new_[10494]_ , \new_[10495]_ ,
    \new_[10496]_ , \new_[10497]_ , \new_[10498]_ , \new_[10499]_ ,
    \new_[10500]_ , \new_[10501]_ , \new_[10502]_ , \new_[10503]_ ,
    \new_[10504]_ , \new_[10505]_ , \new_[10506]_ , \new_[10507]_ ,
    \new_[10508]_ , \new_[10509]_ , \new_[10510]_ , \new_[10511]_ ,
    \new_[10512]_ , \new_[10513]_ , \new_[10514]_ , \new_[10515]_ ,
    \new_[10516]_ , \new_[10517]_ , \new_[10518]_ , \new_[10519]_ ,
    \new_[10520]_ , \new_[10521]_ , \new_[10522]_ , \new_[10523]_ ,
    \new_[10524]_ , \new_[10525]_ , \new_[10526]_ , \new_[10527]_ ,
    \new_[10528]_ , \new_[10529]_ , \new_[10530]_ , \new_[10531]_ ,
    \new_[10532]_ , \new_[10533]_ , \new_[10534]_ , \new_[10535]_ ,
    \new_[10536]_ , \new_[10537]_ , \new_[10538]_ , \new_[10539]_ ,
    \new_[10540]_ , \new_[10541]_ , \new_[10542]_ , \new_[10543]_ ,
    \new_[10544]_ , \new_[10545]_ , \new_[10546]_ , \new_[10547]_ ,
    \new_[10548]_ , \new_[10549]_ , \new_[10550]_ , \new_[10551]_ ,
    \new_[10552]_ , \new_[10553]_ , \new_[10554]_ , \new_[10555]_ ,
    \new_[10556]_ , \new_[10557]_ , \new_[10558]_ , \new_[10559]_ ,
    \new_[10560]_ , \new_[10561]_ , \new_[10562]_ , \new_[10563]_ ,
    \new_[10564]_ , \new_[10565]_ , \new_[10566]_ , \new_[10567]_ ,
    \new_[10568]_ , \new_[10569]_ , \new_[10570]_ , \new_[10571]_ ,
    \new_[10572]_ , \new_[10573]_ , \new_[10574]_ , \new_[10575]_ ,
    \new_[10576]_ , \new_[10577]_ , \new_[10578]_ , \new_[10579]_ ,
    \new_[10580]_ , \new_[10581]_ , \new_[10582]_ , \new_[10583]_ ,
    \new_[10584]_ , \new_[10585]_ , \new_[10586]_ , \new_[10587]_ ,
    \new_[10588]_ , \new_[10589]_ , \new_[10590]_ , \new_[10591]_ ,
    \new_[10592]_ , \new_[10593]_ , \new_[10594]_ , \new_[10595]_ ,
    \new_[10596]_ , \new_[10597]_ , \new_[10598]_ , \new_[10599]_ ,
    \new_[10600]_ , \new_[10601]_ , \new_[10602]_ , \new_[10603]_ ,
    \new_[10604]_ , \new_[10605]_ , \new_[10606]_ , \new_[10607]_ ,
    \new_[10608]_ , \new_[10609]_ , \new_[10610]_ , \new_[10611]_ ,
    \new_[10612]_ , \new_[10613]_ , \new_[10614]_ , \new_[10615]_ ,
    \new_[10616]_ , \new_[10617]_ , \new_[10618]_ , \new_[10619]_ ,
    \new_[10620]_ , \new_[10621]_ , \new_[10622]_ , \new_[10623]_ ,
    \new_[10624]_ , \new_[10625]_ , \new_[10626]_ , \new_[10627]_ ,
    \new_[10628]_ , \new_[10629]_ , \new_[10630]_ , \new_[10631]_ ,
    \new_[10632]_ , \new_[10633]_ , \new_[10634]_ , \new_[10635]_ ,
    \new_[10636]_ , \new_[10637]_ , \new_[10638]_ , \new_[10639]_ ,
    \new_[10640]_ , \new_[10641]_ , \new_[10642]_ , \new_[10643]_ ,
    \new_[10644]_ , \new_[10645]_ , \new_[10646]_ , \new_[10647]_ ,
    \new_[10648]_ , \new_[10649]_ , \new_[10650]_ , \new_[10651]_ ,
    \new_[10652]_ , \new_[10653]_ , \new_[10654]_ , \new_[10655]_ ,
    \new_[10656]_ , \new_[10657]_ , \new_[10658]_ , \new_[10659]_ ,
    \new_[10660]_ , \new_[10661]_ , \new_[10662]_ , \new_[10663]_ ,
    \new_[10664]_ , \new_[10665]_ , \new_[10666]_ , \new_[10667]_ ,
    \new_[10668]_ , \new_[10669]_ , \new_[10670]_ , \new_[10671]_ ,
    \new_[10672]_ , \new_[10673]_ , \new_[10674]_ , \new_[10675]_ ,
    \new_[10676]_ , \new_[10677]_ , \new_[10678]_ , \new_[10679]_ ,
    \new_[10680]_ , \new_[10681]_ , \new_[10682]_ , \new_[10683]_ ,
    \new_[10684]_ , \new_[10685]_ , \new_[10686]_ , \new_[10687]_ ,
    \new_[10688]_ , \new_[10689]_ , \new_[10690]_ , \new_[10691]_ ,
    \new_[10692]_ , \new_[10693]_ , \new_[10694]_ , \new_[10695]_ ,
    \new_[10696]_ , \new_[10697]_ , \new_[10698]_ , \new_[10699]_ ,
    \new_[10700]_ , \new_[10701]_ , \new_[10702]_ , \new_[10703]_ ,
    \new_[10704]_ , \new_[10705]_ , \new_[10706]_ , \new_[10707]_ ,
    \new_[10708]_ , \new_[10709]_ , \new_[10710]_ , \new_[10711]_ ,
    \new_[10712]_ , \new_[10715]_ , \new_[10716]_ , \new_[10717]_ ,
    \new_[10718]_ , \new_[10719]_ , \new_[10720]_ , \new_[10721]_ ,
    \new_[10722]_ , \new_[10723]_ , \new_[10724]_ , \new_[10725]_ ,
    \new_[10726]_ , \new_[10727]_ , \new_[10728]_ , \new_[10729]_ ,
    \new_[10730]_ , \new_[10731]_ , \new_[10732]_ , \new_[10733]_ ,
    \new_[10734]_ , \new_[10735]_ , \new_[10736]_ , \new_[10737]_ ,
    \new_[10738]_ , \new_[10739]_ , \new_[10740]_ , \new_[10741]_ ,
    \new_[10742]_ , \new_[10743]_ , \new_[10744]_ , \new_[10745]_ ,
    \new_[10746]_ , \new_[10747]_ , \new_[10748]_ , \new_[10749]_ ,
    \new_[10750]_ , \new_[10751]_ , \new_[10752]_ , \new_[10753]_ ,
    \new_[10754]_ , \new_[10755]_ , \new_[10756]_ , \new_[10757]_ ,
    \new_[10758]_ , \new_[10759]_ , \new_[10760]_ , \new_[10761]_ ,
    \new_[10762]_ , \new_[10763]_ , \new_[10764]_ , \new_[10765]_ ,
    \new_[10766]_ , \new_[10767]_ , \new_[10768]_ , \new_[10769]_ ,
    \new_[10770]_ , \new_[10771]_ , \new_[10772]_ , \new_[10773]_ ,
    \new_[10774]_ , \new_[10775]_ , \new_[10776]_ , \new_[10777]_ ,
    \new_[10778]_ , \new_[10779]_ , \new_[10780]_ , \new_[10781]_ ,
    \new_[10782]_ , \new_[10783]_ , \new_[10784]_ , \new_[10785]_ ,
    \new_[10786]_ , \new_[10787]_ , \new_[10788]_ , \new_[10789]_ ,
    \new_[10790]_ , \new_[10791]_ , \new_[10792]_ , \new_[10793]_ ,
    \new_[10794]_ , \new_[10795]_ , \new_[10796]_ , \new_[10797]_ ,
    \new_[10798]_ , \new_[10799]_ , \new_[10800]_ , \new_[10801]_ ,
    \new_[10802]_ , \new_[10803]_ , \new_[10804]_ , \new_[10805]_ ,
    \new_[10806]_ , \new_[10807]_ , \new_[10808]_ , \new_[10809]_ ,
    \new_[10810]_ , \new_[10811]_ , \new_[10812]_ , \new_[10813]_ ,
    \new_[10814]_ , \new_[10815]_ , \new_[10816]_ , \new_[10817]_ ,
    \new_[10818]_ , \new_[10819]_ , \new_[10820]_ , \new_[10821]_ ,
    \new_[10822]_ , \new_[10823]_ , \new_[10824]_ , \new_[10825]_ ,
    \new_[10826]_ , \new_[10827]_ , \new_[10828]_ , \new_[10829]_ ,
    \new_[10830]_ , \new_[10831]_ , \new_[10832]_ , \new_[10833]_ ,
    \new_[10834]_ , \new_[10835]_ , \new_[10836]_ , \new_[10837]_ ,
    \new_[10838]_ , \new_[10839]_ , \new_[10840]_ , \new_[10841]_ ,
    \new_[10842]_ , \new_[10843]_ , \new_[10844]_ , \new_[10845]_ ,
    \new_[10846]_ , \new_[10847]_ , \new_[10848]_ , \new_[10849]_ ,
    \new_[10850]_ , \new_[10851]_ , \new_[10852]_ , \new_[10853]_ ,
    \new_[10854]_ , \new_[10855]_ , \new_[10856]_ , \new_[10857]_ ,
    \new_[10858]_ , \new_[10859]_ , \new_[10860]_ , \new_[10861]_ ,
    \new_[10862]_ , \new_[10863]_ , \new_[10864]_ , \new_[10865]_ ,
    \new_[10866]_ , \new_[10867]_ , \new_[10868]_ , \new_[10869]_ ,
    \new_[10870]_ , \new_[10871]_ , \new_[10872]_ , \new_[10873]_ ,
    \new_[10874]_ , \new_[10875]_ , \new_[10876]_ , \new_[10877]_ ,
    \new_[10878]_ , \new_[10879]_ , \new_[10880]_ , \new_[10881]_ ,
    \new_[10882]_ , \new_[10883]_ , \new_[10884]_ , \new_[10885]_ ,
    \new_[10886]_ , \new_[10887]_ , \new_[10888]_ , \new_[10889]_ ,
    \new_[10890]_ , \new_[10891]_ , \new_[10892]_ , \new_[10893]_ ,
    \new_[10894]_ , \new_[10895]_ , \new_[10896]_ , \new_[10897]_ ,
    \new_[10898]_ , \new_[10899]_ , \new_[10900]_ , \new_[10901]_ ,
    \new_[10902]_ , \new_[10903]_ , \new_[10904]_ , \new_[10905]_ ,
    \new_[10906]_ , \new_[10907]_ , \new_[10908]_ , \new_[10909]_ ,
    \new_[10910]_ , \new_[10911]_ , \new_[10912]_ , \new_[10913]_ ,
    \new_[10914]_ , \new_[10915]_ , \new_[10916]_ , \new_[10917]_ ,
    \new_[10918]_ , \new_[10919]_ , \new_[10920]_ , \new_[10921]_ ,
    \new_[10922]_ , \new_[10923]_ , \new_[10924]_ , \new_[10925]_ ,
    \new_[10926]_ , \new_[10927]_ , \new_[10928]_ , \new_[10929]_ ,
    \new_[10930]_ , \new_[10931]_ , \new_[10932]_ , \new_[10933]_ ,
    \new_[10934]_ , \new_[10935]_ , \new_[10936]_ , \new_[10937]_ ,
    \new_[10938]_ , \new_[10939]_ , \new_[10940]_ , \new_[10941]_ ,
    \new_[10942]_ , \new_[10943]_ , \new_[10944]_ , \new_[10945]_ ,
    \new_[10946]_ , \new_[10947]_ , \new_[10948]_ , \new_[10949]_ ,
    \new_[10950]_ , \new_[10951]_ , \new_[10952]_ , \new_[10953]_ ,
    \new_[10954]_ , \new_[10955]_ , \new_[10956]_ , \new_[10957]_ ,
    \new_[10958]_ , \new_[10959]_ , \new_[10960]_ , \new_[10961]_ ,
    \new_[10962]_ , \new_[10963]_ , \new_[10964]_ , \new_[10965]_ ,
    \new_[10966]_ , \new_[10967]_ , \new_[10968]_ , \new_[10969]_ ,
    \new_[10970]_ , \new_[10971]_ , \new_[10972]_ , \new_[10973]_ ,
    \new_[10974]_ , \new_[10975]_ , \new_[10976]_ , \new_[10977]_ ,
    \new_[10978]_ , \new_[10979]_ , \new_[10980]_ , \new_[10981]_ ,
    \new_[10982]_ , \new_[10983]_ , \new_[10984]_ , \new_[10985]_ ,
    \new_[10986]_ , \new_[10987]_ , \new_[10988]_ , \new_[10989]_ ,
    \new_[10990]_ , \new_[10991]_ , \new_[10992]_ , \new_[10993]_ ,
    \new_[10994]_ , \new_[10995]_ , \new_[10996]_ , \new_[10997]_ ,
    \new_[10998]_ , \new_[10999]_ , \new_[11000]_ , \new_[11001]_ ,
    \new_[11002]_ , \new_[11003]_ , \new_[11004]_ , \new_[11005]_ ,
    \new_[11006]_ , \new_[11007]_ , \new_[11008]_ , \new_[11009]_ ,
    \new_[11010]_ , \new_[11011]_ , \new_[11012]_ , \new_[11013]_ ,
    \new_[11014]_ , \new_[11015]_ , \new_[11016]_ , \new_[11017]_ ,
    \new_[11018]_ , \new_[11019]_ , \new_[11020]_ , \new_[11021]_ ,
    \new_[11022]_ , \new_[11023]_ , \new_[11024]_ , \new_[11025]_ ,
    \new_[11026]_ , \new_[11027]_ , \new_[11028]_ , \new_[11029]_ ,
    \new_[11030]_ , \new_[11031]_ , \new_[11032]_ , \new_[11033]_ ,
    \new_[11034]_ , \new_[11035]_ , \new_[11036]_ , \new_[11037]_ ,
    \new_[11038]_ , \new_[11039]_ , \new_[11040]_ , \new_[11041]_ ,
    \new_[11042]_ , \new_[11043]_ , \new_[11044]_ , \new_[11045]_ ,
    \new_[11046]_ , \new_[11047]_ , \new_[11048]_ , \new_[11049]_ ,
    \new_[11050]_ , \new_[11051]_ , \new_[11052]_ , \new_[11053]_ ,
    \new_[11054]_ , \new_[11055]_ , \new_[11056]_ , \new_[11057]_ ,
    \new_[11058]_ , \new_[11059]_ , \new_[11060]_ , \new_[11061]_ ,
    \new_[11062]_ , \new_[11063]_ , \new_[11064]_ , \new_[11065]_ ,
    \new_[11066]_ , \new_[11067]_ , \new_[11068]_ , \new_[11069]_ ,
    \new_[11070]_ , \new_[11071]_ , \new_[11072]_ , \new_[11073]_ ,
    \new_[11074]_ , \new_[11075]_ , \new_[11076]_ , \new_[11077]_ ,
    \new_[11078]_ , \new_[11079]_ , \new_[11080]_ , \new_[11081]_ ,
    \new_[11082]_ , \new_[11083]_ , \new_[11084]_ , \new_[11085]_ ,
    \new_[11086]_ , \new_[11087]_ , \new_[11088]_ , \new_[11089]_ ,
    \new_[11090]_ , \new_[11091]_ , \new_[11092]_ , \new_[11093]_ ,
    \new_[11094]_ , \new_[11095]_ , \new_[11096]_ , \new_[11097]_ ,
    \new_[11098]_ , \new_[11099]_ , \new_[11100]_ , \new_[11101]_ ,
    \new_[11102]_ , \new_[11103]_ , \new_[11104]_ , \new_[11105]_ ,
    \new_[11106]_ , \new_[11107]_ , \new_[11108]_ , \new_[11109]_ ,
    \new_[11110]_ , \new_[11111]_ , \new_[11112]_ , \new_[11113]_ ,
    \new_[11114]_ , \new_[11115]_ , \new_[11116]_ , \new_[11117]_ ,
    \new_[11118]_ , \new_[11119]_ , \new_[11120]_ , \new_[11121]_ ,
    \new_[11122]_ , \new_[11123]_ , \new_[11124]_ , \new_[11125]_ ,
    \new_[11126]_ , \new_[11127]_ , \new_[11128]_ , \new_[11129]_ ,
    \new_[11130]_ , \new_[11131]_ , \new_[11132]_ , \new_[11133]_ ,
    \new_[11134]_ , \new_[11135]_ , \new_[11136]_ , \new_[11137]_ ,
    \new_[11138]_ , \new_[11139]_ , \new_[11140]_ , \new_[11141]_ ,
    \new_[11142]_ , \new_[11143]_ , \new_[11144]_ , \new_[11145]_ ,
    \new_[11146]_ , \new_[11147]_ , \new_[11148]_ , \new_[11149]_ ,
    \new_[11150]_ , \new_[11151]_ , \new_[11152]_ , \new_[11153]_ ,
    \new_[11154]_ , \new_[11155]_ , \new_[11156]_ , \new_[11157]_ ,
    \new_[11158]_ , \new_[11159]_ , \new_[11160]_ , \new_[11161]_ ,
    \new_[11162]_ , \new_[11163]_ , \new_[11164]_ , \new_[11165]_ ,
    \new_[11166]_ , \new_[11167]_ , \new_[11168]_ , \new_[11169]_ ,
    \new_[11170]_ , \new_[11171]_ , \new_[11172]_ , \new_[11173]_ ,
    \new_[11174]_ , \new_[11175]_ , \new_[11176]_ , \new_[11177]_ ,
    \new_[11178]_ , \new_[11179]_ , \new_[11180]_ , \new_[11181]_ ,
    \new_[11182]_ , \new_[11183]_ , \new_[11184]_ , \new_[11185]_ ,
    \new_[11186]_ , \new_[11187]_ , \new_[11188]_ , \new_[11189]_ ,
    \new_[11190]_ , \new_[11191]_ , \new_[11192]_ , \new_[11193]_ ,
    \new_[11194]_ , \new_[11195]_ , \new_[11196]_ , \new_[11197]_ ,
    \new_[11198]_ , \new_[11199]_ , \new_[11200]_ , \new_[11201]_ ,
    \new_[11202]_ , \new_[11203]_ , \new_[11204]_ , \new_[11205]_ ,
    \new_[11206]_ , \new_[11207]_ , \new_[11208]_ , \new_[11209]_ ,
    \new_[11210]_ , \new_[11211]_ , \new_[11212]_ , \new_[11213]_ ,
    \new_[11214]_ , \new_[11215]_ , \new_[11216]_ , \new_[11217]_ ,
    \new_[11218]_ , \new_[11219]_ , \new_[11220]_ , \new_[11221]_ ,
    \new_[11222]_ , \new_[11223]_ , \new_[11224]_ , \new_[11225]_ ,
    \new_[11226]_ , \new_[11227]_ , \new_[11228]_ , \new_[11229]_ ,
    \new_[11230]_ , \new_[11231]_ , \new_[11232]_ , \new_[11233]_ ,
    \new_[11234]_ , \new_[11235]_ , \new_[11236]_ , \new_[11237]_ ,
    \new_[11238]_ , \new_[11239]_ , \new_[11240]_ , \new_[11241]_ ,
    \new_[11242]_ , \new_[11243]_ , \new_[11244]_ , \new_[11245]_ ,
    \new_[11246]_ , \new_[11247]_ , \new_[11248]_ , \new_[11249]_ ,
    \new_[11250]_ , \new_[11251]_ , \new_[11252]_ , \new_[11253]_ ,
    \new_[11254]_ , \new_[11255]_ , \new_[11256]_ , \new_[11257]_ ,
    \new_[11258]_ , \new_[11259]_ , \new_[11260]_ , \new_[11261]_ ,
    \new_[11262]_ , \new_[11263]_ , \new_[11264]_ , \new_[11265]_ ,
    \new_[11266]_ , \new_[11267]_ , \new_[11268]_ , \new_[11269]_ ,
    \new_[11270]_ , \new_[11271]_ , \new_[11272]_ , \new_[11273]_ ,
    \new_[11274]_ , \new_[11275]_ , \new_[11276]_ , \new_[11277]_ ,
    \new_[11278]_ , \new_[11279]_ , \new_[11280]_ , \new_[11281]_ ,
    \new_[11282]_ , \new_[11283]_ , \new_[11284]_ , \new_[11285]_ ,
    \new_[11286]_ , \new_[11287]_ , \new_[11288]_ , \new_[11289]_ ,
    \new_[11290]_ , \new_[11291]_ , \new_[11292]_ , \new_[11293]_ ,
    \new_[11294]_ , \new_[11295]_ , \new_[11296]_ , \new_[11297]_ ,
    \new_[11298]_ , \new_[11299]_ , \new_[11300]_ , \new_[11301]_ ,
    \new_[11302]_ , \new_[11303]_ , \new_[11304]_ , \new_[11305]_ ,
    \new_[11306]_ , \new_[11307]_ , \new_[11308]_ , \new_[11309]_ ,
    \new_[11310]_ , \new_[11311]_ , \new_[11312]_ , \new_[11313]_ ,
    \new_[11314]_ , \new_[11315]_ , \new_[11316]_ , \new_[11317]_ ,
    \new_[11318]_ , \new_[11319]_ , \new_[11320]_ , \new_[11321]_ ,
    \new_[11322]_ , \new_[11323]_ , \new_[11324]_ , \new_[11325]_ ,
    \new_[11326]_ , \new_[11327]_ , \new_[11328]_ , \new_[11329]_ ,
    \new_[11330]_ , \new_[11331]_ , \new_[11332]_ , \new_[11333]_ ,
    \new_[11334]_ , \new_[11335]_ , \new_[11336]_ , \new_[11337]_ ,
    \new_[11338]_ , \new_[11339]_ , \new_[11340]_ , \new_[11341]_ ,
    \new_[11342]_ , \new_[11343]_ , \new_[11344]_ , \new_[11345]_ ,
    \new_[11346]_ , \new_[11347]_ , \new_[11348]_ , \new_[11349]_ ,
    \new_[11350]_ , \new_[11351]_ , \new_[11352]_ , \new_[11353]_ ,
    \new_[11354]_ , \new_[11355]_ , \new_[11356]_ , \new_[11357]_ ,
    \new_[11358]_ , \new_[11359]_ , \new_[11360]_ , \new_[11361]_ ,
    \new_[11362]_ , \new_[11363]_ , \new_[11364]_ , \new_[11365]_ ,
    \new_[11366]_ , \new_[11367]_ , \new_[11368]_ , \new_[11369]_ ,
    \new_[11370]_ , \new_[11371]_ , \new_[11372]_ , \new_[11373]_ ,
    \new_[11374]_ , \new_[11375]_ , \new_[11376]_ , \new_[11377]_ ,
    \new_[11378]_ , \new_[11379]_ , \new_[11380]_ , \new_[11381]_ ,
    \new_[11382]_ , \new_[11383]_ , \new_[11384]_ , \new_[11385]_ ,
    \new_[11386]_ , \new_[11387]_ , \new_[11388]_ , \new_[11389]_ ,
    \new_[11390]_ , \new_[11391]_ , \new_[11392]_ , \new_[11393]_ ,
    \new_[11394]_ , \new_[11395]_ , \new_[11396]_ , \new_[11397]_ ,
    \new_[11398]_ , \new_[11399]_ , \new_[11400]_ , \new_[11401]_ ,
    \new_[11402]_ , \new_[11403]_ , \new_[11404]_ , \new_[11405]_ ,
    \new_[11406]_ , \new_[11407]_ , \new_[11408]_ , \new_[11409]_ ,
    \new_[11410]_ , \new_[11411]_ , \new_[11412]_ , \new_[11413]_ ,
    \new_[11414]_ , \new_[11415]_ , \new_[11416]_ , \new_[11417]_ ,
    \new_[11418]_ , \new_[11419]_ , \new_[11420]_ , \new_[11421]_ ,
    \new_[11422]_ , \new_[11423]_ , \new_[11424]_ , \new_[11425]_ ,
    \new_[11426]_ , \new_[11427]_ , \new_[11428]_ , \new_[11429]_ ,
    \new_[11430]_ , \new_[11431]_ , \new_[11433]_ , \new_[11434]_ ,
    \new_[11435]_ , \new_[11436]_ , \new_[11437]_ , \new_[11438]_ ,
    \new_[11439]_ , \new_[11440]_ , \new_[11441]_ , \new_[11442]_ ,
    \new_[11443]_ , \new_[11444]_ , \new_[11445]_ , \new_[11446]_ ,
    \new_[11447]_ , \new_[11448]_ , \new_[11449]_ , \new_[11450]_ ,
    \new_[11452]_ , \new_[11453]_ , \new_[11454]_ , \new_[11456]_ ,
    \new_[11457]_ , \new_[11458]_ , \new_[11459]_ , \new_[11460]_ ,
    \new_[11461]_ , \new_[11462]_ , \new_[11463]_ , \new_[11464]_ ,
    \new_[11465]_ , \new_[11466]_ , \new_[11467]_ , \new_[11468]_ ,
    \new_[11469]_ , \new_[11470]_ , \new_[11471]_ , \new_[11472]_ ,
    \new_[11473]_ , \new_[11474]_ , \new_[11475]_ , \new_[11476]_ ,
    \new_[11477]_ , \new_[11478]_ , \new_[11479]_ , \new_[11480]_ ,
    \new_[11481]_ , \new_[11482]_ , \new_[11483]_ , \new_[11484]_ ,
    \new_[11485]_ , \new_[11486]_ , \new_[11487]_ , \new_[11488]_ ,
    \new_[11489]_ , \new_[11490]_ , \new_[11491]_ , \new_[11492]_ ,
    \new_[11493]_ , \new_[11494]_ , \new_[11495]_ , \new_[11496]_ ,
    \new_[11497]_ , \new_[11498]_ , \new_[11499]_ , \new_[11500]_ ,
    \new_[11501]_ , \new_[11502]_ , \new_[11503]_ , \new_[11504]_ ,
    \new_[11505]_ , \new_[11506]_ , \new_[11507]_ , \new_[11508]_ ,
    \new_[11509]_ , \new_[11510]_ , \new_[11511]_ , \new_[11512]_ ,
    \new_[11513]_ , \new_[11514]_ , \new_[11515]_ , \new_[11516]_ ,
    \new_[11517]_ , \new_[11518]_ , \new_[11519]_ , \new_[11520]_ ,
    \new_[11521]_ , \new_[11522]_ , \new_[11523]_ , \new_[11524]_ ,
    \new_[11525]_ , \new_[11526]_ , \new_[11527]_ , \new_[11528]_ ,
    \new_[11529]_ , \new_[11530]_ , \new_[11531]_ , \new_[11532]_ ,
    \new_[11533]_ , \new_[11534]_ , \new_[11535]_ , \new_[11536]_ ,
    \new_[11537]_ , \new_[11538]_ , \new_[11539]_ , \new_[11540]_ ,
    \new_[11541]_ , \new_[11542]_ , \new_[11543]_ , \new_[11544]_ ,
    \new_[11545]_ , \new_[11546]_ , \new_[11547]_ , \new_[11548]_ ,
    \new_[11549]_ , \new_[11550]_ , \new_[11551]_ , \new_[11552]_ ,
    \new_[11553]_ , \new_[11554]_ , \new_[11555]_ , \new_[11556]_ ,
    \new_[11557]_ , \new_[11558]_ , \new_[11559]_ , \new_[11560]_ ,
    \new_[11561]_ , \new_[11562]_ , \new_[11563]_ , \new_[11564]_ ,
    \new_[11565]_ , \new_[11566]_ , \new_[11567]_ , \new_[11568]_ ,
    \new_[11569]_ , \new_[11570]_ , \new_[11571]_ , \new_[11572]_ ,
    \new_[11573]_ , \new_[11574]_ , \new_[11575]_ , \new_[11576]_ ,
    \new_[11577]_ , \new_[11578]_ , \new_[11579]_ , \new_[11580]_ ,
    \new_[11581]_ , \new_[11582]_ , \new_[11583]_ , \new_[11584]_ ,
    \new_[11585]_ , \new_[11586]_ , \new_[11587]_ , \new_[11588]_ ,
    \new_[11589]_ , \new_[11590]_ , \new_[11591]_ , \new_[11592]_ ,
    \new_[11593]_ , \new_[11594]_ , \new_[11595]_ , \new_[11596]_ ,
    \new_[11597]_ , \new_[11598]_ , \new_[11599]_ , \new_[11600]_ ,
    \new_[11601]_ , \new_[11602]_ , \new_[11603]_ , \new_[11604]_ ,
    \new_[11605]_ , \new_[11606]_ , \new_[11607]_ , \new_[11608]_ ,
    \new_[11609]_ , \new_[11610]_ , \new_[11611]_ , \new_[11612]_ ,
    \new_[11613]_ , \new_[11614]_ , \new_[11615]_ , \new_[11616]_ ,
    \new_[11617]_ , \new_[11618]_ , \new_[11619]_ , \new_[11620]_ ,
    \new_[11621]_ , \new_[11622]_ , \new_[11623]_ , \new_[11624]_ ,
    \new_[11625]_ , \new_[11626]_ , \new_[11627]_ , \new_[11628]_ ,
    \new_[11629]_ , \new_[11630]_ , \new_[11631]_ , \new_[11632]_ ,
    \new_[11633]_ , \new_[11634]_ , \new_[11635]_ , \new_[11636]_ ,
    \new_[11637]_ , \new_[11638]_ , \new_[11639]_ , \new_[11640]_ ,
    \new_[11641]_ , \new_[11642]_ , \new_[11643]_ , \new_[11644]_ ,
    \new_[11645]_ , \new_[11646]_ , \new_[11647]_ , \new_[11648]_ ,
    \new_[11649]_ , \new_[11650]_ , \new_[11651]_ , \new_[11652]_ ,
    \new_[11653]_ , \new_[11654]_ , \new_[11655]_ , \new_[11656]_ ,
    \new_[11657]_ , \new_[11658]_ , \new_[11659]_ , \new_[11660]_ ,
    \new_[11661]_ , \new_[11662]_ , \new_[11663]_ , \new_[11664]_ ,
    \new_[11665]_ , \new_[11666]_ , \new_[11667]_ , \new_[11668]_ ,
    \new_[11669]_ , \new_[11670]_ , \new_[11671]_ , \new_[11672]_ ,
    \new_[11673]_ , \new_[11674]_ , \new_[11675]_ , \new_[11676]_ ,
    \new_[11677]_ , \new_[11678]_ , \new_[11679]_ , \new_[11680]_ ,
    \new_[11681]_ , \new_[11682]_ , \new_[11683]_ , \new_[11684]_ ,
    \new_[11685]_ , \new_[11686]_ , \new_[11687]_ , \new_[11688]_ ,
    \new_[11689]_ , \new_[11690]_ , \new_[11691]_ , \new_[11692]_ ,
    \new_[11693]_ , \new_[11694]_ , \new_[11695]_ , \new_[11696]_ ,
    \new_[11697]_ , \new_[11698]_ , \new_[11699]_ , \new_[11700]_ ,
    \new_[11701]_ , \new_[11702]_ , \new_[11703]_ , \new_[11704]_ ,
    \new_[11705]_ , \new_[11706]_ , \new_[11707]_ , \new_[11708]_ ,
    \new_[11709]_ , \new_[11710]_ , \new_[11711]_ , \new_[11712]_ ,
    \new_[11713]_ , \new_[11714]_ , \new_[11715]_ , \new_[11716]_ ,
    \new_[11717]_ , \new_[11718]_ , \new_[11719]_ , \new_[11720]_ ,
    \new_[11721]_ , \new_[11722]_ , \new_[11723]_ , \new_[11724]_ ,
    \new_[11725]_ , \new_[11726]_ , \new_[11727]_ , \new_[11728]_ ,
    \new_[11729]_ , \new_[11730]_ , \new_[11731]_ , \new_[11732]_ ,
    \new_[11733]_ , \new_[11734]_ , \new_[11735]_ , \new_[11736]_ ,
    \new_[11737]_ , \new_[11738]_ , \new_[11739]_ , \new_[11740]_ ,
    \new_[11741]_ , \new_[11742]_ , \new_[11743]_ , \new_[11744]_ ,
    \new_[11745]_ , \new_[11746]_ , \new_[11747]_ , \new_[11748]_ ,
    \new_[11749]_ , \new_[11750]_ , \new_[11751]_ , \new_[11752]_ ,
    \new_[11753]_ , \new_[11754]_ , \new_[11755]_ , \new_[11756]_ ,
    \new_[11757]_ , \new_[11758]_ , \new_[11759]_ , \new_[11760]_ ,
    \new_[11761]_ , \new_[11762]_ , \new_[11763]_ , \new_[11764]_ ,
    \new_[11765]_ , \new_[11766]_ , \new_[11767]_ , \new_[11768]_ ,
    \new_[11769]_ , \new_[11770]_ , \new_[11771]_ , \new_[11772]_ ,
    \new_[11773]_ , \new_[11774]_ , \new_[11775]_ , \new_[11776]_ ,
    \new_[11777]_ , \new_[11778]_ , \new_[11779]_ , \new_[11780]_ ,
    \new_[11781]_ , \new_[11782]_ , \new_[11783]_ , \new_[11784]_ ,
    \new_[11785]_ , \new_[11786]_ , \new_[11787]_ , \new_[11788]_ ,
    \new_[11789]_ , \new_[11790]_ , \new_[11791]_ , \new_[11792]_ ,
    \new_[11793]_ , \new_[11794]_ , \new_[11795]_ , \new_[11796]_ ,
    \new_[11797]_ , \new_[11798]_ , \new_[11799]_ , \new_[11800]_ ,
    \new_[11801]_ , \new_[11802]_ , \new_[11803]_ , \new_[11804]_ ,
    \new_[11805]_ , \new_[11806]_ , \new_[11807]_ , \new_[11808]_ ,
    \new_[11809]_ , \new_[11810]_ , \new_[11811]_ , \new_[11812]_ ,
    \new_[11813]_ , \new_[11814]_ , \new_[11815]_ , \new_[11816]_ ,
    \new_[11817]_ , \new_[11818]_ , \new_[11819]_ , \new_[11820]_ ,
    \new_[11821]_ , \new_[11822]_ , \new_[11823]_ , \new_[11824]_ ,
    \new_[11825]_ , \new_[11826]_ , \new_[11827]_ , \new_[11828]_ ,
    \new_[11829]_ , \new_[11830]_ , \new_[11831]_ , \new_[11832]_ ,
    \new_[11833]_ , \new_[11834]_ , \new_[11835]_ , \new_[11836]_ ,
    \new_[11837]_ , \new_[11838]_ , \new_[11839]_ , \new_[11840]_ ,
    \new_[11841]_ , \new_[11842]_ , \new_[11843]_ , \new_[11844]_ ,
    \new_[11845]_ , \new_[11846]_ , \new_[11847]_ , \new_[11848]_ ,
    \new_[11849]_ , \new_[11850]_ , \new_[11851]_ , \new_[11852]_ ,
    \new_[11853]_ , \new_[11854]_ , \new_[11855]_ , \new_[11856]_ ,
    \new_[11857]_ , \new_[11858]_ , \new_[11859]_ , \new_[11860]_ ,
    \new_[11861]_ , \new_[11862]_ , \new_[11863]_ , \new_[11864]_ ,
    \new_[11865]_ , \new_[11866]_ , \new_[11867]_ , \new_[11868]_ ,
    \new_[11869]_ , \new_[11870]_ , \new_[11871]_ , \new_[11872]_ ,
    \new_[11873]_ , \new_[11874]_ , \new_[11875]_ , \new_[11876]_ ,
    \new_[11877]_ , \new_[11878]_ , \new_[11879]_ , \new_[11880]_ ,
    \new_[11881]_ , \new_[11882]_ , \new_[11883]_ , \new_[11884]_ ,
    \new_[11885]_ , \new_[11886]_ , \new_[11887]_ , \new_[11888]_ ,
    \new_[11889]_ , \new_[11890]_ , \new_[11891]_ , \new_[11892]_ ,
    \new_[11893]_ , \new_[11894]_ , \new_[11895]_ , \new_[11896]_ ,
    \new_[11897]_ , \new_[11898]_ , \new_[11899]_ , \new_[11900]_ ,
    \new_[11901]_ , \new_[11902]_ , \new_[11903]_ , \new_[11904]_ ,
    \new_[11905]_ , \new_[11906]_ , \new_[11907]_ , \new_[11908]_ ,
    \new_[11909]_ , \new_[11910]_ , \new_[11911]_ , \new_[11912]_ ,
    \new_[11913]_ , \new_[11914]_ , \new_[11915]_ , \new_[11916]_ ,
    \new_[11917]_ , \new_[11918]_ , \new_[11919]_ , \new_[11920]_ ,
    \new_[11921]_ , \new_[11922]_ , \new_[11923]_ , \new_[11924]_ ,
    \new_[11925]_ , \new_[11926]_ , \new_[11927]_ , \new_[11928]_ ,
    \new_[11929]_ , \new_[11930]_ , \new_[11931]_ , \new_[11932]_ ,
    \new_[11933]_ , \new_[11934]_ , \new_[11935]_ , \new_[11936]_ ,
    \new_[11937]_ , \new_[11938]_ , \new_[11939]_ , \new_[11940]_ ,
    \new_[11941]_ , \new_[11942]_ , \new_[11943]_ , \new_[11944]_ ,
    \new_[11945]_ , \new_[11946]_ , \new_[11947]_ , \new_[11948]_ ,
    \new_[11949]_ , \new_[11950]_ , \new_[11951]_ , \new_[11952]_ ,
    \new_[11953]_ , \new_[11954]_ , \new_[11955]_ , \new_[11956]_ ,
    \new_[11957]_ , \new_[11958]_ , \new_[11959]_ , \new_[11960]_ ,
    \new_[11961]_ , \new_[11962]_ , \new_[11963]_ , \new_[11964]_ ,
    \new_[11965]_ , \new_[11966]_ , \new_[11967]_ , \new_[11968]_ ,
    \new_[11969]_ , \new_[11970]_ , \new_[11971]_ , \new_[11972]_ ,
    \new_[11973]_ , \new_[11974]_ , \new_[11975]_ , \new_[11976]_ ,
    \new_[11977]_ , \new_[11978]_ , \new_[11979]_ , \new_[11980]_ ,
    \new_[11981]_ , \new_[11982]_ , \new_[11983]_ , \new_[11984]_ ,
    \new_[11985]_ , \new_[11986]_ , \new_[11987]_ , \new_[11988]_ ,
    \new_[11989]_ , \new_[11990]_ , \new_[11991]_ , \new_[11992]_ ,
    \new_[11993]_ , \new_[11994]_ , \new_[11995]_ , \new_[11996]_ ,
    \new_[11997]_ , \new_[11998]_ , \new_[11999]_ , \new_[12000]_ ,
    \new_[12001]_ , \new_[12002]_ , \new_[12005]_ , \new_[12006]_ ,
    \new_[12009]_ , \new_[12010]_ , \new_[12011]_ , \new_[12012]_ ,
    \new_[12013]_ , \new_[12014]_ , \new_[12015]_ , \new_[12016]_ ,
    \new_[12017]_ , \new_[12018]_ , \new_[12019]_ , \new_[12020]_ ,
    \new_[12021]_ , \new_[12022]_ , \new_[12023]_ , \new_[12024]_ ,
    \new_[12025]_ , \new_[12026]_ , \new_[12027]_ , \new_[12028]_ ,
    \new_[12029]_ , \new_[12030]_ , \new_[12031]_ , \new_[12032]_ ,
    \new_[12033]_ , \new_[12034]_ , \new_[12035]_ , \new_[12036]_ ,
    \new_[12037]_ , \new_[12038]_ , \new_[12039]_ , \new_[12040]_ ,
    \new_[12041]_ , \new_[12042]_ , \new_[12043]_ , \new_[12044]_ ,
    \new_[12045]_ , \new_[12046]_ , \new_[12047]_ , \new_[12048]_ ,
    \new_[12049]_ , \new_[12050]_ , \new_[12051]_ , \new_[12052]_ ,
    \new_[12053]_ , \new_[12054]_ , \new_[12055]_ , \new_[12056]_ ,
    \new_[12057]_ , \new_[12058]_ , \new_[12059]_ , \new_[12060]_ ,
    \new_[12061]_ , \new_[12062]_ , \new_[12063]_ , \new_[12064]_ ,
    \new_[12065]_ , \new_[12066]_ , \new_[12067]_ , \new_[12068]_ ,
    \new_[12069]_ , \new_[12070]_ , \new_[12071]_ , \new_[12072]_ ,
    \new_[12073]_ , \new_[12074]_ , \new_[12075]_ , \new_[12076]_ ,
    \new_[12077]_ , \new_[12078]_ , \new_[12079]_ , \new_[12080]_ ,
    \new_[12081]_ , \new_[12082]_ , \new_[12083]_ , \new_[12084]_ ,
    \new_[12085]_ , \new_[12086]_ , \new_[12087]_ , \new_[12088]_ ,
    \new_[12089]_ , \new_[12090]_ , \new_[12091]_ , \new_[12092]_ ,
    \new_[12093]_ , \new_[12094]_ , \new_[12095]_ , \new_[12096]_ ,
    \new_[12097]_ , \new_[12098]_ , \new_[12100]_ , \new_[12101]_ ,
    \new_[12102]_ , \new_[12103]_ , \new_[12104]_ , \new_[12105]_ ,
    \new_[12106]_ , \new_[12107]_ , \new_[12108]_ , \new_[12109]_ ,
    \new_[12110]_ , \new_[12111]_ , \new_[12112]_ , \new_[12113]_ ,
    \new_[12115]_ , \new_[12116]_ , \new_[12117]_ , \new_[12118]_ ,
    \new_[12119]_ , \new_[12120]_ , \new_[12121]_ , \new_[12122]_ ,
    \new_[12123]_ , \new_[12124]_ , \new_[12125]_ , \new_[12126]_ ,
    \new_[12127]_ , \new_[12128]_ , \new_[12129]_ , \new_[12130]_ ,
    \new_[12131]_ , \new_[12132]_ , \new_[12133]_ , \new_[12134]_ ,
    \new_[12135]_ , \new_[12136]_ , \new_[12137]_ , \new_[12138]_ ,
    \new_[12139]_ , \new_[12140]_ , \new_[12141]_ , \new_[12142]_ ,
    \new_[12143]_ , \new_[12144]_ , \new_[12145]_ , \new_[12146]_ ,
    \new_[12147]_ , \new_[12148]_ , \new_[12149]_ , \new_[12150]_ ,
    \new_[12151]_ , \new_[12152]_ , \new_[12153]_ , \new_[12154]_ ,
    \new_[12155]_ , \new_[12156]_ , \new_[12157]_ , \new_[12158]_ ,
    \new_[12159]_ , \new_[12160]_ , \new_[12161]_ , \new_[12162]_ ,
    \new_[12163]_ , \new_[12164]_ , \new_[12165]_ , \new_[12166]_ ,
    \new_[12167]_ , \new_[12168]_ , \new_[12169]_ , \new_[12170]_ ,
    \new_[12171]_ , \new_[12172]_ , \new_[12173]_ , \new_[12174]_ ,
    \new_[12175]_ , \new_[12176]_ , \new_[12177]_ , \new_[12178]_ ,
    \new_[12179]_ , \new_[12180]_ , \new_[12181]_ , \new_[12182]_ ,
    \new_[12183]_ , \new_[12184]_ , \new_[12185]_ , \new_[12186]_ ,
    \new_[12187]_ , \new_[12188]_ , \new_[12189]_ , \new_[12190]_ ,
    \new_[12191]_ , \new_[12192]_ , \new_[12193]_ , \new_[12194]_ ,
    \new_[12195]_ , \new_[12196]_ , \new_[12197]_ , \new_[12198]_ ,
    \new_[12199]_ , \new_[12200]_ , \new_[12201]_ , \new_[12202]_ ,
    \new_[12203]_ , \new_[12204]_ , \new_[12205]_ , \new_[12206]_ ,
    \new_[12207]_ , \new_[12208]_ , \new_[12209]_ , \new_[12210]_ ,
    \new_[12211]_ , \new_[12212]_ , \new_[12213]_ , \new_[12214]_ ,
    \new_[12215]_ , \new_[12216]_ , \new_[12217]_ , \new_[12218]_ ,
    \new_[12219]_ , \new_[12220]_ , \new_[12221]_ , \new_[12222]_ ,
    \new_[12223]_ , \new_[12224]_ , \new_[12225]_ , \new_[12226]_ ,
    \new_[12227]_ , \new_[12228]_ , \new_[12229]_ , \new_[12230]_ ,
    \new_[12231]_ , \new_[12232]_ , \new_[12233]_ , \new_[12234]_ ,
    \new_[12235]_ , \new_[12236]_ , \new_[12237]_ , \new_[12238]_ ,
    \new_[12239]_ , \new_[12240]_ , \new_[12241]_ , \new_[12242]_ ,
    \new_[12243]_ , \new_[12244]_ , \new_[12245]_ , \new_[12246]_ ,
    \new_[12247]_ , \new_[12248]_ , \new_[12249]_ , \new_[12250]_ ,
    \new_[12251]_ , \new_[12252]_ , \new_[12253]_ , \new_[12254]_ ,
    \new_[12255]_ , \new_[12256]_ , \new_[12257]_ , \new_[12258]_ ,
    \new_[12259]_ , \new_[12260]_ , \new_[12261]_ , \new_[12262]_ ,
    \new_[12263]_ , \new_[12264]_ , \new_[12265]_ , \new_[12266]_ ,
    \new_[12267]_ , \new_[12268]_ , \new_[12269]_ , \new_[12270]_ ,
    \new_[12271]_ , \new_[12272]_ , \new_[12273]_ , \new_[12274]_ ,
    \new_[12275]_ , \new_[12276]_ , \new_[12277]_ , \new_[12278]_ ,
    \new_[12279]_ , \new_[12280]_ , \new_[12281]_ , \new_[12282]_ ,
    \new_[12283]_ , \new_[12284]_ , \new_[12285]_ , \new_[12286]_ ,
    \new_[12287]_ , \new_[12288]_ , \new_[12289]_ , \new_[12290]_ ,
    \new_[12291]_ , \new_[12292]_ , \new_[12293]_ , \new_[12294]_ ,
    \new_[12295]_ , \new_[12296]_ , \new_[12297]_ , \new_[12298]_ ,
    \new_[12299]_ , \new_[12300]_ , \new_[12301]_ , \new_[12302]_ ,
    \new_[12303]_ , \new_[12304]_ , \new_[12305]_ , \new_[12306]_ ,
    \new_[12307]_ , \new_[12308]_ , \new_[12309]_ , \new_[12310]_ ,
    \new_[12311]_ , \new_[12312]_ , \new_[12313]_ , \new_[12314]_ ,
    \new_[12315]_ , \new_[12316]_ , \new_[12317]_ , \new_[12318]_ ,
    \new_[12319]_ , \new_[12320]_ , \new_[12321]_ , \new_[12322]_ ,
    \new_[12323]_ , \new_[12324]_ , \new_[12325]_ , \new_[12326]_ ,
    \new_[12327]_ , \new_[12328]_ , \new_[12329]_ , \new_[12330]_ ,
    \new_[12331]_ , \new_[12332]_ , \new_[12333]_ , \new_[12334]_ ,
    \new_[12335]_ , \new_[12336]_ , \new_[12337]_ , \new_[12338]_ ,
    \new_[12339]_ , \new_[12340]_ , \new_[12341]_ , \new_[12342]_ ,
    \new_[12343]_ , \new_[12344]_ , \new_[12345]_ , \new_[12346]_ ,
    \new_[12347]_ , \new_[12348]_ , \new_[12349]_ , \new_[12350]_ ,
    \new_[12351]_ , \new_[12352]_ , \new_[12353]_ , \new_[12354]_ ,
    \new_[12355]_ , \new_[12356]_ , \new_[12357]_ , \new_[12358]_ ,
    \new_[12359]_ , \new_[12360]_ , \new_[12361]_ , \new_[12362]_ ,
    \new_[12363]_ , \new_[12364]_ , \new_[12365]_ , \new_[12366]_ ,
    \new_[12367]_ , \new_[12368]_ , \new_[12369]_ , \new_[12370]_ ,
    \new_[12371]_ , \new_[12372]_ , \new_[12373]_ , \new_[12374]_ ,
    \new_[12375]_ , \new_[12376]_ , \new_[12377]_ , \new_[12378]_ ,
    \new_[12379]_ , \new_[12380]_ , \new_[12381]_ , \new_[12382]_ ,
    \new_[12383]_ , \new_[12384]_ , \new_[12385]_ , \new_[12386]_ ,
    \new_[12387]_ , \new_[12388]_ , \new_[12389]_ , \new_[12390]_ ,
    \new_[12391]_ , \new_[12392]_ , \new_[12393]_ , \new_[12394]_ ,
    \new_[12395]_ , \new_[12396]_ , \new_[12397]_ , \new_[12398]_ ,
    \new_[12399]_ , \new_[12400]_ , \new_[12401]_ , \new_[12402]_ ,
    \new_[12403]_ , \new_[12404]_ , \new_[12405]_ , \new_[12406]_ ,
    \new_[12407]_ , \new_[12408]_ , \new_[12409]_ , \new_[12410]_ ,
    \new_[12411]_ , \new_[12412]_ , \new_[12413]_ , \new_[12414]_ ,
    \new_[12415]_ , \new_[12416]_ , \new_[12417]_ , \new_[12418]_ ,
    \new_[12419]_ , \new_[12420]_ , \new_[12421]_ , \new_[12422]_ ,
    \new_[12423]_ , \new_[12424]_ , \new_[12425]_ , \new_[12426]_ ,
    \new_[12427]_ , \new_[12428]_ , \new_[12429]_ , \new_[12430]_ ,
    \new_[12431]_ , \new_[12432]_ , \new_[12433]_ , \new_[12434]_ ,
    \new_[12435]_ , \new_[12436]_ , \new_[12437]_ , \new_[12438]_ ,
    \new_[12439]_ , \new_[12440]_ , \new_[12441]_ , \new_[12442]_ ,
    \new_[12443]_ , \new_[12444]_ , \new_[12445]_ , \new_[12446]_ ,
    \new_[12447]_ , \new_[12448]_ , \new_[12449]_ , \new_[12450]_ ,
    \new_[12451]_ , \new_[12452]_ , \new_[12453]_ , \new_[12454]_ ,
    \new_[12455]_ , \new_[12456]_ , \new_[12457]_ , \new_[12458]_ ,
    \new_[12459]_ , \new_[12460]_ , \new_[12461]_ , \new_[12462]_ ,
    \new_[12463]_ , \new_[12464]_ , \new_[12465]_ , \new_[12466]_ ,
    \new_[12467]_ , \new_[12468]_ , \new_[12469]_ , \new_[12470]_ ,
    \new_[12471]_ , \new_[12472]_ , \new_[12473]_ , \new_[12474]_ ,
    \new_[12475]_ , \new_[12476]_ , \new_[12477]_ , \new_[12478]_ ,
    \new_[12479]_ , \new_[12480]_ , \new_[12481]_ , \new_[12482]_ ,
    \new_[12483]_ , \new_[12484]_ , \new_[12485]_ , \new_[12486]_ ,
    \new_[12487]_ , \new_[12488]_ , \new_[12489]_ , \new_[12490]_ ,
    \new_[12491]_ , \new_[12492]_ , \new_[12493]_ , \new_[12494]_ ,
    \new_[12495]_ , \new_[12496]_ , \new_[12497]_ , \new_[12498]_ ,
    \new_[12499]_ , \new_[12500]_ , \new_[12501]_ , \new_[12502]_ ,
    \new_[12503]_ , \new_[12504]_ , \new_[12505]_ , \new_[12506]_ ,
    \new_[12507]_ , \new_[12508]_ , \new_[12509]_ , \new_[12510]_ ,
    \new_[12511]_ , \new_[12512]_ , \new_[12513]_ , \new_[12514]_ ,
    \new_[12515]_ , \new_[12516]_ , \new_[12517]_ , \new_[12518]_ ,
    \new_[12519]_ , \new_[12520]_ , \new_[12521]_ , \new_[12522]_ ,
    \new_[12523]_ , \new_[12524]_ , \new_[12525]_ , \new_[12526]_ ,
    \new_[12527]_ , \new_[12528]_ , \new_[12529]_ , \new_[12530]_ ,
    \new_[12531]_ , \new_[12533]_ , \new_[12534]_ , \new_[12535]_ ,
    \new_[12543]_ , \new_[12544]_ , \new_[12545]_ , \new_[12546]_ ,
    \new_[12547]_ , \new_[12548]_ , \new_[12549]_ , \new_[12550]_ ,
    \new_[12551]_ , \new_[12552]_ , \new_[12553]_ , \new_[12554]_ ,
    \new_[12555]_ , \new_[12556]_ , \new_[12557]_ , \new_[12558]_ ,
    \new_[12559]_ , \new_[12560]_ , \new_[12561]_ , \new_[12562]_ ,
    \new_[12563]_ , \new_[12564]_ , \new_[12565]_ , \new_[12566]_ ,
    \new_[12567]_ , \new_[12568]_ , \new_[12569]_ , \new_[12570]_ ,
    \new_[12571]_ , \new_[12572]_ , \new_[12573]_ , \new_[12574]_ ,
    \new_[12575]_ , \new_[12576]_ , \new_[12577]_ , \new_[12578]_ ,
    \new_[12579]_ , \new_[12580]_ , \new_[12581]_ , \new_[12582]_ ,
    \new_[12583]_ , \new_[12584]_ , \new_[12585]_ , \new_[12586]_ ,
    \new_[12587]_ , \new_[12588]_ , \new_[12589]_ , \new_[12590]_ ,
    \new_[12591]_ , \new_[12592]_ , \new_[12593]_ , \new_[12594]_ ,
    \new_[12595]_ , \new_[12596]_ , \new_[12597]_ , \new_[12598]_ ,
    \new_[12599]_ , \new_[12600]_ , \new_[12601]_ , \new_[12602]_ ,
    \new_[12603]_ , \new_[12604]_ , \new_[12605]_ , \new_[12606]_ ,
    \new_[12607]_ , \new_[12608]_ , \new_[12609]_ , \new_[12610]_ ,
    \new_[12611]_ , \new_[12612]_ , \new_[12613]_ , \new_[12614]_ ,
    \new_[12615]_ , \new_[12616]_ , \new_[12617]_ , \new_[12618]_ ,
    \new_[12619]_ , \new_[12620]_ , \new_[12621]_ , \new_[12622]_ ,
    \new_[12623]_ , \new_[12624]_ , \new_[12625]_ , \new_[12626]_ ,
    \new_[12627]_ , \new_[12628]_ , \new_[12629]_ , \new_[12630]_ ,
    \new_[12631]_ , \new_[12632]_ , \new_[12633]_ , \new_[12635]_ ,
    \new_[12636]_ , \new_[12637]_ , \new_[12638]_ , \new_[12639]_ ,
    \new_[12640]_ , \new_[12641]_ , \new_[12642]_ , \new_[12643]_ ,
    \new_[12644]_ , \new_[12645]_ , \new_[12647]_ , \new_[12648]_ ,
    \new_[12649]_ , \new_[12650]_ , \new_[12651]_ , \new_[12652]_ ,
    \new_[12653]_ , \new_[12654]_ , \new_[12655]_ , \new_[12656]_ ,
    \new_[12657]_ , \new_[12658]_ , \new_[12659]_ , \new_[12660]_ ,
    \new_[12662]_ , \new_[12663]_ , \new_[12664]_ , \new_[12665]_ ,
    \new_[12666]_ , \new_[12667]_ , \new_[12670]_ , \new_[12671]_ ,
    \new_[12672]_ , \new_[12676]_ , \new_[12678]_ , \new_[12679]_ ,
    \new_[12680]_ , \new_[12681]_ , \new_[12682]_ , \new_[12684]_ ,
    \new_[12685]_ , \new_[12686]_ , \new_[12687]_ , \new_[12688]_ ,
    \new_[12689]_ , \new_[12690]_ , \new_[12691]_ , \new_[12692]_ ,
    \new_[12693]_ , \new_[12694]_ , \new_[12696]_ , \new_[12697]_ ,
    \new_[12698]_ , \new_[12699]_ , \new_[12700]_ , \new_[12701]_ ,
    \new_[12702]_ , \new_[12703]_ , \new_[12704]_ , \new_[12705]_ ,
    \new_[12706]_ , \new_[12707]_ , \new_[12708]_ , \new_[12709]_ ,
    \new_[12710]_ , \new_[12711]_ , \new_[12712]_ , \new_[12713]_ ,
    \new_[12714]_ , \new_[12715]_ , \new_[12716]_ , \new_[12717]_ ,
    \new_[12718]_ , \new_[12719]_ , \new_[12720]_ , \new_[12721]_ ,
    \new_[12722]_ , \new_[12723]_ , \new_[12724]_ , \new_[12725]_ ,
    \new_[12726]_ , \new_[12727]_ , \new_[12728]_ , \new_[12729]_ ,
    \new_[12730]_ , \new_[12731]_ , \new_[12732]_ , \new_[12733]_ ,
    \new_[12734]_ , \new_[12735]_ , \new_[12736]_ , \new_[12737]_ ,
    \new_[12738]_ , \new_[12739]_ , \new_[12740]_ , \new_[12741]_ ,
    \new_[12742]_ , \new_[12743]_ , \new_[12744]_ , \new_[12745]_ ,
    \new_[12746]_ , \new_[12747]_ , \new_[12748]_ , \new_[12749]_ ,
    \new_[12750]_ , \new_[12751]_ , \new_[12752]_ , \new_[12753]_ ,
    \new_[12754]_ , \new_[12755]_ , \new_[12756]_ , \new_[12757]_ ,
    \new_[12758]_ , \new_[12759]_ , \new_[12760]_ , \new_[12761]_ ,
    \new_[12762]_ , \new_[12763]_ , \new_[12764]_ , \new_[12765]_ ,
    \new_[12766]_ , \new_[12767]_ , \new_[12768]_ , \new_[12769]_ ,
    \new_[12770]_ , \new_[12771]_ , \new_[12772]_ , \new_[12773]_ ,
    \new_[12774]_ , \new_[12775]_ , \new_[12776]_ , \new_[12777]_ ,
    \new_[12778]_ , \new_[12779]_ , \new_[12780]_ , \new_[12781]_ ,
    \new_[12782]_ , \new_[12783]_ , \new_[12784]_ , \new_[12785]_ ,
    \new_[12786]_ , \new_[12787]_ , \new_[12788]_ , \new_[12789]_ ,
    \new_[12790]_ , \new_[12791]_ , \new_[12792]_ , \new_[12793]_ ,
    \new_[12794]_ , \new_[12795]_ , \new_[12796]_ , \new_[12797]_ ,
    \new_[12798]_ , \new_[12799]_ , \new_[12800]_ , \new_[12801]_ ,
    \new_[12803]_ , \new_[12804]_ , \new_[12805]_ , \new_[12806]_ ,
    \new_[12807]_ , \new_[12808]_ , \new_[12809]_ , \new_[12810]_ ,
    \new_[12811]_ , \new_[12812]_ , \new_[12813]_ , \new_[12814]_ ,
    \new_[12815]_ , \new_[12816]_ , \new_[12817]_ , \new_[12818]_ ,
    \new_[12819]_ , \new_[12820]_ , \new_[12821]_ , \new_[12822]_ ,
    \new_[12823]_ , \new_[12824]_ , \new_[12825]_ , \new_[12826]_ ,
    \new_[12827]_ , \new_[12828]_ , \new_[12829]_ , \new_[12830]_ ,
    \new_[12831]_ , \new_[12832]_ , \new_[12833]_ , \new_[12834]_ ,
    \new_[12835]_ , \new_[12836]_ , \new_[12837]_ , \new_[12838]_ ,
    \new_[12839]_ , \new_[12840]_ , \new_[12841]_ , \new_[12842]_ ,
    \new_[12843]_ , \new_[12844]_ , \new_[12845]_ , \new_[12846]_ ,
    \new_[12847]_ , \new_[12848]_ , \new_[12849]_ , \new_[12850]_ ,
    \new_[12851]_ , \new_[12852]_ , \new_[12853]_ , \new_[12854]_ ,
    \new_[12855]_ , \new_[12856]_ , \new_[12857]_ , \new_[12858]_ ,
    \new_[12859]_ , \new_[12860]_ , \new_[12861]_ , \new_[12862]_ ,
    \new_[12863]_ , \new_[12864]_ , \new_[12865]_ , \new_[12866]_ ,
    \new_[12867]_ , \new_[12868]_ , \new_[12869]_ , \new_[12870]_ ,
    \new_[12871]_ , \new_[12872]_ , \new_[12873]_ , \new_[12874]_ ,
    \new_[12875]_ , \new_[12876]_ , \new_[12877]_ , \new_[12878]_ ,
    \new_[12879]_ , \new_[12880]_ , \new_[12881]_ , \new_[12882]_ ,
    \new_[12883]_ , \new_[12884]_ , \new_[12885]_ , \new_[12886]_ ,
    \new_[12887]_ , \new_[12888]_ , \new_[12889]_ , \new_[12890]_ ,
    \new_[12891]_ , \new_[12892]_ , \new_[12893]_ , \new_[12894]_ ,
    \new_[12895]_ , \new_[12896]_ , \new_[12897]_ , \new_[12898]_ ,
    \new_[12899]_ , \new_[12900]_ , \new_[12901]_ , \new_[12902]_ ,
    \new_[12903]_ , \new_[12904]_ , \new_[12905]_ , \new_[12906]_ ,
    \new_[12907]_ , \new_[12908]_ , \new_[12909]_ , \new_[12910]_ ,
    \new_[12911]_ , \new_[12912]_ , \new_[12913]_ , \new_[12914]_ ,
    \new_[12915]_ , \new_[12916]_ , \new_[12917]_ , \new_[12918]_ ,
    \new_[12919]_ , \new_[12920]_ , \new_[12921]_ , \new_[12922]_ ,
    \new_[12923]_ , \new_[12924]_ , \new_[12925]_ , \new_[12926]_ ,
    \new_[12927]_ , \new_[12928]_ , \new_[12929]_ , \new_[12930]_ ,
    \new_[12931]_ , \new_[12932]_ , \new_[12933]_ , \new_[12934]_ ,
    \new_[12935]_ , \new_[12936]_ , \new_[12937]_ , \new_[12938]_ ,
    \new_[12939]_ , \new_[12941]_ , \new_[12942]_ , \new_[12943]_ ,
    \new_[12944]_ , \new_[12945]_ , \new_[12946]_ , \new_[12947]_ ,
    \new_[12948]_ , \new_[12949]_ , \new_[12950]_ , \new_[12951]_ ,
    \new_[12952]_ , \new_[12953]_ , \new_[12954]_ , \new_[12955]_ ,
    \new_[12956]_ , \new_[12957]_ , \new_[12958]_ , \new_[12959]_ ,
    \new_[12960]_ , \new_[12961]_ , \new_[12962]_ , \new_[12963]_ ,
    \new_[12964]_ , \new_[12965]_ , \new_[12966]_ , \new_[12967]_ ,
    \new_[12968]_ , \new_[12969]_ , \new_[12970]_ , \new_[12971]_ ,
    \new_[12972]_ , \new_[12973]_ , \new_[12974]_ , \new_[12975]_ ,
    \new_[12976]_ , \new_[12977]_ , \new_[12978]_ , \new_[12979]_ ,
    \new_[12980]_ , \new_[12981]_ , \new_[12982]_ , \new_[12983]_ ,
    \new_[12984]_ , \new_[12985]_ , \new_[12986]_ , \new_[12987]_ ,
    \new_[12988]_ , \new_[12989]_ , \new_[12990]_ , \new_[12991]_ ,
    \new_[12992]_ , \new_[12993]_ , \new_[12994]_ , \new_[12995]_ ,
    \new_[12996]_ , \new_[12997]_ , \new_[12998]_ , \new_[12999]_ ,
    \new_[13000]_ , \new_[13001]_ , \new_[13002]_ , \new_[13003]_ ,
    \new_[13004]_ , \new_[13005]_ , \new_[13006]_ , \new_[13007]_ ,
    \new_[13008]_ , \new_[13009]_ , \new_[13010]_ , \new_[13011]_ ,
    \new_[13012]_ , \new_[13013]_ , \new_[13014]_ , \new_[13015]_ ,
    \new_[13016]_ , \new_[13017]_ , \new_[13018]_ , \new_[13019]_ ,
    \new_[13020]_ , \new_[13021]_ , \new_[13022]_ , \new_[13023]_ ,
    \new_[13024]_ , \new_[13025]_ , \new_[13026]_ , \new_[13027]_ ,
    \new_[13028]_ , \new_[13029]_ , \new_[13030]_ , \new_[13031]_ ,
    \new_[13032]_ , \new_[13033]_ , \new_[13034]_ , \new_[13035]_ ,
    \new_[13036]_ , \new_[13037]_ , \new_[13038]_ , \new_[13039]_ ,
    \new_[13040]_ , \new_[13041]_ , \new_[13042]_ , \new_[13043]_ ,
    \new_[13044]_ , \new_[13045]_ , \new_[13046]_ , \new_[13047]_ ,
    \new_[13048]_ , \new_[13049]_ , \new_[13050]_ , \new_[13051]_ ,
    \new_[13052]_ , \new_[13053]_ , \new_[13054]_ , \new_[13055]_ ,
    \new_[13056]_ , \new_[13057]_ , \new_[13058]_ , \new_[13059]_ ,
    \new_[13060]_ , \new_[13061]_ , \new_[13063]_ , \new_[13064]_ ,
    \new_[13065]_ , \new_[13066]_ , \new_[13067]_ , \new_[13068]_ ,
    \new_[13069]_ , \new_[13070]_ , \new_[13071]_ , \new_[13072]_ ,
    \new_[13073]_ , \new_[13074]_ , \new_[13075]_ , \new_[13076]_ ,
    \new_[13077]_ , \new_[13078]_ , \new_[13079]_ , \new_[13080]_ ,
    \new_[13081]_ , \new_[13082]_ , \new_[13083]_ , \new_[13084]_ ,
    \new_[13085]_ , \new_[13086]_ , \new_[13087]_ , \new_[13088]_ ,
    \new_[13089]_ , \new_[13090]_ , \new_[13091]_ , \new_[13092]_ ,
    \new_[13093]_ , \new_[13094]_ , \new_[13095]_ , \new_[13096]_ ,
    \new_[13097]_ , \new_[13098]_ , \new_[13099]_ , \new_[13100]_ ,
    \new_[13101]_ , \new_[13102]_ , \new_[13103]_ , \new_[13104]_ ,
    \new_[13105]_ , \new_[13106]_ , \new_[13107]_ , \new_[13108]_ ,
    \new_[13109]_ , \new_[13110]_ , \new_[13111]_ , \new_[13112]_ ,
    \new_[13113]_ , \new_[13114]_ , \new_[13115]_ , \new_[13116]_ ,
    \new_[13117]_ , \new_[13118]_ , \new_[13119]_ , \new_[13120]_ ,
    \new_[13121]_ , \new_[13122]_ , \new_[13123]_ , \new_[13124]_ ,
    \new_[13125]_ , \new_[13126]_ , \new_[13127]_ , \new_[13128]_ ,
    \new_[13129]_ , \new_[13130]_ , \new_[13131]_ , \new_[13132]_ ,
    \new_[13133]_ , \new_[13134]_ , \new_[13135]_ , \new_[13136]_ ,
    \new_[13137]_ , \new_[13138]_ , \new_[13139]_ , \new_[13140]_ ,
    \new_[13141]_ , \new_[13142]_ , \new_[13143]_ , \new_[13144]_ ,
    \new_[13145]_ , \new_[13146]_ , \new_[13147]_ , \new_[13148]_ ,
    \new_[13149]_ , \new_[13150]_ , \new_[13151]_ , \new_[13152]_ ,
    \new_[13153]_ , \new_[13154]_ , \new_[13155]_ , \new_[13156]_ ,
    \new_[13157]_ , \new_[13158]_ , \new_[13159]_ , \new_[13160]_ ,
    \new_[13161]_ , \new_[13162]_ , \new_[13163]_ , \new_[13164]_ ,
    \new_[13165]_ , \new_[13166]_ , \new_[13167]_ , \new_[13168]_ ,
    \new_[13169]_ , \new_[13170]_ , \new_[13171]_ , \new_[13172]_ ,
    \new_[13173]_ , \new_[13174]_ , \new_[13175]_ , \new_[13176]_ ,
    \new_[13177]_ , \new_[13178]_ , \new_[13179]_ , \new_[13180]_ ,
    \new_[13181]_ , \new_[13182]_ , \new_[13183]_ , \new_[13184]_ ,
    \new_[13185]_ , \new_[13186]_ , \new_[13187]_ , \new_[13188]_ ,
    \new_[13189]_ , \new_[13190]_ , \new_[13191]_ , \new_[13192]_ ,
    \new_[13193]_ , \new_[13194]_ , \new_[13195]_ , \new_[13196]_ ,
    \new_[13197]_ , \new_[13198]_ , \new_[13199]_ , \new_[13200]_ ,
    \new_[13201]_ , \new_[13202]_ , \new_[13203]_ , \new_[13204]_ ,
    \new_[13205]_ , \new_[13206]_ , \new_[13207]_ , \new_[13208]_ ,
    \new_[13209]_ , \new_[13210]_ , \new_[13211]_ , \new_[13212]_ ,
    \new_[13213]_ , \new_[13214]_ , \new_[13215]_ , \new_[13216]_ ,
    \new_[13217]_ , \new_[13218]_ , \new_[13219]_ , \new_[13220]_ ,
    \new_[13221]_ , \new_[13222]_ , \new_[13223]_ , \new_[13224]_ ,
    \new_[13225]_ , \new_[13226]_ , \new_[13227]_ , \new_[13228]_ ,
    \new_[13229]_ , \new_[13230]_ , \new_[13231]_ , \new_[13232]_ ,
    \new_[13233]_ , \new_[13234]_ , \new_[13235]_ , \new_[13236]_ ,
    \new_[13237]_ , \new_[13238]_ , \new_[13239]_ , \new_[13240]_ ,
    \new_[13241]_ , \new_[13242]_ , \new_[13243]_ , \new_[13244]_ ,
    \new_[13245]_ , \new_[13246]_ , \new_[13247]_ , \new_[13248]_ ,
    \new_[13249]_ , \new_[13250]_ , \new_[13251]_ , \new_[13252]_ ,
    \new_[13253]_ , \new_[13254]_ , \new_[13255]_ , \new_[13256]_ ,
    \new_[13257]_ , \new_[13258]_ , \new_[13259]_ , \new_[13260]_ ,
    \new_[13261]_ , \new_[13262]_ , \new_[13263]_ , \new_[13264]_ ,
    \new_[13265]_ , \new_[13266]_ , \new_[13267]_ , \new_[13268]_ ,
    \new_[13269]_ , \new_[13270]_ , \new_[13271]_ , \new_[13272]_ ,
    \new_[13273]_ , \new_[13274]_ , \new_[13275]_ , \new_[13276]_ ,
    \new_[13277]_ , \new_[13278]_ , \new_[13279]_ , \new_[13280]_ ,
    \new_[13281]_ , \new_[13282]_ , \new_[13283]_ , \new_[13284]_ ,
    \new_[13285]_ , \new_[13286]_ , \new_[13287]_ , \new_[13288]_ ,
    \new_[13289]_ , \new_[13290]_ , \new_[13291]_ , \new_[13292]_ ,
    \new_[13293]_ , \new_[13294]_ , \new_[13295]_ , \new_[13296]_ ,
    \new_[13297]_ , \new_[13298]_ , \new_[13299]_ , \new_[13300]_ ,
    \new_[13301]_ , \new_[13302]_ , \new_[13303]_ , \new_[13304]_ ,
    \new_[13305]_ , \new_[13306]_ , \new_[13307]_ , \new_[13308]_ ,
    \new_[13309]_ , \new_[13310]_ , \new_[13311]_ , \new_[13312]_ ,
    \new_[13313]_ , \new_[13314]_ , \new_[13315]_ , \new_[13316]_ ,
    \new_[13317]_ , \new_[13318]_ , \new_[13319]_ , \new_[13320]_ ,
    \new_[13321]_ , \new_[13322]_ , \new_[13323]_ , \new_[13324]_ ,
    \new_[13325]_ , \new_[13326]_ , \new_[13327]_ , \new_[13328]_ ,
    \new_[13329]_ , \new_[13330]_ , \new_[13331]_ , \new_[13332]_ ,
    \new_[13333]_ , \new_[13334]_ , \new_[13335]_ , \new_[13336]_ ,
    \new_[13337]_ , \new_[13338]_ , \new_[13339]_ , \new_[13340]_ ,
    \new_[13341]_ , \new_[13342]_ , \new_[13343]_ , \new_[13344]_ ,
    \new_[13345]_ , \new_[13346]_ , \new_[13347]_ , \new_[13348]_ ,
    \new_[13349]_ , \new_[13350]_ , \new_[13351]_ , \new_[13352]_ ,
    \new_[13353]_ , \new_[13354]_ , \new_[13355]_ , \new_[13356]_ ,
    \new_[13357]_ , \new_[13358]_ , \new_[13359]_ , \new_[13360]_ ,
    \new_[13361]_ , \new_[13362]_ , \new_[13363]_ , \new_[13364]_ ,
    \new_[13365]_ , \new_[13366]_ , \new_[13367]_ , \new_[13368]_ ,
    \new_[13369]_ , \new_[13370]_ , \new_[13371]_ , \new_[13372]_ ,
    \new_[13373]_ , \new_[13374]_ , \new_[13375]_ , \new_[13376]_ ,
    \new_[13377]_ , \new_[13378]_ , \new_[13379]_ , \new_[13380]_ ,
    \new_[13381]_ , \new_[13382]_ , \new_[13383]_ , \new_[13384]_ ,
    \new_[13385]_ , \new_[13386]_ , \new_[13387]_ , \new_[13388]_ ,
    \new_[13389]_ , \new_[13390]_ , \new_[13391]_ , \new_[13392]_ ,
    \new_[13393]_ , \new_[13394]_ , \new_[13395]_ , \new_[13396]_ ,
    \new_[13397]_ , \new_[13398]_ , \new_[13399]_ , \new_[13400]_ ,
    \new_[13401]_ , \new_[13402]_ , \new_[13403]_ , \new_[13404]_ ,
    \new_[13405]_ , \new_[13406]_ , \new_[13407]_ , \new_[13408]_ ,
    \new_[13409]_ , \new_[13410]_ , \new_[13411]_ , \new_[13412]_ ,
    \new_[13413]_ , \new_[13414]_ , \new_[13415]_ , \new_[13416]_ ,
    \new_[13417]_ , \new_[13418]_ , \new_[13419]_ , \new_[13420]_ ,
    \new_[13421]_ , \new_[13422]_ , \new_[13423]_ , \new_[13424]_ ,
    \new_[13425]_ , \new_[13426]_ , \new_[13427]_ , \new_[13428]_ ,
    \new_[13429]_ , \new_[13430]_ , \new_[13431]_ , \new_[13432]_ ,
    \new_[13433]_ , \new_[13434]_ , \new_[13435]_ , \new_[13436]_ ,
    \new_[13437]_ , \new_[13438]_ , \new_[13439]_ , \new_[13440]_ ,
    \new_[13441]_ , \new_[13442]_ , \new_[13443]_ , \new_[13444]_ ,
    \new_[13445]_ , \new_[13446]_ , \new_[13447]_ , \new_[13448]_ ,
    \new_[13449]_ , \new_[13450]_ , \new_[13451]_ , \new_[13452]_ ,
    \new_[13453]_ , \new_[13454]_ , \new_[13455]_ , \new_[13456]_ ,
    \new_[13457]_ , \new_[13458]_ , \new_[13459]_ , \new_[13460]_ ,
    \new_[13461]_ , \new_[13462]_ , \new_[13463]_ , \new_[13464]_ ,
    \new_[13465]_ , \new_[13466]_ , \new_[13467]_ , \new_[13468]_ ,
    \new_[13469]_ , \new_[13470]_ , \new_[13471]_ , \new_[13472]_ ,
    \new_[13473]_ , \new_[13474]_ , \new_[13475]_ , \new_[13476]_ ,
    \new_[13477]_ , \new_[13478]_ , \new_[13479]_ , \new_[13480]_ ,
    \new_[13481]_ , \new_[13482]_ , \new_[13483]_ , \new_[13484]_ ,
    \new_[13485]_ , \new_[13486]_ , \new_[13487]_ , \new_[13488]_ ,
    \new_[13489]_ , \new_[13490]_ , \new_[13491]_ , \new_[13492]_ ,
    \new_[13493]_ , \new_[13494]_ , \new_[13495]_ , \new_[13496]_ ,
    \new_[13497]_ , \new_[13498]_ , \new_[13499]_ , \new_[13500]_ ,
    \new_[13501]_ , \new_[13502]_ , \new_[13503]_ , \new_[13504]_ ,
    \new_[13505]_ , \new_[13506]_ , \new_[13507]_ , \new_[13508]_ ,
    \new_[13509]_ , \new_[13510]_ , \new_[13511]_ , \new_[13512]_ ,
    \new_[13513]_ , \new_[13514]_ , \new_[13515]_ , \new_[13516]_ ,
    \new_[13517]_ , \new_[13518]_ , \new_[13519]_ , \new_[13520]_ ,
    \new_[13521]_ , \new_[13522]_ , \new_[13523]_ , \new_[13524]_ ,
    \new_[13525]_ , \new_[13526]_ , \new_[13527]_ , \new_[13528]_ ,
    \new_[13529]_ , \new_[13530]_ , \new_[13531]_ , \new_[13532]_ ,
    \new_[13533]_ , \new_[13534]_ , \new_[13535]_ , \new_[13536]_ ,
    \new_[13537]_ , \new_[13538]_ , \new_[13539]_ , \new_[13540]_ ,
    \new_[13541]_ , \new_[13542]_ , \new_[13543]_ , \new_[13544]_ ,
    \new_[13545]_ , \new_[13546]_ , \new_[13547]_ , \new_[13548]_ ,
    \new_[13549]_ , \new_[13550]_ , \new_[13551]_ , \new_[13552]_ ,
    \new_[13553]_ , \new_[13554]_ , \new_[13555]_ , \new_[13556]_ ,
    \new_[13557]_ , \new_[13558]_ , \new_[13559]_ , \new_[13560]_ ,
    \new_[13561]_ , \new_[13562]_ , \new_[13563]_ , \new_[13564]_ ,
    \new_[13565]_ , \new_[13566]_ , \new_[13567]_ , \new_[13568]_ ,
    \new_[13569]_ , \new_[13570]_ , \new_[13571]_ , \new_[13572]_ ,
    \new_[13573]_ , \new_[13574]_ , \new_[13575]_ , \new_[13576]_ ,
    \new_[13577]_ , \new_[13578]_ , \new_[13579]_ , \new_[13580]_ ,
    \new_[13581]_ , \new_[13582]_ , \new_[13583]_ , \new_[13584]_ ,
    \new_[13585]_ , \new_[13586]_ , \new_[13587]_ , \new_[13588]_ ,
    \new_[13589]_ , \new_[13590]_ , \new_[13591]_ , \new_[13592]_ ,
    \new_[13593]_ , \new_[13594]_ , \new_[13595]_ , \new_[13596]_ ,
    \new_[13597]_ , \new_[13598]_ , \new_[13599]_ , \new_[13600]_ ,
    \new_[13601]_ , \new_[13602]_ , \new_[13603]_ , \new_[13604]_ ,
    \new_[13605]_ , \new_[13606]_ , \new_[13607]_ , \new_[13608]_ ,
    \new_[13609]_ , \new_[13610]_ , \new_[13611]_ , \new_[13612]_ ,
    \new_[13613]_ , \new_[13614]_ , \new_[13615]_ , \new_[13616]_ ,
    \new_[13617]_ , \new_[13618]_ , \new_[13619]_ , \new_[13620]_ ,
    \new_[13621]_ , \new_[13622]_ , \new_[13623]_ , \new_[13624]_ ,
    \new_[13625]_ , \new_[13626]_ , \new_[13627]_ , \new_[13628]_ ,
    \new_[13629]_ , \new_[13630]_ , \new_[13631]_ , \new_[13632]_ ,
    \new_[13633]_ , \new_[13634]_ , \new_[13635]_ , \new_[13636]_ ,
    \new_[13637]_ , \new_[13638]_ , \new_[13639]_ , \new_[13640]_ ,
    \new_[13641]_ , \new_[13642]_ , \new_[13643]_ , \new_[13644]_ ,
    \new_[13645]_ , \new_[13646]_ , \new_[13647]_ , \new_[13648]_ ,
    \new_[13649]_ , \new_[13650]_ , \new_[13651]_ , \new_[13652]_ ,
    \new_[13653]_ , \new_[13654]_ , \new_[13655]_ , \new_[13656]_ ,
    \new_[13657]_ , \new_[13658]_ , \new_[13659]_ , \new_[13660]_ ,
    \new_[13661]_ , \new_[13662]_ , \new_[13663]_ , \new_[13664]_ ,
    \new_[13665]_ , \new_[13666]_ , \new_[13667]_ , \new_[13668]_ ,
    \new_[13669]_ , \new_[13670]_ , \new_[13671]_ , \new_[13672]_ ,
    \new_[13673]_ , \new_[13674]_ , \new_[13675]_ , \new_[13676]_ ,
    \new_[13677]_ , \new_[13678]_ , \new_[13679]_ , \new_[13680]_ ,
    \new_[13681]_ , \new_[13682]_ , \new_[13683]_ , \new_[13684]_ ,
    \new_[13685]_ , \new_[13686]_ , \new_[13687]_ , \new_[13688]_ ,
    \new_[13689]_ , \new_[13690]_ , \new_[13691]_ , \new_[13692]_ ,
    \new_[13693]_ , \new_[13694]_ , \new_[13695]_ , \new_[13696]_ ,
    \new_[13697]_ , \new_[13698]_ , \new_[13699]_ , \new_[13700]_ ,
    \new_[13701]_ , \new_[13702]_ , \new_[13703]_ , \new_[13704]_ ,
    \new_[13705]_ , \new_[13706]_ , \new_[13707]_ , \new_[13708]_ ,
    \new_[13709]_ , \new_[13710]_ , \new_[13711]_ , \new_[13712]_ ,
    \new_[13713]_ , \new_[13714]_ , \new_[13715]_ , \new_[13716]_ ,
    \new_[13717]_ , \new_[13718]_ , \new_[13719]_ , \new_[13720]_ ,
    \new_[13721]_ , \new_[13722]_ , \new_[13723]_ , \new_[13724]_ ,
    \new_[13725]_ , \new_[13726]_ , \new_[13727]_ , \new_[13728]_ ,
    \new_[13729]_ , \new_[13730]_ , \new_[13731]_ , \new_[13732]_ ,
    \new_[13733]_ , \new_[13734]_ , \new_[13735]_ , \new_[13736]_ ,
    \new_[13737]_ , \new_[13738]_ , \new_[13739]_ , \new_[13740]_ ,
    \new_[13741]_ , \new_[13742]_ , \new_[13743]_ , \new_[13744]_ ,
    \new_[13745]_ , \new_[13746]_ , \new_[13747]_ , \new_[13748]_ ,
    \new_[13749]_ , \new_[13750]_ , \new_[13751]_ , \new_[13752]_ ,
    \new_[13753]_ , \new_[13754]_ , \new_[13755]_ , \new_[13756]_ ,
    \new_[13757]_ , \new_[13758]_ , \new_[13759]_ , \new_[13760]_ ,
    \new_[13761]_ , \new_[13762]_ , \new_[13763]_ , \new_[13764]_ ,
    \new_[13765]_ , \new_[13766]_ , \new_[13767]_ , \new_[13768]_ ,
    \new_[13769]_ , \new_[13770]_ , \new_[13771]_ , \new_[13772]_ ,
    \new_[13773]_ , \new_[13774]_ , \new_[13775]_ , \new_[13776]_ ,
    \new_[13777]_ , \new_[13778]_ , \new_[13780]_ , \new_[13781]_ ,
    \new_[13782]_ , \new_[13783]_ , \new_[13784]_ , \new_[13785]_ ,
    \new_[13786]_ , \new_[13787]_ , \new_[13788]_ , \new_[13789]_ ,
    \new_[13790]_ , \new_[13791]_ , \new_[13792]_ , \new_[13793]_ ,
    \new_[13794]_ , \new_[13795]_ , \new_[13796]_ , \new_[13797]_ ,
    \new_[13798]_ , \new_[13799]_ , \new_[13800]_ , \new_[13801]_ ,
    \new_[13802]_ , \new_[13803]_ , \new_[13804]_ , \new_[13805]_ ,
    \new_[13806]_ , \new_[13807]_ , \new_[13808]_ , \new_[13809]_ ,
    \new_[13810]_ , \new_[13811]_ , \new_[13812]_ , \new_[13813]_ ,
    \new_[13814]_ , \new_[13815]_ , \new_[13816]_ , \new_[13817]_ ,
    \new_[13818]_ , \new_[13819]_ , \new_[13820]_ , \new_[13821]_ ,
    \new_[13822]_ , \new_[13823]_ , \new_[13824]_ , \new_[13825]_ ,
    \new_[13826]_ , \new_[13827]_ , \new_[13828]_ , \new_[13829]_ ,
    \new_[13830]_ , \new_[13831]_ , \new_[13832]_ , \new_[13833]_ ,
    \new_[13834]_ , \new_[13835]_ , \new_[13836]_ , \new_[13837]_ ,
    \new_[13838]_ , \new_[13839]_ , \new_[13840]_ , \new_[13841]_ ,
    \new_[13842]_ , \new_[13843]_ , \new_[13844]_ , \new_[13845]_ ,
    \new_[13846]_ , \new_[13847]_ , \new_[13848]_ , \new_[13849]_ ,
    \new_[13850]_ , \new_[13851]_ , \new_[13852]_ , \new_[13853]_ ,
    \new_[13854]_ , \new_[13855]_ , \new_[13856]_ , \new_[13857]_ ,
    \new_[13858]_ , \new_[13859]_ , \new_[13860]_ , \new_[13861]_ ,
    \new_[13862]_ , \new_[13863]_ , \new_[13864]_ , \new_[13865]_ ,
    \new_[13866]_ , \new_[13867]_ , \new_[13868]_ , \new_[13869]_ ,
    \new_[13870]_ , \new_[13871]_ , \new_[13872]_ , \new_[13873]_ ,
    \new_[13874]_ , \new_[13875]_ , \new_[13876]_ , \new_[13877]_ ,
    \new_[13878]_ , \new_[13879]_ , \new_[13880]_ , \new_[13881]_ ,
    \new_[13882]_ , \new_[13883]_ , \new_[13885]_ , \new_[13886]_ ,
    \new_[13887]_ , \new_[13888]_ , \new_[13889]_ , \new_[13890]_ ,
    \new_[13891]_ , \new_[13892]_ , \new_[13893]_ , \new_[13894]_ ,
    \new_[13895]_ , \new_[13896]_ , \new_[13897]_ , \new_[13898]_ ,
    \new_[13899]_ , \new_[13900]_ , \new_[13901]_ , \new_[13902]_ ,
    \new_[13903]_ , \new_[13904]_ , \new_[13905]_ , \new_[13906]_ ,
    \new_[13907]_ , \new_[13908]_ , \new_[13910]_ , \new_[13911]_ ,
    \new_[13912]_ , \new_[13914]_ , \new_[13915]_ , \new_[13916]_ ,
    \new_[13917]_ , \new_[13918]_ , \new_[13919]_ , \new_[13920]_ ,
    \new_[13921]_ , \new_[13922]_ , \new_[13923]_ , \new_[13924]_ ,
    \new_[13925]_ , \new_[13926]_ , \new_[13927]_ , \new_[13928]_ ,
    \new_[13929]_ , \new_[13930]_ , \new_[13931]_ , \new_[13932]_ ,
    \new_[13933]_ , \new_[13934]_ , \new_[13935]_ , \new_[13936]_ ,
    \new_[13937]_ , \new_[13938]_ , \new_[13939]_ , \new_[13940]_ ,
    \new_[13941]_ , \new_[13942]_ , \new_[13943]_ , \new_[13944]_ ,
    \new_[13945]_ , \new_[13946]_ , \new_[13947]_ , \new_[13948]_ ,
    \new_[13949]_ , \new_[13950]_ , \new_[13951]_ , \new_[13952]_ ,
    \new_[13953]_ , \new_[13954]_ , \new_[13955]_ , \new_[13956]_ ,
    \new_[13957]_ , \new_[13958]_ , \new_[13959]_ , \new_[13960]_ ,
    \new_[13961]_ , \new_[13962]_ , \new_[13963]_ , \new_[13964]_ ,
    \new_[13965]_ , \new_[13966]_ , \new_[13967]_ , \new_[13968]_ ,
    \new_[13969]_ , \new_[13970]_ , \new_[13971]_ , \new_[13972]_ ,
    \new_[13973]_ , \new_[13974]_ , \new_[13975]_ , \new_[13976]_ ,
    \new_[13977]_ , \new_[13978]_ , \new_[13979]_ , \new_[13980]_ ,
    \new_[13981]_ , \new_[13982]_ , \new_[13983]_ , \new_[13984]_ ,
    \new_[13985]_ , \new_[13986]_ , \new_[13987]_ , \new_[13988]_ ,
    \new_[13989]_ , \new_[13990]_ , \new_[13991]_ , \new_[13992]_ ,
    \new_[13993]_ , \new_[13994]_ , \new_[13995]_ , \new_[13996]_ ,
    \new_[13997]_ , \new_[13998]_ , \new_[13999]_ , \new_[14000]_ ,
    \new_[14001]_ , \new_[14002]_ , \new_[14003]_ , \new_[14004]_ ,
    \new_[14005]_ , \new_[14006]_ , \new_[14007]_ , \new_[14008]_ ,
    \new_[14009]_ , \new_[14010]_ , \new_[14011]_ , \new_[14012]_ ,
    \new_[14013]_ , \new_[14014]_ , \new_[14015]_ , \new_[14016]_ ,
    \new_[14017]_ , \new_[14018]_ , \new_[14019]_ , \new_[14021]_ ,
    \new_[14022]_ , \new_[14023]_ , \new_[14026]_ , \new_[14027]_ ,
    \new_[14028]_ , \new_[14030]_ , \new_[14031]_ , \new_[14032]_ ,
    \new_[14033]_ , \new_[14034]_ , \new_[14035]_ , \new_[14036]_ ,
    \new_[14037]_ , \new_[14038]_ , \new_[14039]_ , \new_[14040]_ ,
    \new_[14041]_ , \new_[14042]_ , \new_[14043]_ , \new_[14044]_ ,
    \new_[14045]_ , \new_[14046]_ , \new_[14047]_ , \new_[14048]_ ,
    \new_[14049]_ , \new_[14050]_ , \new_[14051]_ , \new_[14052]_ ,
    \new_[14053]_ , \new_[14054]_ , \new_[14055]_ , \new_[14056]_ ,
    \new_[14057]_ , \new_[14058]_ , \new_[14059]_ , \new_[14060]_ ,
    \new_[14061]_ , \new_[14062]_ , \new_[14063]_ , \new_[14064]_ ,
    \new_[14065]_ , \new_[14066]_ , \new_[14067]_ , \new_[14068]_ ,
    \new_[14069]_ , \new_[14070]_ , \new_[14071]_ , \new_[14072]_ ,
    \new_[14073]_ , \new_[14074]_ , \new_[14075]_ , \new_[14076]_ ,
    \new_[14077]_ , \new_[14078]_ , \new_[14079]_ , \new_[14080]_ ,
    \new_[14081]_ , \new_[14082]_ , \new_[14083]_ , \new_[14084]_ ,
    \new_[14085]_ , \new_[14086]_ , \new_[14087]_ , \new_[14088]_ ,
    \new_[14089]_ , \new_[14090]_ , \new_[14091]_ , \new_[14093]_ ,
    \new_[14094]_ , \new_[14095]_ , \new_[14096]_ , \new_[14097]_ ,
    \new_[14098]_ , \new_[14099]_ , \new_[14100]_ , \new_[14101]_ ,
    \new_[14102]_ , \new_[14103]_ , \new_[14104]_ , \new_[14105]_ ,
    \new_[14106]_ , \new_[14107]_ , \new_[14108]_ , \new_[14109]_ ,
    \new_[14110]_ , \new_[14111]_ , \new_[14112]_ , \new_[14113]_ ,
    \new_[14114]_ , \new_[14115]_ , \new_[14116]_ , \new_[14117]_ ,
    \new_[14118]_ , \new_[14119]_ , \new_[14120]_ , \new_[14121]_ ,
    \new_[14122]_ , \new_[14123]_ , \new_[14124]_ , \new_[14125]_ ,
    \new_[14126]_ , \new_[14127]_ , \new_[14128]_ , \new_[14129]_ ,
    \new_[14130]_ , \new_[14131]_ , \new_[14132]_ , \new_[14133]_ ,
    \new_[14134]_ , \new_[14135]_ , \new_[14136]_ , \new_[14137]_ ,
    \new_[14138]_ , \new_[14139]_ , \new_[14140]_ , \new_[14141]_ ,
    \new_[14142]_ , \new_[14143]_ , \new_[14144]_ , \new_[14145]_ ,
    \new_[14146]_ , \new_[14147]_ , \new_[14148]_ , \new_[14149]_ ,
    \new_[14150]_ , \new_[14151]_ , \new_[14152]_ , \new_[14153]_ ,
    \new_[14154]_ , \new_[14155]_ , \new_[14156]_ , \new_[14157]_ ,
    \new_[14158]_ , \new_[14159]_ , \new_[14160]_ , \new_[14161]_ ,
    \new_[14162]_ , \new_[14163]_ , \new_[14164]_ , \new_[14165]_ ,
    \new_[14166]_ , \new_[14167]_ , \new_[14168]_ , \new_[14169]_ ,
    \new_[14170]_ , \new_[14171]_ , \new_[14172]_ , \new_[14173]_ ,
    \new_[14174]_ , \new_[14175]_ , \new_[14176]_ , \new_[14177]_ ,
    \new_[14178]_ , \new_[14179]_ , \new_[14180]_ , \new_[14181]_ ,
    \new_[14182]_ , \new_[14183]_ , \new_[14184]_ , \new_[14185]_ ,
    \new_[14186]_ , \new_[14187]_ , \new_[14188]_ , \new_[14189]_ ,
    \new_[14190]_ , \new_[14191]_ , \new_[14192]_ , \new_[14193]_ ,
    \new_[14194]_ , n266, n271, n276, n281, n286, n291, n296, n301, n306,
    n311, n316, n321, n326, n331, n336, n341, n346, n351, n356, n361, n366,
    n371, n376, n381, n386, n391, n396, n401, n406, n411, n416, n421, n426,
    n431, n436, n441, n446, n451, n456, n461, n466, n471, n476, n481, n486,
    n491, n496, n501, n506, n511, n516, n521, n526, n531, n536, n541, n546,
    n551, n556, n561, n566, n571, n576, n581, n586, n591, n596, n601, n606,
    n611, n616, n621, n626, n631, n636, n641, n646, n651, n656, n661, n666,
    n671, n676, n681, n686, n691, n696, n701, n706, n711, n716, n721, n726,
    n731, n736, n741, n746, n751, n756, n761, n766, n771, n776, n781, n786,
    n791, n796, n801, n806, n811, n816, n821, n826, n831, n836, n841, n846,
    n851, n856, n861, n866, n871, n876, n881, n886, n891, n896, n901, n906,
    n911, n916, n921, n926, n931, n936, n941, n946, n951, n956, n961, n966,
    n971, n976, n981, n986, n991, n996, n1001, n1006, n1011, n1016, n1021,
    n1026, n1031, n1036, n1041, n1046, n1051, n1056, n1061, n1066, n1071,
    n1076, n1081, n1086, n1091, n1096, n1101, n1106, n1111, n1116, n1121,
    n1126, n1131, n1136, n1141, n1146, n1151, n1156, n1161, n1166, n1171,
    n1176, n1181, n1186, n1191, n1196, n1201, n1206, n1211, n1216, n1221,
    n1226, n1231, n1236, n1241, n1246, n1251, n1256, n1261, n1266, n1271,
    n1276, n1281, n1286, n1291, n1296, n1301, n1306, n1311, n1316, n1321,
    n1326, n1331, n1336, n1341, n1346, n1351, n1356, n1361, n1366, n1371,
    n1376, n1381, n1386, n1391, n1396, n1401, n1406, n1411, n1416, n1421,
    n1426, n1431, n1436, n1441, n1446, n1451, n1456, n1461, n1466, n1471,
    n1476, n1481, n1486, n1491, n1496, n1501, n1506, n1511, n1516, n1521,
    n1526, n1531, n1536, n1541, n1546, n1551, n1556, n1561, n1566, n1571,
    n1576, n1581, n1586, n1591, n1596, n1601, n1606, n1611, n1616, n1621,
    n1626, n1631, n1636, n1641, n1646, n1651, n1656, n1661, n1666, n1671,
    n1676, n1681, n1686, n1691, n1696, n1701, n1706, n1711, n1716, n1721,
    n1726, n1731, n1736, n1741, n1746, n1751, n1756, n1761, n1766, n1771,
    n1776, n1781, n1786, n1791, n1796, n1801, n1806, n1811, n1816, n1821,
    n1826, n1831, n1836, n1841, n1846, n1851, n1856, n1861, n1866, n1871,
    n1876, n1881, n1886, n1891, n1896, n1901, n1906, n1911, n1916, n1921,
    n1926, n1931, n1936, n1941, n1946, n1951, n1956, n1961, n1966, n1971,
    n1976, n1981, n1986, n1991, n1996, n2001, n2006, n2011, n2016, n2021,
    n2026, n2031, n2036, n2041, n2046, n2051, n2056, n2061, n2066, n2071,
    n2076, n2081, n2086, n2091, n2096, n2101, n2106, n2111, n2116, n2121,
    n2126, n2131, n2136, n2141, n2146, n2151, n2156, n2161, n2166, n2171,
    n2176, n2181, n2186, n2191, n2196, n2201, n2206, n2211, n2216, n2221,
    n2226, n2231, n2236, n2241, n2246, n2251, n2256, n2261, n2266, n2271,
    n2276, n2281, n2286, n2291, n2296, n2301, n2306, n2311, n2316, n2321,
    n2326, n2331, n2336, n2341, n2346, n2351, n2356, n2361, n2366, n2371,
    n2376, n2381, n2386, n2391, n2396, n2401, n2406, n2411, n2416, n2421,
    n2426, n2431, n2436, n2441, n2446, n2451, n2456, n2461, n2466, n2471,
    n2476, n2481, n2486, n2491, n2496, n2501, n2506, n2511, n2516, n2521,
    n2526, n2531, n2536, n2541, n2546, n2551, n2556, n2561, n2566, n2571,
    n2576, n2581, n2586, n2591, n2596, n2601, n2606, n2611, n2616, n2621,
    n2626, n2631, n2636, n2641, n2646, n2651, n2656, n2661, n2666, n2671,
    n2676, n2681, n2686, n2691, n2696, n2701, n2706, n2711, n2716, n2721,
    n2726, n2731, n2736, n2741, n2746, n2751, n2756, n2761, n2766, n2771,
    n2776, n2781, n2786, n2791, n2796, n2801, n2806, n2811, n2816, n2821,
    n2826, n2831, n2836, n2841, n2846, n2851, n2856, n2861, n2866, n2871,
    n2876, n2881, n2886, n2891, n2896, n2901, n2906, n2911, n2916, n2921,
    n2926, n2931, n2936, n2941, n2946, n2951, n2956, n2961, n2966, n2971,
    n2976, n2981, n2986, n2991, n2996, n3001, n3006, n3011, n3016, n3021,
    n3026, n3031, n3036, n3041, n3046, n3051, n3056, n3061, n3066, n3071,
    n3076, n3081, n3086, n3091, n3096, n3101, n3106, n3111, n3116, n3121,
    n3126, n3131, n3136, n3141, n3146, n3151, n3156, n3161, n3166, n3171,
    n3176, n3181, n3186, n3191, n3196, n3201, n3206, n3211, n3216, n3221,
    n3226, n3231, n3236, n3241, n3246, n3251, n3256, n3261, n3266, n3271,
    n3276, n3281, n3286, n3291, n3296, n3301, n3306, n3311, n3316, n3321,
    n3326, n3331, n3336, n3341, n3346, n3351, n3356, n3361, n3366, n3371,
    n3376, n3381, n3386, n3391, n3396, n3401, n3406, n3411, n3416, n3421,
    n3426, n3431, n3436, n3441, n3446, n3451, n3456, n3461, n3466, n3471,
    n3476, n3481, n3486, n3491, n3496, n3501, n3506, n3511, n3516, n3521,
    n3526, n3531, n3536, n3541, n3546, n3551, n3556, n3561, n3566, n3571,
    n3576, n3581, n3586, n3591, n3596, n3601, n3606, n3611, n3616, n3621,
    n3626, n3631, n3636, n3641, n3646, n3651, n3656, n3661, n3666, n3671,
    n3676, n3681, n3686, n3691, n3696, n3701, n3706, n3711, n3716, n3721,
    n3726, n3731, n3736, n3741, n3746, n3751, n3756, n3761, n3766, n3771,
    n3776, n3781, n3786, n3791, n3796, n3801, n3806, n3811, n3816, n3821,
    n3826, n3831, n3836, n3841, n3846, n3851, n3856, n3861, n3866, n3871,
    n3876, n3881, n3886, n3891, n3896, n3901, n3906, n3911, n3916, n3921,
    n3926, n3931, n3936, n3941, n3946, n3951, n3956, n3961, n3966, n3971,
    n3976, n3981, n3986, n3991, n3996, n4001, n4006, n4011, n4016, n4021,
    n4026, n4031, n4036, n4041, n4046, n4051, n4056, n4061, n4066, n4071,
    n4076, n4081, n4086, n4091, n4096, n4101, n4106, n4111, n4116, n4121,
    n4126, n4131, n4136, n4141, n4146, n4151, n4156, n4161, n4166, n4171,
    n4176, n4181, n4186, n4191, n4196, n4201, n4206, n4211, n4216, n4221,
    n4226, n4231, n4236, n4241, n4246, n4251, n4256, n4261, n4266, n4271,
    n4276, n4281, n4286, n4291, n4296, n4301, n4306, n4311, n4316, n4321,
    n4326, n4331, n4336, n4341, n4346, n4351, n4356, n4361, n4366, n4371,
    n4376, n4381, n4386, n4391, n4396, n4401, n4406, n4411, n4416, n4421,
    n4426, n4431, n4436, n4441, n4446, n4451, n4456, n4461, n4466, n4471,
    n4476, n4481, n4486, n4491, n4496, n4501, n4506, n4511, n4516, n4521,
    n4526, n4531, n4536, n4541, n4546, n4551, n4556, n4561, n4566, n4571,
    n4576, n4581, n4586, n4591, n4596, n4601, n4606, n4611, n4616, n4621,
    n4626, n4631, n4636, n4641, n4646, n4651, n4656, n4661, n4666, n4671,
    n4676, n4681, n4686, n4691, n4696, n4701, n4706, n4711, n4716, n4721,
    n4726, n4731, n4736, n4741, n4746, n4751, n4756, n4761, n4766, n4771,
    n4776, n4781, n4786, n4791, n4796, n4801, n4806, n4811, n4816, n4821,
    n4826, n4831, n4836, n4841, n4846, n4851, n4856, n4861, n4866, n4871,
    n4876, n4881, n4886, n4891, n4896, n4901, n4906, n4911, n4916, n4921,
    n4926, n4931, n4936, n4941, n4946, n4951, n4956, n4961, n4966, n4971,
    n4976, n4981, n4986, n4991, n4996, n5001, n5006, n5011, n5016, n5021,
    n5026, n5031, n5036, n5041, n5046, n5051, n5056, n5061, n5066, n5071,
    n5076, n5081, n5086, n5091, n5096, n5101, n5106, n5111, n5116, n5121,
    n5126, n5131, n5136, n5141, n5146, n5151, n5156, n5161, n5166, n5171,
    n5176, n5181, n5186, n5191, n5196, n5201, n5206, n5211, n5216, n5221,
    n5226, n5231, n5236, n5241, n5246, n5251, n5256, n5261, n5266, n5271,
    n5276, n5281, n5286, n5291, n5296, n5301, n5306, n5311, n5316, n5321,
    n5326, n5331, n5336, n5341, n5346, n5351, n5356, n5361, n5366, n5371,
    n5376, n5381, n5386, n5391, n5396, n5401, n5406, n5411, n5416, n5421,
    n5426, n5431, n5436, n5441, n5446, n5451, n5456, n5461, n5466, n5471,
    n5476, n5481, n5486, n5491, n5496, n5501, n5506, n5511, n5516, n5521,
    n5526, n5531, n5536, n5541, n5546, n5551, n5556, n5561, n5566, n5571,
    n5576, n5581, n5586, n5591, n5596, n5601, n5606, n5611, n5616, n5621,
    n5626, n5631, n5636, n5641, n5646, n5651, n5656, n5661, n5666, n5671,
    n5676, n5681, n5686, n5691, n5696, n5701, n5706, n5711, n5716, n5721,
    n5726, n5731, n5736, n5741, n5746, n5751, n5756, n5761, n5766, n5771,
    n5776, n5781, n5786, n5791, n5796, n5801, n5806, n5811, n5816, n5821,
    n5826, n5831, n5836, n5841, n5846, n5851, n5856, n5861, n5866, n5871,
    n5876, n5881, n5886, n5891, n5896, n5901, n5906, n5911, n5916, n5921,
    n5926, n5931, n5936, n5941, n5946, n5951, n5956, n5961, n5966, n5971,
    n5976, n5981, n5986, n5991, n5996, n6001, n6006, n6011, n6016, n6021,
    n6026, n6031, n6036, n6041, n6046, n6051, n6056, n6061, n6066, n6071,
    n6076, n6081, n6086, n6091, n6096, n6101, n6106, n6111, n6116, n6121,
    n6126, n6131, n6136, n6141, n6146, n6151, n6156, n6161, n6166, n6171,
    n6176, n6181, n6186, n6191, n6196, n6201, n6206, n6211, n6216, n6221,
    n6226, n6231, n6236, n6241, n6246, n6251, n6256, n6261, n6266, n6271,
    n6276, n6281, n6286, n6291, n6296, n6301, n6306, n6311, n6316, n6321,
    n6326, n6331, n6336, n6341, n6346, n6351, n6356, n6361, n6366, n6371,
    n6376, n6381, n6386, n6391, n6396, n6401, n6406, n6411, n6416, n6421,
    n6426, n6431, n6436, n6441, n6446, n6451, n6456, n6461, n6466, n6471,
    n6476, n6481, n6486, n6491, n6496, n6501, n6506, n6511, n6516, n6521,
    n6526, n6531, n6536, n6541, n6546, n6551, n6556, n6561, n6566, n6571,
    n6576, n6581, n6586, n6591, n6596, n6601, n6606, n6611, n6616, n6621,
    n6626, n6631, n6636, n6641, n6646, n6651, n6656, n6661, n6666, n6671,
    n6676, n6681, n6686, n6691, n6696, n6701, n6706, n6711, n6716, n6721,
    n6726, n6731, n6736, n6741, n6746, n6751, n6756, n6761, n6766, n6771,
    n6776, n6781, n6786, n6791, n6796, n6801, n6806, n6811, n6816, n6821,
    n6826, n6831, n6836, n6841, n6846, n6851, n6856, n6861, n6866, n6871,
    n6876, n6881, n6886, n6891, n6896, n6901, n6906, n6911, n6916, n6921,
    n6926, n6931, n6936, n6941, n6946, n6951, n6956, n6961, n6966, n6971,
    n6976, n6981, n6986, n6991, n6996, n7001, n7006, n7011, n7016, n7021,
    n7026, n7031, n7036, n7041, n7046, n7051, n7056, n7061, n7066, n7071,
    n7076, n7081, n7086, n7091, n7096, n7101, n7106, n7111, n7116, n7121,
    n7126, n7131, n7136, n7141, n7146, n7151, n7156, n7161, n7166, n7171,
    n7176, n7181, n7186, n7191, n7196, n7201, n7206, n7211, n7216, n7221,
    n7226, n7231, n7236, n7241, n7246, n7251, n7256, n7261, n7266, n7271,
    n7276, n7281, n7286, n7291, n7296, n7301, n7306, n7311, n7316, n7321,
    n7326, n7331, n7336, n7341, n7346, n7351, n7356, n7361, n7366, n7371,
    n7376, n7381, n7386, n7391, n7396, n7401, n7406, n7411, n7416, n7421,
    n7426, n7431, n7436, n7441, n7446, n7451, n7456, n7461, n7466, n7471,
    n7476, n7481, n7486, n7491, n7496, n7501, n7506, n7511, n7516, n7521,
    n7526, n7531, n7536, n7541, n7546, n7551, n7556, n7561, n7566, n7571,
    n7576, n7581, n7586, n7591, n7596, n7601, n7606, n7611, n7616, n7621,
    n7626, n7631, n7636, n7641, n7646, n7651, n7656, n7661, n7666, n7671,
    n7676, n7681, n7686, n7691, n7696, n7701, n7706, n7711, n7716, n7721,
    n7726, n7731, n7736, n7741, n7746, n7751, n7756, n7761, n7766, n7771,
    n7776, n7781, n7786, n7791, n7796, n7801, n7806, n7811, n7816, n7821,
    n7826, n7831, n7836, n7841, n7846, n7851, n7856, n7861, n7866, n7871,
    n7876, n7881, n7886, n7891, n7896, n7901, n7906, n7911, n7916, n7921,
    n7926, n7931, n7936, n7941, n7946, n7951, n7956, n7961, n7966, n7971,
    n7976, n7981, n7986, n7991, n7996, n8001, n8006, n8011, n8016, n8021,
    n8026, n8031, n8036, n8041, n8046, n8051, n8056, n8061, n8066, n8071,
    n8076, n8081, n8086, n8091, n8096, n8101, n8106, n8111, n8116, n8121,
    n8126, n8131, n8136, n8141, n8146, n8151, n8156, n8161, n8166, n8171,
    n8176, n8181, n8186, n8191, n8196, n8201, n8206, n8211, n8216, n8221,
    n8226, n8231, n8236, n8241, n8246, n8251, n8256, n8261, n8266, n8271,
    n8276, n8281, n8286, n8291, n8296, n8301, n8306, n8311, n8316, n8321,
    n8326, n8331, n8336, n8341, n8346, n8351, n8356, n8361, n8366, n8371,
    n8376, n8381, n8386, n8391, n8396, n8401, n8406, n8411, n8416, n8421,
    n8426, n8431, n8436, n8441, n8446, n8451, n8456, n8461, n8466, n8471,
    n8476, n8481, n8486, n8491, n8496, n8501, n8506, n8511, n8516, n8521,
    n8526, n8531, n8536, n8541, n8546, n8551, n8556, n8561, n8566, n8571,
    n8576, n8581, n8586, n8591, n8596, n8601, n8606, n8611, n8616, n8621,
    n8626, n8631, n8636, n8641, n8646, n8651, n8656, n8661, n8666, n8671,
    n8676, n8681, n8686, n8691, n8696, n8701, n8706, n8711, n8716, n8721,
    n8726, n8731, n8736, n8741, n8746, n8751, n8756, n8761, n8766, n8771,
    n8776, n8781, n8786, n8791, n8796, n8801, n8806, n8811, n8816, n8821,
    n8826, n8831, n8836, n8841, n8846, n8851, n8856, n8861, n8866, n8871,
    n8876, n8881, n8886, n8891, n8896, n8901, n8906, n8911, n8916, n8921,
    n8926, n8931, n8936, n8941, n8946, n8951, n8956, n8961, n8966, n8971,
    n8976, n8981, n8986, n8991, n8996, n9001, n9006, n9011, n9016, n9021,
    n9026, n9031, n9036, n9041, n9046, n9051, n9056, n9061, n9066, n9071,
    n9076, n9081, n9086, n9091, n9096, n9101, n9106, n9111, n9116, n9121,
    n9126, n9131, n9136, n9141, n9146, n9151, n9156, n9161, n9166, n9171,
    n9176, n9181, n9186, n9191, n9196, n9201, n9206, n9211, n9216, n9221,
    n9226, n9231, n9236, n9241, n9246, n9251, n9256, n9261, n9266, n9271,
    n9276, n9281, n9286, n9291, n9296, n9301, n9306, n9311, n9316, n9321,
    n9326, n9331, n9336, n9341, n9346, n9351, n9356, n9361, n9366, n9371,
    n9376, n9381, n9386, n9391, n9396, n9401, n9406, n9411, n9416, n9421,
    n9426, n9431, n9436, n9441, n9446, n9451, n9456, n9461, n9466, n9471,
    n9476, n9481, n9486, n9491, n9496, n9501, n9506, n9511, n9516, n9521,
    n9526, n9531, n9536, n9541, n9546, n9551, n9556, n9561, n9566, n9571,
    n9576, n9581, n9586, n9591, n9596, n9601, n9606, n9611, n9616, n9621,
    n9626, n9631, n9636, n9641, n9646, n9651, n9656, n9661, n9666, n9671,
    n9676, n9681, n9686, n9691, n9696, n9701, n9706, n9711, n9716, n9721,
    n9726, n9731, n9736, n9741, n9746, n9751, n9756, n9761, n9766, n9771,
    n9776, n9781, n9786, n9791, n9796, n9801, n9806, n9811, n9816, n9821,
    n9826, n9831, n9836, n9841, n9846, n9851, n9856, n9861, n9866, n9871,
    n9876, n9881, n9886, n9891, n9896, n9901, n9906, n9911, n9916, n9921,
    n9926, n9931, n9936, n9941, n9946, n9951, n9956, n9961, n9966, n9971,
    n9976, n9981, n9986, n9991, n9996, n10001, n10006, n10011, n10016,
    n10021, n10026, n10031, n10036, n10041, n10046, n10051, n10056, n10061,
    n10066, n10071, n10076, n10081, n10086, n10091, n10096, n10101, n10106,
    n10111, n10116, n10121, n10126, n10131, n10136, n10141, n10146, n10151,
    n10156, n10161, n10166, n10171, n10176, n10181, n10186, n10191, n10196,
    n10201, n10206, n10211, n10216, n10221, n10226, n10231, n10236, n10241,
    n10246, n10251, n10256, n10261, n10266, n10271, n10276, n10281, n10286,
    n10291, n10296, n10301, n10306, n10311, n10316, n10321, n10326, n10331,
    n10336, n10341, n10346, n10351, n10356, n10361, n10366, n10371, n10376,
    n10381, n10386, n10391, n10396, n10401, n10406, n10411, n10416, n10421,
    n10426, n10431, n10436, n10441, n10446, n10451, n10456, n10461, n10466,
    n10471, n10476, n10481, n10486, n10491, n10496, n10501, n10506, n10511,
    n10516, n10521, n10526, n10531, n10536, n10541, n10546, n10551, n10556,
    n10561, n10566, n10571, n10576, n10581, n10586, n10591, n10596, n10601,
    n10606, n10611, n10616, n10621, n10626, n10631, n10636, n10641, n10646,
    n10651, n10656, n10661, n10666, n10671, n10676, n10681, n10686, n10691,
    n10696, n10701, n10706, n10711, n10716, n10721, n10726, n10731, n10736,
    n10741, n10746, n10751, n10756, n10761, n10766, n10771, n10776, n10781,
    n10786, n10791, n10796, n10801, n10806, n10811, n10816, n10821, n10826,
    n10831, n10836, n10841, n10846, n10851, n10856, n10861, n10866, n10871,
    n10876, n10881, n10886, n10891, n10896, n10901, n10906, n10911, n10916,
    n10921, n10926, n10931, n10936, n10941, n10946, n10951, n10956, n10961,
    n10966, n10971, n10976, n10981, n10986, n10991, n10996, n11001, n11006,
    n11011, n11016, n11021, n11026, n11031, n11036, n11041, n11046, n11051,
    n11056, n11061, n11066, n11071, n11076, n11081, n11086, n11091, n11096,
    n11101, n11106, n11111, n11116, n11121, n11126, n11131, n11136, n11141,
    n11146, n11151, n11156, n11161, n11166, n11171, n11176, n11181, n11186,
    n11191, n11196, n11201, n11206, n11211, n11216, n11221, n11226, n11231,
    n11236, n11241, n11246, n11251, n11256;
  assign \new_[2331]_  = 1'b0;
  assign wb_err_o = \new_[2331]_ ;
  assign sdata_pad_o = \\u0_slt0_r_reg[15] ;
  assign n266 = ~\new_[7960]_  | ~\new_[2336]_  | ~\new_[7934]_ ;
  assign \new_[2336]_  = ~\new_[7963]_  & (~\new_[2337]_  | ~\new_[8483]_ );
  assign \new_[2337]_  = \\u0_slt0_r_reg[14] ;
  assign n271 = \new_[4591]_  ? \new_[7966]_  : \new_[2339]_ ;
  assign \new_[2339]_  = \\u0_slt0_r_reg[13] ;
  assign n276 = \new_[4648]_  ? \new_[7966]_  : \new_[2341]_ ;
  assign \new_[2341]_  = \\u0_slt0_r_reg[12] ;
  assign n281 = \new_[4586]_  ? \new_[7966]_  : \new_[2343]_ ;
  assign \new_[2343]_  = \\u0_slt0_r_reg[11] ;
  assign n286 = \new_[4587]_  ? \new_[7966]_  : \new_[2345]_ ;
  assign \new_[2345]_  = \\u0_slt0_r_reg[10] ;
  assign n291 = \new_[2347]_  & \new_[8483]_ ;
  assign \new_[2347]_  = \\u0_slt0_r_reg[9] ;
  assign n296 = \new_[4588]_  ? \new_[7937]_  : \new_[2349]_ ;
  assign \new_[2349]_  = \\u0_slt0_r_reg[8] ;
  assign n301 = \new_[4589]_  ? \new_[7966]_  : \new_[2351]_ ;
  assign \new_[2351]_  = \\u0_slt0_r_reg[7] ;
  assign n306 = \new_[4581]_  ? \new_[7966]_  : \new_[2353]_ ;
  assign \new_[2353]_  = \\u0_slt0_r_reg[6] ;
  assign n311 = ~\new_[2355]_  | ~\new_[7960]_ ;
  assign \new_[2355]_  = ~\new_[2356]_  | ~\new_[8483]_ ;
  assign \new_[2356]_  = \\u0_slt0_r_reg[5] ;
  assign n316 = \new_[2358]_  & \new_[7962]_ ;
  assign \new_[2358]_  = \\u0_slt0_r_reg[4] ;
  assign n321 = \new_[2360]_  & \new_[8483]_ ;
  assign \new_[2360]_  = \\u0_slt0_r_reg[3] ;
  assign n326 = \new_[2362]_  & \new_[7962]_ ;
  assign \new_[2362]_  = \\u0_slt0_r_reg[2] ;
  assign n331 = \new_[2364]_  & \new_[8483]_ ;
  assign \new_[2364]_  = \\u0_slt0_r_reg[1] ;
  assign n336 = \new_[2366]_  & \new_[7962]_ ;
  assign \new_[2366]_  = \\u0_slt0_r_reg[0] ;
  assign n341 = \new_[2368]_  & \new_[7962]_ ;
  assign \new_[2368]_  = \\u0_slt1_r_reg[19] ;
  assign n346 = \new_[5055]_  ? \new_[7966]_  : \new_[2370]_ ;
  assign \new_[2370]_  = \\u0_slt1_r_reg[18] ;
  assign n351 = \new_[4894]_  ? \new_[7966]_  : \new_[2372]_ ;
  assign \new_[2372]_  = \\u0_slt1_r_reg[17] ;
  assign n356 = \new_[5054]_  ? \new_[7937]_  : \new_[2374]_ ;
  assign \new_[2374]_  = \\u0_slt1_r_reg[16] ;
  assign n361 = \new_[5053]_  ? \new_[8483]_  : \new_[2376]_ ;
  assign \new_[2376]_  = \\u0_slt1_r_reg[15] ;
  assign n366 = \new_[5052]_  ? \new_[8483]_  : \new_[2378]_ ;
  assign \new_[2378]_  = \\u0_slt1_r_reg[14] ;
  assign n371 = \new_[5688]_  ? \new_[8483]_  : \new_[2380]_ ;
  assign \new_[2380]_  = \\u0_slt1_r_reg[13] ;
  assign n376 = \new_[5051]_  ? \new_[7966]_  : \new_[2382]_ ;
  assign \new_[2382]_  = \\u0_slt1_r_reg[12] ;
  assign n381 = \new_[5050]_  ? \new_[7966]_  : \new_[2384]_ ;
  assign \new_[2384]_  = \\u0_slt1_r_reg[11] ;
  assign n386 = \new_[2386]_  & \new_[7962]_ ;
  assign \new_[2386]_  = \\u0_slt1_r_reg[10] ;
  assign n391 = \new_[2388]_  & \new_[7962]_ ;
  assign \new_[2388]_  = \\u0_slt1_r_reg[9] ;
  assign n396 = \new_[2390]_  & \new_[7962]_ ;
  assign \new_[2390]_  = \\u0_slt1_r_reg[8] ;
  assign n401 = \new_[2392]_  & \new_[8483]_ ;
  assign \new_[2392]_  = \\u0_slt1_r_reg[7] ;
  assign n406 = \new_[2394]_  & \new_[7962]_ ;
  assign \new_[2394]_  = \\u0_slt1_r_reg[6] ;
  assign n411 = \new_[2396]_  & \new_[7962]_ ;
  assign \new_[2396]_  = \\u0_slt1_r_reg[5] ;
  assign n416 = \new_[2398]_  & \new_[7962]_ ;
  assign \new_[2398]_  = \\u0_slt1_r_reg[4] ;
  assign n421 = \new_[2400]_  & \new_[7962]_ ;
  assign \new_[2400]_  = \\u0_slt1_r_reg[3] ;
  assign n426 = \new_[2402]_  & \new_[7962]_ ;
  assign \new_[2402]_  = \\u0_slt1_r_reg[2] ;
  assign n431 = \new_[2404]_  & \new_[7962]_ ;
  assign \new_[2404]_  = \\u0_slt1_r_reg[1] ;
  assign n436 = \new_[2406]_  & \new_[7962]_ ;
  assign \new_[2406]_  = \\u0_slt1_r_reg[0] ;
  assign n441 = \new_[2408]_  & \new_[7962]_ ;
  assign \new_[2408]_  = \\u0_slt2_r_reg[19] ;
  assign n446 = \new_[13632]_  ? \new_[7966]_  : \new_[2410]_ ;
  assign \new_[2410]_  = \\u0_slt2_r_reg[18] ;
  assign n451 = \new_[13614]_  ? \new_[7937]_  : \new_[2412]_ ;
  assign \new_[2412]_  = \\u0_slt2_r_reg[17] ;
  assign n456 = \new_[13611]_  ? \new_[7966]_  : \new_[2414]_ ;
  assign \new_[2414]_  = \\u0_slt2_r_reg[16] ;
  assign n461 = \new_[13324]_  ? \new_[8501]_  : \new_[2416]_ ;
  assign \new_[2416]_  = \\u0_slt2_r_reg[15] ;
  assign n466 = \new_[13689]_  ? \new_[7937]_  : \new_[2418]_ ;
  assign \new_[2418]_  = \\u0_slt2_r_reg[14] ;
  assign n471 = \new_[13813]_  ? \new_[7937]_  : \new_[2420]_ ;
  assign \new_[2420]_  = \\u0_slt2_r_reg[13] ;
  assign n476 = \new_[13730]_  ? \new_[7937]_  : \new_[2422]_ ;
  assign \new_[2422]_  = \\u0_slt2_r_reg[12] ;
  assign n481 = \new_[13505]_  ? \new_[7937]_  : \new_[2424]_ ;
  assign \new_[2424]_  = \\u0_slt2_r_reg[11] ;
  assign n486 = \new_[13269]_  ? \new_[7962]_  : \new_[2426]_ ;
  assign \new_[2426]_  = \\u0_slt2_r_reg[10] ;
  assign n491 = \new_[13671]_  ? \new_[7966]_  : \new_[2428]_ ;
  assign \new_[2428]_  = \\u0_slt2_r_reg[9] ;
  assign n496 = \new_[13370]_  ? \new_[7937]_  : \new_[2430]_ ;
  assign \new_[2430]_  = \\u0_slt2_r_reg[8] ;
  assign n501 = \new_[13704]_  ? \new_[7937]_  : \new_[2432]_ ;
  assign \new_[2432]_  = \\u0_slt2_r_reg[7] ;
  assign n506 = \new_[13790]_  ? \new_[7937]_  : \new_[2434]_ ;
  assign \new_[2434]_  = \\u0_slt2_r_reg[6] ;
  assign n511 = \new_[13382]_  ? \new_[7937]_  : \new_[2436]_ ;
  assign \new_[2436]_  = \\u0_slt2_r_reg[5] ;
  assign n516 = \new_[13509]_  ? \new_[7937]_  : \new_[2438]_ ;
  assign \new_[2438]_  = \\u0_slt2_r_reg[4] ;
  assign n521 = \new_[13218]_  ? \new_[7937]_  : \new_[2440]_ ;
  assign \new_[2440]_  = \\u0_slt2_r_reg[3] ;
  assign n526 = \new_[2442]_  & \new_[7962]_ ;
  assign \new_[2442]_  = \\u0_slt2_r_reg[2] ;
  assign n531 = \new_[2444]_  & \new_[8483]_ ;
  assign \new_[2444]_  = \\u0_slt2_r_reg[1] ;
  assign n536 = \new_[2446]_  & \new_[8483]_ ;
  assign \new_[2446]_  = \\u0_slt2_r_reg[0] ;
  assign n541 = \new_[2448]_  & \new_[7962]_ ;
  assign \new_[2448]_  = \\u0_slt3_r_reg[19] ;
  assign n546 = \new_[13339]_  ? \new_[7966]_  : \new_[2450]_ ;
  assign \new_[2450]_  = \\u0_slt3_r_reg[18] ;
  assign n551 = \new_[13855]_  ? \new_[7966]_  : \new_[2452]_ ;
  assign \new_[2452]_  = \\u0_slt3_r_reg[17] ;
  assign n556 = \new_[13733]_  ? \new_[7937]_  : \new_[2454]_ ;
  assign \new_[2454]_  = \\u0_slt3_r_reg[16] ;
  assign n561 = \new_[13415]_  ? \new_[7962]_  : \new_[2456]_ ;
  assign \new_[2456]_  = \\u0_slt3_r_reg[15] ;
  assign n566 = \new_[13413]_  ? \new_[7962]_  : \new_[2458]_ ;
  assign \new_[2458]_  = \\u0_slt3_r_reg[14] ;
  assign n571 = \new_[13442]_  ? \new_[8483]_  : \new_[2460]_ ;
  assign \new_[2460]_  = \\u0_slt3_r_reg[13] ;
  assign n576 = \new_[13579]_  ? \new_[8483]_  : \new_[2462]_ ;
  assign \new_[2462]_  = \\u0_slt3_r_reg[12] ;
  assign n581 = \new_[13657]_  ? \new_[7937]_  : \new_[2464]_ ;
  assign \new_[2464]_  = \\u0_slt3_r_reg[11] ;
  assign n586 = \new_[13207]_  ? \new_[7962]_  : \new_[2466]_ ;
  assign \new_[2466]_  = \\u0_slt3_r_reg[10] ;
  assign n591 = \new_[13220]_  ? \new_[7962]_  : \new_[2468]_ ;
  assign \new_[2468]_  = \\u0_slt3_r_reg[9] ;
  assign n596 = \new_[13299]_  ? \new_[8501]_  : \new_[2470]_ ;
  assign \new_[2470]_  = \\u0_slt3_r_reg[8] ;
  assign n601 = \new_[13771]_  ? \new_[7937]_  : \new_[2472]_ ;
  assign \new_[2472]_  = \\u0_slt3_r_reg[7] ;
  assign n606 = \new_[13506]_  ? \new_[7937]_  : \new_[2474]_ ;
  assign \new_[2474]_  = \\u0_slt3_r_reg[6] ;
  assign n611 = \new_[13548]_  ? \new_[7937]_  : \new_[2476]_ ;
  assign \new_[2476]_  = \\u0_slt3_r_reg[5] ;
  assign n616 = \new_[13562]_  ? \new_[7937]_  : \new_[2478]_ ;
  assign \new_[2478]_  = \\u0_slt3_r_reg[4] ;
  assign n621 = \new_[13280]_  ? \new_[7966]_  : \new_[2480]_ ;
  assign \new_[2480]_  = \\u0_slt3_r_reg[3] ;
  assign n626 = \new_[13647]_  ? \new_[7966]_  : \new_[2482]_ ;
  assign \new_[2482]_  = \\u0_slt3_r_reg[2] ;
  assign n631 = \new_[13529]_  ? \new_[7966]_  : \new_[2484]_ ;
  assign \new_[2484]_  = \\u0_slt3_r_reg[1] ;
  assign n636 = \new_[13525]_  ? \new_[7937]_  : \new_[2486]_ ;
  assign \new_[2486]_  = \\u0_slt3_r_reg[0] ;
  assign n641 = \new_[13471]_  ? \new_[7937]_  : \new_[2488]_ ;
  assign \new_[2488]_  = \\u0_slt4_r_reg[19] ;
  assign n646 = \new_[13260]_  ? \new_[7966]_  : \new_[2490]_ ;
  assign \new_[2490]_  = \\u0_slt4_r_reg[18] ;
  assign n651 = \new_[13392]_  ? \new_[8501]_  : \new_[2492]_ ;
  assign \new_[2492]_  = \\u0_slt4_r_reg[17] ;
  assign n656 = \new_[13210]_  ? \new_[8501]_  : \new_[2494]_ ;
  assign \new_[2494]_  = \\u0_slt4_r_reg[16] ;
  assign n661 = \new_[13477]_  ? \new_[7937]_  : \new_[2496]_ ;
  assign \new_[2496]_  = \\u0_slt4_r_reg[15] ;
  assign n666 = \new_[13486]_  ? \new_[7937]_  : \new_[2498]_ ;
  assign \new_[2498]_  = \\u0_slt4_r_reg[14] ;
  assign n671 = \new_[13743]_  ? \new_[8501]_  : \new_[2500]_ ;
  assign \new_[2500]_  = \\u0_slt4_r_reg[13] ;
  assign n676 = \new_[13338]_  ? \new_[7937]_  : \new_[2502]_ ;
  assign \new_[2502]_  = \\u0_slt4_r_reg[12] ;
  assign n681 = \new_[13335]_  ? \new_[8483]_  : \new_[2504]_ ;
  assign \new_[2504]_  = \\u0_slt4_r_reg[11] ;
  assign n686 = \new_[13352]_  ? \new_[7966]_  : \new_[2506]_ ;
  assign \new_[2506]_  = \\u0_slt4_r_reg[10] ;
  assign n691 = \new_[13353]_  ? \new_[8501]_  : \new_[2508]_ ;
  assign \new_[2508]_  = \\u0_slt4_r_reg[9] ;
  assign n696 = \new_[13214]_  ? \new_[7937]_  : \new_[2510]_ ;
  assign \new_[2510]_  = \\u0_slt4_r_reg[8] ;
  assign n701 = \new_[13219]_  ? \new_[7937]_  : \new_[2512]_ ;
  assign \new_[2512]_  = \\u0_slt4_r_reg[7] ;
  assign n706 = \new_[13275]_  ? \new_[8483]_  : \new_[2514]_ ;
  assign \new_[2514]_  = \\u0_slt4_r_reg[6] ;
  assign n711 = \new_[13251]_  ? \new_[7966]_  : \new_[2516]_ ;
  assign \new_[2516]_  = \\u0_slt4_r_reg[5] ;
  assign n716 = \new_[13235]_  ? \new_[8483]_  : \new_[2518]_ ;
  assign \new_[2518]_  = \\u0_slt4_r_reg[4] ;
  assign n721 = \new_[13247]_  ? \new_[7937]_  : \new_[2520]_ ;
  assign \new_[2520]_  = \\u0_slt4_r_reg[3] ;
  assign n726 = \new_[13661]_  ? \new_[7966]_  : \new_[2522]_ ;
  assign \new_[2522]_  = \\u0_slt4_r_reg[2] ;
  assign n731 = \new_[13201]_  ? \new_[8501]_  : \new_[2524]_ ;
  assign \new_[2524]_  = \\u0_slt4_r_reg[1] ;
  assign n736 = \new_[13334]_  ? \new_[8483]_  : \new_[2526]_ ;
  assign \new_[2526]_  = \\u0_slt4_r_reg[0] ;
  assign n741 = \new_[13209]_  ? \new_[8483]_  : \new_[2528]_ ;
  assign \new_[2528]_  = \\u0_slt5_r_reg[19] ;
  assign n746 = \new_[2530]_  & \new_[7962]_ ;
  assign \new_[2530]_  = \\u0_slt5_r_reg[18] ;
  assign n751 = \new_[2532]_  & \new_[7962]_ ;
  assign \new_[2532]_  = \\u0_slt5_r_reg[17] ;
  assign n756 = \new_[2534]_  & \new_[7962]_ ;
  assign \new_[2534]_  = \\u0_slt5_r_reg[16] ;
  assign n761 = \new_[2536]_  & \new_[7962]_ ;
  assign \new_[2536]_  = \\u0_slt5_r_reg[15] ;
  assign n766 = \new_[2538]_  & \new_[7962]_ ;
  assign \new_[2538]_  = \\u0_slt5_r_reg[14] ;
  assign n771 = \new_[2540]_  & \new_[7962]_ ;
  assign \new_[2540]_  = \\u0_slt5_r_reg[13] ;
  assign n776 = \new_[2542]_  & \new_[7962]_ ;
  assign \new_[2542]_  = \\u0_slt5_r_reg[12] ;
  assign n781 = \new_[2544]_  & \new_[7962]_ ;
  assign \new_[2544]_  = \\u0_slt5_r_reg[11] ;
  assign n786 = \new_[2546]_  & \new_[7962]_ ;
  assign \new_[2546]_  = \\u0_slt5_r_reg[10] ;
  assign n791 = \new_[2548]_  & \new_[7962]_ ;
  assign \new_[2548]_  = \\u0_slt5_r_reg[9] ;
  assign n796 = \new_[2550]_  & \new_[7962]_ ;
  assign \new_[2550]_  = \\u0_slt5_r_reg[8] ;
  assign n801 = \new_[2552]_  & \new_[8483]_ ;
  assign \new_[2552]_  = \\u0_slt5_r_reg[7] ;
  assign n806 = \new_[2554]_  & \new_[8483]_ ;
  assign \new_[2554]_  = \\u0_slt5_r_reg[6] ;
  assign n811 = \new_[2556]_  & \new_[7962]_ ;
  assign \new_[2556]_  = \\u0_slt5_r_reg[5] ;
  assign n816 = \new_[2558]_  & \new_[7962]_ ;
  assign \new_[2558]_  = \\u0_slt5_r_reg[4] ;
  assign n821 = \new_[2560]_  & \new_[7962]_ ;
  assign \new_[2560]_  = \\u0_slt5_r_reg[3] ;
  assign n826 = \new_[2562]_  & \new_[7962]_ ;
  assign \new_[2562]_  = \\u0_slt5_r_reg[2] ;
  assign n831 = \new_[2564]_  & \new_[7962]_ ;
  assign \new_[2564]_  = \\u0_slt5_r_reg[1] ;
  assign n836 = \new_[2566]_  & \new_[7962]_ ;
  assign \new_[2566]_  = \\u0_slt5_r_reg[0] ;
  assign n841 = \new_[2568]_  & \new_[7962]_ ;
  assign \new_[2568]_  = \\u0_slt6_r_reg[19] ;
  assign n846 = \new_[13744]_  ? \new_[7937]_  : \new_[2570]_ ;
  assign \new_[2570]_  = \\u0_slt6_r_reg[18] ;
  assign n851 = \new_[13721]_  ? \new_[7966]_  : \new_[2572]_ ;
  assign \new_[2572]_  = \\u0_slt6_r_reg[17] ;
  assign n856 = \new_[13728]_  ? \new_[7937]_  : \new_[2574]_ ;
  assign \new_[2574]_  = \\u0_slt6_r_reg[16] ;
  assign n861 = \new_[13729]_  ? \new_[7937]_  : \new_[2576]_ ;
  assign \new_[2576]_  = \\u0_slt6_r_reg[15] ;
  assign n866 = \new_[13749]_  ? \new_[7966]_  : \new_[2578]_ ;
  assign \new_[2578]_  = \\u0_slt6_r_reg[14] ;
  assign n871 = \new_[13454]_  ? \new_[8483]_  : \new_[2580]_ ;
  assign \new_[2580]_  = \\u0_slt6_r_reg[13] ;
  assign n876 = \new_[13387]_  ? \new_[7937]_  : \new_[2582]_ ;
  assign \new_[2582]_  = \\u0_slt6_r_reg[12] ;
  assign n881 = \new_[13770]_  ? \new_[7937]_  : \new_[2584]_ ;
  assign \new_[2584]_  = \\u0_slt6_r_reg[11] ;
  assign n886 = \new_[13404]_  ? \new_[7966]_  : \new_[2586]_ ;
  assign \new_[2586]_  = \\u0_slt6_r_reg[10] ;
  assign n891 = \new_[13399]_  ? \new_[7937]_  : \new_[2588]_ ;
  assign \new_[2588]_  = \\u0_slt6_r_reg[9] ;
  assign n896 = \new_[13447]_  ? \new_[8501]_  : \new_[2590]_ ;
  assign \new_[2590]_  = \\u0_slt6_r_reg[8] ;
  assign n901 = \new_[13444]_  ? \new_[7937]_  : \new_[2592]_ ;
  assign \new_[2592]_  = \\u0_slt6_r_reg[7] ;
  assign n906 = \new_[13643]_  ? \new_[8501]_  : \new_[2594]_ ;
  assign \new_[2594]_  = \\u0_slt6_r_reg[6] ;
  assign n911 = \new_[13496]_  ? \new_[7937]_  : \new_[2596]_ ;
  assign \new_[2596]_  = \\u0_slt6_r_reg[5] ;
  assign n916 = \new_[13451]_  ? \new_[7937]_  : \new_[2598]_ ;
  assign \new_[2598]_  = \\u0_slt6_r_reg[4] ;
  assign n921 = \new_[13383]_  ? \new_[7966]_  : \new_[2600]_ ;
  assign \new_[2600]_  = \\u0_slt6_r_reg[3] ;
  assign n926 = \new_[13405]_  ? \new_[7966]_  : \new_[2602]_ ;
  assign \new_[2602]_  = \\u0_slt6_r_reg[2] ;
  assign n931 = \new_[13433]_  ? \new_[7937]_  : \new_[2604]_ ;
  assign \new_[2604]_  = \\u0_slt6_r_reg[1] ;
  assign n936 = \new_[13850]_  ? \new_[7937]_  : \new_[2606]_ ;
  assign \new_[2606]_  = \\u0_slt6_r_reg[0] ;
  assign n941 = \new_[13515]_  ? \new_[7966]_  : \new_[2608]_ ;
  assign \new_[2608]_  = \\u0_slt7_r_reg[19] ;
  assign n946 = \new_[13388]_  ? \new_[7966]_  : \new_[2610]_ ;
  assign \new_[2610]_  = \\u0_slt7_r_reg[18] ;
  assign n951 = \new_[13206]_  ? \new_[7937]_  : \new_[2612]_ ;
  assign \new_[2612]_  = \\u0_slt7_r_reg[17] ;
  assign n956 = \new_[13648]_  ? \new_[7937]_  : \new_[2614]_ ;
  assign \new_[2614]_  = \\u0_slt7_r_reg[16] ;
  assign n961 = \new_[13469]_  ? \new_[7966]_  : \new_[2616]_ ;
  assign \new_[2616]_  = \\u0_slt7_r_reg[15] ;
  assign n966 = \new_[13697]_  ? \new_[7966]_  : \new_[2618]_ ;
  assign \new_[2618]_  = \\u0_slt7_r_reg[14] ;
  assign n971 = \new_[13595]_  ? \new_[7937]_  : \new_[2620]_ ;
  assign \new_[2620]_  = \\u0_slt7_r_reg[13] ;
  assign n976 = \new_[13462]_  ? \new_[7937]_  : \new_[2622]_ ;
  assign \new_[2622]_  = \\u0_slt7_r_reg[12] ;
  assign n981 = \new_[13198]_  ? \new_[7966]_  : \new_[2624]_ ;
  assign \new_[2624]_  = \\u0_slt7_r_reg[11] ;
  assign n986 = \new_[13507]_  ? \new_[7966]_  : \new_[2626]_ ;
  assign \new_[2626]_  = \\u0_slt7_r_reg[10] ;
  assign n991 = \new_[13225]_  ? \new_[7937]_  : \new_[2628]_ ;
  assign \new_[2628]_  = \\u0_slt7_r_reg[9] ;
  assign n996 = \new_[13244]_  ? \new_[7966]_  : \new_[2630]_ ;
  assign \new_[2630]_  = \\u0_slt7_r_reg[8] ;
  assign n1001 = \new_[13445]_  ? \new_[7937]_  : \new_[2632]_ ;
  assign \new_[2632]_  = \\u0_slt7_r_reg[7] ;
  assign n1006 = \new_[13255]_  ? \new_[7937]_  : \new_[2634]_ ;
  assign \new_[2634]_  = \\u0_slt7_r_reg[6] ;
  assign n1011 = \new_[13531]_  ? \new_[7937]_  : \new_[2636]_ ;
  assign \new_[2636]_  = \\u0_slt7_r_reg[5] ;
  assign n1016 = \new_[13561]_  ? \new_[8501]_  : \new_[2638]_ ;
  assign \new_[2638]_  = \\u0_slt7_r_reg[4] ;
  assign n1021 = \new_[13331]_  ? \new_[7966]_  : \new_[2640]_ ;
  assign \new_[2640]_  = \\u0_slt7_r_reg[3] ;
  assign n1026 = \new_[13745]_  ? \new_[7966]_  : \new_[2642]_ ;
  assign \new_[2642]_  = \\u0_slt7_r_reg[2] ;
  assign n1031 = \new_[13541]_  ? \new_[7962]_  : \new_[2644]_ ;
  assign \new_[2644]_  = \\u0_slt7_r_reg[1] ;
  assign n1036 = \new_[13846]_  ? \new_[7966]_  : \new_[2646]_ ;
  assign \new_[2646]_  = \\u0_slt7_r_reg[0] ;
  assign n1041 = \new_[13598]_  ? \new_[7937]_  : \new_[2648]_ ;
  assign \new_[2648]_  = \\u0_slt8_r_reg[19] ;
  assign n1046 = \new_[13343]_  ? \new_[7937]_  : \new_[2650]_ ;
  assign \new_[2650]_  = \\u0_slt8_r_reg[18] ;
  assign n1051 = \new_[13767]_  ? \new_[7962]_  : \new_[2652]_ ;
  assign \new_[2652]_  = \\u0_slt8_r_reg[17] ;
  assign n1056 = \new_[13492]_  ? \new_[8501]_  : \new_[2654]_ ;
  assign \new_[2654]_  = \\u0_slt8_r_reg[16] ;
  assign n1061 = \new_[13775]_  ? \new_[7937]_  : \new_[2656]_ ;
  assign \new_[2656]_  = \\u0_slt8_r_reg[15] ;
  assign n1066 = \new_[13493]_  ? \new_[7962]_  : \new_[2658]_ ;
  assign \new_[2658]_  = \\u0_slt8_r_reg[14] ;
  assign n1071 = \new_[13508]_  ? \new_[7937]_  : \new_[2660]_ ;
  assign \new_[2660]_  = \\u0_slt8_r_reg[13] ;
  assign n1076 = \new_[13780]_  ? \new_[8501]_  : \new_[2662]_ ;
  assign \new_[2662]_  = \\u0_slt8_r_reg[12] ;
  assign n1081 = \new_[13547]_  ? \new_[7937]_  : \new_[2664]_ ;
  assign \new_[2664]_  = \\u0_slt8_r_reg[11] ;
  assign n1086 = \new_[13608]_  ? \new_[7937]_  : \new_[2666]_ ;
  assign \new_[2666]_  = \\u0_slt8_r_reg[10] ;
  assign n1091 = \new_[13642]_  ? \new_[7966]_  : \new_[2668]_ ;
  assign \new_[2668]_  = \\u0_slt8_r_reg[9] ;
  assign n1096 = \new_[13230]_  ? \new_[7937]_  : \new_[2670]_ ;
  assign \new_[2670]_  = \\u0_slt8_r_reg[8] ;
  assign n1101 = \new_[13243]_  ? \new_[7966]_  : \new_[2672]_ ;
  assign \new_[2672]_  = \\u0_slt8_r_reg[7] ;
  assign n1106 = \new_[13259]_  ? \new_[7937]_  : \new_[2674]_ ;
  assign \new_[2674]_  = \\u0_slt8_r_reg[6] ;
  assign n1111 = \new_[13272]_  ? \new_[7966]_  : \new_[2676]_ ;
  assign \new_[2676]_  = \\u0_slt8_r_reg[5] ;
  assign n1116 = \new_[13416]_  ? \new_[7966]_  : \new_[2678]_ ;
  assign \new_[2678]_  = \\u0_slt8_r_reg[4] ;
  assign n1121 = \new_[13602]_  ? \new_[7966]_  : \new_[2680]_ ;
  assign \new_[2680]_  = \\u0_slt8_r_reg[3] ;
  assign n1126 = \new_[13739]_  ? \new_[7937]_  : \new_[2682]_ ;
  assign \new_[2682]_  = \\u0_slt8_r_reg[2] ;
  assign n1131 = \new_[13317]_  ? \new_[7937]_  : \new_[2684]_ ;
  assign \new_[2684]_  = \\u0_slt8_r_reg[1] ;
  assign n1136 = \new_[13812]_  ? \new_[7966]_  : \new_[2686]_ ;
  assign \new_[2686]_  = \\u0_slt8_r_reg[0] ;
  assign n1141 = \new_[13428]_  ? \new_[7966]_  : \new_[2688]_ ;
  assign \new_[2688]_  = \\u0_slt9_r_reg[19] ;
  assign n1146 = \new_[13231]_  ? \new_[7937]_  : \new_[2690]_ ;
  assign \new_[2690]_  = \\u0_slt9_r_reg[18] ;
  assign n1151 = \new_[13853]_  ? \new_[7937]_  : \new_[2692]_ ;
  assign \new_[2692]_  = \\u0_slt9_r_reg[17] ;
  assign n1156 = \new_[13669]_  ? \new_[8483]_  : \new_[2694]_ ;
  assign \new_[2694]_  = \\u0_slt9_r_reg[16] ;
  assign n1161 = \new_[13552]_  ? \new_[7962]_  : \new_[2696]_ ;
  assign \new_[2696]_  = \\u0_slt9_r_reg[15] ;
  assign n1166 = \new_[13391]_  ? \new_[7937]_  : \new_[2698]_ ;
  assign \new_[2698]_  = \\u0_slt9_r_reg[14] ;
  assign n1171 = \new_[13449]_  ? \new_[7966]_  : \new_[2700]_ ;
  assign \new_[2700]_  = \\u0_slt9_r_reg[13] ;
  assign n1176 = \new_[13559]_  ? \new_[7966]_  : \new_[2702]_ ;
  assign \new_[2702]_  = \\u0_slt9_r_reg[12] ;
  assign n1181 = \new_[13665]_  ? \new_[8483]_  : \new_[2704]_ ;
  assign \new_[2704]_  = \\u0_slt9_r_reg[11] ;
  assign n1186 = \new_[13385]_  ? \new_[8501]_  : \new_[2706]_ ;
  assign \new_[2706]_  = \\u0_slt9_r_reg[10] ;
  assign n1191 = \new_[13377]_  ? \new_[8501]_  : \new_[2708]_ ;
  assign \new_[2708]_  = \\u0_slt9_r_reg[9] ;
  assign n1196 = \new_[13599]_  ? \new_[7966]_  : \new_[2710]_ ;
  assign \new_[2710]_  = \\u0_slt9_r_reg[8] ;
  assign n1201 = \new_[13651]_  ? \new_[7966]_  : \new_[2712]_ ;
  assign \new_[2712]_  = \\u0_slt9_r_reg[7] ;
  assign n1206 = \new_[13585]_  ? \new_[8501]_  : \new_[2714]_ ;
  assign \new_[2714]_  = \\u0_slt9_r_reg[6] ;
  assign \new_[2715]_  = \\u1_slt2_reg[19] ;
  assign \new_[2716]_  = \\u1_slt3_reg[19] ;
  assign \new_[2717]_  = \\u1_slt4_reg[19] ;
  assign \new_[2718]_  = \\u1_slt6_reg[19] ;
  assign n1211 = \new_[13249]_  ? \new_[8501]_  : \new_[2730]_ ;
  assign n1216 = \new_[2745]_  ? \new_[8996]_  : \new_[2715]_ ;
  assign n1221 = \new_[2745]_  ? \new_[9002]_  : \new_[2716]_ ;
  assign n1226 = \new_[2745]_  ? \new_[9000]_  : \new_[2717]_ ;
  assign n1231 = \new_[2745]_  ? \new_[9001]_  : \new_[2718]_ ;
  assign \new_[2724]_  = \\u1_slt2_reg[18] ;
  assign \new_[2725]_  = \\u1_slt3_reg[18] ;
  assign \new_[2726]_  = \\u1_slt4_reg[18] ;
  assign \new_[2727]_  = \\u1_slt6_reg[18] ;
  assign \dma_req_o[1]  = u16_u1_dma_req_reg;
  assign \dma_req_o[3]  = u16_u3_dma_req_reg;
  assign \new_[2730]_  = \\u0_slt9_r_reg[5] ;
  assign \dma_req_o[0]  = u16_u0_dma_req_reg;
  assign \dma_req_o[2]  = u16_u2_dma_req_reg;
  assign \dma_req_o[4]  = u16_u4_dma_req_reg;
  assign \dma_req_o[5]  = u16_u5_dma_req_reg;
  assign \new_[2735]_  = \\u1_slt2_reg[17] ;
  assign \new_[2736]_  = \\u1_slt3_reg[17] ;
  assign \new_[2737]_  = \\u1_slt4_reg[17] ;
  assign \new_[2738]_  = \\u1_slt6_reg[17] ;
  assign n1236 = n1311 ? \new_[8996]_  : \new_[2724]_ ;
  assign n1241 = n1311 ? \new_[9002]_  : \new_[2725]_ ;
  assign n1246 = n1311 ? \new_[9000]_  : \new_[2726]_ ;
  assign n1251 = n1311 ? \new_[9001]_  : \new_[2727]_ ;
  assign n1256 = ~\new_[2773]_  | (~\dma_ack_i[1]  & ~\new_[13421]_ );
  assign n1261 = ~\new_[2774]_  | (~\dma_ack_i[3]  & ~\new_[13720]_ );
  assign \new_[2745]_  = \\u1_sr_reg[19] ;
  assign \new_[2746]_  = \\u1_slt2_reg[16] ;
  assign \new_[2747]_  = \\u1_slt3_reg[16] ;
  assign \new_[2748]_  = \\u1_slt4_reg[16] ;
  assign \new_[2749]_  = \\u1_slt6_reg[16] ;
  assign \new_[2750]_  = \\u4_rp_reg[2] ;
  assign \new_[2751]_  = \\u5_rp_reg[2] ;
  assign \new_[2752]_  = \\u8_rp_reg[2] ;
  assign \new_[2753]_  = \\u3_rp_reg[2] ;
  assign \new_[2754]_  = \\u6_rp_reg[2] ;
  assign \new_[2755]_  = \\u7_rp_reg[2] ;
  assign \new_[2756]_  = \\u8_rp_reg[3] ;
  assign \new_[2757]_  = \\u3_rp_reg[3] ;
  assign \new_[2758]_  = \\u6_rp_reg[3] ;
  assign \new_[2759]_  = \\u7_rp_reg[3] ;
  assign n1271 = ~\new_[2802]_  | (~\dma_ack_i[0]  & ~\new_[13434]_ );
  assign n1276 = ~\new_[2803]_  | (~\dma_ack_i[2]  & ~\new_[13740]_ );
  assign n1281 = ~\new_[2804]_  | (~\dma_ack_i[4]  & ~\new_[13441]_ );
  assign n1286 = ~\new_[2805]_  | (~\dma_ack_i[5]  & ~\new_[13407]_ );
  assign n1266 = \new_[13264]_  ? \new_[7937]_  : \new_[2896]_ ;
  assign n1291 = n1406 ? \new_[8996]_  : \new_[2735]_ ;
  assign n1296 = n1406 ? \new_[9002]_  : \new_[2736]_ ;
  assign n1301 = n1406 ? \new_[9000]_  : \new_[2737]_ ;
  assign n1306 = n1406 ? \new_[9001]_  : \new_[2738]_ ;
  assign \new_[2769]_  = \\u8_rp_reg[1] ;
  assign \new_[2770]_  = \\u3_rp_reg[1] ;
  assign \new_[2771]_  = \\u7_rp_reg[1] ;
  assign \new_[2772]_  = \\u6_rp_reg[1] ;
  assign \new_[2773]_  = ~n1911 | ~\new_[2897]_ ;
  assign \new_[2774]_  = ~n1916 | ~\new_[2898]_ ;
  assign n1311 = \\u1_sr_reg[18] ;
  assign n1346 = ~\new_[14093]_  & ~\new_[2910]_ ;
  assign n1351 = ~\new_[2911]_  & ~\new_[12811]_ ;
  assign n1356 = ~\new_[12042]_  & ~\new_[2912]_ ;
  assign n1361 = ~\new_[13168]_  & ~\new_[2913]_ ;
  assign n1371 = ~\new_[12039]_  & ~\new_[2914]_ ;
  assign n1376 = ~\new_[12042]_  & ~\new_[2917]_ ;
  assign n1381 = ~\new_[12409]_  & ~\new_[2920]_ ;
  assign \new_[2783]_  = \\u13_ints_r_reg[11] ;
  assign \new_[2784]_  = \\u13_ints_r_reg[5] ;
  assign \new_[2785]_  = \\u1_slt3_reg[15] ;
  assign \new_[2786]_  = \\u1_slt0_reg[15] ;
  assign \new_[2787]_  = \\u1_slt6_reg[15] ;
  assign \new_[2788]_  = \\u1_slt2_reg[15] ;
  assign \new_[2789]_  = \\u1_slt4_reg[15] ;
  assign \new_[2790]_  = \\u4_rp_reg[1] ;
  assign \new_[2791]_  = \\u4_rp_reg[3] ;
  assign \new_[2792]_  = \\u5_rp_reg[1] ;
  assign \new_[2793]_  = \\u5_rp_reg[3] ;
  assign \new_[2794]_  = ~\\u6_dout_reg[2] ;
  assign \new_[2795]_  = ~\\u6_dout_reg[3] ;
  assign \new_[2796]_  = ~\\u7_dout_reg[2] ;
  assign \new_[2797]_  = ~\\u7_dout_reg[3] ;
  assign \new_[2798]_  = ~\\u3_dout_reg[2] ;
  assign \new_[2799]_  = ~\\u3_dout_reg[3] ;
  assign \new_[2800]_  = ~\\u8_dout_reg[2] ;
  assign \new_[2801]_  = ~\\u8_dout_reg[3] ;
  assign \new_[2802]_  = ~n1971 | ~\new_[2930]_ ;
  assign \new_[2803]_  = ~n1976 | ~\new_[2931]_ ;
  assign \new_[2804]_  = ~n1981 | ~\new_[2932]_ ;
  assign \new_[2805]_  = ~n1986 | ~\new_[2933]_ ;
  assign n1316 = n1921 ? \new_[8996]_  : \new_[2746]_ ;
  assign n1321 = n1921 ? \new_[9002]_  : \new_[2747]_ ;
  assign n1326 = n1921 ? \new_[9000]_  : \new_[2748]_ ;
  assign n1331 = n1921 ? \new_[9001]_  : \new_[2749]_ ;
  assign n1336 = \new_[2904]_  & \new_[12886]_ ;
  assign n1341 = \new_[2905]_  & \new_[12691]_ ;
  assign n1386 = ~\new_[14093]_  & (~\new_[3143]_  | ~\new_[4006]_ );
  assign n1391 = ~\new_[12811]_  & (~\new_[4007]_  | ~\new_[3144]_ );
  assign n1401 = ~\new_[12042]_  & (~\new_[3146]_  | ~\new_[4008]_ );
  assign n1396 = ~\new_[12409]_  & (~\new_[3147]_  | ~\new_[4009]_ );
  assign \new_[2816]_  = \\u13_ints_r_reg[14] ;
  assign \new_[2817]_  = \\u13_ints_r_reg[17] ;
  assign \new_[2818]_  = \\u13_ints_r_reg[2] ;
  assign \new_[2819]_  = \\u13_ints_r_reg[8] ;
  assign \new_[2820]_  = ~\\u6_dout_reg[0] ;
  assign \new_[2821]_  = ~\\u6_dout_reg[1] ;
  assign \new_[2822]_  = ~\\u7_dout_reg[0] ;
  assign \new_[2823]_  = ~\\u7_dout_reg[1] ;
  assign \new_[2824]_  = ~\\u3_dout_reg[0] ;
  assign \new_[2825]_  = ~\\u8_dout_reg[0] ;
  assign \new_[2826]_  = ~\\u3_dout_reg[1] ;
  assign \new_[2827]_  = ~\\u8_dout_reg[1] ;
  assign \new_[2828]_  = \\u8_rp_reg[0] ;
  assign \new_[2829]_  = \\u3_rp_reg[0] ;
  assign \new_[2830]_  = \\u6_rp_reg[0] ;
  assign \new_[2831]_  = \\u7_rp_reg[0] ;
  assign \new_[2832]_  = ~\\u6_dout_reg[12] ;
  assign \new_[2833]_  = ~\\u6_dout_reg[13] ;
  assign \new_[2834]_  = ~\\u6_dout_reg[14] ;
  assign \new_[2835]_  = ~\\u6_dout_reg[15] ;
  assign \new_[2836]_  = ~\\u6_dout_reg[10] ;
  assign \new_[2837]_  = ~\\u6_dout_reg[11] ;
  assign \new_[2838]_  = ~\\u6_dout_reg[18] ;
  assign \new_[2839]_  = ~\\u6_dout_reg[19] ;
  assign \new_[2840]_  = ~\\u6_dout_reg[16] ;
  assign \new_[2841]_  = ~\\u6_dout_reg[17] ;
  assign \new_[2842]_  = ~\\u6_dout_reg[4] ;
  assign \new_[2843]_  = ~\\u6_dout_reg[5] ;
  assign \new_[2844]_  = ~\\u6_dout_reg[6] ;
  assign \new_[2845]_  = ~\\u6_dout_reg[7] ;
  assign \new_[2846]_  = ~\\u6_dout_reg[8] ;
  assign \new_[2847]_  = ~\\u6_dout_reg[9] ;
  assign \new_[2848]_  = ~\\u7_dout_reg[10] ;
  assign \new_[2849]_  = ~\\u7_dout_reg[11] ;
  assign \new_[2850]_  = ~\\u7_dout_reg[12] ;
  assign \new_[2851]_  = ~\\u7_dout_reg[13] ;
  assign \new_[2852]_  = ~\\u7_dout_reg[14] ;
  assign \new_[2853]_  = ~\\u7_dout_reg[17] ;
  assign \new_[2854]_  = ~\\u7_dout_reg[15] ;
  assign \new_[2855]_  = ~\\u7_dout_reg[19] ;
  assign \new_[2856]_  = ~\\u7_dout_reg[16] ;
  assign \new_[2857]_  = ~\\u7_dout_reg[18] ;
  assign \new_[2858]_  = ~\\u7_dout_reg[4] ;
  assign \new_[2859]_  = ~\\u7_dout_reg[5] ;
  assign \new_[2860]_  = ~\\u7_dout_reg[6] ;
  assign \new_[2861]_  = ~\\u7_dout_reg[7] ;
  assign \new_[2862]_  = ~\\u7_dout_reg[8] ;
  assign \new_[2863]_  = ~\\u7_dout_reg[9] ;
  assign \new_[2864]_  = ~\\u3_dout_reg[10] ;
  assign \new_[2865]_  = ~\\u3_dout_reg[11] ;
  assign \new_[2866]_  = ~\\u3_dout_reg[13] ;
  assign \new_[2867]_  = ~\\u3_dout_reg[14] ;
  assign \new_[2868]_  = ~\\u3_dout_reg[15] ;
  assign \new_[2869]_  = ~\\u3_dout_reg[16] ;
  assign \new_[2870]_  = ~\\u3_dout_reg[17] ;
  assign \new_[2871]_  = ~\\u3_dout_reg[18] ;
  assign \new_[2872]_  = ~\\u8_dout_reg[10] ;
  assign \new_[2873]_  = ~\\u3_dout_reg[19] ;
  assign \new_[2874]_  = ~\\u8_dout_reg[11] ;
  assign \new_[2875]_  = ~\\u8_dout_reg[12] ;
  assign \new_[2876]_  = ~\\u3_dout_reg[12] ;
  assign \new_[2877]_  = ~\\u8_dout_reg[13] ;
  assign \new_[2878]_  = ~\\u8_dout_reg[14] ;
  assign \new_[2879]_  = ~\\u3_dout_reg[4] ;
  assign \new_[2880]_  = ~\\u8_dout_reg[16] ;
  assign \new_[2881]_  = ~\\u3_dout_reg[6] ;
  assign \new_[2882]_  = ~\\u8_dout_reg[17] ;
  assign \new_[2883]_  = ~\\u3_dout_reg[7] ;
  assign \new_[2884]_  = ~\\u8_dout_reg[18] ;
  assign \new_[2885]_  = ~\\u3_dout_reg[8] ;
  assign \new_[2886]_  = ~\\u8_dout_reg[15] ;
  assign \new_[2887]_  = ~\\u3_dout_reg[5] ;
  assign \new_[2888]_  = ~\\u8_dout_reg[19] ;
  assign \new_[2889]_  = ~\\u3_dout_reg[9] ;
  assign \new_[2890]_  = ~\\u8_dout_reg[4] ;
  assign \new_[2891]_  = ~\\u8_dout_reg[5] ;
  assign \new_[2892]_  = ~\\u8_dout_reg[6] ;
  assign \new_[2893]_  = ~\\u8_dout_reg[7] ;
  assign \new_[2894]_  = ~\\u8_dout_reg[8] ;
  assign \new_[2895]_  = ~\\u8_dout_reg[9] ;
  assign \new_[2896]_  = \\u0_slt9_r_reg[4] ;
  assign \new_[2897]_  = u16_u1_dma_req_r1_reg;
  assign \new_[2898]_  = u16_u3_dma_req_r1_reg;
  assign n1406 = \\u1_sr_reg[17] ;
  assign n1451 = \new_[3177]_  & \new_[12886]_ ;
  assign n1461 = \new_[3178]_  & \new_[12691]_ ;
  assign n1446 = \new_[3181]_  & \new_[12886]_ ;
  assign n1456 = \new_[3182]_  & \new_[12691]_ ;
  assign \new_[2904]_  = ~\new_[3164]_  | (~\new_[9155]_  & ~\new_[4658]_ );
  assign \new_[2905]_  = ~\new_[3167]_  | (~\new_[9700]_  & ~\new_[4659]_ );
  assign n1466 = ~\new_[3165]_  & ~\new_[12074]_ ;
  assign n1471 = ~\new_[3166]_  & ~\new_[12074]_ ;
  assign n1476 = ~\new_[3168]_  & ~\new_[12409]_ ;
  assign n1481 = ~\new_[3169]_  & ~\new_[12409]_ ;
  assign \new_[2910]_  = ~\new_[3351]_  & (~\new_[9153]_  | ~\new_[14097]_ );
  assign \new_[2911]_  = ~\new_[3353]_  & (~\new_[9154]_  | ~\new_[4515]_ );
  assign \new_[2912]_  = ~\new_[3137]_  & (~\new_[8932]_  | ~\new_[4527]_ );
  assign \new_[2913]_  = ~\new_[3140]_  & (~\new_[9156]_  | ~\new_[4528]_ );
  assign \new_[2914]_  = ~\new_[3354]_  & (~\new_[9660]_  | ~\new_[4515]_ );
  assign n1486 = ~\new_[3170]_  & ~\new_[12811]_ ;
  assign n1491 = ~\new_[3171]_  & ~\new_[12811]_ ;
  assign \new_[2917]_  = ~\new_[3139]_  & (~\new_[9663]_  | ~\new_[4527]_ );
  assign n1496 = ~\new_[3172]_  & ~\new_[12402]_ ;
  assign n1501 = ~\new_[3173]_  & ~\new_[12402]_ ;
  assign \new_[2920]_  = ~\new_[3142]_  & (~\new_[10308]_  | ~\new_[4528]_ );
  assign \dma_req_o[8]  = u16_u8_dma_req_reg;
  assign \new_[2922]_  = \\u1_slt3_reg[14] ;
  assign \new_[2923]_  = \\u1_slt4_reg[14] ;
  assign \new_[2924]_  = \\u1_slt6_reg[14] ;
  assign \new_[2925]_  = \\u1_slt2_reg[14] ;
  assign \new_[2926]_  = ~\\u4_dout_reg[3] ;
  assign \new_[2927]_  = ~\\u5_dout_reg[3] ;
  assign \new_[2928]_  = ~\\u5_dout_reg[2] ;
  assign \new_[2929]_  = ~\\u4_dout_reg[2] ;
  assign \new_[2930]_  = u16_u0_dma_req_r1_reg;
  assign \new_[2931]_  = u16_u2_dma_req_r1_reg;
  assign \new_[2932]_  = u16_u4_dma_req_r1_reg;
  assign \new_[2933]_  = u16_u5_dma_req_r1_reg;
  assign n1411 = \new_[3342]_  & \new_[9077]_ ;
  assign n1416 = \new_[3343]_  & \new_[9077]_ ;
  assign n1426 = \new_[2786]_  ? \new_[9006]_  : n2546;
  assign n1436 = n2546 ? \new_[8996]_  : \new_[2788]_ ;
  assign n1421 = n2546 ? \new_[9002]_  : \new_[2785]_ ;
  assign n1441 = n2546 ? \new_[9000]_  : \new_[2789]_ ;
  assign n1431 = n2546 ? \new_[9001]_  : \new_[2787]_ ;
  assign n1576 = ~\new_[3644]_  & ~\new_[12074]_ ;
  assign n1581 = ~\new_[3645]_  & ~\new_[12409]_ ;
  assign n1526 = (~\new_[3658]_  & ~\new_[8876]_ ) | (~\new_[2820]_  & ~\new_[4144]_ );
  assign n1531 = (~\new_[3658]_  & ~\new_[8729]_ ) | (~\new_[4144]_  & ~\new_[2821]_ );
  assign n1536 = (~\new_[3662]_  & ~\new_[8736]_ ) | (~\new_[2822]_  & ~\new_[4151]_ );
  assign n1541 = (~\new_[3662]_  & ~\new_[8718]_ ) | (~\new_[4151]_  & ~\new_[2823]_ );
  assign n1546 = (~\new_[3665]_  & ~\new_[8745]_ ) | (~\new_[2824]_  & ~\new_[4157]_ );
  assign n1551 = (~\new_[3666]_  & ~\new_[8914]_ ) | (~\new_[2825]_  & ~\new_[4160]_ );
  assign \new_[2949]_  = ~\\u4_dout_reg[4] ;
  assign n1556 = (~\new_[3665]_  & ~\new_[8754]_ ) | (~\new_[4157]_  & ~\new_[2826]_ );
  assign n1561 = (~\new_[3666]_  & ~\new_[8760]_ ) | (~\new_[4160]_  & ~\new_[2827]_ );
  assign \new_[2952]_  = \\u11_wp_reg[3] ;
  assign n1606 = ~\new_[12074]_  & (~\new_[3895]_  | ~\new_[3800]_ );
  assign n1611 = ~\new_[12853]_  & (~\new_[3897]_  | ~\new_[3801]_ );
  assign n1586 = ~\new_[12042]_  & (~\new_[3898]_  | ~\new_[3802]_ );
  assign n1591 = ~\new_[12073]_  & (~\new_[3899]_  | ~\new_[3803]_ );
  assign n1596 = ~\new_[12073]_  & (~\new_[3901]_  | ~\new_[3804]_ );
  assign n1601 = ~\new_[12853]_  & (~\new_[3902]_  | ~\new_[3805]_ );
  assign n1626 = ~\new_[12074]_  & (~\new_[3903]_  | ~\new_[3806]_ );
  assign n1631 = ~\new_[12073]_  & (~\new_[3904]_  | ~\new_[3807]_ );
  assign n1616 = ~\new_[12073]_  & (~\new_[3809]_  | ~\new_[3905]_ );
  assign n1621 = ~\new_[12853]_  & (~\new_[3906]_  | ~\new_[3810]_ );
  assign n1636 = ~\new_[12073]_  & (~\new_[3908]_  | ~\new_[3813]_ );
  assign n1641 = ~\new_[12073]_  & (~\new_[3909]_  | ~\new_[3814]_ );
  assign n1646 = ~\new_[12073]_  & (~\new_[3910]_  | ~\new_[3815]_ );
  assign n1651 = ~\new_[12073]_  & (~\new_[3911]_  | ~\new_[3816]_ );
  assign n1656 = ~\new_[12853]_  & (~\new_[3912]_  | ~\new_[3817]_ );
  assign n1661 = ~\new_[12074]_  & (~\new_[3914]_  | ~\new_[3818]_ );
  assign n1666 = ~\new_[12458]_  & (~\new_[3819]_  | ~\new_[4181]_ );
  assign n1671 = ~\new_[13168]_  & (~\new_[3820]_  | ~\new_[4182]_ );
  assign n1676 = ~\new_[12409]_  & (~\new_[3821]_  | ~\new_[4183]_ );
  assign n1681 = ~\new_[13168]_  & (~\new_[3822]_  | ~\new_[4185]_ );
  assign n1686 = ~\new_[12458]_  & (~\new_[3823]_  | ~\new_[4186]_ );
  assign n1696 = ~\new_[12409]_  & (~\new_[3824]_  | ~\new_[4187]_ );
  assign n1706 = ~\new_[12322]_  & (~\new_[3825]_  | ~\new_[4188]_ );
  assign n1691 = ~\new_[13168]_  & (~\new_[3826]_  | ~\new_[4189]_ );
  assign n1711 = ~\new_[12409]_  & (~\new_[3827]_  | ~\new_[4190]_ );
  assign n1701 = ~\new_[12409]_  & (~\new_[3828]_  | ~\new_[4192]_ );
  assign n1716 = ~\new_[12458]_  & (~\new_[13938]_  | ~\new_[3831]_ );
  assign n1721 = ~\new_[12458]_  & (~\new_[13957]_  | ~\new_[3832]_ );
  assign n1726 = ~\new_[12322]_  & (~\new_[4194]_  | ~\new_[3833]_ );
  assign n1731 = ~\new_[12322]_  & (~\new_[3834]_  | ~\new_[14055]_ );
  assign n1736 = ~\new_[12322]_  & (~\new_[4196]_  | ~\new_[3835]_ );
  assign n1741 = ~\new_[13168]_  & (~\new_[3836]_  | ~\new_[4197]_ );
  assign n1746 = ~\new_[12811]_  & (~\new_[3915]_  | ~\new_[3837]_ );
  assign n1751 = ~\new_[12811]_  & (~\new_[14082]_  | ~\new_[3838]_ );
  assign n1806 = ~\new_[12811]_  & (~\new_[3917]_  | ~\new_[3839]_ );
  assign n1756 = ~\new_[12811]_  & (~\new_[13914]_  | ~\new_[3840]_ );
  assign n1761 = ~\new_[12811]_  & (~\new_[3841]_  | ~\new_[3918]_ );
  assign n1766 = ~\new_[12811]_  & (~\new_[3843]_  | ~\new_[14156]_ );
  assign n1771 = ~\new_[12811]_  & (~\new_[3844]_  | ~\new_[14141]_ );
  assign n1776 = ~\new_[12039]_  & (~\new_[14043]_  | ~\new_[3845]_ );
  assign n1781 = ~\new_[12039]_  & (~\new_[3846]_  | ~\new_[3921]_ );
  assign n1786 = ~\new_[12403]_  & (~\new_[3922]_  | ~\new_[3847]_ );
  assign n1791 = ~\new_[12811]_  & (~\new_[3848]_  | ~\new_[3924]_ );
  assign n1796 = ~\new_[12330]_  & (~\new_[3925]_  | ~\new_[3849]_ );
  assign n1801 = ~\new_[14093]_  & (~\new_[3926]_  | ~\new_[3850]_ );
  assign n1811 = ~\new_[12329]_  & (~\new_[3928]_  | ~\new_[3852]_ );
  assign n1816 = ~\new_[12329]_  & (~\new_[3929]_  | ~\new_[3854]_ );
  assign n1821 = ~\new_[12811]_  & (~\new_[3930]_  | ~\new_[3855]_ );
  assign n1856 = ~\new_[12330]_  & (~\new_[3931]_  | ~\new_[3856]_ );
  assign n1861 = ~\new_[12811]_  & (~\new_[3932]_  | ~\new_[3857]_ );
  assign n1826 = ~\new_[12403]_  & (~\new_[3933]_  | ~\new_[3858]_ );
  assign n1836 = ~\new_[12404]_  & (~\new_[3934]_  | ~\new_[3859]_ );
  assign n1831 = ~\new_[12039]_  & (~\new_[3935]_  | ~\new_[3860]_ );
  assign n1841 = ~\new_[12039]_  & (~\new_[3936]_  | ~\new_[3808]_ );
  assign n1846 = ~\new_[12404]_  & (~\new_[3938]_  | ~\new_[3861]_ );
  assign n1851 = ~\new_[12811]_  & (~\new_[3939]_  | ~\new_[3862]_ );
  assign n1866 = ~\new_[12330]_  & (~\new_[3940]_  | ~\new_[3863]_ );
  assign n1871 = ~\new_[12811]_  & (~\new_[3942]_  | ~\new_[3864]_ );
  assign n1876 = ~\new_[12329]_  & (~\new_[3943]_  | ~\new_[3867]_ );
  assign n1881 = ~\new_[12329]_  & (~\new_[3944]_  | ~\new_[3868]_ );
  assign n1886 = ~\new_[12404]_  & (~\new_[3946]_  | ~\new_[3869]_ );
  assign n1891 = ~\new_[12404]_  & (~\new_[3947]_  | ~\new_[3870]_ );
  assign n1896 = ~\new_[12330]_  & (~\new_[3948]_  | ~\new_[3798]_ );
  assign n1901 = ~\new_[12403]_  & (~\new_[3950]_  | ~\new_[3871]_ );
  assign \dma_req_o[6]  = u16_u6_dma_req_reg;
  assign \dma_req_o[7]  = u16_u7_dma_req_reg;
  assign \new_[3019]_  = ~\\u5_dout_reg[0] ;
  assign \new_[3020]_  = ~\\u5_dout_reg[1] ;
  assign \new_[3021]_  = ~\\u4_dout_reg[1] ;
  assign \new_[3022]_  = ~\\u4_dout_reg[0] ;
  assign \new_[3023]_  = \\u4_rp_reg[0] ;
  assign \new_[3024]_  = \\u5_rp_reg[0] ;
  assign \new_[3025]_  = ~\\u11_mem_reg[0][18] ;
  assign \new_[3026]_  = ~\\u11_mem_reg[0][19] ;
  assign \new_[3027]_  = ~\\u11_mem_reg[1][18] ;
  assign \new_[3028]_  = ~\\u11_mem_reg[1][19] ;
  assign \new_[3029]_  = ~\\u11_mem_reg[1][20] ;
  assign \new_[3030]_  = ~\\u11_mem_reg[1][21] ;
  assign \new_[3031]_  = ~\\u11_mem_reg[1][22] ;
  assign \new_[3032]_  = ~\\u11_mem_reg[1][23] ;
  assign \new_[3033]_  = ~\\u11_mem_reg[1][24] ;
  assign \new_[3034]_  = ~\\u11_mem_reg[1][25] ;
  assign \new_[3035]_  = ~\\u11_mem_reg[1][26] ;
  assign \new_[3036]_  = ~\\u11_mem_reg[1][27] ;
  assign \new_[3037]_  = ~\\u11_mem_reg[1][28] ;
  assign \new_[3038]_  = ~\\u11_mem_reg[1][29] ;
  assign \new_[3039]_  = ~\\u11_mem_reg[1][30] ;
  assign \new_[3040]_  = ~\\u11_mem_reg[1][31] ;
  assign \new_[3041]_  = ~\\u11_mem_reg[2][18] ;
  assign \new_[3042]_  = ~\\u11_mem_reg[2][19] ;
  assign \new_[3043]_  = ~\\u11_mem_reg[2][20] ;
  assign \new_[3044]_  = ~\\u11_mem_reg[2][21] ;
  assign \new_[3045]_  = ~\\u11_mem_reg[2][22] ;
  assign \new_[3046]_  = ~\\u11_mem_reg[2][23] ;
  assign \new_[3047]_  = ~\\u11_mem_reg[2][24] ;
  assign \new_[3048]_  = ~\\u11_mem_reg[2][25] ;
  assign \new_[3049]_  = ~\\u11_mem_reg[2][26] ;
  assign \new_[3050]_  = ~\\u11_mem_reg[2][27] ;
  assign \new_[3051]_  = ~\\u11_mem_reg[2][28] ;
  assign \new_[3052]_  = ~\\u11_mem_reg[2][29] ;
  assign \new_[3053]_  = ~\\u11_mem_reg[2][30] ;
  assign \new_[3054]_  = ~\\u11_mem_reg[2][31] ;
  assign \new_[3055]_  = ~\\u11_mem_reg[3][18] ;
  assign \new_[3056]_  = ~\\u11_mem_reg[3][19] ;
  assign \new_[3057]_  = ~\\u11_mem_reg[3][20] ;
  assign \new_[3058]_  = ~\\u11_mem_reg[3][21] ;
  assign \new_[3059]_  = ~\\u11_mem_reg[3][22] ;
  assign \new_[3060]_  = ~\\u11_mem_reg[3][23] ;
  assign \new_[3061]_  = ~\\u11_mem_reg[3][24] ;
  assign \new_[3062]_  = ~\\u11_mem_reg[3][25] ;
  assign \new_[3063]_  = ~\\u11_mem_reg[3][26] ;
  assign \new_[3064]_  = ~\\u11_mem_reg[3][27] ;
  assign \new_[3065]_  = ~\\u11_mem_reg[3][28] ;
  assign \new_[3066]_  = ~\\u11_mem_reg[3][29] ;
  assign \new_[3067]_  = ~\\u11_mem_reg[3][30] ;
  assign \new_[3068]_  = ~\\u11_mem_reg[3][31] ;
  assign \new_[3069]_  = ~\\u11_mem_reg[3][7] ;
  assign \new_[3070]_  = ~\\u11_mem_reg[1][12] ;
  assign \new_[3071]_  = ~\\u11_mem_reg[1][13] ;
  assign \new_[3072]_  = ~\\u11_mem_reg[1][16] ;
  assign \new_[3073]_  = ~\\u11_mem_reg[2][17] ;
  assign \new_[3074]_  = ~\\u11_mem_reg[2][1] ;
  assign \new_[3075]_  = ~\\u11_mem_reg[2][7] ;
  assign \new_[3076]_  = ~\\u11_mem_reg[2][8] ;
  assign \new_[3077]_  = ~\\u11_mem_reg[3][16] ;
  assign \new_[3078]_  = ~\\u11_mem_reg[3][17] ;
  assign \new_[3079]_  = ~\\u11_mem_reg[3][5] ;
  assign \new_[3080]_  = ~\\u11_mem_reg[3][6] ;
  assign \new_[3081]_  = \\u11_wp_reg[1] ;
  assign \new_[3082]_  = \\u11_wp_reg[2] ;
  assign \new_[3083]_  = ~\\u4_dout_reg[10] ;
  assign \new_[3084]_  = ~\\u4_dout_reg[13] ;
  assign \new_[3085]_  = ~\\u4_dout_reg[14] ;
  assign \new_[3086]_  = ~\\u4_dout_reg[15] ;
  assign \new_[3087]_  = ~\\u4_dout_reg[16] ;
  assign \new_[3088]_  = ~\\u4_dout_reg[11] ;
  assign \new_[3089]_  = ~\\u4_dout_reg[18] ;
  assign \new_[3090]_  = ~\\u4_dout_reg[12] ;
  assign \new_[3091]_  = ~\\u4_dout_reg[19] ;
  assign \new_[3092]_  = ~\\u4_dout_reg[17] ;
  assign \new_[3093]_  = ~\\u4_dout_reg[5] ;
  assign \new_[3094]_  = ~\\u4_dout_reg[6] ;
  assign \new_[3095]_  = ~\\u4_dout_reg[7] ;
  assign \new_[3096]_  = ~\\u4_dout_reg[8] ;
  assign \new_[3097]_  = ~\\u4_dout_reg[9] ;
  assign \new_[3098]_  = ~\\u5_dout_reg[10] ;
  assign \new_[3099]_  = ~\\u5_dout_reg[11] ;
  assign \new_[3100]_  = ~\\u5_dout_reg[12] ;
  assign \new_[3101]_  = ~\\u5_dout_reg[14] ;
  assign \new_[3102]_  = ~\\u5_dout_reg[15] ;
  assign \new_[3103]_  = ~\\u5_dout_reg[16] ;
  assign \new_[3104]_  = ~\\u5_dout_reg[18] ;
  assign \new_[3105]_  = ~\\u5_dout_reg[19] ;
  assign \new_[3106]_  = ~\\u5_dout_reg[4] ;
  assign \new_[3107]_  = ~\\u5_dout_reg[5] ;
  assign \new_[3108]_  = ~\\u5_dout_reg[6] ;
  assign \new_[3109]_  = ~\\u5_dout_reg[8] ;
  assign \new_[3110]_  = ~\\u5_dout_reg[9] ;
  assign \new_[3111]_  = ~\\u11_mem_reg[0][0] ;
  assign \new_[3112]_  = ~\\u11_mem_reg[0][10] ;
  assign \new_[3113]_  = ~\\u11_mem_reg[0][11] ;
  assign \new_[3114]_  = ~\\u11_mem_reg[0][12] ;
  assign \new_[3115]_  = ~\\u11_mem_reg[0][13] ;
  assign \new_[3116]_  = ~\\u11_mem_reg[0][14] ;
  assign \new_[3117]_  = ~\\u11_mem_reg[0][15] ;
  assign \new_[3118]_  = ~\\u11_mem_reg[0][1] ;
  assign \new_[3119]_  = u15_crac_rd_reg;
  assign \new_[3120]_  = ~\\u17_int_set_reg[1] ;
  assign \new_[3121]_  = ~\\u20_int_set_reg[1] ;
  assign \new_[3122]_  = ~\\u21_int_set_reg[1] ;
  assign \new_[3123]_  = ~\\u22_int_set_reg[1] ;
  assign n1506 = \new_[3627]_  & \new_[9077]_ ;
  assign n1511 = \new_[3628]_  & \new_[9077]_ ;
  assign n1516 = \new_[3629]_  & \new_[9077]_ ;
  assign n1521 = \new_[3630]_  & \new_[9077]_ ;
  assign \new_[3128]_  = ~\\u5_dout_reg[7] ;
  assign n1911 = ~\new_[3646]_  & ~\dma_ack_i[1] ;
  assign \new_[3130]_  = ~\\u5_dout_reg[17] ;
  assign n1916 = ~\new_[3647]_  & ~\dma_ack_i[3] ;
  assign n1906 = \new_[13350]_  ? \new_[7937]_  : \new_[3650]_ ;
  assign n1921 = \\u1_sr_reg[16] ;
  assign \new_[3134]_  = ~\\u5_dout_reg[13] ;
  assign n1566 = ~\new_[3634]_  & ~\new_[12402]_ ;
  assign n1571 = ~\new_[3635]_  & ~\new_[12811]_ ;
  assign \new_[3137]_  = ~\new_[3678]_  & ~\new_[4527]_ ;
  assign \new_[3138]_  = ~\\u10_mem_reg[0][18] ;
  assign \new_[3139]_  = ~\new_[3792]_  & ~\new_[4527]_ ;
  assign \new_[3140]_  = ~\new_[3679]_  & ~\new_[4528]_ ;
  assign \new_[3141]_  = ~\\u10_mem_reg[3][28] ;
  assign \new_[3142]_  = ~\new_[3793]_  & ~\new_[4528]_ ;
  assign \new_[3143]_  = \new_[3999]_  | \new_[14097]_ ;
  assign \new_[3144]_  = \new_[4000]_  | \new_[4515]_ ;
  assign \new_[3145]_  = ~\\u10_mem_reg[3][24] ;
  assign \new_[3146]_  = \new_[4001]_  | \new_[4527]_ ;
  assign \new_[3147]_  = \new_[4002]_  | \new_[4528]_ ;
  assign \new_[3148]_  = ~\\u9_mem_reg[3][30] ;
  assign \new_[3149]_  = ~\\u9_mem_reg[3][26] ;
  assign \new_[3150]_  = \\u10_wp_reg[3] ;
  assign \new_[3151]_  = ~\\u9_mem_reg[3][22] ;
  assign \new_[3152]_  = ~\\u9_mem_reg[2][28] ;
  assign \new_[3153]_  = ~\\u9_mem_reg[2][24] ;
  assign \new_[3154]_  = ~\\u9_mem_reg[2][20] ;
  assign n1966 = ~\new_[3667]_  & ~\new_[12040]_ ;
  assign n1951 = ~\new_[3668]_  & ~\new_[12040]_ ;
  assign \new_[3157]_  = ~\\u9_mem_reg[1][28] ;
  assign \new_[3158]_  = ~\\u9_mem_reg[1][25] ;
  assign \new_[3159]_  = ~\\u9_mem_reg[1][22] ;
  assign n1961 = ~\new_[3669]_  & ~\new_[11421]_ ;
  assign \new_[3161]_  = ~\\u10_mem_reg[2][24] ;
  assign n1956 = ~\new_[3670]_  & ~\new_[11421]_ ;
  assign \new_[3163]_  = ~\\u11_mem_reg[3][14] ;
  assign \new_[3164]_  = ~\new_[4066]_  | ~\new_[4658]_  | ~\new_[4358]_ ;
  assign \new_[3165]_  = ~\new_[3811]_  & (~\new_[13541]_  | ~\new_[4623]_ );
  assign \new_[3166]_  = ~\new_[3812]_  & (~\new_[13745]_  | ~\new_[4623]_ );
  assign \new_[3167]_  = ~\new_[4067]_  | ~\new_[4659]_  | ~\new_[4360]_ ;
  assign \new_[3168]_  = ~\new_[3829]_  & (~\new_[13317]_  | ~\new_[4476]_ );
  assign \new_[3169]_  = ~\new_[3830]_  & (~\new_[13739]_  | ~\new_[4476]_ );
  assign \new_[3170]_  = ~\new_[3851]_  & (~\new_[13529]_  | ~\new_[4472]_ );
  assign \new_[3171]_  = ~\new_[3853]_  & (~\new_[13647]_  | ~\new_[4472]_ );
  assign \new_[3172]_  = ~\new_[3865]_  & (~\new_[13369]_  | ~\new_[4624]_ );
  assign \new_[3173]_  = ~\new_[3866]_  & (~\new_[13361]_  | ~\new_[4624]_ );
  assign \new_[3174]_  = ~\\u11_mem_reg[3][0] ;
  assign \new_[3175]_  = ~\\u11_mem_reg[3][13] ;
  assign \new_[3176]_  = ~\\u10_mem_reg[1][0] ;
  assign \new_[3177]_  = \new_[8827]_  ? \new_[4658]_  : \new_[4088]_ ;
  assign \new_[3178]_  = \new_[9078]_  ? \new_[4659]_  : \new_[4089]_ ;
  assign \new_[3179]_  = ~\\u11_mem_reg[1][15] ;
  assign \new_[3180]_  = ~\\u11_mem_reg[1][6] ;
  assign \new_[3181]_  = \new_[12011]_  ? \new_[4658]_  : \new_[4277]_ ;
  assign \new_[3182]_  = \new_[12672]_  ? \new_[4659]_  : \new_[4278]_ ;
  assign \new_[3183]_  = \\u1_slt2_reg[13] ;
  assign \new_[3184]_  = \\u1_slt4_reg[13] ;
  assign \new_[3185]_  = \\u1_slt6_reg[13] ;
  assign \new_[3186]_  = \\u1_slt3_reg[13] ;
  assign \new_[3187]_  = ~\\u10_mem_reg[2][18] ;
  assign \new_[3188]_  = ~\\u10_mem_reg[2][19] ;
  assign \new_[3189]_  = ~\\u10_mem_reg[2][20] ;
  assign \new_[3190]_  = ~\\u10_mem_reg[2][21] ;
  assign \new_[3191]_  = ~\\u10_mem_reg[2][22] ;
  assign \new_[3192]_  = ~\\u9_mem_reg[0][18] ;
  assign \new_[3193]_  = ~\\u9_mem_reg[0][19] ;
  assign \new_[3194]_  = ~\\u10_mem_reg[2][23] ;
  assign \new_[3195]_  = ~\\u10_mem_reg[2][25] ;
  assign \new_[3196]_  = ~\\u10_mem_reg[2][26] ;
  assign \new_[3197]_  = ~\\u10_mem_reg[2][27] ;
  assign \new_[3198]_  = ~\\u9_mem_reg[1][18] ;
  assign \new_[3199]_  = ~\\u9_mem_reg[1][19] ;
  assign \new_[3200]_  = ~\\u9_mem_reg[1][20] ;
  assign \new_[3201]_  = ~\\u9_mem_reg[1][21] ;
  assign \new_[3202]_  = ~\\u10_mem_reg[2][28] ;
  assign \new_[3203]_  = ~\\u9_mem_reg[1][23] ;
  assign \new_[3204]_  = ~\\u9_mem_reg[1][24] ;
  assign \new_[3205]_  = ~\\u9_mem_reg[1][26] ;
  assign \new_[3206]_  = ~\\u10_mem_reg[2][29] ;
  assign \new_[3207]_  = ~\\u9_mem_reg[1][27] ;
  assign \new_[3208]_  = ~\\u9_mem_reg[1][29] ;
  assign \new_[3209]_  = ~\\u9_mem_reg[1][30] ;
  assign \new_[3210]_  = ~\\u9_mem_reg[1][31] ;
  assign \new_[3211]_  = ~\\u10_mem_reg[2][30] ;
  assign \new_[3212]_  = ~\\u9_mem_reg[2][18] ;
  assign \new_[3213]_  = ~\\u9_mem_reg[2][19] ;
  assign \new_[3214]_  = ~\\u10_mem_reg[2][31] ;
  assign \new_[3215]_  = ~\\u9_mem_reg[2][21] ;
  assign \new_[3216]_  = ~\\u9_mem_reg[2][22] ;
  assign \new_[3217]_  = ~\\u9_mem_reg[2][23] ;
  assign \new_[3218]_  = ~\\u9_mem_reg[2][25] ;
  assign \new_[3219]_  = ~\\u9_mem_reg[2][26] ;
  assign \new_[3220]_  = ~\\u9_mem_reg[2][27] ;
  assign \new_[3221]_  = ~\\u9_mem_reg[2][29] ;
  assign \new_[3222]_  = ~\\u9_mem_reg[2][30] ;
  assign \new_[3223]_  = ~\\u9_mem_reg[2][31] ;
  assign \new_[3224]_  = ~\\u9_mem_reg[3][18] ;
  assign \new_[3225]_  = ~\\u9_mem_reg[3][19] ;
  assign \new_[3226]_  = ~\\u9_mem_reg[3][20] ;
  assign \new_[3227]_  = ~\\u9_mem_reg[3][21] ;
  assign \new_[3228]_  = ~\\u9_mem_reg[3][23] ;
  assign \new_[3229]_  = ~\\u9_mem_reg[3][24] ;
  assign \new_[3230]_  = ~\\u9_mem_reg[3][25] ;
  assign \new_[3231]_  = ~\\u9_mem_reg[3][27] ;
  assign \new_[3232]_  = ~\\u9_mem_reg[3][28] ;
  assign \new_[3233]_  = ~\\u9_mem_reg[3][29] ;
  assign \new_[3234]_  = ~\\u9_mem_reg[3][31] ;
  assign \new_[3235]_  = ~\\u10_mem_reg[3][18] ;
  assign \new_[3236]_  = ~\\u10_mem_reg[3][19] ;
  assign \new_[3237]_  = ~\\u10_mem_reg[3][20] ;
  assign \new_[3238]_  = ~\\u10_mem_reg[3][21] ;
  assign \new_[3239]_  = ~\\u10_mem_reg[3][22] ;
  assign \new_[3240]_  = ~\\u10_mem_reg[3][23] ;
  assign \new_[3241]_  = ~\\u10_mem_reg[3][25] ;
  assign \new_[3242]_  = ~\\u10_mem_reg[3][26] ;
  assign \new_[3243]_  = ~\\u10_mem_reg[3][27] ;
  assign \new_[3244]_  = ~\\u10_mem_reg[3][29] ;
  assign \new_[3245]_  = ~\\u10_mem_reg[3][30] ;
  assign \new_[3246]_  = ~\\u10_mem_reg[3][31] ;
  assign \new_[3247]_  = ~\\u10_mem_reg[0][19] ;
  assign \new_[3248]_  = ~\\u10_mem_reg[1][18] ;
  assign \new_[3249]_  = ~\\u10_mem_reg[1][19] ;
  assign \new_[3250]_  = ~\\u10_mem_reg[1][21] ;
  assign \new_[3251]_  = ~\\u10_mem_reg[1][22] ;
  assign \new_[3252]_  = ~\\u10_mem_reg[1][23] ;
  assign \new_[3253]_  = ~\\u10_mem_reg[1][24] ;
  assign \new_[3254]_  = ~\\u10_mem_reg[1][25] ;
  assign \new_[3255]_  = ~\\u10_mem_reg[1][26] ;
  assign \new_[3256]_  = ~\\u10_mem_reg[1][27] ;
  assign \new_[3257]_  = ~\\u10_mem_reg[1][28] ;
  assign \new_[3258]_  = ~\\u10_mem_reg[1][29] ;
  assign \new_[3259]_  = ~\\u10_mem_reg[1][20] ;
  assign \new_[3260]_  = ~\\u10_mem_reg[1][30] ;
  assign \new_[3261]_  = ~\\u10_mem_reg[1][31] ;
  assign \new_[3262]_  = ~\\u11_mem_reg[3][8] ;
  assign \new_[3263]_  = ~\\u11_mem_reg[3][9] ;
  assign \new_[3264]_  = ~\\u10_mem_reg[2][1] ;
  assign \new_[3265]_  = ~\\u10_mem_reg[2][5] ;
  assign \new_[3266]_  = ~\\u10_mem_reg[2][6] ;
  assign \new_[3267]_  = ~\\u10_mem_reg[3][3] ;
  assign \new_[3268]_  = ~\\u10_mem_reg[2][9] ;
  assign \new_[3269]_  = ~\\u11_mem_reg[1][0] ;
  assign \new_[3270]_  = ~\\u11_mem_reg[1][10] ;
  assign \new_[3271]_  = ~\\u11_mem_reg[1][11] ;
  assign \new_[3272]_  = ~\\u10_mem_reg[3][2] ;
  assign \new_[3273]_  = ~\\u10_mem_reg[3][9] ;
  assign \new_[3274]_  = ~\\u11_mem_reg[1][14] ;
  assign \new_[3275]_  = ~\\u11_mem_reg[1][1] ;
  assign \new_[3276]_  = ~\\u11_mem_reg[1][2] ;
  assign \new_[3277]_  = ~\\u11_mem_reg[1][3] ;
  assign \new_[3278]_  = ~\\u11_mem_reg[1][4] ;
  assign \new_[3279]_  = ~\\u11_mem_reg[1][5] ;
  assign \new_[3280]_  = ~\\u11_mem_reg[1][7] ;
  assign \new_[3281]_  = ~\\u11_mem_reg[1][8] ;
  assign \new_[3282]_  = ~\\u11_mem_reg[1][9] ;
  assign \new_[3283]_  = ~\\u11_mem_reg[2][0] ;
  assign \new_[3284]_  = ~\\u11_mem_reg[2][10] ;
  assign \new_[3285]_  = ~\\u11_mem_reg[2][11] ;
  assign \new_[3286]_  = ~\\u11_mem_reg[2][13] ;
  assign \new_[3287]_  = ~\\u11_mem_reg[2][14] ;
  assign \new_[3288]_  = ~\\u11_mem_reg[2][15] ;
  assign \new_[3289]_  = ~\\u11_mem_reg[2][16] ;
  assign \new_[3290]_  = ~\\u11_mem_reg[1][17] ;
  assign \new_[3291]_  = ~\\u11_mem_reg[2][12] ;
  assign \new_[3292]_  = ~\\u11_mem_reg[2][2] ;
  assign \new_[3293]_  = ~\\u11_mem_reg[2][3] ;
  assign \new_[3294]_  = ~\\u11_mem_reg[2][6] ;
  assign \new_[3295]_  = ~\\u11_mem_reg[2][4] ;
  assign \new_[3296]_  = ~\\u11_mem_reg[2][5] ;
  assign \new_[3297]_  = ~\\u11_mem_reg[2][9] ;
  assign \new_[3298]_  = ~\\u11_mem_reg[3][11] ;
  assign \new_[3299]_  = ~\\u11_mem_reg[3][12] ;
  assign \new_[3300]_  = ~\\u11_mem_reg[3][15] ;
  assign \new_[3301]_  = ~\\u11_mem_reg[3][10] ;
  assign \new_[3302]_  = ~\\u11_mem_reg[3][2] ;
  assign \new_[3303]_  = ~\\u11_mem_reg[3][3] ;
  assign \new_[3304]_  = ~\\u11_mem_reg[3][4] ;
  assign \new_[3305]_  = ~\\u11_mem_reg[3][1] ;
  assign \new_[3306]_  = \\u10_wp_reg[1] ;
  assign \new_[3307]_  = \\u10_wp_reg[2] ;
  assign \new_[3308]_  = ~\\u10_mem_reg[0][2] ;
  assign \new_[3309]_  = ~\\u11_mem_reg[0][5] ;
  assign \new_[3310]_  = ~\\u10_mem_reg[0][13] ;
  assign \new_[3311]_  = ~\\u10_mem_reg[0][12] ;
  assign \new_[3312]_  = ~\\u11_mem_reg[0][16] ;
  assign \new_[3313]_  = ~\\u11_mem_reg[0][20] ;
  assign \new_[3314]_  = ~\\u11_mem_reg[0][21] ;
  assign \new_[3315]_  = ~\\u11_mem_reg[0][22] ;
  assign \new_[3316]_  = ~\\u11_mem_reg[0][23] ;
  assign \new_[3317]_  = ~\\u11_mem_reg[0][24] ;
  assign \new_[3318]_  = ~\\u11_mem_reg[0][25] ;
  assign \new_[3319]_  = ~\\u10_mem_reg[0][21] ;
  assign \new_[3320]_  = ~\\u11_mem_reg[0][26] ;
  assign \new_[3321]_  = ~\\u11_mem_reg[0][27] ;
  assign \new_[3322]_  = ~\\u10_mem_reg[0][22] ;
  assign \new_[3323]_  = ~\\u11_mem_reg[0][28] ;
  assign \new_[3324]_  = ~\\u11_mem_reg[0][29] ;
  assign \new_[3325]_  = ~\\u11_mem_reg[0][2] ;
  assign \new_[3326]_  = ~\\u11_mem_reg[0][30] ;
  assign \new_[3327]_  = ~\\u11_mem_reg[0][31] ;
  assign \new_[3328]_  = ~\\u11_mem_reg[0][3] ;
  assign \new_[3329]_  = ~\\u10_mem_reg[0][25] ;
  assign \new_[3330]_  = ~\\u11_mem_reg[0][4] ;
  assign \new_[3331]_  = ~\\u10_mem_reg[0][26] ;
  assign \new_[3332]_  = ~\\u10_mem_reg[0][27] ;
  assign \new_[3333]_  = ~\\u11_mem_reg[0][6] ;
  assign \new_[3334]_  = ~\\u10_mem_reg[0][28] ;
  assign \new_[3335]_  = ~\\u11_mem_reg[0][7] ;
  assign \new_[3336]_  = ~\\u11_mem_reg[0][8] ;
  assign \new_[3337]_  = ~\\u10_mem_reg[0][29] ;
  assign \new_[3338]_  = ~\\u11_mem_reg[0][9] ;
  assign \new_[3339]_  = ~\\u10_mem_reg[0][5] ;
  assign \new_[3340]_  = \\u11_wp_reg[0] ;
  assign \new_[3341]_  = ~\\u25_int_set_reg[2] ;
  assign \new_[3342]_  = \new_[2783]_  | \new_[3961]_ ;
  assign \new_[3343]_  = \new_[2784]_  | \new_[3962]_ ;
  assign \new_[3344]_  = ~\\u10_mem_reg[0][1] ;
  assign n1971 = ~\new_[3995]_  & ~\dma_ack_i[0] ;
  assign n1976 = ~\new_[3996]_  & ~\dma_ack_i[2] ;
  assign n1981 = ~\new_[3997]_  & ~\dma_ack_i[4] ;
  assign n1986 = ~\new_[3998]_  & ~\dma_ack_i[5] ;
  assign \new_[3349]_  = ~\\u11_mem_reg[0][17] ;
  assign n1946 = n3466 ? \new_[8996]_  : \new_[2925]_ ;
  assign \new_[3351]_  = ~\new_[3676]_  & ~\new_[14097]_ ;
  assign n1931 = n3466 ? \new_[9002]_  : \new_[2922]_ ;
  assign \new_[3353]_  = ~\new_[3677]_  & ~\new_[4515]_ ;
  assign \new_[3354]_  = ~\new_[3791]_  & ~\new_[4515]_ ;
  assign n1936 = n3466 ? \new_[9000]_  : \new_[2923]_ ;
  assign n1941 = n3466 ? \new_[9001]_  : \new_[2924]_ ;
  assign \new_[3357]_  = ~\\u10_mem_reg[3][17] ;
  assign n2546 = \\u1_sr_reg[15] ;
  assign n2026 = (~\new_[4384]_  & ~\new_[8462]_ ) | (~\new_[3022]_  & ~\new_[4514]_ );
  assign n2021 = (~\new_[4384]_  & ~\new_[8459]_ ) | (~\new_[4514]_  & ~\new_[3021]_ );
  assign n2011 = (~\new_[4385]_  & ~\new_[8859]_ ) | (~\new_[3019]_  & ~\new_[4513]_ );
  assign n2016 = (~\new_[4385]_  & ~\new_[8872]_ ) | (~\new_[4513]_  & ~\new_[3020]_ );
  assign \new_[3363]_  = ~\\u10_mem_reg[0][11] ;
  assign \new_[3364]_  = ~\\u9_mem_reg[0][4] ;
  assign n2326 = \new_[4059]_  & \new_[13876]_ ;
  assign n2331 = ~\new_[11721]_  & (~\new_[4465]_  | ~\new_[4413]_ );
  assign n2356 = ~\new_[11721]_  & (~\new_[4470]_  | ~\new_[4414]_ );
  assign n2366 = ~\new_[12040]_  & (~\new_[4469]_  | ~\new_[4446]_ );
  assign n2336 = ~\new_[12517]_  & (~\new_[4464]_  | ~\new_[4415]_ );
  assign n2341 = ~\new_[12517]_  & (~\new_[4457]_  | ~\new_[4448]_ );
  assign n2346 = ~\new_[12040]_  & (~\new_[4468]_  | ~\new_[4447]_ );
  assign n2351 = ~\new_[12517]_  & (~\new_[4471]_  | ~\new_[4416]_ );
  assign n2376 = ~\new_[12517]_  & (~\new_[4458]_  | ~\new_[4417]_ );
  assign \new_[3374]_  = \\u9_wp_reg[3] ;
  assign n2361 = ~\new_[11721]_  & (~\new_[4459]_  | ~\new_[4418]_ );
  assign n2371 = ~\new_[12517]_  & (~\new_[4460]_  | ~\new_[4419]_ );
  assign \new_[3377]_  = ~\\u9_mem_reg[0][8] ;
  assign n1991 = ~\new_[12517]_  & (~\new_[13943]_  | ~\new_[4422]_ );
  assign n2381 = ~\new_[12040]_  & (~\new_[13948]_  | ~\new_[4423]_ );
  assign n2386 = ~\new_[12040]_  & (~\new_[4461]_  | ~\new_[4424]_ );
  assign n2391 = ~\new_[11721]_  & (~\new_[4462]_  | ~\new_[4425]_ );
  assign n2396 = ~\new_[12517]_  & (~\new_[4463]_  | ~\new_[4426]_ );
  assign n2401 = ~\new_[12517]_  & (~\new_[13920]_  | ~\new_[4427]_ );
  assign n2406 = ~\new_[12710]_  & (~\new_[4428]_  | ~\new_[4529]_ );
  assign n2411 = ~\new_[12710]_  & (~\new_[4429]_  | ~\new_[4530]_ );
  assign n2416 = ~\new_[11422]_  & (~\new_[4430]_  | ~\new_[4531]_ );
  assign n2551 = ~\new_[11116]_  & (~\new_[4431]_  | ~\new_[4532]_ );
  assign n2421 = ~\new_[11422]_  & (~\new_[4432]_  | ~\new_[4533]_ );
  assign n2426 = ~\new_[12710]_  & (~\new_[4433]_  | ~\new_[4534]_ );
  assign n2431 = ~\new_[12710]_  & (~\new_[4434]_  | ~\new_[4535]_ );
  assign n2541 = ~\new_[11116]_  & (~\new_[4435]_  | ~\new_[4536]_ );
  assign n2436 = ~\new_[12710]_  & (~\new_[4537]_  | ~\new_[4436]_ );
  assign n2441 = ~\new_[11422]_  & (~\new_[4437]_  | ~\new_[4538]_ );
  assign n2446 = ~\new_[11422]_  & (~\new_[14099]_  | ~\new_[4440]_ );
  assign n2451 = ~\new_[12710]_  & (~\new_[4540]_  | ~\new_[4441]_ );
  assign n2456 = ~\new_[12710]_  & (~\new_[14070]_  | ~\new_[4442]_ );
  assign n2536 = ~\new_[11116]_  & (~\new_[4541]_  | ~\new_[4443]_ );
  assign n2461 = ~\new_[11116]_  & (~\new_[4444]_  | ~\new_[4542]_ );
  assign n2466 = ~\new_[12710]_  & (~\new_[4445]_  | ~\new_[4543]_ );
  assign n2516 = ~\new_[3659]_ ;
  assign n2521 = ~\new_[3660]_ ;
  assign n2526 = ~\new_[3661]_ ;
  assign n2531 = ~\new_[3663]_ ;
  assign \new_[3404]_  = ~\\u10_mem_reg[1][8] ;
  assign \new_[3405]_  = ~\\u9_mem_reg[0][2] ;
  assign \new_[3406]_  = ~\\u9_mem_reg[0][26] ;
  assign \new_[3407]_  = ~\\u10_mem_reg[1][6] ;
  assign \new_[3408]_  = ~\\u9_mem_reg[0][17] ;
  assign \new_[3409]_  = ~\\u9_mem_reg[0][13] ;
  assign n2511 = ~\new_[3671]_ ;
  assign \new_[3411]_  = ~\\u10_mem_reg[1][1] ;
  assign \new_[3412]_  = ~\\u10_mem_reg[1][15] ;
  assign \new_[3413]_  = ~\\u10_mem_reg[1][13] ;
  assign \new_[3414]_  = ~\\u10_mem_reg[1][10] ;
  assign \new_[3415]_  = ~\\u10_mem_reg[3][8] ;
  assign n2321 = \new_[4062]_  & \new_[13876]_ ;
  assign n1996 = \new_[4063]_  & \new_[13876]_ ;
  assign n2041 = ~\new_[4011]_  | (~\new_[9086]_  & ~\new_[4454]_ );
  assign n2046 = ~\new_[4012]_  | (~\new_[9092]_  & ~\new_[4453]_ );
  assign n2051 = ~\new_[4013]_  | (~\new_[9094]_  & ~\new_[4453]_ );
  assign n2056 = ~\new_[4014]_  | (~\new_[9098]_  & ~\new_[4453]_ );
  assign n2061 = ~\new_[4015]_  | (~\new_[9217]_  & ~\new_[4454]_ );
  assign n2066 = ~\new_[4016]_  | (~\new_[9225]_  & ~\new_[4454]_ );
  assign n2071 = ~\new_[4017]_  | (~\new_[9219]_  & ~\new_[4454]_ );
  assign n2076 = ~\new_[4018]_  | (~\new_[9221]_  & ~\new_[4453]_ );
  assign n2081 = ~\new_[4019]_  | (~\new_[9222]_  & ~\new_[4453]_ );
  assign n2086 = ~\new_[4020]_  | (~\new_[9247]_  & ~\new_[4454]_ );
  assign n2091 = ~\new_[4021]_  | (~\new_[9223]_  & ~\new_[4453]_ );
  assign n2096 = ~\new_[4022]_  | (~\new_[9228]_  & ~\new_[4454]_ );
  assign n2101 = ~\new_[4023]_  | (~\new_[9227]_  & ~\new_[4454]_ );
  assign n2106 = ~\new_[4024]_  | (~\new_[9224]_  & ~\new_[4454]_ );
  assign n2111 = ~\new_[4025]_  | (~\new_[9215]_  & ~\new_[4453]_ );
  assign n2116 = ~\new_[4026]_  | (~\new_[9191]_  & ~\new_[4453]_ );
  assign n2121 = ~\new_[4027]_  | (~\new_[9095]_  & ~\new_[4454]_ );
  assign n2126 = ~\new_[4028]_  | (~\new_[9096]_  & ~\new_[4453]_ );
  assign n2131 = ~\new_[4029]_  | (~\new_[9216]_  & ~\new_[4454]_ );
  assign n2136 = ~\new_[4030]_  | (~\new_[9229]_  & ~\new_[4454]_ );
  assign n2141 = ~\new_[4031]_  | (~\new_[9230]_  & ~\new_[4454]_ );
  assign n2146 = ~\new_[4032]_  | (~\new_[9231]_  & ~\new_[4454]_ );
  assign n2151 = ~\new_[4033]_  | (~\new_[9226]_  & ~\new_[4454]_ );
  assign n2156 = ~\new_[4034]_  | (~\new_[9232]_  & ~\new_[4454]_ );
  assign n2161 = ~\new_[4035]_  | (~\new_[9233]_  & ~\new_[4454]_ );
  assign n2166 = ~\new_[4036]_  | (~\new_[9234]_  & ~\new_[4454]_ );
  assign n2171 = ~\new_[4037]_  | (~\new_[9235]_  & ~\new_[4453]_ );
  assign n2176 = ~\new_[4038]_  | (~\new_[9238]_  & ~\new_[4454]_ );
  assign n2181 = ~\new_[4039]_  | (~\new_[9239]_  & ~\new_[4454]_ );
  assign n2186 = ~\new_[4040]_  | (~\new_[9237]_  & ~\new_[4454]_ );
  assign \new_[3448]_  = ~\\u10_mem_reg[0][23] ;
  assign \new_[3449]_  = \\u11_din_tmp1_reg[8] ;
  assign \new_[3450]_  = ~\\u9_mem_reg[2][12] ;
  assign \new_[3451]_  = ~\\u10_mem_reg[3][13] ;
  assign \new_[3452]_  = ~\\u10_mem_reg[3][0] ;
  assign \new_[3453]_  = ~\\u9_mem_reg[3][4] ;
  assign \new_[3454]_  = ~\\u9_mem_reg[3][1] ;
  assign \new_[3455]_  = ~\\u9_mem_reg[3][15] ;
  assign \new_[3456]_  = ~\\u9_mem_reg[2][5] ;
  assign \new_[3457]_  = ~\\u9_mem_reg[2][2] ;
  assign \new_[3458]_  = ~\\u10_mem_reg[1][9] ;
  assign \new_[3459]_  = ~\\u10_mem_reg[2][0] ;
  assign \new_[3460]_  = ~\\u10_mem_reg[2][11] ;
  assign \new_[3461]_  = ~\\u10_mem_reg[2][12] ;
  assign \new_[3462]_  = ~\\u10_mem_reg[2][13] ;
  assign \new_[3463]_  = ~\\u10_mem_reg[2][14] ;
  assign \new_[3464]_  = ~\\u10_mem_reg[2][15] ;
  assign \new_[3465]_  = ~\\u10_mem_reg[2][16] ;
  assign \new_[3466]_  = ~\\u10_mem_reg[2][10] ;
  assign \new_[3467]_  = ~\\u9_mem_reg[1][0] ;
  assign \new_[3468]_  = ~\\u9_mem_reg[1][10] ;
  assign \new_[3469]_  = ~\\u9_mem_reg[1][12] ;
  assign \new_[3470]_  = ~\\u9_mem_reg[1][13] ;
  assign \new_[3471]_  = ~\\u9_mem_reg[1][14] ;
  assign \new_[3472]_  = ~\\u9_mem_reg[1][16] ;
  assign \new_[3473]_  = ~\\u9_mem_reg[1][17] ;
  assign \new_[3474]_  = ~\\u9_mem_reg[1][1] ;
  assign \new_[3475]_  = ~\\u9_mem_reg[1][2] ;
  assign \new_[3476]_  = ~\\u9_mem_reg[1][3] ;
  assign \new_[3477]_  = ~\\u9_mem_reg[1][4] ;
  assign \new_[3478]_  = ~\\u9_mem_reg[1][5] ;
  assign \new_[3479]_  = ~\\u9_mem_reg[1][6] ;
  assign \new_[3480]_  = ~\\u9_mem_reg[1][7] ;
  assign \new_[3481]_  = ~\\u9_mem_reg[1][8] ;
  assign \new_[3482]_  = ~\\u9_mem_reg[2][0] ;
  assign \new_[3483]_  = ~\\u9_mem_reg[2][10] ;
  assign \new_[3484]_  = ~\\u9_mem_reg[2][11] ;
  assign \new_[3485]_  = ~\\u9_mem_reg[2][14] ;
  assign \new_[3486]_  = ~\\u9_mem_reg[2][15] ;
  assign \new_[3487]_  = ~\\u9_mem_reg[2][16] ;
  assign \new_[3488]_  = ~\\u9_mem_reg[2][17] ;
  assign \new_[3489]_  = ~\\u9_mem_reg[2][1] ;
  assign \new_[3490]_  = ~\\u10_mem_reg[2][3] ;
  assign \new_[3491]_  = ~\\u9_mem_reg[2][3] ;
  assign \new_[3492]_  = ~\\u10_mem_reg[2][4] ;
  assign \new_[3493]_  = ~\\u9_mem_reg[2][4] ;
  assign \new_[3494]_  = ~\\u9_mem_reg[2][6] ;
  assign \new_[3495]_  = ~\\u9_mem_reg[2][7] ;
  assign \new_[3496]_  = ~\\u9_mem_reg[2][8] ;
  assign \new_[3497]_  = ~\\u9_mem_reg[3][0] ;
  assign \new_[3498]_  = ~\\u9_mem_reg[3][10] ;
  assign \new_[3499]_  = ~\\u9_mem_reg[3][11] ;
  assign \new_[3500]_  = ~\\u9_mem_reg[3][12] ;
  assign \new_[3501]_  = ~\\u9_mem_reg[3][13] ;
  assign \new_[3502]_  = ~\\u9_mem_reg[3][14] ;
  assign \new_[3503]_  = ~\\u9_mem_reg[2][13] ;
  assign \new_[3504]_  = ~\\u9_mem_reg[3][16] ;
  assign \new_[3505]_  = ~\\u9_mem_reg[3][17] ;
  assign \new_[3506]_  = ~\\u10_mem_reg[2][7] ;
  assign \new_[3507]_  = ~\\u9_mem_reg[3][2] ;
  assign \new_[3508]_  = ~\\u9_mem_reg[3][3] ;
  assign \new_[3509]_  = ~\\u9_mem_reg[3][5] ;
  assign \new_[3510]_  = ~\\u9_mem_reg[3][6] ;
  assign \new_[3511]_  = ~\\u9_mem_reg[3][7] ;
  assign \new_[3512]_  = ~\\u10_mem_reg[2][8] ;
  assign \new_[3513]_  = ~\\u9_mem_reg[3][9] ;
  assign \new_[3514]_  = ~\\u9_mem_reg[3][8] ;
  assign \new_[3515]_  = ~\\u10_mem_reg[3][10] ;
  assign \new_[3516]_  = ~\\u10_mem_reg[3][11] ;
  assign \new_[3517]_  = ~\\u10_mem_reg[3][12] ;
  assign \new_[3518]_  = ~\\u10_mem_reg[3][14] ;
  assign \new_[3519]_  = ~\\u10_mem_reg[3][15] ;
  assign \new_[3520]_  = ~\\u10_mem_reg[3][16] ;
  assign \new_[3521]_  = ~\\u10_mem_reg[3][1] ;
  assign \new_[3522]_  = ~\\u10_mem_reg[3][4] ;
  assign \new_[3523]_  = ~\\u10_mem_reg[3][5] ;
  assign \new_[3524]_  = ~\\u10_mem_reg[3][6] ;
  assign \new_[3525]_  = ~\\u10_mem_reg[3][7] ;
  assign n2191 = ~\new_[4041]_  | (~\new_[8843]_  & ~\new_[4453]_ );
  assign \new_[3527]_  = ~\\u10_mem_reg[1][11] ;
  assign \new_[3528]_  = ~\\u10_mem_reg[1][12] ;
  assign \new_[3529]_  = ~\\u10_mem_reg[1][14] ;
  assign \new_[3530]_  = ~\\u10_mem_reg[1][17] ;
  assign \new_[3531]_  = ~\\u10_mem_reg[1][16] ;
  assign \new_[3532]_  = ~\\u9_mem_reg[1][9] ;
  assign \new_[3533]_  = ~\\u10_mem_reg[1][3] ;
  assign \new_[3534]_  = ~\\u10_mem_reg[1][4] ;
  assign \new_[3535]_  = ~\\u10_mem_reg[1][5] ;
  assign \new_[3536]_  = ~\\u10_mem_reg[1][2] ;
  assign \new_[3537]_  = ~\\u10_mem_reg[2][2] ;
  assign \new_[3538]_  = ~\\u10_mem_reg[1][7] ;
  assign n2196 = ~\new_[4042]_  | (~\new_[8842]_  & ~\new_[4453]_ );
  assign \new_[3540]_  = \\u9_wp_reg[2] ;
  assign \new_[3541]_  = ~\\u9_mem_reg[1][15] ;
  assign \new_[3542]_  = ~\\u9_mem_reg[1][11] ;
  assign \new_[3543]_  = ~\\u10_mem_reg[2][17] ;
  assign \new_[3544]_  = ~\\u10_mem_reg[0][24] ;
  assign n2201 = ~\new_[4043]_  | (~\new_[8960]_  & ~\new_[4453]_ );
  assign \new_[3546]_  = \\u11_din_tmp1_reg[4] ;
  assign \new_[3547]_  = ~\\u10_mem_reg[0][8] ;
  assign \new_[3548]_  = ~\\u10_mem_reg[0][4] ;
  assign \new_[3549]_  = ~\\u9_mem_reg[0][0] ;
  assign \new_[3550]_  = ~\\u9_mem_reg[0][10] ;
  assign \new_[3551]_  = ~\\u9_mem_reg[0][11] ;
  assign \new_[3552]_  = ~\\u9_mem_reg[0][12] ;
  assign \new_[3553]_  = ~\\u9_mem_reg[0][14] ;
  assign \new_[3554]_  = ~\\u9_mem_reg[0][15] ;
  assign \new_[3555]_  = ~\\u9_mem_reg[0][16] ;
  assign \new_[3556]_  = ~\\u9_mem_reg[0][1] ;
  assign \new_[3557]_  = ~\\u9_mem_reg[0][20] ;
  assign \new_[3558]_  = ~\\u9_mem_reg[0][21] ;
  assign \new_[3559]_  = ~\\u9_mem_reg[0][22] ;
  assign \new_[3560]_  = ~\\u9_mem_reg[0][23] ;
  assign \new_[3561]_  = ~\\u9_mem_reg[0][24] ;
  assign \new_[3562]_  = ~\\u9_mem_reg[0][25] ;
  assign \new_[3563]_  = ~\\u9_mem_reg[0][27] ;
  assign \new_[3564]_  = ~\\u9_mem_reg[0][28] ;
  assign \new_[3565]_  = ~\\u9_mem_reg[0][29] ;
  assign \new_[3566]_  = ~\\u9_mem_reg[0][30] ;
  assign \new_[3567]_  = ~\\u9_mem_reg[0][31] ;
  assign \new_[3568]_  = ~\\u9_mem_reg[0][3] ;
  assign \new_[3569]_  = ~\\u9_mem_reg[0][5] ;
  assign \new_[3570]_  = ~\\u9_mem_reg[0][6] ;
  assign \new_[3571]_  = ~\\u9_mem_reg[0][7] ;
  assign \new_[3572]_  = ~\\u9_mem_reg[0][9] ;
  assign \new_[3573]_  = ~\\u10_mem_reg[0][0] ;
  assign \new_[3574]_  = ~\\u10_mem_reg[0][10] ;
  assign n2206 = ~\new_[4044]_  | (~\new_[8944]_  & ~\new_[4454]_ );
  assign \new_[3576]_  = ~\\u10_mem_reg[0][14] ;
  assign \new_[3577]_  = ~\\u10_mem_reg[0][15] ;
  assign \new_[3578]_  = ~\\u10_mem_reg[0][16] ;
  assign \new_[3579]_  = ~\\u10_mem_reg[0][17] ;
  assign n2211 = ~\new_[4045]_  | (~\new_[8963]_  & ~\new_[4454]_ );
  assign \new_[3581]_  = ~\\u10_mem_reg[0][31] ;
  assign \new_[3582]_  = ~\\u10_mem_reg[0][3] ;
  assign \new_[3583]_  = ~\\u10_mem_reg[0][30] ;
  assign \new_[3584]_  = ~\\u10_mem_reg[0][6] ;
  assign \new_[3585]_  = ~\\u10_mem_reg[0][7] ;
  assign \new_[3586]_  = ~\\u10_mem_reg[0][9] ;
  assign \new_[3587]_  = \\u10_wp_reg[0] ;
  assign \new_[3588]_  = \\u11_din_tmp1_reg[0] ;
  assign \new_[3589]_  = \\u11_din_tmp1_reg[10] ;
  assign \new_[3590]_  = \\u11_din_tmp1_reg[11] ;
  assign \new_[3591]_  = \\u11_din_tmp1_reg[12] ;
  assign \new_[3592]_  = \\u11_din_tmp1_reg[13] ;
  assign \new_[3593]_  = \\u11_din_tmp1_reg[14] ;
  assign \new_[3594]_  = \\u11_din_tmp1_reg[15] ;
  assign \new_[3595]_  = \\u11_din_tmp1_reg[1] ;
  assign \new_[3596]_  = \\u11_din_tmp1_reg[2] ;
  assign \new_[3597]_  = \\u11_din_tmp1_reg[3] ;
  assign \new_[3598]_  = \\u11_din_tmp1_reg[5] ;
  assign \new_[3599]_  = \\u11_din_tmp1_reg[6] ;
  assign \new_[3600]_  = \\u11_din_tmp1_reg[7] ;
  assign \new_[3601]_  = \\u11_din_tmp1_reg[9] ;
  assign \new_[3602]_  = ~\\u9_mem_reg[2][9] ;
  assign \new_[3603]_  = ~\\u18_int_set_reg[1] ;
  assign \new_[3604]_  = ~\\u19_int_set_reg[1] ;
  assign \new_[3605]_  = ~\\u24_int_set_reg[2] ;
  assign \new_[3606]_  = u15_crac_wr_reg;
  assign \new_[3607]_  = \\u13_ints_r_reg[1] ;
  assign n2216 = ~\new_[4046]_  | (~\new_[8962]_  & ~\new_[4453]_ );
  assign n2221 = ~\new_[4047]_  | (~\new_[8959]_  & ~\new_[4454]_ );
  assign n2226 = ~\new_[4048]_  | (~\new_[8961]_  & ~\new_[4454]_ );
  assign n2231 = ~\new_[4049]_  | (~\new_[8957]_  & ~\new_[4454]_ );
  assign n2236 = ~\new_[4050]_  | (~\new_[8956]_  & ~\new_[4454]_ );
  assign n2241 = ~\new_[4051]_  | (~\new_[8958]_  & ~\new_[4454]_ );
  assign n2246 = ~\new_[4052]_  | (~\new_[8945]_  & ~\new_[4454]_ );
  assign n2251 = ~\new_[4053]_  | (~\new_[8953]_  & ~\new_[4453]_ );
  assign n2256 = ~\new_[4054]_  | (~\new_[8946]_  & ~\new_[4453]_ );
  assign n2266 = \new_[8237]_  ? \new_[4452]_  : \new_[13736]_ ;
  assign n2271 = \new_[8238]_  ? \new_[4454]_  : \new_[13737]_ ;
  assign n2276 = \new_[8522]_  ? \new_[4616]_  : \new_[13727]_ ;
  assign \new_[3620]_  = ~\\u10_mem_reg[0][20] ;
  assign n2281 = \new_[8526]_  ? \new_[4452]_  : \new_[13680]_ ;
  assign n2286 = \new_[8259]_  ? \new_[4452]_  : \new_[13613]_ ;
  assign n2291 = \new_[8230]_  ? \new_[4452]_  : \new_[13777]_ ;
  assign n2296 = \new_[8268]_  ? \new_[4452]_  : \new_[13192]_ ;
  assign n2301 = \new_[8511]_  ? \new_[4452]_  : \new_[13236]_ ;
  assign n2306 = \new_[8509]_  ? \new_[4452]_  : \new_[13652]_ ;
  assign \new_[3627]_  = \new_[2816]_  | \new_[4245]_ ;
  assign \new_[3628]_  = \new_[2817]_  | \new_[4246]_ ;
  assign \new_[3629]_  = \new_[2818]_  | \new_[4247]_ ;
  assign \new_[3630]_  = \new_[2819]_  | \new_[4249]_ ;
  assign n2311 = \new_[8220]_  ? \new_[4452]_  : \new_[13274]_ ;
  assign n2316 = \new_[8184]_  ? \new_[4616]_  : \new_[13304]_ ;
  assign n2261 = \new_[8197]_  ? \new_[4616]_  : \new_[13342]_ ;
  assign \new_[3634]_  = \new_[2828]_  ^ \new_[4450]_ ;
  assign \new_[3635]_  = \new_[13140]_  ^ \new_[4451]_ ;
  assign n2471 = \new_[8293]_  ? \new_[4454]_  : \new_[13658]_ ;
  assign n2476 = \new_[8295]_  ? \new_[4454]_  : \new_[13674]_ ;
  assign n2481 = \new_[8296]_  ? \new_[4454]_  : \new_[13686]_ ;
  assign n2491 = \new_[8298]_  ? \new_[4616]_  : \new_[13742]_ ;
  assign n2486 = \new_[8297]_  ? \new_[4616]_  : \new_[13212]_ ;
  assign n2496 = \new_[8299]_  ? \new_[4616]_  : \new_[13534]_ ;
  assign n2501 = \new_[8300]_  ? \new_[4616]_  : \new_[13540]_ ;
  assign n2506 = \new_[8288]_  ? \new_[4616]_  : \new_[13682]_ ;
  assign \new_[3644]_  = \new_[13154]_  ^ \new_[4455]_ ;
  assign \new_[3645]_  = \new_[2831]_  ^ \new_[4456]_ ;
  assign \new_[3646]_  = ~\new_[4003]_  & (~\new_[4730]_  | ~\new_[12730]_ );
  assign \new_[3647]_  = ~\new_[4004]_  & (~\new_[4731]_  | ~\new_[13048]_ );
  assign n2031 = \new_[4237]_  & \new_[12325]_ ;
  assign n2036 = \new_[4238]_  & \new_[12691]_ ;
  assign \new_[3650]_  = \\u0_slt9_r_reg[3] ;
  assign n3016 = ~\new_[4376]_  | (~\new_[9734]_  & ~\new_[4518]_ );
  assign n2656 = n4466 ? \new_[8996]_  : \new_[3183]_ ;
  assign n2671 = n4466 ? \new_[9002]_  : \new_[3186]_ ;
  assign n2661 = n4466 ? \new_[9000]_  : \new_[3184]_ ;
  assign n3276 = \new_[4394]_  & \new_[13873]_ ;
  assign n2666 = n4466 ? \new_[9001]_  : \new_[3185]_ ;
  assign \new_[3657]_  = \\u10_din_tmp1_reg[13] ;
  assign \new_[3658]_  = ~\new_[12993]_  | ~\new_[12591]_  | ~\new_[4475]_ ;
  assign \new_[3659]_  = ~\new_[13629]_  & (~\new_[6829]_  | ~\new_[14161]_ );
  assign \new_[3660]_  = ~\new_[13789]_  & (~\new_[6561]_  | ~\new_[4475]_ );
  assign \new_[3661]_  = ~\new_[13597]_  & (~\new_[6833]_  | ~\new_[13962]_ );
  assign \new_[3662]_  = ~\new_[12686]_  | ~\new_[12544]_  | ~\new_[14061]_ ;
  assign \new_[3663]_  = ~\new_[13822]_  & (~\new_[6834]_  | ~\new_[4478]_ );
  assign n3446 = ~\new_[4058]_ ;
  assign \new_[3665]_  = ~\new_[13012]_  | ~\new_[13935]_  | ~\new_[14161]_ ;
  assign \new_[3666]_  = ~\new_[12519]_  | ~\new_[12583]_  | ~\new_[4478]_ ;
  assign \new_[3667]_  = ~\new_[4420]_  & (~\new_[13201]_  | ~\new_[13927]_ );
  assign \new_[3668]_  = ~\new_[4421]_  & (~\new_[13661]_  | ~\new_[13927]_ );
  assign \new_[3669]_  = ~\new_[4438]_  & (~\new_[13433]_  | ~\new_[4622]_ );
  assign \new_[3670]_  = ~\new_[4439]_  & (~\new_[13405]_  | ~\new_[4622]_ );
  assign \new_[3671]_  = (~\new_[4545]_  | ~\new_[3119]_ ) & (~\new_[5055]_  | ~\new_[6835]_ );
  assign \new_[3672]_  = \\u1_slt6_reg[12] ;
  assign n3271 = \new_[4397]_  & \new_[13873]_ ;
  assign n2581 = \new_[4398]_  & \new_[13873]_ ;
  assign n3441 = ~\new_[4286]_  | ~\new_[4449]_ ;
  assign \new_[3676]_  = ~\new_[4392]_  & (~\new_[13902]_  | ~\new_[13989]_ );
  assign \new_[3677]_  = ~\new_[4393]_  & (~\new_[14001]_  | ~\new_[13091]_ );
  assign \new_[3678]_  = ~\new_[4395]_  & (~\new_[13900]_  | ~\new_[13104]_ );
  assign \new_[3679]_  = ~\new_[4396]_  & (~\new_[13898]_  | ~\new_[13151]_ );
  assign n2676 = ~\new_[4288]_  | (~\new_[9087]_  & ~\new_[4518]_ );
  assign n2681 = ~\new_[4290]_  | (~\new_[9088]_  & ~\new_[4519]_ );
  assign n2686 = ~\new_[4291]_  | (~\new_[9192]_  & ~\new_[4519]_ );
  assign n2691 = ~\new_[4292]_  | (~\new_[9715]_  & ~\new_[4519]_ );
  assign n2696 = ~\new_[4293]_  | (~\new_[9193]_  & ~\new_[4518]_ );
  assign n2711 = ~\new_[4294]_  | (~\new_[9246]_  & ~\new_[4519]_ );
  assign n2701 = ~\new_[4295]_  | (~\new_[8692]_  & ~\new_[4595]_ );
  assign n2706 = ~\new_[4296]_  | (~\new_[8693]_  & ~\new_[4595]_ );
  assign n2621 = ~\new_[4297]_  | (~\new_[9194]_  & ~\new_[4519]_ );
  assign n2716 = ~\new_[4298]_  | (~\new_[9195]_  & ~\new_[4519]_ );
  assign n2721 = ~\new_[4299]_  | (~\new_[9736]_  & ~\new_[4519]_ );
  assign n2726 = ~\new_[4301]_  | (~\new_[9737]_  & ~\new_[4518]_ );
  assign n2751 = ~\new_[4302]_  | (~\new_[9741]_  & ~\new_[4519]_ );
  assign n2731 = ~\new_[4303]_  | (~\new_[8694]_  & ~\new_[4595]_ );
  assign n2736 = ~\new_[4365]_  | (~\new_[8697]_  & ~\new_[4595]_ );
  assign n2741 = ~\new_[4304]_  | (~\new_[9717]_  & ~\new_[4595]_ );
  assign n2746 = ~\new_[4305]_  | (~\new_[9718]_  & ~\new_[4655]_ );
  assign n2771 = ~\new_[4308]_  | (~\new_[9213]_  & ~\new_[4519]_ );
  assign n2616 = ~\new_[4306]_  | (~\new_[9714]_  & ~\new_[4655]_ );
  assign n2756 = ~\new_[4307]_  | (~\new_[9719]_  & ~\new_[4595]_ );
  assign n2761 = ~\new_[4361]_  | (~\new_[9740]_  & ~\new_[4595]_ );
  assign n2611 = ~\new_[4309]_  | (~\new_[9720]_  & ~\new_[4595]_ );
  assign n2766 = ~\new_[4310]_  | (~\new_[9742]_  & ~\new_[4655]_ );
  assign n2776 = ~\new_[4311]_  | (~\new_[9721]_  & ~\new_[4595]_ );
  assign n2606 = ~\new_[4312]_  | (~\new_[9722]_  & ~\new_[4655]_ );
  assign n2781 = ~\new_[4313]_  | (~\new_[9723]_  & ~\new_[4595]_ );
  assign n2786 = ~\new_[4314]_  | (~\new_[9724]_  & ~\new_[4655]_ );
  assign n2791 = ~\new_[4315]_  | (~\new_[9725]_  & ~\new_[4595]_ );
  assign n2796 = ~\new_[4316]_  | (~\new_[9220]_  & ~\new_[4519]_ );
  assign n2811 = ~\new_[4317]_  | (~\new_[9214]_  & ~\new_[4518]_ );
  assign n2801 = ~\new_[4318]_  | (~\new_[8695]_  & ~\new_[4598]_ );
  assign n2806 = ~\new_[4319]_  | (~\new_[8696]_  & ~\new_[4595]_ );
  assign n2601 = ~\new_[4320]_  | (~\new_[9727]_  & ~\new_[4655]_ );
  assign n2816 = ~\new_[4321]_  | (~\new_[9743]_  & ~\new_[4655]_ );
  assign n2821 = ~\new_[4322]_  | (~\new_[9728]_  & ~\new_[4595]_ );
  assign n2826 = ~\new_[4323]_  | (~\new_[9738]_  & ~\new_[4655]_ );
  assign n2596 = ~\new_[4324]_  | (~\new_[9729]_  & ~\new_[4595]_ );
  assign n2831 = ~\new_[4362]_  | (~\new_[9739]_  & ~\new_[4655]_ );
  assign n2836 = ~\new_[4325]_  | (~\new_[9730]_  & ~\new_[4595]_ );
  assign n2841 = ~\new_[4326]_  | (~\new_[9745]_  & ~\new_[4655]_ );
  assign n2591 = ~\new_[4327]_  | (~\new_[9731]_  & ~\new_[4595]_ );
  assign n2846 = ~\new_[4328]_  | (~\new_[9732]_  & ~\new_[4598]_ );
  assign n2851 = ~\new_[4329]_  | (~\new_[9735]_  & ~\new_[4598]_ );
  assign n2856 = ~\new_[4330]_  | (~\new_[9733]_  & ~\new_[4655]_ );
  assign n2861 = ~\new_[4331]_  | (~\new_[8453]_  & ~\new_[4655]_ );
  assign n2866 = ~\new_[4332]_  | (~\new_[8454]_  & ~\new_[4595]_ );
  assign n2871 = ~\new_[4333]_  | (~\new_[9240]_  & ~\new_[4595]_ );
  assign n2876 = ~\new_[4334]_  | (~\new_[9196]_  & ~\new_[4595]_ );
  assign n2586 = ~\new_[4335]_  | (~\new_[9212]_  & ~\new_[4598]_ );
  assign n2881 = ~\new_[4336]_  | (~\new_[9197]_  & ~\new_[4595]_ );
  assign n2886 = ~\new_[4337]_  | (~\new_[9218]_  & ~\new_[4595]_ );
  assign n2891 = ~\new_[4338]_  | (~\new_[9236]_  & ~\new_[4595]_ );
  assign n2576 = ~\new_[4359]_  | (~\new_[9198]_  & ~\new_[4595]_ );
  assign n2896 = ~\new_[4339]_  | (~\new_[9199]_  & ~\new_[4655]_ );
  assign n2901 = ~\new_[4340]_  | (~\new_[9210]_  & ~\new_[4655]_ );
  assign n2906 = ~\new_[4341]_  | (~\new_[9211]_  & ~\new_[4655]_ );
  assign n2571 = ~\new_[4342]_  | (~\new_[9200]_  & ~\new_[4595]_ );
  assign n2911 = ~\new_[4343]_  | (~\new_[9208]_  & ~\new_[4655]_ );
  assign n2916 = ~\new_[4344]_  | (~\new_[8844]_  & ~\new_[4519]_ );
  assign n2921 = ~\new_[4345]_  | (~\new_[8845]_  & ~\new_[4519]_ );
  assign n2926 = ~\new_[4346]_  | (~\new_[8947]_  & ~\new_[4518]_ );
  assign n2931 = ~\new_[4347]_  | (~\new_[9201]_  & ~\new_[4519]_ );
  assign n2936 = ~\new_[4348]_  | (~\new_[8948]_  & ~\new_[4519]_ );
  assign n2941 = ~\new_[4349]_  | (~\new_[8949]_  & ~\new_[4518]_ );
  assign n2566 = ~\new_[4350]_  | (~\new_[8950]_  & ~\new_[4518]_ );
  assign n2946 = ~\new_[4351]_  | (~\new_[8951]_  & ~\new_[4518]_ );
  assign n2951 = ~\new_[4352]_  | (~\new_[9204]_  & ~\new_[4518]_ );
  assign n2956 = ~\new_[4353]_  | (~\new_[9205]_  & ~\new_[4519]_ );
  assign n2561 = ~\new_[4354]_  | (~\new_[9207]_  & ~\new_[4519]_ );
  assign n2961 = ~\new_[4355]_  | (~\new_[8952]_  & ~\new_[4519]_ );
  assign n2966 = ~\new_[4356]_  | (~\new_[8954]_  & ~\new_[4519]_ );
  assign n2971 = ~\new_[4357]_  | (~\new_[8955]_  & ~\new_[4518]_ );
  assign n2556 = ~\new_[4363]_  | (~\new_[9091]_  & ~\new_[4518]_ );
  assign n2976 = ~\new_[4364]_  | (~\new_[9093]_  & ~\new_[4519]_ );
  assign n2981 = ~\new_[4368]_  | (~\new_[9097]_  & ~\new_[4519]_ );
  assign n2986 = ~\new_[4369]_  | (~\new_[9089]_  & ~\new_[4519]_ );
  assign n3036 = ~\new_[4370]_  | (~\new_[9241]_  & ~\new_[4519]_ );
  assign n2991 = ~\new_[4371]_  | (~\new_[9744]_  & ~\new_[4518]_ );
  assign n2996 = ~\new_[4372]_  | (~\new_[9242]_  & ~\new_[4518]_ );
  assign n3001 = ~\new_[4373]_  | (~\new_[9243]_  & ~\new_[4519]_ );
  assign \new_[3760]_  = \\u13_ints_r_reg[26] ;
  assign \new_[3761]_  = \\u1_slt0_reg[12] ;
  assign \new_[3762]_  = \\u1_slt2_reg[12] ;
  assign \new_[3763]_  = \\u1_slt3_reg[12] ;
  assign \new_[3764]_  = \\u1_slt4_reg[12] ;
  assign n3006 = ~\new_[4374]_  | (~\new_[9244]_  & ~\new_[4519]_ );
  assign \new_[3766]_  = \\u10_din_tmp1_reg[11] ;
  assign n3011 = ~\new_[4375]_  | (~\new_[9206]_  & ~\new_[4519]_ );
  assign n3031 = ~\new_[4379]_  | (~\new_[9245]_  & ~\new_[4519]_ );
  assign n3021 = ~\new_[4377]_  | (~\new_[9726]_  & ~\new_[4518]_ );
  assign n3026 = ~\new_[4378]_  | (~\new_[9716]_  & ~\new_[4518]_ );
  assign \new_[3771]_  = \\u9_wp_reg[0] ;
  assign n3046 = ~\new_[4381]_  | (~\new_[9209]_  & ~\new_[4519]_ );
  assign \new_[3773]_  = \\u10_din_tmp1_reg[5] ;
  assign \new_[3774]_  = \\u10_din_tmp1_reg[3] ;
  assign n3041 = ~\new_[4380]_  | (~\new_[9202]_  & ~\new_[4519]_ );
  assign \new_[3776]_  = \\u10_din_tmp1_reg[1] ;
  assign \new_[3777]_  = \\u10_din_tmp1_reg[2] ;
  assign \new_[3778]_  = \\u10_din_tmp1_reg[4] ;
  assign \new_[3779]_  = \\u10_din_tmp1_reg[6] ;
  assign \new_[3780]_  = \\u10_din_tmp1_reg[8] ;
  assign \new_[3781]_  = \\u10_din_tmp1_reg[9] ;
  assign \new_[3782]_  = \\u10_din_tmp1_reg[7] ;
  assign \new_[3783]_  = \\u10_din_tmp1_reg[0] ;
  assign \new_[3784]_  = \\u10_din_tmp1_reg[10] ;
  assign \new_[3785]_  = \\u10_din_tmp1_reg[15] ;
  assign \new_[3786]_  = \\u10_din_tmp1_reg[14] ;
  assign \new_[3787]_  = \\u10_din_tmp1_reg[12] ;
  assign \new_[3788]_  = u15_rdd1_reg;
  assign \new_[3789]_  = ~u15_rdd2_reg;
  assign \new_[3790]_  = ~\new_[4382]_  & (~\new_[13902]_  | ~\new_[2756]_ );
  assign \new_[3791]_  = ~\new_[4383]_  & (~\new_[14001]_  | ~\new_[2757]_ );
  assign \new_[3792]_  = ~\new_[4389]_  & (~\new_[13900]_  | ~\new_[2758]_ );
  assign \new_[3793]_  = ~\new_[4391]_  & (~\new_[13898]_  | ~\new_[2759]_ );
  assign n3051 = \new_[8188]_  ? \new_[4521]_  : \new_[13348]_ ;
  assign n3056 = \new_[8505]_  ? \new_[4521]_  : \new_[13191]_ ;
  assign n3061 = \new_[8508]_  ? \new_[4519]_  : \new_[13543]_ ;
  assign n3066 = \new_[8198]_  ? \new_[4661]_  : \new_[13806]_ ;
  assign \new_[3798]_  = ~\new_[13651]_  | ~\new_[4477]_ ;
  assign n3071 = \new_[8202]_  ? \new_[4661]_  : \new_[13240]_ ;
  assign \new_[3800]_  = ~\new_[13225]_  | ~\new_[4474]_ ;
  assign \new_[3801]_  = ~\new_[13507]_  | ~\new_[4474]_ ;
  assign \new_[3802]_  = ~\new_[13198]_  | ~\new_[4474]_ ;
  assign \new_[3803]_  = ~\new_[13462]_  | ~\new_[4474]_ ;
  assign \new_[3804]_  = ~\new_[13595]_  | ~\new_[4474]_ ;
  assign \new_[3805]_  = ~\new_[13697]_  | ~\new_[4474]_ ;
  assign \new_[3806]_  = ~\new_[13469]_  | ~\new_[4474]_ ;
  assign \new_[3807]_  = ~\new_[13648]_  | ~\new_[4474]_ ;
  assign \new_[3808]_  = ~\new_[13506]_  | ~\new_[4472]_ ;
  assign \new_[3809]_  = ~\new_[13206]_  | ~\new_[4474]_ ;
  assign \new_[3810]_  = ~\new_[13388]_  | ~\new_[4474]_ ;
  assign \new_[3811]_  = ~\new_[4623]_  & (~\new_[8083]_  | ~\new_[8620]_ );
  assign \new_[3812]_  = ~\new_[4623]_  & (~\new_[8372]_  | ~\new_[8373]_ );
  assign \new_[3813]_  = ~\new_[13331]_  | ~\new_[4474]_ ;
  assign \new_[3814]_  = ~\new_[13561]_  | ~\new_[4474]_ ;
  assign \new_[3815]_  = ~\new_[13531]_  | ~\new_[4474]_ ;
  assign \new_[3816]_  = ~\new_[13255]_  | ~\new_[4474]_ ;
  assign \new_[3817]_  = ~\new_[13445]_  | ~\new_[4474]_ ;
  assign \new_[3818]_  = ~\new_[13244]_  | ~\new_[4474]_ ;
  assign \new_[3819]_  = ~\new_[13642]_  | ~\new_[4476]_ ;
  assign \new_[3820]_  = ~\new_[13608]_  | ~\new_[4476]_ ;
  assign \new_[3821]_  = ~\new_[13547]_  | ~\new_[4476]_ ;
  assign \new_[3822]_  = ~\new_[13780]_  | ~\new_[4476]_ ;
  assign \new_[3823]_  = ~\new_[13508]_  | ~\new_[4476]_ ;
  assign \new_[3824]_  = ~\new_[13493]_  | ~\new_[4476]_ ;
  assign \new_[3825]_  = ~\new_[13775]_  | ~\new_[4476]_ ;
  assign \new_[3826]_  = ~\new_[13492]_  | ~\new_[4476]_ ;
  assign \new_[3827]_  = ~\new_[13767]_  | ~\new_[4476]_ ;
  assign \new_[3828]_  = ~\new_[13343]_  | ~\new_[4476]_ ;
  assign \new_[3829]_  = ~\new_[4476]_  & (~\new_[8384]_  | ~\new_[8385]_ );
  assign \new_[3830]_  = ~\new_[4476]_  & (~\new_[8357]_  | ~\new_[8371]_ );
  assign \new_[3831]_  = ~\new_[13602]_  | ~\new_[4476]_ ;
  assign \new_[3832]_  = ~\new_[13416]_  | ~\new_[4476]_ ;
  assign \new_[3833]_  = ~\new_[13272]_  | ~\new_[4476]_ ;
  assign \new_[3834]_  = ~\new_[13259]_  | ~\new_[4476]_ ;
  assign \new_[3835]_  = ~\new_[13243]_  | ~\new_[4476]_ ;
  assign \new_[3836]_  = ~\new_[13230]_  | ~\new_[4476]_ ;
  assign \new_[3837]_  = ~\new_[13220]_  | ~\new_[4472]_ ;
  assign \new_[3838]_  = ~\new_[13207]_  | ~\new_[4472]_ ;
  assign \new_[3839]_  = ~\new_[13657]_  | ~\new_[4472]_ ;
  assign \new_[3840]_  = ~\new_[13579]_  | ~\new_[4472]_ ;
  assign \new_[3841]_  = ~\new_[13442]_  | ~\new_[4472]_ ;
  assign n3081 = \new_[8513]_  ? \new_[4517]_  : \new_[13241]_ ;
  assign \new_[3843]_  = ~\new_[13413]_  | ~\new_[4472]_ ;
  assign \new_[3844]_  = ~\new_[13415]_  | ~\new_[4472]_ ;
  assign \new_[3845]_  = ~\new_[13733]_  | ~\new_[4472]_ ;
  assign \new_[3846]_  = ~\new_[13855]_  | ~\new_[4472]_ ;
  assign \new_[3847]_  = ~\new_[13377]_  | ~\new_[4477]_ ;
  assign \new_[3848]_  = ~\new_[13339]_  | ~\new_[4472]_ ;
  assign \new_[3849]_  = ~\new_[13385]_  | ~\new_[4477]_ ;
  assign \new_[3850]_  = ~\new_[13665]_  | ~\new_[4477]_ ;
  assign \new_[3851]_  = ~\new_[4472]_  & (~\new_[8394]_  | ~\new_[8410]_ );
  assign \new_[3852]_  = ~\new_[13559]_  | ~\new_[4477]_ ;
  assign \new_[3853]_  = ~\new_[4472]_  & (~\new_[8397]_  | ~\new_[8398]_ );
  assign \new_[3854]_  = ~\new_[13449]_  | ~\new_[4477]_ ;
  assign \new_[3855]_  = ~\new_[13280]_  | ~\new_[4472]_ ;
  assign \new_[3856]_  = ~\new_[13391]_  | ~\new_[4477]_ ;
  assign \new_[3857]_  = ~\new_[13562]_  | ~\new_[4472]_ ;
  assign \new_[3858]_  = ~\new_[13552]_  | ~\new_[4477]_ ;
  assign \new_[3859]_  = ~\new_[13669]_  | ~\new_[4477]_ ;
  assign \new_[3860]_  = ~\new_[13548]_  | ~\new_[4472]_ ;
  assign \new_[3861]_  = ~\new_[13853]_  | ~\new_[4477]_ ;
  assign \new_[3862]_  = ~\new_[13771]_  | ~\new_[4472]_ ;
  assign \new_[3863]_  = ~\new_[13231]_  | ~\new_[4477]_ ;
  assign \new_[3864]_  = ~\new_[13299]_  | ~\new_[4472]_ ;
  assign \new_[3865]_  = ~\new_[4624]_  & (~\new_[8406]_  | ~\new_[8642]_ );
  assign \new_[3866]_  = ~\new_[4624]_  & (~\new_[8364]_  | ~\new_[8362]_ );
  assign \new_[3867]_  = ~\new_[13350]_  | ~\new_[4477]_ ;
  assign \new_[3868]_  = ~\new_[13264]_  | ~\new_[4477]_ ;
  assign \new_[3869]_  = ~\new_[13249]_  | ~\new_[4477]_ ;
  assign \new_[3870]_  = ~\new_[13585]_  | ~\new_[4477]_ ;
  assign \new_[3871]_  = ~\new_[13599]_  | ~\new_[4477]_ ;
  assign n3101 = \new_[8213]_  ? \new_[4517]_  : \new_[13590]_ ;
  assign n3076 = \new_[8214]_  ? \new_[4517]_  : \new_[13557]_ ;
  assign n3106 = \new_[8519]_  ? \new_[4517]_  : \new_[13856]_ ;
  assign n3086 = \new_[8234]_  ? \new_[4520]_  : \new_[13696]_ ;
  assign n3091 = \new_[8235]_  ? \new_[4520]_  : \new_[13751]_ ;
  assign n3096 = \new_[8236]_  ? \new_[4520]_  : \new_[13843]_ ;
  assign n3111 = \new_[8239]_  ? \new_[4520]_  : \new_[13423]_ ;
  assign n2646 = \new_[8241]_  ? \new_[4520]_  : \new_[13390]_ ;
  assign n3191 = \new_[8523]_  ? \new_[4520]_  : \new_[13741]_ ;
  assign n3116 = \new_[8242]_  ? \new_[4662]_  : \new_[13426]_ ;
  assign n3121 = \new_[8243]_  ? \new_[4662]_  : \new_[13430]_ ;
  assign n3126 = \new_[8245]_  ? \new_[4520]_  : \new_[13431]_ ;
  assign n3131 = \new_[8246]_  ? \new_[4520]_  : \new_[13367]_ ;
  assign n3136 = \new_[8224]_  ? \new_[4520]_  : \new_[13345]_ ;
  assign n2651 = \new_[8247]_  ? \new_[4520]_  : \new_[13510]_ ;
  assign n3141 = \new_[8223]_  ? \new_[4521]_  : \new_[13752]_ ;
  assign n3146 = \new_[8248]_  ? \new_[4521]_  : \new_[13440]_ ;
  assign n2641 = \new_[8525]_  ? \new_[4517]_  : \new_[13654]_ ;
  assign n3151 = \new_[8524]_  ? \new_[4520]_  : \new_[13645]_ ;
  assign n3156 = \new_[8249]_  ? \new_[4520]_  : \new_[13754]_ ;
  assign n3161 = \new_[8250]_  ? \new_[4521]_  : \new_[13646]_ ;
  assign n3166 = \new_[8252]_  ? \new_[4521]_  : \new_[13448]_ ;
  assign n3196 = \new_[8253]_  ? \new_[4521]_  : \new_[13840]_ ;
  assign \new_[3895]_  = ~\new_[4475]_  | (~\new_[7732]_  & ~\new_[7773]_ );
  assign n3171 = \new_[8178]_  ? \new_[4521]_  : \new_[13837]_ ;
  assign \new_[3897]_  = ~\new_[4475]_  | (~\new_[7733]_  & ~\new_[7775]_ );
  assign \new_[3898]_  = ~\new_[4475]_  | (~\new_[7734]_  & ~\new_[7776]_ );
  assign \new_[3899]_  = ~\new_[4475]_  | (~\new_[7672]_  & ~\new_[8024]_ );
  assign n3176 = \new_[8255]_  ? \new_[4521]_  : \new_[13664]_ ;
  assign \new_[3901]_  = ~\new_[4475]_  | (~\new_[7673]_  & ~\new_[7777]_ );
  assign \new_[3902]_  = ~\new_[4475]_  | (~\new_[7735]_  & ~\new_[7961]_ );
  assign \new_[3903]_  = ~\new_[4475]_  | (~\new_[7674]_  & ~\new_[7884]_ );
  assign \new_[3904]_  = ~\new_[4475]_  | (~\new_[7736]_  & ~\new_[7779]_ );
  assign \new_[3905]_  = ~\new_[4475]_  | (~\new_[7737]_  & ~\new_[7895]_ );
  assign \new_[3906]_  = ~\new_[4475]_  | (~\new_[7738]_  & ~\new_[7780]_ );
  assign n3181 = \new_[8257]_  ? \new_[4520]_  : \new_[13580]_ ;
  assign \new_[3908]_  = ~\new_[4475]_  | (~\new_[7739]_  & ~\new_[7781]_ );
  assign \new_[3909]_  = ~\new_[4475]_  | (~\new_[7675]_  & ~\new_[7896]_ );
  assign \new_[3910]_  = ~\new_[4475]_  | (~\new_[7676]_  & ~\new_[7981]_ );
  assign \new_[3911]_  = ~\new_[4475]_  | (~\new_[7677]_  & ~\new_[7982]_ );
  assign \new_[3912]_  = ~\new_[4475]_  | (~\new_[7741]_  & ~\new_[7983]_ );
  assign n3186 = \new_[8521]_  ? \new_[4520]_  : \new_[13627]_ ;
  assign \new_[3914]_  = ~\new_[4475]_  | (~\new_[7742]_  & ~\new_[7782]_ );
  assign \new_[3915]_  = ~\new_[4473]_  | (~\new_[7722]_  & ~\new_[7873]_ );
  assign n3201 = \new_[8262]_  ? \new_[4520]_  : \new_[13556]_ ;
  assign \new_[3917]_  = ~\new_[4473]_  | (~\new_[7752]_  & ~\new_[7905]_ );
  assign \new_[3918]_  = ~\new_[14161]_  | (~\new_[7753]_  & ~\new_[7906]_ );
  assign n3206 = \new_[8263]_  ? \new_[4520]_  : \new_[13476]_ ;
  assign n3216 = \new_[8265]_  ? \new_[4520]_  : \new_[13623]_ ;
  assign \new_[3921]_  = ~\new_[4473]_  | (~\new_[7754]_  & ~\new_[7908]_ );
  assign \new_[3922]_  = ~\new_[4478]_  | (~\new_[7755]_  & ~\new_[7985]_ );
  assign n3221 = \new_[8266]_  ? \new_[4520]_  : \new_[13768]_ ;
  assign \new_[3924]_  = ~\new_[4473]_  | (~\new_[7756]_  & ~\new_[7909]_ );
  assign \new_[3925]_  = ~\new_[4478]_  | (~\new_[7848]_  & ~\new_[7910]_ );
  assign \new_[3926]_  = ~\new_[4478]_  | (~\new_[7849]_  & ~\new_[7911]_ );
  assign n3211 = \new_[8267]_  ? \new_[4520]_  : \new_[13772]_ ;
  assign \new_[3928]_  = ~\new_[4478]_  | (~\new_[7757]_  & ~\new_[7986]_ );
  assign \new_[3929]_  = ~\new_[4478]_  | (~\new_[7847]_  & ~\new_[7907]_ );
  assign \new_[3930]_  = ~\new_[4473]_  | (~\new_[7758]_  & ~\new_[7912]_ );
  assign \new_[3931]_  = ~\new_[4478]_  | (~\new_[7850]_  & ~\new_[7987]_ );
  assign \new_[3932]_  = ~\new_[4473]_  | (~\new_[7743]_  & ~\new_[13904]_ );
  assign \new_[3933]_  = ~\new_[4478]_  | (~\new_[7759]_  & ~\new_[7913]_ );
  assign \new_[3934]_  = ~\new_[4478]_  | (~\new_[7851]_  & ~\new_[7988]_ );
  assign \new_[3935]_  = ~\new_[14161]_  | (~\new_[7760]_  & ~\new_[7914]_ );
  assign \new_[3936]_  = ~\new_[14161]_  | (~\new_[7761]_  & ~\new_[7915]_ );
  assign n3226 = \new_[8531]_  ? \new_[4521]_  : \new_[13660]_ ;
  assign \new_[3938]_  = ~\new_[4478]_  | (~\new_[7846]_  & ~\new_[7916]_ );
  assign \new_[3939]_  = ~\new_[4473]_  | (~\new_[7762]_  & ~\new_[7917]_ );
  assign \new_[3940]_  = ~\new_[4478]_  | (~\new_[7852]_  & ~\new_[7989]_ );
  assign n2631 = \new_[8221]_  ? \new_[4521]_  : \new_[13631]_ ;
  assign \new_[3942]_  = ~\new_[4473]_  | (~\new_[7763]_  & ~\new_[7918]_ );
  assign \new_[3943]_  = ~\new_[4478]_  | (~\new_[7764]_  & ~\new_[7919]_ );
  assign \new_[3944]_  = ~\new_[4478]_  | (~\new_[7765]_  & ~\new_[7920]_ );
  assign n3246 = \new_[8269]_  ? \new_[4521]_  : \new_[13684]_ ;
  assign \new_[3946]_  = ~\new_[4478]_  | (~\new_[7766]_  & ~\new_[7990]_ );
  assign \new_[3947]_  = ~\new_[4478]_  | (~\new_[7719]_  & ~\new_[7991]_ );
  assign \new_[3948]_  = ~\new_[4478]_  | (~\new_[7795]_  & ~\new_[7992]_ );
  assign n3231 = \new_[8270]_  ? \new_[4521]_  : \new_[13782]_ ;
  assign \new_[3950]_  = ~\new_[4478]_  | (~\new_[7854]_  & ~\new_[7921]_ );
  assign n3236 = \new_[8205]_  ? \new_[4521]_  : \new_[13814]_ ;
  assign n2636 = \new_[8271]_  ? \new_[4521]_  : \new_[13807]_ ;
  assign n2626 = \new_[8272]_  ? \new_[4521]_  : \new_[13630]_ ;
  assign n3241 = \new_[8273]_  ? \new_[4521]_  : \new_[13662]_ ;
  assign n3266 = \new_[8276]_  ? \new_[4520]_  : \new_[13635]_ ;
  assign n3251 = \new_[8233]_  ? \new_[4520]_  : \new_[13265]_ ;
  assign n3256 = \new_[8274]_  ? \new_[4520]_  : \new_[13821]_ ;
  assign n3261 = \new_[8264]_  ? \new_[4520]_  : \new_[13351]_ ;
  assign n3296 = \new_[8291]_  ? \new_[4519]_  : \new_[13533]_ ;
  assign n3291 = \new_[8292]_  ? \new_[4519]_  : \new_[13213]_ ;
  assign \new_[3961]_  = \\u20_int_set_reg[0] ;
  assign \new_[3962]_  = \\u18_int_set_reg[0] ;
  assign n3301 = \new_[8538]_  ? \new_[4520]_  : \new_[13464]_ ;
  assign n3456 = \new_[8539]_  ? \new_[4520]_  : \new_[13567]_ ;
  assign n3451 = \new_[8540]_  ? \new_[4519]_  : \new_[13817]_ ;
  assign n3306 = \new_[8772]_  ? \new_[4520]_  : \new_[13716]_ ;
  assign n3311 = \new_[8767]_  ? \new_[4521]_  : \new_[13594]_ ;
  assign n3316 = \new_[8773]_  ? \new_[4521]_  : \new_[13808]_ ;
  assign n3321 = \new_[8774]_  ? \new_[4662]_  : \new_[13596]_ ;
  assign n3326 = \new_[8765]_  ? \new_[4662]_  : \new_[13836]_ ;
  assign n3331 = \new_[8775]_  ? \new_[4521]_  : \new_[13262]_ ;
  assign n3336 = \new_[8975]_  ? \new_[4661]_  : \new_[13732]_ ;
  assign n3341 = \new_[8776]_  ? \new_[4521]_  : \new_[13323]_ ;
  assign n3346 = \new_[8769]_  ? \new_[4520]_  : \new_[13706]_ ;
  assign n3351 = \new_[8768]_  ? \new_[4661]_  : \new_[13472]_ ;
  assign n3356 = \new_[8781]_  ? \new_[4520]_  : \new_[13291]_ ;
  assign n3361 = \new_[8771]_  ? \new_[4521]_  : \new_[13641]_ ;
  assign n3366 = \new_[8301]_  ? \new_[4521]_  : \new_[13748]_ ;
  assign n3371 = \new_[8778]_  ? \new_[4520]_  : \new_[13702]_ ;
  assign n3376 = \new_[8770]_  ? \new_[4520]_  : \new_[13475]_ ;
  assign n3386 = \new_[8780]_  ? \new_[4661]_  : \new_[13488]_ ;
  assign n3381 = \new_[8302]_  ? \new_[4520]_  : \new_[13412]_ ;
  assign n3391 = \new_[8303]_  ? \new_[4520]_  : \new_[13834]_ ;
  assign n3396 = \new_[8976]_  ? \new_[4661]_  : \new_[13610]_ ;
  assign n3286 = \new_[8304]_  ? \new_[4521]_  : \new_[13490]_ ;
  assign n3401 = \new_[8977]_  ? \new_[4661]_  : \new_[13735]_ ;
  assign n3406 = \new_[8305]_  ? \new_[4521]_  : \new_[13266]_ ;
  assign n3411 = \new_[8978]_  ? \new_[4661]_  : \new_[13393]_ ;
  assign n3416 = \new_[8306]_  ? \new_[4521]_  : \new_[13719]_ ;
  assign n3421 = \new_[8307]_  ? \new_[4521]_  : \new_[13778]_ ;
  assign n3426 = \new_[8784]_  ? \new_[4517]_  : \new_[13288]_ ;
  assign n3431 = \new_[8541]_  ? \new_[4521]_  : \new_[13731]_ ;
  assign n3281 = \new_[8308]_  ? \new_[4517]_  : \new_[13466]_ ;
  assign n3436 = \new_[8311]_  ? \new_[4517]_  : \new_[13607]_ ;
  assign \new_[3995]_  = ~\new_[4282]_  & (~\new_[4786]_  | ~\new_[12765]_ );
  assign \new_[3996]_  = ~\new_[4283]_  & (~\new_[4788]_  | ~\new_[12632]_ );
  assign \new_[3997]_  = ~\new_[4284]_  & (~\new_[4790]_  | ~\new_[12772]_ );
  assign \new_[3998]_  = ~\new_[4285]_  & (~\new_[4791]_  | ~\new_[12865]_ );
  assign \new_[3999]_  = ~\new_[4287]_  & (~\new_[13902]_  | ~\new_[12896]_ );
  assign \new_[4000]_  = ~\new_[4300]_  & (~\new_[14001]_  | ~\new_[12623]_ );
  assign \new_[4001]_  = ~\new_[4366]_  & (~\new_[13900]_  | ~\new_[13870]_ );
  assign \new_[4002]_  = ~\new_[4367]_  & (~\new_[13898]_  | ~\new_[12549]_ );
  assign \new_[4003]_  = ~\new_[4508]_  | (~\new_[4782]_  & ~\new_[12744]_ );
  assign \new_[4004]_  = ~\new_[4509]_  | (~\new_[4783]_  & ~\new_[13052]_ );
  assign n4316 = ~\new_[4539]_  & ~\new_[8829]_ ;
  assign \new_[4006]_  = ~\new_[12350]_  | ~\new_[14097]_ ;
  assign \new_[4007]_  = ~\new_[12010]_  | ~\new_[4515]_ ;
  assign \new_[4008]_  = ~\new_[12012]_  | ~\new_[4527]_ ;
  assign \new_[4009]_  = ~\new_[12013]_  | ~\new_[4528]_ ;
  assign n3996 = \new_[4506]_  & \new_[13866]_ ;
  assign \new_[4011]_  = ~\new_[13332]_  | ~\new_[4522]_ ;
  assign \new_[4012]_  = ~\new_[13359]_  | ~\new_[4522]_ ;
  assign \new_[4013]_  = ~\new_[13522]_  | ~\new_[4522]_ ;
  assign \new_[4014]_  = ~\new_[13341]_  | ~\new_[4522]_ ;
  assign \new_[4015]_  = ~\new_[13838]_  | ~\new_[4525]_ ;
  assign \new_[4016]_  = ~\new_[13303]_  | ~\new_[4525]_ ;
  assign \new_[4017]_  = ~\new_[13287]_  | ~\new_[4525]_ ;
  assign \new_[4018]_  = ~\new_[13282]_  | ~\new_[4522]_ ;
  assign \new_[4019]_  = ~\new_[13261]_  | ~\new_[4522]_ ;
  assign \new_[4020]_  = ~\new_[13245]_  | ~\new_[4525]_ ;
  assign \new_[4021]_  = ~\new_[13239]_  | ~\new_[4524]_ ;
  assign \new_[4022]_  = ~\new_[13295]_  | ~\new_[4525]_ ;
  assign \new_[4023]_  = ~\new_[13211]_  | ~\new_[4524]_ ;
  assign \new_[4024]_  = ~\new_[13196]_  | ~\new_[4524]_ ;
  assign \new_[4025]_  = ~\new_[13242]_  | ~\new_[4525]_ ;
  assign \new_[4026]_  = ~\new_[13865]_  | ~\new_[4525]_ ;
  assign \new_[4027]_  = ~\new_[13705]_  | ~\new_[4522]_ ;
  assign \new_[4028]_  = ~\new_[13402]_  | ~\new_[4522]_ ;
  assign \new_[4029]_  = ~\new_[13773]_  | ~\new_[4525]_ ;
  assign \new_[4030]_  = ~\new_[13859]_  | ~\new_[4524]_ ;
  assign \new_[4031]_  = ~\new_[13419]_  | ~\new_[4524]_ ;
  assign \new_[4032]_  = ~\new_[13422]_  | ~\new_[4524]_ ;
  assign \new_[4033]_  = ~\new_[13424]_  | ~\new_[4524]_ ;
  assign \new_[4034]_  = ~\new_[13435]_  | ~\new_[4525]_ ;
  assign \new_[4035]_  = ~\new_[13389]_  | ~\new_[4524]_ ;
  assign \new_[4036]_  = ~\new_[13495]_  | ~\new_[4524]_ ;
  assign \new_[4037]_  = ~\new_[13588]_  | ~\new_[4525]_ ;
  assign \new_[4038]_  = ~\new_[13708]_  | ~\new_[4524]_ ;
  assign \new_[4039]_  = ~\new_[13587]_  | ~\new_[4524]_ ;
  assign \new_[4040]_  = ~\new_[13712]_  | ~\new_[4524]_ ;
  assign \new_[4041]_  = ~\new_[13593]_  | ~\new_[4522]_ ;
  assign \new_[4042]_  = ~\new_[13694]_  | ~\new_[4522]_ ;
  assign \new_[4043]_  = ~\new_[13616]_  | ~\new_[4525]_ ;
  assign \new_[4044]_  = ~\new_[13860]_  | ~\new_[4525]_ ;
  assign \new_[4045]_  = ~\new_[13763]_  | ~\new_[4525]_ ;
  assign \new_[4046]_  = ~\new_[13847]_  | ~\new_[4522]_ ;
  assign \new_[4047]_  = ~\new_[13258]_  | ~\new_[4524]_ ;
  assign \new_[4048]_  = ~\new_[13252]_  | ~\new_[4524]_ ;
  assign \new_[4049]_  = ~\new_[13427]_  | ~\new_[4524]_ ;
  assign \new_[4050]_  = ~\new_[13776]_  | ~\new_[4524]_ ;
  assign \new_[4051]_  = ~\new_[13764]_  | ~\new_[4525]_ ;
  assign \new_[4052]_  = ~\new_[13204]_  | ~\new_[4522]_ ;
  assign \new_[4053]_  = ~\new_[13238]_  | ~\new_[4525]_ ;
  assign \new_[4054]_  = ~\new_[13849]_  | ~\new_[4525]_ ;
  assign n4296 = ~\new_[4387]_ ;
  assign n4301 = ~\new_[4388]_ ;
  assign n4306 = ~\new_[4390]_ ;
  assign \new_[4058]_  = ~\new_[13571]_  & (~\new_[4709]_  | ~\new_[8503]_ );
  assign \new_[4059]_  = ~\new_[4511]_  | (~\new_[9648]_  & ~\new_[4778]_ );
  assign n3466 = \\u1_sr_reg[14] ;
  assign n4311 = ~\new_[4546]_  | (~\new_[5055]_  & ~\new_[6562]_ );
  assign \new_[4062]_  = \new_[3081]_  ? \new_[4709]_  : \new_[10314]_ ;
  assign \new_[4063]_  = ~\new_[4512]_  | (~\new_[8790]_  & ~\new_[4778]_ );
  assign n3481 = \new_[4507]_  & \new_[13866]_ ;
  assign n4216 = ~\new_[4503]_  | ~\new_[4516]_ ;
  assign \new_[4066]_  = ~\new_[4606]_  | ~\new_[13929]_  | ~\new_[13977]_ ;
  assign \new_[4067]_  = ~\new_[4607]_  | ~\new_[13973]_  | ~\new_[12019]_ ;
  assign \new_[4068]_  = \\u13_ints_r_reg[23] ;
  assign \new_[4069]_  = \\u13_ints_r_reg[20] ;
  assign \new_[4070]_  = \\u9_wp_reg[1] ;
  assign \new_[4071]_  = \\u9_din_tmp1_reg[9] ;
  assign \new_[4072]_  = \\u9_din_tmp1_reg[3] ;
  assign \new_[4073]_  = \\u9_din_tmp1_reg[10] ;
  assign \new_[4074]_  = \\u9_din_tmp1_reg[14] ;
  assign \new_[4075]_  = \\u9_din_tmp1_reg[0] ;
  assign \new_[4076]_  = \\u9_din_tmp1_reg[11] ;
  assign \new_[4077]_  = \\u9_din_tmp1_reg[12] ;
  assign \new_[4078]_  = \\u9_din_tmp1_reg[13] ;
  assign \new_[4079]_  = \\u9_din_tmp1_reg[15] ;
  assign \new_[4080]_  = \\u9_din_tmp1_reg[1] ;
  assign \new_[4081]_  = \\u9_din_tmp1_reg[2] ;
  assign \new_[4082]_  = \\u9_din_tmp1_reg[5] ;
  assign \new_[4083]_  = \\u9_din_tmp1_reg[6] ;
  assign \new_[4084]_  = \\u9_din_tmp1_reg[4] ;
  assign \new_[4085]_  = \\u9_din_tmp1_reg[8] ;
  assign \new_[4086]_  = \\u9_din_tmp1_reg[7] ;
  assign \new_[4087]_  = u15_rdd3_reg;
  assign \new_[4088]_  = \new_[2791]_  ? \new_[4606]_  : \new_[8980]_ ;
  assign \new_[4089]_  = \new_[2793]_  ? \new_[4607]_  : \new_[9813]_ ;
  assign n3601 = \new_[8520]_  ? \new_[4608]_  : \new_[13603]_ ;
  assign n3636 = \new_[8203]_  ? \new_[4608]_  : \new_[13750]_ ;
  assign n3606 = \new_[8179]_  ? \new_[4608]_  : \new_[13273]_ ;
  assign n3611 = \new_[8180]_  ? \new_[4608]_  : \new_[13711]_ ;
  assign n3616 = \new_[8181]_  ? \new_[4608]_  : \new_[13414]_ ;
  assign n3621 = \new_[8182]_  ? \new_[4609]_  : \new_[13766]_ ;
  assign n3626 = \new_[8183]_  ? \new_[4608]_  : \new_[13232]_ ;
  assign n3631 = \new_[8506]_  ? \new_[4609]_  : \new_[13792]_ ;
  assign n4011 = \new_[8507]_  ? \new_[4609]_  : \new_[13347]_ ;
  assign n3641 = \new_[8008]_  ? \new_[4600]_  : \new_[13583]_ ;
  assign n3646 = \new_[8185]_  ? \new_[4600]_  : \new_[13514]_ ;
  assign n4006 = \new_[8222]_  ? \new_[4603]_  : \new_[13494]_ ;
  assign n3651 = \new_[8226]_  ? \new_[4596]_  : \new_[13318]_ ;
  assign n3656 = \new_[8229]_  ? \new_[4596]_  : \new_[13675]_ ;
  assign n3661 = \new_[8186]_  ? \new_[4601]_  : \new_[13577]_ ;
  assign n4001 = \new_[8231]_  ? \new_[4596]_  : \new_[13294]_ ;
  assign n3666 = \new_[8036]_  ? \new_[4604]_  : \new_[13628]_ ;
  assign n3671 = \new_[8009]_  ? \new_[4604]_  : \new_[13409]_ ;
  assign n3676 = \new_[8011]_  ? \new_[4601]_  : \new_[13819]_ ;
  assign n3986 = \new_[8187]_  ? \new_[4609]_  : \new_[13722]_ ;
  assign n3681 = \new_[8038]_  ? \new_[4601]_  : \new_[13436]_ ;
  assign n3686 = \new_[8012]_  ? \new_[4596]_  : \new_[13638]_ ;
  assign n3691 = \new_[8039]_  ? \new_[4596]_  : \new_[13439]_ ;
  assign n3696 = \new_[8013]_  ? \new_[4596]_  : \new_[13845]_ ;
  assign n3701 = \new_[8014]_  ? \new_[4596]_  : \new_[13420]_ ;
  assign n3706 = \new_[8015]_  ? \new_[4601]_  : \new_[13246]_ ;
  assign n3711 = \new_[8227]_  ? \new_[4601]_  : \new_[13717]_ ;
  assign n3961 = \new_[8016]_  ? \new_[4603]_  : \new_[13453]_ ;
  assign n3716 = \new_[8041]_  ? \new_[4601]_  : \new_[13663]_ ;
  assign n3721 = \new_[8189]_  ? \new_[4600]_  : \new_[13586]_ ;
  assign n3726 = \new_[8190]_  ? \new_[4600]_  : \new_[13284]_ ;
  assign n3556 = \new_[8244]_  ? \new_[4600]_  : \new_[13854]_ ;
  assign n3821 = \new_[8191]_  ? \new_[4603]_  : \new_[13621]_ ;
  assign n3731 = \new_[8192]_  ? \new_[4603]_  : \new_[13679]_ ;
  assign n3736 = \new_[8193]_  ? \new_[4603]_  : \new_[13257]_ ;
  assign n3741 = \new_[8040]_  ? \new_[4603]_  : \new_[13333]_ ;
  assign n3746 = \new_[8017]_  ? \new_[4602]_  : \new_[13830]_ ;
  assign n3751 = \new_[8037]_  ? \new_[4602]_  : \new_[13521]_ ;
  assign n3756 = \new_[8194]_  ? \new_[4608]_  : \new_[13858]_ ;
  assign n3591 = \new_[8018]_  ? \new_[4602]_  : \new_[13406]_ ;
  assign n3766 = \new_[8195]_  ? \new_[4608]_  : \new_[13553]_ ;
  assign n3761 = \new_[8034]_  ? \new_[4602]_  : \new_[13542]_ ;
  assign n3771 = \new_[8019]_  ? \new_[4600]_  : \new_[13544]_ ;
  assign n3586 = \new_[8029]_  ? \new_[4600]_  : \new_[13499]_ ;
  assign n3776 = \new_[8030]_  ? \new_[4603]_  : \new_[13310]_ ;
  assign n3781 = \new_[8020]_  ? \new_[4603]_  : \new_[13591]_ ;
  assign n3786 = \new_[8196]_  ? \new_[4603]_  : \new_[13713]_ ;
  assign n4291 = \new_[8032]_  ? \new_[4602]_  : \new_[13699]_ ;
  assign n3791 = \new_[8021]_  ? \new_[4602]_  : \new_[13800]_ ;
  assign n3796 = \new_[8199]_  ? \new_[4595]_  : \new_[13362]_ ;
  assign n3801 = \new_[8200]_  ? \new_[4595]_  : \new_[13468]_ ;
  assign n3806 = \new_[8201]_  ? \new_[4600]_  : \new_[13328]_ ;
  assign n3811 = \new_[8261]_  ? \new_[4600]_  : \new_[13327]_ ;
  assign n3816 = \new_[8240]_  ? \new_[4595]_  : \new_[13329]_ ;
  assign \new_[4144]_  = ~\new_[4623]_  | ~\new_[12993]_ ;
  assign n3581 = \new_[8212]_  ? \new_[4595]_  : \new_[13528]_ ;
  assign n3826 = \new_[8022]_  ? \new_[4600]_  : \new_[13690]_ ;
  assign n3831 = \new_[8010]_  ? \new_[4600]_  : \new_[13346]_ ;
  assign n3576 = \new_[8023]_  ? \new_[4601]_  : \new_[13512]_ ;
  assign n3836 = \new_[8204]_  ? \new_[4609]_  : \new_[13340]_ ;
  assign n3841 = \new_[8025]_  ? \new_[4601]_  : \new_[13746]_ ;
  assign \new_[4151]_  = ~\new_[4476]_  | ~\new_[12686]_ ;
  assign n3846 = \new_[8033]_  ? \new_[4602]_  : \new_[13290]_ ;
  assign n3866 = \new_[8512]_  ? \new_[4609]_  : \new_[13263]_ ;
  assign n3571 = \new_[8031]_  ? \new_[4602]_  : \new_[13216]_ ;
  assign n3851 = \new_[8026]_  ? \new_[4596]_  : \new_[13268]_ ;
  assign n3856 = \new_[8035]_  ? \new_[4596]_  : \new_[13386]_ ;
  assign \new_[4157]_  = ~\new_[14162]_  | ~\new_[13012]_ ;
  assign n3861 = \new_[8027]_  ? \new_[4601]_  : \new_[13637]_ ;
  assign n3876 = \new_[8219]_  ? \new_[4600]_  : \new_[13381]_ ;
  assign \new_[4160]_  = ~\new_[4624]_  | ~\new_[12519]_ ;
  assign n3871 = \new_[8028]_  ? \new_[4600]_  : \new_[13376]_ ;
  assign n3566 = \new_[8517]_  ? \new_[4608]_  : \new_[13233]_ ;
  assign n3881 = \new_[8206]_  ? \new_[4608]_  : \new_[13267]_ ;
  assign n3886 = \new_[8207]_  ? \new_[4608]_  : \new_[13226]_ ;
  assign n3891 = \new_[8208]_  ? \new_[4608]_  : \new_[13215]_ ;
  assign n3561 = \new_[8209]_  ? \new_[4706]_  : \new_[13443]_ ;
  assign n3896 = \new_[8210]_  ? \new_[4706]_  : \new_[13640]_ ;
  assign n3901 = \new_[8211]_  ? \new_[4706]_  : \new_[13644]_ ;
  assign n3906 = \new_[8514]_  ? \new_[4706]_  : \new_[13380]_ ;
  assign n3461 = \new_[8515]_  ? \new_[4608]_  : \new_[13691]_ ;
  assign n3911 = \new_[8516]_  ? \new_[4608]_  : \new_[13394]_ ;
  assign n3916 = \new_[8215]_  ? \new_[4608]_  : \new_[13536]_ ;
  assign n3921 = \new_[8216]_  ? \new_[4608]_  : \new_[13498]_ ;
  assign n3926 = \new_[8217]_  ? \new_[4608]_  : \new_[13487]_ ;
  assign n3931 = \new_[8218]_  ? \new_[4608]_  : \new_[13502]_ ;
  assign n3541 = \new_[8518]_  ? \new_[4608]_  : \new_[13411]_ ;
  assign n3536 = \new_[8251]_  ? \new_[4609]_  : \new_[13446]_ ;
  assign n3936 = \new_[8254]_  ? \new_[4609]_  : \new_[13224]_ ;
  assign n3941 = \new_[8256]_  ? \new_[4609]_  : \new_[13667]_ ;
  assign n3531 = \new_[8258]_  ? \new_[4609]_  : \new_[13760]_ ;
  assign \new_[4181]_  = ~\new_[13962]_  | (~\new_[14123]_  & ~\new_[7897]_ );
  assign \new_[4182]_  = ~\new_[13962]_  | (~\new_[14128]_  & ~\new_[7898]_ );
  assign \new_[4183]_  = ~\new_[14060]_  | (~\new_[7744]_  & ~\new_[7899]_ );
  assign n3946 = \new_[8228]_  ? \new_[4609]_  : \new_[13762]_ ;
  assign \new_[4185]_  = ~\new_[14060]_  | (~\new_[7740]_  & ~\new_[7900]_ );
  assign \new_[4186]_  = ~\new_[13962]_  | (~\new_[7745]_  & ~\new_[7901]_ );
  assign \new_[4187]_  = ~\new_[14060]_  | (~\new_[14049]_  & ~\new_[7902]_ );
  assign \new_[4188]_  = ~\new_[14060]_  | (~\new_[7746]_  & ~\new_[7783]_ );
  assign \new_[4189]_  = ~\new_[14060]_  | (~\new_[7747]_  & ~\new_[7784]_ );
  assign \new_[4190]_  = ~\new_[14060]_  | (~\new_[7748]_  & ~\new_[7785]_ );
  assign n3526 = \new_[8260]_  ? \new_[4609]_  : \new_[13786]_ ;
  assign \new_[4192]_  = ~\new_[14060]_  | (~\new_[7749]_  & ~\new_[7786]_ );
  assign n3956 = \new_[8528]_  ? \new_[4609]_  : \new_[13470]_ ;
  assign \new_[4194]_  = ~\new_[13962]_  | (~\new_[7767]_  & ~\new_[7903]_ );
  assign n3951 = \new_[8529]_  ? \new_[4609]_  : \new_[13687]_ ;
  assign \new_[4196]_  = ~\new_[13962]_  | (~\new_[7751]_  & ~\new_[7904]_ );
  assign \new_[4197]_  = ~\new_[13962]_  | (~\new_[7678]_  & ~\new_[7984]_ );
  assign n3521 = \new_[8530]_  ? \new_[4609]_  : \new_[13473]_ ;
  assign n3981 = \new_[8232]_  ? \new_[4609]_  : \new_[13397]_ ;
  assign n3966 = \new_[8275]_  ? \new_[4608]_  : \new_[13784]_ ;
  assign n3971 = \new_[8225]_  ? \new_[4608]_  : \new_[13195]_ ;
  assign n3976 = \new_[8277]_  ? \new_[4608]_  : \new_[13250]_ ;
  assign n3506 = \new_[8278]_  ? \new_[4608]_  : \new_[13513]_ ;
  assign n3991 = \new_[8279]_  ? \new_[4609]_  : \new_[13653]_ ;
  assign n3491 = \new_[8532]_  ? \new_[4609]_  : \new_[13276]_ ;
  assign n3596 = \new_[8504]_  ? \new_[4609]_  : \new_[13759]_ ;
  assign n4036 = \new_[8042]_  ? \new_[4596]_  : \new_[13479]_ ;
  assign n4041 = \new_[8280]_  ? \new_[4596]_  : \new_[13312]_ ;
  assign n4046 = \new_[8281]_  ? \new_[4596]_  : \new_[13410]_ ;
  assign n4051 = \new_[8282]_  ? \new_[4601]_  : \new_[13527]_ ;
  assign n3516 = \new_[8286]_  ? \new_[4601]_  : \new_[13222]_ ;
  assign n4056 = \new_[8283]_  ? \new_[4600]_  : \new_[13256]_ ;
  assign n4061 = \new_[8284]_  ? \new_[4600]_  : \new_[13356]_ ;
  assign n4066 = \new_[8043]_  ? \new_[4604]_  : \new_[13517]_ ;
  assign n3511 = \new_[8044]_  ? \new_[4604]_  : \new_[13848]_ ;
  assign n4071 = \new_[8045]_  ? \new_[4601]_  : \new_[13432]_ ;
  assign n4076 = \new_[8965]_  ? \new_[4601]_  : \new_[13851]_ ;
  assign n4081 = \new_[8966]_  ? \new_[4604]_  : \new_[13852]_ ;
  assign n4086 = \new_[8979]_  ? \new_[4604]_  : \new_[13203]_ ;
  assign n4091 = \new_[8967]_  ? \new_[4596]_  : \new_[13785]_ ;
  assign n4096 = \new_[8968]_  ? \new_[4596]_  : \new_[13636]_ ;
  assign n4101 = \new_[8969]_  ? \new_[4604]_  : \new_[13491]_ ;
  assign n3501 = \new_[8970]_  ? \new_[4604]_  : \new_[13418]_ ;
  assign n4106 = \new_[8971]_  ? \new_[4596]_  : \new_[13349]_ ;
  assign n4111 = \new_[8972]_  ? \new_[4596]_  : \new_[13581]_ ;
  assign n4116 = \new_[8973]_  ? \new_[4603]_  : \new_[13659]_ ;
  assign n3496 = \new_[8046]_  ? \new_[4603]_  : \new_[13504]_ ;
  assign n4121 = \new_[8974]_  ? \new_[4603]_  : \new_[13503]_ ;
  assign n4126 = \new_[8964]_  ? \new_[4603]_  : \new_[13484]_ ;
  assign n4131 = \new_[8047]_  ? \new_[4603]_  : \new_[13774]_ ;
  assign n3476 = \new_[8048]_  ? \new_[4603]_  : \new_[13485]_ ;
  assign n4136 = \new_[8049]_  ? \new_[4603]_  : \new_[13400]_ ;
  assign n4141 = \new_[8050]_  ? \new_[4601]_  : \new_[13842]_ ;
  assign n4146 = \new_[8051]_  ? \new_[4601]_  : \new_[13202]_ ;
  assign n3486 = \new_[8285]_  ? \new_[4601]_  : \new_[13497]_ ;
  assign n4151 = \new_[8052]_  ? \new_[4600]_  : \new_[13862]_ ;
  assign \new_[4237]_  = ~\new_[4504]_  | (~\new_[4658]_  & ~\new_[3023]_ );
  assign \new_[4238]_  = ~\new_[4505]_  | (~\new_[4659]_  & ~\new_[13075]_ );
  assign n4156 = \new_[8535]_  ? \new_[4608]_  : \new_[13864]_ ;
  assign n4161 = \new_[8289]_  ? \new_[4608]_  : \new_[13355]_ ;
  assign n3471 = \new_[8290]_  ? \new_[4608]_  : \new_[13296]_ ;
  assign n4166 = \new_[8294]_  ? \new_[4609]_  : \new_[13524]_ ;
  assign n4171 = \new_[8287]_  ? \new_[4609]_  : \new_[13530]_ ;
  assign n4176 = \new_[8536]_  ? \new_[4609]_  : \new_[13831]_ ;
  assign \new_[4245]_  = \\u21_int_set_reg[0] ;
  assign \new_[4246]_  = \\u22_int_set_reg[0] ;
  assign \new_[4247]_  = \\u17_int_set_reg[0] ;
  assign n4181 = \new_[8537]_  ? \new_[4609]_  : \new_[13565]_ ;
  assign \new_[4249]_  = \\u19_int_set_reg[0] ;
  assign n4321 = \new_[8766]_  ? \new_[4609]_  : \new_[13841]_ ;
  assign n3546 = \new_[8777]_  ? \new_[4608]_  : \new_[13725]_ ;
  assign n4016 = \new_[8779]_  ? \new_[4608]_  : \new_[13205]_ ;
  assign n4196 = \new_[8782]_  ? \new_[4609]_  : \new_[13373]_ ;
  assign n4186 = \new_[8783]_  ? \new_[4609]_  : \new_[13336]_ ;
  assign n4191 = \new_[8309]_  ? \new_[4609]_  : \new_[13673]_ ;
  assign n4031 = \new_[8310]_  ? \new_[4609]_  : \new_[13625]_ ;
  assign n4201 = \new_[8313]_  ? \new_[4608]_  : \new_[13458]_ ;
  assign n4206 = \new_[8312]_  ? \new_[4608]_  : \new_[13221]_ ;
  assign n4026 = \new_[8542]_  ? \new_[4608]_  : \new_[13795]_ ;
  assign n4211 = \new_[8534]_  ? \new_[4608]_  : \new_[13793]_ ;
  assign n4221 = \new_[3588]_  ? \new_[4594]_  : \new_[7688]_ ;
  assign n4226 = \new_[3589]_  ? \new_[4594]_  : \new_[2924]_ ;
  assign n4231 = \new_[3590]_  ? \new_[4594]_  : \new_[2787]_ ;
  assign n4236 = \new_[3591]_  ? \new_[4594]_  : \new_[2749]_ ;
  assign n4241 = \new_[3592]_  ? \new_[4594]_  : \new_[2738]_ ;
  assign n4246 = \new_[3593]_  ? \new_[4594]_  : \new_[2727]_ ;
  assign n4251 = \new_[3594]_  ? \new_[4594]_  : \new_[2718]_ ;
  assign n4256 = \new_[3595]_  ? \new_[4594]_  : \new_[7503]_ ;
  assign n4261 = \new_[3596]_  ? \new_[4594]_  : \new_[6809]_ ;
  assign n4266 = \new_[3597]_  ? \new_[4594]_  : \new_[5888]_ ;
  assign n4021 = \new_[3546]_  ? \new_[4594]_  : \new_[4813]_ ;
  assign n4271 = \new_[3598]_  ? \new_[4594]_  : \new_[4720]_ ;
  assign n4276 = \new_[3599]_  ? \new_[4594]_  : \new_[4576]_ ;
  assign n4281 = \new_[3600]_  ? \new_[4594]_  : \new_[4410]_ ;
  assign n3551 = \new_[3449]_  ? \new_[4594]_  : \new_[3672]_ ;
  assign n4286 = \new_[3601]_  ? \new_[4594]_  : \new_[3185]_ ;
  assign \new_[4277]_  = \new_[12698]_  ^ \new_[4606]_ ;
  assign \new_[4278]_  = \new_[12994]_  ^ \new_[4607]_ ;
  assign \new_[4279]_  = u16_u8_dma_req_r1_reg;
  assign n4461 = ~\new_[4667]_  | ~\new_[4564]_  | ~\new_[4735]_ ;
  assign n4456 = ~\new_[4668]_  | ~\new_[4565]_  | ~\new_[4736]_ ;
  assign \new_[4282]_  = ~\new_[4575]_  | (~\new_[4924]_  & ~\new_[12750]_ );
  assign \new_[4283]_  = ~\new_[4577]_  | (~\new_[4925]_  & ~\new_[12770]_ );
  assign \new_[4284]_  = ~\new_[4579]_  | (~\new_[4926]_  & ~\new_[12752]_ );
  assign \new_[4285]_  = ~\new_[4580]_  | (~\new_[4927]_  & ~\new_[12737]_ );
  assign \new_[4286]_  = ~\new_[4778]_  | ~\new_[3340]_  | ~\new_[13876]_ ;
  assign \new_[4287]_  = ~\new_[13903]_  & ~\new_[12896]_ ;
  assign \new_[4288]_  = ~\new_[13277]_  | ~\new_[4610]_ ;
  assign n4341 = \new_[4574]_  & \new_[9077]_ ;
  assign \new_[4290]_  = ~\new_[13465]_  | ~\new_[4610]_ ;
  assign \new_[4291]_  = ~\new_[13753]_  | ~\new_[4610]_ ;
  assign \new_[4292]_  = ~\new_[13829]_  | ~\new_[4613]_ ;
  assign \new_[4293]_  = ~\new_[13805]_  | ~\new_[4613]_ ;
  assign \new_[4294]_  = ~\new_[13253]_  | ~\new_[4613]_ ;
  assign \new_[4295]_  = ~\new_[13279]_  | ~\new_[4704]_ ;
  assign \new_[4296]_  = ~\new_[13618]_  | ~\new_[4704]_ ;
  assign \new_[4297]_  = ~\new_[13861]_  | ~\new_[4612]_ ;
  assign \new_[4298]_  = ~\new_[13429]_  | ~\new_[4613]_ ;
  assign \new_[4299]_  = ~\new_[13237]_  | ~\new_[4613]_ ;
  assign \new_[4300]_  = ~\new_[14001]_  & ~\new_[12623]_ ;
  assign \new_[4301]_  = ~\new_[13634]_  | ~\new_[4613]_ ;
  assign \new_[4302]_  = ~\new_[13293]_  | ~\new_[4612]_ ;
  assign \new_[4303]_  = ~\new_[13558]_  | ~\new_[4597]_ ;
  assign \new_[4304]_  = ~\new_[13271]_  | ~\new_[4599]_ ;
  assign \new_[4305]_  = ~\new_[13417]_  | ~\new_[4599]_ ;
  assign \new_[4306]_  = ~\new_[13398]_  | ~\new_[4599]_ ;
  assign \new_[4307]_  = ~\new_[13302]_  | ~\new_[4599]_ ;
  assign \new_[4308]_  = ~\new_[13826]_  | ~\new_[4613]_ ;
  assign \new_[4309]_  = ~\new_[13825]_  | ~\new_[4599]_ ;
  assign \new_[4310]_  = ~\new_[13193]_  | ~\new_[4599]_ ;
  assign \new_[4311]_  = ~\new_[13568]_  | ~\new_[4599]_ ;
  assign \new_[4312]_  = ~\new_[13378]_  | ~\new_[4599]_ ;
  assign \new_[4313]_  = ~\new_[13555]_  | ~\new_[4599]_ ;
  assign \new_[4314]_  = ~\new_[13364]_  | ~\new_[4597]_ ;
  assign \new_[4315]_  = ~\new_[13452]_  | ~\new_[4599]_ ;
  assign \new_[4316]_  = ~\new_[13450]_  | ~\new_[4613]_ ;
  assign \new_[4317]_  = ~\new_[13368]_  | ~\new_[4613]_ ;
  assign \new_[4318]_  = ~\new_[13194]_  | ~\new_[4597]_ ;
  assign \new_[4319]_  = ~\new_[13681]_  | ~\new_[4597]_ ;
  assign \new_[4320]_  = ~\new_[13804]_  | ~\new_[4599]_ ;
  assign \new_[4321]_  = ~\new_[13835]_  | ~\new_[4599]_ ;
  assign \new_[4322]_  = ~\new_[13566]_  | ~\new_[4597]_ ;
  assign \new_[4323]_  = ~\new_[13401]_  | ~\new_[4597]_ ;
  assign \new_[4324]_  = ~\new_[13283]_  | ~\new_[4597]_ ;
  assign \new_[4325]_  = ~\new_[13254]_  | ~\new_[4597]_ ;
  assign \new_[4326]_  = ~\new_[13286]_  | ~\new_[4597]_ ;
  assign \new_[4327]_  = ~\new_[13289]_  | ~\new_[4599]_ ;
  assign \new_[4328]_  = ~\new_[13229]_  | ~\new_[4599]_ ;
  assign \new_[4329]_  = ~\new_[13227]_  | ~\new_[4599]_ ;
  assign \new_[4330]_  = ~\new_[13292]_  | ~\new_[4597]_ ;
  assign \new_[4331]_  = ~\new_[13670]_  | ~\new_[4597]_ ;
  assign \new_[4332]_  = ~\new_[13672]_  | ~\new_[4704]_ ;
  assign \new_[4333]_  = ~\new_[13633]_  | ~\new_[4703]_ ;
  assign \new_[4334]_  = ~\new_[13297]_  | ~\new_[4598]_ ;
  assign \new_[4335]_  = ~\new_[13298]_  | ~\new_[4703]_ ;
  assign \new_[4336]_  = ~\new_[13685]_  | ~\new_[4598]_ ;
  assign \new_[4337]_  = ~\new_[13301]_  | ~\new_[4598]_ ;
  assign \new_[4338]_  = ~\new_[13839]_  | ~\new_[4598]_ ;
  assign \new_[4339]_  = ~\new_[13305]_  | ~\new_[4598]_ ;
  assign \new_[4340]_  = ~\new_[13609]_  | ~\new_[4703]_ ;
  assign \new_[4341]_  = ~\new_[13307]_  | ~\new_[4703]_ ;
  assign \new_[4342]_  = ~\new_[13693]_  | ~\new_[4598]_ ;
  assign \new_[4343]_  = ~\new_[13309]_  | ~\new_[4598]_ ;
  assign \new_[4344]_  = ~\new_[13371]_  | ~\new_[4610]_ ;
  assign \new_[4345]_  = ~\new_[13311]_  | ~\new_[4610]_ ;
  assign \new_[4346]_  = ~\new_[13313]_  | ~\new_[4613]_ ;
  assign \new_[4347]_  = ~\new_[13578]_  | ~\new_[4610]_ ;
  assign \new_[4348]_  = ~\new_[13319]_  | ~\new_[4613]_ ;
  assign \new_[4349]_  = ~\new_[13572]_  | ~\new_[4612]_ ;
  assign \new_[4350]_  = ~\new_[13321]_  | ~\new_[4613]_ ;
  assign \new_[4351]_  = ~\new_[13363]_  | ~\new_[4613]_ ;
  assign \new_[4352]_  = ~\new_[13564]_  | ~\new_[4612]_ ;
  assign \new_[4353]_  = ~\new_[13325]_  | ~\new_[4613]_ ;
  assign \new_[4354]_  = ~\new_[13511]_  | ~\new_[4613]_ ;
  assign \new_[4355]_  = ~\new_[13560]_  | ~\new_[4613]_ ;
  assign \new_[4356]_  = ~\new_[13360]_  | ~\new_[4613]_ ;
  assign \new_[4357]_  = ~\new_[13549]_  | ~\new_[4613]_ ;
  assign \new_[4358]_  = \new_[4606]_  | \new_[13142]_ ;
  assign \new_[4359]_  = ~\new_[13374]_  | ~\new_[4598]_ ;
  assign \new_[4360]_  = \new_[4607]_  | \new_[13113]_ ;
  assign \new_[4361]_  = ~\new_[13781]_  | ~\new_[4597]_ ;
  assign \new_[4362]_  = ~\new_[13285]_  | ~\new_[4599]_ ;
  assign \new_[4363]_  = ~\new_[13357]_  | ~\new_[4610]_ ;
  assign \new_[4364]_  = ~\new_[13326]_  | ~\new_[4610]_ ;
  assign \new_[4365]_  = ~\new_[13516]_  | ~\new_[4704]_ ;
  assign \new_[4366]_  = ~\new_[13901]_  & ~\new_[13870]_ ;
  assign \new_[4367]_  = ~\new_[13899]_  & ~\new_[12549]_ ;
  assign \new_[4368]_  = ~\new_[13358]_  | ~\new_[4610]_ ;
  assign \new_[4369]_  = ~\new_[13755]_  | ~\new_[4610]_ ;
  assign \new_[4370]_  = ~\new_[13761]_  | ~\new_[4613]_ ;
  assign \new_[4371]_  = ~\new_[13474]_  | ~\new_[4613]_ ;
  assign \new_[4372]_  = ~\new_[13765]_  | ~\new_[4613]_ ;
  assign \new_[4373]_  = ~\new_[13501]_  | ~\new_[4610]_ ;
  assign \new_[4374]_  = ~\new_[13787]_  | ~\new_[4612]_ ;
  assign \new_[4375]_  = ~\new_[13676]_  | ~\new_[4613]_ ;
  assign \new_[4376]_  = ~\new_[13668]_  | ~\new_[4612]_ ;
  assign \new_[4377]_  = ~\new_[13678]_  | ~\new_[4612]_ ;
  assign \new_[4378]_  = ~\new_[13535]_  | ~\new_[4610]_ ;
  assign \new_[4379]_  = ~\new_[13438]_  | ~\new_[4612]_ ;
  assign \new_[4380]_  = ~\new_[13576]_  | ~\new_[4613]_ ;
  assign \new_[4381]_  = ~\new_[13649]_  | ~\new_[4613]_ ;
  assign \new_[4382]_  = ~\new_[13903]_  & (~\new_[11625]_  | ~\new_[10487]_ );
  assign \new_[4383]_  = ~\new_[14001]_  & (~\new_[11147]_  | ~\new_[10868]_ );
  assign \new_[4384]_  = ~\new_[12886]_  | ~\new_[14081]_  | ~\new_[13955]_ ;
  assign \new_[4385]_  = ~\new_[12691]_  | ~\new_[12501]_  | ~\new_[14107]_ ;
  assign \new_[4386]_  = \\u1_slt4_reg[11] ;
  assign \new_[4387]_  = ~\new_[13199]_  & (~\new_[6560]_  | ~\new_[13955]_ );
  assign \new_[4388]_  = ~\new_[13815]_  & (~\new_[6831]_  | ~\new_[14106]_ );
  assign \new_[4389]_  = ~\new_[13901]_  & (~\new_[11631]_  | ~\new_[10809]_ );
  assign \new_[4390]_  = ~\new_[13322]_  & (~\new_[4781]_  | ~\new_[8995]_ );
  assign \new_[4391]_  = ~\new_[13899]_  & (~\new_[12307]_  | ~\new_[11679]_ );
  assign \new_[4392]_  = ~\new_[13903]_  & (~\new_[12267]_  | ~\new_[13995]_ );
  assign \new_[4393]_  = ~\new_[14001]_  & (~\new_[11523]_  | ~\new_[12016]_ );
  assign \new_[4394]_  = ~\new_[4592]_  | (~\new_[8998]_  & ~\new_[4887]_ );
  assign \new_[4395]_  = ~\new_[13901]_  & (~\new_[12534]_  | ~\new_[12437]_ );
  assign \new_[4396]_  = ~\new_[13899]_  & (~\new_[14137]_  | ~\new_[12021]_ );
  assign \new_[4397]_  = \new_[12991]_  ? \new_[4781]_  : \new_[9090]_ ;
  assign \new_[4398]_  = ~\new_[4593]_  | (~\new_[8485]_  & ~\new_[4887]_ );
  assign n4346 = \new_[3761]_  ? \new_[9006]_  : n4646;
  assign n4351 = n4646 ? \new_[8996]_  : \new_[3762]_ ;
  assign n4356 = n4646 ? \new_[9002]_  : \new_[3763]_ ;
  assign n4361 = n4646 ? \new_[9000]_  : \new_[3764]_ ;
  assign n4336 = n4646 ? \new_[9001]_  : \new_[3672]_ ;
  assign n4326 = \new_[13361]_  ? \new_[7937]_  : \new_[4629]_ ;
  assign n4371 = ~\new_[4572]_  | ~\new_[4605]_ ;
  assign \new_[4406]_  = \\u1_slt0_reg[11] ;
  assign \new_[4407]_  = \\u1_slt1_reg[11] ;
  assign \new_[4408]_  = \\u1_slt2_reg[11] ;
  assign \new_[4409]_  = \\u1_slt3_reg[11] ;
  assign \new_[4410]_  = \\u1_slt6_reg[11] ;
  assign \new_[4411]_  = ~\\u23_int_set_reg[2] ;
  assign \new_[4412]_  = u15_crac_rd_done_reg;
  assign \new_[4413]_  = ~\new_[13353]_  | ~\new_[4619]_ ;
  assign \new_[4414]_  = ~\new_[13352]_  | ~\new_[4620]_ ;
  assign \new_[4415]_  = ~\new_[13338]_  | ~\new_[4620]_ ;
  assign \new_[4416]_  = ~\new_[13477]_  | ~\new_[4620]_ ;
  assign \new_[4417]_  = ~\new_[13210]_  | ~\new_[4620]_ ;
  assign \new_[4418]_  = ~\new_[13392]_  | ~\new_[4619]_ ;
  assign \new_[4419]_  = ~\new_[13260]_  | ~\new_[4619]_ ;
  assign \new_[4420]_  = ~\new_[13927]_  & (~\new_[8072]_  | ~\new_[8073]_ );
  assign \new_[4421]_  = ~\new_[13927]_  & (~\new_[8074]_  | ~\new_[8075]_ );
  assign \new_[4422]_  = ~\new_[13247]_  | ~\new_[4619]_ ;
  assign \new_[4423]_  = ~\new_[13235]_  | ~\new_[4620]_ ;
  assign \new_[4424]_  = ~\new_[13251]_  | ~\new_[4620]_ ;
  assign \new_[4425]_  = ~\new_[13275]_  | ~\new_[4620]_ ;
  assign \new_[4426]_  = ~\new_[13219]_  | ~\new_[4619]_ ;
  assign \new_[4427]_  = ~\new_[13214]_  | ~\new_[4620]_ ;
  assign \new_[4428]_  = ~\new_[13399]_  | ~\new_[4622]_ ;
  assign \new_[4429]_  = ~\new_[13404]_  | ~\new_[4622]_ ;
  assign \new_[4430]_  = ~\new_[13770]_  | ~\new_[4622]_ ;
  assign \new_[4431]_  = ~\new_[13387]_  | ~\new_[4622]_ ;
  assign \new_[4432]_  = ~\new_[13454]_  | ~\new_[4622]_ ;
  assign \new_[4433]_  = ~\new_[13749]_  | ~\new_[4622]_ ;
  assign \new_[4434]_  = ~\new_[13729]_  | ~\new_[4622]_ ;
  assign \new_[4435]_  = ~\new_[13728]_  | ~\new_[4622]_ ;
  assign \new_[4436]_  = ~\new_[13721]_  | ~\new_[4622]_ ;
  assign \new_[4437]_  = ~\new_[13744]_  | ~\new_[4622]_ ;
  assign \new_[4438]_  = ~\new_[4622]_  & (~\new_[8606]_  | ~\new_[8607]_ );
  assign \new_[4439]_  = ~\new_[4622]_  & (~\new_[8608]_  | ~\new_[8609]_ );
  assign \new_[4440]_  = ~\new_[13383]_  | ~\new_[4622]_ ;
  assign \new_[4441]_  = ~\new_[13451]_  | ~\new_[4622]_ ;
  assign \new_[4442]_  = ~\new_[13496]_  | ~\new_[4622]_ ;
  assign \new_[4443]_  = ~\new_[13643]_  | ~\new_[4622]_ ;
  assign \new_[4444]_  = ~\new_[13444]_  | ~\new_[4622]_ ;
  assign \new_[4445]_  = ~\new_[13447]_  | ~\new_[4622]_ ;
  assign \new_[4446]_  = ~\new_[13335]_  | ~\new_[4619]_ ;
  assign \new_[4447]_  = ~\new_[13486]_  | ~\new_[4619]_ ;
  assign \new_[4448]_  = ~\new_[13743]_  | ~\new_[4619]_ ;
  assign \new_[4449]_  = ~\new_[13876]_  | ~\new_[4709]_  | ~\new_[9781]_ ;
  assign \new_[4450]_  = ~\new_[14097]_ ;
  assign \new_[4451]_  = ~\new_[4515]_ ;
  assign \new_[4452]_  = ~\new_[4523]_ ;
  assign \new_[4453]_  = ~\new_[4523]_ ;
  assign \new_[4454]_  = ~\new_[4526]_ ;
  assign \new_[4455]_  = ~\new_[4527]_ ;
  assign \new_[4456]_  = ~\new_[4528]_ ;
  assign \new_[4457]_  = ~\new_[4621]_  | (~\new_[7718]_  & ~\new_[7770]_ );
  assign \new_[4458]_  = ~\new_[4621]_  | (~\new_[7666]_  & ~\new_[7788]_ );
  assign \new_[4459]_  = ~\new_[13955]_  | (~\new_[7667]_  & ~\new_[7691]_ );
  assign \new_[4460]_  = ~\new_[13955]_  | (~\new_[7668]_  & ~\new_[7771]_ );
  assign \new_[4461]_  = ~\new_[4621]_  | (~\new_[7669]_  & ~\new_[7866]_ );
  assign \new_[4462]_  = ~\new_[4621]_  | (~\new_[7670]_  & ~\new_[7772]_ );
  assign \new_[4463]_  = ~\new_[13955]_  | (~\new_[7721]_  & ~\new_[7867]_ );
  assign \new_[4464]_  = ~\new_[4621]_  | (~\new_[7723]_  & ~\new_[7769]_ );
  assign \new_[4465]_  = ~\new_[4621]_  | (~\new_[7716]_  & ~\new_[7864]_ );
  assign n4446 = ~\new_[13174]_  | ~\new_[4618]_ ;
  assign n4451 = ~\new_[4618]_  | (~\new_[12900]_  & ~\new_[3789]_ );
  assign \new_[4468]_  = ~\new_[13955]_  | (~\new_[7671]_  & ~\new_[14006]_ );
  assign \new_[4469]_  = ~\new_[13955]_  | (~\new_[7717]_  & ~\new_[7924]_ );
  assign \new_[4470]_  = ~\new_[4621]_  | (~\new_[7665]_  & ~\new_[7768]_ );
  assign \new_[4471]_  = ~\new_[4621]_  | (~\new_[7720]_  & ~\new_[7787]_ );
  assign \new_[4472]_  = ~\new_[14161]_ ;
  assign \new_[4473]_  = ~\new_[14162]_ ;
  assign \new_[4474]_  = ~\new_[4475]_ ;
  assign \new_[4475]_  = ~\new_[4623]_ ;
  assign \new_[4476]_  = ~\new_[14061]_ ;
  assign \new_[4477]_  = ~\new_[4478]_ ;
  assign \new_[4478]_  = ~\new_[4624]_ ;
  assign n4391 = \new_[3777]_  ? \new_[4653]_  : \new_[6794]_ ;
  assign n4381 = \new_[3774]_  ? \new_[4653]_  : \new_[5855]_ ;
  assign n4396 = \new_[3778]_  ? \new_[4653]_  : \new_[4816]_ ;
  assign n4376 = \new_[3773]_  ? \new_[4653]_  : \new_[4687]_ ;
  assign n4401 = \new_[3779]_  ? \new_[4653]_  : \new_[4584]_ ;
  assign n4416 = \new_[3782]_  ? \new_[4653]_  : \new_[4386]_ ;
  assign n4406 = \new_[3780]_  ? \new_[4653]_  : \new_[3764]_ ;
  assign n4411 = \new_[3781]_  ? \new_[4653]_  : \new_[3184]_ ;
  assign n4421 = \new_[3783]_  ? \new_[4653]_  : \new_[7687]_ ;
  assign n4426 = \new_[3784]_  ? \new_[4653]_  : \new_[2923]_ ;
  assign n4366 = \new_[3766]_  ? \new_[4653]_  : \new_[2789]_ ;
  assign n4441 = \new_[3787]_  ? \new_[4653]_  : \new_[2748]_ ;
  assign n4331 = \new_[3657]_  ? \new_[4653]_  : \new_[2737]_ ;
  assign n4436 = \new_[3786]_  ? \new_[4653]_  : \new_[2726]_ ;
  assign n4431 = \new_[3785]_  ? \new_[4653]_  : \new_[2717]_ ;
  assign n4386 = \new_[3776]_  ? \new_[4653]_  : \new_[7501]_ ;
  assign \new_[4495]_  = u16_u6_dma_req_r1_reg;
  assign \new_[4496]_  = u16_u7_dma_req_r1_reg;
  assign n4581 = ~\new_[4722]_  | ~\new_[4625]_  | ~\new_[4807]_ ;
  assign n4586 = ~\new_[4723]_  | ~\new_[4626]_  | ~\new_[4808]_ ;
  assign n4571 = ~\new_[4669]_  | ~\new_[4627]_  | ~\new_[4809]_ ;
  assign n4576 = ~\new_[4670]_  | ~\new_[4628]_  | ~\new_[4810]_ ;
  assign n4476 = \new_[4634]_  & \new_[9077]_ ;
  assign n4471 = \new_[4635]_  & \new_[9077]_ ;
  assign \new_[4503]_  = ~\new_[4887]_  | ~\new_[3587]_  | ~\new_[13873]_ ;
  assign \new_[4504]_  = ~\new_[4658]_  | ~\new_[3023]_ ;
  assign \new_[4505]_  = ~\new_[4659]_  | ~\new_[13075]_ ;
  assign \new_[4506]_  = ~\new_[4649]_  | (~\new_[9647]_  & ~\new_[5749]_ );
  assign \new_[4507]_  = ~\new_[4650]_  | (~\new_[8484]_  & ~\new_[5749]_ );
  assign \new_[4508]_  = (~\new_[4677]_  | ~\new_[12964]_ ) & (~\new_[12915]_  | ~\new_[14193]_ );
  assign \new_[4509]_  = (~\new_[4678]_  | ~\new_[13146]_ ) & (~\new_[12971]_  | ~\new_[5878]_ );
  assign n4481 = \new_[4636]_  & \new_[13866]_ ;
  assign \new_[4511]_  = ~\new_[13096]_  | ~\new_[4778]_ ;
  assign \new_[4512]_  = ~\new_[2952]_  | ~\new_[4778]_ ;
  assign \new_[4513]_  = ~\new_[4622]_  | ~\new_[12691]_ ;
  assign \new_[4514]_  = ~\new_[13927]_  | ~\new_[12886]_ ;
  assign \new_[4515]_  = \new_[14161]_  & \new_[14088]_ ;
  assign \new_[4516]_  = ~\new_[13873]_  | ~\new_[4781]_  | ~\new_[9268]_ ;
  assign \new_[4517]_  = ~\new_[4611]_ ;
  assign \new_[4518]_  = ~\new_[4611]_ ;
  assign \new_[4519]_  = ~\new_[4614]_ ;
  assign \new_[4520]_  = ~\new_[4615]_ ;
  assign \new_[4521]_  = ~\new_[4615]_ ;
  assign \new_[4522]_  = \new_[4616]_ ;
  assign \new_[4523]_  = ~\new_[4616]_ ;
  assign \new_[4524]_  = ~\new_[4663]_ ;
  assign \new_[4525]_  = ~\new_[4663]_ ;
  assign \new_[4526]_  = ~\new_[4524]_ ;
  assign \new_[4527]_  = \new_[4665]_  & \new_[13079]_ ;
  assign \new_[4528]_  = \new_[14062]_  & \new_[14131]_ ;
  assign \new_[4529]_  = ~\new_[14106]_  | (~\new_[7724]_  & ~\new_[7967]_ );
  assign \new_[4530]_  = ~\new_[14106]_  | (~\new_[7725]_  & ~\new_[7868]_ );
  assign \new_[4531]_  = ~\new_[14106]_  | (~\new_[7840]_  & ~\new_[7971]_ );
  assign \new_[4532]_  = ~\new_[14106]_  | (~\new_[7726]_  & ~\new_[7968]_ );
  assign \new_[4533]_  = ~\new_[14106]_  | (~\new_[7841]_  & ~\new_[7804]_ );
  assign \new_[4534]_  = ~\new_[14106]_  | (~\new_[7842]_  & ~\new_[7969]_ );
  assign \new_[4535]_  = ~\new_[14106]_  | (~\new_[7843]_  & ~\new_[7794]_ );
  assign \new_[4536]_  = ~\new_[14106]_  | (~\new_[7844]_  & ~\new_[7970]_ );
  assign \new_[4537]_  = ~\new_[14106]_  | (~\new_[7727]_  & ~\new_[7869]_ );
  assign \new_[4538]_  = ~\new_[14106]_  | (~\new_[7728]_  & ~\new_[7870]_ );
  assign \new_[4539]_  = ~\new_[3607]_  & (~\new_[3606]_  | ~\new_[4679]_ );
  assign \new_[4540]_  = ~\new_[14106]_  | (~\new_[7845]_  & ~\new_[7871]_ );
  assign \new_[4541]_  = ~\new_[14106]_  | (~\new_[7729]_  & ~\new_[7923]_ );
  assign \new_[4542]_  = ~\new_[14106]_  | (~\new_[7730]_  & ~\new_[7872]_ );
  assign \new_[4543]_  = ~\new_[14106]_  | (~\new_[7731]_  & ~\new_[7853]_ );
  assign n4566 = ~\new_[12942]_  | (~\new_[4680]_  & ~\new_[3789]_ );
  assign \new_[4545]_  = ~\new_[3788]_  | ~\new_[4638]_ ;
  assign \new_[4546]_  = ~\new_[3606]_  | ~\new_[4637]_ ;
  assign n4506 = \new_[4075]_  ? \new_[4695]_  : \new_[7686]_ ;
  assign n4496 = \new_[4073]_  ? \new_[4695]_  : \new_[2922]_ ;
  assign n4511 = \new_[4076]_  ? \new_[4695]_  : \new_[2785]_ ;
  assign n4516 = \new_[4077]_  ? \new_[4695]_  : \new_[2747]_ ;
  assign n4521 = \new_[4078]_  ? \new_[4695]_  : \new_[2736]_ ;
  assign n4501 = \new_[4074]_  ? \new_[4695]_  : \new_[2725]_ ;
  assign n4526 = \new_[4079]_  ? \new_[4695]_  : \new_[2716]_ ;
  assign n4531 = \new_[4080]_  ? \new_[4695]_  : \new_[7502]_ ;
  assign n4536 = \new_[4081]_  ? \new_[4695]_  : \new_[6791]_ ;
  assign n4491 = \new_[4072]_  ? \new_[4695]_  : \new_[5856]_ ;
  assign n4551 = \new_[4084]_  ? \new_[4695]_  : \new_[4817]_ ;
  assign n4541 = \new_[4082]_  ? \new_[4695]_  : \new_[4688]_ ;
  assign n4546 = \new_[4083]_  ? \new_[4695]_  : \new_[4585]_ ;
  assign n4561 = \new_[4086]_  ? \new_[4695]_  : \new_[4409]_ ;
  assign n4556 = \new_[4085]_  ? \new_[4695]_  : \new_[3763]_ ;
  assign n4486 = \new_[4071]_  ? \new_[4695]_  : \new_[3186]_ ;
  assign n4466 = \\u1_sr_reg[13] ;
  assign \new_[4564]_  = ~\new_[4675]_  & (~\new_[12730]_  | ~\new_[4784]_ );
  assign \new_[4565]_  = ~\new_[4676]_  & (~\new_[13048]_  | ~\new_[4785]_ );
  assign n4601 = \new_[4406]_  ? \new_[9006]_  : n4721;
  assign n4606 = n4721 ? \new_[8805]_  : \new_[4407]_ ;
  assign n4611 = n4721 ? \new_[8996]_  : \new_[4408]_ ;
  assign n4616 = n4721 ? \new_[9002]_  : \new_[4409]_ ;
  assign n4596 = n4721 ? \new_[9000]_  : \new_[4386]_ ;
  assign n4621 = n4721 ? \new_[9001]_  : \new_[4410]_ ;
  assign \new_[4572]_  = ~\new_[5749]_  | ~\new_[13866]_  | ~\new_[3771]_ ;
  assign n4626 = ~\new_[4632]_ ;
  assign \new_[4574]_  = \new_[3760]_  | \new_[4674]_ ;
  assign \new_[4575]_  = (~\new_[4747]_  | ~\new_[12898]_ ) & (~\new_[12981]_  | ~\new_[14194]_ );
  assign \new_[4576]_  = \\u1_slt6_reg[10] ;
  assign \new_[4577]_  = (~\new_[4748]_  | ~\new_[12725]_ ) & (~\new_[12901]_  | ~\new_[6444]_ );
  assign \new_[4578]_  = \\u1_slt2_reg[10] ;
  assign \new_[4579]_  = (~\new_[4749]_  | ~\new_[12983]_ ) & (~\new_[12966]_  | ~\new_[6445]_ );
  assign \new_[4580]_  = (~\new_[4750]_  | ~\new_[12921]_ ) & (~\new_[13032]_  | ~\new_[6446]_ );
  assign \new_[4581]_  = u14_u4_en_out_l_reg;
  assign \new_[4582]_  = u2_sync_resume_reg;
  assign \new_[4583]_  = \\u1_slt1_reg[10] ;
  assign \new_[4584]_  = \\u1_slt4_reg[10] ;
  assign \new_[4585]_  = \\u1_slt3_reg[10] ;
  assign \new_[4586]_  = u14_u0_en_out_l_reg;
  assign \new_[4587]_  = u14_u1_en_out_l_reg;
  assign \new_[4588]_  = u14_u2_en_out_l_reg;
  assign \new_[4589]_  = u14_u3_en_out_l_reg;
  assign \new_[4590]_  = u14_u5_en_out_l_reg;
  assign \new_[4591]_  = u14_crac_valid_r_reg;
  assign \new_[4592]_  = ~\new_[3307]_  | ~\new_[4887]_ ;
  assign \new_[4593]_  = ~\new_[3150]_  | ~\new_[4887]_ ;
  assign \new_[4594]_  = ~\new_[4651]_ ;
  assign \new_[4595]_  = ~\new_[4654]_ ;
  assign \new_[4596]_  = ~\new_[4657]_ ;
  assign \new_[4597]_  = ~\new_[4657]_ ;
  assign \new_[4598]_  = ~\new_[4656]_ ;
  assign \new_[4599]_  = ~\new_[4656]_ ;
  assign \new_[4600]_  = ~\new_[4656]_ ;
  assign \new_[4601]_  = ~\new_[4656]_ ;
  assign \new_[4602]_  = ~\new_[4657]_ ;
  assign \new_[4603]_  = ~\new_[4657]_ ;
  assign \new_[4604]_  = ~\new_[4657]_ ;
  assign \new_[4605]_  = ~\new_[13866]_  | ~\new_[4886]_  | ~\new_[9780]_ ;
  assign \new_[4606]_  = ~\new_[4713]_  & ~\new_[13953]_ ;
  assign \new_[4607]_  = ~\new_[14104]_  & ~\new_[4715]_ ;
  assign \new_[4608]_  = ~\new_[4660]_ ;
  assign \new_[4609]_  = ~\new_[4660]_ ;
  assign \new_[4610]_  = \new_[4661]_ ;
  assign \new_[4611]_  = ~\new_[4661]_ ;
  assign \new_[4612]_  = ~\new_[4707]_ ;
  assign \new_[4613]_  = ~\new_[4707]_ ;
  assign \new_[4614]_  = ~\new_[4612]_ ;
  assign \new_[4615]_  = ~\new_[4662]_ ;
  assign \new_[4616]_  = ~\new_[4663]_ ;
  assign n4631 = ~\new_[4680]_  & ~\new_[13395]_ ;
  assign \new_[4618]_  = ~\new_[4679]_  | ~\new_[3119]_ ;
  assign \new_[4619]_  = ~\new_[13955]_ ;
  assign \new_[4620]_  = ~\new_[13955]_ ;
  assign \new_[4621]_  = ~\new_[13927]_ ;
  assign \new_[4622]_  = ~\new_[14107]_ ;
  assign \new_[4623]_  = ~\new_[4665]_ ;
  assign \new_[4624]_  = ~\new_[4666]_ ;
  assign \new_[4625]_  = ~\new_[4743]_  & (~\new_[12765]_  | ~\new_[4928]_ );
  assign \new_[4626]_  = ~\new_[4744]_  & (~\new_[12632]_  | ~\new_[4930]_ );
  assign \new_[4627]_  = ~\new_[4745]_  & (~\new_[12772]_  | ~\new_[4931]_ );
  assign \new_[4628]_  = ~\new_[4746]_  & (~\new_[12865]_  | ~\new_[4932]_ );
  assign \new_[4629]_  = \\u0_slt9_r_reg[2] ;
  assign n4646 = \\u1_sr_reg[12] ;
  assign \new_[4631]_  = \\u26_ps_cnt_reg[5] ;
  assign \new_[4632]_  = ~\new_[13306]_  & (~\new_[8803]_  | ~\new_[4886]_ );
  assign \new_[4633]_  = \\u26_ps_cnt_reg[2] ;
  assign \new_[4634]_  = \new_[4069]_  | \new_[4733]_ ;
  assign \new_[4635]_  = \new_[4068]_  | \new_[4734]_ ;
  assign \new_[4636]_  = \new_[13141]_  ? \new_[4886]_  : \new_[10313]_ ;
  assign \new_[4637]_  = ~\new_[4679]_ ;
  assign \new_[4638]_  = ~\new_[4680]_ ;
  assign \new_[4639]_  = \\u26_ps_cnt_reg[0] ;
  assign \new_[4640]_  = \\u26_ps_cnt_reg[1] ;
  assign \new_[4641]_  = \\u26_ps_cnt_reg[4] ;
  assign \new_[4642]_  = \\u26_ps_cnt_reg[3] ;
  assign \wb_data_o[1]  = \\u12_wb_data_o_reg[1] ;
  assign \new_[4644]_  = ~\\u17_int_set_reg[2] ;
  assign \new_[4645]_  = ~\\u18_int_set_reg[2] ;
  assign \new_[4646]_  = ~\\u21_int_set_reg[2] ;
  assign \new_[4647]_  = ~\\u20_int_set_reg[2] ;
  assign \new_[4648]_  = u14_crac_wr_r_reg;
  assign \new_[4649]_  = ~\new_[3540]_  | ~\new_[5749]_ ;
  assign \new_[4650]_  = ~\new_[5749]_  | ~\new_[3374]_ ;
  assign \new_[4651]_  = \new_[3340]_  | \new_[4778]_ ;
  assign \new_[4652]_  = ~\\u22_int_set_reg[2] ;
  assign \new_[4653]_  = ~\new_[4696]_ ;
  assign \new_[4654]_  = ~\new_[4703]_ ;
  assign \new_[4655]_  = ~\new_[4705]_ ;
  assign \new_[4656]_  = ~\new_[4704]_ ;
  assign \new_[4657]_  = ~\new_[4704]_ ;
  assign \new_[4658]_  = ~\new_[13956]_  | ~\new_[13953]_ ;
  assign \new_[4659]_  = ~\new_[14108]_  | ~\new_[14104]_ ;
  assign \new_[4660]_  = ~\new_[4706]_ ;
  assign \new_[4661]_  = ~\new_[4707]_ ;
  assign \new_[4662]_  = \new_[4708]_ ;
  assign \new_[4663]_  = ~\new_[4708]_ ;
  assign \new_[4664]_  = ~\\u19_int_set_reg[2] ;
  assign \new_[4665]_  = ~\new_[4716]_ ;
  assign \new_[4666]_  = ~\new_[4717]_ ;
  assign \new_[4667]_  = ~\new_[12964]_  | (~\new_[8626]_  & ~\new_[4784]_ );
  assign \new_[4668]_  = ~\new_[13146]_  | (~\new_[8628]_  & ~\new_[4785]_ );
  assign \new_[4669]_  = ~\new_[12983]_  | (~\new_[8629]_  & ~\new_[4931]_ );
  assign \new_[4670]_  = ~\new_[12921]_  | (~\new_[9081]_  & ~\new_[4932]_ );
  assign \new_[4671]_  = ~\new_[4806]_  & (~\new_[7519]_  | ~\new_[12766]_ );
  assign \new_[4672]_  = \\u1_slt2_reg[9] ;
  assign \new_[4673]_  = u14_u3_full_empty_r_reg;
  assign \new_[4674]_  = \\u25_int_set_reg[0] ;
  assign \new_[4675]_  = ~\new_[4792]_  & ~\new_[12744]_ ;
  assign \new_[4676]_  = ~\new_[4793]_  & ~\new_[13052]_ ;
  assign \new_[4677]_  = ~\new_[4787]_  | (~\new_[12604]_  & ~\new_[10320]_ );
  assign \new_[4678]_  = ~\new_[4789]_  | (~\new_[12648]_  & ~\new_[10318]_ );
  assign \new_[4679]_  = \new_[4812]_  & \new_[13885]_ ;
  assign \new_[4680]_  = \new_[4812]_  | \new_[13885]_ ;
  assign \new_[4681]_  = u14_u0_full_empty_r_reg;
  assign \new_[4682]_  = u14_u1_full_empty_r_reg;
  assign \new_[4683]_  = u14_u2_full_empty_r_reg;
  assign \new_[4684]_  = u14_u5_full_empty_r_reg;
  assign \new_[4685]_  = \\u1_slt0_reg[9] ;
  assign \new_[4686]_  = u14_u4_full_empty_r_reg;
  assign \new_[4687]_  = \\u1_slt4_reg[9] ;
  assign \new_[4688]_  = \\u1_slt3_reg[9] ;
  assign \new_[4689]_  = \\u8_wp_reg[0] ;
  assign \new_[4690]_  = \\u3_wp_reg[0] ;
  assign \new_[4691]_  = \\u4_wp_reg[0] ;
  assign \new_[4692]_  = \\u5_wp_reg[0] ;
  assign \new_[4693]_  = \\u6_wp_reg[0] ;
  assign \new_[4694]_  = \\u7_wp_reg[0] ;
  assign \new_[4695]_  = ~\new_[4775]_ ;
  assign \new_[4696]_  = \new_[3587]_  | \new_[4887]_ ;
  assign n4686 = \new_[4888]_  | n5641;
  assign n4691 = \new_[4889]_  | n5646;
  assign n4696 = \new_[4890]_  | n5651;
  assign n4701 = \new_[4891]_  | n5656;
  assign n4661 = \new_[4892]_  | n5661;
  assign n4706 = \new_[4893]_  | n5666;
  assign \new_[4703]_  = ~\new_[4776]_ ;
  assign \new_[4704]_  = ~\new_[4776]_ ;
  assign \new_[4705]_  = \new_[4776]_ ;
  assign \new_[4706]_  = \new_[4777]_ ;
  assign \new_[4707]_  = ~\new_[4777]_ ;
  assign \new_[4708]_  = ~\new_[12408]_  | ~\new_[4885]_ ;
  assign \new_[4709]_  = ~\new_[4778]_ ;
  assign n4671 = n4891 ? \new_[8805]_  : \new_[4583]_ ;
  assign n4711 = ~\new_[5020]_  | ~\new_[5021]_  | ~\new_[5019]_ ;
  assign n4656 = n4891 ? \new_[8996]_  : \new_[4578]_ ;
  assign \new_[4713]_  = ~\new_[13956]_ ;
  assign n4681 = n4891 ? \new_[9002]_  : \new_[4585]_ ;
  assign \new_[4715]_  = ~\new_[14108]_ ;
  assign \new_[4716]_  = ~\new_[4779]_ ;
  assign \new_[4717]_  = ~\new_[4780]_ ;
  assign n4676 = n4891 ? \new_[9000]_  : \new_[4584]_ ;
  assign n4651 = n4891 ? \new_[9001]_  : \new_[4576]_ ;
  assign \new_[4720]_  = \\u1_slt6_reg[9] ;
  assign n4666 = ~\new_[4811]_  & (~\new_[13171]_  | ~\new_[13170]_ );
  assign \new_[4722]_  = ~\new_[12898]_  | (~\new_[8622]_  & ~\new_[4928]_ );
  assign \new_[4723]_  = ~\new_[12725]_  | (~\new_[9080]_  & ~\new_[4930]_ );
  assign \new_[4724]_  = ~\new_[4988]_  & (~\new_[7603]_  | ~\new_[12734]_ );
  assign \new_[4725]_  = ~\new_[4989]_  & (~\new_[7604]_  | ~\new_[12754]_ );
  assign ac97_reset_pad_o_ = u26_ac97_rst__reg;
  assign n4721 = \\u1_sr_reg[11] ;
  assign \new_[4728]_  = \\u26_cnt_reg[2] ;
  assign n4756 = ~\new_[8168]_  | ~\new_[5713]_ ;
  assign \new_[4730]_  = ~\new_[4787]_ ;
  assign \new_[4731]_  = ~\new_[4789]_ ;
  assign n4716 = \new_[13369]_  ? \new_[7937]_  : \new_[5886]_ ;
  assign \new_[4733]_  = \\u23_int_set_reg[0] ;
  assign \new_[4734]_  = \\u24_int_set_reg[0] ;
  assign \new_[4735]_  = ~\new_[5879]_  | ~\new_[5078]_  | ~\new_[5077]_ ;
  assign \new_[4736]_  = ~\new_[5880]_  | ~\new_[5091]_  | ~\new_[5090]_ ;
  assign n4736 = ~\new_[4934]_  & ~\new_[4639]_ ;
  assign n4741 = ~\new_[12346]_  & ~\new_[4934]_ ;
  assign n4731 = ~\new_[10509]_  & ~\new_[4934]_ ;
  assign n4751 = ~\new_[11429]_  & ~\new_[4934]_ ;
  assign n4746 = ~\new_[10395]_  & ~\new_[4934]_ ;
  assign n4726 = ~\new_[9668]_  & ~\new_[4934]_ ;
  assign \new_[4743]_  = ~\new_[4956]_  & ~\new_[12750]_ ;
  assign \new_[4744]_  = ~\new_[4957]_  & ~\new_[12770]_ ;
  assign \new_[4745]_  = ~\new_[4959]_  & ~\new_[12752]_ ;
  assign \new_[4746]_  = ~\new_[4960]_  & ~\new_[12737]_ ;
  assign \new_[4747]_  = ~\new_[4946]_  | (~\new_[12607]_  & ~\new_[10319]_ );
  assign \new_[4748]_  = ~\new_[4947]_  | (~\new_[12529]_  & ~\new_[12085]_ );
  assign \new_[4749]_  = ~\new_[4949]_  | (~\new_[12917]_  & ~\new_[10321]_ );
  assign \new_[4750]_  = ~\new_[4950]_  | (~\new_[12979]_  & ~\new_[12086]_ );
  assign n4781 = ~\new_[5022]_  | ~\new_[5021]_ ;
  assign \new_[4752]_  = u14_u8_en_out_l_reg;
  assign \new_[4753]_  = \\u5_wp_reg[1] ;
  assign \new_[4754]_  = \\u6_wp_reg[2] ;
  assign \new_[4755]_  = \\u26_cnt_reg[0] ;
  assign \new_[4756]_  = \\u26_cnt_reg[1] ;
  assign \new_[4757]_  = \\u8_wp_reg[2] ;
  assign \new_[4758]_  = \\u3_wp_reg[2] ;
  assign \new_[4759]_  = \\u5_wp_reg[2] ;
  assign \new_[4760]_  = \\u7_wp_reg[2] ;
  assign \new_[4761]_  = u14_u6_en_out_l_reg;
  assign \new_[4762]_  = u14_u7_en_out_l_reg;
  assign \new_[4763]_  = \\u8_wp_reg[1] ;
  assign \new_[4764]_  = \\u3_wp_reg[1] ;
  assign \new_[4765]_  = \\u4_wp_reg[1] ;
  assign \new_[4766]_  = \\u6_wp_reg[1] ;
  assign \new_[4767]_  = \\u7_wp_reg[1] ;
  assign \new_[4768]_  = \\u4_wp_reg[2] ;
  assign n4761 = ~\new_[5739]_  | ~\new_[4644]_ ;
  assign n4766 = ~\new_[5741]_  | ~\new_[4645]_ ;
  assign n4791 = ~\new_[5742]_  | ~\new_[4664]_ ;
  assign n4776 = ~\new_[5745]_  | ~\new_[4647]_ ;
  assign n4771 = ~\new_[5746]_  | ~\new_[4646]_ ;
  assign n4786 = ~\new_[5747]_  | ~\new_[4652]_ ;
  assign \new_[4775]_  = \new_[3771]_  | \new_[5749]_ ;
  assign \new_[4776]_  = ~\new_[4879]_ ;
  assign \new_[4777]_  = ~\new_[12407]_  | ~\new_[5750]_ ;
  assign \new_[4778]_  = ~\new_[4885]_ ;
  assign \new_[4779]_  = ~\new_[4983]_  & ~\new_[6787]_ ;
  assign \new_[4780]_  = ~\new_[4985]_  & ~\new_[6789]_ ;
  assign \new_[4781]_  = ~\new_[4887]_ ;
  assign \new_[4782]_  = ~\new_[14193]_  & (~\new_[7694]_  | ~\new_[12815]_ );
  assign \new_[4783]_  = ~\new_[5878]_  & (~\new_[7801]_  | ~\new_[12783]_ );
  assign \new_[4784]_  = \new_[5879]_  | \new_[7692]_ ;
  assign \new_[4785]_  = \new_[5880]_  | \new_[7797]_ ;
  assign \new_[4786]_  = ~\new_[4946]_ ;
  assign \new_[4787]_  = ~\new_[5877]_  & (~\new_[12815]_  | ~\new_[7805]_ );
  assign \new_[4788]_  = ~\new_[4947]_ ;
  assign \new_[4789]_  = ~\new_[5878]_  & (~\new_[12783]_  | ~\new_[7941]_ );
  assign \new_[4790]_  = ~\new_[4949]_ ;
  assign \new_[4791]_  = ~\new_[4950]_ ;
  assign \new_[4792]_  = ~\new_[5879]_  & (~\new_[9675]_  | ~\new_[7692]_ );
  assign \new_[4793]_  = ~\new_[5880]_  & (~\new_[9672]_  | ~\new_[7797]_ );
  assign n4806 = ~\new_[6810]_  | ~\new_[5769]_  | ~\new_[12035]_ ;
  assign n4811 = \new_[4681]_  ? \new_[13885]_  : \new_[6829]_ ;
  assign n4816 = \new_[4682]_  ? \new_[13885]_  : \new_[6560]_ ;
  assign n4821 = \new_[4683]_  ? \new_[13885]_  : \new_[6831]_ ;
  assign n4801 = \new_[4673]_  ? \new_[13885]_  : \new_[6561]_ ;
  assign n4836 = \new_[4686]_  ? \new_[13885]_  : \new_[6833]_ ;
  assign n4826 = \new_[4684]_  ? \new_[13885]_  : \new_[6834]_ ;
  assign n4831 = \new_[4685]_  ? \new_[9006]_  : n9106;
  assign n4796 = n9106 ? \new_[8996]_  : \new_[4672]_ ;
  assign n4846 = n9106 ? \new_[9002]_  : \new_[4688]_ ;
  assign n4841 = n9106 ? \new_[9000]_  : \new_[4687]_ ;
  assign n4881 = n9106 ? \new_[9001]_  : \new_[4720]_ ;
  assign \new_[4806]_  = ~\new_[5768]_  | (~\new_[7597]_  & ~\new_[12872]_ );
  assign \new_[4807]_  = ~\new_[6447]_  | ~\new_[5095]_  | ~\new_[5042]_ ;
  assign \new_[4808]_  = ~\new_[6448]_  | ~\new_[5085]_  | ~\new_[5084]_ ;
  assign \new_[4809]_  = ~\new_[6449]_  | ~\new_[5850]_  | ~\new_[5876]_ ;
  assign \new_[4810]_  = ~\new_[6450]_  | ~\new_[5845]_  | ~\new_[5844]_ ;
  assign \new_[4811]_  = ~\new_[4582]_  & (~\new_[6442]_  | ~suspended_o);
  assign \new_[4812]_  = u15_valid_r_reg;
  assign \new_[4813]_  = \\u1_slt6_reg[8] ;
  assign \new_[4814]_  = \\u1_slt2_reg[8] ;
  assign \new_[4815]_  = \\u1_slt1_reg[8] ;
  assign \new_[4816]_  = \\u1_slt4_reg[8] ;
  assign \new_[4817]_  = \\u1_slt3_reg[8] ;
  assign \new_[4818]_  = \\u4_mem_reg[0][13] ;
  assign \new_[4819]_  = \\u4_mem_reg[0][14] ;
  assign \new_[4820]_  = \\u4_mem_reg[0][16] ;
  assign \new_[4821]_  = \\u4_mem_reg[0][19] ;
  assign \new_[4822]_  = \\u4_mem_reg[0][22] ;
  assign \new_[4823]_  = \\u4_mem_reg[0][24] ;
  assign \new_[4824]_  = \\u4_mem_reg[0][31] ;
  assign \new_[4825]_  = \\u4_mem_reg[0][4] ;
  assign \new_[4826]_  = \\u4_mem_reg[0][7] ;
  assign \new_[4827]_  = \\u4_mem_reg[0][9] ;
  assign \new_[4828]_  = \\u5_mem_reg[0][13] ;
  assign \new_[4829]_  = \\u5_mem_reg[0][14] ;
  assign \new_[4830]_  = \\u5_mem_reg[0][16] ;
  assign \new_[4831]_  = \\u5_mem_reg[0][19] ;
  assign \new_[4832]_  = \\u5_mem_reg[0][22] ;
  assign \new_[4833]_  = \\u5_mem_reg[0][24] ;
  assign \new_[4834]_  = \\u5_mem_reg[0][31] ;
  assign \new_[4835]_  = \\u5_mem_reg[0][4] ;
  assign \new_[4836]_  = \\u5_mem_reg[0][7] ;
  assign \new_[4837]_  = \\u5_mem_reg[0][9] ;
  assign \new_[4838]_  = \\u6_mem_reg[0][13] ;
  assign \new_[4839]_  = \\u6_mem_reg[0][14] ;
  assign \new_[4840]_  = \\u6_mem_reg[0][16] ;
  assign \new_[4841]_  = \\u6_mem_reg[0][19] ;
  assign \new_[4842]_  = \\u6_mem_reg[0][22] ;
  assign \new_[4843]_  = \\u6_mem_reg[0][24] ;
  assign \new_[4844]_  = \\u6_mem_reg[0][31] ;
  assign \new_[4845]_  = \\u6_mem_reg[0][4] ;
  assign \new_[4846]_  = \\u6_mem_reg[0][7] ;
  assign \new_[4847]_  = \\u6_mem_reg[0][9] ;
  assign \new_[4848]_  = \\u7_mem_reg[0][13] ;
  assign \new_[4849]_  = \\u7_mem_reg[0][14] ;
  assign \new_[4850]_  = \\u7_mem_reg[0][16] ;
  assign \new_[4851]_  = \\u7_mem_reg[0][19] ;
  assign \new_[4852]_  = \\u7_mem_reg[0][22] ;
  assign \new_[4853]_  = \\u7_mem_reg[0][24] ;
  assign \new_[4854]_  = \\u7_mem_reg[0][31] ;
  assign \new_[4855]_  = \\u7_mem_reg[0][4] ;
  assign \new_[4856]_  = \\u7_mem_reg[0][7] ;
  assign \new_[4857]_  = \\u7_mem_reg[0][9] ;
  assign \new_[4858]_  = \\u3_mem_reg[0][11] ;
  assign \new_[4859]_  = \\u3_mem_reg[0][12] ;
  assign \new_[4860]_  = \\u3_mem_reg[0][15] ;
  assign \new_[4861]_  = \\u8_mem_reg[0][0] ;
  assign \new_[4862]_  = \\u8_mem_reg[0][11] ;
  assign \new_[4863]_  = \\u8_mem_reg[0][12] ;
  assign \new_[4864]_  = \\u8_mem_reg[0][17] ;
  assign \new_[4865]_  = \\u3_mem_reg[0][1] ;
  assign \new_[4866]_  = \\u3_mem_reg[0][21] ;
  assign \new_[4867]_  = \\u8_mem_reg[0][26] ;
  assign \new_[4868]_  = \\u8_mem_reg[0][28] ;
  assign \new_[4869]_  = \\u8_mem_reg[0][29] ;
  assign \new_[4870]_  = \\u8_mem_reg[0][30] ;
  assign \new_[4871]_  = \\u3_mem_reg[0][27] ;
  assign \new_[4872]_  = \\u8_mem_reg[0][4] ;
  assign \new_[4873]_  = \\u8_mem_reg[0][5] ;
  assign \new_[4874]_  = \\u3_mem_reg[0][2] ;
  assign \new_[4875]_  = \\u3_mem_reg[0][29] ;
  assign \new_[4876]_  = \\u3_mem_reg[0][6] ;
  assign \new_[4877]_  = \\u3_mem_reg[0][5] ;
  assign n4851 = ~\new_[5831]_  & ~\new_[12402]_ ;
  assign \new_[4879]_  = ~\new_[12266]_  | ~\new_[5887]_ ;
  assign n4856 = ~\new_[5834]_  & ~\new_[12811]_ ;
  assign n4861 = ~\new_[5832]_  & ~\new_[12040]_ ;
  assign n4866 = ~\new_[5833]_  & ~\new_[11421]_ ;
  assign n4871 = ~\new_[5835]_  & ~\new_[12074]_ ;
  assign n4876 = ~\new_[5836]_  & ~\new_[12409]_ ;
  assign \new_[4885]_  = ~\new_[7420]_  & ~\new_[5837]_ ;
  assign \new_[4886]_  = ~\new_[5749]_ ;
  assign \new_[4887]_  = ~\new_[5750]_ ;
  assign \new_[4888]_  = ~\new_[12684]_  & (~\new_[6429]_  | ~\new_[12392]_ );
  assign \new_[4889]_  = ~\new_[12699]_  & (~\new_[6431]_  | ~\new_[12438]_ );
  assign \new_[4890]_  = ~\new_[12700]_  & (~\new_[6433]_  | ~\new_[12394]_ );
  assign \new_[4891]_  = ~\new_[12682]_  & (~\new_[6435]_  | ~\new_[12400]_ );
  assign \new_[4892]_  = ~\new_[12701]_  & (~\new_[6437]_  | ~\new_[12622]_ );
  assign \new_[4893]_  = ~\new_[12702]_  & (~\new_[6439]_  | ~\new_[12592]_ );
  assign \new_[4894]_  = \\u13_crac_r_reg[6] ;
  assign \new_[4895]_  = \\u3_mem_reg[0][17] ;
  assign \new_[4896]_  = \\u8_mem_reg[2][18] ;
  assign \new_[4897]_  = \\u7_mem_reg[0][20] ;
  assign \new_[4898]_  = \\u8_mem_reg[2][25] ;
  assign \new_[4899]_  = \\u8_mem_reg[2][28] ;
  assign \new_[4900]_  = \\u4_mem_reg[2][16] ;
  assign \new_[4901]_  = \\u5_mem_reg[1][26] ;
  assign \new_[4902]_  = \\u13_occ0_r_reg[11] ;
  assign \new_[4903]_  = \\u5_mem_reg[1][22] ;
  assign \new_[4904]_  = \\u5_mem_reg[1][15] ;
  assign \new_[4905]_  = \\u5_mem_reg[1][19] ;
  assign \new_[4906]_  = \\u5_mem_reg[1][11] ;
  assign \new_[4907]_  = \\u3_mem_reg[1][22] ;
  assign \new_[4908]_  = \\u8_mem_reg[2][20] ;
  assign \new_[4909]_  = \\u4_mem_reg[3][9] ;
  assign \new_[4910]_  = \\u4_mem_reg[3][5] ;
  assign \new_[4911]_  = \\u4_mem_reg[3][30] ;
  assign \new_[4912]_  = \\u8_mem_reg[0][15] ;
  assign \new_[4913]_  = \\u3_mem_reg[0][16] ;
  assign \new_[4914]_  = \\u4_mem_reg[3][23] ;
  assign \new_[4915]_  = \\u4_mem_reg[3][27] ;
  assign \new_[4916]_  = \\u8_mem_reg[1][6] ;
  assign \new_[4917]_  = \\u13_occ0_r_reg[8] ;
  assign \new_[4918]_  = \\u13_icc_r_reg[8] ;
  assign \new_[4919]_  = \\u8_mem_reg[2][13] ;
  assign \new_[4920]_  = \\u3_mem_reg[1][19] ;
  assign \new_[4921]_  = \\u4_mem_reg[2][9] ;
  assign \new_[4922]_  = \\u4_mem_reg[3][16] ;
  assign \new_[4923]_  = \\u4_mem_reg[3][12] ;
  assign \new_[4924]_  = ~\new_[14194]_  & (~\new_[7800]_  | ~\new_[12724]_ );
  assign \new_[4925]_  = ~\new_[6444]_  & (~\new_[7695]_  | ~\new_[12782]_ );
  assign \new_[4926]_  = ~\new_[6445]_  & (~\new_[7802]_  | ~\new_[12820]_ );
  assign \new_[4927]_  = ~\new_[6446]_  & (~\new_[7803]_  | ~\new_[12723]_ );
  assign \new_[4928]_  = \new_[6447]_  | \new_[7796]_ ;
  assign \new_[4929]_  = \\u4_mem_reg[2][5] ;
  assign \new_[4930]_  = \new_[6448]_  | \new_[7693]_ ;
  assign \new_[4931]_  = \new_[6449]_  | \new_[7798]_ ;
  assign \new_[4932]_  = \new_[6450]_  | \new_[7799]_ ;
  assign n4926 = \new_[8801]_  & \new_[6441]_ ;
  assign \new_[4934]_  = ~\new_[12077]_  | ~\new_[6441]_ ;
  assign \new_[4935]_  = \\u3_mem_reg[1][15] ;
  assign \new_[4936]_  = \\u4_mem_reg[2][30] ;
  assign \new_[4937]_  = \\u4_mem_reg[2][27] ;
  assign \new_[4938]_  = \\u4_mem_reg[2][23] ;
  assign n4931 = \new_[8795]_  & \new_[6441]_ ;
  assign n4896 = \new_[8796]_  & \new_[6441]_ ;
  assign \new_[4941]_  = \\u7_mem_reg[0][30] ;
  assign \new_[4942]_  = \\u3_mem_reg[2][2] ;
  assign \new_[4943]_  = \\u8_mem_reg[1][21] ;
  assign n4886 = \new_[12118]_  & \new_[6441]_ ;
  assign \new_[4945]_  = \\u3_mem_reg[1][11] ;
  assign \new_[4946]_  = ~\new_[6443]_  & (~\new_[12724]_  | ~\new_[7938]_ );
  assign \new_[4947]_  = ~\new_[6444]_  & (~\new_[12782]_  | ~\new_[7806]_ );
  assign \new_[4948]_  = \\u8_mem_reg[1][3] ;
  assign \new_[4949]_  = ~\new_[6445]_  & (~\new_[12820]_  | ~\new_[7942]_ );
  assign \new_[4950]_  = ~\new_[6446]_  & (~\new_[12723]_  | ~\new_[7943]_ );
  assign \new_[4951]_  = \\u4_mem_reg[2][12] ;
  assign \new_[4952]_  = \\u4_mem_reg[1][30] ;
  assign \new_[4953]_  = \\u4_mem_reg[1][9] ;
  assign \new_[4954]_  = \\u4_mem_reg[1][5] ;
  assign n4901 = ~\new_[7427]_  | ~\new_[6289]_  | ~\new_[12033]_ ;
  assign \new_[4956]_  = ~\new_[6447]_  & (~\new_[9674]_  | ~\new_[7796]_ );
  assign \new_[4957]_  = ~\new_[6448]_  & (~\new_[11443]_  | ~\new_[7693]_ );
  assign n4906 = ~\new_[7428]_  | ~\new_[6292]_  | ~\new_[12034]_ ;
  assign \new_[4959]_  = ~\new_[6449]_  & (~\new_[9676]_  | ~\new_[7798]_ );
  assign \new_[4960]_  = ~\new_[6450]_  & (~\new_[11428]_  | ~\new_[7799]_ );
  assign \new_[4961]_  = \\u4_mem_reg[1][27] ;
  assign \new_[4962]_  = \\u8_mem_reg[1][28] ;
  assign \new_[4963]_  = \\u3_mem_reg[0][13] ;
  assign \new_[4964]_  = \\u8_mem_reg[1][25] ;
  assign \new_[4965]_  = \\u4_mem_reg[1][23] ;
  assign \new_[4966]_  = \\u4_mem_reg[1][16] ;
  assign \new_[4967]_  = \\u7_mem_reg[0][6] ;
  assign \new_[4968]_  = \\u7_mem_reg[1][25] ;
  assign \new_[4969]_  = \\u3_mem_reg[3][3] ;
  assign \new_[4970]_  = \\u4_mem_reg[1][12] ;
  assign \new_[4971]_  = \\u7_mem_reg[3][3] ;
  assign \new_[4972]_  = \\u8_mem_reg[1][14] ;
  assign \new_[4973]_  = \\u8_mem_reg[1][18] ;
  assign \new_[4974]_  = \\u3_mem_reg[3][6] ;
  assign \new_[4975]_  = \\u3_mem_reg[3][22] ;
  assign \new_[4976]_  = \\u3_mem_reg[3][30] ;
  assign \new_[4977]_  = \\u3_mem_reg[3][27] ;
  assign \new_[4978]_  = \\u7_mem_reg[0][23] ;
  assign \new_[4979]_  = \\u3_mem_reg[3][19] ;
  assign \new_[4980]_  = u14_u0_en_out_l2_reg;
  assign \new_[4981]_  = u14_u1_en_out_l2_reg;
  assign \new_[4982]_  = u14_u2_en_out_l2_reg;
  assign \new_[4983]_  = u14_u3_en_out_l2_reg;
  assign \new_[4984]_  = u14_u4_en_out_l2_reg;
  assign \new_[4985]_  = u14_u5_en_out_l2_reg;
  assign \new_[4986]_  = \\u6_mem_reg[0][12] ;
  assign \new_[4987]_  = \\u8_mem_reg[1][10] ;
  assign \new_[4988]_  = ~\new_[6237]_  | (~\new_[7689]_  & ~\new_[12801]_ );
  assign \new_[4989]_  = ~\new_[6241]_  | (~\new_[7690]_  & ~\new_[12755]_ );
  assign \new_[4990]_  = \\u7_mem_reg[3][7] ;
  assign \new_[4991]_  = \\u3_mem_reg[3][15] ;
  assign \new_[4992]_  = \\u3_mem_reg[3][11] ;
  assign \new_[4993]_  = \\u3_mem_reg[2][8] ;
  assign \new_[4994]_  = \\u7_mem_reg[0][12] ;
  assign \new_[4995]_  = \\u7_mem_reg[3][14] ;
  assign \new_[4996]_  = \\u7_mem_reg[3][25] ;
  assign \new_[4997]_  = \\u7_mem_reg[3][29] ;
  assign \new_[4998]_  = \\u3_mem_reg[2][26] ;
  assign \new_[4999]_  = \\u3_mem_reg[2][22] ;
  assign \new_[5000]_  = \\u3_mem_reg[2][18] ;
  assign \new_[5001]_  = \\u8_mem_reg[3][8] ;
  assign \new_[5002]_  = \\u8_mem_reg[3][6] ;
  assign \new_[5003]_  = \\u7_mem_reg[3][21] ;
  assign \new_[5004]_  = \\u7_mem_reg[3][18] ;
  assign \new_[5005]_  = \\u8_mem_reg[3][3] ;
  assign \new_[5006]_  = \\u3_mem_reg[2][11] ;
  assign \new_[5007]_  = \\u8_mem_reg[3][28] ;
  assign \new_[5008]_  = \\u7_mem_reg[0][17] ;
  assign \new_[5009]_  = \\u7_mem_reg[0][0] ;
  assign \new_[5010]_  = \\u8_mem_reg[3][22] ;
  assign \new_[5011]_  = \\u8_mem_reg[3][25] ;
  assign \new_[5012]_  = \\u7_mem_reg[2][25] ;
  assign \new_[5013]_  = \\u7_mem_reg[2][7] ;
  assign \new_[5014]_  = \\u7_mem_reg[3][10] ;
  assign \new_[5015]_  = \\u8_mem_reg[3][18] ;
  assign \new_[5016]_  = \\u3_mem_reg[1][3] ;
  assign \new_[5017]_  = \\u8_mem_reg[3][15] ;
  assign \new_[5018]_  = \\u8_mem_reg[3][10] ;
  assign \new_[5019]_  = \new_[13833]_  | \new_[13885]_ ;
  assign \new_[5020]_  = ~\new_[4591]_  | ~\new_[13885]_ ;
  assign \new_[5021]_  = \new_[13344]_  | \new_[13885]_ ;
  assign \new_[5022]_  = ~\new_[4648]_  | ~\new_[13885]_ ;
  assign \new_[5023]_  = \\u7_mem_reg[2][3] ;
  assign \new_[5024]_  = \\u7_mem_reg[2][29] ;
  assign \new_[5025]_  = \\u3_mem_reg[1][2] ;
  assign \new_[5026]_  = \\u7_mem_reg[2][21] ;
  assign \new_[5027]_  = \\u7_mem_reg[2][18] ;
  assign \new_[5028]_  = \\u6_mem_reg[0][30] ;
  assign \new_[5029]_  = \\u6_mem_reg[0][6] ;
  assign \new_[5030]_  = \\u7_mem_reg[2][14] ;
  assign \new_[5031]_  = \\u7_mem_reg[2][10] ;
  assign \new_[5032]_  = \\u8_mem_reg[2][6] ;
  assign \new_[5033]_  = \\u6_mem_reg[0][28] ;
  assign \new_[5034]_  = \\u7_mem_reg[1][7] ;
  assign \new_[5035]_  = \\u6_mem_reg[3][8] ;
  assign \new_[5036]_  = ~\\u13_crac_dout_r_reg[3] ;
  assign \new_[5037]_  = ~\\u13_crac_dout_r_reg[9] ;
  assign \new_[5038]_  = \\u7_mem_reg[1][3] ;
  assign \new_[5039]_  = \\u13_icc_r_reg[22] ;
  assign \new_[5040]_  = ~\\u13_crac_dout_r_reg[14] ;
  assign \new_[5041]_  = \\u13_occ0_r_reg[2] ;
  assign \new_[5042]_  = \\u13_occ0_r_reg[4] ;
  assign \new_[5043]_  = \\u13_intm_r_reg[7] ;
  assign \new_[5044]_  = \\u13_intm_r_reg[22] ;
  assign \new_[5045]_  = \\u13_icc_r_reg[11] ;
  assign \new_[5046]_  = \\u7_mem_reg[1][29] ;
  assign \new_[5047]_  = \\u6_mem_reg[0][23] ;
  assign \new_[5048]_  = \\u13_icc_r_reg[15] ;
  assign \new_[5049]_  = \\u13_icc_r_reg[19] ;
  assign \new_[5050]_  = \\u13_crac_r_reg[0] ;
  assign \new_[5051]_  = \\u13_crac_r_reg[1] ;
  assign \new_[5052]_  = \\u13_crac_r_reg[3] ;
  assign \new_[5053]_  = \\u13_crac_r_reg[4] ;
  assign \new_[5054]_  = \\u13_crac_r_reg[5] ;
  assign \new_[5055]_  = \\u13_crac_r_reg[7] ;
  assign \new_[5056]_  = \\u13_icc_r_reg[0] ;
  assign \new_[5057]_  = \\u13_icc_r_reg[10] ;
  assign \new_[5058]_  = \\u13_icc_r_reg[12] ;
  assign \new_[5059]_  = \\u13_icc_r_reg[13] ;
  assign \new_[5060]_  = \\u13_icc_r_reg[14] ;
  assign \new_[5061]_  = \\u13_icc_r_reg[16] ;
  assign \new_[5062]_  = \\u13_icc_r_reg[17] ;
  assign \new_[5063]_  = \\u13_icc_r_reg[18] ;
  assign \new_[5064]_  = \\u13_icc_r_reg[1] ;
  assign \new_[5065]_  = \\u13_icc_r_reg[20] ;
  assign \new_[5066]_  = \\u13_icc_r_reg[21] ;
  assign \new_[5067]_  = \\u13_icc_r_reg[23] ;
  assign \new_[5068]_  = \\u13_icc_r_reg[2] ;
  assign \new_[5069]_  = \\u13_icc_r_reg[3] ;
  assign \new_[5070]_  = \\u13_icc_r_reg[4] ;
  assign \new_[5071]_  = \\u13_icc_r_reg[5] ;
  assign \new_[5072]_  = \\u13_icc_r_reg[6] ;
  assign \new_[5073]_  = \\u13_icc_r_reg[7] ;
  assign \new_[5074]_  = \\u13_icc_r_reg[9] ;
  assign \new_[5075]_  = \\u13_occ0_r_reg[0] ;
  assign \new_[5076]_  = \\u13_occ0_r_reg[10] ;
  assign \new_[5077]_  = \\u13_occ0_r_reg[12] ;
  assign \new_[5078]_  = \\u13_occ0_r_reg[13] ;
  assign \new_[5079]_  = \\u13_occ0_r_reg[14] ;
  assign \new_[5080]_  = \\u13_occ0_r_reg[16] ;
  assign \new_[5081]_  = \\u13_occ0_r_reg[17] ;
  assign \new_[5082]_  = \\u13_occ0_r_reg[18] ;
  assign \new_[5083]_  = \\u13_occ0_r_reg[1] ;
  assign \new_[5084]_  = \\u13_occ0_r_reg[20] ;
  assign \new_[5085]_  = \\u13_occ0_r_reg[21] ;
  assign \new_[5086]_  = \\u13_occ0_r_reg[23] ;
  assign \new_[5087]_  = \\u13_occ0_r_reg[24] ;
  assign \new_[5088]_  = \\u13_occ0_r_reg[25] ;
  assign \new_[5089]_  = \\u13_occ0_r_reg[27] ;
  assign \new_[5090]_  = \\u13_occ0_r_reg[28] ;
  assign \new_[5091]_  = \\u13_occ0_r_reg[29] ;
  assign \new_[5092]_  = \\u13_occ0_r_reg[30] ;
  assign \new_[5093]_  = \\u13_occ0_r_reg[31] ;
  assign \new_[5094]_  = \\u13_occ0_r_reg[3] ;
  assign \new_[5095]_  = \\u13_occ0_r_reg[5] ;
  assign \new_[5096]_  = \\u13_occ0_r_reg[6] ;
  assign \new_[5097]_  = \\u13_occ0_r_reg[7] ;
  assign \new_[5098]_  = \\u13_occ0_r_reg[9] ;
  assign \new_[5099]_  = \\u13_intm_r_reg[0] ;
  assign \new_[5100]_  = \\u13_intm_r_reg[10] ;
  assign \new_[5101]_  = \\u13_intm_r_reg[11] ;
  assign \new_[5102]_  = \\u13_intm_r_reg[12] ;
  assign \new_[5103]_  = \\u13_intm_r_reg[13] ;
  assign \new_[5104]_  = \\u13_intm_r_reg[14] ;
  assign \new_[5105]_  = \\u13_intm_r_reg[16] ;
  assign \new_[5106]_  = \\u13_intm_r_reg[17] ;
  assign \new_[5107]_  = \\u13_intm_r_reg[18] ;
  assign \new_[5108]_  = \\u13_intm_r_reg[19] ;
  assign \new_[5109]_  = \\u13_intm_r_reg[1] ;
  assign \new_[5110]_  = \\u13_intm_r_reg[20] ;
  assign \new_[5111]_  = \\u13_intm_r_reg[21] ;
  assign \new_[5112]_  = \\u13_intm_r_reg[23] ;
  assign \new_[5113]_  = \\u13_intm_r_reg[24] ;
  assign \new_[5114]_  = \\u13_intm_r_reg[25] ;
  assign \new_[5115]_  = \\u13_intm_r_reg[27] ;
  assign \new_[5116]_  = \\u13_intm_r_reg[28] ;
  assign \new_[5117]_  = \\u13_intm_r_reg[2] ;
  assign \new_[5118]_  = \\u13_intm_r_reg[5] ;
  assign \new_[5119]_  = \\u13_intm_r_reg[6] ;
  assign \new_[5120]_  = \\u13_intm_r_reg[9] ;
  assign \new_[5121]_  = \\u13_intm_r_reg[4] ;
  assign \new_[5122]_  = \\u13_intm_r_reg[15] ;
  assign \new_[5123]_  = ~\\u13_crac_dout_r_reg[0] ;
  assign \new_[5124]_  = ~\\u13_crac_dout_r_reg[10] ;
  assign \new_[5125]_  = ~\\u13_crac_dout_r_reg[11] ;
  assign \new_[5126]_  = ~\\u13_crac_dout_r_reg[12] ;
  assign \new_[5127]_  = ~\\u13_crac_dout_r_reg[13] ;
  assign \new_[5128]_  = ~\\u13_crac_dout_r_reg[15] ;
  assign \new_[5129]_  = ~\\u13_crac_dout_r_reg[1] ;
  assign \new_[5130]_  = ~\\u13_crac_dout_r_reg[2] ;
  assign \new_[5131]_  = ~\\u13_crac_dout_r_reg[4] ;
  assign \new_[5132]_  = ~\\u13_crac_dout_r_reg[5] ;
  assign \new_[5133]_  = ~\\u13_crac_dout_r_reg[6] ;
  assign \new_[5134]_  = ~\\u13_crac_dout_r_reg[8] ;
  assign \new_[5135]_  = \\u8_mem_reg[2][4] ;
  assign \new_[5136]_  = \\u3_mem_reg[1][28] ;
  assign \new_[5137]_  = \\u8_mem_reg[2][5] ;
  assign \new_[5138]_  = \\u3_mem_reg[1][29] ;
  assign \new_[5139]_  = \\u8_mem_reg[2][7] ;
  assign \new_[5140]_  = \\u8_mem_reg[2][8] ;
  assign \new_[5141]_  = \\u8_mem_reg[2][9] ;
  assign \new_[5142]_  = \\u8_mem_reg[3][0] ;
  assign \new_[5143]_  = \\u3_mem_reg[1][30] ;
  assign \new_[5144]_  = \\u8_mem_reg[3][11] ;
  assign \new_[5145]_  = \\u3_mem_reg[1][31] ;
  assign \new_[5146]_  = \\u8_mem_reg[3][12] ;
  assign \new_[5147]_  = \\u8_mem_reg[3][13] ;
  assign \new_[5148]_  = \\u3_mem_reg[1][4] ;
  assign \new_[5149]_  = \\u8_mem_reg[3][14] ;
  assign \new_[5150]_  = \\u8_mem_reg[3][16] ;
  assign \new_[5151]_  = \\u8_mem_reg[3][17] ;
  assign \new_[5152]_  = \\u3_mem_reg[1][5] ;
  assign \new_[5153]_  = \\u8_mem_reg[3][19] ;
  assign \new_[5154]_  = \\u3_mem_reg[1][6] ;
  assign \new_[5155]_  = \\u8_mem_reg[3][1] ;
  assign \new_[5156]_  = \\u3_mem_reg[1][7] ;
  assign \new_[5157]_  = \\u8_mem_reg[3][20] ;
  assign \new_[5158]_  = \\u8_mem_reg[3][21] ;
  assign \new_[5159]_  = \\u3_mem_reg[1][8] ;
  assign \new_[5160]_  = \\u8_mem_reg[3][23] ;
  assign \new_[5161]_  = \\u8_mem_reg[3][24] ;
  assign \new_[5162]_  = \\u3_mem_reg[1][9] ;
  assign \new_[5163]_  = \\u8_mem_reg[3][26] ;
  assign \new_[5164]_  = \\u3_mem_reg[2][0] ;
  assign \new_[5165]_  = \\u8_mem_reg[3][27] ;
  assign \new_[5166]_  = \\u3_mem_reg[2][10] ;
  assign \new_[5167]_  = \\u8_mem_reg[3][29] ;
  assign \new_[5168]_  = \\u8_mem_reg[3][2] ;
  assign \new_[5169]_  = \\u8_mem_reg[3][30] ;
  assign \new_[5170]_  = \\u8_mem_reg[3][31] ;
  assign \new_[5171]_  = \\u3_mem_reg[2][12] ;
  assign \new_[5172]_  = \\u8_mem_reg[3][4] ;
  assign \new_[5173]_  = \\u3_mem_reg[2][13] ;
  assign \new_[5174]_  = \\u8_mem_reg[3][5] ;
  assign \new_[5175]_  = \\u3_mem_reg[2][14] ;
  assign \new_[5176]_  = \\u8_mem_reg[3][7] ;
  assign \new_[5177]_  = \\u3_mem_reg[2][15] ;
  assign \new_[5178]_  = \\u8_mem_reg[3][9] ;
  assign \new_[5179]_  = \\u3_mem_reg[2][16] ;
  assign \new_[5180]_  = \\u3_mem_reg[2][17] ;
  assign \new_[5181]_  = \\u3_mem_reg[2][19] ;
  assign \new_[5182]_  = \\u3_mem_reg[2][1] ;
  assign \new_[5183]_  = \\u3_mem_reg[2][21] ;
  assign \new_[5184]_  = \\u3_mem_reg[2][23] ;
  assign \new_[5185]_  = \\u3_mem_reg[2][24] ;
  assign \new_[5186]_  = \\u3_mem_reg[2][25] ;
  assign \new_[5187]_  = \\u3_mem_reg[2][27] ;
  assign \new_[5188]_  = \\u3_mem_reg[2][28] ;
  assign \new_[5189]_  = \\u3_mem_reg[2][29] ;
  assign \new_[5190]_  = \\u3_mem_reg[2][30] ;
  assign \new_[5191]_  = \\u3_mem_reg[2][31] ;
  assign \new_[5192]_  = \\u3_mem_reg[2][3] ;
  assign \new_[5193]_  = \\u3_mem_reg[2][4] ;
  assign \new_[5194]_  = \\u3_mem_reg[2][5] ;
  assign \new_[5195]_  = \\u3_mem_reg[2][6] ;
  assign \new_[5196]_  = \\u3_mem_reg[2][7] ;
  assign \new_[5197]_  = \\u3_mem_reg[2][9] ;
  assign \new_[5198]_  = \\u3_mem_reg[3][0] ;
  assign \new_[5199]_  = \\u3_mem_reg[3][10] ;
  assign \new_[5200]_  = \\u3_mem_reg[3][12] ;
  assign \new_[5201]_  = \\u3_mem_reg[3][13] ;
  assign \new_[5202]_  = \\u3_mem_reg[3][14] ;
  assign \new_[5203]_  = \\u3_mem_reg[3][16] ;
  assign \new_[5204]_  = \\u3_mem_reg[3][17] ;
  assign \new_[5205]_  = \\u3_mem_reg[3][18] ;
  assign \new_[5206]_  = \\u3_mem_reg[3][1] ;
  assign \new_[5207]_  = \\u3_mem_reg[3][20] ;
  assign \new_[5208]_  = \\u3_mem_reg[3][21] ;
  assign \new_[5209]_  = \\u3_mem_reg[3][23] ;
  assign \new_[5210]_  = \\u3_mem_reg[3][24] ;
  assign \new_[5211]_  = \\u3_mem_reg[3][26] ;
  assign \new_[5212]_  = \\u3_mem_reg[3][28] ;
  assign \new_[5213]_  = \\u3_mem_reg[3][29] ;
  assign \new_[5214]_  = \\u3_mem_reg[3][2] ;
  assign \new_[5215]_  = \\u3_mem_reg[3][31] ;
  assign \new_[5216]_  = \\u3_mem_reg[3][4] ;
  assign \new_[5217]_  = \\u3_mem_reg[3][5] ;
  assign \new_[5218]_  = \\u3_mem_reg[3][7] ;
  assign \new_[5219]_  = \\u3_mem_reg[3][9] ;
  assign \new_[5220]_  = \\u3_mem_reg[3][25] ;
  assign \new_[5221]_  = \\u4_mem_reg[1][0] ;
  assign \new_[5222]_  = \\u4_mem_reg[1][10] ;
  assign \new_[5223]_  = \\u4_mem_reg[1][11] ;
  assign \new_[5224]_  = \\u4_mem_reg[1][13] ;
  assign \new_[5225]_  = \\u4_mem_reg[1][14] ;
  assign \new_[5226]_  = \\u4_mem_reg[1][15] ;
  assign \new_[5227]_  = \\u4_mem_reg[1][17] ;
  assign \new_[5228]_  = \\u4_mem_reg[1][18] ;
  assign \new_[5229]_  = \\u4_mem_reg[1][19] ;
  assign \new_[5230]_  = \\u4_mem_reg[1][1] ;
  assign \new_[5231]_  = \\u4_mem_reg[1][20] ;
  assign \new_[5232]_  = \\u4_mem_reg[1][21] ;
  assign \new_[5233]_  = \\u4_mem_reg[1][22] ;
  assign \new_[5234]_  = \\u4_mem_reg[1][24] ;
  assign \new_[5235]_  = \\u4_mem_reg[1][25] ;
  assign \new_[5236]_  = \\u4_mem_reg[1][26] ;
  assign \new_[5237]_  = \\u4_mem_reg[1][28] ;
  assign \new_[5238]_  = \\u4_mem_reg[1][29] ;
  assign \new_[5239]_  = \\u4_mem_reg[1][2] ;
  assign \new_[5240]_  = \\u4_mem_reg[1][31] ;
  assign \new_[5241]_  = \\u4_mem_reg[1][3] ;
  assign \new_[5242]_  = \\u4_mem_reg[1][4] ;
  assign \new_[5243]_  = \\u4_mem_reg[1][6] ;
  assign \new_[5244]_  = \\u4_mem_reg[1][7] ;
  assign \new_[5245]_  = \\u4_mem_reg[1][8] ;
  assign \new_[5246]_  = \\u4_mem_reg[2][0] ;
  assign \new_[5247]_  = \\u4_mem_reg[2][10] ;
  assign \new_[5248]_  = \\u4_mem_reg[2][11] ;
  assign \new_[5249]_  = \\u4_mem_reg[2][13] ;
  assign \new_[5250]_  = \\u4_mem_reg[2][14] ;
  assign \new_[5251]_  = \\u4_mem_reg[2][15] ;
  assign \new_[5252]_  = \\u4_mem_reg[2][17] ;
  assign \new_[5253]_  = \\u4_mem_reg[2][18] ;
  assign \new_[5254]_  = \\u4_mem_reg[2][19] ;
  assign \new_[5255]_  = \\u4_mem_reg[2][1] ;
  assign \new_[5256]_  = \\u4_mem_reg[2][20] ;
  assign \new_[5257]_  = \\u4_mem_reg[2][21] ;
  assign \new_[5258]_  = \\u4_mem_reg[2][22] ;
  assign \new_[5259]_  = \\u4_mem_reg[2][24] ;
  assign \new_[5260]_  = \\u4_mem_reg[2][25] ;
  assign \new_[5261]_  = \\u4_mem_reg[2][26] ;
  assign \new_[5262]_  = \\u4_mem_reg[2][28] ;
  assign \new_[5263]_  = \\u4_mem_reg[2][29] ;
  assign \new_[5264]_  = \\u4_mem_reg[2][2] ;
  assign \new_[5265]_  = \\u4_mem_reg[2][31] ;
  assign \new_[5266]_  = \\u4_mem_reg[2][3] ;
  assign \new_[5267]_  = \\u4_mem_reg[2][4] ;
  assign \new_[5268]_  = \\u4_mem_reg[2][6] ;
  assign \new_[5269]_  = \\u4_mem_reg[2][7] ;
  assign \new_[5270]_  = \\u4_mem_reg[2][8] ;
  assign \new_[5271]_  = \\u4_mem_reg[3][0] ;
  assign \new_[5272]_  = \\u4_mem_reg[3][10] ;
  assign \new_[5273]_  = \\u4_mem_reg[3][11] ;
  assign \new_[5274]_  = \\u4_mem_reg[3][13] ;
  assign \new_[5275]_  = \\u4_mem_reg[3][14] ;
  assign \new_[5276]_  = \\u4_mem_reg[3][15] ;
  assign \new_[5277]_  = \\u4_mem_reg[3][17] ;
  assign \new_[5278]_  = \\u4_mem_reg[3][18] ;
  assign \new_[5279]_  = \\u4_mem_reg[3][19] ;
  assign \new_[5280]_  = \\u4_mem_reg[3][1] ;
  assign \new_[5281]_  = \\u4_mem_reg[3][20] ;
  assign \new_[5282]_  = \\u4_mem_reg[3][21] ;
  assign \new_[5283]_  = \\u4_mem_reg[3][22] ;
  assign \new_[5284]_  = \\u4_mem_reg[3][24] ;
  assign \new_[5285]_  = \\u4_mem_reg[3][25] ;
  assign \new_[5286]_  = \\u4_mem_reg[3][26] ;
  assign \new_[5287]_  = \\u4_mem_reg[3][28] ;
  assign \new_[5288]_  = \\u4_mem_reg[3][29] ;
  assign \new_[5289]_  = \\u4_mem_reg[3][2] ;
  assign \new_[5290]_  = \\u4_mem_reg[3][31] ;
  assign \new_[5291]_  = \\u4_mem_reg[3][3] ;
  assign \new_[5292]_  = \\u4_mem_reg[3][4] ;
  assign \new_[5293]_  = \\u4_mem_reg[3][6] ;
  assign \new_[5294]_  = \\u4_mem_reg[3][7] ;
  assign \new_[5295]_  = \\u4_mem_reg[3][8] ;
  assign \new_[5296]_  = \\u3_mem_reg[2][20] ;
  assign \new_[5297]_  = \\u5_mem_reg[1][0] ;
  assign \new_[5298]_  = \\u5_mem_reg[1][10] ;
  assign \new_[5299]_  = \\u5_mem_reg[1][12] ;
  assign \new_[5300]_  = \\u5_mem_reg[1][13] ;
  assign \new_[5301]_  = \\u5_mem_reg[1][14] ;
  assign \new_[5302]_  = \\u7_mem_reg[1][14] ;
  assign \new_[5303]_  = \\u5_mem_reg[1][16] ;
  assign \new_[5304]_  = \\u5_mem_reg[1][17] ;
  assign \new_[5305]_  = \\u5_mem_reg[1][18] ;
  assign \new_[5306]_  = \\u5_mem_reg[1][1] ;
  assign \new_[5307]_  = \\u5_mem_reg[1][20] ;
  assign \new_[5308]_  = \\u5_mem_reg[1][21] ;
  assign \new_[5309]_  = \\u5_mem_reg[1][23] ;
  assign \new_[5310]_  = \\u5_mem_reg[1][24] ;
  assign \new_[5311]_  = \\u5_mem_reg[1][25] ;
  assign \new_[5312]_  = \\u5_mem_reg[1][27] ;
  assign \new_[5313]_  = \\u5_mem_reg[1][28] ;
  assign \new_[5314]_  = \\u5_mem_reg[1][29] ;
  assign \new_[5315]_  = \\u5_mem_reg[1][30] ;
  assign \new_[5316]_  = \\u5_mem_reg[1][31] ;
  assign \new_[5317]_  = \\u5_mem_reg[1][3] ;
  assign \new_[5318]_  = \\u5_mem_reg[1][5] ;
  assign \new_[5319]_  = \\u5_mem_reg[1][6] ;
  assign \new_[5320]_  = \\u5_mem_reg[1][7] ;
  assign \new_[5321]_  = \\u5_mem_reg[1][9] ;
  assign \new_[5322]_  = \\u5_mem_reg[2][0] ;
  assign \new_[5323]_  = \\u5_mem_reg[2][10] ;
  assign \new_[5324]_  = \\u5_mem_reg[2][12] ;
  assign \new_[5325]_  = \\u5_mem_reg[2][13] ;
  assign \new_[5326]_  = \\u5_mem_reg[2][14] ;
  assign \new_[5327]_  = \\u5_mem_reg[2][16] ;
  assign \new_[5328]_  = \\u5_mem_reg[2][17] ;
  assign \new_[5329]_  = \\u5_mem_reg[2][18] ;
  assign \new_[5330]_  = \\u5_mem_reg[2][1] ;
  assign \new_[5331]_  = \\u5_mem_reg[2][20] ;
  assign \new_[5332]_  = \\u5_mem_reg[2][21] ;
  assign \new_[5333]_  = \\u5_mem_reg[2][23] ;
  assign \new_[5334]_  = \\u5_mem_reg[2][24] ;
  assign \new_[5335]_  = \\u5_mem_reg[2][25] ;
  assign \new_[5336]_  = \\u5_mem_reg[2][27] ;
  assign \new_[5337]_  = \\u5_mem_reg[2][28] ;
  assign \new_[5338]_  = \\u5_mem_reg[2][29] ;
  assign \new_[5339]_  = \\u5_mem_reg[2][30] ;
  assign \new_[5340]_  = \\u5_mem_reg[2][31] ;
  assign \new_[5341]_  = \\u5_mem_reg[2][3] ;
  assign \new_[5342]_  = \\u5_mem_reg[2][4] ;
  assign \new_[5343]_  = \\u5_mem_reg[2][5] ;
  assign \new_[5344]_  = \\u5_mem_reg[2][6] ;
  assign \new_[5345]_  = \\u5_mem_reg[2][7] ;
  assign \new_[5346]_  = \\u5_mem_reg[2][9] ;
  assign \new_[5347]_  = \\u5_mem_reg[3][0] ;
  assign \new_[5348]_  = \\u5_mem_reg[3][10] ;
  assign \new_[5349]_  = \\u5_mem_reg[3][12] ;
  assign \new_[5350]_  = \\u5_mem_reg[3][13] ;
  assign \new_[5351]_  = \\u5_mem_reg[3][14] ;
  assign \new_[5352]_  = \\u5_mem_reg[3][16] ;
  assign \new_[5353]_  = \\u5_mem_reg[3][17] ;
  assign \new_[5354]_  = \\u5_mem_reg[3][18] ;
  assign \new_[5355]_  = \\u5_mem_reg[3][1] ;
  assign \new_[5356]_  = \\u5_mem_reg[3][20] ;
  assign \new_[5357]_  = \\u5_mem_reg[3][21] ;
  assign \new_[5358]_  = \\u6_mem_reg[0][17] ;
  assign \new_[5359]_  = \\u5_mem_reg[3][23] ;
  assign \new_[5360]_  = \\u5_mem_reg[3][24] ;
  assign \new_[5361]_  = \\u5_mem_reg[3][25] ;
  assign \new_[5362]_  = \\u5_mem_reg[3][27] ;
  assign \new_[5363]_  = \\u5_mem_reg[3][28] ;
  assign \new_[5364]_  = \\u5_mem_reg[3][29] ;
  assign \new_[5365]_  = \\u5_mem_reg[3][30] ;
  assign \new_[5366]_  = \\u5_mem_reg[3][31] ;
  assign \new_[5367]_  = \\u5_mem_reg[3][3] ;
  assign \new_[5368]_  = \\u5_mem_reg[3][5] ;
  assign \new_[5369]_  = \\u5_mem_reg[3][6] ;
  assign \new_[5370]_  = \\u5_mem_reg[3][7] ;
  assign \new_[5371]_  = \\u5_mem_reg[3][9] ;
  assign \new_[5372]_  = \\u6_mem_reg[1][0] ;
  assign \new_[5373]_  = \\u6_mem_reg[1][10] ;
  assign \new_[5374]_  = \\u6_mem_reg[1][12] ;
  assign \new_[5375]_  = \\u6_mem_reg[1][13] ;
  assign \new_[5376]_  = \\u6_mem_reg[1][14] ;
  assign \new_[5377]_  = \\u6_mem_reg[1][16] ;
  assign \new_[5378]_  = \\u6_mem_reg[1][17] ;
  assign \new_[5379]_  = \\u6_mem_reg[1][18] ;
  assign \new_[5380]_  = \\u6_mem_reg[1][19] ;
  assign \new_[5381]_  = \\u6_mem_reg[1][1] ;
  assign \new_[5382]_  = \\u6_mem_reg[1][20] ;
  assign \new_[5383]_  = \\u6_mem_reg[1][21] ;
  assign \new_[5384]_  = \\u6_mem_reg[1][23] ;
  assign \new_[5385]_  = \\u6_mem_reg[1][24] ;
  assign \new_[5386]_  = \\u6_mem_reg[1][25] ;
  assign \new_[5387]_  = \\u6_mem_reg[1][27] ;
  assign \new_[5388]_  = \\u6_mem_reg[1][28] ;
  assign \new_[5389]_  = \\u6_mem_reg[1][29] ;
  assign \new_[5390]_  = \\u6_mem_reg[1][30] ;
  assign \new_[5391]_  = \\u6_mem_reg[1][31] ;
  assign \new_[5392]_  = \\u6_mem_reg[1][3] ;
  assign \new_[5393]_  = \\u6_mem_reg[1][5] ;
  assign \new_[5394]_  = \\u6_mem_reg[1][6] ;
  assign \new_[5395]_  = \\u6_mem_reg[1][7] ;
  assign \new_[5396]_  = \\u6_mem_reg[1][9] ;
  assign \new_[5397]_  = \\u6_mem_reg[2][0] ;
  assign \new_[5398]_  = \\u6_mem_reg[2][10] ;
  assign \new_[5399]_  = \\u6_mem_reg[2][12] ;
  assign \new_[5400]_  = \\u6_mem_reg[2][13] ;
  assign \new_[5401]_  = \\u6_mem_reg[2][14] ;
  assign \new_[5402]_  = \\u6_mem_reg[2][16] ;
  assign \new_[5403]_  = \\u6_mem_reg[2][17] ;
  assign \new_[5404]_  = \\u6_mem_reg[2][18] ;
  assign \new_[5405]_  = \\u6_mem_reg[2][1] ;
  assign \new_[5406]_  = \\u6_mem_reg[2][20] ;
  assign \new_[5407]_  = \\u6_mem_reg[2][21] ;
  assign \new_[5408]_  = \\u6_mem_reg[2][23] ;
  assign \new_[5409]_  = \\u6_mem_reg[2][24] ;
  assign \new_[5410]_  = \\u6_mem_reg[2][25] ;
  assign \new_[5411]_  = \\u6_mem_reg[2][27] ;
  assign \new_[5412]_  = \\u6_mem_reg[2][28] ;
  assign \new_[5413]_  = \\u6_mem_reg[2][29] ;
  assign \new_[5414]_  = \\u6_mem_reg[2][30] ;
  assign \new_[5415]_  = \\u6_mem_reg[2][31] ;
  assign \new_[5416]_  = \\u6_mem_reg[2][3] ;
  assign \new_[5417]_  = \\u6_mem_reg[2][5] ;
  assign \new_[5418]_  = \\u6_mem_reg[2][6] ;
  assign \new_[5419]_  = \\u6_mem_reg[2][7] ;
  assign \new_[5420]_  = \\u6_mem_reg[2][9] ;
  assign \new_[5421]_  = \\u6_mem_reg[3][0] ;
  assign \new_[5422]_  = \\u6_mem_reg[3][10] ;
  assign \new_[5423]_  = \\u6_mem_reg[3][12] ;
  assign \new_[5424]_  = \\u6_mem_reg[3][13] ;
  assign \new_[5425]_  = \\u6_mem_reg[3][14] ;
  assign \new_[5426]_  = \\u6_mem_reg[3][16] ;
  assign \new_[5427]_  = \\u6_mem_reg[3][17] ;
  assign \new_[5428]_  = \\u6_mem_reg[3][18] ;
  assign \new_[5429]_  = \\u6_mem_reg[3][1] ;
  assign \new_[5430]_  = \\u6_mem_reg[3][20] ;
  assign \new_[5431]_  = \\u6_mem_reg[3][21] ;
  assign \new_[5432]_  = \\u6_mem_reg[3][23] ;
  assign \new_[5433]_  = \\u6_mem_reg[3][24] ;
  assign \new_[5434]_  = \\u6_mem_reg[3][25] ;
  assign \new_[5435]_  = \\u6_mem_reg[3][27] ;
  assign \new_[5436]_  = \\u6_mem_reg[3][28] ;
  assign \new_[5437]_  = \\u6_mem_reg[3][29] ;
  assign \new_[5438]_  = \\u6_mem_reg[3][30] ;
  assign \new_[5439]_  = \\u6_mem_reg[3][31] ;
  assign \new_[5440]_  = \\u6_mem_reg[3][3] ;
  assign \new_[5441]_  = \\u6_mem_reg[3][5] ;
  assign \new_[5442]_  = \\u6_mem_reg[3][6] ;
  assign \new_[5443]_  = \\u6_mem_reg[3][7] ;
  assign \new_[5444]_  = \\u6_mem_reg[3][9] ;
  assign \new_[5445]_  = \\u3_mem_reg[3][8] ;
  assign \new_[5446]_  = \\u7_mem_reg[1][0] ;
  assign \new_[5447]_  = \\u7_mem_reg[1][11] ;
  assign \new_[5448]_  = \\u7_mem_reg[1][12] ;
  assign \new_[5449]_  = \\u7_mem_reg[1][13] ;
  assign \new_[5450]_  = \\u7_mem_reg[1][15] ;
  assign \new_[5451]_  = \\u7_mem_reg[1][16] ;
  assign \new_[5452]_  = \\u7_mem_reg[1][17] ;
  assign \new_[5453]_  = \\u7_mem_reg[1][18] ;
  assign \new_[5454]_  = \\u7_mem_reg[1][19] ;
  assign \new_[5455]_  = \\u7_mem_reg[1][1] ;
  assign \new_[5456]_  = \\u7_mem_reg[1][20] ;
  assign \new_[5457]_  = \\u7_mem_reg[1][22] ;
  assign \new_[5458]_  = \\u7_mem_reg[1][23] ;
  assign \new_[5459]_  = \\u7_mem_reg[1][24] ;
  assign \new_[5460]_  = \\u7_mem_reg[1][26] ;
  assign \new_[5461]_  = \\u7_mem_reg[1][27] ;
  assign \new_[5462]_  = \\u7_mem_reg[1][28] ;
  assign \new_[5463]_  = \\u7_mem_reg[1][2] ;
  assign \new_[5464]_  = \\u7_mem_reg[1][30] ;
  assign \new_[5465]_  = \\u7_mem_reg[1][31] ;
  assign \new_[5466]_  = \\u7_mem_reg[1][4] ;
  assign \new_[5467]_  = \\u7_mem_reg[1][5] ;
  assign \new_[5468]_  = \\u7_mem_reg[1][6] ;
  assign \new_[5469]_  = \\u7_mem_reg[1][8] ;
  assign \new_[5470]_  = \\u7_mem_reg[1][9] ;
  assign \new_[5471]_  = \\u7_mem_reg[2][0] ;
  assign \new_[5472]_  = \\u7_mem_reg[2][11] ;
  assign \new_[5473]_  = \\u7_mem_reg[2][12] ;
  assign \new_[5474]_  = \\u7_mem_reg[2][13] ;
  assign \new_[5475]_  = \\u7_mem_reg[2][15] ;
  assign \new_[5476]_  = \\u7_mem_reg[2][16] ;
  assign \new_[5477]_  = \\u7_mem_reg[2][17] ;
  assign \new_[5478]_  = \\u7_mem_reg[2][19] ;
  assign \new_[5479]_  = \\u7_mem_reg[2][1] ;
  assign \new_[5480]_  = \\u7_mem_reg[2][20] ;
  assign \new_[5481]_  = \\u7_mem_reg[2][22] ;
  assign \new_[5482]_  = \\u7_mem_reg[2][23] ;
  assign \new_[5483]_  = \\u7_mem_reg[2][24] ;
  assign \new_[5484]_  = \\u7_mem_reg[2][26] ;
  assign \new_[5485]_  = \\u7_mem_reg[2][27] ;
  assign \new_[5486]_  = \\u7_mem_reg[2][28] ;
  assign \new_[5487]_  = \\u7_mem_reg[2][2] ;
  assign \new_[5488]_  = \\u7_mem_reg[2][30] ;
  assign \new_[5489]_  = \\u7_mem_reg[2][31] ;
  assign \new_[5490]_  = \\u7_mem_reg[2][4] ;
  assign \new_[5491]_  = \\u7_mem_reg[2][5] ;
  assign \new_[5492]_  = \\u7_mem_reg[2][6] ;
  assign \new_[5493]_  = \\u7_mem_reg[2][8] ;
  assign \new_[5494]_  = \\u7_mem_reg[2][9] ;
  assign \new_[5495]_  = \\u7_mem_reg[3][0] ;
  assign \new_[5496]_  = \\u7_mem_reg[3][11] ;
  assign \new_[5497]_  = \\u7_mem_reg[3][12] ;
  assign \new_[5498]_  = \\u7_mem_reg[3][13] ;
  assign \new_[5499]_  = \\u7_mem_reg[3][15] ;
  assign \new_[5500]_  = \\u7_mem_reg[3][16] ;
  assign \new_[5501]_  = \\u7_mem_reg[3][17] ;
  assign \new_[5502]_  = \\u7_mem_reg[3][19] ;
  assign \new_[5503]_  = \\u7_mem_reg[3][1] ;
  assign \new_[5504]_  = \\u7_mem_reg[3][20] ;
  assign \new_[5505]_  = \\u6_mem_reg[0][20] ;
  assign \new_[5506]_  = \\u7_mem_reg[3][22] ;
  assign \new_[5507]_  = \\u7_mem_reg[3][23] ;
  assign \new_[5508]_  = \\u7_mem_reg[3][24] ;
  assign \new_[5509]_  = \\u7_mem_reg[3][26] ;
  assign \new_[5510]_  = \\u7_mem_reg[3][27] ;
  assign \new_[5511]_  = \\u7_mem_reg[3][28] ;
  assign \new_[5512]_  = \\u7_mem_reg[3][2] ;
  assign \new_[5513]_  = \\u7_mem_reg[3][30] ;
  assign \new_[5514]_  = \\u7_mem_reg[3][31] ;
  assign \new_[5515]_  = \\u7_mem_reg[3][4] ;
  assign \new_[5516]_  = \\u7_mem_reg[3][5] ;
  assign \new_[5517]_  = \\u7_mem_reg[3][6] ;
  assign \new_[5518]_  = \\u7_mem_reg[3][8] ;
  assign \new_[5519]_  = \\u7_mem_reg[3][9] ;
  assign \new_[5520]_  = \\u8_mem_reg[1][0] ;
  assign \new_[5521]_  = \\u8_mem_reg[1][11] ;
  assign \new_[5522]_  = \\u8_mem_reg[1][12] ;
  assign \new_[5523]_  = \\u8_mem_reg[1][13] ;
  assign \new_[5524]_  = \\u8_mem_reg[1][15] ;
  assign \new_[5525]_  = \\u8_mem_reg[1][16] ;
  assign \new_[5526]_  = \\u8_mem_reg[1][17] ;
  assign \new_[5527]_  = \\u8_mem_reg[1][19] ;
  assign \new_[5528]_  = \\u8_mem_reg[1][1] ;
  assign \new_[5529]_  = \\u8_mem_reg[1][20] ;
  assign \new_[5530]_  = \\u8_mem_reg[1][22] ;
  assign \new_[5531]_  = \\u8_mem_reg[1][23] ;
  assign \new_[5532]_  = \\u8_mem_reg[1][24] ;
  assign \new_[5533]_  = \\u8_mem_reg[1][26] ;
  assign \new_[5534]_  = \\u3_mem_reg[1][0] ;
  assign \new_[5535]_  = \\u8_mem_reg[1][27] ;
  assign \new_[5536]_  = \\u3_mem_reg[1][10] ;
  assign \new_[5537]_  = \\u8_mem_reg[1][29] ;
  assign \new_[5538]_  = \\u8_mem_reg[1][2] ;
  assign \new_[5539]_  = \\u8_mem_reg[1][30] ;
  assign \new_[5540]_  = \\u8_mem_reg[1][31] ;
  assign \new_[5541]_  = \\u3_mem_reg[1][12] ;
  assign \new_[5542]_  = \\u8_mem_reg[1][4] ;
  assign \new_[5543]_  = \\u3_mem_reg[1][13] ;
  assign \new_[5544]_  = \\u8_mem_reg[1][5] ;
  assign \new_[5545]_  = \\u3_mem_reg[1][14] ;
  assign \new_[5546]_  = \\u8_mem_reg[1][7] ;
  assign \new_[5547]_  = \\u8_mem_reg[1][8] ;
  assign \new_[5548]_  = \\u8_mem_reg[1][9] ;
  assign \new_[5549]_  = \\u8_mem_reg[2][0] ;
  assign \new_[5550]_  = \\u3_mem_reg[1][16] ;
  assign \new_[5551]_  = \\u8_mem_reg[2][10] ;
  assign \new_[5552]_  = \\u8_mem_reg[2][11] ;
  assign \new_[5553]_  = \\u3_mem_reg[1][17] ;
  assign \new_[5554]_  = \\u8_mem_reg[2][12] ;
  assign \new_[5555]_  = \\u3_mem_reg[1][18] ;
  assign \new_[5556]_  = \\u8_mem_reg[2][14] ;
  assign \new_[5557]_  = \\u8_mem_reg[2][15] ;
  assign \new_[5558]_  = \\u8_mem_reg[2][16] ;
  assign \new_[5559]_  = \\u8_mem_reg[2][17] ;
  assign \new_[5560]_  = \\u3_mem_reg[1][1] ;
  assign \new_[5561]_  = \\u8_mem_reg[2][19] ;
  assign \new_[5562]_  = \\u3_mem_reg[1][20] ;
  assign \new_[5563]_  = \\u8_mem_reg[2][1] ;
  assign \new_[5564]_  = \\u3_mem_reg[1][21] ;
  assign \new_[5565]_  = \\u8_mem_reg[2][21] ;
  assign \new_[5566]_  = \\u8_mem_reg[2][22] ;
  assign \new_[5567]_  = \\u8_mem_reg[2][23] ;
  assign \new_[5568]_  = \\u8_mem_reg[2][24] ;
  assign \new_[5569]_  = \\u3_mem_reg[1][23] ;
  assign \new_[5570]_  = \\u8_mem_reg[2][26] ;
  assign \new_[5571]_  = \\u3_mem_reg[1][24] ;
  assign \new_[5572]_  = \\u8_mem_reg[2][27] ;
  assign \new_[5573]_  = \\u3_mem_reg[1][25] ;
  assign \new_[5574]_  = \\u8_mem_reg[2][29] ;
  assign \new_[5575]_  = \\u8_mem_reg[2][2] ;
  assign \new_[5576]_  = \\u8_mem_reg[2][30] ;
  assign \new_[5577]_  = \\u8_mem_reg[2][31] ;
  assign \new_[5578]_  = \\u3_mem_reg[1][27] ;
  assign \new_[5579]_  = \\u4_mem_reg[0][0] ;
  assign \new_[5580]_  = \\u4_mem_reg[0][10] ;
  assign \new_[5581]_  = \\u4_mem_reg[0][11] ;
  assign \new_[5582]_  = \\u4_mem_reg[0][15] ;
  assign \new_[5583]_  = \\u4_mem_reg[0][18] ;
  assign \new_[5584]_  = \\u4_mem_reg[0][1] ;
  assign \new_[5585]_  = \\u4_mem_reg[0][21] ;
  assign \new_[5586]_  = \\u4_mem_reg[0][25] ;
  assign \new_[5587]_  = \\u4_mem_reg[0][27] ;
  assign \new_[5588]_  = \\u4_mem_reg[0][28] ;
  assign \new_[5589]_  = \\u4_mem_reg[0][26] ;
  assign \new_[5590]_  = \\u4_mem_reg[0][2] ;
  assign \new_[5591]_  = \\u4_mem_reg[0][29] ;
  assign \new_[5592]_  = \\u4_mem_reg[0][3] ;
  assign \new_[5593]_  = \\u4_mem_reg[0][5] ;
  assign \new_[5594]_  = \\u4_mem_reg[0][8] ;
  assign \new_[5595]_  = \\u5_mem_reg[0][10] ;
  assign \new_[5596]_  = \\u5_mem_reg[0][11] ;
  assign \new_[5597]_  = \\u5_mem_reg[0][15] ;
  assign \new_[5598]_  = \\u5_mem_reg[0][18] ;
  assign \new_[5599]_  = \\u5_mem_reg[0][1] ;
  assign \new_[5600]_  = \\u5_mem_reg[0][21] ;
  assign \new_[5601]_  = \\u13_intm_r_reg[8] ;
  assign \new_[5602]_  = \\u5_mem_reg[0][26] ;
  assign \new_[5603]_  = \\u5_mem_reg[0][27] ;
  assign \new_[5604]_  = \\u5_mem_reg[0][25] ;
  assign \new_[5605]_  = \\u5_mem_reg[0][2] ;
  assign \new_[5606]_  = \\u5_mem_reg[0][29] ;
  assign \new_[5607]_  = \\u5_mem_reg[0][3] ;
  assign \new_[5608]_  = \\u5_mem_reg[0][5] ;
  assign \new_[5609]_  = \\u5_mem_reg[0][8] ;
  assign \new_[5610]_  = \\u6_mem_reg[0][10] ;
  assign \new_[5611]_  = \\u6_mem_reg[0][11] ;
  assign \new_[5612]_  = \\u6_mem_reg[0][15] ;
  assign \new_[5613]_  = \\u7_mem_reg[1][21] ;
  assign \new_[5614]_  = \\u6_mem_reg[0][18] ;
  assign \new_[5615]_  = \\u6_mem_reg[0][1] ;
  assign \new_[5616]_  = \\u6_mem_reg[0][21] ;
  assign \new_[5617]_  = \\u6_mem_reg[0][26] ;
  assign \new_[5618]_  = \\u6_mem_reg[0][27] ;
  assign \new_[5619]_  = \\u6_mem_reg[0][25] ;
  assign \new_[5620]_  = \\u6_mem_reg[0][2] ;
  assign \new_[5621]_  = \\u6_mem_reg[0][29] ;
  assign \new_[5622]_  = \\u6_mem_reg[0][3] ;
  assign \new_[5623]_  = \\u6_mem_reg[0][5] ;
  assign \new_[5624]_  = \\u6_mem_reg[0][8] ;
  assign \new_[5625]_  = \\u7_mem_reg[0][10] ;
  assign \new_[5626]_  = \\u7_mem_reg[0][11] ;
  assign \new_[5627]_  = \\u7_mem_reg[0][15] ;
  assign \new_[5628]_  = \\u7_mem_reg[0][18] ;
  assign \new_[5629]_  = \\u7_mem_reg[0][1] ;
  assign \new_[5630]_  = \\u7_mem_reg[0][21] ;
  assign \new_[5631]_  = \\u7_mem_reg[0][25] ;
  assign \new_[5632]_  = \\u7_mem_reg[0][27] ;
  assign \new_[5633]_  = \\u7_mem_reg[0][28] ;
  assign \new_[5634]_  = \\u7_mem_reg[0][26] ;
  assign \new_[5635]_  = \\u7_mem_reg[0][2] ;
  assign \new_[5636]_  = \\u7_mem_reg[0][29] ;
  assign \new_[5637]_  = \\u7_mem_reg[0][3] ;
  assign \new_[5638]_  = \\u7_mem_reg[0][5] ;
  assign \new_[5639]_  = \\u7_mem_reg[0][8] ;
  assign \new_[5640]_  = \\u3_mem_reg[0][10] ;
  assign \new_[5641]_  = \\u8_mem_reg[0][10] ;
  assign \new_[5642]_  = \\u8_mem_reg[0][13] ;
  assign \new_[5643]_  = \\u3_mem_reg[0][18] ;
  assign \new_[5644]_  = \\u8_mem_reg[0][14] ;
  assign \new_[5645]_  = \\u3_mem_reg[0][19] ;
  assign \new_[5646]_  = \\u8_mem_reg[0][18] ;
  assign \new_[5647]_  = \\u8_mem_reg[0][19] ;
  assign \new_[5648]_  = \\u3_mem_reg[0][20] ;
  assign \new_[5649]_  = \\u8_mem_reg[0][20] ;
  assign \new_[5650]_  = \\u8_mem_reg[0][21] ;
  assign \new_[5651]_  = \\u3_mem_reg[0][22] ;
  assign \new_[5652]_  = \\u8_mem_reg[0][23] ;
  assign \new_[5653]_  = \\u8_mem_reg[0][24] ;
  assign \new_[5654]_  = \\u8_mem_reg[0][25] ;
  assign \new_[5655]_  = \\u3_mem_reg[0][24] ;
  assign \new_[5656]_  = \\u3_mem_reg[0][25] ;
  assign \new_[5657]_  = \\u3_mem_reg[0][26] ;
  assign \new_[5658]_  = \\u3_mem_reg[0][28] ;
  assign \new_[5659]_  = \\u8_mem_reg[0][7] ;
  assign \new_[5660]_  = \\u8_mem_reg[0][8] ;
  assign \new_[5661]_  = \\u8_mem_reg[0][6] ;
  assign \new_[5662]_  = \\u8_mem_reg[0][9] ;
  assign \new_[5663]_  = \\u3_mem_reg[0][30] ;
  assign \new_[5664]_  = \\u3_mem_reg[0][3] ;
  assign \new_[5665]_  = \\u3_mem_reg[0][8] ;
  assign \new_[5666]_  = \\u7_mem_reg[1][10] ;
  assign \new_[5667]_  = ~\\u13_crac_dout_r_reg[7] ;
  assign \new_[5668]_  = \\u6_mem_reg[2][22] ;
  assign \new_[5669]_  = \\u6_mem_reg[0][0] ;
  assign \new_[5670]_  = \\u6_mem_reg[3][4] ;
  assign \new_[5671]_  = \\u13_intm_r_reg[26] ;
  assign \new_[5672]_  = \\u6_mem_reg[3][2] ;
  assign \new_[5673]_  = \\u13_occ0_r_reg[22] ;
  assign \new_[5674]_  = \\u6_mem_reg[3][26] ;
  assign \new_[5675]_  = \\u6_mem_reg[3][22] ;
  assign \new_[5676]_  = \\u6_mem_reg[3][15] ;
  assign \new_[5677]_  = \\u5_mem_reg[0][6] ;
  assign \new_[5678]_  = \\u6_mem_reg[3][19] ;
  assign n4891 = \\u1_sr_reg[10] ;
  assign n4936 = ~\new_[6568]_  & ~\new_[12403]_ ;
  assign n4991 = ~\new_[6570]_  & ~\new_[12040]_ ;
  assign n4946 = ~\new_[6571]_  & ~\new_[11421]_ ;
  assign n4941 = ~\new_[6569]_  & ~\new_[12811]_ ;
  assign n4921 = ~\new_[6572]_  & ~\new_[12074]_ ;
  assign n4951 = ~\new_[6573]_  & ~\new_[13168]_ ;
  assign \new_[5686]_  = \\u5_mem_reg[0][30] ;
  assign \new_[5687]_  = \\u5_mem_reg[0][23] ;
  assign \new_[5688]_  = \\u13_crac_r_reg[2] ;
  assign \new_[5689]_  = \\u6_mem_reg[2][4] ;
  assign \new_[5690]_  = \\u6_mem_reg[3][11] ;
  assign \new_[5691]_  = \\u6_mem_reg[2][8] ;
  assign \new_[5692]_  = \\u6_mem_reg[2][2] ;
  assign \new_[5693]_  = \\u3_mem_reg[0][9] ;
  assign \new_[5694]_  = \\u13_occ0_r_reg[26] ;
  assign \new_[5695]_  = \\u5_mem_reg[0][28] ;
  assign \new_[5696]_  = \\u13_intm_r_reg[3] ;
  assign \new_[5697]_  = \\u6_mem_reg[2][26] ;
  assign n4956 = \new_[6565]_  | n9671;
  assign n4961 = \new_[6566]_  | n9646;
  assign n4911 = \new_[6567]_  | n9436;
  assign \new_[5701]_  = \\u3_mem_reg[0][4] ;
  assign \new_[5702]_  = \\u5_mem_reg[0][20] ;
  assign \new_[5703]_  = \\u8_mem_reg[0][31] ;
  assign \new_[5704]_  = \\u6_mem_reg[2][15] ;
  assign \new_[5705]_  = \\u6_mem_reg[1][15] ;
  assign n4966 = ~\new_[6836]_  | ~\new_[6422]_ ;
  assign n4976 = ~\new_[6838]_  | ~\new_[6423]_ ;
  assign \new_[5708]_  = \\u6_mem_reg[2][19] ;
  assign n4916 = ~\new_[6839]_  | ~\new_[6424]_ ;
  assign n4971 = ~\new_[6837]_  | ~\new_[6425]_ ;
  assign n4981 = ~\new_[6840]_  | ~\new_[6426]_ ;
  assign n4986 = ~\new_[6841]_  | ~\new_[6427]_ ;
  assign \new_[5713]_  = ~\new_[6564]_  & (~\new_[8549]_  | ~\new_[9782]_ );
  assign \new_[5714]_  = \\u6_mem_reg[2][11] ;
  assign \new_[5715]_  = \\u5_mem_reg[0][17] ;
  assign \new_[5716]_  = \\u13_occ0_r_reg[19] ;
  assign \new_[5717]_  = \\u5_mem_reg[0][12] ;
  assign \new_[5718]_  = \\u6_mem_reg[1][26] ;
  assign \new_[5719]_  = \\u4_mem_reg[0][6] ;
  assign \new_[5720]_  = \\u6_mem_reg[1][4] ;
  assign \new_[5721]_  = \\u6_mem_reg[1][8] ;
  assign \new_[5722]_  = \\u6_mem_reg[1][2] ;
  assign \new_[5723]_  = \\u5_mem_reg[0][0] ;
  assign \new_[5724]_  = \\u6_mem_reg[1][22] ;
  assign \new_[5725]_  = \\u8_mem_reg[0][3] ;
  assign \new_[5726]_  = \\u4_mem_reg[0][30] ;
  assign \new_[5727]_  = \\u8_mem_reg[0][16] ;
  assign \new_[5728]_  = \\u5_mem_reg[3][8] ;
  assign \new_[5729]_  = \\u6_mem_reg[1][11] ;
  assign \new_[5730]_  = \\u5_mem_reg[3][4] ;
  assign \new_[5731]_  = \\u8_mem_reg[0][2] ;
  assign \new_[5732]_  = \\u5_mem_reg[2][8] ;
  assign \new_[5733]_  = \\u4_mem_reg[0][23] ;
  assign \new_[5734]_  = \\u3_mem_reg[0][23] ;
  assign \new_[5735]_  = \\u4_mem_reg[0][17] ;
  assign \new_[5736]_  = \\u5_mem_reg[3][19] ;
  assign \new_[5737]_  = \\u5_mem_reg[3][26] ;
  assign \new_[5738]_  = \\u5_mem_reg[3][2] ;
  assign \new_[5739]_  = ~\new_[12848]_  | ~\new_[7451]_  | ~n10961 | ~\new_[12070]_ ;
  assign \new_[5740]_  = \\u5_mem_reg[3][22] ;
  assign \new_[5741]_  = ~\new_[12709]_  | ~\new_[7552]_  | ~n10966 | ~\new_[11413]_ ;
  assign \new_[5742]_  = ~\new_[12735]_  | ~\new_[7561]_  | ~n11056 | ~\new_[11414]_ ;
  assign \new_[5743]_  = \\u5_mem_reg[3][15] ;
  assign \new_[5744]_  = \\u8_mem_reg[0][27] ;
  assign \new_[5745]_  = ~\new_[12484]_  | ~\new_[7528]_  | ~n10956 | ~\new_[12097]_ ;
  assign \new_[5746]_  = ~\new_[12345]_  | ~\new_[7575]_  | ~n10971 | ~\new_[12006]_ ;
  assign \new_[5747]_  = ~\new_[12344]_  | ~\new_[7588]_  | ~n11061 | ~\new_[11999]_ ;
  assign \new_[5748]_  = \\u4_mem_reg[0][20] ;
  assign \new_[5749]_  = ~\new_[5887]_ ;
  assign \new_[5750]_  = ~\new_[7465]_  & ~\new_[6421]_ ;
  assign \new_[5751]_  = \\u5_mem_reg[3][11] ;
  assign \new_[5752]_  = \\u5_mem_reg[2][2] ;
  assign \new_[5753]_  = \\u4_mem_reg[0][12] ;
  assign \new_[5754]_  = \\u5_mem_reg[2][26] ;
  assign \new_[5755]_  = \\u8_mem_reg[0][22] ;
  assign \new_[5756]_  = \\u13_occ0_r_reg[15] ;
  assign \new_[5757]_  = \\u5_mem_reg[1][2] ;
  assign \new_[5758]_  = \\u5_mem_reg[2][11] ;
  assign \new_[5759]_  = \\u3_mem_reg[1][26] ;
  assign \new_[5760]_  = \\u5_mem_reg[2][19] ;
  assign \new_[5761]_  = \\u5_mem_reg[2][22] ;
  assign \new_[5762]_  = \\u5_mem_reg[2][15] ;
  assign \new_[5763]_  = \\u8_mem_reg[2][3] ;
  assign \new_[5764]_  = \\u5_mem_reg[1][8] ;
  assign \new_[5765]_  = \\u5_mem_reg[1][4] ;
  assign \new_[5766]_  = \\u8_mem_reg[0][1] ;
  assign \new_[5767]_  = \\u13_occ1_r_reg[11] ;
  assign \new_[5768]_  = (~\new_[7437]_  | ~\new_[13018]_ ) & (~\new_[13057]_  | ~\new_[12638]_ );
  assign \new_[5769]_  = ~\new_[6812]_  & (~\new_[12766]_  | ~\new_[7513]_ );
  assign n5226 = \new_[4858]_  ? \new_[7451]_  : \new_[10540]_ ;
  assign n5026 = \new_[4818]_  ? \new_[7552]_  : \new_[10549]_ ;
  assign n5031 = \new_[4819]_  ? \new_[7552]_  : \new_[10550]_ ;
  assign n5036 = \new_[4820]_  ? \new_[7552]_  : \new_[10553]_ ;
  assign n5041 = \new_[4821]_  ? \new_[7552]_  : \new_[10558]_ ;
  assign n5046 = \new_[4822]_  ? \new_[7552]_  : \new_[10562]_ ;
  assign n5051 = \new_[4823]_  ? \new_[7552]_  : \new_[10565]_ ;
  assign \new_[5777]_  = \\u3_mem_reg[0][0] ;
  assign n5056 = \new_[4824]_  ? \new_[7552]_  : \new_[10573]_ ;
  assign n5061 = \new_[4825]_  ? \new_[7552]_  : \new_[10575]_ ;
  assign n5066 = \new_[4826]_  ? \new_[7552]_  : \new_[10577]_ ;
  assign n5071 = \new_[4827]_  ? \new_[7552]_  : \new_[10579]_ ;
  assign n5076 = \new_[4828]_  ? \new_[7561]_  : \new_[10659]_ ;
  assign n5081 = \new_[4829]_  ? \new_[7561]_  : \new_[10589]_ ;
  assign n5086 = \new_[4830]_  ? \new_[7561]_  : \new_[10591]_ ;
  assign n5091 = \new_[4831]_  ? \new_[7561]_  : \new_[10594]_ ;
  assign n5096 = \new_[4832]_  ? \new_[7561]_  : \new_[10598]_ ;
  assign n5101 = \new_[4833]_  ? \new_[7561]_  : \new_[10600]_ ;
  assign n5106 = \new_[4834]_  ? \new_[7561]_  : \new_[10609]_ ;
  assign n5111 = \new_[4835]_  ? \new_[7561]_  : \new_[10611]_ ;
  assign n5116 = \new_[4836]_  ? \new_[7561]_  : \new_[10612]_ ;
  assign n5121 = \new_[4837]_  ? \new_[7561]_  : \new_[10614]_ ;
  assign n5306 = \new_[4874]_  ? \new_[7451]_  : \new_[10533]_ ;
  assign n5126 = \new_[4838]_  ? \new_[7528]_  : \new_[10622]_ ;
  assign n5131 = \new_[4839]_  ? \new_[7528]_  : \new_[10709]_ ;
  assign n5136 = \new_[4840]_  ? \new_[7528]_  : \new_[10625]_ ;
  assign n5141 = \new_[4841]_  ? \new_[7528]_  : \new_[10703]_ ;
  assign n5146 = \new_[4842]_  ? \new_[7528]_  : \new_[10670]_ ;
  assign n5151 = \new_[4843]_  ? \new_[7528]_  : \new_[10667]_ ;
  assign n5156 = \new_[4844]_  ? \new_[7528]_  : \new_[10632]_ ;
  assign n5161 = \new_[4845]_  ? \new_[7528]_  : \new_[10642]_ ;
  assign n5166 = \new_[4846]_  ? \new_[7528]_  : \new_[10634]_ ;
  assign n5171 = \new_[4847]_  ? \new_[7528]_  : \new_[10636]_ ;
  assign n5176 = \new_[4848]_  ? \new_[7575]_  : \new_[10643]_ ;
  assign n5181 = \new_[4849]_  ? \new_[7575]_  : \new_[10618]_ ;
  assign n5186 = \new_[4850]_  ? \new_[7575]_  : \new_[10552]_ ;
  assign n5191 = \new_[4851]_  ? \new_[7575]_  : \new_[11424]_ ;
  assign n5196 = \new_[4852]_  ? \new_[7575]_  : \new_[10647]_ ;
  assign n5201 = \new_[4853]_  ? \new_[7575]_  : \new_[10648]_ ;
  assign n5206 = \new_[4854]_  ? \new_[7575]_  : \new_[10651]_ ;
  assign n5211 = \new_[4855]_  ? \new_[7575]_  : \new_[10663]_ ;
  assign n5216 = \new_[4856]_  ? \new_[7575]_  : \new_[10660]_ ;
  assign n5221 = \new_[4857]_  ? \new_[7575]_  : \new_[10657]_ ;
  assign n5231 = \new_[4859]_  ? \new_[7451]_  : \new_[10539]_ ;
  assign n5236 = \new_[4860]_  ? \new_[7451]_  : \new_[10544]_ ;
  assign n5241 = \new_[4861]_  ? \new_[7588]_  : \new_[10676]_ ;
  assign n5246 = \new_[4862]_  ? \new_[7588]_  : \new_[10537]_ ;
  assign n5251 = \new_[4863]_  ? \new_[7588]_  : \new_[10535]_ ;
  assign n5261 = \new_[4865]_  ? \new_[7451]_  : \new_[10682]_ ;
  assign n5256 = \new_[4864]_  ? \new_[7588]_  : \new_[10529]_ ;
  assign n5266 = \new_[4866]_  ? \new_[7451]_  : \new_[10685]_ ;
  assign n5271 = \new_[4867]_  ? \new_[7588]_  : \new_[10689]_ ;
  assign n5276 = \new_[4868]_  ? \new_[7588]_  : \new_[10617]_ ;
  assign n5281 = \new_[4869]_  ? \new_[7588]_  : \new_[10691]_ ;
  assign n5286 = \new_[4870]_  ? \new_[7588]_  : \new_[10582]_ ;
  assign n5291 = \new_[4871]_  ? \new_[7451]_  : \new_[10693]_ ;
  assign n5296 = \new_[4872]_  ? \new_[7588]_  : \new_[10520]_ ;
  assign n5301 = \new_[4873]_  ? \new_[7588]_  : \new_[10695]_ ;
  assign n5311 = \new_[4875]_  ? \new_[7451]_  : \new_[10696]_ ;
  assign n5321 = \new_[4877]_  ? \new_[7451]_  : \new_[10564]_ ;
  assign n5316 = \new_[4876]_  ? \new_[7451]_  : \new_[10702]_ ;
  assign \new_[5831]_  = ~\new_[6760]_  & (~\new_[4689]_  | ~\new_[7616]_ );
  assign \new_[5832]_  = ~\new_[6777]_  & (~\new_[13124]_  | ~\new_[7610]_ );
  assign \new_[5833]_  = ~\new_[6778]_  & (~\new_[13083]_  | ~\new_[7612]_ );
  assign \new_[5834]_  = ~\new_[6765]_  & (~\new_[13161]_  | ~\new_[7609]_ );
  assign \new_[5835]_  = ~\new_[6779]_  & (~\new_[13158]_  | ~\new_[7605]_ );
  assign \new_[5836]_  = ~\new_[6780]_  & (~\new_[13092]_  | ~\new_[7614]_ );
  assign \new_[5837]_  = u14_u8_en_out_l2_reg;
  assign \wb_data_o[4]  = \\u12_wb_data_o_reg[4] ;
  assign \wb_data_o[6]  = \\u12_wb_data_o_reg[6] ;
  assign \wb_data_o[10]  = \\u12_wb_data_o_reg[10] ;
  assign \new_[5841]_  = \\u13_occ1_r_reg[8] ;
  assign \new_[5842]_  = \\u13_occ1_r_reg[0] ;
  assign \new_[5843]_  = \\u13_occ1_r_reg[10] ;
  assign \new_[5844]_  = \\u13_occ1_r_reg[12] ;
  assign \new_[5845]_  = \\u13_occ1_r_reg[13] ;
  assign \new_[5846]_  = \\u13_occ1_r_reg[14] ;
  assign \new_[5847]_  = \\u13_occ1_r_reg[1] ;
  assign \new_[5848]_  = \\u13_occ1_r_reg[2] ;
  assign \new_[5849]_  = \\u13_occ1_r_reg[3] ;
  assign \new_[5850]_  = \\u13_occ1_r_reg[5] ;
  assign \new_[5851]_  = \\u13_occ1_r_reg[6] ;
  assign \new_[5852]_  = \\u13_occ1_r_reg[7] ;
  assign \new_[5853]_  = \\u1_slt1_reg[7] ;
  assign \new_[5854]_  = \\u1_slt2_reg[7] ;
  assign \new_[5855]_  = \\u1_slt4_reg[7] ;
  assign \new_[5856]_  = \\u1_slt3_reg[7] ;
  assign \new_[5857]_  = \\u3_mem_reg[0][14] ;
  assign \new_[5858]_  = \\u3_mem_reg[0][7] ;
  assign \new_[5859]_  = u14_u6_full_empty_r_reg;
  assign \new_[5860]_  = u14_u8_full_empty_r_reg;
  assign \wb_data_o[0]  = \\u12_wb_data_o_reg[0] ;
  assign \wb_data_o[14]  = \\u12_wb_data_o_reg[14] ;
  assign \wb_data_o[13]  = \\u12_wb_data_o_reg[13] ;
  assign \wb_data_o[12]  = \\u12_wb_data_o_reg[12] ;
  assign \wb_data_o[11]  = \\u12_wb_data_o_reg[11] ;
  assign \wb_data_o[9]  = \\u12_wb_data_o_reg[9] ;
  assign \wb_data_o[7]  = \\u12_wb_data_o_reg[7] ;
  assign \wb_data_o[15]  = \\u12_wb_data_o_reg[15] ;
  assign \wb_data_o[5]  = \\u12_wb_data_o_reg[5] ;
  assign \wb_data_o[3]  = \\u12_wb_data_o_reg[3] ;
  assign \wb_data_o[8]  = \\u12_wb_data_o_reg[8] ;
  assign \wb_data_o[2]  = \\u12_wb_data_o_reg[2] ;
  assign \new_[5873]_  = \\u13_occ1_r_reg[9] ;
  assign \new_[5874]_  = \\u13_occ1_r_reg[15] ;
  assign \new_[5875]_  = \\u3_mem_reg[0][31] ;
  assign \new_[5876]_  = \\u13_occ1_r_reg[4] ;
  assign \new_[5877]_  = ~\new_[13077]_  & ~\new_[6830]_ ;
  assign \new_[5878]_  = ~\new_[14185]_  & ~\new_[6832]_ ;
  assign \new_[5879]_  = ~\new_[6830]_  & ~\new_[13518]_ ;
  assign \new_[5880]_  = ~\new_[6832]_  & ~\new_[13223]_ ;
  assign n5011 = n9666 ? \new_[8805]_  : \new_[4815]_ ;
  assign n5006 = n9666 ? \new_[8996]_  : \new_[4814]_ ;
  assign n5021 = n9666 ? \new_[9002]_  : \new_[4817]_ ;
  assign n5016 = n9666 ? \new_[9000]_  : \new_[4816]_ ;
  assign n5001 = n9666 ? \new_[9001]_  : \new_[4813]_ ;
  assign \new_[5886]_  = \\u0_slt9_r_reg[1] ;
  assign \new_[5887]_  = n9671 & \new_[6759]_ ;
  assign \new_[5888]_  = \\u1_slt6_reg[7] ;
  assign n7091 = ~\new_[7018]_  | (~\new_[9407]_  & ~\new_[7549]_ );
  assign n5466 = ~\new_[7020]_  | (~\new_[9409]_  & ~\new_[7549]_ );
  assign n7096 = ~\new_[7021]_  | (~\new_[9410]_  & ~\new_[7547]_ );
  assign n7101 = ~\new_[7022]_  | (~\new_[9411]_  & ~\new_[7547]_ );
  assign n7106 = ~\new_[7023]_  | (~\new_[9413]_  & ~\new_[7547]_ );
  assign n7111 = ~\new_[7024]_  | (~\new_[9414]_  & ~\new_[7547]_ );
  assign n7116 = ~\new_[7025]_  | (~\new_[9415]_  & ~\new_[7553]_ );
  assign n7121 = ~\new_[7026]_  | (~\new_[9416]_  & ~\new_[7553]_ );
  assign n7126 = ~\new_[7027]_  | (~\new_[9417]_  & ~\new_[7553]_ );
  assign n5426 = ~\new_[7028]_  | (~\new_[9418]_  & ~\new_[7553]_ );
  assign n7131 = ~\new_[7029]_  | (~\new_[9419]_  & ~\new_[7548]_ );
  assign n7136 = ~\new_[7030]_  | (~\new_[9420]_  & ~\new_[7548]_ );
  assign n7141 = ~\new_[7031]_  | (~\new_[9421]_  & ~\new_[7546]_ );
  assign n5431 = ~\new_[7032]_  | (~\new_[9423]_  & ~\new_[7546]_ );
  assign n7146 = ~\new_[7033]_  | (~\new_[9424]_  & ~\new_[7546]_ );
  assign n7151 = ~\new_[7034]_  | (~\new_[9425]_  & ~\new_[7546]_ );
  assign n7156 = ~\new_[7035]_  | (~\new_[9427]_  & ~\new_[7548]_ );
  assign n5411 = ~\new_[7036]_  | (~\new_[9428]_  & ~\new_[7548]_ );
  assign n7161 = ~\new_[7037]_  | (~\new_[9430]_  & ~\new_[7550]_ );
  assign n7166 = ~\new_[7039]_  | (~\new_[9431]_  & ~\new_[7550]_ );
  assign n7171 = ~\new_[7040]_  | (~\new_[9433]_  & ~\new_[7549]_ );
  assign n5406 = ~\new_[7041]_  | (~\new_[9434]_  & ~\new_[7549]_ );
  assign n7176 = ~\new_[7042]_  | (~\new_[9436]_  & ~\new_[7550]_ );
  assign n7181 = ~\new_[7043]_  | (~\new_[9437]_  & ~\new_[7550]_ );
  assign n7186 = ~\new_[7044]_  | (~\new_[9439]_  & ~\new_[7549]_ );
  assign n5401 = ~\new_[7045]_  | (~\new_[9440]_  & ~\new_[7549]_ );
  assign n6586 = ~\new_[6877]_  | (~\new_[10045]_  & ~\new_[7542]_ );
  assign n7196 = ~\new_[7051]_  | (~\new_[9454]_  & ~\new_[7564]_ );
  assign n7201 = ~\new_[7052]_  | (~\new_[9455]_  & ~\new_[7564]_ );
  assign n5386 = ~\new_[7053]_  | (~\new_[9456]_  & ~\new_[7559]_ );
  assign n7206 = ~\new_[7054]_  | (~\new_[9478]_  & ~\new_[7559]_ );
  assign n7211 = ~\new_[7055]_  | (~\new_[9459]_  & ~\new_[7559]_ );
  assign n7216 = ~\new_[7056]_  | (~\new_[9460]_  & ~\new_[7564]_ );
  assign n5376 = ~\new_[7057]_  | (~\new_[9462]_  & ~\new_[7564]_ );
  assign n7226 = ~\new_[7058]_  | (~\new_[9463]_  & ~\new_[7559]_ );
  assign n7231 = ~\new_[7059]_  | (~\new_[9464]_  & ~\new_[7559]_ );
  assign n7236 = ~\new_[7060]_  | (~\new_[9466]_  & ~\new_[7559]_ );
  assign n5381 = ~\new_[7061]_  | (~\new_[9467]_  & ~\new_[7559]_ );
  assign n7241 = ~\new_[7062]_  | (~\new_[9468]_  & ~\new_[7564]_ );
  assign n7246 = ~\new_[7063]_  | (~\new_[9469]_  & ~\new_[7554]_ );
  assign n7251 = ~\new_[7064]_  | (~\new_[9470]_  & ~\new_[7563]_ );
  assign n5371 = ~\new_[7065]_  | (~\new_[9471]_  & ~\new_[7564]_ );
  assign n7256 = ~\new_[7066]_  | (~\new_[9472]_  & ~\new_[7560]_ );
  assign n7261 = ~\new_[7067]_  | (~\new_[9473]_  & ~\new_[7560]_ );
  assign n7266 = ~\new_[7068]_  | (~\new_[9474]_  & ~\new_[7562]_ );
  assign n5361 = ~\new_[7069]_  | (~\new_[9475]_  & ~\new_[7563]_ );
  assign n7271 = ~\new_[7070]_  | (~\new_[9476]_  & ~\new_[7560]_ );
  assign n7276 = ~\new_[7071]_  | (~\new_[9477]_  & ~\new_[7562]_ );
  assign n7281 = ~\new_[7072]_  | (~\new_[9479]_  & ~\new_[7560]_ );
  assign n9376 = ~\new_[7073]_  | (~\new_[9480]_  & ~\new_[7564]_ );
  assign n7286 = ~\new_[7074]_  | (~\new_[9482]_  & ~\new_[7554]_ );
  assign n7291 = ~\new_[7075]_  | (~\new_[9483]_  & ~\new_[7559]_ );
  assign n7296 = ~\new_[7076]_  | (~\new_[9484]_  & ~\new_[7556]_ );
  assign n9416 = ~\new_[7077]_  | (~\new_[9485]_  & ~\new_[7564]_ );
  assign n7301 = ~\new_[7078]_  | (~\new_[9486]_  & ~\new_[7564]_ );
  assign n7306 = ~\new_[7079]_  | (~\new_[9487]_  & ~\new_[7555]_ );
  assign n7311 = ~\new_[7080]_  | (~\new_[9488]_  & ~\new_[7559]_ );
  assign n9411 = ~\new_[7081]_  | (~\new_[9371]_  & ~\new_[7564]_ );
  assign n7316 = ~\new_[7082]_  | (~\new_[9490]_  & ~\new_[7564]_ );
  assign n7321 = ~\new_[7084]_  | (~\new_[10050]_  & ~\new_[7564]_ );
  assign n7326 = ~\new_[7085]_  | (~\new_[10051]_  & ~\new_[7560]_ );
  assign n9381 = ~\new_[7086]_  | (~\new_[10052]_  & ~\new_[7559]_ );
  assign n7331 = ~\new_[7087]_  | (~\new_[10053]_  & ~\new_[7559]_ );
  assign n7336 = ~\new_[7088]_  | (~\new_[9900]_  & ~\new_[7560]_ );
  assign n7341 = ~\new_[7089]_  | (~\new_[10054]_  & ~\new_[7559]_ );
  assign n9401 = ~\new_[7090]_  | (~\new_[10055]_  & ~\new_[7562]_ );
  assign n7346 = ~\new_[7091]_  | (~\new_[10056]_  & ~\new_[7559]_ );
  assign n7351 = ~\new_[7092]_  | (~\new_[10057]_  & ~\new_[7563]_ );
  assign n7356 = ~\new_[7093]_  | (~\new_[10058]_  & ~\new_[7559]_ );
  assign n9391 = ~\new_[7094]_  | (~\new_[10151]_  & ~\new_[7560]_ );
  assign n7361 = ~\new_[7095]_  | (~\new_[10059]_  & ~\new_[7555]_ );
  assign n7366 = ~\new_[7096]_  | (~\new_[10060]_  & ~\new_[7562]_ );
  assign n7371 = ~\new_[7097]_  | (~\new_[10062]_  & ~\new_[7560]_ );
  assign n9396 = ~\new_[7098]_  | (~\new_[10063]_  & ~\new_[7559]_ );
  assign n7376 = ~\new_[7099]_  | (~\new_[10138]_  & ~\new_[7564]_ );
  assign n7381 = ~\new_[7100]_  | (~\new_[10064]_  & ~\new_[7563]_ );
  assign n7386 = ~\new_[7101]_  | (~\new_[10065]_  & ~\new_[7563]_ );
  assign n9361 = ~\new_[7102]_  | (~\new_[10066]_  & ~\new_[7554]_ );
  assign n7391 = ~\new_[7103]_  | (~\new_[10067]_  & ~\new_[7556]_ );
  assign n7396 = ~\new_[7104]_  | (~\new_[10068]_  & ~\new_[7555]_ );
  assign n7401 = ~\new_[7105]_  | (~\new_[10070]_  & ~\new_[7563]_ );
  assign n9351 = ~\new_[7106]_  | (~\new_[10127]_  & ~\new_[7564]_ );
  assign n7406 = ~\new_[7107]_  | (~\new_[10126]_  & ~\new_[7564]_ );
  assign n7411 = ~\new_[7108]_  | (~\new_[10071]_  & ~\new_[7554]_ );
  assign n7416 = ~\new_[7109]_  | (~\new_[10072]_  & ~\new_[7564]_ );
  assign n7421 = ~\new_[7110]_  | (~\new_[10121]_  & ~\new_[7555]_ );
  assign n7426 = ~\new_[7111]_  | (~\new_[10119]_  & ~\new_[7556]_ );
  assign n7431 = ~\new_[7112]_  | (~\new_[10073]_  & ~\new_[7556]_ );
  assign n7436 = ~\new_[7113]_  | (~\new_[10074]_  & ~\new_[7563]_ );
  assign n9291 = ~\new_[7114]_  | (~\new_[10075]_  & ~\new_[7563]_ );
  assign n7441 = ~\new_[7115]_  | (~\new_[10076]_  & ~\new_[7559]_ );
  assign n7446 = ~\new_[7116]_  | (~\new_[9498]_  & ~\new_[7554]_ );
  assign n7451 = ~\new_[7117]_  | (~\new_[9499]_  & ~\new_[7554]_ );
  assign n9346 = ~\new_[7118]_  | (~\new_[9500]_  & ~\new_[7554]_ );
  assign n7456 = ~\new_[7119]_  | (~\new_[9501]_  & ~\new_[7554]_ );
  assign n7461 = ~\new_[7120]_  | (~\new_[9502]_  & ~\new_[7557]_ );
  assign n7466 = ~\new_[7121]_  | (~\new_[9503]_  & ~\new_[7557]_ );
  assign n9331 = ~\new_[7122]_  | (~\new_[9504]_  & ~\new_[7557]_ );
  assign n7471 = ~\new_[7123]_  | (~\new_[9505]_  & ~\new_[7557]_ );
  assign n7476 = ~\new_[7124]_  | (~\new_[9506]_  & ~\new_[7558]_ );
  assign n7481 = ~\new_[7125]_  | (~\new_[9508]_  & ~\new_[7558]_ );
  assign n9311 = ~\new_[7126]_  | (~\new_[9509]_  & ~\new_[7558]_ );
  assign n7486 = ~\new_[7127]_  | (~\new_[9511]_  & ~\new_[7558]_ );
  assign n7491 = ~\new_[7128]_  | (~\new_[9512]_  & ~\new_[7562]_ );
  assign n7496 = ~\new_[7129]_  | (~\new_[9513]_  & ~\new_[7562]_ );
  assign n9326 = ~\new_[7130]_  | (~\new_[9514]_  & ~\new_[7562]_ );
  assign n7506 = ~\new_[7131]_  | (~\new_[9515]_  & ~\new_[7562]_ );
  assign n7511 = ~\new_[7132]_  | (~\new_[9516]_  & ~\new_[7557]_ );
  assign n7516 = ~\new_[7133]_  | (~\new_[9517]_  & ~\new_[7557]_ );
  assign n9316 = ~\new_[7134]_  | (~\new_[9518]_  & ~\new_[7555]_ );
  assign n7521 = ~\new_[7135]_  | (~\new_[9519]_  & ~\new_[7555]_ );
  assign n7526 = ~\new_[7136]_  | (~\new_[9520]_  & ~\new_[7555]_ );
  assign n7531 = ~\new_[7137]_  | (~\new_[9521]_  & ~\new_[7555]_ );
  assign n9321 = ~\new_[7138]_  | (~\new_[9522]_  & ~\new_[7557]_ );
  assign n7536 = ~\new_[7139]_  | (~\new_[9524]_  & ~\new_[7557]_ );
  assign n7541 = ~\new_[7140]_  | (~\new_[9526]_  & ~\new_[7558]_ );
  assign n7546 = ~\new_[7141]_  | (~\new_[9527]_  & ~\new_[7558]_ );
  assign n9281 = ~\new_[7142]_  | (~\new_[9528]_  & ~\new_[7556]_ );
  assign n7551 = ~\new_[7143]_  | (~\new_[9529]_  & ~\new_[7556]_ );
  assign n7556 = ~\new_[7144]_  | (~\new_[9547]_  & ~\new_[7558]_ );
  assign n7561 = ~\new_[7145]_  | (~\new_[9530]_  & ~\new_[7558]_ );
  assign n9271 = ~\new_[7146]_  | (~\new_[9532]_  & ~\new_[7556]_ );
  assign n7566 = ~\new_[7147]_  | (~\new_[9533]_  & ~\new_[7556]_ );
  assign n5741 = ~\new_[7150]_  | (~\new_[10501]_  & ~\new_[7584]_ );
  assign n5551 = ~\new_[7380]_  | (~\new_[10108]_  & ~\new_[7579]_ );
  assign n7191 = ~\new_[7152]_  | (~\new_[10081]_  & ~\new_[7542]_ );
  assign n6561 = ~\new_[7254]_  | (~\new_[10508]_  & ~\new_[7580]_ );
  assign n7571 = ~\new_[7155]_  | (~\new_[9549]_  & ~\new_[7531]_ );
  assign n7576 = ~\new_[7156]_  | (~\new_[9567]_  & ~\new_[7531]_ );
  assign n9276 = ~\new_[7157]_  | (~\new_[9550]_  & ~\new_[7527]_ );
  assign n7581 = ~\new_[7158]_  | (~\new_[9564]_  & ~\new_[7527]_ );
  assign n7586 = ~\new_[7159]_  | (~\new_[9551]_  & ~\new_[7527]_ );
  assign n7591 = ~\new_[7160]_  | (~\new_[9559]_  & ~\new_[7531]_ );
  assign n9191 = ~\new_[7161]_  | (~\new_[9556]_  & ~\new_[7531]_ );
  assign n7596 = ~\new_[7162]_  | (~\new_[9553]_  & ~\new_[7527]_ );
  assign n7601 = ~\new_[7163]_  | (~\new_[9552]_  & ~\new_[7527]_ );
  assign n7606 = ~\new_[7164]_  | (~\new_[9531]_  & ~\new_[7527]_ );
  assign n7611 = ~\new_[7165]_  | (~\new_[9525]_  & ~\new_[7527]_ );
  assign n7616 = ~\new_[7167]_  | (~\new_[9554]_  & ~\new_[7531]_ );
  assign n7621 = ~\new_[7168]_  | (~\new_[9555]_  & ~\new_[7520]_ );
  assign n7626 = ~\new_[7169]_  | (~\new_[9497]_  & ~\new_[7530]_ );
  assign n9251 = ~\new_[7170]_  | (~\new_[9496]_  & ~\new_[7531]_ );
  assign n7631 = ~\new_[7171]_  | (~\new_[9493]_  & ~\new_[7526]_ );
  assign n7636 = ~\new_[7172]_  | (~\new_[9557]_  & ~\new_[7526]_ );
  assign n7641 = ~\new_[7173]_  | (~\new_[9492]_  & ~\new_[7529]_ );
  assign n9221 = ~\new_[7174]_  | (~\new_[9489]_  & ~\new_[7530]_ );
  assign n7646 = ~\new_[7175]_  | (~\new_[9481]_  & ~\new_[7521]_ );
  assign n7651 = ~\new_[7176]_  | (~\new_[9558]_  & ~\new_[7529]_ );
  assign n7656 = ~\new_[7178]_  | (~\new_[9449]_  & ~\new_[7521]_ );
  assign n9241 = ~\new_[7179]_  | (~\new_[9560]_  & ~\new_[7531]_ );
  assign n7661 = ~\new_[7180]_  | (~\new_[9372]_  & ~\new_[7520]_ );
  assign n7666 = ~\new_[7181]_  | (~\new_[9561]_  & ~\new_[7527]_ );
  assign n7671 = ~\new_[7182]_  | (~\new_[9562]_  & ~\new_[7523]_ );
  assign n9231 = ~\new_[7183]_  | (~\new_[9408]_  & ~\new_[7531]_ );
  assign n7676 = ~\new_[7184]_  | (~\new_[9400]_  & ~\new_[7531]_ );
  assign n7681 = ~\new_[7185]_  | (~\new_[9563]_  & ~\new_[7526]_ );
  assign n7686 = ~\new_[7186]_  | (~\new_[9396]_  & ~\new_[7527]_ );
  assign n9236 = ~\new_[7187]_  | (~\new_[9397]_  & ~\new_[7531]_ );
  assign n7691 = ~\new_[7188]_  | (~\new_[9591]_  & ~\new_[7531]_ );
  assign n7696 = ~\new_[7189]_  | (~\new_[9989]_  & ~\new_[7531]_ );
  assign n7701 = ~\new_[7190]_  | (~\new_[10089]_  & ~\new_[7526]_ );
  assign n9201 = ~\new_[7192]_  | (~\new_[9964]_  & ~\new_[7527]_ );
  assign n7706 = ~\new_[7193]_  | (~\new_[9957]_  & ~\new_[7527]_ );
  assign n7711 = ~\new_[7194]_  | (~\new_[9945]_  & ~\new_[7526]_ );
  assign n7716 = ~\new_[7195]_  | (~\new_[10090]_  & ~\new_[7527]_ );
  assign n9186 = ~\new_[7196]_  | (~\new_[9936]_  & ~\new_[7529]_ );
  assign n7721 = ~\new_[7197]_  | (~\new_[10091]_  & ~\new_[7527]_ );
  assign n7726 = ~\new_[7198]_  | (~\new_[9932]_  & ~\new_[7530]_ );
  assign n7731 = ~\new_[7199]_  | (~\new_[9924]_  & ~\new_[7527]_ );
  assign n9196 = ~\new_[7200]_  | (~\new_[9917]_  & ~\new_[7521]_ );
  assign n7736 = ~\new_[7201]_  | (~\new_[10092]_  & ~\new_[7526]_ );
  assign n7741 = ~\new_[7202]_  | (~\new_[9915]_  & ~\new_[7529]_ );
  assign n7746 = ~\new_[7203]_  | (~\new_[9909]_  & ~\new_[7521]_ );
  assign n9051 = ~\new_[7204]_  | (~\new_[9906]_  & ~\new_[7527]_ );
  assign n7751 = ~\new_[7205]_  | (~\new_[10093]_  & ~\new_[7531]_ );
  assign n7756 = ~\new_[7206]_  | (~\new_[9902]_  & ~\new_[7530]_ );
  assign n7761 = ~\new_[7207]_  | (~\new_[10095]_  & ~\new_[7530]_ );
  assign n9166 = ~\new_[7208]_  | (~\new_[9899]_  & ~\new_[7520]_ );
  assign n7766 = ~\new_[7209]_  | (~\new_[9898]_  & ~\new_[7523]_ );
  assign n7771 = ~\new_[7210]_  | (~\new_[9896]_  & ~\new_[7526]_ );
  assign n7776 = ~\new_[7211]_  | (~\new_[10069]_  & ~\new_[7530]_ );
  assign n9141 = ~\new_[7212]_  | (~\new_[10104]_  & ~\new_[7531]_ );
  assign n7781 = ~\new_[7213]_  | (~\new_[10031]_  & ~\new_[7531]_ );
  assign n7786 = ~\new_[7214]_  | (~\new_[10032]_  & ~\new_[7520]_ );
  assign n7791 = ~\new_[7215]_  | (~\new_[10097]_  & ~\new_[7531]_ );
  assign n9126 = ~\new_[7216]_  | (~\new_[9975]_  & ~\new_[7526]_ );
  assign n7796 = ~\new_[7217]_  | (~\new_[10029]_  & ~\new_[7523]_ );
  assign n7801 = ~\new_[7218]_  | (~\new_[10027]_  & ~\new_[7523]_ );
  assign n7806 = ~\new_[7219]_  | (~\new_[10025]_  & ~\new_[7530]_ );
  assign n9136 = ~\new_[7220]_  | (~\new_[10015]_  & ~\new_[7530]_ );
  assign n7811 = ~\new_[7221]_  | (~\new_[10105]_  & ~\new_[7527]_ );
  assign n7816 = ~\new_[7222]_  | (~\new_[9569]_  & ~\new_[7520]_ );
  assign n7821 = ~\new_[7223]_  | (~\new_[9570]_  & ~\new_[7520]_ );
  assign n9131 = ~\new_[7224]_  | (~\new_[9571]_  & ~\new_[7520]_ );
  assign n7826 = ~\new_[7225]_  | (~\new_[9510]_  & ~\new_[7520]_ );
  assign n7831 = ~\new_[7226]_  | (~\new_[9572]_  & ~\new_[7524]_ );
  assign n7836 = ~\new_[7227]_  | (~\new_[9573]_  & ~\new_[7524]_ );
  assign n9091 = ~\new_[7228]_  | (~\new_[9574]_  & ~\new_[7524]_ );
  assign n7841 = ~\new_[7229]_  | (~\new_[9465]_  & ~\new_[7524]_ );
  assign n7846 = ~\new_[7230]_  | (~\new_[9461]_  & ~\new_[7522]_ );
  assign n7851 = ~\new_[7231]_  | (~\new_[9458]_  & ~\new_[7522]_ );
  assign n9101 = ~\new_[7232]_  | (~\new_[9575]_  & ~\new_[7522]_ );
  assign n7856 = ~\new_[7233]_  | (~\new_[9453]_  & ~\new_[7522]_ );
  assign n7861 = ~\new_[7234]_  | (~\new_[9452]_  & ~\new_[7529]_ );
  assign n7866 = ~\new_[7235]_  | (~\new_[9576]_  & ~\new_[7529]_ );
  assign n9086 = ~\new_[7236]_  | (~\new_[9451]_  & ~\new_[7529]_ );
  assign n7871 = ~\new_[7237]_  | (~\new_[9450]_  & ~\new_[7529]_ );
  assign n7876 = ~\new_[7238]_  | (~\new_[9448]_  & ~\new_[7524]_ );
  assign n7881 = ~\new_[7239]_  | (~\new_[9447]_  & ~\new_[7524]_ );
  assign n9081 = ~\new_[7240]_  | (~\new_[9577]_  & ~\new_[7521]_ );
  assign n7886 = ~\new_[7241]_  | (~\new_[9444]_  & ~\new_[7521]_ );
  assign n7891 = ~\new_[7242]_  | (~\new_[9494]_  & ~\new_[7521]_ );
  assign n7896 = ~\new_[7243]_  | (~\new_[9443]_  & ~\new_[7521]_ );
  assign n9071 = ~\new_[7244]_  | (~\new_[9578]_  & ~\new_[7524]_ );
  assign n7901 = ~\new_[7245]_  | (~\new_[9442]_  & ~\new_[7524]_ );
  assign n7906 = ~\new_[7246]_  | (~\new_[9441]_  & ~\new_[7525]_ );
  assign n7911 = ~\new_[7247]_  | (~\new_[9399]_  & ~\new_[7525]_ );
  assign n9061 = ~\new_[7248]_  | (~\new_[9580]_  & ~\new_[7523]_ );
  assign n7916 = ~\new_[7249]_  | (~\new_[9405]_  & ~\new_[7523]_ );
  assign n7921 = ~\new_[7250]_  | (~\new_[9581]_  & ~\new_[7525]_ );
  assign n7926 = ~\new_[7251]_  | (~\new_[9582]_  & ~\new_[7525]_ );
  assign n5886 = ~\new_[7252]_  | (~\new_[9583]_  & ~\new_[7523]_ );
  assign n7931 = ~\new_[7253]_  | (~\new_[9445]_  & ~\new_[7523]_ );
  assign n5436 = ~\new_[7388]_  | (~\new_[10087]_  & ~\new_[7587]_ );
  assign n6641 = ~\new_[6886]_  | (~\new_[10084]_  & ~\new_[7545]_ );
  assign n6571 = ~\new_[6875]_  | (~\new_[10506]_  & ~\new_[7583]_ );
  assign n5586 = ~\new_[6926]_  | (~\new_[9394]_  & ~\new_[7540]_ );
  assign n5736 = ~\new_[6879]_  | (~\new_[10502]_  & ~\new_[7585]_ );
  assign n8436 = ~\new_[7387]_  | (~\new_[9630]_  & ~\new_[7544]_ );
  assign n7941 = ~\new_[7259]_  | (~\new_[9595]_  & ~\new_[7578]_ );
  assign n9041 = ~\new_[7260]_  | (~\new_[9592]_  & ~\new_[7578]_ );
  assign n7946 = ~\new_[7261]_  | (~\new_[9579]_  & ~\new_[7573]_ );
  assign n8556 = ~\new_[7408]_  | (~\new_[9639]_  & ~\new_[7542]_ );
  assign n7951 = ~\new_[7262]_  | (~\new_[9593]_  & ~\new_[7573]_ );
  assign n7956 = ~\new_[7263]_  | (~\new_[9568]_  & ~\new_[7573]_ );
  assign n7221 = ~\new_[7264]_  | (~\new_[9594]_  & ~\new_[7578]_ );
  assign n7961 = ~\new_[7265]_  | (~\new_[9398]_  & ~\new_[7578]_ );
  assign n7966 = ~\new_[7266]_  | (~\new_[9596]_  & ~\new_[7573]_ );
  assign n7971 = ~\new_[7267]_  | (~\new_[9597]_  & ~\new_[7573]_ );
  assign n7976 = ~\new_[7268]_  | (~\new_[9382]_  & ~\new_[7573]_ );
  assign n7981 = ~\new_[7269]_  | (~\new_[9565]_  & ~\new_[7573]_ );
  assign n7986 = ~\new_[7270]_  | (~\new_[9422]_  & ~\new_[7578]_ );
  assign n7991 = ~\new_[7271]_  | (~\new_[9507]_  & ~\new_[7565]_ );
  assign n8776 = ~\new_[7272]_  | (~\new_[9598]_  & ~\new_[7577]_ );
  assign n7996 = ~\new_[7273]_  | (~\new_[9534]_  & ~\new_[7578]_ );
  assign n8001 = ~\new_[7274]_  | (~\new_[9600]_  & ~\new_[7572]_ );
  assign n8006 = ~\new_[7275]_  | (~\new_[9523]_  & ~\new_[7572]_ );
  assign n5581 = ~\new_[7276]_  | (~\new_[9601]_  & ~\new_[7576]_ );
  assign n8011 = ~\new_[7278]_  | (~\new_[9586]_  & ~\new_[7577]_ );
  assign n8016 = ~\new_[7279]_  | (~\new_[9602]_  & ~\new_[7574]_ );
  assign n8021 = ~\new_[7281]_  | (~\new_[9495]_  & ~\new_[7576]_ );
  assign n5941 = ~\new_[7282]_  | (~\new_[9603]_  & ~\new_[7574]_ );
  assign n8026 = ~\new_[7284]_  | (~\new_[9391]_  & ~\new_[7578]_ );
  assign n8031 = ~\new_[7285]_  | (~\new_[9604]_  & ~\new_[7565]_ );
  assign n8036 = ~\new_[7083]_  | (~\new_[9491]_  & ~\new_[7573]_ );
  assign n5901 = ~\new_[7286]_  | (~\new_[9605]_  & ~\new_[7568]_ );
  assign n8041 = ~\new_[7287]_  | (~\new_[9392]_  & ~\new_[7578]_ );
  assign n8046 = ~\new_[7288]_  | (~\new_[9546]_  & ~\new_[7578]_ );
  assign n8051 = ~\new_[7289]_  | (~\new_[9435]_  & ~\new_[7572]_ );
  assign n5881 = ~\new_[7290]_  | (~\new_[9606]_  & ~\new_[7573]_ );
  assign n8056 = ~\new_[7291]_  | (~\new_[9426]_  & ~\new_[7578]_ );
  assign n6746 = ~\new_[6914]_  | (~\new_[9457]_  & ~\new_[7540]_ );
  assign n8061 = ~\new_[7292]_  | (~\new_[9607]_  & ~\new_[7578]_ );
  assign n8066 = ~\new_[7293]_  | (~\new_[10026]_  & ~\new_[7578]_ );
  assign n5866 = ~\new_[7294]_  | (~\new_[10024]_  & ~\new_[7572]_ );
  assign n8071 = ~\new_[7295]_  | (~\new_[10109]_  & ~\new_[7573]_ );
  assign n8076 = ~\new_[7296]_  | (~\new_[10006]_  & ~\new_[7573]_ );
  assign n8081 = ~\new_[7297]_  | (~\new_[10110]_  & ~\new_[7572]_ );
  assign n5861 = ~\new_[7298]_  | (~\new_[10111]_  & ~\new_[7573]_ );
  assign n8086 = ~\new_[7299]_  | (~\new_[10112]_  & ~\new_[7576]_ );
  assign n8091 = ~\new_[7300]_  | (~\new_[9980]_  & ~\new_[7573]_ );
  assign n8096 = ~\new_[7301]_  | (~\new_[10113]_  & ~\new_[7577]_ );
  assign n5846 = ~\new_[7302]_  | (~\new_[9966]_  & ~\new_[7573]_ );
  assign n8101 = ~\new_[7303]_  | (~\new_[10114]_  & ~\new_[7574]_ );
  assign n8106 = ~\new_[6925]_  | (~\new_[9938]_  & ~\new_[7572]_ );
  assign n8111 = ~\new_[7304]_  | (~\new_[9934]_  & ~\new_[7576]_ );
  assign n5841 = ~\new_[7305]_  | (~\new_[9929]_  & ~\new_[7574]_ );
  assign n8116 = ~\new_[7306]_  | (~\new_[9931]_  & ~\new_[7573]_ );
  assign n8121 = ~\new_[7307]_  | (~\new_[9923]_  & ~\new_[7578]_ );
  assign n8126 = ~\new_[7308]_  | (~\new_[9952]_  & ~\new_[7577]_ );
  assign n5791 = ~\new_[7309]_  | (~\new_[10115]_  & ~\new_[7577]_ );
  assign n8131 = ~\new_[7310]_  | (~\new_[10116]_  & ~\new_[7565]_ );
  assign n8136 = ~\new_[7311]_  | (~\new_[9911]_  & ~\new_[7568]_ );
  assign n8141 = ~\new_[7312]_  | (~\new_[10118]_  & ~\new_[7572]_ );
  assign n5831 = ~\new_[6866]_  | (~\new_[9905]_  & ~\new_[7577]_ );
  assign n8146 = ~\new_[7313]_  | (~\new_[9903]_  & ~\new_[7578]_ );
  assign n8151 = ~\new_[7314]_  | (~\new_[9901]_  & ~\new_[7578]_ );
  assign n8156 = ~\new_[7316]_  | (~\new_[10120]_  & ~\new_[7565]_ );
  assign n5826 = ~\new_[7317]_  | (~\new_[9897]_  & ~\new_[7578]_ );
  assign n8161 = ~\new_[7318]_  | (~\new_[10088]_  & ~\new_[7572]_ );
  assign n8166 = ~\new_[7319]_  | (~\new_[10061]_  & ~\new_[7568]_ );
  assign n8171 = ~\new_[7320]_  | (~\new_[10122]_  & ~\new_[7568]_ );
  assign n5796 = ~\new_[7321]_  | (~\new_[10135]_  & ~\new_[7577]_ );
  assign n8176 = ~\new_[7322]_  | (~\new_[10133]_  & ~\new_[7577]_ );
  assign n8181 = ~\new_[7323]_  | (~\new_[10124]_  & ~\new_[7573]_ );
  assign n8186 = ~\new_[7324]_  | (~\new_[9622]_  & ~\new_[7565]_ );
  assign n5801 = ~\new_[7325]_  | (~\new_[9609]_  & ~\new_[7565]_ );
  assign n8191 = ~\new_[7326]_  | (~\new_[9590]_  & ~\new_[7565]_ );
  assign n8196 = ~\new_[7327]_  | (~\new_[9610]_  & ~\new_[7565]_ );
  assign n8201 = ~\new_[7328]_  | (~\new_[9623]_  & ~\new_[7570]_ );
  assign n5706 = ~\new_[7329]_  | (~\new_[9611]_  & ~\new_[7570]_ );
  assign n8206 = ~\new_[7330]_  | (~\new_[9548]_  & ~\new_[7570]_ );
  assign n8211 = ~\new_[7331]_  | (~\new_[9536]_  & ~\new_[7570]_ );
  assign n8216 = ~\new_[7332]_  | (~\new_[9429]_  & ~\new_[7567]_ );
  assign n5751 = ~\new_[7333]_  | (~\new_[9545]_  & ~\new_[7567]_ );
  assign n8221 = ~\new_[7334]_  | (~\new_[9446]_  & ~\new_[7567]_ );
  assign n8226 = ~\new_[7335]_  | (~\new_[9613]_  & ~\new_[7567]_ );
  assign n8231 = ~\new_[7336]_  | (~\new_[9356]_  & ~\new_[7576]_ );
  assign n5746 = ~\new_[7337]_  | (~\new_[9614]_  & ~\new_[7576]_ );
  assign n8241 = ~\new_[7338]_  | (~\new_[9432]_  & ~\new_[7576]_ );
  assign n8246 = ~\new_[7339]_  | (~\new_[9615]_  & ~\new_[7576]_ );
  assign n8251 = ~\new_[7340]_  | (~\new_[9599]_  & ~\new_[7569]_ );
  assign n5711 = ~\new_[7341]_  | (~\new_[9616]_  & ~\new_[7569]_ );
  assign n8256 = ~\new_[7342]_  | (~\new_[9635]_  & ~\new_[7566]_ );
  assign n8261 = ~\new_[7343]_  | (~\new_[9538]_  & ~\new_[7566]_ );
  assign n8266 = ~\new_[7344]_  | (~\new_[9621]_  & ~\new_[7566]_ );
  assign n5716 = ~\new_[7345]_  | (~\new_[9617]_  & ~\new_[7566]_ );
  assign n8271 = ~\new_[7346]_  | (~\new_[9588]_  & ~\new_[7569]_ );
  assign n8276 = ~\new_[7348]_  | (~\new_[9618]_  & ~\new_[7569]_ );
  assign n8281 = ~\new_[7349]_  | (~\new_[9585]_  & ~\new_[7571]_ );
  assign n5596 = ~\new_[7350]_  | (~\new_[9619]_  & ~\new_[7571]_ );
  assign n8286 = ~\new_[7351]_  | (~\new_[9540]_  & ~\new_[7568]_ );
  assign n8291 = ~\new_[7352]_  | (~\new_[9566]_  & ~\new_[7568]_ );
  assign n8296 = ~\new_[7353]_  | (~\new_[9612]_  & ~\new_[7571]_ );
  assign n5681 = ~\new_[7354]_  | (~\new_[9541]_  & ~\new_[7571]_ );
  assign n8301 = ~\new_[7355]_  | (~\new_[9367]_  & ~\new_[7568]_ );
  assign n8306 = ~\new_[7356]_  | (~\new_[9620]_  & ~\new_[7568]_ );
  assign n6611 = ~\new_[7359]_  | (~\new_[9949]_  & ~\new_[7542]_ );
  assign n8311 = ~\new_[7014]_  | (~\new_[10018]_  & ~\new_[7580]_ );
  assign n5676 = ~\new_[7361]_  | (~\new_[10098]_  & ~\new_[7590]_ );
  assign n8316 = ~\new_[7362]_  | (~\new_[10139]_  & ~\new_[7581]_ );
  assign n8321 = ~\new_[7047]_  | (~\new_[10042]_  & ~\new_[7581]_ );
  assign n8326 = ~\new_[7363]_  | (~\new_[10140]_  & ~\new_[7582]_ );
  assign n5601 = ~\new_[7364]_  | (~\new_[10039]_  & ~\new_[7591]_ );
  assign n8331 = ~\new_[7365]_  | (~\new_[10141]_  & ~\new_[7591]_ );
  assign n8336 = ~\new_[7148]_  | (~\new_[10049]_  & ~\new_[7585]_ );
  assign n8341 = ~\new_[7366]_  | (~\new_[10142]_  & ~\new_[7585]_ );
  assign n5606 = ~\new_[7368]_  | (~\new_[10046]_  & ~\new_[7591]_ );
  assign n8346 = ~\new_[7370]_  | (~\new_[10143]_  & ~\new_[7591]_ );
  assign n8351 = ~\new_[7050]_  | (~\new_[10044]_  & ~\new_[7586]_ );
  assign n8356 = ~\new_[7371]_  | (~\new_[10144]_  & ~\new_[7590]_ );
  assign n5511 = ~\new_[7372]_  | (~\new_[10043]_  & ~\new_[7582]_ );
  assign n8361 = ~\new_[7373]_  | (~\new_[10145]_  & ~\new_[7582]_ );
  assign n8366 = ~\new_[7046]_  | (~\new_[10033]_  & ~\new_[7591]_ );
  assign n8371 = ~\new_[7374]_  | (~\new_[10146]_  & ~\new_[7590]_ );
  assign n5561 = ~\new_[7375]_  | (~\new_[10030]_  & ~\new_[7590]_ );
  assign n8381 = ~\new_[7376]_  | (~\new_[9627]_  & ~\new_[7543]_ );
  assign n8376 = ~\new_[7377]_  | (~\new_[10147]_  & ~\new_[7583]_ );
  assign \new_[6237]_  = (~\new_[7504]_  | ~\new_[12914]_ ) & (~\new_[12956]_  | ~\new_[12636]_ );
  assign n8386 = ~\new_[7378]_  | (~\new_[10047]_  & ~\new_[7583]_ );
  assign n8391 = ~\new_[7379]_  | (~\new_[9628]_  & ~\new_[7543]_ );
  assign n8396 = ~\new_[7412]_  | (~\new_[10137]_  & ~\new_[7585]_ );
  assign \new_[6241]_  = (~\new_[7505]_  | ~\new_[12985]_ ) & (~\new_[13055]_  | ~\new_[12637]_ );
  assign n5516 = ~\new_[7038]_  | (~\new_[9629]_  & ~\new_[7543]_ );
  assign n8401 = ~\new_[7381]_  | (~\new_[10148]_  & ~\new_[7585]_ );
  assign n8406 = ~\new_[7382]_  | (~\new_[10037]_  & ~\new_[7587]_ );
  assign n8416 = ~\new_[7383]_  | (~\new_[9368]_  & ~\new_[7543]_ );
  assign n6431 = ~\new_[6849]_  | (~\new_[10517]_  & ~\new_[7581]_ );
  assign n5521 = ~\new_[6884]_  | (~\new_[10028]_  & ~\new_[7584]_ );
  assign n8426 = ~\new_[7385]_  | (~\new_[9369]_  & ~\new_[7542]_ );
  assign n8431 = ~\new_[7386]_  | (~\new_[9933]_  & ~\new_[7589]_ );
  assign n8441 = ~\new_[7255]_  | (~\new_[10125]_  & ~\new_[7587]_ );
  assign n5481 = ~\new_[7256]_  | (~\new_[9584]_  & ~\new_[7532]_ );
  assign n8446 = ~\new_[7389]_  | (~\new_[10153]_  & ~\new_[7587]_ );
  assign n8451 = ~\new_[7390]_  | (~\new_[10152]_  & ~\new_[7589]_ );
  assign n8461 = ~\new_[7391]_  | (~\new_[9631]_  & ~\new_[7542]_ );
  assign n8456 = ~\new_[7392]_  | (~\new_[10099]_  & ~\new_[7590]_ );
  assign n8466 = ~\new_[7393]_  | (~\new_[10154]_  & ~\new_[7579]_ );
  assign n8476 = ~\new_[7191]_  | (~\new_[9632]_  & ~\new_[7542]_ );
  assign n8471 = ~\new_[7177]_  | (~\new_[10096]_  & ~\new_[7579]_ );
  assign n8481 = ~\new_[7394]_  | (~\new_[10083]_  & ~\new_[7584]_ );
  assign n8486 = ~\new_[7395]_  | (~\new_[9535]_  & ~\new_[7545]_ );
  assign n5451 = ~\new_[6883]_  | (~\new_[10077]_  & ~\new_[7579]_ );
  assign n8491 = ~\new_[7397]_  | (~\new_[9940]_  & ~\new_[7583]_ );
  assign n5456 = ~\new_[7398]_  | (~\new_[9633]_  & ~\new_[7543]_ );
  assign n8496 = ~\new_[7399]_  | (~\new_[9939]_  & ~\new_[7583]_ );
  assign n8501 = ~\new_[7400]_  | (~\new_[9937]_  & ~\new_[7587]_ );
  assign n8506 = ~\new_[6927]_  | (~\new_[9935]_  & ~\new_[7587]_ );
  assign n5336 = ~\new_[7402]_  | (~\new_[10155]_  & ~\new_[7587]_ );
  assign n8521 = ~\new_[7048]_  | (~\new_[9636]_  & ~\new_[7543]_ );
  assign n8516 = ~\new_[7396]_  | (~\new_[10157]_  & ~\new_[7590]_ );
  assign n8526 = ~\new_[7403]_  | (~\new_[10149]_  & ~\new_[7586]_ );
  assign n8531 = ~\new_[7404]_  | (~\new_[9625]_  & ~\new_[7543]_ );
  assign n5396 = ~\new_[7360]_  | (~\new_[10136]_  & ~\new_[7586]_ );
  assign n8536 = ~\new_[7405]_  | (~\new_[10034]_  & ~\new_[7586]_ );
  assign n5391 = ~\new_[7406]_  | (~\new_[9637]_  & ~\new_[7542]_ );
  assign n8541 = ~\new_[7277]_  | (~\new_[10129]_  & ~\new_[7586]_ );
  assign n8546 = ~\new_[7407]_  | (~\new_[10040]_  & ~\new_[7580]_ );
  assign n8551 = ~\new_[7315]_  | (~\new_[10123]_  & ~\new_[7590]_ );
  assign n5346 = ~\new_[7409]_  | (~\new_[10156]_  & ~\new_[7580]_ );
  assign n8566 = ~\new_[7283]_  | (~\new_[9640]_  & ~\new_[7532]_ );
  assign n8561 = ~\new_[7280]_  | (~\new_[10101]_  & ~\new_[7580]_ );
  assign n8571 = ~\new_[7410]_  | (~\new_[10106]_  & ~\new_[7581]_ );
  assign n8576 = ~\new_[7411]_  | (~\new_[9393]_  & ~\new_[7542]_ );
  assign n5351 = ~\new_[7019]_  | (~\new_[9996]_  & ~\new_[7581]_ );
  assign n8581 = ~\new_[7413]_  | (~\new_[9956]_  & ~\new_[7586]_ );
  assign n9386 = ~\new_[7414]_  | (~\new_[9641]_  & ~\new_[7542]_ );
  assign n8586 = ~\new_[7415]_  | (~\new_[9954]_  & ~\new_[7586]_ );
  assign n8591 = ~\new_[7416]_  | (~\new_[9951]_  & ~\new_[7582]_ );
  assign n8596 = ~\new_[6941]_  | (~\new_[9950]_  & ~\new_[7591]_ );
  assign \new_[6289]_  = ~\new_[7429]_  & (~\new_[12734]_  | ~\new_[7599]_ );
  assign n6391 = ~\new_[6935]_  | (~\new_[9355]_  & ~\new_[7544]_ );
  assign n6386 = ~\new_[6936]_  | (~\new_[9946]_  & ~\new_[7591]_ );
  assign \new_[6292]_  = ~\new_[7430]_  & (~\new_[12754]_  | ~\new_[7601]_ );
  assign n8966 = \new_[5651]_  ? \new_[7451]_  : \new_[10522]_ ;
  assign n9001 = \new_[5658]_  ? \new_[7451]_  : \new_[10694]_ ;
  assign n8936 = \new_[5645]_  ? \new_[7451]_  : \new_[10531]_ ;
  assign n8611 = \new_[5580]_  ? \new_[7552]_  : \new_[10546]_ ;
  assign n8606 = \new_[5579]_  ? \new_[7552]_  : \new_[10545]_ ;
  assign n8616 = \new_[5581]_  ? \new_[7552]_  : \new_[10547]_ ;
  assign n9356 = \new_[5753]_  ? \new_[7552]_  : \new_[10548]_ ;
  assign n8621 = \new_[5582]_  ? \new_[7552]_  : \new_[10551]_ ;
  assign n9306 = \new_[5735]_  ? \new_[7552]_  : \new_[10555]_ ;
  assign n8626 = \new_[5583]_  ? \new_[7552]_  : \new_[10557]_ ;
  assign n8631 = \new_[5584]_  ? \new_[7552]_  : \new_[10559]_ ;
  assign n9341 = \new_[5748]_  ? \new_[7552]_  : \new_[10560]_ ;
  assign n8636 = \new_[5585]_  ? \new_[7552]_  : \new_[10561]_ ;
  assign n9296 = \new_[5733]_  ? \new_[7552]_  : \new_[10563]_ ;
  assign n8641 = \new_[5586]_  ? \new_[7552]_  : \new_[10566]_ ;
  assign n8656 = \new_[5589]_  ? \new_[7552]_  : \new_[10567]_ ;
  assign n8646 = \new_[5587]_  ? \new_[7552]_  : \new_[10568]_ ;
  assign n8651 = \new_[5588]_  ? \new_[7552]_  : \new_[10569]_ ;
  assign n8666 = \new_[5591]_  ? \new_[7552]_  : \new_[10570]_ ;
  assign n8661 = \new_[5590]_  ? \new_[7552]_  : \new_[10571]_ ;
  assign n9261 = \new_[5726]_  ? \new_[7552]_  : \new_[10572]_ ;
  assign n8671 = \new_[5592]_  ? \new_[7552]_  : \new_[10574]_ ;
  assign n8676 = \new_[5593]_  ? \new_[7552]_  : \new_[10554]_ ;
  assign n9226 = \new_[5719]_  ? \new_[7552]_  : \new_[10576]_ ;
  assign n8681 = \new_[5594]_  ? \new_[7552]_  : \new_[10578]_ ;
  assign n8996 = \new_[5657]_  ? \new_[7451]_  : \new_[10692]_ ;
  assign n9246 = \new_[5723]_  ? \new_[7561]_  : \new_[10585]_ ;
  assign n8686 = \new_[5595]_  ? \new_[7561]_  : \new_[10586]_ ;
  assign n8691 = \new_[5596]_  ? \new_[7561]_  : \new_[10587]_ ;
  assign n9216 = \new_[5717]_  ? \new_[7561]_  : \new_[10588]_ ;
  assign n8696 = \new_[5597]_  ? \new_[7561]_  : \new_[10590]_ ;
  assign n9206 = \new_[5715]_  ? \new_[7561]_  : \new_[10592]_ ;
  assign n8701 = \new_[5598]_  ? \new_[7561]_  : \new_[10593]_ ;
  assign n8706 = \new_[5599]_  ? \new_[7561]_  : \new_[10595]_ ;
  assign n9176 = \new_[5702]_  ? \new_[7561]_  : \new_[10596]_ ;
  assign n8711 = \new_[5600]_  ? \new_[7561]_  : \new_[10597]_ ;
  assign n9116 = \new_[5687]_  ? \new_[7561]_  : \new_[10599]_ ;
  assign n8731 = \new_[5604]_  ? \new_[7561]_  : \new_[10601]_ ;
  assign n8721 = \new_[5602]_  ? \new_[7561]_  : \new_[10603]_ ;
  assign n8726 = \new_[5603]_  ? \new_[7561]_  : \new_[10637]_ ;
  assign n9156 = \new_[5695]_  ? \new_[7561]_  : \new_[10604]_ ;
  assign n8741 = \new_[5606]_  ? \new_[7561]_  : \new_[10605]_ ;
  assign n8736 = \new_[5605]_  ? \new_[7561]_  : \new_[10607]_ ;
  assign n9111 = \new_[5686]_  ? \new_[7561]_  : \new_[10608]_ ;
  assign n8746 = \new_[5607]_  ? \new_[7561]_  : \new_[10610]_ ;
  assign n8751 = \new_[5608]_  ? \new_[7561]_  : \new_[10615]_ ;
  assign n9096 = \new_[5677]_  ? \new_[7561]_  : \new_[10616]_ ;
  assign n8756 = \new_[5609]_  ? \new_[7561]_  : \new_[10613]_ ;
  assign n9056 = \new_[5669]_  ? \new_[7528]_  : \new_[10619]_ ;
  assign n8761 = \new_[5610]_  ? \new_[7528]_  : \new_[10620]_ ;
  assign n8766 = \new_[5611]_  ? \new_[7528]_  : \new_[10711]_ ;
  assign n5671 = \new_[4986]_  ? \new_[7528]_  : \new_[10621]_ ;
  assign n8771 = \new_[5612]_  ? \new_[7528]_  : \new_[10624]_ ;
  assign n7501 = \new_[5358]_  ? \new_[7528]_  : \new_[10700]_ ;
  assign n8781 = \new_[5614]_  ? \new_[7528]_  : \new_[10626]_ ;
  assign n8786 = \new_[5615]_  ? \new_[7528]_  : \new_[10654]_ ;
  assign n8236 = \new_[5505]_  ? \new_[7528]_  : \new_[10672]_ ;
  assign n8791 = \new_[5616]_  ? \new_[7528]_  : \new_[10673]_ ;
  assign n5946 = \new_[5047]_  ? \new_[7528]_  : \new_[10627]_ ;
  assign n8806 = \new_[5619]_  ? \new_[7528]_  : \new_[10666]_ ;
  assign n8796 = \new_[5617]_  ? \new_[7528]_  : \new_[10628]_ ;
  assign n8801 = \new_[5618]_  ? \new_[7528]_  : \new_[10664]_ ;
  assign n5876 = \new_[5033]_  ? \new_[7528]_  : \new_[10661]_ ;
  assign n8816 = \new_[5621]_  ? \new_[7528]_  : \new_[10652]_ ;
  assign n8811 = \new_[5620]_  ? \new_[7528]_  : \new_[10630]_ ;
  assign n5851 = \new_[5028]_  ? \new_[7528]_  : \new_[10631]_ ;
  assign n8821 = \new_[5622]_  ? \new_[7528]_  : \new_[10655]_ ;
  assign n8826 = \new_[5623]_  ? \new_[7528]_  : \new_[10633]_ ;
  assign n5856 = \new_[5029]_  ? \new_[7528]_  : \new_[10639]_ ;
  assign n8831 = \new_[5624]_  ? \new_[7528]_  : \new_[10635]_ ;
  assign n5776 = \new_[5009]_  ? \new_[7575]_  : \new_[10602]_ ;
  assign n8836 = \new_[5625]_  ? \new_[7575]_  : \new_[10623]_ ;
  assign n8841 = \new_[5626]_  ? \new_[7575]_  : \new_[10543]_ ;
  assign n5701 = \new_[4994]_  ? \new_[7575]_  : \new_[10556]_ ;
  assign n8846 = \new_[5627]_  ? \new_[7575]_  : \new_[10644]_ ;
  assign n5771 = \new_[5008]_  ? \new_[7575]_  : \new_[10645]_ ;
  assign n8851 = \new_[5628]_  ? \new_[7575]_  : \new_[10712]_ ;
  assign n8856 = \new_[5629]_  ? \new_[7575]_  : \new_[10710]_ ;
  assign n5341 = \new_[4897]_  ? \new_[7575]_  : \new_[10646]_ ;
  assign n8861 = \new_[5630]_  ? \new_[7575]_  : \new_[10708]_ ;
  assign n5631 = \new_[4978]_  ? \new_[7575]_  : \new_[10707]_ ;
  assign n8866 = \new_[5631]_  ? \new_[7575]_  : \new_[10705]_ ;
  assign n8881 = \new_[5634]_  ? \new_[7575]_  : \new_[10649]_ ;
  assign n8871 = \new_[5632]_  ? \new_[7575]_  : \new_[10674]_ ;
  assign n8876 = \new_[5633]_  ? \new_[7575]_  : \new_[10650]_ ;
  assign n8891 = \new_[5636]_  ? \new_[7575]_  : \new_[10671]_ ;
  assign n8886 = \new_[5635]_  ? \new_[7575]_  : \new_[10669]_ ;
  assign n5501 = \new_[4941]_  ? \new_[7575]_  : \new_[10668]_ ;
  assign n8896 = \new_[5637]_  ? \new_[7575]_  : \new_[10665]_ ;
  assign n8901 = \new_[5638]_  ? \new_[7575]_  : \new_[10662]_ ;
  assign n5576 = \new_[4967]_  ? \new_[7575]_  : \new_[10653]_ ;
  assign n8906 = \new_[5639]_  ? \new_[7575]_  : \new_[10658]_ ;
  assign n8911 = \new_[5640]_  ? \new_[7451]_  : \new_[10541]_ ;
  assign n5556 = \new_[4963]_  ? \new_[7451]_  : \new_[10675]_ ;
  assign n5421 = \new_[4913]_  ? \new_[7608]_  : \new_[10677]_ ;
  assign n8916 = \new_[5641]_  ? \new_[7588]_  : \new_[10678]_ ;
  assign n5331 = \new_[4895]_  ? \new_[7451]_  : \new_[10536]_ ;
  assign n8926 = \new_[5643]_  ? \new_[7451]_  : \new_[10679]_ ;
  assign n8921 = \new_[5642]_  ? \new_[7588]_  : \new_[10534]_ ;
  assign n8931 = \new_[5644]_  ? \new_[7588]_  : \new_[10680]_ ;
  assign n5416 = \new_[4912]_  ? \new_[7588]_  : \new_[10530]_ ;
  assign n9266 = \new_[5727]_  ? \new_[7588]_  : \new_[10681]_ ;
  assign n8941 = \new_[5646]_  ? \new_[7588]_  : \new_[10683]_ ;
  assign n8951 = \new_[5648]_  ? \new_[7451]_  : \new_[10684]_ ;
  assign n8946 = \new_[5647]_  ? \new_[7588]_  : \new_[10528]_ ;
  assign n9421 = \new_[5766]_  ? \new_[7588]_  : \new_[10527]_ ;
  assign n8956 = \new_[5649]_  ? \new_[7588]_  : \new_[10526]_ ;
  assign n8961 = \new_[5650]_  ? \new_[7588]_  : \new_[10525]_ ;
  assign n9366 = \new_[5755]_  ? \new_[7588]_  : \new_[10523]_ ;
  assign n8971 = \new_[5652]_  ? \new_[7588]_  : \new_[10521]_ ;
  assign n9301 = \new_[5734]_  ? \new_[7451]_  : \new_[10686]_ ;
  assign n8976 = \new_[5653]_  ? \new_[7588]_  : \new_[10519]_ ;
  assign n8981 = \new_[5654]_  ? \new_[7588]_  : \new_[10688]_ ;
  assign n8986 = \new_[5655]_  ? \new_[7451]_  : \new_[10656]_ ;
  assign n9336 = \new_[5744]_  ? \new_[7588]_  : \new_[10640]_ ;
  assign n8991 = \new_[5656]_  ? \new_[7451]_  : \new_[10690]_ ;
  assign n9286 = \new_[5731]_  ? \new_[7588]_  : \new_[10583]_ ;
  assign n9181 = \new_[5703]_  ? \new_[7588]_  : \new_[10532]_ ;
  assign n9256 = \new_[5725]_  ? \new_[7588]_  : \new_[10524]_ ;
  assign n9016 = \new_[5661]_  ? \new_[7588]_  : \new_[10581]_ ;
  assign n9006 = \new_[5659]_  ? \new_[7588]_  : \new_[10706]_ ;
  assign n9011 = \new_[5660]_  ? \new_[7588]_  : \new_[10641]_ ;
  assign n9021 = \new_[5662]_  ? \new_[7588]_  : \new_[10697]_ ;
  assign n9026 = \new_[5663]_  ? \new_[7451]_  : \new_[10698]_ ;
  assign n9031 = \new_[5664]_  ? \new_[7608]_  : \new_[10584]_ ;
  assign n9171 = \new_[5701]_  ? \new_[7451]_  : \new_[10701]_ ;
  assign n9036 = \new_[5665]_  ? \new_[7451]_  : \new_[10704]_ ;
  assign n9146 = \new_[5693]_  ? \new_[7451]_  : \new_[10580]_ ;
  assign \new_[6421]_  = u14_u7_en_out_l2_reg;
  assign \new_[6422]_  = ~\new_[12519]_  | ~\new_[7588]_  | ~\new_[12340]_ ;
  assign \new_[6423]_  = ~\new_[12886]_  | ~\new_[7552]_  | ~\new_[12342]_ ;
  assign \new_[6424]_  = ~\new_[12691]_  | ~\new_[7561]_  | ~\new_[11800]_ ;
  assign \new_[6425]_  = ~\new_[13012]_  | ~\new_[7451]_  | ~\new_[11813]_ ;
  assign \new_[6426]_  = ~\new_[12993]_  | ~\new_[7528]_  | ~\new_[11956]_ ;
  assign \new_[6427]_  = ~\new_[12686]_  | ~\new_[7575]_  | ~\new_[11889]_ ;
  assign n5641 = ~\new_[13886]_ ;
  assign \new_[6429]_  = \new_[12811]_  | \new_[13885]_ ;
  assign n5646 = ~\new_[6785]_ ;
  assign \new_[6431]_  = \new_[12718]_  | \new_[13885]_ ;
  assign n5651 = ~\new_[6786]_ ;
  assign \new_[6433]_  = \new_[12710]_  | \new_[13885]_ ;
  assign n5656 = ~\new_[6787]_ ;
  assign \new_[6435]_  = \new_[12853]_  | \new_[13885]_ ;
  assign n5661 = ~\new_[6788]_ ;
  assign \new_[6437]_  = \new_[13168]_  | \new_[13885]_ ;
  assign n5666 = ~\new_[6789]_ ;
  assign \new_[6439]_  = \new_[13885]_  | \new_[14093]_ ;
  assign \new_[6440]_  = u14_u7_full_empty_r_reg;
  assign \new_[6441]_  = ~u13_ac97_rst_force_reg;
  assign \new_[6442]_  = u13_resume_req_reg;
  assign \new_[6443]_  = ~\new_[13014]_  & ~\new_[7431]_ ;
  assign \new_[6444]_  = ~\new_[14187]_  & ~\new_[7432]_ ;
  assign \new_[6445]_  = ~\new_[12917]_  & ~\new_[7433]_ ;
  assign \new_[6446]_  = ~\new_[12979]_  & ~\new_[7434]_ ;
  assign \new_[6447]_  = ~\new_[7431]_  & ~\new_[13605]_ ;
  assign \new_[6448]_  = ~\new_[7432]_  & ~\new_[13437]_ ;
  assign \new_[6449]_  = ~\new_[7433]_  & ~\new_[13168]_ ;
  assign \new_[6450]_  = ~\new_[7434]_  & ~\new_[14093]_ ;
  assign n6326 = \new_[13218]_  ? n9791 : \new_[13166]_ ;
  assign n6331 = \new_[13813]_  ? n9791 : \new_[13162]_ ;
  assign n6336 = \new_[13689]_  ? n9791 : \new_[13111]_ ;
  assign n6341 = \new_[13324]_  ? n9791 : \new_[13090]_ ;
  assign n6346 = \new_[13611]_  ? n9791 : \new_[13122]_ ;
  assign n5911 = \new_[13614]_  ? n9791 : \new_[13187]_ ;
  assign n6351 = \new_[13632]_  ? n9791 : \new_[13133]_ ;
  assign n6356 = \new_[13509]_  ? n9791 : \new_[13189]_ ;
  assign n6361 = \new_[13382]_  ? n9791 : \new_[13177]_ ;
  assign n6366 = \new_[13704]_  ? n9791 : \new_[13087]_ ;
  assign n5891 = \new_[13790]_  ? n9791 : \new_[13183]_ ;
  assign n6371 = \new_[13370]_  ? n9791 : \new_[13172]_ ;
  assign n6376 = \new_[13671]_  ? n9791 : \new_[13163]_ ;
  assign n9046 = \new_[13269]_  ? n9791 : \new_[13086]_ ;
  assign n6381 = \new_[13505]_  ? n9791 : \new_[13184]_ ;
  assign n5896 = \new_[13730]_  ? n9791 : \new_[13179]_ ;
  assign n5961 = \new_[5050]_  ? n9791 : \new_[13185]_ ;
  assign n9121 = \new_[5688]_  ? n9791 : \new_[13173]_ ;
  assign n5966 = \new_[5051]_  ? n9791 : \new_[13182]_ ;
  assign n5971 = \new_[5052]_  ? n9791 : \new_[13136]_ ;
  assign n5976 = \new_[5053]_  ? n9791 : \new_[13164]_ ;
  assign n5981 = \new_[5054]_  ? n9791 : \new_[13167]_ ;
  assign n5326 = \new_[4894]_  ? n9791 : \new_[13128]_ ;
  assign n5986 = \new_[5055]_  ? n9791 : \new_[13117]_ ;
  assign n5991 = \new_[13866]_  ? \new_[7441]_  : \new_[13166]_ ;
  assign n5996 = \new_[13157]_  ? \new_[7441]_  : \new_[13162]_ ;
  assign n5936 = \new_[13108]_  ? \new_[7441]_  : \new_[13111]_ ;
  assign n6001 = \new_[5058]_  ? \new_[7441]_  : \new_[13090]_ ;
  assign n6006 = \new_[5059]_  ? \new_[7441]_  : \new_[13122]_ ;
  assign n6011 = \new_[13088]_  ? \new_[7441]_  : \new_[13187]_ ;
  assign n5951 = \new_[5048]_  ? \new_[7441]_  : \new_[13133]_ ;
  assign n6016 = \new_[13876]_  ? \new_[7441]_  : \new_[13185]_ ;
  assign n6021 = \new_[5062]_  ? \new_[7441]_  : \new_[13182]_ ;
  assign n6026 = \new_[13155]_  ? \new_[7441]_  : \new_[13173]_ ;
  assign n5956 = \new_[13098]_  ? \new_[7441]_  : \new_[13136]_ ;
  assign n6031 = \new_[5064]_  ? \new_[7441]_  : \new_[13189]_ ;
  assign n6036 = \new_[5065]_  ? \new_[7441]_  : \new_[13164]_ ;
  assign n6041 = \new_[5066]_  ? \new_[7441]_  : \new_[13167]_ ;
  assign n5906 = \new_[5039]_  ? \new_[7441]_  : \new_[13128]_ ;
  assign n6046 = \new_[5067]_  ? \new_[7441]_  : \new_[13106]_ ;
  assign n6051 = \new_[13130]_  ? \new_[7441]_  : \new_[13177]_ ;
  assign n6056 = \new_[13129]_  ? \new_[7441]_  : \new_[13183]_ ;
  assign n6061 = \new_[5070]_  ? \new_[7441]_  : \new_[13087]_ ;
  assign n6066 = \new_[5071]_  ? \new_[7441]_  : \new_[13172]_ ;
  assign n6071 = \new_[13181]_  ? \new_[7441]_  : \new_[13163]_ ;
  assign n6076 = \new_[5073]_  ? \new_[7441]_  : \new_[13086]_ ;
  assign n5446 = \new_[13873]_  ? \new_[7441]_  : \new_[13184]_ ;
  assign n6081 = \new_[5074]_  ? \new_[7441]_  : \new_[13179]_ ;
  assign n6086 = \new_[13166]_  ? \new_[7443]_  : \new_[13012]_ ;
  assign n6091 = \new_[13162]_  ? \new_[7443]_  : \new_[5076]_ ;
  assign n5366 = \new_[13111]_  ? \new_[7443]_  : \new_[4902]_ ;
  assign n6096 = \new_[13090]_  ? \new_[7443]_  : \new_[5077]_ ;
  assign n6101 = \new_[13122]_  ? \new_[7443]_  : \new_[5078]_ ;
  assign n6106 = \new_[13187]_  ? \new_[7443]_  : \new_[5079]_ ;
  assign n9371 = \new_[13133]_  ? \new_[7443]_  : \new_[5756]_ ;
  assign n6111 = \new_[13185]_  ? \new_[7443]_  : \new_[12691]_ ;
  assign n6116 = \new_[13182]_  ? \new_[7443]_  : \new_[5081]_ ;
  assign n6121 = \new_[13173]_  ? \new_[7443]_  : \new_[5082]_ ;
  assign n9211 = \new_[13136]_  ? \new_[7443]_  : \new_[5716]_ ;
  assign n6126 = \new_[13189]_  ? \new_[7443]_  : \new_[5083]_ ;
  assign n6131 = \new_[13164]_  ? \new_[7443]_  : \new_[5084]_ ;
  assign n6136 = \new_[13167]_  ? \new_[7443]_  : \new_[5085]_ ;
  assign n9076 = \new_[13128]_  ? \new_[7443]_  : \new_[13085]_ ;
  assign n6141 = \new_[13106]_  ? \new_[7443]_  : \new_[5086]_ ;
  assign n6146 = \new_[13094]_  ? \new_[7443]_  : \new_[12993]_ ;
  assign n6151 = \new_[13176]_  ? \new_[7443]_  : \new_[5088]_ ;
  assign n9151 = \new_[13095]_  ? \new_[7443]_  : \new_[5694]_ ;
  assign n6156 = \new_[13156]_  ? \new_[7443]_  : \new_[5089]_ ;
  assign n6161 = \new_[13159]_  ? \new_[7443]_  : \new_[5090]_ ;
  assign n6166 = \new_[13123]_  ? \new_[7443]_  : \new_[5091]_ ;
  assign n5916 = \new_[13177]_  ? \new_[7443]_  : \new_[5041]_ ;
  assign n6171 = \new_[13132]_  ? \new_[7443]_  : \new_[5092]_ ;
  assign n6176 = \new_[13117]_  ? \new_[7443]_  : \new_[5093]_ ;
  assign n6181 = \new_[13183]_  ? \new_[7443]_  : \new_[5094]_ ;
  assign n5921 = \new_[13087]_  ? \new_[7443]_  : \new_[5042]_ ;
  assign n6186 = \new_[13172]_  ? \new_[7443]_  : \new_[5095]_ ;
  assign n6191 = \new_[13163]_  ? \new_[7443]_  : \new_[5096]_ ;
  assign n6196 = \new_[13086]_  ? \new_[7443]_  : \new_[5097]_ ;
  assign n5441 = \new_[13184]_  ? \new_[7443]_  : \new_[12886]_ ;
  assign n6201 = \new_[13179]_  ? \new_[7443]_  : \new_[5098]_ ;
  assign n6206 = \new_[5099]_  ? \new_[7442]_  : \new_[13166]_ ;
  assign n6211 = \new_[5100]_  ? \new_[7442]_  : \new_[13162]_ ;
  assign n6216 = \new_[5101]_  ? \new_[7442]_  : \new_[13111]_ ;
  assign n6221 = \new_[5102]_  ? \new_[7442]_  : \new_[13090]_ ;
  assign n6226 = \new_[5103]_  ? \new_[7442]_  : \new_[13122]_ ;
  assign n6231 = \new_[5104]_  ? \new_[7442]_  : \new_[13187]_ ;
  assign n6321 = \new_[5122]_  ? \new_[7442]_  : \new_[13133]_ ;
  assign n6236 = \new_[5105]_  ? \new_[7442]_  : \new_[13185]_ ;
  assign n6241 = \new_[5106]_  ? \new_[7442]_  : \new_[13182]_ ;
  assign n6246 = \new_[5107]_  ? \new_[7442]_  : \new_[13173]_ ;
  assign n6251 = \new_[5108]_  ? \new_[7442]_  : \new_[13136]_ ;
  assign n6256 = \new_[5109]_  ? \new_[7442]_  : \new_[13189]_ ;
  assign n6261 = \new_[5110]_  ? \new_[7442]_  : \new_[13164]_ ;
  assign n6266 = \new_[5111]_  ? \new_[7442]_  : \new_[13167]_ ;
  assign n5931 = \new_[5044]_  ? \new_[7442]_  : \new_[13128]_ ;
  assign n6271 = \new_[5112]_  ? \new_[7442]_  : \new_[13106]_ ;
  assign n6276 = \new_[5113]_  ? \new_[7442]_  : \new_[13094]_ ;
  assign n6281 = \new_[5114]_  ? \new_[7442]_  : \new_[13176]_ ;
  assign n9066 = \new_[5671]_  ? \new_[7442]_  : \new_[13095]_ ;
  assign n6286 = \new_[5115]_  ? \new_[7442]_  : \new_[13156]_ ;
  assign n6291 = \new_[5116]_  ? \new_[7442]_  : \new_[13159]_ ;
  assign n6296 = \new_[5117]_  ? \new_[7442]_  : \new_[13177]_ ;
  assign n9161 = \new_[5696]_  ? \new_[7442]_  : \new_[13183]_ ;
  assign n6316 = \new_[5121]_  ? \new_[7442]_  : \new_[13087]_ ;
  assign n6301 = \new_[5118]_  ? \new_[7442]_  : \new_[13172]_ ;
  assign n6306 = \new_[5119]_  ? \new_[7442]_  : \new_[13163]_ ;
  assign n5926 = \new_[5043]_  ? \new_[7442]_  : \new_[13086]_ ;
  assign n8716 = \new_[5601]_  ? \new_[7442]_  : \new_[13184]_ ;
  assign n6311 = \new_[5120]_  ? \new_[7442]_  : \new_[13179]_ ;
  assign \new_[6560]_  = ~\new_[6830]_ ;
  assign \new_[6561]_  = ~\new_[6832]_ ;
  assign \new_[6562]_  = ~\new_[6835]_ ;
  assign n9106 = \\u1_sr_reg[9] ;
  assign \new_[6564]_  = ~\new_[8413]_  & (~\new_[7481]_  | ~\new_[9752]_ );
  assign \new_[6565]_  = ~\new_[12479]_  & (~\new_[12435]_  | ~\new_[7461]_ );
  assign \new_[6566]_  = ~\new_[12480]_  & (~\new_[12605]_  | ~\new_[7462]_ );
  assign \new_[6567]_  = ~\new_[12453]_  & (~\new_[12612]_  | ~\new_[7463]_ );
  assign \new_[6568]_  = (~\new_[11524]_  | ~\new_[7588]_ ) & (~\new_[7616]_  | ~\new_[4757]_ );
  assign \new_[6569]_  = (~\new_[10094]_  | ~\new_[7608]_ ) & (~\new_[7533]_  | ~\new_[4758]_ );
  assign \new_[6570]_  = (~\new_[10035]_  | ~\new_[7552]_ ) & (~\new_[7610]_  | ~\new_[4768]_ );
  assign \new_[6571]_  = (~\new_[10078]_  | ~\new_[7561]_ ) & (~\new_[7612]_  | ~\new_[4759]_ );
  assign \new_[6572]_  = (~\new_[10041]_  | ~\new_[7528]_ ) & (~\new_[7605]_  | ~\new_[4754]_ );
  assign \new_[6573]_  = (~\new_[10128]_  | ~\new_[7575]_ ) & (~\new_[7614]_  | ~\new_[4760]_ );
  assign n6396 = ~\new_[6843]_  | (~\new_[9944]_  & ~\new_[7584]_ );
  assign n6401 = ~\new_[6844]_  | (~\new_[9388]_  & ~\new_[7542]_ );
  assign n5871 = ~\new_[6933]_  | (~\new_[9943]_  & ~\new_[7589]_ );
  assign n6406 = ~\new_[6845]_  | (~\new_[9942]_  & ~\new_[7586]_ );
  assign n5836 = ~\new_[6846]_  | (~\new_[9357]_  & ~\new_[7543]_ );
  assign n6411 = ~\new_[6931]_  | (~\new_[9941]_  & ~\new_[7591]_ );
  assign n6416 = ~\new_[6847]_  | (~\new_[9910]_  & ~\new_[7584]_ );
  assign n6476 = ~\new_[6857]_  | (~\new_[10494]_  & ~\new_[7589]_ );
  assign n6421 = ~\new_[6890]_  | (~\new_[10480]_  & ~\new_[7589]_ );
  assign n5821 = ~\new_[7149]_  | (~\new_[10507]_  & ~\new_[7584]_ );
  assign n6436 = ~\new_[7369]_  | (~\new_[9359]_  & ~\new_[7542]_ );
  assign n6441 = ~\new_[7367]_  | (~\new_[10516]_  & ~\new_[7585]_ );
  assign n5811 = ~\new_[6850]_  | (~\new_[9360]_  & ~\new_[7543]_ );
  assign n6446 = ~\new_[6851]_  | (~\new_[10477]_  & ~\new_[7582]_ );
  assign n6456 = ~\new_[6852]_  | (~\new_[10513]_  & ~\new_[7582]_ );
  assign n5816 = ~\new_[6853]_  | (~\new_[10482]_  & ~\new_[7579]_ );
  assign n6451 = ~\new_[7358]_  | (~\new_[9361]_  & ~\new_[7543]_ );
  assign n6461 = ~\new_[7347]_  | (~\new_[10511]_  & ~\new_[7580]_ );
  assign n6471 = ~\new_[6854]_  | (~\new_[9362]_  & ~\new_[7532]_ );
  assign n6466 = ~\new_[6855]_  | (~\new_[10515]_  & ~\new_[7581]_ );
  assign n5806 = ~\new_[6856]_  | (~\new_[10492]_  & ~\new_[7581]_ );
  assign n6481 = ~\new_[7166]_  | (~\new_[9363]_  & ~\new_[7532]_ );
  assign n6486 = ~\new_[6953]_  | (~\new_[10493]_  & ~\new_[7589]_ );
  assign n6491 = ~\new_[6944]_  | (~\new_[9364]_  & ~\new_[7545]_ );
  assign n6496 = ~\new_[6858]_  | (~\new_[10478]_  & ~\new_[7584]_ );
  assign n6501 = ~\new_[6859]_  | (~\new_[10490]_  & ~\new_[7580]_ );
  assign n6506 = ~\new_[6939]_  | (~\new_[9365]_  & ~\new_[7545]_ );
  assign n5781 = ~\new_[6860]_  | (~\new_[10486]_  & ~\new_[7583]_ );
  assign n6511 = ~\new_[6861]_  | (~\new_[10485]_  & ~\new_[7583]_ );
  assign n6521 = ~\new_[6934]_  | (~\new_[9366]_  & ~\new_[7532]_ );
  assign n6516 = ~\new_[6862]_  | (~\new_[10484]_  & ~\new_[7583]_ );
  assign n5786 = ~\new_[6863]_  | (~\new_[10483]_  & ~\new_[7579]_ );
  assign n6531 = ~\new_[6932]_  | (~\new_[9904]_  & ~\new_[7533]_ );
  assign n6536 = ~\new_[6865]_  | (~\new_[10481]_  & ~\new_[7579]_ );
  assign n6541 = ~\new_[6867]_  | (~\new_[10079]_  & ~\new_[7533]_ );
  assign n6546 = ~\new_[6868]_  | (~\new_[10505]_  & ~\new_[7585]_ );
  assign n5761 = ~\new_[6869]_  | (~\new_[9907]_  & ~\new_[7545]_ );
  assign n6551 = ~\new_[6870]_  | (~\new_[10504]_  & ~\new_[7585]_ );
  assign n6556 = ~\new_[6871]_  | (~\new_[10500]_  & ~\new_[7579]_ );
  assign n6566 = ~\new_[6872]_  | (~\new_[9908]_  & ~\new_[7544]_ );
  assign n5756 = ~\new_[6873]_  | (~\new_[10497]_  & ~\new_[7580]_ );
  assign n6576 = ~\new_[6874]_  | (~\new_[10102]_  & ~\new_[7542]_ );
  assign n6581 = ~\new_[6876]_  | (~\new_[10503]_  & ~\new_[7582]_ );
  assign n6591 = ~\new_[7154]_  | (~\new_[10499]_  & ~\new_[7582]_ );
  assign n6596 = ~\new_[6878]_  | (~\new_[9912]_  & ~\new_[7543]_ );
  assign n6601 = ~\new_[7151]_  | (~\new_[10488]_  & ~\new_[7581]_ );
  assign n6606 = ~\new_[7258]_  | (~\new_[10131]_  & ~\new_[7532]_ );
  assign n8421 = ~\new_[6882]_  | (~\new_[10150]_  & ~\new_[7587]_ );
  assign n5731 = ~\new_[6880]_  | (~\new_[9947]_  & ~\new_[7542]_ );
  assign n6616 = ~\new_[6881]_  | (~\new_[10080]_  & ~\new_[7543]_ );
  assign n6621 = ~\new_[7257]_  | (~\new_[9914]_  & ~\new_[7532]_ );
  assign n6426 = ~\new_[6848]_  | (~\new_[9358]_  & ~\new_[7543]_ );
  assign n6626 = ~\new_[7049]_  | (~\new_[9959]_  & ~\new_[7544]_ );
  assign n5726 = ~\new_[6943]_  | (~\new_[9916]_  & ~\new_[7543]_ );
  assign n6636 = ~\new_[6885]_  | (~\new_[10107]_  & ~\new_[7533]_ );
  assign n5721 = ~\new_[6887]_  | (~\new_[9918]_  & ~\new_[7532]_ );
  assign n6646 = ~\new_[6888]_  | (~\new_[10086]_  & ~\new_[7542]_ );
  assign n6651 = ~\new_[6889]_  | (~\new_[9919]_  & ~\new_[7533]_ );
  assign n6656 = ~\new_[6891]_  | (~\new_[9920]_  & ~\new_[7545]_ );
  assign n5506 = ~\new_[6892]_  | (~\new_[9921]_  & ~\new_[7532]_ );
  assign n6661 = ~\new_[6893]_  | (~\new_[10038]_  & ~\new_[7544]_ );
  assign n6666 = ~\new_[6894]_  | (~\new_[9953]_  & ~\new_[7532]_ );
  assign n6671 = ~\new_[6895]_  | (~\new_[10036]_  & ~\new_[7532]_ );
  assign n6676 = ~\new_[6896]_  | (~\new_[10134]_  & ~\new_[7542]_ );
  assign n6681 = ~\new_[6897]_  | (~\new_[10103]_  & ~\new_[7543]_ );
  assign n6686 = ~\new_[6898]_  | (~\new_[9926]_  & ~\new_[7544]_ );
  assign n6691 = ~\new_[6899]_  | (~\new_[9927]_  & ~\new_[7545]_ );
  assign n5696 = ~\new_[6900]_  | (~\new_[9922]_  & ~\new_[7544]_ );
  assign n6696 = ~\new_[6901]_  | (~\new_[9928]_  & ~\new_[7545]_ );
  assign n6701 = ~\new_[6902]_  | (~\new_[9638]_  & ~\new_[7534]_ );
  assign n6706 = ~\new_[6903]_  | (~\new_[9624]_  & ~\new_[7534]_ );
  assign n5691 = ~\new_[6904]_  | (~\new_[9626]_  & ~\new_[7540]_ );
  assign n6711 = ~\new_[6905]_  | (~\new_[9608]_  & ~\new_[7537]_ );
  assign n6716 = ~\new_[6906]_  | (~\new_[9373]_  & ~\new_[7537]_ );
  assign n6721 = ~\new_[6907]_  | (~\new_[9542]_  & ~\new_[7536]_ );
  assign n5686 = ~\new_[6908]_  | (~\new_[9374]_  & ~\new_[7536]_ );
  assign n6726 = ~\new_[6909]_  | (~\new_[9375]_  & ~\new_[7536]_ );
  assign n6731 = ~\new_[6910]_  | (~\new_[9376]_  & ~\new_[7536]_ );
  assign n6736 = ~\new_[6911]_  | (~\new_[9587]_  & ~\new_[7541]_ );
  assign n5636 = ~\new_[6912]_  | (~\new_[9377]_  & ~\new_[7541]_ );
  assign n6741 = ~\new_[6913]_  | (~\new_[9378]_  & ~\new_[7538]_ );
  assign n6751 = ~\new_[6915]_  | (~\new_[9539]_  & ~\new_[7538]_ );
  assign n5616 = ~\new_[6916]_  | (~\new_[9412]_  & ~\new_[7539]_ );
  assign n6756 = ~\new_[6942]_  | (~\new_[9379]_  & ~\new_[7539]_ );
  assign n6761 = ~\new_[6940]_  | (~\new_[9390]_  & ~\new_[7538]_ );
  assign n6766 = ~\new_[6918]_  | (~\new_[9381]_  & ~\new_[7538]_ );
  assign n5626 = ~\new_[6919]_  | (~\new_[9387]_  & ~\new_[7539]_ );
  assign n5766 = ~\new_[6923]_  | (~\new_[10479]_  & ~\new_[7589]_ );
  assign n6771 = ~\new_[6920]_  | (~\new_[9370]_  & ~\new_[7539]_ );
  assign n6776 = ~\new_[6922]_  | (~\new_[9438]_  & ~\new_[7537]_ );
  assign n6781 = ~\new_[6921]_  | (~\new_[9383]_  & ~\new_[7537]_ );
  assign n5621 = ~\new_[7357]_  | (~\new_[9380]_  & ~\new_[7541]_ );
  assign n6786 = ~\new_[6924]_  | (~\new_[9544]_  & ~\new_[7541]_ );
  assign n6791 = ~\new_[6945]_  | (~\new_[9543]_  & ~\new_[7535]_ );
  assign n6796 = ~\new_[6938]_  | (~\new_[9385]_  & ~\new_[7535]_ );
  assign n8511 = ~\new_[7401]_  | (~\new_[9634]_  & ~\new_[7532]_ );
  assign n5611 = ~\new_[6928]_  | (~\new_[9389]_  & ~\new_[7535]_ );
  assign n6801 = ~\new_[6929]_  | (~\new_[9386]_  & ~\new_[7535]_ );
  assign n7936 = ~\new_[6930]_  | (~\new_[9589]_  & ~\new_[7534]_ );
  assign n6806 = ~\new_[7153]_  | (~\new_[9384]_  & ~\new_[7534]_ );
  assign n8411 = ~\new_[7384]_  | (~\new_[9913]_  & ~\new_[7589]_ );
  assign n6526 = ~\new_[6864]_  | (~\new_[10491]_  & ~\new_[7584]_ );
  assign n9406 = ~\new_[7418]_  | (~\new_[9948]_  & ~\new_[7590]_ );
  assign n6811 = ~\new_[6917]_  | (~\new_[9537]_  & ~\new_[7540]_ );
  assign n8601 = ~\new_[7417]_  | (~\new_[9642]_  & ~\new_[7543]_ );
  assign n6631 = ~\new_[6937]_  | (~\new_[10082]_  & ~\new_[7544]_ );
  assign n6816 = ~\new_[6946]_  | (~\new_[9960]_  & ~\new_[7551]_ );
  assign n6821 = ~\new_[6947]_  | (~\new_[10048]_  & ~\new_[7549]_ );
  assign n6826 = ~\new_[6948]_  | (~\new_[9961]_  & ~\new_[7551]_ );
  assign n5591 = ~\new_[6949]_  | (~\new_[9962]_  & ~\new_[7547]_ );
  assign n6831 = ~\new_[6950]_  | (~\new_[9963]_  & ~\new_[7551]_ );
  assign n6836 = ~\new_[6951]_  | (~\new_[9965]_  & ~\new_[7551]_ );
  assign n6841 = ~\new_[6952]_  | (~\new_[9967]_  & ~\new_[7549]_ );
  assign n5571 = ~\new_[6954]_  | (~\new_[9958]_  & ~\new_[7551]_ );
  assign n6846 = ~\new_[6955]_  | (~\new_[9968]_  & ~\new_[7551]_ );
  assign n6851 = ~\new_[6956]_  | (~\new_[9969]_  & ~\new_[7547]_ );
  assign n6856 = ~\new_[6957]_  | (~\new_[9970]_  & ~\new_[7547]_ );
  assign n6861 = ~\new_[6958]_  | (~\new_[9971]_  & ~\new_[7551]_ );
  assign n6866 = ~\new_[6959]_  | (~\new_[9972]_  & ~\new_[7550]_ );
  assign n6871 = ~\new_[6960]_  | (~\new_[9973]_  & ~\new_[7551]_ );
  assign n6876 = ~\new_[6961]_  | (~\new_[9974]_  & ~\new_[7549]_ );
  assign n5566 = ~\new_[6962]_  | (~\new_[9976]_  & ~\new_[7549]_ );
  assign n6881 = ~\new_[6963]_  | (~\new_[9955]_  & ~\new_[7549]_ );
  assign n6886 = ~\new_[6964]_  | (~\new_[9977]_  & ~\new_[7553]_ );
  assign n6891 = ~\new_[6965]_  | (~\new_[9978]_  & ~\new_[7551]_ );
  assign n5546 = ~\new_[6966]_  | (~\new_[9979]_  & ~\new_[7546]_ );
  assign n6896 = ~\new_[6967]_  | (~\new_[9930]_  & ~\new_[7553]_ );
  assign n6901 = ~\new_[6968]_  | (~\new_[9925]_  & ~\new_[7546]_ );
  assign n6906 = ~\new_[6969]_  | (~\new_[9981]_  & ~\new_[7551]_ );
  assign n5531 = ~\new_[6970]_  | (~\new_[9982]_  & ~\new_[7550]_ );
  assign n6911 = ~\new_[6971]_  | (~\new_[9983]_  & ~\new_[7551]_ );
  assign n6916 = ~\new_[6972]_  | (~\new_[9984]_  & ~\new_[7551]_ );
  assign n6921 = ~\new_[6973]_  | (~\new_[9985]_  & ~\new_[7548]_ );
  assign n5541 = ~\new_[6974]_  | (~\new_[9986]_  & ~\new_[7548]_ );
  assign n6926 = ~\new_[6975]_  | (~\new_[10130]_  & ~\new_[7551]_ );
  assign n6931 = ~\new_[6976]_  | (~\new_[9987]_  & ~\new_[7553]_ );
  assign n6936 = ~\new_[6977]_  | (~\new_[9988]_  & ~\new_[7551]_ );
  assign n5536 = ~\new_[6978]_  | (~\new_[10132]_  & ~\new_[7549]_ );
  assign n6941 = ~\new_[6979]_  | (~\new_[9990]_  & ~\new_[7551]_ );
  assign n6946 = ~\new_[6980]_  | (~\new_[9991]_  & ~\new_[7549]_ );
  assign n6951 = ~\new_[6981]_  | (~\new_[9992]_  & ~\new_[7553]_ );
  assign n5526 = ~\new_[6982]_  | (~\new_[10117]_  & ~\new_[7553]_ );
  assign n6956 = ~\new_[6983]_  | (~\new_[9993]_  & ~\new_[7549]_ );
  assign n6961 = ~\new_[6984]_  | (~\new_[9994]_  & ~\new_[7551]_ );
  assign n6966 = ~\new_[6985]_  | (~\new_[9995]_  & ~\new_[7553]_ );
  assign n5356 = ~\new_[6986]_  | (~\new_[9997]_  & ~\new_[7551]_ );
  assign n6971 = ~\new_[6987]_  | (~\new_[9998]_  & ~\new_[7551]_ );
  assign n6976 = ~\new_[6988]_  | (~\new_[9999]_  & ~\new_[7551]_ );
  assign n6981 = ~\new_[6989]_  | (~\new_[10000]_  & ~\new_[7546]_ );
  assign n6986 = ~\new_[6990]_  | (~\new_[10001]_  & ~\new_[7551]_ );
  assign n6991 = ~\new_[6991]_  | (~\new_[10100]_  & ~\new_[7553]_ );
  assign n6996 = ~\new_[6992]_  | (~\new_[10002]_  & ~\new_[7546]_ );
  assign n7001 = ~\new_[6993]_  | (~\new_[10003]_  & ~\new_[7547]_ );
  assign n5496 = ~\new_[6994]_  | (~\new_[10004]_  & ~\new_[7551]_ );
  assign n7006 = ~\new_[6995]_  | (~\new_[10005]_  & ~\new_[7551]_ );
  assign n7011 = ~\new_[6996]_  | (~\new_[10007]_  & ~\new_[7551]_ );
  assign n7016 = ~\new_[6997]_  | (~\new_[10008]_  & ~\new_[7550]_ );
  assign n5491 = ~\new_[6998]_  | (~\new_[10009]_  & ~\new_[7551]_ );
  assign n7021 = ~\new_[6999]_  | (~\new_[10010]_  & ~\new_[7551]_ );
  assign n7026 = ~\new_[7000]_  | (~\new_[10011]_  & ~\new_[7551]_ );
  assign n7031 = ~\new_[7001]_  | (~\new_[10012]_  & ~\new_[7551]_ );
  assign n5486 = ~\new_[7002]_  | (~\new_[10013]_  & ~\new_[7548]_ );
  assign n7036 = ~\new_[7003]_  | (~\new_[10014]_  & ~\new_[7550]_ );
  assign n7041 = ~\new_[7004]_  | (~\new_[10016]_  & ~\new_[7548]_ );
  assign n7046 = ~\new_[7005]_  | (~\new_[10017]_  & ~\new_[7551]_ );
  assign n5476 = ~\new_[7006]_  | (~\new_[10019]_  & ~\new_[7551]_ );
  assign n7051 = ~\new_[7007]_  | (~\new_[10020]_  & ~\new_[7551]_ );
  assign n7056 = ~\new_[7008]_  | (~\new_[10021]_  & ~\new_[7551]_ );
  assign n7061 = ~\new_[7009]_  | (~\new_[10022]_  & ~\new_[7551]_ );
  assign n5461 = ~\new_[7010]_  | (~\new_[10023]_  & ~\new_[7553]_ );
  assign n7066 = ~\new_[7011]_  | (~\new_[9395]_  & ~\new_[7553]_ );
  assign n7071 = ~\new_[7012]_  | (~\new_[9401]_  & ~\new_[7553]_ );
  assign n7076 = ~\new_[7013]_  | (~\new_[9402]_  & ~\new_[7553]_ );
  assign n5471 = ~\new_[7015]_  | (~\new_[9403]_  & ~\new_[7553]_ );
  assign n7081 = ~\new_[7016]_  | (~\new_[9404]_  & ~\new_[7549]_ );
  assign n7086 = ~\new_[7017]_  | (~\new_[9406]_  & ~\new_[7549]_ );
  assign n9516 = n9796 ? \new_[8805]_  : \new_[5853]_ ;
  assign n9521 = n9796 ? \new_[8996]_  : \new_[5854]_ ;
  assign n9531 = n9796 ? \new_[9002]_  : \new_[5856]_ ;
  assign n9526 = n9796 ? \new_[9000]_  : \new_[5855]_ ;
  assign n9641 = n9796 ? \new_[9001]_  : \new_[5888]_ ;
  assign n9431 = \new_[5777]_  ? \new_[7608]_  : \new_[10542]_ ;
  assign n9536 = \new_[5857]_  ? \new_[7608]_  : \new_[10538]_ ;
  assign n9626 = \new_[5875]_  ? \new_[7608]_  : \new_[10699]_ ;
  assign n9541 = \new_[5858]_  ? \new_[7608]_  : \new_[10638]_ ;
  assign \new_[6759]_  = ~u14_u6_en_out_l2_reg;
  assign \new_[6760]_  = ~\new_[4689]_  & ~\new_[7616]_ ;
  assign n9556 = ~\new_[8150]_  | ~\new_[7466]_ ;
  assign n9451 = ~\new_[8172]_  | ~\new_[7480]_ ;
  assign n9576 = ~\new_[8151]_  | ~\new_[7467]_ ;
  assign n9571 = ~\new_[8170]_  | ~\new_[7468]_ ;
  assign \new_[6765]_  = ~\new_[13161]_  & ~\new_[7609]_ ;
  assign n9566 = ~\new_[8171]_  | ~\new_[7478]_ ;
  assign n9561 = ~\new_[8152]_  | ~\new_[7479]_ ;
  assign n9591 = ~\new_[8153]_  | ~\new_[7469]_ ;
  assign n9611 = ~\new_[8112]_  | ~\new_[7470]_ ;
  assign n9601 = ~\new_[8160]_  | ~\new_[7471]_ ;
  assign n9441 = ~\new_[8162]_  | ~\new_[7472]_ ;
  assign n9596 = ~\new_[8163]_  | ~\new_[7473]_ ;
  assign n9446 = ~\new_[8470]_  | ~\new_[7474]_ ;
  assign n9586 = ~\new_[8165]_  | ~\new_[7475]_ ;
  assign n9606 = ~\new_[8166]_  | ~\new_[7476]_ ;
  assign n9581 = ~\new_[8167]_  | ~\new_[7477]_ ;
  assign \new_[6777]_  = ~\new_[13124]_  & ~\new_[7610]_ ;
  assign \new_[6778]_  = ~\new_[13083]_  & ~\new_[7612]_ ;
  assign \new_[6779]_  = ~\new_[13158]_  & ~\new_[7605]_ ;
  assign \new_[6780]_  = ~\new_[13092]_  & ~\new_[7614]_ ;
  assign n9546 = \new_[8803]_  ? \new_[7595]_  : \new_[5859]_ ;
  assign n9551 = \new_[8503]_  ? \new_[7596]_  : \new_[5860]_ ;
  assign n9636 = \new_[13715]_  ? \new_[7937]_  : \new_[7594]_ ;
  assign n9436 = ~\new_[7420]_ ;
  assign \new_[6785]_  = ~\new_[7421]_ ;
  assign \new_[6786]_  = ~\new_[7422]_ ;
  assign \new_[6787]_  = ~\new_[7423]_ ;
  assign \new_[6788]_  = ~\new_[7424]_ ;
  assign \new_[6789]_  = ~\new_[7425]_ ;
  assign \wb_data_o[31]  = \\u12_wb_data_o_reg[31] ;
  assign \new_[6791]_  = \\u1_slt3_reg[6] ;
  assign \new_[6792]_  = \\u1_slt1_reg[6] ;
  assign \new_[6793]_  = \\u1_slt2_reg[6] ;
  assign \new_[6794]_  = \\u1_slt4_reg[6] ;
  assign \wb_data_o[23]  = \\u12_wb_data_o_reg[23] ;
  assign \wb_data_o[22]  = \\u12_wb_data_o_reg[22] ;
  assign \wb_data_o[21]  = \\u12_wb_data_o_reg[21] ;
  assign \wb_data_o[16]  = \\u12_wb_data_o_reg[16] ;
  assign \wb_data_o[20]  = \\u12_wb_data_o_reg[20] ;
  assign \wb_data_o[19]  = \\u12_wb_data_o_reg[19] ;
  assign \wb_data_o[17]  = \\u12_wb_data_o_reg[17] ;
  assign \wb_data_o[24]  = \\u12_wb_data_o_reg[24] ;
  assign \wb_data_o[30]  = \\u12_wb_data_o_reg[30] ;
  assign \wb_data_o[28]  = \\u12_wb_data_o_reg[28] ;
  assign \wb_data_o[27]  = \\u12_wb_data_o_reg[27] ;
  assign \wb_data_o[26]  = \\u12_wb_data_o_reg[26] ;
  assign \wb_data_o[29]  = \\u12_wb_data_o_reg[29] ;
  assign \wb_data_o[25]  = \\u12_wb_data_o_reg[25] ;
  assign \new_[6809]_  = \\u1_slt6_reg[6] ;
  assign \new_[6810]_  = ~\new_[13018]_  | (~\new_[9082]_  & ~\new_[7513]_ );
  assign \wb_data_o[18]  = \\u12_wb_data_o_reg[18] ;
  assign \new_[6812]_  = ~\new_[12872]_  & (~\new_[7514]_  | ~\new_[13007]_ );
  assign n9461 = \new_[13166]_  ? \new_[7512]_  : \new_[12686]_ ;
  assign n9466 = \new_[13162]_  ? \new_[7512]_  : \new_[5843]_ ;
  assign n9426 = \new_[13111]_  ? \new_[7512]_  : \new_[5767]_ ;
  assign n9471 = \new_[13090]_  ? \new_[7512]_  : \new_[5844]_ ;
  assign n9476 = \new_[13122]_  ? \new_[7512]_  : \new_[5845]_ ;
  assign n9481 = \new_[13187]_  ? \new_[7512]_  : \new_[13126]_ ;
  assign n9621 = \new_[13133]_  ? \new_[7512]_  : \new_[5874]_ ;
  assign n9486 = \new_[13189]_  ? \new_[7512]_  : \new_[5847]_ ;
  assign n9491 = \new_[13177]_  ? \new_[7512]_  : \new_[13110]_ ;
  assign n9496 = \new_[13183]_  ? \new_[7512]_  : \new_[13082]_ ;
  assign n9631 = \new_[13087]_  ? \new_[7512]_  : \new_[5876]_ ;
  assign n9501 = \new_[13172]_  ? \new_[7512]_  : \new_[5850]_ ;
  assign n9506 = \new_[13163]_  ? \new_[7512]_  : \new_[13137]_ ;
  assign n9511 = \new_[13086]_  ? \new_[7512]_  : \new_[5852]_ ;
  assign n9456 = \new_[13184]_  ? \new_[7512]_  : \new_[12519]_ ;
  assign n9616 = \new_[13179]_  ? \new_[7512]_  : \new_[5873]_ ;
  assign \new_[6829]_  = ~\new_[7431]_ ;
  assign \new_[6830]_  = ~u4_empty_reg;
  assign \new_[6831]_  = ~\new_[7432]_ ;
  assign \new_[6832]_  = ~u6_empty_reg;
  assign \new_[6833]_  = ~\new_[7433]_ ;
  assign \new_[6834]_  = ~\new_[7434]_ ;
  assign \new_[6835]_  = u15_crac_we_r_reg;
  assign \new_[6836]_  = ~\new_[7616]_  | ~\new_[12519]_  | ~\new_[4763]_ ;
  assign \new_[6837]_  = ~\new_[7533]_  | ~\new_[13012]_  | ~\new_[13127]_ ;
  assign \new_[6838]_  = ~\new_[7610]_  | ~\new_[12886]_  | ~\new_[13144]_ ;
  assign \new_[6839]_  = ~\new_[7612]_  | ~\new_[12691]_  | ~\new_[13175]_ ;
  assign \new_[6840]_  = ~\new_[7605]_  | ~\new_[12993]_  | ~\new_[13169]_ ;
  assign \new_[6841]_  = ~\new_[7614]_  | ~\new_[12686]_  | ~\new_[13105]_ ;
  assign n9666 = \\u1_sr_reg[8] ;
  assign \new_[6843]_  = ~\new_[5137]_  | ~\new_[7616]_ ;
  assign \new_[6844]_  = ~\new_[5138]_  | ~\new_[7533]_ ;
  assign \new_[6845]_  = ~\new_[5139]_  | ~\new_[7616]_ ;
  assign \new_[6846]_  = ~\new_[5025]_  | ~\new_[7533]_ ;
  assign \new_[6847]_  = ~\new_[5141]_  | ~\new_[7616]_ ;
  assign \new_[6848]_  = ~\new_[5143]_  | ~\new_[7533]_ ;
  assign \new_[6849]_  = ~\new_[5144]_  | ~\new_[7616]_ ;
  assign \new_[6850]_  = ~\new_[5016]_  | ~\new_[7533]_ ;
  assign \new_[6851]_  = ~\new_[5147]_  | ~\new_[7616]_ ;
  assign \new_[6852]_  = ~\new_[5149]_  | ~\new_[7616]_ ;
  assign \new_[6853]_  = ~\new_[5017]_  | ~\new_[7616]_ ;
  assign \new_[6854]_  = ~\new_[5152]_  | ~\new_[7533]_ ;
  assign \new_[6855]_  = ~\new_[5151]_  | ~\new_[7616]_ ;
  assign \new_[6856]_  = ~\new_[5015]_  | ~\new_[7616]_ ;
  assign \new_[6857]_  = ~\new_[5153]_  | ~\new_[7616]_ ;
  assign \new_[6858]_  = ~\new_[5157]_  | ~\new_[7616]_ ;
  assign \new_[6859]_  = ~\new_[5158]_  | ~\new_[7616]_ ;
  assign \new_[6860]_  = ~\new_[5010]_  | ~\new_[7616]_ ;
  assign \new_[6861]_  = ~\new_[5160]_  | ~\new_[7616]_ ;
  assign \new_[6862]_  = ~\new_[5161]_  | ~\new_[7616]_ ;
  assign \new_[6863]_  = ~\new_[5011]_  | ~\new_[7616]_ ;
  assign \new_[6864]_  = ~\new_[5163]_  | ~\new_[7616]_ ;
  assign \new_[6865]_  = ~\new_[5165]_  | ~\new_[7616]_ ;
  assign \new_[6866]_  = ~\new_[5024]_  | ~\new_[7614]_ ;
  assign \new_[6867]_  = ~\new_[5166]_  | ~\new_[7609]_ ;
  assign \new_[6868]_  = ~\new_[5167]_  | ~\new_[7616]_ ;
  assign \new_[6869]_  = ~\new_[5006]_  | ~\new_[7609]_ ;
  assign \new_[6870]_  = ~\new_[5168]_  | ~\new_[7616]_ ;
  assign \new_[6871]_  = ~\new_[5169]_  | ~\new_[7616]_ ;
  assign \new_[6872]_  = ~\new_[5171]_  | ~\new_[7533]_ ;
  assign \new_[6873]_  = ~\new_[5005]_  | ~\new_[7616]_ ;
  assign \new_[6874]_  = ~\new_[5173]_  | ~\new_[7533]_ ;
  assign \new_[6875]_  = ~\new_[5172]_  | ~\new_[7616]_ ;
  assign \new_[6876]_  = ~\new_[5174]_  | ~\new_[7616]_ ;
  assign \new_[6877]_  = ~\new_[5175]_  | ~\new_[7609]_ ;
  assign \new_[6878]_  = ~\new_[5177]_  | ~\new_[7533]_ ;
  assign \new_[6879]_  = ~\new_[5001]_  | ~\new_[7616]_ ;
  assign \new_[6880]_  = ~\new_[5000]_  | ~\new_[7533]_ ;
  assign \new_[6881]_  = ~\new_[5181]_  | ~\new_[7609]_ ;
  assign \new_[6882]_  = ~\new_[5542]_  | ~\new_[7616]_ ;
  assign \new_[6883]_  = ~\new_[4919]_  | ~\new_[7616]_ ;
  assign \new_[6884]_  = ~\new_[4948]_  | ~\new_[7616]_ ;
  assign \new_[6885]_  = ~\new_[5185]_  | ~\new_[7533]_ ;
  assign \new_[6886]_  = ~\new_[5186]_  | ~\new_[7609]_ ;
  assign \new_[6887]_  = ~\new_[4998]_  | ~\new_[7533]_ ;
  assign \new_[6888]_  = ~\new_[5187]_  | ~\new_[7609]_ ;
  assign \new_[6889]_  = ~\new_[5188]_  | ~\new_[7609]_ ;
  assign \new_[6890]_  = ~\new_[5142]_  | ~\new_[7616]_ ;
  assign \new_[6891]_  = ~\new_[5189]_  | ~\new_[7609]_ ;
  assign \new_[6892]_  = ~\new_[4942]_  | ~\new_[7533]_ ;
  assign \new_[6893]_  = ~\new_[5190]_  | ~\new_[7609]_ ;
  assign \new_[6894]_  = ~\new_[5191]_  | ~\new_[7533]_ ;
  assign \new_[6895]_  = ~\new_[5192]_  | ~\new_[7533]_ ;
  assign \new_[6896]_  = ~\new_[5193]_  | ~\new_[7609]_ ;
  assign \new_[6897]_  = ~\new_[5194]_  | ~\new_[7609]_ ;
  assign \new_[6898]_  = ~\new_[5195]_  | ~\new_[7533]_ ;
  assign \new_[6899]_  = ~\new_[5196]_  | ~\new_[7533]_ ;
  assign \new_[6900]_  = ~\new_[4993]_  | ~\new_[7609]_ ;
  assign \new_[6901]_  = ~\new_[5197]_  | ~\new_[7533]_ ;
  assign \new_[6902]_  = ~\new_[5198]_  | ~\new_[7533]_ ;
  assign \new_[6903]_  = ~\new_[5199]_  | ~\new_[7533]_ ;
  assign \new_[6904]_  = ~\new_[4992]_  | ~\new_[7533]_ ;
  assign \new_[6905]_  = ~\new_[5200]_  | ~\new_[7532]_ ;
  assign \new_[6906]_  = ~\new_[5201]_  | ~\new_[7532]_ ;
  assign \new_[6907]_  = ~\new_[5202]_  | ~\new_[7533]_ ;
  assign \new_[6908]_  = ~\new_[4991]_  | ~\new_[7533]_ ;
  assign \new_[6909]_  = ~\new_[5203]_  | ~\new_[7532]_ ;
  assign \new_[6910]_  = ~\new_[5204]_  | ~\new_[7532]_ ;
  assign \new_[6911]_  = ~\new_[5205]_  | ~\new_[7533]_ ;
  assign \new_[6912]_  = ~\new_[4979]_  | ~\new_[7533]_ ;
  assign \new_[6913]_  = ~\new_[5206]_  | ~\new_[7533]_ ;
  assign \new_[6914]_  = ~\new_[5207]_  | ~\new_[7533]_ ;
  assign \new_[6915]_  = ~\new_[5208]_  | ~\new_[7533]_ ;
  assign \new_[6916]_  = ~\new_[4975]_  | ~\new_[7533]_ ;
  assign \new_[6917]_  = ~\new_[5220]_  | ~\new_[7533]_ ;
  assign \new_[6918]_  = ~\new_[5211]_  | ~\new_[7609]_ ;
  assign \new_[6919]_  = ~\new_[4977]_  | ~\new_[7609]_ ;
  assign \new_[6920]_  = ~\new_[5212]_  | ~\new_[7533]_ ;
  assign \new_[6921]_  = ~\new_[5214]_  | ~\new_[7609]_ ;
  assign \new_[6922]_  = ~\new_[5213]_  | ~\new_[7533]_ ;
  assign \new_[6923]_  = ~\new_[5007]_  | ~\new_[7616]_ ;
  assign \new_[6924]_  = ~\new_[5215]_  | ~\new_[7609]_ ;
  assign \new_[6925]_  = ~\new_[5479]_  | ~\new_[7614]_ ;
  assign \new_[6926]_  = ~\new_[4969]_  | ~\new_[7533]_ ;
  assign \new_[6927]_  = ~\new_[5559]_  | ~\new_[7616]_ ;
  assign \new_[6928]_  = ~\new_[4974]_  | ~\new_[7609]_ ;
  assign \new_[6929]_  = ~\new_[5218]_  | ~\new_[7609]_ ;
  assign \new_[6930]_  = ~\new_[5445]_  | ~\new_[7609]_ ;
  assign \new_[6931]_  = ~\new_[5140]_  | ~\new_[7616]_ ;
  assign \new_[6932]_  = ~\new_[5164]_  | ~\new_[7533]_ ;
  assign \new_[6933]_  = ~\new_[5032]_  | ~\new_[7616]_ ;
  assign \new_[6934]_  = ~\new_[5162]_  | ~\new_[7533]_ ;
  assign \new_[6935]_  = ~\new_[5136]_  | ~\new_[7533]_ ;
  assign \new_[6936]_  = ~\new_[5135]_  | ~\new_[7616]_ ;
  assign \new_[6937]_  = ~\new_[5184]_  | ~\new_[7533]_ ;
  assign \new_[6938]_  = ~\new_[5217]_  | ~\new_[7609]_ ;
  assign \new_[6939]_  = ~\new_[5159]_  | ~\new_[7609]_ ;
  assign \new_[6940]_  = ~\new_[5210]_  | ~\new_[7532]_ ;
  assign \new_[6941]_  = ~\new_[5577]_  | ~\new_[7616]_ ;
  assign \new_[6942]_  = ~\new_[5209]_  | ~\new_[7532]_ ;
  assign \new_[6943]_  = ~\new_[4999]_  | ~\new_[7533]_ ;
  assign \new_[6944]_  = ~\new_[5156]_  | ~\new_[7609]_ ;
  assign \new_[6945]_  = ~\new_[5216]_  | ~\new_[7533]_ ;
  assign \new_[6946]_  = ~\new_[5221]_  | ~\new_[7610]_ ;
  assign \new_[6947]_  = ~\new_[5222]_  | ~\new_[7610]_ ;
  assign \new_[6948]_  = ~\new_[5223]_  | ~\new_[7610]_ ;
  assign \new_[6949]_  = ~\new_[4970]_  | ~\new_[7610]_ ;
  assign \new_[6950]_  = ~\new_[5224]_  | ~\new_[7610]_ ;
  assign \new_[6951]_  = ~\new_[5225]_  | ~\new_[7610]_ ;
  assign \new_[6952]_  = ~\new_[5226]_  | ~\new_[7610]_ ;
  assign \new_[6953]_  = ~\new_[5155]_  | ~\new_[7616]_ ;
  assign \new_[6954]_  = ~\new_[4966]_  | ~\new_[7610]_ ;
  assign \new_[6955]_  = ~\new_[5227]_  | ~\new_[7610]_ ;
  assign \new_[6956]_  = ~\new_[5228]_  | ~\new_[7610]_ ;
  assign \new_[6957]_  = ~\new_[5229]_  | ~\new_[7610]_ ;
  assign \new_[6958]_  = ~\new_[5230]_  | ~\new_[7610]_ ;
  assign \new_[6959]_  = ~\new_[5231]_  | ~\new_[7610]_ ;
  assign \new_[6960]_  = ~\new_[5232]_  | ~\new_[7610]_ ;
  assign \new_[6961]_  = ~\new_[5233]_  | ~\new_[7610]_ ;
  assign \new_[6962]_  = ~\new_[4965]_  | ~\new_[7610]_ ;
  assign \new_[6963]_  = ~\new_[5234]_  | ~\new_[7610]_ ;
  assign \new_[6964]_  = ~\new_[5235]_  | ~\new_[7610]_ ;
  assign \new_[6965]_  = ~\new_[5236]_  | ~\new_[7610]_ ;
  assign \new_[6966]_  = ~\new_[4961]_  | ~\new_[7610]_ ;
  assign \new_[6967]_  = ~\new_[5237]_  | ~\new_[7610]_ ;
  assign \new_[6968]_  = ~\new_[5238]_  | ~\new_[7610]_ ;
  assign \new_[6969]_  = ~\new_[5239]_  | ~\new_[7610]_ ;
  assign \new_[6970]_  = ~\new_[4952]_  | ~\new_[7610]_ ;
  assign \new_[6971]_  = ~\new_[5240]_  | ~\new_[7610]_ ;
  assign \new_[6972]_  = ~\new_[5241]_  | ~\new_[7610]_ ;
  assign \new_[6973]_  = ~\new_[5242]_  | ~\new_[7610]_ ;
  assign \new_[6974]_  = ~\new_[4954]_  | ~\new_[7610]_ ;
  assign \new_[6975]_  = ~\new_[5243]_  | ~\new_[7610]_ ;
  assign \new_[6976]_  = ~\new_[5244]_  | ~\new_[7610]_ ;
  assign \new_[6977]_  = ~\new_[5245]_  | ~\new_[7610]_ ;
  assign \new_[6978]_  = ~\new_[4953]_  | ~\new_[7610]_ ;
  assign \new_[6979]_  = ~\new_[5246]_  | ~\new_[7610]_ ;
  assign \new_[6980]_  = ~\new_[5247]_  | ~\new_[7610]_ ;
  assign \new_[6981]_  = ~\new_[5248]_  | ~\new_[7610]_ ;
  assign \new_[6982]_  = ~\new_[4951]_  | ~\new_[7610]_ ;
  assign \new_[6983]_  = ~\new_[5249]_  | ~\new_[7610]_ ;
  assign \new_[6984]_  = ~\new_[5250]_  | ~\new_[7610]_ ;
  assign \new_[6985]_  = ~\new_[5251]_  | ~\new_[7610]_ ;
  assign \new_[6986]_  = ~\new_[4900]_  | ~\new_[7610]_ ;
  assign \new_[6987]_  = ~\new_[5252]_  | ~\new_[7610]_ ;
  assign \new_[6988]_  = ~\new_[5253]_  | ~\new_[7610]_ ;
  assign \new_[6989]_  = ~\new_[5254]_  | ~\new_[7610]_ ;
  assign \new_[6990]_  = ~\new_[5255]_  | ~\new_[7610]_ ;
  assign \new_[6991]_  = ~\new_[5256]_  | ~\new_[7610]_ ;
  assign \new_[6992]_  = ~\new_[5257]_  | ~\new_[7610]_ ;
  assign \new_[6993]_  = ~\new_[5258]_  | ~\new_[7610]_ ;
  assign \new_[6994]_  = ~\new_[4938]_  | ~\new_[7610]_ ;
  assign \new_[6995]_  = ~\new_[5259]_  | ~\new_[7610]_ ;
  assign \new_[6996]_  = ~\new_[5260]_  | ~\new_[7610]_ ;
  assign \new_[6997]_  = ~\new_[5261]_  | ~\new_[7610]_ ;
  assign \new_[6998]_  = ~\new_[4937]_  | ~\new_[7610]_ ;
  assign \new_[6999]_  = ~\new_[5262]_  | ~\new_[7610]_ ;
  assign \new_[7000]_  = ~\new_[5263]_  | ~\new_[7610]_ ;
  assign \new_[7001]_  = ~\new_[5264]_  | ~\new_[7610]_ ;
  assign \new_[7002]_  = ~\new_[4936]_  | ~\new_[7610]_ ;
  assign \new_[7003]_  = ~\new_[5265]_  | ~\new_[7610]_ ;
  assign \new_[7004]_  = ~\new_[5266]_  | ~\new_[7610]_ ;
  assign \new_[7005]_  = ~\new_[5267]_  | ~\new_[7610]_ ;
  assign \new_[7006]_  = ~\new_[4929]_  | ~\new_[7610]_ ;
  assign \new_[7007]_  = ~\new_[5268]_  | ~\new_[7610]_ ;
  assign \new_[7008]_  = ~\new_[5269]_  | ~\new_[7610]_ ;
  assign \new_[7009]_  = ~\new_[5270]_  | ~\new_[7610]_ ;
  assign \new_[7010]_  = ~\new_[4921]_  | ~\new_[7610]_ ;
  assign \new_[7011]_  = ~\new_[5271]_  | ~\new_[7610]_ ;
  assign \new_[7012]_  = ~\new_[5272]_  | ~\new_[7610]_ ;
  assign \new_[7013]_  = ~\new_[5273]_  | ~\new_[7610]_ ;
  assign \new_[7014]_  = ~\new_[5520]_  | ~\new_[7616]_ ;
  assign \new_[7015]_  = ~\new_[4923]_  | ~\new_[7610]_ ;
  assign \new_[7016]_  = ~\new_[5274]_  | ~\new_[7610]_ ;
  assign \new_[7017]_  = ~\new_[5275]_  | ~\new_[7610]_ ;
  assign \new_[7018]_  = ~\new_[5276]_  | ~\new_[7610]_ ;
  assign \new_[7019]_  = ~\new_[4899]_  | ~\new_[7616]_ ;
  assign \new_[7020]_  = ~\new_[4922]_  | ~\new_[7610]_ ;
  assign \new_[7021]_  = ~\new_[5277]_  | ~\new_[7610]_ ;
  assign \new_[7022]_  = ~\new_[5278]_  | ~\new_[7610]_ ;
  assign \new_[7023]_  = ~\new_[5279]_  | ~\new_[7610]_ ;
  assign \new_[7024]_  = ~\new_[5280]_  | ~\new_[7610]_ ;
  assign \new_[7025]_  = ~\new_[5281]_  | ~\new_[7610]_ ;
  assign \new_[7026]_  = ~\new_[5282]_  | ~\new_[7610]_ ;
  assign \new_[7027]_  = ~\new_[5283]_  | ~\new_[7610]_ ;
  assign \new_[7028]_  = ~\new_[4914]_  | ~\new_[7610]_ ;
  assign \new_[7029]_  = ~\new_[5284]_  | ~\new_[7610]_ ;
  assign \new_[7030]_  = ~\new_[5285]_  | ~\new_[7610]_ ;
  assign \new_[7031]_  = ~\new_[5286]_  | ~\new_[7610]_ ;
  assign \new_[7032]_  = ~\new_[4915]_  | ~\new_[7610]_ ;
  assign \new_[7033]_  = ~\new_[5287]_  | ~\new_[7610]_ ;
  assign \new_[7034]_  = ~\new_[5288]_  | ~\new_[7610]_ ;
  assign \new_[7035]_  = ~\new_[5289]_  | ~\new_[7610]_ ;
  assign \new_[7036]_  = ~\new_[4911]_  | ~\new_[7610]_ ;
  assign \new_[7037]_  = ~\new_[5290]_  | ~\new_[7610]_ ;
  assign \new_[7038]_  = ~\new_[4945]_  | ~\new_[7533]_ ;
  assign \new_[7039]_  = ~\new_[5291]_  | ~\new_[7610]_ ;
  assign \new_[7040]_  = ~\new_[5292]_  | ~\new_[7610]_ ;
  assign \new_[7041]_  = ~\new_[4910]_  | ~\new_[7610]_ ;
  assign \new_[7042]_  = ~\new_[5293]_  | ~\new_[7610]_ ;
  assign \new_[7043]_  = ~\new_[5294]_  | ~\new_[7610]_ ;
  assign \new_[7044]_  = ~\new_[5295]_  | ~\new_[7610]_ ;
  assign \new_[7045]_  = ~\new_[4909]_  | ~\new_[7610]_ ;
  assign \new_[7046]_  = ~\new_[5531]_  | ~\new_[7616]_ ;
  assign \new_[7047]_  = ~\new_[5522]_  | ~\new_[7616]_ ;
  assign \new_[7048]_  = ~\new_[5562]_  | ~\new_[7533]_ ;
  assign \new_[7049]_  = ~\new_[5183]_  | ~\new_[7533]_ ;
  assign \new_[7050]_  = ~\new_[5528]_  | ~\new_[7616]_ ;
  assign \new_[7051]_  = ~\new_[5297]_  | ~\new_[7612]_ ;
  assign \new_[7052]_  = ~\new_[5298]_  | ~\new_[7612]_ ;
  assign \new_[7053]_  = ~\new_[4906]_  | ~\new_[7612]_ ;
  assign \new_[7054]_  = ~\new_[5299]_  | ~\new_[7612]_ ;
  assign \new_[7055]_  = ~\new_[5300]_  | ~\new_[7612]_ ;
  assign \new_[7056]_  = ~\new_[5301]_  | ~\new_[7612]_ ;
  assign \new_[7057]_  = ~\new_[4904]_  | ~\new_[7612]_ ;
  assign \new_[7058]_  = ~\new_[5303]_  | ~\new_[7612]_ ;
  assign \new_[7059]_  = ~\new_[5304]_  | ~\new_[7612]_ ;
  assign \new_[7060]_  = ~\new_[5305]_  | ~\new_[7612]_ ;
  assign \new_[7061]_  = ~\new_[4905]_  | ~\new_[7612]_ ;
  assign \new_[7062]_  = ~\new_[5306]_  | ~\new_[7612]_ ;
  assign \new_[7063]_  = ~\new_[5307]_  | ~\new_[7612]_ ;
  assign \new_[7064]_  = ~\new_[5308]_  | ~\new_[7612]_ ;
  assign \new_[7065]_  = ~\new_[4903]_  | ~\new_[7612]_ ;
  assign \new_[7066]_  = ~\new_[5309]_  | ~\new_[7612]_ ;
  assign \new_[7067]_  = ~\new_[5310]_  | ~\new_[7612]_ ;
  assign \new_[7068]_  = ~\new_[5311]_  | ~\new_[7612]_ ;
  assign \new_[7069]_  = ~\new_[4901]_  | ~\new_[7612]_ ;
  assign \new_[7070]_  = ~\new_[5312]_  | ~\new_[7612]_ ;
  assign \new_[7071]_  = ~\new_[5313]_  | ~\new_[7612]_ ;
  assign \new_[7072]_  = ~\new_[5314]_  | ~\new_[7612]_ ;
  assign \new_[7073]_  = ~\new_[5757]_  | ~\new_[7612]_ ;
  assign \new_[7074]_  = ~\new_[5315]_  | ~\new_[7612]_ ;
  assign \new_[7075]_  = ~\new_[5316]_  | ~\new_[7612]_ ;
  assign \new_[7076]_  = ~\new_[5317]_  | ~\new_[7612]_ ;
  assign \new_[7077]_  = ~\new_[5765]_  | ~\new_[7612]_ ;
  assign \new_[7078]_  = ~\new_[5318]_  | ~\new_[7612]_ ;
  assign \new_[7079]_  = ~\new_[5319]_  | ~\new_[7612]_ ;
  assign \new_[7080]_  = ~\new_[5320]_  | ~\new_[7612]_ ;
  assign \new_[7081]_  = ~\new_[5764]_  | ~\new_[7612]_ ;
  assign \new_[7082]_  = ~\new_[5321]_  | ~\new_[7612]_ ;
  assign \new_[7083]_  = ~\new_[5465]_  | ~\new_[7614]_ ;
  assign \new_[7084]_  = ~\new_[5322]_  | ~\new_[7612]_ ;
  assign \new_[7085]_  = ~\new_[5323]_  | ~\new_[7612]_ ;
  assign \new_[7086]_  = ~\new_[5758]_  | ~\new_[7612]_ ;
  assign \new_[7087]_  = ~\new_[5324]_  | ~\new_[7612]_ ;
  assign \new_[7088]_  = ~\new_[5325]_  | ~\new_[7612]_ ;
  assign \new_[7089]_  = ~\new_[5326]_  | ~\new_[7612]_ ;
  assign \new_[7090]_  = ~\new_[5762]_  | ~\new_[7612]_ ;
  assign \new_[7091]_  = ~\new_[5327]_  | ~\new_[7612]_ ;
  assign \new_[7092]_  = ~\new_[5328]_  | ~\new_[7612]_ ;
  assign \new_[7093]_  = ~\new_[5329]_  | ~\new_[7612]_ ;
  assign \new_[7094]_  = ~\new_[5760]_  | ~\new_[7612]_ ;
  assign \new_[7095]_  = ~\new_[5330]_  | ~\new_[7612]_ ;
  assign \new_[7096]_  = ~\new_[5331]_  | ~\new_[7612]_ ;
  assign \new_[7097]_  = ~\new_[5332]_  | ~\new_[7612]_ ;
  assign \new_[7098]_  = ~\new_[5761]_  | ~\new_[7612]_ ;
  assign \new_[7099]_  = ~\new_[5333]_  | ~\new_[7612]_ ;
  assign \new_[7100]_  = ~\new_[5334]_  | ~\new_[7612]_ ;
  assign \new_[7101]_  = ~\new_[5335]_  | ~\new_[7612]_ ;
  assign \new_[7102]_  = ~\new_[5754]_  | ~\new_[7612]_ ;
  assign \new_[7103]_  = ~\new_[5336]_  | ~\new_[7612]_ ;
  assign \new_[7104]_  = ~\new_[5337]_  | ~\new_[7612]_ ;
  assign \new_[7105]_  = ~\new_[5338]_  | ~\new_[7612]_ ;
  assign \new_[7106]_  = ~\new_[5752]_  | ~\new_[7612]_ ;
  assign \new_[7107]_  = ~\new_[5339]_  | ~\new_[7612]_ ;
  assign \new_[7108]_  = ~\new_[5340]_  | ~\new_[7612]_ ;
  assign \new_[7109]_  = ~\new_[5341]_  | ~\new_[7612]_ ;
  assign \new_[7110]_  = ~\new_[5342]_  | ~\new_[7612]_ ;
  assign \new_[7111]_  = ~\new_[5343]_  | ~\new_[7612]_ ;
  assign \new_[7112]_  = ~\new_[5344]_  | ~\new_[7612]_ ;
  assign \new_[7113]_  = ~\new_[5345]_  | ~\new_[7612]_ ;
  assign \new_[7114]_  = ~\new_[5732]_  | ~\new_[7612]_ ;
  assign \new_[7115]_  = ~\new_[5346]_  | ~\new_[7612]_ ;
  assign \new_[7116]_  = ~\new_[5347]_  | ~\new_[7612]_ ;
  assign \new_[7117]_  = ~\new_[5348]_  | ~\new_[7612]_ ;
  assign \new_[7118]_  = ~\new_[5751]_  | ~\new_[7612]_ ;
  assign \new_[7119]_  = ~\new_[5349]_  | ~\new_[7612]_ ;
  assign \new_[7120]_  = ~\new_[5350]_  | ~\new_[7612]_ ;
  assign \new_[7121]_  = ~\new_[5351]_  | ~\new_[7612]_ ;
  assign \new_[7122]_  = ~\new_[5743]_  | ~\new_[7612]_ ;
  assign \new_[7123]_  = ~\new_[5352]_  | ~\new_[7612]_ ;
  assign \new_[7124]_  = ~\new_[5353]_  | ~\new_[7612]_ ;
  assign \new_[7125]_  = ~\new_[5354]_  | ~\new_[7612]_ ;
  assign \new_[7126]_  = ~\new_[5736]_  | ~\new_[7612]_ ;
  assign \new_[7127]_  = ~\new_[5355]_  | ~\new_[7612]_ ;
  assign \new_[7128]_  = ~\new_[5356]_  | ~\new_[7612]_ ;
  assign \new_[7129]_  = ~\new_[5357]_  | ~\new_[7612]_ ;
  assign \new_[7130]_  = ~\new_[5740]_  | ~\new_[7612]_ ;
  assign \new_[7131]_  = ~\new_[5359]_  | ~\new_[7612]_ ;
  assign \new_[7132]_  = ~\new_[5360]_  | ~\new_[7612]_ ;
  assign \new_[7133]_  = ~\new_[5361]_  | ~\new_[7612]_ ;
  assign \new_[7134]_  = ~\new_[5737]_  | ~\new_[7612]_ ;
  assign \new_[7135]_  = ~\new_[5362]_  | ~\new_[7612]_ ;
  assign \new_[7136]_  = ~\new_[5363]_  | ~\new_[7612]_ ;
  assign \new_[7137]_  = ~\new_[5364]_  | ~\new_[7612]_ ;
  assign \new_[7138]_  = ~\new_[5738]_  | ~\new_[7612]_ ;
  assign \new_[7139]_  = ~\new_[5365]_  | ~\new_[7612]_ ;
  assign \new_[7140]_  = ~\new_[5366]_  | ~\new_[7612]_ ;
  assign \new_[7141]_  = ~\new_[5367]_  | ~\new_[7612]_ ;
  assign \new_[7142]_  = ~\new_[5730]_  | ~\new_[7612]_ ;
  assign \new_[7143]_  = ~\new_[5368]_  | ~\new_[7612]_ ;
  assign \new_[7144]_  = ~\new_[5369]_  | ~\new_[7612]_ ;
  assign \new_[7145]_  = ~\new_[5370]_  | ~\new_[7612]_ ;
  assign \new_[7146]_  = ~\new_[5728]_  | ~\new_[7612]_ ;
  assign \new_[7147]_  = ~\new_[5371]_  | ~\new_[7612]_ ;
  assign \new_[7148]_  = ~\new_[5525]_  | ~\new_[7616]_ ;
  assign \new_[7149]_  = ~\new_[5018]_  | ~\new_[7616]_ ;
  assign \new_[7150]_  = ~\new_[5002]_  | ~\new_[7616]_ ;
  assign \new_[7151]_  = ~\new_[5178]_  | ~\new_[7616]_ ;
  assign \new_[7152]_  = ~\new_[5296]_  | ~\new_[7609]_ ;
  assign \new_[7153]_  = ~\new_[5219]_  | ~\new_[7533]_ ;
  assign \new_[7154]_  = ~\new_[5176]_  | ~\new_[7616]_ ;
  assign \new_[7155]_  = ~\new_[5372]_  | ~\new_[7605]_ ;
  assign \new_[7156]_  = ~\new_[5373]_  | ~\new_[7605]_ ;
  assign \new_[7157]_  = ~\new_[5729]_  | ~\new_[7605]_ ;
  assign \new_[7158]_  = ~\new_[5374]_  | ~\new_[7605]_ ;
  assign \new_[7159]_  = ~\new_[5375]_  | ~\new_[7605]_ ;
  assign \new_[7160]_  = ~\new_[5376]_  | ~\new_[7605]_ ;
  assign \new_[7161]_  = ~\new_[5705]_  | ~\new_[7605]_ ;
  assign \new_[7162]_  = ~\new_[5377]_  | ~\new_[7605]_ ;
  assign \new_[7163]_  = ~\new_[5378]_  | ~\new_[7605]_ ;
  assign \new_[7164]_  = ~\new_[5379]_  | ~\new_[7605]_ ;
  assign \new_[7165]_  = ~\new_[5380]_  | ~\new_[7605]_ ;
  assign \new_[7166]_  = ~\new_[5154]_  | ~\new_[7533]_ ;
  assign \new_[7167]_  = ~\new_[5381]_  | ~\new_[7605]_ ;
  assign \new_[7168]_  = ~\new_[5382]_  | ~\new_[7605]_ ;
  assign \new_[7169]_  = ~\new_[5383]_  | ~\new_[7605]_ ;
  assign \new_[7170]_  = ~\new_[5724]_  | ~\new_[7605]_ ;
  assign \new_[7171]_  = ~\new_[5384]_  | ~\new_[7605]_ ;
  assign \new_[7172]_  = ~\new_[5385]_  | ~\new_[7605]_ ;
  assign \new_[7173]_  = ~\new_[5386]_  | ~\new_[7605]_ ;
  assign \new_[7174]_  = ~\new_[5718]_  | ~\new_[7605]_ ;
  assign \new_[7175]_  = ~\new_[5387]_  | ~\new_[7605]_ ;
  assign \new_[7176]_  = ~\new_[5388]_  | ~\new_[7605]_ ;
  assign \new_[7177]_  = ~\new_[5552]_  | ~\new_[7616]_ ;
  assign \new_[7178]_  = ~\new_[5389]_  | ~\new_[7605]_ ;
  assign \new_[7179]_  = ~\new_[5722]_  | ~\new_[7605]_ ;
  assign \new_[7180]_  = ~\new_[5390]_  | ~\new_[7605]_ ;
  assign \new_[7181]_  = ~\new_[5391]_  | ~\new_[7605]_ ;
  assign \new_[7182]_  = ~\new_[5392]_  | ~\new_[7605]_ ;
  assign \new_[7183]_  = ~\new_[5720]_  | ~\new_[7605]_ ;
  assign \new_[7184]_  = ~\new_[5393]_  | ~\new_[7605]_ ;
  assign \new_[7185]_  = ~\new_[5394]_  | ~\new_[7605]_ ;
  assign \new_[7186]_  = ~\new_[5395]_  | ~\new_[7605]_ ;
  assign \new_[7187]_  = ~\new_[5721]_  | ~\new_[7605]_ ;
  assign \new_[7188]_  = ~\new_[5396]_  | ~\new_[7605]_ ;
  assign \new_[7189]_  = ~\new_[5397]_  | ~\new_[7605]_ ;
  assign \new_[7190]_  = ~\new_[5398]_  | ~\new_[7605]_ ;
  assign \new_[7191]_  = ~\new_[5553]_  | ~\new_[7533]_ ;
  assign \new_[7192]_  = ~\new_[5714]_  | ~\new_[7605]_ ;
  assign \new_[7193]_  = ~\new_[5399]_  | ~\new_[7605]_ ;
  assign \new_[7194]_  = ~\new_[5400]_  | ~\new_[7605]_ ;
  assign \new_[7195]_  = ~\new_[5401]_  | ~\new_[7605]_ ;
  assign \new_[7196]_  = ~\new_[5704]_  | ~\new_[7605]_ ;
  assign \new_[7197]_  = ~\new_[5402]_  | ~\new_[7605]_ ;
  assign \new_[7198]_  = ~\new_[5403]_  | ~\new_[7605]_ ;
  assign \new_[7199]_  = ~\new_[5404]_  | ~\new_[7605]_ ;
  assign \new_[7200]_  = ~\new_[5708]_  | ~\new_[7605]_ ;
  assign \new_[7201]_  = ~\new_[5405]_  | ~\new_[7605]_ ;
  assign \new_[7202]_  = ~\new_[5406]_  | ~\new_[7605]_ ;
  assign \new_[7203]_  = ~\new_[5407]_  | ~\new_[7605]_ ;
  assign \new_[7204]_  = ~\new_[5668]_  | ~\new_[7605]_ ;
  assign \new_[7205]_  = ~\new_[5408]_  | ~\new_[7605]_ ;
  assign \new_[7206]_  = ~\new_[5409]_  | ~\new_[7605]_ ;
  assign \new_[7207]_  = ~\new_[5410]_  | ~\new_[7605]_ ;
  assign \new_[7208]_  = ~\new_[5697]_  | ~\new_[7605]_ ;
  assign \new_[7209]_  = ~\new_[5411]_  | ~\new_[7605]_ ;
  assign \new_[7210]_  = ~\new_[5412]_  | ~\new_[7605]_ ;
  assign \new_[7211]_  = ~\new_[5413]_  | ~\new_[7605]_ ;
  assign \new_[7212]_  = ~\new_[5692]_  | ~\new_[7605]_ ;
  assign \new_[7213]_  = ~\new_[5414]_  | ~\new_[7605]_ ;
  assign \new_[7214]_  = ~\new_[5415]_  | ~\new_[7605]_ ;
  assign \new_[7215]_  = ~\new_[5416]_  | ~\new_[7605]_ ;
  assign \new_[7216]_  = ~\new_[5689]_  | ~\new_[7605]_ ;
  assign \new_[7217]_  = ~\new_[5417]_  | ~\new_[7605]_ ;
  assign \new_[7218]_  = ~\new_[5418]_  | ~\new_[7605]_ ;
  assign \new_[7219]_  = ~\new_[5419]_  | ~\new_[7605]_ ;
  assign \new_[7220]_  = ~\new_[5691]_  | ~\new_[7605]_ ;
  assign \new_[7221]_  = ~\new_[5420]_  | ~\new_[7605]_ ;
  assign \new_[7222]_  = ~\new_[5421]_  | ~\new_[7605]_ ;
  assign \new_[7223]_  = ~\new_[5422]_  | ~\new_[7605]_ ;
  assign \new_[7224]_  = ~\new_[5690]_  | ~\new_[7605]_ ;
  assign \new_[7225]_  = ~\new_[5423]_  | ~\new_[7605]_ ;
  assign \new_[7226]_  = ~\new_[5424]_  | ~\new_[7605]_ ;
  assign \new_[7227]_  = ~\new_[5425]_  | ~\new_[7605]_ ;
  assign \new_[7228]_  = ~\new_[5676]_  | ~\new_[7605]_ ;
  assign \new_[7229]_  = ~\new_[5426]_  | ~\new_[7605]_ ;
  assign \new_[7230]_  = ~\new_[5427]_  | ~\new_[7605]_ ;
  assign \new_[7231]_  = ~\new_[5428]_  | ~\new_[7605]_ ;
  assign \new_[7232]_  = ~\new_[5678]_  | ~\new_[7605]_ ;
  assign \new_[7233]_  = ~\new_[5429]_  | ~\new_[7605]_ ;
  assign \new_[7234]_  = ~\new_[5430]_  | ~\new_[7605]_ ;
  assign \new_[7235]_  = ~\new_[5431]_  | ~\new_[7605]_ ;
  assign \new_[7236]_  = ~\new_[5675]_  | ~\new_[7605]_ ;
  assign \new_[7237]_  = ~\new_[5432]_  | ~\new_[7605]_ ;
  assign \new_[7238]_  = ~\new_[5433]_  | ~\new_[7605]_ ;
  assign \new_[7239]_  = ~\new_[5434]_  | ~\new_[7605]_ ;
  assign \new_[7240]_  = ~\new_[5674]_  | ~\new_[7605]_ ;
  assign \new_[7241]_  = ~\new_[5435]_  | ~\new_[7605]_ ;
  assign \new_[7242]_  = ~\new_[5436]_  | ~\new_[7605]_ ;
  assign \new_[7243]_  = ~\new_[5437]_  | ~\new_[7605]_ ;
  assign \new_[7244]_  = ~\new_[5672]_  | ~\new_[7605]_ ;
  assign \new_[7245]_  = ~\new_[5438]_  | ~\new_[7605]_ ;
  assign \new_[7246]_  = ~\new_[5439]_  | ~\new_[7605]_ ;
  assign \new_[7247]_  = ~\new_[5440]_  | ~\new_[7605]_ ;
  assign \new_[7248]_  = ~\new_[5670]_  | ~\new_[7605]_ ;
  assign \new_[7249]_  = ~\new_[5441]_  | ~\new_[7605]_ ;
  assign \new_[7250]_  = ~\new_[5442]_  | ~\new_[7605]_ ;
  assign \new_[7251]_  = ~\new_[5443]_  | ~\new_[7605]_ ;
  assign \new_[7252]_  = ~\new_[5035]_  | ~\new_[7605]_ ;
  assign \new_[7253]_  = ~\new_[5444]_  | ~\new_[7605]_ ;
  assign \new_[7254]_  = ~\new_[5170]_  | ~\new_[7616]_ ;
  assign \new_[7255]_  = ~\new_[5546]_  | ~\new_[7616]_ ;
  assign \new_[7256]_  = ~\new_[4935]_  | ~\new_[7533]_ ;
  assign \new_[7257]_  = ~\new_[5182]_  | ~\new_[7533]_ ;
  assign \new_[7258]_  = ~\new_[5179]_  | ~\new_[7609]_ ;
  assign \new_[7259]_  = ~\new_[5446]_  | ~\new_[7614]_ ;
  assign \new_[7260]_  = ~\new_[5666]_  | ~\new_[7614]_ ;
  assign \new_[7261]_  = ~\new_[5447]_  | ~\new_[7614]_ ;
  assign \new_[7262]_  = ~\new_[5448]_  | ~\new_[7614]_ ;
  assign \new_[7263]_  = ~\new_[5449]_  | ~\new_[7614]_ ;
  assign \new_[7264]_  = ~\new_[5302]_  | ~\new_[7614]_ ;
  assign \new_[7265]_  = ~\new_[5450]_  | ~\new_[7614]_ ;
  assign \new_[7266]_  = ~\new_[5451]_  | ~\new_[7614]_ ;
  assign \new_[7267]_  = ~\new_[5452]_  | ~\new_[7614]_ ;
  assign \new_[7268]_  = ~\new_[5453]_  | ~\new_[7614]_ ;
  assign \new_[7269]_  = ~\new_[5454]_  | ~\new_[7614]_ ;
  assign \new_[7270]_  = ~\new_[5455]_  | ~\new_[7614]_ ;
  assign \new_[7271]_  = ~\new_[5456]_  | ~\new_[7614]_ ;
  assign \new_[7272]_  = ~\new_[5613]_  | ~\new_[7614]_ ;
  assign \new_[7273]_  = ~\new_[5457]_  | ~\new_[7614]_ ;
  assign \new_[7274]_  = ~\new_[5458]_  | ~\new_[7614]_ ;
  assign \new_[7275]_  = ~\new_[5459]_  | ~\new_[7614]_ ;
  assign \new_[7276]_  = ~\new_[4968]_  | ~\new_[7614]_ ;
  assign \new_[7277]_  = ~\new_[5566]_  | ~\new_[7616]_ ;
  assign \new_[7278]_  = ~\new_[5460]_  | ~\new_[7614]_ ;
  assign \new_[7279]_  = ~\new_[5461]_  | ~\new_[7614]_ ;
  assign \new_[7280]_  = ~\new_[5570]_  | ~\new_[7616]_ ;
  assign \new_[7281]_  = ~\new_[5462]_  | ~\new_[7614]_ ;
  assign \new_[7282]_  = ~\new_[5046]_  | ~\new_[7614]_ ;
  assign \new_[7283]_  = ~\new_[5571]_  | ~\new_[7533]_ ;
  assign \new_[7284]_  = ~\new_[5463]_  | ~\new_[7614]_ ;
  assign \new_[7285]_  = ~\new_[5464]_  | ~\new_[7614]_ ;
  assign \new_[7286]_  = ~\new_[5038]_  | ~\new_[7614]_ ;
  assign \new_[7287]_  = ~\new_[5466]_  | ~\new_[7614]_ ;
  assign \new_[7288]_  = ~\new_[5467]_  | ~\new_[7614]_ ;
  assign \new_[7289]_  = ~\new_[5468]_  | ~\new_[7614]_ ;
  assign \new_[7290]_  = ~\new_[5034]_  | ~\new_[7614]_ ;
  assign \new_[7291]_  = ~\new_[5469]_  | ~\new_[7614]_ ;
  assign \new_[7292]_  = ~\new_[5470]_  | ~\new_[7614]_ ;
  assign \new_[7293]_  = ~\new_[5471]_  | ~\new_[7614]_ ;
  assign \new_[7294]_  = ~\new_[5031]_  | ~\new_[7614]_ ;
  assign \new_[7295]_  = ~\new_[5472]_  | ~\new_[7614]_ ;
  assign \new_[7296]_  = ~\new_[5473]_  | ~\new_[7614]_ ;
  assign \new_[7297]_  = ~\new_[5474]_  | ~\new_[7614]_ ;
  assign \new_[7298]_  = ~\new_[5030]_  | ~\new_[7614]_ ;
  assign \new_[7299]_  = ~\new_[5475]_  | ~\new_[7614]_ ;
  assign \new_[7300]_  = ~\new_[5476]_  | ~\new_[7614]_ ;
  assign \new_[7301]_  = ~\new_[5477]_  | ~\new_[7614]_ ;
  assign \new_[7302]_  = ~\new_[5027]_  | ~\new_[7614]_ ;
  assign \new_[7303]_  = ~\new_[5478]_  | ~\new_[7614]_ ;
  assign \new_[7304]_  = ~\new_[5480]_  | ~\new_[7614]_ ;
  assign \new_[7305]_  = ~\new_[5026]_  | ~\new_[7614]_ ;
  assign \new_[7306]_  = ~\new_[5481]_  | ~\new_[7614]_ ;
  assign \new_[7307]_  = ~\new_[5482]_  | ~\new_[7614]_ ;
  assign \new_[7308]_  = ~\new_[5483]_  | ~\new_[7614]_ ;
  assign \new_[7309]_  = ~\new_[5012]_  | ~\new_[7614]_ ;
  assign \new_[7310]_  = ~\new_[5484]_  | ~\new_[7614]_ ;
  assign \new_[7311]_  = ~\new_[5485]_  | ~\new_[7614]_ ;
  assign \new_[7312]_  = ~\new_[5486]_  | ~\new_[7614]_ ;
  assign \new_[7313]_  = ~\new_[5487]_  | ~\new_[7614]_ ;
  assign \new_[7314]_  = ~\new_[5488]_  | ~\new_[7614]_ ;
  assign \new_[7315]_  = ~\new_[5568]_  | ~\new_[7616]_ ;
  assign \new_[7316]_  = ~\new_[5489]_  | ~\new_[7614]_ ;
  assign \new_[7317]_  = ~\new_[5023]_  | ~\new_[7614]_ ;
  assign \new_[7318]_  = ~\new_[5490]_  | ~\new_[7614]_ ;
  assign \new_[7319]_  = ~\new_[5491]_  | ~\new_[7614]_ ;
  assign \new_[7320]_  = ~\new_[5492]_  | ~\new_[7614]_ ;
  assign \new_[7321]_  = ~\new_[5013]_  | ~\new_[7614]_ ;
  assign \new_[7322]_  = ~\new_[5493]_  | ~\new_[7614]_ ;
  assign \new_[7323]_  = ~\new_[5494]_  | ~\new_[7614]_ ;
  assign \new_[7324]_  = ~\new_[5495]_  | ~\new_[7614]_ ;
  assign \new_[7325]_  = ~\new_[5014]_  | ~\new_[7614]_ ;
  assign \new_[7326]_  = ~\new_[5496]_  | ~\new_[7614]_ ;
  assign \new_[7327]_  = ~\new_[5497]_  | ~\new_[7614]_ ;
  assign \new_[7328]_  = ~\new_[5498]_  | ~\new_[7614]_ ;
  assign \new_[7329]_  = ~\new_[4995]_  | ~\new_[7614]_ ;
  assign \new_[7330]_  = ~\new_[5499]_  | ~\new_[7614]_ ;
  assign \new_[7331]_  = ~\new_[5500]_  | ~\new_[7614]_ ;
  assign \new_[7332]_  = ~\new_[5501]_  | ~\new_[7614]_ ;
  assign \new_[7333]_  = ~\new_[5004]_  | ~\new_[7614]_ ;
  assign \new_[7334]_  = ~\new_[5502]_  | ~\new_[7614]_ ;
  assign \new_[7335]_  = ~\new_[5503]_  | ~\new_[7614]_ ;
  assign \new_[7336]_  = ~\new_[5504]_  | ~\new_[7614]_ ;
  assign \new_[7337]_  = ~\new_[5003]_  | ~\new_[7614]_ ;
  assign \new_[7338]_  = ~\new_[5506]_  | ~\new_[7614]_ ;
  assign \new_[7339]_  = ~\new_[5507]_  | ~\new_[7614]_ ;
  assign \new_[7340]_  = ~\new_[5508]_  | ~\new_[7614]_ ;
  assign \new_[7341]_  = ~\new_[4996]_  | ~\new_[7614]_ ;
  assign \new_[7342]_  = ~\new_[5509]_  | ~\new_[7614]_ ;
  assign \new_[7343]_  = ~\new_[5510]_  | ~\new_[7614]_ ;
  assign \new_[7344]_  = ~\new_[5511]_  | ~\new_[7614]_ ;
  assign \new_[7345]_  = ~\new_[4997]_  | ~\new_[7614]_ ;
  assign \new_[7346]_  = ~\new_[5512]_  | ~\new_[7614]_ ;
  assign \new_[7347]_  = ~\new_[5150]_  | ~\new_[7616]_ ;
  assign \new_[7348]_  = ~\new_[5513]_  | ~\new_[7614]_ ;
  assign \new_[7349]_  = ~\new_[5514]_  | ~\new_[7614]_ ;
  assign \new_[7350]_  = ~\new_[4971]_  | ~\new_[7614]_ ;
  assign \new_[7351]_  = ~\new_[5515]_  | ~\new_[7614]_ ;
  assign \new_[7352]_  = ~\new_[5516]_  | ~\new_[7614]_ ;
  assign \new_[7353]_  = ~\new_[5517]_  | ~\new_[7614]_ ;
  assign \new_[7354]_  = ~\new_[4990]_  | ~\new_[7614]_ ;
  assign \new_[7355]_  = ~\new_[5518]_  | ~\new_[7614]_ ;
  assign \new_[7356]_  = ~\new_[5519]_  | ~\new_[7614]_ ;
  assign \new_[7357]_  = ~\new_[4976]_  | ~\new_[7532]_ ;
  assign \new_[7358]_  = ~\new_[5148]_  | ~\new_[7609]_ ;
  assign \new_[7359]_  = ~\new_[5180]_  | ~\new_[7533]_ ;
  assign \new_[7360]_  = ~\new_[4908]_  | ~\new_[7616]_ ;
  assign \new_[7361]_  = ~\new_[4987]_  | ~\new_[7616]_ ;
  assign \new_[7362]_  = ~\new_[5521]_  | ~\new_[7616]_ ;
  assign \new_[7363]_  = ~\new_[5523]_  | ~\new_[7616]_ ;
  assign \new_[7364]_  = ~\new_[4972]_  | ~\new_[7616]_ ;
  assign \new_[7365]_  = ~\new_[5524]_  | ~\new_[7616]_ ;
  assign \new_[7366]_  = ~\new_[5526]_  | ~\new_[7616]_ ;
  assign \new_[7367]_  = ~\new_[5146]_  | ~\new_[7616]_ ;
  assign \new_[7368]_  = ~\new_[4973]_  | ~\new_[7616]_ ;
  assign \new_[7369]_  = ~\new_[5145]_  | ~\new_[7533]_ ;
  assign \new_[7370]_  = ~\new_[5527]_  | ~\new_[7616]_ ;
  assign \new_[7371]_  = ~\new_[5529]_  | ~\new_[7616]_ ;
  assign \new_[7372]_  = ~\new_[4943]_  | ~\new_[7616]_ ;
  assign \new_[7373]_  = ~\new_[5530]_  | ~\new_[7616]_ ;
  assign \new_[7374]_  = ~\new_[5532]_  | ~\new_[7616]_ ;
  assign \new_[7375]_  = ~\new_[4964]_  | ~\new_[7616]_ ;
  assign \new_[7376]_  = ~\new_[5534]_  | ~\new_[7609]_ ;
  assign \new_[7377]_  = ~\new_[5533]_  | ~\new_[7616]_ ;
  assign \new_[7378]_  = ~\new_[5535]_  | ~\new_[7616]_ ;
  assign \new_[7379]_  = ~\new_[5536]_  | ~\new_[7533]_ ;
  assign \new_[7380]_  = ~\new_[4962]_  | ~\new_[7616]_ ;
  assign \new_[7381]_  = ~\new_[5538]_  | ~\new_[7616]_ ;
  assign \new_[7382]_  = ~\new_[5539]_  | ~\new_[7616]_ ;
  assign \new_[7383]_  = ~\new_[5541]_  | ~\new_[7533]_ ;
  assign \new_[7384]_  = ~\new_[5540]_  | ~\new_[7616]_ ;
  assign \new_[7385]_  = ~\new_[5543]_  | ~\new_[7533]_ ;
  assign \new_[7386]_  = ~\new_[5544]_  | ~\new_[7616]_ ;
  assign \new_[7387]_  = ~\new_[5545]_  | ~\new_[7609]_ ;
  assign \new_[7388]_  = ~\new_[4916]_  | ~\new_[7616]_ ;
  assign \new_[7389]_  = ~\new_[5547]_  | ~\new_[7616]_ ;
  assign \new_[7390]_  = ~\new_[5548]_  | ~\new_[7616]_ ;
  assign \new_[7391]_  = ~\new_[5550]_  | ~\new_[7609]_ ;
  assign \new_[7392]_  = ~\new_[5549]_  | ~\new_[7616]_ ;
  assign \new_[7393]_  = ~\new_[5551]_  | ~\new_[7616]_ ;
  assign \new_[7394]_  = ~\new_[5554]_  | ~\new_[7616]_ ;
  assign \new_[7395]_  = ~\new_[5555]_  | ~\new_[7609]_ ;
  assign \new_[7396]_  = ~\new_[5561]_  | ~\new_[7616]_ ;
  assign \new_[7397]_  = ~\new_[5556]_  | ~\new_[7616]_ ;
  assign \new_[7398]_  = ~\new_[4920]_  | ~\new_[7609]_ ;
  assign \new_[7399]_  = ~\new_[5557]_  | ~\new_[7616]_ ;
  assign \new_[7400]_  = ~\new_[5558]_  | ~\new_[7616]_ ;
  assign \new_[7401]_  = ~\new_[5560]_  | ~\new_[7533]_ ;
  assign \new_[7402]_  = ~\new_[4896]_  | ~\new_[7616]_ ;
  assign \new_[7403]_  = ~\new_[5563]_  | ~\new_[7616]_ ;
  assign \new_[7404]_  = ~\new_[5564]_  | ~\new_[7533]_ ;
  assign \new_[7405]_  = ~\new_[5565]_  | ~\new_[7616]_ ;
  assign \new_[7406]_  = ~\new_[4907]_  | ~\new_[7609]_ ;
  assign \new_[7407]_  = ~\new_[5567]_  | ~\new_[7616]_ ;
  assign \new_[7408]_  = ~\new_[5569]_  | ~\new_[7533]_ ;
  assign \new_[7409]_  = ~\new_[4898]_  | ~\new_[7616]_ ;
  assign \new_[7410]_  = ~\new_[5572]_  | ~\new_[7616]_ ;
  assign \new_[7411]_  = ~\new_[5573]_  | ~\new_[7533]_ ;
  assign \new_[7412]_  = ~\new_[5537]_  | ~\new_[7616]_ ;
  assign \new_[7413]_  = ~\new_[5574]_  | ~\new_[7616]_ ;
  assign \new_[7414]_  = ~\new_[5759]_  | ~\new_[7533]_ ;
  assign \new_[7415]_  = ~\new_[5575]_  | ~\new_[7616]_ ;
  assign \new_[7416]_  = ~\new_[5576]_  | ~\new_[7616]_ ;
  assign \new_[7417]_  = ~\new_[5578]_  | ~\new_[7609]_ ;
  assign \new_[7418]_  = ~\new_[5763]_  | ~\new_[7616]_ ;
  assign n9651 = \new_[8995]_  ? \new_[7638]_  : \new_[6440]_ ;
  assign \new_[7420]_  = ~\new_[7459]_ ;
  assign \new_[7421]_  = ~\new_[13320]_  & ~\new_[14004]_ ;
  assign \new_[7422]_  = ~\new_[13769]_  & ~\new_[14004]_ ;
  assign \new_[7423]_  = ~\new_[13824]_  & ~\new_[14004]_ ;
  assign \new_[7424]_  = ~\new_[13575]_  & ~\new_[14004]_ ;
  assign \new_[7425]_  = ~\new_[13574]_  & ~\new_[14004]_ ;
  assign n9646 = ~\new_[7465]_ ;
  assign \new_[7427]_  = ~\new_[12914]_  | (~\new_[8832]_  & ~\new_[7599]_ );
  assign \new_[7428]_  = ~\new_[12985]_  | (~\new_[8833]_  & ~\new_[7601]_ );
  assign \new_[7429]_  = ~\new_[12801]_  & (~\new_[7600]_  | ~\new_[13005]_ );
  assign \new_[7430]_  = ~\new_[12755]_  & (~\new_[7602]_  | ~\new_[13006]_ );
  assign \new_[7431]_  = ~u3_empty_reg;
  assign \new_[7432]_  = ~u5_empty_reg;
  assign \new_[7433]_  = ~u7_empty_reg;
  assign \new_[7434]_  = ~u8_empty_reg;
  assign n9656 = \new_[7507]_  & \new_[13166]_ ;
  assign n9661 = \new_[7507]_  & \new_[13189]_ ;
  assign \new_[7437]_  = \new_[9079]_  | \new_[7519]_ ;
  assign \new_[7438]_  = \\u10_rp_reg[2] ;
  assign \new_[7439]_  = \\u11_rp_reg[2] ;
  assign n9791 = ~\new_[7508]_ ;
  assign \new_[7441]_  = ~\new_[7509]_ ;
  assign \new_[7442]_  = ~\new_[7510]_ ;
  assign \new_[7443]_  = ~\new_[7511]_ ;
  assign n9781 = ~\new_[7626]_  & ~\new_[9710]_ ;
  assign n9786 = ~\new_[7628]_  & ~\new_[9711]_ ;
  assign n9696 = n9906 ? \new_[9000]_  : \new_[6794]_ ;
  assign n9691 = n9906 ? \new_[8996]_  : \new_[6793]_ ;
  assign n9681 = n9906 ? \new_[9002]_  : \new_[6791]_ ;
  assign n9771 = n9906 ? \new_[9001]_  : \new_[6809]_ ;
  assign n9686 = n9906 ? \new_[8805]_  : \new_[6792]_ ;
  assign \new_[7451]_  = ~\new_[7609]_ ;
  assign n9716 = ~\new_[8173]_  | ~\new_[7662]_ ;
  assign n9731 = ~\new_[8169]_  | ~\new_[7663]_ ;
  assign n9726 = ~\new_[8154]_  | ~\new_[7658]_ ;
  assign n9721 = ~\new_[7856]_  | ~\new_[7659]_ ;
  assign n9711 = ~\new_[8164]_  | ~\new_[7660]_ ;
  assign n9706 = ~\new_[8161]_  | ~\new_[7661]_ ;
  assign n9701 = ~\new_[7664]_  | ~\new_[8155]_ ;
  assign \new_[7459]_  = ~\new_[7639]_  & ~\new_[13810]_ ;
  assign n9671 = ~\new_[7637]_  & ~\new_[13316]_ ;
  assign \new_[7461]_  = \new_[13867]_  | \new_[7637]_ ;
  assign \new_[7462]_  = ~\new_[13873]_  | ~\new_[7816]_ ;
  assign \new_[7463]_  = \new_[13877]_  | \new_[7639]_ ;
  assign n9776 = ~\new_[8104]_  | ~\new_[7657]_ ;
  assign \new_[7465]_  = ~\new_[7593]_ ;
  assign \new_[7466]_  = ~\new_[7641]_  & (~\new_[8811]_  | ~\new_[9782]_ );
  assign \new_[7467]_  = ~\new_[7642]_  & (~\new_[8810]_  | ~\new_[9782]_ );
  assign \new_[7468]_  = ~\new_[7643]_  & (~\new_[8813]_  | ~\new_[9782]_ );
  assign \new_[7469]_  = ~\new_[7640]_  & (~\new_[8545]_  | ~\new_[9782]_ );
  assign \new_[7470]_  = ~\new_[7646]_  & (~\new_[8819]_  | ~\new_[9782]_ );
  assign \new_[7471]_  = ~\new_[7647]_  & (~\new_[8821]_  | ~\new_[9782]_ );
  assign \new_[7472]_  = ~\new_[7648]_  & (~\new_[8822]_  | ~\new_[9782]_ );
  assign \new_[7473]_  = ~\new_[7649]_  & (~\new_[9049]_  | ~\new_[9782]_ );
  assign \new_[7474]_  = ~\new_[7650]_  & (~\new_[8823]_  | ~\new_[9782]_ );
  assign \new_[7475]_  = ~\new_[7651]_  & (~\new_[8824]_  | ~\new_[9782]_ );
  assign \new_[7476]_  = ~\new_[7652]_  & (~\new_[8825]_  | ~\new_[9782]_ );
  assign \new_[7477]_  = ~\new_[7653]_  & (~\new_[9782]_  | ~\new_[8826]_ );
  assign \new_[7478]_  = ~\new_[7644]_  & (~\new_[8814]_  | ~\new_[9782]_ );
  assign \new_[7479]_  = ~\new_[7645]_  & (~\new_[8544]_  | ~\new_[10402]_ );
  assign \new_[7480]_  = ~\new_[7654]_  & (~\new_[8812]_  | ~\new_[9782]_ );
  assign \new_[7481]_  = ~\new_[7655]_  & (~\new_[10819]_  | ~\new_[5083]_ );
  assign n9736 = ~\new_[7679]_  | ~\new_[8174]_ ;
  assign n9766 = ~\new_[7598]_  | ~\new_[7964]_ ;
  assign n9756 = ~\new_[7681]_  | ~\new_[8156]_ ;
  assign n9751 = ~\new_[7682]_  | ~\new_[8157]_ ;
  assign n9746 = ~\new_[7683]_  | ~\new_[8158]_ ;
  assign n9761 = ~\new_[7685]_  | ~\new_[8113]_ ;
  assign n9741 = ~\new_[7684]_  | ~\new_[8106]_ ;
  assign n9676 = ~\new_[8159]_  | ~\new_[7680]_ ;
  assign \new_[7490]_  = \\u23_int_set_reg[1] ;
  assign \new_[7491]_  = \\u24_int_set_reg[1] ;
  assign \new_[7492]_  = \\u11_rp_reg[1] ;
  assign \new_[7493]_  = \\u9_rp_reg[1] ;
  assign \new_[7494]_  = \\u10_rp_reg[1] ;
  assign \new_[7495]_  = \\u11_rp_reg[0] ;
  assign \new_[7496]_  = \\u9_rp_reg[0] ;
  assign \new_[7497]_  = \\u9_rp_reg[2] ;
  assign \new_[7498]_  = \\u10_rp_reg[0] ;
  assign \new_[7499]_  = \\u1_slt1_reg[5] ;
  assign \new_[7500]_  = \\u1_slt2_reg[5] ;
  assign \new_[7501]_  = \\u1_slt4_reg[5] ;
  assign \new_[7502]_  = \\u1_slt3_reg[5] ;
  assign \new_[7503]_  = \\u1_slt6_reg[5] ;
  assign \new_[7504]_  = \new_[8830]_  | \new_[7603]_ ;
  assign \new_[7505]_  = \new_[8831]_  | \new_[7604]_ ;
  assign \new_[7506]_  = \\u25_int_set_reg[1] ;
  assign \new_[7507]_  = \new_[7702]_  & \new_[13125]_ ;
  assign \new_[7508]_  = ~\new_[7703]_  | ~\new_[13103]_ ;
  assign \new_[7509]_  = ~\new_[12831]_  | ~\new_[7704]_ ;
  assign \new_[7510]_  = ~\new_[7703]_  | ~\new_[12926]_ ;
  assign \new_[7511]_  = \new_[7705]_  & \new_[13125]_ ;
  assign \new_[7512]_  = ~\new_[13015]_  | ~\new_[7704]_ ;
  assign \new_[7513]_  = ~\new_[13007]_  | ~\new_[7708]_ ;
  assign \new_[7514]_  = \new_[10317]_  | \new_[7708]_ ;
  assign n9806 = ~\new_[7706]_  & ~\new_[11453]_ ;
  assign n9811 = ~\new_[9712]_  & ~\new_[7709]_ ;
  assign n9801 = ~\new_[7710]_  & ~\new_[9713]_ ;
  assign n9816 = ~\new_[7711]_  & ~\new_[10396]_ ;
  assign \new_[7519]_  = \new_[12638]_  | \new_[7707]_ ;
  assign \new_[7520]_  = ~\new_[7606]_ ;
  assign \new_[7521]_  = ~\new_[7606]_ ;
  assign \new_[7522]_  = ~\new_[7606]_ ;
  assign \new_[7523]_  = ~\new_[7606]_ ;
  assign \new_[7524]_  = ~\new_[7606]_ ;
  assign \new_[7525]_  = ~\new_[7606]_ ;
  assign \new_[7526]_  = ~\new_[7606]_ ;
  assign \new_[7527]_  = ~\new_[7606]_ ;
  assign \new_[7528]_  = ~\new_[7605]_ ;
  assign \new_[7529]_  = ~\new_[7606]_ ;
  assign \new_[7530]_  = ~\new_[7606]_ ;
  assign \new_[7531]_  = ~\new_[7606]_ ;
  assign \new_[7532]_  = ~\new_[7608]_ ;
  assign \new_[7533]_  = ~\new_[7608]_ ;
  assign \new_[7534]_  = ~\new_[7607]_ ;
  assign \new_[7535]_  = ~\new_[7607]_ ;
  assign \new_[7536]_  = ~\new_[7607]_ ;
  assign \new_[7537]_  = ~\new_[7607]_ ;
  assign \new_[7538]_  = ~\new_[7607]_ ;
  assign \new_[7539]_  = ~\new_[7607]_ ;
  assign \new_[7540]_  = ~\new_[7607]_ ;
  assign \new_[7541]_  = ~\new_[7607]_ ;
  assign \new_[7542]_  = ~\new_[7608]_ ;
  assign \new_[7543]_  = ~\new_[7607]_ ;
  assign \new_[7544]_  = ~\new_[7607]_ ;
  assign \new_[7545]_  = ~\new_[7607]_ ;
  assign \new_[7546]_  = ~\new_[7611]_ ;
  assign \new_[7547]_  = ~\new_[7611]_ ;
  assign \new_[7548]_  = ~\new_[7611]_ ;
  assign \new_[7549]_  = ~\new_[7611]_ ;
  assign \new_[7550]_  = ~\new_[7611]_ ;
  assign \new_[7551]_  = ~\new_[7611]_ ;
  assign \new_[7552]_  = ~\new_[7610]_ ;
  assign \new_[7553]_  = ~\new_[7611]_ ;
  assign \new_[7554]_  = ~\new_[7613]_ ;
  assign \new_[7555]_  = ~\new_[7613]_ ;
  assign \new_[7556]_  = ~\new_[7613]_ ;
  assign \new_[7557]_  = ~\new_[7613]_ ;
  assign \new_[7558]_  = ~\new_[7613]_ ;
  assign \new_[7559]_  = ~\new_[7613]_ ;
  assign \new_[7560]_  = ~\new_[7613]_ ;
  assign \new_[7561]_  = ~\new_[7612]_ ;
  assign \new_[7562]_  = ~\new_[7613]_ ;
  assign \new_[7563]_  = ~\new_[7613]_ ;
  assign \new_[7564]_  = ~\new_[7613]_ ;
  assign \new_[7565]_  = ~\new_[7615]_ ;
  assign \new_[7566]_  = ~\new_[7615]_ ;
  assign \new_[7567]_  = ~\new_[7615]_ ;
  assign \new_[7568]_  = ~\new_[7615]_ ;
  assign \new_[7569]_  = ~\new_[7615]_ ;
  assign \new_[7570]_  = ~\new_[7615]_ ;
  assign \new_[7571]_  = ~\new_[7615]_ ;
  assign \new_[7572]_  = ~\new_[7615]_ ;
  assign \new_[7573]_  = ~\new_[7615]_ ;
  assign \new_[7574]_  = ~\new_[7615]_ ;
  assign \new_[7575]_  = ~\new_[7614]_ ;
  assign \new_[7576]_  = ~\new_[7615]_ ;
  assign \new_[7577]_  = ~\new_[7615]_ ;
  assign \new_[7578]_  = ~\new_[7615]_ ;
  assign \new_[7579]_  = ~\new_[7617]_ ;
  assign \new_[7580]_  = ~\new_[7617]_ ;
  assign \new_[7581]_  = ~\new_[7617]_ ;
  assign \new_[7582]_  = ~\new_[7617]_ ;
  assign \new_[7583]_  = ~\new_[7617]_ ;
  assign \new_[7584]_  = ~\new_[7617]_ ;
  assign \new_[7585]_  = ~\new_[7617]_ ;
  assign \new_[7586]_  = ~\new_[7617]_ ;
  assign \new_[7587]_  = ~\new_[7617]_ ;
  assign \new_[7588]_  = ~\new_[7616]_ ;
  assign \new_[7589]_  = ~\new_[7617]_ ;
  assign \new_[7590]_  = ~\new_[7617]_ ;
  assign \new_[7591]_  = ~\new_[7617]_ ;
  assign n9796 = \\u1_sr_reg[7] ;
  assign \new_[7593]_  = ~\new_[7714]_  & ~\new_[13314]_ ;
  assign \new_[7594]_  = \\u0_slt9_r_reg[0] ;
  assign \new_[7595]_  = ~\new_[7637]_ ;
  assign \new_[7596]_  = ~\new_[7639]_ ;
  assign \new_[7597]_  = ~\new_[12638]_  & (~\new_[7812]_  | ~\new_[12862]_ );
  assign \new_[7598]_  = ~\new_[7863]_  & (~\new_[9016]_  | ~\new_[9784]_ );
  assign \new_[7599]_  = ~\new_[13005]_  | ~\new_[7810]_ ;
  assign \new_[7600]_  = \new_[9677]_  | \new_[7810]_ ;
  assign \new_[7601]_  = ~\new_[13006]_  | ~\new_[7811]_ ;
  assign \new_[7602]_  = \new_[9673]_  | \new_[7811]_ ;
  assign \new_[7603]_  = \new_[12636]_  | \new_[7808]_ ;
  assign \new_[7604]_  = \new_[12637]_  | \new_[7809]_ ;
  assign \new_[7605]_  = ~\new_[7696]_ ;
  assign \new_[7606]_  = \new_[7696]_ ;
  assign \new_[7607]_  = \new_[7697]_ ;
  assign \new_[7608]_  = \new_[7697]_ ;
  assign \new_[7609]_  = ~\new_[7697]_ ;
  assign \new_[7610]_  = ~\new_[7698]_ ;
  assign \new_[7611]_  = \new_[7698]_ ;
  assign \new_[7612]_  = ~\new_[7699]_ ;
  assign \new_[7613]_  = \new_[7699]_ ;
  assign \new_[7614]_  = ~\new_[7700]_ ;
  assign \new_[7615]_  = \new_[7700]_ ;
  assign \new_[7616]_  = ~\new_[7701]_ ;
  assign \new_[7617]_  = \new_[7701]_ ;
  assign n9846 = ~\new_[7818]_  & ~\new_[13867]_ ;
  assign n9851 = ~\new_[7820]_  & ~\new_[13874]_ ;
  assign n9841 = ~\new_[7817]_  & ~\new_[13877]_ ;
  assign n9866 = ~\new_[7823]_  & ~\new_[13867]_ ;
  assign n9826 = ~\new_[7824]_  & ~\new_[13877]_ ;
  assign n9821 = ~\new_[7825]_  & ~\new_[13874]_ ;
  assign n9856 = ~\new_[7829]_  & ~\new_[13877]_ ;
  assign n9861 = ~\new_[7827]_  & ~\new_[13867]_ ;
  assign \new_[7626]_  = ~\new_[12337]_  | ~\new_[8314]_  | ~\new_[7965]_ ;
  assign n9871 = ~\new_[7828]_  & ~\new_[13874]_ ;
  assign \new_[7628]_  = ~\new_[11713]_  | ~\new_[7922]_  | ~\new_[8533]_ ;
  assign n9831 = \new_[7821]_  | \new_[7490]_ ;
  assign n9836 = \new_[7822]_  | \new_[7491]_ ;
  assign n9886 = n9976 ? \new_[9000]_  : \new_[7501]_ ;
  assign n9896 = n9976 ? \new_[9001]_  : \new_[7503]_ ;
  assign n9881 = n9976 ? \new_[8996]_  : \new_[7500]_ ;
  assign n9876 = n9976 ? \new_[8805]_  : \new_[7499]_ ;
  assign n9891 = n9976 ? \new_[9002]_  : \new_[7502]_ ;
  assign \new_[7636]_  = valid_s_reg;
  assign \new_[7637]_  = ~\\in_valid_s_reg[0] ;
  assign \new_[7638]_  = ~\new_[7714]_ ;
  assign \new_[7639]_  = ~\new_[7715]_ ;
  assign \new_[7640]_  = ~\new_[8413]_  & (~\new_[7996]_  | ~\new_[9774]_ );
  assign \new_[7641]_  = ~\new_[8413]_  & (~\new_[7993]_  | ~\new_[9746]_ );
  assign \new_[7642]_  = ~\new_[8413]_  & (~\new_[7994]_  | ~\new_[9775]_ );
  assign \new_[7643]_  = ~\new_[8413]_  & (~\new_[8005]_  | ~\new_[9748]_ );
  assign \new_[7644]_  = ~\new_[8413]_  & (~\new_[7995]_  | ~\new_[9749]_ );
  assign \new_[7645]_  = ~\new_[8413]_  & (~\new_[8007]_  | ~\new_[9776]_ );
  assign \new_[7646]_  = ~\new_[8413]_  & (~\new_[7997]_  | ~\new_[9764]_ );
  assign \new_[7647]_  = ~\new_[8413]_  & (~\new_[7998]_  | ~\new_[9765]_ );
  assign \new_[7648]_  = ~\new_[8413]_  & (~\new_[7999]_  | ~\new_[9766]_ );
  assign \new_[7649]_  = ~\new_[8413]_  & (~\new_[8000]_  | ~\new_[9768]_ );
  assign \new_[7650]_  = ~\new_[8413]_  & (~\new_[8001]_  | ~\new_[9769]_ );
  assign \new_[7651]_  = ~\new_[8413]_  & (~\new_[8002]_  | ~\new_[9770]_ );
  assign \new_[7652]_  = ~\new_[8413]_  & (~\new_[8003]_  | ~\new_[9771]_ );
  assign \new_[7653]_  = ~\new_[8413]_  & (~\new_[8004]_  | ~\new_[9772]_ );
  assign \new_[7654]_  = ~\new_[8413]_  & (~\new_[8006]_  | ~\new_[9747]_ );
  assign \new_[7655]_  = ~\new_[9250]_  | ~\new_[7855]_ ;
  assign \new_[7656]_  = \\u1_slt2_reg[4] ;
  assign \new_[7657]_  = ~\new_[7833]_  & (~\new_[8547]_  | ~\new_[9782]_ );
  assign \new_[7658]_  = ~\new_[7834]_  & (~\new_[8548]_  | ~\new_[9782]_ );
  assign \new_[7659]_  = ~\new_[7835]_  & (~\new_[9011]_  | ~\new_[9784]_ );
  assign \new_[7660]_  = ~\new_[7836]_  & (~\new_[8551]_  | ~\new_[9782]_ );
  assign \new_[7661]_  = ~\new_[7837]_  & (~\new_[8552]_  | ~\new_[9782]_ );
  assign \new_[7662]_  = ~\new_[7838]_  & (~\new_[9017]_  | ~\new_[9784]_ );
  assign \new_[7663]_  = ~\new_[7832]_  & (~\new_[8546]_  | ~\new_[9782]_ );
  assign \new_[7664]_  = ~\new_[7839]_  & (~\new_[8553]_  | ~\new_[9782]_ );
  assign \new_[7665]_  = ~\new_[13952]_  & (~\new_[8066]_  | ~\new_[8421]_ );
  assign \new_[7666]_  = ~\new_[12792]_  & (~\new_[8061]_  | ~\new_[8430]_ );
  assign \new_[7667]_  = ~\new_[12792]_  & (~\new_[8056]_  | ~\new_[8426]_ );
  assign \new_[7668]_  = ~\new_[12792]_  & (~\new_[8057]_  | ~\new_[8427]_ );
  assign \new_[7669]_  = ~\new_[13952]_  & (~\new_[8058]_  | ~\new_[8076]_ );
  assign \new_[7670]_  = ~\new_[13952]_  & (~\new_[8059]_  | ~\new_[8077]_ );
  assign \new_[7671]_  = ~\new_[13952]_  & (~\new_[8065]_  | ~\new_[8424]_ );
  assign \new_[7672]_  = ~\new_[12629]_  & (~\new_[8062]_  | ~\new_[8438]_ );
  assign \new_[7673]_  = ~\new_[12629]_  & (~\new_[8060]_  | ~\new_[8439]_ );
  assign \new_[7674]_  = ~\new_[12629]_  & (~\new_[8063]_  | ~\new_[8440]_ );
  assign \new_[7675]_  = ~\new_[12629]_  & (~\new_[8090]_  | ~\new_[8330]_ );
  assign \new_[7676]_  = ~\new_[12629]_  & (~\new_[8627]_  | ~\new_[8064]_ );
  assign \new_[7677]_  = ~\new_[12629]_  & (~\new_[8084]_  | ~\new_[8331]_ );
  assign \new_[7678]_  = ~\new_[14133]_  & (~\new_[8576]_  | ~\new_[8091]_ );
  assign \new_[7679]_  = ~\new_[7859]_  & (~\new_[9015]_  | ~\new_[9784]_ );
  assign \new_[7680]_  = ~\new_[7858]_  & (~\new_[9042]_  | ~\new_[9782]_ );
  assign \new_[7681]_  = ~\new_[7931]_  & (~\new_[9035]_  | ~\new_[9782]_ );
  assign \new_[7682]_  = ~\new_[7860]_  & (~\new_[8816]_  | ~\new_[9782]_ );
  assign \new_[7683]_  = ~\new_[7861]_  & (~\new_[8817]_  | ~\new_[9782]_ );
  assign \new_[7684]_  = ~\new_[7819]_  & (~\new_[8820]_  | ~\new_[10402]_ );
  assign \new_[7685]_  = ~\new_[7862]_  & (~\new_[8818]_  | ~\new_[9782]_ );
  assign \new_[7686]_  = \\u1_slt3_reg[4] ;
  assign \new_[7687]_  = \\u1_slt4_reg[4] ;
  assign \new_[7688]_  = \\u1_slt6_reg[4] ;
  assign \new_[7689]_  = ~\new_[12636]_  & (~\new_[7945]_  | ~\new_[12824]_ );
  assign \new_[7690]_  = ~\new_[12637]_  & (~\new_[7946]_  | ~\new_[12844]_ );
  assign \new_[7691]_  = ~\new_[8070]_  | (~\new_[8752]_  & ~\new_[13928]_ );
  assign \new_[7692]_  = ~\new_[7939]_  & ~\new_[13518]_ ;
  assign \new_[7693]_  = ~\new_[7940]_  & ~\new_[13437]_ ;
  assign \new_[7694]_  = ~\new_[10320]_  & ~\new_[7939]_ ;
  assign \new_[7695]_  = ~\new_[12085]_  & ~\new_[7940]_ ;
  assign \new_[7696]_  = u12_o7_we_reg;
  assign \new_[7697]_  = u12_o3_we_reg;
  assign \new_[7698]_  = u12_o4_we_reg;
  assign \new_[7699]_  = u12_o6_we_reg;
  assign \new_[7700]_  = u12_o8_we_reg;
  assign \new_[7701]_  = u12_o9_we_reg;
  assign \new_[7702]_  = ~\new_[13084]_  & ~\new_[7947]_ ;
  assign \new_[7703]_  = ~\new_[7947]_  & ~\new_[13109]_ ;
  assign \new_[7704]_  = ~\new_[7947]_  & ~\wb_addr_i[4] ;
  assign \new_[7705]_  = ~\new_[13058]_  & ~\new_[7947]_ ;
  assign \new_[7706]_  = ~\new_[11683]_  | ~\new_[8543]_  | ~\new_[8094]_ ;
  assign \new_[7707]_  = \new_[12862]_  & \new_[7948]_ ;
  assign \new_[7708]_  = ~\new_[7948]_  | ~\new_[13876]_ ;
  assign \new_[7709]_  = ~\new_[12103]_  | ~\new_[8053]_  | ~\new_[8786]_ ;
  assign \new_[7710]_  = ~\new_[11753]_  | ~\new_[8054]_  | ~\new_[8479]_ ;
  assign \new_[7711]_  = ~\new_[11681]_  | ~\new_[8055]_  | ~\new_[8502]_ ;
  assign n9901 = \new_[7957]_  | \new_[7506]_ ;
  assign n9906 = \\u1_sr_reg[6] ;
  assign \new_[7714]_  = ~\new_[7816]_ ;
  assign \new_[7715]_  = \\in_valid_s_reg[2] ;
  assign \new_[7716]_  = ~\new_[12792]_  & (~\new_[8327]_  | ~\new_[8419]_ );
  assign \new_[7717]_  = ~\new_[12792]_  & (~\new_[8326]_  | ~\new_[8422]_ );
  assign \new_[7718]_  = ~\new_[13952]_  & (~\new_[8328]_  | ~\new_[8420]_ );
  assign \new_[7719]_  = ~\new_[12650]_  & (~\new_[8590]_  | ~\new_[8317]_ );
  assign \new_[7720]_  = ~\new_[12792]_  & (~\new_[8315]_  | ~\new_[8425]_ );
  assign \new_[7721]_  = ~\new_[13952]_  & (~\new_[8318]_  | ~\new_[8428]_ );
  assign \new_[7722]_  = ~\new_[12599]_  & (~\new_[8332]_  | ~\new_[8680]_ );
  assign \new_[7723]_  = ~\new_[12792]_  & (~\new_[8320]_  | ~\new_[8423]_ );
  assign \new_[7724]_  = ~\new_[12615]_  & (~\new_[8321]_  | ~\new_[8663]_ );
  assign \new_[7725]_  = ~\new_[12615]_  & (~\new_[8322]_  | ~\new_[8664]_ );
  assign \new_[7726]_  = ~\new_[12615]_  & (~\new_[8324]_  | ~\new_[8666]_ );
  assign \new_[7727]_  = ~\new_[12615]_  & (~\new_[8325]_  | ~\new_[8452]_ );
  assign \new_[7728]_  = ~\new_[14103]_  & (~\new_[8562]_  | ~\new_[8432]_ );
  assign \new_[7729]_  = ~\new_[14103]_  & (~\new_[8416]_  | ~\new_[8564]_ );
  assign \new_[7730]_  = ~\new_[14103]_  & (~\new_[8585]_  | ~\new_[8434]_ );
  assign \new_[7731]_  = ~\new_[12615]_  & (~\new_[8354]_  | ~\new_[8673]_ );
  assign \new_[7732]_  = ~\new_[12629]_  & (~\new_[8565]_  | ~\new_[8435]_ );
  assign \new_[7733]_  = ~\new_[12629]_  & (~\new_[8566]_  | ~\new_[8436]_ );
  assign \new_[7734]_  = ~\new_[12629]_  & (~\new_[8567]_  | ~\new_[8437]_ );
  assign \new_[7735]_  = ~\new_[12629]_  & (~\new_[8568]_  | ~\new_[8418]_ );
  assign \new_[7736]_  = ~\new_[12629]_  & (~\new_[8569]_  | ~\new_[8417]_ );
  assign \new_[7737]_  = ~\new_[12629]_  & (~\new_[8554]_  | ~\new_[8441]_ );
  assign \new_[7738]_  = ~\new_[12629]_  & (~\new_[8570]_  | ~\new_[8445]_ );
  assign \new_[7739]_  = ~\new_[12629]_  & (~\new_[8571]_  | ~\new_[8374]_ );
  assign \new_[7740]_  = ~\new_[14133]_  & (~\new_[8572]_  | ~\new_[8442]_ );
  assign \new_[7741]_  = ~\new_[12629]_  & (~\new_[8573]_  | ~\new_[8443]_ );
  assign \new_[7742]_  = ~\new_[12629]_  & (~\new_[8574]_  | ~\new_[8444]_ );
  assign \new_[7743]_  = ~\new_[12599]_  & (~\new_[8414]_  | ~\new_[8346]_ );
  assign \new_[7744]_  = ~\new_[14133]_  & (~\new_[8333]_  | ~\new_[8450]_ );
  assign \new_[7745]_  = ~\new_[14133]_  & (~\new_[8334]_  | ~\new_[8431]_ );
  assign \new_[7746]_  = ~\new_[14133]_  & (~\new_[8335]_  | ~\new_[8433]_ );
  assign \new_[7747]_  = ~\new_[14133]_  & (~\new_[8336]_  | ~\new_[8446]_ );
  assign \new_[7748]_  = ~\new_[14133]_  & (~\new_[8337]_  | ~\new_[8447]_ );
  assign \new_[7749]_  = ~\new_[14133]_  & (~\new_[8329]_  | ~\new_[8448]_ );
  assign n9911 = ~\new_[7962]_  & ~\new_[2825]_ ;
  assign \new_[7751]_  = ~\new_[14133]_  & (~\new_[8338]_  | ~\new_[8449]_ );
  assign \new_[7752]_  = ~\new_[12599]_  & (~\new_[8316]_  | ~\new_[8681]_ );
  assign \new_[7753]_  = ~\new_[12599]_  & (~\new_[8340]_  | ~\new_[8682]_ );
  assign \new_[7754]_  = ~\new_[12599]_  & (~\new_[8342]_  | ~\new_[8646]_ );
  assign \new_[7755]_  = ~\new_[12603]_  & (~\new_[8577]_  | ~\new_[8451]_ );
  assign \new_[7756]_  = ~\new_[12599]_  & (~\new_[8343]_  | ~\new_[8684]_ );
  assign \new_[7757]_  = ~\new_[12603]_  & (~\new_[8344]_  | ~\new_[8688]_ );
  assign \new_[7758]_  = ~\new_[12599]_  & (~\new_[8399]_  | ~\new_[8345]_ );
  assign \new_[7759]_  = ~\new_[12603]_  & (~\new_[8339]_  | ~\new_[8689]_ );
  assign \new_[7760]_  = ~\new_[12599]_  & (~\new_[8377]_  | ~\new_[8347]_ );
  assign \new_[7761]_  = ~\new_[12599]_  & (~\new_[8403]_  | ~\new_[8348]_ );
  assign \new_[7762]_  = ~\new_[12599]_  & (~\new_[8349]_  | ~\new_[8677]_ );
  assign \new_[7763]_  = ~\new_[12599]_  & (~\new_[8350]_  | ~\new_[8671]_ );
  assign \new_[7764]_  = ~\new_[12650]_  & (~\new_[8583]_  | ~\new_[8408]_ );
  assign \new_[7765]_  = ~\new_[12650]_  & (~\new_[8594]_  | ~\new_[8351]_ );
  assign \new_[7766]_  = ~\new_[12650]_  & (~\new_[8409]_  | ~\new_[8352]_ );
  assign \new_[7767]_  = ~\new_[14133]_  & (~\new_[8353]_  | ~\new_[8411]_ );
  assign \new_[7768]_  = ~\new_[8068]_  | (~\new_[8700]_  & ~\new_[13928]_ );
  assign \new_[7769]_  = ~\new_[8069]_  | (~\new_[8466]_  & ~\new_[13928]_ );
  assign \new_[7770]_  = ~\new_[8086]_  | (~\new_[8701]_  & ~\new_[13928]_ );
  assign \new_[7771]_  = ~\new_[8071]_  | (~\new_[8458]_  & ~\new_[13928]_ );
  assign \new_[7772]_  = ~\new_[8078]_  | (~\new_[8711]_  & ~\new_[13928]_ );
  assign \new_[7773]_  = ~\new_[8080]_  | (~\new_[8878]_  & ~\new_[12448]_ );
  assign \new_[7774]_  = \\u2_to_cnt_reg[5] ;
  assign \new_[7775]_  = ~\new_[8615]_  | (~\new_[8464]_  & ~\new_[12448]_ );
  assign \new_[7776]_  = ~\new_[8081]_  | (~\new_[8463]_  & ~\new_[12448]_ );
  assign \new_[7777]_  = ~\new_[8617]_  | (~\new_[8465]_  & ~\new_[12448]_ );
  assign int_o = u13_int_reg;
  assign \new_[7779]_  = ~\new_[8067]_  | (~\new_[8884]_  & ~\new_[12448]_ );
  assign \new_[7780]_  = ~\new_[8082]_  | (~\new_[8455]_  & ~\new_[12448]_ );
  assign \new_[7781]_  = ~\new_[8621]_  | (~\new_[8469]_  & ~\new_[12448]_ );
  assign \new_[7782]_  = ~\new_[8085]_  | (~\new_[8879]_  & ~\new_[12448]_ );
  assign \new_[7783]_  = ~\new_[8087]_  | (~\new_[8703]_  & ~\new_[12579]_ );
  assign \new_[7784]_  = ~\new_[8088]_  | (~\new_[8742]_  & ~\new_[12579]_ );
  assign \new_[7785]_  = ~\new_[8383]_  | (~\new_[8467]_  & ~\new_[12579]_ );
  assign \new_[7786]_  = ~\new_[8089]_  | (~\new_[8468]_  & ~\new_[12579]_ );
  assign \new_[7787]_  = ~\new_[8396]_  | (~\new_[8456]_  & ~\new_[13928]_ );
  assign \new_[7788]_  = ~\new_[8079]_  | (~\new_[8457]_  & ~\new_[13928]_ );
  assign \new_[7789]_  = \\u13_ints_r_reg[21] ;
  assign \new_[7790]_  = \\u1_slt3_reg[0] ;
  assign \new_[7791]_  = \\u13_ints_r_reg[0] ;
  assign \new_[7792]_  = \\u13_ints_r_reg[27] ;
  assign \new_[7793]_  = \\u13_ints_r_reg[15] ;
  assign \new_[7794]_  = ~\new_[8365]_  | (~\new_[8719]_  & ~\new_[12774]_ );
  assign \new_[7795]_  = ~\new_[12603]_  & (~\new_[8556]_  | ~\new_[8649]_ );
  assign \new_[7796]_  = ~\new_[8117]_  & ~\new_[13605]_ ;
  assign \new_[7797]_  = ~\new_[8118]_  & ~\new_[13223]_ ;
  assign \new_[7798]_  = ~\new_[8119]_  & ~\new_[13168]_ ;
  assign \new_[7799]_  = ~\new_[8120]_  & ~\new_[14093]_ ;
  assign \new_[7800]_  = ~\new_[10319]_  & ~\new_[8117]_ ;
  assign \new_[7801]_  = ~\new_[10318]_  & ~\new_[8118]_ ;
  assign \new_[7802]_  = ~\new_[10321]_  & ~\new_[8119]_ ;
  assign \new_[7803]_  = ~\new_[12086]_  & ~\new_[8120]_ ;
  assign \new_[7804]_  = ~\new_[8601]_  | (~\new_[8719]_  & ~\new_[12869]_ );
  assign \new_[7805]_  = ~\new_[7939]_ ;
  assign \new_[7806]_  = ~\new_[7940]_ ;
  assign \new_[7807]_  = \\u2_cnt_reg[7] ;
  assign \new_[7808]_  = \new_[12824]_  & \new_[8136]_ ;
  assign \new_[7809]_  = \new_[12844]_  & \new_[8135]_ ;
  assign \new_[7810]_  = ~\new_[8136]_  | ~\new_[13866]_ ;
  assign \new_[7811]_  = ~\new_[8135]_  | ~\new_[13873]_ ;
  assign \new_[7812]_  = ~\new_[10317]_  & ~\new_[8134]_ ;
  assign n9931 = n10226 ? \new_[9002]_  : \new_[7686]_ ;
  assign n9936 = n10226 ? \new_[9000]_  : \new_[7687]_ ;
  assign n9941 = n10226 ? \new_[9001]_  : \new_[7688]_ ;
  assign \new_[7816]_  = \\in_valid_s_reg[1] ;
  assign \new_[7817]_  = ~\new_[8100]_  & (~\new_[7492]_  | ~\new_[8804]_ );
  assign \new_[7818]_  = ~\new_[8148]_  & (~\new_[8806]_  | ~\new_[7493]_ );
  assign \new_[7819]_  = ~\new_[9797]_  & ~\new_[8413]_ ;
  assign \new_[7820]_  = ~\new_[8149]_  & (~\new_[7494]_  | ~\new_[8787]_ );
  assign \new_[7821]_  = ~\new_[8139]_  & ~\new_[8806]_ ;
  assign \new_[7822]_  = ~\new_[8138]_  & ~\new_[8787]_ ;
  assign \new_[7823]_  = ~\new_[8143]_  & (~\new_[8806]_  | ~\new_[7497]_ );
  assign \new_[7824]_  = ~\new_[8141]_  & (~\new_[7439]_  | ~\new_[8804]_ );
  assign \new_[7825]_  = ~\new_[8145]_  & (~\new_[7438]_  | ~\new_[8787]_ );
  assign n9926 = n10226 ? \new_[8996]_  : \new_[7656]_ ;
  assign \new_[7827]_  = ~\new_[8142]_  & (~\new_[8806]_  | ~\new_[7496]_ );
  assign \new_[7828]_  = ~\new_[8144]_  & (~\new_[13188]_  | ~\new_[8787]_ );
  assign \new_[7829]_  = ~\new_[8146]_  & (~\new_[7495]_  | ~\new_[8804]_ );
  assign n9916 = valid_s1_reg;
  assign n9921 = \\in_valid_s1_reg[0] ;
  assign \new_[7832]_  = ~\new_[8413]_  & (~\new_[8835]_  | ~\new_[9751]_ );
  assign \new_[7833]_  = ~\new_[8413]_  & (~\new_[8841]_  | ~\new_[9773]_ );
  assign \new_[7834]_  = ~\new_[8413]_  & (~\new_[8836]_  | ~\new_[9777]_ );
  assign \new_[7835]_  = ~\new_[8413]_  & (~\new_[8652]_  | ~\new_[9754]_ );
  assign \new_[7836]_  = ~\new_[8413]_  & (~\new_[8837]_  | ~\new_[9756]_ );
  assign \new_[7837]_  = ~\new_[8413]_  & (~\new_[8838]_  | ~\new_[9758]_ );
  assign \new_[7838]_  = ~\new_[8413]_  & (~\new_[8840]_  | ~\new_[9759]_ );
  assign \new_[7839]_  = ~\new_[8413]_  & (~\new_[8839]_  | ~\new_[10407]_ );
  assign \new_[7840]_  = ~\new_[12615]_  & (~\new_[8557]_  | ~\new_[8665]_ );
  assign \new_[7841]_  = ~\new_[14103]_  & (~\new_[8558]_  | ~\new_[8667]_ );
  assign \new_[7842]_  = ~\new_[14103]_  & (~\new_[8559]_  | ~\new_[8668]_ );
  assign \new_[7843]_  = ~\new_[12615]_  & (~\new_[8560]_  | ~\new_[8669]_ );
  assign \new_[7844]_  = ~\new_[12615]_  & (~\new_[8561]_  | ~\new_[8670]_ );
  assign \new_[7845]_  = ~\new_[14103]_  & (~\new_[8596]_  | ~\new_[8563]_ );
  assign \new_[7846]_  = ~\new_[12603]_  & (~\new_[8575]_  | ~\new_[8678]_ );
  assign \new_[7847]_  = ~\new_[12650]_  & (~\new_[8579]_  | ~\new_[8687]_ );
  assign \new_[7848]_  = ~\new_[12603]_  & (~\new_[8578]_  | ~\new_[8685]_ );
  assign \new_[7849]_  = ~\new_[12650]_  & (~\new_[8584]_  | ~\new_[8686]_ );
  assign \new_[7850]_  = ~\new_[12650]_  & (~\new_[8580]_  | ~\new_[8651]_ );
  assign \new_[7851]_  = ~\new_[12603]_  & (~\new_[8581]_  | ~\new_[8679]_ );
  assign \new_[7852]_  = ~\new_[12650]_  & (~\new_[8582]_  | ~\new_[8690]_ );
  assign \new_[7853]_  = ~\new_[8366]_  | (~\new_[8716]_  & ~\new_[12774]_ );
  assign \new_[7854]_  = ~\new_[12603]_  & (~\new_[8555]_  | ~\new_[8648]_ );
  assign \new_[7855]_  = (~\new_[8593]_  | ~\new_[13125]_ ) & (~\new_[3607]_  | ~\new_[12509]_ );
  assign \new_[7856]_  = (~\new_[12117]_  | ~\new_[9051]_ ) & (~\new_[8550]_  | ~\new_[10402]_ );
  assign \new_[7857]_  = \\u2_to_cnt_reg[3] ;
  assign \new_[7858]_  = ~\new_[8413]_  & ~\new_[9255]_ ;
  assign \new_[7859]_  = ~\new_[8413]_  & (~\new_[11458]_  | ~\new_[9761]_ );
  assign \new_[7860]_  = ~\new_[8413]_  & (~\new_[11460]_  | ~\new_[9253]_ );
  assign \new_[7861]_  = ~\new_[8413]_  & (~\new_[11461]_  | ~\new_[9763]_ );
  assign \new_[7862]_  = ~\new_[9794]_  & ~\new_[8413]_ ;
  assign \new_[7863]_  = ~\new_[8413]_  & (~\new_[11440]_  | ~\new_[9762]_ );
  assign \new_[7864]_  = ~\new_[8367]_  | (~\new_[8731]_  & ~\new_[13928]_ );
  assign \new_[7865]_  = \\u2_res_cnt_reg[3] ;
  assign \new_[7866]_  = ~\new_[8361]_  | (~\new_[8710]_  & ~\new_[13928]_ );
  assign \new_[7867]_  = ~\new_[8363]_  | (~\new_[8699]_  & ~\new_[13928]_ );
  assign \new_[7868]_  = ~\new_[8598]_  | (~\new_[8717]_  & ~\new_[12774]_ );
  assign \new_[7869]_  = ~\new_[8604]_  | (~\new_[8720]_  & ~\new_[12774]_ );
  assign \new_[7870]_  = ~\new_[8605]_  | (~\new_[8721]_  & ~\new_[12869]_ );
  assign \new_[7871]_  = ~\new_[8611]_  | (~\new_[8722]_  & ~\new_[12869]_ );
  assign \new_[7872]_  = ~\new_[8613]_  | (~\new_[8715]_  & ~\new_[12774]_ );
  assign \new_[7873]_  = ~\new_[8368]_  | (~\new_[8723]_  & ~\new_[12363]_ );
  assign \new_[7874]_  = \\u2_to_cnt_reg[4] ;
  assign \new_[7875]_  = \\u1_slt3_reg[2] ;
  assign \new_[7876]_  = \\u1_slt3_reg[1] ;
  assign \new_[7877]_  = \\u1_slt4_reg[1] ;
  assign \new_[7878]_  = \\u1_slt6_reg[1] ;
  assign \new_[7879]_  = \\u1_slt6_reg[2] ;
  assign wb_ack_o = u12_wb_ack_o_reg;
  assign \new_[7881]_  = \\u13_ints_r_reg[10] ;
  assign \new_[7882]_  = \\u13_ints_r_reg[12] ;
  assign \new_[7883]_  = \\u13_ints_r_reg[13] ;
  assign \new_[7884]_  = ~\new_[8370]_  | (~\new_[8883]_  & ~\new_[12448]_ );
  assign \new_[7885]_  = \\u13_ints_r_reg[16] ;
  assign \new_[7886]_  = \\u13_ints_r_reg[18] ;
  assign \new_[7887]_  = \\u13_ints_r_reg[19] ;
  assign \new_[7888]_  = \\u13_ints_r_reg[22] ;
  assign \new_[7889]_  = \\u13_ints_r_reg[24] ;
  assign \new_[7890]_  = \\u13_ints_r_reg[25] ;
  assign \new_[7891]_  = \\u13_ints_r_reg[28] ;
  assign \new_[7892]_  = \\u13_ints_r_reg[3] ;
  assign \new_[7893]_  = \\u13_ints_r_reg[4] ;
  assign \new_[7894]_  = \\u13_ints_r_reg[7] ;
  assign \new_[7895]_  = ~\new_[8619]_  | (~\new_[8727]_  & ~\new_[12448]_ );
  assign \new_[7896]_  = ~\new_[8623]_  | (~\new_[8730]_  & ~\new_[12448]_ );
  assign \new_[7897]_  = ~\new_[8378]_  | (~\new_[8738]_  & ~\new_[12579]_ );
  assign \new_[7898]_  = ~\new_[8379]_  | (~\new_[8896]_  & ~\new_[12579]_ );
  assign \new_[7899]_  = ~\new_[8380]_  | (~\new_[8739]_  & ~\new_[12579]_ );
  assign \new_[7900]_  = ~\new_[8369]_  | (~\new_[8759]_  & ~\new_[12579]_ );
  assign \new_[7901]_  = ~\new_[8381]_  | (~\new_[8740]_  & ~\new_[12579]_ );
  assign \new_[7902]_  = ~\new_[8382]_  | (~\new_[8741]_  & ~\new_[12579]_ );
  assign \new_[7903]_  = ~\new_[8387]_  | (~\new_[8737]_  & ~\new_[12854]_ );
  assign \new_[7904]_  = ~\new_[8388]_  | (~\new_[8738]_  & ~\new_[12854]_ );
  assign \new_[7905]_  = ~\new_[8390]_  | (~\new_[8746]_  & ~\new_[12363]_ );
  assign \new_[7906]_  = ~\new_[8391]_  | (~\new_[8749]_  & ~\new_[12363]_ );
  assign \new_[7907]_  = ~\new_[8636]_  | (~\new_[8755]_  & ~\new_[12665]_ );
  assign \new_[7908]_  = ~\new_[8393]_  | (~\new_[8735]_  & ~\new_[12363]_ );
  assign \new_[7909]_  = ~\new_[8358]_  | (~\new_[8753]_  & ~\new_[12363]_ );
  assign \new_[7910]_  = ~\new_[8638]_  | (~\new_[8764]_  & ~\new_[12665]_ );
  assign \new_[7911]_  = ~\new_[8395]_  | (~\new_[8917]_  & ~\new_[12665]_ );
  assign \new_[7912]_  = ~\new_[8400]_  | (~\new_[8762]_  & ~\new_[12363]_ );
  assign \new_[7913]_  = ~\new_[8401]_  | (~\new_[8922]_  & ~\new_[12665]_ );
  assign \new_[7914]_  = ~\new_[8402]_  | (~\new_[8751]_  & ~\new_[12363]_ );
  assign \new_[7915]_  = ~\new_[8404]_  | (~\new_[8757]_  & ~\new_[12363]_ );
  assign \new_[7916]_  = ~\new_[8375]_  | (~\new_[8758]_  & ~\new_[12665]_ );
  assign \new_[7917]_  = ~\new_[8405]_  | (~\new_[8732]_  & ~\new_[12363]_ );
  assign \new_[7918]_  = ~\new_[8407]_  | (~\new_[8747]_  & ~\new_[12363]_ );
  assign \new_[7919]_  = ~\new_[8643]_  | (~\new_[8761]_  & ~\new_[12665]_ );
  assign \new_[7920]_  = ~\new_[8592]_  | (~\new_[8714]_  & ~\new_[12665]_ );
  assign \new_[7921]_  = ~\new_[8359]_  | (~\new_[8847]_  & ~\new_[12665]_ );
  assign \new_[7922]_  = ~\new_[8355]_  | (~\new_[8932]_  & ~\new_[13169]_ );
  assign \new_[7923]_  = ~\new_[8415]_  | (~\new_[8722]_  & ~\new_[12774]_ );
  assign \new_[7924]_  = ~\new_[8356]_  | (~\new_[8713]_  & ~\new_[13928]_ );
  assign \new_[7925]_  = \\u13_ints_r_reg[6] ;
  assign \new_[7926]_  = \\u1_slt6_reg[3] ;
  assign \new_[7927]_  = \\u1_slt6_reg[0] ;
  assign \new_[7928]_  = \\u1_slt4_reg[3] ;
  assign \new_[7929]_  = \\u1_slt3_reg[3] ;
  assign \new_[7930]_  = \\u13_ints_r_reg[9] ;
  assign \new_[7931]_  = ~\new_[8413]_  & (~\new_[11459]_  | ~\new_[9252]_ );
  assign \new_[7932]_  = \\u1_slt4_reg[2] ;
  assign \new_[7933]_  = \\u1_slt4_reg[0] ;
  assign \new_[7934]_  = \new_[12627]_  | \new_[8483]_ ;
  assign \new_[7935]_  = \\u2_cnt_reg[1] ;
  assign \new_[7936]_  = \\u2_to_cnt_reg[2] ;
  assign \new_[7937]_  = ~\new_[8115]_ ;
  assign \new_[7938]_  = ~\new_[8117]_ ;
  assign \new_[7939]_  = \\u4_status_reg[1] ;
  assign \new_[7940]_  = \\u5_status_reg[1] ;
  assign \new_[7941]_  = ~\new_[8118]_ ;
  assign \new_[7942]_  = ~\new_[8119]_ ;
  assign \new_[7943]_  = ~\new_[8120]_ ;
  assign n9986 = ~\new_[8494]_  & ~\new_[9656]_ ;
  assign \new_[7945]_  = ~\new_[9677]_  & ~\new_[8488]_ ;
  assign \new_[7946]_  = ~\new_[9673]_  & ~\new_[8487]_ ;
  assign \new_[7947]_  = ~u12_rf_we_reg;
  assign \new_[7948]_  = ~\new_[8134]_ ;
  assign n9951 = ~\new_[8497]_  & ~\new_[12602]_ ;
  assign n9956 = ~\new_[12439]_  & ~\new_[8498]_ ;
  assign n9961 = ~\new_[8497]_  & ~\new_[12516]_ ;
  assign n9966 = ~\new_[8497]_  & ~\new_[12722]_ ;
  assign n9971 = ~\new_[8498]_  & ~\new_[12382]_ ;
  assign n9991 = ~\new_[12929]_  | ~\new_[8478]_  | ~\new_[12930]_ ;
  assign n9946 = ~\new_[8499]_  & ~\new_[12439]_ ;
  assign \new_[7956]_  = \\u2_res_cnt_reg[0] ;
  assign \new_[7957]_  = ~\new_[8495]_  & ~\new_[8804]_ ;
  assign n9981 = \\in_valid_s1_reg[2] ;
  assign n9976 = \\u1_sr_reg[5] ;
  assign \new_[7960]_  = \new_[8483]_  | \new_[13574]_ ;
  assign \new_[7961]_  = ~\new_[8618]_  | (~\new_[8882]_  & ~\new_[12448]_ );
  assign \new_[7962]_  = ~\new_[8116]_ ;
  assign \new_[7963]_  = ~\new_[8483]_  & (~\new_[13152]_  | ~\new_[12973]_ );
  assign \new_[7964]_  = (~\new_[12117]_  | ~\new_[9056]_ ) & (~\new_[8815]_  | ~\new_[10402]_ );
  assign \new_[7965]_  = \new_[13757]_  ^ \new_[8827]_ ;
  assign \new_[7966]_  = ~\new_[8147]_ ;
  assign \new_[7967]_  = ~\new_[8597]_  | (~\new_[8861]_  & ~\new_[12774]_ );
  assign \new_[7968]_  = ~\new_[8600]_  | (~\new_[8865]_  & ~\new_[12774]_ );
  assign \new_[7969]_  = ~\new_[8602]_  | (~\new_[8868]_  & ~\new_[12869]_ );
  assign \new_[7970]_  = ~\new_[8603]_  | (~\new_[8868]_  & ~\new_[12774]_ );
  assign \new_[7971]_  = ~\new_[8599]_  | (~\new_[8862]_  & ~\new_[12774]_ );
  assign \new_[7972]_  = \\u2_cnt_reg[4] ;
  assign \new_[7973]_  = \\u2_cnt_reg[3] ;
  assign \new_[7974]_  = \\u2_to_cnt_reg[0] ;
  assign \new_[7975]_  = \\u2_to_cnt_reg[1] ;
  assign \new_[7976]_  = \\u2_cnt_reg[5] ;
  assign \new_[7977]_  = \\u2_cnt_reg[6] ;
  assign \new_[7978]_  = \\u2_cnt_reg[0] ;
  assign \new_[7979]_  = \\u2_cnt_reg[2] ;
  assign sync_pad_o = \new_[4582]_  | \new_[8496]_ ;
  assign \new_[7981]_  = ~\new_[8624]_  | (~\new_[8887]_  & ~\new_[12448]_ );
  assign \new_[7982]_  = ~\new_[8625]_  | (~\new_[8888]_  & ~\new_[12448]_ );
  assign \new_[7983]_  = ~\new_[8614]_  | (~\new_[8877]_  & ~\new_[12448]_ );
  assign \new_[7984]_  = ~\new_[8635]_  | (~\new_[8896]_  & ~\new_[12854]_ );
  assign \new_[7985]_  = ~\new_[8637]_  | (~\new_[8916]_  & ~\new_[12665]_ );
  assign \new_[7986]_  = ~\new_[8640]_  | (~\new_[8920]_  & ~\new_[13037]_ );
  assign \new_[7987]_  = ~\new_[8639]_  | (~\new_[8924]_  & ~\new_[13037]_ );
  assign \new_[7988]_  = ~\new_[8630]_  | (~\new_[8910]_  & ~\new_[12665]_ );
  assign \new_[7989]_  = ~\new_[8641]_  | (~\new_[8891]_  & ~\new_[13037]_ );
  assign \new_[7990]_  = ~\new_[8591]_  | (~\new_[8928]_  & ~\new_[12665]_ );
  assign \new_[7991]_  = ~\new_[8644]_  | (~\new_[8929]_  & ~\new_[13037]_ );
  assign \new_[7992]_  = ~\new_[8589]_  | (~\new_[8858]_  & ~\new_[12665]_ );
  assign \new_[7993]_  = ~\new_[8650]_  & (~\new_[10819]_  | ~\new_[13012]_ );
  assign \new_[7994]_  = ~\new_[8647]_  & (~\new_[10819]_  | ~\new_[4902]_ );
  assign \new_[7995]_  = ~\new_[8672]_  & (~\new_[10819]_  | ~\new_[5078]_ );
  assign \new_[7996]_  = ~\new_[8674]_  & (~\new_[10819]_  | ~\new_[5756]_ );
  assign \new_[7997]_  = ~\new_[8653]_  & (~\new_[10819]_  | ~\new_[5041]_ );
  assign \new_[7998]_  = ~\new_[8655]_  & (~\new_[10819]_  | ~\new_[5094]_ );
  assign \new_[7999]_  = ~\new_[8656]_  & (~\new_[10819]_  | ~\new_[5042]_ );
  assign \new_[8000]_  = ~\new_[8657]_  & (~\new_[10819]_  | ~\new_[5095]_ );
  assign \new_[8001]_  = ~\new_[8658]_  & (~\new_[10819]_  | ~\new_[5096]_ );
  assign \new_[8002]_  = ~\new_[8659]_  & (~\new_[10819]_  | ~\new_[5097]_ );
  assign \new_[8003]_  = ~\new_[8660]_  & (~\new_[10819]_  | ~\new_[12886]_ );
  assign \new_[8004]_  = ~\new_[8661]_  & (~\new_[10819]_  | ~\new_[5098]_ );
  assign \new_[8005]_  = ~\new_[8676]_  & (~\new_[10819]_  | ~\new_[5077]_ );
  assign \new_[8006]_  = ~\new_[8654]_  & (~\new_[10819]_  | ~\new_[5076]_ );
  assign \new_[8007]_  = ~\new_[8662]_  & (~\new_[10819]_  | ~\new_[5079]_ );
  assign \new_[8008]_  = \new_[13583]_  ? \new_[12733]_  : \new_[8942]_ ;
  assign \new_[8009]_  = \new_[13409]_  ? \new_[12662]_  : \new_[8935]_ ;
  assign \new_[8010]_  = \new_[8935]_  ? \new_[12434]_  : \new_[13346]_ ;
  assign \new_[8011]_  = \new_[13819]_  ? \new_[12889]_  : \new_[8933]_ ;
  assign \new_[8012]_  = \new_[13638]_  ? \new_[12662]_  : \new_[8938]_ ;
  assign \new_[8013]_  = \new_[13845]_  ? \new_[12733]_  : \new_[8941]_ ;
  assign \new_[8014]_  = \new_[13420]_  ? \new_[12733]_  : \new_[8939]_ ;
  assign \new_[8015]_  = \new_[13246]_  ? \new_[12662]_  : \new_[8940]_ ;
  assign \new_[8016]_  = \new_[13453]_  ? \new_[12662]_  : \new_[8937]_ ;
  assign \new_[8017]_  = \new_[13830]_  ? \new_[12578]_  : \new_[8935]_ ;
  assign \new_[8018]_  = \new_[13406]_  ? \new_[12967]_  : \new_[8934]_ ;
  assign \new_[8019]_  = \new_[13544]_  ? \new_[12967]_  : \new_[8943]_ ;
  assign \new_[8020]_  = \new_[13591]_  ? \new_[12578]_  : \new_[8940]_ ;
  assign \new_[8021]_  = \new_[8942]_  ? \new_[12513]_  : \new_[13800]_ ;
  assign \new_[8022]_  = \new_[8936]_  ? \new_[12434]_  : \new_[13690]_ ;
  assign \new_[8023]_  = \new_[8933]_  ? \new_[12434]_  : \new_[13512]_ ;
  assign \new_[8024]_  = ~\new_[8616]_  | (~\new_[8881]_  & ~\new_[12448]_ );
  assign \new_[8025]_  = \new_[8934]_  ? \new_[12434]_  : \new_[13746]_ ;
  assign \new_[8026]_  = \new_[8941]_  ? \new_[12434]_  : \new_[13268]_ ;
  assign \new_[8027]_  = \new_[8940]_  ? \new_[12434]_  : \new_[13637]_ ;
  assign \new_[8028]_  = \new_[8937]_  ? \new_[12434]_  : \new_[13376]_ ;
  assign \new_[8029]_  = \new_[13499]_  ? \new_[12578]_  : \new_[8941]_ ;
  assign \new_[8030]_  = \new_[13310]_  ? \new_[12578]_  : \new_[8939]_ ;
  assign \new_[8031]_  = \new_[8943]_  ? \new_[12434]_  : \new_[13216]_ ;
  assign \new_[8032]_  = \new_[13699]_  ? \new_[12578]_  : \new_[8937]_ ;
  assign \new_[8033]_  = \new_[8938]_  ? \new_[12434]_  : \new_[13290]_ ;
  assign \new_[8034]_  = \new_[13542]_  ? \new_[12967]_  : \new_[8938]_ ;
  assign \new_[8035]_  = \new_[8939]_  ? \new_[12434]_  : \new_[13386]_ ;
  assign \new_[8036]_  = \new_[13628]_  ? \new_[12662]_  : \new_[8936]_ ;
  assign \new_[8037]_  = \new_[13521]_  ? \new_[12578]_  : \new_[8933]_ ;
  assign \new_[8038]_  = \new_[13436]_  ? \new_[12662]_  : \new_[8934]_ ;
  assign \new_[8039]_  = \new_[13439]_  ? \new_[12889]_  : \new_[8943]_ ;
  assign \new_[8040]_  = \new_[13333]_  ? \new_[12578]_  : \new_[8936]_ ;
  assign \new_[8041]_  = \new_[13663]_  ? \new_[12578]_  : \new_[8942]_ ;
  assign \new_[8042]_  = \new_[13479]_  ? \new_[12027]_  : \new_[8942]_ ;
  assign \new_[8043]_  = \new_[13517]_  ? \new_[12027]_  : \new_[8936]_ ;
  assign \new_[8044]_  = \new_[13848]_  ? \new_[12027]_  : \new_[8935]_ ;
  assign \new_[8045]_  = \new_[13432]_  ? \new_[12027]_  : \new_[8933]_ ;
  assign \new_[8046]_  = \new_[13504]_  ? \new_[12027]_  : \new_[8934]_ ;
  assign \new_[8047]_  = \new_[13774]_  ? \new_[12027]_  : \new_[8938]_ ;
  assign \new_[8048]_  = \new_[13485]_  ? \new_[12027]_  : \new_[8943]_ ;
  assign \new_[8049]_  = \new_[13400]_  ? \new_[12027]_  : \new_[8941]_ ;
  assign \new_[8050]_  = \new_[13842]_  ? \new_[12027]_  : \new_[8939]_ ;
  assign \new_[8051]_  = \new_[13202]_  ? \new_[12027]_  : \new_[8940]_ ;
  assign \new_[8052]_  = \new_[13862]_  ? \new_[12027]_  : \new_[8937]_ ;
  assign \new_[8053]_  = ~\new_[8587]_  | (~\new_[9156]_  & ~\new_[13105]_ );
  assign \new_[8054]_  = ~\new_[8588]_  | (~\new_[9154]_  & ~\new_[13127]_ );
  assign \new_[8055]_  = ~\new_[8586]_  | (~\new_[9153]_  & ~\new_[4763]_ );
  assign \new_[8056]_  = ~\new_[8702]_  | ~\new_[13622]_ ;
  assign \new_[8057]_  = ~\new_[14008]_  | ~\new_[13622]_ ;
  assign \new_[8058]_  = ~\new_[8708]_  | ~\new_[13622]_ ;
  assign \new_[8059]_  = ~\new_[8709]_  | ~\new_[13677]_ ;
  assign \new_[8060]_  = ~\new_[13794]_  | ~\new_[13963]_ ;
  assign \new_[8061]_  = ~\new_[14167]_  | ~\new_[13622]_ ;
  assign \new_[8062]_  = ~\new_[8725]_  | ~\new_[13794]_ ;
  assign \new_[8063]_  = ~\new_[8726]_  | ~\new_[13794]_ ;
  assign \new_[8064]_  = ~\new_[8763]_  | ~\new_[13794]_ ;
  assign \new_[8065]_  = ~\new_[8733]_  | ~\new_[13622]_ ;
  assign \new_[8066]_  = ~\new_[13925]_  | ~\new_[13622]_ ;
  assign \new_[8067]_  = ~\new_[8698]_  | ~\new_[12591]_ ;
  assign \new_[8068]_  = ~\new_[8733]_  | ~\new_[14081]_ ;
  assign \new_[8069]_  = ~\new_[14167]_  | ~\new_[14081]_ ;
  assign \new_[8070]_  = ~\new_[8705]_  | ~\new_[14081]_ ;
  assign \new_[8071]_  = ~\new_[8706]_  | ~\new_[14081]_ ;
  assign \new_[8072]_  = ~\new_[8708]_  | ~\new_[14081]_ ;
  assign \new_[8073]_  = ~\new_[8724]_  | ~\new_[14010]_ ;
  assign \new_[8074]_  = ~\new_[8707]_  | ~\new_[14010]_ ;
  assign \new_[8075]_  = ~\new_[8709]_  | ~\new_[14081]_ ;
  assign \new_[8076]_  = ~\new_[8705]_  | ~\new_[3023]_ ;
  assign \new_[8077]_  = ~\new_[8706]_  | ~\new_[3023]_ ;
  assign \new_[8078]_  = ~\new_[13925]_  | ~\new_[14081]_ ;
  assign \new_[8079]_  = ~\new_[14081]_  | ~\new_[8704]_ ;
  assign \new_[8080]_  = ~\new_[13963]_  | ~\new_[12591]_ ;
  assign \new_[8081]_  = ~\new_[8726]_  | ~\new_[12591]_ ;
  assign \new_[8082]_  = ~\new_[8728]_  | ~\new_[12591]_ ;
  assign \new_[8083]_  = ~\new_[8763]_  | ~\new_[12591]_ ;
  assign \new_[8084]_  = ~\new_[8728]_  | ~\new_[13154]_ ;
  assign \new_[8085]_  = ~\new_[8725]_  | ~\new_[12591]_ ;
  assign \new_[8086]_  = ~\new_[14081]_  | ~\new_[8702]_ ;
  assign \new_[8087]_  = ~\new_[12544]_  | ~\new_[8743]_ ;
  assign \new_[8088]_  = ~\new_[12544]_  | ~\new_[8756]_ ;
  assign \new_[8089]_  = ~\new_[14038]_  | ~\new_[12544]_ ;
  assign \new_[8090]_  = ~\new_[8698]_  | ~\new_[13154]_ ;
  assign \new_[8091]_  = ~\new_[8734]_  | ~\new_[12717]_ ;
  assign n10136 = ~\new_[13019]_  & ~\new_[8829]_ ;
  assign n10131 = ~\new_[12903]_  & ~\new_[8829]_ ;
  assign \new_[8094]_  = \new_[13723]_  ^ \new_[9078]_ ;
  assign n10011 = ~\new_[13099]_  & ~\new_[8829]_ ;
  assign n10126 = ~\new_[13024]_  & ~\new_[8829]_ ;
  assign n9996 = ~\new_[13138]_  & ~\new_[8829]_ ;
  assign n10121 = ~\new_[13107]_  & ~\new_[8829]_ ;
  assign \new_[8099]_  = \\u2_res_cnt_reg[2] ;
  assign \new_[8100]_  = ~\new_[8804]_  & (~\new_[12906]_  | ~\new_[13056]_ );
  assign n10116 = ~\new_[12916]_  & ~\new_[8829]_ ;
  assign n10111 = ~\new_[13045]_  & ~\new_[9661]_ ;
  assign n10101 = ~\new_[12960]_  & ~\new_[8829]_ ;
  assign \new_[8104]_  = (~\new_[12117]_  | ~\new_[9047]_ ) & (~\new_[9009]_  | ~\new_[9784]_ );
  assign n10016 = ~\new_[12984]_  & ~\new_[8829]_ ;
  assign \new_[8106]_  = (~\new_[12117]_  | ~\new_[9062]_ ) & (~\new_[9024]_  | ~\new_[9784]_ );
  assign n10091 = ~\new_[12974]_  & ~\new_[9661]_ ;
  assign n10096 = ~\new_[13033]_  & ~\new_[9661]_ ;
  assign n10086 = ~\new_[12963]_  & ~\new_[8829]_ ;
  assign n10006 = ~\new_[12721]_  & ~\new_[8829]_ ;
  assign n10031 = u2_valid_reg;
  assign \new_[8112]_  = (~\new_[12117]_  | ~\new_[9061]_ ) & (~\new_[9023]_  | ~\new_[9784]_ );
  assign \new_[8113]_  = (~\new_[12117]_  | ~\new_[9060]_ ) & (~\new_[9022]_  | ~\new_[9784]_ );
  assign \new_[8114]_  = \\u2_res_cnt_reg[1] ;
  assign \new_[8115]_  = ~\new_[8788]_ ;
  assign \new_[8116]_  = ~\new_[8483]_ ;
  assign \new_[8117]_  = \\u3_status_reg[1] ;
  assign \new_[8118]_  = \\u6_status_reg[1] ;
  assign \new_[8119]_  = \\u7_status_reg[1] ;
  assign \new_[8120]_  = \\u8_status_reg[1] ;
  assign n10051 = ~\new_[8802]_  & ~\new_[9656]_ ;
  assign n10061 = n10976 ? \new_[9002]_  : \new_[7876]_ ;
  assign n10001 = n11071 ? \new_[9002]_  : \new_[7790]_ ;
  assign n10056 = n10671 ? \new_[9002]_  : \new_[7875]_ ;
  assign n10171 = n10336 ? \new_[9002]_  : \new_[7929]_ ;
  assign n10186 = n11071 ? \new_[9000]_  : \new_[7933]_ ;
  assign n10066 = n10976 ? \new_[9000]_  : \new_[7877]_ ;
  assign n10181 = n10671 ? \new_[9000]_  : \new_[7932]_ ;
  assign n10166 = n10336 ? \new_[9000]_  : \new_[7928]_ ;
  assign n10161 = n11071 ? \new_[9001]_  : \new_[7927]_ ;
  assign n10071 = n10976 ? \new_[9001]_  : \new_[7878]_ ;
  assign n10076 = n10671 ? \new_[9001]_  : \new_[7879]_ ;
  assign n10156 = n10336 ? \new_[9001]_  : \new_[7926]_ ;
  assign \new_[8134]_  = \\u11_status_reg[1] ;
  assign \new_[8135]_  = ~\new_[8487]_ ;
  assign \new_[8136]_  = ~\new_[8488]_ ;
  assign n10081 = ~\new_[8491]_ ;
  assign \new_[8138]_  = ~u10_empty_reg;
  assign \new_[8139]_  = ~u9_empty_reg;
  assign n10026 = \\in_valid_s1_reg[1] ;
  assign \new_[8141]_  = ~\new_[12641]_  & ~\new_[8804]_ ;
  assign \new_[8142]_  = ~\new_[8806]_  & ~\new_[7496]_ ;
  assign \new_[8143]_  = ~\new_[12630]_  & ~\new_[8806]_ ;
  assign \new_[8144]_  = ~\new_[13188]_  & ~\new_[8787]_ ;
  assign \new_[8145]_  = ~\new_[12666]_  & ~\new_[8787]_ ;
  assign \new_[8146]_  = ~\new_[7495]_  & ~\new_[8804]_ ;
  assign \new_[8147]_  = ~\new_[8501]_ ;
  assign \new_[8148]_  = ~\new_[8806]_  & (~\new_[12945]_  | ~\new_[13059]_ );
  assign \new_[8149]_  = ~\new_[8787]_  & (~\new_[12864]_  | ~\new_[12707]_ );
  assign \new_[8150]_  = (~\new_[12117]_  | ~\new_[9037]_ ) & (~\new_[9073]_  | ~\new_[9784]_ );
  assign \new_[8151]_  = (~\new_[12117]_  | ~\new_[9039]_ ) & (~\new_[9007]_  | ~\new_[9784]_ );
  assign \new_[8152]_  = (~\new_[12117]_  | ~\new_[9043]_ ) & (~\new_[9008]_  | ~\new_[9784]_ );
  assign \new_[8153]_  = (~\new_[12117]_  | ~\new_[9044]_ ) & (~\new_[9071]_  | ~\new_[9784]_ );
  assign \new_[8154]_  = (~\new_[12117]_  | ~\new_[9048]_ ) & (~\new_[9010]_  | ~\new_[9784]_ );
  assign \new_[8155]_  = (~\new_[12117]_  | ~\new_[9054]_ ) & (~\new_[9014]_  | ~\new_[9784]_ );
  assign \new_[8156]_  = (~\new_[12117]_  | ~\new_[9057]_ ) & (~\new_[9019]_  | ~\new_[9784]_ );
  assign \new_[8157]_  = (~\new_[12117]_  | ~\new_[9058]_ ) & (~\new_[9020]_  | ~\new_[9784]_ );
  assign \new_[8158]_  = (~\new_[12117]_  | ~\new_[9059]_ ) & (~\new_[9021]_  | ~\new_[9784]_ );
  assign \new_[8159]_  = (~\new_[12117]_  | ~\new_[9063]_ ) & (~\new_[9025]_  | ~\new_[9784]_ );
  assign \new_[8160]_  = (~\new_[12117]_  | ~\new_[9064]_ ) & (~\new_[9026]_  | ~\new_[9784]_ );
  assign \new_[8161]_  = (~\new_[12117]_  | ~\new_[9053]_ ) & (~\new_[9013]_  | ~\new_[9784]_ );
  assign \new_[8162]_  = (~\new_[12117]_  | ~\new_[9065]_ ) & (~\new_[9028]_  | ~\new_[9784]_ );
  assign \new_[8163]_  = (~\new_[12117]_  | ~\new_[9066]_ ) & (~\new_[9029]_  | ~\new_[9784]_ );
  assign \new_[8164]_  = (~\new_[12117]_  | ~\new_[9052]_ ) & (~\new_[9012]_  | ~\new_[9784]_ );
  assign \new_[8165]_  = (~\new_[12117]_  | ~\new_[9068]_ ) & (~\new_[9031]_  | ~\new_[9784]_ );
  assign \new_[8166]_  = (~\new_[12117]_  | ~\new_[9069]_ ) & (~\new_[9032]_  | ~\new_[9784]_ );
  assign \new_[8167]_  = (~\new_[12117]_  | ~\new_[9070]_ ) & (~\new_[9784]_  | ~\new_[9033]_ );
  assign \new_[8168]_  = (~\new_[12117]_  | ~\new_[9050]_ ) & (~\new_[9076]_  | ~\new_[9784]_ );
  assign \new_[8169]_  = (~\new_[12117]_  | ~\new_[9046]_ ) & (~\new_[9072]_  | ~\new_[9784]_ );
  assign \new_[8170]_  = (~\new_[12117]_  | ~\new_[9040]_ ) & (~\new_[9074]_  | ~\new_[9784]_ );
  assign \new_[8171]_  = (~\new_[12117]_  | ~\new_[9041]_ ) & (~\new_[9036]_  | ~\new_[9784]_ );
  assign \new_[8172]_  = (~\new_[12117]_  | ~\new_[9038]_ ) & (~\new_[9075]_  | ~\new_[9784]_ );
  assign \new_[8173]_  = (~\new_[12117]_  | ~\new_[9045]_ ) & (~\new_[9018]_  | ~\new_[10402]_ );
  assign \new_[8174]_  = (~\new_[12117]_  | ~\new_[9055]_ ) & (~\new_[9034]_  | ~\new_[10402]_ );
  assign n10106 = ~\new_[13022]_  & ~\new_[8829]_ ;
  assign n10036 = \\u2_in_valid_reg[0] ;
  assign n10141 = ~\new_[12922]_  & ~\new_[8829]_ ;
  assign \new_[8178]_  = \new_[13837]_  ? \new_[12758]_  : \new_[9174]_ ;
  assign \new_[8179]_  = \new_[13273]_  ? \new_[12951]_  : \new_[9167]_ ;
  assign \new_[8180]_  = \new_[13711]_  ? \new_[12574]_  : \new_[9168]_ ;
  assign \new_[8181]_  = \new_[13414]_  ? \new_[12574]_  : \new_[9169]_ ;
  assign \new_[8182]_  = \new_[13766]_  ? \new_[12574]_  : \new_[9177]_ ;
  assign \new_[8183]_  = \new_[13232]_  ? \new_[12574]_  : \new_[9172]_ ;
  assign \new_[8184]_  = \new_[9182]_  ? \new_[12828]_  : \new_[13304]_ ;
  assign \new_[8185]_  = \new_[13514]_  ? \new_[12662]_  : \new_[9164]_ ;
  assign \new_[8186]_  = \new_[13577]_  ? \new_[12662]_  : \new_[9160]_ ;
  assign \new_[8187]_  = \new_[13722]_  ? \new_[12574]_  : \new_[9185]_ ;
  assign \new_[8188]_  = \new_[9184]_  ? \new_[12828]_  : \new_[13348]_ ;
  assign \new_[8189]_  = \new_[13586]_  ? \new_[12967]_  : \new_[9164]_ ;
  assign \new_[8190]_  = \new_[13284]_  ? \new_[12578]_  : \new_[9163]_ ;
  assign \new_[8191]_  = \new_[13621]_  ? \new_[12578]_  : \new_[9161]_ ;
  assign \new_[8192]_  = \new_[13679]_  ? \new_[12578]_  : \new_[9160]_ ;
  assign \new_[8193]_  = \new_[13257]_  ? \new_[12578]_  : \new_[9159]_ ;
  assign \new_[8194]_  = \new_[13858]_  ? \new_[12574]_  : \new_[9157]_ ;
  assign \new_[8195]_  = \new_[13553]_  ? \new_[12574]_  : \new_[9186]_ ;
  assign \new_[8196]_  = \new_[13713]_  ? \new_[12578]_  : \new_[9158]_ ;
  assign \new_[8197]_  = \new_[9183]_  ? \new_[12828]_  : \new_[13342]_ ;
  assign \new_[8198]_  = \new_[13806]_  ? \new_[12574]_  : \new_[9187]_ ;
  assign \new_[8199]_  = \new_[9164]_  ? \new_[12434]_  : \new_[13362]_ ;
  assign \new_[8200]_  = \new_[9163]_  ? \new_[12434]_  : \new_[13468]_ ;
  assign \new_[8201]_  = \new_[9162]_  ? \new_[12434]_  : \new_[13328]_ ;
  assign \new_[8202]_  = \new_[13240]_  ? \new_[12574]_  : \new_[9188]_ ;
  assign \new_[8203]_  = \new_[13750]_  ? \new_[12951]_  : \new_[9166]_ ;
  assign \new_[8204]_  = \new_[13340]_  ? \new_[12574]_  : \new_[9189]_ ;
  assign \new_[8205]_  = \new_[9173]_  ? \new_[12828]_  : \new_[13814]_ ;
  assign \new_[8206]_  = \new_[9166]_  ? \new_[12432]_  : \new_[13267]_ ;
  assign \new_[8207]_  = \new_[9167]_  ? \new_[12432]_  : \new_[13226]_ ;
  assign \new_[8208]_  = \new_[9168]_  ? \new_[12432]_  : \new_[13215]_ ;
  assign \new_[8209]_  = \new_[9169]_  ? \new_[12432]_  : \new_[13443]_ ;
  assign \new_[8210]_  = \new_[9177]_  ? \new_[12432]_  : \new_[13640]_ ;
  assign \new_[8211]_  = \new_[9172]_  ? \new_[12432]_  : \new_[13644]_ ;
  assign \new_[8212]_  = \new_[9159]_  ? \new_[12434]_  : \new_[13528]_ ;
  assign \new_[8213]_  = \new_[9185]_  ? \new_[12432]_  : \new_[13590]_ ;
  assign \new_[8214]_  = \new_[9157]_  ? \new_[12432]_  : \new_[13557]_ ;
  assign \new_[8215]_  = \new_[9186]_  ? \new_[12432]_  : \new_[13536]_ ;
  assign \new_[8216]_  = \new_[9187]_  ? \new_[12432]_  : \new_[13498]_ ;
  assign \new_[8217]_  = \new_[9188]_  ? \new_[12432]_  : \new_[13487]_ ;
  assign \new_[8218]_  = \new_[9189]_  ? \new_[12432]_  : \new_[13502]_ ;
  assign \new_[8219]_  = \new_[9158]_  ? \new_[12513]_  : \new_[13381]_ ;
  assign \new_[8220]_  = \new_[9181]_  ? \new_[12828]_  : \new_[13274]_ ;
  assign \new_[8221]_  = \new_[9170]_  ? \new_[12828]_  : \new_[13631]_ ;
  assign \new_[8222]_  = \new_[13494]_  ? \new_[12662]_  : \new_[9163]_ ;
  assign \new_[8223]_  = \new_[13752]_  ? \new_[12996]_  : \new_[9183]_ ;
  assign \new_[8224]_  = \new_[13345]_  ? \new_[12626]_  : \new_[9181]_ ;
  assign \new_[8225]_  = \new_[13195]_  ? \new_[12924]_  : \new_[9186]_ ;
  assign \new_[8226]_  = \new_[13318]_  ? \new_[12662]_  : \new_[9162]_ ;
  assign \new_[8227]_  = \new_[13717]_  ? \new_[12733]_  : \new_[9158]_ ;
  assign \new_[8228]_  = \new_[13762]_  ? \new_[12663]_  : \new_[9177]_ ;
  assign \new_[8229]_  = \new_[13675]_  ? \new_[12662]_  : \new_[9161]_ ;
  assign \new_[8230]_  = \new_[13777]_  ? \new_[12642]_  : \new_[9183]_ ;
  assign \new_[8231]_  = \new_[13294]_  ? \new_[12662]_  : \new_[9159]_ ;
  assign \new_[8232]_  = \new_[13397]_  ? \new_[12663]_  : \new_[9185]_ ;
  assign \new_[8233]_  = \new_[9178]_  ? \new_[12828]_  : \new_[13265]_ ;
  assign \new_[8234]_  = \new_[13696]_  ? \new_[12626]_  : \new_[9170]_ ;
  assign \new_[8235]_  = \new_[13751]_  ? \new_[12626]_  : \new_[9171]_ ;
  assign \new_[8236]_  = \new_[13843]_  ? \new_[12626]_  : \new_[9165]_ ;
  assign \new_[8237]_  = \new_[13736]_  ? \new_[12626]_  : \new_[9173]_ ;
  assign \new_[8238]_  = \new_[13737]_  ? \new_[12996]_  : \new_[9174]_ ;
  assign \new_[8239]_  = \new_[13423]_  ? \new_[12996]_  : \new_[9175]_ ;
  assign \new_[8240]_  = \new_[9160]_  ? \new_[12434]_  : \new_[13329]_ ;
  assign \new_[8241]_  = \new_[13390]_  ? \new_[12626]_  : \new_[9190]_ ;
  assign \new_[8242]_  = \new_[13426]_  ? \new_[12626]_  : \new_[9176]_ ;
  assign \new_[8243]_  = \new_[13430]_  ? \new_[12626]_  : \new_[9178]_ ;
  assign \new_[8244]_  = \new_[13854]_  ? \new_[12578]_  : \new_[9162]_ ;
  assign \new_[8245]_  = \new_[13431]_  ? \new_[12996]_  : \new_[9179]_ ;
  assign \new_[8246]_  = \new_[13367]_  ? \new_[12626]_  : \new_[9180]_ ;
  assign \new_[8247]_  = \new_[13510]_  ? \new_[12626]_  : \new_[9182]_ ;
  assign \new_[8248]_  = \new_[13440]_  ? \new_[12626]_  : \new_[9184]_ ;
  assign \new_[8249]_  = \new_[13754]_  ? \new_[12642]_  : \new_[9170]_ ;
  assign \new_[8250]_  = \new_[13646]_  ? \new_[12642]_  : \new_[9171]_ ;
  assign \new_[8251]_  = \new_[13446]_  ? \new_[12663]_  : \new_[9166]_ ;
  assign \new_[8252]_  = \new_[13448]_  ? \new_[12642]_  : \new_[9165]_ ;
  assign \new_[8253]_  = \new_[13840]_  ? \new_[12758]_  : \new_[9173]_ ;
  assign \new_[8254]_  = \new_[13224]_  ? \new_[12837]_  : \new_[9167]_ ;
  assign \new_[8255]_  = \new_[13664]_  ? \new_[12758]_  : \new_[9175]_ ;
  assign \new_[8256]_  = \new_[13667]_  ? \new_[12837]_  : \new_[9168]_ ;
  assign \new_[8257]_  = \new_[13580]_  ? \new_[12642]_  : \new_[9190]_ ;
  assign \new_[8258]_  = \new_[13760]_  ? \new_[12663]_  : \new_[9169]_ ;
  assign \new_[8259]_  = \new_[13613]_  ? \new_[13013]_  : \new_[9176]_ ;
  assign \new_[8260]_  = \new_[13786]_  ? \new_[12663]_  : \new_[9172]_ ;
  assign \new_[8261]_  = \new_[9161]_  ? \new_[12434]_  : \new_[13327]_ ;
  assign \new_[8262]_  = \new_[13556]_  ? \new_[13013]_  : \new_[9178]_ ;
  assign \new_[8263]_  = \new_[13476]_  ? \new_[12642]_  : \new_[9179]_ ;
  assign \new_[8264]_  = \new_[9180]_  ? \new_[12828]_  : \new_[13351]_ ;
  assign \new_[8265]_  = \new_[13623]_  ? \new_[12758]_  : \new_[9180]_ ;
  assign \new_[8266]_  = \new_[13768]_  ? \new_[12642]_  : \new_[9181]_ ;
  assign \new_[8267]_  = \new_[13772]_  ? \new_[12642]_  : \new_[9182]_ ;
  assign \new_[8268]_  = \new_[13192]_  ? \new_[12642]_  : \new_[9184]_ ;
  assign \new_[8269]_  = \new_[9171]_  ? \new_[12828]_  : \new_[13684]_ ;
  assign \new_[8270]_  = \new_[9165]_  ? \new_[12828]_  : \new_[13782]_ ;
  assign \new_[8271]_  = \new_[9174]_  ? \new_[12828]_  : \new_[13807]_ ;
  assign \new_[8272]_  = \new_[9175]_  ? \new_[12828]_  : \new_[13630]_ ;
  assign \new_[8273]_  = \new_[9190]_  ? \new_[12828]_  : \new_[13662]_ ;
  assign \new_[8274]_  = \new_[9179]_  ? \new_[12828]_  : \new_[13821]_ ;
  assign \new_[8275]_  = \new_[13784]_  ? \new_[12837]_  : \new_[9157]_ ;
  assign \new_[8276]_  = \new_[9176]_  ? \new_[12828]_  : \new_[13635]_ ;
  assign \new_[8277]_  = \new_[13250]_  ? \new_[12924]_  : \new_[9187]_ ;
  assign \new_[8278]_  = \new_[13513]_  ? \new_[12663]_  : \new_[9188]_ ;
  assign \new_[8279]_  = \new_[13653]_  ? \new_[12663]_  : \new_[9189]_ ;
  assign \new_[8280]_  = \new_[13312]_  ? \new_[12027]_  : \new_[9164]_ ;
  assign \new_[8281]_  = \new_[13410]_  ? \new_[12027]_  : \new_[9163]_ ;
  assign \new_[8282]_  = \new_[13527]_  ? \new_[12027]_  : \new_[9162]_ ;
  assign \new_[8283]_  = \new_[13256]_  ? \new_[12027]_  : \new_[9160]_ ;
  assign \new_[8284]_  = \new_[13356]_  ? \new_[12027]_  : \new_[9159]_ ;
  assign \new_[8285]_  = \new_[13497]_  ? \new_[12027]_  : \new_[9158]_ ;
  assign \new_[8286]_  = \new_[13222]_  ? \new_[12027]_  : \new_[9161]_ ;
  assign \new_[8287]_  = \new_[13530]_  ? \new_[12028]_  : \new_[9172]_ ;
  assign \new_[8288]_  = \new_[13682]_  ? \new_[12030]_  : \new_[9176]_ ;
  assign \new_[8289]_  = \new_[13355]_  ? \new_[12028]_  : \new_[9166]_ ;
  assign \new_[8290]_  = \new_[13296]_  ? \new_[12028]_  : \new_[9167]_ ;
  assign \new_[8291]_  = \new_[13533]_  ? \new_[12028]_  : \new_[9168]_ ;
  assign \new_[8292]_  = \new_[13213]_  ? \new_[12028]_  : \new_[9169]_ ;
  assign \new_[8293]_  = \new_[13658]_  ? \new_[12030]_  : \new_[9170]_ ;
  assign \new_[8294]_  = \new_[13524]_  ? \new_[12028]_  : \new_[9177]_ ;
  assign \new_[8295]_  = \new_[13674]_  ? \new_[12030]_  : \new_[9171]_ ;
  assign \new_[8296]_  = \new_[13686]_  ? \new_[12030]_  : \new_[9165]_ ;
  assign \new_[8297]_  = \new_[13212]_  ? \new_[12030]_  : \new_[9173]_ ;
  assign \new_[8298]_  = \new_[13742]_  ? \new_[12030]_  : \new_[9174]_ ;
  assign \new_[8299]_  = \new_[13534]_  ? \new_[12030]_  : \new_[9175]_ ;
  assign \new_[8300]_  = \new_[13540]_  ? \new_[12030]_  : \new_[9190]_ ;
  assign \new_[8301]_  = \new_[13748]_  ? \new_[12030]_  : \new_[9178]_ ;
  assign \new_[8302]_  = \new_[13412]_  ? \new_[12030]_  : \new_[9179]_ ;
  assign \new_[8303]_  = \new_[13834]_  ? \new_[12030]_  : \new_[9180]_ ;
  assign \new_[8304]_  = \new_[13490]_  ? \new_[12030]_  : \new_[9181]_ ;
  assign \new_[8305]_  = \new_[13266]_  ? \new_[12030]_  : \new_[9182]_ ;
  assign \new_[8306]_  = \new_[13719]_  ? \new_[12030]_  : \new_[9183]_ ;
  assign \new_[8307]_  = \new_[13778]_  ? \new_[12030]_  : \new_[9184]_ ;
  assign \new_[8308]_  = \new_[13466]_  ? \new_[12028]_  : \new_[9185]_ ;
  assign \new_[8309]_  = \new_[13673]_  ? \new_[12028]_  : \new_[9157]_ ;
  assign \new_[8310]_  = \new_[13625]_  ? \new_[12028]_  : \new_[9186]_ ;
  assign \new_[8311]_  = \new_[13607]_  ? \new_[12028]_  : \new_[9187]_ ;
  assign \new_[8312]_  = \new_[13221]_  ? \new_[12028]_  : \new_[9189]_ ;
  assign \new_[8313]_  = \new_[13458]_  ? \new_[12028]_  : \new_[9188]_ ;
  assign \new_[8314]_  = \new_[13144]_  ^ \new_[9155]_ ;
  assign \new_[8315]_  = ~\new_[8850]_  | ~\new_[13622]_ ;
  assign \new_[8316]_  = ~\new_[8875]_  | ~\new_[13500]_ ;
  assign \new_[8317]_  = ~\new_[8857]_  | ~\new_[13738]_ ;
  assign \new_[8318]_  = ~\new_[14076]_  | ~\new_[13622]_ ;
  assign \new_[8319]_  = ~\new_[8854]_  | ~\new_[13622]_ ;
  assign \new_[8320]_  = ~\new_[13622]_  | ~\new_[8848]_ ;
  assign \new_[8321]_  = ~\new_[8860]_  | ~\new_[12895]_ ;
  assign \new_[8322]_  = ~\new_[8863]_  | ~\new_[12895]_ ;
  assign \new_[8323]_  = ~\new_[8909]_  | ~\new_[13500]_ ;
  assign \new_[8324]_  = ~\new_[8864]_  | ~\new_[12895]_ ;
  assign \new_[8325]_  = ~\new_[8867]_  | ~\new_[12895]_ ;
  assign \new_[8326]_  = ~\new_[8889]_  | ~\new_[13622]_ ;
  assign \new_[8327]_  = ~\new_[8846]_  | ~\new_[13622]_ ;
  assign \new_[8328]_  = ~\new_[8856]_  | ~\new_[13622]_ ;
  assign \new_[8329]_  = ~\new_[8900]_  | ~\new_[14127]_ ;
  assign \new_[8330]_  = ~\new_[8885]_  | ~\new_[13794]_ ;
  assign \new_[8331]_  = ~\new_[8886]_  | ~\new_[13794]_ ;
  assign \new_[8332]_  = ~\new_[8890]_  | ~\new_[13500]_ ;
  assign \new_[8333]_  = ~\new_[8894]_  | ~\new_[14127]_ ;
  assign \new_[8334]_  = ~\new_[8895]_  | ~\new_[14127]_ ;
  assign \new_[8335]_  = ~\new_[8897]_  | ~\new_[14127]_ ;
  assign \new_[8336]_  = ~\new_[8898]_  | ~\new_[14127]_ ;
  assign \new_[8337]_  = ~\new_[8853]_  | ~\new_[14127]_ ;
  assign \new_[8338]_  = ~\new_[14064]_  | ~\new_[14127]_ ;
  assign \new_[8339]_  = ~\new_[8921]_  | ~\new_[13738]_ ;
  assign \new_[8340]_  = ~\new_[8907]_  | ~\new_[13500]_ ;
  assign \new_[8341]_  = ~\new_[14109]_  | ~\new_[13500]_ ;
  assign \new_[8342]_  = ~\new_[14176]_  | ~\new_[13500]_ ;
  assign \new_[8343]_  = ~\new_[13937]_  | ~\new_[13500]_ ;
  assign \new_[8344]_  = ~\new_[8931]_  | ~\new_[13738]_ ;
  assign \new_[8345]_  = ~\new_[8906]_  | ~\new_[13500]_ ;
  assign \new_[8346]_  = ~\new_[8919]_  | ~\new_[13500]_ ;
  assign \new_[8347]_  = ~\new_[8930]_  | ~\new_[13500]_ ;
  assign \new_[8348]_  = ~\new_[13908]_  | ~\new_[13500]_ ;
  assign \new_[8349]_  = ~\new_[8911]_  | ~\new_[13500]_ ;
  assign \new_[8350]_  = ~\new_[13906]_  | ~\new_[13500]_ ;
  assign \new_[8351]_  = ~\new_[8926]_  | ~\new_[13738]_ ;
  assign \new_[8352]_  = ~\new_[8927]_  | ~\new_[13738]_ ;
  assign \new_[8353]_  = ~\new_[8901]_  | ~\new_[14127]_ ;
  assign \new_[8354]_  = ~\new_[8873]_  | ~\new_[12895]_ ;
  assign \new_[8355]_  = ~\new_[8932]_  | ~\new_[13169]_ ;
  assign \new_[8356]_  = ~\new_[8850]_  | ~\new_[14081]_ ;
  assign \new_[8357]_  = ~\new_[8866]_  | ~\new_[12860]_ ;
  assign \new_[8358]_  = ~\new_[8918]_  | ~\new_[13935]_ ;
  assign \new_[8359]_  = ~\new_[8931]_  | ~\new_[12583]_ ;
  assign \new_[8360]_  = ~\new_[8854]_  | ~\new_[14081]_ ;
  assign \new_[8361]_  = ~\new_[8846]_  | ~\new_[14081]_ ;
  assign \new_[8362]_  = ~\new_[8926]_  | ~\new_[12843]_ ;
  assign \new_[8363]_  = ~\new_[8889]_  | ~\new_[14081]_ ;
  assign \new_[8364]_  = ~\new_[8857]_  | ~\new_[12583]_ ;
  assign \new_[8365]_  = ~\new_[8869]_  | ~\new_[12874]_ ;
  assign \new_[8366]_  = ~\new_[8864]_  | ~\new_[12863]_ ;
  assign \new_[8367]_  = ~\new_[8856]_  | ~\new_[14081]_ ;
  assign \new_[8368]_  = ~\new_[8907]_  | ~\new_[13935]_ ;
  assign \new_[8369]_  = ~\new_[8898]_  | ~\new_[12544]_ ;
  assign \new_[8370]_  = ~\new_[14011]_  | ~\new_[12591]_ ;
  assign \new_[8371]_  = ~\new_[8902]_  | ~\new_[12544]_ ;
  assign \new_[8372]_  = ~\new_[8886]_  | ~\new_[12591]_ ;
  assign \new_[8373]_  = ~\new_[8885]_  | ~\new_[12584]_ ;
  assign \new_[8374]_  = ~\new_[14011]_  | ~\new_[13154]_ ;
  assign \new_[8375]_  = ~\new_[8925]_  | ~\new_[12583]_ ;
  assign \new_[8376]_  = ~\new_[13934]_  | ~\new_[13935]_ ;
  assign \new_[8377]_  = ~\new_[8899]_  | ~\new_[13140]_ ;
  assign \new_[8378]_  = ~\new_[8895]_  | ~\new_[12544]_ ;
  assign \new_[8379]_  = ~\new_[14054]_  | ~\new_[12544]_ ;
  assign \new_[8380]_  = ~\new_[8897]_  | ~\new_[12544]_ ;
  assign \new_[8381]_  = ~\new_[8853]_  | ~\new_[12544]_ ;
  assign \new_[8382]_  = ~\new_[8900]_  | ~\new_[12544]_ ;
  assign \new_[8383]_  = ~\new_[8880]_  | ~\new_[12544]_ ;
  assign \new_[8384]_  = ~\new_[8901]_  | ~\new_[12544]_ ;
  assign \new_[8385]_  = ~\new_[8893]_  | ~\new_[12860]_ ;
  assign \new_[8386]_  = ~\new_[8902]_  | ~\new_[12860]_ ;
  assign \new_[8387]_  = ~\new_[14064]_  | ~\new_[12860]_ ;
  assign \new_[8388]_  = ~\new_[13891]_  | ~\new_[12860]_ ;
  assign \new_[8389]_  = ~\new_[8909]_  | ~\new_[13935]_ ;
  assign \new_[8390]_  = ~\new_[14109]_  | ~\new_[13935]_ ;
  assign \new_[8391]_  = ~\new_[14176]_  | ~\new_[13935]_ ;
  assign \new_[8392]_  = ~\new_[8913]_  | ~\new_[13935]_ ;
  assign \new_[8393]_  = ~\new_[8899]_  | ~\new_[13935]_ ;
  assign \new_[8394]_  = ~\new_[8930]_  | ~\new_[13935]_ ;
  assign \new_[8395]_  = ~\new_[8921]_  | ~\new_[12583]_ ;
  assign \new_[8396]_  = ~\new_[8912]_  | ~\new_[14081]_ ;
  assign \new_[8397]_  = ~\new_[13908]_  | ~\new_[13935]_ ;
  assign \new_[8398]_  = ~\new_[8919]_  | ~\new_[14145]_ ;
  assign \new_[8399]_  = ~\new_[8892]_  | ~\new_[13140]_ ;
  assign \new_[8400]_  = ~\new_[8911]_  | ~\new_[13935]_ ;
  assign \new_[8401]_  = ~\new_[8923]_  | ~\new_[12583]_ ;
  assign \new_[8402]_  = ~\new_[8890]_  | ~\new_[13935]_ ;
  assign \new_[8403]_  = ~\new_[8918]_  | ~\new_[13140]_ ;
  assign \new_[8404]_  = ~\new_[8908]_  | ~\new_[13935]_ ;
  assign \new_[8405]_  = ~\new_[8875]_  | ~\new_[13935]_ ;
  assign \new_[8406]_  = ~\new_[8927]_  | ~\new_[12583]_ ;
  assign \new_[8407]_  = ~\new_[8855]_  | ~\new_[13935]_ ;
  assign \new_[8408]_  = ~\new_[8923]_  | ~\new_[13135]_ ;
  assign \new_[8409]_  = ~\new_[8925]_  | ~\new_[13135]_ ;
  assign \new_[8410]_  = ~\new_[8906]_  | ~\new_[14145]_ ;
  assign \new_[8411]_  = ~\new_[8880]_  | ~\new_[12717]_ ;
  assign \new_[8412]_  = ~\new_[14064]_  | ~\new_[12544]_ ;
  assign \new_[8413]_  = ~\new_[8645]_ ;
  assign \new_[8414]_  = ~\new_[8913]_  | ~\new_[13140]_ ;
  assign \new_[8415]_  = ~\new_[8863]_  | ~\new_[12863]_ ;
  assign \new_[8416]_  = ~\new_[8871]_  | ~\new_[3024]_ ;
  assign \new_[8417]_  = ~\new_[13154]_  | (~\new_[9828]_  & ~\new_[9315]_ );
  assign \new_[8418]_  = ~\new_[13154]_  | (~\new_[9874]_  & ~\new_[9312]_ );
  assign \new_[8419]_  = ~\new_[12995]_  | (~\new_[9881]_  & ~\new_[9319]_ );
  assign \new_[8420]_  = ~\new_[13186]_  | (~\new_[9824]_  & ~\new_[8989]_ );
  assign \new_[8421]_  = ~\new_[13186]_  | (~\new_[9882]_  & ~\new_[8981]_ );
  assign \new_[8422]_  = ~\new_[13186]_  | (~\new_[9865]_  & ~\new_[9303]_ );
  assign \new_[8423]_  = ~\new_[12995]_  | (~\new_[9848]_  & ~\new_[9291]_ );
  assign \new_[8424]_  = ~\new_[3023]_  | (~\new_[9292]_  & ~\new_[9863]_ );
  assign \new_[8425]_  = ~\new_[3023]_  | (~\new_[9294]_  & ~\new_[9323]_ );
  assign \new_[8426]_  = ~\new_[13186]_  | (~\new_[9843]_  & ~\new_[9293]_ );
  assign \new_[8427]_  = ~\new_[12995]_  | (~\new_[9844]_  & ~\new_[9295]_ );
  assign \new_[8428]_  = ~\new_[3023]_  | (~\new_[9845]_  & ~\new_[9296]_ );
  assign \new_[8429]_  = ~\new_[3023]_  | (~\new_[9846]_  & ~\new_[9297]_ );
  assign \new_[8430]_  = ~\new_[12995]_  | (~\new_[9856]_  & ~\new_[9302]_ );
  assign \new_[8431]_  = ~\new_[12717]_  | (~\new_[9301]_  & ~\new_[8983]_ );
  assign \new_[8432]_  = ~\new_[8905]_  | ~\new_[3024]_ ;
  assign \new_[8433]_  = ~\new_[12717]_  | (~\new_[9300]_  & ~\new_[8985]_ );
  assign \new_[8434]_  = ~\new_[8874]_  | ~\new_[3024]_ ;
  assign \new_[8435]_  = ~\new_[13154]_  | (~\new_[9306]_  & ~\new_[9868]_ );
  assign \new_[8436]_  = ~\new_[13154]_  | (~\new_[9307]_  & ~\new_[9871]_ );
  assign \new_[8437]_  = ~\new_[13154]_  | (~\new_[9308]_  & ~\new_[9872]_ );
  assign \new_[8438]_  = ~\new_[13154]_  | (~\new_[9309]_  & ~\new_[9849]_ );
  assign \new_[8439]_  = ~\new_[13154]_  | (~\new_[9311]_  & ~\new_[9873]_ );
  assign \new_[8440]_  = ~\new_[13154]_  | (~\new_[9314]_  & ~\new_[9875]_ );
  assign \new_[8441]_  = ~\new_[13154]_  | (~\new_[9877]_  & ~\new_[9316]_ );
  assign \new_[8442]_  = ~\new_[12717]_  | (~\new_[8982]_  & ~\new_[9310]_ );
  assign \new_[8443]_  = ~\new_[13154]_  | (~\new_[9842]_  & ~\new_[9318]_ );
  assign \new_[8444]_  = ~\new_[13154]_  | (~\new_[9299]_  & ~\new_[9866]_ );
  assign \new_[8445]_  = ~\new_[13154]_  | (~\new_[9878]_  & ~\new_[9317]_ );
  assign \new_[8446]_  = ~\new_[12717]_  | (~\new_[8992]_  & ~\new_[8986]_ );
  assign \new_[8447]_  = ~\new_[12717]_  | (~\new_[8988]_  & ~\new_[8987]_ );
  assign \new_[8448]_  = ~\new_[12717]_  | (~\new_[9305]_  & ~\new_[9313]_ );
  assign \new_[8449]_  = ~\new_[8904]_  | ~\new_[12717]_ ;
  assign \new_[8450]_  = ~\new_[12717]_  | (~\new_[8991]_  & ~\new_[8990]_ );
  assign \new_[8451]_  = ~\new_[8915]_  | ~\new_[13135]_ ;
  assign \new_[8452]_  = ~\new_[8870]_  | ~\new_[3024]_ ;
  assign \new_[8453]_  = ~\new_[8851]_  & (~\new_[13670]_  | ~\new_[12513]_ );
  assign \new_[8454]_  = ~\new_[8852]_  & (~\new_[13672]_  | ~\new_[12513]_ );
  assign \new_[8455]_  = ~\new_[8698]_ ;
  assign \new_[8456]_  = ~\new_[8702]_ ;
  assign \new_[8457]_  = ~\new_[14008]_ ;
  assign \new_[8458]_  = ~\new_[8704]_ ;
  assign \new_[8459]_  = ~\new_[8707]_ ;
  assign \new_[8460]_  = ~\new_[8708]_ ;
  assign \new_[8461]_  = ~\new_[8709]_ ;
  assign \new_[8462]_  = ~\new_[8724]_ ;
  assign \new_[8463]_  = ~\new_[13963]_ ;
  assign \new_[8464]_  = ~\new_[8725]_ ;
  assign \new_[8465]_  = ~\new_[8726]_ ;
  assign \new_[8466]_  = ~\new_[8733]_ ;
  assign \new_[8467]_  = ~\new_[8743]_ ;
  assign \new_[8468]_  = ~\new_[8756]_ ;
  assign \new_[8469]_  = ~\new_[8763]_ ;
  assign \new_[8470]_  = (~\new_[12117]_  | ~\new_[9067]_ ) & (~\new_[9030]_  | ~\new_[9784]_ );
  assign n10046 = \new_[8791]_  & \new_[4582]_ ;
  assign n10021 = ~\new_[8789]_  | ~\new_[9101]_ ;
  assign n10041 = ~\new_[8792]_  & ~\new_[9656]_ ;
  assign n10176 = ~\new_[12987]_  & ~\new_[8829]_ ;
  assign n10146 = ~\new_[13068]_  & ~\new_[9661]_ ;
  assign n10151 = ~\new_[13073]_  & ~\new_[9661]_ ;
  assign \new_[8477]_  = u12_we1_reg;
  assign \new_[8478]_  = ~\new_[9003]_  & ~\new_[12468]_ ;
  assign \new_[8479]_  = \new_[13537]_  ^ \new_[9660]_ ;
  assign n10226 = \\u1_sr_reg[4] ;
  assign n10221 = \\u2_in_valid_reg[2] ;
  assign n10231 = ~\new_[8997]_  | ~\new_[9101]_ ;
  assign \new_[8483]_  = \new_[8788]_ ;
  assign \new_[8484]_  = ~\new_[9697]_  & (~\new_[9650]_  | ~\new_[12594]_ );
  assign \new_[8485]_  = ~\new_[10355]_  & (~\new_[9651]_  | ~\new_[12618]_ );
  assign n10196 = ~\new_[8999]_  & ~\new_[9656]_ ;
  assign \new_[8487]_  = \\u10_status_reg[1] ;
  assign \new_[8488]_  = \\u9_status_reg[1] ;
  assign n10216 = \new_[8993]_  & \new_[4582]_ ;
  assign n10236 = ~\new_[11430]_  | ~\new_[9101]_ ;
  assign \new_[8491]_  = ~wb_stb_i | ~\new_[13384]_  | ~\new_[9269]_  | ~wb_cyc_i;
  assign n10201 = n10966 ^ \new_[9654]_ ;
  assign n10206 = n11056 ^ \new_[9655]_ ;
  assign \new_[8494]_  = (~n10936 | ~\new_[7774]_ ) & (~\new_[12119]_  | ~\new_[9645]_ );
  assign \new_[8495]_  = ~u11_empty_reg;
  assign \new_[8496]_  = u2_sync_beat_reg;
  assign \new_[8497]_  = ~\new_[9298]_  | ~\new_[13112]_ ;
  assign \new_[8498]_  = ~\new_[9298]_  | ~\new_[12926]_ ;
  assign \new_[8499]_  = ~\new_[9298]_  | ~\new_[12831]_ ;
  assign n10211 = \new_[9290]_  & \new_[12483]_ ;
  assign \new_[8501]_  = \new_[8788]_ ;
  assign \new_[8502]_  = \new_[13461]_  ^ \new_[14096]_ ;
  assign \new_[8503]_  = u11_full_reg;
  assign \new_[8504]_  = \new_[13759]_  ? \new_[12837]_  : \new_[9701]_ ;
  assign \new_[8505]_  = \new_[9708]_  ? \new_[12828]_  : \new_[13191]_ ;
  assign \new_[8506]_  = \new_[13792]_  ? \new_[12574]_  : \new_[9703]_ ;
  assign \new_[8507]_  = \new_[13347]_  ? \new_[12951]_  : \new_[9704]_ ;
  assign \new_[8508]_  = \new_[13543]_  ? \new_[12951]_  : \new_[9706]_ ;
  assign \new_[8509]_  = \new_[9705]_  ? \new_[12828]_  : \new_[13652]_ ;
  assign n10246 = ~\new_[9099]_  & ~\new_[9656]_ ;
  assign \new_[8511]_  = \new_[9707]_  ? \new_[12828]_  : \new_[13236]_ ;
  assign \new_[8512]_  = \new_[13263]_  ? \new_[12574]_  : \new_[9709]_ ;
  assign \new_[8513]_  = \new_[13241]_  ? \new_[12574]_  : \new_[9701]_ ;
  assign \new_[8514]_  = \new_[9703]_  ? \new_[12432]_  : \new_[13380]_ ;
  assign \new_[8515]_  = \new_[9704]_  ? \new_[12432]_  : \new_[13691]_ ;
  assign \new_[8516]_  = \new_[9706]_  ? \new_[12432]_  : \new_[13394]_ ;
  assign \new_[8517]_  = \new_[9702]_  ? \new_[12432]_  : \new_[13233]_ ;
  assign \new_[8518]_  = \new_[9709]_  ? \new_[12432]_  : \new_[13411]_ ;
  assign \new_[8519]_  = \new_[9701]_  ? \new_[12432]_  : \new_[13856]_ ;
  assign \new_[8520]_  = \new_[13603]_  ? \new_[12574]_  : \new_[9702]_ ;
  assign \new_[8521]_  = \new_[13627]_  ? \new_[12642]_  : \new_[9707]_ ;
  assign \new_[8522]_  = \new_[13727]_  ? \new_[12626]_  : \new_[9707]_ ;
  assign \new_[8523]_  = \new_[13741]_  ? \new_[12626]_  : \new_[9705]_ ;
  assign \new_[8524]_  = \new_[13645]_  ? \new_[12626]_  : \new_[9708]_ ;
  assign \new_[8525]_  = \new_[13654]_  ? \new_[12663]_  : \new_[9702]_ ;
  assign \new_[8526]_  = \new_[13680]_  ? \new_[12642]_  : \new_[9705]_ ;
  assign n10241 = ~\new_[9100]_  & ~\new_[9656]_ ;
  assign \new_[8528]_  = \new_[13470]_  ? \new_[12663]_  : \new_[9703]_ ;
  assign \new_[8529]_  = \new_[13687]_  ? \new_[12663]_  : \new_[9704]_ ;
  assign \new_[8530]_  = \new_[13473]_  ? \new_[12663]_  : \new_[9706]_ ;
  assign \new_[8531]_  = \new_[13660]_  ? \new_[12642]_  : \new_[9708]_ ;
  assign \new_[8532]_  = \new_[13276]_  ? \new_[12663]_  : \new_[9709]_ ;
  assign \new_[8533]_  = \new_[13482]_  ^ \new_[9663]_ ;
  assign \new_[8534]_  = \new_[13793]_  ? \new_[12028]_  : \new_[9701]_ ;
  assign \new_[8535]_  = \new_[13864]_  ? \new_[12028]_  : \new_[9702]_ ;
  assign \new_[8536]_  = \new_[13831]_  ? \new_[12028]_  : \new_[9703]_ ;
  assign \new_[8537]_  = \new_[13565]_  ? \new_[12028]_  : \new_[9704]_ ;
  assign \new_[8538]_  = \new_[13464]_  ? \new_[12030]_  : \new_[9707]_ ;
  assign \new_[8539]_  = \new_[13567]_  ? \new_[12030]_  : \new_[9705]_ ;
  assign \new_[8540]_  = \new_[13817]_  ? \new_[12028]_  : \new_[9706]_ ;
  assign \new_[8541]_  = \new_[13731]_  ? \new_[12030]_  : \new_[9708]_ ;
  assign \new_[8542]_  = \new_[13795]_  ? \new_[12028]_  : \new_[9709]_ ;
  assign \new_[8543]_  = \new_[13175]_  ^ \new_[9700]_ ;
  assign \new_[8544]_  = \\u10_dout_reg[14] ;
  assign \new_[8545]_  = \\u10_dout_reg[15] ;
  assign \new_[8546]_  = \\u10_dout_reg[17] ;
  assign \new_[8547]_  = \\u10_dout_reg[18] ;
  assign \new_[8548]_  = \\u10_dout_reg[19] ;
  assign \new_[8549]_  = \\u10_dout_reg[1] ;
  assign \new_[8550]_  = \\u10_dout_reg[20] ;
  assign \new_[8551]_  = \\u10_dout_reg[21] ;
  assign \new_[8552]_  = \\u10_dout_reg[22] ;
  assign \new_[8553]_  = \\u10_dout_reg[23] ;
  assign \new_[8554]_  = ~\new_[13794]_  | ~\new_[14116]_ ;
  assign \new_[8555]_  = ~\new_[9152]_  | ~\new_[13738]_ ;
  assign \new_[8556]_  = ~\new_[9151]_  | ~\new_[13738]_ ;
  assign \new_[8557]_  = ~\new_[9115]_  | ~\new_[12895]_ ;
  assign \new_[8558]_  = ~\new_[9116]_  | ~\new_[12895]_ ;
  assign \new_[8559]_  = ~\new_[9117]_  | ~\new_[12895]_ ;
  assign \new_[8560]_  = ~\new_[9118]_  | ~\new_[12895]_ ;
  assign \new_[8561]_  = ~\new_[9119]_  | ~\new_[12895]_ ;
  assign \new_[8562]_  = ~\new_[9120]_  | ~\new_[12895]_ ;
  assign \new_[8563]_  = ~\new_[9122]_  | ~\new_[12895]_ ;
  assign \new_[8564]_  = ~\new_[9124]_  | ~\new_[13425]_ ;
  assign \new_[8565]_  = ~\new_[9129]_  | ~\new_[13794]_ ;
  assign \new_[8566]_  = ~\new_[9131]_  | ~\new_[13794]_ ;
  assign \new_[8567]_  = ~\new_[9130]_  | ~\new_[13794]_ ;
  assign \new_[8568]_  = ~\new_[9132]_  | ~\new_[13794]_ ;
  assign \new_[8569]_  = ~\new_[13794]_  | ~\new_[9134]_ ;
  assign \new_[8570]_  = ~\new_[9135]_  | ~\new_[13794]_ ;
  assign \new_[8571]_  = ~\new_[13794]_  | ~\new_[9128]_ ;
  assign \new_[8572]_  = ~\new_[9141]_  | ~\new_[14127]_ ;
  assign \new_[8573]_  = ~\new_[9137]_  | ~\new_[13794]_ ;
  assign \new_[8574]_  = ~\new_[9138]_  | ~\new_[13794]_ ;
  assign \new_[8575]_  = ~\new_[9149]_  | ~\new_[13738]_ ;
  assign \new_[8576]_  = ~\new_[9142]_  | ~\new_[14127]_ ;
  assign \new_[8577]_  = ~\new_[9113]_  | ~\new_[13738]_ ;
  assign \new_[8578]_  = ~\new_[9102]_  | ~\new_[13738]_ ;
  assign \new_[8579]_  = ~\new_[9147]_  | ~\new_[13738]_ ;
  assign \new_[8580]_  = ~\new_[9148]_  | ~\new_[13738]_ ;
  assign \new_[8581]_  = ~\new_[9150]_  | ~\new_[13738]_ ;
  assign \new_[8582]_  = ~\new_[9143]_  | ~\new_[13738]_ ;
  assign \new_[8583]_  = ~\new_[9145]_  | ~\new_[13738]_ ;
  assign \new_[8584]_  = ~\new_[9146]_  | ~\new_[13738]_ ;
  assign \new_[8585]_  = ~\new_[9103]_  | ~\new_[13425]_ ;
  assign \new_[8586]_  = ~\new_[9153]_  | ~\new_[4763]_ ;
  assign \new_[8587]_  = ~\new_[9156]_  | ~\new_[13105]_ ;
  assign \new_[8588]_  = ~\new_[9154]_  | ~\new_[13127]_ ;
  assign \new_[8589]_  = ~\new_[9146]_  | ~\new_[12583]_ ;
  assign \new_[8590]_  = ~\new_[9133]_  | ~\new_[13135]_ ;
  assign \new_[8591]_  = ~\new_[9113]_  | ~\new_[12583]_ ;
  assign \new_[8592]_  = ~\new_[9152]_  | ~\new_[12583]_ ;
  assign \new_[8593]_  = ~\new_[13084]_  & ~\new_[9101]_ ;
  assign \new_[8594]_  = ~\new_[9139]_  | ~\new_[13135]_ ;
  assign n10256 = ~\new_[9670]_  | ~\new_[9101]_ ;
  assign \new_[8596]_  = ~\new_[9121]_  | ~\new_[3024]_ ;
  assign \new_[8597]_  = ~\new_[9116]_  | ~\new_[12863]_ ;
  assign \new_[8598]_  = ~\new_[9117]_  | ~\new_[12863]_ ;
  assign \new_[8599]_  = ~\new_[9118]_  | ~\new_[12874]_ ;
  assign \new_[8600]_  = ~\new_[9119]_  | ~\new_[12874]_ ;
  assign \new_[8601]_  = ~\new_[9118]_  | ~\new_[13035]_ ;
  assign \new_[8602]_  = ~\new_[9119]_  | ~\new_[13035]_ ;
  assign \new_[8603]_  = ~\new_[9121]_  | ~\new_[12863]_ ;
  assign \new_[8604]_  = ~\new_[14147]_  | ~\new_[12863]_ ;
  assign \new_[8605]_  = ~\new_[9121]_  | ~\new_[13035]_ ;
  assign \new_[8606]_  = ~\new_[9123]_  | ~\new_[12501]_ ;
  assign \new_[8607]_  = ~\new_[9114]_  | ~\new_[13035]_ ;
  assign \new_[8608]_  = ~\new_[9124]_  | ~\new_[12501]_ ;
  assign \new_[8609]_  = ~\new_[9122]_  | ~\new_[13035]_ ;
  assign \new_[8610]_  = ~\new_[9123]_  | ~\new_[13035]_ ;
  assign \new_[8611]_  = ~\new_[9124]_  | ~\new_[13035]_ ;
  assign \new_[8612]_  = ~\new_[9103]_  | ~\new_[13035]_ ;
  assign \new_[8613]_  = ~\new_[9115]_  | ~\new_[12874]_ ;
  assign \new_[8614]_  = ~\new_[12591]_  | ~\new_[9130]_ ;
  assign \new_[8615]_  = ~\new_[12591]_  | ~\new_[9132]_ ;
  assign \new_[8616]_  = ~\new_[12591]_  | ~\new_[9134]_ ;
  assign \new_[8617]_  = ~\new_[14116]_  | ~\new_[12591]_ ;
  assign \new_[8618]_  = ~\new_[12591]_  | ~\new_[9135]_ ;
  assign \new_[8619]_  = ~\new_[9136]_  | ~\new_[12591]_ ;
  assign \new_[8620]_  = ~\new_[9128]_  | ~\new_[12584]_ ;
  assign \new_[8621]_  = ~\new_[12591]_  | ~\new_[9137]_ ;
  assign \new_[8622]_  = ~\new_[10319]_  & ~\new_[12811]_ ;
  assign \new_[8623]_  = ~\new_[12591]_  | ~\new_[9138]_ ;
  assign \new_[8624]_  = ~\new_[12591]_  | ~\new_[9129]_ ;
  assign \new_[8625]_  = ~\new_[12591]_  | ~\new_[9131]_ ;
  assign \new_[8626]_  = ~\new_[10320]_  & ~\new_[12718]_ ;
  assign \new_[8627]_  = ~\new_[9136]_  | ~\new_[13154]_ ;
  assign \new_[8628]_  = ~\new_[10318]_  & ~\new_[12853]_ ;
  assign \new_[8629]_  = ~\new_[10321]_  & ~\new_[13168]_ ;
  assign \new_[8630]_  = ~\new_[9139]_  | ~\new_[12583]_ ;
  assign n10261 = ~\new_[7978]_  | ~\new_[9101]_ ;
  assign n10191 = ~\new_[12002]_  | ~\new_[9101]_ ;
  assign n10266 = ~\new_[12265]_  | ~\new_[9101]_ ;
  assign \new_[8634]_  = ~\new_[9140]_  | ~\new_[12544]_ ;
  assign \new_[8635]_  = ~\new_[9140]_  | ~\new_[12860]_ ;
  assign \new_[8636]_  = ~\new_[9149]_  | ~\new_[12583]_ ;
  assign \new_[8637]_  = ~\new_[9147]_  | ~\new_[12583]_ ;
  assign \new_[8638]_  = ~\new_[9148]_  | ~\new_[12583]_ ;
  assign \new_[8639]_  = ~\new_[9143]_  | ~\new_[12583]_ ;
  assign \new_[8640]_  = ~\new_[9150]_  | ~\new_[12583]_ ;
  assign \new_[8641]_  = ~\new_[9133]_  | ~\new_[12583]_ ;
  assign \new_[8642]_  = ~\new_[9145]_  | ~\new_[12843]_ ;
  assign \new_[8643]_  = ~\new_[9151]_  | ~\new_[12583]_ ;
  assign \new_[8644]_  = ~\new_[9102]_  | ~\new_[12583]_ ;
  assign \new_[8645]_  = \new_[9125]_  & \new_[12455]_ ;
  assign \new_[8646]_  = ~\new_[13140]_  | (~\new_[9330]_  & ~\new_[9331]_ );
  assign \new_[8647]_  = ~\new_[9266]_  | ~\new_[10405]_ ;
  assign \new_[8648]_  = ~\new_[13135]_  | (~\new_[9841]_  & ~\new_[9352]_ );
  assign \new_[8649]_  = ~\new_[13135]_  | (~\new_[9350]_  & ~\new_[9351]_ );
  assign \new_[8650]_  = ~\new_[9249]_  | ~\new_[10403]_ ;
  assign \new_[8651]_  = ~\new_[13135]_  | (~\new_[9892]_  & ~\new_[9342]_ );
  assign \new_[8652]_  = ~\new_[9251]_  & (~\new_[11697]_  | ~\new_[5065]_ );
  assign \new_[8653]_  = ~\new_[9254]_  | ~\new_[10408]_ ;
  assign \new_[8654]_  = ~\new_[9248]_  | ~\new_[10404]_ ;
  assign \new_[8655]_  = ~\new_[9256]_  | ~\new_[10409]_ ;
  assign \new_[8656]_  = ~\new_[9257]_  | ~\new_[11462]_ ;
  assign \new_[8657]_  = ~\new_[9258]_  | ~\new_[10411]_ ;
  assign \new_[8658]_  = ~\new_[9259]_  | ~\new_[11463]_ ;
  assign \new_[8659]_  = ~\new_[9260]_  | ~\new_[11464]_ ;
  assign \new_[8660]_  = ~\new_[9261]_  | ~\new_[10412]_ ;
  assign \new_[8661]_  = ~\new_[9262]_  | ~\new_[10413]_ ;
  assign \new_[8662]_  = ~\new_[9267]_  | ~\new_[11438]_ ;
  assign \new_[8663]_  = ~\new_[3024]_  | (~\new_[10455]_  & ~\new_[9852]_ );
  assign \new_[8664]_  = ~\new_[3024]_  | (~\new_[10456]_  & ~\new_[9853]_ );
  assign \new_[8665]_  = ~\new_[13075]_  | (~\new_[9880]_  & ~\new_[9854]_ );
  assign \new_[8666]_  = ~\new_[13075]_  | (~\new_[10457]_  & ~\new_[9855]_ );
  assign \new_[8667]_  = ~\new_[13075]_  | (~\new_[10458]_  & ~\new_[9857]_ );
  assign \new_[8668]_  = ~\new_[13075]_  | (~\new_[9858]_  & ~\new_[9859]_ );
  assign \new_[8669]_  = ~\new_[13075]_  | (~\new_[9869]_  & ~\new_[9860]_ );
  assign \new_[8670]_  = ~\new_[13075]_  | (~\new_[9861]_  & ~\new_[9862]_ );
  assign \new_[8671]_  = ~\new_[13140]_  | (~\new_[9348]_  & ~\new_[9349]_ );
  assign \new_[8672]_  = ~\new_[9264]_  | ~\new_[10406]_ ;
  assign \new_[8673]_  = ~\new_[13075]_  | (~\new_[9864]_  & ~\new_[9332]_ );
  assign \new_[8674]_  = ~\new_[9265]_  | ~\new_[11465]_ ;
  assign \new_[8675]_  = ~\new_[13140]_  | (~\new_[9327]_  & ~\new_[9353]_ );
  assign \new_[8676]_  = ~\new_[9263]_  | ~\new_[10416]_ ;
  assign \new_[8677]_  = ~\new_[13140]_  | (~\new_[9345]_  & ~\new_[9347]_ );
  assign \new_[8678]_  = ~\new_[13135]_  | (~\new_[9344]_  & ~\new_[9870]_ );
  assign \new_[8679]_  = ~\new_[13135]_  | (~\new_[9876]_  & ~\new_[9343]_ );
  assign \new_[8680]_  = ~\new_[13140]_  | (~\new_[9321]_  & ~\new_[9322]_ );
  assign \new_[8681]_  = ~\new_[13140]_  | (~\new_[9830]_  & ~\new_[9324]_ );
  assign \new_[8682]_  = ~\new_[13140]_  | (~\new_[9336]_  & ~\new_[9320]_ );
  assign \new_[8683]_  = ~\new_[13140]_  | (~\new_[9325]_  & ~\new_[9326]_ );
  assign \new_[8684]_  = ~\new_[13140]_  | (~\new_[9334]_  & ~\new_[9335]_ );
  assign \new_[8685]_  = ~\new_[13135]_  | (~\new_[9829]_  & ~\new_[9337]_ );
  assign \new_[8686]_  = ~\new_[13135]_  | (~\new_[9338]_  & ~\new_[9339]_ );
  assign \new_[8687]_  = ~\new_[13135]_  | (~\new_[9341]_  & ~\new_[9333]_ );
  assign \new_[8688]_  = ~\new_[13135]_  | (~\new_[9893]_  & ~\new_[9340]_ );
  assign \new_[8689]_  = ~\new_[13135]_  | (~\new_[9894]_  & ~\new_[9354]_ );
  assign \new_[8690]_  = ~\new_[13135]_  | (~\new_[9879]_  & ~\new_[9346]_ );
  assign n10251 = ~\new_[9669]_  | ~\new_[9101]_ ;
  assign \new_[8692]_  = \new_[3192]_  ? \new_[12027]_  : \new_[9827]_ ;
  assign \new_[8693]_  = \new_[3193]_  ? \new_[12027]_  : \new_[9833]_ ;
  assign \new_[8694]_  = \new_[3198]_  ? \new_[12733]_  : \new_[9827]_ ;
  assign \new_[8695]_  = \new_[3212]_  ? \new_[12760]_  : \new_[9827]_ ;
  assign \new_[8696]_  = \new_[3213]_  ? \new_[12760]_  : \new_[9833]_ ;
  assign \new_[8697]_  = \new_[3199]_  ? \new_[12733]_  : \new_[9833]_ ;
  assign \new_[8698]_  = ~\new_[11577]_  | ~\new_[10173]_  | ~\new_[10757]_  | ~\new_[11088]_ ;
  assign \new_[8699]_  = ~\new_[8846]_ ;
  assign \new_[8700]_  = ~\new_[8848]_ ;
  assign \new_[8701]_  = ~\new_[8850]_ ;
  assign \new_[8702]_  = ~\new_[10190]_  | ~\new_[11221]_  | ~\new_[11018]_  | ~\new_[10162]_ ;
  assign \new_[8703]_  = ~\new_[8853]_ ;
  assign \new_[8704]_  = ~\new_[10163]_  | ~\new_[11639]_  | ~\new_[10177]_  | ~\new_[10751]_ ;
  assign \new_[8705]_  = ~\new_[10170]_  | ~\new_[11720]_  | ~\new_[10254]_  | ~\new_[11161]_ ;
  assign \new_[8706]_  = ~\new_[10164]_  | ~\new_[11640]_  | ~\new_[10252]_  | ~\new_[10836]_ ;
  assign \new_[8707]_  = ~\new_[10165]_  | ~\new_[11704]_  | ~\new_[10217]_  | ~\new_[11045]_ ;
  assign \new_[8708]_  = ~\new_[10166]_  | ~\new_[11668]_  | ~\new_[10219]_  | ~\new_[12315]_ ;
  assign \new_[8709]_  = ~\new_[10167]_  | ~\new_[11677]_  | ~\new_[10204]_  | ~\new_[10841]_ ;
  assign \new_[8710]_  = ~\new_[14076]_ ;
  assign \new_[8711]_  = ~\new_[8854]_ ;
  assign \new_[8712]_  = ~\new_[8855]_ ;
  assign \new_[8713]_  = ~\new_[8856]_ ;
  assign \new_[8714]_  = ~\new_[8857]_ ;
  assign \new_[8715]_  = ~\new_[8860]_ ;
  assign \new_[8716]_  = ~\new_[8863]_ ;
  assign \new_[8717]_  = ~\new_[8864]_ ;
  assign \new_[8718]_  = ~\new_[8866]_ ;
  assign \new_[8719]_  = ~\new_[8867]_ ;
  assign \new_[8720]_  = ~\new_[8869]_ ;
  assign \new_[8721]_  = ~\new_[8871]_ ;
  assign \new_[8722]_  = ~\new_[8873]_ ;
  assign \new_[8723]_  = ~\new_[8875]_ ;
  assign \new_[8724]_  = ~\new_[10172]_  | ~\new_[12113]_  | ~\new_[11071]_  | ~\new_[10279]_ ;
  assign \new_[8725]_  = ~\new_[12050]_  | ~\new_[10175]_  | ~\new_[11059]_  | ~\new_[11204]_ ;
  assign \new_[8726]_  = ~\new_[11553]_  | ~\new_[10238]_  | ~\new_[11065]_  | ~\new_[10926]_ ;
  assign \new_[8727]_  = ~\new_[14011]_ ;
  assign \new_[8728]_  = ~\new_[11579]_  | ~\new_[10244]_  | ~\new_[11094]_  | ~\new_[10779]_ ;
  assign \new_[8729]_  = ~\new_[8885]_ ;
  assign \new_[8730]_  = ~\new_[8886]_ ;
  assign \new_[8731]_  = ~\new_[8889]_ ;
  assign \new_[8732]_  = ~\new_[8890]_ ;
  assign \new_[8733]_  = ~\new_[10215]_  | ~\new_[12095]_  | ~\new_[11153]_  | ~\new_[10168]_ ;
  assign \new_[8734]_  = ~\new_[10795]_  | ~\new_[10198]_  | ~\new_[12406]_  | ~\new_[11135]_ ;
  assign \new_[8735]_  = ~\new_[8892]_ ;
  assign \new_[8736]_  = ~\new_[8893]_ ;
  assign \new_[8737]_  = ~\new_[13891]_ ;
  assign \new_[8738]_  = ~\new_[8894]_ ;
  assign \new_[8739]_  = ~\new_[8895]_ ;
  assign \new_[8740]_  = ~\new_[8897]_ ;
  assign \new_[8741]_  = ~\new_[8898]_ ;
  assign \new_[8742]_  = ~\new_[8900]_ ;
  assign \new_[8743]_  = ~\new_[12385]_  | ~\new_[10216]_  | ~\new_[10174]_  | ~\new_[11780]_ ;
  assign \new_[8744]_  = ~\new_[8901]_ ;
  assign \new_[8745]_  = ~\new_[8906]_ ;
  assign \new_[8746]_  = ~\new_[8907]_ ;
  assign \new_[8747]_  = ~\new_[8908]_ ;
  assign \new_[8748]_  = ~\new_[8909]_ ;
  assign \new_[8749]_  = ~\new_[14109]_ ;
  assign \new_[8750]_  = ~\new_[13937]_ ;
  assign \new_[8751]_  = ~\new_[8911]_ ;
  assign \new_[8752]_  = ~\new_[8912]_ ;
  assign \new_[8753]_  = ~\new_[8913]_ ;
  assign \new_[8754]_  = ~\new_[8919]_ ;
  assign \new_[8755]_  = ~\new_[8921]_ ;
  assign \new_[8756]_  = ~\new_[12390]_  | ~\new_[10273]_  | ~\new_[10191]_  | ~\new_[11652]_ ;
  assign \new_[8757]_  = ~\new_[13906]_ ;
  assign \new_[8758]_  = ~\new_[8923]_ ;
  assign \new_[8759]_  = ~\new_[14054]_ ;
  assign \new_[8760]_  = ~\new_[8926]_ ;
  assign \new_[8761]_  = ~\new_[8927]_ ;
  assign \new_[8762]_  = ~\new_[8930]_ ;
  assign \new_[8763]_  = ~\new_[11581]_  | ~\new_[11726]_  | ~\new_[10228]_  | ~\new_[11017]_ ;
  assign \new_[8764]_  = ~\new_[8931]_ ;
  assign \new_[8765]_  = ~\new_[9277]_  | (~\new_[3317]_  & ~\new_[12030]_ );
  assign \new_[8766]_  = ~\new_[9276]_  | (~\new_[3620]_  & ~\new_[12028]_ );
  assign \new_[8767]_  = ~\new_[9274]_  | (~\new_[3314]_  & ~\new_[12030]_ );
  assign \new_[8768]_  = ~\new_[9281]_  | (~\new_[3322]_  & ~\new_[12028]_ );
  assign \new_[8769]_  = ~\new_[9280]_  | (~\new_[3321]_  & ~\new_[12030]_ );
  assign \new_[8770]_  = ~\new_[9272]_  | (~\new_[3327]_  & ~\new_[12030]_ );
  assign \new_[8771]_  = ~\new_[9283]_  | (~\new_[3324]_  & ~\new_[12647]_ );
  assign \new_[8772]_  = ~\new_[9271]_  | (~\new_[3313]_  & ~\new_[12647]_ );
  assign \new_[8773]_  = ~\new_[9270]_  | (~\new_[3315]_  & ~\new_[12030]_ );
  assign \new_[8774]_  = ~\new_[9275]_  | (~\new_[3316]_  & ~\new_[12030]_ );
  assign \new_[8775]_  = ~\new_[9278]_  | (~\new_[3318]_  & ~\new_[12030]_ );
  assign \new_[8776]_  = ~\new_[9279]_  | (~\new_[3320]_  & ~\new_[12030]_ );
  assign \new_[8777]_  = ~\new_[9284]_  | (~\new_[3448]_  & ~\new_[12028]_ );
  assign \new_[8778]_  = ~\new_[9273]_  | (~\new_[3326]_  & ~\new_[12030]_ );
  assign \new_[8779]_  = ~\new_[9285]_  | (~\new_[3544]_  & ~\new_[12653]_ );
  assign \new_[8780]_  = ~\new_[9286]_  | (~\new_[3329]_  & ~\new_[12653]_ );
  assign \new_[8781]_  = ~\new_[9282]_  | (~\new_[3323]_  & ~\new_[12030]_ );
  assign \new_[8782]_  = ~\new_[9289]_  | (~\new_[3583]_  & ~\new_[12028]_ );
  assign \new_[8783]_  = ~\new_[9288]_  | (~\new_[3581]_  & ~\new_[12028]_ );
  assign \new_[8784]_  = ~\new_[9287]_  | (~\new_[3337]_  & ~\new_[12028]_ );
  assign n10306 = \new_[12347]_  ^ \new_[10316]_ ;
  assign \new_[8786]_  = \new_[13791]_  ^ \new_[10308]_ ;
  assign \new_[8787]_  = ~u12_i4_re_reg;
  assign \new_[8788]_  = ~u2_ld_reg;
  assign \new_[8789]_  = \new_[7807]_  ^ \new_[10290]_ ;
  assign \new_[8790]_  = ~\new_[11447]_  & (~\new_[10291]_  | ~\new_[12679]_ );
  assign \new_[8791]_  = \new_[10292]_  ? \new_[12077]_  : \new_[7865]_ ;
  assign \new_[8792]_  = (~n10936 | ~\new_[7857]_ ) & (~\new_[12119]_  | ~\new_[10293]_ );
  assign n10271 = \new_[9649]_  & \new_[4582]_ ;
  assign n10281 = \new_[9652]_  & \new_[4582]_ ;
  assign \new_[8795]_  = \new_[4756]_  ? \new_[10315]_  : \new_[12880]_ ;
  assign \new_[8796]_  = \new_[4728]_  ? \new_[10315]_  : \new_[12082]_ ;
  assign n10301 = n11061 ^ \new_[10298]_ ;
  assign n10286 = n10961 ^ \new_[10299]_ ;
  assign n10291 = n10956 ^ \new_[10300]_ ;
  assign n10296 = n10971 ^ \new_[10301]_ ;
  assign \new_[8801]_  = \new_[4755]_  ^ \new_[10315]_ ;
  assign \new_[8802]_  = (~n10936 | ~\new_[7874]_ ) & (~\new_[12119]_  | ~\new_[10302]_ );
  assign \new_[8803]_  = u9_full_reg;
  assign \new_[8804]_  = ~u12_i6_re_reg;
  assign \new_[8805]_  = ~\\u2_out_le_reg[1] ;
  assign \new_[8806]_  = ~u12_i3_re_reg;
  assign n10316 = ~\new_[9666]_  & ~\new_[11434]_ ;
  assign n10311 = ~\new_[9662]_  & ~\new_[11435]_ ;
  assign n10321 = \\u2_in_valid_reg[1] ;
  assign \new_[8810]_  = \\u10_dout_reg[11] ;
  assign \new_[8811]_  = \\u10_dout_reg[0] ;
  assign \new_[8812]_  = \\u10_dout_reg[10] ;
  assign \new_[8813]_  = \\u10_dout_reg[12] ;
  assign \new_[8814]_  = \\u10_dout_reg[13] ;
  assign \new_[8815]_  = \\u10_dout_reg[25] ;
  assign \new_[8816]_  = \\u10_dout_reg[27] ;
  assign \new_[8817]_  = \\u10_dout_reg[28] ;
  assign \new_[8818]_  = \\u10_dout_reg[29] ;
  assign \new_[8819]_  = \\u10_dout_reg[2] ;
  assign \new_[8820]_  = \\u10_dout_reg[30] ;
  assign \new_[8821]_  = \\u10_dout_reg[3] ;
  assign \new_[8822]_  = \\u10_dout_reg[4] ;
  assign \new_[8823]_  = \\u10_dout_reg[6] ;
  assign \new_[8824]_  = \\u10_dout_reg[7] ;
  assign \new_[8825]_  = \\u10_dout_reg[8] ;
  assign \new_[8826]_  = \\u10_dout_reg[9] ;
  assign \new_[8827]_  = ~\new_[10437]_  | ~\new_[9644]_ ;
  assign n10276 = ~\new_[12507]_  & (~\new_[10417]_  | ~\new_[12907]_ );
  assign \new_[8829]_  = ~\new_[9077]_ ;
  assign \new_[8830]_  = ~\new_[13027]_  & ~\new_[9677]_ ;
  assign \new_[8831]_  = ~\new_[13038]_  & ~\new_[9673]_ ;
  assign \new_[8832]_  = ~\new_[9677]_  & ~\new_[13867]_ ;
  assign \new_[8833]_  = ~\new_[9673]_  & ~\new_[13874]_ ;
  assign n10326 = ~\new_[9085]_ ;
  assign \new_[8835]_  = ~\new_[9779]_  & (~\new_[11697]_  | ~\new_[5062]_ );
  assign \new_[8836]_  = \new_[10414]_  & \new_[9767]_ ;
  assign \new_[8837]_  = ~\new_[9755]_  & (~\new_[11697]_  | ~\new_[5066]_ );
  assign \new_[8838]_  = ~\new_[9757]_  & (~\new_[11697]_  | ~\new_[5039]_ );
  assign \new_[8839]_  = ~\new_[9760]_  & (~\new_[11697]_  | ~\new_[5067]_ );
  assign \new_[8840]_  = \new_[10410]_  & \new_[9750]_ ;
  assign \new_[8841]_  = \new_[10415]_  & \new_[9778]_ ;
  assign \new_[8842]_  = ~\new_[9699]_  & (~\new_[13694]_  | ~\new_[12828]_ );
  assign \new_[8843]_  = ~\new_[9698]_  & (~\new_[13593]_  | ~\new_[12828]_ );
  assign \new_[8844]_  = ~\new_[9682]_  & (~\new_[13371]_  | ~\new_[12432]_ );
  assign \new_[8845]_  = ~\new_[9683]_  & (~\new_[13311]_  | ~\new_[12432]_ );
  assign \new_[8846]_  = ~\new_[10735]_  | ~\new_[11275]_  | ~\new_[11145]_  | ~\new_[10259]_ ;
  assign \new_[8847]_  = ~\new_[9102]_ ;
  assign \new_[8848]_  = ~\new_[10736]_  | ~\new_[11415]_  | ~\new_[11255]_  | ~\new_[10249]_ ;
  assign \new_[8849]_  = ~\new_[9103]_ ;
  assign \new_[8850]_  = ~\new_[10725]_  | ~\new_[10937]_  | ~\new_[11188]_  | ~\new_[10223]_ ;
  assign \new_[8851]_  = ~\new_[9827]_  & ~\new_[12513]_ ;
  assign \new_[8852]_  = ~\new_[9833]_  & ~\new_[12513]_ ;
  assign \new_[8853]_  = ~\new_[12287]_  | ~\new_[11042]_  | ~\new_[10281]_  | ~\new_[11522]_ ;
  assign \new_[8854]_  = ~\new_[11425]_  | ~\new_[10845]_  | ~\new_[11005]_  | ~\new_[10199]_ ;
  assign \new_[8855]_  = ~\new_[11554]_  | ~\new_[10878]_  | ~\new_[10774]_  | ~\new_[10884]_ ;
  assign \new_[8856]_  = ~\new_[10737]_  | ~\new_[10996]_  | ~\new_[10849]_  | ~\new_[10257]_ ;
  assign \new_[8857]_  = ~\new_[11552]_  | ~\new_[11259]_  | ~\new_[10879]_  | ~\new_[11196]_ ;
  assign \new_[8858]_  = ~\new_[9113]_ ;
  assign \new_[8859]_  = ~\new_[9114]_ ;
  assign \new_[8860]_  = ~\new_[12419]_  | ~\new_[10924]_  | ~\new_[10923]_  | ~\new_[11729]_ ;
  assign \new_[8861]_  = ~\new_[9115]_ ;
  assign \new_[8862]_  = ~\new_[9116]_ ;
  assign \new_[8863]_  = ~\new_[12268]_  | ~\new_[10932]_  | ~\new_[11660]_  | ~\new_[10931]_ ;
  assign \new_[8864]_  = ~\new_[12420]_  | ~\new_[10974]_  | ~\new_[11648]_  | ~\new_[10933]_ ;
  assign \new_[8865]_  = ~\new_[9117]_ ;
  assign \new_[8866]_  = ~\new_[12398]_  | ~\new_[11112]_  | ~\new_[10276]_  | ~\new_[11661]_ ;
  assign \new_[8867]_  = ~\new_[12273]_  | ~\new_[10949]_  | ~\new_[10948]_  | ~\new_[11630]_ ;
  assign \new_[8868]_  = ~\new_[9120]_ ;
  assign \new_[8869]_  = ~\new_[11589]_  | ~\new_[11708]_  | ~\new_[10959]_  | ~\new_[10958]_ ;
  assign \new_[8870]_  = ~\new_[11754]_  | ~\new_[11267]_  | ~\new_[10728]_  | ~\new_[10963]_ ;
  assign \new_[8871]_  = ~\new_[11563]_  | ~\new_[10967]_  | ~\new_[11740]_  | ~\new_[10966]_ ;
  assign \new_[8872]_  = ~\new_[9122]_ ;
  assign \new_[8873]_  = ~\new_[12413]_  | ~\new_[11477]_  | ~\new_[10978]_  | ~\new_[11644]_ ;
  assign \new_[8874]_  = ~\new_[12110]_  | ~\new_[10907]_  | ~\new_[10743]_  | ~\new_[10981]_ ;
  assign \new_[8875]_  = ~\new_[11593]_  | ~\new_[11016]_  | ~\new_[11202]_  | ~\new_[11205]_ ;
  assign \new_[8876]_  = ~\new_[9128]_ ;
  assign \new_[8877]_  = ~\new_[9129]_ ;
  assign \new_[8878]_  = ~\new_[9130]_ ;
  assign \new_[8879]_  = ~\new_[9131]_ ;
  assign \new_[8880]_  = ~\new_[12290]_  | ~\new_[10754]_  | ~\new_[11001]_  | ~\new_[11736]_ ;
  assign \new_[8881]_  = ~\new_[9132]_ ;
  assign \new_[8882]_  = ~\new_[9134]_ ;
  assign \new_[8883]_  = ~\new_[14116]_ ;
  assign \new_[8884]_  = ~\new_[9135]_ ;
  assign \new_[8885]_  = ~\new_[11580]_  | ~\new_[10241]_  | ~\new_[11095]_  | ~\new_[12372]_ ;
  assign \new_[8886]_  = ~\new_[11618]_  | ~\new_[10245]_  | ~\new_[11097]_  | ~\new_[11269]_ ;
  assign \new_[8887]_  = ~\new_[9137]_ ;
  assign \new_[8888]_  = ~\new_[9138]_ ;
  assign \new_[8889]_  = ~\new_[10740]_  | ~\new_[11634]_  | ~\new_[10979]_  | ~\new_[10178]_ ;
  assign \new_[8890]_  = ~\new_[12279]_  | ~\new_[11246]_  | ~\new_[11123]_  | ~\new_[10908]_ ;
  assign \new_[8891]_  = ~\new_[9139]_ ;
  assign \new_[8892]_  = ~\new_[12405]_  | ~\new_[11138]_  | ~\new_[10985]_  | ~\new_[11265]_ ;
  assign \new_[8893]_  = ~\new_[12401]_  | ~\new_[11162]_  | ~\new_[10213]_  | ~\new_[10844]_ ;
  assign \new_[8894]_  = ~\new_[12282]_  | ~\new_[10510]_  | ~\new_[10221]_  | ~\new_[10992]_ ;
  assign \new_[8895]_  = ~\new_[12270]_  | ~\new_[10980]_  | ~\new_[10266]_  | ~\new_[11700]_ ;
  assign \new_[8896]_  = ~\new_[9141]_ ;
  assign \new_[8897]_  = ~\new_[12281]_  | ~\new_[11037]_  | ~\new_[10269]_  | ~\new_[11687]_ ;
  assign \new_[8898]_  = ~\new_[12274]_  | ~\new_[11057]_  | ~\new_[10232]_  | ~\new_[11172]_ ;
  assign \new_[8899]_  = ~\new_[11590]_  | ~\new_[11228]_  | ~\new_[10772]_  | ~\new_[10761]_ ;
  assign \new_[8900]_  = ~\new_[12278]_  | ~\new_[11175]_  | ~\new_[10271]_  | ~\new_[11654]_ ;
  assign \new_[8901]_  = ~\new_[12467]_  | ~\new_[10916]_  | ~\new_[10202]_  | ~\new_[12309]_ ;
  assign \new_[8902]_  = ~\new_[12280]_  | ~\new_[11185]_  | ~\new_[10208]_  | ~\new_[11692]_ ;
  assign \new_[8903]_  = ~\new_[9142]_ ;
  assign \new_[8904]_  = ~\new_[10719]_  | ~\new_[10775]_  | ~\new_[12293]_  | ~\new_[10746]_ ;
  assign \new_[8905]_  = ~\new_[12218]_  | ~\new_[11100]_  | ~\new_[10729]_  | ~\new_[10964]_ ;
  assign \new_[8906]_  = ~\new_[12295]_  | ~\new_[11233]_  | ~\new_[10828]_  | ~\new_[11013]_ ;
  assign \new_[8907]_  = ~\new_[12296]_  | ~\new_[10965]_  | ~\new_[10750]_  | ~\new_[11276]_ ;
  assign \new_[8908]_  = ~\new_[12423]_  | ~\new_[10906]_  | ~\new_[10914]_  | ~\new_[11134]_ ;
  assign \new_[8909]_  = ~\new_[11599]_  | ~\new_[10874]_  | ~\new_[10925]_  | ~\new_[11474]_ ;
  assign \new_[8910]_  = ~\new_[9143]_ ;
  assign \new_[8911]_  = ~\new_[12292]_  | ~\new_[11252]_  | ~\new_[11182]_  | ~\new_[11084]_ ;
  assign \new_[8912]_  = ~\new_[10730]_  | ~\new_[11737]_  | ~\new_[11227]_  | ~\new_[10253]_ ;
  assign \new_[8913]_  = ~\new_[12299]_  | ~\new_[11038]_  | ~\new_[10846]_  | ~\new_[10971]_ ;
  assign \new_[8914]_  = ~\new_[9145]_ ;
  assign \new_[8915]_  = ~\new_[11739]_  | ~\new_[10827]_  | ~\new_[11558]_  | ~\new_[10832]_ ;
  assign \new_[8916]_  = ~\new_[9146]_ ;
  assign \new_[8917]_  = ~\new_[9147]_ ;
  assign \new_[8918]_  = ~\new_[11603]_  | ~\new_[10951]_  | ~\new_[10783]_  | ~\new_[11232]_ ;
  assign \new_[8919]_  = ~\new_[12297]_  | ~\new_[11031]_  | ~\new_[10984]_  | ~\new_[12318]_ ;
  assign \new_[8920]_  = ~\new_[9148]_ ;
  assign \new_[8921]_  = ~\new_[11604]_  | ~\new_[10847]_  | ~\new_[10839]_  | ~\new_[11755]_ ;
  assign \new_[8922]_  = ~\new_[9149]_ ;
  assign \new_[8923]_  = ~\new_[11596]_  | ~\new_[11249]_  | ~\new_[10875]_  | ~\new_[12313]_ ;
  assign \new_[8924]_  = ~\new_[9150]_ ;
  assign \new_[8925]_  = ~\new_[12037]_  | ~\new_[11274]_  | ~\new_[11637]_  | ~\new_[10476]_ ;
  assign \new_[8926]_  = ~\new_[11566]_  | ~\new_[11277]_  | ~\new_[10936]_  | ~\new_[11051]_ ;
  assign \new_[8927]_  = ~\new_[11611]_  | ~\new_[11208]_  | ~\new_[10920]_  | ~\new_[11536]_ ;
  assign \new_[8928]_  = ~\new_[9151]_ ;
  assign \new_[8929]_  = ~\new_[9152]_ ;
  assign \new_[8930]_  = ~\new_[12388]_  | ~\new_[10826]_  | ~\new_[11022]_  | ~\new_[11210]_ ;
  assign \new_[8931]_  = ~\new_[11624]_  | ~\new_[11278]_  | ~\new_[11280]_  | ~\new_[12046]_ ;
  assign \new_[8932]_  = ~\new_[9643]_  | ~\new_[12534]_ ;
  assign \new_[8933]_  = ~\new_[9834]_  | ~\new_[10863]_ ;
  assign \new_[8934]_  = ~\new_[9835]_  | ~\new_[10848]_ ;
  assign \new_[8935]_  = ~\new_[9832]_  | ~\new_[11723]_ ;
  assign \new_[8936]_  = ~\new_[9831]_  | ~\new_[11635]_ ;
  assign \new_[8937]_  = ~\new_[9840]_  | ~\new_[11728]_ ;
  assign \new_[8938]_  = ~\new_[9836]_  | ~\new_[10973]_ ;
  assign \new_[8939]_  = ~\new_[9838]_  | ~\new_[10866]_ ;
  assign \new_[8940]_  = ~\new_[9839]_  | ~\new_[10753]_ ;
  assign \new_[8941]_  = ~\new_[9867]_  | ~\new_[11190]_ ;
  assign \new_[8942]_  = ~\new_[9847]_  | ~\new_[10904]_ ;
  assign \new_[8943]_  = ~\new_[9837]_  | ~\new_[10818]_ ;
  assign \new_[8944]_  = ~\new_[9785]_  & (~\new_[13860]_  | ~\new_[12828]_ );
  assign \new_[8945]_  = ~\new_[9821]_  & (~\new_[13204]_  | ~\new_[12828]_ );
  assign \new_[8946]_  = ~\new_[9822]_  & (~\new_[13849]_  | ~\new_[12828]_ );
  assign \new_[8947]_  = ~\new_[9793]_  & (~\new_[13313]_  | ~\new_[12432]_ );
  assign \new_[8948]_  = ~\new_[9795]_  & (~\new_[13319]_  | ~\new_[12432]_ );
  assign \new_[8949]_  = ~\new_[9796]_  & (~\new_[13572]_  | ~\new_[12432]_ );
  assign \new_[8950]_  = ~\new_[9798]_  & (~\new_[13321]_  | ~\new_[12432]_ );
  assign \new_[8951]_  = ~\new_[9799]_  & (~\new_[13363]_  | ~\new_[12432]_ );
  assign \new_[8952]_  = ~\new_[9801]_  & (~\new_[13560]_  | ~\new_[12432]_ );
  assign \new_[8953]_  = ~\new_[9814]_  & (~\new_[13238]_  | ~\new_[12828]_ );
  assign \new_[8954]_  = ~\new_[9802]_  & (~\new_[13360]_  | ~\new_[12432]_ );
  assign \new_[8955]_  = ~\new_[9803]_  & (~\new_[13549]_  | ~\new_[12432]_ );
  assign \new_[8956]_  = ~\new_[9817]_  & (~\new_[13776]_  | ~\new_[12828]_ );
  assign \new_[8957]_  = ~\new_[9806]_  & (~\new_[13427]_  | ~\new_[12828]_ );
  assign \new_[8958]_  = ~\new_[9808]_  & (~\new_[13764]_  | ~\new_[12828]_ );
  assign \new_[8959]_  = ~\new_[9820]_  & (~\new_[13258]_  | ~\new_[12828]_ );
  assign \new_[8960]_  = ~\new_[9819]_  & (~\new_[13616]_  | ~\new_[12828]_ );
  assign \new_[8961]_  = ~\new_[9809]_  & (~\new_[13252]_  | ~\new_[12828]_ );
  assign \new_[8962]_  = ~\new_[9807]_  & (~\new_[13847]_  | ~\new_[12828]_ );
  assign \new_[8963]_  = ~\new_[9804]_  & (~\new_[13763]_  | ~\new_[12828]_ );
  assign \new_[8964]_  = ~\new_[9811]_  | (~\new_[3567]_  & ~\new_[12027]_ );
  assign \new_[8965]_  = ~\new_[9812]_  | (~\new_[3557]_  & ~\new_[12027]_ );
  assign \new_[8966]_  = ~\new_[9786]_  | (~\new_[3558]_  & ~\new_[12027]_ );
  assign \new_[8967]_  = ~\new_[9787]_  | (~\new_[3560]_  & ~\new_[12027]_ );
  assign \new_[8968]_  = ~\new_[9783]_  | (~\new_[3561]_  & ~\new_[12655]_ );
  assign \new_[8969]_  = ~\new_[9800]_  | (~\new_[3562]_  & ~\new_[12655]_ );
  assign \new_[8970]_  = ~\new_[9788]_  | (~\new_[3406]_  & ~\new_[12027]_ );
  assign \new_[8971]_  = ~\new_[9792]_  | (~\new_[3563]_  & ~\new_[12027]_ );
  assign \new_[8972]_  = ~\new_[9790]_  | (~\new_[3564]_  & ~\new_[12027]_ );
  assign \new_[8973]_  = ~\new_[9791]_  | (~\new_[3565]_  & ~\new_[12027]_ );
  assign \new_[8974]_  = ~\new_[9789]_  | (~\new_[3566]_  & ~\new_[12027]_ );
  assign \new_[8975]_  = ~\new_[9815]_  | (~\new_[3319]_  & ~\new_[12028]_ );
  assign \new_[8976]_  = ~\new_[9816]_  | (~\new_[3331]_  & ~\new_[12028]_ );
  assign \new_[8977]_  = ~\new_[9810]_  | (~\new_[3332]_  & ~\new_[12028]_ );
  assign \new_[8978]_  = ~\new_[9805]_  | (~\new_[3334]_  & ~\new_[12028]_ );
  assign \new_[8979]_  = ~\new_[9818]_  | (~\new_[3559]_  & ~\new_[12027]_ );
  assign \new_[8980]_  = ~\new_[9644]_  | (~\new_[12029]_  & ~\new_[2791]_ );
  assign \new_[8981]_  = ~\new_[10212]_  | ~\new_[10953]_ ;
  assign \new_[8982]_  = ~\new_[12269]_  | ~\new_[10270]_ ;
  assign \new_[8983]_  = ~\new_[10200]_  | ~\new_[10840]_ ;
  assign \new_[8984]_  = ~\new_[12276]_  | ~\new_[10256]_ ;
  assign \new_[8985]_  = ~\new_[10193]_  | ~\new_[11179]_ ;
  assign \new_[8986]_  = ~\new_[10272]_  | ~\new_[11531]_ ;
  assign \new_[8987]_  = ~\new_[10209]_  | ~\new_[10934]_ ;
  assign \new_[8988]_  = ~\new_[12289]_  | ~\new_[10278]_ ;
  assign \new_[8989]_  = ~\new_[10230]_  | ~\new_[10752]_ ;
  assign \new_[8990]_  = ~\new_[10194]_  | ~\new_[11099]_ ;
  assign \new_[8991]_  = ~\new_[12286]_  | ~\new_[10268]_ ;
  assign \new_[8992]_  = ~\new_[12386]_  | ~\new_[10251]_ ;
  assign \new_[8993]_  = ~\new_[10297]_  | (~\new_[12077]_  & ~\new_[7956]_ );
  assign n10351 = \new_[12000]_  ^ \new_[11442]_ ;
  assign \new_[8995]_  = u10_full_reg;
  assign \new_[8996]_  = ~\\u2_out_le_reg[2] ;
  assign \new_[8997]_  = \new_[7972]_  ^ \new_[11427]_ ;
  assign \new_[8998]_  = ~\new_[10436]_  & (~\new_[12257]_  | ~\new_[12618]_ );
  assign \new_[8999]_  = (~n10936 | ~\new_[7936]_ ) & (~\new_[12119]_  | ~\new_[12083]_ );
  assign \new_[9000]_  = ~\\u2_out_le_reg[4] ;
  assign \new_[9001]_  = ~\\u2_out_le_reg[5] ;
  assign \new_[9002]_  = ~\\u2_out_le_reg[3] ;
  assign \new_[9003]_  = ~\new_[13047]_  | ~\new_[10306]_  | ~\new_[12928]_ ;
  assign n10366 = ~\new_[10303]_  & ~\new_[12347]_ ;
  assign n10361 = ~\new_[10394]_  | ~\new_[10309]_ ;
  assign \new_[9006]_  = \\u2_out_le_reg[0] ;
  assign \new_[9007]_  = \\u9_dout_reg[11] ;
  assign \new_[9008]_  = \\u9_dout_reg[14] ;
  assign \new_[9009]_  = \\u9_dout_reg[18] ;
  assign \new_[9010]_  = \\u9_dout_reg[19] ;
  assign \new_[9011]_  = \\u9_dout_reg[20] ;
  assign \new_[9012]_  = \\u9_dout_reg[21] ;
  assign \new_[9013]_  = \\u9_dout_reg[22] ;
  assign \new_[9014]_  = \\u9_dout_reg[23] ;
  assign \new_[9015]_  = \\u9_dout_reg[24] ;
  assign \new_[9016]_  = \\u9_dout_reg[25] ;
  assign \new_[9017]_  = \\u9_dout_reg[16] ;
  assign \new_[9018]_  = \\u10_dout_reg[16] ;
  assign \new_[9019]_  = \\u9_dout_reg[26] ;
  assign \new_[9020]_  = \\u9_dout_reg[27] ;
  assign \new_[9021]_  = \\u9_dout_reg[28] ;
  assign \new_[9022]_  = \\u9_dout_reg[29] ;
  assign \new_[9023]_  = \\u9_dout_reg[2] ;
  assign \new_[9024]_  = \\u9_dout_reg[30] ;
  assign \new_[9025]_  = \\u9_dout_reg[31] ;
  assign \new_[9026]_  = \\u9_dout_reg[3] ;
  assign n10336 = \\u1_sr_reg[3] ;
  assign \new_[9028]_  = \\u9_dout_reg[4] ;
  assign \new_[9029]_  = \\u9_dout_reg[5] ;
  assign \new_[9030]_  = \\u9_dout_reg[6] ;
  assign \new_[9031]_  = \\u9_dout_reg[7] ;
  assign \new_[9032]_  = \\u9_dout_reg[8] ;
  assign \new_[9033]_  = \\u9_dout_reg[9] ;
  assign \new_[9034]_  = \\u10_dout_reg[24] ;
  assign \new_[9035]_  = \\u10_dout_reg[26] ;
  assign \new_[9036]_  = \\u9_dout_reg[13] ;
  assign \new_[9037]_  = \\u11_dout_reg[0] ;
  assign \new_[9038]_  = \\u11_dout_reg[10] ;
  assign \new_[9039]_  = \\u11_dout_reg[11] ;
  assign \new_[9040]_  = \\u11_dout_reg[12] ;
  assign \new_[9041]_  = \\u11_dout_reg[13] ;
  assign \new_[9042]_  = \\u10_dout_reg[31] ;
  assign \new_[9043]_  = \\u11_dout_reg[14] ;
  assign \new_[9044]_  = \\u11_dout_reg[15] ;
  assign \new_[9045]_  = \\u11_dout_reg[16] ;
  assign \new_[9046]_  = \\u11_dout_reg[17] ;
  assign \new_[9047]_  = \\u11_dout_reg[18] ;
  assign \new_[9048]_  = \\u11_dout_reg[19] ;
  assign \new_[9049]_  = \\u10_dout_reg[5] ;
  assign \new_[9050]_  = \\u11_dout_reg[1] ;
  assign \new_[9051]_  = \\u11_dout_reg[20] ;
  assign \new_[9052]_  = \\u11_dout_reg[21] ;
  assign \new_[9053]_  = \\u11_dout_reg[22] ;
  assign \new_[9054]_  = \\u11_dout_reg[23] ;
  assign \new_[9055]_  = \\u11_dout_reg[24] ;
  assign \new_[9056]_  = \\u11_dout_reg[25] ;
  assign \new_[9057]_  = \\u11_dout_reg[26] ;
  assign \new_[9058]_  = \\u11_dout_reg[27] ;
  assign \new_[9059]_  = \\u11_dout_reg[28] ;
  assign \new_[9060]_  = \\u11_dout_reg[29] ;
  assign \new_[9061]_  = \\u11_dout_reg[2] ;
  assign \new_[9062]_  = \\u11_dout_reg[30] ;
  assign \new_[9063]_  = \\u11_dout_reg[31] ;
  assign \new_[9064]_  = \\u11_dout_reg[3] ;
  assign \new_[9065]_  = \\u11_dout_reg[4] ;
  assign \new_[9066]_  = \\u11_dout_reg[5] ;
  assign \new_[9067]_  = \\u11_dout_reg[6] ;
  assign \new_[9068]_  = \\u11_dout_reg[7] ;
  assign \new_[9069]_  = \\u11_dout_reg[8] ;
  assign \new_[9070]_  = \\u11_dout_reg[9] ;
  assign \new_[9071]_  = \\u9_dout_reg[15] ;
  assign \new_[9072]_  = \\u9_dout_reg[17] ;
  assign \new_[9073]_  = \\u9_dout_reg[0] ;
  assign \new_[9074]_  = \\u9_dout_reg[12] ;
  assign \new_[9075]_  = \\u9_dout_reg[10] ;
  assign \new_[9076]_  = \\u9_dout_reg[1] ;
  assign \new_[9077]_  = ~\new_[9661]_ ;
  assign \new_[9078]_  = ~\new_[10438]_  | ~\new_[11532]_ ;
  assign \new_[9079]_  = ~\new_[13070]_  & ~\new_[10317]_ ;
  assign \new_[9080]_  = ~\new_[12085]_  & ~\new_[12710]_ ;
  assign \new_[9081]_  = ~\new_[12086]_  & ~\new_[14093]_ ;
  assign \new_[9082]_  = ~\new_[10317]_  & ~\new_[13877]_ ;
  assign n10341 = \new_[10390]_  & \new_[7807]_ ;
  assign n10346 = \new_[11441]_  ^ \new_[12001]_ ;
  assign \new_[9085]_  = ~\new_[7807]_  & (~\new_[11468]_  | ~\new_[7977]_ );
  assign \new_[9086]_  = \new_[3025]_  ? \new_[12030]_  : \new_[11506]_ ;
  assign \new_[9087]_  = \new_[3187]_  ? \new_[12871]_  : \new_[11500]_ ;
  assign \new_[9088]_  = \new_[3188]_  ? \new_[12871]_  : \new_[11508]_ ;
  assign \new_[9089]_  = \new_[3249]_  ? \new_[12837]_  : \new_[11508]_ ;
  assign \new_[9090]_  = ~\new_[10354]_  | (~\new_[12618]_  & ~\new_[12991]_ );
  assign \new_[9091]_  = \new_[3138]_  ? \new_[12028]_  : \new_[11500]_ ;
  assign \new_[9092]_  = \new_[3026]_  ? \new_[12030]_  : \new_[11507]_ ;
  assign \new_[9093]_  = \new_[3247]_  ? \new_[12028]_  : \new_[11508]_ ;
  assign \new_[9094]_  = \new_[3027]_  ? \new_[12716]_  : \new_[11506]_ ;
  assign \new_[9095]_  = \new_[3041]_  ? \new_[12758]_  : \new_[11506]_ ;
  assign \new_[9096]_  = \new_[3042]_  ? \new_[12758]_  : \new_[11507]_ ;
  assign \new_[9097]_  = \new_[3248]_  ? \new_[12837]_  : \new_[11500]_ ;
  assign \new_[9098]_  = \new_[3028]_  ? \new_[12716]_  : \new_[11507]_ ;
  assign \new_[9099]_  = (~n10936 | ~\new_[7975]_ ) & (~\new_[12119]_  | ~\new_[12878]_ );
  assign \new_[9100]_  = \new_[7974]_  ^ n10936;
  assign \new_[9101]_  = ~suspended_o;
  assign \new_[9102]_  = ~\new_[11602]_  | ~\new_[11629]_  | ~\new_[10801]_  | ~\new_[10802]_ ;
  assign \new_[9103]_  = ~\new_[12412]_  | ~\new_[10890]_  | ~\new_[11675]_  | ~\new_[10976]_ ;
  assign n10376 = ~\new_[12171]_  | ~\new_[10445]_ ;
  assign n10381 = ~\new_[10311]_  | ~\new_[12487]_ ;
  assign n10386 = ~\new_[12175]_  | ~\new_[10447]_ ;
  assign n10391 = ~\new_[10448]_  | ~\new_[12488]_ ;
  assign n10396 = ~\new_[12177]_  | ~\new_[10449]_ ;
  assign n10401 = ~\new_[10450]_  | ~\new_[12489]_ ;
  assign n10406 = ~\new_[10451]_  | ~\new_[12490]_ ;
  assign n10411 = ~\new_[11478]_  | ~\new_[10453]_ ;
  assign n10416 = ~\new_[10454]_  | ~\new_[12491]_ ;
  assign \new_[9113]_  = ~\new_[12038]_  | ~\new_[11511]_  | ~\new_[11418]_  | ~\new_[11061]_ ;
  assign \new_[9114]_  = ~\new_[12422]_  | ~\new_[10921]_  | ~\new_[11658]_  | ~\new_[10922]_ ;
  assign \new_[9115]_  = ~\new_[12271]_  | ~\new_[11521]_  | ~\new_[10928]_  | ~\new_[10929]_ ;
  assign \new_[9116]_  = ~\new_[12410]_  | ~\new_[11659]_  | ~\new_[11223]_  | ~\new_[10930]_ ;
  assign \new_[9117]_  = ~\new_[12272]_  | ~\new_[11519]_  | ~\new_[11132]_  | ~\new_[10935]_ ;
  assign \new_[9118]_  = ~\new_[12421]_  | ~\new_[10939]_  | ~\new_[10940]_  | ~\new_[11664]_ ;
  assign \new_[9119]_  = ~\new_[12277]_  | ~\new_[10944]_  | ~\new_[11186]_  | ~\new_[11741]_ ;
  assign \new_[9120]_  = ~\new_[12416]_  | ~\new_[11667]_  | ~\new_[11262]_  | ~\new_[10956]_ ;
  assign \new_[9121]_  = ~\new_[12414]_  | ~\new_[11114]_  | ~\new_[11264]_  | ~\new_[11670]_ ;
  assign \new_[9122]_  = ~\new_[11587]_  | ~\new_[11096]_  | ~\new_[11671]_  | ~\new_[10969]_ ;
  assign \new_[9123]_  = ~\new_[12415]_  | ~\new_[10970]_  | ~\new_[11646]_  | ~\new_[12426]_ ;
  assign \new_[9124]_  = ~\new_[11564]_  | ~\new_[10993]_  | ~\new_[11672]_  | ~\new_[10975]_ ;
  assign \new_[9125]_  = ~\new_[10402]_  & ~\new_[10418]_ ;
  assign n10356 = ~\new_[10307]_  & ~\new_[11436]_ ;
  assign n10371 = ~\new_[11475]_  | ~\new_[10444]_ ;
  assign \new_[9128]_  = ~\new_[11569]_  | ~\new_[11756]_  | ~\new_[11052]_  | ~\new_[10185]_ ;
  assign \new_[9129]_  = ~\new_[12043]_  | ~\new_[11529]_  | ~\new_[11055]_  | ~\new_[10224]_ ;
  assign \new_[9130]_  = ~\new_[11571]_  | ~\new_[11695]_  | ~\new_[11217]_  | ~\new_[10222]_ ;
  assign \new_[9131]_  = ~\new_[11572]_  | ~\new_[12093]_  | ~\new_[11448]_  | ~\new_[10211]_ ;
  assign \new_[9132]_  = ~\new_[11556]_  | ~\new_[11699]_  | ~\new_[10892]_  | ~\new_[10236]_ ;
  assign \new_[9133]_  = ~\new_[11567]_  | ~\new_[11694]_  | ~\new_[11070]_  | ~\new_[11256]_ ;
  assign \new_[9134]_  = ~\new_[11574]_  | ~\new_[11703]_  | ~\new_[10687]_  | ~\new_[10169]_ ;
  assign \new_[9135]_  = ~\new_[11575]_  | ~\new_[11717]_  | ~\new_[10796]_  | ~\new_[10234]_ ;
  assign \new_[9136]_  = ~\new_[11588]_  | ~\new_[11709]_  | ~\new_[10243]_  | ~\new_[11032]_ ;
  assign \new_[9137]_  = ~\new_[11582]_  | ~\new_[11707]_  | ~\new_[11012]_  | ~\new_[10284]_ ;
  assign \new_[9138]_  = ~\new_[11598]_  | ~\new_[11712]_  | ~\new_[11008]_  | ~\new_[10225]_ ;
  assign \new_[9139]_  = ~\new_[11609]_  | ~\new_[11730]_  | ~\new_[11129]_  | ~\new_[11160]_ ;
  assign \new_[9140]_  = ~\new_[12283]_  | ~\new_[12094]_  | ~\new_[11164]_  | ~\new_[11033]_ ;
  assign \new_[9141]_  = ~\new_[12285]_  | ~\new_[11520]_  | ~\new_[11167]_  | ~\new_[11048]_ ;
  assign \new_[9142]_  = ~\new_[12301]_  | ~\new_[11537]_  | ~\new_[11047]_  | ~\new_[11187]_ ;
  assign \new_[9143]_  = ~\new_[11608]_  | ~\new_[11746]_  | ~\new_[11006]_  | ~\new_[11053]_ ;
  assign \new_[9144]_  = u12_re2_reg;
  assign \new_[9145]_  = ~\new_[11601]_  | ~\new_[11738]_  | ~\new_[11226]_  | ~\new_[11101]_ ;
  assign \new_[9146]_  = ~\new_[11551]_  | ~\new_[11647]_  | ~\new_[11287]_  | ~\new_[10952]_ ;
  assign \new_[9147]_  = ~\new_[11549]_  | ~\new_[11636]_  | ~\new_[10791]_  | ~\new_[10792]_ ;
  assign \new_[9148]_  = ~\new_[11621]_  | ~\new_[11682]_  | ~\new_[11271]_  | ~\new_[11234]_ ;
  assign \new_[9149]_  = ~\new_[12031]_  | ~\new_[11834]_  | ~\new_[11417]_  | ~\new_[10856]_ ;
  assign \new_[9150]_  = ~\new_[11605]_  | ~\new_[12044]_  | ~\new_[11239]_  | ~\new_[11243]_ ;
  assign \new_[9151]_  = ~\new_[11613]_  | ~\new_[12005]_  | ~\new_[11125]_  | ~\new_[11014]_ ;
  assign \new_[9152]_  = ~\new_[11614]_  | ~\new_[11686]_  | ~\new_[10860]_  | ~\new_[11263]_ ;
  assign \new_[9153]_  = ~\new_[10158]_  | ~\new_[12267]_ ;
  assign \new_[9154]_  = ~\new_[10160]_  | ~\new_[11523]_ ;
  assign \new_[9155]_  = ~\new_[10159]_  & ~\new_[13930]_ ;
  assign \new_[9156]_  = ~\new_[10161]_  | ~\new_[14137]_ ;
  assign \new_[9157]_  = ~\new_[9889]_  | ~\new_[12024]_ ;
  assign \new_[9158]_  = ~\new_[10443]_  | ~\new_[12009]_ ;
  assign \new_[9159]_  = ~\new_[10442]_  | ~\new_[10786]_ ;
  assign \new_[9160]_  = ~\new_[10441]_  | ~\new_[11067]_ ;
  assign \new_[9161]_  = ~\new_[10440]_  | ~\new_[10955]_ ;
  assign \new_[9162]_  = ~\new_[10439]_  | ~\new_[10865]_ ;
  assign \new_[9163]_  = ~\new_[11476]_  | ~\new_[10195]_ ;
  assign \new_[9164]_  = ~\new_[11426]_  | ~\new_[10180]_ ;
  assign \new_[9165]_  = ~\new_[10464]_  | ~\new_[11702]_ ;
  assign \new_[9166]_  = ~\new_[10452]_  | ~\new_[11701]_ ;
  assign \new_[9167]_  = ~\new_[10459]_  | ~\new_[11633]_ ;
  assign \new_[9168]_  = ~\new_[10460]_  | ~\new_[11742]_ ;
  assign \new_[9169]_  = ~\new_[10461]_  | ~\new_[12106]_ ;
  assign \new_[9170]_  = ~\new_[10462]_  | ~\new_[11711]_ ;
  assign \new_[9171]_  = ~\new_[10463]_  | ~\new_[11715]_ ;
  assign \new_[9172]_  = ~\new_[10465]_  | ~\new_[11643]_ ;
  assign \new_[9173]_  = ~\new_[10466]_  | ~\new_[12254]_ ;
  assign \new_[9174]_  = ~\new_[10467]_  | ~\new_[11757]_ ;
  assign \new_[9175]_  = ~\new_[10468]_  | ~\new_[11693]_ ;
  assign \new_[9176]_  = ~\new_[10470]_  | ~\new_[11657]_ ;
  assign \new_[9177]_  = ~\new_[10469]_  | ~\new_[11714]_ ;
  assign \new_[9178]_  = ~\new_[10471]_  | ~\new_[11538]_ ;
  assign \new_[9179]_  = ~\new_[10472]_  | ~\new_[11655]_ ;
  assign \new_[9180]_  = ~\new_[9883]_  | ~\new_[11732]_ ;
  assign \new_[9181]_  = ~\new_[9884]_  | ~\new_[11685]_ ;
  assign \new_[9182]_  = ~\new_[9885]_  | ~\new_[11731]_ ;
  assign \new_[9183]_  = ~\new_[9886]_  | ~\new_[11734]_ ;
  assign \new_[9184]_  = ~\new_[9887]_  | ~\new_[11735]_ ;
  assign \new_[9185]_  = ~\new_[9888]_  | ~\new_[11691]_ ;
  assign \new_[9186]_  = ~\new_[9890]_  | ~\new_[11743]_ ;
  assign \new_[9187]_  = ~\new_[10446]_  | ~\new_[11676]_ ;
  assign \new_[9188]_  = ~\new_[9895]_  | ~\new_[11651]_ ;
  assign \new_[9189]_  = ~\new_[9891]_  | ~\new_[12105]_ ;
  assign \new_[9190]_  = ~\new_[10294]_  | ~\new_[11745]_ ;
  assign \new_[9191]_  = \new_[3040]_  ? \new_[12626]_  : \new_[11087]_ ;
  assign \new_[9192]_  = \new_[3189]_  ? \new_[12574]_  : \new_[11439]_ ;
  assign \new_[9193]_  = \new_[3191]_  ? \new_[12871]_  : \new_[11028]_ ;
  assign \new_[9194]_  = \new_[3161]_  ? \new_[12574]_  : \new_[10804]_ ;
  assign \new_[9195]_  = \new_[3195]_  ? \new_[12574]_  : \new_[11154]_ ;
  assign \new_[9196]_  = ~\new_[10305]_  & (~\new_[13297]_  | ~\new_[12513]_ );
  assign \new_[9197]_  = ~\new_[10430]_  & (~\new_[13685]_  | ~\new_[12513]_ );
  assign \new_[9198]_  = ~\new_[10419]_  & (~\new_[13374]_  | ~\new_[12513]_ );
  assign \new_[9199]_  = ~\new_[10428]_  & (~\new_[13305]_  | ~\new_[12513]_ );
  assign \new_[9200]_  = ~\new_[10426]_  & (~\new_[13693]_  | ~\new_[12513]_ );
  assign \new_[9201]_  = ~\new_[10422]_  & (~\new_[13578]_  | ~\new_[12432]_ );
  assign \new_[9202]_  = \new_[3260]_  ? \new_[12663]_  : \new_[11258]_ ;
  assign n10331 = \new_[12456]_  & \new_[10310]_ ;
  assign \new_[9204]_  = ~\new_[10423]_  & (~\new_[13564]_  | ~\new_[12432]_ );
  assign \new_[9205]_  = ~\new_[10424]_  & (~\new_[13325]_  | ~\new_[12432]_ );
  assign \new_[9206]_  = \new_[3254]_  ? \new_[12663]_  : \new_[11154]_ ;
  assign \new_[9207]_  = ~\new_[10425]_  & (~\new_[13511]_  | ~\new_[12432]_ );
  assign \new_[9208]_  = ~\new_[10427]_  & (~\new_[13309]_  | ~\new_[12513]_ );
  assign \new_[9209]_  = \new_[3261]_  ? \new_[12663]_  : \new_[10876]_ ;
  assign \new_[9210]_  = ~\new_[10420]_  & (~\new_[13609]_  | ~\new_[12513]_ );
  assign \new_[9211]_  = ~\new_[10421]_  & (~\new_[13307]_  | ~\new_[12513]_ );
  assign \new_[9212]_  = ~\new_[10429]_  & (~\new_[13298]_  | ~\new_[12513]_ );
  assign \new_[9213]_  = \new_[3206]_  ? \new_[12574]_  : \new_[11106]_ ;
  assign \new_[9214]_  = \new_[3214]_  ? \new_[12871]_  : \new_[10876]_ ;
  assign \new_[9215]_  = \new_[3039]_  ? \new_[12716]_  : \new_[11484]_ ;
  assign \new_[9216]_  = \new_[3043]_  ? \new_[12642]_  : \new_[10769]_ ;
  assign \new_[9217]_  = \new_[3029]_  ? \new_[12716]_  : \new_[10769]_ ;
  assign \new_[9218]_  = ~\new_[10431]_  & (~\new_[13301]_  | ~\new_[12513]_ );
  assign \new_[9219]_  = \new_[3031]_  ? \new_[12626]_  : \new_[10790]_ ;
  assign \new_[9220]_  = \new_[3211]_  ? \new_[12574]_  : \new_[11258]_ ;
  assign \new_[9221]_  = \new_[3032]_  ? \new_[12626]_  : \new_[10770]_ ;
  assign \new_[9222]_  = \new_[3033]_  ? \new_[12626]_  : \new_[11139]_ ;
  assign \new_[9223]_  = \new_[3035]_  ? \new_[12626]_  : \new_[10873]_ ;
  assign \new_[9224]_  = \new_[3038]_  ? \new_[12626]_  : \new_[10869]_ ;
  assign \new_[9225]_  = \new_[3030]_  ? \new_[12626]_  : \new_[10629]_ ;
  assign \new_[9226]_  = \new_[3047]_  ? \new_[12758]_  : \new_[11139]_ ;
  assign \new_[9227]_  = \new_[3037]_  ? \new_[12716]_  : \new_[11011]_ ;
  assign \new_[9228]_  = \new_[3036]_  ? \new_[12626]_  : \new_[11089]_ ;
  assign \new_[9229]_  = \new_[3044]_  ? \new_[12758]_  : \new_[10629]_ ;
  assign \new_[9230]_  = \new_[3045]_  ? \new_[12642]_  : \new_[10790]_ ;
  assign \new_[9231]_  = \new_[3046]_  ? \new_[12642]_  : \new_[10770]_ ;
  assign \new_[9232]_  = \new_[3048]_  ? \new_[12642]_  : \new_[10915]_ ;
  assign \new_[9233]_  = \new_[3049]_  ? \new_[12642]_  : \new_[10873]_ ;
  assign \new_[9234]_  = \new_[3050]_  ? \new_[12642]_  : \new_[11089]_ ;
  assign \new_[9235]_  = \new_[3051]_  ? \new_[12642]_  : \new_[11011]_ ;
  assign \new_[9236]_  = ~\new_[10432]_  & (~\new_[13839]_  | ~\new_[12513]_ );
  assign \new_[9237]_  = \new_[3054]_  ? \new_[12758]_  : \new_[11087]_ ;
  assign \new_[9238]_  = \new_[3052]_  ? \new_[12642]_  : \new_[10869]_ ;
  assign \new_[9239]_  = \new_[3053]_  ? \new_[12758]_  : \new_[11484]_ ;
  assign \new_[9240]_  = ~\new_[10433]_  & (~\new_[13633]_  | ~\new_[12513]_ );
  assign \new_[9241]_  = \new_[3259]_  ? \new_[12663]_  : \new_[11439]_ ;
  assign \new_[9242]_  = \new_[3251]_  ? \new_[12663]_  : \new_[11028]_ ;
  assign \new_[9243]_  = \new_[3252]_  ? \new_[12837]_  : \new_[11416]_ ;
  assign \new_[9244]_  = \new_[3253]_  ? \new_[12663]_  : \new_[10804]_ ;
  assign \new_[9245]_  = \new_[3258]_  ? \new_[12837]_  : \new_[11106]_ ;
  assign \new_[9246]_  = \new_[3194]_  ? \new_[12871]_  : \new_[11416]_ ;
  assign \new_[9247]_  = \new_[3034]_  ? \new_[12716]_  : \new_[10915]_ ;
  assign \new_[9248]_  = (~\new_[12308]_  | ~\new_[5100]_ ) & (~\new_[12500]_  | ~\new_[12057]_ );
  assign \new_[9249]_  = (~\new_[12308]_  | ~\new_[5099]_ ) & (~\new_[12500]_  | ~\new_[12069]_ );
  assign \new_[9250]_  = (~\new_[12308]_  | ~\new_[5109]_ ) & (~\new_[12500]_  | ~\new_[12045]_ );
  assign \new_[9251]_  = ~\new_[9753]_ ;
  assign \new_[9252]_  = (~\new_[12308]_  | ~\new_[5671]_ ) & (~\new_[10819]_  | ~\new_[5694]_ );
  assign \new_[9253]_  = (~\new_[12308]_  | ~\new_[5115]_ ) & (~\new_[10819]_  | ~\new_[5089]_ );
  assign \new_[9254]_  = (~\new_[12308]_  | ~\new_[5117]_ ) & (~\new_[12500]_  | ~\new_[12066]_ );
  assign \new_[9255]_  = (~\new_[12500]_  | ~\new_[5055]_ ) & (~\new_[10819]_  | ~\new_[5093]_ );
  assign \new_[9256]_  = (~\new_[12308]_  | ~\new_[5696]_ ) & (~\new_[12500]_  | ~\new_[12104]_ );
  assign \new_[9257]_  = (~\new_[12308]_  | ~\new_[5121]_ ) & (~\new_[12500]_  | ~\new_[12059]_ );
  assign \new_[9258]_  = (~\new_[12308]_  | ~\new_[5118]_ ) & (~\new_[12500]_  | ~\new_[12075]_ );
  assign \new_[9259]_  = (~\new_[12308]_  | ~\new_[5119]_ ) & (~\new_[12500]_  | ~\new_[11528]_ );
  assign \new_[9260]_  = (~\new_[12308]_  | ~\new_[5043]_ ) & (~\new_[12500]_  | ~\new_[12048]_ );
  assign \new_[9261]_  = (~\new_[12308]_  | ~\new_[5601]_ ) & (~\new_[12500]_  | ~\new_[12060]_ );
  assign \new_[9262]_  = (~\new_[12308]_  | ~\new_[5120]_ ) & (~\new_[12500]_  | ~\new_[11710]_ );
  assign \new_[9263]_  = (~\new_[12308]_  | ~\new_[5102]_ ) & (~\new_[12500]_  | ~\new_[12020]_ );
  assign \new_[9264]_  = (~\new_[12308]_  | ~\new_[5103]_ ) & (~\new_[12500]_  | ~\new_[12065]_ );
  assign \new_[9265]_  = (~\new_[12308]_  | ~\new_[5122]_ ) & (~\new_[12500]_  | ~\new_[12058]_ );
  assign \new_[9266]_  = (~\new_[12308]_  | ~\new_[5101]_ ) & (~\new_[12500]_  | ~\new_[12062]_ );
  assign \new_[9267]_  = (~\new_[12308]_  | ~\new_[5104]_ ) & (~\new_[12500]_  | ~\new_[12051]_ );
  assign \new_[9268]_  = ~\new_[9823]_ ;
  assign \new_[9269]_  = ~\new_[12704]_  | ~\new_[10310]_ ;
  assign \new_[9270]_  = ~\new_[12647]_  | ~\new_[10186]_ ;
  assign \new_[9271]_  = ~\new_[12647]_  | ~\new_[10181]_ ;
  assign \new_[9272]_  = ~\new_[12647]_  | ~\new_[10240]_ ;
  assign \new_[9273]_  = ~\new_[12647]_  | ~\new_[10218]_ ;
  assign \new_[9274]_  = ~\new_[12647]_  | ~\new_[10207]_ ;
  assign \new_[9275]_  = ~\new_[12647]_  | ~\new_[10182]_ ;
  assign \new_[9276]_  = ~\new_[12653]_  | ~\new_[10283]_ ;
  assign \new_[9277]_  = ~\new_[12647]_  | ~\new_[10260]_ ;
  assign \new_[9278]_  = ~\new_[12647]_  | ~\new_[10210]_ ;
  assign \new_[9279]_  = ~\new_[12647]_  | ~\new_[10205]_ ;
  assign \new_[9280]_  = ~\new_[12647]_  | ~\new_[10288]_ ;
  assign \new_[9281]_  = ~\new_[12653]_  | ~\new_[10229]_ ;
  assign \new_[9282]_  = ~\new_[12647]_  | ~\new_[10265]_ ;
  assign \new_[9283]_  = ~\new_[12647]_  | ~\new_[10203]_ ;
  assign \new_[9284]_  = ~\new_[12653]_  | ~\new_[10187]_ ;
  assign \new_[9285]_  = ~\new_[12653]_  | ~\new_[10188]_ ;
  assign \new_[9286]_  = ~\new_[12653]_  | ~\new_[10263]_ ;
  assign \new_[9287]_  = ~\new_[12653]_  | ~\new_[10248]_ ;
  assign \new_[9288]_  = ~\new_[12653]_  | ~\new_[10206]_ ;
  assign \new_[9289]_  = ~\new_[12653]_  | ~\new_[10286]_ ;
  assign \new_[9290]_  = ~\new_[10310]_  & ~\new_[13112]_ ;
  assign \new_[9291]_  = ~\new_[10285]_  | ~\new_[11023]_ ;
  assign \new_[9292]_  = ~\new_[10282]_  | ~\new_[10771]_ ;
  assign \new_[9293]_  = ~\new_[10197]_  | ~\new_[11181]_ ;
  assign \new_[9294]_  = ~\new_[10246]_  | ~\new_[11203]_ ;
  assign \new_[9295]_  = ~\new_[10262]_  | ~\new_[11107]_ ;
  assign \new_[9296]_  = ~\new_[10258]_  | ~\new_[10852]_ ;
  assign \new_[9297]_  = ~\new_[10196]_  | ~\new_[10855]_ ;
  assign \new_[9298]_  = ~\new_[10310]_  & ~\wb_addr_i[6] ;
  assign \new_[9299]_  = ~\new_[10247]_  | ~\new_[11105]_ ;
  assign \new_[9300]_  = ~\new_[12288]_  | ~\new_[10184]_ ;
  assign \new_[9301]_  = ~\new_[12418]_  | ~\new_[10233]_ ;
  assign \new_[9302]_  = ~\new_[10264]_  | ~\new_[10814]_ ;
  assign \new_[9303]_  = ~\new_[10226]_  | ~\new_[11367]_ ;
  assign \new_[9304]_  = ~\new_[10214]_  | ~\new_[10990]_ ;
  assign \new_[9305]_  = ~\new_[12275]_  | ~\new_[10274]_ ;
  assign \new_[9306]_  = ~\new_[10227]_  | ~\new_[11000]_ ;
  assign \new_[9307]_  = ~\new_[10235]_  | ~\new_[10905]_ ;
  assign \new_[9308]_  = ~\new_[10237]_  | ~\new_[11063]_ ;
  assign \new_[9309]_  = ~\new_[10192]_  | ~\new_[10803]_ ;
  assign \new_[9310]_  = ~\new_[10277]_  | ~\new_[12253]_ ;
  assign \new_[9311]_  = ~\new_[10239]_  | ~\new_[11074]_ ;
  assign \new_[9312]_  = ~\new_[10189]_  | ~\new_[11076]_ ;
  assign \new_[9313]_  = ~\new_[10275]_  | ~\new_[11163]_ ;
  assign \new_[9314]_  = ~\new_[10250]_  | ~\new_[10781]_ ;
  assign \new_[9315]_  = ~\new_[10176]_  | ~\new_[11086]_ ;
  assign \new_[9316]_  = ~\new_[10242]_  | ~\new_[10749]_ ;
  assign \new_[9317]_  = ~\new_[10201]_  | ~\new_[11140]_ ;
  assign \new_[9318]_  = ~\new_[10255]_  | ~\new_[11102]_ ;
  assign \new_[9319]_  = ~\new_[10183]_  | ~\new_[11049]_ ;
  assign \new_[9320]_  = ~\new_[11216]_  | ~\new_[11268]_ ;
  assign \new_[9321]_  = ~\new_[11568]_  | ~\new_[10889]_ ;
  assign \new_[9322]_  = ~\new_[10861]_  | ~\new_[11174]_ ;
  assign \new_[9323]_  = ~\new_[10724]_  | ~\new_[10831]_ ;
  assign \new_[9324]_  = ~\new_[10763]_  | ~\new_[10776]_ ;
  assign \new_[9325]_  = ~\new_[11565]_  | ~\new_[10881]_ ;
  assign \new_[9326]_  = ~\new_[11192]_  | ~\new_[10825]_ ;
  assign \new_[9327]_  = ~\new_[11616]_  | ~\new_[10983]_ ;
  assign \new_[9328]_  = ~\new_[12092]_  | ~\new_[10765]_ ;
  assign \new_[9329]_  = ~\new_[11098]_  | ~\new_[11130]_ ;
  assign \new_[9330]_  = ~\new_[11543]_  | ~\new_[11035]_ ;
  assign \new_[9331]_  = ~\new_[11253]_  | ~\new_[11149]_ ;
  assign \new_[9332]_  = ~\new_[11238]_  | ~\new_[10518]_ ;
  assign \new_[9333]_  = ~\new_[10498]_  | ~\new_[11021]_ ;
  assign \new_[9334]_  = ~\new_[11550]_  | ~\new_[11230]_ ;
  assign \new_[9335]_  = ~\new_[11131]_  | ~\new_[10808]_ ;
  assign \new_[9336]_  = ~\new_[11600]_  | ~\new_[11279]_ ;
  assign \new_[9337]_  = ~\new_[10816]_  | ~\new_[10789]_ ;
  assign \new_[9338]_  = ~\new_[11619]_  | ~\new_[11235]_ ;
  assign \new_[9339]_  = ~\new_[11272]_  | ~\new_[11002]_ ;
  assign \new_[9340]_  = ~\new_[11257]_  | ~\new_[11248]_ ;
  assign \new_[9341]_  = ~\new_[12091]_  | ~\new_[10800]_ ;
  assign \new_[9342]_  = ~\new_[11212]_  | ~\new_[11194]_ ;
  assign \new_[9343]_  = ~\new_[11004]_  | ~\new_[11159]_ ;
  assign \new_[9344]_  = ~\new_[11540]_  | ~\new_[10495]_ ;
  assign \new_[9345]_  = ~\new_[11586]_  | ~\new_[11254]_ ;
  assign \new_[9346]_  = ~\new_[11073]_  | ~\new_[11079]_ ;
  assign \new_[9347]_  = ~\new_[10821]_  | ~\new_[11066]_ ;
  assign \new_[9348]_  = ~\new_[11561]_  | ~\new_[11214]_ ;
  assign \new_[9349]_  = ~\new_[10962]_  | ~\new_[10745]_ ;
  assign \new_[9350]_  = ~\new_[11615]_  | ~\new_[11092]_ ;
  assign \new_[9351]_  = ~\new_[10977]_  | ~\new_[11111]_ ;
  assign \new_[9352]_  = ~\new_[10911]_  | ~\new_[10780]_ ;
  assign \new_[9353]_  = ~\new_[11046]_  | ~\new_[11224]_ ;
  assign \new_[9354]_  = ~\new_[11281]_  | ~\new_[11137]_ ;
  assign \new_[9355]_  = ~\new_[11330]_  & (~\new_[5136]_  | ~\new_[12582]_ );
  assign \new_[9356]_  = ~\new_[10824]_  & (~\new_[5504]_  | ~\new_[12706]_ );
  assign \new_[9357]_  = ~\new_[11398]_  & (~\new_[5025]_  | ~\new_[12582]_ );
  assign \new_[9358]_  = ~\new_[11405]_  & (~\new_[5143]_  | ~\new_[12582]_ );
  assign \new_[9359]_  = ~\new_[11351]_  & (~\new_[5145]_  | ~\new_[12582]_ );
  assign \new_[9360]_  = ~\new_[11319]_  & (~\new_[5016]_  | ~\new_[12582]_ );
  assign \new_[9361]_  = ~\new_[11358]_  & (~\new_[5148]_  | ~\new_[12582]_ );
  assign \new_[9362]_  = ~\new_[11381]_  & (~\new_[5152]_  | ~\new_[12693]_ );
  assign \new_[9363]_  = ~\new_[11327]_  & (~\new_[5154]_  | ~\new_[12582]_ );
  assign \new_[9364]_  = ~\new_[11408]_  & (~\new_[5156]_  | ~\new_[12582]_ );
  assign \new_[9365]_  = ~\new_[11323]_  & (~\new_[5159]_  | ~\new_[12693]_ );
  assign \new_[9366]_  = ~\new_[11382]_  & (~\new_[5162]_  | ~\new_[12693]_ );
  assign \new_[9367]_  = ~\new_[11080]_  & (~\new_[5518]_  | ~\new_[12706]_ );
  assign \new_[9368]_  = ~\new_[11289]_  & (~\new_[5541]_  | ~\new_[12693]_ );
  assign \new_[9369]_  = ~\new_[11383]_  & (~\new_[5543]_  | ~\new_[12693]_ );
  assign \new_[9370]_  = ~\new_[10858]_  & (~\new_[5212]_  | ~\new_[12784]_ );
  assign \new_[9371]_  = ~\new_[11328]_  & (~\new_[5764]_  | ~\new_[12577]_ );
  assign \new_[9372]_  = ~\new_[11333]_  & (~\new_[5390]_  | ~\new_[12587]_ );
  assign \new_[9373]_  = ~\new_[11148]_  & (~\new_[5201]_  | ~\new_[12784]_ );
  assign \new_[9374]_  = ~\new_[11273]_  & (~\new_[4991]_  | ~\new_[12611]_ );
  assign \new_[9375]_  = ~\new_[11241]_  & (~\new_[5203]_  | ~\new_[12784]_ );
  assign \new_[9376]_  = ~\new_[11009]_  & (~\new_[5204]_  | ~\new_[12784]_ );
  assign \new_[9377]_  = ~\new_[11222]_  & (~\new_[4979]_  | ~\new_[12611]_ );
  assign \new_[9378]_  = ~\new_[10812]_  & (~\new_[5206]_  | ~\new_[12784]_ );
  assign \new_[9379]_  = ~\new_[10830]_  & (~\new_[5209]_  | ~\new_[12784]_ );
  assign \new_[9380]_  = ~\new_[10837]_  & (~\new_[4976]_  | ~\new_[12784]_ );
  assign \new_[9381]_  = ~\new_[10787]_  & (~\new_[5211]_  | ~\new_[12611]_ );
  assign \new_[9382]_  = ~\new_[11356]_  & (~\new_[5453]_  | ~\new_[12689]_ );
  assign \new_[9383]_  = ~\new_[11078]_  & (~\new_[5214]_  | ~\new_[12611]_ );
  assign \new_[9384]_  = ~\new_[10755]_  & (~\new_[5219]_  | ~\new_[12611]_ );
  assign \new_[9385]_  = ~\new_[11244]_  & (~\new_[5217]_  | ~\new_[12611]_ );
  assign \new_[9386]_  = ~\new_[10850]_  & (~\new_[5218]_  | ~\new_[12784]_ );
  assign \new_[9387]_  = ~\new_[10496]_  & (~\new_[4977]_  | ~\new_[12611]_ );
  assign \new_[9388]_  = ~\new_[11311]_  & (~\new_[5138]_  | ~\new_[12693]_ );
  assign \new_[9389]_  = ~\new_[10811]_  & (~\new_[4974]_  | ~\new_[12784]_ );
  assign \new_[9390]_  = ~\new_[11183]_  & (~\new_[5210]_  | ~\new_[12784]_ );
  assign \new_[9391]_  = ~\new_[11322]_  & (~\new_[5463]_  | ~\new_[12689]_ );
  assign \new_[9392]_  = ~\new_[11346]_  & (~\new_[5466]_  | ~\new_[12689]_ );
  assign \new_[9393]_  = ~\new_[11288]_  & (~\new_[5573]_  | ~\new_[12582]_ );
  assign \new_[9394]_  = ~\new_[11251]_  & (~\new_[4969]_  | ~\new_[12784]_ );
  assign \new_[9395]_  = ~\new_[10891]_  & (~\new_[5271]_  | ~\new_[12692]_ );
  assign \new_[9396]_  = ~\new_[11375]_  & (~\new_[5395]_  | ~\new_[12587]_ );
  assign \new_[9397]_  = ~\new_[11403]_  & (~\new_[5721]_  | ~\new_[12660]_ );
  assign \new_[9398]_  = ~\new_[11390]_  & (~\new_[5450]_  | ~\new_[12689]_ );
  assign \new_[9399]_  = ~\new_[10758]_  & (~\new_[5440]_  | ~\new_[12676]_ );
  assign \new_[9400]_  = ~\new_[11338]_  & (~\new_[5393]_  | ~\new_[12587]_ );
  assign \new_[9401]_  = ~\new_[11242]_  & (~\new_[5272]_  | ~\new_[12692]_ );
  assign \new_[9402]_  = ~\new_[10871]_  & (~\new_[5273]_  | ~\new_[12788]_ );
  assign \new_[9403]_  = ~\new_[10894]_  & (~\new_[4923]_  | ~\new_[12692]_ );
  assign \new_[9404]_  = ~\new_[10895]_  & (~\new_[5274]_  | ~\new_[12788]_ );
  assign \new_[9405]_  = ~\new_[10760]_  & (~\new_[5441]_  | ~\new_[12676]_ );
  assign \new_[9406]_  = ~\new_[10514]_  & (~\new_[5275]_  | ~\new_[12788]_ );
  assign \new_[9407]_  = ~\new_[10896]_  & (~\new_[5276]_  | ~\new_[12692]_ );
  assign \new_[9408]_  = ~\new_[11316]_  & (~\new_[5720]_  | ~\new_[12587]_ );
  assign \new_[9409]_  = ~\new_[10806]_  & (~\new_[4922]_  | ~\new_[12692]_ );
  assign \new_[9410]_  = ~\new_[10897]_  & (~\new_[5277]_  | ~\new_[12788]_ );
  assign \new_[9411]_  = ~\new_[10898]_  & (~\new_[5278]_  | ~\new_[12788]_ );
  assign \new_[9412]_  = ~\new_[11177]_  & (~\new_[4975]_  | ~\new_[12784]_ );
  assign \new_[9413]_  = ~\new_[10773]_  & (~\new_[5279]_  | ~\new_[12692]_ );
  assign \new_[9414]_  = ~\new_[11189]_  & (~\new_[5280]_  | ~\new_[12788]_ );
  assign \new_[9415]_  = ~\new_[10756]_  & (~\new_[5281]_  | ~\new_[12692]_ );
  assign \new_[9416]_  = ~\new_[10901]_  & (~\new_[5282]_  | ~\new_[12692]_ );
  assign \new_[9417]_  = ~\new_[11180]_  & (~\new_[5283]_  | ~\new_[12788]_ );
  assign \new_[9418]_  = ~\new_[10902]_  & (~\new_[4914]_  | ~\new_[12788]_ );
  assign \new_[9419]_  = ~\new_[10982]_  & (~\new_[5284]_  | ~\new_[12788]_ );
  assign \new_[9420]_  = ~\new_[10903]_  & (~\new_[5285]_  | ~\new_[12788]_ );
  assign \new_[9421]_  = ~\new_[11201]_  & (~\new_[5286]_  | ~\new_[12788]_ );
  assign \new_[9422]_  = ~\new_[11387]_  & (~\new_[5455]_  | ~\new_[12681]_ );
  assign \new_[9423]_  = ~\new_[10938]_  & (~\new_[4915]_  | ~\new_[12692]_ );
  assign \new_[9424]_  = ~\new_[11173]_  & (~\new_[5287]_  | ~\new_[12692]_ );
  assign \new_[9425]_  = ~\new_[10759]_  & (~\new_[5288]_  | ~\new_[12692]_ );
  assign \new_[9426]_  = ~\new_[11308]_  & (~\new_[5469]_  | ~\new_[12689]_ );
  assign \new_[9427]_  = ~\new_[11247]_  & (~\new_[5289]_  | ~\new_[12788]_ );
  assign \new_[9428]_  = ~\new_[11260]_  & (~\new_[4911]_  | ~\new_[12692]_ );
  assign \new_[9429]_  = ~\new_[10999]_  & (~\new_[5501]_  | ~\new_[12794]_ );
  assign \new_[9430]_  = ~\new_[10913]_  & (~\new_[5290]_  | ~\new_[12692]_ );
  assign \new_[9431]_  = ~\new_[10912]_  & (~\new_[5291]_  | ~\new_[12692]_ );
  assign \new_[9432]_  = ~\new_[10734]_  & (~\new_[5506]_  | ~\new_[12706]_ );
  assign \new_[9433]_  = ~\new_[11178]_  & (~\new_[5292]_  | ~\new_[12692]_ );
  assign \new_[9434]_  = ~\new_[10744]_  & (~\new_[4910]_  | ~\new_[12692]_ );
  assign \new_[9435]_  = ~\new_[11331]_  & (~\new_[5468]_  | ~\new_[12681]_ );
  assign \new_[9436]_  = ~\new_[11170]_  & (~\new_[5293]_  | ~\new_[12788]_ );
  assign \new_[9437]_  = ~\new_[11305]_  & (~\new_[5294]_  | ~\new_[12788]_ );
  assign \new_[9438]_  = ~\new_[10788]_  & (~\new_[5213]_  | ~\new_[12611]_ );
  assign \new_[9439]_  = ~\new_[11143]_  & (~\new_[5295]_  | ~\new_[12788]_ );
  assign \new_[9440]_  = ~\new_[11127]_  & (~\new_[4909]_  | ~\new_[12788]_ );
  assign \new_[9441]_  = ~\new_[11117]_  & (~\new_[5439]_  | ~\new_[12786]_ );
  assign \new_[9442]_  = ~\new_[11136]_  & (~\new_[5438]_  | ~\new_[12676]_ );
  assign \new_[9443]_  = ~\new_[10945]_  & (~\new_[5437]_  | ~\new_[12676]_ );
  assign \new_[9444]_  = ~\new_[10957]_  & (~\new_[5435]_  | ~\new_[12786]_ );
  assign \new_[9445]_  = ~\new_[11326]_  & (~\new_[5444]_  | ~\new_[12676]_ );
  assign \new_[9446]_  = ~\new_[10941]_  & (~\new_[5502]_  | ~\new_[12706]_ );
  assign \new_[9447]_  = ~\new_[10986]_  & (~\new_[5434]_  | ~\new_[12676]_ );
  assign \new_[9448]_  = ~\new_[10989]_  & (~\new_[5433]_  | ~\new_[12786]_ );
  assign \new_[9449]_  = ~\new_[11370]_  & (~\new_[5389]_  | ~\new_[12587]_ );
  assign \new_[9450]_  = ~\new_[10950]_  & (~\new_[5432]_  | ~\new_[12786]_ );
  assign \new_[9451]_  = ~\new_[10994]_  & (~\new_[5675]_  | ~\new_[12786]_ );
  assign \new_[9452]_  = ~\new_[10987]_  & (~\new_[5430]_  | ~\new_[12786]_ );
  assign \new_[9453]_  = ~\new_[10998]_  & (~\new_[5429]_  | ~\new_[12676]_ );
  assign \new_[9454]_  = ~\new_[11312]_  & (~\new_[5297]_  | ~\new_[12577]_ );
  assign \new_[9455]_  = ~\new_[11334]_  & (~\new_[5298]_  | ~\new_[12577]_ );
  assign \new_[9456]_  = ~\new_[11359]_  & (~\new_[4906]_  | ~\new_[12577]_ );
  assign \new_[9457]_  = ~\new_[10810]_  & (~\new_[5207]_  | ~\new_[12611]_ );
  assign \new_[9458]_  = ~\new_[10870]_  & (~\new_[5428]_  | ~\new_[12786]_ );
  assign \new_[9459]_  = ~\new_[11354]_  & (~\new_[5300]_  | ~\new_[12577]_ );
  assign \new_[9460]_  = ~\new_[11321]_  & (~\new_[5301]_  | ~\new_[12577]_ );
  assign \new_[9461]_  = ~\new_[10859]_  & (~\new_[5427]_  | ~\new_[12676]_ );
  assign \new_[9462]_  = ~\new_[11341]_  & (~\new_[4904]_  | ~\new_[12639]_ );
  assign \new_[9463]_  = ~\new_[11324]_  & (~\new_[5303]_  | ~\new_[12577]_ );
  assign \new_[9464]_  = ~\new_[11353]_  & (~\new_[5304]_  | ~\new_[12639]_ );
  assign \new_[9465]_  = ~\new_[10900]_  & (~\new_[5426]_  | ~\new_[12676]_ );
  assign \new_[9466]_  = ~\new_[11394]_  & (~\new_[5305]_  | ~\new_[12639]_ );
  assign \new_[9467]_  = ~\new_[11314]_  & (~\new_[4905]_  | ~\new_[12639]_ );
  assign \new_[9468]_  = ~\new_[11399]_  & (~\new_[5306]_  | ~\new_[12639]_ );
  assign \new_[9469]_  = ~\new_[11325]_  & (~\new_[5307]_  | ~\new_[12639]_ );
  assign \new_[9470]_  = ~\new_[11337]_  & (~\new_[5308]_  | ~\new_[12639]_ );
  assign \new_[9471]_  = ~\new_[11393]_  & (~\new_[4903]_  | ~\new_[12577]_ );
  assign \new_[9472]_  = ~\new_[11377]_  & (~\new_[5309]_  | ~\new_[12577]_ );
  assign \new_[9473]_  = ~\new_[11391]_  & (~\new_[5310]_  | ~\new_[12577]_ );
  assign \new_[9474]_  = ~\new_[11329]_  & (~\new_[5311]_  | ~\new_[12639]_ );
  assign \new_[9475]_  = ~\new_[11395]_  & (~\new_[4901]_  | ~\new_[12577]_ );
  assign \new_[9476]_  = ~\new_[11293]_  & (~\new_[5312]_  | ~\new_[12639]_ );
  assign \new_[9477]_  = ~\new_[11307]_  & (~\new_[5313]_  | ~\new_[12639]_ );
  assign \new_[9478]_  = ~\new_[11299]_  & (~\new_[5299]_  | ~\new_[12577]_ );
  assign \new_[9479]_  = ~\new_[11309]_  & (~\new_[5314]_  | ~\new_[12577]_ );
  assign \new_[9480]_  = ~\new_[11388]_  & (~\new_[5757]_  | ~\new_[12639]_ );
  assign \new_[9481]_  = ~\new_[11332]_  & (~\new_[5387]_  | ~\new_[12660]_ );
  assign \new_[9482]_  = ~\new_[11290]_  & (~\new_[5315]_  | ~\new_[12639]_ );
  assign \new_[9483]_  = ~\new_[11357]_  & (~\new_[5316]_  | ~\new_[12639]_ );
  assign \new_[9484]_  = ~\new_[11313]_  & (~\new_[5317]_  | ~\new_[12639]_ );
  assign \new_[9485]_  = ~\new_[11166]_  & (~\new_[5765]_  | ~\new_[12639]_ );
  assign \new_[9486]_  = ~\new_[11342]_  & (~\new_[5318]_  | ~\new_[12639]_ );
  assign \new_[9487]_  = ~\new_[11335]_  & (~\new_[5319]_  | ~\new_[12577]_ );
  assign \new_[9488]_  = ~\new_[11286]_  & (~\new_[5320]_  | ~\new_[12639]_ );
  assign \new_[9489]_  = ~\new_[11392]_  & (~\new_[5718]_  | ~\new_[12587]_ );
  assign \new_[9490]_  = ~\new_[11349]_  & (~\new_[5321]_  | ~\new_[12577]_ );
  assign \new_[9491]_  = ~\new_[11285]_  & (~\new_[5465]_  | ~\new_[12689]_ );
  assign \new_[9492]_  = ~\new_[11296]_  & (~\new_[5386]_  | ~\new_[12660]_ );
  assign \new_[9493]_  = ~\new_[11409]_  & (~\new_[5384]_  | ~\new_[12587]_ );
  assign \new_[9494]_  = ~\new_[10946]_  & (~\new_[5436]_  | ~\new_[12676]_ );
  assign \new_[9495]_  = ~\new_[11344]_  & (~\new_[5462]_  | ~\new_[12681]_ );
  assign \new_[9496]_  = ~\new_[11315]_  & (~\new_[5724]_  | ~\new_[12660]_ );
  assign \new_[9497]_  = ~\new_[11400]_  & (~\new_[5383]_  | ~\new_[12660]_ );
  assign \new_[9498]_  = ~\new_[11115]_  & (~\new_[5347]_  | ~\new_[12649]_ );
  assign \new_[9499]_  = ~\new_[11081]_  & (~\new_[5348]_  | ~\new_[12649]_ );
  assign \new_[9500]_  = ~\new_[11200]_  & (~\new_[5751]_  | ~\new_[12817]_ );
  assign \new_[9501]_  = ~\new_[11345]_  & (~\new_[5349]_  | ~\new_[12649]_ );
  assign \new_[9502]_  = ~\new_[11197]_  & (~\new_[5350]_  | ~\new_[12817]_ );
  assign \new_[9503]_  = ~\new_[11195]_  & (~\new_[5351]_  | ~\new_[12817]_ );
  assign \new_[9504]_  = ~\new_[11191]_  & (~\new_[5743]_  | ~\new_[12649]_ );
  assign \new_[9505]_  = ~\new_[11007]_  & (~\new_[5352]_  | ~\new_[12649]_ );
  assign \new_[9506]_  = ~\new_[11024]_  & (~\new_[5353]_  | ~\new_[12817]_ );
  assign \new_[9507]_  = ~\new_[11348]_  & (~\new_[5456]_  | ~\new_[12689]_ );
  assign \new_[9508]_  = ~\new_[11168]_  & (~\new_[5354]_  | ~\new_[12817]_ );
  assign \new_[9509]_  = ~\new_[11025]_  & (~\new_[5736]_  | ~\new_[12649]_ );
  assign \new_[9510]_  = ~\new_[11146]_  & (~\new_[5423]_  | ~\new_[12676]_ );
  assign \new_[9511]_  = ~\new_[11158]_  & (~\new_[5355]_  | ~\new_[12817]_ );
  assign \new_[9512]_  = ~\new_[10797]_  & (~\new_[5356]_  | ~\new_[12649]_ );
  assign \new_[9513]_  = ~\new_[11091]_  & (~\new_[5357]_  | ~\new_[12649]_ );
  assign \new_[9514]_  = ~\new_[11026]_  & (~\new_[5740]_  | ~\new_[12817]_ );
  assign \new_[9515]_  = ~\new_[11029]_  & (~\new_[5359]_  | ~\new_[12817]_ );
  assign \new_[9516]_  = ~\new_[11030]_  & (~\new_[5360]_  | ~\new_[12817]_ );
  assign \new_[9517]_  = ~\new_[11133]_  & (~\new_[5361]_  | ~\new_[12817]_ );
  assign \new_[9518]_  = ~\new_[11128]_  & (~\new_[5737]_  | ~\new_[12817]_ );
  assign \new_[9519]_  = ~\new_[10867]_  & (~\new_[5362]_  | ~\new_[12649]_ );
  assign \new_[9520]_  = ~\new_[11034]_  & (~\new_[5363]_  | ~\new_[12649]_ );
  assign \new_[9521]_  = ~\new_[11126]_  & (~\new_[5364]_  | ~\new_[12649]_ );
  assign \new_[9522]_  = ~\new_[10862]_  & (~\new_[5738]_  | ~\new_[12817]_ );
  assign \new_[9523]_  = ~\new_[11318]_  & (~\new_[5459]_  | ~\new_[12689]_ );
  assign \new_[9524]_  = ~\new_[11120]_  & (~\new_[5365]_  | ~\new_[12649]_ );
  assign \new_[9525]_  = ~\new_[11295]_  & (~\new_[5380]_  | ~\new_[12660]_ );
  assign \new_[9526]_  = ~\new_[11039]_  & (~\new_[5366]_  | ~\new_[12649]_ );
  assign \new_[9527]_  = ~\new_[11040]_  & (~\new_[5367]_  | ~\new_[12649]_ );
  assign \new_[9528]_  = ~\new_[11041]_  & (~\new_[5730]_  | ~\new_[12649]_ );
  assign \new_[9529]_  = ~\new_[11113]_  & (~\new_[5368]_  | ~\new_[12649]_ );
  assign \new_[9530]_  = ~\new_[11043]_  & (~\new_[5370]_  | ~\new_[12817]_ );
  assign \new_[9531]_  = ~\new_[11306]_  & (~\new_[5379]_  | ~\new_[12660]_ );
  assign \new_[9532]_  = ~\new_[11270]_  & (~\new_[5728]_  | ~\new_[12817]_ );
  assign \new_[9533]_  = ~\new_[11085]_  & (~\new_[5371]_  | ~\new_[12817]_ );
  assign \new_[9534]_  = ~\new_[11317]_  & (~\new_[5457]_  | ~\new_[12681]_ );
  assign \new_[9535]_  = ~\new_[11406]_  & (~\new_[5555]_  | ~\new_[12582]_ );
  assign \new_[9536]_  = ~\new_[10793]_  & (~\new_[5500]_  | ~\new_[12794]_ );
  assign \new_[9537]_  = ~\new_[10785]_  & (~\new_[5220]_  | ~\new_[12611]_ );
  assign \new_[9538]_  = ~\new_[11245]_  & (~\new_[5510]_  | ~\new_[12706]_ );
  assign \new_[9539]_  = ~\new_[11171]_  & (~\new_[5208]_  | ~\new_[12611]_ );
  assign \new_[9540]_  = ~\new_[11220]_  & (~\new_[5515]_  | ~\new_[12706]_ );
  assign \new_[9541]_  = ~\new_[10794]_  & (~\new_[4990]_  | ~\new_[12706]_ );
  assign \new_[9542]_  = ~\new_[10778]_  & (~\new_[5202]_  | ~\new_[12784]_ );
  assign \new_[9543]_  = ~\new_[10838]_  & (~\new_[5216]_  | ~\new_[12611]_ );
  assign \new_[9544]_  = ~\new_[10877]_  & (~\new_[5215]_  | ~\new_[12611]_ );
  assign \new_[9545]_  = ~\new_[10972]_  & (~\new_[5004]_  | ~\new_[12794]_ );
  assign \new_[9546]_  = ~\new_[11372]_  & (~\new_[5467]_  | ~\new_[12681]_ );
  assign \new_[9547]_  = ~\new_[11110]_  & (~\new_[5369]_  | ~\new_[12817]_ );
  assign \new_[9548]_  = ~\new_[10762]_  & (~\new_[5499]_  | ~\new_[12794]_ );
  assign \new_[9549]_  = ~\new_[11385]_  & (~\new_[5372]_  | ~\new_[12587]_ );
  assign \new_[9550]_  = ~\new_[11407]_  & (~\new_[5729]_  | ~\new_[12587]_ );
  assign \new_[9551]_  = ~\new_[11379]_  & (~\new_[5375]_  | ~\new_[12660]_ );
  assign \new_[9552]_  = ~\new_[11347]_  & (~\new_[5378]_  | ~\new_[12587]_ );
  assign \new_[9553]_  = ~\new_[11320]_  & (~\new_[5377]_  | ~\new_[12587]_ );
  assign \new_[9554]_  = ~\new_[11363]_  & (~\new_[5381]_  | ~\new_[12660]_ );
  assign \new_[9555]_  = ~\new_[11396]_  & (~\new_[5382]_  | ~\new_[12660]_ );
  assign \new_[9556]_  = ~\new_[11378]_  & (~\new_[5705]_  | ~\new_[12587]_ );
  assign \new_[9557]_  = ~\new_[11298]_  & (~\new_[5385]_  | ~\new_[12587]_ );
  assign \new_[9558]_  = ~\new_[11291]_  & (~\new_[5388]_  | ~\new_[12660]_ );
  assign \new_[9559]_  = ~\new_[11380]_  & (~\new_[5376]_  | ~\new_[12660]_ );
  assign \new_[9560]_  = ~\new_[11292]_  & (~\new_[5722]_  | ~\new_[12660]_ );
  assign \new_[9561]_  = ~\new_[11340]_  & (~\new_[5391]_  | ~\new_[12660]_ );
  assign \new_[9562]_  = ~\new_[11304]_  & (~\new_[5392]_  | ~\new_[12660]_ );
  assign \new_[9563]_  = ~\new_[11352]_  & (~\new_[5394]_  | ~\new_[12660]_ );
  assign \new_[9564]_  = ~\new_[11284]_  & (~\new_[5374]_  | ~\new_[12587]_ );
  assign \new_[9565]_  = ~\new_[11373]_  & (~\new_[5454]_  | ~\new_[12681]_ );
  assign \new_[9566]_  = ~\new_[11109]_  & (~\new_[5516]_  | ~\new_[12794]_ );
  assign \new_[9567]_  = ~\new_[11384]_  & (~\new_[5373]_  | ~\new_[12660]_ );
  assign \new_[9568]_  = ~\new_[11303]_  & (~\new_[5449]_  | ~\new_[12689]_ );
  assign \new_[9569]_  = ~\new_[11169]_  & (~\new_[5421]_  | ~\new_[12786]_ );
  assign \new_[9570]_  = ~\new_[11211]_  & (~\new_[5422]_  | ~\new_[12786]_ );
  assign \new_[9571]_  = ~\new_[11103]_  & (~\new_[5690]_  | ~\new_[12786]_ );
  assign \new_[9572]_  = ~\new_[11184]_  & (~\new_[5424]_  | ~\new_[12786]_ );
  assign \new_[9573]_  = ~\new_[10880]_  & (~\new_[5425]_  | ~\new_[12676]_ );
  assign \new_[9574]_  = ~\new_[10822]_  & (~\new_[5676]_  | ~\new_[12786]_ );
  assign \new_[9575]_  = ~\new_[11036]_  & (~\new_[5678]_  | ~\new_[12786]_ );
  assign \new_[9576]_  = ~\new_[10995]_  & (~\new_[5431]_  | ~\new_[12676]_ );
  assign \new_[9577]_  = ~\new_[10864]_  & (~\new_[5674]_  | ~\new_[12676]_ );
  assign \new_[9578]_  = ~\new_[10909]_  & (~\new_[5672]_  | ~\new_[12786]_ );
  assign \new_[9579]_  = ~\new_[11339]_  & (~\new_[5447]_  | ~\new_[12689]_ );
  assign \new_[9580]_  = ~\new_[10968]_  & (~\new_[5670]_  | ~\new_[12786]_ );
  assign \new_[9581]_  = ~\new_[10887]_  & (~\new_[5442]_  | ~\new_[12786]_ );
  assign \new_[9582]_  = ~\new_[11156]_  & (~\new_[5443]_  | ~\new_[12676]_ );
  assign \new_[9583]_  = ~\new_[11108]_  & (~\new_[5035]_  | ~\new_[12676]_ );
  assign \new_[9584]_  = ~\new_[11343]_  & (~\new_[4935]_  | ~\new_[12582]_ );
  assign \new_[9585]_  = ~\new_[10886]_  & (~\new_[5514]_  | ~\new_[12794]_ );
  assign \new_[9586]_  = ~\new_[11362]_  & (~\new_[5460]_  | ~\new_[12681]_ );
  assign \new_[9587]_  = ~\new_[11225]_  & (~\new_[5205]_  | ~\new_[12784]_ );
  assign \new_[9588]_  = ~\new_[10853]_  & (~\new_[5512]_  | ~\new_[12706]_ );
  assign \new_[9589]_  = ~\new_[10882]_  & (~\new_[5445]_  | ~\new_[12611]_ );
  assign \new_[9590]_  = ~\new_[11069]_  & (~\new_[5496]_  | ~\new_[12794]_ );
  assign \new_[9591]_  = ~\new_[11401]_  & (~\new_[5396]_  | ~\new_[12587]_ );
  assign \new_[9592]_  = ~\new_[11374]_  & (~\new_[5666]_  | ~\new_[12689]_ );
  assign \new_[9593]_  = ~\new_[11366]_  & (~\new_[5448]_  | ~\new_[12689]_ );
  assign \new_[9594]_  = ~\new_[11368]_  & (~\new_[5302]_  | ~\new_[12681]_ );
  assign \new_[9595]_  = ~\new_[11389]_  & (~\new_[5446]_  | ~\new_[12681]_ );
  assign \new_[9596]_  = ~\new_[11386]_  & (~\new_[5451]_  | ~\new_[12681]_ );
  assign \new_[9597]_  = ~\new_[11364]_  & (~\new_[5452]_  | ~\new_[12689]_ );
  assign \new_[9598]_  = ~\new_[11350]_  & (~\new_[5613]_  | ~\new_[12681]_ );
  assign \new_[9599]_  = ~\new_[11050]_  & (~\new_[5508]_  | ~\new_[12706]_ );
  assign \new_[9600]_  = ~\new_[11410]_  & (~\new_[5458]_  | ~\new_[12681]_ );
  assign \new_[9601]_  = ~\new_[11282]_  & (~\new_[4968]_  | ~\new_[12681]_ );
  assign \new_[9602]_  = ~\new_[11404]_  & (~\new_[5461]_  | ~\new_[12681]_ );
  assign \new_[9603]_  = ~\new_[11360]_  & (~\new_[5046]_  | ~\new_[12681]_ );
  assign \new_[9604]_  = ~\new_[11412]_  & (~\new_[5464]_  | ~\new_[12681]_ );
  assign \new_[9605]_  = ~\new_[11310]_  & (~\new_[5038]_  | ~\new_[12689]_ );
  assign \new_[9606]_  = ~\new_[11361]_  & (~\new_[5034]_  | ~\new_[12681]_ );
  assign \new_[9607]_  = ~\new_[11376]_  & (~\new_[5470]_  | ~\new_[12689]_ );
  assign \new_[9608]_  = ~\new_[11215]_  & (~\new_[5200]_  | ~\new_[12611]_ );
  assign \new_[9609]_  = ~\new_[10893]_  & (~\new_[5014]_  | ~\new_[12706]_ );
  assign \new_[9610]_  = ~\new_[10748]_  & (~\new_[5497]_  | ~\new_[12706]_ );
  assign \new_[9611]_  = ~\new_[11199]_  & (~\new_[4995]_  | ~\new_[12706]_ );
  assign \new_[9612]_  = ~\new_[10843]_  & (~\new_[5517]_  | ~\new_[12794]_ );
  assign \new_[9613]_  = ~\new_[10823]_  & (~\new_[5503]_  | ~\new_[12794]_ );
  assign \new_[9614]_  = ~\new_[11072]_  & (~\new_[5003]_  | ~\new_[12794]_ );
  assign \new_[9615]_  = ~\new_[10885]_  & (~\new_[5507]_  | ~\new_[12794]_ );
  assign \new_[9616]_  = ~\new_[11157]_  & (~\new_[4996]_  | ~\new_[12706]_ );
  assign \new_[9617]_  = ~\new_[10817]_  & (~\new_[4997]_  | ~\new_[12794]_ );
  assign \new_[9618]_  = ~\new_[11122]_  & (~\new_[5513]_  | ~\new_[12794]_ );
  assign \new_[9619]_  = ~\new_[10799]_  & (~\new_[4971]_  | ~\new_[12706]_ );
  assign \new_[9620]_  = ~\new_[10798]_  & (~\new_[5519]_  | ~\new_[12794]_ );
  assign \new_[9621]_  = ~\new_[10991]_  & (~\new_[5511]_  | ~\new_[12794]_ );
  assign \new_[9622]_  = ~\new_[11236]_  & (~\new_[5495]_  | ~\new_[12794]_ );
  assign \new_[9623]_  = ~\new_[10872]_  & (~\new_[5498]_  | ~\new_[12706]_ );
  assign \new_[9624]_  = ~\new_[11060]_  & (~\new_[5199]_  | ~\new_[12611]_ );
  assign \new_[9625]_  = ~\new_[11371]_  & (~\new_[5564]_  | ~\new_[12693]_ );
  assign \new_[9626]_  = ~\new_[11266]_  & (~\new_[4992]_  | ~\new_[12784]_ );
  assign \new_[9627]_  = ~\new_[10820]_  & (~\new_[5534]_  | ~\new_[12693]_ );
  assign \new_[9628]_  = ~\new_[11411]_  & (~\new_[5536]_  | ~\new_[12693]_ );
  assign \new_[9629]_  = ~\new_[11369]_  & (~\new_[4945]_  | ~\new_[12693]_ );
  assign \new_[9630]_  = ~\new_[11336]_  & (~\new_[5545]_  | ~\new_[12582]_ );
  assign \new_[9631]_  = ~\new_[11283]_  & (~\new_[5550]_  | ~\new_[12582]_ );
  assign \new_[9632]_  = ~\new_[11302]_  & (~\new_[5553]_  | ~\new_[12693]_ );
  assign \new_[9633]_  = ~\new_[11297]_  & (~\new_[4920]_  | ~\new_[12693]_ );
  assign \new_[9634]_  = ~\new_[11301]_  & (~\new_[5560]_  | ~\new_[12693]_ );
  assign \new_[9635]_  = ~\new_[11218]_  & (~\new_[5509]_  | ~\new_[12706]_ );
  assign \new_[9636]_  = ~\new_[11300]_  & (~\new_[5562]_  | ~\new_[12693]_ );
  assign \new_[9637]_  = ~\new_[11402]_  & (~\new_[4907]_  | ~\new_[12693]_ );
  assign \new_[9638]_  = ~\new_[11193]_  & (~\new_[5198]_  | ~\new_[12784]_ );
  assign \new_[9639]_  = ~\new_[11294]_  & (~\new_[5569]_  | ~\new_[12693]_ );
  assign \new_[9640]_  = ~\new_[11397]_  & (~\new_[5571]_  | ~\new_[12582]_ );
  assign \new_[9641]_  = ~\new_[11365]_  & (~\new_[5759]_  | ~\new_[12693]_ );
  assign \new_[9642]_  = ~\new_[11355]_  & (~\new_[5578]_  | ~\new_[12582]_ );
  assign \new_[9643]_  = (~\new_[12026]_  | ~\new_[13154]_ ) & (~\new_[13794]_  | ~\new_[13104]_ );
  assign \new_[9644]_  = ~\new_[14175]_  | ~\new_[2791]_ ;
  assign \new_[9645]_  = ~\new_[11437]_  | (~\new_[12262]_  & ~\new_[7774]_ );
  assign n10431 = ~\new_[11433]_  & ~\new_[12000]_ ;
  assign \new_[9647]_  = ~\new_[11469]_  & (~\new_[12259]_  | ~\new_[12594]_ );
  assign \new_[9648]_  = ~\new_[11470]_  & (~\new_[12498]_  | ~\new_[12679]_ );
  assign \new_[9649]_  = \new_[12084]_  ? \new_[12077]_  : \new_[8099]_ ;
  assign \new_[9650]_  = \new_[3374]_  ^ \new_[12258]_ ;
  assign \new_[9651]_  = \new_[3150]_  ^ \new_[12256]_ ;
  assign \new_[9652]_  = \new_[12876]_  ? \new_[12077]_  : \new_[8114]_ ;
  assign \new_[9653]_  = u12_re1_reg;
  assign \new_[9654]_  = \new_[12369]_  ^ \new_[12111]_ ;
  assign \new_[9655]_  = \new_[12873]_  ^ \new_[12112]_ ;
  assign \new_[9656]_  = u2_bit_clk_e_reg;
  assign n10451 = \new_[11452]_  | \new_[7807]_ ;
  assign n10446 = ~\new_[11466]_  & ~\new_[12088]_ ;
  assign n10421 = ~\new_[10807]_  & ~\new_[12088]_ ;
  assign \new_[9660]_  = ~\new_[11473]_  | ~\new_[10868]_ ;
  assign \new_[9661]_  = ~\new_[11445]_  & ~\new_[12120]_ ;
  assign \new_[9662]_  = ~n10941 | ~\new_[12870]_ ;
  assign \new_[9663]_  = ~\new_[11472]_  | ~\new_[10809]_ ;
  assign n10426 = ~\new_[10309]_ ;
  assign n10441 = ~\new_[12957]_  & ~\new_[11449]_ ;
  assign \new_[9666]_  = ~n10946 | ~\new_[12478]_ ;
  assign n10436 = ~\new_[11444]_  & ~\new_[11457]_ ;
  assign \new_[9668]_  = \new_[4631]_  ^ \new_[12121]_ ;
  assign \new_[9669]_  = \new_[7976]_  ^ \new_[12122]_ ;
  assign \new_[9670]_  = ~\new_[11450]_  & (~\new_[12485]_  | ~\new_[7977]_ );
  assign suspended_o = u2_suspended_reg;
  assign \new_[9672]_  = ~\new_[10318]_ ;
  assign \new_[9673]_  = \\u10_status_reg[0] ;
  assign \new_[9674]_  = ~\new_[10319]_ ;
  assign \new_[9675]_  = ~\new_[10320]_ ;
  assign \new_[9676]_  = ~\new_[10321]_ ;
  assign \new_[9677]_  = \\u9_status_reg[0] ;
  assign n10461 = ~\new_[12049]_  | ~\new_[10474]_ ;
  assign n10456 = ~\new_[12061]_  | ~\new_[11479]_ ;
  assign n10471 = ~\new_[12198]_  | ~\new_[11480]_ ;
  assign n10476 = ~\new_[11496]_  | ~\new_[10475]_ ;
  assign \new_[9682]_  = ~\new_[11500]_  & ~\new_[12432]_ ;
  assign \new_[9683]_  = ~\new_[11508]_  & ~\new_[12432]_ ;
  assign n10481 = ~\new_[11482]_  | ~\new_[11483]_ ;
  assign n10486 = ~\new_[11431]_  | ~\new_[12492]_ ;
  assign n10491 = ~\new_[11485]_  | ~\new_[12493]_ ;
  assign n10496 = ~\new_[11487]_  | ~\new_[11488]_ ;
  assign n10506 = ~\new_[11486]_  | ~\new_[12486]_ ;
  assign n10511 = ~\new_[11492]_  | ~\new_[12494]_ ;
  assign n10516 = ~\new_[11493]_  | ~\new_[12495]_ ;
  assign n10521 = ~\new_[11494]_  | ~\new_[12427]_ ;
  assign n10526 = ~\new_[11495]_  | ~\new_[12496]_ ;
  assign n10531 = ~\new_[11497]_  | ~\new_[12224]_ ;
  assign n10536 = ~\new_[11498]_  | ~\new_[11499]_ ;
  assign n10466 = ~\new_[11490]_  | ~\new_[11510]_ ;
  assign n10501 = ~\new_[11489]_  | ~\new_[12450]_ ;
  assign \new_[9697]_  = ~\new_[10489]_  & ~\new_[12594]_ ;
  assign \new_[9698]_  = ~\new_[11506]_  & ~\new_[12828]_ ;
  assign \new_[9699]_  = ~\new_[11507]_  & ~\new_[12828]_ ;
  assign \new_[9700]_  = ~\new_[10715]_  & ~\new_[14188]_ ;
  assign \new_[9701]_  = ~\new_[11481]_  | ~\new_[11678]_ ;
  assign \new_[9702]_  = ~\new_[11501]_  | ~\new_[11748]_ ;
  assign \new_[9703]_  = ~\new_[11502]_  | ~\new_[11716]_ ;
  assign \new_[9704]_  = ~\new_[11503]_  | ~\new_[11719]_ ;
  assign \new_[9705]_  = ~\new_[11505]_  | ~\new_[11783]_ ;
  assign \new_[9706]_  = ~\new_[11509]_  | ~\new_[11632]_ ;
  assign \new_[9707]_  = ~\new_[11504]_  | ~\new_[11207]_ ;
  assign \new_[9708]_  = ~\new_[10473]_  | ~\new_[11118]_ ;
  assign \new_[9709]_  = ~\new_[11491]_  | ~\new_[11744]_ ;
  assign \new_[9710]_  = \new_[13124]_  ^ \new_[12011]_ ;
  assign \new_[9711]_  = \new_[13158]_  ^ \new_[12012]_ ;
  assign \new_[9712]_  = \new_[13092]_  ^ \new_[12013]_ ;
  assign \new_[9713]_  = \new_[13161]_  ^ \new_[12010]_ ;
  assign \new_[9714]_  = \new_[3159]_  ? \new_[12662]_  : \new_[11706]_ ;
  assign \new_[9715]_  = \new_[3190]_  ? \new_[12871]_  : \new_[11727]_ ;
  assign \new_[9716]_  = \new_[3257]_  ? \new_[12663]_  : \new_[11673]_ ;
  assign \new_[9717]_  = \new_[3200]_  ? \new_[12733]_  : \new_[11626]_ ;
  assign \new_[9718]_  = \new_[3201]_  ? \new_[12733]_  : \new_[11749]_ ;
  assign \new_[9719]_  = \new_[3203]_  ? \new_[12662]_  : \new_[12015]_ ;
  assign \new_[9720]_  = \new_[3158]_  ? \new_[12662]_  : \new_[11696]_ ;
  assign \new_[9721]_  = \new_[3207]_  ? \new_[12662]_  : \new_[11688]_ ;
  assign \new_[9722]_  = \new_[3157]_  ? \new_[12662]_  : \new_[12101]_ ;
  assign \new_[9723]_  = \new_[3208]_  ? \new_[12662]_  : \new_[12080]_ ;
  assign \new_[9724]_  = \new_[3209]_  ? \new_[12662]_  : \new_[11641]_ ;
  assign \new_[9725]_  = \new_[3210]_  ? \new_[12733]_  : \new_[11698]_ ;
  assign \new_[9726]_  = \new_[3256]_  ? \new_[12837]_  : \new_[11705]_ ;
  assign \new_[9727]_  = \new_[3154]_  ? \new_[12578]_  : \new_[11626]_ ;
  assign \new_[9728]_  = \new_[3216]_  ? \new_[12760]_  : \new_[11706]_ ;
  assign \new_[9729]_  = \new_[3153]_  ? \new_[12760]_  : \new_[11747]_ ;
  assign \new_[9730]_  = \new_[3219]_  ? \new_[12578]_  : \new_[11890]_ ;
  assign \new_[9731]_  = \new_[3152]_  ? \new_[12578]_  : \new_[12101]_ ;
  assign \new_[9732]_  = \new_[3221]_  ? \new_[12578]_  : \new_[12080]_ ;
  assign \new_[9733]_  = \new_[3223]_  ? \new_[12578]_  : \new_[11698]_ ;
  assign \new_[9734]_  = \new_[3255]_  ? \new_[12837]_  : \new_[11722]_ ;
  assign \new_[9735]_  = \new_[3222]_  ? \new_[12578]_  : \new_[11641]_ ;
  assign \new_[9736]_  = \new_[3196]_  ? \new_[12574]_  : \new_[11722]_ ;
  assign \new_[9737]_  = \new_[3197]_  ? \new_[12574]_  : \new_[11705]_ ;
  assign \new_[9738]_  = \new_[3217]_  ? \new_[12578]_  : \new_[12015]_ ;
  assign \new_[9739]_  = \new_[3218]_  ? \new_[12760]_  : \new_[11696]_ ;
  assign \new_[9740]_  = \new_[3204]_  ? \new_[12662]_  : \new_[11747]_ ;
  assign \new_[9741]_  = \new_[3202]_  ? \new_[12574]_  : \new_[11673]_ ;
  assign \new_[9742]_  = \new_[3205]_  ? \new_[12733]_  : \new_[11890]_ ;
  assign \new_[9743]_  = \new_[3215]_  ? \new_[12578]_  : \new_[11749]_ ;
  assign \new_[9744]_  = \new_[3250]_  ? \new_[12663]_  : \new_[11727]_ ;
  assign \new_[9745]_  = \new_[3220]_  ? \new_[12760]_  : \new_[11688]_ ;
  assign \new_[9746]_  = (~\new_[12473]_  | ~\new_[12686]_ ) & (~\new_[11697]_  | ~\new_[13866]_ );
  assign \new_[9747]_  = (~\new_[12473]_  | ~\new_[5843]_ ) & (~\new_[11697]_  | ~\new_[13157]_ );
  assign \new_[9748]_  = (~\new_[12473]_  | ~\new_[5844]_ ) & (~\new_[11697]_  | ~\new_[5058]_ );
  assign \new_[9749]_  = (~\new_[12473]_  | ~\new_[5845]_ ) & (~\new_[11697]_  | ~\new_[5059]_ );
  assign \new_[9750]_  = (~\new_[11697]_  | ~\new_[13876]_ ) & (~\new_[10819]_  | ~\new_[13017]_ );
  assign \new_[9751]_  = (~\new_[12308]_  | ~\new_[5106]_ ) & (~\new_[2817]_  | ~\new_[12304]_ );
  assign \new_[9752]_  = (~\new_[12473]_  | ~\new_[5847]_ ) & (~\new_[11697]_  | ~\new_[5064]_ );
  assign \new_[9753]_  = (~\new_[12500]_  | ~\new_[5053]_ ) & (~\new_[10819]_  | ~\new_[5084]_ );
  assign \new_[9754]_  = (~\new_[12308]_  | ~\new_[5110]_ ) & (~\new_[4069]_  | ~\new_[12304]_ );
  assign \new_[9755]_  = ~\new_[10397]_ ;
  assign \new_[9756]_  = (~\new_[12308]_  | ~\new_[5111]_ ) & (~\new_[7789]_  | ~\new_[12304]_ );
  assign \new_[9757]_  = ~\new_[10398]_ ;
  assign \new_[9758]_  = (~\new_[12308]_  | ~\new_[5044]_ ) & (~\new_[7888]_  | ~\new_[12304]_ );
  assign \new_[9759]_  = (~\new_[12308]_  | ~\new_[5105]_ ) & (~\new_[7885]_  | ~\new_[12304]_ );
  assign \new_[9760]_  = ~\new_[10399]_ ;
  assign \new_[9761]_  = (~\new_[12308]_  | ~\new_[5113]_ ) & (~\new_[10819]_  | ~\new_[12993]_ );
  assign \new_[9762]_  = (~\new_[12308]_  | ~\new_[5114]_ ) & (~\new_[10819]_  | ~\new_[5088]_ );
  assign \new_[9763]_  = (~\new_[12308]_  | ~\new_[5116]_ ) & (~\new_[10819]_  | ~\new_[5090]_ );
  assign \new_[9764]_  = (~\new_[12473]_  | ~\new_[13110]_ ) & (~\new_[11697]_  | ~\new_[13130]_ );
  assign \new_[9765]_  = (~\new_[12473]_  | ~\new_[13082]_ ) & (~\new_[11697]_  | ~\new_[13129]_ );
  assign \new_[9766]_  = (~\new_[12473]_  | ~\new_[5876]_ ) & (~\new_[11697]_  | ~\new_[5070]_ );
  assign \new_[9767]_  = (~\new_[11697]_  | ~\new_[13098]_ ) & (~\new_[10819]_  | ~\new_[5716]_ );
  assign \new_[9768]_  = (~\new_[12473]_  | ~\new_[5850]_ ) & (~\new_[11697]_  | ~\new_[5071]_ );
  assign \new_[9769]_  = (~\new_[12473]_  | ~\new_[13137]_ ) & (~\new_[11697]_  | ~\new_[13181]_ );
  assign \new_[9770]_  = (~\new_[12473]_  | ~\new_[5852]_ ) & (~\new_[11697]_  | ~\new_[5073]_ );
  assign \new_[9771]_  = (~\new_[12473]_  | ~\new_[12519]_ ) & (~\new_[11697]_  | ~\new_[13873]_ );
  assign \new_[9772]_  = (~\new_[12473]_  | ~\new_[5873]_ ) & (~\new_[11697]_  | ~\new_[5074]_ );
  assign \new_[9773]_  = (~\new_[12308]_  | ~\new_[5107]_ ) & (~\new_[7886]_  | ~\new_[12304]_ );
  assign \new_[9774]_  = (~\new_[12473]_  | ~\new_[5874]_ ) & (~\new_[11697]_  | ~\new_[5048]_ );
  assign \new_[9775]_  = (~\new_[12473]_  | ~\new_[5767]_ ) & (~\new_[11697]_  | ~\new_[13108]_ );
  assign \new_[9776]_  = (~\new_[12473]_  | ~\new_[13126]_ ) & (~\new_[11697]_  | ~\new_[13088]_ );
  assign \new_[9777]_  = (~\new_[12308]_  | ~\new_[5108]_ ) & (~\new_[7887]_  | ~\new_[12304]_ );
  assign \new_[9778]_  = (~\new_[11697]_  | ~\new_[13155]_ ) & (~\new_[10819]_  | ~\new_[5082]_ );
  assign \new_[9779]_  = ~\new_[10401]_ ;
  assign \new_[9780]_  = ~\new_[10435]_ ;
  assign \new_[9781]_  = ~\new_[10434]_ ;
  assign \new_[9782]_  = \new_[10402]_ ;
  assign \new_[9783]_  = ~\new_[12655]_  | ~\new_[11209]_ ;
  assign \new_[9784]_  = \new_[10418]_ ;
  assign \new_[9785]_  = ~\new_[10629]_  & ~\new_[12828]_ ;
  assign \new_[9786]_  = ~\new_[12655]_  | ~\new_[11231]_ ;
  assign \new_[9787]_  = ~\new_[12655]_  | ~\new_[10782]_ ;
  assign \new_[9788]_  = ~\new_[12655]_  | ~\new_[10815]_ ;
  assign \new_[9789]_  = ~\new_[12655]_  | ~\new_[10854]_ ;
  assign \new_[9790]_  = ~\new_[12655]_  | ~\new_[11019]_ ;
  assign \new_[9791]_  = ~\new_[12655]_  | ~\new_[10918]_ ;
  assign \new_[9792]_  = ~\new_[12655]_  | ~\new_[11020]_ ;
  assign \new_[9793]_  = ~\new_[11439]_  & ~\new_[12432]_ ;
  assign \new_[9794]_  = ~\new_[10819]_  | ~\new_[5091]_ ;
  assign \new_[9795]_  = ~\new_[11028]_  & ~\new_[12432]_ ;
  assign \new_[9796]_  = ~\new_[11416]_  & ~\new_[12432]_ ;
  assign \new_[9797]_  = ~\new_[10819]_  | ~\new_[5092]_ ;
  assign \new_[9798]_  = ~\new_[10804]_  & ~\new_[12432]_ ;
  assign \new_[9799]_  = ~\new_[11154]_  & ~\new_[12432]_ ;
  assign \new_[9800]_  = ~\new_[12655]_  | ~\new_[11058]_ ;
  assign \new_[9801]_  = ~\new_[11106]_  & ~\new_[12432]_ ;
  assign \new_[9802]_  = ~\new_[11258]_  & ~\new_[12432]_ ;
  assign \new_[9803]_  = ~\new_[10876]_  & ~\new_[12432]_ ;
  assign \new_[9804]_  = ~\new_[10790]_  & ~\new_[12828]_ ;
  assign \new_[9805]_  = ~\new_[12653]_  | ~\new_[11165]_ ;
  assign \new_[9806]_  = ~\new_[10873]_  & ~\new_[12828]_ ;
  assign \new_[9807]_  = ~\new_[10770]_  & ~\new_[12828]_ ;
  assign \new_[9808]_  = ~\new_[11011]_  & ~\new_[12828]_ ;
  assign \new_[9809]_  = ~\new_[10915]_  & ~\new_[12828]_ ;
  assign \new_[9810]_  = ~\new_[12653]_  | ~\new_[11082]_ ;
  assign \new_[9811]_  = ~\new_[12655]_  | ~\new_[11144]_ ;
  assign \new_[9812]_  = ~\new_[12655]_  | ~\new_[10768]_ ;
  assign \new_[9813]_  = ~\new_[11532]_  | (~\new_[12727]_  & ~\new_[2793]_ );
  assign \new_[9814]_  = ~\new_[11484]_  & ~\new_[12828]_ ;
  assign \new_[9815]_  = ~\new_[12653]_  | ~\new_[11141]_ ;
  assign \new_[9816]_  = ~\new_[12653]_  | ~\new_[11240]_ ;
  assign \new_[9817]_  = ~\new_[11089]_  & ~\new_[12828]_ ;
  assign \new_[9818]_  = ~\new_[12655]_  | ~\new_[11083]_ ;
  assign \new_[9819]_  = ~\new_[10769]_  & ~\new_[12828]_ ;
  assign \new_[9820]_  = ~\new_[11139]_  & ~\new_[12828]_ ;
  assign \new_[9821]_  = ~\new_[10869]_  & ~\new_[12828]_ ;
  assign \new_[9822]_  = ~\new_[11087]_  & ~\new_[12828]_ ;
  assign \new_[9823]_  = \new_[10723]_  & \new_[12407]_ ;
  assign \new_[9824]_  = ~\new_[10718]_  | ~\new_[10764]_ ;
  assign \new_[9825]_  = ~\new_[10747]_  | ~\new_[10805]_ ;
  assign \new_[9826]_  = ~\new_[11545]_  | ~\new_[11419]_ ;
  assign \new_[9827]_  = (~\new_[2725]_  | ~\new_[12025]_ ) & (~\new_[6791]_  | ~\new_[12594]_ );
  assign \new_[9828]_  = ~\new_[11576]_  | ~\new_[10766]_ ;
  assign \new_[9829]_  = ~\new_[11546]_  | ~\new_[11420]_ ;
  assign \new_[9830]_  = ~\new_[11547]_  | ~\new_[11423]_ ;
  assign \new_[9831]_  = (~\new_[2747]_  | ~\new_[12590]_ ) & (~\new_[2725]_  | ~\new_[12589]_ );
  assign \new_[9832]_  = (~\new_[2736]_  | ~\new_[12590]_ ) & (~\new_[2716]_  | ~\new_[12589]_ );
  assign \new_[9833]_  = (~\new_[2716]_  | ~\new_[12025]_ ) & (~\new_[5856]_  | ~\new_[12594]_ );
  assign \new_[9834]_  = (~\new_[7876]_  | ~\new_[12590]_ ) & (~\new_[4080]_  | ~\new_[12594]_ );
  assign \new_[9835]_  = (~\new_[7875]_  | ~\new_[12590]_ ) & (~\new_[4081]_  | ~\new_[12594]_ );
  assign \new_[9836]_  = (~\new_[7929]_  | ~\new_[12025]_ ) & (~\new_[4072]_  | ~\new_[12595]_ );
  assign \new_[9837]_  = (~\new_[7686]_  | ~\new_[12590]_ ) & (~\new_[4084]_  | ~\new_[12595]_ );
  assign \new_[9838]_  = (~\new_[6791]_  | ~\new_[12590]_ ) & (~\new_[4083]_  | ~\new_[12595]_ );
  assign \new_[9839]_  = (~\new_[5856]_  | ~\new_[12590]_ ) & (~\new_[4086]_  | ~\new_[12595]_ );
  assign \new_[9840]_  = (~\new_[12441]_  | ~\new_[4409]_ ) & (~\new_[12590]_  | ~\new_[4688]_ );
  assign \new_[9841]_  = ~\new_[11620]_  | ~\new_[11261]_ ;
  assign \new_[9842]_  = ~\new_[11584]_  | ~\new_[10910]_ ;
  assign \new_[9843]_  = ~\new_[11446]_  | ~\new_[10829]_ ;
  assign \new_[9844]_  = ~\new_[10720]_  | ~\new_[10835]_ ;
  assign \new_[9845]_  = ~\new_[10738]_  | ~\new_[10851]_ ;
  assign \new_[9846]_  = ~\new_[10721]_  | ~\new_[10899]_ ;
  assign \new_[9847]_  = (~\new_[7790]_  | ~\new_[12590]_ ) & (~\new_[4075]_  | ~\new_[12594]_ );
  assign \new_[9848]_  = ~\new_[10722]_  | ~\new_[10883]_ ;
  assign \new_[9849]_  = ~\new_[11573]_  | ~\new_[11068]_ ;
  assign \new_[9850]_  = ~\new_[11206]_  | ~\new_[11003]_ ;
  assign \new_[9851]_  = ~\new_[11557]_  | ~\new_[11152]_ ;
  assign \new_[9852]_  = ~\new_[10927]_  | ~\new_[11237]_ ;
  assign \new_[9853]_  = ~\new_[11077]_  | ~\new_[10512]_ ;
  assign \new_[9854]_  = ~\new_[10988]_  | ~\new_[11075]_ ;
  assign \new_[9855]_  = ~\new_[10942]_  | ~\new_[10943]_ ;
  assign \new_[9856]_  = ~\new_[10717]_  | ~\new_[10767]_ ;
  assign \new_[9857]_  = ~\new_[11027]_  | ~\new_[10947]_ ;
  assign \new_[9858]_  = ~\new_[10741]_  | ~\new_[11750]_ ;
  assign \new_[9859]_  = ~\new_[11062]_  | ~\new_[10954]_ ;
  assign \new_[9860]_  = ~\new_[10919]_  | ~\new_[11151]_ ;
  assign \new_[9861]_  = ~\new_[10733]_  | ~\new_[11669]_ ;
  assign \new_[9862]_  = ~\new_[10960]_  | ~\new_[10961]_ ;
  assign \new_[9863]_  = ~\new_[10731]_  | ~\new_[11150]_ ;
  assign \new_[9864]_  = ~\new_[10742]_  | ~\new_[11684]_ ;
  assign \new_[9865]_  = ~\new_[10732]_  | ~\new_[11229]_ ;
  assign \new_[9866]_  = ~\new_[11592]_  | ~\new_[11104]_ ;
  assign \new_[9867]_  = (~\new_[7502]_  | ~\new_[12590]_ ) & (~\new_[4082]_  | ~\new_[12594]_ );
  assign \new_[9868]_  = ~\new_[11570]_  | ~\new_[11219]_ ;
  assign \new_[9869]_  = ~\new_[10727]_  | ~\new_[11724]_ ;
  assign \new_[9870]_  = ~\new_[11121]_  | ~\new_[10857]_ ;
  assign \new_[9871]_  = ~\new_[11542]_  | ~\new_[11056]_ ;
  assign \new_[9872]_  = ~\new_[11555]_  | ~\new_[11176]_ ;
  assign \new_[9873]_  = ~\new_[11562]_  | ~\new_[10813]_ ;
  assign \new_[9874]_  = ~\new_[11607]_  | ~\new_[10777]_ ;
  assign \new_[9875]_  = ~\new_[11548]_  | ~\new_[10784]_ ;
  assign \new_[9876]_  = ~\new_[11595]_  | ~\new_[11064]_ ;
  assign \new_[9877]_  = ~\new_[11544]_  | ~\new_[11090]_ ;
  assign \new_[9878]_  = ~\new_[11578]_  | ~\new_[11093]_ ;
  assign \new_[9879]_  = ~\new_[11610]_  | ~\new_[11015]_ ;
  assign \new_[9880]_  = ~\new_[10726]_  | ~\new_[11518]_ ;
  assign \new_[9881]_  = ~\new_[10716]_  | ~\new_[11124]_ ;
  assign \new_[9882]_  = ~\new_[10739]_  | ~\new_[11044]_ ;
  assign \new_[9883]_  = (~\new_[3546]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[6809]_ );
  assign \new_[9884]_  = (~\new_[3598]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[5888]_ );
  assign \new_[9885]_  = (~\new_[3599]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[4813]_ );
  assign \new_[9886]_  = (~\new_[3600]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[4720]_ );
  assign \new_[9887]_  = (~\new_[3449]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[4576]_ );
  assign \new_[9888]_  = (~\new_[3777]_  | ~\new_[12264]_ ) & (~\new_[12696]_  | ~\new_[7687]_ );
  assign \new_[9889]_  = (~\new_[3774]_  | ~\new_[12264]_ ) & (~\new_[12696]_  | ~\new_[7501]_ );
  assign \new_[9890]_  = (~\new_[3778]_  | ~\new_[12264]_ ) & (~\new_[12696]_  | ~\new_[6794]_ );
  assign \new_[9891]_  = (~\new_[3782]_  | ~\new_[12264]_ ) & (~\new_[12696]_  | ~\new_[4687]_ );
  assign \new_[9892]_  = ~\new_[11606]_  | ~\new_[11627]_ ;
  assign \new_[9893]_  = ~\new_[11612]_  | ~\new_[11680]_ ;
  assign \new_[9894]_  = ~\new_[11585]_  | ~\new_[12017]_ ;
  assign \new_[9895]_  = (~\new_[3779]_  | ~\new_[12264]_ ) & (~\new_[12696]_  | ~\new_[4816]_ );
  assign \new_[9896]_  = ~\new_[11761]_  & (~\new_[5412]_  | ~\new_[12745]_ );
  assign \new_[9897]_  = ~\new_[11913]_  & (~\new_[5023]_  | ~\new_[12748]_ );
  assign \new_[9898]_  = ~\new_[11867]_  & (~\new_[5411]_  | ~\new_[12745]_ );
  assign \new_[9899]_  = ~\new_[11809]_  & (~\new_[5697]_  | ~\new_[12711]_ );
  assign \new_[9900]_  = ~\new_[12063]_  & (~\new_[5325]_  | ~\new_[12756]_ );
  assign \new_[9901]_  = ~\new_[11762]_  & (~\new_[5488]_  | ~\new_[12748]_ );
  assign \new_[9902]_  = ~\new_[11764]_  & (~\new_[5409]_  | ~\new_[12745]_ );
  assign \new_[9903]_  = ~\new_[11777]_  & (~\new_[5487]_  | ~\new_[12748]_ );
  assign \new_[9904]_  = ~\new_[11853]_  & (~\new_[5164]_  | ~\new_[12759]_ );
  assign \new_[9905]_  = ~\new_[11765]_  & (~\new_[5024]_  | ~\new_[12748]_ );
  assign \new_[9906]_  = ~\new_[11791]_  & (~\new_[5668]_  | ~\new_[12745]_ );
  assign \new_[9907]_  = ~\new_[11871]_  & (~\new_[5006]_  | ~\new_[12759]_ );
  assign \new_[9908]_  = ~\new_[11835]_  & (~\new_[5171]_  | ~\new_[12759]_ );
  assign \new_[9909]_  = ~\new_[12102]_  & (~\new_[5407]_  | ~\new_[12745]_ );
  assign \new_[9910]_  = ~\new_[11784]_  & (~\new_[5141]_  | ~\new_[12749]_ );
  assign \new_[9911]_  = ~\new_[11980]_  & (~\new_[5485]_  | ~\new_[12790]_ );
  assign \new_[9912]_  = ~\new_[11869]_  & (~\new_[5177]_  | ~\new_[12759]_ );
  assign \new_[9913]_  = ~\new_[11638]_  & (~\new_[5540]_  | ~\new_[12742]_ );
  assign \new_[9914]_  = ~\new_[11965]_  & (~\new_[5182]_  | ~\new_[12759]_ );
  assign \new_[9915]_  = ~\new_[11769]_  & (~\new_[5406]_  | ~\new_[12745]_ );
  assign \new_[9916]_  = ~\new_[11820]_  & (~\new_[4999]_  | ~\new_[12759]_ );
  assign \new_[9917]_  = ~\new_[11663]_  & (~\new_[5708]_  | ~\new_[12745]_ );
  assign \new_[9918]_  = ~\new_[11957]_  & (~\new_[4998]_  | ~\new_[12741]_ );
  assign \new_[9919]_  = ~\new_[11785]_  & (~\new_[5188]_  | ~\new_[12759]_ );
  assign \new_[9920]_  = ~\new_[11718]_  & (~\new_[5189]_  | ~\new_[12741]_ );
  assign \new_[9921]_  = ~\new_[11832]_  & (~\new_[4942]_  | ~\new_[12741]_ );
  assign \new_[9922]_  = ~\new_[11904]_  & (~\new_[4993]_  | ~\new_[12741]_ );
  assign \new_[9923]_  = ~\new_[11961]_  & (~\new_[5482]_  | ~\new_[12748]_ );
  assign \new_[9924]_  = ~\new_[11751]_  & (~\new_[5404]_  | ~\new_[12745]_ );
  assign \new_[9925]_  = ~\new_[11931]_  & (~\new_[5238]_  | ~\new_[12851]_ );
  assign \new_[9926]_  = ~\new_[11825]_  & (~\new_[5195]_  | ~\new_[12741]_ );
  assign \new_[9927]_  = ~\new_[11987]_  & (~\new_[5196]_  | ~\new_[12741]_ );
  assign \new_[9928]_  = ~\new_[11908]_  & (~\new_[5197]_  | ~\new_[12741]_ );
  assign \new_[9929]_  = ~\new_[11983]_  & (~\new_[5026]_  | ~\new_[12790]_ );
  assign \new_[9930]_  = ~\new_[11821]_  & (~\new_[5237]_  | ~\new_[12851]_ );
  assign \new_[9931]_  = ~\new_[11781]_  & (~\new_[5481]_  | ~\new_[12748]_ );
  assign \new_[9932]_  = ~\new_[11905]_  & (~\new_[5403]_  | ~\new_[12711]_ );
  assign \new_[9933]_  = ~\new_[12014]_  & (~\new_[5544]_  | ~\new_[12742]_ );
  assign \new_[9934]_  = ~\new_[11964]_  & (~\new_[5480]_  | ~\new_[12790]_ );
  assign \new_[9935]_  = ~\new_[11926]_  & (~\new_[5559]_  | ~\new_[12749]_ );
  assign \new_[9936]_  = ~\new_[11945]_  & (~\new_[5704]_  | ~\new_[12711]_ );
  assign \new_[9937]_  = ~\new_[11816]_  & (~\new_[5558]_  | ~\new_[12749]_ );
  assign \new_[9938]_  = ~\new_[11929]_  & (~\new_[5479]_  | ~\new_[12748]_ );
  assign \new_[9939]_  = ~\new_[12036]_  & (~\new_[5557]_  | ~\new_[12769]_ );
  assign \new_[9940]_  = ~\new_[11937]_  & (~\new_[5556]_  | ~\new_[12749]_ );
  assign \new_[9941]_  = ~\new_[11794]_  & (~\new_[5140]_  | ~\new_[12749]_ );
  assign \new_[9942]_  = ~\new_[11811]_  & (~\new_[5139]_  | ~\new_[12769]_ );
  assign \new_[9943]_  = ~\new_[11801]_  & (~\new_[5032]_  | ~\new_[12749]_ );
  assign \new_[9944]_  = ~\new_[12098]_  & (~\new_[5137]_  | ~\new_[12769]_ );
  assign \new_[9945]_  = ~\new_[11976]_  & (~\new_[5400]_  | ~\new_[12711]_ );
  assign \new_[9946]_  = ~\new_[11807]_  & (~\new_[5135]_  | ~\new_[12749]_ );
  assign \new_[9947]_  = ~\new_[11946]_  & (~\new_[5000]_  | ~\new_[12759]_ );
  assign \new_[9948]_  = ~\new_[11819]_  & (~\new_[5763]_  | ~\new_[12769]_ );
  assign \new_[9949]_  = ~\new_[11874]_  & (~\new_[5180]_  | ~\new_[12759]_ );
  assign \new_[9950]_  = ~\new_[11947]_  & (~\new_[5577]_  | ~\new_[12749]_ );
  assign \new_[9951]_  = ~\new_[11812]_  & (~\new_[5576]_  | ~\new_[12769]_ );
  assign \new_[9952]_  = ~\new_[11854]_  & (~\new_[5483]_  | ~\new_[12748]_ );
  assign \new_[9953]_  = ~\new_[11850]_  & (~\new_[5191]_  | ~\new_[12759]_ );
  assign \new_[9954]_  = ~\new_[11928]_  & (~\new_[5575]_  | ~\new_[12769]_ );
  assign \new_[9955]_  = ~\new_[11844]_  & (~\new_[5234]_  | ~\new_[12866]_ );
  assign \new_[9956]_  = ~\new_[11827]_  & (~\new_[5574]_  | ~\new_[12749]_ );
  assign \new_[9957]_  = ~\new_[11828]_  & (~\new_[5399]_  | ~\new_[12711]_ );
  assign \new_[9958]_  = ~\new_[11879]_  & (~\new_[4966]_  | ~\new_[12851]_ );
  assign \new_[9959]_  = ~\new_[11788]_  & (~\new_[5183]_  | ~\new_[12741]_ );
  assign \new_[9960]_  = ~\new_[11843]_  & (~\new_[5221]_  | ~\new_[12851]_ );
  assign \new_[9961]_  = ~\new_[11773]_  & (~\new_[5223]_  | ~\new_[12866]_ );
  assign \new_[9962]_  = ~\new_[12109]_  & (~\new_[4970]_  | ~\new_[12851]_ );
  assign \new_[9963]_  = ~\new_[11796]_  & (~\new_[5224]_  | ~\new_[12851]_ );
  assign \new_[9964]_  = ~\new_[11802]_  & (~\new_[5714]_  | ~\new_[12711]_ );
  assign \new_[9965]_  = ~\new_[11967]_  & (~\new_[5225]_  | ~\new_[12866]_ );
  assign \new_[9966]_  = ~\new_[11930]_  & (~\new_[5027]_  | ~\new_[12790]_ );
  assign \new_[9967]_  = ~\new_[11971]_  & (~\new_[5226]_  | ~\new_[12851]_ );
  assign \new_[9968]_  = ~\new_[11985]_  & (~\new_[5227]_  | ~\new_[12851]_ );
  assign \new_[9969]_  = ~\new_[11818]_  & (~\new_[5228]_  | ~\new_[12866]_ );
  assign \new_[9970]_  = ~\new_[11810]_  & (~\new_[5229]_  | ~\new_[12866]_ );
  assign \new_[9971]_  = ~\new_[11793]_  & (~\new_[5230]_  | ~\new_[12851]_ );
  assign \new_[9972]_  = ~\new_[11772]_  & (~\new_[5231]_  | ~\new_[12866]_ );
  assign \new_[9973]_  = ~\new_[11881]_  & (~\new_[5232]_  | ~\new_[12851]_ );
  assign \new_[9974]_  = ~\new_[11883]_  & (~\new_[5233]_  | ~\new_[12866]_ );
  assign \new_[9975]_  = ~\new_[11860]_  & (~\new_[5689]_  | ~\new_[12745]_ );
  assign \new_[9976]_  = ~\new_[11875]_  & (~\new_[4965]_  | ~\new_[12866]_ );
  assign \new_[9977]_  = ~\new_[11846]_  & (~\new_[5235]_  | ~\new_[12866]_ );
  assign \new_[9978]_  = ~\new_[11966]_  & (~\new_[5236]_  | ~\new_[12851]_ );
  assign \new_[9979]_  = ~\new_[11872]_  & (~\new_[4961]_  | ~\new_[12851]_ );
  assign \new_[9980]_  = ~\new_[11805]_  & (~\new_[5476]_  | ~\new_[12790]_ );
  assign \new_[9981]_  = ~\new_[11826]_  & (~\new_[5239]_  | ~\new_[12851]_ );
  assign \new_[9982]_  = ~\new_[11539]_  & (~\new_[4952]_  | ~\new_[12851]_ );
  assign \new_[9983]_  = ~\new_[11838]_  & (~\new_[5240]_  | ~\new_[12866]_ );
  assign \new_[9984]_  = ~\new_[11527]_  & (~\new_[5241]_  | ~\new_[12866]_ );
  assign \new_[9985]_  = ~\new_[11849]_  & (~\new_[5242]_  | ~\new_[12866]_ );
  assign \new_[9986]_  = ~\new_[11894]_  & (~\new_[4954]_  | ~\new_[12866]_ );
  assign \new_[9987]_  = ~\new_[11988]_  & (~\new_[5244]_  | ~\new_[12866]_ );
  assign \new_[9988]_  = ~\new_[11970]_  & (~\new_[5245]_  | ~\new_[12866]_ );
  assign \new_[9989]_  = ~\new_[11911]_  & (~\new_[5397]_  | ~\new_[12745]_ );
  assign \new_[9990]_  = ~\new_[11852]_  & (~\new_[5246]_  | ~\new_[12797]_ );
  assign \new_[9991]_  = ~\new_[11981]_  & (~\new_[5247]_  | ~\new_[12797]_ );
  assign \new_[9992]_  = ~\new_[11833]_  & (~\new_[5248]_  | ~\new_[12797]_ );
  assign \new_[9993]_  = ~\new_[11804]_  & (~\new_[5249]_  | ~\new_[12797]_ );
  assign \new_[9994]_  = ~\new_[11847]_  & (~\new_[5250]_  | ~\new_[12797]_ );
  assign \new_[9995]_  = ~\new_[11790]_  & (~\new_[5251]_  | ~\new_[12797]_ );
  assign \new_[9996]_  = ~\new_[11941]_  & (~\new_[4899]_  | ~\new_[12769]_ );
  assign \new_[9997]_  = ~\new_[11848]_  & (~\new_[4900]_  | ~\new_[12797]_ );
  assign \new_[9998]_  = ~\new_[11952]_  & (~\new_[5252]_  | ~\new_[12797]_ );
  assign \new_[9999]_  = ~\new_[11855]_  & (~\new_[5253]_  | ~\new_[12797]_ );
  assign \new_[10000]_  = ~\new_[11959]_  & (~\new_[5254]_  | ~\new_[12797]_ );
  assign \new_[10001]_  = ~\new_[12076]_  & (~\new_[5255]_  | ~\new_[12797]_ );
  assign \new_[10002]_  = ~\new_[11938]_  & (~\new_[5257]_  | ~\new_[12797]_ );
  assign \new_[10003]_  = ~\new_[11939]_  & (~\new_[5258]_  | ~\new_[12797]_ );
  assign \new_[10004]_  = ~\new_[11856]_  & (~\new_[4938]_  | ~\new_[12797]_ );
  assign \new_[10005]_  = ~\new_[11932]_  & (~\new_[5259]_  | ~\new_[12797]_ );
  assign \new_[10006]_  = ~\new_[11936]_  & (~\new_[5473]_  | ~\new_[12790]_ );
  assign \new_[10007]_  = ~\new_[11526]_  & (~\new_[5260]_  | ~\new_[12797]_ );
  assign \new_[10008]_  = ~\new_[11893]_  & (~\new_[5261]_  | ~\new_[12797]_ );
  assign \new_[10009]_  = ~\new_[11958]_  & (~\new_[4937]_  | ~\new_[12797]_ );
  assign \new_[10010]_  = ~\new_[11920]_  & (~\new_[5262]_  | ~\new_[12797]_ );
  assign \new_[10011]_  = ~\new_[11910]_  & (~\new_[5263]_  | ~\new_[12797]_ );
  assign \new_[10012]_  = ~\new_[11775]_  & (~\new_[5264]_  | ~\new_[12797]_ );
  assign \new_[10013]_  = ~\new_[11533]_  & (~\new_[4936]_  | ~\new_[12797]_ );
  assign \new_[10014]_  = ~\new_[12214]_  & (~\new_[5265]_  | ~\new_[12797]_ );
  assign \new_[10015]_  = ~\new_[11863]_  & (~\new_[5691]_  | ~\new_[12745]_ );
  assign \new_[10016]_  = ~\new_[11774]_  & (~\new_[5266]_  | ~\new_[12797]_ );
  assign \new_[10017]_  = ~\new_[11878]_  & (~\new_[5267]_  | ~\new_[12797]_ );
  assign \new_[10018]_  = ~\new_[11862]_  & (~\new_[5520]_  | ~\new_[12742]_ );
  assign \new_[10019]_  = ~\new_[11870]_  & (~\new_[4929]_  | ~\new_[12797]_ );
  assign \new_[10020]_  = ~\new_[11622]_  & (~\new_[5268]_  | ~\new_[12797]_ );
  assign \new_[10021]_  = ~\new_[11859]_  & (~\new_[5269]_  | ~\new_[12797]_ );
  assign \new_[10022]_  = ~\new_[11955]_  & (~\new_[5270]_  | ~\new_[12797]_ );
  assign \new_[10023]_  = ~\new_[11771]_  & (~\new_[4921]_  | ~\new_[12797]_ );
  assign \new_[10024]_  = ~\new_[11864]_  & (~\new_[5031]_  | ~\new_[12748]_ );
  assign \new_[10025]_  = ~\new_[12184]_  & (~\new_[5419]_  | ~\new_[12711]_ );
  assign \new_[10026]_  = ~\new_[11896]_  & (~\new_[5471]_  | ~\new_[12748]_ );
  assign \new_[10027]_  = ~\new_[11900]_  & (~\new_[5418]_  | ~\new_[12711]_ );
  assign \new_[10028]_  = ~\new_[11885]_  & (~\new_[4948]_  | ~\new_[12742]_ );
  assign \new_[10029]_  = ~\new_[11768]_  & (~\new_[5417]_  | ~\new_[12711]_ );
  assign \new_[10030]_  = ~\new_[11814]_  & (~\new_[4964]_  | ~\new_[12742]_ );
  assign \new_[10031]_  = ~\new_[11940]_  & (~\new_[5414]_  | ~\new_[12711]_ );
  assign \new_[10032]_  = ~\new_[11822]_  & (~\new_[5415]_  | ~\new_[12745]_ );
  assign \new_[10033]_  = ~\new_[11888]_  & (~\new_[5531]_  | ~\new_[12742]_ );
  assign \new_[10034]_  = ~\new_[11808]_  & (~\new_[5565]_  | ~\new_[12769]_ );
  assign \new_[10035]_  = \new_[13757]_  ^ \new_[12788]_ ;
  assign \new_[10036]_  = ~\new_[11831]_  & (~\new_[5192]_  | ~\new_[12759]_ );
  assign \new_[10037]_  = ~\new_[11925]_  & (~\new_[5539]_  | ~\new_[12791]_ );
  assign \new_[10038]_  = ~\new_[11865]_  & (~\new_[5190]_  | ~\new_[12741]_ );
  assign \new_[10039]_  = ~\new_[11942]_  & (~\new_[4972]_  | ~\new_[12742]_ );
  assign \new_[10040]_  = ~\new_[11882]_  & (~\new_[5567]_  | ~\new_[12749]_ );
  assign \new_[10041]_  = \new_[13482]_  ^ \new_[12786]_ ;
  assign \new_[10042]_  = ~\new_[11907]_  & (~\new_[5522]_  | ~\new_[12791]_ );
  assign \new_[10043]_  = ~\new_[11873]_  & (~\new_[4943]_  | ~\new_[12791]_ );
  assign \new_[10044]_  = ~\new_[11948]_  & (~\new_[5528]_  | ~\new_[12791]_ );
  assign \new_[10045]_  = ~\new_[11918]_  & (~\new_[5175]_  | ~\new_[12741]_ );
  assign \new_[10046]_  = ~\new_[11891]_  & (~\new_[4973]_  | ~\new_[12791]_ );
  assign \new_[10047]_  = ~\new_[11767]_  & (~\new_[5535]_  | ~\new_[12791]_ );
  assign \new_[10048]_  = ~\new_[11824]_  & (~\new_[5222]_  | ~\new_[12866]_ );
  assign \new_[10049]_  = ~\new_[11766]_  & (~\new_[5525]_  | ~\new_[12791]_ );
  assign \new_[10050]_  = ~\new_[11770]_  & (~\new_[5322]_  | ~\new_[12756]_ );
  assign \new_[10051]_  = ~\new_[11993]_  & (~\new_[5323]_  | ~\new_[12756]_ );
  assign \new_[10052]_  = ~\new_[11924]_  & (~\new_[5758]_  | ~\new_[12756]_ );
  assign \new_[10053]_  = ~\new_[11763]_  & (~\new_[5324]_  | ~\new_[12756]_ );
  assign \new_[10054]_  = ~\new_[11995]_  & (~\new_[5326]_  | ~\new_[12756]_ );
  assign \new_[10055]_  = ~\new_[11782]_  & (~\new_[5762]_  | ~\new_[12803]_ );
  assign \new_[10056]_  = ~\new_[11806]_  & (~\new_[5327]_  | ~\new_[12756]_ );
  assign \new_[10057]_  = ~\new_[11897]_  & (~\new_[5328]_  | ~\new_[12803]_ );
  assign \new_[10058]_  = ~\new_[11758]_  & (~\new_[5329]_  | ~\new_[12803]_ );
  assign \new_[10059]_  = ~\new_[11845]_  & (~\new_[5330]_  | ~\new_[12803]_ );
  assign \new_[10060]_  = ~\new_[11887]_  & (~\new_[5331]_  | ~\new_[12803]_ );
  assign \new_[10061]_  = ~\new_[11902]_  & (~\new_[5491]_  | ~\new_[12790]_ );
  assign \new_[10062]_  = ~\new_[11974]_  & (~\new_[5332]_  | ~\new_[12803]_ );
  assign \new_[10063]_  = ~\new_[11898]_  & (~\new_[5761]_  | ~\new_[12803]_ );
  assign \new_[10064]_  = ~\new_[11892]_  & (~\new_[5334]_  | ~\new_[12756]_ );
  assign \new_[10065]_  = ~\new_[11989]_  & (~\new_[5335]_  | ~\new_[12756]_ );
  assign \new_[10066]_  = ~\new_[11921]_  & (~\new_[5754]_  | ~\new_[12756]_ );
  assign \new_[10067]_  = ~\new_[11979]_  & (~\new_[5336]_  | ~\new_[12803]_ );
  assign \new_[10068]_  = ~\new_[11977]_  & (~\new_[5337]_  | ~\new_[12756]_ );
  assign \new_[10069]_  = ~\new_[11975]_  & (~\new_[5413]_  | ~\new_[12745]_ );
  assign \new_[10070]_  = ~\new_[11836]_  & (~\new_[5338]_  | ~\new_[12803]_ );
  assign \new_[10071]_  = ~\new_[11759]_  & (~\new_[5340]_  | ~\new_[12803]_ );
  assign \new_[10072]_  = ~\new_[11817]_  & (~\new_[5341]_  | ~\new_[12756]_ );
  assign \new_[10073]_  = ~\new_[11919]_  & (~\new_[5344]_  | ~\new_[12756]_ );
  assign \new_[10074]_  = ~\new_[11917]_  & (~\new_[5345]_  | ~\new_[12803]_ );
  assign \new_[10075]_  = ~\new_[11534]_  & (~\new_[5732]_  | ~\new_[12803]_ );
  assign \new_[10076]_  = ~\new_[11949]_  & (~\new_[5346]_  | ~\new_[12803]_ );
  assign \new_[10077]_  = ~\new_[11689]_  & (~\new_[4919]_  | ~\new_[12749]_ );
  assign \new_[10078]_  = \new_[13723]_  ^ \new_[12817]_ ;
  assign \new_[10079]_  = ~\new_[11922]_  & (~\new_[5166]_  | ~\new_[12759]_ );
  assign \new_[10080]_  = ~\new_[11990]_  & (~\new_[5181]_  | ~\new_[12759]_ );
  assign \new_[10081]_  = ~\new_[11760]_  & (~\new_[5296]_  | ~\new_[12741]_ );
  assign \new_[10082]_  = ~\new_[11927]_  & (~\new_[5184]_  | ~\new_[12741]_ );
  assign \new_[10083]_  = ~\new_[11962]_  & (~\new_[5554]_  | ~\new_[12749]_ );
  assign \new_[10084]_  = ~\new_[11866]_  & (~\new_[5186]_  | ~\new_[12741]_ );
  assign n10626 = ~\new_[11514]_  | ~\new_[12174]_ ;
  assign \new_[10086]_  = ~\new_[11973]_  & (~\new_[5187]_  | ~\new_[12741]_ );
  assign \new_[10087]_  = ~\new_[11786]_  & (~\new_[4916]_  | ~\new_[12742]_ );
  assign \new_[10088]_  = ~\new_[11776]_  & (~\new_[5490]_  | ~\new_[12748]_ );
  assign \new_[10089]_  = ~\new_[11868]_  & (~\new_[5398]_  | ~\new_[12711]_ );
  assign \new_[10090]_  = ~\new_[11960]_  & (~\new_[5401]_  | ~\new_[12711]_ );
  assign \new_[10091]_  = ~\new_[11789]_  & (~\new_[5402]_  | ~\new_[12711]_ );
  assign \new_[10092]_  = ~\new_[11934]_  & (~\new_[5405]_  | ~\new_[12711]_ );
  assign \new_[10093]_  = ~\new_[11815]_  & (~\new_[5408]_  | ~\new_[12711]_ );
  assign \new_[10094]_  = \new_[13537]_  ^ \new_[12784]_ ;
  assign \new_[10095]_  = ~\new_[11969]_  & (~\new_[5410]_  | ~\new_[12711]_ );
  assign \new_[10096]_  = ~\new_[11823]_  & (~\new_[5552]_  | ~\new_[12749]_ );
  assign \new_[10097]_  = ~\new_[11991]_  & (~\new_[5416]_  | ~\new_[12745]_ );
  assign \new_[10098]_  = ~\new_[11837]_  & (~\new_[4987]_  | ~\new_[12742]_ );
  assign \new_[10099]_  = ~\new_[11861]_  & (~\new_[5549]_  | ~\new_[12749]_ );
  assign \new_[10100]_  = ~\new_[11953]_  & (~\new_[5256]_  | ~\new_[13066]_ );
  assign \new_[10101]_  = ~\new_[11944]_  & (~\new_[5570]_  | ~\new_[12769]_ );
  assign \new_[10102]_  = ~\new_[11858]_  & (~\new_[5173]_  | ~\new_[12741]_ );
  assign \new_[10103]_  = ~\new_[11906]_  & (~\new_[5194]_  | ~\new_[12741]_ );
  assign \new_[10104]_  = ~\new_[11954]_  & (~\new_[5692]_  | ~\new_[12711]_ );
  assign \new_[10105]_  = ~\new_[11797]_  & (~\new_[5420]_  | ~\new_[12745]_ );
  assign \new_[10106]_  = ~\new_[12041]_  & (~\new_[5572]_  | ~\new_[12749]_ );
  assign \new_[10107]_  = ~\new_[11840]_  & (~\new_[5185]_  | ~\new_[12759]_ );
  assign \new_[10108]_  = ~\new_[11982]_  & (~\new_[4962]_  | ~\new_[12742]_ );
  assign \new_[10109]_  = ~\new_[11880]_  & (~\new_[5472]_  | ~\new_[12748]_ );
  assign \new_[10110]_  = ~\new_[11935]_  & (~\new_[5474]_  | ~\new_[12790]_ );
  assign \new_[10111]_  = ~\new_[11884]_  & (~\new_[5030]_  | ~\new_[12790]_ );
  assign \new_[10112]_  = ~\new_[11792]_  & (~\new_[5475]_  | ~\new_[12790]_ );
  assign \new_[10113]_  = ~\new_[11842]_  & (~\new_[5477]_  | ~\new_[12748]_ );
  assign \new_[10114]_  = ~\new_[11984]_  & (~\new_[5478]_  | ~\new_[12790]_ );
  assign \new_[10115]_  = ~\new_[11903]_  & (~\new_[5012]_  | ~\new_[12790]_ );
  assign \new_[10116]_  = ~\new_[11951]_  & (~\new_[5484]_  | ~\new_[12790]_ );
  assign \new_[10117]_  = ~\new_[11916]_  & (~\new_[4951]_  | ~\new_[12797]_ );
  assign \new_[10118]_  = ~\new_[11899]_  & (~\new_[5486]_  | ~\new_[12790]_ );
  assign \new_[10119]_  = ~\new_[11830]_  & (~\new_[5343]_  | ~\new_[12803]_ );
  assign \new_[10120]_  = ~\new_[11909]_  & (~\new_[5489]_  | ~\new_[12790]_ );
  assign \new_[10121]_  = ~\new_[11829]_  & (~\new_[5342]_  | ~\new_[12803]_ );
  assign \new_[10122]_  = ~\new_[11933]_  & (~\new_[5492]_  | ~\new_[12790]_ );
  assign \new_[10123]_  = ~\new_[12078]_  & (~\new_[5568]_  | ~\new_[12769]_ );
  assign \new_[10124]_  = ~\new_[11914]_  & (~\new_[5494]_  | ~\new_[12748]_ );
  assign \new_[10125]_  = ~\new_[11895]_  & (~\new_[5546]_  | ~\new_[12791]_ );
  assign \new_[10126]_  = ~\new_[11803]_  & (~\new_[5339]_  | ~\new_[12803]_ );
  assign \new_[10127]_  = ~\new_[11798]_  & (~\new_[5752]_  | ~\new_[12756]_ );
  assign \new_[10128]_  = \new_[13791]_  ^ \new_[12794]_ ;
  assign \new_[10129]_  = ~\new_[11997]_  & (~\new_[5566]_  | ~\new_[12769]_ );
  assign \new_[10130]_  = ~\new_[11530]_  & (~\new_[5243]_  | ~\new_[12678]_ );
  assign \new_[10131]_  = ~\new_[11994]_  & (~\new_[5179]_  | ~\new_[12741]_ );
  assign \new_[10132]_  = ~\new_[11851]_  & (~\new_[4953]_  | ~\new_[12851]_ );
  assign \new_[10133]_  = ~\new_[11795]_  & (~\new_[5493]_  | ~\new_[12790]_ );
  assign \new_[10134]_  = ~\new_[11978]_  & (~\new_[5193]_  | ~\new_[12759]_ );
  assign \new_[10135]_  = ~\new_[11986]_  & (~\new_[5013]_  | ~\new_[12748]_ );
  assign \new_[10136]_  = ~\new_[11799]_  & (~\new_[4908]_  | ~\new_[12769]_ );
  assign \new_[10137]_  = ~\new_[11943]_  & (~\new_[5537]_  | ~\new_[12742]_ );
  assign \new_[10138]_  = ~\new_[11992]_  & (~\new_[5333]_  | ~\new_[12803]_ );
  assign \new_[10139]_  = ~\new_[11963]_  & (~\new_[5521]_  | ~\new_[12791]_ );
  assign \new_[10140]_  = ~\new_[11841]_  & (~\new_[5523]_  | ~\new_[12791]_ );
  assign \new_[10141]_  = ~\new_[11968]_  & (~\new_[5524]_  | ~\new_[12742]_ );
  assign \new_[10142]_  = ~\new_[11778]_  & (~\new_[5526]_  | ~\new_[12742]_ );
  assign \new_[10143]_  = ~\new_[11839]_  & (~\new_[5527]_  | ~\new_[12791]_ );
  assign \new_[10144]_  = ~\new_[11972]_  & (~\new_[5529]_  | ~\new_[12791]_ );
  assign \new_[10145]_  = ~\new_[11901]_  & (~\new_[5530]_  | ~\new_[12791]_ );
  assign \new_[10146]_  = ~\new_[11857]_  & (~\new_[5532]_  | ~\new_[12791]_ );
  assign \new_[10147]_  = ~\new_[11923]_  & (~\new_[5533]_  | ~\new_[12791]_ );
  assign \new_[10148]_  = ~\new_[11912]_  & (~\new_[5538]_  | ~\new_[12791]_ );
  assign \new_[10149]_  = ~\new_[11915]_  & (~\new_[5563]_  | ~\new_[12769]_ );
  assign \new_[10150]_  = ~\new_[11998]_  & (~\new_[5542]_  | ~\new_[12742]_ );
  assign \new_[10151]_  = ~\new_[11996]_  & (~\new_[5760]_  | ~\new_[12756]_ );
  assign \new_[10152]_  = ~\new_[11876]_  & (~\new_[5548]_  | ~\new_[12791]_ );
  assign \new_[10153]_  = ~\new_[11877]_  & (~\new_[5547]_  | ~\new_[12742]_ );
  assign \new_[10154]_  = ~\new_[11950]_  & (~\new_[5551]_  | ~\new_[12769]_ );
  assign \new_[10155]_  = ~\new_[11886]_  & (~\new_[4896]_  | ~\new_[12769]_ );
  assign \new_[10156]_  = ~\new_[11787]_  & (~\new_[4898]_  | ~\new_[12769]_ );
  assign \new_[10157]_  = ~\new_[11779]_  & (~\new_[5561]_  | ~\new_[12769]_ );
  assign \new_[10158]_  = (~\new_[13992]_  | ~\new_[13135]_ ) & (~\new_[13738]_  | ~\new_[13989]_ );
  assign \new_[10159]_  = ~\new_[12761]_  | (~\new_[13980]_  & ~\new_[13677]_ );
  assign \new_[10160]_  = (~\new_[12354]_  | ~\new_[13140]_ ) & (~\new_[13500]_  | ~\new_[13091]_ );
  assign \new_[10161]_  = (~\new_[12447]_  | ~\new_[2831]_ ) & (~\new_[14127]_  | ~\new_[13151]_ );
  assign \new_[10162]_  = ~\new_[5275]_  | ~\new_[14172]_ ;
  assign \new_[10163]_  = ~\new_[5277]_  | ~\new_[12055]_ ;
  assign \new_[10164]_  = ~\new_[5279]_  | ~\new_[14172]_ ;
  assign \new_[10165]_  = ~\new_[5280]_  | ~\new_[12055]_ ;
  assign \new_[10166]_  = ~\new_[5289]_  | ~\new_[12055]_ ;
  assign \new_[10167]_  = ~\new_[5291]_  | ~\new_[12055]_ ;
  assign \new_[10168]_  = ~\new_[5273]_  | ~\new_[14172]_ ;
  assign \new_[10169]_  = ~\new_[5375]_  | ~\new_[12026]_ ;
  assign \new_[10170]_  = ~\new_[5278]_  | ~\new_[14172]_ ;
  assign \new_[10171]_  = ~\new_[5294]_  | ~\new_[14172]_ ;
  assign \new_[10172]_  = ~\new_[5271]_  | ~\new_[14172]_ ;
  assign \new_[10173]_  = ~\new_[5378]_  | ~\new_[13968]_ ;
  assign \new_[10174]_  = ~\new_[5451]_  | ~\new_[12022]_ ;
  assign \new_[10175]_  = ~\new_[5396]_  | ~\new_[13968]_ ;
  assign \new_[10176]_  = ~\new_[5389]_  | ~\new_[12026]_ ;
  assign \new_[10177]_  = ~\new_[5227]_  | ~\new_[13978]_ ;
  assign \new_[10178]_  = ~\new_[5245]_  | ~\new_[13986]_ ;
  assign \new_[10179]_  = ~\new_[5458]_  | ~\new_[12023]_ ;
  assign \new_[10180]_  = ~\new_[4585]_  | ~\new_[12025]_ ;
  assign \new_[10181]_  = ~\new_[10769]_ ;
  assign \new_[10182]_  = ~\new_[10770]_ ;
  assign \new_[10183]_  = ~\new_[5233]_  | ~\new_[13984]_ ;
  assign \new_[10184]_  = ~\new_[5486]_  | ~\new_[14136]_ ;
  assign \new_[10185]_  = ~\new_[5372]_  | ~\new_[13968]_ ;
  assign \new_[10186]_  = ~\new_[10790]_ ;
  assign \new_[10187]_  = ~\new_[11416]_ ;
  assign \new_[10188]_  = ~\new_[10804]_ ;
  assign \new_[10189]_  = ~\new_[5387]_  | ~\new_[13968]_ ;
  assign \new_[10190]_  = ~\new_[5225]_  | ~\new_[13981]_ ;
  assign \new_[10191]_  = ~\new_[5452]_  | ~\new_[12022]_ ;
  assign \new_[10192]_  = ~\new_[5386]_  | ~\new_[12026]_ ;
  assign \new_[10193]_  = ~\new_[5462]_  | ~\new_[12022]_ ;
  assign \new_[10194]_  = ~\new_[5459]_  | ~\new_[12023]_ ;
  assign \new_[10195]_  = ~\new_[4409]_  | ~\new_[12025]_ ;
  assign \new_[10196]_  = ~\new_[5232]_  | ~\new_[13982]_ ;
  assign \new_[10197]_  = ~\new_[4952]_  | ~\new_[13983]_ ;
  assign \new_[10198]_  = ~\new_[5613]_  | ~\new_[13897]_ ;
  assign \new_[10199]_  = ~\new_[4954]_  | ~\new_[13976]_ ;
  assign \new_[10200]_  = ~\new_[5460]_  | ~\new_[12022]_ ;
  assign \new_[10201]_  = ~\new_[5391]_  | ~\new_[13968]_ ;
  assign \new_[10202]_  = ~\new_[5463]_  | ~\new_[12022]_ ;
  assign \new_[10203]_  = ~\new_[10869]_ ;
  assign \new_[10204]_  = ~\new_[5241]_  | ~\new_[13978]_ ;
  assign \new_[10205]_  = ~\new_[10873]_ ;
  assign \new_[10206]_  = ~\new_[10876]_ ;
  assign \new_[10207]_  = ~\new_[10629]_ ;
  assign \new_[10208]_  = ~\new_[5038]_  | ~\new_[12022]_ ;
  assign \new_[10209]_  = ~\new_[5464]_  | ~\new_[12023]_ ;
  assign \new_[10210]_  = ~\new_[10915]_ ;
  assign \new_[10211]_  = ~\new_[5395]_  | ~\new_[12026]_ ;
  assign \new_[10212]_  = ~\new_[4965]_  | ~\new_[13983]_ ;
  assign \new_[10213]_  = ~\new_[5446]_  | ~\new_[12023]_ ;
  assign \new_[10214]_  = ~\new_[5461]_  | ~\new_[12023]_ ;
  assign \new_[10215]_  = ~\new_[13981]_  | ~\new_[5223]_ ;
  assign \new_[10216]_  = ~\new_[5476]_  | ~\new_[14134]_ ;
  assign \new_[10217]_  = ~\new_[5230]_  | ~\new_[13986]_ ;
  assign \new_[10218]_  = ~\new_[11484]_ ;
  assign \new_[10219]_  = ~\new_[5239]_  | ~\new_[13978]_ ;
  assign \new_[10220]_  = ~\new_[5457]_  | ~\new_[12023]_ ;
  assign \new_[10221]_  = ~\new_[5469]_  | ~\new_[12023]_ ;
  assign \new_[10222]_  = ~\new_[5721]_  | ~\new_[12026]_ ;
  assign \new_[10223]_  = ~\new_[4970]_  | ~\new_[13975]_ ;
  assign \new_[10224]_  = ~\new_[5394]_  | ~\new_[13968]_ ;
  assign \new_[10225]_  = ~\new_[5393]_  | ~\new_[12026]_ ;
  assign \new_[10226]_  = ~\new_[5234]_  | ~\new_[13982]_ ;
  assign \new_[10227]_  = ~\new_[5724]_  | ~\new_[12026]_ ;
  assign \new_[10228]_  = ~\new_[5722]_  | ~\new_[13968]_ ;
  assign \new_[10229]_  = ~\new_[11028]_ ;
  assign \new_[10230]_  = ~\new_[5236]_  | ~\new_[13984]_ ;
  assign \new_[10231]_  = ~\new_[5481]_  | ~\new_[14135]_ ;
  assign \new_[10232]_  = ~\new_[5449]_  | ~\new_[13897]_ ;
  assign \new_[10233]_  = ~\new_[5484]_  | ~\new_[14136]_ ;
  assign \new_[10234]_  = ~\new_[5705]_  | ~\new_[12026]_ ;
  assign \new_[10235]_  = ~\new_[5384]_  | ~\new_[12026]_ ;
  assign \new_[10236]_  = ~\new_[5729]_  | ~\new_[13968]_ ;
  assign \new_[10237]_  = ~\new_[5385]_  | ~\new_[12026]_ ;
  assign \new_[10238]_  = ~\new_[5374]_  | ~\new_[13968]_ ;
  assign \new_[10239]_  = ~\new_[5718]_  | ~\new_[12026]_ ;
  assign \new_[10240]_  = ~\new_[11087]_ ;
  assign \new_[10241]_  = ~\new_[5381]_  | ~\new_[13968]_ ;
  assign \new_[10242]_  = ~\new_[5390]_  | ~\new_[13968]_ ;
  assign \new_[10243]_  = ~\new_[5379]_  | ~\new_[12026]_ ;
  assign \new_[10244]_  = ~\new_[5380]_  | ~\new_[13968]_ ;
  assign \new_[10245]_  = ~\new_[5392]_  | ~\new_[13968]_ ;
  assign \new_[10246]_  = ~\new_[5237]_  | ~\new_[13983]_ ;
  assign \new_[10247]_  = ~\new_[5383]_  | ~\new_[12026]_ ;
  assign \new_[10248]_  = ~\new_[11106]_ ;
  assign \new_[10249]_  = ~\new_[4953]_  | ~\new_[13976]_ ;
  assign \new_[10250]_  = ~\new_[5388]_  | ~\new_[12026]_ ;
  assign \new_[10251]_  = ~\new_[5024]_  | ~\new_[14136]_ ;
  assign \new_[10252]_  = ~\new_[5229]_  | ~\new_[13978]_ ;
  assign \new_[10253]_  = ~\new_[4966]_  | ~\new_[13975]_ ;
  assign \new_[10254]_  = ~\new_[5228]_  | ~\new_[13975]_ ;
  assign \new_[10255]_  = ~\new_[5382]_  | ~\new_[13968]_ ;
  assign \new_[10256]_  = ~\new_[5485]_  | ~\new_[14136]_ ;
  assign \new_[10257]_  = ~\new_[5222]_  | ~\new_[13975]_ ;
  assign \new_[10258]_  = ~\new_[5231]_  | ~\new_[13982]_ ;
  assign \new_[10259]_  = ~\new_[5243]_  | ~\new_[13982]_ ;
  assign \new_[10260]_  = ~\new_[11139]_ ;
  assign \new_[10261]_  = ~\new_[5244]_  | ~\new_[13987]_ ;
  assign \new_[10262]_  = ~\new_[5240]_  | ~\new_[13984]_ ;
  assign \new_[10263]_  = ~\new_[11154]_ ;
  assign \new_[10264]_  = ~\new_[5238]_  | ~\new_[13983]_ ;
  assign \new_[10265]_  = ~\new_[11011]_ ;
  assign \new_[10266]_  = ~\new_[5666]_  | ~\new_[12023]_ ;
  assign \new_[10267]_  = ~\new_[5482]_  | ~\new_[14135]_ ;
  assign \new_[10268]_  = ~\new_[5483]_  | ~\new_[14136]_ ;
  assign \new_[10269]_  = ~\new_[5448]_  | ~\new_[12023]_ ;
  assign \new_[10270]_  = ~\new_[5012]_  | ~\new_[14136]_ ;
  assign \new_[10271]_  = ~\new_[5450]_  | ~\new_[12023]_ ;
  assign \new_[10272]_  = ~\new_[5046]_  | ~\new_[12023]_ ;
  assign \new_[10273]_  = ~\new_[5477]_  | ~\new_[14134]_ ;
  assign \new_[10274]_  = ~\new_[5489]_  | ~\new_[14136]_ ;
  assign \new_[10275]_  = ~\new_[5465]_  | ~\new_[12022]_ ;
  assign \new_[10276]_  = ~\new_[5455]_  | ~\new_[12023]_ ;
  assign \new_[10277]_  = ~\new_[4968]_  | ~\new_[12022]_ ;
  assign \new_[10278]_  = ~\new_[5488]_  | ~\new_[14136]_ ;
  assign \new_[10279]_  = ~\new_[5221]_  | ~\new_[13976]_ ;
  assign \new_[10280]_  = ~\new_[5447]_  | ~\new_[12023]_ ;
  assign \new_[10281]_  = ~\new_[5302]_  | ~\new_[13897]_ ;
  assign \new_[10282]_  = ~\new_[4961]_  | ~\new_[13984]_ ;
  assign \new_[10283]_  = ~\new_[11439]_ ;
  assign \new_[10284]_  = ~\new_[5720]_  | ~\new_[12026]_ ;
  assign \new_[10285]_  = ~\new_[5235]_  | ~\new_[13975]_ ;
  assign \new_[10286]_  = ~\new_[11258]_ ;
  assign n10561 = ~\new_[12081]_  & ~\new_[12333]_ ;
  assign \new_[10288]_  = ~\new_[11089]_ ;
  assign n10541 = ~\new_[12452]_  & ~\new_[12001]_ ;
  assign \new_[10290]_  = ~\new_[7972]_  | ~\new_[7977]_  | ~\new_[12072]_  | ~\new_[7976]_ ;
  assign \new_[10291]_  = \new_[2952]_  ^ \new_[12497]_ ;
  assign \new_[10292]_  = \new_[7865]_  ^ \new_[12462]_ ;
  assign \new_[10293]_  = \new_[7857]_  ^ \new_[12463]_ ;
  assign \new_[10294]_  = (~\new_[3594]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[2738]_ );
  assign n10551 = ~\new_[12079]_  & ~\new_[12319]_ ;
  assign n10556 = ~\new_[7976]_  & ~\new_[12520]_  & ~\new_[12471]_ ;
  assign \new_[10297]_  = ~\new_[12077]_  | ~\new_[7956]_ ;
  assign \new_[10298]_  = \new_[12773]_  ^ \new_[12451]_ ;
  assign \new_[10299]_  = \new_[12366]_  ^ \new_[12474]_ ;
  assign \new_[10300]_  = \new_[12370]_  ^ \new_[12475]_ ;
  assign \new_[10301]_  = \new_[12368]_  ^ \new_[12476]_ ;
  assign \new_[10302]_  = \new_[7874]_  ^ \new_[12460]_ ;
  assign \new_[10303]_  = ~\new_[12100]_  | ~\new_[12859]_ ;
  assign n10921 = ~\new_[13160]_  & ~\new_[12089]_ ;
  assign \new_[10305]_  = ~\new_[11749]_  & ~\new_[12513]_ ;
  assign \new_[10306]_  = ~\new_[12107]_  & ~\new_[12108]_ ;
  assign \new_[10307]_  = ~n10951 | ~\new_[12100]_ ;
  assign \new_[10308]_  = ~\new_[12123]_  | ~\new_[11679]_ ;
  assign \new_[10309]_  = ~\new_[12507]_  | ~\new_[13726]_  | ~\new_[11617]_  | ~\new_[13300]_ ;
  assign \new_[10310]_  = ~\new_[8477]_  | ~\new_[12713]_  | ~\new_[12465]_ ;
  assign \new_[10311]_  = ~\new_[11628]_  & (~\new_[13347]_  | ~\new_[13076]_ );
  assign n10546 = ~\new_[12115]_  & ~\new_[12471]_ ;
  assign \new_[10313]_  = ~\new_[12090]_  | (~\new_[12594]_  & ~\new_[13141]_ );
  assign \new_[10314]_  = ~\new_[12087]_  | (~\new_[12679]_  & ~\new_[3081]_ );
  assign \new_[10315]_  = ~\new_[12077]_  & ~\new_[12670]_ ;
  assign \new_[10316]_  = \new_[12580]_  ^ \new_[12349]_ ;
  assign \new_[10317]_  = \\u11_status_reg[0] ;
  assign \new_[10318]_  = \\u6_status_reg[0] ;
  assign \new_[10319]_  = \\u3_status_reg[0] ;
  assign \new_[10320]_  = \\u4_status_reg[0] ;
  assign \new_[10321]_  = \\u7_status_reg[0] ;
  assign n10671 = \\u1_sr_reg[2] ;
  assign n10901 = ~\new_[12124]_  | ~\new_[12125]_ ;
  assign n10911 = ~\new_[12169]_  | ~\new_[12056]_ ;
  assign n10571 = ~\new_[12127]_  | ~\new_[12128]_ ;
  assign n10906 = ~\new_[12250]_  | ~\new_[12129]_ ;
  assign n10716 = ~\new_[12052]_  | ~\new_[12130]_ ;
  assign n10576 = ~\new_[12210]_  | ~\new_[12168]_ ;
  assign n10891 = ~\new_[12131]_  | ~\new_[12132]_ ;
  assign n10621 = ~\new_[12067]_  | ~\new_[12134]_ ;
  assign n10896 = ~\new_[12135]_  | ~\new_[12136]_ ;
  assign n10581 = ~\new_[12126]_  | ~\new_[12137]_ ;
  assign n10586 = ~\new_[12138]_  | ~\new_[12068]_ ;
  assign n10916 = ~\new_[12139]_  | ~\new_[12140]_ ;
  assign n10591 = ~\new_[12141]_  | ~\new_[12142]_ ;
  assign n10596 = ~\new_[12180]_  | ~\new_[12143]_ ;
  assign n10601 = ~\new_[12144]_  | ~\new_[12145]_ ;
  assign n10606 = ~\new_[12255]_  | ~\new_[12146]_ ;
  assign n10611 = ~\new_[12147]_  | ~\new_[12167]_ ;
  assign n10631 = ~\new_[12165]_  | ~\new_[12149]_ ;
  assign n10636 = ~\new_[12150]_  | ~\new_[12151]_ ;
  assign n10641 = ~\new_[12152]_  | ~\new_[12153]_ ;
  assign n10646 = ~\new_[11516]_  | ~\new_[12154]_ ;
  assign n10651 = ~\new_[12155]_  | ~\new_[12156]_ ;
  assign n10656 = ~\new_[11512]_  | ~\new_[12053]_ ;
  assign n10661 = ~\new_[12157]_  | ~\new_[11513]_ ;
  assign n10666 = ~\new_[12158]_  | ~\new_[12159]_ ;
  assign n10681 = ~\new_[12183]_  | ~\new_[12161]_ ;
  assign n10686 = ~\new_[12172]_  | ~\new_[12173]_ ;
  assign n10691 = ~\new_[12162]_  | ~\new_[12170]_ ;
  assign n10616 = ~\new_[12166]_  | ~\new_[12148]_ ;
  assign n10871 = ~\new_[12246]_  | ~\new_[12247]_ ;
  assign n10706 = ~\new_[12178]_  | ~\new_[12179]_ ;
  assign \new_[10354]_  = ~\new_[12545]_  | ~\new_[12618]_ ;
  assign \new_[10355]_  = ~\new_[11525]_  & ~\new_[12618]_ ;
  assign n10711 = ~\new_[12181]_  | ~\new_[12182]_ ;
  assign n10676 = ~\new_[12187]_  | ~\new_[12160]_ ;
  assign n10721 = ~\new_[12185]_  | ~\new_[12186]_ ;
  assign n10726 = ~\new_[12064]_  | ~\new_[12202]_ ;
  assign n10731 = ~\new_[12188]_  | ~\new_[12189]_ ;
  assign n10736 = ~\new_[12190]_  | ~\new_[12032]_ ;
  assign n10741 = ~\new_[12191]_  | ~\new_[12192]_ ;
  assign n10751 = ~\new_[12194]_  | ~\new_[12195]_ ;
  assign n10756 = ~\new_[12196]_  | ~\new_[12197]_ ;
  assign n10761 = ~\new_[12199]_  | ~\new_[12200]_ ;
  assign n10766 = ~\new_[12201]_  | ~\new_[12203]_ ;
  assign n10771 = ~\new_[12204]_  | ~\new_[12205]_ ;
  assign n10781 = ~\new_[12206]_  | ~\new_[12209]_ ;
  assign n10776 = ~\new_[12207]_  | ~\new_[12208]_ ;
  assign n10786 = ~\new_[12211]_  | ~\new_[12212]_ ;
  assign n10791 = ~\new_[12213]_  | ~\new_[12215]_ ;
  assign n10796 = ~\new_[12216]_  | ~\new_[12217]_ ;
  assign n10801 = ~\new_[12133]_  | ~\new_[12219]_ ;
  assign n10806 = ~\new_[12220]_  | ~\new_[12221]_ ;
  assign n10811 = ~\new_[12222]_  | ~\new_[12223]_ ;
  assign n10816 = ~\new_[12225]_  | ~\new_[12226]_ ;
  assign n10821 = ~\new_[12227]_  | ~\new_[12228]_ ;
  assign n10826 = ~\new_[12230]_  | ~\new_[12054]_ ;
  assign n10831 = ~\new_[12231]_  | ~\new_[12232]_ ;
  assign n10836 = ~\new_[12233]_  | ~\new_[12234]_ ;
  assign n10841 = ~\new_[12235]_  | ~\new_[12236]_ ;
  assign n10846 = ~\new_[12237]_  | ~\new_[12238]_ ;
  assign n10851 = ~\new_[12239]_  | ~\new_[12229]_ ;
  assign n10856 = ~\new_[12240]_  | ~\new_[12241]_ ;
  assign n10861 = ~\new_[12242]_  | ~\new_[12243]_ ;
  assign n10866 = ~\new_[12244]_  | ~\new_[12245]_ ;
  assign n10876 = ~\new_[12248]_  | ~\new_[12176]_ ;
  assign n10881 = ~\new_[12249]_  | ~\new_[12071]_ ;
  assign n10886 = ~\new_[12251]_  | ~\new_[12252]_ ;
  assign \new_[10390]_  = ~\new_[13726]_  | ~\new_[13796]_  | ~\new_[11597]_  | ~\new_[13455]_ ;
  assign n10696 = ~\new_[11515]_  | ~\new_[12163]_ ;
  assign n10746 = ~\new_[12047]_  | ~\new_[12193]_ ;
  assign n10701 = ~\new_[11517]_  | ~\new_[12164]_ ;
  assign \new_[10394]_  = ~\new_[12907]_  | ~\new_[12116]_  | ~\new_[12975]_ ;
  assign \new_[10395]_  = \new_[4641]_  ^ \new_[12343]_ ;
  assign \new_[10396]_  = \new_[4689]_  ^ \new_[12350]_ ;
  assign \new_[10397]_  = (~\new_[12500]_  | ~\new_[5054]_ ) & (~\new_[10819]_  | ~\new_[5085]_ );
  assign \new_[10398]_  = (~\new_[12500]_  | ~\new_[4894]_ ) & (~\new_[10819]_  | ~\new_[13085]_ );
  assign \new_[10399]_  = (~\new_[10819]_  | ~\new_[5086]_ ) & (~\new_[4068]_  | ~\new_[12509]_ );
  assign n10566 = ~\new_[11454]_ ;
  assign \new_[10401]_  = (~\new_[12500]_  | ~\new_[5051]_ ) & (~\new_[10819]_  | ~\new_[5081]_ );
  assign \new_[10402]_  = ~\new_[11456]_ ;
  assign \new_[10403]_  = ~\new_[7791]_  | ~\new_[12018]_ ;
  assign \new_[10404]_  = ~\new_[7881]_  | ~\new_[12018]_ ;
  assign \new_[10405]_  = ~\new_[2783]_  | ~\new_[12018]_ ;
  assign \new_[10406]_  = ~\new_[7883]_  | ~\new_[12018]_ ;
  assign \new_[10407]_  = ~\new_[12308]_  | ~\new_[5112]_ ;
  assign \new_[10408]_  = ~\new_[2818]_  | ~\new_[12018]_ ;
  assign \new_[10409]_  = ~\new_[7892]_  | ~\new_[12018]_ ;
  assign \new_[10410]_  = ~\new_[12500]_  | ~\new_[5050]_ ;
  assign \new_[10411]_  = ~\new_[2784]_  | ~\new_[12018]_ ;
  assign \new_[10412]_  = ~\new_[2819]_  | ~\new_[12018]_ ;
  assign \new_[10413]_  = ~\new_[12018]_  | ~\new_[7930]_ ;
  assign \new_[10414]_  = ~\new_[12500]_  | ~\new_[5052]_ ;
  assign \new_[10415]_  = ~\new_[12500]_  | ~\new_[5688]_ ;
  assign \new_[10416]_  = ~\new_[7882]_  | ~\new_[12018]_ ;
  assign \new_[10417]_  = \new_[11597]_  | \new_[13726]_ ;
  assign \new_[10418]_  = ~\new_[11467]_ ;
  assign \new_[10419]_  = ~\new_[11890]_  & ~\new_[12513]_ ;
  assign \new_[10420]_  = ~\new_[12101]_  & ~\new_[12513]_ ;
  assign \new_[10421]_  = ~\new_[12080]_  & ~\new_[12513]_ ;
  assign \new_[10422]_  = ~\new_[11727]_  & ~\new_[12432]_ ;
  assign \new_[10423]_  = ~\new_[11722]_  & ~\new_[12432]_ ;
  assign \new_[10424]_  = ~\new_[11705]_  & ~\new_[12432]_ ;
  assign \new_[10425]_  = ~\new_[11673]_  & ~\new_[12432]_ ;
  assign \new_[10426]_  = ~\new_[11641]_  & ~\new_[12513]_ ;
  assign \new_[10427]_  = ~\new_[11698]_  & ~\new_[12513]_ ;
  assign \new_[10428]_  = ~\new_[11688]_  & ~\new_[12513]_ ;
  assign \new_[10429]_  = ~\new_[11706]_  & ~\new_[12513]_ ;
  assign \new_[10430]_  = ~\new_[12015]_  & ~\new_[12513]_ ;
  assign \new_[10431]_  = ~\new_[11747]_  & ~\new_[12513]_ ;
  assign \new_[10432]_  = ~\new_[11696]_  & ~\new_[12513]_ ;
  assign \new_[10433]_  = ~\new_[11626]_  & ~\new_[12513]_ ;
  assign \new_[10434]_  = \new_[11583]_  & \new_[12408]_ ;
  assign \new_[10435]_  = \new_[11623]_  & \new_[12266]_ ;
  assign \new_[10436]_  = ~\new_[12535]_  & ~\new_[12618]_ ;
  assign \new_[10437]_  = (~\new_[12946]_  | ~\new_[12341]_ ) & (~\new_[13677]_  | ~\new_[2791]_ );
  assign \new_[10438]_  = (~\new_[12887]_  | ~\new_[12396]_ ) & (~\new_[13425]_  | ~\new_[2793]_ );
  assign \new_[10439]_  = (~\new_[4077]_  | ~\new_[12594]_ ) & (~\new_[3763]_  | ~\new_[12380]_ );
  assign \new_[10440]_  = (~\new_[4078]_  | ~\new_[12594]_ ) & (~\new_[3186]_  | ~\new_[12380]_ );
  assign \new_[10441]_  = (~\new_[4074]_  | ~\new_[12594]_ ) & (~\new_[2922]_  | ~\new_[12380]_ );
  assign \new_[10442]_  = (~\new_[4079]_  | ~\new_[12594]_ ) & (~\new_[2785]_  | ~\new_[12380]_ );
  assign \new_[10443]_  = (~\new_[4585]_  | ~\new_[12441]_ ) & (~\new_[4817]_  | ~\new_[12380]_ );
  assign \new_[10444]_  = ~\new_[11725]_  & (~\new_[12982]_  | ~\new_[13524]_ );
  assign \new_[10445]_  = ~\new_[11642]_  & (~\new_[13644]_  | ~\new_[13011]_ );
  assign \new_[10446]_  = (~\new_[3773]_  | ~\new_[12264]_ ) & (~\new_[12696]_  | ~\new_[5855]_ );
  assign \new_[10447]_  = ~\new_[11645]_  & (~\new_[13371]_  | ~\new_[13011]_ );
  assign \new_[10448]_  = ~\new_[11674]_  & (~\new_[13465]_  | ~\new_[13076]_ );
  assign \new_[10449]_  = ~\new_[11649]_  & (~\new_[13394]_  | ~\new_[13011]_ );
  assign \new_[10450]_  = ~\new_[11650]_  & (~\new_[13753]_  | ~\new_[13076]_ );
  assign \new_[10451]_  = ~\new_[11535]_  & (~\new_[13829]_  | ~\new_[13076]_ );
  assign \new_[10452]_  = (~\new_[3784]_  | ~\new_[12264]_ ) & (~\new_[12696]_  | ~\new_[3764]_ );
  assign \new_[10453]_  = ~\new_[11653]_  & (~\new_[13319]_  | ~\new_[13011]_ );
  assign \new_[10454]_  = ~\new_[11656]_  & (~\new_[13253]_  | ~\new_[13076]_ );
  assign \new_[10455]_  = ~\new_[11591]_  | ~\new_[11733]_ ;
  assign \new_[10456]_  = ~\new_[11559]_  | ~\new_[11662]_ ;
  assign \new_[10457]_  = ~\new_[11594]_  | ~\new_[11665]_ ;
  assign \new_[10458]_  = ~\new_[11560]_  | ~\new_[11666]_ ;
  assign \new_[10459]_  = (~\new_[3766]_  | ~\new_[12264]_ ) & (~\new_[12696]_  | ~\new_[3184]_ );
  assign \new_[10460]_  = (~\new_[3787]_  | ~\new_[12264]_ ) & (~\new_[12696]_  | ~\new_[2923]_ );
  assign \new_[10461]_  = (~\new_[3657]_  | ~\new_[12264]_ ) & (~\new_[12696]_  | ~\new_[2789]_ );
  assign \new_[10462]_  = (~\new_[3588]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[7879]_ );
  assign \new_[10463]_  = (~\new_[3589]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[3672]_ );
  assign \new_[10464]_  = (~\new_[3590]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[3185]_ );
  assign \new_[10465]_  = (~\new_[3785]_  | ~\new_[12264]_ ) & (~\new_[12696]_  | ~\new_[2737]_ );
  assign \new_[10466]_  = (~\new_[3591]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[2924]_ );
  assign \new_[10467]_  = (~\new_[3592]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[2787]_ );
  assign \new_[10468]_  = (~\new_[3593]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[2749]_ );
  assign \new_[10469]_  = (~\new_[3786]_  | ~\new_[12264]_ ) & (~\new_[12696]_  | ~\new_[2748]_ );
  assign \new_[10470]_  = (~\new_[3595]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[7926]_ );
  assign \new_[10471]_  = (~\new_[3596]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[7688]_ );
  assign \new_[10472]_  = (~\new_[3597]_  | ~\new_[12399]_ ) & (~\new_[12667]_  | ~\new_[7503]_ );
  assign \new_[10473]_  = (~\new_[12667]_  | ~\new_[4410]_ ) & (~\new_[12586]_  | ~\new_[4720]_ );
  assign \new_[10474]_  = (~\new_[13654]_  | ~\new_[13001]_ ) & (~\new_[13233]_  | ~\new_[13011]_ );
  assign \new_[10475]_  = (~\new_[13760]_  | ~\new_[13001]_ ) & (~\new_[13443]_  | ~\new_[13011]_ );
  assign \new_[10476]_  = ~\new_[13882]_  | ~\new_[5646]_ ;
  assign \new_[10477]_  = ~\new_[12338]_  & (~\new_[5147]_  | ~\new_[12818]_ );
  assign \new_[10478]_  = ~\new_[12302]_  & (~\new_[5157]_  | ~\new_[12818]_ );
  assign \new_[10479]_  = ~\new_[12457]_  & (~\new_[5007]_  | ~\new_[12818]_ );
  assign \new_[10480]_  = ~\new_[12303]_  & (~\new_[5142]_  | ~\new_[12818]_ );
  assign \new_[10481]_  = ~\new_[12328]_  & (~\new_[5165]_  | ~\new_[12818]_ );
  assign \new_[10482]_  = ~\new_[12367]_  & (~\new_[5017]_  | ~\new_[12818]_ );
  assign \new_[10483]_  = ~\new_[12310]_  & (~\new_[5011]_  | ~\new_[12818]_ );
  assign \new_[10484]_  = ~\new_[12311]_  & (~\new_[5161]_  | ~\new_[12818]_ );
  assign \new_[10485]_  = ~\new_[12336]_  & (~\new_[5160]_  | ~\new_[12818]_ );
  assign \new_[10486]_  = ~\new_[12324]_  & (~\new_[5010]_  | ~\new_[12818]_ );
  assign \new_[10487]_  = ~\new_[12397]_  | ~\new_[2756]_ ;
  assign \new_[10488]_  = ~\new_[12332]_  & (~\new_[5178]_  | ~\new_[12818]_ );
  assign \new_[10489]_  = \new_[3374]_  ^ \new_[12654]_ ;
  assign \new_[10490]_  = ~\new_[12314]_  & (~\new_[5158]_  | ~\new_[12818]_ );
  assign \new_[10491]_  = ~\new_[12261]_  & (~\new_[5163]_  | ~\new_[12818]_ );
  assign \new_[10492]_  = ~\new_[12472]_  & (~\new_[5015]_  | ~\new_[12818]_ );
  assign \new_[10493]_  = ~\new_[12316]_  & (~\new_[5155]_  | ~\new_[12818]_ );
  assign \new_[10494]_  = ~\new_[12321]_  & (~\new_[5153]_  | ~\new_[12818]_ );
  assign \new_[10495]_  = ~\new_[5576]_  | ~\new_[12352]_ ;
  assign \new_[10496]_  = ~\new_[12391]_  & ~\new_[13008]_ ;
  assign \new_[10497]_  = ~\new_[12326]_  & (~\new_[5005]_  | ~\new_[12818]_ );
  assign \new_[10498]_  = ~\new_[5533]_  | ~\new_[13992]_ ;
  assign \new_[10499]_  = ~\new_[12323]_  & (~\new_[5176]_  | ~\new_[12818]_ );
  assign \new_[10500]_  = ~\new_[12331]_  & (~\new_[5169]_  | ~\new_[12818]_ );
  assign \new_[10501]_  = ~\new_[12317]_  & (~\new_[5002]_  | ~\new_[12818]_ );
  assign \new_[10502]_  = ~\new_[12327]_  & (~\new_[5001]_  | ~\new_[12818]_ );
  assign \new_[10503]_  = ~\new_[12305]_  & (~\new_[5174]_  | ~\new_[12818]_ );
  assign \new_[10504]_  = ~\new_[12312]_  & (~\new_[5168]_  | ~\new_[12818]_ );
  assign \new_[10505]_  = ~\new_[12470]_  & (~\new_[5167]_  | ~\new_[12818]_ );
  assign \new_[10506]_  = ~\new_[12373]_  & (~\new_[5172]_  | ~\new_[12818]_ );
  assign \new_[10507]_  = ~\new_[12306]_  & (~\new_[5018]_  | ~\new_[12818]_ );
  assign \new_[10508]_  = ~\new_[12334]_  & (~\new_[5170]_  | ~\new_[12818]_ );
  assign \new_[10509]_  = ~\new_[12320]_  & (~\new_[12959]_  | ~\new_[4633]_ );
  assign \new_[10510]_  = ~\new_[5493]_  | ~\new_[14135]_ ;
  assign \new_[10511]_  = ~\new_[12424]_  & (~\new_[5150]_  | ~\new_[12818]_ );
  assign \new_[10512]_  = ~\new_[14152]_  | ~\new_[5687]_ ;
  assign \new_[10513]_  = ~\new_[12335]_  & (~\new_[5149]_  | ~\new_[12818]_ );
  assign \new_[10514]_  = ~\new_[12395]_  & ~\new_[13060]_ ;
  assign \new_[10515]_  = ~\new_[12339]_  & (~\new_[5151]_  | ~\new_[12818]_ );
  assign \new_[10516]_  = ~\new_[12260]_  & (~\new_[5146]_  | ~\new_[12818]_ );
  assign \new_[10517]_  = ~\new_[12351]_  & (~\new_[5144]_  | ~\new_[12818]_ );
  assign \new_[10518]_  = ~\new_[14152]_  | ~\new_[5600]_ ;
  assign \new_[10519]_  = \new_[5653]_  ? \new_[12601]_  : \new_[13094]_ ;
  assign \new_[10520]_  = \new_[4872]_  ? \new_[12601]_  : \new_[13087]_ ;
  assign \new_[10521]_  = \new_[5652]_  ? \new_[12601]_  : \new_[13106]_ ;
  assign \new_[10522]_  = \new_[5651]_  ? \new_[13009]_  : \new_[13128]_ ;
  assign \new_[10523]_  = \new_[5755]_  ? \new_[12601]_  : \new_[13128]_ ;
  assign \new_[10524]_  = \new_[5725]_  ? \new_[12601]_  : \new_[13183]_ ;
  assign \new_[10525]_  = \new_[5650]_  ? \new_[12601]_  : \new_[13167]_ ;
  assign \new_[10526]_  = \new_[5649]_  ? \new_[12601]_  : \new_[13164]_ ;
  assign \new_[10527]_  = \new_[5766]_  ? \new_[12601]_  : \new_[13189]_ ;
  assign \new_[10528]_  = \new_[5647]_  ? \new_[12601]_  : \new_[13136]_ ;
  assign \new_[10529]_  = \new_[4864]_  ? \new_[12601]_  : \new_[13182]_ ;
  assign \new_[10530]_  = \new_[4912]_  ? \new_[12601]_  : \new_[13133]_ ;
  assign \new_[10531]_  = \new_[5645]_  ? \new_[12606]_  : \new_[13136]_ ;
  assign \new_[10532]_  = \new_[5703]_  ? \new_[12601]_  : \new_[13117]_ ;
  assign \new_[10533]_  = \new_[4874]_  ? \new_[13009]_  : \new_[13177]_ ;
  assign \new_[10534]_  = \new_[5642]_  ? \new_[12601]_  : \new_[13122]_ ;
  assign \new_[10535]_  = \new_[4863]_  ? \new_[12601]_  : \new_[13090]_ ;
  assign \new_[10536]_  = \new_[4895]_  ? \new_[12606]_  : \new_[13182]_ ;
  assign \new_[10537]_  = \new_[4862]_  ? \new_[12601]_  : \new_[13111]_ ;
  assign \new_[10538]_  = \new_[5857]_  ? \new_[12606]_  : \new_[13187]_ ;
  assign \new_[10539]_  = \new_[4859]_  ? \new_[12606]_  : \new_[13090]_ ;
  assign \new_[10540]_  = \new_[4858]_  ? \new_[12606]_  : \new_[13111]_ ;
  assign \new_[10541]_  = \new_[5640]_  ? \new_[12606]_  : \new_[13162]_ ;
  assign \new_[10542]_  = \new_[5777]_  ? \new_[12606]_  : \new_[13166]_ ;
  assign \new_[10543]_  = \new_[5626]_  ? \new_[12953]_  : \new_[13111]_ ;
  assign \new_[10544]_  = \new_[4860]_  ? \new_[12606]_  : \new_[13133]_ ;
  assign \new_[10545]_  = \new_[5579]_  ? \new_[12521]_  : \new_[13166]_ ;
  assign \new_[10546]_  = \new_[5580]_  ? \new_[12521]_  : \new_[13162]_ ;
  assign \new_[10547]_  = \new_[5581]_  ? \new_[12521]_  : \new_[13111]_ ;
  assign \new_[10548]_  = \new_[5753]_  ? \new_[12521]_  : \new_[13090]_ ;
  assign \new_[10549]_  = \new_[4818]_  ? \new_[12521]_  : \new_[13122]_ ;
  assign \new_[10550]_  = \new_[4819]_  ? \new_[12521]_  : \new_[13187]_ ;
  assign \new_[10551]_  = \new_[5582]_  ? \new_[12521]_  : \new_[13133]_ ;
  assign \new_[10552]_  = \new_[4850]_  ? \new_[12616]_  : \new_[13185]_ ;
  assign \new_[10553]_  = \new_[4820]_  ? \new_[12521]_  : \new_[13185]_ ;
  assign \new_[10554]_  = \new_[5593]_  ? \new_[12521]_  : \new_[13172]_ ;
  assign \new_[10555]_  = \new_[5735]_  ? \new_[12899]_  : \new_[13182]_ ;
  assign \new_[10556]_  = \new_[4994]_  ? \new_[12953]_  : \new_[13090]_ ;
  assign \new_[10557]_  = \new_[5583]_  ? \new_[12521]_  : \new_[13173]_ ;
  assign \new_[10558]_  = \new_[4821]_  ? \new_[12521]_  : \new_[13136]_ ;
  assign \new_[10559]_  = \new_[5584]_  ? \new_[12521]_  : \new_[13189]_ ;
  assign \new_[10560]_  = \new_[5748]_  ? \new_[12521]_  : \new_[13164]_ ;
  assign \new_[10561]_  = \new_[5585]_  ? \new_[12521]_  : \new_[13167]_ ;
  assign \new_[10562]_  = \new_[4822]_  ? \new_[12521]_  : \new_[13128]_ ;
  assign \new_[10563]_  = \new_[5733]_  ? \new_[12521]_  : \new_[13106]_ ;
  assign \new_[10564]_  = \new_[4877]_  ? \new_[12606]_  : \new_[13172]_ ;
  assign \new_[10565]_  = \new_[4823]_  ? \new_[12521]_  : \new_[13094]_ ;
  assign \new_[10566]_  = \new_[5586]_  ? \new_[12899]_  : \new_[13176]_ ;
  assign \new_[10567]_  = \new_[5589]_  ? \new_[12521]_  : \new_[13095]_ ;
  assign \new_[10568]_  = \new_[5587]_  ? \new_[12521]_  : \new_[13156]_ ;
  assign \new_[10569]_  = \new_[5588]_  ? \new_[12899]_  : \new_[13159]_ ;
  assign \new_[10570]_  = \new_[5591]_  ? \new_[12521]_  : \new_[13123]_ ;
  assign \new_[10571]_  = \new_[5590]_  ? \new_[12899]_  : \new_[13177]_ ;
  assign \new_[10572]_  = \new_[5726]_  ? \new_[12521]_  : \new_[13132]_ ;
  assign \new_[10573]_  = \new_[4824]_  ? \new_[12521]_  : \new_[13117]_ ;
  assign \new_[10574]_  = \new_[5592]_  ? \new_[12521]_  : \new_[13183]_ ;
  assign \new_[10575]_  = \new_[4825]_  ? \new_[12521]_  : \new_[13087]_ ;
  assign \new_[10576]_  = \new_[5719]_  ? \new_[12521]_  : \new_[13163]_ ;
  assign \new_[10577]_  = \new_[4826]_  ? \new_[12521]_  : \new_[13086]_ ;
  assign \new_[10578]_  = \new_[5594]_  ? \new_[12521]_  : \new_[13184]_ ;
  assign \new_[10579]_  = \new_[4827]_  ? \new_[12521]_  : \new_[13179]_ ;
  assign \new_[10580]_  = \new_[5693]_  ? \new_[13009]_  : \new_[13179]_ ;
  assign \new_[10581]_  = \new_[5661]_  ? \new_[12601]_  : \new_[13163]_ ;
  assign \new_[10582]_  = \new_[4870]_  ? \new_[12601]_  : \new_[13132]_ ;
  assign \new_[10583]_  = \new_[5731]_  ? \new_[12601]_  : \new_[13177]_ ;
  assign \new_[10584]_  = \new_[5664]_  ? \new_[12606]_  : \new_[13183]_ ;
  assign \new_[10585]_  = \new_[5723]_  ? \new_[12598]_  : \new_[13166]_ ;
  assign \new_[10586]_  = \new_[5595]_  ? \new_[12598]_  : \new_[13162]_ ;
  assign \new_[10587]_  = \new_[5596]_  ? \new_[12598]_  : \new_[13111]_ ;
  assign \new_[10588]_  = \new_[5717]_  ? \new_[12598]_  : \new_[13090]_ ;
  assign \new_[10589]_  = \new_[4829]_  ? \new_[12598]_  : \new_[13187]_ ;
  assign \new_[10590]_  = \new_[5597]_  ? \new_[12598]_  : \new_[13133]_ ;
  assign \new_[10591]_  = \new_[4830]_  ? \new_[12598]_  : \new_[13185]_ ;
  assign \new_[10592]_  = \new_[5715]_  ? \new_[12598]_  : \new_[13182]_ ;
  assign \new_[10593]_  = \new_[5598]_  ? \new_[12598]_  : \new_[13173]_ ;
  assign \new_[10594]_  = \new_[4831]_  ? \new_[12598]_  : \new_[13136]_ ;
  assign \new_[10595]_  = \new_[5599]_  ? \new_[12598]_  : \new_[13189]_ ;
  assign \new_[10596]_  = \new_[5702]_  ? \new_[12598]_  : \new_[13164]_ ;
  assign \new_[10597]_  = \new_[5600]_  ? \new_[12598]_  : \new_[13167]_ ;
  assign \new_[10598]_  = \new_[4832]_  ? \new_[12598]_  : \new_[13128]_ ;
  assign \new_[10599]_  = \new_[5687]_  ? \new_[12598]_  : \new_[13106]_ ;
  assign \new_[10600]_  = \new_[4833]_  ? \new_[12598]_  : \new_[13094]_ ;
  assign \new_[10601]_  = \new_[5604]_  ? \new_[12920]_  : \new_[13176]_ ;
  assign \new_[10602]_  = \new_[5009]_  ? \new_[12616]_  : \new_[13166]_ ;
  assign \new_[10603]_  = \new_[5602]_  ? \new_[12598]_  : \new_[13095]_ ;
  assign \new_[10604]_  = \new_[5695]_  ? \new_[12598]_  : \new_[13159]_ ;
  assign \new_[10605]_  = \new_[5606]_  ? \new_[12920]_  : \new_[13123]_ ;
  assign \new_[10606]_  = ~\new_[5016]_  | ~\new_[12354]_ ;
  assign \new_[10607]_  = \new_[5605]_  ? \new_[12920]_  : \new_[13177]_ ;
  assign \new_[10608]_  = \new_[5686]_  ? \new_[12598]_  : \new_[13132]_ ;
  assign \new_[10609]_  = \new_[4834]_  ? \new_[12598]_  : \new_[13117]_ ;
  assign \new_[10610]_  = \new_[5607]_  ? \new_[12598]_  : \new_[13183]_ ;
  assign \new_[10611]_  = \new_[4835]_  ? \new_[12598]_  : \new_[13087]_ ;
  assign \new_[10612]_  = \new_[4836]_  ? \new_[12598]_  : \new_[13086]_ ;
  assign \new_[10613]_  = \new_[5609]_  ? \new_[12920]_  : \new_[13184]_ ;
  assign \new_[10614]_  = \new_[4837]_  ? \new_[12598]_  : \new_[13179]_ ;
  assign \new_[10615]_  = \new_[5608]_  ? \new_[12598]_  : \new_[13172]_ ;
  assign \new_[10616]_  = \new_[5677]_  ? \new_[12598]_  : \new_[13163]_ ;
  assign \new_[10617]_  = \new_[4868]_  ? \new_[12601]_  : \new_[13159]_ ;
  assign \new_[10618]_  = \new_[4849]_  ? \new_[12616]_  : \new_[13187]_ ;
  assign \new_[10619]_  = \new_[5669]_  ? \new_[12685]_  : \new_[13166]_ ;
  assign \new_[10620]_  = \new_[5610]_  ? \new_[12902]_  : \new_[13162]_ ;
  assign \new_[10621]_  = \new_[4986]_  ? \new_[12685]_  : \new_[13090]_ ;
  assign \new_[10622]_  = \new_[4838]_  ? \new_[12685]_  : \new_[13122]_ ;
  assign \new_[10623]_  = \new_[5625]_  ? \new_[12616]_  : \new_[13162]_ ;
  assign \new_[10624]_  = \new_[5612]_  ? \new_[12685]_  : \new_[13133]_ ;
  assign \new_[10625]_  = \new_[4840]_  ? \new_[12685]_  : \new_[13185]_ ;
  assign \new_[10626]_  = \new_[5614]_  ? \new_[12685]_  : \new_[13173]_ ;
  assign \new_[10627]_  = \new_[5047]_  ? \new_[12685]_  : \new_[13106]_ ;
  assign \new_[10628]_  = \new_[5617]_  ? \new_[12685]_  : \new_[13095]_ ;
  assign \new_[10629]_  = ~\new_[12399]_  | ~\new_[4720]_ ;
  assign \new_[10630]_  = \new_[5620]_  ? \new_[12685]_  : \new_[13177]_ ;
  assign \new_[10631]_  = \new_[5028]_  ? \new_[12685]_  : \new_[13132]_ ;
  assign \new_[10632]_  = \new_[4844]_  ? \new_[12685]_  : \new_[13117]_ ;
  assign \new_[10633]_  = \new_[5623]_  ? \new_[12685]_  : \new_[13172]_ ;
  assign \new_[10634]_  = \new_[4846]_  ? \new_[12902]_  : \new_[13086]_ ;
  assign \new_[10635]_  = \new_[5624]_  ? \new_[12902]_  : \new_[13184]_ ;
  assign \new_[10636]_  = \new_[4847]_  ? \new_[12685]_  : \new_[13179]_ ;
  assign \new_[10637]_  = \new_[5603]_  ? \new_[12598]_  : \new_[13156]_ ;
  assign \new_[10638]_  = \new_[5858]_  ? \new_[12606]_  : \new_[13086]_ ;
  assign \new_[10639]_  = \new_[5029]_  ? \new_[12685]_  : \new_[13163]_ ;
  assign \new_[10640]_  = \new_[5744]_  ? \new_[12601]_  : \new_[13156]_ ;
  assign \new_[10641]_  = \new_[5660]_  ? \new_[12601]_  : \new_[13184]_ ;
  assign \new_[10642]_  = \new_[4845]_  ? \new_[12685]_  : \new_[13087]_ ;
  assign \new_[10643]_  = \new_[4848]_  ? \new_[12616]_  : \new_[13122]_ ;
  assign \new_[10644]_  = \new_[5627]_  ? \new_[12616]_  : \new_[13133]_ ;
  assign \new_[10645]_  = \new_[5008]_  ? \new_[12616]_  : \new_[13182]_ ;
  assign \new_[10646]_  = \new_[4897]_  ? \new_[12953]_  : \new_[13164]_ ;
  assign \new_[10647]_  = \new_[4852]_  ? \new_[12616]_  : \new_[13128]_ ;
  assign \new_[10648]_  = \new_[4853]_  ? \new_[12616]_  : \new_[13094]_ ;
  assign \new_[10649]_  = \new_[5634]_  ? \new_[12616]_  : \new_[13095]_ ;
  assign \new_[10650]_  = \new_[5633]_  ? \new_[12616]_  : \new_[13159]_ ;
  assign \new_[10651]_  = \new_[4854]_  ? \new_[12616]_  : \new_[13117]_ ;
  assign \new_[10652]_  = \new_[5621]_  ? \new_[12685]_  : \new_[13123]_ ;
  assign \new_[10653]_  = \new_[4967]_  ? \new_[12616]_  : \new_[13163]_ ;
  assign \new_[10654]_  = \new_[5615]_  ? \new_[12685]_  : \new_[13189]_ ;
  assign \new_[10655]_  = \new_[5622]_  ? \new_[12685]_  : \new_[13183]_ ;
  assign \new_[10656]_  = \new_[5655]_  ? \new_[12606]_  : \new_[13094]_ ;
  assign \new_[10657]_  = \new_[4857]_  ? \new_[12616]_  : \new_[13179]_ ;
  assign \new_[10658]_  = \new_[5639]_  ? \new_[12616]_  : \new_[13184]_ ;
  assign \new_[10659]_  = \new_[4828]_  ? \new_[12598]_  : \new_[13122]_ ;
  assign \new_[10660]_  = \new_[4856]_  ? \new_[12616]_  : \new_[13086]_ ;
  assign \new_[10661]_  = \new_[5033]_  ? \new_[12685]_  : \new_[13159]_ ;
  assign \new_[10662]_  = \new_[5638]_  ? \new_[12616]_  : \new_[13172]_ ;
  assign \new_[10663]_  = \new_[4855]_  ? \new_[12616]_  : \new_[13087]_ ;
  assign \new_[10664]_  = \new_[5618]_  ? \new_[12685]_  : \new_[13156]_ ;
  assign \new_[10665]_  = \new_[5637]_  ? \new_[12616]_  : \new_[13183]_ ;
  assign \new_[10666]_  = \new_[5619]_  ? \new_[12685]_  : \new_[13176]_ ;
  assign \new_[10667]_  = \new_[4843]_  ? \new_[12685]_  : \new_[13094]_ ;
  assign \new_[10668]_  = \new_[4941]_  ? \new_[12616]_  : \new_[13132]_ ;
  assign \new_[10669]_  = \new_[5635]_  ? \new_[12616]_  : \new_[13177]_ ;
  assign \new_[10670]_  = \new_[4842]_  ? \new_[12685]_  : \new_[13128]_ ;
  assign \new_[10671]_  = \new_[5636]_  ? \new_[12616]_  : \new_[13123]_ ;
  assign \new_[10672]_  = \new_[5505]_  ? \new_[12685]_  : \new_[13164]_ ;
  assign \new_[10673]_  = \new_[5616]_  ? \new_[12685]_  : \new_[13167]_ ;
  assign \new_[10674]_  = \new_[5632]_  ? \new_[12616]_  : \new_[13156]_ ;
  assign \new_[10675]_  = \new_[4963]_  ? \new_[12606]_  : \new_[13122]_ ;
  assign \new_[10676]_  = \new_[4861]_  ? \new_[12601]_  : \new_[13166]_ ;
  assign \new_[10677]_  = \new_[4913]_  ? \new_[12606]_  : \new_[13185]_ ;
  assign \new_[10678]_  = \new_[5641]_  ? \new_[12601]_  : \new_[13162]_ ;
  assign \new_[10679]_  = \new_[5643]_  ? \new_[12606]_  : \new_[13173]_ ;
  assign \new_[10680]_  = \new_[5644]_  ? \new_[12601]_  : \new_[13187]_ ;
  assign \new_[10681]_  = \new_[5727]_  ? \new_[12601]_  : \new_[13185]_ ;
  assign \new_[10682]_  = \new_[4865]_  ? \new_[12606]_  : \new_[13189]_ ;
  assign \new_[10683]_  = \new_[5646]_  ? \new_[12601]_  : \new_[13173]_ ;
  assign \new_[10684]_  = \new_[5648]_  ? \new_[12606]_  : \new_[13164]_ ;
  assign \new_[10685]_  = \new_[4866]_  ? \new_[12606]_  : \new_[13167]_ ;
  assign \new_[10686]_  = \new_[5734]_  ? \new_[12606]_  : \new_[13106]_ ;
  assign \new_[10687]_  = ~\new_[13972]_  | ~\new_[4838]_ ;
  assign \new_[10688]_  = \new_[5654]_  ? \new_[12601]_  : \new_[13176]_ ;
  assign \new_[10689]_  = \new_[4867]_  ? \new_[12601]_  : \new_[13095]_ ;
  assign \new_[10690]_  = \new_[5656]_  ? \new_[12606]_  : \new_[13176]_ ;
  assign \new_[10691]_  = \new_[4869]_  ? \new_[12601]_  : \new_[13123]_ ;
  assign \new_[10692]_  = \new_[5657]_  ? \new_[12606]_  : \new_[13095]_ ;
  assign \new_[10693]_  = \new_[4871]_  ? \new_[12606]_  : \new_[13156]_ ;
  assign \new_[10694]_  = \new_[5658]_  ? \new_[12606]_  : \new_[13159]_ ;
  assign \new_[10695]_  = \new_[4873]_  ? \new_[12601]_  : \new_[13172]_ ;
  assign \new_[10696]_  = \new_[4875]_  ? \new_[12606]_  : \new_[13123]_ ;
  assign \new_[10697]_  = \new_[5662]_  ? \new_[12601]_  : \new_[13179]_ ;
  assign \new_[10698]_  = \new_[5663]_  ? \new_[12606]_  : \new_[13132]_ ;
  assign \new_[10699]_  = \new_[5875]_  ? \new_[12606]_  : \new_[13117]_ ;
  assign \new_[10700]_  = \new_[5358]_  ? \new_[12685]_  : \new_[13182]_ ;
  assign \new_[10701]_  = \new_[5701]_  ? \new_[12606]_  : \new_[13087]_ ;
  assign \new_[10702]_  = \new_[4876]_  ? \new_[13009]_  : \new_[13163]_ ;
  assign \new_[10703]_  = \new_[4841]_  ? \new_[12685]_  : \new_[13136]_ ;
  assign \new_[10704]_  = \new_[5665]_  ? \new_[12606]_  : \new_[13184]_ ;
  assign \new_[10705]_  = \new_[5631]_  ? \new_[12616]_  : \new_[13176]_ ;
  assign \new_[10706]_  = \new_[5659]_  ? \new_[12601]_  : \new_[13086]_ ;
  assign \new_[10707]_  = \new_[4978]_  ? \new_[12616]_  : \new_[13106]_ ;
  assign \new_[10708]_  = \new_[5630]_  ? \new_[12616]_  : \new_[13167]_ ;
  assign \new_[10709]_  = \new_[4839]_  ? \new_[12685]_  : \new_[13187]_ ;
  assign \new_[10710]_  = \new_[5629]_  ? \new_[12953]_  : \new_[13189]_ ;
  assign \new_[10711]_  = \new_[5611]_  ? \new_[12902]_  : \new_[13111]_ ;
  assign \new_[10712]_  = \new_[5628]_  ? \new_[12616]_  : \new_[13173]_ ;
  assign n10946 = ~\new_[12000]_ ;
  assign n10941 = ~\new_[12001]_ ;
  assign \new_[10715]_  = ~\new_[12768]_  | (~\new_[12671]_  & ~\new_[13425]_ );
  assign \new_[10716]_  = ~\new_[5283]_  | ~\new_[12341]_ ;
  assign \new_[10717]_  = ~\new_[5288]_  | ~\new_[12341]_ ;
  assign \new_[10718]_  = ~\new_[5286]_  | ~\new_[12341]_ ;
  assign \new_[10719]_  = ~\new_[5480]_  | ~\new_[14138]_ ;
  assign \new_[10720]_  = ~\new_[5290]_  | ~\new_[12341]_ ;
  assign \new_[10721]_  = ~\new_[5282]_  | ~\new_[12341]_ ;
  assign \new_[10722]_  = ~\new_[5285]_  | ~\new_[12341]_ ;
  assign \new_[10723]_  = ~\new_[3587]_  | ~\new_[12263]_ ;
  assign \new_[10724]_  = ~\new_[5287]_  | ~\new_[12341]_ ;
  assign \new_[10725]_  = ~\new_[4923]_  | ~\new_[12431]_ ;
  assign \new_[10726]_  = ~\new_[5360]_  | ~\new_[12396]_ ;
  assign \new_[10727]_  = ~\new_[5363]_  | ~\new_[12396]_ ;
  assign \new_[10728]_  = ~\new_[5365]_  | ~\new_[12396]_ ;
  assign \new_[10729]_  = ~\new_[5366]_  | ~\new_[12396]_ ;
  assign \new_[10730]_  = ~\new_[4922]_  | ~\new_[12431]_ ;
  assign \new_[10731]_  = ~\new_[4915]_  | ~\new_[12341]_ ;
  assign \new_[10732]_  = ~\new_[5284]_  | ~\new_[12341]_ ;
  assign \new_[10733]_  = ~\new_[5364]_  | ~\new_[12396]_ ;
  assign \new_[10734]_  = ~\new_[12794]_  & ~\new_[12910]_ ;
  assign \new_[10735]_  = ~\new_[5293]_  | ~\new_[12431]_ ;
  assign \new_[10736]_  = ~\new_[4909]_  | ~\new_[12431]_ ;
  assign \new_[10737]_  = ~\new_[5272]_  | ~\new_[12431]_ ;
  assign \new_[10738]_  = ~\new_[5281]_  | ~\new_[12341]_ ;
  assign \new_[10739]_  = ~\new_[4914]_  | ~\new_[12341]_ ;
  assign \new_[10740]_  = ~\new_[5295]_  | ~\new_[12431]_ ;
  assign \new_[10741]_  = ~\new_[5362]_  | ~\new_[12396]_ ;
  assign \new_[10742]_  = ~\new_[5357]_  | ~\new_[12396]_ ;
  assign \new_[10743]_  = ~\new_[5356]_  | ~\new_[12396]_ ;
  assign \new_[10744]_  = ~\new_[12395]_  & ~\new_[13020]_ ;
  assign \new_[10745]_  = ~\new_[14189]_  | ~\new_[4866]_ ;
  assign \new_[10746]_  = ~\new_[5456]_  | ~\new_[12447]_ ;
  assign \new_[10747]_  = ~\new_[5573]_  | ~\new_[12354]_ ;
  assign \new_[10748]_  = ~\new_[12469]_  & ~\new_[13003]_ ;
  assign \new_[10749]_  = ~\new_[14019]_  | ~\new_[5028]_ ;
  assign \new_[10750]_  = ~\new_[14190]_  | ~\new_[5640]_ ;
  assign \new_[10751]_  = ~\new_[14191]_  | ~\new_[5735]_ ;
  assign \new_[10752]_  = ~\new_[14033]_  | ~\new_[5589]_ ;
  assign \new_[10753]_  = ~\new_[12441]_  | ~\new_[4688]_ ;
  assign \new_[10754]_  = ~\new_[5027]_  | ~\new_[14135]_ ;
  assign \new_[10755]_  = ~\new_[12391]_  & ~\new_[12938]_ ;
  assign \new_[10756]_  = ~\new_[12395]_  & ~\new_[13053]_ ;
  assign \new_[10757]_  = ~\new_[5403]_  | ~\new_[12446]_ ;
  assign \new_[10758]_  = ~\new_[12393]_  & ~\new_[12913]_ ;
  assign \new_[10759]_  = ~\new_[12395]_  & ~\new_[12738]_ ;
  assign \new_[10760]_  = ~\new_[12393]_  & ~\new_[13020]_ ;
  assign \new_[10761]_  = ~\new_[14190]_  | ~\new_[5643]_ ;
  assign \new_[10762]_  = ~\new_[12469]_  & ~\new_[12998]_ ;
  assign \new_[10763]_  = ~\new_[5571]_  | ~\new_[12354]_ ;
  assign \new_[10764]_  = ~\new_[5261]_  | ~\new_[13930]_ ;
  assign \new_[10765]_  = ~\new_[5189]_  | ~\new_[12361]_ ;
  assign \new_[10766]_  = ~\new_[5413]_  | ~\new_[12378]_ ;
  assign \new_[10767]_  = ~\new_[5263]_  | ~\new_[13932]_ ;
  assign \new_[10768]_  = ~\new_[11626]_ ;
  assign \new_[10769]_  = ~\new_[12399]_  | ~\new_[4813]_ ;
  assign \new_[10770]_  = ~\new_[12399]_  | ~\new_[4410]_ ;
  assign \new_[10771]_  = ~\new_[14191]_  | ~\new_[5587]_ ;
  assign \new_[10772]_  = ~\new_[5555]_  | ~\new_[12354]_ ;
  assign \new_[10773]_  = ~\new_[12395]_  & ~\new_[12884]_ ;
  assign \new_[10774]_  = ~\new_[5162]_  | ~\new_[12354]_ ;
  assign \new_[10775]_  = ~\new_[12425]_  | ~\new_[4897]_ ;
  assign \new_[10776]_  = ~\new_[14189]_  | ~\new_[5655]_ ;
  assign \new_[10777]_  = ~\new_[5411]_  | ~\new_[12378]_ ;
  assign \new_[10778]_  = ~\new_[12391]_  & ~\new_[13060]_ ;
  assign \new_[10779]_  = ~\new_[5708]_  | ~\new_[12446]_ ;
  assign \new_[10780]_  = ~\new_[13882]_  | ~\new_[5650]_ ;
  assign \new_[10781]_  = ~\new_[14019]_  | ~\new_[5033]_ ;
  assign \new_[10782]_  = ~\new_[12015]_ ;
  assign \new_[10783]_  = ~\new_[4920]_  | ~\new_[12354]_ ;
  assign \new_[10784]_  = ~\new_[5412]_  | ~\new_[12378]_ ;
  assign \new_[10785]_  = ~\new_[12784]_  & ~\new_[12935]_ ;
  assign \new_[10786]_  = ~\new_[2736]_  | ~\new_[12441]_ ;
  assign \new_[10787]_  = ~\new_[12784]_  & ~\new_[13004]_ ;
  assign \new_[10788]_  = ~\new_[12391]_  & ~\new_[12738]_ ;
  assign \new_[10789]_  = ~\new_[13882]_  | ~\new_[5652]_ ;
  assign \new_[10790]_  = ~\new_[12399]_  | ~\new_[4576]_ ;
  assign \new_[10791]_  = ~\new_[13880]_  | ~\new_[5641]_ ;
  assign \new_[10792]_  = ~\new_[4987]_  | ~\new_[13993]_ ;
  assign \new_[10793]_  = ~\new_[12469]_  & ~\new_[12923]_ ;
  assign \new_[10794]_  = ~\new_[12469]_  & ~\new_[13054]_ ;
  assign \new_[10795]_  = ~\new_[5026]_  | ~\new_[14138]_ ;
  assign \new_[10796]_  = ~\new_[13972]_  | ~\new_[5612]_ ;
  assign \new_[10797]_  = ~\new_[12430]_  & ~\new_[13053]_ ;
  assign \new_[10798]_  = ~\new_[12794]_  & ~\new_[12938]_ ;
  assign \new_[10799]_  = ~\new_[12469]_  & ~\new_[12913]_ ;
  assign \new_[10800]_  = ~\new_[5570]_  | ~\new_[12352]_ ;
  assign \new_[10801]_  = ~\new_[13880]_  | ~\new_[5659]_ ;
  assign \new_[10802]_  = ~\new_[5546]_  | ~\new_[13993]_ ;
  assign \new_[10803]_  = ~\new_[14019]_  | ~\new_[5619]_ ;
  assign \new_[10804]_  = ~\new_[12264]_  | ~\new_[3764]_ ;
  assign \new_[10805]_  = ~\new_[14190]_  | ~\new_[5656]_ ;
  assign \new_[10806]_  = ~\new_[12395]_  & ~\new_[12923]_ ;
  assign \new_[10807]_  = \new_[12382]_  | \new_[12533]_ ;
  assign \new_[10808]_  = ~\new_[14189]_  | ~\new_[5875]_ ;
  assign \new_[10809]_  = ~\new_[12389]_  | ~\new_[2758]_ ;
  assign \new_[10810]_  = ~\new_[12391]_  & ~\new_[13053]_ ;
  assign \new_[10811]_  = ~\new_[12784]_  & ~\new_[13034]_ ;
  assign \new_[10812]_  = ~\new_[12391]_  & ~\new_[12939]_ ;
  assign \new_[10813]_  = ~\new_[5697]_  | ~\new_[12378]_ ;
  assign \new_[10814]_  = ~\new_[14033]_  | ~\new_[5591]_ ;
  assign \new_[10815]_  = ~\new_[11890]_ ;
  assign \new_[10816]_  = ~\new_[5531]_  | ~\new_[13992]_ ;
  assign \new_[10817]_  = ~\new_[12469]_  & ~\new_[12738]_ ;
  assign \new_[10818]_  = ~\new_[6791]_  | ~\new_[12441]_ ;
  assign \new_[10819]_  = ~\new_[12511]_ ;
  assign \new_[10820]_  = ~\new_[12466]_  & ~\new_[13046]_ ;
  assign \new_[10821]_  = ~\new_[5562]_  | ~\new_[12354]_ ;
  assign \new_[10822]_  = ~\new_[12393]_  & ~\new_[12998]_ ;
  assign \new_[10823]_  = ~\new_[12469]_  & ~\new_[12939]_ ;
  assign \new_[10824]_  = ~\new_[12469]_  & ~\new_[13053]_ ;
  assign \new_[10825]_  = ~\new_[14190]_  | ~\new_[4871]_ ;
  assign \new_[10826]_  = ~\new_[4942]_  | ~\new_[14115]_ ;
  assign \new_[10827]_  = ~\new_[5530]_  | ~\new_[13992]_ ;
  assign \new_[10828]_  = ~\new_[5534]_  | ~\new_[12354]_ ;
  assign \new_[10829]_  = ~\new_[4936]_  | ~\new_[13930]_ ;
  assign \new_[10830]_  = ~\new_[12391]_  & ~\new_[12941]_ ;
  assign \new_[10831]_  = ~\new_[5262]_  | ~\new_[13932]_ ;
  assign \new_[10832]_  = ~\new_[13882]_  | ~\new_[5755]_ ;
  assign \new_[10833]_  = ~\new_[4935]_  | ~\new_[12354]_ ;
  assign \new_[10834]_  = ~\new_[5173]_  | ~\new_[14115]_ ;
  assign \new_[10835]_  = ~\new_[5265]_  | ~\new_[13931]_ ;
  assign \new_[10836]_  = ~\new_[14033]_  | ~\new_[4821]_ ;
  assign \new_[10837]_  = ~\new_[12391]_  & ~\new_[12739]_ ;
  assign \new_[10838]_  = ~\new_[12784]_  & ~\new_[12934]_ ;
  assign \new_[10839]_  = ~\new_[13880]_  | ~\new_[4863]_ ;
  assign \new_[10840]_  = ~\new_[12425]_  | ~\new_[5634]_ ;
  assign \new_[10841]_  = ~\new_[14192]_  | ~\new_[5592]_ ;
  assign \new_[10842]_  = ~\new_[5192]_  | ~\new_[14115]_ ;
  assign \new_[10843]_  = ~\new_[12794]_  & ~\new_[13034]_ ;
  assign \new_[10844]_  = ~\new_[12425]_  | ~\new_[5009]_ ;
  assign \new_[10845]_  = ~\new_[4929]_  | ~\new_[13931]_ ;
  assign \new_[10846]_  = ~\new_[5553]_  | ~\new_[12354]_ ;
  assign \new_[10847]_  = ~\new_[5522]_  | ~\new_[13994]_ ;
  assign \new_[10848]_  = ~\new_[7686]_  | ~\new_[12441]_ ;
  assign \new_[10849]_  = ~\new_[14033]_  | ~\new_[5580]_ ;
  assign \new_[10850]_  = ~\new_[12391]_  & ~\new_[13054]_ ;
  assign \new_[10851]_  = ~\new_[5256]_  | ~\new_[13931]_ ;
  assign \new_[10852]_  = ~\new_[14033]_  | ~\new_[5748]_ ;
  assign \new_[10853]_  = ~\new_[12469]_  & ~\new_[12937]_ ;
  assign \new_[10854]_  = ~\new_[11641]_ ;
  assign \new_[10855]_  = ~\new_[14192]_  | ~\new_[5585]_ ;
  assign \new_[10856]_  = ~\new_[4972]_  | ~\new_[13993]_ ;
  assign \new_[10857]_  = ~\new_[13880]_  | ~\new_[4870]_ ;
  assign \new_[10858]_  = ~\new_[12391]_  & ~\new_[12905]_ ;
  assign \new_[10859]_  = ~\new_[12393]_  & ~\new_[12989]_ ;
  assign \new_[10860]_  = ~\new_[5544]_  | ~\new_[13992]_ ;
  assign \new_[10861]_  = ~\new_[4907]_  | ~\new_[12354]_ ;
  assign \new_[10862]_  = ~\new_[12430]_  & ~\new_[12937]_ ;
  assign \new_[10863]_  = ~\new_[7929]_  | ~\new_[12441]_ ;
  assign \new_[10864]_  = ~\new_[12786]_  & ~\new_[13004]_ ;
  assign \new_[10865]_  = ~\new_[2922]_  | ~\new_[12441]_ ;
  assign \new_[10866]_  = ~\new_[4817]_  | ~\new_[12441]_ ;
  assign \new_[10867]_  = ~\new_[12430]_  & ~\new_[13008]_ ;
  assign \new_[10868]_  = ~\new_[12381]_  | ~\new_[2757]_ ;
  assign \new_[10869]_  = ~\new_[12399]_  | ~\new_[2738]_ ;
  assign \new_[10870]_  = ~\new_[12393]_  & ~\new_[13043]_ ;
  assign \new_[10871]_  = ~\new_[12395]_  & ~\new_[12897]_ ;
  assign \new_[10872]_  = ~\new_[12794]_  & ~\new_[12999]_ ;
  assign \new_[10873]_  = ~\new_[12399]_  | ~\new_[2924]_ ;
  assign \new_[10874]_  = ~\new_[5006]_  | ~\new_[14115]_ ;
  assign \new_[10875]_  = ~\new_[5558]_  | ~\new_[12353]_ ;
  assign \new_[10876]_  = ~\new_[12264]_  | ~\new_[2717]_ ;
  assign \new_[10877]_  = ~\new_[12784]_  & ~\new_[13042]_ ;
  assign \new_[10878]_  = ~\new_[5197]_  | ~\new_[14115]_ ;
  assign \new_[10879]_  = ~\new_[5763]_  | ~\new_[12353]_ ;
  assign \new_[10880]_  = ~\new_[12393]_  & ~\new_[13060]_ ;
  assign \new_[10881]_  = ~\new_[5187]_  | ~\new_[12361]_ ;
  assign \new_[10882]_  = ~\new_[12784]_  & ~\new_[13026]_ ;
  assign \new_[10883]_  = ~\new_[5260]_  | ~\new_[13931]_ ;
  assign \new_[10884]_  = ~\new_[14164]_  | ~\new_[5693]_ ;
  assign \new_[10885]_  = ~\new_[12794]_  & ~\new_[12941]_ ;
  assign \new_[10886]_  = ~\new_[12469]_  & ~\new_[13042]_ ;
  assign \new_[10887]_  = ~\new_[12393]_  & ~\new_[13034]_ ;
  assign \new_[10888]_  = ~\new_[12354]_  | ~\new_[5543]_ ;
  assign \new_[10889]_  = ~\new_[4999]_  | ~\new_[12361]_ ;
  assign \new_[10890]_  = ~\new_[5765]_  | ~\new_[12377]_ ;
  assign \new_[10891]_  = ~\new_[12395]_  & ~\new_[13046]_ ;
  assign \new_[10892]_  = ~\new_[13972]_  | ~\new_[5611]_ ;
  assign \new_[10893]_  = ~\new_[12469]_  & ~\new_[12881]_ ;
  assign \new_[10894]_  = ~\new_[12788]_  & ~\new_[13003]_ ;
  assign \new_[10895]_  = ~\new_[12395]_  & ~\new_[12999]_ ;
  assign \new_[10896]_  = ~\new_[12395]_  & ~\new_[12998]_ ;
  assign \new_[10897]_  = ~\new_[12395]_  & ~\new_[12989]_ ;
  assign \new_[10898]_  = ~\new_[12395]_  & ~\new_[13043]_ ;
  assign \new_[10899]_  = ~\new_[5257]_  | ~\new_[13932]_ ;
  assign \new_[10900]_  = ~\new_[12393]_  & ~\new_[12923]_ ;
  assign \new_[10901]_  = ~\new_[12788]_  & ~\new_[12936]_ ;
  assign \new_[10902]_  = ~\new_[12788]_  & ~\new_[12941]_ ;
  assign \new_[10903]_  = ~\new_[12395]_  & ~\new_[12935]_ ;
  assign \new_[10904]_  = ~\new_[7875]_  | ~\new_[12441]_ ;
  assign \new_[10905]_  = ~\new_[14019]_  | ~\new_[5047]_ ;
  assign \new_[10906]_  = ~\new_[5196]_  | ~\new_[12360]_ ;
  assign \new_[10907]_  = ~\new_[5307]_  | ~\new_[12377]_ ;
  assign \new_[10908]_  = ~\new_[14164]_  | ~\new_[4876]_ ;
  assign \new_[10909]_  = ~\new_[12393]_  & ~\new_[12937]_ ;
  assign \new_[10910]_  = ~\new_[5406]_  | ~\new_[12378]_ ;
  assign \new_[10911]_  = ~\new_[4943]_  | ~\new_[13992]_ ;
  assign \new_[10912]_  = ~\new_[12395]_  & ~\new_[12913]_ ;
  assign \new_[10913]_  = ~\new_[12788]_  & ~\new_[13042]_ ;
  assign \new_[10914]_  = ~\new_[5156]_  | ~\new_[12354]_ ;
  assign \new_[10915]_  = ~\new_[12399]_  | ~\new_[3185]_ ;
  assign \new_[10916]_  = ~\new_[5487]_  | ~\new_[14138]_ ;
  assign \new_[10917]_  = ~\new_[5194]_  | ~\new_[14115]_ ;
  assign \new_[10918]_  = ~\new_[12080]_ ;
  assign \new_[10919]_  = ~\new_[5313]_  | ~\new_[12417]_ ;
  assign \new_[10920]_  = ~\new_[5538]_  | ~\new_[13992]_ ;
  assign \new_[10921]_  = ~\new_[5297]_  | ~\new_[12377]_ ;
  assign \new_[10922]_  = ~\new_[12384]_  | ~\new_[5723]_ ;
  assign \new_[10923]_  = ~\new_[5319]_  | ~\new_[12375]_ ;
  assign \new_[10924]_  = ~\new_[12383]_  | ~\new_[5677]_ ;
  assign \new_[10925]_  = ~\new_[14190]_  | ~\new_[4858]_ ;
  assign \new_[10926]_  = ~\new_[5399]_  | ~\new_[12446]_ ;
  assign \new_[10927]_  = ~\new_[4903]_  | ~\new_[12376]_ ;
  assign \new_[10928]_  = ~\new_[5764]_  | ~\new_[12377]_ ;
  assign \new_[10929]_  = ~\new_[12384]_  | ~\new_[5609]_ ;
  assign \new_[10930]_  = ~\new_[12384]_  | ~\new_[5595]_ ;
  assign \new_[10931]_  = ~\new_[5320]_  | ~\new_[12375]_ ;
  assign \new_[10932]_  = ~\new_[12383]_  | ~\new_[4836]_ ;
  assign \new_[10933]_  = ~\new_[12384]_  | ~\new_[4837]_ ;
  assign \new_[10934]_  = ~\new_[12425]_  | ~\new_[4941]_ ;
  assign \new_[10935]_  = ~\new_[12384]_  | ~\new_[5596]_ ;
  assign \new_[10936]_  = ~\new_[5563]_  | ~\new_[12353]_ ;
  assign \new_[10937]_  = ~\new_[4951]_  | ~\new_[13930]_ ;
  assign \new_[10938]_  = ~\new_[12395]_  & ~\new_[13008]_ ;
  assign \new_[10939]_  = ~\new_[5299]_  | ~\new_[12377]_ ;
  assign \new_[10940]_  = ~\new_[12384]_  | ~\new_[5717]_ ;
  assign \new_[10941]_  = ~\new_[12794]_  & ~\new_[12884]_ ;
  assign \new_[10942]_  = ~\new_[5311]_  | ~\new_[12376]_ ;
  assign \new_[10943]_  = ~\new_[14152]_  | ~\new_[5604]_ ;
  assign \new_[10944]_  = ~\new_[5300]_  | ~\new_[12377]_ ;
  assign \new_[10945]_  = ~\new_[12393]_  & ~\new_[12738]_ ;
  assign \new_[10946]_  = ~\new_[12393]_  & ~\new_[12905]_ ;
  assign \new_[10947]_  = ~\new_[14152]_  | ~\new_[5602]_ ;
  assign \new_[10948]_  = ~\new_[5301]_  | ~\new_[12375]_ ;
  assign \new_[10949]_  = ~\new_[12384]_  | ~\new_[4829]_ ;
  assign \new_[10950]_  = ~\new_[12393]_  & ~\new_[12941]_ ;
  assign \new_[10951]_  = ~\new_[5181]_  | ~\new_[14115]_ ;
  assign \new_[10952]_  = ~\new_[5547]_  | ~\new_[13993]_ ;
  assign \new_[10953]_  = ~\new_[14192]_  | ~\new_[5733]_ ;
  assign \new_[10954]_  = ~\new_[14152]_  | ~\new_[5603]_ ;
  assign \new_[10955]_  = ~\new_[2785]_  | ~\new_[12441]_ ;
  assign \new_[10956]_  = ~\new_[4904]_  | ~\new_[12377]_ ;
  assign \new_[10957]_  = ~\new_[12393]_  & ~\new_[13008]_ ;
  assign \new_[10958]_  = ~\new_[5303]_  | ~\new_[12375]_ ;
  assign \new_[10959]_  = ~\new_[12384]_  | ~\new_[4830]_ ;
  assign \new_[10960]_  = ~\new_[5314]_  | ~\new_[12376]_ ;
  assign \new_[10961]_  = ~\new_[14152]_  | ~\new_[5606]_ ;
  assign \new_[10962]_  = ~\new_[5564]_  | ~\new_[12354]_ ;
  assign \new_[10963]_  = ~\new_[14152]_  | ~\new_[5686]_ ;
  assign \new_[10964]_  = ~\new_[5316]_  | ~\new_[12417]_ ;
  assign \new_[10965]_  = ~\new_[5166]_  | ~\new_[12360]_ ;
  assign \new_[10966]_  = ~\new_[4905]_  | ~\new_[12417]_ ;
  assign \new_[10967]_  = ~\new_[12384]_  | ~\new_[4831]_ ;
  assign \new_[10968]_  = ~\new_[12786]_  & ~\new_[12934]_ ;
  assign \new_[10969]_  = ~\new_[12383]_  | ~\new_[5599]_ ;
  assign \new_[10970]_  = ~\new_[5757]_  | ~\new_[12377]_ ;
  assign \new_[10971]_  = ~\new_[14164]_  | ~\new_[4895]_ ;
  assign \new_[10972]_  = ~\new_[12469]_  & ~\new_[13043]_ ;
  assign \new_[10973]_  = ~\new_[7502]_  | ~\new_[12441]_ ;
  assign \new_[10974]_  = ~\new_[5321]_  | ~\new_[12840]_ ;
  assign \new_[10975]_  = ~\new_[12383]_  | ~\new_[5607]_ ;
  assign \new_[10976]_  = ~\new_[12384]_  | ~\new_[4835]_ ;
  assign \new_[10977]_  = ~\new_[5529]_  | ~\new_[13992]_ ;
  assign \new_[10978]_  = ~\new_[5318]_  | ~\new_[12375]_ ;
  assign \new_[10979]_  = ~\new_[14033]_  | ~\new_[5594]_ ;
  assign \new_[10980]_  = ~\new_[5031]_  | ~\new_[14134]_ ;
  assign \new_[10981]_  = ~\new_[14152]_  | ~\new_[5702]_ ;
  assign \new_[10982]_  = ~\new_[12395]_  & ~\new_[13041]_ ;
  assign \new_[10983]_  = ~\new_[5188]_  | ~\new_[12361]_ ;
  assign \new_[10984]_  = ~\new_[5560]_  | ~\new_[12354]_ ;
  assign \new_[10985]_  = ~\new_[5550]_  | ~\new_[12354]_ ;
  assign \new_[10986]_  = ~\new_[12786]_  & ~\new_[12935]_ ;
  assign \new_[10987]_  = ~\new_[12786]_  & ~\new_[13053]_ ;
  assign \new_[10988]_  = ~\new_[5310]_  | ~\new_[12376]_ ;
  assign \new_[10989]_  = ~\new_[12393]_  & ~\new_[13041]_ ;
  assign \new_[10990]_  = ~\new_[12425]_  | ~\new_[5632]_ ;
  assign \new_[10991]_  = ~\new_[12469]_  & ~\new_[12905]_ ;
  assign \new_[10992]_  = ~\new_[12425]_  | ~\new_[5639]_ ;
  assign \new_[10993]_  = ~\new_[5317]_  | ~\new_[12377]_ ;
  assign \new_[10994]_  = ~\new_[12393]_  & ~\new_[12910]_ ;
  assign \new_[10995]_  = ~\new_[12393]_  & ~\new_[12936]_ ;
  assign \new_[10996]_  = ~\new_[5247]_  | ~\new_[13930]_ ;
  assign \new_[10997]_  = ~\new_[14190]_  | ~\new_[4877]_ ;
  assign \new_[10998]_  = ~\new_[12393]_  & ~\new_[12939]_ ;
  assign \new_[10999]_  = ~\new_[12469]_  & ~\new_[12989]_ ;
  assign \new_[11000]_  = ~\new_[14019]_  | ~\new_[4842]_ ;
  assign \new_[11001]_  = ~\new_[5453]_  | ~\new_[12447]_ ;
  assign \new_[11002]_  = ~\new_[13879]_  | ~\new_[5653]_ ;
  assign \new_[11003]_  = ~\new_[14189]_  | ~\new_[5734]_ ;
  assign \new_[11004]_  = ~\new_[5537]_  | ~\new_[13992]_ ;
  assign \new_[11005]_  = ~\new_[14033]_  | ~\new_[5593]_ ;
  assign \new_[11006]_  = ~\new_[13880]_  | ~\new_[4912]_ ;
  assign \new_[11007]_  = ~\new_[12430]_  & ~\new_[12923]_ ;
  assign \new_[11008]_  = ~\new_[13972]_  | ~\new_[5623]_ ;
  assign \new_[11009]_  = ~\new_[12784]_  & ~\new_[12989]_ ;
  assign \new_[11010]_  = ~\new_[14164]_  | ~\new_[5664]_ ;
  assign \new_[11011]_  = ~\new_[12399]_  | ~\new_[2749]_ ;
  assign \new_[11012]_  = ~\new_[13972]_  | ~\new_[4845]_ ;
  assign \new_[11013]_  = ~\new_[14190]_  | ~\new_[5777]_ ;
  assign \new_[11014]_  = ~\new_[5542]_  | ~\new_[13993]_ ;
  assign \new_[11015]_  = ~\new_[5577]_  | ~\new_[12352]_ ;
  assign \new_[11016]_  = ~\new_[4993]_  | ~\new_[14115]_ ;
  assign \new_[11017]_  = ~\new_[14019]_  | ~\new_[5620]_ ;
  assign \new_[11018]_  = ~\new_[14192]_  | ~\new_[4819]_ ;
  assign \new_[11019]_  = ~\new_[12101]_ ;
  assign \new_[11020]_  = ~\new_[11688]_ ;
  assign \new_[11021]_  = ~\new_[13880]_  | ~\new_[4867]_ ;
  assign \new_[11022]_  = ~\new_[5025]_  | ~\new_[12354]_ ;
  assign \new_[11023]_  = ~\new_[14033]_  | ~\new_[5586]_ ;
  assign \new_[11024]_  = ~\new_[12430]_  & ~\new_[12989]_ ;
  assign \new_[11025]_  = ~\new_[12430]_  & ~\new_[12884]_ ;
  assign \new_[11026]_  = ~\new_[12430]_  & ~\new_[12910]_ ;
  assign \new_[11027]_  = ~\new_[4901]_  | ~\new_[12376]_ ;
  assign \new_[11028]_  = ~\new_[12264]_  | ~\new_[4584]_ ;
  assign \new_[11029]_  = ~\new_[12430]_  & ~\new_[12941]_ ;
  assign \new_[11030]_  = ~\new_[12817]_  & ~\new_[13041]_ ;
  assign \new_[11031]_  = ~\new_[5182]_  | ~\new_[14115]_ ;
  assign \new_[11032]_  = ~\new_[14019]_  | ~\new_[5614]_ ;
  assign \new_[11033]_  = ~\new_[5034]_  | ~\new_[12447]_ ;
  assign \new_[11034]_  = ~\new_[12817]_  & ~\new_[12905]_ ;
  assign \new_[11035]_  = ~\new_[5190]_  | ~\new_[12361]_ ;
  assign \new_[11036]_  = ~\new_[12393]_  & ~\new_[12884]_ ;
  assign \new_[11037]_  = ~\new_[5473]_  | ~\new_[14135]_ ;
  assign \new_[11038]_  = ~\new_[5180]_  | ~\new_[14115]_ ;
  assign \new_[11039]_  = ~\new_[12430]_  & ~\new_[13042]_ ;
  assign \new_[11040]_  = ~\new_[12817]_  & ~\new_[12913]_ ;
  assign \new_[11041]_  = ~\new_[12817]_  & ~\new_[12934]_ ;
  assign \new_[11042]_  = ~\new_[5030]_  | ~\new_[14135]_ ;
  assign \new_[11043]_  = ~\new_[12430]_  & ~\new_[13054]_ ;
  assign \new_[11044]_  = ~\new_[4938]_  | ~\new_[13932]_ ;
  assign \new_[11045]_  = ~\new_[14191]_  | ~\new_[5584]_ ;
  assign \new_[11046]_  = ~\new_[5136]_  | ~\new_[12354]_ ;
  assign \new_[11047]_  = ~\new_[5491]_  | ~\new_[14138]_ ;
  assign \new_[11048]_  = ~\new_[5470]_  | ~\new_[12447]_ ;
  assign \new_[11049]_  = ~\new_[14191]_  | ~\new_[4822]_ ;
  assign \new_[11050]_  = ~\new_[12469]_  & ~\new_[13041]_ ;
  assign \new_[11051]_  = ~\new_[5528]_  | ~\new_[13993]_ ;
  assign \new_[11052]_  = ~\new_[13972]_  | ~\new_[5669]_ ;
  assign \new_[11053]_  = ~\new_[5524]_  | ~\new_[13993]_ ;
  assign \new_[11054]_  = ~\new_[5472]_  | ~\new_[14138]_ ;
  assign \new_[11055]_  = ~\new_[13972]_  | ~\new_[5029]_ ;
  assign \new_[11056]_  = ~\new_[5408]_  | ~\new_[12378]_ ;
  assign \new_[11057]_  = ~\new_[5474]_  | ~\new_[14134]_ ;
  assign \new_[11058]_  = ~\new_[11696]_ ;
  assign \new_[11059]_  = ~\new_[5420]_  | ~\new_[12446]_ ;
  assign \new_[11060]_  = ~\new_[12391]_  & ~\new_[12881]_ ;
  assign \new_[11061]_  = ~\new_[4916]_  | ~\new_[13993]_ ;
  assign \new_[11062]_  = ~\new_[5312]_  | ~\new_[12376]_ ;
  assign \new_[11063]_  = ~\new_[14019]_  | ~\new_[4843]_ ;
  assign \new_[11064]_  = ~\new_[5574]_  | ~\new_[12352]_ ;
  assign \new_[11065]_  = ~\new_[13972]_  | ~\new_[4986]_ ;
  assign \new_[11066]_  = ~\new_[14189]_  | ~\new_[5648]_ ;
  assign \new_[11067]_  = ~\new_[2747]_  | ~\new_[12441]_ ;
  assign \new_[11068]_  = ~\new_[5410]_  | ~\new_[12378]_ ;
  assign \new_[11069]_  = ~\new_[12469]_  & ~\new_[12897]_ ;
  assign \new_[11070]_  = ~\new_[5527]_  | ~\new_[13992]_ ;
  assign \new_[11071]_  = ~\new_[14192]_  | ~\new_[5579]_ ;
  assign \new_[11072]_  = ~\new_[12794]_  & ~\new_[12936]_ ;
  assign \new_[11073]_  = ~\new_[5540]_  | ~\new_[13992]_ ;
  assign \new_[11074]_  = ~\new_[14019]_  | ~\new_[5617]_ ;
  assign \new_[11075]_  = ~\new_[14152]_  | ~\new_[4833]_ ;
  assign \new_[11076]_  = ~\new_[13972]_  | ~\new_[5618]_ ;
  assign \new_[11077]_  = ~\new_[5309]_  | ~\new_[12376]_ ;
  assign \new_[11078]_  = ~\new_[12391]_  & ~\new_[12937]_ ;
  assign \new_[11079]_  = ~\new_[13879]_  | ~\new_[5703]_ ;
  assign \new_[11080]_  = ~\new_[12469]_  & ~\new_[13026]_ ;
  assign \new_[11081]_  = ~\new_[12430]_  & ~\new_[12881]_ ;
  assign \new_[11082]_  = ~\new_[11705]_ ;
  assign \new_[11083]_  = ~\new_[11706]_ ;
  assign \new_[11084]_  = ~\new_[5148]_  | ~\new_[14181]_ ;
  assign \new_[11085]_  = ~\new_[12430]_  & ~\new_[12938]_ ;
  assign \new_[11086]_  = ~\new_[13972]_  | ~\new_[5621]_ ;
  assign \new_[11087]_  = ~\new_[12399]_  | ~\new_[2718]_ ;
  assign \new_[11088]_  = ~\new_[14019]_  | ~\new_[5358]_ ;
  assign \new_[11089]_  = ~\new_[12399]_  | ~\new_[2787]_ ;
  assign \new_[11090]_  = ~\new_[5414]_  | ~\new_[12378]_ ;
  assign \new_[11091]_  = ~\new_[12430]_  & ~\new_[12936]_ ;
  assign \new_[11092]_  = ~\new_[4908]_  | ~\new_[12352]_ ;
  assign \new_[11093]_  = ~\new_[5415]_  | ~\new_[12378]_ ;
  assign \new_[11094]_  = ~\new_[13972]_  | ~\new_[4841]_ ;
  assign \new_[11095]_  = ~\new_[5405]_  | ~\new_[12446]_ ;
  assign \new_[11096]_  = ~\new_[5306]_  | ~\new_[12377]_ ;
  assign \new_[11097]_  = ~\new_[5416]_  | ~\new_[12446]_ ;
  assign \new_[11098]_  = ~\new_[5138]_  | ~\new_[12354]_ ;
  assign \new_[11099]_  = ~\new_[12425]_  | ~\new_[4853]_ ;
  assign \new_[11100]_  = ~\new_[12384]_  | ~\new_[4834]_ ;
  assign \new_[11101]_  = ~\new_[5520]_  | ~\new_[13993]_ ;
  assign \new_[11102]_  = ~\new_[14019]_  | ~\new_[5505]_ ;
  assign \new_[11103]_  = ~\new_[12393]_  & ~\new_[12897]_ ;
  assign \new_[11104]_  = ~\new_[5407]_  | ~\new_[12378]_ ;
  assign \new_[11105]_  = ~\new_[13972]_  | ~\new_[5616]_ ;
  assign \new_[11106]_  = ~\new_[12264]_  | ~\new_[2737]_ ;
  assign \new_[11107]_  = ~\new_[14033]_  | ~\new_[4824]_ ;
  assign \new_[11108]_  = ~\new_[12786]_  & ~\new_[13026]_ ;
  assign \new_[11109]_  = ~\new_[12469]_  & ~\new_[13020]_ ;
  assign \new_[11110]_  = ~\new_[12817]_  & ~\new_[13034]_ ;
  assign \new_[11111]_  = ~\new_[13882]_  | ~\new_[5649]_ ;
  assign \new_[11112]_  = ~\new_[5479]_  | ~\new_[14135]_ ;
  assign \new_[11113]_  = ~\new_[12430]_  & ~\new_[13020]_ ;
  assign \new_[11114]_  = ~\new_[5304]_  | ~\new_[12377]_ ;
  assign \new_[11115]_  = ~\new_[12430]_  & ~\new_[13046]_ ;
  assign \new_[11116]_  = ~\new_[12691]_ ;
  assign \new_[11117]_  = ~\new_[12393]_  & ~\new_[13042]_ ;
  assign \new_[11118]_  = ~\new_[3601]_  | ~\new_[12399]_ ;
  assign \new_[11119]_  = ~\new_[5177]_  | ~\new_[12360]_ ;
  assign \new_[11120]_  = ~\new_[12430]_  & ~\new_[12739]_ ;
  assign \new_[11121]_  = ~\new_[5539]_  | ~\new_[13992]_ ;
  assign \new_[11122]_  = ~\new_[12469]_  & ~\new_[12739]_ ;
  assign \new_[11123]_  = ~\new_[5154]_  | ~\new_[12354]_ ;
  assign \new_[11124]_  = ~\new_[5258]_  | ~\new_[13932]_ ;
  assign \new_[11125]_  = ~\new_[13879]_  | ~\new_[4872]_ ;
  assign \new_[11126]_  = ~\new_[12430]_  & ~\new_[12738]_ ;
  assign \new_[11127]_  = ~\new_[12788]_  & ~\new_[12938]_ ;
  assign \new_[11128]_  = ~\new_[12430]_  & ~\new_[13004]_ ;
  assign \new_[11129]_  = ~\new_[13879]_  | ~\new_[4864]_ ;
  assign \new_[11130]_  = ~\new_[14189]_  | ~\new_[4875]_ ;
  assign \new_[11131]_  = ~\new_[5145]_  | ~\new_[12354]_ ;
  assign \new_[11132]_  = ~\new_[4906]_  | ~\new_[12377]_ ;
  assign \new_[11133]_  = ~\new_[12430]_  & ~\new_[12935]_ ;
  assign \new_[11134]_  = ~\new_[14164]_  | ~\new_[5858]_ ;
  assign \new_[11135]_  = ~\new_[12425]_  | ~\new_[5630]_ ;
  assign \new_[11136]_  = ~\new_[12393]_  & ~\new_[12739]_ ;
  assign \new_[11137]_  = ~\new_[13880]_  | ~\new_[4868]_ ;
  assign \new_[11138]_  = ~\new_[5179]_  | ~\new_[14115]_ ;
  assign \new_[11139]_  = ~\new_[12399]_  | ~\new_[3672]_ ;
  assign \new_[11140]_  = ~\new_[13972]_  | ~\new_[4844]_ ;
  assign \new_[11141]_  = ~\new_[11727]_ ;
  assign \new_[11142]_  = ~\new_[12425]_  | ~\new_[4852]_ ;
  assign \new_[11143]_  = ~\new_[12788]_  & ~\new_[13026]_ ;
  assign \new_[11144]_  = ~\new_[11698]_ ;
  assign \new_[11145]_  = ~\new_[14191]_  | ~\new_[5719]_ ;
  assign \new_[11146]_  = ~\new_[12393]_  & ~\new_[13003]_ ;
  assign \new_[11147]_  = \new_[12776]_  | \new_[2757]_ ;
  assign \new_[11148]_  = ~\new_[12784]_  & ~\new_[12999]_ ;
  assign \new_[11149]_  = ~\new_[14189]_  | ~\new_[5663]_ ;
  assign \new_[11150]_  = ~\new_[4937]_  | ~\new_[13931]_ ;
  assign \new_[11151]_  = ~\new_[14152]_  | ~\new_[5695]_ ;
  assign \new_[11152]_  = ~\new_[5184]_  | ~\new_[12361]_ ;
  assign \new_[11153]_  = ~\new_[14033]_  | ~\new_[5581]_ ;
  assign \new_[11154]_  = ~\new_[12264]_  | ~\new_[3184]_ ;
  assign \new_[11155]_  = ~\new_[14033]_  | ~\new_[4826]_ ;
  assign \new_[11156]_  = ~\new_[12393]_  & ~\new_[13054]_ ;
  assign \new_[11157]_  = ~\new_[12794]_  & ~\new_[12935]_ ;
  assign \new_[11158]_  = ~\new_[12817]_  & ~\new_[12939]_ ;
  assign \new_[11159]_  = ~\new_[13879]_  | ~\new_[4869]_ ;
  assign \new_[11160]_  = ~\new_[5526]_  | ~\new_[13993]_ ;
  assign \new_[11161]_  = ~\new_[14033]_  | ~\new_[5583]_ ;
  assign \new_[11162]_  = ~\new_[5471]_  | ~\new_[14134]_ ;
  assign \new_[11163]_  = ~\new_[12425]_  | ~\new_[4854]_ ;
  assign \new_[11164]_  = ~\new_[5013]_  | ~\new_[14138]_ ;
  assign \new_[11165]_  = ~\new_[11673]_ ;
  assign \new_[11166]_  = ~\new_[12364]_  & ~\new_[12934]_ ;
  assign \new_[11167]_  = ~\new_[5494]_  | ~\new_[14138]_ ;
  assign \new_[11168]_  = ~\new_[12817]_  & ~\new_[13043]_ ;
  assign \new_[11169]_  = ~\new_[12393]_  & ~\new_[13046]_ ;
  assign \new_[11170]_  = ~\new_[12788]_  & ~\new_[13034]_ ;
  assign \new_[11171]_  = ~\new_[12391]_  & ~\new_[12936]_ ;
  assign \new_[11172]_  = ~\new_[12425]_  | ~\new_[4848]_ ;
  assign \new_[11173]_  = ~\new_[12788]_  & ~\new_[12905]_ ;
  assign \new_[11174]_  = ~\new_[14189]_  | ~\new_[5651]_ ;
  assign \new_[11175]_  = ~\new_[5475]_  | ~\new_[14135]_ ;
  assign \new_[11176]_  = ~\new_[5409]_  | ~\new_[12378]_ ;
  assign \new_[11177]_  = ~\new_[12391]_  & ~\new_[12910]_ ;
  assign \new_[11178]_  = ~\new_[12395]_  & ~\new_[12934]_ ;
  assign \new_[11179]_  = ~\new_[12425]_  | ~\new_[5633]_ ;
  assign \new_[11180]_  = ~\new_[12395]_  & ~\new_[12910]_ ;
  assign \new_[11181]_  = ~\new_[14191]_  | ~\new_[5726]_ ;
  assign \new_[11182]_  = ~\new_[14190]_  | ~\new_[5701]_ ;
  assign \new_[11183]_  = ~\new_[12391]_  & ~\new_[13041]_ ;
  assign \new_[11184]_  = ~\new_[12786]_  & ~\new_[12999]_ ;
  assign \new_[11185]_  = ~\new_[5023]_  | ~\new_[14135]_ ;
  assign \new_[11186]_  = ~\new_[12384]_  | ~\new_[4828]_ ;
  assign \new_[11187]_  = ~\new_[5467]_  | ~\new_[12447]_ ;
  assign \new_[11188]_  = ~\new_[14033]_  | ~\new_[5753]_ ;
  assign \new_[11189]_  = ~\new_[12395]_  & ~\new_[12939]_ ;
  assign \new_[11190]_  = ~\new_[5856]_  | ~\new_[12441]_ ;
  assign \new_[11191]_  = ~\new_[12817]_  & ~\new_[12998]_ ;
  assign \new_[11192]_  = ~\new_[5578]_  | ~\new_[12354]_ ;
  assign \new_[11193]_  = ~\new_[12391]_  & ~\new_[13046]_ ;
  assign \new_[11194]_  = ~\new_[13880]_  | ~\new_[5744]_ ;
  assign \new_[11195]_  = ~\new_[12430]_  & ~\new_[13060]_ ;
  assign \new_[11196]_  = ~\new_[4948]_  | ~\new_[13994]_ ;
  assign \new_[11197]_  = ~\new_[12430]_  & ~\new_[12999]_ ;
  assign \new_[11198]_  = ~\new_[14190]_  | ~\new_[4860]_ ;
  assign \new_[11199]_  = ~\new_[12469]_  & ~\new_[13060]_ ;
  assign \new_[11200]_  = ~\new_[12430]_  & ~\new_[12897]_ ;
  assign \new_[11201]_  = ~\new_[12395]_  & ~\new_[13004]_ ;
  assign \new_[11202]_  = ~\new_[5159]_  | ~\new_[12354]_ ;
  assign \new_[11203]_  = ~\new_[14191]_  | ~\new_[5588]_ ;
  assign \new_[11204]_  = ~\new_[14019]_  | ~\new_[4847]_ ;
  assign \new_[11205]_  = ~\new_[14190]_  | ~\new_[5665]_ ;
  assign \new_[11206]_  = ~\new_[5569]_  | ~\new_[12354]_ ;
  assign \new_[11207]_  = ~\new_[12399]_  | ~\new_[7688]_ ;
  assign \new_[11208]_  = ~\new_[13879]_  | ~\new_[5731]_ ;
  assign \new_[11209]_  = ~\new_[11747]_ ;
  assign \new_[11210]_  = ~\new_[14164]_  | ~\new_[4874]_ ;
  assign \new_[11211]_  = ~\new_[12786]_  & ~\new_[12881]_ ;
  assign \new_[11212]_  = ~\new_[5535]_  | ~\new_[13992]_ ;
  assign \new_[11213]_  = ~\new_[14164]_  | ~\new_[4963]_ ;
  assign \new_[11214]_  = ~\new_[5183]_  | ~\new_[12361]_ ;
  assign \new_[11215]_  = ~\new_[12391]_  & ~\new_[13003]_ ;
  assign \new_[11216]_  = ~\new_[5759]_  | ~\new_[12354]_ ;
  assign \new_[11217]_  = ~\new_[13972]_  | ~\new_[5624]_ ;
  assign \new_[11218]_  = ~\new_[12469]_  & ~\new_[13004]_ ;
  assign \new_[11219]_  = ~\new_[5668]_  | ~\new_[12378]_ ;
  assign \new_[11220]_  = ~\new_[12469]_  & ~\new_[12934]_ ;
  assign \new_[11221]_  = ~\new_[5250]_  | ~\new_[13932]_ ;
  assign \new_[11222]_  = ~\new_[12391]_  & ~\new_[12884]_ ;
  assign \new_[11223]_  = ~\new_[5298]_  | ~\new_[12377]_ ;
  assign \new_[11224]_  = ~\new_[14190]_  | ~\new_[5658]_ ;
  assign \new_[11225]_  = ~\new_[12391]_  & ~\new_[13043]_ ;
  assign \new_[11226]_  = ~\new_[13880]_  | ~\new_[4861]_ ;
  assign \new_[11227]_  = ~\new_[14191]_  | ~\new_[4820]_ ;
  assign \new_[11228]_  = ~\new_[5000]_  | ~\new_[14115]_ ;
  assign \new_[11229]_  = ~\new_[5259]_  | ~\new_[13932]_ ;
  assign \new_[11230]_  = ~\new_[5191]_  | ~\new_[12361]_ ;
  assign \new_[11231]_  = ~\new_[11749]_ ;
  assign \new_[11232]_  = ~\new_[14189]_  | ~\new_[5645]_ ;
  assign \new_[11233]_  = ~\new_[5164]_  | ~\new_[14115]_ ;
  assign \new_[11234]_  = ~\new_[5521]_  | ~\new_[13993]_ ;
  assign \new_[11235]_  = ~\new_[5568]_  | ~\new_[12352]_ ;
  assign \new_[11236]_  = ~\new_[12469]_  & ~\new_[13046]_ ;
  assign \new_[11237]_  = ~\new_[14152]_  | ~\new_[4832]_ ;
  assign \new_[11238]_  = ~\new_[5308]_  | ~\new_[12376]_ ;
  assign \new_[11239]_  = ~\new_[13880]_  | ~\new_[5642]_ ;
  assign \new_[11240]_  = ~\new_[11722]_ ;
  assign \new_[11241]_  = ~\new_[12391]_  & ~\new_[12923]_ ;
  assign \new_[11242]_  = ~\new_[12395]_  & ~\new_[12881]_ ;
  assign \new_[11243]_  = ~\new_[5523]_  | ~\new_[13993]_ ;
  assign \new_[11244]_  = ~\new_[12391]_  & ~\new_[13020]_ ;
  assign \new_[11245]_  = ~\new_[12469]_  & ~\new_[13008]_ ;
  assign \new_[11246]_  = ~\new_[5195]_  | ~\new_[12360]_ ;
  assign \new_[11247]_  = ~\new_[12395]_  & ~\new_[12937]_ ;
  assign \new_[11248]_  = ~\new_[13882]_  | ~\new_[5654]_ ;
  assign \new_[11249]_  = ~\new_[5525]_  | ~\new_[13994]_ ;
  assign \new_[11250]_  = ~\new_[5152]_  | ~\new_[12354]_ ;
  assign \new_[11251]_  = ~\new_[12391]_  & ~\new_[12913]_ ;
  assign \new_[11252]_  = ~\new_[5193]_  | ~\new_[12360]_ ;
  assign \new_[11253]_  = ~\new_[5143]_  | ~\new_[12354]_ ;
  assign \new_[11254]_  = ~\new_[5296]_  | ~\new_[12361]_ ;
  assign \new_[11255]_  = ~\new_[14192]_  | ~\new_[4827]_ ;
  assign \new_[11256]_  = ~\new_[13880]_  | ~\new_[5647]_ ;
  assign \new_[11257]_  = ~\new_[4964]_  | ~\new_[13992]_ ;
  assign \new_[11258]_  = ~\new_[12264]_  | ~\new_[2726]_ ;
  assign \new_[11259]_  = ~\new_[13879]_  | ~\new_[5725]_ ;
  assign \new_[11260]_  = ~\new_[12395]_  & ~\new_[12739]_ ;
  assign \new_[11261]_  = ~\new_[5565]_  | ~\new_[12352]_ ;
  assign \new_[11262]_  = ~\new_[12384]_  | ~\new_[5597]_ ;
  assign \new_[11263]_  = ~\new_[13879]_  | ~\new_[4873]_ ;
  assign \new_[11264]_  = ~\new_[12384]_  | ~\new_[5715]_ ;
  assign \new_[11265]_  = ~\new_[14164]_  | ~\new_[4913]_ ;
  assign \new_[11266]_  = ~\new_[12391]_  & ~\new_[12897]_ ;
  assign \new_[11267]_  = ~\new_[5315]_  | ~\new_[12377]_ ;
  assign \new_[11268]_  = ~\new_[14189]_  | ~\new_[5657]_ ;
  assign \new_[11269]_  = ~\new_[14019]_  | ~\new_[5622]_ ;
  assign \new_[11270]_  = ~\new_[12430]_  & ~\new_[13026]_ ;
  assign \new_[11271]_  = ~\new_[13880]_  | ~\new_[4862]_ ;
  assign \new_[11272]_  = ~\new_[5532]_  | ~\new_[13992]_ ;
  assign \new_[11273]_  = ~\new_[12391]_  & ~\new_[12998]_ ;
  assign \new_[11274]_  = ~\new_[4973]_  | ~\new_[13992]_ ;
  assign \new_[11275]_  = ~\new_[5268]_  | ~\new_[13930]_ ;
  assign \new_[11276]_  = ~\new_[5536]_  | ~\new_[14181]_ ;
  assign \new_[11277]_  = ~\new_[13882]_  | ~\new_[5766]_ ;
  assign \new_[11278]_  = ~\new_[5548]_  | ~\new_[13994]_ ;
  assign \new_[11279]_  = ~\new_[4998]_  | ~\new_[12361]_ ;
  assign \new_[11280]_  = ~\new_[13880]_  | ~\new_[5662]_ ;
  assign \new_[11281]_  = ~\new_[4962]_  | ~\new_[13992]_ ;
  assign \new_[11282]_  = ~\new_[12357]_  & ~\new_[12935]_ ;
  assign \new_[11283]_  = ~\new_[12464]_  & ~\new_[12923]_ ;
  assign \new_[11284]_  = ~\new_[12379]_  & ~\new_[13003]_ ;
  assign \new_[11285]_  = ~\new_[12357]_  & ~\new_[13042]_ ;
  assign \new_[11286]_  = ~\new_[12365]_  & ~\new_[13054]_ ;
  assign \new_[11287]_  = ~\new_[13880]_  | ~\new_[5660]_ ;
  assign \new_[11288]_  = ~\new_[12464]_  & ~\new_[12935]_ ;
  assign \new_[11289]_  = ~\new_[12464]_  & ~\new_[13003]_ ;
  assign \new_[11290]_  = ~\new_[12365]_  & ~\new_[12739]_ ;
  assign \new_[11291]_  = ~\new_[12379]_  & ~\new_[12905]_ ;
  assign \new_[11292]_  = ~\new_[12379]_  & ~\new_[12937]_ ;
  assign \new_[11293]_  = ~\new_[12365]_  & ~\new_[13008]_ ;
  assign \new_[11294]_  = ~\new_[12743]_  & ~\new_[12941]_ ;
  assign \new_[11295]_  = ~\new_[12445]_  & ~\new_[12884]_ ;
  assign \new_[11296]_  = ~\new_[12379]_  & ~\new_[12935]_ ;
  assign \new_[11297]_  = ~\new_[12464]_  & ~\new_[12884]_ ;
  assign \new_[11298]_  = ~\new_[12442]_  & ~\new_[13041]_ ;
  assign \new_[11299]_  = ~\new_[12428]_  & ~\new_[13003]_ ;
  assign \new_[11300]_  = ~\new_[12743]_  & ~\new_[13053]_ ;
  assign \new_[11301]_  = ~\new_[12371]_  & ~\new_[12939]_ ;
  assign \new_[11302]_  = ~\new_[12461]_  & ~\new_[12989]_ ;
  assign \new_[11303]_  = ~\new_[12357]_  & ~\new_[12999]_ ;
  assign \new_[11304]_  = ~\new_[12443]_  & ~\new_[12913]_ ;
  assign \new_[11305]_  = ~\new_[12395]_  & ~\new_[13054]_ ;
  assign \new_[11306]_  = ~\new_[12379]_  & ~\new_[13043]_ ;
  assign \new_[11307]_  = ~\new_[12365]_  & ~\new_[12905]_ ;
  assign \new_[11308]_  = ~\new_[12812]_  & ~\new_[13026]_ ;
  assign \new_[11309]_  = ~\new_[12449]_  & ~\new_[12738]_ ;
  assign \new_[11310]_  = ~\new_[12357]_  & ~\new_[12913]_ ;
  assign \new_[11311]_  = ~\new_[12459]_  & ~\new_[12738]_ ;
  assign \new_[11312]_  = ~\new_[12374]_  & ~\new_[13046]_ ;
  assign \new_[11313]_  = ~\new_[12364]_  & ~\new_[12913]_ ;
  assign \new_[11314]_  = ~\new_[12364]_  & ~\new_[12884]_ ;
  assign \new_[11315]_  = ~\new_[12834]_  & ~\new_[12910]_ ;
  assign \new_[11316]_  = ~\new_[12834]_  & ~\new_[12934]_ ;
  assign \new_[11317]_  = ~\new_[12355]_  & ~\new_[12910]_ ;
  assign \new_[11318]_  = ~\new_[12812]_  & ~\new_[13041]_ ;
  assign \new_[11319]_  = ~\new_[12459]_  & ~\new_[12913]_ ;
  assign \new_[11320]_  = ~\new_[12834]_  & ~\new_[12923]_ ;
  assign \new_[11321]_  = ~\new_[12364]_  & ~\new_[13060]_ ;
  assign \new_[11322]_  = ~\new_[12358]_  & ~\new_[12937]_ ;
  assign \new_[11323]_  = ~\new_[12466]_  & ~\new_[13026]_ ;
  assign \new_[11324]_  = ~\new_[12850]_  & ~\new_[12923]_ ;
  assign \new_[11325]_  = ~\new_[12850]_  & ~\new_[13053]_ ;
  assign \new_[11326]_  = ~\new_[12786]_  & ~\new_[12938]_ ;
  assign \new_[11327]_  = ~\new_[12371]_  & ~\new_[13034]_ ;
  assign \new_[11328]_  = ~\new_[12428]_  & ~\new_[13026]_ ;
  assign \new_[11329]_  = ~\new_[12374]_  & ~\new_[12935]_ ;
  assign \new_[11330]_  = ~\new_[12743]_  & ~\new_[12905]_ ;
  assign \new_[11331]_  = ~\new_[12359]_  & ~\new_[13034]_ ;
  assign \new_[11332]_  = ~\new_[12444]_  & ~\new_[13008]_ ;
  assign \new_[11333]_  = ~\new_[12443]_  & ~\new_[12739]_ ;
  assign \new_[11334]_  = ~\new_[12449]_  & ~\new_[12881]_ ;
  assign \new_[11335]_  = ~\new_[12364]_  & ~\new_[13034]_ ;
  assign \new_[11336]_  = ~\new_[12743]_  & ~\new_[13060]_ ;
  assign \new_[11337]_  = ~\new_[12364]_  & ~\new_[12936]_ ;
  assign \new_[11338]_  = ~\new_[12834]_  & ~\new_[13020]_ ;
  assign \new_[11339]_  = ~\new_[12359]_  & ~\new_[12897]_ ;
  assign \new_[11340]_  = ~\new_[12442]_  & ~\new_[13042]_ ;
  assign \new_[11341]_  = ~\new_[12428]_  & ~\new_[12998]_ ;
  assign \new_[11342]_  = ~\new_[12850]_  & ~\new_[13020]_ ;
  assign \new_[11343]_  = ~\new_[12461]_  & ~\new_[12998]_ ;
  assign \new_[11344]_  = ~\new_[12356]_  & ~\new_[12905]_ ;
  assign \new_[11345]_  = ~\new_[12430]_  & ~\new_[13003]_ ;
  assign \new_[11346]_  = ~\new_[12355]_  & ~\new_[12934]_ ;
  assign \new_[11347]_  = ~\new_[12379]_  & ~\new_[12989]_ ;
  assign \new_[11348]_  = ~\new_[12812]_  & ~\new_[13053]_ ;
  assign \new_[11349]_  = ~\new_[12364]_  & ~\new_[12938]_ ;
  assign \new_[11350]_  = ~\new_[12359]_  & ~\new_[12936]_ ;
  assign \new_[11351]_  = ~\new_[12459]_  & ~\new_[13042]_ ;
  assign \new_[11352]_  = ~\new_[12834]_  & ~\new_[13034]_ ;
  assign \new_[11353]_  = ~\new_[12850]_  & ~\new_[12989]_ ;
  assign \new_[11354]_  = ~\new_[12850]_  & ~\new_[12999]_ ;
  assign \new_[11355]_  = ~\new_[12371]_  & ~\new_[13008]_ ;
  assign \new_[11356]_  = ~\new_[12358]_  & ~\new_[13043]_ ;
  assign \new_[11357]_  = ~\new_[12449]_  & ~\new_[13042]_ ;
  assign \new_[11358]_  = ~\new_[12743]_  & ~\new_[12934]_ ;
  assign \new_[11359]_  = ~\new_[12364]_  & ~\new_[12897]_ ;
  assign \new_[11360]_  = ~\new_[12359]_  & ~\new_[12738]_ ;
  assign \new_[11361]_  = ~\new_[12356]_  & ~\new_[13054]_ ;
  assign \new_[11362]_  = ~\new_[12812]_  & ~\new_[13004]_ ;
  assign \new_[11363]_  = ~\new_[12834]_  & ~\new_[12939]_ ;
  assign \new_[11364]_  = ~\new_[12355]_  & ~\new_[12989]_ ;
  assign \new_[11365]_  = ~\new_[12371]_  & ~\new_[13004]_ ;
  assign \new_[11366]_  = ~\new_[12356]_  & ~\new_[13003]_ ;
  assign \new_[11367]_  = ~\new_[14033]_  | ~\new_[4823]_ ;
  assign \new_[11368]_  = ~\new_[12356]_  & ~\new_[13060]_ ;
  assign \new_[11369]_  = ~\new_[12371]_  & ~\new_[12897]_ ;
  assign \new_[11370]_  = ~\new_[12445]_  & ~\new_[12738]_ ;
  assign \new_[11371]_  = ~\new_[12466]_  & ~\new_[12936]_ ;
  assign \new_[11372]_  = ~\new_[12355]_  & ~\new_[13020]_ ;
  assign \new_[11373]_  = ~\new_[12358]_  & ~\new_[12884]_ ;
  assign \new_[11374]_  = ~\new_[12358]_  & ~\new_[12881]_ ;
  assign \new_[11375]_  = ~\new_[12444]_  & ~\new_[13054]_ ;
  assign \new_[11376]_  = ~\new_[12355]_  & ~\new_[12938]_ ;
  assign \new_[11377]_  = ~\new_[12850]_  & ~\new_[12941]_ ;
  assign \new_[11378]_  = ~\new_[12834]_  & ~\new_[12998]_ ;
  assign \new_[11379]_  = ~\new_[12834]_  & ~\new_[12999]_ ;
  assign \new_[11380]_  = ~\new_[12444]_  & ~\new_[13060]_ ;
  assign \new_[11381]_  = ~\new_[12461]_  & ~\new_[13020]_ ;
  assign \new_[11382]_  = ~\new_[12466]_  & ~\new_[12938]_ ;
  assign \new_[11383]_  = ~\new_[12459]_  & ~\new_[12999]_ ;
  assign \new_[11384]_  = ~\new_[12379]_  & ~\new_[12881]_ ;
  assign \new_[11385]_  = ~\new_[12379]_  & ~\new_[13046]_ ;
  assign \new_[11386]_  = ~\new_[12812]_  & ~\new_[12923]_ ;
  assign \new_[11387]_  = ~\new_[12355]_  & ~\new_[12939]_ ;
  assign \new_[11388]_  = ~\new_[12374]_  & ~\new_[12937]_ ;
  assign \new_[11389]_  = ~\new_[12812]_  & ~\new_[13046]_ ;
  assign \new_[11390]_  = ~\new_[12355]_  & ~\new_[12998]_ ;
  assign \new_[11391]_  = ~\new_[12374]_  & ~\new_[13041]_ ;
  assign \new_[11392]_  = ~\new_[12445]_  & ~\new_[13004]_ ;
  assign \new_[11393]_  = ~\new_[12850]_  & ~\new_[12910]_ ;
  assign \new_[11394]_  = ~\new_[12850]_  & ~\new_[13043]_ ;
  assign \new_[11395]_  = ~\new_[12449]_  & ~\new_[13004]_ ;
  assign \new_[11396]_  = ~\new_[12444]_  & ~\new_[13053]_ ;
  assign \new_[11397]_  = ~\new_[12461]_  & ~\new_[13041]_ ;
  assign \new_[11398]_  = ~\new_[12371]_  & ~\new_[12937]_ ;
  assign \new_[11399]_  = ~\new_[12428]_  & ~\new_[12939]_ ;
  assign \new_[11400]_  = ~\new_[12443]_  & ~\new_[12936]_ ;
  assign \new_[11401]_  = ~\new_[12442]_  & ~\new_[12938]_ ;
  assign \new_[11402]_  = ~\new_[12371]_  & ~\new_[12910]_ ;
  assign \new_[11403]_  = ~\new_[12443]_  & ~\new_[13026]_ ;
  assign \new_[11404]_  = ~\new_[12812]_  & ~\new_[13008]_ ;
  assign \new_[11405]_  = ~\new_[12743]_  & ~\new_[12739]_ ;
  assign \new_[11406]_  = ~\new_[12371]_  & ~\new_[13043]_ ;
  assign \new_[11407]_  = ~\new_[12442]_  & ~\new_[12897]_ ;
  assign \new_[11408]_  = ~\new_[12743]_  & ~\new_[13054]_ ;
  assign \new_[11409]_  = ~\new_[12445]_  & ~\new_[12941]_ ;
  assign \new_[11410]_  = ~\new_[12355]_  & ~\new_[12941]_ ;
  assign \new_[11411]_  = ~\new_[12743]_  & ~\new_[12881]_ ;
  assign \new_[11412]_  = ~\new_[12812]_  & ~\new_[12739]_ ;
  assign \new_[11413]_  = \new_[13144]_  ^ \new_[12893]_ ;
  assign \new_[11414]_  = \new_[12892]_  ^ \new_[13175]_ ;
  assign \new_[11415]_  = ~\new_[4921]_  | ~\new_[13930]_ ;
  assign \new_[11416]_  = ~\new_[12264]_  | ~\new_[4386]_ ;
  assign \new_[11417]_  = ~\new_[13880]_  | ~\new_[5644]_ ;
  assign \new_[11418]_  = ~\new_[13880]_  | ~\new_[5661]_ ;
  assign \new_[11419]_  = ~\new_[5186]_  | ~\new_[12361]_ ;
  assign \new_[11420]_  = ~\new_[5567]_  | ~\new_[12352]_ ;
  assign \new_[11421]_  = ~\new_[12691]_ ;
  assign \new_[11422]_  = ~\new_[12691]_ ;
  assign \new_[11423]_  = ~\new_[5185]_  | ~\new_[12361]_ ;
  assign \new_[11424]_  = \new_[4851]_  ? \new_[12616]_  : \new_[13136]_ ;
  assign \new_[11425]_  = ~\new_[4910]_  | ~\new_[12431]_ ;
  assign \new_[11426]_  = (~\new_[4073]_  | ~\new_[12594]_ ) & (~\new_[3763]_  | ~\new_[12589]_ );
  assign \new_[11427]_  = ~\new_[12072]_ ;
  assign \new_[11428]_  = ~\new_[12086]_ ;
  assign \new_[11429]_  = \new_[4642]_  ^ \new_[12620]_ ;
  assign \new_[11430]_  = \new_[7973]_  ^ \new_[12506]_ ;
  assign \new_[11431]_  = (~\new_[13678]_  | ~\new_[12560]_ ) & (~\new_[13634]_  | ~\new_[12779]_ );
  assign n10936 = ~\new_[12119]_ ;
  assign \new_[11433]_  = ~\new_[12478]_  | ~\new_[12868]_ ;
  assign \new_[11434]_  = \new_[12868]_  | \new_[12266]_ ;
  assign \new_[11435]_  = \new_[12849]_  | \new_[12407]_ ;
  assign \new_[11436]_  = \new_[12859]_  | \new_[12408]_ ;
  assign \new_[11437]_  = ~\new_[12262]_  | ~\new_[7774]_ ;
  assign \new_[11438]_  = ~\new_[2816]_  | ~\new_[12509]_ ;
  assign \new_[11439]_  = ~\new_[12264]_  | ~\new_[4816]_ ;
  assign \new_[11440]_  = ~\new_[7890]_  | ~\new_[12304]_ ;
  assign \new_[11441]_  = \new_[12885]_  ^ \new_[12571]_ ;
  assign \new_[11442]_  = \new_[12547]_  ^ \new_[12575]_ ;
  assign \new_[11443]_  = ~\new_[12085]_ ;
  assign \new_[11444]_  = ~\new_[12482]_  | ~\wb_addr_i[6] ;
  assign \new_[11445]_  = ~\new_[12482]_  | ~\new_[12483]_ ;
  assign \new_[11446]_  = ~\new_[4911]_  | ~\new_[12341]_ ;
  assign \new_[11447]_  = ~\new_[12680]_  & ~\new_[12679]_ ;
  assign \new_[11448]_  = ~\new_[13972]_  | ~\new_[4846]_ ;
  assign \new_[11449]_  = ~\new_[13726]_  | ~\new_[12907]_  | ~\new_[7979]_  | ~\new_[12600]_ ;
  assign \new_[11450]_  = ~\new_[12485]_  & ~\new_[7977]_ ;
  assign n10926 = ~\new_[13160]_  & ~\new_[12477]_ ;
  assign \new_[11452]_  = ~\new_[12955]_  & (~\new_[12614]_  | ~\new_[13726]_ );
  assign \new_[11453]_  = \new_[13083]_  ^ \new_[12672]_ ;
  assign \new_[11454]_  = ~\new_[7978]_  | ~\new_[13455]_  | ~\new_[12614]_  | ~\new_[12522]_ ;
  assign n10931 = \new_[12503]_  ^ \new_[13139]_ ;
  assign \new_[11456]_  = ~\new_[12348]_  | ~\new_[13084]_ ;
  assign \new_[11457]_  = ~\new_[13058]_  | ~\new_[13538]_  | ~\new_[13125]_ ;
  assign \new_[11458]_  = ~\new_[7889]_  | ~\new_[12304]_ ;
  assign \new_[11459]_  = ~\new_[3760]_  | ~\new_[12304]_ ;
  assign \new_[11460]_  = ~\new_[7792]_  | ~\new_[12304]_ ;
  assign \new_[11461]_  = ~\new_[7891]_  | ~\new_[12304]_ ;
  assign \new_[11462]_  = ~\new_[7893]_  | ~\new_[12509]_ ;
  assign \new_[11463]_  = ~\new_[7925]_  | ~\new_[12509]_ ;
  assign \new_[11464]_  = ~\new_[7894]_  | ~\new_[12509]_ ;
  assign \new_[11465]_  = ~\new_[7793]_  | ~\new_[12509]_ ;
  assign \new_[11466]_  = ~\new_[12304]_  | ~\new_[13112]_ ;
  assign \new_[11467]_  = ~\new_[12348]_  | ~\new_[13058]_ ;
  assign \new_[11468]_  = ~\new_[12291]_  | ~\new_[12975]_ ;
  assign \new_[11469]_  = ~\new_[12527]_  & ~\new_[12594]_ ;
  assign \new_[11470]_  = ~\new_[12510]_  & ~\new_[12679]_ ;
  assign \new_[11471]_  = (~\new_[12997]_  | ~\new_[12644]_ ) & (~\new_[13738]_  | ~\new_[2756]_ );
  assign \new_[11472]_  = (~\new_[12949]_  | ~\new_[12610]_ ) & (~\new_[13794]_  | ~\new_[2758]_ );
  assign \new_[11473]_  = (~\new_[12988]_  | ~\new_[12657]_ ) & (~\new_[13500]_  | ~\new_[2757]_ );
  assign \new_[11474]_  = ~\new_[4945]_  | ~\new_[14181]_ ;
  assign \new_[11475]_  = (~\new_[13766]_  | ~\new_[13076]_ ) & (~\new_[13640]_  | ~\new_[13011]_ );
  assign \new_[11476]_  = (~\new_[4076]_  | ~\new_[12594]_ ) & (~\new_[3186]_  | ~\new_[12589]_ );
  assign \new_[11477]_  = ~\new_[12384]_  | ~\new_[5608]_ ;
  assign \new_[11478]_  = (~\new_[12982]_  | ~\new_[13472]_ ) & (~\new_[13805]_  | ~\new_[12572]_ );
  assign \new_[11479]_  = (~\new_[13273]_  | ~\new_[13076]_ ) & (~\new_[13226]_  | ~\new_[13011]_ );
  assign \new_[11480]_  = (~\new_[13711]_  | ~\new_[13076]_ ) & (~\new_[13215]_  | ~\new_[13011]_ );
  assign \new_[11481]_  = (~\new_[12696]_  | ~\new_[4386]_ ) & (~\new_[12581]_  | ~\new_[4687]_ );
  assign \new_[11482]_  = (~\new_[12982]_  | ~\new_[13488]_ ) & (~\new_[13429]_  | ~\new_[12572]_ );
  assign \new_[11483]_  = (~\new_[13676]_  | ~\new_[13001]_ ) & (~\new_[13363]_  | ~\new_[13011]_ );
  assign \new_[11484]_  = ~\new_[12399]_  | ~\new_[2727]_ ;
  assign \new_[11485]_  = (~\new_[13535]_  | ~\new_[12560]_ ) & (~\new_[13293]_  | ~\new_[12779]_ );
  assign \new_[11486]_  = (~\new_[13576]_  | ~\new_[12560]_ ) & (~\new_[13450]_  | ~\new_[12572]_ );
  assign \new_[11487]_  = (~\new_[12982]_  | ~\new_[13288]_ ) & (~\new_[13438]_  | ~\new_[13001]_ );
  assign \new_[11488]_  = (~\new_[13826]_  | ~\new_[13076]_ ) & (~\new_[13560]_  | ~\new_[13011]_ );
  assign \new_[11489]_  = (~\new_[13397]_  | ~\new_[12560]_ ) & (~\new_[13722]_  | ~\new_[12572]_ );
  assign \new_[11490]_  = (~\new_[12982]_  | ~\new_[13355]_ ) & (~\new_[13750]_  | ~\new_[12572]_ );
  assign \new_[11491]_  = (~\new_[3780]_  | ~\new_[12618]_ ) & (~\new_[12696]_  | ~\new_[4584]_ );
  assign \new_[11492]_  = (~\new_[13784]_  | ~\new_[12560]_ ) & (~\new_[13858]_  | ~\new_[12779]_ );
  assign \new_[11493]_  = (~\new_[13195]_  | ~\new_[12560]_ ) & (~\new_[13553]_  | ~\new_[12572]_ );
  assign \new_[11494]_  = (~\new_[13513]_  | ~\new_[12560]_ ) & (~\new_[13240]_  | ~\new_[12779]_ );
  assign \new_[11495]_  = (~\new_[13653]_  | ~\new_[12560]_ ) & (~\new_[13340]_  | ~\new_[12779]_ );
  assign \new_[11496]_  = (~\new_[12982]_  | ~\new_[13213]_ ) & (~\new_[13414]_  | ~\new_[12572]_ );
  assign \new_[11497]_  = (~\new_[12982]_  | ~\new_[13795]_ ) & (~\new_[13263]_  | ~\new_[12572]_ );
  assign \new_[11498]_  = (~\new_[12982]_  | ~\new_[13793]_ ) & (~\new_[13759]_  | ~\new_[13001]_ );
  assign \new_[11499]_  = (~\new_[13241]_  | ~\new_[13076]_ ) & (~\new_[13856]_  | ~\new_[13011]_ );
  assign \new_[11500]_  = (~\new_[12581]_  | ~\new_[2726]_ ) & (~\new_[12618]_  | ~\new_[6794]_ );
  assign \new_[11501]_  = (~\new_[3783]_  | ~\new_[12618]_ ) & (~\new_[12696]_  | ~\new_[7932]_ );
  assign \new_[11502]_  = (~\new_[12696]_  | ~\new_[2726]_ ) & (~\new_[12581]_  | ~\new_[2748]_ );
  assign \new_[11503]_  = (~\new_[12696]_  | ~\new_[2717]_ ) & (~\new_[12581]_  | ~\new_[2737]_ );
  assign \new_[11504]_  = (~\new_[12667]_  | ~\new_[2727]_ ) & (~\new_[12586]_  | ~\new_[2749]_ );
  assign \new_[11505]_  = (~\new_[12667]_  | ~\new_[2718]_ ) & (~\new_[12586]_  | ~\new_[2738]_ );
  assign \new_[11506]_  = (~\new_[12586]_  | ~\new_[2727]_ ) & (~\new_[12679]_  | ~\new_[6809]_ );
  assign \new_[11507]_  = (~\new_[12586]_  | ~\new_[2718]_ ) & (~\new_[12679]_  | ~\new_[5888]_ );
  assign \new_[11508]_  = (~\new_[12581]_  | ~\new_[2717]_ ) & (~\new_[12618]_  | ~\new_[5855]_ );
  assign \new_[11509]_  = (~\new_[3776]_  | ~\new_[12618]_ ) & (~\new_[12696]_  | ~\new_[7928]_ );
  assign \new_[11510]_  = (~\new_[13446]_  | ~\new_[13001]_ ) & (~\new_[13267]_  | ~\new_[13011]_ );
  assign \new_[11511]_  = ~\new_[5032]_  | ~\new_[12553]_ ;
  assign \new_[11512]_  = (~\new_[12778]_  | ~\new_[13503]_ ) & (~\new_[13364]_  | ~\new_[12805]_ );
  assign \new_[11513]_  = (~\new_[13292]_  | ~\new_[12763]_ ) & (~\new_[13309]_  | ~\new_[13023]_ );
  assign \new_[11514]_  = (~\new_[12982]_  | ~\new_[13831]_ ) & (~\new_[13470]_  | ~\new_[12747]_ );
  assign \new_[11515]_  = (~\new_[12778]_  | ~\new_[13497]_ ) & (~\new_[13717]_  | ~\new_[12805]_ );
  assign \new_[11516]_  = (~\new_[12778]_  | ~\new_[13659]_ ) & (~\new_[13229]_  | ~\new_[12763]_ );
  assign \new_[11517]_  = (~\new_[12778]_  | ~\new_[13862]_ ) & (~\new_[13453]_  | ~\new_[12805]_ );
  assign \new_[11518]_  = ~\new_[5334]_  | ~\new_[14188]_ ;
  assign \new_[11519]_  = ~\new_[5758]_  | ~\new_[14188]_ ;
  assign \new_[11520]_  = ~\new_[12608]_  | ~\new_[4857]_ ;
  assign \new_[11521]_  = ~\new_[5732]_  | ~\new_[14188]_ ;
  assign \new_[11522]_  = ~\new_[12635]_  | ~\new_[4849]_ ;
  assign \new_[11523]_  = ~\new_[12361]_ ;
  assign \new_[11524]_  = \new_[13461]_  ^ \new_[13102]_ ;
  assign \new_[11525]_  = \new_[3150]_  ^ \new_[12780]_ ;
  assign \new_[11526]_  = ~\new_[12687]_  & ~\new_[12935]_ ;
  assign \new_[11527]_  = ~\new_[12678]_  & ~\new_[12913]_ ;
  assign \new_[11528]_  = \\u15_crac_din_reg[6] ;
  assign \new_[11529]_  = ~\new_[5418]_  | ~\new_[12585]_ ;
  assign \new_[11530]_  = ~\new_[12678]_  & ~\new_[13034]_ ;
  assign \new_[11531]_  = ~\new_[12608]_  | ~\new_[5636]_ ;
  assign \new_[11532]_  = ~\new_[12727]_  | ~\new_[2793]_ ;
  assign \new_[11533]_  = ~\new_[12687]_  & ~\new_[12739]_ ;
  assign \new_[11534]_  = ~\new_[12948]_  & ~\new_[13026]_ ;
  assign \new_[11535]_  = ~\new_[3250]_  & ~\new_[12707]_ ;
  assign \new_[11536]_  = ~\new_[5575]_  | ~\new_[12554]_ ;
  assign \new_[11537]_  = ~\new_[12608]_  | ~\new_[5638]_ ;
  assign \new_[11538]_  = ~\new_[12586]_  | ~\new_[7879]_ ;
  assign \new_[11539]_  = ~\new_[12678]_  & ~\new_[12739]_ ;
  assign \new_[11540]_  = ~\new_[5169]_  | ~\new_[12644]_ ;
  assign \new_[11541]_  = ~\new_[5201]_  | ~\new_[12657]_ ;
  assign \new_[11542]_  = ~\new_[5432]_  | ~\new_[12610]_ ;
  assign \new_[11543]_  = ~\new_[4976]_  | ~\new_[12657]_ ;
  assign \new_[11544]_  = ~\new_[5438]_  | ~\new_[12610]_ ;
  assign \new_[11545]_  = ~\new_[5220]_  | ~\new_[12657]_ ;
  assign \new_[11546]_  = ~\new_[5160]_  | ~\new_[12644]_ ;
  assign \new_[11547]_  = ~\new_[5210]_  | ~\new_[12657]_ ;
  assign \new_[11548]_  = ~\new_[5436]_  | ~\new_[12610]_ ;
  assign \new_[11549]_  = ~\new_[5018]_  | ~\new_[12644]_ ;
  assign \new_[11550]_  = ~\new_[5215]_  | ~\new_[12657]_ ;
  assign \new_[11551]_  = ~\new_[5001]_  | ~\new_[12644]_ ;
  assign \new_[11552]_  = ~\new_[5005]_  | ~\new_[12644]_ ;
  assign \new_[11553]_  = ~\new_[5423]_  | ~\new_[14118]_ ;
  assign \new_[11554]_  = ~\new_[5219]_  | ~\new_[12657]_ ;
  assign \new_[11555]_  = ~\new_[5433]_  | ~\new_[12610]_ ;
  assign \new_[11556]_  = ~\new_[5690]_  | ~\new_[12593]_ ;
  assign \new_[11557]_  = ~\new_[5209]_  | ~\new_[12657]_ ;
  assign \new_[11558]_  = ~\new_[5010]_  | ~\new_[12644]_ ;
  assign \new_[11559]_  = ~\new_[5359]_  | ~\new_[12396]_ ;
  assign \new_[11560]_  = ~\new_[5737]_  | ~\new_[12396]_ ;
  assign \new_[11561]_  = ~\new_[5208]_  | ~\new_[12657]_ ;
  assign \new_[11562]_  = ~\new_[5674]_  | ~\new_[12610]_ ;
  assign \new_[11563]_  = ~\new_[5736]_  | ~\new_[12396]_ ;
  assign \new_[11564]_  = ~\new_[5367]_  | ~\new_[12396]_ ;
  assign \new_[11565]_  = ~\new_[4977]_  | ~\new_[12657]_ ;
  assign \new_[11566]_  = ~\new_[5155]_  | ~\new_[12644]_ ;
  assign \new_[11567]_  = ~\new_[5153]_  | ~\new_[12644]_ ;
  assign \new_[11568]_  = ~\new_[4975]_  | ~\new_[12657]_ ;
  assign \new_[11569]_  = ~\new_[5421]_  | ~\new_[12593]_ ;
  assign \new_[11570]_  = ~\new_[5675]_  | ~\new_[12610]_ ;
  assign \new_[11571]_  = ~\new_[5035]_  | ~\new_[12593]_ ;
  assign \new_[11572]_  = ~\new_[5443]_  | ~\new_[12593]_ ;
  assign \new_[11573]_  = ~\new_[5434]_  | ~\new_[12610]_ ;
  assign \new_[11574]_  = ~\new_[5424]_  | ~\new_[12593]_ ;
  assign \new_[11575]_  = ~\new_[5676]_  | ~\new_[12593]_ ;
  assign \new_[11576]_  = ~\new_[5437]_  | ~\new_[12610]_ ;
  assign \new_[11577]_  = ~\new_[5427]_  | ~\new_[12593]_ ;
  assign \new_[11578]_  = ~\new_[5439]_  | ~\new_[12610]_ ;
  assign \new_[11579]_  = ~\new_[5678]_  | ~\new_[12593]_ ;
  assign \new_[11580]_  = ~\new_[5429]_  | ~\new_[14118]_ ;
  assign \new_[11581]_  = ~\new_[5672]_  | ~\new_[14118]_ ;
  assign \new_[11582]_  = ~\new_[5670]_  | ~\new_[12593]_ ;
  assign \new_[11583]_  = \new_[13217]_  | \new_[12679]_ ;
  assign \new_[11584]_  = ~\new_[5430]_  | ~\new_[12610]_ ;
  assign \new_[11585]_  = ~\new_[5007]_  | ~\new_[12644]_ ;
  assign \new_[11586]_  = ~\new_[5207]_  | ~\new_[12657]_ ;
  assign \new_[11587]_  = ~\new_[5355]_  | ~\new_[12396]_ ;
  assign \new_[11588]_  = ~\new_[5428]_  | ~\new_[12593]_ ;
  assign \new_[11589]_  = ~\new_[5352]_  | ~\new_[12396]_ ;
  assign \new_[11590]_  = ~\new_[5205]_  | ~\new_[12657]_ ;
  assign \new_[11591]_  = ~\new_[5740]_  | ~\new_[12396]_ ;
  assign \new_[11592]_  = ~\new_[5431]_  | ~\new_[12610]_ ;
  assign \new_[11593]_  = ~\new_[5445]_  | ~\new_[12657]_ ;
  assign \new_[11594]_  = ~\new_[5361]_  | ~\new_[12396]_ ;
  assign \new_[11595]_  = ~\new_[5167]_  | ~\new_[12644]_ ;
  assign \new_[11596]_  = ~\new_[5150]_  | ~\new_[12644]_ ;
  assign \new_[11597]_  = ~\new_[12596]_  | ~\new_[7973]_ ;
  assign \new_[11598]_  = ~\new_[5441]_  | ~\new_[14118]_ ;
  assign \new_[11599]_  = ~\new_[4992]_  | ~\new_[12657]_ ;
  assign \new_[11600]_  = ~\new_[5211]_  | ~\new_[12657]_ ;
  assign \new_[11601]_  = ~\new_[5142]_  | ~\new_[12644]_ ;
  assign \new_[11602]_  = ~\new_[5176]_  | ~\new_[12644]_ ;
  assign \new_[11603]_  = ~\new_[4979]_  | ~\new_[12657]_ ;
  assign \new_[11604]_  = ~\new_[5146]_  | ~\new_[12644]_ ;
  assign \new_[11605]_  = ~\new_[5147]_  | ~\new_[12644]_ ;
  assign \new_[11606]_  = ~\new_[5165]_  | ~\new_[12644]_ ;
  assign \new_[11607]_  = ~\new_[5435]_  | ~\new_[12610]_ ;
  assign \new_[11608]_  = ~\new_[5017]_  | ~\new_[12644]_ ;
  assign \new_[11609]_  = ~\new_[5151]_  | ~\new_[12644]_ ;
  assign \new_[11610]_  = ~\new_[5170]_  | ~\new_[12644]_ ;
  assign \new_[11611]_  = ~\new_[5168]_  | ~\new_[12644]_ ;
  assign \new_[11612]_  = ~\new_[5011]_  | ~\new_[12644]_ ;
  assign \new_[11613]_  = ~\new_[5172]_  | ~\new_[12644]_ ;
  assign \new_[11614]_  = ~\new_[5174]_  | ~\new_[12644]_ ;
  assign \new_[11615]_  = ~\new_[5157]_  | ~\new_[12644]_ ;
  assign \new_[11616]_  = ~\new_[5212]_  | ~\new_[12657]_ ;
  assign \new_[11617]_  = ~\new_[7978]_  & ~\new_[12596]_ ;
  assign \new_[11618]_  = ~\new_[5440]_  | ~\new_[14118]_ ;
  assign \new_[11619]_  = ~\new_[5161]_  | ~\new_[12644]_ ;
  assign \new_[11620]_  = ~\new_[5158]_  | ~\new_[12644]_ ;
  assign \new_[11621]_  = ~\new_[5144]_  | ~\new_[12644]_ ;
  assign \new_[11622]_  = ~\new_[12645]_  & ~\new_[13034]_ ;
  assign \new_[11623]_  = \new_[13756]_  | \new_[12594]_ ;
  assign \new_[11624]_  = ~\new_[5178]_  | ~\new_[12644]_ ;
  assign \new_[11625]_  = ~\new_[12644]_  | ~\new_[13857]_ ;
  assign \new_[11626]_  = ~\new_[4817]_  | ~\new_[12594]_ ;
  assign \new_[11627]_  = ~\new_[5572]_  | ~\new_[12554]_ ;
  assign \new_[11628]_  = ~\new_[3530]_  & ~\new_[12707]_ ;
  assign \new_[11629]_  = ~\new_[5139]_  | ~\new_[12553]_ ;
  assign \new_[11630]_  = ~\new_[5326]_  | ~\new_[14188]_ ;
  assign \new_[11631]_  = ~\new_[12610]_  | ~\new_[13532]_ ;
  assign \new_[11632]_  = ~\new_[12581]_  | ~\new_[7877]_ ;
  assign \new_[11633]_  = ~\new_[12581]_  | ~\new_[4386]_ ;
  assign \new_[11634]_  = ~\new_[5270]_  | ~\new_[13930]_ ;
  assign \new_[11635]_  = ~\new_[7686]_  | ~\new_[12594]_ ;
  assign \new_[11636]_  = ~\new_[5551]_  | ~\new_[12553]_ ;
  assign \new_[11637]_  = ~\new_[4896]_  | ~\new_[12554]_ ;
  assign \new_[11638]_  = ~\new_[13042]_  & ~\new_[12550]_ ;
  assign \new_[11639]_  = ~\new_[5252]_  | ~\new_[13930]_ ;
  assign \new_[11640]_  = ~\new_[5254]_  | ~\new_[13930]_ ;
  assign \new_[11641]_  = ~\new_[2725]_  | ~\new_[12594]_ ;
  assign \new_[11642]_  = ~\new_[3412]_  & ~\new_[12707]_ ;
  assign \new_[11643]_  = ~\new_[12581]_  | ~\new_[2789]_ ;
  assign \new_[11644]_  = ~\new_[5343]_  | ~\new_[14188]_ ;
  assign \new_[11645]_  = ~\new_[3248]_  & ~\new_[12707]_ ;
  assign \new_[11646]_  = ~\new_[5752]_  | ~\new_[14188]_ ;
  assign \new_[11647]_  = ~\new_[5140]_  | ~\new_[12553]_ ;
  assign \new_[11648]_  = ~\new_[5346]_  | ~\new_[14188]_ ;
  assign \new_[11649]_  = ~\new_[3411]_  & ~\new_[12707]_ ;
  assign \new_[11650]_  = ~\new_[3259]_  & ~\new_[12707]_ ;
  assign \new_[11651]_  = ~\new_[12581]_  | ~\new_[6794]_ ;
  assign \new_[11652]_  = ~\new_[12608]_  | ~\new_[5008]_ ;
  assign \new_[11653]_  = ~\new_[3251]_  & ~\new_[12707]_ ;
  assign \new_[11654]_  = ~\new_[12635]_  | ~\new_[5627]_ ;
  assign \new_[11655]_  = ~\new_[12586]_  | ~\new_[7926]_ ;
  assign \new_[11656]_  = ~\new_[3252]_  & ~\new_[12707]_ ;
  assign \new_[11657]_  = ~\new_[12586]_  | ~\new_[7878]_ ;
  assign \new_[11658]_  = ~\new_[5322]_  | ~\new_[14188]_ ;
  assign \new_[11659]_  = ~\new_[5323]_  | ~\new_[14188]_ ;
  assign \new_[11660]_  = ~\new_[5345]_  | ~\new_[14188]_ ;
  assign \new_[11661]_  = ~\new_[12635]_  | ~\new_[5629]_ ;
  assign \new_[11662]_  = ~\new_[5333]_  | ~\new_[14188]_ ;
  assign \new_[11663]_  = ~\new_[12556]_  & ~\new_[12884]_ ;
  assign \new_[11664]_  = ~\new_[5324]_  | ~\new_[14188]_ ;
  assign \new_[11665]_  = ~\new_[5335]_  | ~\new_[14188]_ ;
  assign \new_[11666]_  = ~\new_[5754]_  | ~\new_[14188]_ ;
  assign \new_[11667]_  = ~\new_[5762]_  | ~\new_[14188]_ ;
  assign \new_[11668]_  = ~\new_[5264]_  | ~\new_[13930]_ ;
  assign \new_[11669]_  = ~\new_[5338]_  | ~\new_[14188]_ ;
  assign \new_[11670]_  = ~\new_[5328]_  | ~\new_[14188]_ ;
  assign \new_[11671]_  = ~\new_[5330]_  | ~\new_[14188]_ ;
  assign \new_[11672]_  = ~\new_[5341]_  | ~\new_[14188]_ ;
  assign \new_[11673]_  = ~\new_[12618]_  | ~\new_[2748]_ ;
  assign \new_[11674]_  = ~\new_[3249]_  & ~\new_[12707]_ ;
  assign \new_[11675]_  = ~\new_[5342]_  | ~\new_[14188]_ ;
  assign \new_[11676]_  = ~\new_[12581]_  | ~\new_[7501]_ ;
  assign \new_[11677]_  = ~\new_[5266]_  | ~\new_[13930]_ ;
  assign \new_[11678]_  = ~\new_[3781]_  | ~\new_[12618]_ ;
  assign \new_[11679]_  = ~\new_[12651]_  | ~\new_[2759]_ ;
  assign \new_[11680]_  = ~\new_[4898]_  | ~\new_[12554]_ ;
  assign \new_[11681]_  = \new_[12650]_  | \new_[13738]_ ;
  assign \new_[11682]_  = ~\new_[5552]_  | ~\new_[12553]_ ;
  assign \new_[11683]_  = \new_[14103]_  | \new_[13425]_ ;
  assign \new_[11684]_  = ~\new_[5332]_  | ~\new_[14188]_ ;
  assign \new_[11685]_  = ~\new_[12586]_  | ~\new_[7503]_ ;
  assign \new_[11686]_  = ~\new_[5137]_  | ~\new_[12553]_ ;
  assign \new_[11687]_  = ~\new_[12635]_  | ~\new_[4994]_ ;
  assign \new_[11688]_  = ~\new_[2785]_  | ~\new_[12594]_ ;
  assign \new_[11689]_  = ~\new_[12999]_  & ~\new_[12568]_ ;
  assign \new_[11690]_  = ~\new_[12635]_  | ~\new_[5626]_ ;
  assign \new_[11691]_  = ~\new_[12581]_  | ~\new_[7932]_ ;
  assign \new_[11692]_  = ~\new_[12608]_  | ~\new_[5637]_ ;
  assign \new_[11693]_  = ~\new_[12586]_  | ~\new_[2924]_ ;
  assign \new_[11694]_  = ~\new_[5561]_  | ~\new_[12554]_ ;
  assign \new_[11695]_  = ~\new_[5691]_  | ~\new_[12585]_ ;
  assign \new_[11696]_  = ~\new_[3186]_  | ~\new_[12594]_ ;
  assign \new_[11697]_  = ~\new_[12481]_ ;
  assign \new_[11698]_  = ~\new_[2716]_  | ~\new_[12594]_ ;
  assign \new_[11699]_  = ~\new_[5714]_  | ~\new_[12585]_ ;
  assign \new_[11700]_  = ~\new_[12635]_  | ~\new_[5625]_ ;
  assign \new_[11701]_  = ~\new_[12581]_  | ~\new_[4584]_ ;
  assign \new_[11702]_  = ~\new_[12586]_  | ~\new_[4410]_ ;
  assign \new_[11703]_  = ~\new_[5400]_  | ~\new_[12585]_ ;
  assign \new_[11704]_  = ~\new_[5255]_  | ~\new_[13931]_ ;
  assign \new_[11705]_  = ~\new_[12618]_  | ~\new_[2789]_ ;
  assign \new_[11706]_  = ~\new_[4585]_  | ~\new_[12594]_ ;
  assign \new_[11707]_  = ~\new_[5689]_  | ~\new_[12585]_ ;
  assign \new_[11708]_  = ~\new_[5327]_  | ~\new_[14188]_ ;
  assign \new_[11709]_  = ~\new_[5404]_  | ~\new_[12585]_ ;
  assign \new_[11710]_  = \\u15_crac_din_reg[9] ;
  assign \new_[11711]_  = ~\new_[12586]_  | ~\new_[7927]_ ;
  assign \new_[11712]_  = ~\new_[5417]_  | ~\new_[12585]_ ;
  assign \new_[11713]_  = \new_[12629]_  | \new_[13794]_ ;
  assign \new_[11714]_  = ~\new_[12581]_  | ~\new_[2923]_ ;
  assign \new_[11715]_  = ~\new_[12586]_  | ~\new_[4576]_ ;
  assign \new_[11716]_  = ~\new_[12618]_  | ~\new_[7687]_ ;
  assign \new_[11717]_  = ~\new_[5704]_  | ~\new_[12585]_ ;
  assign \new_[11718]_  = ~\new_[12576]_  & ~\new_[12738]_ ;
  assign \new_[11719]_  = ~\new_[12618]_  | ~\new_[7501]_ ;
  assign \new_[11720]_  = ~\new_[5253]_  | ~\new_[13930]_ ;
  assign \new_[11721]_  = ~\new_[12886]_ ;
  assign \new_[11722]_  = ~\new_[12618]_  | ~\new_[2923]_ ;
  assign \new_[11723]_  = ~\new_[7502]_  | ~\new_[12594]_ ;
  assign \new_[11724]_  = ~\new_[5337]_  | ~\new_[14188]_ ;
  assign \new_[11725]_  = ~\new_[3529]_  & ~\new_[12707]_ ;
  assign \new_[11726]_  = ~\new_[5692]_  | ~\new_[12585]_ ;
  assign \new_[11727]_  = ~\new_[12618]_  | ~\new_[4687]_ ;
  assign \new_[11728]_  = ~\new_[4071]_  | ~\new_[12594]_ ;
  assign \new_[11729]_  = ~\new_[5344]_  | ~\new_[14188]_ ;
  assign \new_[11730]_  = ~\new_[5559]_  | ~\new_[12553]_ ;
  assign \new_[11731]_  = ~\new_[12586]_  | ~\new_[6809]_ ;
  assign \new_[11732]_  = ~\new_[12586]_  | ~\new_[7688]_ ;
  assign \new_[11733]_  = ~\new_[5761]_  | ~\new_[14188]_ ;
  assign \new_[11734]_  = ~\new_[12586]_  | ~\new_[5888]_ ;
  assign \new_[11735]_  = ~\new_[12586]_  | ~\new_[4813]_ ;
  assign \new_[11736]_  = ~\new_[12608]_  | ~\new_[5628]_ ;
  assign \new_[11737]_  = ~\new_[4900]_  | ~\new_[13931]_ ;
  assign \new_[11738]_  = ~\new_[5549]_  | ~\new_[12553]_ ;
  assign \new_[11739]_  = ~\new_[5566]_  | ~\new_[12554]_ ;
  assign \new_[11740]_  = ~\new_[5760]_  | ~\new_[14188]_ ;
  assign \new_[11741]_  = ~\new_[5325]_  | ~\new_[14188]_ ;
  assign \new_[11742]_  = ~\new_[12581]_  | ~\new_[3764]_ ;
  assign \new_[11743]_  = ~\new_[12581]_  | ~\new_[7687]_ ;
  assign \new_[11744]_  = ~\new_[12581]_  | ~\new_[4816]_ ;
  assign \new_[11745]_  = ~\new_[12586]_  | ~\new_[2787]_ ;
  assign \new_[11746]_  = ~\new_[5557]_  | ~\new_[12553]_ ;
  assign \new_[11747]_  = ~\new_[3763]_  | ~\new_[12594]_ ;
  assign \new_[11748]_  = ~\new_[12581]_  | ~\new_[7933]_ ;
  assign \new_[11749]_  = ~\new_[4688]_  | ~\new_[12594]_ ;
  assign \new_[11750]_  = ~\new_[5336]_  | ~\new_[14188]_ ;
  assign \new_[11751]_  = ~\new_[12697]_  & ~\new_[13043]_ ;
  assign \new_[11752]_  = ~\new_[5269]_  | ~\new_[13931]_ ;
  assign \new_[11753]_  = \new_[12599]_  | \new_[13500]_ ;
  assign \new_[11754]_  = ~\new_[5339]_  | ~\new_[14188]_ ;
  assign \new_[11755]_  = ~\new_[5554]_  | ~\new_[12554]_ ;
  assign \new_[11756]_  = ~\new_[5397]_  | ~\new_[12585]_ ;
  assign \new_[11757]_  = ~\new_[12586]_  | ~\new_[3185]_ ;
  assign \new_[11758]_  = ~\new_[12948]_  & ~\new_[13043]_ ;
  assign \new_[11759]_  = ~\new_[12948]_  & ~\new_[13042]_ ;
  assign \new_[11760]_  = ~\new_[13064]_  & ~\new_[13053]_ ;
  assign \new_[11761]_  = ~\new_[12555]_  & ~\new_[12905]_ ;
  assign \new_[11762]_  = ~\new_[12561]_  & ~\new_[12739]_ ;
  assign \new_[11763]_  = ~\new_[12948]_  & ~\new_[13003]_ ;
  assign \new_[11764]_  = ~\new_[12555]_  & ~\new_[13041]_ ;
  assign \new_[11765]_  = ~\new_[12561]_  & ~\new_[12738]_ ;
  assign \new_[11766]_  = ~\new_[12923]_  & ~\new_[12550]_ ;
  assign \new_[11767]_  = ~\new_[13008]_  & ~\new_[12550]_ ;
  assign \new_[11768]_  = ~\new_[12555]_  & ~\new_[13020]_ ;
  assign \new_[11769]_  = ~\new_[12557]_  & ~\new_[13053]_ ;
  assign \new_[11770]_  = ~\new_[12624]_  & ~\new_[13046]_ ;
  assign \new_[11771]_  = ~\new_[12687]_  & ~\new_[12938]_ ;
  assign \new_[11772]_  = ~\new_[13050]_  & ~\new_[13053]_ ;
  assign \new_[11773]_  = ~\new_[12678]_  & ~\new_[12897]_ ;
  assign \new_[11774]_  = ~\new_[12690]_  & ~\new_[12913]_ ;
  assign \new_[11775]_  = ~\new_[12687]_  & ~\new_[12937]_ ;
  assign \new_[11776]_  = ~\new_[12561]_  & ~\new_[12934]_ ;
  assign \new_[11777]_  = ~\new_[12563]_  & ~\new_[12937]_ ;
  assign \new_[11778]_  = ~\new_[12989]_  & ~\new_[12550]_ ;
  assign \new_[11779]_  = ~\new_[12884]_  & ~\new_[12568]_ ;
  assign \new_[11780]_  = ~\new_[12608]_  | ~\new_[4850]_ ;
  assign \new_[11781]_  = ~\new_[12561]_  & ~\new_[12910]_ ;
  assign \new_[11782]_  = ~\new_[12948]_  & ~\new_[12998]_ ;
  assign \new_[11783]_  = ~\new_[12679]_  | ~\new_[7503]_ ;
  assign \new_[11784]_  = ~\new_[12938]_  & ~\new_[12568]_ ;
  assign \new_[11785]_  = ~\new_[13064]_  & ~\new_[12905]_ ;
  assign \new_[11786]_  = ~\new_[13034]_  & ~\new_[12550]_ ;
  assign \new_[11787]_  = ~\new_[12935]_  & ~\new_[12621]_ ;
  assign \new_[11788]_  = ~\new_[13064]_  & ~\new_[12936]_ ;
  assign \new_[11789]_  = ~\new_[12697]_  & ~\new_[12923]_ ;
  assign \new_[11790]_  = ~\new_[13066]_  & ~\new_[12998]_ ;
  assign \new_[11791]_  = ~\new_[12703]_  & ~\new_[12910]_ ;
  assign \new_[11792]_  = ~\new_[12546]_  & ~\new_[12998]_ ;
  assign \new_[11793]_  = ~\new_[12678]_  & ~\new_[12939]_ ;
  assign \new_[11794]_  = ~\new_[13026]_  & ~\new_[12621]_ ;
  assign \new_[11795]_  = ~\new_[12543]_  & ~\new_[13026]_ ;
  assign \new_[11796]_  = ~\new_[12678]_  & ~\new_[12999]_ ;
  assign \new_[11797]_  = ~\new_[12559]_  & ~\new_[12938]_ ;
  assign \new_[11798]_  = ~\new_[12569]_  & ~\new_[12937]_ ;
  assign \new_[11799]_  = ~\new_[13053]_  & ~\new_[12597]_ ;
  assign \new_[11800]_  = ~\new_[12577]_  | ~\new_[12756]_ ;
  assign \new_[11801]_  = ~\new_[13034]_  & ~\new_[12621]_ ;
  assign \new_[11802]_  = ~\new_[13081]_  & ~\new_[12897]_ ;
  assign \new_[11803]_  = ~\new_[12624]_  & ~\new_[12739]_ ;
  assign \new_[11804]_  = ~\new_[12690]_  & ~\new_[12999]_ ;
  assign \new_[11805]_  = ~\new_[12564]_  & ~\new_[12923]_ ;
  assign \new_[11806]_  = ~\new_[12948]_  & ~\new_[12923]_ ;
  assign \new_[11807]_  = ~\new_[12934]_  & ~\new_[12568]_ ;
  assign \new_[11808]_  = ~\new_[12936]_  & ~\new_[12568]_ ;
  assign \new_[11809]_  = ~\new_[12558]_  & ~\new_[13004]_ ;
  assign \new_[11810]_  = ~\new_[12678]_  & ~\new_[12884]_ ;
  assign \new_[11811]_  = ~\new_[13054]_  & ~\new_[12568]_ ;
  assign \new_[11812]_  = ~\new_[12739]_  & ~\new_[12568]_ ;
  assign \new_[11813]_  = ~\new_[12582]_  | ~\new_[12759]_ ;
  assign \new_[11814]_  = ~\new_[12935]_  & ~\new_[12525]_ ;
  assign \new_[11815]_  = ~\new_[12556]_  & ~\new_[12941]_ ;
  assign \new_[11816]_  = ~\new_[12923]_  & ~\new_[12568]_ ;
  assign \new_[11817]_  = ~\new_[12625]_  & ~\new_[12913]_ ;
  assign \new_[11818]_  = ~\new_[13050]_  & ~\new_[13043]_ ;
  assign \new_[11819]_  = ~\new_[12913]_  & ~\new_[12568]_ ;
  assign \new_[11820]_  = ~\new_[13064]_  & ~\new_[12910]_ ;
  assign \new_[11821]_  = ~\new_[13050]_  & ~\new_[12905]_ ;
  assign \new_[11822]_  = ~\new_[12703]_  & ~\new_[13042]_ ;
  assign \new_[11823]_  = ~\new_[12897]_  & ~\new_[12568]_ ;
  assign \new_[11824]_  = ~\new_[12678]_  & ~\new_[12881]_ ;
  assign \new_[11825]_  = ~\new_[13064]_  & ~\new_[13034]_ ;
  assign \new_[11826]_  = ~\new_[12678]_  & ~\new_[12937]_ ;
  assign \new_[11827]_  = ~\new_[12738]_  & ~\new_[12597]_ ;
  assign \new_[11828]_  = ~\new_[12557]_  & ~\new_[13003]_ ;
  assign \new_[11829]_  = ~\new_[12625]_  & ~\new_[12934]_ ;
  assign \new_[11830]_  = ~\new_[12570]_  & ~\new_[13020]_ ;
  assign \new_[11831]_  = ~\new_[12567]_  & ~\new_[12913]_ ;
  assign \new_[11832]_  = ~\new_[12566]_  & ~\new_[12937]_ ;
  assign \new_[11833]_  = ~\new_[12690]_  & ~\new_[12897]_ ;
  assign \new_[11834]_  = ~\new_[5556]_  | ~\new_[12553]_ ;
  assign \new_[11835]_  = ~\new_[12565]_  & ~\new_[13003]_ ;
  assign \new_[11836]_  = ~\new_[12948]_  & ~\new_[12738]_ ;
  assign \new_[11837]_  = ~\new_[12881]_  & ~\new_[12550]_ ;
  assign \new_[11838]_  = ~\new_[12678]_  & ~\new_[13042]_ ;
  assign \new_[11839]_  = ~\new_[12884]_  & ~\new_[12552]_ ;
  assign \new_[11840]_  = ~\new_[12565]_  & ~\new_[13041]_ ;
  assign \new_[11841]_  = ~\new_[12999]_  & ~\new_[12552]_ ;
  assign \new_[11842]_  = ~\new_[12628]_  & ~\new_[12989]_ ;
  assign \new_[11843]_  = ~\new_[12678]_  & ~\new_[13046]_ ;
  assign \new_[11844]_  = ~\new_[12678]_  & ~\new_[13041]_ ;
  assign \new_[11845]_  = ~\new_[12631]_  & ~\new_[12939]_ ;
  assign \new_[11846]_  = ~\new_[12678]_  & ~\new_[12935]_ ;
  assign \new_[11847]_  = ~\new_[12687]_  & ~\new_[13060]_ ;
  assign \new_[11848]_  = ~\new_[12687]_  & ~\new_[12923]_ ;
  assign \new_[11849]_  = ~\new_[12678]_  & ~\new_[12934]_ ;
  assign \new_[11850]_  = ~\new_[12573]_  & ~\new_[13042]_ ;
  assign \new_[11851]_  = ~\new_[12678]_  & ~\new_[12938]_ ;
  assign \new_[11852]_  = ~\new_[12687]_  & ~\new_[13046]_ ;
  assign \new_[11853]_  = ~\new_[13064]_  & ~\new_[13046]_ ;
  assign \new_[11854]_  = ~\new_[12628]_  & ~\new_[13041]_ ;
  assign \new_[11855]_  = ~\new_[12687]_  & ~\new_[13043]_ ;
  assign \new_[11856]_  = ~\new_[12645]_  & ~\new_[12941]_ ;
  assign \new_[11857]_  = ~\new_[13041]_  & ~\new_[12950]_ ;
  assign \new_[11858]_  = ~\new_[12567]_  & ~\new_[12999]_ ;
  assign \new_[11859]_  = ~\new_[13066]_  & ~\new_[13054]_ ;
  assign \new_[11860]_  = ~\new_[12559]_  & ~\new_[12934]_ ;
  assign \new_[11861]_  = ~\new_[13046]_  & ~\new_[12597]_ ;
  assign \new_[11862]_  = ~\new_[13046]_  & ~\new_[12550]_ ;
  assign \new_[11863]_  = ~\new_[13081]_  & ~\new_[13026]_ ;
  assign \new_[11864]_  = ~\new_[12908]_  & ~\new_[12881]_ ;
  assign \new_[11865]_  = ~\new_[12576]_  & ~\new_[12739]_ ;
  assign \new_[11866]_  = ~\new_[12566]_  & ~\new_[12935]_ ;
  assign \new_[11867]_  = ~\new_[12558]_  & ~\new_[13008]_ ;
  assign \new_[11868]_  = ~\new_[12557]_  & ~\new_[12881]_ ;
  assign \new_[11869]_  = ~\new_[13064]_  & ~\new_[12998]_ ;
  assign \new_[11870]_  = ~\new_[13066]_  & ~\new_[13020]_ ;
  assign \new_[11871]_  = ~\new_[12565]_  & ~\new_[12897]_ ;
  assign \new_[11872]_  = ~\new_[12678]_  & ~\new_[13008]_ ;
  assign \new_[11873]_  = ~\new_[12936]_  & ~\new_[12551]_ ;
  assign \new_[11874]_  = ~\new_[12573]_  & ~\new_[12989]_ ;
  assign \new_[11875]_  = ~\new_[12678]_  & ~\new_[12941]_ ;
  assign \new_[11876]_  = ~\new_[12938]_  & ~\new_[12619]_ ;
  assign \new_[11877]_  = ~\new_[13026]_  & ~\new_[12550]_ ;
  assign \new_[11878]_  = ~\new_[12687]_  & ~\new_[12934]_ ;
  assign \new_[11879]_  = ~\new_[12678]_  & ~\new_[12923]_ ;
  assign \new_[11880]_  = ~\new_[12562]_  & ~\new_[12897]_ ;
  assign \new_[11881]_  = ~\new_[12678]_  & ~\new_[12936]_ ;
  assign \new_[11882]_  = ~\new_[12941]_  & ~\new_[12568]_ ;
  assign \new_[11883]_  = ~\new_[12678]_  & ~\new_[12910]_ ;
  assign \new_[11884]_  = ~\new_[12543]_  & ~\new_[13060]_ ;
  assign \new_[11885]_  = ~\new_[12913]_  & ~\new_[12525]_ ;
  assign \new_[11886]_  = ~\new_[13043]_  & ~\new_[12568]_ ;
  assign \new_[11887]_  = ~\new_[12569]_  & ~\new_[13053]_ ;
  assign \new_[11888]_  = ~\new_[12941]_  & ~\new_[12552]_ ;
  assign \new_[11889]_  = ~\new_[12689]_  | ~\new_[12748]_ ;
  assign \new_[11890]_  = ~\new_[2922]_  | ~\new_[12594]_ ;
  assign \new_[11891]_  = ~\new_[13043]_  & ~\new_[12950]_ ;
  assign \new_[11892]_  = ~\new_[12625]_  & ~\new_[13041]_ ;
  assign \new_[11893]_  = ~\new_[12687]_  & ~\new_[13004]_ ;
  assign \new_[11894]_  = ~\new_[12678]_  & ~\new_[13020]_ ;
  assign \new_[11895]_  = ~\new_[13054]_  & ~\new_[12619]_ ;
  assign \new_[11896]_  = ~\new_[12546]_  & ~\new_[13046]_ ;
  assign \new_[11897]_  = ~\new_[12570]_  & ~\new_[12989]_ ;
  assign \new_[11898]_  = ~\new_[12624]_  & ~\new_[12910]_ ;
  assign \new_[11899]_  = ~\new_[12564]_  & ~\new_[12905]_ ;
  assign \new_[11900]_  = ~\new_[12558]_  & ~\new_[13034]_ ;
  assign \new_[11901]_  = ~\new_[12910]_  & ~\new_[12950]_ ;
  assign \new_[11902]_  = ~\new_[12628]_  & ~\new_[13020]_ ;
  assign \new_[11903]_  = ~\new_[12908]_  & ~\new_[12935]_ ;
  assign \new_[11904]_  = ~\new_[13064]_  & ~\new_[13026]_ ;
  assign \new_[11905]_  = ~\new_[12558]_  & ~\new_[12989]_ ;
  assign \new_[11906]_  = ~\new_[12573]_  & ~\new_[13020]_ ;
  assign \new_[11907]_  = ~\new_[13003]_  & ~\new_[12950]_ ;
  assign \new_[11908]_  = ~\new_[12573]_  & ~\new_[12938]_ ;
  assign \new_[11909]_  = ~\new_[12563]_  & ~\new_[13042]_ ;
  assign \new_[11910]_  = ~\new_[12687]_  & ~\new_[12738]_ ;
  assign \new_[11911]_  = ~\new_[12556]_  & ~\new_[13046]_ ;
  assign \new_[11912]_  = ~\new_[12937]_  & ~\new_[12550]_ ;
  assign \new_[11913]_  = ~\new_[12562]_  & ~\new_[12913]_ ;
  assign \new_[11914]_  = ~\new_[12908]_  & ~\new_[12938]_ ;
  assign \new_[11915]_  = ~\new_[12939]_  & ~\new_[12568]_ ;
  assign \new_[11916]_  = ~\new_[13066]_  & ~\new_[13003]_ ;
  assign \new_[11917]_  = ~\new_[12948]_  & ~\new_[13054]_ ;
  assign \new_[11918]_  = ~\new_[13064]_  & ~\new_[13060]_ ;
  assign \new_[11919]_  = ~\new_[12570]_  & ~\new_[13034]_ ;
  assign \new_[11920]_  = ~\new_[12645]_  & ~\new_[12905]_ ;
  assign \new_[11921]_  = ~\new_[12570]_  & ~\new_[13004]_ ;
  assign \new_[11922]_  = ~\new_[12567]_  & ~\new_[12881]_ ;
  assign \new_[11923]_  = ~\new_[13004]_  & ~\new_[12551]_ ;
  assign \new_[11924]_  = ~\new_[12631]_  & ~\new_[12897]_ ;
  assign \new_[11925]_  = ~\new_[12739]_  & ~\new_[12525]_ ;
  assign \new_[11926]_  = ~\new_[12989]_  & ~\new_[12597]_ ;
  assign \new_[11927]_  = ~\new_[13064]_  & ~\new_[12941]_ ;
  assign \new_[11928]_  = ~\new_[12937]_  & ~\new_[12568]_ ;
  assign \new_[11929]_  = ~\new_[12908]_  & ~\new_[12939]_ ;
  assign \new_[11930]_  = ~\new_[12562]_  & ~\new_[13043]_ ;
  assign \new_[11931]_  = ~\new_[12678]_  & ~\new_[12738]_ ;
  assign \new_[11932]_  = ~\new_[13066]_  & ~\new_[13041]_ ;
  assign \new_[11933]_  = ~\new_[12564]_  & ~\new_[13034]_ ;
  assign \new_[11934]_  = ~\new_[12559]_  & ~\new_[12939]_ ;
  assign \new_[11935]_  = ~\new_[12564]_  & ~\new_[12999]_ ;
  assign \new_[11936]_  = ~\new_[12628]_  & ~\new_[13003]_ ;
  assign \new_[11937]_  = ~\new_[13060]_  & ~\new_[12568]_ ;
  assign \new_[11938]_  = ~\new_[12687]_  & ~\new_[12936]_ ;
  assign \new_[11939]_  = ~\new_[13066]_  & ~\new_[12910]_ ;
  assign \new_[11940]_  = ~\new_[12556]_  & ~\new_[12739]_ ;
  assign \new_[11941]_  = ~\new_[12905]_  & ~\new_[12568]_ ;
  assign \new_[11942]_  = ~\new_[13060]_  & ~\new_[12552]_ ;
  assign \new_[11943]_  = ~\new_[12738]_  & ~\new_[12550]_ ;
  assign \new_[11944]_  = ~\new_[13004]_  & ~\new_[12568]_ ;
  assign \new_[11945]_  = ~\new_[13081]_  & ~\new_[12998]_ ;
  assign \new_[11946]_  = ~\new_[12565]_  & ~\new_[13043]_ ;
  assign \new_[11947]_  = ~\new_[13042]_  & ~\new_[12568]_ ;
  assign \new_[11948]_  = ~\new_[12939]_  & ~\new_[12550]_ ;
  assign \new_[11949]_  = ~\new_[12569]_  & ~\new_[12938]_ ;
  assign \new_[11950]_  = ~\new_[12881]_  & ~\new_[12568]_ ;
  assign \new_[11951]_  = ~\new_[12563]_  & ~\new_[13004]_ ;
  assign \new_[11952]_  = ~\new_[12645]_  & ~\new_[12989]_ ;
  assign \new_[11953]_  = ~\new_[13066]_  & ~\new_[13053]_ ;
  assign \new_[11954]_  = ~\new_[12559]_  & ~\new_[12937]_ ;
  assign \new_[11955]_  = ~\new_[12687]_  & ~\new_[13026]_ ;
  assign \new_[11956]_  = ~\new_[12587]_  | ~\new_[12745]_ ;
  assign \new_[11957]_  = ~\new_[13064]_  & ~\new_[13004]_ ;
  assign \new_[11958]_  = ~\new_[12687]_  & ~\new_[13008]_ ;
  assign \new_[11959]_  = ~\new_[12687]_  & ~\new_[12884]_ ;
  assign \new_[11960]_  = ~\new_[12703]_  & ~\new_[13060]_ ;
  assign \new_[11961]_  = ~\new_[12562]_  & ~\new_[12941]_ ;
  assign \new_[11962]_  = ~\new_[13003]_  & ~\new_[12568]_ ;
  assign \new_[11963]_  = ~\new_[12897]_  & ~\new_[12550]_ ;
  assign \new_[11964]_  = ~\new_[12543]_  & ~\new_[13053]_ ;
  assign \new_[11965]_  = ~\new_[12566]_  & ~\new_[12939]_ ;
  assign \new_[11966]_  = ~\new_[12678]_  & ~\new_[13004]_ ;
  assign \new_[11967]_  = ~\new_[12678]_  & ~\new_[13060]_ ;
  assign \new_[11968]_  = ~\new_[12998]_  & ~\new_[12619]_ ;
  assign \new_[11969]_  = ~\new_[12697]_  & ~\new_[12935]_ ;
  assign \new_[11970]_  = ~\new_[13050]_  & ~\new_[13026]_ ;
  assign \new_[11971]_  = ~\new_[12678]_  & ~\new_[12998]_ ;
  assign \new_[11972]_  = ~\new_[13053]_  & ~\new_[12551]_ ;
  assign \new_[11973]_  = ~\new_[12566]_  & ~\new_[13008]_ ;
  assign \new_[11974]_  = ~\new_[12625]_  & ~\new_[12936]_ ;
  assign \new_[11975]_  = ~\new_[12703]_  & ~\new_[12738]_ ;
  assign \new_[11976]_  = ~\new_[12697]_  & ~\new_[12999]_ ;
  assign \new_[11977]_  = ~\new_[12948]_  & ~\new_[12905]_ ;
  assign \new_[11978]_  = ~\new_[12576]_  & ~\new_[12934]_ ;
  assign \new_[11979]_  = ~\new_[12948]_  & ~\new_[13008]_ ;
  assign \new_[11980]_  = ~\new_[12546]_  & ~\new_[13008]_ ;
  assign \new_[11981]_  = ~\new_[12690]_  & ~\new_[12881]_ ;
  assign \new_[11982]_  = ~\new_[12905]_  & ~\new_[12525]_ ;
  assign \new_[11983]_  = ~\new_[12543]_  & ~\new_[12936]_ ;
  assign \new_[11984]_  = ~\new_[12546]_  & ~\new_[12884]_ ;
  assign \new_[11985]_  = ~\new_[12678]_  & ~\new_[12989]_ ;
  assign \new_[11986]_  = ~\new_[12563]_  & ~\new_[13054]_ ;
  assign \new_[11987]_  = ~\new_[12567]_  & ~\new_[13054]_ ;
  assign \new_[11988]_  = ~\new_[12678]_  & ~\new_[13054]_ ;
  assign \new_[11989]_  = ~\new_[12948]_  & ~\new_[12935]_ ;
  assign \new_[11990]_  = ~\new_[13064]_  & ~\new_[12884]_ ;
  assign \new_[11991]_  = ~\new_[12557]_  & ~\new_[12913]_ ;
  assign \new_[11992]_  = ~\new_[12631]_  & ~\new_[12941]_ ;
  assign \new_[11993]_  = ~\new_[12631]_  & ~\new_[12881]_ ;
  assign \new_[11994]_  = ~\new_[12576]_  & ~\new_[12923]_ ;
  assign \new_[11995]_  = ~\new_[12569]_  & ~\new_[13060]_ ;
  assign \new_[11996]_  = ~\new_[12624]_  & ~\new_[12884]_ ;
  assign \new_[11997]_  = ~\new_[12910]_  & ~\new_[12568]_ ;
  assign \new_[11998]_  = ~\new_[12934]_  & ~\new_[12619]_ ;
  assign \new_[11999]_  = \new_[4763]_  ^ \new_[13990]_ ;
  assign \new_[12000]_  = ~\new_[12656]_  & (~\new_[7496]_  | ~\new_[13141]_ );
  assign \new_[12001]_  = ~\new_[12530]_  & (~\new_[13188]_  | ~\new_[12991]_ );
  assign \new_[12002]_  = ~\new_[12806]_  & (~\new_[13480]_  | ~\new_[7935]_ );
  assign n10971 = \new_[13092]_  ^ \new_[12883]_ ;
  assign n10966 = \new_[13124]_  ^ \new_[12894]_ ;
  assign \new_[12005]_  = ~\new_[5135]_  | ~\new_[12553]_ ;
  assign \new_[12006]_  = \new_[13105]_  ^ \new_[12796]_ ;
  assign n10956 = \new_[13158]_  ^ \new_[13869]_ ;
  assign n10961 = \new_[13161]_  ^ \new_[12990]_ ;
  assign \new_[12009]_  = ~\new_[4085]_  | ~\new_[12594]_ ;
  assign \new_[12010]_  = \new_[13500]_  ^ \new_[12990]_ ;
  assign \new_[12011]_  = \new_[12894]_  ^ \new_[13622]_ ;
  assign \new_[12012]_  = \new_[13794]_  ^ \new_[13869]_ ;
  assign \new_[12013]_  = \new_[14127]_  ^ \new_[12883]_ ;
  assign \new_[12014]_  = ~\new_[13020]_  & ~\new_[12551]_ ;
  assign \new_[12015]_  = ~\new_[4409]_  | ~\new_[12594]_ ;
  assign \new_[12016]_  = ~\new_[12354]_ ;
  assign \new_[12017]_  = ~\new_[4899]_  | ~\new_[12554]_ ;
  assign \new_[12018]_  = ~\new_[12362]_ ;
  assign \new_[12019]_  = ~\new_[12417]_ ;
  assign \new_[12020]_  = \\u15_crac_din_reg[12] ;
  assign \new_[12021]_  = ~\new_[12447]_ ;
  assign \new_[12022]_  = ~\new_[13895]_ ;
  assign \new_[12023]_  = ~\new_[13895]_ ;
  assign \new_[12024]_  = ~\new_[12581]_  | ~\new_[7928]_ ;
  assign \new_[12025]_  = ~\new_[12440]_ ;
  assign \new_[12026]_  = ~\new_[12437]_ ;
  assign \new_[12027]_  = ~\new_[12436]_ ;
  assign \new_[12028]_  = ~\new_[12433]_ ;
  assign \new_[12029]_  = ~\new_[12341]_ ;
  assign \new_[12030]_  = ~\new_[12429]_ ;
  assign \new_[12031]_  = ~\new_[5149]_  | ~\new_[12644]_ ;
  assign \new_[12032]_  = (~\new_[13840]_  | ~\new_[12842]_ ) & (~\new_[13814]_  | ~\new_[12918]_ );
  assign \new_[12033]_  = ~\new_[12808]_  | ~\new_[5071]_  | ~\new_[5070]_ ;
  assign \new_[12034]_  = ~\new_[12809]_  | ~\new_[5059]_  | ~\new_[5058]_ ;
  assign \new_[12035]_  = ~\new_[12810]_  | ~\new_[5066]_  | ~\new_[5065]_ ;
  assign \new_[12036]_  = ~\new_[12998]_  & ~\new_[12568]_ ;
  assign \new_[12037]_  = ~\new_[5015]_  | ~\new_[12644]_ ;
  assign \new_[12038]_  = ~\new_[5002]_  | ~\new_[12644]_ ;
  assign \new_[12039]_  = ~\new_[13012]_ ;
  assign \new_[12040]_  = ~\new_[12325]_ ;
  assign \new_[12041]_  = ~\new_[13008]_  & ~\new_[12568]_ ;
  assign \new_[12042]_  = ~\new_[12993]_ ;
  assign \new_[12043]_  = ~\new_[5442]_  | ~\new_[12593]_ ;
  assign \new_[12044]_  = ~\new_[4919]_  | ~\new_[12553]_ ;
  assign \new_[12045]_  = \\u15_crac_din_reg[1] ;
  assign \new_[12046]_  = ~\new_[5141]_  | ~\new_[12554]_ ;
  assign \new_[12047]_  = (~\new_[12982]_  | ~\new_[13336]_ ) & (~\new_[13368]_  | ~\new_[12779]_ );
  assign \new_[12048]_  = \\u15_crac_din_reg[7] ;
  assign \new_[12049]_  = (~\new_[12982]_  | ~\new_[13864]_ ) & (~\new_[13603]_  | ~\new_[12779]_ );
  assign \new_[12050]_  = ~\new_[5444]_  | ~\new_[14118]_ ;
  assign \new_[12051]_  = \\u15_crac_din_reg[14] ;
  assign \new_[12052]_  = (~\new_[12778]_  | ~\new_[13222]_ ) & (~\new_[13675]_  | ~\new_[12805]_ );
  assign \new_[12053]_  = (~\new_[13227]_  | ~\new_[12763]_ ) & (~\new_[13693]_  | ~\new_[13023]_ );
  assign \new_[12054]_  = (~\new_[13495]_  | ~\new_[12842]_ ) & (~\new_[13776]_  | ~\new_[12918]_ );
  assign \new_[12055]_  = ~\new_[14175]_ ;
  assign \new_[12056]_  = (~\new_[13514]_  | ~\new_[12805]_ ) & (~\new_[13362]_  | ~\new_[13023]_ );
  assign \new_[12057]_  = \\u15_crac_din_reg[10] ;
  assign \new_[12058]_  = \\u15_crac_din_reg[15] ;
  assign \new_[12059]_  = \\u15_crac_din_reg[4] ;
  assign \new_[12060]_  = \\u15_crac_din_reg[8] ;
  assign \new_[12061]_  = (~\new_[12982]_  | ~\new_[13296]_ ) & (~\new_[13224]_  | ~\new_[12747]_ );
  assign \new_[12062]_  = \\u15_crac_din_reg[11] ;
  assign \new_[12063]_  = ~\new_[12948]_  & ~\new_[12999]_ ;
  assign \new_[12064]_  = (~\new_[12777]_  | ~\new_[13674]_ ) & (~\new_[13751]_  | ~\new_[12740]_ );
  assign \new_[12065]_  = \\u15_crac_din_reg[13] ;
  assign \new_[12066]_  = \\u15_crac_din_reg[2] ;
  assign \new_[12067]_  = (~\new_[13628]_  | ~\new_[12805]_ ) & (~\new_[13333]_  | ~\new_[12763]_ );
  assign \new_[12068]_  = ~\new_[12512]_  & (~\new_[13672]_  | ~\new_[13023]_ );
  assign \new_[12069]_  = \\u15_crac_din_reg[0] ;
  assign \new_[12070]_  = \new_[13127]_  ^ \new_[12855]_ ;
  assign \new_[12071]_  = (~\new_[13192]_  | ~\new_[12842]_ ) & (~\new_[13348]_  | ~\new_[12918]_ );
  assign \new_[12072]_  = ~\new_[12506]_  & ~\new_[13300]_ ;
  assign \new_[12073]_  = ~\new_[12454]_ ;
  assign \new_[12074]_  = ~\new_[12454]_ ;
  assign \new_[12075]_  = \\u15_crac_din_reg[5] ;
  assign \new_[12076]_  = ~\new_[12687]_  & ~\new_[12939]_ ;
  assign \new_[12077]_  = ~\new_[4641]_  | ~\new_[4631]_  | ~\new_[12694]_  | ~\new_[13747]_ ;
  assign \new_[12078]_  = ~\new_[13041]_  & ~\new_[12568]_ ;
  assign \new_[12079]_  = ~\new_[13656]_  | ~\new_[12947]_  | ~\new_[12806]_ ;
  assign \new_[12080]_  = ~\new_[2736]_  | ~\new_[12594]_ ;
  assign \new_[12081]_  = ~\new_[7979]_  | ~\new_[12947]_  | ~\new_[12806]_ ;
  assign \new_[12082]_  = \new_[4728]_  ^ \new_[12879]_ ;
  assign \new_[12083]_  = \new_[7936]_  ^ \new_[12877]_ ;
  assign \new_[12084]_  = \new_[8099]_  ^ \new_[12875]_ ;
  assign \new_[12085]_  = \\u5_status_reg[0] ;
  assign \new_[12086]_  = \\u8_status_reg[0] ;
  assign \new_[12087]_  = ~\new_[12846]_  | ~\new_[12679]_ ;
  assign \new_[12088]_  = \new_[12704]_  | \wb_addr_i[6] ;
  assign \new_[12089]_  = \new_[12704]_  | wb_we_i;
  assign \new_[12090]_  = ~\new_[12531]_  | ~\new_[12594]_ ;
  assign \new_[12091]_  = ~\new_[5163]_  | ~\new_[12644]_ ;
  assign \new_[12092]_  = ~\new_[5213]_  | ~\new_[12657]_ ;
  assign \new_[12093]_  = ~\new_[5419]_  | ~\new_[12585]_ ;
  assign \new_[12094]_  = ~\new_[12608]_  | ~\new_[4856]_ ;
  assign \new_[12095]_  = ~\new_[5248]_  | ~\new_[13930]_ ;
  assign \new_[12096]_  = ~\new_[12608]_  | ~\new_[4978]_ ;
  assign \new_[12097]_  = \new_[13169]_  ^ \new_[12799]_ ;
  assign \new_[12098]_  = ~\new_[13020]_  & ~\new_[12621]_ ;
  assign n10951 = ~\new_[12347]_ ;
  assign \new_[12100]_  = ~\new_[12609]_  | (~\new_[7492]_  & ~\new_[13096]_ );
  assign \new_[12101]_  = ~\new_[2747]_  | ~\new_[12594]_ ;
  assign \new_[12102]_  = ~\new_[13081]_  & ~\new_[12936]_ ;
  assign \new_[12103]_  = \new_[14133]_  | \new_[14127]_ ;
  assign \new_[12104]_  = \\u15_crac_din_reg[3] ;
  assign \new_[12105]_  = ~\new_[12581]_  | ~\new_[5855]_ ;
  assign \new_[12106]_  = ~\new_[12581]_  | ~\new_[3184]_ ;
  assign \new_[12107]_  = ~\new_[13072]_  | ~\new_[12931]_  | ~\new_[12882]_  | ~\new_[13069]_ ;
  assign \new_[12108]_  = ~\new_[12933]_  | ~\new_[13051]_  | ~\new_[12927]_  | ~\new_[13061]_ ;
  assign \new_[12109]_  = ~\new_[12678]_  & ~\new_[13003]_ ;
  assign \new_[12110]_  = ~\new_[5331]_  | ~\new_[14188]_ ;
  assign \new_[12111]_  = \new_[13144]_  ^ \new_[13142]_ ;
  assign \new_[12112]_  = \new_[13175]_  ^ \new_[13113]_ ;
  assign \new_[12113]_  = ~\new_[5246]_  | ~\new_[13930]_ ;
  assign n10976 = \\u1_sr_reg[1] ;
  assign \new_[12115]_  = ~\new_[12522]_  | ~\new_[7976]_ ;
  assign \new_[12116]_  = ~\new_[12614]_  | ~\new_[13480]_ ;
  assign \new_[12117]_  = ~\new_[12455]_ ;
  assign \new_[12118]_  = \new_[12670]_  | ac97_reset_pad_o_;
  assign \new_[12119]_  = ~\new_[7974]_  | ~\new_[13624]_  | ~\new_[12658]_  | ~\new_[13554]_ ;
  assign \new_[12120]_  = ~\new_[12509]_  | ~\new_[13538]_ ;
  assign \new_[12121]_  = ~\new_[12972]_  | ~\new_[4639]_  | ~\new_[4642]_  | ~\new_[4640]_ ;
  assign \new_[12122]_  = ~\new_[7972]_  | ~\new_[12505]_  | ~\new_[7978]_ ;
  assign \new_[12123]_  = (~\new_[12992]_  | ~\new_[12781]_ ) & (~\new_[14127]_  | ~\new_[2759]_ );
  assign \new_[12124]_  = (~\new_[12778]_  | ~\new_[13479]_ ) & (~\new_[13583]_  | ~\new_[12805]_ );
  assign \new_[12125]_  = ~\new_[12515]_  & (~\new_[13800]_  | ~\new_[13023]_ );
  assign \new_[12126]_  = (~\new_[12778]_  | ~\new_[13279]_ ) & (~\new_[13194]_  | ~\new_[12763]_ );
  assign \new_[12127]_  = (~\new_[12778]_  | ~\new_[13410]_ ) & (~\new_[13494]_  | ~\new_[12805]_ );
  assign \new_[12128]_  = (~\new_[13284]_  | ~\new_[12763]_ ) & (~\new_[13468]_  | ~\new_[13023]_ );
  assign \new_[12129]_  = (~\new_[13854]_  | ~\new_[12763]_ ) & (~\new_[13328]_  | ~\new_[13023]_ );
  assign \new_[12130]_  = (~\new_[13621]_  | ~\new_[12763]_ ) & (~\new_[13327]_  | ~\new_[13023]_ );
  assign \new_[12131]_  = (~\new_[12778]_  | ~\new_[13356]_ ) & (~\new_[13294]_  | ~\new_[12805]_ );
  assign \new_[12132]_  = (~\new_[13257]_  | ~\new_[12763]_ ) & (~\new_[13528]_  | ~\new_[13023]_ );
  assign \new_[12133]_  = (~\new_[12777]_  | ~\new_[13808]_ ) & (~\new_[13287]_  | ~\new_[12740]_ );
  assign \new_[12134]_  = (~\new_[12778]_  | ~\new_[13517]_ ) & (~\new_[13690]_  | ~\new_[13023]_ );
  assign \new_[12135]_  = (~\new_[12778]_  | ~\new_[13848]_ ) & (~\new_[13409]_  | ~\new_[12805]_ );
  assign \new_[12136]_  = (~\new_[13830]_  | ~\new_[12763]_ ) & (~\new_[13346]_  | ~\new_[13023]_ );
  assign \new_[12137]_  = (~\new_[13558]_  | ~\new_[12805]_ ) & (~\new_[13670]_  | ~\new_[13023]_ );
  assign \new_[12138]_  = (~\new_[12778]_  | ~\new_[13618]_ ) & (~\new_[13516]_  | ~\new_[12805]_ );
  assign \new_[12139]_  = (~\new_[12778]_  | ~\new_[13432]_ ) & (~\new_[13819]_  | ~\new_[12805]_ );
  assign \new_[12140]_  = (~\new_[13521]_  | ~\new_[12763]_ ) & (~\new_[13512]_  | ~\new_[13023]_ );
  assign \new_[12141]_  = (~\new_[13271]_  | ~\new_[12805]_ ) & (~\new_[13804]_  | ~\new_[12763]_ );
  assign \new_[12142]_  = (~\new_[12778]_  | ~\new_[13851]_ ) & (~\new_[13633]_  | ~\new_[13023]_ );
  assign \new_[12143]_  = (~\new_[13835]_  | ~\new_[12763]_ ) & (~\new_[13297]_  | ~\new_[13023]_ );
  assign \new_[12144]_  = (~\new_[12778]_  | ~\new_[13203]_ ) & (~\new_[13398]_  | ~\new_[12805]_ );
  assign \new_[12145]_  = (~\new_[13566]_  | ~\new_[12763]_ ) & (~\new_[13298]_  | ~\new_[13023]_ );
  assign \new_[12146]_  = (~\new_[13302]_  | ~\new_[12805]_ ) & (~\new_[13685]_  | ~\new_[13023]_ );
  assign \new_[12147]_  = (~\new_[12778]_  | ~\new_[13636]_ ) & (~\new_[13781]_  | ~\new_[12805]_ );
  assign \new_[12148]_  = (~\new_[13825]_  | ~\new_[12805]_ ) & (~\new_[13839]_  | ~\new_[13023]_ );
  assign \new_[12149]_  = (~\new_[13254]_  | ~\new_[12763]_ ) & (~\new_[13374]_  | ~\new_[13023]_ );
  assign \new_[12150]_  = (~\new_[12778]_  | ~\new_[13349]_ ) & (~\new_[13568]_  | ~\new_[12805]_ );
  assign \new_[12151]_  = (~\new_[13286]_  | ~\new_[12763]_ ) & (~\new_[13305]_  | ~\new_[13023]_ );
  assign \new_[12152]_  = (~\new_[12778]_  | ~\new_[13581]_ ) & (~\new_[13378]_  | ~\new_[12805]_ );
  assign \new_[12153]_  = (~\new_[13289]_  | ~\new_[12763]_ ) & (~\new_[13609]_  | ~\new_[13023]_ );
  assign \new_[12154]_  = (~\new_[13555]_  | ~\new_[12805]_ ) & (~\new_[13307]_  | ~\new_[13023]_ );
  assign \new_[12155]_  = (~\new_[12778]_  | ~\new_[13504]_ ) & (~\new_[13436]_  | ~\new_[12805]_ );
  assign \new_[12156]_  = (~\new_[13406]_  | ~\new_[12763]_ ) & (~\new_[13746]_  | ~\new_[13023]_ );
  assign \new_[12157]_  = (~\new_[12778]_  | ~\new_[13484]_ ) & (~\new_[13452]_  | ~\new_[12805]_ );
  assign \new_[12158]_  = (~\new_[12778]_  | ~\new_[13774]_ ) & (~\new_[13638]_  | ~\new_[12805]_ );
  assign \new_[12159]_  = (~\new_[13542]_  | ~\new_[12763]_ ) & (~\new_[13290]_  | ~\new_[13023]_ );
  assign \new_[12160]_  = (~\new_[13544]_  | ~\new_[12763]_ ) & (~\new_[13216]_  | ~\new_[13023]_ );
  assign \new_[12161]_  = (~\new_[13499]_  | ~\new_[12763]_ ) & (~\new_[13268]_  | ~\new_[13023]_ );
  assign \new_[12162]_  = (~\new_[12778]_  | ~\new_[13202]_ ) & (~\new_[13591]_  | ~\new_[12763]_ );
  assign \new_[12163]_  = (~\new_[13713]_  | ~\new_[12763]_ ) & (~\new_[13381]_  | ~\new_[13023]_ );
  assign \new_[12164]_  = (~\new_[13699]_  | ~\new_[12763]_ ) & (~\new_[13376]_  | ~\new_[13023]_ );
  assign \new_[12165]_  = (~\new_[12778]_  | ~\new_[13418]_ ) & (~\new_[13193]_  | ~\new_[12805]_ );
  assign \new_[12166]_  = (~\new_[12778]_  | ~\new_[13491]_ ) & (~\new_[13285]_  | ~\new_[12763]_ );
  assign \new_[12167]_  = (~\new_[13283]_  | ~\new_[12763]_ ) & (~\new_[13301]_  | ~\new_[13023]_ );
  assign \new_[12168]_  = (~\new_[13679]_  | ~\new_[12763]_ ) & (~\new_[13329]_  | ~\new_[13023]_ );
  assign \new_[12169]_  = (~\new_[12778]_  | ~\new_[13312]_ ) & (~\new_[13586]_  | ~\new_[12763]_ );
  assign \new_[12170]_  = (~\new_[13246]_  | ~\new_[12805]_ ) & (~\new_[13637]_  | ~\new_[13023]_ );
  assign \new_[12171]_  = (~\new_[12982]_  | ~\new_[13530]_ ) & (~\new_[13232]_  | ~\new_[12779]_ );
  assign \new_[12172]_  = (~\new_[13420]_  | ~\new_[12805]_ ) & (~\new_[13310]_  | ~\new_[12763]_ );
  assign \new_[12173]_  = (~\new_[12778]_  | ~\new_[13842]_ ) & (~\new_[13386]_  | ~\new_[13023]_ );
  assign \new_[12174]_  = (~\new_[13792]_  | ~\new_[12779]_ ) & (~\new_[13380]_  | ~\new_[13011]_ );
  assign \new_[12175]_  = (~\new_[12982]_  | ~\new_[13357]_ ) & (~\new_[13277]_  | ~\new_[12779]_ );
  assign \new_[12176]_  = (~\new_[13752]_  | ~\new_[12740]_ ) & (~\new_[13342]_  | ~\new_[12918]_ );
  assign \new_[12177]_  = (~\new_[12982]_  | ~\new_[13817]_ ) & (~\new_[13543]_  | ~\new_[12779]_ );
  assign \new_[12178]_  = (~\new_[12982]_  | ~\new_[13205]_ ) & (~\new_[13787]_  | ~\new_[12747]_ );
  assign \new_[12179]_  = (~\new_[13861]_  | ~\new_[12779]_ ) & (~\new_[13321]_  | ~\new_[13011]_ );
  assign \new_[12180]_  = (~\new_[12778]_  | ~\new_[13852]_ ) & (~\new_[13417]_  | ~\new_[12805]_ );
  assign \new_[12181]_  = (~\new_[12982]_  | ~\new_[13610]_ ) & (~\new_[13668]_  | ~\new_[12747]_ );
  assign \new_[12182]_  = (~\new_[13237]_  | ~\new_[12779]_ ) & (~\new_[13564]_  | ~\new_[13011]_ );
  assign \new_[12183]_  = (~\new_[12778]_  | ~\new_[13400]_ ) & (~\new_[13845]_  | ~\new_[12805]_ );
  assign \new_[12184]_  = ~\new_[12555]_  & ~\new_[13054]_ ;
  assign \new_[12185]_  = (~\new_[12777]_  | ~\new_[13658]_ ) & (~\new_[13696]_  | ~\new_[12740]_ );
  assign \new_[12186]_  = ~\new_[12518]_  & (~\new_[13631]_  | ~\new_[12918]_ );
  assign \new_[12187]_  = (~\new_[12778]_  | ~\new_[13485]_ ) & (~\new_[13439]_  | ~\new_[12805]_ );
  assign \new_[12188]_  = (~\new_[12777]_  | ~\new_[13686]_ ) & (~\new_[13843]_  | ~\new_[12740]_ );
  assign \new_[12189]_  = ~\new_[12705]_  & (~\new_[13782]_  | ~\new_[12918]_ );
  assign \new_[12190]_  = (~\new_[12777]_  | ~\new_[13212]_ ) & (~\new_[13736]_  | ~\new_[12740]_ );
  assign \new_[12191]_  = (~\new_[12777]_  | ~\new_[13742]_ ) & (~\new_[13737]_  | ~\new_[12740]_ );
  assign \new_[12192]_  = ~\new_[12523]_  & (~\new_[13807]_  | ~\new_[12918]_ );
  assign \new_[12193]_  = (~\new_[13649]_  | ~\new_[12747]_ ) & (~\new_[13549]_  | ~\new_[13011]_ );
  assign \new_[12194]_  = (~\new_[12777]_  | ~\new_[13534]_ ) & (~\new_[13664]_  | ~\new_[12842]_ );
  assign \new_[12195]_  = (~\new_[13423]_  | ~\new_[12740]_ ) & (~\new_[13630]_  | ~\new_[12918]_ );
  assign \new_[12196]_  = (~\new_[12777]_  | ~\new_[13540]_ ) & (~\new_[13390]_  | ~\new_[12740]_ );
  assign \new_[12197]_  = (~\new_[13580]_  | ~\new_[12842]_ ) & (~\new_[13662]_  | ~\new_[12918]_ );
  assign \new_[12198]_  = (~\new_[12982]_  | ~\new_[13533]_ ) & (~\new_[13667]_  | ~\new_[12747]_ );
  assign \new_[12199]_  = (~\new_[12777]_  | ~\new_[13464]_ ) & (~\new_[13727]_  | ~\new_[12740]_ );
  assign \new_[12200]_  = (~\new_[13627]_  | ~\new_[12842]_ ) & (~\new_[13236]_  | ~\new_[12918]_ );
  assign \new_[12201]_  = (~\new_[12777]_  | ~\new_[13567]_ ) & (~\new_[13741]_  | ~\new_[12740]_ );
  assign \new_[12202]_  = (~\new_[13646]_  | ~\new_[12842]_ ) & (~\new_[13684]_  | ~\new_[12918]_ );
  assign \new_[12203]_  = (~\new_[13680]_  | ~\new_[12842]_ ) & (~\new_[13652]_  | ~\new_[12918]_ );
  assign \new_[12204]_  = (~\new_[12777]_  | ~\new_[13332]_ ) & (~\new_[13522]_  | ~\new_[12740]_ );
  assign \new_[12205]_  = (~\new_[13705]_  | ~\new_[12842]_ ) & (~\new_[13593]_  | ~\new_[12918]_ );
  assign \new_[12206]_  = (~\new_[12982]_  | ~\new_[13607]_ ) & (~\new_[13806]_  | ~\new_[12779]_ );
  assign \new_[12207]_  = (~\new_[12777]_  | ~\new_[13359]_ ) & (~\new_[13341]_  | ~\new_[12740]_ );
  assign \new_[12208]_  = (~\new_[13402]_  | ~\new_[12842]_ ) & (~\new_[13694]_  | ~\new_[12918]_ );
  assign \new_[12209]_  = (~\new_[13250]_  | ~\new_[12747]_ ) & (~\new_[13498]_  | ~\new_[13011]_ );
  assign \new_[12210]_  = (~\new_[12778]_  | ~\new_[13256]_ ) & (~\new_[13577]_  | ~\new_[12805]_ );
  assign \new_[12211]_  = (~\new_[12777]_  | ~\new_[13682]_ ) & (~\new_[13426]_  | ~\new_[12740]_ );
  assign \new_[12212]_  = (~\new_[13613]_  | ~\new_[12842]_ ) & (~\new_[13635]_  | ~\new_[12918]_ );
  assign \new_[12213]_  = (~\new_[12777]_  | ~\new_[13716]_ ) & (~\new_[13838]_  | ~\new_[12740]_ );
  assign \new_[12214]_  = ~\new_[12687]_  & ~\new_[13042]_ ;
  assign \new_[12215]_  = (~\new_[13773]_  | ~\new_[12842]_ ) & (~\new_[13616]_  | ~\new_[12918]_ );
  assign \new_[12216]_  = (~\new_[12777]_  | ~\new_[13594]_ ) & (~\new_[13859]_  | ~\new_[12842]_ );
  assign \new_[12217]_  = (~\new_[13303]_  | ~\new_[12740]_ ) & (~\new_[13860]_  | ~\new_[12918]_ );
  assign \new_[12218]_  = ~\new_[5340]_  | ~\new_[14188]_ ;
  assign \new_[12219]_  = (~\new_[13419]_  | ~\new_[12842]_ ) & (~\new_[13763]_  | ~\new_[12918]_ );
  assign \new_[12220]_  = (~\new_[12777]_  | ~\new_[13596]_ ) & (~\new_[13282]_  | ~\new_[12740]_ );
  assign \new_[12221]_  = (~\new_[13422]_  | ~\new_[12842]_ ) & (~\new_[13847]_  | ~\new_[12918]_ );
  assign \new_[12222]_  = (~\new_[12777]_  | ~\new_[13836]_ ) & (~\new_[13261]_  | ~\new_[12740]_ );
  assign \new_[12223]_  = (~\new_[13424]_  | ~\new_[12842]_ ) & (~\new_[13258]_  | ~\new_[12918]_ );
  assign \new_[12224]_  = (~\new_[13276]_  | ~\new_[12747]_ ) & (~\new_[13411]_  | ~\new_[13011]_ );
  assign \new_[12225]_  = (~\new_[12777]_  | ~\new_[13262]_ ) & (~\new_[13245]_  | ~\new_[12740]_ );
  assign \new_[12226]_  = (~\new_[13435]_  | ~\new_[12842]_ ) & (~\new_[13252]_  | ~\new_[12918]_ );
  assign \new_[12227]_  = (~\new_[12777]_  | ~\new_[13323]_ ) & (~\new_[13239]_  | ~\new_[12740]_ );
  assign \new_[12228]_  = (~\new_[13389]_  | ~\new_[12842]_ ) & (~\new_[13427]_  | ~\new_[12918]_ );
  assign \new_[12229]_  = (~\new_[13712]_  | ~\new_[12842]_ ) & (~\new_[13849]_  | ~\new_[12918]_ );
  assign \new_[12230]_  = (~\new_[12777]_  | ~\new_[13706]_ ) & (~\new_[13295]_  | ~\new_[12740]_ );
  assign \new_[12231]_  = (~\new_[12777]_  | ~\new_[13291]_ ) & (~\new_[13211]_  | ~\new_[12740]_ );
  assign \new_[12232]_  = (~\new_[13588]_  | ~\new_[12842]_ ) & (~\new_[13764]_  | ~\new_[12918]_ );
  assign \new_[12233]_  = (~\new_[12777]_  | ~\new_[13641]_ ) & (~\new_[13196]_  | ~\new_[12740]_ );
  assign \new_[12234]_  = (~\new_[13708]_  | ~\new_[12842]_ ) & (~\new_[13204]_  | ~\new_[12918]_ );
  assign \new_[12235]_  = (~\new_[12777]_  | ~\new_[13748]_ ) & (~\new_[13430]_  | ~\new_[12740]_ );
  assign \new_[12236]_  = (~\new_[13556]_  | ~\new_[12842]_ ) & (~\new_[13265]_  | ~\new_[12918]_ );
  assign \new_[12237]_  = (~\new_[12777]_  | ~\new_[13702]_ ) & (~\new_[13242]_  | ~\new_[12740]_ );
  assign \new_[12238]_  = (~\new_[13587]_  | ~\new_[12842]_ ) & (~\new_[13238]_  | ~\new_[12918]_ );
  assign \new_[12239]_  = (~\new_[12777]_  | ~\new_[13475]_ ) & (~\new_[13865]_  | ~\new_[12740]_ );
  assign \new_[12240]_  = (~\new_[12777]_  | ~\new_[13412]_ ) & (~\new_[13431]_  | ~\new_[12740]_ );
  assign \new_[12241]_  = (~\new_[13476]_  | ~\new_[12842]_ ) & (~\new_[13821]_  | ~\new_[12918]_ );
  assign \new_[12242]_  = (~\new_[12777]_  | ~\new_[13834]_ ) & (~\new_[13367]_  | ~\new_[12740]_ );
  assign \new_[12243]_  = (~\new_[13623]_  | ~\new_[12842]_ ) & (~\new_[13351]_  | ~\new_[12918]_ );
  assign \new_[12244]_  = (~\new_[12777]_  | ~\new_[13490]_ ) & (~\new_[13345]_  | ~\new_[12740]_ );
  assign \new_[12245]_  = (~\new_[13768]_  | ~\new_[12842]_ ) & (~\new_[13274]_  | ~\new_[12918]_ );
  assign \new_[12246]_  = (~\new_[12777]_  | ~\new_[13266]_ ) & (~\new_[13510]_  | ~\new_[12740]_ );
  assign \new_[12247]_  = (~\new_[13772]_  | ~\new_[12842]_ ) & (~\new_[13304]_  | ~\new_[12918]_ );
  assign \new_[12248]_  = (~\new_[12777]_  | ~\new_[13719]_ ) & (~\new_[13777]_  | ~\new_[12842]_ );
  assign \new_[12249]_  = (~\new_[12777]_  | ~\new_[13778]_ ) & (~\new_[13440]_  | ~\new_[12740]_ );
  assign \new_[12250]_  = (~\new_[12778]_  | ~\new_[13527]_ ) & (~\new_[13318]_  | ~\new_[12805]_ );
  assign \new_[12251]_  = (~\new_[12777]_  | ~\new_[13731]_ ) & (~\new_[13645]_  | ~\new_[12740]_ );
  assign \new_[12252]_  = (~\new_[13660]_  | ~\new_[12842]_ ) & (~\new_[13191]_  | ~\new_[12918]_ );
  assign \new_[12253]_  = ~\new_[12608]_  | ~\new_[5631]_ ;
  assign \new_[12254]_  = ~\new_[12586]_  | ~\new_[3672]_ ;
  assign \new_[12255]_  = (~\new_[12778]_  | ~\new_[13785]_ ) & (~\new_[13401]_  | ~\new_[12763]_ );
  assign \new_[12256]_  = \new_[12969]_  & \new_[3307]_ ;
  assign \new_[12257]_  = \new_[12969]_  ^ \new_[3307]_ ;
  assign \new_[12258]_  = \new_[13028]_  & \new_[3540]_ ;
  assign \new_[12259]_  = \new_[13028]_  ^ \new_[3540]_ ;
  assign \new_[12260]_  = ~\new_[13003]_  & ~\new_[12819]_ ;
  assign \new_[12261]_  = ~\new_[13004]_  & ~\new_[12819]_ ;
  assign \new_[12262]_  = ~\new_[7874]_  | ~\new_[12877]_  | ~\new_[12912]_ ;
  assign \new_[12263]_  = ~\new_[12618]_ ;
  assign \new_[12264]_  = ~\new_[12617]_ ;
  assign \new_[12265]_  = \new_[13656]_  ^ \new_[12968]_ ;
  assign \new_[12266]_  = ~\new_[13756]_  | ~\new_[12829]_ ;
  assign \new_[12267]_  = ~\new_[12554]_ ;
  assign \new_[12268]_  = ~\new_[5370]_  | ~\new_[12789]_ ;
  assign \new_[12269]_  = ~\new_[4996]_  | ~\new_[12781]_ ;
  assign \new_[12270]_  = ~\new_[5014]_  | ~\new_[12821]_ ;
  assign \new_[12271]_  = ~\new_[5728]_  | ~\new_[12789]_ ;
  assign \new_[12272]_  = ~\new_[5751]_  | ~\new_[12789]_ ;
  assign \new_[12273]_  = ~\new_[5351]_  | ~\new_[12789]_ ;
  assign \new_[12274]_  = ~\new_[5498]_  | ~\new_[12821]_ ;
  assign \new_[12275]_  = ~\new_[5514]_  | ~\new_[12781]_ ;
  assign \new_[12276]_  = ~\new_[5510]_  | ~\new_[12781]_ ;
  assign \new_[12277]_  = ~\new_[5350]_  | ~\new_[12789]_ ;
  assign \new_[12278]_  = ~\new_[5499]_  | ~\new_[12821]_ ;
  assign \new_[12279]_  = ~\new_[4974]_  | ~\new_[12830]_ ;
  assign \new_[12280]_  = ~\new_[4971]_  | ~\new_[12821]_ ;
  assign \new_[12281]_  = ~\new_[5497]_  | ~\new_[12821]_ ;
  assign \new_[12282]_  = ~\new_[5518]_  | ~\new_[12821]_ ;
  assign \new_[12283]_  = ~\new_[4990]_  | ~\new_[12821]_ ;
  assign \new_[12284]_  = ~\new_[5507]_  | ~\new_[12781]_ ;
  assign \new_[12285]_  = ~\new_[5519]_  | ~\new_[12821]_ ;
  assign \new_[12286]_  = ~\new_[5508]_  | ~\new_[12781]_ ;
  assign \new_[12287]_  = ~\new_[4995]_  | ~\new_[12821]_ ;
  assign \new_[12288]_  = ~\new_[5511]_  | ~\new_[12781]_ ;
  assign \new_[12289]_  = ~\new_[5513]_  | ~\new_[12781]_ ;
  assign \new_[12290]_  = ~\new_[5004]_  | ~\new_[12821]_ ;
  assign \new_[12291]_  = ~\new_[12505]_ ;
  assign \new_[12292]_  = ~\new_[5216]_  | ~\new_[12830]_ ;
  assign \new_[12293]_  = ~\new_[5504]_  | ~\new_[12781]_ ;
  assign \new_[12294]_  = ~\new_[4991]_  | ~\new_[12830]_ ;
  assign \new_[12295]_  = ~\new_[5198]_  | ~\new_[12830]_ ;
  assign \new_[12296]_  = ~\new_[5199]_  | ~\new_[12830]_ ;
  assign \new_[12297]_  = ~\new_[5206]_  | ~\new_[12830]_ ;
  assign \new_[12298]_  = ~\new_[4969]_  | ~\new_[12830]_ ;
  assign \new_[12299]_  = ~\new_[5204]_  | ~\new_[12830]_ ;
  assign \new_[12300]_  = ~\new_[5217]_  | ~\new_[12830]_ ;
  assign \new_[12301]_  = ~\new_[5516]_  | ~\new_[12821]_ ;
  assign \new_[12302]_  = ~\new_[13053]_  & ~\new_[12819]_ ;
  assign \new_[12303]_  = ~\new_[13046]_  & ~\new_[12819]_ ;
  assign \new_[12304]_  = \new_[12509]_ ;
  assign \new_[12305]_  = ~\new_[13020]_  & ~\new_[12819]_ ;
  assign \new_[12306]_  = ~\new_[12881]_  & ~\new_[12819]_ ;
  assign \new_[12307]_  = ~\new_[12781]_  | ~\new_[13365]_ ;
  assign \new_[12308]_  = ~\new_[12548]_ ;
  assign \new_[12309]_  = ~\new_[12883]_  | ~\new_[5635]_  | ~\new_[12796]_ ;
  assign \new_[12310]_  = ~\new_[12935]_  & ~\new_[12819]_ ;
  assign \new_[12311]_  = ~\new_[13041]_  & ~\new_[12819]_ ;
  assign \new_[12312]_  = ~\new_[12937]_  & ~\new_[12819]_ ;
  assign \new_[12313]_  = ~\new_[13270]_  | ~\new_[5727]_  | ~\new_[13990]_ ;
  assign \new_[12314]_  = ~\new_[12936]_  & ~\new_[12819]_ ;
  assign \new_[12315]_  = ~\new_[12894]_  | ~\new_[5590]_  | ~\new_[12893]_ ;
  assign \new_[12316]_  = ~\new_[12939]_  & ~\new_[12819]_ ;
  assign \new_[12317]_  = ~\new_[13034]_  & ~\new_[12819]_ ;
  assign \new_[12318]_  = ~\new_[12990]_  | ~\new_[4865]_  | ~\new_[12855]_ ;
  assign \new_[12319]_  = ~\new_[13197]_  | ~\new_[13300]_  | ~\new_[7976]_ ;
  assign \new_[12320]_  = ~\new_[12959]_  & ~\new_[4633]_ ;
  assign \new_[12321]_  = ~\new_[12884]_  & ~\new_[12819]_ ;
  assign \new_[12322]_  = ~\new_[12686]_ ;
  assign \new_[12323]_  = ~\new_[13054]_  & ~\new_[12819]_ ;
  assign \new_[12324]_  = ~\new_[12910]_  & ~\new_[12819]_ ;
  assign \new_[12325]_  = ~\new_[12517]_ ;
  assign \new_[12326]_  = ~\new_[12913]_  & ~\new_[12819]_ ;
  assign \new_[12327]_  = ~\new_[13026]_  & ~\new_[12819]_ ;
  assign \new_[12328]_  = ~\new_[13008]_  & ~\new_[12819]_ ;
  assign \new_[12329]_  = ~\new_[12519]_ ;
  assign \new_[12330]_  = ~\new_[12519]_ ;
  assign \new_[12331]_  = ~\new_[12739]_  & ~\new_[12819]_ ;
  assign \new_[12332]_  = ~\new_[12938]_  & ~\new_[12819]_ ;
  assign \new_[12333]_  = ~\new_[13197]_  | ~\new_[7973]_  | ~\new_[13455]_ ;
  assign \new_[12334]_  = ~\new_[13042]_  & ~\new_[12819]_ ;
  assign \new_[12335]_  = ~\new_[13060]_  & ~\new_[12819]_ ;
  assign \new_[12336]_  = ~\new_[12941]_  & ~\new_[12819]_ ;
  assign \new_[12337]_  = \new_[13952]_  | \new_[13622]_ ;
  assign \new_[12338]_  = ~\new_[12999]_  & ~\new_[12819]_ ;
  assign \new_[12339]_  = ~\new_[12989]_  & ~\new_[12819]_ ;
  assign \new_[12340]_  = ~\new_[12742]_  | ~\new_[12749]_ ;
  assign \new_[12341]_  = \new_[14173]_ ;
  assign \new_[12342]_  = ~\new_[12851]_  | ~\new_[12797]_ ;
  assign \new_[12343]_  = \new_[12785]_  | \new_[12959]_ ;
  assign \new_[12344]_  = (~\new_[13857]_  | ~\new_[13461]_ ) & (~\new_[2756]_  | ~\new_[4757]_ );
  assign \new_[12345]_  = (~\new_[13365]_  | ~\new_[13791]_ ) & (~\new_[2759]_  | ~\new_[4760]_ );
  assign \new_[12346]_  = ~\new_[12852]_  & (~\new_[4640]_  | ~\new_[13650]_ );
  assign \new_[12347]_  = ~\new_[12775]_  & (~\new_[7495]_  | ~\new_[3081]_ );
  assign \new_[12348]_  = ~\new_[12499]_ ;
  assign \new_[12349]_  = \new_[7492]_  ^ \new_[13096]_ ;
  assign \new_[12350]_  = \new_[13190]_  ^ \new_[13738]_ ;
  assign \new_[12351]_  = ~\new_[12897]_  & ~\new_[12819]_ ;
  assign \new_[12352]_  = ~\new_[12504]_ ;
  assign \new_[12353]_  = ~\new_[12504]_ ;
  assign \new_[12354]_  = ~\new_[12502]_ ;
  assign \new_[12355]_  = ~\new_[12508]_ ;
  assign \new_[12356]_  = ~\new_[12508]_ ;
  assign \new_[12357]_  = ~\new_[12508]_ ;
  assign \new_[12358]_  = ~\new_[12508]_ ;
  assign \new_[12359]_  = ~\new_[12508]_ ;
  assign \new_[12360]_  = ~\new_[12643]_ ;
  assign \new_[12361]_  = ~\new_[12643]_ ;
  assign \new_[12362]_  = ~\new_[12509]_ ;
  assign \new_[12363]_  = ~\new_[14145]_ ;
  assign \new_[12364]_  = ~\new_[12640]_ ;
  assign \new_[12365]_  = ~\new_[12640]_ ;
  assign \new_[12366]_  = ~\new_[12990]_  & ~\new_[13161]_ ;
  assign \new_[12367]_  = ~\new_[12998]_  & ~\new_[12819]_ ;
  assign \new_[12368]_  = ~\new_[12883]_  & ~\new_[13092]_ ;
  assign \new_[12369]_  = ~\new_[12894]_  & ~\new_[13124]_ ;
  assign \new_[12370]_  = ~\new_[13869]_  & ~\new_[13158]_ ;
  assign \new_[12371]_  = ~\new_[12688]_ ;
  assign \new_[12372]_  = ~\new_[13869]_  | ~\new_[5615]_  | ~\new_[12799]_ ;
  assign \new_[12373]_  = ~\new_[12934]_  & ~\new_[12819]_ ;
  assign \new_[12374]_  = ~\new_[12640]_ ;
  assign \new_[12375]_  = ~\new_[12671]_ ;
  assign \new_[12376]_  = ~\new_[12671]_ ;
  assign \new_[12377]_  = ~\new_[12671]_ ;
  assign \new_[12378]_  = ~\new_[12534]_ ;
  assign \new_[12379]_  = ~\new_[12588]_ ;
  assign \new_[12380]_  = \new_[12590]_ ;
  assign \new_[12381]_  = ~\new_[12657]_ ;
  assign \new_[12382]_  = ~\new_[13112]_  | ~\wb_addr_i[4] ;
  assign \new_[12383]_  = ~\new_[14155]_ ;
  assign \new_[12384]_  = ~\new_[12514]_ ;
  assign \new_[12385]_  = ~\new_[5500]_  | ~\new_[12781]_ ;
  assign \new_[12386]_  = ~\new_[4997]_  | ~\new_[12781]_ ;
  assign \new_[12387]_  = ~\new_[5496]_  | ~\new_[12821]_ ;
  assign \new_[12388]_  = ~\new_[5214]_  | ~\new_[12830]_ ;
  assign \new_[12389]_  = ~\new_[12593]_ ;
  assign \new_[12390]_  = ~\new_[5501]_  | ~\new_[12781]_ ;
  assign \new_[12391]_  = ~\new_[12526]_ ;
  assign \new_[12392]_  = \new_[13823]_  | \new_[12811]_ ;
  assign \new_[12393]_  = ~\new_[12524]_ ;
  assign \new_[12394]_  = \new_[13769]_  | \new_[12710]_ ;
  assign \new_[12395]_  = ~\new_[12613]_ ;
  assign \new_[12396]_  = ~\new_[12727]_ ;
  assign \new_[12397]_  = ~\new_[12644]_ ;
  assign \new_[12398]_  = ~\new_[5503]_  | ~\new_[12821]_ ;
  assign \new_[12399]_  = ~\new_[12664]_ ;
  assign \new_[12400]_  = \new_[13824]_  | \new_[12853]_ ;
  assign \new_[12401]_  = ~\new_[5495]_  | ~\new_[12821]_ ;
  assign \new_[12402]_  = ~\new_[12519]_ ;
  assign \new_[12403]_  = ~\new_[12519]_ ;
  assign \new_[12404]_  = ~\new_[12519]_ ;
  assign \new_[12405]_  = ~\new_[5203]_  | ~\new_[12830]_ ;
  assign \new_[12406]_  = ~\new_[5003]_  | ~\new_[12781]_ ;
  assign \new_[12407]_  = ~\new_[13330]_  | ~\new_[12793]_ ;
  assign \new_[12408]_  = ~\new_[13217]_  | ~\new_[12839]_ ;
  assign \new_[12409]_  = ~\new_[12686]_ ;
  assign \new_[12410]_  = ~\new_[5348]_  | ~\new_[12789]_ ;
  assign \new_[12411]_  = ~\new_[5506]_  | ~\new_[12781]_ ;
  assign \new_[12412]_  = ~\new_[5730]_  | ~\new_[12789]_ ;
  assign \new_[12413]_  = ~\new_[5368]_  | ~\new_[12789]_ ;
  assign \new_[12414]_  = ~\new_[5353]_  | ~\new_[12789]_ ;
  assign \new_[12415]_  = ~\new_[5738]_  | ~\new_[12789]_ ;
  assign \new_[12416]_  = ~\new_[5743]_  | ~\new_[12789]_ ;
  assign \new_[12417]_  = ~\new_[12671]_ ;
  assign \new_[12418]_  = ~\new_[5509]_  | ~\new_[12781]_ ;
  assign \new_[12419]_  = ~\new_[5369]_  | ~\new_[12789]_ ;
  assign \new_[12420]_  = ~\new_[5371]_  | ~\new_[12789]_ ;
  assign \new_[12421]_  = ~\new_[5349]_  | ~\new_[12789]_ ;
  assign \new_[12422]_  = ~\new_[5347]_  | ~\new_[12789]_ ;
  assign \new_[12423]_  = ~\new_[5218]_  | ~\new_[12830]_ ;
  assign \new_[12424]_  = ~\new_[12923]_  & ~\new_[12819]_ ;
  assign \new_[12425]_  = ~\new_[12633]_ ;
  assign \new_[12426]_  = ~\new_[14037]_  | ~\new_[5605]_  | ~\new_[12892]_ ;
  assign \new_[12427]_  = (~\new_[12982]_  | ~\new_[13458]_ ) & (~\new_[13487]_  | ~\new_[13011]_ );
  assign \new_[12428]_  = ~\new_[12640]_ ;
  assign \new_[12429]_  = ~\new_[12816]_ ;
  assign \new_[12430]_  = ~\new_[12528]_ ;
  assign \new_[12431]_  = \new_[14173]_ ;
  assign \new_[12432]_  = ~\new_[12652]_ ;
  assign \new_[12433]_  = ~\new_[12822]_ ;
  assign \new_[12434]_  = ~\new_[12726]_ ;
  assign \new_[12435]_  = \new_[13867]_  | \new_[13316]_ ;
  assign \new_[12436]_  = ~\new_[12826]_ ;
  assign \new_[12437]_  = ~\new_[13971]_ ;
  assign \new_[12438]_  = \new_[13320]_  | \new_[12718]_ ;
  assign \new_[12439]_  = ~\new_[13112]_  | ~\new_[13109]_ ;
  assign \new_[12440]_  = ~\new_[12590]_ ;
  assign \new_[12441]_  = ~\new_[12659]_ ;
  assign \new_[12442]_  = ~\new_[12588]_ ;
  assign \new_[12443]_  = ~\new_[12588]_ ;
  assign \new_[12444]_  = ~\new_[12588]_ ;
  assign \new_[12445]_  = ~\new_[12588]_ ;
  assign \new_[12446]_  = ~\new_[12534]_ ;
  assign \new_[12447]_  = \new_[13896]_ ;
  assign \new_[12448]_  = ~\new_[12584]_ ;
  assign \new_[12449]_  = ~\new_[12640]_ ;
  assign \new_[12450]_  = (~\new_[12982]_  | ~\new_[13466]_ ) & (~\new_[13590]_  | ~\new_[13011]_ );
  assign \new_[12451]_  = \new_[4763]_  ^ \new_[13989]_ ;
  assign \new_[12452]_  = ~\new_[12870]_  | ~\new_[12849]_ ;
  assign \new_[12453]_  = ~\new_[12858]_  | ~\new_[2786]_ ;
  assign \new_[12454]_  = \new_[12993]_ ;
  assign \new_[12455]_  = ~\new_[13538]_  | ~\new_[12714]_  | ~\wb_addr_i[6] ;
  assign \new_[12456]_  = \new_[12867]_  & \new_[12713]_ ;
  assign \new_[12457]_  = ~\new_[12905]_  & ~\new_[12819]_ ;
  assign \new_[12458]_  = ~\new_[12686]_ ;
  assign \new_[12459]_  = ~\new_[12688]_ ;
  assign \new_[12460]_  = \new_[12877]_  & \new_[12912]_ ;
  assign \new_[12461]_  = ~\new_[12688]_ ;
  assign \new_[12462]_  = \new_[12875]_  & \new_[8099]_ ;
  assign \new_[12463]_  = \new_[12877]_  & \new_[7936]_ ;
  assign \new_[12464]_  = ~\new_[12688]_ ;
  assign \new_[12465]_  = ~u12_we2_reg;
  assign \new_[12466]_  = ~\new_[12688]_ ;
  assign \new_[12467]_  = ~\new_[5512]_  | ~\new_[12821]_ ;
  assign \new_[12468]_  = ~\new_[12932]_  | ~\new_[13049]_  | ~\new_[13147]_ ;
  assign \new_[12469]_  = ~\new_[12708]_ ;
  assign \new_[12470]_  = ~\new_[12738]_  & ~\new_[12819]_ ;
  assign \new_[12471]_  = ~\new_[7973]_  | ~\new_[12806]_  | ~\new_[13656]_ ;
  assign \new_[12472]_  = ~\new_[13043]_  & ~\new_[12819]_ ;
  assign \new_[12473]_  = ~\new_[12516]_ ;
  assign \new_[12474]_  = \new_[13127]_  ^ \new_[13091]_ ;
  assign \new_[12475]_  = \new_[13169]_  ^ \new_[13104]_ ;
  assign \new_[12476]_  = \new_[13105]_  ^ \new_[13151]_ ;
  assign \new_[12477]_  = ~\new_[12867]_  | ~\new_[13114]_ ;
  assign \new_[12478]_  = ~\new_[12720]_  | (~\new_[7493]_  & ~\new_[3540]_ );
  assign \new_[12479]_  = ~\new_[12825]_  | ~\new_[2786]_ ;
  assign \new_[12480]_  = ~\new_[12728]_  | ~\new_[2786]_ ;
  assign \new_[12481]_  = ~\new_[12831]_  | ~\new_[13109]_ ;
  assign \new_[12482]_  = ~\new_[12704]_ ;
  assign \new_[12483]_  = ~\wb_addr_i[6]  & (~\new_[13112]_  | ~\new_[12977]_ );
  assign \new_[12484]_  = (~\new_[13532]_  | ~\new_[13482]_ ) & (~\new_[2758]_  | ~\new_[4754]_ );
  assign \new_[12485]_  = ~\new_[7976]_  | ~\new_[7972]_  | ~\new_[12968]_  | ~\new_[12970]_ ;
  assign \new_[12486]_  = (~\new_[12982]_  | ~\new_[13373]_ ) & (~\new_[13360]_  | ~\new_[13011]_ );
  assign \new_[12487]_  = (~\new_[12982]_  | ~\new_[13565]_ ) & (~\new_[13691]_  | ~\new_[13011]_ );
  assign \new_[12488]_  = (~\new_[12982]_  | ~\new_[13326]_ ) & (~\new_[13311]_  | ~\new_[13011]_ );
  assign \new_[12489]_  = (~\new_[12982]_  | ~\new_[13841]_ ) & (~\new_[13313]_  | ~\new_[13011]_ );
  assign \new_[12490]_  = (~\new_[12982]_  | ~\new_[13732]_ ) & (~\new_[13578]_  | ~\new_[13011]_ );
  assign \new_[12491]_  = (~\new_[12982]_  | ~\new_[13725]_ ) & (~\new_[13572]_  | ~\new_[13011]_ );
  assign \new_[12492]_  = (~\new_[12982]_  | ~\new_[13735]_ ) & (~\new_[13325]_  | ~\new_[13011]_ );
  assign \new_[12493]_  = (~\new_[12982]_  | ~\new_[13393]_ ) & (~\new_[13511]_  | ~\new_[13011]_ );
  assign \new_[12494]_  = (~\new_[12982]_  | ~\new_[13673]_ ) & (~\new_[13557]_  | ~\new_[13011]_ );
  assign \new_[12495]_  = (~\new_[12982]_  | ~\new_[13625]_ ) & (~\new_[13536]_  | ~\new_[13011]_ );
  assign \new_[12496]_  = (~\new_[12982]_  | ~\new_[13221]_ ) & (~\new_[13502]_  | ~\new_[13011]_ );
  assign \new_[12497]_  = \new_[13100]_  & \new_[13096]_ ;
  assign \new_[12498]_  = \new_[13100]_  ^ \new_[13096]_ ;
  assign \new_[12499]_  = ~\wb_addr_i[4]  | ~\new_[13036]_  | ~\wb_addr_i[3] ;
  assign \new_[12500]_  = ~\new_[12722]_ ;
  assign \new_[12501]_  = ~\new_[12869]_ ;
  assign \new_[12502]_  = ~\new_[14182]_ ;
  assign \new_[12503]_  = ~u2_bit_clk_r1_reg;
  assign \new_[12504]_  = ~\new_[12712]_ ;
  assign \new_[12505]_  = \new_[12970]_  & \new_[7935]_ ;
  assign \new_[12506]_  = ~\new_[12968]_  | ~\new_[7979]_ ;
  assign \new_[12507]_  = \new_[13455]_  & \new_[12907]_ ;
  assign \new_[12508]_  = ~\new_[12812]_ ;
  assign \new_[12509]_  = \new_[13015]_  & \wb_addr_i[4] ;
  assign \new_[12510]_  = ~\new_[12996]_  & ~\new_[13013]_ ;
  assign \new_[12511]_  = ~\new_[12926]_  | ~\new_[13109]_ ;
  assign \new_[12512]_  = ~\new_[3213]_  & ~\new_[13059]_ ;
  assign \new_[12513]_  = ~\new_[12726]_ ;
  assign \new_[12514]_  = ~\new_[14153]_ ;
  assign \new_[12515]_  = ~\new_[3482]_  & ~\new_[13059]_ ;
  assign \new_[12516]_  = ~\new_[13015]_  | ~\new_[13109]_ ;
  assign \new_[12517]_  = ~\new_[12886]_ ;
  assign \new_[12518]_  = ~\new_[3283]_  & ~\new_[13056]_ ;
  assign \new_[12519]_  = ~\new_[14093]_ ;
  assign \new_[12520]_  = ~\new_[13796]_  | ~\new_[13726]_  | ~\new_[7807]_ ;
  assign \new_[12521]_  = ~\new_[12841]_ ;
  assign \new_[12522]_  = \new_[7972]_  & \new_[12907]_ ;
  assign \new_[12523]_  = ~\new_[3286]_  & ~\new_[13056]_ ;
  assign \new_[12524]_  = ~\new_[12786]_ ;
  assign \new_[12525]_  = ~\new_[12798]_ ;
  assign \new_[12526]_  = ~\new_[12784]_ ;
  assign \new_[12527]_  = ~\new_[12889]_  & ~\new_[12967]_ ;
  assign \new_[12528]_  = ~\new_[12817]_ ;
  assign \new_[12529]_  = ~\new_[12782]_ ;
  assign \new_[12530]_  = ~\new_[13188]_  & ~\new_[12991]_ ;
  assign \new_[12531]_  = \new_[3771]_  ^ \new_[13141]_ ;
  assign n10996 = \new_[12045]_  ? \new_[4412]_  : \new_[7500]_ ;
  assign \new_[12533]_  = ~\new_[12831]_ ;
  assign \new_[12534]_  = ~\new_[12835]_ ;
  assign \new_[12535]_  = ~\new_[12924]_  & ~\new_[12951]_ ;
  assign n11056 = \new_[13083]_  ^ \new_[14037]_ ;
  assign n11061 = \new_[13190]_  ^ \new_[4689]_ ;
  assign n11051 = \new_[12075]_  ? \new_[4412]_  : \new_[4672]_ ;
  assign n10981 = \new_[11528]_  ? \new_[4412]_  : \new_[4578]_ ;
  assign n11041 = \new_[12066]_  ? \new_[4412]_  : \new_[6793]_ ;
  assign n10991 = \new_[12020]_  ? \new_[4412]_  : \new_[2746]_ ;
  assign n11036 = \new_[12065]_  ? \new_[4412]_  : \new_[2735]_ ;
  assign \new_[12543]_  = ~\new_[12715]_ ;
  assign \new_[12544]_  = ~\new_[12854]_ ;
  assign \new_[12545]_  = \new_[3587]_  ^ \new_[3306]_ ;
  assign \new_[12546]_  = ~\new_[12715]_ ;
  assign \new_[12547]_  = \new_[7493]_  ^ \new_[3540]_ ;
  assign \new_[12548]_  = ~\new_[12926]_  | ~\wb_addr_i[4] ;
  assign \new_[12549]_  = ~\new_[12883]_ ;
  assign \new_[12550]_  = ~\new_[12798]_ ;
  assign \new_[12551]_  = ~\new_[12798]_ ;
  assign \new_[12552]_  = ~\new_[12798]_ ;
  assign \new_[12553]_  = \new_[12712]_ ;
  assign \new_[12554]_  = \new_[12712]_ ;
  assign \new_[12555]_  = ~\new_[12746]_ ;
  assign \new_[12556]_  = ~\new_[12746]_ ;
  assign \new_[12557]_  = ~\new_[12746]_ ;
  assign \new_[12558]_  = ~\new_[12746]_ ;
  assign \new_[12559]_  = ~\new_[12746]_ ;
  assign \new_[12560]_  = ~\new_[12707]_ ;
  assign \new_[12561]_  = ~\new_[12715]_ ;
  assign \new_[12562]_  = ~\new_[12715]_ ;
  assign \new_[12563]_  = ~\new_[12715]_ ;
  assign \new_[12564]_  = ~\new_[12715]_ ;
  assign \new_[12565]_  = ~\new_[12800]_ ;
  assign \new_[12566]_  = ~\new_[12800]_ ;
  assign \new_[12567]_  = ~\new_[12800]_ ;
  assign \new_[12568]_  = ~\new_[12751]_ ;
  assign \new_[12569]_  = ~\new_[12804]_ ;
  assign \new_[12570]_  = ~\new_[12804]_ ;
  assign \new_[12571]_  = ~\new_[13546]_  | ~\new_[12991]_ ;
  assign \new_[12572]_  = ~\new_[12864]_ ;
  assign \new_[12573]_  = ~\new_[12800]_ ;
  assign \new_[12574]_  = ~\new_[12845]_ ;
  assign \new_[12575]_  = ~\new_[13714]_  | ~\new_[13141]_ ;
  assign \new_[12576]_  = ~\new_[12800]_ ;
  assign \new_[12577]_  = \new_[12850]_ ;
  assign \new_[12578]_  = ~\new_[12857]_ ;
  assign \new_[12579]_  = ~\new_[12860]_ ;
  assign \new_[12580]_  = ~\new_[13828]_  | ~\new_[3081]_ ;
  assign \new_[12581]_  = ~\new_[12753]_ ;
  assign \new_[12582]_  = \new_[12743]_ ;
  assign \new_[12583]_  = ~\new_[12762]_ ;
  assign \new_[12584]_  = ~\new_[12836]_ ;
  assign \new_[12585]_  = \new_[12835]_ ;
  assign \new_[12586]_  = ~\new_[12732]_ ;
  assign \new_[12587]_  = \new_[12834]_ ;
  assign \new_[12588]_  = ~\new_[12834]_ ;
  assign \new_[12589]_  = \new_[12833]_ ;
  assign \new_[12590]_  = ~\new_[12731]_ ;
  assign \new_[12591]_  = ~\new_[12832]_ ;
  assign \new_[12592]_  = \new_[13574]_  | \new_[14093]_ ;
  assign \new_[12593]_  = ~\new_[14119]_ ;
  assign \new_[12594]_  = ~\new_[12729]_ ;
  assign \new_[12595]_  = \new_[12829]_ ;
  assign \new_[12596]_  = ~\new_[13656]_  | ~\new_[13403]_ ;
  assign \new_[12597]_  = ~\new_[12751]_ ;
  assign \new_[12598]_  = ~\new_[12827]_ ;
  assign \new_[12599]_  = ~\new_[14087]_ ;
  assign \new_[12600]_  = ~\new_[13480]_  & ~\new_[13455]_ ;
  assign \new_[12601]_  = ~\new_[12823]_ ;
  assign \new_[12602]_  = ~\new_[12714]_ ;
  assign \new_[12603]_  = ~\new_[12919]_ ;
  assign \new_[12604]_  = ~\new_[12815]_ ;
  assign \new_[12605]_  = \new_[13874]_  | \new_[13314]_ ;
  assign \new_[12606]_  = ~\new_[12814]_ ;
  assign \new_[12607]_  = ~\new_[12724]_ ;
  assign \new_[12608]_  = \new_[12807]_ ;
  assign \new_[12609]_  = ~\new_[7492]_  | ~\new_[13096]_ ;
  assign \new_[12610]_  = ~\new_[14119]_ ;
  assign \new_[12611]_  = \new_[12784]_ ;
  assign \new_[12612]_  = \new_[13877]_  | \new_[13810]_ ;
  assign \new_[12613]_  = ~\new_[12788]_ ;
  assign \new_[12614]_  = ~\new_[12957]_  & ~\new_[7979]_ ;
  assign \new_[12615]_  = ~\new_[14104]_ ;
  assign \new_[12616]_  = ~\new_[12787]_ ;
  assign \new_[12617]_  = ~\new_[12847]_ ;
  assign \new_[12618]_  = \new_[12847]_ ;
  assign \new_[12619]_  = ~\new_[12798]_ ;
  assign \new_[12620]_  = \new_[12959]_  | \new_[13747]_ ;
  assign \new_[12621]_  = ~\new_[12751]_ ;
  assign \new_[12622]_  = \new_[13575]_  | \new_[13168]_ ;
  assign \new_[12623]_  = ~\new_[12990]_ ;
  assign \new_[12624]_  = ~\new_[12804]_ ;
  assign \new_[12625]_  = ~\new_[12804]_ ;
  assign \new_[12626]_  = ~\new_[12719]_ ;
  assign \new_[12627]_  = \new_[12978]_  & \new_[13769]_ ;
  assign \new_[12628]_  = ~\new_[12715]_ ;
  assign \new_[12629]_  = ~\new_[13079]_ ;
  assign \new_[12630]_  = \new_[7497]_  ^ \new_[13145]_ ;
  assign \new_[12631]_  = ~\new_[12804]_ ;
  assign \new_[12632]_  = ~\new_[5085]_  & ~\new_[13459]_ ;
  assign \new_[12633]_  = ~\new_[12807]_ ;
  assign n11016 = \new_[12058]_  ? \new_[4412]_  : \new_[2715]_ ;
  assign \new_[12635]_  = \new_[12807]_ ;
  assign \new_[12636]_  = ~\new_[13027]_  & ~\new_[13758]_ ;
  assign \new_[12637]_  = ~\new_[13038]_  & ~\new_[13456]_ ;
  assign \new_[12638]_  = ~\new_[13070]_  & ~\new_[13457]_ ;
  assign \new_[12639]_  = \new_[12850]_ ;
  assign \new_[12640]_  = ~\new_[12850]_ ;
  assign \new_[12641]_  = \new_[7439]_  ^ \new_[13101]_ ;
  assign \new_[12642]_  = ~\new_[12813]_ ;
  assign \new_[12643]_  = ~\new_[14114]_ ;
  assign \new_[12644]_  = ~\new_[12861]_ ;
  assign \new_[12645]_  = ~\new_[12757]_ ;
  assign n11046 = \new_[12069]_  ? \new_[4412]_  : \new_[7656]_ ;
  assign \new_[12647]_  = \new_[12816]_ ;
  assign \new_[12648]_  = ~\new_[12783]_ ;
  assign \new_[12649]_  = \new_[12817]_ ;
  assign \new_[12650]_  = ~\new_[12919]_ ;
  assign \new_[12651]_  = ~\new_[12781]_ ;
  assign \new_[12652]_  = ~\new_[12780]_ ;
  assign \new_[12653]_  = \new_[12822]_ ;
  assign \new_[12654]_  = ~\new_[12726]_ ;
  assign \new_[12655]_  = \new_[12826]_ ;
  assign \new_[12656]_  = ~\new_[7496]_  & ~\new_[13141]_ ;
  assign \new_[12657]_  = ~\new_[12776]_ ;
  assign \new_[12658]_  = ~\new_[12954]_  & ~\new_[7975]_ ;
  assign \new_[12659]_  = ~\new_[12833]_ ;
  assign \new_[12660]_  = \new_[12834]_ ;
  assign n11066 = \new_[12104]_  ? \new_[4412]_  : \new_[5854]_ ;
  assign \new_[12662]_  = ~\new_[12771]_ ;
  assign \new_[12663]_  = ~\new_[12838]_ ;
  assign \new_[12664]_  = ~\new_[12795]_ ;
  assign \new_[12665]_  = ~\new_[12843]_ ;
  assign \new_[12666]_  = \new_[7438]_  ^ \new_[13131]_ ;
  assign \new_[12667]_  = ~\new_[12764]_ ;
  assign n11026 = \new_[12060]_  ? \new_[4412]_  : \new_[3762]_ ;
  assign n11021 = \new_[12059]_  ? \new_[4412]_  : \new_[4814]_ ;
  assign \new_[12670]_  = ~\new_[12944]_  & ~\new_[4755]_ ;
  assign \new_[12671]_  = ~\new_[12840]_ ;
  assign \new_[12672]_  = \new_[14037]_  ^ \new_[13425]_ ;
  assign n11011 = \new_[12057]_  ? \new_[4412]_  : \new_[2925]_ ;
  assign n11006 = \new_[12051]_  ? \new_[4412]_  : \new_[2724]_ ;
  assign n11031 = \new_[12062]_  ? \new_[4412]_  : \new_[2788]_ ;
  assign \new_[12676]_  = \new_[12786]_ ;
  assign n10986 = \new_[11710]_  ? \new_[4412]_  : \new_[3183]_ ;
  assign \new_[12678]_  = ~\new_[12736]_ ;
  assign \new_[12679]_  = \new_[12795]_ ;
  assign \new_[12680]_  = \new_[2952]_  ^ \new_[13150]_ ;
  assign \new_[12681]_  = \new_[12812]_ ;
  assign \new_[12682]_  = ~\new_[13065]_  | ~\new_[2786]_ ;
  assign n11001 = \new_[12048]_  ? \new_[4412]_  : \new_[4408]_ ;
  assign \new_[12684]_  = ~\new_[13002]_  | ~\new_[2786]_ ;
  assign \new_[12685]_  = ~\new_[12856]_ ;
  assign \new_[12686]_  = ~\new_[13168]_ ;
  assign \new_[12687]_  = ~\new_[12757]_ ;
  assign \new_[12688]_  = ~\new_[12743]_ ;
  assign \new_[12689]_  = \new_[12812]_ ;
  assign \new_[12690]_  = ~\new_[12757]_ ;
  assign \new_[12691]_  = ~\new_[12710]_ ;
  assign \new_[12692]_  = \new_[12788]_ ;
  assign \new_[12693]_  = \new_[12743]_ ;
  assign \new_[12694]_  = ~\new_[4642]_  & ~\new_[12925]_ ;
  assign n11071 = \\u1_sr_reg[0] ;
  assign \new_[12696]_  = ~\new_[12767]_ ;
  assign \new_[12697]_  = ~\new_[12746]_ ;
  assign \new_[12698]_  = ~\new_[12894]_ ;
  assign \new_[12699]_  = ~\new_[13016]_  | ~\new_[2786]_ ;
  assign \new_[12700]_  = ~\new_[13080]_  | ~\new_[2786]_ ;
  assign \new_[12701]_  = ~\new_[13074]_  | ~\new_[2786]_ ;
  assign \new_[12702]_  = ~\new_[13063]_  | ~\new_[2786]_ ;
  assign \new_[12703]_  = ~\new_[12746]_ ;
  assign \new_[12704]_  = ~\new_[9653]_  | ~\new_[13044]_  | ~\new_[13114]_ ;
  assign \new_[12705]_  = ~\new_[3285]_  & ~\new_[13056]_ ;
  assign \new_[12706]_  = \new_[12794]_ ;
  assign \new_[12707]_  = ~\new_[13001]_ ;
  assign \new_[12708]_  = ~\new_[12794]_ ;
  assign \new_[12709]_  = ~\new_[13149]_  & (~\new_[2791]_  | ~\new_[4768]_ );
  assign \new_[12710]_  = ~\new_[13017]_ ;
  assign \new_[12711]_  = \new_[13081]_ ;
  assign \new_[12712]_  = ~\new_[12943]_ ;
  assign \new_[12713]_  = \new_[13148]_  & wb_cyc_i;
  assign \new_[12714]_  = \new_[13103]_  & \new_[13109]_ ;
  assign \new_[12715]_  = ~\new_[12908]_ ;
  assign \new_[12716]_  = \new_[12996]_ ;
  assign \new_[12717]_  = ~\new_[14127]_ ;
  assign \new_[12718]_  = ~\new_[12886]_ ;
  assign \new_[12719]_  = ~\new_[12996]_ ;
  assign \new_[12720]_  = ~\new_[7493]_  | ~\new_[3540]_ ;
  assign \new_[12721]_  = ~\new_[7791]_  & ~\new_[4412]_ ;
  assign \new_[12722]_  = ~\new_[13103]_  | ~\wb_addr_i[4] ;
  assign \new_[12723]_  = ~\new_[12979]_ ;
  assign \new_[12724]_  = ~\new_[13014]_ ;
  assign \new_[12725]_  = ~\new_[5085]_  & ~\new_[5084]_ ;
  assign \new_[12726]_  = \new_[4070]_  & \new_[3540]_ ;
  assign \new_[12727]_  = ~\new_[13040]_ ;
  assign \new_[12728]_  = ~\new_[6440]_  & (~\new_[5074]_  | ~\new_[13570]_ );
  assign \new_[12729]_  = \new_[12961]_ ;
  assign \new_[12730]_  = ~\new_[5078]_  & ~\new_[13308]_ ;
  assign \new_[12731]_  = ~\new_[5069]_  | ~\new_[13818]_ ;
  assign \new_[12732]_  = ~\new_[13797]_  | ~\new_[13098]_ ;
  assign \new_[12733]_  = \new_[12889]_ ;
  assign \new_[12734]_  = ~\new_[5071]_  & ~\new_[13523]_ ;
  assign \new_[12735]_  = ~\new_[13178]_  & (~\new_[2793]_  | ~\new_[4759]_ );
  assign \new_[12736]_  = ~\new_[13050]_ ;
  assign \new_[12737]_  = ~\new_[5845]_  | ~\new_[13460]_ ;
  assign \new_[12738]_  = ~\new_[13123]_ ;
  assign \new_[12739]_  = ~\new_[13132]_ ;
  assign \new_[12740]_  = ~\new_[12906]_ ;
  assign \new_[12741]_  = \new_[13064]_ ;
  assign \new_[12742]_  = \new_[12950]_ ;
  assign \new_[12743]_  = ~\new_[13161]_  | ~\new_[13606]_ ;
  assign \new_[12744]_  = ~\new_[5078]_  | ~\new_[13308]_ ;
  assign \new_[12745]_  = \new_[13081]_ ;
  assign \new_[12746]_  = ~\new_[13081]_ ;
  assign \new_[12747]_  = \new_[13001]_ ;
  assign \new_[12748]_  = \new_[12908]_ ;
  assign \new_[12749]_  = \new_[12976]_ ;
  assign \new_[12750]_  = ~\new_[5095]_  | ~\new_[13695]_ ;
  assign \new_[12751]_  = ~\new_[12976]_ ;
  assign \new_[12752]_  = ~\new_[5850]_  | ~\new_[13604]_ ;
  assign \new_[12753]_  = ~\new_[13701]_  | ~\new_[13108]_ ;
  assign \new_[12754]_  = ~\new_[5059]_  & ~\new_[13783]_ ;
  assign \new_[12755]_  = ~\new_[5059]_  | ~\new_[13783]_ ;
  assign \new_[12756]_  = \new_[12948]_ ;
  assign \new_[12757]_  = ~\new_[13066]_ ;
  assign \new_[12758]_  = \new_[13013]_ ;
  assign \new_[12759]_  = \new_[13064]_ ;
  assign \new_[12760]_  = \new_[12967]_ ;
  assign \new_[12761]_  = ~\new_[13677]_  | ~\new_[13142]_ ;
  assign \new_[12762]_  = ~\new_[13481]_  | ~\new_[5767]_ ;
  assign \new_[12763]_  = ~\new_[13059]_ ;
  assign \new_[12764]_  = ~\new_[13155]_  | ~\new_[13801]_ ;
  assign \new_[12765]_  = ~\new_[5095]_  & ~\new_[13695]_ ;
  assign \new_[12766]_  = ~\new_[5066]_  & ~\new_[13539]_ ;
  assign \new_[12767]_  = ~\new_[13157]_  | ~\new_[13700]_ ;
  assign \new_[12768]_  = ~\new_[13425]_  | ~\new_[13113]_ ;
  assign \new_[12769]_  = \new_[12976]_ ;
  assign \new_[12770]_  = ~\new_[5085]_  | ~\new_[13459]_ ;
  assign \new_[12771]_  = ~\new_[12889]_ ;
  assign \new_[12772]_  = ~\new_[5850]_  & ~\new_[13604]_ ;
  assign \new_[12773]_  = ~\new_[13190]_  & ~\new_[4689]_ ;
  assign \new_[12774]_  = ~\new_[13035]_ ;
  assign \new_[12775]_  = ~\new_[7495]_  & ~\new_[3081]_ ;
  assign \new_[12776]_  = ~\new_[12958]_ ;
  assign \new_[12777]_  = ~\new_[13030]_ ;
  assign \new_[12778]_  = ~\new_[13029]_ ;
  assign \new_[12779]_  = \new_[13076]_ ;
  assign \new_[12780]_  = ~\new_[3306]_  | ~\new_[3307]_ ;
  assign \new_[12781]_  = \new_[12891]_ ;
  assign \new_[12782]_  = ~\new_[14186]_ ;
  assign \new_[12783]_  = ~\new_[14184]_ ;
  assign \new_[12784]_  = ~\new_[12911]_ ;
  assign \new_[12785]_  = ~\new_[4642]_  | ~\new_[4633]_ ;
  assign \new_[12786]_  = ~\new_[12952]_ ;
  assign \new_[12787]_  = ~\new_[12953]_ ;
  assign \new_[12788]_  = ~\new_[12909]_ ;
  assign \new_[12789]_  = \new_[13040]_ ;
  assign \new_[12790]_  = \new_[12908]_ ;
  assign \new_[12791]_  = \new_[12950]_ ;
  assign \new_[12792]_  = ~\new_[13953]_ ;
  assign \new_[12793]_  = ~\new_[13010]_ ;
  assign \new_[12794]_  = ~\new_[12904]_ ;
  assign \new_[12795]_  = ~\new_[12986]_ ;
  assign \new_[12796]_  = ~\new_[13151]_ ;
  assign \new_[12797]_  = \new_[13066]_ ;
  assign \new_[12798]_  = ~\new_[12950]_ ;
  assign \new_[12799]_  = ~\new_[13104]_ ;
  assign \new_[12800]_  = ~\new_[13064]_ ;
  assign \new_[12801]_  = ~\new_[5071]_  | ~\new_[13523]_ ;
  assign n11076 = \new_[13120]_  & \new_[13148]_ ;
  assign \new_[12803]_  = \new_[12948]_ ;
  assign \new_[12804]_  = ~\new_[12948]_ ;
  assign \new_[12805]_  = ~\new_[12945]_ ;
  assign \new_[12806]_  = ~\new_[13480]_  & ~\new_[7935]_ ;
  assign \new_[12807]_  = ~\new_[13078]_ ;
  assign \new_[12808]_  = ~\new_[13005]_ ;
  assign \new_[12809]_  = ~\new_[13006]_ ;
  assign \new_[12810]_  = ~\new_[13007]_ ;
  assign \new_[12811]_  = ~\new_[13012]_ ;
  assign \new_[12812]_  = ~\new_[13180]_  | ~\new_[13379]_ ;
  assign \new_[12813]_  = ~\new_[13013]_ ;
  assign \new_[12814]_  = ~\new_[13009]_ ;
  assign \new_[12815]_  = ~\new_[13077]_ ;
  assign \new_[12816]_  = ~\new_[3081]_  & ~\new_[13096]_ ;
  assign \new_[12817]_  = ~\new_[13021]_ ;
  assign \new_[12818]_  = ~\new_[12888]_ ;
  assign \new_[12819]_  = ~\new_[12888]_ ;
  assign \new_[12820]_  = ~\new_[12917]_ ;
  assign \new_[12821]_  = \new_[12891]_ ;
  assign \new_[12822]_  = ~\new_[3306]_  & ~\new_[3307]_ ;
  assign \new_[12823]_  = ~\new_[13025]_ ;
  assign \new_[12824]_  = ~\new_[13027]_ ;
  assign \new_[12825]_  = ~\new_[5859]_  & (~\new_[5064]_  | ~\new_[13520]_ );
  assign \new_[12826]_  = ~\new_[13141]_  & ~\new_[3540]_ ;
  assign \new_[12827]_  = ~\new_[12920]_ ;
  assign \new_[12828]_  = ~\new_[12962]_ ;
  assign \new_[12829]_  = ~\new_[12961]_ ;
  assign \new_[12830]_  = \new_[12958]_ ;
  assign \new_[12831]_  = \new_[13084]_  & \wb_addr_i[3] ;
  assign \new_[12832]_  = \new_[5694]_  | \new_[13315]_ ;
  assign \new_[12833]_  = ~\new_[13129]_  & ~\new_[13818]_ ;
  assign \new_[12834]_  = ~\new_[13121]_  | ~\new_[13615]_ ;
  assign \new_[12835]_  = ~\new_[12890]_ ;
  assign \new_[12836]_  = ~\new_[5694]_  | ~\new_[13315]_ ;
  assign \new_[12837]_  = \new_[12924]_ ;
  assign \new_[12838]_  = ~\new_[12924]_ ;
  assign \new_[12839]_  = ~\new_[12986]_ ;
  assign \new_[12840]_  = ~\new_[13039]_ ;
  assign \new_[12841]_  = ~\new_[12899]_ ;
  assign \new_[12842]_  = ~\new_[13056]_ ;
  assign \new_[12843]_  = ~\new_[13037]_ ;
  assign \new_[12844]_  = ~\new_[13038]_ ;
  assign \new_[12845]_  = ~\new_[12951]_ ;
  assign \new_[12846]_  = \new_[3340]_  ^ \new_[3081]_ ;
  assign \new_[12847]_  = ~\new_[13010]_ ;
  assign \new_[12848]_  = ~\new_[13119]_  & (~\new_[2757]_  | ~\new_[4758]_ );
  assign \new_[12849]_  = ~\new_[13097]_  & (~\new_[7438]_  | ~\new_[3150]_ );
  assign \new_[12850]_  = ~\new_[13083]_  | ~\new_[13375]_ ;
  assign \new_[12851]_  = \new_[13050]_ ;
  assign \new_[12852]_  = ~\new_[12925]_ ;
  assign \new_[12853]_  = ~\new_[12993]_ ;
  assign \new_[12854]_  = ~\new_[13278]_  | ~\new_[13082]_ ;
  assign \new_[12855]_  = ~\new_[13091]_ ;
  assign \new_[12856]_  = ~\new_[12902]_ ;
  assign \new_[12857]_  = ~\new_[12967]_ ;
  assign \new_[12858]_  = ~\new_[5860]_  & (~\new_[5062]_  | ~\new_[13550]_ );
  assign \new_[12859]_  = ~\new_[13089]_  & (~\new_[7439]_  | ~\new_[2952]_ );
  assign \new_[12860]_  = ~\new_[13278]_  & ~\new_[13082]_ ;
  assign \new_[12861]_  = ~\new_[12980]_ ;
  assign \new_[12862]_  = ~\new_[13070]_ ;
  assign \new_[12863]_  = ~\new_[13071]_ ;
  assign \new_[12864]_  = ~\new_[13076]_ ;
  assign \new_[12865]_  = ~\new_[5845]_  & ~\new_[13460]_ ;
  assign \new_[12866]_  = \new_[13050]_ ;
  assign \new_[12867]_  = ~\new_[13165]_  & ~\wb_addr_i[30] ;
  assign \new_[12868]_  = ~\new_[13118]_  & (~\new_[7497]_  | ~\new_[3374]_ );
  assign \new_[12869]_  = \new_[13071]_ ;
  assign \new_[12870]_  = ~\new_[13116]_  | (~\new_[7494]_  & ~\new_[3307]_ );
  assign \new_[12871]_  = \new_[12951]_ ;
  assign \new_[12872]_  = ~\new_[5066]_  | ~\new_[13539]_ ;
  assign \new_[12873]_  = ~\new_[14037]_  & ~\new_[13083]_ ;
  assign \new_[12874]_  = ~\new_[13071]_ ;
  assign \new_[12875]_  = \new_[8114]_  & \new_[7956]_ ;
  assign \new_[12876]_  = \new_[8114]_  ^ \new_[7956]_ ;
  assign \new_[12877]_  = \new_[7974]_  & \new_[7975]_ ;
  assign \new_[12878]_  = \new_[7974]_  ^ \new_[7975]_ ;
  assign \new_[12879]_  = \new_[4755]_  & \new_[4756]_ ;
  assign \new_[12880]_  = \new_[4755]_  ^ \new_[4756]_ ;
  assign \new_[12881]_  = ~\new_[13162]_ ;
  assign \new_[12882]_  = (~\new_[5109]_  | ~\new_[3607]_ ) & (~\new_[5696]_  | ~\new_[7892]_ );
  assign \new_[12883]_  = ~\new_[13998]_ ;
  assign \new_[12884]_  = ~\new_[13136]_ ;
  assign \new_[12885]_  = \new_[7494]_  ^ \new_[3307]_ ;
  assign \new_[12886]_  = ~\new_[13518]_ ;
  assign \new_[12887]_  = ~\new_[13425]_  & ~\new_[2793]_ ;
  assign \new_[12888]_  = ~\new_[13102]_ ;
  assign \new_[12889]_  = ~\new_[13718]_  & ~\new_[3540]_ ;
  assign \new_[12890]_  = ~\new_[2754]_  | ~\new_[13872]_ ;
  assign \new_[12891]_  = ~\new_[14000]_  & ~\new_[13999]_ ;
  assign \new_[12892]_  = ~\new_[13113]_ ;
  assign \new_[12893]_  = ~\new_[13142]_ ;
  assign \new_[12894]_  = ~\new_[13134]_ ;
  assign \new_[12895]_  = ~\new_[13075]_ ;
  assign \new_[12896]_  = ~\new_[13190]_ ;
  assign \new_[12897]_  = ~\new_[13111]_ ;
  assign \new_[12898]_  = \new_[13703]_  & \new_[13695]_ ;
  assign \new_[12899]_  = \new_[13467]_  & \new_[13688]_ ;
  assign \new_[12900]_  = ~\new_[13626]_  & ~\new_[13395]_ ;
  assign \new_[12901]_  = ~\new_[13698]_  & ~\new_[13459]_ ;
  assign \new_[12902]_  = \new_[13396]_  & \new_[13615]_ ;
  assign \new_[12903]_  = ~\new_[7891]_  & ~\new_[13571]_ ;
  assign \new_[12904]_  = ~\new_[13379]_  & ~\new_[13803]_ ;
  assign \new_[12905]_  = ~\new_[13159]_ ;
  assign \new_[12906]_  = ~\new_[13863]_  | ~\new_[7495]_ ;
  assign \new_[12907]_  = \new_[13197]_  & \new_[13796]_ ;
  assign \new_[12908]_  = ~\new_[13803]_  | ~\new_[4767]_ ;
  assign \new_[12909]_  = ~\new_[13467]_  & ~\new_[13688]_ ;
  assign \new_[12910]_  = ~\new_[13128]_ ;
  assign \new_[12911]_  = ~\new_[13228]_  & ~\new_[13606]_ ;
  assign \new_[12912]_  = ~\new_[13624]_  & ~\new_[13563]_ ;
  assign \new_[12913]_  = ~\new_[13183]_ ;
  assign \new_[12914]_  = \new_[13519]_  & \new_[13523]_ ;
  assign \new_[12915]_  = ~\new_[13639]_  & ~\new_[13308]_ ;
  assign \new_[12916]_  = ~\new_[7888]_  & ~\new_[13306]_ ;
  assign \new_[12917]_  = \new_[13200]_  | \new_[13710]_ ;
  assign \new_[12918]_  = ~\new_[13101]_ ;
  assign \new_[12919]_  = \new_[13481]_  & \new_[13707]_ ;
  assign \new_[12920]_  = \new_[13366]_  & \new_[13375]_ ;
  assign \new_[12921]_  = \new_[13809]_  & \new_[13460]_ ;
  assign \new_[12922]_  = ~\new_[7893]_  & ~\new_[13234]_ ;
  assign \new_[12923]_  = ~\new_[13185]_ ;
  assign \new_[12924]_  = ~\new_[13208]_  & ~\new_[3307]_ ;
  assign \new_[12925]_  = ~\new_[13526]_  | ~\new_[4639]_ ;
  assign \new_[12926]_  = ~\new_[13281]_  & ~\wb_addr_i[3] ;
  assign \new_[12927]_  = (~\new_[5104]_  | ~\new_[2816]_ ) & (~\new_[5105]_  | ~\new_[7885]_ );
  assign \new_[12928]_  = (~\new_[5115]_  | ~\new_[7792]_ ) & (~\new_[5116]_  | ~\new_[7891]_ );
  assign \new_[12929]_  = (~\new_[5111]_  | ~\new_[7789]_ ) & (~\new_[5044]_  | ~\new_[7888]_ );
  assign \new_[12930]_  = (~\new_[5112]_  | ~\new_[4068]_ ) & (~\new_[5113]_  | ~\new_[7889]_ );
  assign \new_[12931]_  = (~\new_[5118]_  | ~\new_[2784]_ ) & (~\new_[5119]_  | ~\new_[7925]_ );
  assign \new_[12932]_  = (~\new_[5108]_  | ~\new_[7887]_ ) & (~\new_[5110]_  | ~\new_[4069]_ );
  assign \new_[12933]_  = (~\new_[5101]_  | ~\new_[2783]_ ) & (~\new_[5102]_  | ~\new_[7882]_ );
  assign \new_[12934]_  = ~\new_[13087]_ ;
  assign \new_[12935]_  = ~\new_[13176]_ ;
  assign \new_[12936]_  = ~\new_[13167]_ ;
  assign \new_[12937]_  = ~\new_[13177]_ ;
  assign \new_[12938]_  = ~\new_[13179]_ ;
  assign \new_[12939]_  = ~\new_[13189]_ ;
  assign n11081 = ~\new_[13139]_ ;
  assign \new_[12941]_  = ~\new_[13106]_ ;
  assign \new_[12942]_  = ~\new_[13626]_  | ~\new_[4087]_ ;
  assign \new_[12943]_  = ~\new_[13988]_  | ~\new_[13270]_ ;
  assign \new_[12944]_  = ~\new_[13832]_  | ~\new_[4728]_ ;
  assign \new_[12945]_  = ~\new_[13816]_  | ~\new_[7496]_ ;
  assign \new_[12946]_  = ~\new_[13677]_  & ~\new_[2791]_ ;
  assign \new_[12947]_  = ~\new_[7972]_  & ~\new_[13796]_ ;
  assign \new_[12948]_  = ~\new_[13366]_  | ~\new_[4753]_ ;
  assign \new_[12949]_  = ~\new_[13794]_  & ~\new_[2758]_ ;
  assign \new_[12950]_  = ~\new_[4689]_  | ~\new_[13612]_ ;
  assign \new_[12951]_  = \new_[13208]_  & \new_[3307]_ ;
  assign \new_[12952]_  = ~\new_[13615]_  & ~\new_[13396]_ ;
  assign \new_[12953]_  = \new_[13803]_  & \new_[13379]_ ;
  assign \new_[12954]_  = ~\new_[13563]_  | ~\new_[7774]_ ;
  assign \new_[12955]_  = \new_[13455]_  | \new_[13796]_ ;
  assign \new_[12956]_  = ~\new_[13519]_  & ~\new_[13523]_ ;
  assign \new_[12957]_  = ~\new_[13403]_  | ~\new_[13300]_ ;
  assign \new_[12958]_  = ~\new_[13802]_  & ~\new_[13478]_ ;
  assign \new_[12959]_  = \new_[13526]_  | \new_[13650]_ ;
  assign \new_[12960]_  = ~\new_[7885]_  & ~\new_[13551]_ ;
  assign \new_[12961]_  = ~\new_[13788]_  | ~\new_[13818]_ ;
  assign \new_[12962]_  = ~\new_[13150]_ ;
  assign \new_[12963]_  = ~\new_[7881]_  & ~\new_[13248]_ ;
  assign \new_[12964]_  = \new_[13639]_  & \new_[13308]_ ;
  assign \new_[12965]_  = ~\new_[13270]_  | ~\new_[13991]_ ;
  assign \new_[12966]_  = ~\new_[13827]_  & ~\new_[13604]_ ;
  assign \new_[12967]_  = \new_[13718]_  & \new_[3540]_ ;
  assign \new_[12968]_  = ~\new_[13480]_  & ~\new_[13403]_ ;
  assign \new_[12969]_  = ~\new_[13330]_  & ~\new_[13208]_ ;
  assign \new_[12970]_  = ~\new_[13656]_  & ~\new_[13300]_ ;
  assign \new_[12971]_  = ~\new_[13617]_  & ~\new_[13372]_ ;
  assign \new_[12972]_  = ~\new_[13747]_  & ~\new_[13619]_ ;
  assign \new_[12973]_  = \new_[13823]_  & \new_[13320]_ ;
  assign \new_[12974]_  = ~\new_[7882]_  & ~\new_[13789]_ ;
  assign \new_[12975]_  = \new_[13455]_  & \new_[13726]_ ;
  assign \new_[12976]_  = ~\new_[13811]_  | ~\new_[4763]_ ;
  assign \new_[12977]_  = ~\new_[13125]_ ;
  assign \new_[12978]_  = \new_[13824]_  & \new_[13575]_ ;
  assign \new_[12979]_  = \new_[13724]_  | \new_[14094]_ ;
  assign \new_[12980]_  = ~\new_[13991]_  & ~\new_[13483]_ ;
  assign \new_[12981]_  = ~\new_[13703]_  & ~\new_[13695]_ ;
  assign \new_[12982]_  = ~\new_[13115]_ ;
  assign \new_[12983]_  = \new_[13827]_  & \new_[13604]_ ;
  assign \new_[12984]_  = ~\new_[7793]_  & ~\new_[13597]_ ;
  assign \new_[12985]_  = \new_[13709]_  & \new_[13783]_ ;
  assign \new_[12986]_  = ~\new_[13797]_  | ~\new_[13801]_ ;
  assign \new_[12987]_  = ~\new_[7930]_  & ~\new_[13815]_ ;
  assign \new_[12988]_  = ~\new_[13500]_  & ~\new_[2757]_ ;
  assign \new_[12989]_  = ~\new_[13182]_ ;
  assign \new_[12990]_  = ~\new_[13143]_ ;
  assign \new_[12991]_  = \new_[3306]_ ;
  assign \new_[12992]_  = ~\new_[14127]_  & ~\new_[2759]_ ;
  assign \new_[12993]_  = ~\new_[13223]_ ;
  assign \new_[12994]_  = ~\new_[14037]_ ;
  assign \new_[12995]_  = ~\new_[13622]_ ;
  assign \new_[12996]_  = \new_[3081]_  & \new_[13666]_ ;
  assign \new_[12997]_  = ~\new_[13738]_  & ~\new_[2756]_ ;
  assign \new_[12998]_  = ~\new_[13133]_ ;
  assign \new_[12999]_  = ~\new_[13122]_ ;
  assign \new_[13000]_  = ~\new_[13991]_  | ~\new_[2769]_ ;
  assign \new_[13001]_  = ~\new_[7494]_  & ~\new_[13546]_ ;
  assign \new_[13002]_  = ~\new_[4681]_  & (~\new_[5083]_  | ~\new_[4407]_ );
  assign \new_[13003]_  = ~\new_[13090]_ ;
  assign \new_[13004]_  = ~\new_[13095]_ ;
  assign \new_[13005]_  = \new_[13758]_  | \new_[13867]_ ;
  assign \new_[13006]_  = \new_[13874]_  | \new_[13456]_ ;
  assign \new_[13007]_  = \new_[13877]_  | \new_[13457]_ ;
  assign \new_[13008]_  = ~\new_[13156]_ ;
  assign \new_[13009]_  = \new_[13228]_  & \new_[13606]_ ;
  assign \new_[13010]_  = ~\new_[13701]_  | ~\new_[13700]_ ;
  assign \new_[13011]_  = ~\new_[13131]_ ;
  assign \new_[13012]_  = ~\new_[13605]_ ;
  assign \new_[13013]_  = ~\new_[3081]_  & ~\new_[13666]_ ;
  assign \new_[13014]_  = \new_[13573]_  | \new_[13605]_ ;
  assign \new_[13015]_  = \new_[13281]_  & \wb_addr_i[3] ;
  assign \new_[13016]_  = ~\new_[4682]_  & (~\new_[5098]_  | ~\new_[4583]_ );
  assign \new_[13017]_  = ~\new_[13437]_ ;
  assign \new_[13018]_  = \new_[13734]_  & \new_[13539]_ ;
  assign \new_[13019]_  = ~\new_[7892]_  & ~\new_[13629]_ ;
  assign \new_[13020]_  = ~\new_[13172]_ ;
  assign \new_[13021]_  = ~\new_[13375]_  & ~\new_[13366]_ ;
  assign \new_[13022]_  = ~\new_[7886]_  & ~\new_[13822]_ ;
  assign \new_[13023]_  = ~\new_[13145]_ ;
  assign \new_[13024]_  = ~\new_[7890]_  & ~\new_[13322]_ ;
  assign \new_[13025]_  = \new_[13811]_  & \new_[13612]_ ;
  assign \new_[13026]_  = ~\new_[13184]_ ;
  assign \new_[13027]_  = \new_[13692]_  | \new_[13868]_ ;
  assign \new_[13028]_  = ~\new_[13756]_  & ~\new_[13718]_ ;
  assign \new_[13029]_  = ~\new_[13816]_  | ~\new_[13714]_ ;
  assign \new_[13030]_  = ~\new_[13863]_  | ~\new_[13828]_ ;
  assign \new_[13031]_  = ~\new_[13683]_  | ~\new_[13478]_ ;
  assign \new_[13032]_  = ~\new_[13809]_  & ~\new_[13460]_ ;
  assign \new_[13033]_  = ~\new_[7883]_  & ~\new_[13620]_ ;
  assign \new_[13034]_  = ~\new_[13163]_ ;
  assign \new_[13035]_  = \new_[5082]_  & \new_[13489]_ ;
  assign \new_[13036]_  = ~\wb_addr_i[6]  & ~\new_[13538]_ ;
  assign \new_[13037]_  = \new_[13481]_  | \new_[5767]_ ;
  assign \new_[13038]_  = \new_[13582]_  | \new_[13875]_ ;
  assign \new_[13039]_  = ~\new_[14090]_  | ~\new_[2792]_ ;
  assign \new_[13040]_  = ~\new_[14090]_  & ~\new_[14091]_ ;
  assign \new_[13041]_  = ~\new_[13094]_ ;
  assign \new_[13042]_  = ~\new_[13117]_ ;
  assign \new_[13043]_  = ~\new_[13173]_ ;
  assign \new_[13044]_  = ~\new_[13160]_ ;
  assign \new_[13045]_  = ~\new_[7887]_  & ~\new_[13545]_ ;
  assign \new_[13046]_  = ~\new_[13166]_ ;
  assign \new_[13047]_  = (~\new_[5114]_  | ~\new_[7890]_ ) & (~\new_[5671]_  | ~\new_[3760]_ );
  assign \new_[13048]_  = ~\new_[5091]_  & ~\new_[13372]_ ;
  assign \new_[13049]_  = (~\new_[5106]_  | ~\new_[2817]_ ) & (~\new_[5107]_  | ~\new_[7886]_ );
  assign \new_[13050]_  = ~\new_[4691]_  | ~\new_[13688]_ ;
  assign \new_[13051]_  = (~\new_[5100]_  | ~\new_[7881]_ ) & (~\new_[5120]_  | ~\new_[7930]_ );
  assign \new_[13052]_  = ~\new_[5091]_  | ~\new_[13372]_ ;
  assign \new_[13053]_  = ~\new_[13164]_ ;
  assign \new_[13054]_  = ~\new_[13086]_ ;
  assign \new_[13055]_  = ~\new_[13709]_  & ~\new_[13783]_ ;
  assign \new_[13056]_  = ~\new_[7492]_  | ~\new_[13828]_ ;
  assign \new_[13057]_  = ~\new_[13734]_  & ~\new_[13539]_ ;
  assign \new_[13058]_  = ~\new_[13084]_ ;
  assign \new_[13059]_  = ~\new_[7493]_  | ~\new_[13714]_ ;
  assign \new_[13060]_  = ~\new_[13187]_ ;
  assign \new_[13061]_  = (~\new_[5103]_  | ~\new_[7883]_ ) & (~\new_[5122]_  | ~\new_[7793]_ );
  assign n11086 = u1_sdata_in_r_reg;
  assign \new_[13063]_  = ~\new_[4684]_  & (~\new_[5873]_  | ~\new_[7499]_ );
  assign \new_[13064]_  = ~\new_[13228]_  | ~\new_[4764]_ ;
  assign \new_[13065]_  = ~\new_[4673]_  & (~\new_[5088]_  | ~\new_[5853]_ );
  assign \new_[13066]_  = ~\new_[13467]_  | ~\new_[4765]_ ;
  assign \new_[13067]_  = ~\new_[2750]_  | ~\new_[13844]_ ;
  assign \new_[13068]_  = ~\new_[7894]_  & ~\new_[13337]_ ;
  assign \new_[13069]_  = (~\new_[5117]_  | ~\new_[2818]_ ) & (~\new_[5121]_  | ~\new_[7893]_ );
  assign \new_[13070]_  = \new_[13878]_  | \new_[13592]_ ;
  assign \new_[13071]_  = ~\new_[13820]_  | ~\new_[5716]_ ;
  assign \new_[13072]_  = (~\new_[5043]_  | ~\new_[7894]_ ) & (~\new_[5601]_  | ~\new_[2819]_ );
  assign \new_[13073]_  = ~\new_[7925]_  & ~\new_[13199]_ ;
  assign \new_[13074]_  = ~\new_[4686]_  & (~\new_[5847]_  | ~\new_[6792]_ );
  assign \new_[13075]_  = ~\new_[13425]_ ;
  assign \new_[13076]_  = \new_[7494]_  & \new_[13546]_ ;
  assign \new_[13077]_  = \new_[13799]_  | \new_[13518]_ ;
  assign \new_[13078]_  = ~\new_[14000]_  | ~\new_[13999]_ ;
  assign \new_[13079]_  = \new_[13354]_  & \new_[13315]_ ;
  assign \new_[13080]_  = ~\new_[4683]_  & (~\new_[5081]_  | ~\new_[4815]_ );
  assign \new_[13081]_  = ~\new_[13396]_  | ~\new_[4766]_ ;
  assign \new_[13082]_  = ~\new_[13601]_ ;
  assign \new_[13083]_  = ~\new_[13366]_ ;
  assign \new_[13084]_  = ~\new_[13281]_ ;
  assign \new_[13085]_  = ~\new_[13655]_ ;
  assign \new_[13086]_  = \\u12_dout_reg[7] ;
  assign \new_[13087]_  = \\u12_dout_reg[4] ;
  assign \new_[13088]_  = ~\new_[13582]_ ;
  assign \new_[13089]_  = ~\new_[7439]_  & ~\new_[2952]_ ;
  assign \new_[13090]_  = \\u12_dout_reg[12] ;
  assign \new_[13091]_  = ~\new_[13683]_ ;
  assign \new_[13092]_  = ~\new_[13803]_ ;
  assign \new_[13093]_  = ~\new_[13844]_ ;
  assign \new_[13094]_  = \\u12_dout_reg[24] ;
  assign \new_[13095]_  = \\u12_dout_reg[26] ;
  assign \new_[13096]_  = ~\new_[13666]_ ;
  assign \new_[13097]_  = ~\new_[7438]_  & ~\new_[3150]_ ;
  assign \new_[13098]_  = ~\new_[13801]_ ;
  assign \new_[13099]_  = ~\new_[7792]_  & ~\new_[7506]_ ;
  assign \new_[13100]_  = \new_[3340]_  & \new_[3081]_ ;
  assign \new_[13101]_  = ~\new_[7492]_  | ~\new_[7495]_ ;
  assign \new_[13102]_  = ~\new_[4689]_  | ~\new_[4763]_ ;
  assign \new_[13103]_  = ~\wb_addr_i[2]  & ~\wb_addr_i[3] ;
  assign \new_[13104]_  = ~\new_[13589]_ ;
  assign \new_[13105]_  = ~\new_[13379]_ ;
  assign \new_[13106]_  = \\u12_dout_reg[23] ;
  assign \new_[13107]_  = ~\new_[7889]_  & ~\new_[7491]_ ;
  assign \new_[13108]_  = ~\new_[13700]_ ;
  assign \new_[13109]_  = ~\wb_addr_i[4] ;
  assign \new_[13110]_  = ~\new_[13278]_ ;
  assign \new_[13111]_  = \\u12_dout_reg[11] ;
  assign \new_[13112]_  = ~\new_[13538]_ ;
  assign \new_[13113]_  = ~\new_[14090]_ ;
  assign \new_[13114]_  = ~wb_we_i & ~\new_[9144]_ ;
  assign \new_[13115]_  = \new_[7494]_  | \new_[7498]_ ;
  assign \new_[13116]_  = ~\new_[7494]_  | ~\new_[3307]_ ;
  assign \new_[13117]_  = \\u12_dout_reg[31] ;
  assign \new_[13118]_  = ~\new_[7497]_  & ~\new_[3374]_ ;
  assign \new_[13119]_  = ~\new_[2757]_  & ~\new_[4758]_ ;
  assign \new_[13120]_  = \new_[8477]_  & wb_cyc_i;
  assign \new_[13121]_  = ~\new_[13396]_ ;
  assign \new_[13122]_  = \\u12_dout_reg[13] ;
  assign \new_[13123]_  = \\u12_dout_reg[29] ;
  assign \new_[13124]_  = ~\new_[13467]_ ;
  assign \new_[13125]_  = ~\wb_addr_i[3]  & ~\wb_addr_i[4] ;
  assign \new_[13126]_  = ~\new_[13724]_ ;
  assign \new_[13127]_  = ~\new_[13606]_ ;
  assign \new_[13128]_  = \\u12_dout_reg[22] ;
  assign \new_[13129]_  = ~\new_[13788]_ ;
  assign \new_[13130]_  = ~\new_[13818]_ ;
  assign \new_[13131]_  = ~\new_[7494]_  | ~\new_[7498]_ ;
  assign \new_[13132]_  = \\u12_dout_reg[30] ;
  assign \new_[13133]_  = \\u12_dout_reg[15] ;
  assign \new_[13134]_  = ~\new_[13844]_ ;
  assign \new_[13135]_  = ~\new_[13738]_ ;
  assign \new_[13136]_  = \\u12_dout_reg[19] ;
  assign \new_[13137]_  = ~\new_[13200]_ ;
  assign \new_[13138]_  = ~\new_[7789]_  & ~\new_[7490]_ ;
  assign \new_[13139]_  = ~u2_bit_clk_r_reg;
  assign \new_[13140]_  = ~\new_[13500]_ ;
  assign \new_[13141]_  = ~\new_[13718]_ ;
  assign \new_[13142]_  = ~\new_[13600]_ ;
  assign \new_[13143]_  = ~\new_[13478]_ ;
  assign \new_[13144]_  = ~\new_[13688]_ ;
  assign \new_[13145]_  = ~\new_[7493]_  | ~\new_[7496]_ ;
  assign \new_[13146]_  = ~\new_[5091]_  & ~\new_[5090]_ ;
  assign \new_[13147]_  = ~\new_[5099]_  | ~\new_[7791]_ ;
  assign \new_[13148]_  = wb_we_i & wb_stb_i;
  assign \new_[13149]_  = ~\new_[2791]_  & ~\new_[4768]_ ;
  assign \new_[13150]_  = ~\new_[3081]_  | ~\new_[3082]_ ;
  assign \new_[13151]_  = ~\new_[14000]_ ;
  assign \new_[13152]_  = ~\new_[4591]_  & ~\new_[4648]_ ;
  assign \new_[13153]_  = ~\new_[14000]_ ;
  assign \new_[13154]_  = ~\new_[13794]_ ;
  assign \new_[13155]_  = ~\new_[13797]_ ;
  assign \new_[13156]_  = \\u12_dout_reg[27] ;
  assign \new_[13157]_  = ~\new_[13701]_ ;
  assign \new_[13158]_  = ~\new_[13396]_ ;
  assign \new_[13159]_  = \\u12_dout_reg[28] ;
  assign \new_[13160]_  = ~wb_cyc_i | ~wb_stb_i;
  assign \new_[13161]_  = ~\new_[13228]_ ;
  assign \new_[13162]_  = \\u12_dout_reg[10] ;
  assign \new_[13163]_  = \\u12_dout_reg[6] ;
  assign \new_[13164]_  = \\u12_dout_reg[20] ;
  assign \new_[13165]_  = \wb_addr_i[31]  | \wb_addr_i[29] ;
  assign \new_[13166]_  = \\u12_dout_reg[0] ;
  assign \new_[13167]_  = \\u12_dout_reg[21] ;
  assign \new_[13168]_  = \new_[13710]_ ;
  assign \new_[13169]_  = ~\new_[13615]_ ;
  assign \new_[13170]_  = \new_[7956]_  & \new_[8099]_ ;
  assign \new_[13171]_  = ~\new_[8114]_  & ~\new_[7865]_ ;
  assign \new_[13172]_  = \\u12_dout_reg[5] ;
  assign \new_[13173]_  = \\u12_dout_reg[18] ;
  assign \new_[13174]_  = ~\new_[3788]_  | ~\new_[3119]_ ;
  assign \new_[13175]_  = ~\new_[13375]_ ;
  assign \new_[13176]_  = \\u12_dout_reg[25] ;
  assign \new_[13177]_  = \\u12_dout_reg[2] ;
  assign \new_[13178]_  = ~\new_[2793]_  & ~\new_[4759]_ ;
  assign \new_[13179]_  = \\u12_dout_reg[9] ;
  assign \new_[13180]_  = ~\new_[13803]_ ;
  assign \new_[13181]_  = ~\new_[13692]_ ;
  assign \new_[13182]_  = \\u12_dout_reg[17] ;
  assign \new_[13183]_  = \\u12_dout_reg[3] ;
  assign \new_[13184]_  = \\u12_dout_reg[8] ;
  assign \new_[13185]_  = \\u12_dout_reg[16] ;
  assign \new_[13186]_  = ~\new_[13677]_ ;
  assign \new_[13187]_  = \\u12_dout_reg[14] ;
  assign \new_[13188]_  = ~\new_[13546]_ ;
  assign \new_[13189]_  = \\u12_dout_reg[1] ;
  assign \new_[13190]_  = \new_[13270]_ ;
  assign \new_[13191]_  = ~\new_[3263]_ ;
  assign \new_[13192]_  = ~\new_[3076]_ ;
  assign \new_[13193]_  = ~\new_[3205]_ ;
  assign \new_[13194]_  = ~\new_[3212]_ ;
  assign \new_[13195]_  = ~\new_[3534]_ ;
  assign \new_[13196]_  = ~\new_[3038]_ ;
  assign \new_[13197]_  = ~\new_[7807]_ ;
  assign \new_[13198]_  = ~\new_[2832]_ ;
  assign \new_[13199]_  = ~\new_[3603]_ ;
  assign \new_[13200]_  = ~\new_[5851]_ ;
  assign \new_[13201]_  = ~\new_[2929]_ ;
  assign \new_[13202]_  = ~\new_[3571]_ ;
  assign \new_[13203]_  = ~\new_[3559]_ ;
  assign \new_[13204]_  = ~\new_[3066]_ ;
  assign \new_[13205]_  = ~\new_[3544]_ ;
  assign \new_[13206]_  = ~\new_[2838]_ ;
  assign \new_[13207]_  = ~\new_[2865]_ ;
  assign \new_[13208]_  = ~\new_[3306]_ ;
  assign \new_[13209]_  = ~\new_[3022]_ ;
  assign \new_[13210]_  = ~\new_[3092]_ ;
  assign \new_[13211]_  = ~\new_[3037]_ ;
  assign \new_[13212]_  = ~\new_[3114]_ ;
  assign \new_[13213]_  = ~\new_[3310]_ ;
  assign \new_[13214]_  = ~\new_[3097]_ ;
  assign \new_[13215]_  = ~\new_[3517]_ ;
  assign \new_[13216]_  = ~\new_[3453]_ ;
  assign \new_[13217]_  = ~\new_[3340]_ ;
  assign \new_[13218]_  = ~\new_[5123]_ ;
  assign \new_[13219]_  = ~\new_[3096]_ ;
  assign \new_[13220]_  = ~\new_[2864]_ ;
  assign \new_[13221]_  = ~\new_[3585]_ ;
  assign \new_[13222]_  = ~\new_[3409]_ ;
  assign \new_[13223]_  = ~\new_[5087]_ ;
  assign \new_[13224]_  = ~\new_[3527]_ ;
  assign \new_[13225]_  = ~\new_[2836]_ ;
  assign \new_[13226]_  = ~\new_[3516]_ ;
  assign \new_[13227]_  = ~\new_[3222]_ ;
  assign \new_[13228]_  = ~\new_[4690]_ ;
  assign \new_[13229]_  = ~\new_[3221]_ ;
  assign \new_[13230]_  = ~\new_[2863]_ ;
  assign \new_[13231]_  = ~\new_[2888]_ ;
  assign \new_[13232]_  = ~\new_[3464]_ ;
  assign \new_[13233]_  = ~\new_[3452]_ ;
  assign \new_[13234]_  = ~\new_[4644]_ ;
  assign \new_[13235]_  = ~\new_[3093]_ ;
  assign \new_[13236]_  = ~\new_[3077]_ ;
  assign \new_[13237]_  = ~\new_[3196]_ ;
  assign \new_[13238]_  = ~\new_[3067]_ ;
  assign \new_[13239]_  = ~\new_[3035]_ ;
  assign \new_[13240]_  = ~\new_[3266]_ ;
  assign \new_[13241]_  = ~\new_[3268]_ ;
  assign \new_[13242]_  = ~\new_[3039]_ ;
  assign \new_[13243]_  = ~\new_[2862]_ ;
  assign \new_[13244]_  = ~\new_[2847]_ ;
  assign \new_[13245]_  = ~\new_[3034]_ ;
  assign \new_[13246]_  = ~\new_[3480]_ ;
  assign \new_[13247]_  = ~\new_[2949]_ ;
  assign \new_[13248]_  = ~\new_[4664]_ ;
  assign \new_[13249]_  = ~\new_[2892]_ ;
  assign \new_[13250]_  = ~\new_[3535]_ ;
  assign \new_[13251]_  = ~\new_[3094]_ ;
  assign \new_[13252]_  = ~\new_[3062]_ ;
  assign \new_[13253]_  = ~\new_[3194]_ ;
  assign \new_[13254]_  = ~\new_[3219]_ ;
  assign \new_[13255]_  = ~\new_[2845]_ ;
  assign \new_[13256]_  = ~\new_[3553]_ ;
  assign \new_[13257]_  = ~\new_[3486]_ ;
  assign \new_[13258]_  = ~\new_[3061]_ ;
  assign \new_[13259]_  = ~\new_[2861]_ ;
  assign \new_[13260]_  = ~\new_[3091]_ ;
  assign \new_[13261]_  = ~\new_[3033]_ ;
  assign \new_[13262]_  = ~\new_[3318]_ ;
  assign \new_[13263]_  = ~\new_[3512]_ ;
  assign \new_[13264]_  = ~\new_[2891]_ ;
  assign \new_[13265]_  = ~\new_[3302]_ ;
  assign \new_[13266]_  = ~\new_[3333]_ ;
  assign \new_[13267]_  = ~\new_[3515]_ ;
  assign \new_[13268]_  = ~\new_[3509]_ ;
  assign \new_[13269]_  = ~\new_[5667]_ ;
  assign \new_[13270]_  = ~\new_[2769]_ ;
  assign \new_[13271]_  = ~\new_[3200]_ ;
  assign \new_[13272]_  = ~\new_[2860]_ ;
  assign \new_[13273]_  = ~\new_[3460]_ ;
  assign \new_[13274]_  = ~\new_[3079]_ ;
  assign \new_[13275]_  = ~\new_[3095]_ ;
  assign \new_[13276]_  = ~\new_[3404]_ ;
  assign \new_[13277]_  = ~\new_[3187]_ ;
  assign \new_[13278]_  = ~\new_[5848]_ ;
  assign \new_[13279]_  = ~\new_[3192]_ ;
  assign \new_[13280]_  = ~\new_[2879]_ ;
  assign \new_[13281]_  = ~\wb_addr_i[2] ;
  assign \new_[13282]_  = ~\new_[3032]_ ;
  assign \new_[13283]_  = ~\new_[3153]_ ;
  assign \new_[13284]_  = ~\new_[3484]_ ;
  assign \new_[13285]_  = ~\new_[3218]_ ;
  assign \new_[13286]_  = ~\new_[3220]_ ;
  assign \new_[13287]_  = ~\new_[3031]_ ;
  assign \new_[13288]_  = ~\new_[3337]_ ;
  assign \new_[13289]_  = ~\new_[3152]_ ;
  assign \new_[13290]_  = ~\new_[3508]_ ;
  assign \new_[13291]_  = ~\new_[3323]_ ;
  assign \new_[13292]_  = ~\new_[3223]_ ;
  assign \new_[13293]_  = ~\new_[3202]_ ;
  assign \new_[13294]_  = ~\new_[3541]_ ;
  assign \new_[13295]_  = ~\new_[3036]_ ;
  assign \new_[13296]_  = ~\new_[3363]_ ;
  assign \new_[13297]_  = ~\new_[3227]_ ;
  assign \new_[13298]_  = ~\new_[3151]_ ;
  assign \new_[13299]_  = ~\new_[2889]_ ;
  assign \new_[13300]_  = ~\new_[7973]_ ;
  assign \new_[13301]_  = ~\new_[3229]_ ;
  assign \new_[13302]_  = ~\new_[3203]_ ;
  assign \new_[13303]_  = ~\new_[3030]_ ;
  assign \new_[13304]_  = ~\new_[3080]_ ;
  assign \new_[13305]_  = ~\new_[3231]_ ;
  assign \new_[13306]_  = ~\new_[4411]_ ;
  assign \new_[13307]_  = ~\new_[3233]_ ;
  assign \new_[13308]_  = ~\new_[5077]_ ;
  assign \new_[13309]_  = ~\new_[3234]_ ;
  assign \new_[13310]_  = ~\new_[3494]_ ;
  assign \new_[13311]_  = ~\new_[3236]_ ;
  assign \new_[13312]_  = ~\new_[3550]_ ;
  assign \new_[13313]_  = ~\new_[3237]_ ;
  assign \new_[13314]_  = ~\new_[4762]_ ;
  assign \new_[13315]_  = ~\new_[5089]_ ;
  assign \new_[13316]_  = ~\new_[4761]_ ;
  assign \new_[13317]_  = ~\new_[2796]_ ;
  assign \new_[13318]_  = ~\new_[3469]_ ;
  assign \new_[13319]_  = ~\new_[3239]_ ;
  assign \new_[13320]_  = ~\new_[4587]_ ;
  assign \new_[13321]_  = ~\new_[3145]_ ;
  assign \new_[13322]_  = ~\new_[3605]_ ;
  assign \new_[13323]_  = ~\new_[3320]_ ;
  assign \new_[13324]_  = ~\new_[5126]_ ;
  assign \new_[13325]_  = ~\new_[3243]_ ;
  assign \new_[13326]_  = ~\new_[3247]_ ;
  assign \new_[13327]_  = ~\new_[3501]_ ;
  assign \new_[13328]_  = ~\new_[3500]_ ;
  assign \new_[13329]_  = ~\new_[3502]_ ;
  assign \new_[13330]_  = ~\new_[3587]_ ;
  assign \new_[13331]_  = ~\new_[2842]_ ;
  assign \new_[13332]_  = ~\new_[3025]_ ;
  assign \new_[13333]_  = ~\new_[3487]_ ;
  assign \new_[13334]_  = ~\new_[3021]_ ;
  assign \new_[13335]_  = ~\new_[3090]_ ;
  assign \new_[13336]_  = ~\new_[3581]_ ;
  assign \new_[13337]_  = ~\new_[4645]_ ;
  assign \new_[13338]_  = ~\new_[3084]_ ;
  assign \new_[13339]_  = ~\new_[2873]_ ;
  assign \new_[13340]_  = ~\new_[3506]_ ;
  assign \new_[13341]_  = ~\new_[3028]_ ;
  assign \new_[13342]_  = ~\new_[3069]_ ;
  assign \new_[13343]_  = ~\new_[2855]_ ;
  assign \new_[13344]_  = ~\new_[3606]_ ;
  assign \new_[13345]_  = ~\new_[3279]_ ;
  assign \new_[13346]_  = ~\new_[3505]_ ;
  assign \new_[13347]_  = ~\new_[3543]_ ;
  assign \new_[13348]_  = ~\new_[3262]_ ;
  assign \new_[13349]_  = ~\new_[3563]_ ;
  assign \new_[13350]_  = ~\new_[2890]_ ;
  assign \new_[13351]_  = ~\new_[3304]_ ;
  assign \new_[13352]_  = ~\new_[3088]_ ;
  assign \new_[13353]_  = ~\new_[3083]_ ;
  assign \new_[13354]_  = ~\new_[5694]_ ;
  assign \new_[13355]_  = ~\new_[3574]_ ;
  assign \new_[13356]_  = ~\new_[3554]_ ;
  assign \new_[13357]_  = ~\new_[3138]_ ;
  assign \new_[13358]_  = ~\new_[3248]_ ;
  assign \new_[13359]_  = ~\new_[3026]_ ;
  assign \new_[13360]_  = ~\new_[3245]_ ;
  assign \new_[13361]_  = ~\new_[2801]_ ;
  assign \new_[13362]_  = ~\new_[3498]_ ;
  assign \new_[13363]_  = ~\new_[3241]_ ;
  assign \new_[13364]_  = ~\new_[3209]_ ;
  assign \new_[13365]_  = ~\new_[2759]_ ;
  assign \new_[13366]_  = ~\new_[4692]_ ;
  assign \new_[13367]_  = ~\new_[3278]_ ;
  assign \new_[13368]_  = ~\new_[3214]_ ;
  assign \new_[13369]_  = ~\new_[2800]_ ;
  assign \new_[13370]_  = ~\new_[5132]_ ;
  assign \new_[13371]_  = ~\new_[3235]_ ;
  assign \new_[13372]_  = ~\new_[5090]_ ;
  assign \new_[13373]_  = ~\new_[3583]_ ;
  assign \new_[13374]_  = ~\new_[3149]_ ;
  assign \new_[13375]_  = ~\new_[4753]_ ;
  assign \new_[13376]_  = ~\new_[3513]_ ;
  assign \new_[13377]_  = ~\new_[2872]_ ;
  assign \new_[13378]_  = ~\new_[3157]_ ;
  assign \new_[13379]_  = ~\new_[4767]_ ;
  assign \new_[13380]_  = ~\new_[3520]_ ;
  assign \new_[13381]_  = ~\new_[3514]_ ;
  assign \new_[13382]_  = ~\new_[5130]_ ;
  assign \new_[13383]_  = ~\new_[3106]_ ;
  assign \new_[13384]_  = ~wb_ack_o;
  assign \new_[13385]_  = ~\new_[2874]_ ;
  assign \new_[13386]_  = ~\new_[3510]_ ;
  assign \new_[13387]_  = ~\new_[3134]_ ;
  assign \new_[13388]_  = ~\new_[2839]_ ;
  assign \new_[13389]_  = ~\new_[3049]_ ;
  assign \new_[13390]_  = ~\new_[3179]_ ;
  assign \new_[13391]_  = ~\new_[2886]_ ;
  assign \new_[13392]_  = ~\new_[3089]_ ;
  assign \new_[13393]_  = ~\new_[3334]_ ;
  assign \new_[13394]_  = ~\new_[3521]_ ;
  assign \new_[13395]_  = ~\new_[4087]_ ;
  assign \new_[13396]_  = ~\new_[4693]_ ;
  assign \new_[13397]_  = ~\new_[3536]_ ;
  assign \new_[13398]_  = ~\new_[3159]_ ;
  assign \new_[13399]_  = ~\new_[3098]_ ;
  assign \new_[13400]_  = ~\new_[3569]_ ;
  assign \new_[13401]_  = ~\new_[3217]_ ;
  assign \new_[13402]_  = ~\new_[3042]_ ;
  assign \new_[13403]_  = ~\new_[7935]_ ;
  assign \new_[13404]_  = ~\new_[3099]_ ;
  assign \new_[13405]_  = ~\new_[2927]_ ;
  assign \new_[13406]_  = ~\new_[3457]_ ;
  assign \new_[13407]_  = ~\dma_req_o[5] ;
  assign \new_[13408]_  = ~\new_[4902]_ ;
  assign \new_[13409]_  = ~\new_[3473]_ ;
  assign \new_[13410]_  = ~\new_[3551]_ ;
  assign \new_[13411]_  = ~\new_[3415]_ ;
  assign \new_[13412]_  = ~\new_[3328]_ ;
  assign \new_[13413]_  = ~\new_[2868]_ ;
  assign \new_[13414]_  = ~\new_[3462]_ ;
  assign \new_[13415]_  = ~\new_[2869]_ ;
  assign \new_[13416]_  = ~\new_[2859]_ ;
  assign \new_[13417]_  = ~\new_[3201]_ ;
  assign \new_[13418]_  = ~\new_[3406]_ ;
  assign \new_[13419]_  = ~\new_[3045]_ ;
  assign \new_[13420]_  = ~\new_[3479]_ ;
  assign \new_[13421]_  = ~\dma_req_o[1] ;
  assign \new_[13422]_  = ~\new_[3046]_ ;
  assign \new_[13423]_  = ~\new_[3274]_ ;
  assign \new_[13424]_  = ~\new_[3047]_ ;
  assign \new_[13425]_  = ~\new_[3024]_ ;
  assign \new_[13426]_  = ~\new_[3275]_ ;
  assign \new_[13427]_  = ~\new_[3063]_ ;
  assign \new_[13428]_  = ~\new_[2822]_ ;
  assign \new_[13429]_  = ~\new_[3195]_ ;
  assign \new_[13430]_  = ~\new_[3276]_ ;
  assign \new_[13431]_  = ~\new_[3277]_ ;
  assign \new_[13432]_  = ~\new_[3556]_ ;
  assign \new_[13433]_  = ~\new_[2928]_ ;
  assign \new_[13434]_  = ~\dma_req_o[0] ;
  assign \new_[13435]_  = ~\new_[3048]_ ;
  assign \new_[13436]_  = ~\new_[3475]_ ;
  assign \new_[13437]_  = ~\new_[5080]_ ;
  assign \new_[13438]_  = ~\new_[3258]_ ;
  assign \new_[13439]_  = ~\new_[3477]_ ;
  assign \new_[13440]_  = ~\new_[3281]_ ;
  assign \new_[13441]_  = ~\dma_req_o[4] ;
  assign \new_[13442]_  = ~\new_[2867]_ ;
  assign \new_[13443]_  = ~\new_[3451]_ ;
  assign \new_[13444]_  = ~\new_[3109]_ ;
  assign \new_[13445]_  = ~\new_[2846]_ ;
  assign \new_[13446]_  = ~\new_[3414]_ ;
  assign \new_[13447]_  = ~\new_[3110]_ ;
  assign \new_[13448]_  = ~\new_[3285]_ ;
  assign \new_[13449]_  = ~\new_[2878]_ ;
  assign \new_[13450]_  = ~\new_[3211]_ ;
  assign \new_[13451]_  = ~\new_[3107]_ ;
  assign \new_[13452]_  = ~\new_[3210]_ ;
  assign \new_[13453]_  = ~\new_[3532]_ ;
  assign \new_[13454]_  = ~\new_[3101]_ ;
  assign \new_[13455]_  = ~\new_[7976]_ ;
  assign \new_[13456]_  = ~\new_[8995]_ ;
  assign \new_[13457]_  = ~\new_[8503]_ ;
  assign \new_[13458]_  = ~\new_[3584]_ ;
  assign \new_[13459]_  = ~\new_[5084]_ ;
  assign \new_[13460]_  = ~\new_[5844]_ ;
  assign \new_[13461]_  = ~\new_[4757]_ ;
  assign \new_[13462]_  = ~\new_[2833]_ ;
  assign \new_[13463]_  = ~\new_[5041]_ ;
  assign \new_[13464]_  = ~\new_[3312]_ ;
  assign \new_[13465]_  = ~\new_[3188]_ ;
  assign \new_[13466]_  = ~\new_[3308]_ ;
  assign \new_[13467]_  = ~\new_[4691]_ ;
  assign \new_[13468]_  = ~\new_[3499]_ ;
  assign \new_[13469]_  = ~\new_[2840]_ ;
  assign \new_[13470]_  = ~\new_[3531]_ ;
  assign \new_[13471]_  = ~\new_[2824]_ ;
  assign \new_[13472]_  = ~\new_[3322]_ ;
  assign \new_[13473]_  = ~\new_[3411]_ ;
  assign \new_[13474]_  = ~\new_[3250]_ ;
  assign \new_[13475]_  = ~\new_[3327]_ ;
  assign \new_[13476]_  = ~\new_[3293]_ ;
  assign \new_[13477]_  = ~\new_[3087]_ ;
  assign \new_[13478]_  = ~\new_[2770]_ ;
  assign \new_[13479]_  = ~\new_[3549]_ ;
  assign \new_[13480]_  = ~\new_[7978]_ ;
  assign \new_[13481]_  = ~\new_[5843]_ ;
  assign \new_[13482]_  = ~\new_[4754]_ ;
  assign \new_[13483]_  = ~\new_[2769]_ ;
  assign \new_[13484]_  = ~\new_[3567]_ ;
  assign \new_[13485]_  = ~\new_[3364]_ ;
  assign \new_[13486]_  = ~\new_[3086]_ ;
  assign \new_[13487]_  = ~\new_[3524]_ ;
  assign \new_[13488]_  = ~\new_[3329]_ ;
  assign \new_[13489]_  = ~\new_[5716]_ ;
  assign \new_[13490]_  = ~\new_[3309]_ ;
  assign \new_[13491]_  = ~\new_[3562]_ ;
  assign \new_[13492]_  = ~\new_[2853]_ ;
  assign \new_[13493]_  = ~\new_[2854]_ ;
  assign \new_[13494]_  = ~\new_[3542]_ ;
  assign \new_[13495]_  = ~\new_[3050]_ ;
  assign \new_[13496]_  = ~\new_[3108]_ ;
  assign \new_[13497]_  = ~\new_[3377]_ ;
  assign \new_[13498]_  = ~\new_[3523]_ ;
  assign \new_[13499]_  = ~\new_[3456]_ ;
  assign \new_[13500]_  = ~\new_[2829]_ ;
  assign \new_[13501]_  = ~\new_[3252]_ ;
  assign \new_[13502]_  = ~\new_[3525]_ ;
  assign \new_[13503]_  = ~\new_[3566]_ ;
  assign \new_[13504]_  = ~\new_[3405]_ ;
  assign \new_[13505]_  = ~\new_[5134]_ ;
  assign \new_[13506]_  = ~\new_[2883]_ ;
  assign \new_[13507]_  = ~\new_[2837]_ ;
  assign \new_[13508]_  = ~\new_[2852]_ ;
  assign \new_[13509]_  = ~\new_[5129]_ ;
  assign \new_[13510]_  = ~\new_[3180]_ ;
  assign \new_[13511]_  = ~\new_[3141]_ ;
  assign \new_[13512]_  = ~\new_[3454]_ ;
  assign \new_[13513]_  = ~\new_[3407]_ ;
  assign \new_[13514]_  = ~\new_[3468]_ ;
  assign \new_[13515]_  = ~\new_[3019]_ ;
  assign \new_[13516]_  = ~\new_[3199]_ ;
  assign \new_[13517]_  = ~\new_[3555]_ ;
  assign \new_[13518]_  = ~\new_[4917]_ ;
  assign \new_[13519]_  = ~\new_[5071]_ ;
  assign \new_[13520]_  = ~\new_[3761]_ ;
  assign \new_[13521]_  = ~\new_[3489]_ ;
  assign \new_[13522]_  = ~\new_[3027]_ ;
  assign \new_[13523]_  = ~\new_[5070]_ ;
  assign \new_[13524]_  = ~\new_[3576]_ ;
  assign \new_[13525]_  = ~\new_[2826]_ ;
  assign \new_[13526]_  = ~\new_[4640]_ ;
  assign \new_[13527]_  = ~\new_[3552]_ ;
  assign \new_[13528]_  = ~\new_[3455]_ ;
  assign \new_[13529]_  = ~\new_[2798]_ ;
  assign \new_[13530]_  = ~\new_[3577]_ ;
  assign \new_[13531]_  = ~\new_[2844]_ ;
  assign \new_[13532]_  = ~\new_[2758]_ ;
  assign \new_[13533]_  = ~\new_[3311]_ ;
  assign \new_[13534]_  = ~\new_[3116]_ ;
  assign \new_[13535]_  = ~\new_[3257]_ ;
  assign \new_[13536]_  = ~\new_[3522]_ ;
  assign \new_[13537]_  = ~\new_[4758]_ ;
  assign \new_[13538]_  = ~\wb_addr_i[5] ;
  assign \new_[13539]_  = ~\new_[5065]_ ;
  assign \new_[13540]_  = ~\new_[3117]_ ;
  assign \new_[13541]_  = ~\new_[2794]_ ;
  assign \new_[13542]_  = ~\new_[3491]_ ;
  assign \new_[13543]_  = ~\new_[3264]_ ;
  assign \new_[13544]_  = ~\new_[3493]_ ;
  assign \new_[13545]_  = ~\new_[4652]_ ;
  assign \new_[13546]_  = ~\new_[7498]_ ;
  assign \new_[13547]_  = ~\new_[2850]_ ;
  assign \new_[13548]_  = ~\new_[2881]_ ;
  assign \new_[13549]_  = ~\new_[3246]_ ;
  assign \new_[13550]_  = ~\new_[4685]_ ;
  assign \new_[13551]_  = ~\new_[4646]_ ;
  assign \new_[13552]_  = ~\new_[2880]_ ;
  assign \new_[13553]_  = ~\new_[3492]_ ;
  assign \new_[13554]_  = ~\new_[7874]_ ;
  assign \new_[13555]_  = ~\new_[3208]_ ;
  assign \new_[13556]_  = ~\new_[3292]_ ;
  assign \new_[13557]_  = ~\new_[3267]_ ;
  assign \new_[13558]_  = ~\new_[3198]_ ;
  assign \new_[13559]_  = ~\new_[2877]_ ;
  assign \new_[13560]_  = ~\new_[3244]_ ;
  assign \new_[13561]_  = ~\new_[2843]_ ;
  assign \new_[13562]_  = ~\new_[2887]_ ;
  assign \new_[13563]_  = ~\new_[7857]_ ;
  assign \new_[13564]_  = ~\new_[3242]_ ;
  assign \new_[13565]_  = ~\new_[3579]_ ;
  assign \new_[13566]_  = ~\new_[3216]_ ;
  assign \new_[13567]_  = ~\new_[3349]_ ;
  assign \new_[13568]_  = ~\new_[3207]_ ;
  assign \new_[13569]_  = ~\new_[5092]_ ;
  assign \new_[13570]_  = ~\new_[4406]_ ;
  assign \new_[13571]_  = ~\new_[3341]_ ;
  assign \new_[13572]_  = ~\new_[3240]_ ;
  assign \new_[13573]_  = ~\new_[5096]_ ;
  assign \new_[13574]_  = ~\new_[4590]_ ;
  assign \new_[13575]_  = ~\new_[4581]_ ;
  assign \new_[13576]_  = ~\new_[3260]_ ;
  assign \new_[13577]_  = ~\new_[3471]_ ;
  assign \new_[13578]_  = ~\new_[3238]_ ;
  assign \new_[13579]_  = ~\new_[2866]_ ;
  assign \new_[13580]_  = ~\new_[3288]_ ;
  assign \new_[13581]_  = ~\new_[3564]_ ;
  assign \new_[13582]_  = ~\new_[5060]_ ;
  assign \new_[13583]_  = ~\new_[3467]_ ;
  assign \new_[13584]_  = ~\new_[2754]_ ;
  assign \new_[13585]_  = ~\new_[2893]_ ;
  assign \new_[13586]_  = ~\new_[3483]_ ;
  assign \new_[13587]_  = ~\new_[3053]_ ;
  assign \new_[13588]_  = ~\new_[3051]_ ;
  assign \new_[13589]_  = ~\new_[2754]_ ;
  assign \new_[13590]_  = ~\new_[3272]_ ;
  assign \new_[13591]_  = ~\new_[3495]_ ;
  assign \new_[13592]_  = ~\new_[5039]_ ;
  assign \new_[13593]_  = ~\new_[3055]_ ;
  assign \new_[13594]_  = ~\new_[3314]_ ;
  assign \new_[13595]_  = ~\new_[2834]_ ;
  assign \new_[13596]_  = ~\new_[3316]_ ;
  assign \new_[13597]_  = ~\new_[3122]_ ;
  assign \new_[13598]_  = ~\new_[2820]_ ;
  assign \new_[13599]_  = ~\new_[2895]_ ;
  assign \new_[13600]_  = ~\new_[2750]_ ;
  assign \new_[13601]_  = ~\new_[5849]_ ;
  assign \new_[13602]_  = ~\new_[2858]_ ;
  assign \new_[13603]_  = ~\new_[3459]_ ;
  assign \new_[13604]_  = ~\new_[5876]_ ;
  assign \new_[13605]_  = ~\new_[5075]_ ;
  assign \new_[13606]_  = ~\new_[4764]_ ;
  assign \new_[13607]_  = ~\new_[3339]_ ;
  assign \new_[13608]_  = ~\new_[2849]_ ;
  assign \new_[13609]_  = ~\new_[3232]_ ;
  assign \new_[13610]_  = ~\new_[3331]_ ;
  assign \new_[13611]_  = ~\new_[5127]_ ;
  assign \new_[13612]_  = ~\new_[4763]_ ;
  assign \new_[13613]_  = ~\new_[3074]_ ;
  assign \new_[13614]_  = ~\new_[5040]_ ;
  assign \new_[13615]_  = ~\new_[4766]_ ;
  assign \new_[13616]_  = ~\new_[3057]_ ;
  assign \new_[13617]_  = ~\new_[5091]_ ;
  assign \new_[13618]_  = ~\new_[3193]_ ;
  assign \new_[13619]_  = ~\new_[4641]_ ;
  assign \new_[13620]_  = ~\new_[4647]_ ;
  assign \new_[13621]_  = ~\new_[3503]_ ;
  assign \new_[13622]_  = ~\new_[3023]_ ;
  assign \new_[13623]_  = ~\new_[3295]_ ;
  assign \new_[13624]_  = ~\new_[7936]_ ;
  assign \new_[13625]_  = ~\new_[3548]_ ;
  assign \new_[13626]_  = ~\new_[4412]_ ;
  assign \new_[13627]_  = ~\new_[3289]_ ;
  assign \new_[13628]_  = ~\new_[3472]_ ;
  assign \new_[13629]_  = ~\new_[3120]_ ;
  assign \new_[13630]_  = ~\new_[3163]_ ;
  assign \new_[13631]_  = ~\new_[3174]_ ;
  assign \new_[13632]_  = ~\new_[5128]_ ;
  assign \new_[13633]_  = ~\new_[3226]_ ;
  assign \new_[13634]_  = ~\new_[3197]_ ;
  assign \new_[13635]_  = ~\new_[3305]_ ;
  assign \new_[13636]_  = ~\new_[3561]_ ;
  assign \new_[13637]_  = ~\new_[3511]_ ;
  assign \new_[13638]_  = ~\new_[3476]_ ;
  assign \new_[13639]_  = ~\new_[5078]_ ;
  assign \new_[13640]_  = ~\new_[3518]_ ;
  assign \new_[13641]_  = ~\new_[3324]_ ;
  assign \new_[13642]_  = ~\new_[2848]_ ;
  assign \new_[13643]_  = ~\new_[3128]_ ;
  assign \new_[13644]_  = ~\new_[3519]_ ;
  assign \new_[13645]_  = ~\new_[3282]_ ;
  assign \new_[13646]_  = ~\new_[3284]_ ;
  assign \new_[13647]_  = ~\new_[2799]_ ;
  assign \new_[13648]_  = ~\new_[2841]_ ;
  assign \new_[13649]_  = ~\new_[3261]_ ;
  assign \new_[13650]_  = ~\new_[4639]_ ;
  assign \new_[13651]_  = ~\new_[2894]_ ;
  assign \new_[13652]_  = ~\new_[3078]_ ;
  assign \new_[13653]_  = ~\new_[3538]_ ;
  assign \new_[13654]_  = ~\new_[3176]_ ;
  assign \new_[13655]_  = ~\new_[5673]_ ;
  assign \new_[13656]_  = ~\new_[7979]_ ;
  assign \new_[13657]_  = ~\new_[2876]_ ;
  assign \new_[13658]_  = ~\new_[3111]_ ;
  assign \new_[13659]_  = ~\new_[3565]_ ;
  assign \new_[13660]_  = ~\new_[3297]_ ;
  assign \new_[13661]_  = ~\new_[2926]_ ;
  assign \new_[13662]_  = ~\new_[3300]_ ;
  assign \new_[13663]_  = ~\new_[3482]_ ;
  assign \new_[13664]_  = ~\new_[3287]_ ;
  assign \new_[13665]_  = ~\new_[2875]_ ;
  assign \new_[13666]_  = ~\new_[3082]_ ;
  assign \new_[13667]_  = ~\new_[3528]_ ;
  assign \new_[13668]_  = ~\new_[3255]_ ;
  assign \new_[13669]_  = ~\new_[2882]_ ;
  assign \new_[13670]_  = ~\new_[3224]_ ;
  assign \new_[13671]_  = ~\new_[5133]_ ;
  assign \new_[13672]_  = ~\new_[3225]_ ;
  assign \new_[13673]_  = ~\new_[3582]_ ;
  assign \new_[13674]_  = ~\new_[3112]_ ;
  assign \new_[13675]_  = ~\new_[3470]_ ;
  assign \new_[13676]_  = ~\new_[3254]_ ;
  assign \new_[13677]_  = ~\new_[3023]_ ;
  assign \new_[13678]_  = ~\new_[3256]_ ;
  assign \new_[13679]_  = ~\new_[3485]_ ;
  assign \new_[13680]_  = ~\new_[3073]_ ;
  assign \new_[13681]_  = ~\new_[3213]_ ;
  assign \new_[13682]_  = ~\new_[3118]_ ;
  assign \new_[13683]_  = ~\new_[2753]_ ;
  assign \new_[13684]_  = ~\new_[3301]_ ;
  assign \new_[13685]_  = ~\new_[3228]_ ;
  assign \new_[13686]_  = ~\new_[3113]_ ;
  assign \new_[13687]_  = ~\new_[3530]_ ;
  assign \new_[13688]_  = ~\new_[4765]_ ;
  assign \new_[13689]_  = ~\new_[5125]_ ;
  assign \new_[13690]_  = ~\new_[3504]_ ;
  assign \new_[13691]_  = ~\new_[3357]_ ;
  assign \new_[13692]_  = ~\new_[5072]_ ;
  assign \new_[13693]_  = ~\new_[3148]_ ;
  assign \new_[13694]_  = ~\new_[3056]_ ;
  assign \new_[13695]_  = ~\new_[5042]_ ;
  assign \new_[13696]_  = ~\new_[3269]_ ;
  assign \new_[13697]_  = ~\new_[2835]_ ;
  assign \new_[13698]_  = ~\new_[5085]_ ;
  assign \new_[13699]_  = ~\new_[3602]_ ;
  assign \new_[13700]_  = ~\new_[5045]_ ;
  assign \new_[13701]_  = ~\new_[5057]_ ;
  assign \new_[13702]_  = ~\new_[3326]_ ;
  assign \new_[13703]_  = ~\new_[5095]_ ;
  assign \new_[13704]_  = ~\new_[5131]_ ;
  assign \new_[13705]_  = ~\new_[3041]_ ;
  assign \new_[13706]_  = ~\new_[3321]_ ;
  assign \new_[13707]_  = ~\new_[5767]_ ;
  assign \new_[13708]_  = ~\new_[3052]_ ;
  assign \new_[13709]_  = ~\new_[5059]_ ;
  assign \new_[13710]_  = ~\new_[5842]_ ;
  assign \new_[13711]_  = ~\new_[3461]_ ;
  assign \new_[13712]_  = ~\new_[3054]_ ;
  assign \new_[13713]_  = ~\new_[3496]_ ;
  assign \new_[13714]_  = ~\new_[7496]_ ;
  assign \new_[13715]_  = ~\new_[2827]_ ;
  assign \new_[13716]_  = ~\new_[3313]_ ;
  assign \new_[13717]_  = ~\new_[3481]_ ;
  assign \new_[13718]_  = ~\new_[4070]_ ;
  assign \new_[13719]_  = ~\new_[3335]_ ;
  assign \new_[13720]_  = ~\dma_req_o[3] ;
  assign \new_[13721]_  = ~\new_[3104]_ ;
  assign \new_[13722]_  = ~\new_[3537]_ ;
  assign \new_[13723]_  = ~\new_[4759]_ ;
  assign \new_[13724]_  = ~\new_[5846]_ ;
  assign \new_[13725]_  = ~\new_[3448]_ ;
  assign \new_[13726]_  = ~\new_[7972]_ ;
  assign \new_[13727]_  = ~\new_[3072]_ ;
  assign \new_[13728]_  = ~\new_[3130]_ ;
  assign \new_[13729]_  = ~\new_[3103]_ ;
  assign \new_[13730]_  = ~\new_[5037]_ ;
  assign \new_[13731]_  = ~\new_[3338]_ ;
  assign \new_[13732]_  = ~\new_[3319]_ ;
  assign \new_[13733]_  = ~\new_[2870]_ ;
  assign \new_[13734]_  = ~\new_[5066]_ ;
  assign \new_[13735]_  = ~\new_[3332]_ ;
  assign \new_[13736]_  = ~\new_[3070]_ ;
  assign \new_[13737]_  = ~\new_[3071]_ ;
  assign \new_[13738]_  = ~\new_[2828]_ ;
  assign \new_[13739]_  = ~\new_[2797]_ ;
  assign \new_[13740]_  = ~\dma_req_o[2] ;
  assign \new_[13741]_  = ~\new_[3290]_ ;
  assign \new_[13742]_  = ~\new_[3115]_ ;
  assign \new_[13743]_  = ~\new_[3085]_ ;
  assign \new_[13744]_  = ~\new_[3105]_ ;
  assign \new_[13745]_  = ~\new_[2795]_ ;
  assign \new_[13746]_  = ~\new_[3507]_ ;
  assign \new_[13747]_  = ~\new_[4633]_ ;
  assign \new_[13748]_  = ~\new_[3325]_ ;
  assign \new_[13749]_  = ~\new_[3102]_ ;
  assign \new_[13750]_  = ~\new_[3466]_ ;
  assign \new_[13751]_  = ~\new_[3270]_ ;
  assign \new_[13752]_  = ~\new_[3280]_ ;
  assign \new_[13753]_  = ~\new_[3189]_ ;
  assign \new_[13754]_  = ~\new_[3283]_ ;
  assign \new_[13755]_  = ~\new_[3249]_ ;
  assign \new_[13756]_  = ~\new_[3771]_ ;
  assign \new_[13757]_  = ~\new_[4768]_ ;
  assign \new_[13758]_  = ~\new_[8803]_ ;
  assign \new_[13759]_  = ~\new_[3458]_ ;
  assign \new_[13760]_  = ~\new_[3413]_ ;
  assign \new_[13761]_  = ~\new_[3259]_ ;
  assign \new_[13762]_  = ~\new_[3529]_ ;
  assign \new_[13763]_  = ~\new_[3059]_ ;
  assign \new_[13764]_  = ~\new_[3065]_ ;
  assign \new_[13765]_  = ~\new_[3251]_ ;
  assign \new_[13766]_  = ~\new_[3463]_ ;
  assign \new_[13767]_  = ~\new_[2857]_ ;
  assign \new_[13768]_  = ~\new_[3296]_ ;
  assign \new_[13769]_  = ~\new_[4588]_ ;
  assign \new_[13770]_  = ~\new_[3100]_ ;
  assign \new_[13771]_  = ~\new_[2885]_ ;
  assign \new_[13772]_  = ~\new_[3294]_ ;
  assign \new_[13773]_  = ~\new_[3043]_ ;
  assign \new_[13774]_  = ~\new_[3568]_ ;
  assign \new_[13775]_  = ~\new_[2856]_ ;
  assign \new_[13776]_  = ~\new_[3064]_ ;
  assign \new_[13777]_  = ~\new_[3075]_ ;
  assign \new_[13778]_  = ~\new_[3336]_ ;
  assign \new_[13780]_  = ~\new_[2851]_ ;
  assign \new_[13781]_  = ~\new_[3204]_ ;
  assign \new_[13782]_  = ~\new_[3298]_ ;
  assign \new_[13783]_  = ~\new_[5058]_ ;
  assign \new_[13784]_  = ~\new_[3533]_ ;
  assign \new_[13785]_  = ~\new_[3560]_ ;
  assign \new_[13786]_  = ~\new_[3412]_ ;
  assign \new_[13787]_  = ~\new_[3253]_ ;
  assign \new_[13788]_  = ~\new_[5069]_ ;
  assign \new_[13789]_  = ~\new_[3121]_ ;
  assign \new_[13790]_  = ~\new_[5036]_ ;
  assign \new_[13791]_  = ~\new_[4760]_ ;
  assign \new_[13792]_  = ~\new_[3465]_ ;
  assign \new_[13793]_  = ~\new_[3586]_ ;
  assign \new_[13794]_  = ~\new_[2830]_ ;
  assign \new_[13795]_  = ~\new_[3547]_ ;
  assign \new_[13796]_  = ~\new_[7977]_ ;
  assign \new_[13797]_  = ~\new_[5063]_ ;
  assign \new_[13798]_  = ~\new_[5094]_ ;
  assign \new_[13799]_  = ~\new_[5079]_ ;
  assign \new_[13800]_  = ~\new_[3497]_ ;
  assign \new_[13801]_  = ~\new_[5049]_ ;
  assign \new_[13802]_  = ~\new_[2753]_ ;
  assign \new_[13803]_  = ~\new_[4694]_ ;
  assign \new_[13804]_  = ~\new_[3154]_ ;
  assign \new_[13805]_  = ~\new_[3191]_ ;
  assign \new_[13806]_  = ~\new_[3265]_ ;
  assign \new_[13807]_  = ~\new_[3175]_ ;
  assign \new_[13808]_  = ~\new_[3315]_ ;
  assign \new_[13809]_  = ~\new_[5845]_ ;
  assign \new_[13810]_  = ~\new_[4752]_ ;
  assign \new_[13811]_  = ~\new_[4689]_ ;
  assign \new_[13812]_  = ~\new_[2823]_ ;
  assign \new_[13813]_  = ~\new_[5124]_ ;
  assign \new_[13814]_  = ~\new_[3299]_ ;
  assign \new_[13815]_  = ~\new_[3604]_ ;
  assign \new_[13816]_  = ~\new_[7493]_ ;
  assign \new_[13817]_  = ~\new_[3344]_ ;
  assign \new_[13818]_  = ~\new_[5068]_ ;
  assign \new_[13819]_  = ~\new_[3474]_ ;
  assign \new_[13820]_  = ~\new_[5082]_ ;
  assign \new_[13821]_  = ~\new_[3303]_ ;
  assign \new_[13822]_  = ~\new_[3123]_ ;
  assign \new_[13823]_  = ~\new_[4586]_ ;
  assign \new_[13824]_  = ~\new_[4589]_ ;
  assign \new_[13825]_  = ~\new_[3158]_ ;
  assign \new_[13826]_  = ~\new_[3206]_ ;
  assign \new_[13827]_  = ~\new_[5850]_ ;
  assign \new_[13828]_  = ~\new_[7495]_ ;
  assign \new_[13829]_  = ~\new_[3190]_ ;
  assign \new_[13830]_  = ~\new_[3488]_ ;
  assign \new_[13831]_  = ~\new_[3578]_ ;
  assign \new_[13832]_  = ~\new_[4756]_ ;
  assign \new_[13833]_  = ~\new_[3119]_ ;
  assign \new_[13834]_  = ~\new_[3330]_ ;
  assign \new_[13835]_  = ~\new_[3215]_ ;
  assign \new_[13836]_  = ~\new_[3317]_ ;
  assign \new_[13837]_  = ~\new_[3286]_ ;
  assign \new_[13838]_  = ~\new_[3029]_ ;
  assign \new_[13839]_  = ~\new_[3230]_ ;
  assign \new_[13840]_  = ~\new_[3291]_ ;
  assign \new_[13841]_  = ~\new_[3620]_ ;
  assign \new_[13842]_  = ~\new_[3570]_ ;
  assign \new_[13843]_  = ~\new_[3271]_ ;
  assign \new_[13844]_  = ~\new_[2790]_ ;
  assign \new_[13845]_  = ~\new_[3478]_ ;
  assign \new_[13846]_  = ~\new_[2821]_ ;
  assign \new_[13847]_  = ~\new_[3060]_ ;
  assign \new_[13848]_  = ~\new_[3408]_ ;
  assign \new_[13849]_  = ~\new_[3068]_ ;
  assign \new_[13850]_  = ~\new_[3020]_ ;
  assign \new_[13851]_  = ~\new_[3557]_ ;
  assign \new_[13852]_  = ~\new_[3558]_ ;
  assign \new_[13853]_  = ~\new_[2884]_ ;
  assign \new_[13854]_  = ~\new_[3450]_ ;
  assign \new_[13855]_  = ~\new_[2871]_ ;
  assign \new_[13856]_  = ~\new_[3273]_ ;
  assign \new_[13857]_  = ~\new_[2756]_ ;
  assign \new_[13858]_  = ~\new_[3490]_ ;
  assign \new_[13859]_  = ~\new_[3044]_ ;
  assign \new_[13860]_  = ~\new_[3058]_ ;
  assign \new_[13861]_  = ~\new_[3161]_ ;
  assign \new_[13862]_  = ~\new_[3572]_ ;
  assign \new_[13863]_  = ~\new_[7492]_ ;
  assign \new_[13864]_  = ~\new_[3573]_ ;
  assign \new_[13865]_  = ~\new_[3040]_ ;
  assign \new_[13866]_  = ~\new_[13867]_ ;
  assign \new_[13867]_  = \new_[13868]_ ;
  assign \new_[13868]_  = ~\new_[5056]_ ;
  assign \new_[13869]_  = ~\new_[13870]_ ;
  assign \new_[13870]_  = \new_[13871]_ ;
  assign \new_[13871]_  = ~\new_[13872]_ ;
  assign \new_[13872]_  = ~\new_[2772]_ ;
  assign \new_[13873]_  = ~\new_[13874]_ ;
  assign \new_[13874]_  = \new_[13875]_ ;
  assign \new_[13875]_  = ~\new_[4918]_ ;
  assign \new_[13876]_  = ~\new_[13877]_ ;
  assign \new_[13877]_  = \new_[13878]_ ;
  assign \new_[13878]_  = ~\new_[5061]_ ;
  assign \new_[13879]_  = \new_[13883]_ ;
  assign \new_[13880]_  = ~\new_[13881]_ ;
  assign \new_[13881]_  = ~\new_[13883]_ ;
  assign \new_[13882]_  = \new_[13883]_ ;
  assign \new_[13883]_  = ~\new_[12965]_ ;
  assign n4996 = ~\new_[13885]_ ;
  assign \new_[13885]_  = \new_[14004]_ ;
  assign \new_[13886]_  = \new_[13823]_  | \new_[14005]_ ;
  assign \new_[13887]_  = ~\new_[13888]_  & (~\new_[5582]_  | ~\new_[14192]_ );
  assign \new_[13888]_  = \new_[13931]_  & \new_[5251]_ ;
  assign \new_[13889]_  = (~\new_[5276]_  | ~\new_[14172]_ ) & (~\new_[13987]_  | ~\new_[5226]_ );
  assign \new_[13890]_  = ~\new_[13134]_  | ~\new_[13600]_ ;
  assign \new_[13891]_  = ~\new_[13893]_  | ~\new_[13892]_ ;
  assign \new_[13892]_  = (~\new_[5492]_  | ~\new_[14134]_ ) & (~\new_[12635]_  | ~\new_[4967]_ );
  assign \new_[13893]_  = (~\new_[5517]_  | ~\new_[12821]_ ) & (~\new_[13894]_  | ~\new_[5468]_ );
  assign \new_[13894]_  = ~\new_[13895]_ ;
  assign \new_[13895]_  = ~\new_[13896]_ ;
  assign \new_[13896]_  = ~\new_[13997]_ ;
  assign \new_[13897]_  = ~\new_[13895]_ ;
  assign \new_[13898]_  = \new_[14131]_  | \new_[14063]_ ;
  assign \new_[13899]_  = \new_[14131]_  | \new_[14063]_ ;
  assign \new_[13900]_  = \new_[13079]_  | \new_[4716]_ ;
  assign \new_[13901]_  = \new_[13079]_  | \new_[4716]_ ;
  assign \new_[13902]_  = \new_[12919]_  | \new_[4717]_ ;
  assign \new_[13903]_  = \new_[12919]_  | \new_[4717]_ ;
  assign \new_[13904]_  = ~\new_[13905]_  | ~\new_[13907]_ ;
  assign \new_[13905]_  = ~\new_[13906]_  | ~\new_[13935]_ ;
  assign \new_[13906]_  = ~\new_[12300]_  | ~\new_[10917]_  | ~\new_[11250]_  | ~\new_[10997]_ ;
  assign \new_[13907]_  = ~\new_[13908]_  | ~\new_[14145]_ ;
  assign \new_[13908]_  = ~\new_[12298]_  | ~\new_[10842]_  | ~\new_[10606]_  | ~\new_[11010]_ ;
  assign n1926 = ~\new_[13912]_  | (~\new_[13910]_  & ~\new_[4671]_ );
  assign \new_[13910]_  = ~\new_[4279]_  | ~\new_[13911]_ ;
  assign \new_[13911]_  = ~\dma_ack_i[8] ;
  assign \new_[13912]_  = ~\dma_req_o[8]  | ~\new_[13911]_ ;
  assign n4591 = ~\new_[4671]_  & ~\dma_ack_i[8] ;
  assign \new_[13914]_  = ~\new_[4473]_  | (~\new_[13915]_  & ~\new_[13916]_ );
  assign \new_[13915]_  = ~\new_[8376]_  | (~\new_[8748]_  & ~\new_[12363]_ );
  assign \new_[13916]_  = ~\new_[13917]_  | ~\new_[13918]_ ;
  assign \new_[13917]_  = ~\new_[14087]_  | ~\new_[8855]_  | ~\new_[13500]_ ;
  assign \new_[13918]_  = ~\new_[13919]_  | (~\new_[9825]_  & ~\new_[9826]_ );
  assign \new_[13919]_  = \new_[13140]_  & \new_[14087]_ ;
  assign \new_[13920]_  = ~\new_[13955]_  | (~\new_[13921]_  & ~\new_[13922]_ );
  assign \new_[13921]_  = ~\new_[12792]_  & (~\new_[8319]_  | ~\new_[8429]_ );
  assign \new_[13922]_  = ~\new_[13923]_  | ~\new_[13924]_ ;
  assign \new_[13923]_  = ~\new_[14081]_  | ~\new_[8848]_ ;
  assign \new_[13924]_  = ~\new_[13925]_  | ~\new_[14010]_ ;
  assign \new_[13925]_  = ~\new_[10171]_  | ~\new_[13926]_  | ~\new_[11155]_ ;
  assign \new_[13926]_  = \new_[10261]_  & \new_[11752]_ ;
  assign \new_[13927]_  = ~\new_[13955]_ ;
  assign \new_[13928]_  = ~\new_[14010]_ ;
  assign \new_[13929]_  = ~\new_[13930]_ ;
  assign \new_[13930]_  = ~\new_[13933]_ ;
  assign \new_[13931]_  = ~\new_[13933]_ ;
  assign \new_[13932]_  = ~\new_[13933]_ ;
  assign \new_[13933]_  = \new_[13067]_ ;
  assign \new_[13934]_  = ~\new_[11541]_  | ~\new_[10834]_  | ~\new_[10888]_  | ~\new_[11213]_ ;
  assign \new_[13935]_  = \new_[13936]_ ;
  assign \new_[13936]_  = ~\new_[5041]_  & ~\new_[13798]_ ;
  assign \new_[13937]_  = ~\new_[12294]_  | ~\new_[11119]_  | ~\new_[10833]_  | ~\new_[11198]_ ;
  assign \new_[13938]_  = ~\new_[13962]_  | (~\new_[13939]_  & ~\new_[13942]_ );
  assign \new_[13939]_  = ~\new_[14133]_  & (~\new_[13940]_  | ~\new_[13941]_ );
  assign \new_[13940]_  = ~\new_[8743]_  | ~\new_[2831]_ ;
  assign \new_[13941]_  = ~\new_[14127]_  | ~\new_[8893]_ ;
  assign \new_[13942]_  = ~\new_[8412]_  | (~\new_[8744]_  & ~\new_[12579]_ );
  assign \new_[13943]_  = ~\new_[13955]_  | (~\new_[13944]_  & ~\new_[13947]_ );
  assign \new_[13944]_  = ~\new_[13952]_  & (~\new_[13945]_  | ~\new_[13946]_ );
  assign \new_[13945]_  = ~\new_[13622]_  | ~\new_[8724]_ ;
  assign \new_[13946]_  = ~\new_[3023]_  | ~\new_[8912]_ ;
  assign \new_[13947]_  = ~\new_[14075]_  | (~\new_[8460]_  & ~\new_[13928]_ );
  assign \new_[13948]_  = ~\new_[13955]_  | (~\new_[13949]_  & ~\new_[13954]_ );
  assign \new_[13949]_  = ~\new_[13952]_  & (~\new_[13950]_  | ~\new_[13951]_ );
  assign \new_[13950]_  = ~\new_[8704]_  | ~\new_[3023]_ ;
  assign \new_[13951]_  = ~\new_[13677]_  | ~\new_[8707]_ ;
  assign \new_[13952]_  = ~\new_[13953]_ ;
  assign \new_[13953]_  = ~\new_[5076]_  & ~\new_[4902]_ ;
  assign \new_[13954]_  = ~\new_[8360]_  | (~\new_[8461]_  & ~\new_[13928]_ );
  assign \new_[13955]_  = \new_[13956]_ ;
  assign \new_[13956]_  = ~\new_[4981]_  & ~\new_[6785]_ ;
  assign \new_[13957]_  = ~\new_[13962]_  | (~\new_[13958]_  & ~\new_[13961]_ );
  assign \new_[13958]_  = ~\new_[14133]_  & (~\new_[13959]_  | ~\new_[13960]_ );
  assign \new_[13959]_  = ~\new_[8756]_  | ~\new_[2831]_ ;
  assign \new_[13960]_  = ~\new_[14127]_  | ~\new_[8866]_ ;
  assign \new_[13961]_  = ~\new_[8386]_  | (~\new_[8903]_  & ~\new_[12854]_ );
  assign \new_[13962]_  = \new_[14061]_ ;
  assign \new_[13963]_  = ~\new_[13967]_  | ~\new_[13966]_  | ~\new_[13964]_  | ~\new_[13965]_ ;
  assign \new_[13964]_  = ~\new_[13972]_  | ~\new_[5610]_ ;
  assign \new_[13965]_  = ~\new_[12446]_  | ~\new_[5398]_ ;
  assign \new_[13966]_  = ~\new_[12593]_  | ~\new_[5422]_ ;
  assign \new_[13967]_  = ~\new_[13968]_  | ~\new_[5373]_ ;
  assign \new_[13968]_  = ~\new_[13969]_ ;
  assign \new_[13969]_  = \new_[13970]_ ;
  assign \new_[13970]_  = ~\new_[13871]_  | ~\new_[13589]_ ;
  assign \new_[13971]_  = ~\new_[13970]_ ;
  assign \new_[13972]_  = \new_[14018]_ ;
  assign \new_[13973]_  = ~\new_[14188]_ ;
  assign \new_[13974]_  = ~\new_[14031]_ ;
  assign \new_[13975]_  = ~\new_[13979]_ ;
  assign \new_[13976]_  = ~\new_[13979]_ ;
  assign \new_[13977]_  = ~\new_[13975]_ ;
  assign \new_[13978]_  = ~\new_[13979]_ ;
  assign \new_[13979]_  = ~\new_[13987]_ ;
  assign \new_[13980]_  = ~\new_[13981]_ ;
  assign \new_[13981]_  = \new_[13987]_ ;
  assign \new_[13982]_  = ~\new_[13985]_ ;
  assign \new_[13983]_  = ~\new_[13985]_ ;
  assign \new_[13984]_  = ~\new_[13985]_ ;
  assign \new_[13985]_  = ~\new_[13987]_ ;
  assign \new_[13986]_  = \new_[13987]_ ;
  assign \new_[13987]_  = ~\new_[13890]_ ;
  assign \new_[13988]_  = ~\new_[13991]_ ;
  assign \new_[13989]_  = ~\new_[13990]_ ;
  assign \new_[13990]_  = \new_[13991]_ ;
  assign \new_[13991]_  = ~\new_[2752]_ ;
  assign \new_[13992]_  = ~\new_[13995]_ ;
  assign \new_[13993]_  = ~\new_[13995]_ ;
  assign \new_[13994]_  = ~\new_[13995]_ ;
  assign \new_[13995]_  = ~\new_[13996]_ ;
  assign \new_[13996]_  = ~\new_[13000]_ ;
  assign \new_[13997]_  = ~\new_[13998]_  | ~\new_[14000]_ ;
  assign \new_[13998]_  = ~\new_[13999]_ ;
  assign \new_[13999]_  = ~\new_[2771]_ ;
  assign \new_[14000]_  = ~\new_[2755]_ ;
  assign \new_[14001]_  = \new_[14163]_  | \new_[14088]_ ;
  assign \new_[14002]_  = ~\new_[13823]_  & ~\new_[4980]_ ;
  assign \new_[14003]_  = ~\new_[14004]_ ;
  assign \new_[14004]_  = ~\new_[7636]_ ;
  assign \new_[14005]_  = ~\new_[14003]_ ;
  assign \new_[14006]_  = ~\new_[14007]_  | ~\new_[14009]_ ;
  assign \new_[14007]_  = ~\new_[14081]_  | ~\new_[14008]_ ;
  assign \new_[14008]_  = ~\new_[13889]_  | ~\new_[13887]_ ;
  assign \new_[14009]_  = ~\new_[14167]_  | ~\new_[14010]_ ;
  assign \new_[14010]_  = \new_[13408]_  & \new_[5076]_ ;
  assign \new_[14011]_  = ~\new_[14015]_  | ~\new_[14014]_  | ~\new_[14012]_  | ~\new_[14013]_ ;
  assign \new_[14012]_  = ~\new_[12446]_  | ~\new_[5402]_ ;
  assign \new_[14013]_  = ~\new_[14118]_  | ~\new_[5426]_ ;
  assign \new_[14014]_  = ~\new_[5377]_  | ~\new_[13968]_ ;
  assign \new_[14015]_  = ~\new_[14016]_  | ~\new_[4840]_ ;
  assign \new_[14016]_  = ~\new_[14017]_ ;
  assign \new_[14017]_  = ~\new_[14018]_ ;
  assign \new_[14018]_  = \new_[13589]_  & \new_[13872]_ ;
  assign \new_[14019]_  = ~\new_[14017]_ ;
  assign n2001 = ~\new_[14023]_  | (~\new_[14021]_  & ~\new_[4724]_ );
  assign \new_[14021]_  = ~\new_[4495]_  | ~\new_[14022]_ ;
  assign \new_[14022]_  = ~\dma_ack_i[6] ;
  assign \new_[14023]_  = ~\dma_req_o[6]  | ~\new_[14022]_ ;
  assign n4636 = ~\new_[4724]_  & ~\dma_ack_i[6] ;
  assign n2006 = ~\new_[14028]_  | (~\new_[14026]_  & ~\new_[4725]_ );
  assign \new_[14026]_  = ~\new_[4496]_  | ~\new_[14027]_ ;
  assign \new_[14027]_  = ~\dma_ack_i[7] ;
  assign \new_[14028]_  = ~\dma_req_o[7]  | ~\new_[14027]_ ;
  assign n4641 = ~\new_[4725]_  & ~\dma_ack_i[7] ;
  assign \new_[14030]_  = ~\new_[14031]_ ;
  assign \new_[14031]_  = ~\new_[14032]_ ;
  assign \new_[14032]_  = ~\new_[13600]_  | ~\new_[13844]_ ;
  assign \new_[14033]_  = ~\new_[14030]_ ;
  assign \new_[14034]_  = ~\new_[14035]_  | ~\new_[14036]_ ;
  assign \new_[14035]_  = ~\new_[14090]_ ;
  assign \new_[14036]_  = ~\new_[2792]_ ;
  assign \new_[14037]_  = \new_[14036]_ ;
  assign \new_[14038]_  = ~\new_[14042]_  | ~\new_[14041]_  | ~\new_[14039]_  | ~\new_[14040]_ ;
  assign \new_[14039]_  = ~\new_[12022]_  | ~\new_[5454]_ ;
  assign \new_[14040]_  = ~\new_[12608]_  | ~\new_[4851]_ ;
  assign \new_[14041]_  = ~\new_[12781]_  | ~\new_[5502]_ ;
  assign \new_[14042]_  = ~\new_[14134]_  | ~\new_[5478]_ ;
  assign \new_[14043]_  = ~\new_[4473]_  | (~\new_[14044]_  & ~\new_[14045]_ );
  assign \new_[14044]_  = ~\new_[8392]_  | (~\new_[8750]_  & ~\new_[12363]_ );
  assign \new_[14045]_  = ~\new_[14046]_  | ~\new_[14048]_ ;
  assign \new_[14046]_  = ~\new_[14047]_  | (~\new_[9329]_  & ~\new_[9328]_ );
  assign \new_[14047]_  = \new_[13140]_  & \new_[14087]_ ;
  assign \new_[14048]_  = ~\new_[13934]_  | ~\new_[14087]_  | ~\new_[13500]_ ;
  assign \new_[14049]_  = ~\new_[14050]_  | ~\new_[14052]_ ;
  assign \new_[14050]_  = ~\new_[14051]_  | (~\new_[8984]_  & ~\new_[9304]_ );
  assign \new_[14051]_  = ~\new_[14133]_  & ~\new_[14127]_ ;
  assign \new_[14052]_  = ~\new_[14053]_  | ~\new_[14054]_ ;
  assign \new_[14053]_  = ~\new_[2831]_  & ~\new_[14133]_ ;
  assign \new_[14054]_  = ~\new_[12387]_  | ~\new_[11690]_  | ~\new_[10280]_  | ~\new_[11054]_ ;
  assign \new_[14055]_  = ~\new_[14060]_  | (~\new_[14056]_  & ~\new_[14059]_ );
  assign \new_[14056]_  = ~\new_[14133]_  & (~\new_[14057]_  | ~\new_[14058]_ );
  assign \new_[14057]_  = ~\new_[14127]_  | ~\new_[8902]_ ;
  assign \new_[14058]_  = ~\new_[14038]_  | ~\new_[12717]_ ;
  assign \new_[14059]_  = ~\new_[8634]_  | (~\new_[8903]_  & ~\new_[12579]_ );
  assign \new_[14060]_  = \new_[14061]_ ;
  assign \new_[14061]_  = \new_[14062]_ ;
  assign \new_[14062]_  = ~\new_[14063]_ ;
  assign \new_[14063]_  = \new_[4984]_  | \new_[6788]_ ;
  assign \new_[14064]_  = ~\new_[14068]_  | ~\new_[14067]_  | ~\new_[14065]_  | ~\new_[14066]_ ;
  assign \new_[14065]_  = ~\new_[12023]_  | ~\new_[5466]_ ;
  assign \new_[14066]_  = ~\new_[12635]_  | ~\new_[4855]_ ;
  assign \new_[14067]_  = ~\new_[12821]_  | ~\new_[5515]_ ;
  assign \new_[14068]_  = ~\new_[14134]_  | ~\new_[5490]_ ;
  assign \new_[14069]_  = ~\new_[13153]_  | ~\new_[13999]_ ;
  assign \new_[14070]_  = ~\new_[14106]_  | (~\new_[14071]_  & ~\new_[14074]_ );
  assign \new_[14071]_  = ~\new_[14103]_  & (~\new_[14072]_  | ~\new_[14073]_ );
  assign \new_[14072]_  = ~\new_[3024]_  | ~\new_[14147]_ ;
  assign \new_[14073]_  = ~\new_[9123]_  | ~\new_[13425]_ ;
  assign \new_[14074]_  = ~\new_[8612]_  | (~\new_[8715]_  & ~\new_[12869]_ );
  assign \new_[14075]_  = ~\new_[14076]_  | ~\new_[14081]_ ;
  assign \new_[14076]_  = ~\new_[14080]_  | ~\new_[14079]_  | ~\new_[14077]_  | ~\new_[14078]_ ;
  assign \new_[14077]_  = ~\new_[14033]_  | ~\new_[4825]_ ;
  assign \new_[14078]_  = ~\new_[5242]_  | ~\new_[13976]_ ;
  assign \new_[14079]_  = ~\new_[13931]_  | ~\new_[5267]_ ;
  assign \new_[14080]_  = ~\new_[12431]_  | ~\new_[5292]_ ;
  assign \new_[14081]_  = ~\new_[5076]_  & ~\new_[13408]_ ;
  assign \new_[14082]_  = ~\new_[4473]_  | (~\new_[14083]_  & ~\new_[14084]_ );
  assign \new_[14083]_  = ~\new_[8389]_  | (~\new_[8712]_  & ~\new_[12363]_ );
  assign \new_[14084]_  = ~\new_[14085]_  | ~\new_[14089]_ ;
  assign \new_[14085]_  = ~\new_[14086]_  | (~\new_[9850]_  & ~\new_[9851]_ );
  assign \new_[14086]_  = \new_[13140]_  & \new_[14087]_ ;
  assign \new_[14087]_  = \new_[14088]_ ;
  assign \new_[14088]_  = \new_[13463]_  & \new_[13798]_ ;
  assign \new_[14089]_  = ~\new_[8908]_  | ~\new_[13500]_  | ~\new_[14087]_ ;
  assign \new_[14090]_  = ~\new_[2751]_ ;
  assign \new_[14091]_  = ~\new_[2792]_ ;
  assign n1366 = ~\new_[12402]_  & ~\new_[14095]_ ;
  assign \new_[14093]_  = \new_[14094]_ ;
  assign \new_[14094]_  = ~\new_[5841]_ ;
  assign \new_[14095]_  = ~\new_[14098]_  & (~\new_[14096]_  | ~\new_[14097]_ );
  assign \new_[14096]_  = ~\new_[10487]_  | ~\new_[11471]_ ;
  assign \new_[14097]_  = \new_[4666]_  & \new_[12919]_ ;
  assign \new_[14098]_  = ~\new_[14097]_  & ~\new_[3790]_ ;
  assign \new_[14099]_  = ~\new_[14106]_  | (~\new_[14100]_  & ~\new_[14105]_ );
  assign \new_[14100]_  = ~\new_[14103]_  & (~\new_[14101]_  | ~\new_[14102]_ );
  assign \new_[14101]_  = ~\new_[13425]_  | ~\new_[9114]_ ;
  assign \new_[14102]_  = ~\new_[3024]_  | ~\new_[8869]_ ;
  assign \new_[14103]_  = ~\new_[14104]_ ;
  assign \new_[14104]_  = \new_[13489]_  & \new_[13820]_ ;
  assign \new_[14105]_  = ~\new_[8610]_  | (~\new_[8849]_  & ~\new_[12869]_ );
  assign \new_[14106]_  = \new_[14107]_ ;
  assign \new_[14107]_  = \new_[14108]_ ;
  assign \new_[14108]_  = ~\new_[4982]_  & ~\new_[6786]_ ;
  assign \new_[14109]_  = ~\new_[14113]_  | ~\new_[14112]_  | ~\new_[14110]_  | ~\new_[14111]_ ;
  assign \new_[14110]_  = ~\new_[12354]_  | ~\new_[5541]_ ;
  assign \new_[14111]_  = ~\new_[14189]_  | ~\new_[4859]_ ;
  assign \new_[14112]_  = ~\new_[12830]_  | ~\new_[5200]_ ;
  assign \new_[14113]_  = ~\new_[14115]_  | ~\new_[5171]_ ;
  assign \new_[14114]_  = \new_[13478]_  & \new_[2753]_ ;
  assign \new_[14115]_  = ~\new_[12643]_ ;
  assign \new_[14116]_  = ~\new_[14122]_  | ~\new_[14117]_  | ~\new_[14121]_ ;
  assign \new_[14117]_  = (~\new_[5401]_  | ~\new_[12585]_ ) & (~\new_[14118]_  | ~\new_[5425]_ );
  assign \new_[14118]_  = ~\new_[14119]_ ;
  assign \new_[14119]_  = ~\new_[14120]_ ;
  assign \new_[14120]_  = ~\new_[13872]_  & ~\new_[13584]_ ;
  assign \new_[14121]_  = ~\new_[14019]_  | ~\new_[4839]_ ;
  assign \new_[14122]_  = ~\new_[13968]_  | ~\new_[5376]_ ;
  assign \new_[14123]_  = ~\new_[14124]_  | ~\new_[14126]_ ;
  assign \new_[14124]_  = ~\new_[2831]_  | ~\new_[14125]_  | ~\new_[14131]_ ;
  assign \new_[14125]_  = ~\new_[12411]_  | ~\new_[11142]_  | ~\new_[10231]_  | ~\new_[10220]_ ;
  assign \new_[14126]_  = ~\new_[13891]_  | ~\new_[14127]_  | ~\new_[14131]_ ;
  assign \new_[14127]_  = ~\new_[2831]_ ;
  assign \new_[14128]_  = ~\new_[14129]_  | ~\new_[14132]_ ;
  assign \new_[14129]_  = ~\new_[2831]_  | ~\new_[14130]_  | ~\new_[14131]_ ;
  assign \new_[14130]_  = ~\new_[12284]_  | ~\new_[12096]_  | ~\new_[10267]_  | ~\new_[10179]_ ;
  assign \new_[14131]_  = \new_[13278]_  & \new_[13601]_ ;
  assign \new_[14132]_  = ~\new_[9140]_  | ~\new_[14131]_  | ~\new_[14127]_ ;
  assign \new_[14133]_  = ~\new_[14131]_ ;
  assign \new_[14134]_  = \new_[14140]_ ;
  assign \new_[14135]_  = \new_[14140]_ ;
  assign \new_[14136]_  = ~\new_[14139]_ ;
  assign \new_[14137]_  = ~\new_[14138]_ ;
  assign \new_[14138]_  = ~\new_[14139]_ ;
  assign \new_[14139]_  = ~\new_[14140]_ ;
  assign \new_[14140]_  = ~\new_[14069]_ ;
  assign \new_[14141]_  = ~\new_[4473]_  | (~\new_[14142]_  & ~\new_[14143]_ );
  assign \new_[14142]_  = ~\new_[12599]_  & (~\new_[8341]_  | ~\new_[8675]_ );
  assign \new_[14143]_  = ~\new_[14144]_  | ~\new_[14146]_ ;
  assign \new_[14144]_  = ~\new_[14145]_  | ~\new_[14176]_ ;
  assign \new_[14145]_  = \new_[13798]_  & \new_[5041]_ ;
  assign \new_[14146]_  = ~\new_[8892]_  | ~\new_[13935]_ ;
  assign \new_[14147]_  = ~\new_[14151]_  | ~\new_[14150]_  | ~\new_[14148]_  | ~\new_[14149]_ ;
  assign \new_[14148]_  = ~\new_[12417]_  | ~\new_[5305]_ ;
  assign \new_[14149]_  = ~\new_[14188]_  | ~\new_[5329]_ ;
  assign \new_[14150]_  = ~\new_[12789]_  | ~\new_[5354]_ ;
  assign \new_[14151]_  = ~\new_[14152]_  | ~\new_[5598]_ ;
  assign \new_[14152]_  = \new_[14153]_ ;
  assign \new_[14153]_  = ~\new_[14154]_ ;
  assign \new_[14154]_  = ~\new_[14091]_  | ~\new_[14090]_ ;
  assign \new_[14155]_  = ~\new_[14153]_ ;
  assign \new_[14156]_  = ~\new_[14161]_  | (~\new_[14157]_  & ~\new_[14158]_ );
  assign \new_[14157]_  = ~\new_[12599]_  & (~\new_[8323]_  | ~\new_[8683]_ );
  assign \new_[14158]_  = ~\new_[14159]_  | ~\new_[14160]_ ;
  assign \new_[14159]_  = ~\new_[14145]_  | ~\new_[13934]_ ;
  assign \new_[14160]_  = ~\new_[13935]_  | ~\new_[13937]_ ;
  assign \new_[14161]_  = ~\new_[14162]_ ;
  assign \new_[14162]_  = \new_[14163]_ ;
  assign \new_[14163]_  = ~\new_[14002]_  | ~\new_[14003]_ ;
  assign \new_[14164]_  = \new_[14166]_ ;
  assign \new_[14165]_  = ~\new_[14166]_ ;
  assign \new_[14166]_  = ~\new_[13031]_ ;
  assign \new_[14167]_  = ~\new_[14171]_  | ~\new_[14170]_  | ~\new_[14168]_  | ~\new_[14169]_ ;
  assign \new_[14168]_  = ~\new_[14033]_  | ~\new_[4818]_ ;
  assign \new_[14169]_  = ~\new_[13981]_  | ~\new_[5224]_ ;
  assign \new_[14170]_  = ~\new_[5249]_  | ~\new_[13930]_ ;
  assign \new_[14171]_  = ~\new_[14172]_  | ~\new_[5274]_ ;
  assign \new_[14172]_  = \new_[14173]_ ;
  assign \new_[14173]_  = ~\new_[14174]_ ;
  assign \new_[14174]_  = ~\new_[13093]_  | ~\new_[2750]_ ;
  assign \new_[14175]_  = ~\new_[14173]_ ;
  assign \new_[14176]_  = ~\new_[14180]_  | ~\new_[14179]_  | ~\new_[14177]_  | ~\new_[14178]_ ;
  assign \new_[14177]_  = ~\new_[14189]_  | ~\new_[5857]_ ;
  assign \new_[14178]_  = ~\new_[12360]_  | ~\new_[5175]_ ;
  assign \new_[14179]_  = ~\new_[5202]_  | ~\new_[12657]_ ;
  assign \new_[14180]_  = ~\new_[14181]_  | ~\new_[5545]_ ;
  assign \new_[14181]_  = \new_[14182]_ ;
  assign \new_[14182]_  = ~\new_[14183]_ ;
  assign \new_[14183]_  = ~\new_[13143]_  | ~\new_[13683]_ ;
  assign \new_[14184]_  = \new_[13569]_  | \new_[13223]_ ;
  assign \new_[14185]_  = \new_[13569]_  | \new_[13223]_ ;
  assign \new_[14186]_  = \new_[13655]_  | \new_[13437]_ ;
  assign \new_[14187]_  = \new_[13655]_  | \new_[13437]_ ;
  assign \new_[14188]_  = ~\new_[14034]_ ;
  assign \new_[14189]_  = ~\new_[14165]_ ;
  assign \new_[14190]_  = ~\new_[14165]_ ;
  assign \new_[14191]_  = ~\new_[13974]_ ;
  assign \new_[14192]_  = ~\new_[13974]_ ;
  assign \new_[14193]_  = \new_[5877]_ ;
  assign \new_[14194]_  = \new_[6443]_ ;
  assign n11091 = sdata_pad_i;
  assign n11096 = \wb_data_i[7] ;
  assign n11101 = \wb_data_i[4] ;
  assign n11106 = \wb_data_i[12] ;
  assign n11111 = \wb_data_i[24] ;
  assign n11116 = \wb_data_i[26] ;
  assign n11121 = \wb_data_i[23] ;
  assign n11126 = \wb_data_i[11] ;
  assign n11131 = \wb_data_i[31] ;
  assign n11136 = \wb_data_i[13] ;
  assign n11141 = \wb_data_i[29] ;
  assign n11146 = \wb_data_i[22] ;
  assign n11151 = \wb_data_i[30] ;
  assign n11156 = \wb_data_i[15] ;
  assign n11161 = \wb_data_i[19] ;
  assign n11166 = bit_clk_pad_i;
  assign n11171 = \wb_data_i[27] ;
  assign n11176 = \wb_data_i[28] ;
  assign n11181 = \wb_data_i[10] ;
  assign n11186 = \wb_data_i[6] ;
  assign n11191 = \wb_data_i[20] ;
  assign n11196 = \wb_data_i[0] ;
  assign n11201 = \wb_data_i[21] ;
  assign n11206 = \wb_data_i[5] ;
  assign n11211 = \wb_data_i[18] ;
  assign n11216 = \wb_data_i[25] ;
  assign n11221 = \wb_data_i[2] ;
  assign n11226 = \wb_data_i[9] ;
  assign n11231 = \wb_data_i[17] ;
  assign n11236 = \wb_data_i[3] ;
  assign n11241 = \wb_data_i[8] ;
  assign n11246 = \wb_data_i[16] ;
  assign n11251 = \wb_data_i[14] ;
  assign n11256 = \wb_data_i[1] ;
  always @ (posedge clock) begin
    \\u0_slt0_r_reg[15]  <= n266;
    \\u0_slt0_r_reg[14]  <= n271;
    \\u0_slt0_r_reg[13]  <= n276;
    \\u0_slt0_r_reg[12]  <= n281;
    \\u0_slt0_r_reg[11]  <= n286;
    \\u0_slt0_r_reg[10]  <= n291;
    \\u0_slt0_r_reg[9]  <= n296;
    \\u0_slt0_r_reg[8]  <= n301;
    \\u0_slt0_r_reg[7]  <= n306;
    \\u0_slt0_r_reg[6]  <= n311;
    \\u0_slt0_r_reg[5]  <= n316;
    \\u0_slt0_r_reg[4]  <= n321;
    \\u0_slt0_r_reg[3]  <= n326;
    \\u0_slt0_r_reg[2]  <= n331;
    \\u0_slt0_r_reg[1]  <= n336;
    \\u0_slt0_r_reg[0]  <= n341;
    \\u0_slt1_r_reg[19]  <= n346;
    \\u0_slt1_r_reg[18]  <= n351;
    \\u0_slt1_r_reg[17]  <= n356;
    \\u0_slt1_r_reg[16]  <= n361;
    \\u0_slt1_r_reg[15]  <= n366;
    \\u0_slt1_r_reg[14]  <= n371;
    \\u0_slt1_r_reg[13]  <= n376;
    \\u0_slt1_r_reg[12]  <= n381;
    \\u0_slt1_r_reg[11]  <= n386;
    \\u0_slt1_r_reg[10]  <= n391;
    \\u0_slt1_r_reg[9]  <= n396;
    \\u0_slt1_r_reg[8]  <= n401;
    \\u0_slt1_r_reg[7]  <= n406;
    \\u0_slt1_r_reg[6]  <= n411;
    \\u0_slt1_r_reg[5]  <= n416;
    \\u0_slt1_r_reg[4]  <= n421;
    \\u0_slt1_r_reg[3]  <= n426;
    \\u0_slt1_r_reg[2]  <= n431;
    \\u0_slt1_r_reg[1]  <= n436;
    \\u0_slt1_r_reg[0]  <= n441;
    \\u0_slt2_r_reg[19]  <= n446;
    \\u0_slt2_r_reg[18]  <= n451;
    \\u0_slt2_r_reg[17]  <= n456;
    \\u0_slt2_r_reg[16]  <= n461;
    \\u0_slt2_r_reg[15]  <= n466;
    \\u0_slt2_r_reg[14]  <= n471;
    \\u0_slt2_r_reg[13]  <= n476;
    \\u0_slt2_r_reg[12]  <= n481;
    \\u0_slt2_r_reg[11]  <= n486;
    \\u0_slt2_r_reg[10]  <= n491;
    \\u0_slt2_r_reg[9]  <= n496;
    \\u0_slt2_r_reg[8]  <= n501;
    \\u0_slt2_r_reg[7]  <= n506;
    \\u0_slt2_r_reg[6]  <= n511;
    \\u0_slt2_r_reg[5]  <= n516;
    \\u0_slt2_r_reg[4]  <= n521;
    \\u0_slt2_r_reg[3]  <= n526;
    \\u0_slt2_r_reg[2]  <= n531;
    \\u0_slt2_r_reg[1]  <= n536;
    \\u0_slt2_r_reg[0]  <= n541;
    \\u0_slt3_r_reg[19]  <= n546;
    \\u0_slt3_r_reg[18]  <= n551;
    \\u0_slt3_r_reg[17]  <= n556;
    \\u0_slt3_r_reg[16]  <= n561;
    \\u0_slt3_r_reg[15]  <= n566;
    \\u0_slt3_r_reg[14]  <= n571;
    \\u0_slt3_r_reg[13]  <= n576;
    \\u0_slt3_r_reg[12]  <= n581;
    \\u0_slt3_r_reg[11]  <= n586;
    \\u0_slt3_r_reg[10]  <= n591;
    \\u0_slt3_r_reg[9]  <= n596;
    \\u0_slt3_r_reg[8]  <= n601;
    \\u0_slt3_r_reg[7]  <= n606;
    \\u0_slt3_r_reg[6]  <= n611;
    \\u0_slt3_r_reg[5]  <= n616;
    \\u0_slt3_r_reg[4]  <= n621;
    \\u0_slt3_r_reg[3]  <= n626;
    \\u0_slt3_r_reg[2]  <= n631;
    \\u0_slt3_r_reg[1]  <= n636;
    \\u0_slt3_r_reg[0]  <= n641;
    \\u0_slt4_r_reg[19]  <= n646;
    \\u0_slt4_r_reg[18]  <= n651;
    \\u0_slt4_r_reg[17]  <= n656;
    \\u0_slt4_r_reg[16]  <= n661;
    \\u0_slt4_r_reg[15]  <= n666;
    \\u0_slt4_r_reg[14]  <= n671;
    \\u0_slt4_r_reg[13]  <= n676;
    \\u0_slt4_r_reg[12]  <= n681;
    \\u0_slt4_r_reg[11]  <= n686;
    \\u0_slt4_r_reg[10]  <= n691;
    \\u0_slt4_r_reg[9]  <= n696;
    \\u0_slt4_r_reg[8]  <= n701;
    \\u0_slt4_r_reg[7]  <= n706;
    \\u0_slt4_r_reg[6]  <= n711;
    \\u0_slt4_r_reg[5]  <= n716;
    \\u0_slt4_r_reg[4]  <= n721;
    \\u0_slt4_r_reg[3]  <= n726;
    \\u0_slt4_r_reg[2]  <= n731;
    \\u0_slt4_r_reg[1]  <= n736;
    \\u0_slt4_r_reg[0]  <= n741;
    \\u0_slt5_r_reg[19]  <= n746;
    \\u0_slt5_r_reg[18]  <= n751;
    \\u0_slt5_r_reg[17]  <= n756;
    \\u0_slt5_r_reg[16]  <= n761;
    \\u0_slt5_r_reg[15]  <= n766;
    \\u0_slt5_r_reg[14]  <= n771;
    \\u0_slt5_r_reg[13]  <= n776;
    \\u0_slt5_r_reg[12]  <= n781;
    \\u0_slt5_r_reg[11]  <= n786;
    \\u0_slt5_r_reg[10]  <= n791;
    \\u0_slt5_r_reg[9]  <= n796;
    \\u0_slt5_r_reg[8]  <= n801;
    \\u0_slt5_r_reg[7]  <= n806;
    \\u0_slt5_r_reg[6]  <= n811;
    \\u0_slt5_r_reg[5]  <= n816;
    \\u0_slt5_r_reg[4]  <= n821;
    \\u0_slt5_r_reg[3]  <= n826;
    \\u0_slt5_r_reg[2]  <= n831;
    \\u0_slt5_r_reg[1]  <= n836;
    \\u0_slt5_r_reg[0]  <= n841;
    \\u0_slt6_r_reg[19]  <= n846;
    \\u0_slt6_r_reg[18]  <= n851;
    \\u0_slt6_r_reg[17]  <= n856;
    \\u0_slt6_r_reg[16]  <= n861;
    \\u0_slt6_r_reg[15]  <= n866;
    \\u0_slt6_r_reg[14]  <= n871;
    \\u0_slt6_r_reg[13]  <= n876;
    \\u0_slt6_r_reg[12]  <= n881;
    \\u0_slt6_r_reg[11]  <= n886;
    \\u0_slt6_r_reg[10]  <= n891;
    \\u0_slt6_r_reg[9]  <= n896;
    \\u0_slt6_r_reg[8]  <= n901;
    \\u0_slt6_r_reg[7]  <= n906;
    \\u0_slt6_r_reg[6]  <= n911;
    \\u0_slt6_r_reg[5]  <= n916;
    \\u0_slt6_r_reg[4]  <= n921;
    \\u0_slt6_r_reg[3]  <= n926;
    \\u0_slt6_r_reg[2]  <= n931;
    \\u0_slt6_r_reg[1]  <= n936;
    \\u0_slt6_r_reg[0]  <= n941;
    \\u0_slt7_r_reg[19]  <= n946;
    \\u0_slt7_r_reg[18]  <= n951;
    \\u0_slt7_r_reg[17]  <= n956;
    \\u0_slt7_r_reg[16]  <= n961;
    \\u0_slt7_r_reg[15]  <= n966;
    \\u0_slt7_r_reg[14]  <= n971;
    \\u0_slt7_r_reg[13]  <= n976;
    \\u0_slt7_r_reg[12]  <= n981;
    \\u0_slt7_r_reg[11]  <= n986;
    \\u0_slt7_r_reg[10]  <= n991;
    \\u0_slt7_r_reg[9]  <= n996;
    \\u0_slt7_r_reg[8]  <= n1001;
    \\u0_slt7_r_reg[7]  <= n1006;
    \\u0_slt7_r_reg[6]  <= n1011;
    \\u0_slt7_r_reg[5]  <= n1016;
    \\u0_slt7_r_reg[4]  <= n1021;
    \\u0_slt7_r_reg[3]  <= n1026;
    \\u0_slt7_r_reg[2]  <= n1031;
    \\u0_slt7_r_reg[1]  <= n1036;
    \\u0_slt7_r_reg[0]  <= n1041;
    \\u0_slt8_r_reg[19]  <= n1046;
    \\u0_slt8_r_reg[18]  <= n1051;
    \\u0_slt8_r_reg[17]  <= n1056;
    \\u0_slt8_r_reg[16]  <= n1061;
    \\u0_slt8_r_reg[15]  <= n1066;
    \\u0_slt8_r_reg[14]  <= n1071;
    \\u0_slt8_r_reg[13]  <= n1076;
    \\u0_slt8_r_reg[12]  <= n1081;
    \\u0_slt8_r_reg[11]  <= n1086;
    \\u0_slt8_r_reg[10]  <= n1091;
    \\u0_slt8_r_reg[9]  <= n1096;
    \\u0_slt8_r_reg[8]  <= n1101;
    \\u0_slt8_r_reg[7]  <= n1106;
    \\u0_slt8_r_reg[6]  <= n1111;
    \\u0_slt8_r_reg[5]  <= n1116;
    \\u0_slt8_r_reg[4]  <= n1121;
    \\u0_slt8_r_reg[3]  <= n1126;
    \\u0_slt8_r_reg[2]  <= n1131;
    \\u0_slt8_r_reg[1]  <= n1136;
    \\u0_slt8_r_reg[0]  <= n1141;
    \\u0_slt9_r_reg[19]  <= n1146;
    \\u0_slt9_r_reg[18]  <= n1151;
    \\u0_slt9_r_reg[17]  <= n1156;
    \\u0_slt9_r_reg[16]  <= n1161;
    \\u0_slt9_r_reg[15]  <= n1166;
    \\u0_slt9_r_reg[14]  <= n1171;
    \\u0_slt9_r_reg[13]  <= n1176;
    \\u0_slt9_r_reg[12]  <= n1181;
    \\u0_slt9_r_reg[11]  <= n1186;
    \\u0_slt9_r_reg[10]  <= n1191;
    \\u0_slt9_r_reg[9]  <= n1196;
    \\u0_slt9_r_reg[8]  <= n1201;
    \\u0_slt9_r_reg[7]  <= n1206;
    \\u0_slt9_r_reg[6]  <= n1211;
    \\u1_slt2_reg[19]  <= n1216;
    \\u1_slt3_reg[19]  <= n1221;
    \\u1_slt4_reg[19]  <= n1226;
    \\u1_slt6_reg[19]  <= n1231;
    \\u1_slt2_reg[18]  <= n1236;
    \\u1_slt3_reg[18]  <= n1241;
    \\u1_slt4_reg[18]  <= n1246;
    \\u1_slt6_reg[18]  <= n1251;
    u16_u1_dma_req_reg <= n1256;
    u16_u3_dma_req_reg <= n1261;
    \\u0_slt9_r_reg[5]  <= n1266;
    u16_u0_dma_req_reg <= n1271;
    u16_u2_dma_req_reg <= n1276;
    u16_u4_dma_req_reg <= n1281;
    u16_u5_dma_req_reg <= n1286;
    \\u1_slt2_reg[17]  <= n1291;
    \\u1_slt3_reg[17]  <= n1296;
    \\u1_slt4_reg[17]  <= n1301;
    \\u1_slt6_reg[17]  <= n1306;
    \\u1_sr_reg[19]  <= n1311;
    \\u1_slt2_reg[16]  <= n1316;
    \\u1_slt3_reg[16]  <= n1321;
    \\u1_slt4_reg[16]  <= n1326;
    \\u1_slt6_reg[16]  <= n1331;
    \\u4_rp_reg[2]  <= n1336;
    \\u5_rp_reg[2]  <= n1341;
    \\u8_rp_reg[2]  <= n1346;
    \\u3_rp_reg[2]  <= n1351;
    \\u6_rp_reg[2]  <= n1356;
    \\u7_rp_reg[2]  <= n1361;
    \\u8_rp_reg[3]  <= n1366;
    \\u3_rp_reg[3]  <= n1371;
    \\u6_rp_reg[3]  <= n1376;
    \\u7_rp_reg[3]  <= n1381;
    \\u8_rp_reg[1]  <= n1386;
    \\u3_rp_reg[1]  <= n1391;
    \\u7_rp_reg[1]  <= n1396;
    \\u6_rp_reg[1]  <= n1401;
    \\u1_sr_reg[18]  <= n1406;
    \\u13_ints_r_reg[11]  <= n1411;
    \\u13_ints_r_reg[5]  <= n1416;
    \\u1_slt3_reg[15]  <= n1421;
    \\u1_slt0_reg[15]  <= n1426;
    \\u1_slt6_reg[15]  <= n1431;
    \\u1_slt2_reg[15]  <= n1436;
    \\u1_slt4_reg[15]  <= n1441;
    \\u4_rp_reg[1]  <= n1446;
    \\u4_rp_reg[3]  <= n1451;
    \\u5_rp_reg[1]  <= n1456;
    \\u5_rp_reg[3]  <= n1461;
    \\u6_dout_reg[2]  <= n1466;
    \\u6_dout_reg[3]  <= n1471;
    \\u7_dout_reg[2]  <= n1476;
    \\u7_dout_reg[3]  <= n1481;
    \\u3_dout_reg[2]  <= n1486;
    \\u3_dout_reg[3]  <= n1491;
    \\u8_dout_reg[2]  <= n1496;
    \\u8_dout_reg[3]  <= n1501;
    \\u13_ints_r_reg[14]  <= n1506;
    \\u13_ints_r_reg[17]  <= n1511;
    \\u13_ints_r_reg[2]  <= n1516;
    \\u13_ints_r_reg[8]  <= n1521;
    \\u6_dout_reg[0]  <= n1526;
    \\u6_dout_reg[1]  <= n1531;
    \\u7_dout_reg[0]  <= n1536;
    \\u7_dout_reg[1]  <= n1541;
    \\u3_dout_reg[0]  <= n1546;
    \\u8_dout_reg[0]  <= n1551;
    \\u3_dout_reg[1]  <= n1556;
    \\u8_dout_reg[1]  <= n1561;
    \\u8_rp_reg[0]  <= n1566;
    \\u3_rp_reg[0]  <= n1571;
    \\u6_rp_reg[0]  <= n1576;
    \\u7_rp_reg[0]  <= n1581;
    \\u6_dout_reg[12]  <= n1586;
    \\u6_dout_reg[13]  <= n1591;
    \\u6_dout_reg[14]  <= n1596;
    \\u6_dout_reg[15]  <= n1601;
    \\u6_dout_reg[10]  <= n1606;
    \\u6_dout_reg[11]  <= n1611;
    \\u6_dout_reg[18]  <= n1616;
    \\u6_dout_reg[19]  <= n1621;
    \\u6_dout_reg[16]  <= n1626;
    \\u6_dout_reg[17]  <= n1631;
    \\u6_dout_reg[4]  <= n1636;
    \\u6_dout_reg[5]  <= n1641;
    \\u6_dout_reg[6]  <= n1646;
    \\u6_dout_reg[7]  <= n1651;
    \\u6_dout_reg[8]  <= n1656;
    \\u6_dout_reg[9]  <= n1661;
    \\u7_dout_reg[10]  <= n1666;
    \\u7_dout_reg[11]  <= n1671;
    \\u7_dout_reg[12]  <= n1676;
    \\u7_dout_reg[13]  <= n1681;
    \\u7_dout_reg[14]  <= n1686;
    \\u7_dout_reg[17]  <= n1691;
    \\u7_dout_reg[15]  <= n1696;
    \\u7_dout_reg[19]  <= n1701;
    \\u7_dout_reg[16]  <= n1706;
    \\u7_dout_reg[18]  <= n1711;
    \\u7_dout_reg[4]  <= n1716;
    \\u7_dout_reg[5]  <= n1721;
    \\u7_dout_reg[6]  <= n1726;
    \\u7_dout_reg[7]  <= n1731;
    \\u7_dout_reg[8]  <= n1736;
    \\u7_dout_reg[9]  <= n1741;
    \\u3_dout_reg[10]  <= n1746;
    \\u3_dout_reg[11]  <= n1751;
    \\u3_dout_reg[13]  <= n1756;
    \\u3_dout_reg[14]  <= n1761;
    \\u3_dout_reg[15]  <= n1766;
    \\u3_dout_reg[16]  <= n1771;
    \\u3_dout_reg[17]  <= n1776;
    \\u3_dout_reg[18]  <= n1781;
    \\u8_dout_reg[10]  <= n1786;
    \\u3_dout_reg[19]  <= n1791;
    \\u8_dout_reg[11]  <= n1796;
    \\u8_dout_reg[12]  <= n1801;
    \\u3_dout_reg[12]  <= n1806;
    \\u8_dout_reg[13]  <= n1811;
    \\u8_dout_reg[14]  <= n1816;
    \\u3_dout_reg[4]  <= n1821;
    \\u8_dout_reg[16]  <= n1826;
    \\u3_dout_reg[6]  <= n1831;
    \\u8_dout_reg[17]  <= n1836;
    \\u3_dout_reg[7]  <= n1841;
    \\u8_dout_reg[18]  <= n1846;
    \\u3_dout_reg[8]  <= n1851;
    \\u8_dout_reg[15]  <= n1856;
    \\u3_dout_reg[5]  <= n1861;
    \\u8_dout_reg[19]  <= n1866;
    \\u3_dout_reg[9]  <= n1871;
    \\u8_dout_reg[4]  <= n1876;
    \\u8_dout_reg[5]  <= n1881;
    \\u8_dout_reg[6]  <= n1886;
    \\u8_dout_reg[7]  <= n1891;
    \\u8_dout_reg[8]  <= n1896;
    \\u8_dout_reg[9]  <= n1901;
    \\u0_slt9_r_reg[4]  <= n1906;
    u16_u1_dma_req_r1_reg <= n1911;
    u16_u3_dma_req_r1_reg <= n1916;
    \\u1_sr_reg[17]  <= n1921;
    u16_u8_dma_req_reg <= n1926;
    \\u1_slt3_reg[14]  <= n1931;
    \\u1_slt4_reg[14]  <= n1936;
    \\u1_slt6_reg[14]  <= n1941;
    \\u1_slt2_reg[14]  <= n1946;
    \\u4_dout_reg[3]  <= n1951;
    \\u5_dout_reg[3]  <= n1956;
    \\u5_dout_reg[2]  <= n1961;
    \\u4_dout_reg[2]  <= n1966;
    u16_u0_dma_req_r1_reg <= n1971;
    u16_u2_dma_req_r1_reg <= n1976;
    u16_u4_dma_req_r1_reg <= n1981;
    u16_u5_dma_req_r1_reg <= n1986;
    \\u4_dout_reg[4]  <= n1991;
    \\u11_wp_reg[3]  <= n1996;
    u16_u6_dma_req_reg <= n2001;
    u16_u7_dma_req_reg <= n2006;
    \\u5_dout_reg[0]  <= n2011;
    \\u5_dout_reg[1]  <= n2016;
    \\u4_dout_reg[1]  <= n2021;
    \\u4_dout_reg[0]  <= n2026;
    \\u4_rp_reg[0]  <= n2031;
    \\u5_rp_reg[0]  <= n2036;
    \\u11_mem_reg[0][18]  <= n2041;
    \\u11_mem_reg[0][19]  <= n2046;
    \\u11_mem_reg[1][18]  <= n2051;
    \\u11_mem_reg[1][19]  <= n2056;
    \\u11_mem_reg[1][20]  <= n2061;
    \\u11_mem_reg[1][21]  <= n2066;
    \\u11_mem_reg[1][22]  <= n2071;
    \\u11_mem_reg[1][23]  <= n2076;
    \\u11_mem_reg[1][24]  <= n2081;
    \\u11_mem_reg[1][25]  <= n2086;
    \\u11_mem_reg[1][26]  <= n2091;
    \\u11_mem_reg[1][27]  <= n2096;
    \\u11_mem_reg[1][28]  <= n2101;
    \\u11_mem_reg[1][29]  <= n2106;
    \\u11_mem_reg[1][30]  <= n2111;
    \\u11_mem_reg[1][31]  <= n2116;
    \\u11_mem_reg[2][18]  <= n2121;
    \\u11_mem_reg[2][19]  <= n2126;
    \\u11_mem_reg[2][20]  <= n2131;
    \\u11_mem_reg[2][21]  <= n2136;
    \\u11_mem_reg[2][22]  <= n2141;
    \\u11_mem_reg[2][23]  <= n2146;
    \\u11_mem_reg[2][24]  <= n2151;
    \\u11_mem_reg[2][25]  <= n2156;
    \\u11_mem_reg[2][26]  <= n2161;
    \\u11_mem_reg[2][27]  <= n2166;
    \\u11_mem_reg[2][28]  <= n2171;
    \\u11_mem_reg[2][29]  <= n2176;
    \\u11_mem_reg[2][30]  <= n2181;
    \\u11_mem_reg[2][31]  <= n2186;
    \\u11_mem_reg[3][18]  <= n2191;
    \\u11_mem_reg[3][19]  <= n2196;
    \\u11_mem_reg[3][20]  <= n2201;
    \\u11_mem_reg[3][21]  <= n2206;
    \\u11_mem_reg[3][22]  <= n2211;
    \\u11_mem_reg[3][23]  <= n2216;
    \\u11_mem_reg[3][24]  <= n2221;
    \\u11_mem_reg[3][25]  <= n2226;
    \\u11_mem_reg[3][26]  <= n2231;
    \\u11_mem_reg[3][27]  <= n2236;
    \\u11_mem_reg[3][28]  <= n2241;
    \\u11_mem_reg[3][29]  <= n2246;
    \\u11_mem_reg[3][30]  <= n2251;
    \\u11_mem_reg[3][31]  <= n2256;
    \\u11_mem_reg[3][7]  <= n2261;
    \\u11_mem_reg[1][12]  <= n2266;
    \\u11_mem_reg[1][13]  <= n2271;
    \\u11_mem_reg[1][16]  <= n2276;
    \\u11_mem_reg[2][17]  <= n2281;
    \\u11_mem_reg[2][1]  <= n2286;
    \\u11_mem_reg[2][7]  <= n2291;
    \\u11_mem_reg[2][8]  <= n2296;
    \\u11_mem_reg[3][16]  <= n2301;
    \\u11_mem_reg[3][17]  <= n2306;
    \\u11_mem_reg[3][5]  <= n2311;
    \\u11_mem_reg[3][6]  <= n2316;
    \\u11_wp_reg[1]  <= n2321;
    \\u11_wp_reg[2]  <= n2326;
    \\u4_dout_reg[10]  <= n2331;
    \\u4_dout_reg[13]  <= n2336;
    \\u4_dout_reg[14]  <= n2341;
    \\u4_dout_reg[15]  <= n2346;
    \\u4_dout_reg[16]  <= n2351;
    \\u4_dout_reg[11]  <= n2356;
    \\u4_dout_reg[18]  <= n2361;
    \\u4_dout_reg[12]  <= n2366;
    \\u4_dout_reg[19]  <= n2371;
    \\u4_dout_reg[17]  <= n2376;
    \\u4_dout_reg[5]  <= n2381;
    \\u4_dout_reg[6]  <= n2386;
    \\u4_dout_reg[7]  <= n2391;
    \\u4_dout_reg[8]  <= n2396;
    \\u4_dout_reg[9]  <= n2401;
    \\u5_dout_reg[10]  <= n2406;
    \\u5_dout_reg[11]  <= n2411;
    \\u5_dout_reg[12]  <= n2416;
    \\u5_dout_reg[14]  <= n2421;
    \\u5_dout_reg[15]  <= n2426;
    \\u5_dout_reg[16]  <= n2431;
    \\u5_dout_reg[18]  <= n2436;
    \\u5_dout_reg[19]  <= n2441;
    \\u5_dout_reg[4]  <= n2446;
    \\u5_dout_reg[5]  <= n2451;
    \\u5_dout_reg[6]  <= n2456;
    \\u5_dout_reg[8]  <= n2461;
    \\u5_dout_reg[9]  <= n2466;
    \\u11_mem_reg[0][0]  <= n2471;
    \\u11_mem_reg[0][10]  <= n2476;
    \\u11_mem_reg[0][11]  <= n2481;
    \\u11_mem_reg[0][12]  <= n2486;
    \\u11_mem_reg[0][13]  <= n2491;
    \\u11_mem_reg[0][14]  <= n2496;
    \\u11_mem_reg[0][15]  <= n2501;
    \\u11_mem_reg[0][1]  <= n2506;
    u15_crac_rd_reg <= n2511;
    \\u17_int_set_reg[1]  <= n2516;
    \\u20_int_set_reg[1]  <= n2521;
    \\u21_int_set_reg[1]  <= n2526;
    \\u22_int_set_reg[1]  <= n2531;
    \\u5_dout_reg[7]  <= n2536;
    \\u5_dout_reg[17]  <= n2541;
    \\u1_sr_reg[16]  <= n2546;
    \\u5_dout_reg[13]  <= n2551;
    \\u10_mem_reg[0][18]  <= n2556;
    \\u10_mem_reg[3][28]  <= n2561;
    \\u10_mem_reg[3][24]  <= n2566;
    \\u9_mem_reg[3][30]  <= n2571;
    \\u9_mem_reg[3][26]  <= n2576;
    \\u10_wp_reg[3]  <= n2581;
    \\u9_mem_reg[3][22]  <= n2586;
    \\u9_mem_reg[2][28]  <= n2591;
    \\u9_mem_reg[2][24]  <= n2596;
    \\u9_mem_reg[2][20]  <= n2601;
    \\u9_mem_reg[1][28]  <= n2606;
    \\u9_mem_reg[1][25]  <= n2611;
    \\u9_mem_reg[1][22]  <= n2616;
    \\u10_mem_reg[2][24]  <= n2621;
    \\u11_mem_reg[3][14]  <= n2626;
    \\u11_mem_reg[3][0]  <= n2631;
    \\u11_mem_reg[3][13]  <= n2636;
    \\u10_mem_reg[1][0]  <= n2641;
    \\u11_mem_reg[1][15]  <= n2646;
    \\u11_mem_reg[1][6]  <= n2651;
    \\u1_slt2_reg[13]  <= n2656;
    \\u1_slt4_reg[13]  <= n2661;
    \\u1_slt6_reg[13]  <= n2666;
    \\u1_slt3_reg[13]  <= n2671;
    \\u10_mem_reg[2][18]  <= n2676;
    \\u10_mem_reg[2][19]  <= n2681;
    \\u10_mem_reg[2][20]  <= n2686;
    \\u10_mem_reg[2][21]  <= n2691;
    \\u10_mem_reg[2][22]  <= n2696;
    \\u9_mem_reg[0][18]  <= n2701;
    \\u9_mem_reg[0][19]  <= n2706;
    \\u10_mem_reg[2][23]  <= n2711;
    \\u10_mem_reg[2][25]  <= n2716;
    \\u10_mem_reg[2][26]  <= n2721;
    \\u10_mem_reg[2][27]  <= n2726;
    \\u9_mem_reg[1][18]  <= n2731;
    \\u9_mem_reg[1][19]  <= n2736;
    \\u9_mem_reg[1][20]  <= n2741;
    \\u9_mem_reg[1][21]  <= n2746;
    \\u10_mem_reg[2][28]  <= n2751;
    \\u9_mem_reg[1][23]  <= n2756;
    \\u9_mem_reg[1][24]  <= n2761;
    \\u9_mem_reg[1][26]  <= n2766;
    \\u10_mem_reg[2][29]  <= n2771;
    \\u9_mem_reg[1][27]  <= n2776;
    \\u9_mem_reg[1][29]  <= n2781;
    \\u9_mem_reg[1][30]  <= n2786;
    \\u9_mem_reg[1][31]  <= n2791;
    \\u10_mem_reg[2][30]  <= n2796;
    \\u9_mem_reg[2][18]  <= n2801;
    \\u9_mem_reg[2][19]  <= n2806;
    \\u10_mem_reg[2][31]  <= n2811;
    \\u9_mem_reg[2][21]  <= n2816;
    \\u9_mem_reg[2][22]  <= n2821;
    \\u9_mem_reg[2][23]  <= n2826;
    \\u9_mem_reg[2][25]  <= n2831;
    \\u9_mem_reg[2][26]  <= n2836;
    \\u9_mem_reg[2][27]  <= n2841;
    \\u9_mem_reg[2][29]  <= n2846;
    \\u9_mem_reg[2][30]  <= n2851;
    \\u9_mem_reg[2][31]  <= n2856;
    \\u9_mem_reg[3][18]  <= n2861;
    \\u9_mem_reg[3][19]  <= n2866;
    \\u9_mem_reg[3][20]  <= n2871;
    \\u9_mem_reg[3][21]  <= n2876;
    \\u9_mem_reg[3][23]  <= n2881;
    \\u9_mem_reg[3][24]  <= n2886;
    \\u9_mem_reg[3][25]  <= n2891;
    \\u9_mem_reg[3][27]  <= n2896;
    \\u9_mem_reg[3][28]  <= n2901;
    \\u9_mem_reg[3][29]  <= n2906;
    \\u9_mem_reg[3][31]  <= n2911;
    \\u10_mem_reg[3][18]  <= n2916;
    \\u10_mem_reg[3][19]  <= n2921;
    \\u10_mem_reg[3][20]  <= n2926;
    \\u10_mem_reg[3][21]  <= n2931;
    \\u10_mem_reg[3][22]  <= n2936;
    \\u10_mem_reg[3][23]  <= n2941;
    \\u10_mem_reg[3][25]  <= n2946;
    \\u10_mem_reg[3][26]  <= n2951;
    \\u10_mem_reg[3][27]  <= n2956;
    \\u10_mem_reg[3][29]  <= n2961;
    \\u10_mem_reg[3][30]  <= n2966;
    \\u10_mem_reg[3][31]  <= n2971;
    \\u10_mem_reg[0][19]  <= n2976;
    \\u10_mem_reg[1][18]  <= n2981;
    \\u10_mem_reg[1][19]  <= n2986;
    \\u10_mem_reg[1][21]  <= n2991;
    \\u10_mem_reg[1][22]  <= n2996;
    \\u10_mem_reg[1][23]  <= n3001;
    \\u10_mem_reg[1][24]  <= n3006;
    \\u10_mem_reg[1][25]  <= n3011;
    \\u10_mem_reg[1][26]  <= n3016;
    \\u10_mem_reg[1][27]  <= n3021;
    \\u10_mem_reg[1][28]  <= n3026;
    \\u10_mem_reg[1][29]  <= n3031;
    \\u10_mem_reg[1][20]  <= n3036;
    \\u10_mem_reg[1][30]  <= n3041;
    \\u10_mem_reg[1][31]  <= n3046;
    \\u11_mem_reg[3][8]  <= n3051;
    \\u11_mem_reg[3][9]  <= n3056;
    \\u10_mem_reg[2][1]  <= n3061;
    \\u10_mem_reg[2][5]  <= n3066;
    \\u10_mem_reg[2][6]  <= n3071;
    \\u10_mem_reg[3][3]  <= n3076;
    \\u10_mem_reg[2][9]  <= n3081;
    \\u11_mem_reg[1][0]  <= n3086;
    \\u11_mem_reg[1][10]  <= n3091;
    \\u11_mem_reg[1][11]  <= n3096;
    \\u10_mem_reg[3][2]  <= n3101;
    \\u10_mem_reg[3][9]  <= n3106;
    \\u11_mem_reg[1][14]  <= n3111;
    \\u11_mem_reg[1][1]  <= n3116;
    \\u11_mem_reg[1][2]  <= n3121;
    \\u11_mem_reg[1][3]  <= n3126;
    \\u11_mem_reg[1][4]  <= n3131;
    \\u11_mem_reg[1][5]  <= n3136;
    \\u11_mem_reg[1][7]  <= n3141;
    \\u11_mem_reg[1][8]  <= n3146;
    \\u11_mem_reg[1][9]  <= n3151;
    \\u11_mem_reg[2][0]  <= n3156;
    \\u11_mem_reg[2][10]  <= n3161;
    \\u11_mem_reg[2][11]  <= n3166;
    \\u11_mem_reg[2][13]  <= n3171;
    \\u11_mem_reg[2][14]  <= n3176;
    \\u11_mem_reg[2][15]  <= n3181;
    \\u11_mem_reg[2][16]  <= n3186;
    \\u11_mem_reg[1][17]  <= n3191;
    \\u11_mem_reg[2][12]  <= n3196;
    \\u11_mem_reg[2][2]  <= n3201;
    \\u11_mem_reg[2][3]  <= n3206;
    \\u11_mem_reg[2][6]  <= n3211;
    \\u11_mem_reg[2][4]  <= n3216;
    \\u11_mem_reg[2][5]  <= n3221;
    \\u11_mem_reg[2][9]  <= n3226;
    \\u11_mem_reg[3][11]  <= n3231;
    \\u11_mem_reg[3][12]  <= n3236;
    \\u11_mem_reg[3][15]  <= n3241;
    \\u11_mem_reg[3][10]  <= n3246;
    \\u11_mem_reg[3][2]  <= n3251;
    \\u11_mem_reg[3][3]  <= n3256;
    \\u11_mem_reg[3][4]  <= n3261;
    \\u11_mem_reg[3][1]  <= n3266;
    \\u10_wp_reg[1]  <= n3271;
    \\u10_wp_reg[2]  <= n3276;
    \\u10_mem_reg[0][2]  <= n3281;
    \\u11_mem_reg[0][5]  <= n3286;
    \\u10_mem_reg[0][13]  <= n3291;
    \\u10_mem_reg[0][12]  <= n3296;
    \\u11_mem_reg[0][16]  <= n3301;
    \\u11_mem_reg[0][20]  <= n3306;
    \\u11_mem_reg[0][21]  <= n3311;
    \\u11_mem_reg[0][22]  <= n3316;
    \\u11_mem_reg[0][23]  <= n3321;
    \\u11_mem_reg[0][24]  <= n3326;
    \\u11_mem_reg[0][25]  <= n3331;
    \\u10_mem_reg[0][21]  <= n3336;
    \\u11_mem_reg[0][26]  <= n3341;
    \\u11_mem_reg[0][27]  <= n3346;
    \\u10_mem_reg[0][22]  <= n3351;
    \\u11_mem_reg[0][28]  <= n3356;
    \\u11_mem_reg[0][29]  <= n3361;
    \\u11_mem_reg[0][2]  <= n3366;
    \\u11_mem_reg[0][30]  <= n3371;
    \\u11_mem_reg[0][31]  <= n3376;
    \\u11_mem_reg[0][3]  <= n3381;
    \\u10_mem_reg[0][25]  <= n3386;
    \\u11_mem_reg[0][4]  <= n3391;
    \\u10_mem_reg[0][26]  <= n3396;
    \\u10_mem_reg[0][27]  <= n3401;
    \\u11_mem_reg[0][6]  <= n3406;
    \\u10_mem_reg[0][28]  <= n3411;
    \\u11_mem_reg[0][7]  <= n3416;
    \\u11_mem_reg[0][8]  <= n3421;
    \\u10_mem_reg[0][29]  <= n3426;
    \\u11_mem_reg[0][9]  <= n3431;
    \\u10_mem_reg[0][5]  <= n3436;
    \\u11_wp_reg[0]  <= n3441;
    \\u25_int_set_reg[2]  <= n3446;
    \\u10_mem_reg[0][1]  <= n3451;
    \\u11_mem_reg[0][17]  <= n3456;
    \\u10_mem_reg[3][17]  <= n3461;
    \\u1_sr_reg[15]  <= n3466;
    \\u10_mem_reg[0][11]  <= n3471;
    \\u9_mem_reg[0][4]  <= n3476;
    \\u9_wp_reg[3]  <= n3481;
    \\u9_mem_reg[0][8]  <= n3486;
    \\u10_mem_reg[1][8]  <= n3491;
    \\u9_mem_reg[0][2]  <= n3496;
    \\u9_mem_reg[0][26]  <= n3501;
    \\u10_mem_reg[1][6]  <= n3506;
    \\u9_mem_reg[0][17]  <= n3511;
    \\u9_mem_reg[0][13]  <= n3516;
    \\u10_mem_reg[1][1]  <= n3521;
    \\u10_mem_reg[1][15]  <= n3526;
    \\u10_mem_reg[1][13]  <= n3531;
    \\u10_mem_reg[1][10]  <= n3536;
    \\u10_mem_reg[3][8]  <= n3541;
    \\u10_mem_reg[0][23]  <= n3546;
    \\u11_din_tmp1_reg[8]  <= n3551;
    \\u9_mem_reg[2][12]  <= n3556;
    \\u10_mem_reg[3][13]  <= n3561;
    \\u10_mem_reg[3][0]  <= n3566;
    \\u9_mem_reg[3][4]  <= n3571;
    \\u9_mem_reg[3][1]  <= n3576;
    \\u9_mem_reg[3][15]  <= n3581;
    \\u9_mem_reg[2][5]  <= n3586;
    \\u9_mem_reg[2][2]  <= n3591;
    \\u10_mem_reg[1][9]  <= n3596;
    \\u10_mem_reg[2][0]  <= n3601;
    \\u10_mem_reg[2][11]  <= n3606;
    \\u10_mem_reg[2][12]  <= n3611;
    \\u10_mem_reg[2][13]  <= n3616;
    \\u10_mem_reg[2][14]  <= n3621;
    \\u10_mem_reg[2][15]  <= n3626;
    \\u10_mem_reg[2][16]  <= n3631;
    \\u10_mem_reg[2][10]  <= n3636;
    \\u9_mem_reg[1][0]  <= n3641;
    \\u9_mem_reg[1][10]  <= n3646;
    \\u9_mem_reg[1][12]  <= n3651;
    \\u9_mem_reg[1][13]  <= n3656;
    \\u9_mem_reg[1][14]  <= n3661;
    \\u9_mem_reg[1][16]  <= n3666;
    \\u9_mem_reg[1][17]  <= n3671;
    \\u9_mem_reg[1][1]  <= n3676;
    \\u9_mem_reg[1][2]  <= n3681;
    \\u9_mem_reg[1][3]  <= n3686;
    \\u9_mem_reg[1][4]  <= n3691;
    \\u9_mem_reg[1][5]  <= n3696;
    \\u9_mem_reg[1][6]  <= n3701;
    \\u9_mem_reg[1][7]  <= n3706;
    \\u9_mem_reg[1][8]  <= n3711;
    \\u9_mem_reg[2][0]  <= n3716;
    \\u9_mem_reg[2][10]  <= n3721;
    \\u9_mem_reg[2][11]  <= n3726;
    \\u9_mem_reg[2][14]  <= n3731;
    \\u9_mem_reg[2][15]  <= n3736;
    \\u9_mem_reg[2][16]  <= n3741;
    \\u9_mem_reg[2][17]  <= n3746;
    \\u9_mem_reg[2][1]  <= n3751;
    \\u10_mem_reg[2][3]  <= n3756;
    \\u9_mem_reg[2][3]  <= n3761;
    \\u10_mem_reg[2][4]  <= n3766;
    \\u9_mem_reg[2][4]  <= n3771;
    \\u9_mem_reg[2][6]  <= n3776;
    \\u9_mem_reg[2][7]  <= n3781;
    \\u9_mem_reg[2][8]  <= n3786;
    \\u9_mem_reg[3][0]  <= n3791;
    \\u9_mem_reg[3][10]  <= n3796;
    \\u9_mem_reg[3][11]  <= n3801;
    \\u9_mem_reg[3][12]  <= n3806;
    \\u9_mem_reg[3][13]  <= n3811;
    \\u9_mem_reg[3][14]  <= n3816;
    \\u9_mem_reg[2][13]  <= n3821;
    \\u9_mem_reg[3][16]  <= n3826;
    \\u9_mem_reg[3][17]  <= n3831;
    \\u10_mem_reg[2][7]  <= n3836;
    \\u9_mem_reg[3][2]  <= n3841;
    \\u9_mem_reg[3][3]  <= n3846;
    \\u9_mem_reg[3][5]  <= n3851;
    \\u9_mem_reg[3][6]  <= n3856;
    \\u9_mem_reg[3][7]  <= n3861;
    \\u10_mem_reg[2][8]  <= n3866;
    \\u9_mem_reg[3][9]  <= n3871;
    \\u9_mem_reg[3][8]  <= n3876;
    \\u10_mem_reg[3][10]  <= n3881;
    \\u10_mem_reg[3][11]  <= n3886;
    \\u10_mem_reg[3][12]  <= n3891;
    \\u10_mem_reg[3][14]  <= n3896;
    \\u10_mem_reg[3][15]  <= n3901;
    \\u10_mem_reg[3][16]  <= n3906;
    \\u10_mem_reg[3][1]  <= n3911;
    \\u10_mem_reg[3][4]  <= n3916;
    \\u10_mem_reg[3][5]  <= n3921;
    \\u10_mem_reg[3][6]  <= n3926;
    \\u10_mem_reg[3][7]  <= n3931;
    \\u10_mem_reg[1][11]  <= n3936;
    \\u10_mem_reg[1][12]  <= n3941;
    \\u10_mem_reg[1][14]  <= n3946;
    \\u10_mem_reg[1][17]  <= n3951;
    \\u10_mem_reg[1][16]  <= n3956;
    \\u9_mem_reg[1][9]  <= n3961;
    \\u10_mem_reg[1][3]  <= n3966;
    \\u10_mem_reg[1][4]  <= n3971;
    \\u10_mem_reg[1][5]  <= n3976;
    \\u10_mem_reg[1][2]  <= n3981;
    \\u10_mem_reg[2][2]  <= n3986;
    \\u10_mem_reg[1][7]  <= n3991;
    \\u9_wp_reg[2]  <= n3996;
    \\u9_mem_reg[1][15]  <= n4001;
    \\u9_mem_reg[1][11]  <= n4006;
    \\u10_mem_reg[2][17]  <= n4011;
    \\u10_mem_reg[0][24]  <= n4016;
    \\u11_din_tmp1_reg[4]  <= n4021;
    \\u10_mem_reg[0][8]  <= n4026;
    \\u10_mem_reg[0][4]  <= n4031;
    \\u9_mem_reg[0][0]  <= n4036;
    \\u9_mem_reg[0][10]  <= n4041;
    \\u9_mem_reg[0][11]  <= n4046;
    \\u9_mem_reg[0][12]  <= n4051;
    \\u9_mem_reg[0][14]  <= n4056;
    \\u9_mem_reg[0][15]  <= n4061;
    \\u9_mem_reg[0][16]  <= n4066;
    \\u9_mem_reg[0][1]  <= n4071;
    \\u9_mem_reg[0][20]  <= n4076;
    \\u9_mem_reg[0][21]  <= n4081;
    \\u9_mem_reg[0][22]  <= n4086;
    \\u9_mem_reg[0][23]  <= n4091;
    \\u9_mem_reg[0][24]  <= n4096;
    \\u9_mem_reg[0][25]  <= n4101;
    \\u9_mem_reg[0][27]  <= n4106;
    \\u9_mem_reg[0][28]  <= n4111;
    \\u9_mem_reg[0][29]  <= n4116;
    \\u9_mem_reg[0][30]  <= n4121;
    \\u9_mem_reg[0][31]  <= n4126;
    \\u9_mem_reg[0][3]  <= n4131;
    \\u9_mem_reg[0][5]  <= n4136;
    \\u9_mem_reg[0][6]  <= n4141;
    \\u9_mem_reg[0][7]  <= n4146;
    \\u9_mem_reg[0][9]  <= n4151;
    \\u10_mem_reg[0][0]  <= n4156;
    \\u10_mem_reg[0][10]  <= n4161;
    \\u10_mem_reg[0][14]  <= n4166;
    \\u10_mem_reg[0][15]  <= n4171;
    \\u10_mem_reg[0][16]  <= n4176;
    \\u10_mem_reg[0][17]  <= n4181;
    \\u10_mem_reg[0][31]  <= n4186;
    \\u10_mem_reg[0][3]  <= n4191;
    \\u10_mem_reg[0][30]  <= n4196;
    \\u10_mem_reg[0][6]  <= n4201;
    \\u10_mem_reg[0][7]  <= n4206;
    \\u10_mem_reg[0][9]  <= n4211;
    \\u10_wp_reg[0]  <= n4216;
    \\u11_din_tmp1_reg[0]  <= n4221;
    \\u11_din_tmp1_reg[10]  <= n4226;
    \\u11_din_tmp1_reg[11]  <= n4231;
    \\u11_din_tmp1_reg[12]  <= n4236;
    \\u11_din_tmp1_reg[13]  <= n4241;
    \\u11_din_tmp1_reg[14]  <= n4246;
    \\u11_din_tmp1_reg[15]  <= n4251;
    \\u11_din_tmp1_reg[1]  <= n4256;
    \\u11_din_tmp1_reg[2]  <= n4261;
    \\u11_din_tmp1_reg[3]  <= n4266;
    \\u11_din_tmp1_reg[5]  <= n4271;
    \\u11_din_tmp1_reg[6]  <= n4276;
    \\u11_din_tmp1_reg[7]  <= n4281;
    \\u11_din_tmp1_reg[9]  <= n4286;
    \\u9_mem_reg[2][9]  <= n4291;
    \\u18_int_set_reg[1]  <= n4296;
    \\u19_int_set_reg[1]  <= n4301;
    \\u24_int_set_reg[2]  <= n4306;
    u15_crac_wr_reg <= n4311;
    \\u13_ints_r_reg[1]  <= n4316;
    \\u10_mem_reg[0][20]  <= n4321;
    \\u0_slt9_r_reg[3]  <= n4326;
    \\u10_din_tmp1_reg[13]  <= n4331;
    \\u1_slt6_reg[12]  <= n4336;
    \\u13_ints_r_reg[26]  <= n4341;
    \\u1_slt0_reg[12]  <= n4346;
    \\u1_slt2_reg[12]  <= n4351;
    \\u1_slt3_reg[12]  <= n4356;
    \\u1_slt4_reg[12]  <= n4361;
    \\u10_din_tmp1_reg[11]  <= n4366;
    \\u9_wp_reg[0]  <= n4371;
    \\u10_din_tmp1_reg[5]  <= n4376;
    \\u10_din_tmp1_reg[3]  <= n4381;
    \\u10_din_tmp1_reg[1]  <= n4386;
    \\u10_din_tmp1_reg[2]  <= n4391;
    \\u10_din_tmp1_reg[4]  <= n4396;
    \\u10_din_tmp1_reg[6]  <= n4401;
    \\u10_din_tmp1_reg[8]  <= n4406;
    \\u10_din_tmp1_reg[9]  <= n4411;
    \\u10_din_tmp1_reg[7]  <= n4416;
    \\u10_din_tmp1_reg[0]  <= n4421;
    \\u10_din_tmp1_reg[10]  <= n4426;
    \\u10_din_tmp1_reg[15]  <= n4431;
    \\u10_din_tmp1_reg[14]  <= n4436;
    \\u10_din_tmp1_reg[12]  <= n4441;
    u15_rdd1_reg <= n4446;
    u15_rdd2_reg <= n4451;
    \\u20_int_set_reg[0]  <= n4456;
    \\u18_int_set_reg[0]  <= n4461;
    \\u1_sr_reg[14]  <= n4466;
    \\u13_ints_r_reg[23]  <= n4471;
    \\u13_ints_r_reg[20]  <= n4476;
    \\u9_wp_reg[1]  <= n4481;
    \\u9_din_tmp1_reg[9]  <= n4486;
    \\u9_din_tmp1_reg[3]  <= n4491;
    \\u9_din_tmp1_reg[10]  <= n4496;
    \\u9_din_tmp1_reg[14]  <= n4501;
    \\u9_din_tmp1_reg[0]  <= n4506;
    \\u9_din_tmp1_reg[11]  <= n4511;
    \\u9_din_tmp1_reg[12]  <= n4516;
    \\u9_din_tmp1_reg[13]  <= n4521;
    \\u9_din_tmp1_reg[15]  <= n4526;
    \\u9_din_tmp1_reg[1]  <= n4531;
    \\u9_din_tmp1_reg[2]  <= n4536;
    \\u9_din_tmp1_reg[5]  <= n4541;
    \\u9_din_tmp1_reg[6]  <= n4546;
    \\u9_din_tmp1_reg[4]  <= n4551;
    \\u9_din_tmp1_reg[8]  <= n4556;
    \\u9_din_tmp1_reg[7]  <= n4561;
    u15_rdd3_reg <= n4566;
    \\u21_int_set_reg[0]  <= n4571;
    \\u22_int_set_reg[0]  <= n4576;
    \\u17_int_set_reg[0]  <= n4581;
    \\u19_int_set_reg[0]  <= n4586;
    u16_u8_dma_req_r1_reg <= n4591;
    \\u1_slt4_reg[11]  <= n4596;
    \\u1_slt0_reg[11]  <= n4601;
    \\u1_slt1_reg[11]  <= n4606;
    \\u1_slt2_reg[11]  <= n4611;
    \\u1_slt3_reg[11]  <= n4616;
    \\u1_slt6_reg[11]  <= n4621;
    \\u23_int_set_reg[2]  <= n4626;
    u15_crac_rd_done_reg <= n4631;
    u16_u6_dma_req_r1_reg <= n4636;
    u16_u7_dma_req_r1_reg <= n4641;
    \\u1_sr_reg[13]  <= n4646;
    \\u1_slt6_reg[10]  <= n4651;
    \\u1_slt2_reg[10]  <= n4656;
    u14_u4_en_out_l_reg <= n4661;
    u2_sync_resume_reg <= n4666;
    \\u1_slt1_reg[10]  <= n4671;
    \\u1_slt4_reg[10]  <= n4676;
    \\u1_slt3_reg[10]  <= n4681;
    u14_u0_en_out_l_reg <= n4686;
    u14_u1_en_out_l_reg <= n4691;
    u14_u2_en_out_l_reg <= n4696;
    u14_u3_en_out_l_reg <= n4701;
    u14_u5_en_out_l_reg <= n4706;
    u14_crac_valid_r_reg <= n4711;
    \\u0_slt9_r_reg[2]  <= n4716;
    \\u1_sr_reg[12]  <= n4721;
    \\u26_ps_cnt_reg[5]  <= n4726;
    \\u26_ps_cnt_reg[2]  <= n4731;
    \\u26_ps_cnt_reg[0]  <= n4736;
    \\u26_ps_cnt_reg[1]  <= n4741;
    \\u26_ps_cnt_reg[4]  <= n4746;
    \\u26_ps_cnt_reg[3]  <= n4751;
    \\u12_wb_data_o_reg[1]  <= n4756;
    \\u17_int_set_reg[2]  <= n4761;
    \\u18_int_set_reg[2]  <= n4766;
    \\u21_int_set_reg[2]  <= n4771;
    \\u20_int_set_reg[2]  <= n4776;
    u14_crac_wr_r_reg <= n4781;
    \\u22_int_set_reg[2]  <= n4786;
    \\u19_int_set_reg[2]  <= n4791;
    \\u1_slt2_reg[9]  <= n4796;
    u14_u3_full_empty_r_reg <= n4801;
    \\u25_int_set_reg[0]  <= n4806;
    u14_u0_full_empty_r_reg <= n4811;
    u14_u1_full_empty_r_reg <= n4816;
    u14_u2_full_empty_r_reg <= n4821;
    u14_u5_full_empty_r_reg <= n4826;
    \\u1_slt0_reg[9]  <= n4831;
    u14_u4_full_empty_r_reg <= n4836;
    \\u1_slt4_reg[9]  <= n4841;
    \\u1_slt3_reg[9]  <= n4846;
    \\u8_wp_reg[0]  <= n4851;
    \\u3_wp_reg[0]  <= n4856;
    \\u4_wp_reg[0]  <= n4861;
    \\u5_wp_reg[0]  <= n4866;
    \\u6_wp_reg[0]  <= n4871;
    \\u7_wp_reg[0]  <= n4876;
    \\u1_slt6_reg[9]  <= n4881;
    u26_ac97_rst__reg <= n4886;
    \\u1_sr_reg[11]  <= n4891;
    \\u26_cnt_reg[2]  <= n4896;
    \\u23_int_set_reg[0]  <= n4901;
    \\u24_int_set_reg[0]  <= n4906;
    u14_u8_en_out_l_reg <= n4911;
    \\u5_wp_reg[1]  <= n4916;
    \\u6_wp_reg[2]  <= n4921;
    \\u26_cnt_reg[0]  <= n4926;
    \\u26_cnt_reg[1]  <= n4931;
    \\u8_wp_reg[2]  <= n4936;
    \\u3_wp_reg[2]  <= n4941;
    \\u5_wp_reg[2]  <= n4946;
    \\u7_wp_reg[2]  <= n4951;
    u14_u6_en_out_l_reg <= n4956;
    u14_u7_en_out_l_reg <= n4961;
    \\u8_wp_reg[1]  <= n4966;
    \\u3_wp_reg[1]  <= n4971;
    \\u4_wp_reg[1]  <= n4976;
    \\u6_wp_reg[1]  <= n4981;
    \\u7_wp_reg[1]  <= n4986;
    \\u4_wp_reg[2]  <= n4991;
    u15_valid_r_reg <= n4996;
    \\u1_slt6_reg[8]  <= n5001;
    \\u1_slt2_reg[8]  <= n5006;
    \\u1_slt1_reg[8]  <= n5011;
    \\u1_slt4_reg[8]  <= n5016;
    \\u1_slt3_reg[8]  <= n5021;
    \\u4_mem_reg[0][13]  <= n5026;
    \\u4_mem_reg[0][14]  <= n5031;
    \\u4_mem_reg[0][16]  <= n5036;
    \\u4_mem_reg[0][19]  <= n5041;
    \\u4_mem_reg[0][22]  <= n5046;
    \\u4_mem_reg[0][24]  <= n5051;
    \\u4_mem_reg[0][31]  <= n5056;
    \\u4_mem_reg[0][4]  <= n5061;
    \\u4_mem_reg[0][7]  <= n5066;
    \\u4_mem_reg[0][9]  <= n5071;
    \\u5_mem_reg[0][13]  <= n5076;
    \\u5_mem_reg[0][14]  <= n5081;
    \\u5_mem_reg[0][16]  <= n5086;
    \\u5_mem_reg[0][19]  <= n5091;
    \\u5_mem_reg[0][22]  <= n5096;
    \\u5_mem_reg[0][24]  <= n5101;
    \\u5_mem_reg[0][31]  <= n5106;
    \\u5_mem_reg[0][4]  <= n5111;
    \\u5_mem_reg[0][7]  <= n5116;
    \\u5_mem_reg[0][9]  <= n5121;
    \\u6_mem_reg[0][13]  <= n5126;
    \\u6_mem_reg[0][14]  <= n5131;
    \\u6_mem_reg[0][16]  <= n5136;
    \\u6_mem_reg[0][19]  <= n5141;
    \\u6_mem_reg[0][22]  <= n5146;
    \\u6_mem_reg[0][24]  <= n5151;
    \\u6_mem_reg[0][31]  <= n5156;
    \\u6_mem_reg[0][4]  <= n5161;
    \\u6_mem_reg[0][7]  <= n5166;
    \\u6_mem_reg[0][9]  <= n5171;
    \\u7_mem_reg[0][13]  <= n5176;
    \\u7_mem_reg[0][14]  <= n5181;
    \\u7_mem_reg[0][16]  <= n5186;
    \\u7_mem_reg[0][19]  <= n5191;
    \\u7_mem_reg[0][22]  <= n5196;
    \\u7_mem_reg[0][24]  <= n5201;
    \\u7_mem_reg[0][31]  <= n5206;
    \\u7_mem_reg[0][4]  <= n5211;
    \\u7_mem_reg[0][7]  <= n5216;
    \\u7_mem_reg[0][9]  <= n5221;
    \\u3_mem_reg[0][11]  <= n5226;
    \\u3_mem_reg[0][12]  <= n5231;
    \\u3_mem_reg[0][15]  <= n5236;
    \\u8_mem_reg[0][0]  <= n5241;
    \\u8_mem_reg[0][11]  <= n5246;
    \\u8_mem_reg[0][12]  <= n5251;
    \\u8_mem_reg[0][17]  <= n5256;
    \\u3_mem_reg[0][1]  <= n5261;
    \\u3_mem_reg[0][21]  <= n5266;
    \\u8_mem_reg[0][26]  <= n5271;
    \\u8_mem_reg[0][28]  <= n5276;
    \\u8_mem_reg[0][29]  <= n5281;
    \\u8_mem_reg[0][30]  <= n5286;
    \\u3_mem_reg[0][27]  <= n5291;
    \\u8_mem_reg[0][4]  <= n5296;
    \\u8_mem_reg[0][5]  <= n5301;
    \\u3_mem_reg[0][2]  <= n5306;
    \\u3_mem_reg[0][29]  <= n5311;
    \\u3_mem_reg[0][6]  <= n5316;
    \\u3_mem_reg[0][5]  <= n5321;
    \\u13_crac_r_reg[6]  <= n5326;
    \\u3_mem_reg[0][17]  <= n5331;
    \\u8_mem_reg[2][18]  <= n5336;
    \\u7_mem_reg[0][20]  <= n5341;
    \\u8_mem_reg[2][25]  <= n5346;
    \\u8_mem_reg[2][28]  <= n5351;
    \\u4_mem_reg[2][16]  <= n5356;
    \\u5_mem_reg[1][26]  <= n5361;
    \\u13_occ0_r_reg[11]  <= n5366;
    \\u5_mem_reg[1][22]  <= n5371;
    \\u5_mem_reg[1][15]  <= n5376;
    \\u5_mem_reg[1][19]  <= n5381;
    \\u5_mem_reg[1][11]  <= n5386;
    \\u3_mem_reg[1][22]  <= n5391;
    \\u8_mem_reg[2][20]  <= n5396;
    \\u4_mem_reg[3][9]  <= n5401;
    \\u4_mem_reg[3][5]  <= n5406;
    \\u4_mem_reg[3][30]  <= n5411;
    \\u8_mem_reg[0][15]  <= n5416;
    \\u3_mem_reg[0][16]  <= n5421;
    \\u4_mem_reg[3][23]  <= n5426;
    \\u4_mem_reg[3][27]  <= n5431;
    \\u8_mem_reg[1][6]  <= n5436;
    \\u13_occ0_r_reg[8]  <= n5441;
    \\u13_icc_r_reg[8]  <= n5446;
    \\u8_mem_reg[2][13]  <= n5451;
    \\u3_mem_reg[1][19]  <= n5456;
    \\u4_mem_reg[2][9]  <= n5461;
    \\u4_mem_reg[3][16]  <= n5466;
    \\u4_mem_reg[3][12]  <= n5471;
    \\u4_mem_reg[2][5]  <= n5476;
    \\u3_mem_reg[1][15]  <= n5481;
    \\u4_mem_reg[2][30]  <= n5486;
    \\u4_mem_reg[2][27]  <= n5491;
    \\u4_mem_reg[2][23]  <= n5496;
    \\u7_mem_reg[0][30]  <= n5501;
    \\u3_mem_reg[2][2]  <= n5506;
    \\u8_mem_reg[1][21]  <= n5511;
    \\u3_mem_reg[1][11]  <= n5516;
    \\u8_mem_reg[1][3]  <= n5521;
    \\u4_mem_reg[2][12]  <= n5526;
    \\u4_mem_reg[1][30]  <= n5531;
    \\u4_mem_reg[1][9]  <= n5536;
    \\u4_mem_reg[1][5]  <= n5541;
    \\u4_mem_reg[1][27]  <= n5546;
    \\u8_mem_reg[1][28]  <= n5551;
    \\u3_mem_reg[0][13]  <= n5556;
    \\u8_mem_reg[1][25]  <= n5561;
    \\u4_mem_reg[1][23]  <= n5566;
    \\u4_mem_reg[1][16]  <= n5571;
    \\u7_mem_reg[0][6]  <= n5576;
    \\u7_mem_reg[1][25]  <= n5581;
    \\u3_mem_reg[3][3]  <= n5586;
    \\u4_mem_reg[1][12]  <= n5591;
    \\u7_mem_reg[3][3]  <= n5596;
    \\u8_mem_reg[1][14]  <= n5601;
    \\u8_mem_reg[1][18]  <= n5606;
    \\u3_mem_reg[3][6]  <= n5611;
    \\u3_mem_reg[3][22]  <= n5616;
    \\u3_mem_reg[3][30]  <= n5621;
    \\u3_mem_reg[3][27]  <= n5626;
    \\u7_mem_reg[0][23]  <= n5631;
    \\u3_mem_reg[3][19]  <= n5636;
    u14_u0_en_out_l2_reg <= n5641;
    u14_u1_en_out_l2_reg <= n5646;
    u14_u2_en_out_l2_reg <= n5651;
    u14_u3_en_out_l2_reg <= n5656;
    u14_u4_en_out_l2_reg <= n5661;
    u14_u5_en_out_l2_reg <= n5666;
    \\u6_mem_reg[0][12]  <= n5671;
    \\u8_mem_reg[1][10]  <= n5676;
    \\u7_mem_reg[3][7]  <= n5681;
    \\u3_mem_reg[3][15]  <= n5686;
    \\u3_mem_reg[3][11]  <= n5691;
    \\u3_mem_reg[2][8]  <= n5696;
    \\u7_mem_reg[0][12]  <= n5701;
    \\u7_mem_reg[3][14]  <= n5706;
    \\u7_mem_reg[3][25]  <= n5711;
    \\u7_mem_reg[3][29]  <= n5716;
    \\u3_mem_reg[2][26]  <= n5721;
    \\u3_mem_reg[2][22]  <= n5726;
    \\u3_mem_reg[2][18]  <= n5731;
    \\u8_mem_reg[3][8]  <= n5736;
    \\u8_mem_reg[3][6]  <= n5741;
    \\u7_mem_reg[3][21]  <= n5746;
    \\u7_mem_reg[3][18]  <= n5751;
    \\u8_mem_reg[3][3]  <= n5756;
    \\u3_mem_reg[2][11]  <= n5761;
    \\u8_mem_reg[3][28]  <= n5766;
    \\u7_mem_reg[0][17]  <= n5771;
    \\u7_mem_reg[0][0]  <= n5776;
    \\u8_mem_reg[3][22]  <= n5781;
    \\u8_mem_reg[3][25]  <= n5786;
    \\u7_mem_reg[2][25]  <= n5791;
    \\u7_mem_reg[2][7]  <= n5796;
    \\u7_mem_reg[3][10]  <= n5801;
    \\u8_mem_reg[3][18]  <= n5806;
    \\u3_mem_reg[1][3]  <= n5811;
    \\u8_mem_reg[3][15]  <= n5816;
    \\u8_mem_reg[3][10]  <= n5821;
    \\u7_mem_reg[2][3]  <= n5826;
    \\u7_mem_reg[2][29]  <= n5831;
    \\u3_mem_reg[1][2]  <= n5836;
    \\u7_mem_reg[2][21]  <= n5841;
    \\u7_mem_reg[2][18]  <= n5846;
    \\u6_mem_reg[0][30]  <= n5851;
    \\u6_mem_reg[0][6]  <= n5856;
    \\u7_mem_reg[2][14]  <= n5861;
    \\u7_mem_reg[2][10]  <= n5866;
    \\u8_mem_reg[2][6]  <= n5871;
    \\u6_mem_reg[0][28]  <= n5876;
    \\u7_mem_reg[1][7]  <= n5881;
    \\u6_mem_reg[3][8]  <= n5886;
    \\u13_crac_dout_r_reg[3]  <= n5891;
    \\u13_crac_dout_r_reg[9]  <= n5896;
    \\u7_mem_reg[1][3]  <= n5901;
    \\u13_icc_r_reg[22]  <= n5906;
    \\u13_crac_dout_r_reg[14]  <= n5911;
    \\u13_occ0_r_reg[2]  <= n5916;
    \\u13_occ0_r_reg[4]  <= n5921;
    \\u13_intm_r_reg[7]  <= n5926;
    \\u13_intm_r_reg[22]  <= n5931;
    \\u13_icc_r_reg[11]  <= n5936;
    \\u7_mem_reg[1][29]  <= n5941;
    \\u6_mem_reg[0][23]  <= n5946;
    \\u13_icc_r_reg[15]  <= n5951;
    \\u13_icc_r_reg[19]  <= n5956;
    \\u13_crac_r_reg[0]  <= n5961;
    \\u13_crac_r_reg[1]  <= n5966;
    \\u13_crac_r_reg[3]  <= n5971;
    \\u13_crac_r_reg[4]  <= n5976;
    \\u13_crac_r_reg[5]  <= n5981;
    \\u13_crac_r_reg[7]  <= n5986;
    \\u13_icc_r_reg[0]  <= n5991;
    \\u13_icc_r_reg[10]  <= n5996;
    \\u13_icc_r_reg[12]  <= n6001;
    \\u13_icc_r_reg[13]  <= n6006;
    \\u13_icc_r_reg[14]  <= n6011;
    \\u13_icc_r_reg[16]  <= n6016;
    \\u13_icc_r_reg[17]  <= n6021;
    \\u13_icc_r_reg[18]  <= n6026;
    \\u13_icc_r_reg[1]  <= n6031;
    \\u13_icc_r_reg[20]  <= n6036;
    \\u13_icc_r_reg[21]  <= n6041;
    \\u13_icc_r_reg[23]  <= n6046;
    \\u13_icc_r_reg[2]  <= n6051;
    \\u13_icc_r_reg[3]  <= n6056;
    \\u13_icc_r_reg[4]  <= n6061;
    \\u13_icc_r_reg[5]  <= n6066;
    \\u13_icc_r_reg[6]  <= n6071;
    \\u13_icc_r_reg[7]  <= n6076;
    \\u13_icc_r_reg[9]  <= n6081;
    \\u13_occ0_r_reg[0]  <= n6086;
    \\u13_occ0_r_reg[10]  <= n6091;
    \\u13_occ0_r_reg[12]  <= n6096;
    \\u13_occ0_r_reg[13]  <= n6101;
    \\u13_occ0_r_reg[14]  <= n6106;
    \\u13_occ0_r_reg[16]  <= n6111;
    \\u13_occ0_r_reg[17]  <= n6116;
    \\u13_occ0_r_reg[18]  <= n6121;
    \\u13_occ0_r_reg[1]  <= n6126;
    \\u13_occ0_r_reg[20]  <= n6131;
    \\u13_occ0_r_reg[21]  <= n6136;
    \\u13_occ0_r_reg[23]  <= n6141;
    \\u13_occ0_r_reg[24]  <= n6146;
    \\u13_occ0_r_reg[25]  <= n6151;
    \\u13_occ0_r_reg[27]  <= n6156;
    \\u13_occ0_r_reg[28]  <= n6161;
    \\u13_occ0_r_reg[29]  <= n6166;
    \\u13_occ0_r_reg[30]  <= n6171;
    \\u13_occ0_r_reg[31]  <= n6176;
    \\u13_occ0_r_reg[3]  <= n6181;
    \\u13_occ0_r_reg[5]  <= n6186;
    \\u13_occ0_r_reg[6]  <= n6191;
    \\u13_occ0_r_reg[7]  <= n6196;
    \\u13_occ0_r_reg[9]  <= n6201;
    \\u13_intm_r_reg[0]  <= n6206;
    \\u13_intm_r_reg[10]  <= n6211;
    \\u13_intm_r_reg[11]  <= n6216;
    \\u13_intm_r_reg[12]  <= n6221;
    \\u13_intm_r_reg[13]  <= n6226;
    \\u13_intm_r_reg[14]  <= n6231;
    \\u13_intm_r_reg[16]  <= n6236;
    \\u13_intm_r_reg[17]  <= n6241;
    \\u13_intm_r_reg[18]  <= n6246;
    \\u13_intm_r_reg[19]  <= n6251;
    \\u13_intm_r_reg[1]  <= n6256;
    \\u13_intm_r_reg[20]  <= n6261;
    \\u13_intm_r_reg[21]  <= n6266;
    \\u13_intm_r_reg[23]  <= n6271;
    \\u13_intm_r_reg[24]  <= n6276;
    \\u13_intm_r_reg[25]  <= n6281;
    \\u13_intm_r_reg[27]  <= n6286;
    \\u13_intm_r_reg[28]  <= n6291;
    \\u13_intm_r_reg[2]  <= n6296;
    \\u13_intm_r_reg[5]  <= n6301;
    \\u13_intm_r_reg[6]  <= n6306;
    \\u13_intm_r_reg[9]  <= n6311;
    \\u13_intm_r_reg[4]  <= n6316;
    \\u13_intm_r_reg[15]  <= n6321;
    \\u13_crac_dout_r_reg[0]  <= n6326;
    \\u13_crac_dout_r_reg[10]  <= n6331;
    \\u13_crac_dout_r_reg[11]  <= n6336;
    \\u13_crac_dout_r_reg[12]  <= n6341;
    \\u13_crac_dout_r_reg[13]  <= n6346;
    \\u13_crac_dout_r_reg[15]  <= n6351;
    \\u13_crac_dout_r_reg[1]  <= n6356;
    \\u13_crac_dout_r_reg[2]  <= n6361;
    \\u13_crac_dout_r_reg[4]  <= n6366;
    \\u13_crac_dout_r_reg[5]  <= n6371;
    \\u13_crac_dout_r_reg[6]  <= n6376;
    \\u13_crac_dout_r_reg[8]  <= n6381;
    \\u8_mem_reg[2][4]  <= n6386;
    \\u3_mem_reg[1][28]  <= n6391;
    \\u8_mem_reg[2][5]  <= n6396;
    \\u3_mem_reg[1][29]  <= n6401;
    \\u8_mem_reg[2][7]  <= n6406;
    \\u8_mem_reg[2][8]  <= n6411;
    \\u8_mem_reg[2][9]  <= n6416;
    \\u8_mem_reg[3][0]  <= n6421;
    \\u3_mem_reg[1][30]  <= n6426;
    \\u8_mem_reg[3][11]  <= n6431;
    \\u3_mem_reg[1][31]  <= n6436;
    \\u8_mem_reg[3][12]  <= n6441;
    \\u8_mem_reg[3][13]  <= n6446;
    \\u3_mem_reg[1][4]  <= n6451;
    \\u8_mem_reg[3][14]  <= n6456;
    \\u8_mem_reg[3][16]  <= n6461;
    \\u8_mem_reg[3][17]  <= n6466;
    \\u3_mem_reg[1][5]  <= n6471;
    \\u8_mem_reg[3][19]  <= n6476;
    \\u3_mem_reg[1][6]  <= n6481;
    \\u8_mem_reg[3][1]  <= n6486;
    \\u3_mem_reg[1][7]  <= n6491;
    \\u8_mem_reg[3][20]  <= n6496;
    \\u8_mem_reg[3][21]  <= n6501;
    \\u3_mem_reg[1][8]  <= n6506;
    \\u8_mem_reg[3][23]  <= n6511;
    \\u8_mem_reg[3][24]  <= n6516;
    \\u3_mem_reg[1][9]  <= n6521;
    \\u8_mem_reg[3][26]  <= n6526;
    \\u3_mem_reg[2][0]  <= n6531;
    \\u8_mem_reg[3][27]  <= n6536;
    \\u3_mem_reg[2][10]  <= n6541;
    \\u8_mem_reg[3][29]  <= n6546;
    \\u8_mem_reg[3][2]  <= n6551;
    \\u8_mem_reg[3][30]  <= n6556;
    \\u8_mem_reg[3][31]  <= n6561;
    \\u3_mem_reg[2][12]  <= n6566;
    \\u8_mem_reg[3][4]  <= n6571;
    \\u3_mem_reg[2][13]  <= n6576;
    \\u8_mem_reg[3][5]  <= n6581;
    \\u3_mem_reg[2][14]  <= n6586;
    \\u8_mem_reg[3][7]  <= n6591;
    \\u3_mem_reg[2][15]  <= n6596;
    \\u8_mem_reg[3][9]  <= n6601;
    \\u3_mem_reg[2][16]  <= n6606;
    \\u3_mem_reg[2][17]  <= n6611;
    \\u3_mem_reg[2][19]  <= n6616;
    \\u3_mem_reg[2][1]  <= n6621;
    \\u3_mem_reg[2][21]  <= n6626;
    \\u3_mem_reg[2][23]  <= n6631;
    \\u3_mem_reg[2][24]  <= n6636;
    \\u3_mem_reg[2][25]  <= n6641;
    \\u3_mem_reg[2][27]  <= n6646;
    \\u3_mem_reg[2][28]  <= n6651;
    \\u3_mem_reg[2][29]  <= n6656;
    \\u3_mem_reg[2][30]  <= n6661;
    \\u3_mem_reg[2][31]  <= n6666;
    \\u3_mem_reg[2][3]  <= n6671;
    \\u3_mem_reg[2][4]  <= n6676;
    \\u3_mem_reg[2][5]  <= n6681;
    \\u3_mem_reg[2][6]  <= n6686;
    \\u3_mem_reg[2][7]  <= n6691;
    \\u3_mem_reg[2][9]  <= n6696;
    \\u3_mem_reg[3][0]  <= n6701;
    \\u3_mem_reg[3][10]  <= n6706;
    \\u3_mem_reg[3][12]  <= n6711;
    \\u3_mem_reg[3][13]  <= n6716;
    \\u3_mem_reg[3][14]  <= n6721;
    \\u3_mem_reg[3][16]  <= n6726;
    \\u3_mem_reg[3][17]  <= n6731;
    \\u3_mem_reg[3][18]  <= n6736;
    \\u3_mem_reg[3][1]  <= n6741;
    \\u3_mem_reg[3][20]  <= n6746;
    \\u3_mem_reg[3][21]  <= n6751;
    \\u3_mem_reg[3][23]  <= n6756;
    \\u3_mem_reg[3][24]  <= n6761;
    \\u3_mem_reg[3][26]  <= n6766;
    \\u3_mem_reg[3][28]  <= n6771;
    \\u3_mem_reg[3][29]  <= n6776;
    \\u3_mem_reg[3][2]  <= n6781;
    \\u3_mem_reg[3][31]  <= n6786;
    \\u3_mem_reg[3][4]  <= n6791;
    \\u3_mem_reg[3][5]  <= n6796;
    \\u3_mem_reg[3][7]  <= n6801;
    \\u3_mem_reg[3][9]  <= n6806;
    \\u3_mem_reg[3][25]  <= n6811;
    \\u4_mem_reg[1][0]  <= n6816;
    \\u4_mem_reg[1][10]  <= n6821;
    \\u4_mem_reg[1][11]  <= n6826;
    \\u4_mem_reg[1][13]  <= n6831;
    \\u4_mem_reg[1][14]  <= n6836;
    \\u4_mem_reg[1][15]  <= n6841;
    \\u4_mem_reg[1][17]  <= n6846;
    \\u4_mem_reg[1][18]  <= n6851;
    \\u4_mem_reg[1][19]  <= n6856;
    \\u4_mem_reg[1][1]  <= n6861;
    \\u4_mem_reg[1][20]  <= n6866;
    \\u4_mem_reg[1][21]  <= n6871;
    \\u4_mem_reg[1][22]  <= n6876;
    \\u4_mem_reg[1][24]  <= n6881;
    \\u4_mem_reg[1][25]  <= n6886;
    \\u4_mem_reg[1][26]  <= n6891;
    \\u4_mem_reg[1][28]  <= n6896;
    \\u4_mem_reg[1][29]  <= n6901;
    \\u4_mem_reg[1][2]  <= n6906;
    \\u4_mem_reg[1][31]  <= n6911;
    \\u4_mem_reg[1][3]  <= n6916;
    \\u4_mem_reg[1][4]  <= n6921;
    \\u4_mem_reg[1][6]  <= n6926;
    \\u4_mem_reg[1][7]  <= n6931;
    \\u4_mem_reg[1][8]  <= n6936;
    \\u4_mem_reg[2][0]  <= n6941;
    \\u4_mem_reg[2][10]  <= n6946;
    \\u4_mem_reg[2][11]  <= n6951;
    \\u4_mem_reg[2][13]  <= n6956;
    \\u4_mem_reg[2][14]  <= n6961;
    \\u4_mem_reg[2][15]  <= n6966;
    \\u4_mem_reg[2][17]  <= n6971;
    \\u4_mem_reg[2][18]  <= n6976;
    \\u4_mem_reg[2][19]  <= n6981;
    \\u4_mem_reg[2][1]  <= n6986;
    \\u4_mem_reg[2][20]  <= n6991;
    \\u4_mem_reg[2][21]  <= n6996;
    \\u4_mem_reg[2][22]  <= n7001;
    \\u4_mem_reg[2][24]  <= n7006;
    \\u4_mem_reg[2][25]  <= n7011;
    \\u4_mem_reg[2][26]  <= n7016;
    \\u4_mem_reg[2][28]  <= n7021;
    \\u4_mem_reg[2][29]  <= n7026;
    \\u4_mem_reg[2][2]  <= n7031;
    \\u4_mem_reg[2][31]  <= n7036;
    \\u4_mem_reg[2][3]  <= n7041;
    \\u4_mem_reg[2][4]  <= n7046;
    \\u4_mem_reg[2][6]  <= n7051;
    \\u4_mem_reg[2][7]  <= n7056;
    \\u4_mem_reg[2][8]  <= n7061;
    \\u4_mem_reg[3][0]  <= n7066;
    \\u4_mem_reg[3][10]  <= n7071;
    \\u4_mem_reg[3][11]  <= n7076;
    \\u4_mem_reg[3][13]  <= n7081;
    \\u4_mem_reg[3][14]  <= n7086;
    \\u4_mem_reg[3][15]  <= n7091;
    \\u4_mem_reg[3][17]  <= n7096;
    \\u4_mem_reg[3][18]  <= n7101;
    \\u4_mem_reg[3][19]  <= n7106;
    \\u4_mem_reg[3][1]  <= n7111;
    \\u4_mem_reg[3][20]  <= n7116;
    \\u4_mem_reg[3][21]  <= n7121;
    \\u4_mem_reg[3][22]  <= n7126;
    \\u4_mem_reg[3][24]  <= n7131;
    \\u4_mem_reg[3][25]  <= n7136;
    \\u4_mem_reg[3][26]  <= n7141;
    \\u4_mem_reg[3][28]  <= n7146;
    \\u4_mem_reg[3][29]  <= n7151;
    \\u4_mem_reg[3][2]  <= n7156;
    \\u4_mem_reg[3][31]  <= n7161;
    \\u4_mem_reg[3][3]  <= n7166;
    \\u4_mem_reg[3][4]  <= n7171;
    \\u4_mem_reg[3][6]  <= n7176;
    \\u4_mem_reg[3][7]  <= n7181;
    \\u4_mem_reg[3][8]  <= n7186;
    \\u3_mem_reg[2][20]  <= n7191;
    \\u5_mem_reg[1][0]  <= n7196;
    \\u5_mem_reg[1][10]  <= n7201;
    \\u5_mem_reg[1][12]  <= n7206;
    \\u5_mem_reg[1][13]  <= n7211;
    \\u5_mem_reg[1][14]  <= n7216;
    \\u7_mem_reg[1][14]  <= n7221;
    \\u5_mem_reg[1][16]  <= n7226;
    \\u5_mem_reg[1][17]  <= n7231;
    \\u5_mem_reg[1][18]  <= n7236;
    \\u5_mem_reg[1][1]  <= n7241;
    \\u5_mem_reg[1][20]  <= n7246;
    \\u5_mem_reg[1][21]  <= n7251;
    \\u5_mem_reg[1][23]  <= n7256;
    \\u5_mem_reg[1][24]  <= n7261;
    \\u5_mem_reg[1][25]  <= n7266;
    \\u5_mem_reg[1][27]  <= n7271;
    \\u5_mem_reg[1][28]  <= n7276;
    \\u5_mem_reg[1][29]  <= n7281;
    \\u5_mem_reg[1][30]  <= n7286;
    \\u5_mem_reg[1][31]  <= n7291;
    \\u5_mem_reg[1][3]  <= n7296;
    \\u5_mem_reg[1][5]  <= n7301;
    \\u5_mem_reg[1][6]  <= n7306;
    \\u5_mem_reg[1][7]  <= n7311;
    \\u5_mem_reg[1][9]  <= n7316;
    \\u5_mem_reg[2][0]  <= n7321;
    \\u5_mem_reg[2][10]  <= n7326;
    \\u5_mem_reg[2][12]  <= n7331;
    \\u5_mem_reg[2][13]  <= n7336;
    \\u5_mem_reg[2][14]  <= n7341;
    \\u5_mem_reg[2][16]  <= n7346;
    \\u5_mem_reg[2][17]  <= n7351;
    \\u5_mem_reg[2][18]  <= n7356;
    \\u5_mem_reg[2][1]  <= n7361;
    \\u5_mem_reg[2][20]  <= n7366;
    \\u5_mem_reg[2][21]  <= n7371;
    \\u5_mem_reg[2][23]  <= n7376;
    \\u5_mem_reg[2][24]  <= n7381;
    \\u5_mem_reg[2][25]  <= n7386;
    \\u5_mem_reg[2][27]  <= n7391;
    \\u5_mem_reg[2][28]  <= n7396;
    \\u5_mem_reg[2][29]  <= n7401;
    \\u5_mem_reg[2][30]  <= n7406;
    \\u5_mem_reg[2][31]  <= n7411;
    \\u5_mem_reg[2][3]  <= n7416;
    \\u5_mem_reg[2][4]  <= n7421;
    \\u5_mem_reg[2][5]  <= n7426;
    \\u5_mem_reg[2][6]  <= n7431;
    \\u5_mem_reg[2][7]  <= n7436;
    \\u5_mem_reg[2][9]  <= n7441;
    \\u5_mem_reg[3][0]  <= n7446;
    \\u5_mem_reg[3][10]  <= n7451;
    \\u5_mem_reg[3][12]  <= n7456;
    \\u5_mem_reg[3][13]  <= n7461;
    \\u5_mem_reg[3][14]  <= n7466;
    \\u5_mem_reg[3][16]  <= n7471;
    \\u5_mem_reg[3][17]  <= n7476;
    \\u5_mem_reg[3][18]  <= n7481;
    \\u5_mem_reg[3][1]  <= n7486;
    \\u5_mem_reg[3][20]  <= n7491;
    \\u5_mem_reg[3][21]  <= n7496;
    \\u6_mem_reg[0][17]  <= n7501;
    \\u5_mem_reg[3][23]  <= n7506;
    \\u5_mem_reg[3][24]  <= n7511;
    \\u5_mem_reg[3][25]  <= n7516;
    \\u5_mem_reg[3][27]  <= n7521;
    \\u5_mem_reg[3][28]  <= n7526;
    \\u5_mem_reg[3][29]  <= n7531;
    \\u5_mem_reg[3][30]  <= n7536;
    \\u5_mem_reg[3][31]  <= n7541;
    \\u5_mem_reg[3][3]  <= n7546;
    \\u5_mem_reg[3][5]  <= n7551;
    \\u5_mem_reg[3][6]  <= n7556;
    \\u5_mem_reg[3][7]  <= n7561;
    \\u5_mem_reg[3][9]  <= n7566;
    \\u6_mem_reg[1][0]  <= n7571;
    \\u6_mem_reg[1][10]  <= n7576;
    \\u6_mem_reg[1][12]  <= n7581;
    \\u6_mem_reg[1][13]  <= n7586;
    \\u6_mem_reg[1][14]  <= n7591;
    \\u6_mem_reg[1][16]  <= n7596;
    \\u6_mem_reg[1][17]  <= n7601;
    \\u6_mem_reg[1][18]  <= n7606;
    \\u6_mem_reg[1][19]  <= n7611;
    \\u6_mem_reg[1][1]  <= n7616;
    \\u6_mem_reg[1][20]  <= n7621;
    \\u6_mem_reg[1][21]  <= n7626;
    \\u6_mem_reg[1][23]  <= n7631;
    \\u6_mem_reg[1][24]  <= n7636;
    \\u6_mem_reg[1][25]  <= n7641;
    \\u6_mem_reg[1][27]  <= n7646;
    \\u6_mem_reg[1][28]  <= n7651;
    \\u6_mem_reg[1][29]  <= n7656;
    \\u6_mem_reg[1][30]  <= n7661;
    \\u6_mem_reg[1][31]  <= n7666;
    \\u6_mem_reg[1][3]  <= n7671;
    \\u6_mem_reg[1][5]  <= n7676;
    \\u6_mem_reg[1][6]  <= n7681;
    \\u6_mem_reg[1][7]  <= n7686;
    \\u6_mem_reg[1][9]  <= n7691;
    \\u6_mem_reg[2][0]  <= n7696;
    \\u6_mem_reg[2][10]  <= n7701;
    \\u6_mem_reg[2][12]  <= n7706;
    \\u6_mem_reg[2][13]  <= n7711;
    \\u6_mem_reg[2][14]  <= n7716;
    \\u6_mem_reg[2][16]  <= n7721;
    \\u6_mem_reg[2][17]  <= n7726;
    \\u6_mem_reg[2][18]  <= n7731;
    \\u6_mem_reg[2][1]  <= n7736;
    \\u6_mem_reg[2][20]  <= n7741;
    \\u6_mem_reg[2][21]  <= n7746;
    \\u6_mem_reg[2][23]  <= n7751;
    \\u6_mem_reg[2][24]  <= n7756;
    \\u6_mem_reg[2][25]  <= n7761;
    \\u6_mem_reg[2][27]  <= n7766;
    \\u6_mem_reg[2][28]  <= n7771;
    \\u6_mem_reg[2][29]  <= n7776;
    \\u6_mem_reg[2][30]  <= n7781;
    \\u6_mem_reg[2][31]  <= n7786;
    \\u6_mem_reg[2][3]  <= n7791;
    \\u6_mem_reg[2][5]  <= n7796;
    \\u6_mem_reg[2][6]  <= n7801;
    \\u6_mem_reg[2][7]  <= n7806;
    \\u6_mem_reg[2][9]  <= n7811;
    \\u6_mem_reg[3][0]  <= n7816;
    \\u6_mem_reg[3][10]  <= n7821;
    \\u6_mem_reg[3][12]  <= n7826;
    \\u6_mem_reg[3][13]  <= n7831;
    \\u6_mem_reg[3][14]  <= n7836;
    \\u6_mem_reg[3][16]  <= n7841;
    \\u6_mem_reg[3][17]  <= n7846;
    \\u6_mem_reg[3][18]  <= n7851;
    \\u6_mem_reg[3][1]  <= n7856;
    \\u6_mem_reg[3][20]  <= n7861;
    \\u6_mem_reg[3][21]  <= n7866;
    \\u6_mem_reg[3][23]  <= n7871;
    \\u6_mem_reg[3][24]  <= n7876;
    \\u6_mem_reg[3][25]  <= n7881;
    \\u6_mem_reg[3][27]  <= n7886;
    \\u6_mem_reg[3][28]  <= n7891;
    \\u6_mem_reg[3][29]  <= n7896;
    \\u6_mem_reg[3][30]  <= n7901;
    \\u6_mem_reg[3][31]  <= n7906;
    \\u6_mem_reg[3][3]  <= n7911;
    \\u6_mem_reg[3][5]  <= n7916;
    \\u6_mem_reg[3][6]  <= n7921;
    \\u6_mem_reg[3][7]  <= n7926;
    \\u6_mem_reg[3][9]  <= n7931;
    \\u3_mem_reg[3][8]  <= n7936;
    \\u7_mem_reg[1][0]  <= n7941;
    \\u7_mem_reg[1][11]  <= n7946;
    \\u7_mem_reg[1][12]  <= n7951;
    \\u7_mem_reg[1][13]  <= n7956;
    \\u7_mem_reg[1][15]  <= n7961;
    \\u7_mem_reg[1][16]  <= n7966;
    \\u7_mem_reg[1][17]  <= n7971;
    \\u7_mem_reg[1][18]  <= n7976;
    \\u7_mem_reg[1][19]  <= n7981;
    \\u7_mem_reg[1][1]  <= n7986;
    \\u7_mem_reg[1][20]  <= n7991;
    \\u7_mem_reg[1][22]  <= n7996;
    \\u7_mem_reg[1][23]  <= n8001;
    \\u7_mem_reg[1][24]  <= n8006;
    \\u7_mem_reg[1][26]  <= n8011;
    \\u7_mem_reg[1][27]  <= n8016;
    \\u7_mem_reg[1][28]  <= n8021;
    \\u7_mem_reg[1][2]  <= n8026;
    \\u7_mem_reg[1][30]  <= n8031;
    \\u7_mem_reg[1][31]  <= n8036;
    \\u7_mem_reg[1][4]  <= n8041;
    \\u7_mem_reg[1][5]  <= n8046;
    \\u7_mem_reg[1][6]  <= n8051;
    \\u7_mem_reg[1][8]  <= n8056;
    \\u7_mem_reg[1][9]  <= n8061;
    \\u7_mem_reg[2][0]  <= n8066;
    \\u7_mem_reg[2][11]  <= n8071;
    \\u7_mem_reg[2][12]  <= n8076;
    \\u7_mem_reg[2][13]  <= n8081;
    \\u7_mem_reg[2][15]  <= n8086;
    \\u7_mem_reg[2][16]  <= n8091;
    \\u7_mem_reg[2][17]  <= n8096;
    \\u7_mem_reg[2][19]  <= n8101;
    \\u7_mem_reg[2][1]  <= n8106;
    \\u7_mem_reg[2][20]  <= n8111;
    \\u7_mem_reg[2][22]  <= n8116;
    \\u7_mem_reg[2][23]  <= n8121;
    \\u7_mem_reg[2][24]  <= n8126;
    \\u7_mem_reg[2][26]  <= n8131;
    \\u7_mem_reg[2][27]  <= n8136;
    \\u7_mem_reg[2][28]  <= n8141;
    \\u7_mem_reg[2][2]  <= n8146;
    \\u7_mem_reg[2][30]  <= n8151;
    \\u7_mem_reg[2][31]  <= n8156;
    \\u7_mem_reg[2][4]  <= n8161;
    \\u7_mem_reg[2][5]  <= n8166;
    \\u7_mem_reg[2][6]  <= n8171;
    \\u7_mem_reg[2][8]  <= n8176;
    \\u7_mem_reg[2][9]  <= n8181;
    \\u7_mem_reg[3][0]  <= n8186;
    \\u7_mem_reg[3][11]  <= n8191;
    \\u7_mem_reg[3][12]  <= n8196;
    \\u7_mem_reg[3][13]  <= n8201;
    \\u7_mem_reg[3][15]  <= n8206;
    \\u7_mem_reg[3][16]  <= n8211;
    \\u7_mem_reg[3][17]  <= n8216;
    \\u7_mem_reg[3][19]  <= n8221;
    \\u7_mem_reg[3][1]  <= n8226;
    \\u7_mem_reg[3][20]  <= n8231;
    \\u6_mem_reg[0][20]  <= n8236;
    \\u7_mem_reg[3][22]  <= n8241;
    \\u7_mem_reg[3][23]  <= n8246;
    \\u7_mem_reg[3][24]  <= n8251;
    \\u7_mem_reg[3][26]  <= n8256;
    \\u7_mem_reg[3][27]  <= n8261;
    \\u7_mem_reg[3][28]  <= n8266;
    \\u7_mem_reg[3][2]  <= n8271;
    \\u7_mem_reg[3][30]  <= n8276;
    \\u7_mem_reg[3][31]  <= n8281;
    \\u7_mem_reg[3][4]  <= n8286;
    \\u7_mem_reg[3][5]  <= n8291;
    \\u7_mem_reg[3][6]  <= n8296;
    \\u7_mem_reg[3][8]  <= n8301;
    \\u7_mem_reg[3][9]  <= n8306;
    \\u8_mem_reg[1][0]  <= n8311;
    \\u8_mem_reg[1][11]  <= n8316;
    \\u8_mem_reg[1][12]  <= n8321;
    \\u8_mem_reg[1][13]  <= n8326;
    \\u8_mem_reg[1][15]  <= n8331;
    \\u8_mem_reg[1][16]  <= n8336;
    \\u8_mem_reg[1][17]  <= n8341;
    \\u8_mem_reg[1][19]  <= n8346;
    \\u8_mem_reg[1][1]  <= n8351;
    \\u8_mem_reg[1][20]  <= n8356;
    \\u8_mem_reg[1][22]  <= n8361;
    \\u8_mem_reg[1][23]  <= n8366;
    \\u8_mem_reg[1][24]  <= n8371;
    \\u8_mem_reg[1][26]  <= n8376;
    \\u3_mem_reg[1][0]  <= n8381;
    \\u8_mem_reg[1][27]  <= n8386;
    \\u3_mem_reg[1][10]  <= n8391;
    \\u8_mem_reg[1][29]  <= n8396;
    \\u8_mem_reg[1][2]  <= n8401;
    \\u8_mem_reg[1][30]  <= n8406;
    \\u8_mem_reg[1][31]  <= n8411;
    \\u3_mem_reg[1][12]  <= n8416;
    \\u8_mem_reg[1][4]  <= n8421;
    \\u3_mem_reg[1][13]  <= n8426;
    \\u8_mem_reg[1][5]  <= n8431;
    \\u3_mem_reg[1][14]  <= n8436;
    \\u8_mem_reg[1][7]  <= n8441;
    \\u8_mem_reg[1][8]  <= n8446;
    \\u8_mem_reg[1][9]  <= n8451;
    \\u8_mem_reg[2][0]  <= n8456;
    \\u3_mem_reg[1][16]  <= n8461;
    \\u8_mem_reg[2][10]  <= n8466;
    \\u8_mem_reg[2][11]  <= n8471;
    \\u3_mem_reg[1][17]  <= n8476;
    \\u8_mem_reg[2][12]  <= n8481;
    \\u3_mem_reg[1][18]  <= n8486;
    \\u8_mem_reg[2][14]  <= n8491;
    \\u8_mem_reg[2][15]  <= n8496;
    \\u8_mem_reg[2][16]  <= n8501;
    \\u8_mem_reg[2][17]  <= n8506;
    \\u3_mem_reg[1][1]  <= n8511;
    \\u8_mem_reg[2][19]  <= n8516;
    \\u3_mem_reg[1][20]  <= n8521;
    \\u8_mem_reg[2][1]  <= n8526;
    \\u3_mem_reg[1][21]  <= n8531;
    \\u8_mem_reg[2][21]  <= n8536;
    \\u8_mem_reg[2][22]  <= n8541;
    \\u8_mem_reg[2][23]  <= n8546;
    \\u8_mem_reg[2][24]  <= n8551;
    \\u3_mem_reg[1][23]  <= n8556;
    \\u8_mem_reg[2][26]  <= n8561;
    \\u3_mem_reg[1][24]  <= n8566;
    \\u8_mem_reg[2][27]  <= n8571;
    \\u3_mem_reg[1][25]  <= n8576;
    \\u8_mem_reg[2][29]  <= n8581;
    \\u8_mem_reg[2][2]  <= n8586;
    \\u8_mem_reg[2][30]  <= n8591;
    \\u8_mem_reg[2][31]  <= n8596;
    \\u3_mem_reg[1][27]  <= n8601;
    \\u4_mem_reg[0][0]  <= n8606;
    \\u4_mem_reg[0][10]  <= n8611;
    \\u4_mem_reg[0][11]  <= n8616;
    \\u4_mem_reg[0][15]  <= n8621;
    \\u4_mem_reg[0][18]  <= n8626;
    \\u4_mem_reg[0][1]  <= n8631;
    \\u4_mem_reg[0][21]  <= n8636;
    \\u4_mem_reg[0][25]  <= n8641;
    \\u4_mem_reg[0][27]  <= n8646;
    \\u4_mem_reg[0][28]  <= n8651;
    \\u4_mem_reg[0][26]  <= n8656;
    \\u4_mem_reg[0][2]  <= n8661;
    \\u4_mem_reg[0][29]  <= n8666;
    \\u4_mem_reg[0][3]  <= n8671;
    \\u4_mem_reg[0][5]  <= n8676;
    \\u4_mem_reg[0][8]  <= n8681;
    \\u5_mem_reg[0][10]  <= n8686;
    \\u5_mem_reg[0][11]  <= n8691;
    \\u5_mem_reg[0][15]  <= n8696;
    \\u5_mem_reg[0][18]  <= n8701;
    \\u5_mem_reg[0][1]  <= n8706;
    \\u5_mem_reg[0][21]  <= n8711;
    \\u13_intm_r_reg[8]  <= n8716;
    \\u5_mem_reg[0][26]  <= n8721;
    \\u5_mem_reg[0][27]  <= n8726;
    \\u5_mem_reg[0][25]  <= n8731;
    \\u5_mem_reg[0][2]  <= n8736;
    \\u5_mem_reg[0][29]  <= n8741;
    \\u5_mem_reg[0][3]  <= n8746;
    \\u5_mem_reg[0][5]  <= n8751;
    \\u5_mem_reg[0][8]  <= n8756;
    \\u6_mem_reg[0][10]  <= n8761;
    \\u6_mem_reg[0][11]  <= n8766;
    \\u6_mem_reg[0][15]  <= n8771;
    \\u7_mem_reg[1][21]  <= n8776;
    \\u6_mem_reg[0][18]  <= n8781;
    \\u6_mem_reg[0][1]  <= n8786;
    \\u6_mem_reg[0][21]  <= n8791;
    \\u6_mem_reg[0][26]  <= n8796;
    \\u6_mem_reg[0][27]  <= n8801;
    \\u6_mem_reg[0][25]  <= n8806;
    \\u6_mem_reg[0][2]  <= n8811;
    \\u6_mem_reg[0][29]  <= n8816;
    \\u6_mem_reg[0][3]  <= n8821;
    \\u6_mem_reg[0][5]  <= n8826;
    \\u6_mem_reg[0][8]  <= n8831;
    \\u7_mem_reg[0][10]  <= n8836;
    \\u7_mem_reg[0][11]  <= n8841;
    \\u7_mem_reg[0][15]  <= n8846;
    \\u7_mem_reg[0][18]  <= n8851;
    \\u7_mem_reg[0][1]  <= n8856;
    \\u7_mem_reg[0][21]  <= n8861;
    \\u7_mem_reg[0][25]  <= n8866;
    \\u7_mem_reg[0][27]  <= n8871;
    \\u7_mem_reg[0][28]  <= n8876;
    \\u7_mem_reg[0][26]  <= n8881;
    \\u7_mem_reg[0][2]  <= n8886;
    \\u7_mem_reg[0][29]  <= n8891;
    \\u7_mem_reg[0][3]  <= n8896;
    \\u7_mem_reg[0][5]  <= n8901;
    \\u7_mem_reg[0][8]  <= n8906;
    \\u3_mem_reg[0][10]  <= n8911;
    \\u8_mem_reg[0][10]  <= n8916;
    \\u8_mem_reg[0][13]  <= n8921;
    \\u3_mem_reg[0][18]  <= n8926;
    \\u8_mem_reg[0][14]  <= n8931;
    \\u3_mem_reg[0][19]  <= n8936;
    \\u8_mem_reg[0][18]  <= n8941;
    \\u8_mem_reg[0][19]  <= n8946;
    \\u3_mem_reg[0][20]  <= n8951;
    \\u8_mem_reg[0][20]  <= n8956;
    \\u8_mem_reg[0][21]  <= n8961;
    \\u3_mem_reg[0][22]  <= n8966;
    \\u8_mem_reg[0][23]  <= n8971;
    \\u8_mem_reg[0][24]  <= n8976;
    \\u8_mem_reg[0][25]  <= n8981;
    \\u3_mem_reg[0][24]  <= n8986;
    \\u3_mem_reg[0][25]  <= n8991;
    \\u3_mem_reg[0][26]  <= n8996;
    \\u3_mem_reg[0][28]  <= n9001;
    \\u8_mem_reg[0][7]  <= n9006;
    \\u8_mem_reg[0][8]  <= n9011;
    \\u8_mem_reg[0][6]  <= n9016;
    \\u8_mem_reg[0][9]  <= n9021;
    \\u3_mem_reg[0][30]  <= n9026;
    \\u3_mem_reg[0][3]  <= n9031;
    \\u3_mem_reg[0][8]  <= n9036;
    \\u7_mem_reg[1][10]  <= n9041;
    \\u13_crac_dout_r_reg[7]  <= n9046;
    \\u6_mem_reg[2][22]  <= n9051;
    \\u6_mem_reg[0][0]  <= n9056;
    \\u6_mem_reg[3][4]  <= n9061;
    \\u13_intm_r_reg[26]  <= n9066;
    \\u6_mem_reg[3][2]  <= n9071;
    \\u13_occ0_r_reg[22]  <= n9076;
    \\u6_mem_reg[3][26]  <= n9081;
    \\u6_mem_reg[3][22]  <= n9086;
    \\u6_mem_reg[3][15]  <= n9091;
    \\u5_mem_reg[0][6]  <= n9096;
    \\u6_mem_reg[3][19]  <= n9101;
    \\u1_sr_reg[10]  <= n9106;
    \\u5_mem_reg[0][30]  <= n9111;
    \\u5_mem_reg[0][23]  <= n9116;
    \\u13_crac_r_reg[2]  <= n9121;
    \\u6_mem_reg[2][4]  <= n9126;
    \\u6_mem_reg[3][11]  <= n9131;
    \\u6_mem_reg[2][8]  <= n9136;
    \\u6_mem_reg[2][2]  <= n9141;
    \\u3_mem_reg[0][9]  <= n9146;
    \\u13_occ0_r_reg[26]  <= n9151;
    \\u5_mem_reg[0][28]  <= n9156;
    \\u13_intm_r_reg[3]  <= n9161;
    \\u6_mem_reg[2][26]  <= n9166;
    \\u3_mem_reg[0][4]  <= n9171;
    \\u5_mem_reg[0][20]  <= n9176;
    \\u8_mem_reg[0][31]  <= n9181;
    \\u6_mem_reg[2][15]  <= n9186;
    \\u6_mem_reg[1][15]  <= n9191;
    \\u6_mem_reg[2][19]  <= n9196;
    \\u6_mem_reg[2][11]  <= n9201;
    \\u5_mem_reg[0][17]  <= n9206;
    \\u13_occ0_r_reg[19]  <= n9211;
    \\u5_mem_reg[0][12]  <= n9216;
    \\u6_mem_reg[1][26]  <= n9221;
    \\u4_mem_reg[0][6]  <= n9226;
    \\u6_mem_reg[1][4]  <= n9231;
    \\u6_mem_reg[1][8]  <= n9236;
    \\u6_mem_reg[1][2]  <= n9241;
    \\u5_mem_reg[0][0]  <= n9246;
    \\u6_mem_reg[1][22]  <= n9251;
    \\u8_mem_reg[0][3]  <= n9256;
    \\u4_mem_reg[0][30]  <= n9261;
    \\u8_mem_reg[0][16]  <= n9266;
    \\u5_mem_reg[3][8]  <= n9271;
    \\u6_mem_reg[1][11]  <= n9276;
    \\u5_mem_reg[3][4]  <= n9281;
    \\u8_mem_reg[0][2]  <= n9286;
    \\u5_mem_reg[2][8]  <= n9291;
    \\u4_mem_reg[0][23]  <= n9296;
    \\u3_mem_reg[0][23]  <= n9301;
    \\u4_mem_reg[0][17]  <= n9306;
    \\u5_mem_reg[3][19]  <= n9311;
    \\u5_mem_reg[3][26]  <= n9316;
    \\u5_mem_reg[3][2]  <= n9321;
    \\u5_mem_reg[3][22]  <= n9326;
    \\u5_mem_reg[3][15]  <= n9331;
    \\u8_mem_reg[0][27]  <= n9336;
    \\u4_mem_reg[0][20]  <= n9341;
    \\u5_mem_reg[3][11]  <= n9346;
    \\u5_mem_reg[2][2]  <= n9351;
    \\u4_mem_reg[0][12]  <= n9356;
    \\u5_mem_reg[2][26]  <= n9361;
    \\u8_mem_reg[0][22]  <= n9366;
    \\u13_occ0_r_reg[15]  <= n9371;
    \\u5_mem_reg[1][2]  <= n9376;
    \\u5_mem_reg[2][11]  <= n9381;
    \\u3_mem_reg[1][26]  <= n9386;
    \\u5_mem_reg[2][19]  <= n9391;
    \\u5_mem_reg[2][22]  <= n9396;
    \\u5_mem_reg[2][15]  <= n9401;
    \\u8_mem_reg[2][3]  <= n9406;
    \\u5_mem_reg[1][8]  <= n9411;
    \\u5_mem_reg[1][4]  <= n9416;
    \\u8_mem_reg[0][1]  <= n9421;
    \\u13_occ1_r_reg[11]  <= n9426;
    \\u3_mem_reg[0][0]  <= n9431;
    u14_u8_en_out_l2_reg <= n9436;
    \\u12_wb_data_o_reg[4]  <= n9441;
    \\u12_wb_data_o_reg[6]  <= n9446;
    \\u12_wb_data_o_reg[10]  <= n9451;
    \\u13_occ1_r_reg[8]  <= n9456;
    \\u13_occ1_r_reg[0]  <= n9461;
    \\u13_occ1_r_reg[10]  <= n9466;
    \\u13_occ1_r_reg[12]  <= n9471;
    \\u13_occ1_r_reg[13]  <= n9476;
    \\u13_occ1_r_reg[14]  <= n9481;
    \\u13_occ1_r_reg[1]  <= n9486;
    \\u13_occ1_r_reg[2]  <= n9491;
    \\u13_occ1_r_reg[3]  <= n9496;
    \\u13_occ1_r_reg[5]  <= n9501;
    \\u13_occ1_r_reg[6]  <= n9506;
    \\u13_occ1_r_reg[7]  <= n9511;
    \\u1_slt1_reg[7]  <= n9516;
    \\u1_slt2_reg[7]  <= n9521;
    \\u1_slt4_reg[7]  <= n9526;
    \\u1_slt3_reg[7]  <= n9531;
    \\u3_mem_reg[0][14]  <= n9536;
    \\u3_mem_reg[0][7]  <= n9541;
    u14_u6_full_empty_r_reg <= n9546;
    u14_u8_full_empty_r_reg <= n9551;
    \\u12_wb_data_o_reg[0]  <= n9556;
    \\u12_wb_data_o_reg[14]  <= n9561;
    \\u12_wb_data_o_reg[13]  <= n9566;
    \\u12_wb_data_o_reg[12]  <= n9571;
    \\u12_wb_data_o_reg[11]  <= n9576;
    \\u12_wb_data_o_reg[9]  <= n9581;
    \\u12_wb_data_o_reg[7]  <= n9586;
    \\u12_wb_data_o_reg[15]  <= n9591;
    \\u12_wb_data_o_reg[5]  <= n9596;
    \\u12_wb_data_o_reg[3]  <= n9601;
    \\u12_wb_data_o_reg[8]  <= n9606;
    \\u12_wb_data_o_reg[2]  <= n9611;
    \\u13_occ1_r_reg[9]  <= n9616;
    \\u13_occ1_r_reg[15]  <= n9621;
    \\u3_mem_reg[0][31]  <= n9626;
    \\u13_occ1_r_reg[4]  <= n9631;
    \\u0_slt9_r_reg[1]  <= n9636;
    \\u1_slt6_reg[7]  <= n9641;
    u14_u7_en_out_l2_reg <= n9646;
    u14_u7_full_empty_r_reg <= n9651;
    u13_ac97_rst_force_reg <= n9656;
    u13_resume_req_reg <= n9661;
    \\u1_sr_reg[9]  <= n9666;
    u14_u6_en_out_l2_reg <= n9671;
    \\u12_wb_data_o_reg[31]  <= n9676;
    \\u1_slt3_reg[6]  <= n9681;
    \\u1_slt1_reg[6]  <= n9686;
    \\u1_slt2_reg[6]  <= n9691;
    \\u1_slt4_reg[6]  <= n9696;
    \\u12_wb_data_o_reg[23]  <= n9701;
    \\u12_wb_data_o_reg[22]  <= n9706;
    \\u12_wb_data_o_reg[21]  <= n9711;
    \\u12_wb_data_o_reg[16]  <= n9716;
    \\u12_wb_data_o_reg[20]  <= n9721;
    \\u12_wb_data_o_reg[19]  <= n9726;
    \\u12_wb_data_o_reg[17]  <= n9731;
    \\u12_wb_data_o_reg[24]  <= n9736;
    \\u12_wb_data_o_reg[30]  <= n9741;
    \\u12_wb_data_o_reg[28]  <= n9746;
    \\u12_wb_data_o_reg[27]  <= n9751;
    \\u12_wb_data_o_reg[26]  <= n9756;
    \\u12_wb_data_o_reg[29]  <= n9761;
    \\u12_wb_data_o_reg[25]  <= n9766;
    \\u1_slt6_reg[6]  <= n9771;
    \\u12_wb_data_o_reg[18]  <= n9776;
    u4_empty_reg <= n9781;
    u6_empty_reg <= n9786;
    u15_crac_we_r_reg <= n9791;
    \\u1_sr_reg[8]  <= n9796;
    u3_empty_reg <= n9801;
    u5_empty_reg <= n9806;
    u7_empty_reg <= n9811;
    u8_empty_reg <= n9816;
    \\u10_rp_reg[2]  <= n9821;
    \\u11_rp_reg[2]  <= n9826;
    \\u23_int_set_reg[1]  <= n9831;
    \\u24_int_set_reg[1]  <= n9836;
    \\u11_rp_reg[1]  <= n9841;
    \\u9_rp_reg[1]  <= n9846;
    \\u10_rp_reg[1]  <= n9851;
    \\u11_rp_reg[0]  <= n9856;
    \\u9_rp_reg[0]  <= n9861;
    \\u9_rp_reg[2]  <= n9866;
    \\u10_rp_reg[0]  <= n9871;
    \\u1_slt1_reg[5]  <= n9876;
    \\u1_slt2_reg[5]  <= n9881;
    \\u1_slt4_reg[5]  <= n9886;
    \\u1_slt3_reg[5]  <= n9891;
    \\u1_slt6_reg[5]  <= n9896;
    \\u25_int_set_reg[1]  <= n9901;
    \\u1_sr_reg[7]  <= n9906;
    \\u0_slt9_r_reg[0]  <= n9911;
    valid_s_reg <= n9916;
    \\in_valid_s_reg[0]  <= n9921;
    \\u1_slt2_reg[4]  <= n9926;
    \\u1_slt3_reg[4]  <= n9931;
    \\u1_slt4_reg[4]  <= n9936;
    \\u1_slt6_reg[4]  <= n9941;
    u12_o7_we_reg <= n9946;
    u12_o3_we_reg <= n9951;
    u12_o4_we_reg <= n9956;
    u12_o6_we_reg <= n9961;
    u12_o8_we_reg <= n9966;
    u12_o9_we_reg <= n9971;
    \\u1_sr_reg[6]  <= n9976;
    \\in_valid_s_reg[2]  <= n9981;
    \\u2_to_cnt_reg[5]  <= n9986;
    u13_int_reg <= n9991;
    \\u13_ints_r_reg[21]  <= n9996;
    \\u1_slt3_reg[0]  <= n10001;
    \\u13_ints_r_reg[0]  <= n10006;
    \\u13_ints_r_reg[27]  <= n10011;
    \\u13_ints_r_reg[15]  <= n10016;
    \\u2_cnt_reg[7]  <= n10021;
    \\in_valid_s_reg[1]  <= n10026;
    valid_s1_reg <= n10031;
    \\in_valid_s1_reg[0]  <= n10036;
    \\u2_to_cnt_reg[3]  <= n10041;
    \\u2_res_cnt_reg[3]  <= n10046;
    \\u2_to_cnt_reg[4]  <= n10051;
    \\u1_slt3_reg[2]  <= n10056;
    \\u1_slt3_reg[1]  <= n10061;
    \\u1_slt4_reg[1]  <= n10066;
    \\u1_slt6_reg[1]  <= n10071;
    \\u1_slt6_reg[2]  <= n10076;
    u12_wb_ack_o_reg <= n10081;
    \\u13_ints_r_reg[10]  <= n10086;
    \\u13_ints_r_reg[12]  <= n10091;
    \\u13_ints_r_reg[13]  <= n10096;
    \\u13_ints_r_reg[16]  <= n10101;
    \\u13_ints_r_reg[18]  <= n10106;
    \\u13_ints_r_reg[19]  <= n10111;
    \\u13_ints_r_reg[22]  <= n10116;
    \\u13_ints_r_reg[24]  <= n10121;
    \\u13_ints_r_reg[25]  <= n10126;
    \\u13_ints_r_reg[28]  <= n10131;
    \\u13_ints_r_reg[3]  <= n10136;
    \\u13_ints_r_reg[4]  <= n10141;
    \\u13_ints_r_reg[7]  <= n10146;
    \\u13_ints_r_reg[6]  <= n10151;
    \\u1_slt6_reg[3]  <= n10156;
    \\u1_slt6_reg[0]  <= n10161;
    \\u1_slt4_reg[3]  <= n10166;
    \\u1_slt3_reg[3]  <= n10171;
    \\u13_ints_r_reg[9]  <= n10176;
    \\u1_slt4_reg[2]  <= n10181;
    \\u1_slt4_reg[0]  <= n10186;
    \\u2_cnt_reg[1]  <= n10191;
    \\u2_to_cnt_reg[2]  <= n10196;
    \\u4_status_reg[1]  <= n10201;
    \\u5_status_reg[1]  <= n10206;
    u12_rf_we_reg <= n10211;
    \\u2_res_cnt_reg[0]  <= n10216;
    \\in_valid_s1_reg[2]  <= n10221;
    \\u1_sr_reg[5]  <= n10226;
    \\u2_cnt_reg[4]  <= n10231;
    \\u2_cnt_reg[3]  <= n10236;
    \\u2_to_cnt_reg[0]  <= n10241;
    \\u2_to_cnt_reg[1]  <= n10246;
    \\u2_cnt_reg[5]  <= n10251;
    \\u2_cnt_reg[6]  <= n10256;
    \\u2_cnt_reg[0]  <= n10261;
    \\u2_cnt_reg[2]  <= n10266;
    \\u2_res_cnt_reg[2]  <= n10271;
    u2_valid_reg <= n10276;
    \\u2_res_cnt_reg[1]  <= n10281;
    \\u3_status_reg[1]  <= n10286;
    \\u6_status_reg[1]  <= n10291;
    \\u7_status_reg[1]  <= n10296;
    \\u8_status_reg[1]  <= n10301;
    \\u11_status_reg[1]  <= n10306;
    u10_empty_reg <= n10311;
    u9_empty_reg <= n10316;
    \\in_valid_s1_reg[1]  <= n10321;
    \\u2_in_valid_reg[0]  <= n10326;
    u12_we1_reg <= n10331;
    \\u1_sr_reg[4]  <= n10336;
    \\u2_in_valid_reg[2]  <= n10341;
    \\u10_status_reg[1]  <= n10346;
    \\u9_status_reg[1]  <= n10351;
    u11_empty_reg <= n10356;
    u2_sync_beat_reg <= n10361;
    u11_full_reg <= n10366;
    \\u10_dout_reg[14]  <= n10371;
    \\u10_dout_reg[15]  <= n10376;
    \\u10_dout_reg[17]  <= n10381;
    \\u10_dout_reg[18]  <= n10386;
    \\u10_dout_reg[19]  <= n10391;
    \\u10_dout_reg[1]  <= n10396;
    \\u10_dout_reg[20]  <= n10401;
    \\u10_dout_reg[21]  <= n10406;
    \\u10_dout_reg[22]  <= n10411;
    \\u10_dout_reg[23]  <= n10416;
    u12_i4_re_reg <= n10421;
    u2_ld_reg <= n10426;
    u9_full_reg <= n10431;
    u12_i6_re_reg <= n10436;
    \\u2_out_le_reg[1]  <= n10441;
    u12_i3_re_reg <= n10446;
    \\u2_in_valid_reg[1]  <= n10451;
    \\u10_dout_reg[11]  <= n10456;
    \\u10_dout_reg[0]  <= n10461;
    \\u10_dout_reg[10]  <= n10466;
    \\u10_dout_reg[12]  <= n10471;
    \\u10_dout_reg[13]  <= n10476;
    \\u10_dout_reg[25]  <= n10481;
    \\u10_dout_reg[27]  <= n10486;
    \\u10_dout_reg[28]  <= n10491;
    \\u10_dout_reg[29]  <= n10496;
    \\u10_dout_reg[2]  <= n10501;
    \\u10_dout_reg[30]  <= n10506;
    \\u10_dout_reg[3]  <= n10511;
    \\u10_dout_reg[4]  <= n10516;
    \\u10_dout_reg[6]  <= n10521;
    \\u10_dout_reg[7]  <= n10526;
    \\u10_dout_reg[8]  <= n10531;
    \\u10_dout_reg[9]  <= n10536;
    u10_full_reg <= n10541;
    \\u2_out_le_reg[2]  <= n10546;
    \\u2_out_le_reg[4]  <= n10551;
    \\u2_out_le_reg[5]  <= n10556;
    \\u2_out_le_reg[3]  <= n10561;
    \\u2_out_le_reg[0]  <= n10566;
    \\u9_dout_reg[11]  <= n10571;
    \\u9_dout_reg[14]  <= n10576;
    \\u9_dout_reg[18]  <= n10581;
    \\u9_dout_reg[19]  <= n10586;
    \\u9_dout_reg[20]  <= n10591;
    \\u9_dout_reg[21]  <= n10596;
    \\u9_dout_reg[22]  <= n10601;
    \\u9_dout_reg[23]  <= n10606;
    \\u9_dout_reg[24]  <= n10611;
    \\u9_dout_reg[25]  <= n10616;
    \\u9_dout_reg[16]  <= n10621;
    \\u10_dout_reg[16]  <= n10626;
    \\u9_dout_reg[26]  <= n10631;
    \\u9_dout_reg[27]  <= n10636;
    \\u9_dout_reg[28]  <= n10641;
    \\u9_dout_reg[29]  <= n10646;
    \\u9_dout_reg[2]  <= n10651;
    \\u9_dout_reg[30]  <= n10656;
    \\u9_dout_reg[31]  <= n10661;
    \\u9_dout_reg[3]  <= n10666;
    \\u1_sr_reg[3]  <= n10671;
    \\u9_dout_reg[4]  <= n10676;
    \\u9_dout_reg[5]  <= n10681;
    \\u9_dout_reg[6]  <= n10686;
    \\u9_dout_reg[7]  <= n10691;
    \\u9_dout_reg[8]  <= n10696;
    \\u9_dout_reg[9]  <= n10701;
    \\u10_dout_reg[24]  <= n10706;
    \\u10_dout_reg[26]  <= n10711;
    \\u9_dout_reg[13]  <= n10716;
    \\u11_dout_reg[0]  <= n10721;
    \\u11_dout_reg[10]  <= n10726;
    \\u11_dout_reg[11]  <= n10731;
    \\u11_dout_reg[12]  <= n10736;
    \\u11_dout_reg[13]  <= n10741;
    \\u10_dout_reg[31]  <= n10746;
    \\u11_dout_reg[14]  <= n10751;
    \\u11_dout_reg[15]  <= n10756;
    \\u11_dout_reg[16]  <= n10761;
    \\u11_dout_reg[17]  <= n10766;
    \\u11_dout_reg[18]  <= n10771;
    \\u11_dout_reg[19]  <= n10776;
    \\u10_dout_reg[5]  <= n10781;
    \\u11_dout_reg[1]  <= n10786;
    \\u11_dout_reg[20]  <= n10791;
    \\u11_dout_reg[21]  <= n10796;
    \\u11_dout_reg[22]  <= n10801;
    \\u11_dout_reg[23]  <= n10806;
    \\u11_dout_reg[24]  <= n10811;
    \\u11_dout_reg[25]  <= n10816;
    \\u11_dout_reg[26]  <= n10821;
    \\u11_dout_reg[27]  <= n10826;
    \\u11_dout_reg[28]  <= n10831;
    \\u11_dout_reg[29]  <= n10836;
    \\u11_dout_reg[2]  <= n10841;
    \\u11_dout_reg[30]  <= n10846;
    \\u11_dout_reg[31]  <= n10851;
    \\u11_dout_reg[3]  <= n10856;
    \\u11_dout_reg[4]  <= n10861;
    \\u11_dout_reg[5]  <= n10866;
    \\u11_dout_reg[6]  <= n10871;
    \\u11_dout_reg[7]  <= n10876;
    \\u11_dout_reg[8]  <= n10881;
    \\u11_dout_reg[9]  <= n10886;
    \\u9_dout_reg[15]  <= n10891;
    \\u9_dout_reg[17]  <= n10896;
    \\u9_dout_reg[0]  <= n10901;
    \\u9_dout_reg[12]  <= n10906;
    \\u9_dout_reg[10]  <= n10911;
    \\u9_dout_reg[1]  <= n10916;
    u12_re2_reg <= n10921;
    u12_re1_reg <= n10926;
    u2_bit_clk_e_reg <= n10931;
    u2_suspended_reg <= n10936;
    \\u10_status_reg[0]  <= n10941;
    \\u9_status_reg[0]  <= n10946;
    \\u11_status_reg[0]  <= n10951;
    \\u6_status_reg[0]  <= n10956;
    \\u3_status_reg[0]  <= n10961;
    \\u4_status_reg[0]  <= n10966;
    \\u7_status_reg[0]  <= n10971;
    \\u1_sr_reg[2]  <= n10976;
    \\u15_crac_din_reg[6]  <= n10981;
    \\u15_crac_din_reg[9]  <= n10986;
    \\u15_crac_din_reg[12]  <= n10991;
    \\u15_crac_din_reg[1]  <= n10996;
    \\u15_crac_din_reg[7]  <= n11001;
    \\u15_crac_din_reg[14]  <= n11006;
    \\u15_crac_din_reg[10]  <= n11011;
    \\u15_crac_din_reg[15]  <= n11016;
    \\u15_crac_din_reg[4]  <= n11021;
    \\u15_crac_din_reg[8]  <= n11026;
    \\u15_crac_din_reg[11]  <= n11031;
    \\u15_crac_din_reg[13]  <= n11036;
    \\u15_crac_din_reg[2]  <= n11041;
    \\u15_crac_din_reg[0]  <= n11046;
    \\u15_crac_din_reg[5]  <= n11051;
    \\u5_status_reg[0]  <= n11056;
    \\u8_status_reg[0]  <= n11061;
    \\u15_crac_din_reg[3]  <= n11066;
    \\u1_sr_reg[1]  <= n11071;
    u12_we2_reg <= n11076;
    u2_bit_clk_r1_reg <= n11081;
    \\u1_sr_reg[0]  <= n11086;
    u1_sdata_in_r_reg <= n11091;
    \\u12_dout_reg[7]  <= n11096;
    \\u12_dout_reg[4]  <= n11101;
    \\u12_dout_reg[12]  <= n11106;
    \\u12_dout_reg[24]  <= n11111;
    \\u12_dout_reg[26]  <= n11116;
    \\u12_dout_reg[23]  <= n11121;
    \\u12_dout_reg[11]  <= n11126;
    \\u12_dout_reg[31]  <= n11131;
    \\u12_dout_reg[13]  <= n11136;
    \\u12_dout_reg[29]  <= n11141;
    \\u12_dout_reg[22]  <= n11146;
    \\u12_dout_reg[30]  <= n11151;
    \\u12_dout_reg[15]  <= n11156;
    \\u12_dout_reg[19]  <= n11161;
    u2_bit_clk_r_reg <= n11166;
    \\u12_dout_reg[27]  <= n11171;
    \\u12_dout_reg[28]  <= n11176;
    \\u12_dout_reg[10]  <= n11181;
    \\u12_dout_reg[6]  <= n11186;
    \\u12_dout_reg[20]  <= n11191;
    \\u12_dout_reg[0]  <= n11196;
    \\u12_dout_reg[21]  <= n11201;
    \\u12_dout_reg[5]  <= n11206;
    \\u12_dout_reg[18]  <= n11211;
    \\u12_dout_reg[25]  <= n11216;
    \\u12_dout_reg[2]  <= n11221;
    \\u12_dout_reg[9]  <= n11226;
    \\u12_dout_reg[17]  <= n11231;
    \\u12_dout_reg[3]  <= n11236;
    \\u12_dout_reg[8]  <= n11241;
    \\u12_dout_reg[16]  <= n11246;
    \\u12_dout_reg[14]  <= n11251;
    \\u12_dout_reg[1]  <= n11256;
  end
  initial begin
    u16_u1_dma_req_reg <= 1'b0;
    u16_u3_dma_req_reg <= 1'b0;
    u16_u0_dma_req_reg <= 1'b0;
    u16_u2_dma_req_reg <= 1'b0;
    u16_u4_dma_req_reg <= 1'b0;
    u16_u5_dma_req_reg <= 1'b0;
    \\u13_ints_r_reg[11]  <= 1'b0;
    \\u13_ints_r_reg[5]  <= 1'b0;
    \\u13_ints_r_reg[14]  <= 1'b0;
    \\u13_ints_r_reg[17]  <= 1'b0;
    \\u13_ints_r_reg[2]  <= 1'b0;
    \\u13_ints_r_reg[8]  <= 1'b0;
    u16_u8_dma_req_reg <= 1'b0;
    u16_u6_dma_req_reg <= 1'b0;
    u16_u7_dma_req_reg <= 1'b0;
    u15_crac_rd_reg <= 1'b0;
    \\u17_int_set_reg[1]  <= 1'b0;
    \\u20_int_set_reg[1]  <= 1'b0;
    \\u21_int_set_reg[1]  <= 1'b0;
    \\u22_int_set_reg[1]  <= 1'b0;
    \\u25_int_set_reg[2]  <= 1'b0;
    \\u18_int_set_reg[1]  <= 1'b0;
    \\u19_int_set_reg[1]  <= 1'b0;
    \\u24_int_set_reg[2]  <= 1'b0;
    u15_crac_wr_reg <= 1'b0;
    \\u13_ints_r_reg[1]  <= 1'b0;
    \\u13_ints_r_reg[26]  <= 1'b0;
    u15_rdd1_reg <= 1'b0;
    u15_rdd2_reg <= 1'b0;
    \\u20_int_set_reg[0]  <= 1'b0;
    \\u18_int_set_reg[0]  <= 1'b0;
    \\u13_ints_r_reg[23]  <= 1'b0;
    \\u13_ints_r_reg[20]  <= 1'b0;
    u15_rdd3_reg <= 1'b0;
    \\u21_int_set_reg[0]  <= 1'b0;
    \\u22_int_set_reg[0]  <= 1'b0;
    \\u17_int_set_reg[0]  <= 1'b0;
    \\u19_int_set_reg[0]  <= 1'b0;
    \\u23_int_set_reg[2]  <= 1'b0;
    u2_sync_resume_reg <= 1'b0;
    \\u26_ps_cnt_reg[5]  <= 1'b0;
    \\u26_ps_cnt_reg[2]  <= 1'b0;
    \\u26_ps_cnt_reg[0]  <= 1'b0;
    \\u26_ps_cnt_reg[1]  <= 1'b0;
    \\u26_ps_cnt_reg[4]  <= 1'b0;
    \\u26_ps_cnt_reg[3]  <= 1'b0;
    \\u17_int_set_reg[2]  <= 1'b0;
    \\u18_int_set_reg[2]  <= 1'b0;
    \\u21_int_set_reg[2]  <= 1'b0;
    \\u20_int_set_reg[2]  <= 1'b0;
    \\u22_int_set_reg[2]  <= 1'b0;
    \\u19_int_set_reg[2]  <= 1'b0;
    \\u25_int_set_reg[0]  <= 1'b0;
    u26_ac97_rst__reg <= 1'b0;
    \\u26_cnt_reg[2]  <= 1'b0;
    \\u23_int_set_reg[0]  <= 1'b0;
    \\u24_int_set_reg[0]  <= 1'b0;
    \\u26_cnt_reg[0]  <= 1'b0;
    \\u26_cnt_reg[1]  <= 1'b0;
    \\u13_crac_r_reg[6]  <= 1'b0;
    \\u13_occ0_r_reg[11]  <= 1'b0;
    \\u13_occ0_r_reg[8]  <= 1'b0;
    \\u13_icc_r_reg[8]  <= 1'b0;
    \\u13_icc_r_reg[22]  <= 1'b0;
    \\u13_occ0_r_reg[2]  <= 1'b0;
    \\u13_occ0_r_reg[4]  <= 1'b0;
    \\u13_intm_r_reg[7]  <= 1'b0;
    \\u13_intm_r_reg[22]  <= 1'b0;
    \\u13_icc_r_reg[11]  <= 1'b0;
    \\u13_icc_r_reg[15]  <= 1'b0;
    \\u13_icc_r_reg[19]  <= 1'b0;
    \\u13_crac_r_reg[0]  <= 1'b0;
    \\u13_crac_r_reg[1]  <= 1'b0;
    \\u13_crac_r_reg[3]  <= 1'b0;
    \\u13_crac_r_reg[4]  <= 1'b0;
    \\u13_crac_r_reg[5]  <= 1'b0;
    \\u13_crac_r_reg[7]  <= 1'b0;
    \\u13_icc_r_reg[0]  <= 1'b0;
    \\u13_icc_r_reg[10]  <= 1'b0;
    \\u13_icc_r_reg[12]  <= 1'b0;
    \\u13_icc_r_reg[13]  <= 1'b0;
    \\u13_icc_r_reg[14]  <= 1'b0;
    \\u13_icc_r_reg[16]  <= 1'b0;
    \\u13_icc_r_reg[17]  <= 1'b0;
    \\u13_icc_r_reg[18]  <= 1'b0;
    \\u13_icc_r_reg[1]  <= 1'b0;
    \\u13_icc_r_reg[20]  <= 1'b0;
    \\u13_icc_r_reg[21]  <= 1'b0;
    \\u13_icc_r_reg[23]  <= 1'b0;
    \\u13_icc_r_reg[2]  <= 1'b0;
    \\u13_icc_r_reg[3]  <= 1'b0;
    \\u13_icc_r_reg[4]  <= 1'b0;
    \\u13_icc_r_reg[5]  <= 1'b0;
    \\u13_icc_r_reg[6]  <= 1'b0;
    \\u13_icc_r_reg[7]  <= 1'b0;
    \\u13_icc_r_reg[9]  <= 1'b0;
    \\u13_occ0_r_reg[0]  <= 1'b0;
    \\u13_occ0_r_reg[10]  <= 1'b0;
    \\u13_occ0_r_reg[12]  <= 1'b0;
    \\u13_occ0_r_reg[13]  <= 1'b0;
    \\u13_occ0_r_reg[14]  <= 1'b0;
    \\u13_occ0_r_reg[16]  <= 1'b0;
    \\u13_occ0_r_reg[17]  <= 1'b0;
    \\u13_occ0_r_reg[18]  <= 1'b0;
    \\u13_occ0_r_reg[1]  <= 1'b0;
    \\u13_occ0_r_reg[20]  <= 1'b0;
    \\u13_occ0_r_reg[21]  <= 1'b0;
    \\u13_occ0_r_reg[23]  <= 1'b0;
    \\u13_occ0_r_reg[24]  <= 1'b0;
    \\u13_occ0_r_reg[25]  <= 1'b0;
    \\u13_occ0_r_reg[27]  <= 1'b0;
    \\u13_occ0_r_reg[28]  <= 1'b0;
    \\u13_occ0_r_reg[29]  <= 1'b0;
    \\u13_occ0_r_reg[30]  <= 1'b0;
    \\u13_occ0_r_reg[31]  <= 1'b0;
    \\u13_occ0_r_reg[3]  <= 1'b0;
    \\u13_occ0_r_reg[5]  <= 1'b0;
    \\u13_occ0_r_reg[6]  <= 1'b0;
    \\u13_occ0_r_reg[7]  <= 1'b0;
    \\u13_occ0_r_reg[9]  <= 1'b0;
    \\u13_intm_r_reg[0]  <= 1'b0;
    \\u13_intm_r_reg[10]  <= 1'b0;
    \\u13_intm_r_reg[11]  <= 1'b0;
    \\u13_intm_r_reg[12]  <= 1'b0;
    \\u13_intm_r_reg[13]  <= 1'b0;
    \\u13_intm_r_reg[14]  <= 1'b0;
    \\u13_intm_r_reg[16]  <= 1'b0;
    \\u13_intm_r_reg[17]  <= 1'b0;
    \\u13_intm_r_reg[18]  <= 1'b0;
    \\u13_intm_r_reg[19]  <= 1'b0;
    \\u13_intm_r_reg[1]  <= 1'b0;
    \\u13_intm_r_reg[20]  <= 1'b0;
    \\u13_intm_r_reg[21]  <= 1'b0;
    \\u13_intm_r_reg[23]  <= 1'b0;
    \\u13_intm_r_reg[24]  <= 1'b0;
    \\u13_intm_r_reg[25]  <= 1'b0;
    \\u13_intm_r_reg[27]  <= 1'b0;
    \\u13_intm_r_reg[28]  <= 1'b0;
    \\u13_intm_r_reg[2]  <= 1'b0;
    \\u13_intm_r_reg[5]  <= 1'b0;
    \\u13_intm_r_reg[6]  <= 1'b0;
    \\u13_intm_r_reg[9]  <= 1'b0;
    \\u13_intm_r_reg[4]  <= 1'b0;
    \\u13_intm_r_reg[15]  <= 1'b0;
    \\u13_intm_r_reg[8]  <= 1'b0;
    \\u13_intm_r_reg[26]  <= 1'b0;
    \\u13_occ0_r_reg[22]  <= 1'b0;
    \\u13_crac_r_reg[2]  <= 1'b0;
    \\u13_occ0_r_reg[26]  <= 1'b0;
    \\u13_intm_r_reg[3]  <= 1'b0;
    \\u13_occ0_r_reg[19]  <= 1'b0;
    \\u13_occ0_r_reg[15]  <= 1'b0;
    \\u13_occ1_r_reg[11]  <= 1'b0;
    \\u13_occ1_r_reg[8]  <= 1'b0;
    \\u13_occ1_r_reg[0]  <= 1'b0;
    \\u13_occ1_r_reg[10]  <= 1'b0;
    \\u13_occ1_r_reg[12]  <= 1'b0;
    \\u13_occ1_r_reg[13]  <= 1'b0;
    \\u13_occ1_r_reg[14]  <= 1'b0;
    \\u13_occ1_r_reg[1]  <= 1'b0;
    \\u13_occ1_r_reg[2]  <= 1'b0;
    \\u13_occ1_r_reg[3]  <= 1'b0;
    \\u13_occ1_r_reg[5]  <= 1'b0;
    \\u13_occ1_r_reg[6]  <= 1'b0;
    \\u13_occ1_r_reg[7]  <= 1'b0;
    \\u13_occ1_r_reg[9]  <= 1'b0;
    \\u13_occ1_r_reg[15]  <= 1'b0;
    \\u13_occ1_r_reg[4]  <= 1'b0;
    \\u23_int_set_reg[1]  <= 1'b0;
    \\u24_int_set_reg[1]  <= 1'b0;
    \\u25_int_set_reg[1]  <= 1'b0;
    \\u2_to_cnt_reg[5]  <= 1'b0;
    \\u13_ints_r_reg[21]  <= 1'b0;
    \\u13_ints_r_reg[0]  <= 1'b0;
    \\u13_ints_r_reg[27]  <= 1'b0;
    \\u13_ints_r_reg[15]  <= 1'b0;
    \\u2_cnt_reg[7]  <= 1'b1;
    \\u2_to_cnt_reg[3]  <= 1'b0;
    \\u2_to_cnt_reg[4]  <= 1'b0;
    \\u13_ints_r_reg[10]  <= 1'b0;
    \\u13_ints_r_reg[12]  <= 1'b0;
    \\u13_ints_r_reg[13]  <= 1'b0;
    \\u13_ints_r_reg[16]  <= 1'b0;
    \\u13_ints_r_reg[18]  <= 1'b0;
    \\u13_ints_r_reg[19]  <= 1'b0;
    \\u13_ints_r_reg[22]  <= 1'b0;
    \\u13_ints_r_reg[24]  <= 1'b0;
    \\u13_ints_r_reg[25]  <= 1'b0;
    \\u13_ints_r_reg[28]  <= 1'b0;
    \\u13_ints_r_reg[3]  <= 1'b0;
    \\u13_ints_r_reg[4]  <= 1'b0;
    \\u13_ints_r_reg[7]  <= 1'b0;
    \\u13_ints_r_reg[6]  <= 1'b0;
    \\u13_ints_r_reg[9]  <= 1'b0;
    \\u2_cnt_reg[1]  <= 1'b1;
    \\u2_to_cnt_reg[2]  <= 1'b0;
    \\u2_cnt_reg[4]  <= 1'b1;
    \\u2_cnt_reg[3]  <= 1'b1;
    \\u2_to_cnt_reg[0]  <= 1'b0;
    \\u2_to_cnt_reg[1]  <= 1'b0;
    \\u2_cnt_reg[5]  <= 1'b1;
    \\u2_cnt_reg[6]  <= 1'b1;
    \\u2_cnt_reg[0]  <= 1'b1;
    \\u2_cnt_reg[2]  <= 1'b1;
    \\u15_crac_din_reg[6]  <= 1'b0;
    \\u15_crac_din_reg[9]  <= 1'b0;
    \\u15_crac_din_reg[12]  <= 1'b0;
    \\u15_crac_din_reg[1]  <= 1'b0;
    \\u15_crac_din_reg[7]  <= 1'b0;
    \\u15_crac_din_reg[14]  <= 1'b0;
    \\u15_crac_din_reg[10]  <= 1'b0;
    \\u15_crac_din_reg[15]  <= 1'b0;
    \\u15_crac_din_reg[4]  <= 1'b0;
    \\u15_crac_din_reg[8]  <= 1'b0;
    \\u15_crac_din_reg[11]  <= 1'b0;
    \\u15_crac_din_reg[13]  <= 1'b0;
    \\u15_crac_din_reg[2]  <= 1'b0;
    \\u15_crac_din_reg[0]  <= 1'b0;
    \\u15_crac_din_reg[5]  <= 1'b0;
    \\u15_crac_din_reg[3]  <= 1'b0;
  end
endmodule


