module top ( 
    pv47_3_, pv84_15_, pv84_26_, pv116_20_, pv133_10_, pv15_9_, pv15_14_,
    pv47_4_, pv84_16_, pv84_25_, pv116_9_, pv116_21_, pv119_0_, pv15_13_,
    pv47_5_, pv84_13_, pv84_24_, pv15_12_, pv47_6_, pv84_14_, pv84_23_,
    pv15_6_, pv47_7_, pv47_18_, pv47_29_, pv84_6_, pv84_19_, pv116_6_,
    pv116_11_, pv118_0_, pv15_5_, pv47_8_, pv47_17_, pv84_7_, pv84_29_,
    pv116_5_, pv116_10_, pv15_8_, pv47_9_, pv47_27_, pv84_8_, pv84_17_,
    pv84_28_, pv116_8_, pv15_7_, pv47_19_, pv47_28_, pv84_9_, pv84_18_,
    pv84_27_, pv116_7_, pv118_1_, pv47_14_, pv47_25_, pv116_15_, pv116_28_,
    pv47_13_, pv47_26_, pv84_30_, pv116_14_, pv116_29_, pv122_0_, pv47_16_,
    pv47_23_, pv84_31_, pv116_13_, pv116_26_, pv47_15_, pv47_24_,
    pv116_12_, pv116_27_, pv15_11_, pv47_10_, pv47_21_, pv84_11_, pv84_22_,
    pv116_19_, pv116_24_, pv15_10_, pv47_22_, pv47_31_, pv84_12_, pv84_21_,
    pv116_18_, pv116_25_, pv47_12_, pv47_30_, pv84_20_, pv116_17_,
    pv116_22_, pv116_31_, pv47_11_, pv47_20_, pv84_10_, pv116_16_,
    pv116_23_, pv116_30_, pv133_5_, pv52_0_, pv133_4_, pv133_3_, pv133_2_,
    pv133_1_, pv133_0_, pv15_2_, pv84_2_, pv116_2_, pv121_17_, pv15_1_,
    pv84_3_, pv116_1_, pv15_4_, pv84_4_, pv116_4_, pv15_3_, pv84_5_,
    pv116_3_, pv121_16_, pv133_9_, pv47_0_, pv133_8_, pv15_0_, pv47_1_,
    pv48_0_, pv51_0_, pv84_0_, pv116_0_, pv133_7_, pv47_2_, pv49_0_,
    pv50_0_, pv84_1_, pv133_6_,
    pv150_0_, pv197_21_, pv197_20_, pv197_10_, pv197_11_, pv212_9_,
    pv212_8_, pv142_0_, pv197_7_, pv197_6_, pv165_8_, pv197_9_, pv165_9_,
    pv197_8_, pv149_0_, pv197_3_, pv149_1_, pv197_2_, pv149_2_, pv197_5_,
    pv197_4_, pv145_0_, pv165_2_, pv212_14_, pv145_1_, pv165_3_, pv165_10_,
    pv134_0_, pv165_0_, pv197_1_, pv212_12_, pv146_0_, pv165_1_, pv197_0_,
    pv212_13_, pv165_6_, pv165_13_, pv165_7_, pv165_14_, pv165_4_,
    pv165_11_, pv165_5_, pv165_12_, pv142_1_, pv197_16_, pv197_29_,
    pv212_5_, pv142_2_, pv197_17_, pv197_28_, pv212_4_, pv142_3_, pv143_0_,
    pv197_18_, pv197_27_, pv212_7_, pv136_1_, pv142_4_, pv197_19_,
    pv197_26_, pv212_6_, pv214_0_, pv136_0_, pv142_5_, pv197_12_,
    pv197_25_, pv197_30_, pv212_1_, pv212_10_, pv197_13_, pv197_24_,
    pv197_31_, pv212_0_, pv212_11_, pv197_14_, pv197_23_, pv212_3_,
    pv213_0_, pv197_15_, pv197_22_, pv212_2_  );
  input  pv47_3_, pv84_15_, pv84_26_, pv116_20_, pv133_10_, pv15_9_,
    pv15_14_, pv47_4_, pv84_16_, pv84_25_, pv116_9_, pv116_21_, pv119_0_,
    pv15_13_, pv47_5_, pv84_13_, pv84_24_, pv15_12_, pv47_6_, pv84_14_,
    pv84_23_, pv15_6_, pv47_7_, pv47_18_, pv47_29_, pv84_6_, pv84_19_,
    pv116_6_, pv116_11_, pv118_0_, pv15_5_, pv47_8_, pv47_17_, pv84_7_,
    pv84_29_, pv116_5_, pv116_10_, pv15_8_, pv47_9_, pv47_27_, pv84_8_,
    pv84_17_, pv84_28_, pv116_8_, pv15_7_, pv47_19_, pv47_28_, pv84_9_,
    pv84_18_, pv84_27_, pv116_7_, pv118_1_, pv47_14_, pv47_25_, pv116_15_,
    pv116_28_, pv47_13_, pv47_26_, pv84_30_, pv116_14_, pv116_29_,
    pv122_0_, pv47_16_, pv47_23_, pv84_31_, pv116_13_, pv116_26_, pv47_15_,
    pv47_24_, pv116_12_, pv116_27_, pv15_11_, pv47_10_, pv47_21_, pv84_11_,
    pv84_22_, pv116_19_, pv116_24_, pv15_10_, pv47_22_, pv47_31_, pv84_12_,
    pv84_21_, pv116_18_, pv116_25_, pv47_12_, pv47_30_, pv84_20_,
    pv116_17_, pv116_22_, pv116_31_, pv47_11_, pv47_20_, pv84_10_,
    pv116_16_, pv116_23_, pv116_30_, pv133_5_, pv52_0_, pv133_4_, pv133_3_,
    pv133_2_, pv133_1_, pv133_0_, pv15_2_, pv84_2_, pv116_2_, pv121_17_,
    pv15_1_, pv84_3_, pv116_1_, pv15_4_, pv84_4_, pv116_4_, pv15_3_,
    pv84_5_, pv116_3_, pv121_16_, pv133_9_, pv47_0_, pv133_8_, pv15_0_,
    pv47_1_, pv48_0_, pv51_0_, pv84_0_, pv116_0_, pv133_7_, pv47_2_,
    pv49_0_, pv50_0_, pv84_1_, pv133_6_;
  output pv150_0_, pv197_21_, pv197_20_, pv197_10_, pv197_11_, pv212_9_,
    pv212_8_, pv142_0_, pv197_7_, pv197_6_, pv165_8_, pv197_9_, pv165_9_,
    pv197_8_, pv149_0_, pv197_3_, pv149_1_, pv197_2_, pv149_2_, pv197_5_,
    pv197_4_, pv145_0_, pv165_2_, pv212_14_, pv145_1_, pv165_3_, pv165_10_,
    pv134_0_, pv165_0_, pv197_1_, pv212_12_, pv146_0_, pv165_1_, pv197_0_,
    pv212_13_, pv165_6_, pv165_13_, pv165_7_, pv165_14_, pv165_4_,
    pv165_11_, pv165_5_, pv165_12_, pv142_1_, pv197_16_, pv197_29_,
    pv212_5_, pv142_2_, pv197_17_, pv197_28_, pv212_4_, pv142_3_, pv143_0_,
    pv197_18_, pv197_27_, pv212_7_, pv136_1_, pv142_4_, pv197_19_,
    pv197_26_, pv212_6_, pv214_0_, pv136_0_, pv142_5_, pv197_12_,
    pv197_25_, pv197_30_, pv212_1_, pv212_10_, pv197_13_, pv197_24_,
    pv197_31_, pv212_0_, pv212_11_, pv197_14_, pv197_23_, pv212_3_,
    pv213_0_, pv197_15_, pv197_22_, pv212_2_;
  wire new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_,
    new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n529_, new_n530_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_,
    new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_,
    new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1073_, new_n1074_, new_n1075_,
    new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_,
    new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_,
    new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_,
    new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_,
    new_n1100_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_,
    new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_,
    new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1421_, new_n1422_, new_n1423_,
    new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_,
    new_n1430_, new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_,
    new_n1436_, new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_,
    new_n1442_, new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_,
    new_n1448_, new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1595_, new_n1596_, new_n1597_,
    new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_,
    new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_,
    new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_,
    new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_,
    new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_,
    new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_,
    new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_,
    new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1769_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1809_, new_n1810_, new_n1811_, new_n1812_,
    new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_,
    new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_,
    new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_,
    new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_,
    new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_,
    new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_,
    new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_,
    new_n1855_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_,
    new_n1868_, new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_,
    new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_,
    new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_,
    new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_,
    new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_,
    new_n1924_, new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_,
    new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1936_, new_n1937_,
    new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_,
    new_n1944_, new_n1945_, new_n1947_, new_n1948_, new_n1949_, new_n1950_,
    new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_, new_n1956_,
    new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_, new_n1962_,
    new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_, new_n1968_,
    new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_, new_n1974_,
    new_n1976_, new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_,
    new_n1982_, new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_,
    new_n1988_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_, new_n2088_,
    new_n2089_, new_n2090_, new_n2091_, new_n2093_, new_n2094_, new_n2095_,
    new_n2096_, new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_,
    new_n2102_, new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_,
    new_n2108_, new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_,
    new_n2114_, new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_,
    new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_,
    new_n2145_, new_n2146_, new_n2148_, new_n2149_, new_n2150_, new_n2151_,
    new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_,
    new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_,
    new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_,
    new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_,
    new_n2183_, new_n2184_, new_n2186_, new_n2187_, new_n2188_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_,
    new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_,
    new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_,
    new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_,
    new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2251_, new_n2252_,
    new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_,
    new_n2259_, new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_,
    new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_,
    new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_,
    new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2284_,
    new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_,
    new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_,
    new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_,
    new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_,
    new_n2309_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2337_, new_n2338_, new_n2339_, new_n2340_,
    new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_;
  assign new_n215_ = ~pv133_4_ & ~pv133_1_;
  assign new_n216_ = ~pv133_2_ & new_n215_;
  assign new_n217_ = ~pv133_9_ & new_n216_;
  assign new_n218_ = ~pv133_4_ & ~pv133_6_;
  assign new_n219_ = ~pv133_2_ & new_n218_;
  assign new_n220_ = ~pv133_9_ & new_n219_;
  assign new_n221_ = ~pv133_4_ & pv133_3_;
  assign new_n222_ = ~pv133_9_ & new_n221_;
  assign new_n223_ = ~pv133_6_ & new_n215_;
  assign new_n224_ = ~pv133_9_ & new_n223_;
  assign new_n225_ = pv133_1_ & pv133_8_;
  assign new_n226_ = ~pv133_10_ & new_n225_;
  assign new_n227_ = ~pv133_5_ & ~pv133_0_;
  assign new_n228_ = ~pv133_10_ & new_n227_;
  assign new_n229_ = ~pv133_2_ & ~pv133_6_;
  assign new_n230_ = ~pv133_5_ & new_n229_;
  assign new_n231_ = pv133_1_ & new_n230_;
  assign new_n232_ = ~pv133_10_ & new_n231_;
  assign new_n233_ = ~pv133_0_ & pv133_7_;
  assign new_n234_ = ~pv133_10_ & new_n233_;
  assign new_n235_ = ~new_n226_ & ~new_n228_;
  assign new_n236_ = ~new_n232_ & ~new_n234_;
  assign new_n237_ = new_n235_ & new_n236_;
  assign new_n238_ = pv133_2_ & pv133_1_;
  assign new_n239_ = pv133_3_ & new_n238_;
  assign new_n240_ = ~pv133_10_ & ~new_n239_;
  assign new_n241_ = ~new_n237_ & new_n240_;
  assign new_n242_ = pv47_8_ & new_n241_;
  assign new_n243_ = pv47_16_ & ~new_n240_;
  assign new_n244_ = ~pv133_2_ & pv133_7_;
  assign new_n245_ = ~pv133_1_ & new_n244_;
  assign new_n246_ = ~pv133_10_ & new_n245_;
  assign new_n247_ = ~pv133_1_ & new_n230_;
  assign new_n248_ = ~pv133_10_ & new_n247_;
  assign new_n249_ = ~new_n246_ & ~new_n248_;
  assign new_n250_ = ~pv133_3_ & pv133_2_;
  assign new_n251_ = pv133_1_ & new_n250_;
  assign new_n252_ = ~pv133_10_ & new_n251_;
  assign new_n253_ = pv133_2_ & pv133_8_;
  assign new_n254_ = ~pv133_1_ & new_n253_;
  assign new_n255_ = ~pv133_10_ & new_n254_;
  assign new_n256_ = pv133_2_ & pv133_0_;
  assign new_n257_ = ~pv133_5_ & new_n256_;
  assign new_n258_ = ~pv133_1_ & new_n257_;
  assign new_n259_ = ~pv133_10_ & new_n258_;
  assign new_n260_ = ~pv133_6_ & new_n259_;
  assign new_n261_ = ~new_n252_ & ~new_n255_;
  assign new_n262_ = ~new_n260_ & new_n261_;
  assign new_n263_ = new_n237_ & ~new_n249_;
  assign new_n264_ = new_n262_ & new_n263_;
  assign new_n265_ = new_n240_ & new_n264_;
  assign new_n266_ = pv47_1_ & new_n265_;
  assign new_n267_ = new_n237_ & ~new_n262_;
  assign new_n268_ = new_n240_ & new_n267_;
  assign new_n269_ = pv47_5_ & new_n268_;
  assign new_n270_ = new_n237_ & new_n262_;
  assign new_n271_ = new_n240_ & new_n270_;
  assign new_n272_ = new_n249_ & new_n271_;
  assign new_n273_ = ~new_n269_ & ~new_n272_;
  assign new_n274_ = ~new_n242_ & ~new_n243_;
  assign new_n275_ = ~new_n266_ & new_n274_;
  assign new_n276_ = new_n273_ & new_n275_;
  assign new_n277_ = ~pv133_9_ & pv133_7_;
  assign new_n278_ = ~new_n217_ & ~new_n220_;
  assign new_n279_ = ~new_n222_ & new_n278_;
  assign new_n280_ = ~new_n224_ & new_n279_;
  assign new_n281_ = ~new_n276_ & new_n280_;
  assign new_n282_ = new_n277_ & new_n281_;
  assign new_n283_ = new_n222_ & ~new_n224_;
  assign new_n284_ = ~new_n220_ & new_n283_;
  assign new_n285_ = ~new_n217_ & new_n284_;
  assign new_n286_ = ~new_n276_ & new_n285_;
  assign new_n287_ = ~pv133_10_ & pv133_9_;
  assign new_n288_ = ~new_n217_ & ~new_n224_;
  assign new_n289_ = ~pv133_10_ & new_n288_;
  assign new_n290_ = ~new_n222_ & new_n289_;
  assign new_n291_ = pv116_16_ & new_n290_;
  assign new_n292_ = new_n287_ & new_n291_;
  assign new_n293_ = ~new_n220_ & new_n292_;
  assign new_n294_ = ~new_n277_ & new_n293_;
  assign new_n295_ = ~new_n277_ & new_n288_;
  assign new_n296_ = ~new_n220_ & new_n295_;
  assign new_n297_ = ~new_n276_ & new_n296_;
  assign new_n298_ = ~new_n222_ & new_n297_;
  assign new_n299_ = pv133_10_ & new_n298_;
  assign new_n300_ = new_n278_ & ~new_n287_;
  assign new_n301_ = ~new_n277_ & new_n300_;
  assign new_n302_ = pv84_16_ & new_n301_;
  assign new_n303_ = pv133_2_ & new_n302_;
  assign new_n304_ = pv133_1_ & new_n303_;
  assign new_n305_ = ~pv133_10_ & new_n304_;
  assign new_n306_ = ~pv133_4_ & new_n305_;
  assign new_n307_ = ~pv133_3_ & new_n306_;
  assign new_n308_ = ~pv133_9_ & new_n307_;
  assign new_n309_ = ~pv133_10_ & new_n308_;
  assign new_n310_ = ~pv133_7_ & new_n309_;
  assign new_n311_ = ~new_n224_ & new_n310_;
  assign new_n312_ = ~new_n222_ & new_n311_;
  assign new_n313_ = new_n217_ & ~new_n276_;
  assign new_n314_ = new_n220_ & ~new_n224_;
  assign new_n315_ = ~new_n217_ & new_n314_;
  assign new_n316_ = ~new_n276_ & new_n315_;
  assign new_n317_ = ~new_n217_ & new_n224_;
  assign new_n318_ = ~new_n276_ & new_n317_;
  assign new_n319_ = ~new_n282_ & ~new_n286_;
  assign new_n320_ = ~new_n294_ & ~new_n299_;
  assign new_n321_ = new_n319_ & new_n320_;
  assign new_n322_ = ~new_n312_ & ~new_n313_;
  assign new_n323_ = ~new_n316_ & ~new_n318_;
  assign new_n324_ = new_n322_ & new_n323_;
  assign pv150_0_ = ~new_n321_ | ~new_n324_;
  assign new_n326_ = pv133_5_ & ~pv133_9_;
  assign new_n327_ = ~pv133_1_ & new_n326_;
  assign new_n328_ = ~pv118_0_ & new_n327_;
  assign new_n329_ = pv133_0_ & new_n328_;
  assign new_n330_ = pv133_1_ & new_n221_;
  assign new_n331_ = pv133_2_ & new_n330_;
  assign new_n332_ = ~pv133_9_ & new_n331_;
  assign new_n333_ = ~pv133_6_ & new_n332_;
  assign new_n334_ = pv133_5_ & ~pv133_1_;
  assign new_n335_ = ~pv133_9_ & new_n334_;
  assign new_n336_ = ~pv133_0_ & new_n335_;
  assign new_n337_ = ~pv133_5_ & ~pv133_4_;
  assign new_n338_ = ~pv133_1_ & new_n337_;
  assign new_n339_ = ~pv133_6_ & new_n338_;
  assign new_n340_ = ~pv133_9_ & new_n339_;
  assign new_n341_ = pv84_13_ & new_n241_;
  assign new_n342_ = pv84_21_ & ~new_n240_;
  assign new_n343_ = pv84_6_ & new_n265_;
  assign new_n344_ = pv84_10_ & new_n268_;
  assign new_n345_ = ~new_n272_ & ~new_n344_;
  assign new_n346_ = ~new_n341_ & ~new_n342_;
  assign new_n347_ = ~new_n343_ & new_n346_;
  assign new_n348_ = new_n345_ & new_n347_;
  assign new_n349_ = ~new_n329_ & new_n333_;
  assign new_n350_ = ~new_n336_ & new_n349_;
  assign new_n351_ = ~new_n340_ & new_n350_;
  assign new_n352_ = ~new_n348_ & new_n351_;
  assign new_n353_ = ~new_n329_ & new_n336_;
  assign new_n354_ = ~new_n340_ & new_n353_;
  assign new_n355_ = ~new_n348_ & new_n354_;
  assign new_n356_ = ~pv133_1_ & pv133_7_;
  assign new_n357_ = ~pv133_9_ & new_n356_;
  assign new_n358_ = ~new_n329_ & ~new_n340_;
  assign new_n359_ = ~new_n357_ & new_n358_;
  assign new_n360_ = ~new_n336_ & new_n359_;
  assign new_n361_ = ~new_n348_ & new_n360_;
  assign new_n362_ = ~new_n333_ & new_n361_;
  assign new_n363_ = pv133_10_ & new_n362_;
  assign new_n364_ = ~new_n336_ & ~new_n340_;
  assign new_n365_ = ~new_n333_ & new_n364_;
  assign new_n366_ = ~new_n329_ & new_n365_;
  assign new_n367_ = ~new_n348_ & new_n366_;
  assign new_n368_ = new_n357_ & new_n367_;
  assign new_n369_ = ~pv133_10_ & new_n358_;
  assign new_n370_ = ~new_n333_ & new_n369_;
  assign new_n371_ = pv116_21_ & new_n370_;
  assign new_n372_ = pv133_9_ & new_n371_;
  assign new_n373_ = ~pv133_10_ & new_n372_;
  assign new_n374_ = ~new_n336_ & new_n373_;
  assign new_n375_ = ~new_n357_ & new_n374_;
  assign new_n376_ = new_n329_ & ~new_n340_;
  assign new_n377_ = ~new_n348_ & new_n376_;
  assign new_n378_ = new_n340_ & ~new_n348_;
  assign new_n379_ = ~new_n352_ & ~new_n355_;
  assign new_n380_ = ~new_n363_ & ~new_n368_;
  assign new_n381_ = new_n379_ & new_n380_;
  assign new_n382_ = ~new_n375_ & ~new_n377_;
  assign new_n383_ = ~new_n378_ & new_n382_;
  assign pv197_21_ = ~new_n381_ | ~new_n383_;
  assign new_n385_ = pv84_12_ & new_n241_;
  assign new_n386_ = pv84_20_ & ~new_n240_;
  assign new_n387_ = pv84_5_ & new_n265_;
  assign new_n388_ = pv84_9_ & new_n268_;
  assign new_n389_ = ~new_n272_ & ~new_n388_;
  assign new_n390_ = ~new_n385_ & ~new_n386_;
  assign new_n391_ = ~new_n387_ & new_n390_;
  assign new_n392_ = new_n389_ & new_n391_;
  assign new_n393_ = new_n351_ & ~new_n392_;
  assign new_n394_ = new_n354_ & ~new_n392_;
  assign new_n395_ = new_n360_ & ~new_n392_;
  assign new_n396_ = ~new_n333_ & new_n395_;
  assign new_n397_ = pv133_10_ & new_n396_;
  assign new_n398_ = new_n366_ & ~new_n392_;
  assign new_n399_ = new_n357_ & new_n398_;
  assign new_n400_ = pv116_20_ & new_n370_;
  assign new_n401_ = pv133_9_ & new_n400_;
  assign new_n402_ = ~pv133_10_ & new_n401_;
  assign new_n403_ = ~new_n336_ & new_n402_;
  assign new_n404_ = ~new_n357_ & new_n403_;
  assign new_n405_ = new_n376_ & ~new_n392_;
  assign new_n406_ = new_n340_ & ~new_n392_;
  assign new_n407_ = ~new_n393_ & ~new_n394_;
  assign new_n408_ = ~new_n397_ & ~new_n399_;
  assign new_n409_ = new_n407_ & new_n408_;
  assign new_n410_ = ~new_n404_ & ~new_n405_;
  assign new_n411_ = ~new_n406_ & new_n410_;
  assign pv197_20_ = ~new_n409_ | ~new_n411_;
  assign new_n413_ = pv84_2_ & new_n241_;
  assign new_n414_ = pv84_10_ & ~new_n240_;
  assign new_n415_ = pv47_27_ & new_n265_;
  assign new_n416_ = pv47_31_ & new_n268_;
  assign new_n417_ = ~new_n272_ & ~new_n416_;
  assign new_n418_ = ~new_n413_ & ~new_n414_;
  assign new_n419_ = ~new_n415_ & new_n418_;
  assign new_n420_ = new_n417_ & new_n419_;
  assign new_n421_ = new_n351_ & ~new_n420_;
  assign new_n422_ = new_n354_ & ~new_n420_;
  assign new_n423_ = new_n360_ & ~new_n420_;
  assign new_n424_ = ~new_n333_ & new_n423_;
  assign new_n425_ = pv133_10_ & new_n424_;
  assign new_n426_ = new_n366_ & ~new_n420_;
  assign new_n427_ = new_n357_ & new_n426_;
  assign new_n428_ = pv116_10_ & new_n370_;
  assign new_n429_ = pv133_9_ & new_n428_;
  assign new_n430_ = ~pv133_10_ & new_n429_;
  assign new_n431_ = ~new_n336_ & new_n430_;
  assign new_n432_ = ~new_n357_ & new_n431_;
  assign new_n433_ = new_n376_ & ~new_n420_;
  assign new_n434_ = new_n340_ & ~new_n420_;
  assign new_n435_ = ~new_n421_ & ~new_n422_;
  assign new_n436_ = ~new_n425_ & ~new_n427_;
  assign new_n437_ = new_n435_ & new_n436_;
  assign new_n438_ = ~new_n432_ & ~new_n433_;
  assign new_n439_ = ~new_n434_ & new_n438_;
  assign pv197_10_ = ~new_n437_ | ~new_n439_;
  assign new_n441_ = pv84_3_ & new_n241_;
  assign new_n442_ = pv84_11_ & ~new_n240_;
  assign new_n443_ = pv47_28_ & new_n265_;
  assign new_n444_ = pv84_0_ & new_n268_;
  assign new_n445_ = ~new_n272_ & ~new_n444_;
  assign new_n446_ = ~new_n441_ & ~new_n442_;
  assign new_n447_ = ~new_n443_ & new_n446_;
  assign new_n448_ = new_n445_ & new_n447_;
  assign new_n449_ = new_n351_ & ~new_n448_;
  assign new_n450_ = new_n354_ & ~new_n448_;
  assign new_n451_ = new_n360_ & ~new_n448_;
  assign new_n452_ = ~new_n333_ & new_n451_;
  assign new_n453_ = pv133_10_ & new_n452_;
  assign new_n454_ = new_n366_ & ~new_n448_;
  assign new_n455_ = new_n357_ & new_n454_;
  assign new_n456_ = pv116_11_ & new_n370_;
  assign new_n457_ = pv133_9_ & new_n456_;
  assign new_n458_ = ~pv133_10_ & new_n457_;
  assign new_n459_ = ~new_n336_ & new_n458_;
  assign new_n460_ = ~new_n357_ & new_n459_;
  assign new_n461_ = new_n376_ & ~new_n448_;
  assign new_n462_ = new_n340_ & ~new_n448_;
  assign new_n463_ = ~new_n449_ & ~new_n450_;
  assign new_n464_ = ~new_n453_ & ~new_n455_;
  assign new_n465_ = new_n463_ & new_n464_;
  assign new_n466_ = ~new_n460_ & ~new_n461_;
  assign new_n467_ = ~new_n462_ & new_n466_;
  assign pv197_11_ = ~new_n465_ | ~new_n467_;
  assign new_n469_ = ~pv133_2_ & new_n356_;
  assign new_n470_ = ~pv133_9_ & new_n469_;
  assign new_n471_ = ~pv133_1_ & new_n218_;
  assign new_n472_ = ~pv133_2_ & new_n471_;
  assign new_n473_ = ~pv133_9_ & new_n472_;
  assign new_n474_ = ~pv133_5_ & new_n473_;
  assign new_n475_ = new_n470_ & ~new_n474_;
  assign new_n476_ = pv84_26_ & new_n475_;
  assign new_n477_ = pv84_26_ & new_n474_;
  assign new_n478_ = ~pv133_10_ & ~pv118_0_;
  assign new_n479_ = ~pv133_1_ & new_n478_;
  assign new_n480_ = ~pv133_2_ & new_n479_;
  assign new_n481_ = ~pv118_1_ & new_n480_;
  assign new_n482_ = ~pv133_7_ & new_n481_;
  assign new_n483_ = pv133_5_ & new_n482_;
  assign new_n484_ = ~pv133_9_ & new_n483_;
  assign new_n485_ = ~pv133_10_ & ~new_n470_;
  assign new_n486_ = ~new_n474_ & new_n485_;
  assign new_n487_ = new_n484_ & new_n486_;
  assign new_n488_ = pv133_10_ & ~new_n470_;
  assign new_n489_ = ~new_n474_ & new_n488_;
  assign new_n490_ = pv84_26_ & new_n489_;
  assign new_n491_ = ~pv133_10_ & ~new_n474_;
  assign new_n492_ = ~new_n484_ & new_n491_;
  assign new_n493_ = ~new_n470_ & new_n492_;
  assign new_n494_ = pv116_9_ & new_n493_;
  assign new_n495_ = pv133_9_ & new_n494_;
  assign new_n496_ = ~pv133_10_ & new_n495_;
  assign new_n497_ = ~new_n490_ & ~new_n496_;
  assign new_n498_ = ~new_n476_ & ~new_n477_;
  assign new_n499_ = ~new_n487_ & new_n498_;
  assign pv212_9_ = ~new_n497_ | ~new_n499_;
  assign new_n501_ = pv84_25_ & new_n475_;
  assign new_n502_ = pv84_25_ & new_n474_;
  assign new_n503_ = pv84_25_ & new_n489_;
  assign new_n504_ = pv116_8_ & new_n493_;
  assign new_n505_ = pv133_9_ & new_n504_;
  assign new_n506_ = ~pv133_10_ & new_n505_;
  assign new_n507_ = ~new_n503_ & ~new_n506_;
  assign new_n508_ = ~new_n501_ & ~new_n502_;
  assign new_n509_ = ~new_n487_ & new_n508_;
  assign pv212_8_ = ~new_n507_ | ~new_n509_;
  assign new_n511_ = pv47_3_ & ~new_n240_;
  assign new_n512_ = pv84_3_ & new_n268_;
  assign new_n513_ = pv15_2_ & new_n265_;
  assign new_n514_ = ~new_n511_ & ~new_n512_;
  assign new_n515_ = ~new_n272_ & ~new_n513_;
  assign new_n516_ = new_n514_ & new_n515_;
  assign new_n517_ = ~pv133_9_ & new_n218_;
  assign new_n518_ = ~new_n516_ & new_n517_;
  assign new_n519_ = pv133_10_ & ~new_n277_;
  assign new_n520_ = ~new_n517_ & new_n519_;
  assign new_n521_ = ~new_n516_ & new_n520_;
  assign new_n522_ = new_n277_ & ~new_n517_;
  assign new_n523_ = ~new_n516_ & new_n522_;
  assign new_n524_ = pv133_9_ & ~new_n277_;
  assign new_n525_ = ~pv133_10_ & new_n524_;
  assign new_n526_ = ~new_n517_ & new_n525_;
  assign new_n527_ = pv116_3_ & new_n526_;
  assign new_n528_ = ~pv133_10_ & new_n527_;
  assign new_n529_ = ~new_n518_ & ~new_n521_;
  assign new_n530_ = ~new_n523_ & ~new_n528_;
  assign pv142_0_ = ~new_n529_ | ~new_n530_;
  assign new_n532_ = pv47_31_ & new_n241_;
  assign new_n533_ = pv84_7_ & ~new_n240_;
  assign new_n534_ = pv47_24_ & new_n265_;
  assign new_n535_ = pv47_28_ & new_n268_;
  assign new_n536_ = ~new_n272_ & ~new_n535_;
  assign new_n537_ = ~new_n532_ & ~new_n533_;
  assign new_n538_ = ~new_n534_ & new_n537_;
  assign new_n539_ = new_n536_ & new_n538_;
  assign new_n540_ = new_n351_ & ~new_n539_;
  assign new_n541_ = new_n354_ & ~new_n539_;
  assign new_n542_ = new_n360_ & ~new_n539_;
  assign new_n543_ = ~new_n333_ & new_n542_;
  assign new_n544_ = pv133_10_ & new_n543_;
  assign new_n545_ = new_n366_ & ~new_n539_;
  assign new_n546_ = new_n357_ & new_n545_;
  assign new_n547_ = pv116_7_ & new_n370_;
  assign new_n548_ = pv133_9_ & new_n547_;
  assign new_n549_ = ~pv133_10_ & new_n548_;
  assign new_n550_ = ~new_n336_ & new_n549_;
  assign new_n551_ = ~new_n357_ & new_n550_;
  assign new_n552_ = new_n376_ & ~new_n539_;
  assign new_n553_ = new_n340_ & ~new_n539_;
  assign new_n554_ = ~new_n540_ & ~new_n541_;
  assign new_n555_ = ~new_n544_ & ~new_n546_;
  assign new_n556_ = new_n554_ & new_n555_;
  assign new_n557_ = ~new_n551_ & ~new_n552_;
  assign new_n558_ = ~new_n553_ & new_n557_;
  assign pv197_7_ = ~new_n556_ | ~new_n558_;
  assign new_n560_ = pv47_30_ & new_n241_;
  assign new_n561_ = pv84_6_ & ~new_n240_;
  assign new_n562_ = pv47_23_ & new_n265_;
  assign new_n563_ = pv47_27_ & new_n268_;
  assign new_n564_ = ~new_n272_ & ~new_n563_;
  assign new_n565_ = ~new_n560_ & ~new_n561_;
  assign new_n566_ = ~new_n562_ & new_n565_;
  assign new_n567_ = new_n564_ & new_n566_;
  assign new_n568_ = new_n351_ & ~new_n567_;
  assign new_n569_ = new_n354_ & ~new_n567_;
  assign new_n570_ = new_n360_ & ~new_n567_;
  assign new_n571_ = ~new_n333_ & new_n570_;
  assign new_n572_ = pv133_10_ & new_n571_;
  assign new_n573_ = new_n366_ & ~new_n567_;
  assign new_n574_ = new_n357_ & new_n573_;
  assign new_n575_ = pv116_6_ & new_n370_;
  assign new_n576_ = pv133_9_ & new_n575_;
  assign new_n577_ = ~pv133_10_ & new_n576_;
  assign new_n578_ = ~new_n336_ & new_n577_;
  assign new_n579_ = ~new_n357_ & new_n578_;
  assign new_n580_ = new_n376_ & ~new_n567_;
  assign new_n581_ = new_n340_ & ~new_n567_;
  assign new_n582_ = ~new_n568_ & ~new_n569_;
  assign new_n583_ = ~new_n572_ & ~new_n574_;
  assign new_n584_ = new_n582_ & new_n583_;
  assign new_n585_ = ~new_n579_ & ~new_n580_;
  assign new_n586_ = ~new_n581_ & new_n585_;
  assign pv197_6_ = ~new_n584_ | ~new_n586_;
  assign new_n588_ = pv47_17_ & new_n241_;
  assign new_n589_ = pv47_25_ & ~new_n240_;
  assign new_n590_ = pv47_10_ & new_n265_;
  assign new_n591_ = pv47_14_ & new_n268_;
  assign new_n592_ = ~new_n272_ & ~new_n591_;
  assign new_n593_ = ~new_n588_ & ~new_n589_;
  assign new_n594_ = ~new_n590_ & new_n593_;
  assign new_n595_ = new_n592_ & new_n594_;
  assign new_n596_ = ~new_n220_ & new_n277_;
  assign new_n597_ = ~new_n222_ & new_n596_;
  assign new_n598_ = ~new_n224_ & new_n597_;
  assign new_n599_ = ~new_n595_ & new_n598_;
  assign new_n600_ = ~new_n220_ & new_n222_;
  assign new_n601_ = ~new_n224_ & new_n600_;
  assign new_n602_ = ~new_n595_ & new_n601_;
  assign new_n603_ = ~new_n220_ & ~new_n224_;
  assign new_n604_ = ~pv133_10_ & new_n603_;
  assign new_n605_ = ~new_n222_ & new_n604_;
  assign new_n606_ = pv116_25_ & new_n605_;
  assign new_n607_ = ~new_n277_ & new_n606_;
  assign new_n608_ = new_n287_ & new_n607_;
  assign new_n609_ = ~new_n222_ & ~new_n224_;
  assign new_n610_ = ~new_n277_ & new_n609_;
  assign new_n611_ = ~new_n220_ & new_n610_;
  assign new_n612_ = ~new_n595_ & new_n611_;
  assign new_n613_ = pv133_10_ & new_n612_;
  assign new_n614_ = ~new_n287_ & new_n603_;
  assign new_n615_ = ~new_n277_ & new_n614_;
  assign new_n616_ = pv84_25_ & new_n615_;
  assign new_n617_ = pv133_1_ & new_n616_;
  assign new_n618_ = ~pv133_10_ & new_n617_;
  assign new_n619_ = ~pv133_3_ & new_n618_;
  assign new_n620_ = pv133_2_ & new_n619_;
  assign new_n621_ = ~pv133_4_ & new_n620_;
  assign new_n622_ = ~pv133_7_ & new_n621_;
  assign new_n623_ = ~pv133_9_ & new_n622_;
  assign new_n624_ = ~new_n222_ & new_n623_;
  assign new_n625_ = ~pv133_10_ & new_n624_;
  assign new_n626_ = new_n314_ & ~new_n595_;
  assign new_n627_ = new_n224_ & ~new_n595_;
  assign new_n628_ = ~new_n599_ & ~new_n602_;
  assign new_n629_ = ~new_n608_ & ~new_n613_;
  assign new_n630_ = new_n628_ & new_n629_;
  assign new_n631_ = ~new_n625_ & ~new_n626_;
  assign new_n632_ = ~new_n627_ & new_n631_;
  assign pv165_8_ = ~new_n630_ | ~new_n632_;
  assign new_n634_ = pv84_1_ & new_n241_;
  assign new_n635_ = pv84_9_ & ~new_n240_;
  assign new_n636_ = pv47_26_ & new_n265_;
  assign new_n637_ = pv47_30_ & new_n268_;
  assign new_n638_ = ~new_n272_ & ~new_n637_;
  assign new_n639_ = ~new_n634_ & ~new_n635_;
  assign new_n640_ = ~new_n636_ & new_n639_;
  assign new_n641_ = new_n638_ & new_n640_;
  assign new_n642_ = new_n351_ & ~new_n641_;
  assign new_n643_ = new_n354_ & ~new_n641_;
  assign new_n644_ = new_n360_ & ~new_n641_;
  assign new_n645_ = ~new_n333_ & new_n644_;
  assign new_n646_ = pv133_10_ & new_n645_;
  assign new_n647_ = new_n366_ & ~new_n641_;
  assign new_n648_ = new_n357_ & new_n647_;
  assign new_n649_ = pv116_9_ & new_n370_;
  assign new_n650_ = pv133_9_ & new_n649_;
  assign new_n651_ = ~pv133_10_ & new_n650_;
  assign new_n652_ = ~new_n336_ & new_n651_;
  assign new_n653_ = ~new_n357_ & new_n652_;
  assign new_n654_ = new_n376_ & ~new_n641_;
  assign new_n655_ = new_n340_ & ~new_n641_;
  assign new_n656_ = ~new_n642_ & ~new_n643_;
  assign new_n657_ = ~new_n646_ & ~new_n648_;
  assign new_n658_ = new_n656_ & new_n657_;
  assign new_n659_ = ~new_n653_ & ~new_n654_;
  assign new_n660_ = ~new_n655_ & new_n659_;
  assign pv197_9_ = ~new_n658_ | ~new_n660_;
  assign new_n662_ = pv47_18_ & new_n241_;
  assign new_n663_ = pv47_26_ & ~new_n240_;
  assign new_n664_ = pv47_11_ & new_n265_;
  assign new_n665_ = pv47_15_ & new_n268_;
  assign new_n666_ = ~new_n272_ & ~new_n665_;
  assign new_n667_ = ~new_n662_ & ~new_n663_;
  assign new_n668_ = ~new_n664_ & new_n667_;
  assign new_n669_ = new_n666_ & new_n668_;
  assign new_n670_ = new_n598_ & ~new_n669_;
  assign new_n671_ = new_n601_ & ~new_n669_;
  assign new_n672_ = pv116_26_ & new_n605_;
  assign new_n673_ = ~new_n277_ & new_n672_;
  assign new_n674_ = new_n287_ & new_n673_;
  assign new_n675_ = new_n611_ & ~new_n669_;
  assign new_n676_ = pv133_10_ & new_n675_;
  assign new_n677_ = pv84_26_ & new_n615_;
  assign new_n678_ = pv133_1_ & new_n677_;
  assign new_n679_ = ~pv133_10_ & new_n678_;
  assign new_n680_ = ~pv133_3_ & new_n679_;
  assign new_n681_ = pv133_2_ & new_n680_;
  assign new_n682_ = ~pv133_4_ & new_n681_;
  assign new_n683_ = ~pv133_7_ & new_n682_;
  assign new_n684_ = ~pv133_9_ & new_n683_;
  assign new_n685_ = ~new_n222_ & new_n684_;
  assign new_n686_ = ~pv133_10_ & new_n685_;
  assign new_n687_ = new_n314_ & ~new_n669_;
  assign new_n688_ = new_n224_ & ~new_n669_;
  assign new_n689_ = ~new_n670_ & ~new_n671_;
  assign new_n690_ = ~new_n674_ & ~new_n676_;
  assign new_n691_ = new_n689_ & new_n690_;
  assign new_n692_ = ~new_n686_ & ~new_n687_;
  assign new_n693_ = ~new_n688_ & new_n692_;
  assign pv165_9_ = ~new_n691_ | ~new_n693_;
  assign new_n695_ = pv84_0_ & new_n241_;
  assign new_n696_ = pv84_8_ & ~new_n240_;
  assign new_n697_ = pv47_25_ & new_n265_;
  assign new_n698_ = pv47_29_ & new_n268_;
  assign new_n699_ = ~new_n272_ & ~new_n698_;
  assign new_n700_ = ~new_n695_ & ~new_n696_;
  assign new_n701_ = ~new_n697_ & new_n700_;
  assign new_n702_ = new_n699_ & new_n701_;
  assign new_n703_ = new_n351_ & ~new_n702_;
  assign new_n704_ = new_n354_ & ~new_n702_;
  assign new_n705_ = new_n360_ & ~new_n702_;
  assign new_n706_ = ~new_n333_ & new_n705_;
  assign new_n707_ = pv133_10_ & new_n706_;
  assign new_n708_ = new_n366_ & ~new_n702_;
  assign new_n709_ = new_n357_ & new_n708_;
  assign new_n710_ = pv116_8_ & new_n370_;
  assign new_n711_ = pv133_9_ & new_n710_;
  assign new_n712_ = ~pv133_10_ & new_n711_;
  assign new_n713_ = ~new_n336_ & new_n712_;
  assign new_n714_ = ~new_n357_ & new_n713_;
  assign new_n715_ = new_n376_ & ~new_n702_;
  assign new_n716_ = new_n340_ & ~new_n702_;
  assign new_n717_ = ~new_n703_ & ~new_n704_;
  assign new_n718_ = ~new_n707_ & ~new_n709_;
  assign new_n719_ = new_n717_ & new_n718_;
  assign new_n720_ = ~new_n714_ & ~new_n715_;
  assign new_n721_ = ~new_n716_ & new_n720_;
  assign pv197_8_ = ~new_n719_ | ~new_n721_;
  assign new_n723_ = pv47_5_ & new_n241_;
  assign new_n724_ = pv47_13_ & ~new_n240_;
  assign new_n725_ = pv15_12_ & new_n265_;
  assign new_n726_ = pv47_2_ & new_n268_;
  assign new_n727_ = ~new_n272_ & ~new_n726_;
  assign new_n728_ = ~new_n723_ & ~new_n724_;
  assign new_n729_ = ~new_n725_ & new_n728_;
  assign new_n730_ = new_n727_ & new_n729_;
  assign new_n731_ = new_n598_ & ~new_n730_;
  assign new_n732_ = new_n601_ & ~new_n730_;
  assign new_n733_ = pv116_13_ & new_n605_;
  assign new_n734_ = ~new_n277_ & new_n733_;
  assign new_n735_ = new_n287_ & new_n734_;
  assign new_n736_ = new_n611_ & ~new_n730_;
  assign new_n737_ = pv133_10_ & new_n736_;
  assign new_n738_ = pv84_13_ & new_n615_;
  assign new_n739_ = pv133_1_ & new_n738_;
  assign new_n740_ = ~pv133_10_ & new_n739_;
  assign new_n741_ = ~pv133_3_ & new_n740_;
  assign new_n742_ = pv133_2_ & new_n741_;
  assign new_n743_ = ~pv133_4_ & new_n742_;
  assign new_n744_ = ~pv133_7_ & new_n743_;
  assign new_n745_ = ~pv133_9_ & new_n744_;
  assign new_n746_ = ~new_n222_ & new_n745_;
  assign new_n747_ = ~pv133_10_ & new_n746_;
  assign new_n748_ = new_n314_ & ~new_n730_;
  assign new_n749_ = new_n224_ & ~new_n730_;
  assign new_n750_ = ~new_n731_ & ~new_n732_;
  assign new_n751_ = ~new_n735_ & ~new_n737_;
  assign new_n752_ = new_n750_ & new_n751_;
  assign new_n753_ = ~new_n747_ & ~new_n748_;
  assign new_n754_ = ~new_n749_ & new_n753_;
  assign pv149_0_ = ~new_n752_ | ~new_n754_;
  assign new_n756_ = pv47_27_ & new_n241_;
  assign new_n757_ = pv84_3_ & ~new_n240_;
  assign new_n758_ = pv47_20_ & new_n265_;
  assign new_n759_ = pv47_24_ & new_n268_;
  assign new_n760_ = ~new_n272_ & ~new_n759_;
  assign new_n761_ = ~new_n756_ & ~new_n757_;
  assign new_n762_ = ~new_n758_ & new_n761_;
  assign new_n763_ = new_n760_ & new_n762_;
  assign new_n764_ = new_n351_ & ~new_n763_;
  assign new_n765_ = new_n354_ & ~new_n763_;
  assign new_n766_ = new_n360_ & ~new_n763_;
  assign new_n767_ = ~new_n333_ & new_n766_;
  assign new_n768_ = pv133_10_ & new_n767_;
  assign new_n769_ = new_n366_ & ~new_n763_;
  assign new_n770_ = new_n357_ & new_n769_;
  assign new_n771_ = pv116_3_ & new_n370_;
  assign new_n772_ = pv133_9_ & new_n771_;
  assign new_n773_ = ~pv133_10_ & new_n772_;
  assign new_n774_ = ~new_n336_ & new_n773_;
  assign new_n775_ = ~new_n357_ & new_n774_;
  assign new_n776_ = new_n376_ & ~new_n763_;
  assign new_n777_ = new_n340_ & ~new_n763_;
  assign new_n778_ = ~new_n764_ & ~new_n765_;
  assign new_n779_ = ~new_n768_ & ~new_n770_;
  assign new_n780_ = new_n778_ & new_n779_;
  assign new_n781_ = ~new_n775_ & ~new_n776_;
  assign new_n782_ = ~new_n777_ & new_n781_;
  assign pv197_3_ = ~new_n780_ | ~new_n782_;
  assign new_n784_ = pv47_6_ & new_n241_;
  assign new_n785_ = pv47_14_ & ~new_n240_;
  assign new_n786_ = pv15_13_ & new_n265_;
  assign new_n787_ = pv47_3_ & new_n268_;
  assign new_n788_ = ~new_n272_ & ~new_n787_;
  assign new_n789_ = ~new_n784_ & ~new_n785_;
  assign new_n790_ = ~new_n786_ & new_n789_;
  assign new_n791_ = new_n788_ & new_n790_;
  assign new_n792_ = new_n598_ & ~new_n791_;
  assign new_n793_ = new_n601_ & ~new_n791_;
  assign new_n794_ = pv116_14_ & new_n605_;
  assign new_n795_ = ~new_n277_ & new_n794_;
  assign new_n796_ = new_n287_ & new_n795_;
  assign new_n797_ = new_n611_ & ~new_n791_;
  assign new_n798_ = pv133_10_ & new_n797_;
  assign new_n799_ = pv84_14_ & new_n615_;
  assign new_n800_ = pv133_1_ & new_n799_;
  assign new_n801_ = ~pv133_10_ & new_n800_;
  assign new_n802_ = ~pv133_3_ & new_n801_;
  assign new_n803_ = pv133_2_ & new_n802_;
  assign new_n804_ = ~pv133_4_ & new_n803_;
  assign new_n805_ = ~pv133_7_ & new_n804_;
  assign new_n806_ = ~pv133_9_ & new_n805_;
  assign new_n807_ = ~new_n222_ & new_n806_;
  assign new_n808_ = ~pv133_10_ & new_n807_;
  assign new_n809_ = new_n314_ & ~new_n791_;
  assign new_n810_ = new_n224_ & ~new_n791_;
  assign new_n811_ = ~new_n792_ & ~new_n793_;
  assign new_n812_ = ~new_n796_ & ~new_n798_;
  assign new_n813_ = new_n811_ & new_n812_;
  assign new_n814_ = ~new_n808_ & ~new_n809_;
  assign new_n815_ = ~new_n810_ & new_n814_;
  assign pv149_1_ = ~new_n813_ | ~new_n815_;
  assign new_n817_ = pv47_26_ & new_n241_;
  assign new_n818_ = pv84_2_ & ~new_n240_;
  assign new_n819_ = pv47_19_ & new_n265_;
  assign new_n820_ = pv47_23_ & new_n268_;
  assign new_n821_ = ~new_n272_ & ~new_n820_;
  assign new_n822_ = ~new_n817_ & ~new_n818_;
  assign new_n823_ = ~new_n819_ & new_n822_;
  assign new_n824_ = new_n821_ & new_n823_;
  assign new_n825_ = new_n351_ & ~new_n824_;
  assign new_n826_ = new_n354_ & ~new_n824_;
  assign new_n827_ = new_n360_ & ~new_n824_;
  assign new_n828_ = ~new_n333_ & new_n827_;
  assign new_n829_ = pv133_10_ & new_n828_;
  assign new_n830_ = new_n366_ & ~new_n824_;
  assign new_n831_ = new_n357_ & new_n830_;
  assign new_n832_ = pv116_2_ & new_n370_;
  assign new_n833_ = pv133_9_ & new_n832_;
  assign new_n834_ = ~pv133_10_ & new_n833_;
  assign new_n835_ = ~new_n336_ & new_n834_;
  assign new_n836_ = ~new_n357_ & new_n835_;
  assign new_n837_ = new_n376_ & ~new_n824_;
  assign new_n838_ = new_n340_ & ~new_n824_;
  assign new_n839_ = ~new_n825_ & ~new_n826_;
  assign new_n840_ = ~new_n829_ & ~new_n831_;
  assign new_n841_ = new_n839_ & new_n840_;
  assign new_n842_ = ~new_n836_ & ~new_n837_;
  assign new_n843_ = ~new_n838_ & new_n842_;
  assign pv197_2_ = ~new_n841_ | ~new_n843_;
  assign new_n845_ = pv47_7_ & new_n241_;
  assign new_n846_ = pv47_15_ & ~new_n240_;
  assign new_n847_ = pv15_14_ & new_n265_;
  assign new_n848_ = pv47_4_ & new_n268_;
  assign new_n849_ = ~new_n272_ & ~new_n848_;
  assign new_n850_ = ~new_n845_ & ~new_n846_;
  assign new_n851_ = ~new_n847_ & new_n850_;
  assign new_n852_ = new_n849_ & new_n851_;
  assign new_n853_ = new_n598_ & ~new_n852_;
  assign new_n854_ = new_n601_ & ~new_n852_;
  assign new_n855_ = pv116_15_ & new_n605_;
  assign new_n856_ = ~new_n277_ & new_n855_;
  assign new_n857_ = new_n287_ & new_n856_;
  assign new_n858_ = new_n611_ & ~new_n852_;
  assign new_n859_ = pv133_10_ & new_n858_;
  assign new_n860_ = pv84_15_ & new_n615_;
  assign new_n861_ = pv133_1_ & new_n860_;
  assign new_n862_ = ~pv133_10_ & new_n861_;
  assign new_n863_ = ~pv133_3_ & new_n862_;
  assign new_n864_ = pv133_2_ & new_n863_;
  assign new_n865_ = ~pv133_4_ & new_n864_;
  assign new_n866_ = ~pv133_7_ & new_n865_;
  assign new_n867_ = ~pv133_9_ & new_n866_;
  assign new_n868_ = ~new_n222_ & new_n867_;
  assign new_n869_ = ~pv133_10_ & new_n868_;
  assign new_n870_ = new_n314_ & ~new_n852_;
  assign new_n871_ = new_n224_ & ~new_n852_;
  assign new_n872_ = ~new_n853_ & ~new_n854_;
  assign new_n873_ = ~new_n857_ & ~new_n859_;
  assign new_n874_ = new_n872_ & new_n873_;
  assign new_n875_ = ~new_n869_ & ~new_n870_;
  assign new_n876_ = ~new_n871_ & new_n875_;
  assign pv149_2_ = ~new_n874_ | ~new_n876_;
  assign new_n878_ = pv47_29_ & new_n241_;
  assign new_n879_ = pv84_5_ & ~new_n240_;
  assign new_n880_ = pv47_22_ & new_n265_;
  assign new_n881_ = pv47_26_ & new_n268_;
  assign new_n882_ = ~new_n272_ & ~new_n881_;
  assign new_n883_ = ~new_n878_ & ~new_n879_;
  assign new_n884_ = ~new_n880_ & new_n883_;
  assign new_n885_ = new_n882_ & new_n884_;
  assign new_n886_ = new_n351_ & ~new_n885_;
  assign new_n887_ = new_n354_ & ~new_n885_;
  assign new_n888_ = new_n360_ & ~new_n885_;
  assign new_n889_ = ~new_n333_ & new_n888_;
  assign new_n890_ = pv133_10_ & new_n889_;
  assign new_n891_ = new_n366_ & ~new_n885_;
  assign new_n892_ = new_n357_ & new_n891_;
  assign new_n893_ = pv116_5_ & new_n370_;
  assign new_n894_ = pv133_9_ & new_n893_;
  assign new_n895_ = ~pv133_10_ & new_n894_;
  assign new_n896_ = ~new_n336_ & new_n895_;
  assign new_n897_ = ~new_n357_ & new_n896_;
  assign new_n898_ = new_n376_ & ~new_n885_;
  assign new_n899_ = new_n340_ & ~new_n885_;
  assign new_n900_ = ~new_n886_ & ~new_n887_;
  assign new_n901_ = ~new_n890_ & ~new_n892_;
  assign new_n902_ = new_n900_ & new_n901_;
  assign new_n903_ = ~new_n897_ & ~new_n898_;
  assign new_n904_ = ~new_n899_ & new_n903_;
  assign pv197_5_ = ~new_n902_ | ~new_n904_;
  assign new_n906_ = pv47_28_ & new_n241_;
  assign new_n907_ = pv84_4_ & ~new_n240_;
  assign new_n908_ = pv47_21_ & new_n265_;
  assign new_n909_ = pv47_25_ & new_n268_;
  assign new_n910_ = ~new_n272_ & ~new_n909_;
  assign new_n911_ = ~new_n906_ & ~new_n907_;
  assign new_n912_ = ~new_n908_ & new_n911_;
  assign new_n913_ = new_n910_ & new_n912_;
  assign new_n914_ = new_n351_ & ~new_n913_;
  assign new_n915_ = new_n354_ & ~new_n913_;
  assign new_n916_ = new_n360_ & ~new_n913_;
  assign new_n917_ = ~new_n333_ & new_n916_;
  assign new_n918_ = pv133_10_ & new_n917_;
  assign new_n919_ = new_n366_ & ~new_n913_;
  assign new_n920_ = new_n357_ & new_n919_;
  assign new_n921_ = pv116_4_ & new_n370_;
  assign new_n922_ = pv133_9_ & new_n921_;
  assign new_n923_ = ~pv133_10_ & new_n922_;
  assign new_n924_ = ~new_n336_ & new_n923_;
  assign new_n925_ = ~new_n357_ & new_n924_;
  assign new_n926_ = new_n376_ & ~new_n913_;
  assign new_n927_ = new_n340_ & ~new_n913_;
  assign new_n928_ = ~new_n914_ & ~new_n915_;
  assign new_n929_ = ~new_n918_ & ~new_n920_;
  assign new_n930_ = new_n928_ & new_n929_;
  assign new_n931_ = ~new_n925_ & ~new_n926_;
  assign new_n932_ = ~new_n927_ & new_n931_;
  assign pv197_4_ = ~new_n930_ | ~new_n932_;
  assign new_n934_ = pv47_2_ & new_n241_;
  assign new_n935_ = pv47_10_ & ~new_n240_;
  assign new_n936_ = pv15_9_ & new_n265_;
  assign new_n937_ = ~new_n934_ & ~new_n935_;
  assign new_n938_ = ~new_n936_ & new_n937_;
  assign new_n939_ = new_n345_ & new_n938_;
  assign new_n940_ = new_n517_ & ~new_n939_;
  assign new_n941_ = new_n520_ & ~new_n939_;
  assign new_n942_ = new_n522_ & ~new_n939_;
  assign new_n943_ = pv116_10_ & new_n526_;
  assign new_n944_ = ~pv133_10_ & new_n943_;
  assign new_n945_ = ~new_n940_ & ~new_n941_;
  assign new_n946_ = ~new_n942_ & ~new_n944_;
  assign pv145_0_ = ~new_n945_ | ~new_n946_;
  assign new_n948_ = pv47_11_ & new_n241_;
  assign new_n949_ = pv47_19_ & ~new_n240_;
  assign new_n950_ = pv47_4_ & new_n265_;
  assign new_n951_ = pv47_8_ & new_n268_;
  assign new_n952_ = ~new_n272_ & ~new_n951_;
  assign new_n953_ = ~new_n948_ & ~new_n949_;
  assign new_n954_ = ~new_n950_ & new_n953_;
  assign new_n955_ = new_n952_ & new_n954_;
  assign new_n956_ = new_n598_ & ~new_n955_;
  assign new_n957_ = new_n601_ & ~new_n955_;
  assign new_n958_ = pv116_19_ & new_n605_;
  assign new_n959_ = ~new_n277_ & new_n958_;
  assign new_n960_ = new_n287_ & new_n959_;
  assign new_n961_ = new_n611_ & ~new_n955_;
  assign new_n962_ = pv133_10_ & new_n961_;
  assign new_n963_ = pv84_19_ & new_n615_;
  assign new_n964_ = pv133_1_ & new_n963_;
  assign new_n965_ = ~pv133_10_ & new_n964_;
  assign new_n966_ = ~pv133_3_ & new_n965_;
  assign new_n967_ = pv133_2_ & new_n966_;
  assign new_n968_ = ~pv133_4_ & new_n967_;
  assign new_n969_ = ~pv133_7_ & new_n968_;
  assign new_n970_ = ~pv133_9_ & new_n969_;
  assign new_n971_ = ~new_n222_ & new_n970_;
  assign new_n972_ = ~pv133_10_ & new_n971_;
  assign new_n973_ = new_n314_ & ~new_n955_;
  assign new_n974_ = new_n224_ & ~new_n955_;
  assign new_n975_ = ~new_n956_ & ~new_n957_;
  assign new_n976_ = ~new_n960_ & ~new_n962_;
  assign new_n977_ = new_n975_ & new_n976_;
  assign new_n978_ = ~new_n972_ & ~new_n973_;
  assign new_n979_ = ~new_n974_ & new_n978_;
  assign pv165_2_ = ~new_n977_ | ~new_n979_;
  assign new_n981_ = pv84_31_ & new_n475_;
  assign new_n982_ = pv84_31_ & new_n474_;
  assign new_n983_ = pv84_31_ & new_n489_;
  assign new_n984_ = pv116_14_ & new_n493_;
  assign new_n985_ = pv133_9_ & new_n984_;
  assign new_n986_ = ~pv133_10_ & new_n985_;
  assign new_n987_ = ~new_n983_ & ~new_n986_;
  assign new_n988_ = ~new_n981_ & ~new_n982_;
  assign new_n989_ = ~new_n487_ & new_n988_;
  assign pv212_14_ = ~new_n987_ | ~new_n989_;
  assign new_n991_ = pv47_3_ & new_n241_;
  assign new_n992_ = pv47_11_ & ~new_n240_;
  assign new_n993_ = pv15_10_ & new_n265_;
  assign new_n994_ = pv84_11_ & new_n268_;
  assign new_n995_ = ~new_n272_ & ~new_n994_;
  assign new_n996_ = ~new_n991_ & ~new_n992_;
  assign new_n997_ = ~new_n993_ & new_n996_;
  assign new_n998_ = new_n995_ & new_n997_;
  assign new_n999_ = new_n517_ & ~new_n998_;
  assign new_n1000_ = new_n520_ & ~new_n998_;
  assign new_n1001_ = new_n522_ & ~new_n998_;
  assign new_n1002_ = pv116_11_ & new_n526_;
  assign new_n1003_ = ~pv133_10_ & new_n1002_;
  assign new_n1004_ = ~new_n999_ & ~new_n1000_;
  assign new_n1005_ = ~new_n1001_ & ~new_n1003_;
  assign pv145_1_ = ~new_n1004_ | ~new_n1005_;
  assign new_n1007_ = pv47_12_ & new_n241_;
  assign new_n1008_ = pv47_20_ & ~new_n240_;
  assign new_n1009_ = pv47_5_ & new_n265_;
  assign new_n1010_ = pv47_9_ & new_n268_;
  assign new_n1011_ = ~new_n272_ & ~new_n1010_;
  assign new_n1012_ = ~new_n1007_ & ~new_n1008_;
  assign new_n1013_ = ~new_n1009_ & new_n1012_;
  assign new_n1014_ = new_n1011_ & new_n1013_;
  assign new_n1015_ = new_n598_ & ~new_n1014_;
  assign new_n1016_ = new_n601_ & ~new_n1014_;
  assign new_n1017_ = pv116_20_ & new_n605_;
  assign new_n1018_ = ~new_n277_ & new_n1017_;
  assign new_n1019_ = new_n287_ & new_n1018_;
  assign new_n1020_ = new_n611_ & ~new_n1014_;
  assign new_n1021_ = pv133_10_ & new_n1020_;
  assign new_n1022_ = pv84_20_ & new_n615_;
  assign new_n1023_ = pv133_1_ & new_n1022_;
  assign new_n1024_ = ~pv133_10_ & new_n1023_;
  assign new_n1025_ = ~pv133_3_ & new_n1024_;
  assign new_n1026_ = pv133_2_ & new_n1025_;
  assign new_n1027_ = ~pv133_4_ & new_n1026_;
  assign new_n1028_ = ~pv133_7_ & new_n1027_;
  assign new_n1029_ = ~pv133_9_ & new_n1028_;
  assign new_n1030_ = ~new_n222_ & new_n1029_;
  assign new_n1031_ = ~pv133_10_ & new_n1030_;
  assign new_n1032_ = new_n314_ & ~new_n1014_;
  assign new_n1033_ = new_n224_ & ~new_n1014_;
  assign new_n1034_ = ~new_n1015_ & ~new_n1016_;
  assign new_n1035_ = ~new_n1019_ & ~new_n1021_;
  assign new_n1036_ = new_n1034_ & new_n1035_;
  assign new_n1037_ = ~new_n1031_ & ~new_n1032_;
  assign new_n1038_ = ~new_n1033_ & new_n1037_;
  assign pv165_3_ = ~new_n1036_ | ~new_n1038_;
  assign new_n1040_ = pv47_19_ & new_n241_;
  assign new_n1041_ = pv47_27_ & ~new_n240_;
  assign new_n1042_ = pv47_12_ & new_n265_;
  assign new_n1043_ = pv47_16_ & new_n268_;
  assign new_n1044_ = ~new_n272_ & ~new_n1043_;
  assign new_n1045_ = ~new_n1040_ & ~new_n1041_;
  assign new_n1046_ = ~new_n1042_ & new_n1045_;
  assign new_n1047_ = new_n1044_ & new_n1046_;
  assign new_n1048_ = new_n598_ & ~new_n1047_;
  assign new_n1049_ = new_n601_ & ~new_n1047_;
  assign new_n1050_ = pv116_27_ & new_n605_;
  assign new_n1051_ = ~new_n277_ & new_n1050_;
  assign new_n1052_ = new_n287_ & new_n1051_;
  assign new_n1053_ = new_n611_ & ~new_n1047_;
  assign new_n1054_ = pv133_10_ & new_n1053_;
  assign new_n1055_ = pv84_27_ & new_n615_;
  assign new_n1056_ = pv133_1_ & new_n1055_;
  assign new_n1057_ = ~pv133_10_ & new_n1056_;
  assign new_n1058_ = ~pv133_3_ & new_n1057_;
  assign new_n1059_ = pv133_2_ & new_n1058_;
  assign new_n1060_ = ~pv133_4_ & new_n1059_;
  assign new_n1061_ = ~pv133_7_ & new_n1060_;
  assign new_n1062_ = ~pv133_9_ & new_n1061_;
  assign new_n1063_ = ~new_n222_ & new_n1062_;
  assign new_n1064_ = ~pv133_10_ & new_n1063_;
  assign new_n1065_ = new_n314_ & ~new_n1047_;
  assign new_n1066_ = new_n224_ & ~new_n1047_;
  assign new_n1067_ = ~new_n1048_ & ~new_n1049_;
  assign new_n1068_ = ~new_n1052_ & ~new_n1054_;
  assign new_n1069_ = new_n1067_ & new_n1068_;
  assign new_n1070_ = ~new_n1064_ & ~new_n1065_;
  assign new_n1071_ = ~new_n1066_ & new_n1070_;
  assign pv165_10_ = ~new_n1069_ | ~new_n1071_;
  assign new_n1073_ = ~pv133_9_ & ~pv133_7_;
  assign new_n1074_ = ~pv133_10_ & new_n1073_;
  assign new_n1075_ = ~pv133_2_ & new_n277_;
  assign new_n1076_ = ~pv133_10_ & new_n1075_;
  assign new_n1077_ = ~pv133_10_ & new_n357_;
  assign new_n1078_ = new_n1074_ & ~new_n1076_;
  assign new_n1079_ = ~new_n1077_ & new_n1078_;
  assign new_n1080_ = pv49_0_ & new_n1079_;
  assign new_n1081_ = new_n1076_ & ~new_n1077_;
  assign new_n1082_ = pv48_0_ & new_n1081_;
  assign new_n1083_ = ~new_n1074_ & ~new_n1077_;
  assign new_n1084_ = ~new_n287_ & new_n1083_;
  assign new_n1085_ = ~new_n1076_ & new_n1084_;
  assign new_n1086_ = pv84_0_ & new_n1085_;
  assign new_n1087_ = pv133_10_ & new_n1086_;
  assign new_n1088_ = new_n287_ & ~new_n1076_;
  assign new_n1089_ = ~new_n1074_ & new_n1088_;
  assign new_n1090_ = ~new_n1077_ & new_n1089_;
  assign new_n1091_ = pv116_0_ & new_n1090_;
  assign new_n1092_ = ~new_n287_ & ~new_n1076_;
  assign new_n1093_ = ~new_n1074_ & new_n1092_;
  assign new_n1094_ = ~new_n1077_ & new_n1093_;
  assign new_n1095_ = ~pv133_10_ & new_n1094_;
  assign new_n1096_ = pv48_0_ & new_n1077_;
  assign new_n1097_ = ~new_n1080_ & ~new_n1082_;
  assign new_n1098_ = ~new_n1087_ & new_n1097_;
  assign new_n1099_ = ~new_n1091_ & ~new_n1095_;
  assign new_n1100_ = ~new_n1096_ & new_n1099_;
  assign pv134_0_ = ~new_n1098_ | ~new_n1100_;
  assign new_n1102_ = pv47_9_ & new_n241_;
  assign new_n1103_ = pv47_17_ & ~new_n240_;
  assign new_n1104_ = pv47_2_ & new_n265_;
  assign new_n1105_ = pv47_6_ & new_n268_;
  assign new_n1106_ = ~new_n272_ & ~new_n1105_;
  assign new_n1107_ = ~new_n1102_ & ~new_n1103_;
  assign new_n1108_ = ~new_n1104_ & new_n1107_;
  assign new_n1109_ = new_n1106_ & new_n1108_;
  assign new_n1110_ = new_n598_ & ~new_n1109_;
  assign new_n1111_ = new_n601_ & ~new_n1109_;
  assign new_n1112_ = pv116_17_ & new_n605_;
  assign new_n1113_ = ~new_n277_ & new_n1112_;
  assign new_n1114_ = new_n287_ & new_n1113_;
  assign new_n1115_ = new_n611_ & ~new_n1109_;
  assign new_n1116_ = pv133_10_ & new_n1115_;
  assign new_n1117_ = pv84_17_ & new_n615_;
  assign new_n1118_ = pv133_1_ & new_n1117_;
  assign new_n1119_ = ~pv133_10_ & new_n1118_;
  assign new_n1120_ = ~pv133_3_ & new_n1119_;
  assign new_n1121_ = pv133_2_ & new_n1120_;
  assign new_n1122_ = ~pv133_4_ & new_n1121_;
  assign new_n1123_ = ~pv133_7_ & new_n1122_;
  assign new_n1124_ = ~pv133_9_ & new_n1123_;
  assign new_n1125_ = ~new_n222_ & new_n1124_;
  assign new_n1126_ = ~pv133_10_ & new_n1125_;
  assign new_n1127_ = new_n314_ & ~new_n1109_;
  assign new_n1128_ = new_n224_ & ~new_n1109_;
  assign new_n1129_ = ~new_n1110_ & ~new_n1111_;
  assign new_n1130_ = ~new_n1114_ & ~new_n1116_;
  assign new_n1131_ = new_n1129_ & new_n1130_;
  assign new_n1132_ = ~new_n1126_ & ~new_n1127_;
  assign new_n1133_ = ~new_n1128_ & new_n1132_;
  assign pv165_0_ = ~new_n1131_ | ~new_n1133_;
  assign new_n1135_ = pv47_25_ & new_n241_;
  assign new_n1136_ = pv84_1_ & ~new_n240_;
  assign new_n1137_ = pv47_18_ & new_n265_;
  assign new_n1138_ = pv47_22_ & new_n268_;
  assign new_n1139_ = ~new_n272_ & ~new_n1138_;
  assign new_n1140_ = ~new_n1135_ & ~new_n1136_;
  assign new_n1141_ = ~new_n1137_ & new_n1140_;
  assign new_n1142_ = new_n1139_ & new_n1141_;
  assign new_n1143_ = new_n351_ & ~new_n1142_;
  assign new_n1144_ = new_n354_ & ~new_n1142_;
  assign new_n1145_ = new_n360_ & ~new_n1142_;
  assign new_n1146_ = ~new_n333_ & new_n1145_;
  assign new_n1147_ = pv133_10_ & new_n1146_;
  assign new_n1148_ = new_n366_ & ~new_n1142_;
  assign new_n1149_ = new_n357_ & new_n1148_;
  assign new_n1150_ = pv116_1_ & new_n370_;
  assign new_n1151_ = pv133_9_ & new_n1150_;
  assign new_n1152_ = ~pv133_10_ & new_n1151_;
  assign new_n1153_ = ~new_n336_ & new_n1152_;
  assign new_n1154_ = ~new_n357_ & new_n1153_;
  assign new_n1155_ = new_n376_ & ~new_n1142_;
  assign new_n1156_ = new_n340_ & ~new_n1142_;
  assign new_n1157_ = ~new_n1143_ & ~new_n1144_;
  assign new_n1158_ = ~new_n1147_ & ~new_n1149_;
  assign new_n1159_ = new_n1157_ & new_n1158_;
  assign new_n1160_ = ~new_n1154_ & ~new_n1155_;
  assign new_n1161_ = ~new_n1156_ & new_n1160_;
  assign pv197_1_ = ~new_n1159_ | ~new_n1161_;
  assign new_n1163_ = pv84_29_ & new_n475_;
  assign new_n1164_ = pv84_29_ & new_n474_;
  assign new_n1165_ = pv84_29_ & new_n489_;
  assign new_n1166_ = pv116_12_ & new_n493_;
  assign new_n1167_ = pv133_9_ & new_n1166_;
  assign new_n1168_ = ~pv133_10_ & new_n1167_;
  assign new_n1169_ = ~new_n1165_ & ~new_n1168_;
  assign new_n1170_ = ~new_n1163_ & ~new_n1164_;
  assign new_n1171_ = ~new_n487_ & new_n1170_;
  assign pv212_12_ = ~new_n1169_ | ~new_n1171_;
  assign new_n1173_ = ~pv133_9_ & new_n215_;
  assign new_n1174_ = pv47_4_ & new_n241_;
  assign new_n1175_ = pv47_12_ & ~new_n240_;
  assign new_n1176_ = pv15_11_ & new_n265_;
  assign new_n1177_ = pv47_1_ & new_n268_;
  assign new_n1178_ = ~new_n272_ & ~new_n1177_;
  assign new_n1179_ = ~new_n1174_ & ~new_n1175_;
  assign new_n1180_ = ~new_n1176_ & new_n1179_;
  assign new_n1181_ = new_n1178_ & new_n1180_;
  assign new_n1182_ = new_n597_ & ~new_n1173_;
  assign new_n1183_ = ~new_n1181_ & new_n1182_;
  assign new_n1184_ = new_n600_ & ~new_n1173_;
  assign new_n1185_ = ~new_n1181_ & new_n1184_;
  assign new_n1186_ = ~new_n220_ & ~new_n1173_;
  assign new_n1187_ = ~pv133_10_ & new_n1186_;
  assign new_n1188_ = ~new_n222_ & new_n1187_;
  assign new_n1189_ = pv116_12_ & new_n1188_;
  assign new_n1190_ = ~new_n277_ & new_n1189_;
  assign new_n1191_ = new_n287_ & new_n1190_;
  assign new_n1192_ = ~new_n222_ & ~new_n1173_;
  assign new_n1193_ = ~new_n277_ & new_n1192_;
  assign new_n1194_ = ~new_n220_ & new_n1193_;
  assign new_n1195_ = ~new_n1181_ & new_n1194_;
  assign new_n1196_ = pv133_10_ & new_n1195_;
  assign new_n1197_ = ~new_n287_ & new_n1186_;
  assign new_n1198_ = ~new_n277_ & new_n1197_;
  assign new_n1199_ = pv84_12_ & new_n1198_;
  assign new_n1200_ = pv133_1_ & new_n1199_;
  assign new_n1201_ = ~pv133_10_ & new_n1200_;
  assign new_n1202_ = ~pv133_3_ & new_n1201_;
  assign new_n1203_ = pv133_2_ & new_n1202_;
  assign new_n1204_ = ~pv133_4_ & new_n1203_;
  assign new_n1205_ = ~pv133_7_ & new_n1204_;
  assign new_n1206_ = ~pv133_9_ & new_n1205_;
  assign new_n1207_ = ~new_n222_ & new_n1206_;
  assign new_n1208_ = ~pv133_10_ & new_n1207_;
  assign new_n1209_ = new_n220_ & ~new_n1173_;
  assign new_n1210_ = ~new_n1181_ & new_n1209_;
  assign new_n1211_ = new_n1173_ & ~new_n1181_;
  assign new_n1212_ = ~new_n1183_ & ~new_n1185_;
  assign new_n1213_ = ~new_n1191_ & ~new_n1196_;
  assign new_n1214_ = new_n1212_ & new_n1213_;
  assign new_n1215_ = ~new_n1208_ & ~new_n1210_;
  assign new_n1216_ = ~new_n1211_ & new_n1215_;
  assign pv146_0_ = ~new_n1214_ | ~new_n1216_;
  assign new_n1218_ = pv47_10_ & new_n241_;
  assign new_n1219_ = pv47_18_ & ~new_n240_;
  assign new_n1220_ = pv47_3_ & new_n265_;
  assign new_n1221_ = pv47_7_ & new_n268_;
  assign new_n1222_ = ~new_n272_ & ~new_n1221_;
  assign new_n1223_ = ~new_n1218_ & ~new_n1219_;
  assign new_n1224_ = ~new_n1220_ & new_n1223_;
  assign new_n1225_ = new_n1222_ & new_n1224_;
  assign new_n1226_ = new_n598_ & ~new_n1225_;
  assign new_n1227_ = new_n601_ & ~new_n1225_;
  assign new_n1228_ = pv116_18_ & new_n605_;
  assign new_n1229_ = ~new_n277_ & new_n1228_;
  assign new_n1230_ = new_n287_ & new_n1229_;
  assign new_n1231_ = new_n611_ & ~new_n1225_;
  assign new_n1232_ = pv133_10_ & new_n1231_;
  assign new_n1233_ = pv84_18_ & new_n615_;
  assign new_n1234_ = pv133_1_ & new_n1233_;
  assign new_n1235_ = ~pv133_10_ & new_n1234_;
  assign new_n1236_ = ~pv133_3_ & new_n1235_;
  assign new_n1237_ = pv133_2_ & new_n1236_;
  assign new_n1238_ = ~pv133_4_ & new_n1237_;
  assign new_n1239_ = ~pv133_7_ & new_n1238_;
  assign new_n1240_ = ~pv133_9_ & new_n1239_;
  assign new_n1241_ = ~new_n222_ & new_n1240_;
  assign new_n1242_ = ~pv133_10_ & new_n1241_;
  assign new_n1243_ = new_n314_ & ~new_n1225_;
  assign new_n1244_ = new_n224_ & ~new_n1225_;
  assign new_n1245_ = ~new_n1226_ & ~new_n1227_;
  assign new_n1246_ = ~new_n1230_ & ~new_n1232_;
  assign new_n1247_ = new_n1245_ & new_n1246_;
  assign new_n1248_ = ~new_n1242_ & ~new_n1243_;
  assign new_n1249_ = ~new_n1244_ & new_n1248_;
  assign pv165_1_ = ~new_n1247_ | ~new_n1249_;
  assign new_n1251_ = pv47_24_ & new_n241_;
  assign new_n1252_ = pv84_0_ & ~new_n240_;
  assign new_n1253_ = pv47_17_ & new_n265_;
  assign new_n1254_ = pv47_21_ & new_n268_;
  assign new_n1255_ = ~new_n272_ & ~new_n1254_;
  assign new_n1256_ = ~new_n1251_ & ~new_n1252_;
  assign new_n1257_ = ~new_n1253_ & new_n1256_;
  assign new_n1258_ = new_n1255_ & new_n1257_;
  assign new_n1259_ = new_n351_ & ~new_n1258_;
  assign new_n1260_ = new_n354_ & ~new_n1258_;
  assign new_n1261_ = new_n360_ & ~new_n1258_;
  assign new_n1262_ = ~new_n333_ & new_n1261_;
  assign new_n1263_ = pv133_10_ & new_n1262_;
  assign new_n1264_ = new_n366_ & ~new_n1258_;
  assign new_n1265_ = new_n357_ & new_n1264_;
  assign new_n1266_ = pv116_0_ & new_n370_;
  assign new_n1267_ = pv133_9_ & new_n1266_;
  assign new_n1268_ = ~pv133_10_ & new_n1267_;
  assign new_n1269_ = ~new_n336_ & new_n1268_;
  assign new_n1270_ = ~new_n357_ & new_n1269_;
  assign new_n1271_ = new_n376_ & ~new_n1258_;
  assign new_n1272_ = new_n340_ & ~new_n1258_;
  assign new_n1273_ = ~new_n1259_ & ~new_n1260_;
  assign new_n1274_ = ~new_n1263_ & ~new_n1265_;
  assign new_n1275_ = new_n1273_ & new_n1274_;
  assign new_n1276_ = ~new_n1270_ & ~new_n1271_;
  assign new_n1277_ = ~new_n1272_ & new_n1276_;
  assign pv197_0_ = ~new_n1275_ | ~new_n1277_;
  assign new_n1279_ = pv84_30_ & new_n475_;
  assign new_n1280_ = pv84_30_ & new_n474_;
  assign new_n1281_ = pv84_30_ & new_n489_;
  assign new_n1282_ = pv116_13_ & new_n493_;
  assign new_n1283_ = pv133_9_ & new_n1282_;
  assign new_n1284_ = ~pv133_10_ & new_n1283_;
  assign new_n1285_ = ~new_n1281_ & ~new_n1284_;
  assign new_n1286_ = ~new_n1279_ & ~new_n1280_;
  assign new_n1287_ = ~new_n487_ & new_n1286_;
  assign pv212_13_ = ~new_n1285_ | ~new_n1287_;
  assign new_n1289_ = pv47_15_ & new_n241_;
  assign new_n1290_ = pv47_23_ & ~new_n240_;
  assign new_n1291_ = pv47_8_ & new_n265_;
  assign new_n1292_ = pv47_12_ & new_n268_;
  assign new_n1293_ = ~new_n272_ & ~new_n1292_;
  assign new_n1294_ = ~new_n1289_ & ~new_n1290_;
  assign new_n1295_ = ~new_n1291_ & new_n1294_;
  assign new_n1296_ = new_n1293_ & new_n1295_;
  assign new_n1297_ = new_n598_ & ~new_n1296_;
  assign new_n1298_ = new_n601_ & ~new_n1296_;
  assign new_n1299_ = pv116_23_ & new_n605_;
  assign new_n1300_ = ~new_n277_ & new_n1299_;
  assign new_n1301_ = new_n287_ & new_n1300_;
  assign new_n1302_ = new_n611_ & ~new_n1296_;
  assign new_n1303_ = pv133_10_ & new_n1302_;
  assign new_n1304_ = pv84_23_ & new_n615_;
  assign new_n1305_ = pv133_1_ & new_n1304_;
  assign new_n1306_ = ~pv133_10_ & new_n1305_;
  assign new_n1307_ = ~pv133_3_ & new_n1306_;
  assign new_n1308_ = pv133_2_ & new_n1307_;
  assign new_n1309_ = ~pv133_4_ & new_n1308_;
  assign new_n1310_ = ~pv133_7_ & new_n1309_;
  assign new_n1311_ = ~pv133_9_ & new_n1310_;
  assign new_n1312_ = ~new_n222_ & new_n1311_;
  assign new_n1313_ = ~pv133_10_ & new_n1312_;
  assign new_n1314_ = new_n314_ & ~new_n1296_;
  assign new_n1315_ = new_n224_ & ~new_n1296_;
  assign new_n1316_ = ~new_n1297_ & ~new_n1298_;
  assign new_n1317_ = ~new_n1301_ & ~new_n1303_;
  assign new_n1318_ = new_n1316_ & new_n1317_;
  assign new_n1319_ = ~new_n1313_ & ~new_n1314_;
  assign new_n1320_ = ~new_n1315_ & new_n1319_;
  assign pv165_6_ = ~new_n1318_ | ~new_n1320_;
  assign new_n1322_ = pv47_22_ & new_n241_;
  assign new_n1323_ = pv47_30_ & ~new_n240_;
  assign new_n1324_ = pv47_15_ & new_n265_;
  assign new_n1325_ = pv47_19_ & new_n268_;
  assign new_n1326_ = ~new_n272_ & ~new_n1325_;
  assign new_n1327_ = ~new_n1322_ & ~new_n1323_;
  assign new_n1328_ = ~new_n1324_ & new_n1327_;
  assign new_n1329_ = new_n1326_ & new_n1328_;
  assign new_n1330_ = new_n598_ & ~new_n1329_;
  assign new_n1331_ = new_n601_ & ~new_n1329_;
  assign new_n1332_ = pv116_30_ & new_n605_;
  assign new_n1333_ = ~new_n277_ & new_n1332_;
  assign new_n1334_ = new_n287_ & new_n1333_;
  assign new_n1335_ = new_n611_ & ~new_n1329_;
  assign new_n1336_ = pv133_10_ & new_n1335_;
  assign new_n1337_ = pv84_30_ & new_n615_;
  assign new_n1338_ = pv133_1_ & new_n1337_;
  assign new_n1339_ = ~pv133_10_ & new_n1338_;
  assign new_n1340_ = ~pv133_3_ & new_n1339_;
  assign new_n1341_ = pv133_2_ & new_n1340_;
  assign new_n1342_ = ~pv133_4_ & new_n1341_;
  assign new_n1343_ = ~pv133_7_ & new_n1342_;
  assign new_n1344_ = ~pv133_9_ & new_n1343_;
  assign new_n1345_ = ~new_n222_ & new_n1344_;
  assign new_n1346_ = ~pv133_10_ & new_n1345_;
  assign new_n1347_ = new_n314_ & ~new_n1329_;
  assign new_n1348_ = new_n224_ & ~new_n1329_;
  assign new_n1349_ = ~new_n1330_ & ~new_n1331_;
  assign new_n1350_ = ~new_n1334_ & ~new_n1336_;
  assign new_n1351_ = new_n1349_ & new_n1350_;
  assign new_n1352_ = ~new_n1346_ & ~new_n1347_;
  assign new_n1353_ = ~new_n1348_ & new_n1352_;
  assign pv165_13_ = ~new_n1351_ | ~new_n1353_;
  assign new_n1355_ = pv47_16_ & new_n241_;
  assign new_n1356_ = pv47_24_ & ~new_n240_;
  assign new_n1357_ = pv47_9_ & new_n265_;
  assign new_n1358_ = pv47_13_ & new_n268_;
  assign new_n1359_ = ~new_n272_ & ~new_n1358_;
  assign new_n1360_ = ~new_n1355_ & ~new_n1356_;
  assign new_n1361_ = ~new_n1357_ & new_n1360_;
  assign new_n1362_ = new_n1359_ & new_n1361_;
  assign new_n1363_ = new_n598_ & ~new_n1362_;
  assign new_n1364_ = new_n601_ & ~new_n1362_;
  assign new_n1365_ = pv116_24_ & new_n605_;
  assign new_n1366_ = ~new_n277_ & new_n1365_;
  assign new_n1367_ = new_n287_ & new_n1366_;
  assign new_n1368_ = new_n611_ & ~new_n1362_;
  assign new_n1369_ = pv133_10_ & new_n1368_;
  assign new_n1370_ = pv84_24_ & new_n615_;
  assign new_n1371_ = pv133_1_ & new_n1370_;
  assign new_n1372_ = ~pv133_10_ & new_n1371_;
  assign new_n1373_ = ~pv133_3_ & new_n1372_;
  assign new_n1374_ = pv133_2_ & new_n1373_;
  assign new_n1375_ = ~pv133_4_ & new_n1374_;
  assign new_n1376_ = ~pv133_7_ & new_n1375_;
  assign new_n1377_ = ~pv133_9_ & new_n1376_;
  assign new_n1378_ = ~new_n222_ & new_n1377_;
  assign new_n1379_ = ~pv133_10_ & new_n1378_;
  assign new_n1380_ = new_n314_ & ~new_n1362_;
  assign new_n1381_ = new_n224_ & ~new_n1362_;
  assign new_n1382_ = ~new_n1363_ & ~new_n1364_;
  assign new_n1383_ = ~new_n1367_ & ~new_n1369_;
  assign new_n1384_ = new_n1382_ & new_n1383_;
  assign new_n1385_ = ~new_n1379_ & ~new_n1380_;
  assign new_n1386_ = ~new_n1381_ & new_n1385_;
  assign pv165_7_ = ~new_n1384_ | ~new_n1386_;
  assign new_n1388_ = pv47_23_ & new_n241_;
  assign new_n1389_ = pv47_31_ & ~new_n240_;
  assign new_n1390_ = pv47_16_ & new_n265_;
  assign new_n1391_ = pv47_20_ & new_n268_;
  assign new_n1392_ = ~new_n272_ & ~new_n1391_;
  assign new_n1393_ = ~new_n1388_ & ~new_n1389_;
  assign new_n1394_ = ~new_n1390_ & new_n1393_;
  assign new_n1395_ = new_n1392_ & new_n1394_;
  assign new_n1396_ = new_n598_ & ~new_n1395_;
  assign new_n1397_ = new_n601_ & ~new_n1395_;
  assign new_n1398_ = pv116_31_ & new_n605_;
  assign new_n1399_ = ~new_n277_ & new_n1398_;
  assign new_n1400_ = new_n287_ & new_n1399_;
  assign new_n1401_ = new_n611_ & ~new_n1395_;
  assign new_n1402_ = pv133_10_ & new_n1401_;
  assign new_n1403_ = pv84_31_ & new_n615_;
  assign new_n1404_ = pv133_1_ & new_n1403_;
  assign new_n1405_ = ~pv133_10_ & new_n1404_;
  assign new_n1406_ = ~pv133_3_ & new_n1405_;
  assign new_n1407_ = pv133_2_ & new_n1406_;
  assign new_n1408_ = ~pv133_4_ & new_n1407_;
  assign new_n1409_ = ~pv133_7_ & new_n1408_;
  assign new_n1410_ = ~pv133_9_ & new_n1409_;
  assign new_n1411_ = ~new_n222_ & new_n1410_;
  assign new_n1412_ = ~pv133_10_ & new_n1411_;
  assign new_n1413_ = new_n314_ & ~new_n1395_;
  assign new_n1414_ = new_n224_ & ~new_n1395_;
  assign new_n1415_ = ~new_n1396_ & ~new_n1397_;
  assign new_n1416_ = ~new_n1400_ & ~new_n1402_;
  assign new_n1417_ = new_n1415_ & new_n1416_;
  assign new_n1418_ = ~new_n1412_ & ~new_n1413_;
  assign new_n1419_ = ~new_n1414_ & new_n1418_;
  assign pv165_14_ = ~new_n1417_ | ~new_n1419_;
  assign new_n1421_ = pv47_13_ & new_n241_;
  assign new_n1422_ = pv47_21_ & ~new_n240_;
  assign new_n1423_ = pv47_6_ & new_n265_;
  assign new_n1424_ = pv47_10_ & new_n268_;
  assign new_n1425_ = ~new_n272_ & ~new_n1424_;
  assign new_n1426_ = ~new_n1421_ & ~new_n1422_;
  assign new_n1427_ = ~new_n1423_ & new_n1426_;
  assign new_n1428_ = new_n1425_ & new_n1427_;
  assign new_n1429_ = new_n598_ & ~new_n1428_;
  assign new_n1430_ = new_n601_ & ~new_n1428_;
  assign new_n1431_ = pv116_21_ & new_n605_;
  assign new_n1432_ = ~new_n277_ & new_n1431_;
  assign new_n1433_ = new_n287_ & new_n1432_;
  assign new_n1434_ = new_n611_ & ~new_n1428_;
  assign new_n1435_ = pv133_10_ & new_n1434_;
  assign new_n1436_ = pv84_21_ & new_n615_;
  assign new_n1437_ = pv133_1_ & new_n1436_;
  assign new_n1438_ = ~pv133_10_ & new_n1437_;
  assign new_n1439_ = ~pv133_3_ & new_n1438_;
  assign new_n1440_ = pv133_2_ & new_n1439_;
  assign new_n1441_ = ~pv133_4_ & new_n1440_;
  assign new_n1442_ = ~pv133_7_ & new_n1441_;
  assign new_n1443_ = ~pv133_9_ & new_n1442_;
  assign new_n1444_ = ~new_n222_ & new_n1443_;
  assign new_n1445_ = ~pv133_10_ & new_n1444_;
  assign new_n1446_ = new_n314_ & ~new_n1428_;
  assign new_n1447_ = new_n224_ & ~new_n1428_;
  assign new_n1448_ = ~new_n1429_ & ~new_n1430_;
  assign new_n1449_ = ~new_n1433_ & ~new_n1435_;
  assign new_n1450_ = new_n1448_ & new_n1449_;
  assign new_n1451_ = ~new_n1445_ & ~new_n1446_;
  assign new_n1452_ = ~new_n1447_ & new_n1451_;
  assign pv165_4_ = ~new_n1450_ | ~new_n1452_;
  assign new_n1454_ = pv47_20_ & new_n241_;
  assign new_n1455_ = pv47_28_ & ~new_n240_;
  assign new_n1456_ = pv47_13_ & new_n265_;
  assign new_n1457_ = pv47_17_ & new_n268_;
  assign new_n1458_ = ~new_n272_ & ~new_n1457_;
  assign new_n1459_ = ~new_n1454_ & ~new_n1455_;
  assign new_n1460_ = ~new_n1456_ & new_n1459_;
  assign new_n1461_ = new_n1458_ & new_n1460_;
  assign new_n1462_ = new_n598_ & ~new_n1461_;
  assign new_n1463_ = new_n601_ & ~new_n1461_;
  assign new_n1464_ = pv116_28_ & new_n605_;
  assign new_n1465_ = ~new_n277_ & new_n1464_;
  assign new_n1466_ = new_n287_ & new_n1465_;
  assign new_n1467_ = new_n611_ & ~new_n1461_;
  assign new_n1468_ = pv133_10_ & new_n1467_;
  assign new_n1469_ = pv84_28_ & new_n615_;
  assign new_n1470_ = pv133_1_ & new_n1469_;
  assign new_n1471_ = ~pv133_10_ & new_n1470_;
  assign new_n1472_ = ~pv133_3_ & new_n1471_;
  assign new_n1473_ = pv133_2_ & new_n1472_;
  assign new_n1474_ = ~pv133_4_ & new_n1473_;
  assign new_n1475_ = ~pv133_7_ & new_n1474_;
  assign new_n1476_ = ~pv133_9_ & new_n1475_;
  assign new_n1477_ = ~new_n222_ & new_n1476_;
  assign new_n1478_ = ~pv133_10_ & new_n1477_;
  assign new_n1479_ = new_n314_ & ~new_n1461_;
  assign new_n1480_ = new_n224_ & ~new_n1461_;
  assign new_n1481_ = ~new_n1462_ & ~new_n1463_;
  assign new_n1482_ = ~new_n1466_ & ~new_n1468_;
  assign new_n1483_ = new_n1481_ & new_n1482_;
  assign new_n1484_ = ~new_n1478_ & ~new_n1479_;
  assign new_n1485_ = ~new_n1480_ & new_n1484_;
  assign pv165_11_ = ~new_n1483_ | ~new_n1485_;
  assign new_n1487_ = pv47_14_ & new_n241_;
  assign new_n1488_ = pv47_22_ & ~new_n240_;
  assign new_n1489_ = pv47_7_ & new_n265_;
  assign new_n1490_ = pv47_11_ & new_n268_;
  assign new_n1491_ = ~new_n272_ & ~new_n1490_;
  assign new_n1492_ = ~new_n1487_ & ~new_n1488_;
  assign new_n1493_ = ~new_n1489_ & new_n1492_;
  assign new_n1494_ = new_n1491_ & new_n1493_;
  assign new_n1495_ = new_n598_ & ~new_n1494_;
  assign new_n1496_ = new_n601_ & ~new_n1494_;
  assign new_n1497_ = pv116_22_ & new_n605_;
  assign new_n1498_ = ~new_n277_ & new_n1497_;
  assign new_n1499_ = new_n287_ & new_n1498_;
  assign new_n1500_ = new_n611_ & ~new_n1494_;
  assign new_n1501_ = pv133_10_ & new_n1500_;
  assign new_n1502_ = pv84_22_ & new_n615_;
  assign new_n1503_ = pv133_1_ & new_n1502_;
  assign new_n1504_ = ~pv133_10_ & new_n1503_;
  assign new_n1505_ = ~pv133_3_ & new_n1504_;
  assign new_n1506_ = pv133_2_ & new_n1505_;
  assign new_n1507_ = ~pv133_4_ & new_n1506_;
  assign new_n1508_ = ~pv133_7_ & new_n1507_;
  assign new_n1509_ = ~pv133_9_ & new_n1508_;
  assign new_n1510_ = ~new_n222_ & new_n1509_;
  assign new_n1511_ = ~pv133_10_ & new_n1510_;
  assign new_n1512_ = new_n314_ & ~new_n1494_;
  assign new_n1513_ = new_n224_ & ~new_n1494_;
  assign new_n1514_ = ~new_n1495_ & ~new_n1496_;
  assign new_n1515_ = ~new_n1499_ & ~new_n1501_;
  assign new_n1516_ = new_n1514_ & new_n1515_;
  assign new_n1517_ = ~new_n1511_ & ~new_n1512_;
  assign new_n1518_ = ~new_n1513_ & new_n1517_;
  assign pv165_5_ = ~new_n1516_ | ~new_n1518_;
  assign new_n1520_ = pv47_21_ & new_n241_;
  assign new_n1521_ = pv47_29_ & ~new_n240_;
  assign new_n1522_ = pv47_14_ & new_n265_;
  assign new_n1523_ = pv47_18_ & new_n268_;
  assign new_n1524_ = ~new_n272_ & ~new_n1523_;
  assign new_n1525_ = ~new_n1520_ & ~new_n1521_;
  assign new_n1526_ = ~new_n1522_ & new_n1525_;
  assign new_n1527_ = new_n1524_ & new_n1526_;
  assign new_n1528_ = new_n598_ & ~new_n1527_;
  assign new_n1529_ = new_n601_ & ~new_n1527_;
  assign new_n1530_ = pv116_29_ & new_n605_;
  assign new_n1531_ = ~new_n277_ & new_n1530_;
  assign new_n1532_ = new_n287_ & new_n1531_;
  assign new_n1533_ = new_n611_ & ~new_n1527_;
  assign new_n1534_ = pv133_10_ & new_n1533_;
  assign new_n1535_ = pv84_29_ & new_n615_;
  assign new_n1536_ = pv133_1_ & new_n1535_;
  assign new_n1537_ = ~pv133_10_ & new_n1536_;
  assign new_n1538_ = ~pv133_3_ & new_n1537_;
  assign new_n1539_ = pv133_2_ & new_n1538_;
  assign new_n1540_ = ~pv133_4_ & new_n1539_;
  assign new_n1541_ = ~pv133_7_ & new_n1540_;
  assign new_n1542_ = ~pv133_9_ & new_n1541_;
  assign new_n1543_ = ~new_n222_ & new_n1542_;
  assign new_n1544_ = ~pv133_10_ & new_n1543_;
  assign new_n1545_ = new_n314_ & ~new_n1527_;
  assign new_n1546_ = new_n224_ & ~new_n1527_;
  assign new_n1547_ = ~new_n1528_ & ~new_n1529_;
  assign new_n1548_ = ~new_n1532_ & ~new_n1534_;
  assign new_n1549_ = new_n1547_ & new_n1548_;
  assign new_n1550_ = ~new_n1544_ & ~new_n1545_;
  assign new_n1551_ = ~new_n1546_ & new_n1550_;
  assign pv165_12_ = ~new_n1549_ | ~new_n1551_;
  assign new_n1553_ = pv47_4_ & ~new_n240_;
  assign new_n1554_ = pv84_4_ & new_n268_;
  assign new_n1555_ = pv15_3_ & new_n265_;
  assign new_n1556_ = ~new_n1553_ & ~new_n1554_;
  assign new_n1557_ = ~new_n272_ & ~new_n1555_;
  assign new_n1558_ = new_n1556_ & new_n1557_;
  assign new_n1559_ = new_n517_ & ~new_n1558_;
  assign new_n1560_ = new_n520_ & ~new_n1558_;
  assign new_n1561_ = new_n522_ & ~new_n1558_;
  assign new_n1562_ = pv116_4_ & new_n526_;
  assign new_n1563_ = ~pv133_10_ & new_n1562_;
  assign new_n1564_ = ~new_n1559_ & ~new_n1560_;
  assign new_n1565_ = ~new_n1561_ & ~new_n1563_;
  assign pv142_1_ = ~new_n1564_ | ~new_n1565_;
  assign new_n1567_ = pv84_8_ & new_n241_;
  assign new_n1568_ = pv84_16_ & ~new_n240_;
  assign new_n1569_ = pv84_1_ & new_n265_;
  assign new_n1570_ = pv84_5_ & new_n268_;
  assign new_n1571_ = ~new_n272_ & ~new_n1570_;
  assign new_n1572_ = ~new_n1567_ & ~new_n1568_;
  assign new_n1573_ = ~new_n1569_ & new_n1572_;
  assign new_n1574_ = new_n1571_ & new_n1573_;
  assign new_n1575_ = new_n351_ & ~new_n1574_;
  assign new_n1576_ = new_n354_ & ~new_n1574_;
  assign new_n1577_ = new_n360_ & ~new_n1574_;
  assign new_n1578_ = ~new_n333_ & new_n1577_;
  assign new_n1579_ = pv133_10_ & new_n1578_;
  assign new_n1580_ = new_n366_ & ~new_n1574_;
  assign new_n1581_ = new_n357_ & new_n1580_;
  assign new_n1582_ = pv116_16_ & new_n370_;
  assign new_n1583_ = pv133_9_ & new_n1582_;
  assign new_n1584_ = ~pv133_10_ & new_n1583_;
  assign new_n1585_ = ~new_n336_ & new_n1584_;
  assign new_n1586_ = ~new_n357_ & new_n1585_;
  assign new_n1587_ = new_n376_ & ~new_n1574_;
  assign new_n1588_ = new_n340_ & ~new_n1574_;
  assign new_n1589_ = ~new_n1575_ & ~new_n1576_;
  assign new_n1590_ = ~new_n1579_ & ~new_n1581_;
  assign new_n1591_ = new_n1589_ & new_n1590_;
  assign new_n1592_ = ~new_n1586_ & ~new_n1587_;
  assign new_n1593_ = ~new_n1588_ & new_n1592_;
  assign pv197_16_ = ~new_n1591_ | ~new_n1593_;
  assign new_n1595_ = pv84_21_ & new_n241_;
  assign new_n1596_ = pv84_29_ & ~new_n240_;
  assign new_n1597_ = pv84_14_ & new_n265_;
  assign new_n1598_ = pv84_18_ & new_n268_;
  assign new_n1599_ = ~new_n272_ & ~new_n1598_;
  assign new_n1600_ = ~new_n1595_ & ~new_n1596_;
  assign new_n1601_ = ~new_n1597_ & new_n1600_;
  assign new_n1602_ = new_n1599_ & new_n1601_;
  assign new_n1603_ = new_n351_ & ~new_n1602_;
  assign new_n1604_ = new_n354_ & ~new_n1602_;
  assign new_n1605_ = new_n360_ & ~new_n1602_;
  assign new_n1606_ = ~new_n333_ & new_n1605_;
  assign new_n1607_ = pv133_10_ & new_n1606_;
  assign new_n1608_ = new_n366_ & ~new_n1602_;
  assign new_n1609_ = new_n357_ & new_n1608_;
  assign new_n1610_ = pv116_29_ & new_n370_;
  assign new_n1611_ = pv133_9_ & new_n1610_;
  assign new_n1612_ = ~pv133_10_ & new_n1611_;
  assign new_n1613_ = ~new_n336_ & new_n1612_;
  assign new_n1614_ = ~new_n357_ & new_n1613_;
  assign new_n1615_ = new_n376_ & ~new_n1602_;
  assign new_n1616_ = new_n340_ & ~new_n1602_;
  assign new_n1617_ = ~new_n1603_ & ~new_n1604_;
  assign new_n1618_ = ~new_n1607_ & ~new_n1609_;
  assign new_n1619_ = new_n1617_ & new_n1618_;
  assign new_n1620_ = ~new_n1614_ & ~new_n1615_;
  assign new_n1621_ = ~new_n1616_ & new_n1620_;
  assign pv197_29_ = ~new_n1619_ | ~new_n1621_;
  assign new_n1623_ = pv84_22_ & new_n475_;
  assign new_n1624_ = pv84_22_ & new_n474_;
  assign new_n1625_ = pv84_22_ & new_n489_;
  assign new_n1626_ = pv116_5_ & new_n493_;
  assign new_n1627_ = pv133_9_ & new_n1626_;
  assign new_n1628_ = ~pv133_10_ & new_n1627_;
  assign new_n1629_ = ~new_n1625_ & ~new_n1628_;
  assign new_n1630_ = ~new_n1623_ & ~new_n1624_;
  assign new_n1631_ = ~new_n487_ & new_n1630_;
  assign pv212_5_ = ~new_n1629_ | ~new_n1631_;
  assign new_n1633_ = pv47_5_ & ~new_n240_;
  assign new_n1634_ = pv15_4_ & new_n265_;
  assign new_n1635_ = ~new_n1570_ & ~new_n1633_;
  assign new_n1636_ = ~new_n272_ & ~new_n1634_;
  assign new_n1637_ = new_n1635_ & new_n1636_;
  assign new_n1638_ = new_n517_ & ~new_n1637_;
  assign new_n1639_ = new_n520_ & ~new_n1637_;
  assign new_n1640_ = new_n522_ & ~new_n1637_;
  assign new_n1641_ = pv116_5_ & new_n526_;
  assign new_n1642_ = ~pv133_10_ & new_n1641_;
  assign new_n1643_ = ~new_n1638_ & ~new_n1639_;
  assign new_n1644_ = ~new_n1640_ & ~new_n1642_;
  assign pv142_2_ = ~new_n1643_ | ~new_n1644_;
  assign new_n1646_ = pv84_9_ & new_n241_;
  assign new_n1647_ = pv84_17_ & ~new_n240_;
  assign new_n1648_ = pv84_2_ & new_n265_;
  assign new_n1649_ = pv84_6_ & new_n268_;
  assign new_n1650_ = ~new_n272_ & ~new_n1649_;
  assign new_n1651_ = ~new_n1646_ & ~new_n1647_;
  assign new_n1652_ = ~new_n1648_ & new_n1651_;
  assign new_n1653_ = new_n1650_ & new_n1652_;
  assign new_n1654_ = new_n351_ & ~new_n1653_;
  assign new_n1655_ = new_n354_ & ~new_n1653_;
  assign new_n1656_ = new_n360_ & ~new_n1653_;
  assign new_n1657_ = ~new_n333_ & new_n1656_;
  assign new_n1658_ = pv133_10_ & new_n1657_;
  assign new_n1659_ = new_n366_ & ~new_n1653_;
  assign new_n1660_ = new_n357_ & new_n1659_;
  assign new_n1661_ = pv116_17_ & new_n370_;
  assign new_n1662_ = pv133_9_ & new_n1661_;
  assign new_n1663_ = ~pv133_10_ & new_n1662_;
  assign new_n1664_ = ~new_n336_ & new_n1663_;
  assign new_n1665_ = ~new_n357_ & new_n1664_;
  assign new_n1666_ = new_n376_ & ~new_n1653_;
  assign new_n1667_ = new_n340_ & ~new_n1653_;
  assign new_n1668_ = ~new_n1654_ & ~new_n1655_;
  assign new_n1669_ = ~new_n1658_ & ~new_n1660_;
  assign new_n1670_ = new_n1668_ & new_n1669_;
  assign new_n1671_ = ~new_n1665_ & ~new_n1666_;
  assign new_n1672_ = ~new_n1667_ & new_n1671_;
  assign pv197_17_ = ~new_n1670_ | ~new_n1672_;
  assign new_n1674_ = pv84_20_ & new_n241_;
  assign new_n1675_ = pv84_28_ & ~new_n240_;
  assign new_n1676_ = pv84_13_ & new_n265_;
  assign new_n1677_ = pv84_17_ & new_n268_;
  assign new_n1678_ = ~new_n272_ & ~new_n1677_;
  assign new_n1679_ = ~new_n1674_ & ~new_n1675_;
  assign new_n1680_ = ~new_n1676_ & new_n1679_;
  assign new_n1681_ = new_n1678_ & new_n1680_;
  assign new_n1682_ = new_n351_ & ~new_n1681_;
  assign new_n1683_ = new_n354_ & ~new_n1681_;
  assign new_n1684_ = new_n360_ & ~new_n1681_;
  assign new_n1685_ = ~new_n333_ & new_n1684_;
  assign new_n1686_ = pv133_10_ & new_n1685_;
  assign new_n1687_ = new_n366_ & ~new_n1681_;
  assign new_n1688_ = new_n357_ & new_n1687_;
  assign new_n1689_ = pv116_28_ & new_n370_;
  assign new_n1690_ = pv133_9_ & new_n1689_;
  assign new_n1691_ = ~pv133_10_ & new_n1690_;
  assign new_n1692_ = ~new_n336_ & new_n1691_;
  assign new_n1693_ = ~new_n357_ & new_n1692_;
  assign new_n1694_ = new_n376_ & ~new_n1681_;
  assign new_n1695_ = new_n340_ & ~new_n1681_;
  assign new_n1696_ = ~new_n1682_ & ~new_n1683_;
  assign new_n1697_ = ~new_n1686_ & ~new_n1688_;
  assign new_n1698_ = new_n1696_ & new_n1697_;
  assign new_n1699_ = ~new_n1693_ & ~new_n1694_;
  assign new_n1700_ = ~new_n1695_ & new_n1699_;
  assign pv197_28_ = ~new_n1698_ | ~new_n1700_;
  assign new_n1702_ = pv84_21_ & new_n475_;
  assign new_n1703_ = pv84_21_ & new_n474_;
  assign new_n1704_ = pv84_21_ & new_n489_;
  assign new_n1705_ = pv116_4_ & new_n493_;
  assign new_n1706_ = pv133_9_ & new_n1705_;
  assign new_n1707_ = ~pv133_10_ & new_n1706_;
  assign new_n1708_ = ~new_n1704_ & ~new_n1707_;
  assign new_n1709_ = ~new_n1702_ & ~new_n1703_;
  assign new_n1710_ = ~new_n487_ & new_n1709_;
  assign pv212_4_ = ~new_n1708_ | ~new_n1710_;
  assign new_n1712_ = pv47_6_ & ~new_n240_;
  assign new_n1713_ = pv15_5_ & new_n265_;
  assign new_n1714_ = ~new_n1649_ & ~new_n1712_;
  assign new_n1715_ = ~new_n272_ & ~new_n1713_;
  assign new_n1716_ = new_n1714_ & new_n1715_;
  assign new_n1717_ = new_n517_ & ~new_n1716_;
  assign new_n1718_ = new_n520_ & ~new_n1716_;
  assign new_n1719_ = new_n522_ & ~new_n1716_;
  assign new_n1720_ = pv116_6_ & new_n526_;
  assign new_n1721_ = ~pv133_10_ & new_n1720_;
  assign new_n1722_ = ~new_n1717_ & ~new_n1718_;
  assign new_n1723_ = ~new_n1719_ & ~new_n1721_;
  assign pv142_3_ = ~new_n1722_ | ~new_n1723_;
  assign new_n1725_ = pv47_1_ & new_n241_;
  assign new_n1726_ = pv47_9_ & ~new_n240_;
  assign new_n1727_ = pv15_8_ & new_n265_;
  assign new_n1728_ = ~new_n1725_ & ~new_n1726_;
  assign new_n1729_ = ~new_n1727_ & new_n1728_;
  assign new_n1730_ = new_n389_ & new_n1729_;
  assign new_n1731_ = ~pv133_4_ & ~pv133_9_;
  assign new_n1732_ = ~new_n1730_ & new_n1731_;
  assign new_n1733_ = new_n519_ & ~new_n1731_;
  assign new_n1734_ = ~new_n1730_ & new_n1733_;
  assign new_n1735_ = new_n277_ & ~new_n1731_;
  assign new_n1736_ = ~new_n1730_ & new_n1735_;
  assign new_n1737_ = new_n525_ & ~new_n1731_;
  assign new_n1738_ = pv116_9_ & new_n1737_;
  assign new_n1739_ = ~pv133_10_ & new_n1738_;
  assign new_n1740_ = ~new_n1732_ & ~new_n1734_;
  assign new_n1741_ = ~new_n1736_ & ~new_n1739_;
  assign pv143_0_ = ~new_n1740_ | ~new_n1741_;
  assign new_n1743_ = pv84_10_ & new_n241_;
  assign new_n1744_ = pv84_18_ & ~new_n240_;
  assign new_n1745_ = pv84_3_ & new_n265_;
  assign new_n1746_ = pv84_7_ & new_n268_;
  assign new_n1747_ = ~new_n272_ & ~new_n1746_;
  assign new_n1748_ = ~new_n1743_ & ~new_n1744_;
  assign new_n1749_ = ~new_n1745_ & new_n1748_;
  assign new_n1750_ = new_n1747_ & new_n1749_;
  assign new_n1751_ = new_n351_ & ~new_n1750_;
  assign new_n1752_ = new_n354_ & ~new_n1750_;
  assign new_n1753_ = new_n360_ & ~new_n1750_;
  assign new_n1754_ = ~new_n333_ & new_n1753_;
  assign new_n1755_ = pv133_10_ & new_n1754_;
  assign new_n1756_ = new_n366_ & ~new_n1750_;
  assign new_n1757_ = new_n357_ & new_n1756_;
  assign new_n1758_ = pv116_18_ & new_n370_;
  assign new_n1759_ = pv133_9_ & new_n1758_;
  assign new_n1760_ = ~pv133_10_ & new_n1759_;
  assign new_n1761_ = ~new_n336_ & new_n1760_;
  assign new_n1762_ = ~new_n357_ & new_n1761_;
  assign new_n1763_ = new_n376_ & ~new_n1750_;
  assign new_n1764_ = new_n340_ & ~new_n1750_;
  assign new_n1765_ = ~new_n1751_ & ~new_n1752_;
  assign new_n1766_ = ~new_n1755_ & ~new_n1757_;
  assign new_n1767_ = new_n1765_ & new_n1766_;
  assign new_n1768_ = ~new_n1762_ & ~new_n1763_;
  assign new_n1769_ = ~new_n1764_ & new_n1768_;
  assign pv197_18_ = ~new_n1767_ | ~new_n1769_;
  assign new_n1771_ = pv84_19_ & new_n241_;
  assign new_n1772_ = pv84_27_ & ~new_n240_;
  assign new_n1773_ = pv84_12_ & new_n265_;
  assign new_n1774_ = pv84_16_ & new_n268_;
  assign new_n1775_ = ~new_n272_ & ~new_n1774_;
  assign new_n1776_ = ~new_n1771_ & ~new_n1772_;
  assign new_n1777_ = ~new_n1773_ & new_n1776_;
  assign new_n1778_ = new_n1775_ & new_n1777_;
  assign new_n1779_ = new_n351_ & ~new_n1778_;
  assign new_n1780_ = new_n354_ & ~new_n1778_;
  assign new_n1781_ = new_n360_ & ~new_n1778_;
  assign new_n1782_ = ~new_n333_ & new_n1781_;
  assign new_n1783_ = pv133_10_ & new_n1782_;
  assign new_n1784_ = new_n366_ & ~new_n1778_;
  assign new_n1785_ = new_n357_ & new_n1784_;
  assign new_n1786_ = pv116_27_ & new_n370_;
  assign new_n1787_ = pv133_9_ & new_n1786_;
  assign new_n1788_ = ~pv133_10_ & new_n1787_;
  assign new_n1789_ = ~new_n336_ & new_n1788_;
  assign new_n1790_ = ~new_n357_ & new_n1789_;
  assign new_n1791_ = new_n376_ & ~new_n1778_;
  assign new_n1792_ = new_n340_ & ~new_n1778_;
  assign new_n1793_ = ~new_n1779_ & ~new_n1780_;
  assign new_n1794_ = ~new_n1783_ & ~new_n1785_;
  assign new_n1795_ = new_n1793_ & new_n1794_;
  assign new_n1796_ = ~new_n1790_ & ~new_n1791_;
  assign new_n1797_ = ~new_n1792_ & new_n1796_;
  assign pv197_27_ = ~new_n1795_ | ~new_n1797_;
  assign new_n1799_ = pv84_24_ & new_n475_;
  assign new_n1800_ = pv84_24_ & new_n474_;
  assign new_n1801_ = pv84_24_ & new_n489_;
  assign new_n1802_ = pv116_7_ & new_n493_;
  assign new_n1803_ = pv133_9_ & new_n1802_;
  assign new_n1804_ = ~pv133_10_ & new_n1803_;
  assign new_n1805_ = ~new_n1801_ & ~new_n1804_;
  assign new_n1806_ = ~new_n1799_ & ~new_n1800_;
  assign new_n1807_ = ~new_n487_ & new_n1806_;
  assign pv212_7_ = ~new_n1805_ | ~new_n1807_;
  assign new_n1809_ = ~pv133_8_ & pv133_7_;
  assign new_n1810_ = ~pv133_9_ & new_n1809_;
  assign new_n1811_ = ~pv133_4_ & ~pv133_8_;
  assign new_n1812_ = pv133_1_ & new_n1811_;
  assign new_n1813_ = pv133_2_ & new_n1812_;
  assign new_n1814_ = ~pv133_9_ & new_n1813_;
  assign new_n1815_ = pv47_2_ & ~new_n240_;
  assign new_n1816_ = pv84_2_ & new_n268_;
  assign new_n1817_ = pv15_1_ & new_n265_;
  assign new_n1818_ = ~new_n1815_ & ~new_n1816_;
  assign new_n1819_ = ~new_n272_ & ~new_n1817_;
  assign new_n1820_ = new_n1818_ & new_n1819_;
  assign new_n1821_ = pv133_10_ & ~new_n1810_;
  assign new_n1822_ = ~new_n1814_ & new_n1821_;
  assign new_n1823_ = ~new_n1820_ & new_n1822_;
  assign new_n1824_ = new_n1810_ & ~new_n1814_;
  assign new_n1825_ = ~new_n1820_ & new_n1824_;
  assign new_n1826_ = ~pv133_9_ & pv133_8_;
  assign new_n1827_ = ~pv133_10_ & new_n1826_;
  assign new_n1828_ = ~pv133_1_ & ~pv133_7_;
  assign new_n1829_ = ~pv133_9_ & new_n1828_;
  assign new_n1830_ = ~pv133_10_ & new_n1829_;
  assign new_n1831_ = ~pv133_10_ & ~new_n1814_;
  assign new_n1832_ = ~new_n1827_ & new_n1831_;
  assign new_n1833_ = ~new_n1810_ & new_n1832_;
  assign new_n1834_ = pv52_0_ & new_n1833_;
  assign new_n1835_ = new_n1830_ & new_n1834_;
  assign new_n1836_ = ~pv133_2_ & new_n1073_;
  assign new_n1837_ = ~pv133_10_ & new_n1836_;
  assign new_n1838_ = ~new_n1810_ & ~new_n1814_;
  assign new_n1839_ = ~new_n1837_ & new_n1838_;
  assign new_n1840_ = ~new_n1827_ & new_n1839_;
  assign new_n1841_ = pv116_2_ & new_n1840_;
  assign new_n1842_ = pv133_9_ & new_n1841_;
  assign new_n1843_ = ~pv133_10_ & new_n1842_;
  assign new_n1844_ = ~pv133_10_ & new_n1843_;
  assign new_n1845_ = ~new_n1830_ & new_n1844_;
  assign new_n1846_ = ~new_n1830_ & new_n1838_;
  assign new_n1847_ = ~pv133_10_ & new_n1846_;
  assign new_n1848_ = pv52_0_ & new_n1847_;
  assign new_n1849_ = ~new_n1827_ & new_n1848_;
  assign new_n1850_ = new_n1837_ & new_n1849_;
  assign new_n1851_ = new_n1814_ & ~new_n1820_;
  assign new_n1852_ = ~new_n1823_ & ~new_n1825_;
  assign new_n1853_ = ~new_n1835_ & new_n1852_;
  assign new_n1854_ = ~new_n1845_ & ~new_n1850_;
  assign new_n1855_ = ~new_n1851_ & new_n1854_;
  assign pv136_1_ = ~new_n1853_ | ~new_n1855_;
  assign new_n1857_ = pv47_7_ & ~new_n240_;
  assign new_n1858_ = pv15_6_ & new_n265_;
  assign new_n1859_ = ~new_n1746_ & ~new_n1857_;
  assign new_n1860_ = ~new_n272_ & ~new_n1858_;
  assign new_n1861_ = new_n1859_ & new_n1860_;
  assign new_n1862_ = new_n517_ & ~new_n1861_;
  assign new_n1863_ = new_n520_ & ~new_n1861_;
  assign new_n1864_ = new_n522_ & ~new_n1861_;
  assign new_n1865_ = pv116_7_ & new_n526_;
  assign new_n1866_ = ~pv133_10_ & new_n1865_;
  assign new_n1867_ = ~new_n1862_ & ~new_n1863_;
  assign new_n1868_ = ~new_n1864_ & ~new_n1866_;
  assign pv142_4_ = ~new_n1867_ | ~new_n1868_;
  assign new_n1870_ = pv84_11_ & new_n241_;
  assign new_n1871_ = pv84_19_ & ~new_n240_;
  assign new_n1872_ = pv84_4_ & new_n265_;
  assign new_n1873_ = pv84_8_ & new_n268_;
  assign new_n1874_ = ~new_n272_ & ~new_n1873_;
  assign new_n1875_ = ~new_n1870_ & ~new_n1871_;
  assign new_n1876_ = ~new_n1872_ & new_n1875_;
  assign new_n1877_ = new_n1874_ & new_n1876_;
  assign new_n1878_ = new_n351_ & ~new_n1877_;
  assign new_n1879_ = new_n354_ & ~new_n1877_;
  assign new_n1880_ = new_n360_ & ~new_n1877_;
  assign new_n1881_ = ~new_n333_ & new_n1880_;
  assign new_n1882_ = pv133_10_ & new_n1881_;
  assign new_n1883_ = new_n366_ & ~new_n1877_;
  assign new_n1884_ = new_n357_ & new_n1883_;
  assign new_n1885_ = pv116_19_ & new_n370_;
  assign new_n1886_ = pv133_9_ & new_n1885_;
  assign new_n1887_ = ~pv133_10_ & new_n1886_;
  assign new_n1888_ = ~new_n336_ & new_n1887_;
  assign new_n1889_ = ~new_n357_ & new_n1888_;
  assign new_n1890_ = new_n376_ & ~new_n1877_;
  assign new_n1891_ = new_n340_ & ~new_n1877_;
  assign new_n1892_ = ~new_n1878_ & ~new_n1879_;
  assign new_n1893_ = ~new_n1882_ & ~new_n1884_;
  assign new_n1894_ = new_n1892_ & new_n1893_;
  assign new_n1895_ = ~new_n1889_ & ~new_n1890_;
  assign new_n1896_ = ~new_n1891_ & new_n1895_;
  assign pv197_19_ = ~new_n1894_ | ~new_n1896_;
  assign new_n1898_ = pv84_18_ & new_n241_;
  assign new_n1899_ = pv84_26_ & ~new_n240_;
  assign new_n1900_ = pv84_11_ & new_n265_;
  assign new_n1901_ = pv84_15_ & new_n268_;
  assign new_n1902_ = ~new_n272_ & ~new_n1901_;
  assign new_n1903_ = ~new_n1898_ & ~new_n1899_;
  assign new_n1904_ = ~new_n1900_ & new_n1903_;
  assign new_n1905_ = new_n1902_ & new_n1904_;
  assign new_n1906_ = new_n351_ & ~new_n1905_;
  assign new_n1907_ = new_n354_ & ~new_n1905_;
  assign new_n1908_ = new_n360_ & ~new_n1905_;
  assign new_n1909_ = ~new_n333_ & new_n1908_;
  assign new_n1910_ = pv133_10_ & new_n1909_;
  assign new_n1911_ = new_n366_ & ~new_n1905_;
  assign new_n1912_ = new_n357_ & new_n1911_;
  assign new_n1913_ = pv116_26_ & new_n370_;
  assign new_n1914_ = pv133_9_ & new_n1913_;
  assign new_n1915_ = ~pv133_10_ & new_n1914_;
  assign new_n1916_ = ~new_n336_ & new_n1915_;
  assign new_n1917_ = ~new_n357_ & new_n1916_;
  assign new_n1918_ = new_n376_ & ~new_n1905_;
  assign new_n1919_ = new_n340_ & ~new_n1905_;
  assign new_n1920_ = ~new_n1906_ & ~new_n1907_;
  assign new_n1921_ = ~new_n1910_ & ~new_n1912_;
  assign new_n1922_ = new_n1920_ & new_n1921_;
  assign new_n1923_ = ~new_n1917_ & ~new_n1918_;
  assign new_n1924_ = ~new_n1919_ & new_n1923_;
  assign pv197_26_ = ~new_n1922_ | ~new_n1924_;
  assign new_n1926_ = pv84_23_ & new_n475_;
  assign new_n1927_ = pv84_23_ & new_n474_;
  assign new_n1928_ = pv84_23_ & new_n489_;
  assign new_n1929_ = pv116_6_ & new_n493_;
  assign new_n1930_ = pv133_9_ & new_n1929_;
  assign new_n1931_ = ~pv133_10_ & new_n1930_;
  assign new_n1932_ = ~new_n1928_ & ~new_n1931_;
  assign new_n1933_ = ~new_n1926_ & ~new_n1927_;
  assign new_n1934_ = ~new_n487_ & new_n1933_;
  assign pv212_6_ = ~new_n1932_ | ~new_n1934_;
  assign new_n1936_ = pv133_1_ & ~pv133_9_;
  assign new_n1937_ = pv133_2_ & new_n1936_;
  assign new_n1938_ = ~pv133_10_ & new_n1937_;
  assign new_n1939_ = ~pv133_10_ & new_n277_;
  assign new_n1940_ = new_n1938_ & ~new_n1939_;
  assign new_n1941_ = pv121_17_ & new_n1939_;
  assign new_n1942_ = pv133_10_ & ~new_n1938_;
  assign new_n1943_ = ~new_n1939_ & new_n1942_;
  assign new_n1944_ = pv122_0_ & new_n1943_;
  assign new_n1945_ = ~new_n1940_ & ~new_n1941_;
  assign pv214_0_ = new_n1944_ | ~new_n1945_;
  assign new_n1947_ = ~new_n1810_ & new_n1827_;
  assign new_n1948_ = ~pv133_10_ & new_n1947_;
  assign new_n1949_ = ~new_n1814_ & new_n1948_;
  assign new_n1950_ = pv50_0_ & new_n1949_;
  assign new_n1951_ = pv47_1_ & ~new_n240_;
  assign new_n1952_ = pv84_1_ & new_n268_;
  assign new_n1953_ = pv15_0_ & new_n265_;
  assign new_n1954_ = ~new_n1951_ & ~new_n1952_;
  assign new_n1955_ = ~new_n272_ & ~new_n1953_;
  assign new_n1956_ = new_n1954_ & new_n1955_;
  assign new_n1957_ = new_n1822_ & ~new_n1956_;
  assign new_n1958_ = pv51_0_ & new_n1847_;
  assign new_n1959_ = ~new_n1827_ & new_n1958_;
  assign new_n1960_ = new_n1837_ & new_n1959_;
  assign new_n1961_ = pv51_0_ & new_n1833_;
  assign new_n1962_ = new_n1830_ & new_n1961_;
  assign new_n1963_ = pv116_1_ & new_n1840_;
  assign new_n1964_ = pv133_9_ & new_n1963_;
  assign new_n1965_ = ~pv133_10_ & new_n1964_;
  assign new_n1966_ = ~pv133_10_ & new_n1965_;
  assign new_n1967_ = ~new_n1830_ & new_n1966_;
  assign new_n1968_ = new_n1824_ & ~new_n1956_;
  assign new_n1969_ = new_n1814_ & ~new_n1956_;
  assign new_n1970_ = ~new_n1950_ & ~new_n1957_;
  assign new_n1971_ = ~new_n1960_ & ~new_n1962_;
  assign new_n1972_ = new_n1970_ & new_n1971_;
  assign new_n1973_ = ~new_n1967_ & ~new_n1968_;
  assign new_n1974_ = ~new_n1969_ & new_n1973_;
  assign pv136_0_ = ~new_n1972_ | ~new_n1974_;
  assign new_n1976_ = pv47_0_ & new_n241_;
  assign new_n1977_ = pv47_8_ & ~new_n240_;
  assign new_n1978_ = pv15_7_ & new_n265_;
  assign new_n1979_ = ~new_n1976_ & ~new_n1977_;
  assign new_n1980_ = ~new_n1978_ & new_n1979_;
  assign new_n1981_ = new_n1874_ & new_n1980_;
  assign new_n1982_ = new_n517_ & ~new_n1981_;
  assign new_n1983_ = new_n520_ & ~new_n1981_;
  assign new_n1984_ = new_n522_ & ~new_n1981_;
  assign new_n1985_ = pv116_8_ & new_n526_;
  assign new_n1986_ = ~pv133_10_ & new_n1985_;
  assign new_n1987_ = ~new_n1982_ & ~new_n1983_;
  assign new_n1988_ = ~new_n1984_ & ~new_n1986_;
  assign pv142_5_ = ~new_n1987_ | ~new_n1988_;
  assign new_n1990_ = pv84_4_ & new_n241_;
  assign new_n1991_ = pv84_12_ & ~new_n240_;
  assign new_n1992_ = pv47_29_ & new_n265_;
  assign new_n1993_ = ~new_n272_ & ~new_n1952_;
  assign new_n1994_ = ~new_n1990_ & ~new_n1991_;
  assign new_n1995_ = ~new_n1992_ & new_n1994_;
  assign new_n1996_ = new_n1993_ & new_n1995_;
  assign new_n1997_ = new_n351_ & ~new_n1996_;
  assign new_n1998_ = new_n354_ & ~new_n1996_;
  assign new_n1999_ = new_n360_ & ~new_n1996_;
  assign new_n2000_ = ~new_n333_ & new_n1999_;
  assign new_n2001_ = pv133_10_ & new_n2000_;
  assign new_n2002_ = new_n366_ & ~new_n1996_;
  assign new_n2003_ = new_n357_ & new_n2002_;
  assign new_n2004_ = pv116_12_ & new_n370_;
  assign new_n2005_ = pv133_9_ & new_n2004_;
  assign new_n2006_ = ~pv133_10_ & new_n2005_;
  assign new_n2007_ = ~new_n336_ & new_n2006_;
  assign new_n2008_ = ~new_n357_ & new_n2007_;
  assign new_n2009_ = new_n376_ & ~new_n1996_;
  assign new_n2010_ = new_n340_ & ~new_n1996_;
  assign new_n2011_ = ~new_n1997_ & ~new_n1998_;
  assign new_n2012_ = ~new_n2001_ & ~new_n2003_;
  assign new_n2013_ = new_n2011_ & new_n2012_;
  assign new_n2014_ = ~new_n2008_ & ~new_n2009_;
  assign new_n2015_ = ~new_n2010_ & new_n2014_;
  assign pv197_12_ = ~new_n2013_ | ~new_n2015_;
  assign new_n2017_ = pv84_17_ & new_n241_;
  assign new_n2018_ = pv84_25_ & ~new_n240_;
  assign new_n2019_ = pv84_10_ & new_n265_;
  assign new_n2020_ = pv84_14_ & new_n268_;
  assign new_n2021_ = ~new_n272_ & ~new_n2020_;
  assign new_n2022_ = ~new_n2017_ & ~new_n2018_;
  assign new_n2023_ = ~new_n2019_ & new_n2022_;
  assign new_n2024_ = new_n2021_ & new_n2023_;
  assign new_n2025_ = new_n351_ & ~new_n2024_;
  assign new_n2026_ = new_n354_ & ~new_n2024_;
  assign new_n2027_ = new_n360_ & ~new_n2024_;
  assign new_n2028_ = ~new_n333_ & new_n2027_;
  assign new_n2029_ = pv133_10_ & new_n2028_;
  assign new_n2030_ = new_n366_ & ~new_n2024_;
  assign new_n2031_ = new_n357_ & new_n2030_;
  assign new_n2032_ = pv116_25_ & new_n370_;
  assign new_n2033_ = pv133_9_ & new_n2032_;
  assign new_n2034_ = ~pv133_10_ & new_n2033_;
  assign new_n2035_ = ~new_n336_ & new_n2034_;
  assign new_n2036_ = ~new_n357_ & new_n2035_;
  assign new_n2037_ = new_n376_ & ~new_n2024_;
  assign new_n2038_ = new_n340_ & ~new_n2024_;
  assign new_n2039_ = ~new_n2025_ & ~new_n2026_;
  assign new_n2040_ = ~new_n2029_ & ~new_n2031_;
  assign new_n2041_ = new_n2039_ & new_n2040_;
  assign new_n2042_ = ~new_n2036_ & ~new_n2037_;
  assign new_n2043_ = ~new_n2038_ & new_n2042_;
  assign pv197_25_ = ~new_n2041_ | ~new_n2043_;
  assign new_n2045_ = pv84_22_ & new_n241_;
  assign new_n2046_ = pv84_30_ & ~new_n240_;
  assign new_n2047_ = pv84_15_ & new_n265_;
  assign new_n2048_ = pv84_19_ & new_n268_;
  assign new_n2049_ = ~new_n272_ & ~new_n2048_;
  assign new_n2050_ = ~new_n2045_ & ~new_n2046_;
  assign new_n2051_ = ~new_n2047_ & new_n2050_;
  assign new_n2052_ = new_n2049_ & new_n2051_;
  assign new_n2053_ = new_n351_ & ~new_n2052_;
  assign new_n2054_ = new_n354_ & ~new_n2052_;
  assign new_n2055_ = new_n360_ & ~new_n2052_;
  assign new_n2056_ = ~new_n333_ & new_n2055_;
  assign new_n2057_ = pv133_10_ & new_n2056_;
  assign new_n2058_ = new_n366_ & ~new_n2052_;
  assign new_n2059_ = new_n357_ & new_n2058_;
  assign new_n2060_ = pv116_30_ & new_n370_;
  assign new_n2061_ = pv133_9_ & new_n2060_;
  assign new_n2062_ = ~pv133_10_ & new_n2061_;
  assign new_n2063_ = ~new_n336_ & new_n2062_;
  assign new_n2064_ = ~new_n357_ & new_n2063_;
  assign new_n2065_ = new_n376_ & ~new_n2052_;
  assign new_n2066_ = new_n340_ & ~new_n2052_;
  assign new_n2067_ = ~new_n2053_ & ~new_n2054_;
  assign new_n2068_ = ~new_n2057_ & ~new_n2059_;
  assign new_n2069_ = new_n2067_ & new_n2068_;
  assign new_n2070_ = ~new_n2064_ & ~new_n2065_;
  assign new_n2071_ = ~new_n2066_ & new_n2070_;
  assign pv197_30_ = ~new_n2069_ | ~new_n2071_;
  assign new_n2073_ = pv84_18_ & new_n475_;
  assign new_n2074_ = pv84_18_ & new_n474_;
  assign new_n2075_ = pv84_18_ & new_n489_;
  assign new_n2076_ = pv116_1_ & new_n493_;
  assign new_n2077_ = pv133_9_ & new_n2076_;
  assign new_n2078_ = ~pv133_10_ & new_n2077_;
  assign new_n2079_ = ~new_n2075_ & ~new_n2078_;
  assign new_n2080_ = ~new_n2073_ & ~new_n2074_;
  assign new_n2081_ = ~new_n487_ & new_n2080_;
  assign pv212_1_ = ~new_n2079_ | ~new_n2081_;
  assign new_n2083_ = pv84_27_ & new_n475_;
  assign new_n2084_ = pv84_27_ & new_n474_;
  assign new_n2085_ = pv84_27_ & new_n489_;
  assign new_n2086_ = pv116_10_ & new_n493_;
  assign new_n2087_ = pv133_9_ & new_n2086_;
  assign new_n2088_ = ~pv133_10_ & new_n2087_;
  assign new_n2089_ = ~new_n2085_ & ~new_n2088_;
  assign new_n2090_ = ~new_n2083_ & ~new_n2084_;
  assign new_n2091_ = ~new_n487_ & new_n2090_;
  assign pv212_10_ = ~new_n2089_ | ~new_n2091_;
  assign new_n2093_ = pv84_5_ & new_n241_;
  assign new_n2094_ = pv84_13_ & ~new_n240_;
  assign new_n2095_ = pv47_30_ & new_n265_;
  assign new_n2096_ = ~new_n272_ & ~new_n1816_;
  assign new_n2097_ = ~new_n2093_ & ~new_n2094_;
  assign new_n2098_ = ~new_n2095_ & new_n2097_;
  assign new_n2099_ = new_n2096_ & new_n2098_;
  assign new_n2100_ = new_n351_ & ~new_n2099_;
  assign new_n2101_ = new_n354_ & ~new_n2099_;
  assign new_n2102_ = new_n360_ & ~new_n2099_;
  assign new_n2103_ = ~new_n333_ & new_n2102_;
  assign new_n2104_ = pv133_10_ & new_n2103_;
  assign new_n2105_ = new_n366_ & ~new_n2099_;
  assign new_n2106_ = new_n357_ & new_n2105_;
  assign new_n2107_ = pv116_13_ & new_n370_;
  assign new_n2108_ = pv133_9_ & new_n2107_;
  assign new_n2109_ = ~pv133_10_ & new_n2108_;
  assign new_n2110_ = ~new_n336_ & new_n2109_;
  assign new_n2111_ = ~new_n357_ & new_n2110_;
  assign new_n2112_ = new_n376_ & ~new_n2099_;
  assign new_n2113_ = new_n340_ & ~new_n2099_;
  assign new_n2114_ = ~new_n2100_ & ~new_n2101_;
  assign new_n2115_ = ~new_n2104_ & ~new_n2106_;
  assign new_n2116_ = new_n2114_ & new_n2115_;
  assign new_n2117_ = ~new_n2111_ & ~new_n2112_;
  assign new_n2118_ = ~new_n2113_ & new_n2117_;
  assign pv197_13_ = ~new_n2116_ | ~new_n2118_;
  assign new_n2120_ = pv84_16_ & new_n241_;
  assign new_n2121_ = pv84_24_ & ~new_n240_;
  assign new_n2122_ = pv84_9_ & new_n265_;
  assign new_n2123_ = pv84_13_ & new_n268_;
  assign new_n2124_ = ~new_n272_ & ~new_n2123_;
  assign new_n2125_ = ~new_n2120_ & ~new_n2121_;
  assign new_n2126_ = ~new_n2122_ & new_n2125_;
  assign new_n2127_ = new_n2124_ & new_n2126_;
  assign new_n2128_ = new_n351_ & ~new_n2127_;
  assign new_n2129_ = new_n354_ & ~new_n2127_;
  assign new_n2130_ = new_n360_ & ~new_n2127_;
  assign new_n2131_ = ~new_n333_ & new_n2130_;
  assign new_n2132_ = pv133_10_ & new_n2131_;
  assign new_n2133_ = new_n366_ & ~new_n2127_;
  assign new_n2134_ = new_n357_ & new_n2133_;
  assign new_n2135_ = pv116_24_ & new_n370_;
  assign new_n2136_ = pv133_9_ & new_n2135_;
  assign new_n2137_ = ~pv133_10_ & new_n2136_;
  assign new_n2138_ = ~new_n336_ & new_n2137_;
  assign new_n2139_ = ~new_n357_ & new_n2138_;
  assign new_n2140_ = new_n376_ & ~new_n2127_;
  assign new_n2141_ = new_n340_ & ~new_n2127_;
  assign new_n2142_ = ~new_n2128_ & ~new_n2129_;
  assign new_n2143_ = ~new_n2132_ & ~new_n2134_;
  assign new_n2144_ = new_n2142_ & new_n2143_;
  assign new_n2145_ = ~new_n2139_ & ~new_n2140_;
  assign new_n2146_ = ~new_n2141_ & new_n2145_;
  assign pv197_24_ = ~new_n2144_ | ~new_n2146_;
  assign new_n2148_ = pv84_23_ & new_n241_;
  assign new_n2149_ = pv84_31_ & ~new_n240_;
  assign new_n2150_ = pv84_16_ & new_n265_;
  assign new_n2151_ = pv84_20_ & new_n268_;
  assign new_n2152_ = ~new_n272_ & ~new_n2151_;
  assign new_n2153_ = ~new_n2148_ & ~new_n2149_;
  assign new_n2154_ = ~new_n2150_ & new_n2153_;
  assign new_n2155_ = new_n2152_ & new_n2154_;
  assign new_n2156_ = new_n351_ & ~new_n2155_;
  assign new_n2157_ = new_n354_ & ~new_n2155_;
  assign new_n2158_ = new_n360_ & ~new_n2155_;
  assign new_n2159_ = ~new_n333_ & new_n2158_;
  assign new_n2160_ = pv133_10_ & new_n2159_;
  assign new_n2161_ = new_n366_ & ~new_n2155_;
  assign new_n2162_ = new_n357_ & new_n2161_;
  assign new_n2163_ = pv116_31_ & new_n370_;
  assign new_n2164_ = pv133_9_ & new_n2163_;
  assign new_n2165_ = ~pv133_10_ & new_n2164_;
  assign new_n2166_ = ~new_n336_ & new_n2165_;
  assign new_n2167_ = ~new_n357_ & new_n2166_;
  assign new_n2168_ = new_n376_ & ~new_n2155_;
  assign new_n2169_ = new_n340_ & ~new_n2155_;
  assign new_n2170_ = ~new_n2156_ & ~new_n2157_;
  assign new_n2171_ = ~new_n2160_ & ~new_n2162_;
  assign new_n2172_ = new_n2170_ & new_n2171_;
  assign new_n2173_ = ~new_n2167_ & ~new_n2168_;
  assign new_n2174_ = ~new_n2169_ & new_n2173_;
  assign pv197_31_ = ~new_n2172_ | ~new_n2174_;
  assign new_n2176_ = pv84_17_ & new_n475_;
  assign new_n2177_ = pv84_17_ & new_n474_;
  assign new_n2178_ = pv84_17_ & new_n489_;
  assign new_n2179_ = pv116_0_ & new_n493_;
  assign new_n2180_ = pv133_9_ & new_n2179_;
  assign new_n2181_ = ~pv133_10_ & new_n2180_;
  assign new_n2182_ = ~new_n2178_ & ~new_n2181_;
  assign new_n2183_ = ~new_n2176_ & ~new_n2177_;
  assign new_n2184_ = ~new_n487_ & new_n2183_;
  assign pv212_0_ = ~new_n2182_ | ~new_n2184_;
  assign new_n2186_ = pv84_28_ & new_n475_;
  assign new_n2187_ = pv84_28_ & new_n474_;
  assign new_n2188_ = pv84_28_ & new_n489_;
  assign new_n2189_ = pv116_11_ & new_n493_;
  assign new_n2190_ = pv133_9_ & new_n2189_;
  assign new_n2191_ = ~pv133_10_ & new_n2190_;
  assign new_n2192_ = ~new_n2188_ & ~new_n2191_;
  assign new_n2193_ = ~new_n2186_ & ~new_n2187_;
  assign new_n2194_ = ~new_n487_ & new_n2193_;
  assign pv212_11_ = ~new_n2192_ | ~new_n2194_;
  assign new_n2196_ = pv84_6_ & new_n241_;
  assign new_n2197_ = pv84_14_ & ~new_n240_;
  assign new_n2198_ = pv47_31_ & new_n265_;
  assign new_n2199_ = ~new_n272_ & ~new_n512_;
  assign new_n2200_ = ~new_n2196_ & ~new_n2197_;
  assign new_n2201_ = ~new_n2198_ & new_n2200_;
  assign new_n2202_ = new_n2199_ & new_n2201_;
  assign new_n2203_ = new_n351_ & ~new_n2202_;
  assign new_n2204_ = new_n354_ & ~new_n2202_;
  assign new_n2205_ = new_n360_ & ~new_n2202_;
  assign new_n2206_ = ~new_n333_ & new_n2205_;
  assign new_n2207_ = pv133_10_ & new_n2206_;
  assign new_n2208_ = new_n366_ & ~new_n2202_;
  assign new_n2209_ = new_n357_ & new_n2208_;
  assign new_n2210_ = pv116_14_ & new_n370_;
  assign new_n2211_ = pv133_9_ & new_n2210_;
  assign new_n2212_ = ~pv133_10_ & new_n2211_;
  assign new_n2213_ = ~new_n336_ & new_n2212_;
  assign new_n2214_ = ~new_n357_ & new_n2213_;
  assign new_n2215_ = new_n376_ & ~new_n2202_;
  assign new_n2216_ = new_n340_ & ~new_n2202_;
  assign new_n2217_ = ~new_n2203_ & ~new_n2204_;
  assign new_n2218_ = ~new_n2207_ & ~new_n2209_;
  assign new_n2219_ = new_n2217_ & new_n2218_;
  assign new_n2220_ = ~new_n2214_ & ~new_n2215_;
  assign new_n2221_ = ~new_n2216_ & new_n2220_;
  assign pv197_14_ = ~new_n2219_ | ~new_n2221_;
  assign new_n2223_ = pv84_15_ & new_n241_;
  assign new_n2224_ = pv84_23_ & ~new_n240_;
  assign new_n2225_ = pv84_8_ & new_n265_;
  assign new_n2226_ = pv84_12_ & new_n268_;
  assign new_n2227_ = ~new_n272_ & ~new_n2226_;
  assign new_n2228_ = ~new_n2223_ & ~new_n2224_;
  assign new_n2229_ = ~new_n2225_ & new_n2228_;
  assign new_n2230_ = new_n2227_ & new_n2229_;
  assign new_n2231_ = new_n351_ & ~new_n2230_;
  assign new_n2232_ = new_n354_ & ~new_n2230_;
  assign new_n2233_ = new_n360_ & ~new_n2230_;
  assign new_n2234_ = ~new_n333_ & new_n2233_;
  assign new_n2235_ = pv133_10_ & new_n2234_;
  assign new_n2236_ = new_n366_ & ~new_n2230_;
  assign new_n2237_ = new_n357_ & new_n2236_;
  assign new_n2238_ = pv116_23_ & new_n370_;
  assign new_n2239_ = pv133_9_ & new_n2238_;
  assign new_n2240_ = ~pv133_10_ & new_n2239_;
  assign new_n2241_ = ~new_n336_ & new_n2240_;
  assign new_n2242_ = ~new_n357_ & new_n2241_;
  assign new_n2243_ = new_n376_ & ~new_n2230_;
  assign new_n2244_ = new_n340_ & ~new_n2230_;
  assign new_n2245_ = ~new_n2231_ & ~new_n2232_;
  assign new_n2246_ = ~new_n2235_ & ~new_n2237_;
  assign new_n2247_ = new_n2245_ & new_n2246_;
  assign new_n2248_ = ~new_n2242_ & ~new_n2243_;
  assign new_n2249_ = ~new_n2244_ & new_n2248_;
  assign pv197_23_ = ~new_n2247_ | ~new_n2249_;
  assign new_n2251_ = pv84_20_ & new_n475_;
  assign new_n2252_ = pv84_20_ & new_n474_;
  assign new_n2253_ = pv84_20_ & new_n489_;
  assign new_n2254_ = pv116_3_ & new_n493_;
  assign new_n2255_ = pv133_9_ & new_n2254_;
  assign new_n2256_ = ~pv133_10_ & new_n2255_;
  assign new_n2257_ = ~new_n2253_ & ~new_n2256_;
  assign new_n2258_ = ~new_n2251_ & ~new_n2252_;
  assign new_n2259_ = ~new_n487_ & new_n2258_;
  assign pv212_3_ = ~new_n2257_ | ~new_n2259_;
  assign new_n2261_ = ~pv133_8_ & new_n277_;
  assign new_n2262_ = ~pv133_10_ & new_n2261_;
  assign new_n2263_ = ~pv133_10_ & new_n238_;
  assign new_n2264_ = ~new_n2262_ & ~new_n2263_;
  assign new_n2265_ = ~pv133_10_ & new_n2264_;
  assign new_n2266_ = ~new_n287_ & new_n2265_;
  assign new_n2267_ = ~new_n1830_ & new_n2266_;
  assign new_n2268_ = ~new_n1827_ & new_n2267_;
  assign new_n2269_ = pv121_16_ & new_n2262_;
  assign new_n2270_ = pv133_10_ & ~new_n287_;
  assign new_n2271_ = ~new_n2263_ & new_n2270_;
  assign new_n2272_ = ~new_n2262_ & new_n2271_;
  assign new_n2273_ = pv119_0_ & new_n2272_;
  assign new_n2274_ = new_n1830_ & new_n2266_;
  assign new_n2275_ = ~new_n1827_ & new_n2274_;
  assign new_n2276_ = ~pv133_10_ & ~new_n287_;
  assign new_n2277_ = ~new_n2263_ & new_n2276_;
  assign new_n2278_ = ~new_n2262_ & new_n2277_;
  assign new_n2279_ = new_n1827_ & new_n2278_;
  assign new_n2280_ = ~new_n2275_ & ~new_n2279_;
  assign new_n2281_ = ~new_n2268_ & ~new_n2269_;
  assign new_n2282_ = ~new_n2273_ & new_n2281_;
  assign pv213_0_ = ~new_n2280_ | ~new_n2282_;
  assign new_n2284_ = pv84_7_ & new_n241_;
  assign new_n2285_ = pv84_15_ & ~new_n240_;
  assign new_n2286_ = pv84_0_ & new_n265_;
  assign new_n2287_ = ~new_n272_ & ~new_n1554_;
  assign new_n2288_ = ~new_n2284_ & ~new_n2285_;
  assign new_n2289_ = ~new_n2286_ & new_n2288_;
  assign new_n2290_ = new_n2287_ & new_n2289_;
  assign new_n2291_ = new_n351_ & ~new_n2290_;
  assign new_n2292_ = new_n354_ & ~new_n2290_;
  assign new_n2293_ = new_n360_ & ~new_n2290_;
  assign new_n2294_ = ~new_n333_ & new_n2293_;
  assign new_n2295_ = pv133_10_ & new_n2294_;
  assign new_n2296_ = new_n366_ & ~new_n2290_;
  assign new_n2297_ = new_n357_ & new_n2296_;
  assign new_n2298_ = pv116_15_ & new_n370_;
  assign new_n2299_ = pv133_9_ & new_n2298_;
  assign new_n2300_ = ~pv133_10_ & new_n2299_;
  assign new_n2301_ = ~new_n336_ & new_n2300_;
  assign new_n2302_ = ~new_n357_ & new_n2301_;
  assign new_n2303_ = new_n376_ & ~new_n2290_;
  assign new_n2304_ = new_n340_ & ~new_n2290_;
  assign new_n2305_ = ~new_n2291_ & ~new_n2292_;
  assign new_n2306_ = ~new_n2295_ & ~new_n2297_;
  assign new_n2307_ = new_n2305_ & new_n2306_;
  assign new_n2308_ = ~new_n2302_ & ~new_n2303_;
  assign new_n2309_ = ~new_n2304_ & new_n2308_;
  assign pv197_15_ = ~new_n2307_ | ~new_n2309_;
  assign new_n2311_ = pv84_14_ & new_n241_;
  assign new_n2312_ = pv84_22_ & ~new_n240_;
  assign new_n2313_ = pv84_7_ & new_n265_;
  assign new_n2314_ = ~new_n2311_ & ~new_n2312_;
  assign new_n2315_ = ~new_n2313_ & new_n2314_;
  assign new_n2316_ = new_n995_ & new_n2315_;
  assign new_n2317_ = new_n351_ & ~new_n2316_;
  assign new_n2318_ = new_n354_ & ~new_n2316_;
  assign new_n2319_ = new_n360_ & ~new_n2316_;
  assign new_n2320_ = ~new_n333_ & new_n2319_;
  assign new_n2321_ = pv133_10_ & new_n2320_;
  assign new_n2322_ = new_n366_ & ~new_n2316_;
  assign new_n2323_ = new_n357_ & new_n2322_;
  assign new_n2324_ = pv116_22_ & new_n370_;
  assign new_n2325_ = pv133_9_ & new_n2324_;
  assign new_n2326_ = ~pv133_10_ & new_n2325_;
  assign new_n2327_ = ~new_n336_ & new_n2326_;
  assign new_n2328_ = ~new_n357_ & new_n2327_;
  assign new_n2329_ = new_n376_ & ~new_n2316_;
  assign new_n2330_ = new_n340_ & ~new_n2316_;
  assign new_n2331_ = ~new_n2317_ & ~new_n2318_;
  assign new_n2332_ = ~new_n2321_ & ~new_n2323_;
  assign new_n2333_ = new_n2331_ & new_n2332_;
  assign new_n2334_ = ~new_n2328_ & ~new_n2329_;
  assign new_n2335_ = ~new_n2330_ & new_n2334_;
  assign pv197_22_ = ~new_n2333_ | ~new_n2335_;
  assign new_n2337_ = pv84_19_ & new_n475_;
  assign new_n2338_ = pv84_19_ & new_n474_;
  assign new_n2339_ = pv84_19_ & new_n489_;
  assign new_n2340_ = pv116_2_ & new_n493_;
  assign new_n2341_ = pv133_9_ & new_n2340_;
  assign new_n2342_ = ~pv133_10_ & new_n2341_;
  assign new_n2343_ = ~new_n2339_ & ~new_n2342_;
  assign new_n2344_ = ~new_n2337_ & ~new_n2338_;
  assign new_n2345_ = ~new_n487_ & new_n2344_;
  assign pv212_2_ = ~new_n2343_ | ~new_n2345_;
endmodule

