module top ( 
    ic3_35_, ic7_39_, id4_4_, id22_22_, id26_26_, id21_21_, id27_27_,
    id29_29_, ic4_36_, id5_5_, id20_20_, id28_28_, ic6_38_, id6_6_,
    id17_17_, id31_31_, id18_18_, id23_23_, id25_25_, id30_30_, ic0_32_,
    id7_7_, id19_19_, id24_24_, ic1_33_, ic5_37_, r_40_, id0_0_, id8_8_,
    id14_14_, id16_16_, id1_1_, id9_9_, id15_15_, ic2_34_, id2_2_,
    id13_13_, id10_10_, id12_12_, id3_3_, id11_11_,
    od10_232_, od11_231_, od12_230_, od4_238_, od8_234_, od1_241_,
    od20_222_, od21_221_, od22_220_, od5_237_, od9_233_, od2_240_,
    od23_219_, od24_218_, od25_217_, od26_216_, od27_215_, od28_214_,
    od29_213_, od30_212_, od31_211_, od6_236_, od13_229_, od14_228_,
    od15_227_, od16_226_, od17_225_, od18_224_, od19_223_, od3_239_,
    od7_235_, od0_242_  );
  input  ic3_35_, ic7_39_, id4_4_, id22_22_, id26_26_, id21_21_,
    id27_27_, id29_29_, ic4_36_, id5_5_, id20_20_, id28_28_, ic6_38_,
    id6_6_, id17_17_, id31_31_, id18_18_, id23_23_, id25_25_, id30_30_,
    ic0_32_, id7_7_, id19_19_, id24_24_, ic1_33_, ic5_37_, r_40_, id0_0_,
    id8_8_, id14_14_, id16_16_, id1_1_, id9_9_, id15_15_, ic2_34_, id2_2_,
    id13_13_, id10_10_, id12_12_, id3_3_, id11_11_;
  output od10_232_, od11_231_, od12_230_, od4_238_, od8_234_, od1_241_,
    od20_222_, od21_221_, od22_220_, od5_237_, od9_233_, od2_240_,
    od23_219_, od24_218_, od25_217_, od26_216_, od27_215_, od28_214_,
    od29_213_, od30_212_, od31_211_, od6_236_, od13_229_, od14_228_,
    od15_227_, od16_226_, od17_225_, od18_224_, od19_223_, od3_239_,
    od7_235_, od0_242_;
  wire new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_, new_n80_,
    new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_, new_n87_,
    new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_, new_n94_,
    new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_, new_n101_,
    new_n102_, new_n103_, new_n104_, new_n105_, new_n106_, new_n107_,
    new_n108_, new_n109_, new_n110_, new_n111_, new_n112_, new_n113_,
    new_n114_, new_n115_, new_n116_, new_n117_, new_n118_, new_n119_,
    new_n120_, new_n121_, new_n122_, new_n123_, new_n124_, new_n125_,
    new_n126_, new_n127_, new_n128_, new_n129_, new_n130_, new_n131_,
    new_n132_, new_n133_, new_n134_, new_n135_, new_n136_, new_n137_,
    new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n320_, new_n321_, new_n322_, new_n324_, new_n325_,
    new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n339_,
    new_n340_, new_n341_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n372_,
    new_n373_, new_n374_, new_n376_, new_n377_, new_n378_, new_n380_,
    new_n381_, new_n382_, new_n384_, new_n385_, new_n386_, new_n388_,
    new_n389_, new_n390_, new_n392_, new_n393_, new_n394_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n404_, new_n405_, new_n406_, new_n408_, new_n409_, new_n410_,
    new_n412_, new_n413_, new_n414_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n423_, new_n424_, new_n425_,
    new_n427_, new_n428_, new_n429_, new_n431_, new_n432_, new_n433_,
    new_n435_, new_n436_, new_n437_, new_n439_, new_n440_, new_n441_,
    new_n443_, new_n444_, new_n445_, new_n447_, new_n448_, new_n449_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n458_, new_n459_, new_n460_, new_n462_, new_n463_, new_n464_,
    new_n466_, new_n467_, new_n468_, new_n470_, new_n471_, new_n472_,
    new_n474_, new_n475_, new_n476_, new_n478_, new_n479_, new_n480_;
  assign new_n74_ = id14_14_ & ~id15_15_;
  assign new_n75_ = ~id14_14_ & id15_15_;
  assign new_n76_ = ~new_n74_ & ~new_n75_;
  assign new_n77_ = ~id13_13_ & id12_12_;
  assign new_n78_ = id13_13_ & ~id12_12_;
  assign new_n79_ = ~new_n77_ & ~new_n78_;
  assign new_n80_ = new_n76_ & ~new_n79_;
  assign new_n81_ = ~new_n76_ & new_n79_;
  assign new_n82_ = ~new_n80_ & ~new_n81_;
  assign new_n83_ = id6_6_ & ~id7_7_;
  assign new_n84_ = ~id6_6_ & id7_7_;
  assign new_n85_ = ~new_n83_ & ~new_n84_;
  assign new_n86_ = id4_4_ & ~id5_5_;
  assign new_n87_ = ~id4_4_ & id5_5_;
  assign new_n88_ = ~new_n86_ & ~new_n87_;
  assign new_n89_ = new_n85_ & ~new_n88_;
  assign new_n90_ = ~new_n85_ & new_n88_;
  assign new_n91_ = ~new_n89_ & ~new_n90_;
  assign new_n92_ = new_n82_ & ~new_n91_;
  assign new_n93_ = ~new_n82_ & new_n91_;
  assign new_n94_ = ~new_n92_ & ~new_n93_;
  assign new_n95_ = ic7_39_ & r_40_;
  assign new_n96_ = new_n94_ & new_n95_;
  assign new_n97_ = ~new_n94_ & ~new_n95_;
  assign new_n98_ = ~new_n96_ & ~new_n97_;
  assign new_n99_ = id27_27_ & ~id31_31_;
  assign new_n100_ = ~id27_27_ & id31_31_;
  assign new_n101_ = ~new_n99_ & ~new_n100_;
  assign new_n102_ = ~id23_23_ & id19_19_;
  assign new_n103_ = id23_23_ & ~id19_19_;
  assign new_n104_ = ~new_n102_ & ~new_n103_;
  assign new_n105_ = new_n101_ & ~new_n104_;
  assign new_n106_ = ~new_n101_ & new_n104_;
  assign new_n107_ = ~new_n105_ & ~new_n106_;
  assign new_n108_ = new_n98_ & ~new_n107_;
  assign new_n109_ = ~new_n98_ & new_n107_;
  assign new_n110_ = ~new_n108_ & ~new_n109_;
  assign new_n111_ = ~id31_31_ & id30_30_;
  assign new_n112_ = id31_31_ & ~id30_30_;
  assign new_n113_ = ~new_n111_ & ~new_n112_;
  assign new_n114_ = ~id29_29_ & id28_28_;
  assign new_n115_ = id29_29_ & ~id28_28_;
  assign new_n116_ = ~new_n114_ & ~new_n115_;
  assign new_n117_ = new_n113_ & ~new_n116_;
  assign new_n118_ = ~new_n113_ & new_n116_;
  assign new_n119_ = ~new_n117_ & ~new_n118_;
  assign new_n120_ = id22_22_ & ~id23_23_;
  assign new_n121_ = ~id22_22_ & id23_23_;
  assign new_n122_ = ~new_n120_ & ~new_n121_;
  assign new_n123_ = ~id21_21_ & id20_20_;
  assign new_n124_ = id21_21_ & ~id20_20_;
  assign new_n125_ = ~new_n123_ & ~new_n124_;
  assign new_n126_ = new_n122_ & ~new_n125_;
  assign new_n127_ = ~new_n122_ & new_n125_;
  assign new_n128_ = ~new_n126_ & ~new_n127_;
  assign new_n129_ = new_n119_ & ~new_n128_;
  assign new_n130_ = ~new_n119_ & new_n128_;
  assign new_n131_ = ~new_n129_ & ~new_n130_;
  assign new_n132_ = ic3_35_ & r_40_;
  assign new_n133_ = new_n131_ & new_n132_;
  assign new_n134_ = ~new_n131_ & ~new_n132_;
  assign new_n135_ = ~new_n133_ & ~new_n134_;
  assign new_n136_ = ~id15_15_ & id11_11_;
  assign new_n137_ = id15_15_ & ~id11_11_;
  assign new_n138_ = ~new_n136_ & ~new_n137_;
  assign new_n139_ = ~id7_7_ & id3_3_;
  assign new_n140_ = id7_7_ & ~id3_3_;
  assign new_n141_ = ~new_n139_ & ~new_n140_;
  assign new_n142_ = new_n138_ & ~new_n141_;
  assign new_n143_ = ~new_n138_ & new_n141_;
  assign new_n144_ = ~new_n142_ & ~new_n143_;
  assign new_n145_ = new_n135_ & ~new_n144_;
  assign new_n146_ = ~new_n135_ & new_n144_;
  assign new_n147_ = ~new_n145_ & ~new_n146_;
  assign new_n148_ = id26_26_ & ~id27_27_;
  assign new_n149_ = ~id26_26_ & id27_27_;
  assign new_n150_ = ~new_n148_ & ~new_n149_;
  assign new_n151_ = ~id25_25_ & id24_24_;
  assign new_n152_ = id25_25_ & ~id24_24_;
  assign new_n153_ = ~new_n151_ & ~new_n152_;
  assign new_n154_ = new_n150_ & ~new_n153_;
  assign new_n155_ = ~new_n150_ & new_n153_;
  assign new_n156_ = ~new_n154_ & ~new_n155_;
  assign new_n157_ = new_n119_ & ~new_n156_;
  assign new_n158_ = ~new_n119_ & new_n156_;
  assign new_n159_ = ~new_n157_ & ~new_n158_;
  assign new_n160_ = ic1_33_ & r_40_;
  assign new_n161_ = new_n159_ & new_n160_;
  assign new_n162_ = ~new_n159_ & ~new_n160_;
  assign new_n163_ = ~new_n161_ & ~new_n162_;
  assign new_n164_ = id9_9_ & ~id13_13_;
  assign new_n165_ = ~id9_9_ & id13_13_;
  assign new_n166_ = ~new_n164_ & ~new_n165_;
  assign new_n167_ = ~id5_5_ & id1_1_;
  assign new_n168_ = id5_5_ & ~id1_1_;
  assign new_n169_ = ~new_n167_ & ~new_n168_;
  assign new_n170_ = new_n166_ & ~new_n169_;
  assign new_n171_ = ~new_n166_ & new_n169_;
  assign new_n172_ = ~new_n170_ & ~new_n171_;
  assign new_n173_ = new_n163_ & ~new_n172_;
  assign new_n174_ = ~new_n163_ & new_n172_;
  assign new_n175_ = ~new_n173_ & ~new_n174_;
  assign new_n176_ = id18_18_ & ~id19_19_;
  assign new_n177_ = ~id18_18_ & id19_19_;
  assign new_n178_ = ~new_n176_ & ~new_n177_;
  assign new_n179_ = ~id17_17_ & id16_16_;
  assign new_n180_ = id17_17_ & ~id16_16_;
  assign new_n181_ = ~new_n179_ & ~new_n180_;
  assign new_n182_ = new_n178_ & ~new_n181_;
  assign new_n183_ = ~new_n178_ & new_n181_;
  assign new_n184_ = ~new_n182_ & ~new_n183_;
  assign new_n185_ = new_n156_ & ~new_n184_;
  assign new_n186_ = ~new_n156_ & new_n184_;
  assign new_n187_ = ~new_n185_ & ~new_n186_;
  assign new_n188_ = r_40_ & ic2_34_;
  assign new_n189_ = new_n187_ & new_n188_;
  assign new_n190_ = ~new_n187_ & ~new_n188_;
  assign new_n191_ = ~new_n189_ & ~new_n190_;
  assign new_n192_ = ~id14_14_ & id10_10_;
  assign new_n193_ = id14_14_ & ~id10_10_;
  assign new_n194_ = ~new_n192_ & ~new_n193_;
  assign new_n195_ = ~id6_6_ & id2_2_;
  assign new_n196_ = id6_6_ & ~id2_2_;
  assign new_n197_ = ~new_n195_ & ~new_n196_;
  assign new_n198_ = new_n194_ & ~new_n197_;
  assign new_n199_ = ~new_n194_ & new_n197_;
  assign new_n200_ = ~new_n198_ & ~new_n199_;
  assign new_n201_ = new_n191_ & ~new_n200_;
  assign new_n202_ = ~new_n191_ & new_n200_;
  assign new_n203_ = ~new_n201_ & ~new_n202_;
  assign new_n204_ = new_n128_ & ~new_n184_;
  assign new_n205_ = ~new_n128_ & new_n184_;
  assign new_n206_ = ~new_n204_ & ~new_n205_;
  assign new_n207_ = ic0_32_ & r_40_;
  assign new_n208_ = new_n206_ & new_n207_;
  assign new_n209_ = ~new_n206_ & ~new_n207_;
  assign new_n210_ = ~new_n208_ & ~new_n209_;
  assign new_n211_ = id8_8_ & ~id12_12_;
  assign new_n212_ = ~id8_8_ & id12_12_;
  assign new_n213_ = ~new_n211_ & ~new_n212_;
  assign new_n214_ = ~id4_4_ & id0_0_;
  assign new_n215_ = id4_4_ & ~id0_0_;
  assign new_n216_ = ~new_n214_ & ~new_n215_;
  assign new_n217_ = new_n213_ & ~new_n216_;
  assign new_n218_ = ~new_n213_ & new_n216_;
  assign new_n219_ = ~new_n217_ & ~new_n218_;
  assign new_n220_ = new_n210_ & ~new_n219_;
  assign new_n221_ = ~new_n210_ & new_n219_;
  assign new_n222_ = ~new_n220_ & ~new_n221_;
  assign new_n223_ = new_n147_ & new_n175_;
  assign new_n224_ = new_n203_ & new_n223_;
  assign new_n225_ = ~new_n222_ & new_n224_;
  assign new_n226_ = ~new_n203_ & new_n223_;
  assign new_n227_ = new_n222_ & new_n226_;
  assign new_n228_ = new_n147_ & ~new_n175_;
  assign new_n229_ = new_n203_ & new_n228_;
  assign new_n230_ = new_n222_ & new_n229_;
  assign new_n231_ = ~new_n147_ & new_n175_;
  assign new_n232_ = new_n203_ & new_n231_;
  assign new_n233_ = new_n222_ & new_n232_;
  assign new_n234_ = ~new_n225_ & ~new_n227_;
  assign new_n235_ = ~new_n230_ & new_n234_;
  assign new_n236_ = ~new_n233_ & new_n235_;
  assign new_n237_ = id10_10_ & ~id11_11_;
  assign new_n238_ = ~id10_10_ & id11_11_;
  assign new_n239_ = ~new_n237_ & ~new_n238_;
  assign new_n240_ = id8_8_ & ~id9_9_;
  assign new_n241_ = ~id8_8_ & id9_9_;
  assign new_n242_ = ~new_n240_ & ~new_n241_;
  assign new_n243_ = new_n239_ & ~new_n242_;
  assign new_n244_ = ~new_n239_ & new_n242_;
  assign new_n245_ = ~new_n243_ & ~new_n244_;
  assign new_n246_ = new_n82_ & ~new_n245_;
  assign new_n247_ = ~new_n82_ & new_n245_;
  assign new_n248_ = ~new_n246_ & ~new_n247_;
  assign new_n249_ = ic5_37_ & r_40_;
  assign new_n250_ = new_n248_ & new_n249_;
  assign new_n251_ = ~new_n248_ & ~new_n249_;
  assign new_n252_ = ~new_n250_ & ~new_n251_;
  assign new_n253_ = ~id29_29_ & id25_25_;
  assign new_n254_ = id29_29_ & ~id25_25_;
  assign new_n255_ = ~new_n253_ & ~new_n254_;
  assign new_n256_ = ~id21_21_ & id17_17_;
  assign new_n257_ = id21_21_ & ~id17_17_;
  assign new_n258_ = ~new_n256_ & ~new_n257_;
  assign new_n259_ = new_n255_ & ~new_n258_;
  assign new_n260_ = ~new_n255_ & new_n258_;
  assign new_n261_ = ~new_n259_ & ~new_n260_;
  assign new_n262_ = new_n252_ & ~new_n261_;
  assign new_n263_ = ~new_n252_ & new_n261_;
  assign new_n264_ = ~new_n262_ & ~new_n263_;
  assign new_n265_ = id2_2_ & ~id3_3_;
  assign new_n266_ = ~id2_2_ & id3_3_;
  assign new_n267_ = ~new_n265_ & ~new_n266_;
  assign new_n268_ = id0_0_ & ~id1_1_;
  assign new_n269_ = ~id0_0_ & id1_1_;
  assign new_n270_ = ~new_n268_ & ~new_n269_;
  assign new_n271_ = new_n267_ & ~new_n270_;
  assign new_n272_ = ~new_n267_ & new_n270_;
  assign new_n273_ = ~new_n271_ & ~new_n272_;
  assign new_n274_ = new_n245_ & ~new_n273_;
  assign new_n275_ = ~new_n245_ & new_n273_;
  assign new_n276_ = ~new_n274_ & ~new_n275_;
  assign new_n277_ = ic6_38_ & r_40_;
  assign new_n278_ = new_n276_ & new_n277_;
  assign new_n279_ = ~new_n276_ & ~new_n277_;
  assign new_n280_ = ~new_n278_ & ~new_n279_;
  assign new_n281_ = id26_26_ & ~id30_30_;
  assign new_n282_ = ~id26_26_ & id30_30_;
  assign new_n283_ = ~new_n281_ & ~new_n282_;
  assign new_n284_ = ~id22_22_ & id18_18_;
  assign new_n285_ = id22_22_ & ~id18_18_;
  assign new_n286_ = ~new_n284_ & ~new_n285_;
  assign new_n287_ = new_n283_ & ~new_n286_;
  assign new_n288_ = ~new_n283_ & new_n286_;
  assign new_n289_ = ~new_n287_ & ~new_n288_;
  assign new_n290_ = new_n280_ & ~new_n289_;
  assign new_n291_ = ~new_n280_ & new_n289_;
  assign new_n292_ = ~new_n290_ & ~new_n291_;
  assign new_n293_ = new_n91_ & ~new_n273_;
  assign new_n294_ = ~new_n91_ & new_n273_;
  assign new_n295_ = ~new_n293_ & ~new_n294_;
  assign new_n296_ = ic4_36_ & r_40_;
  assign new_n297_ = new_n295_ & new_n296_;
  assign new_n298_ = ~new_n295_ & ~new_n296_;
  assign new_n299_ = ~new_n297_ & ~new_n298_;
  assign new_n300_ = ~id28_28_ & id24_24_;
  assign new_n301_ = id28_28_ & ~id24_24_;
  assign new_n302_ = ~new_n300_ & ~new_n301_;
  assign new_n303_ = ~id20_20_ & id16_16_;
  assign new_n304_ = id20_20_ & ~id16_16_;
  assign new_n305_ = ~new_n303_ & ~new_n304_;
  assign new_n306_ = new_n302_ & ~new_n305_;
  assign new_n307_ = ~new_n302_ & new_n305_;
  assign new_n308_ = ~new_n306_ & ~new_n307_;
  assign new_n309_ = new_n299_ & ~new_n308_;
  assign new_n310_ = ~new_n299_ & new_n308_;
  assign new_n311_ = ~new_n309_ & ~new_n310_;
  assign new_n312_ = new_n110_ & ~new_n236_;
  assign new_n313_ = ~new_n264_ & new_n312_;
  assign new_n314_ = ~new_n292_ & new_n313_;
  assign new_n315_ = new_n311_ & new_n314_;
  assign new_n316_ = ~new_n203_ & new_n315_;
  assign new_n317_ = id10_10_ & ~new_n316_;
  assign new_n318_ = ~id10_10_ & new_n316_;
  assign od10_232_ = new_n317_ | new_n318_;
  assign new_n320_ = ~new_n147_ & new_n315_;
  assign new_n321_ = id11_11_ & ~new_n320_;
  assign new_n322_ = ~id11_11_ & new_n320_;
  assign od11_231_ = new_n321_ | new_n322_;
  assign new_n324_ = ~new_n110_ & ~new_n236_;
  assign new_n325_ = ~new_n264_ & new_n324_;
  assign new_n326_ = new_n292_ & new_n325_;
  assign new_n327_ = new_n311_ & new_n326_;
  assign new_n328_ = ~new_n222_ & new_n327_;
  assign new_n329_ = id12_12_ & ~new_n328_;
  assign new_n330_ = ~id12_12_ & new_n328_;
  assign od12_230_ = new_n329_ | new_n330_;
  assign new_n332_ = new_n264_ & new_n324_;
  assign new_n333_ = new_n292_ & new_n332_;
  assign new_n334_ = ~new_n311_ & new_n333_;
  assign new_n335_ = ~new_n222_ & new_n334_;
  assign new_n336_ = id4_4_ & ~new_n335_;
  assign new_n337_ = ~id4_4_ & new_n335_;
  assign od4_238_ = new_n336_ | new_n337_;
  assign new_n339_ = ~new_n222_ & new_n315_;
  assign new_n340_ = id8_8_ & ~new_n339_;
  assign new_n341_ = ~id8_8_ & new_n339_;
  assign od8_234_ = new_n340_ | new_n341_;
  assign new_n343_ = new_n264_ & new_n312_;
  assign new_n344_ = ~new_n292_ & new_n343_;
  assign new_n345_ = ~new_n311_ & new_n344_;
  assign new_n346_ = ~new_n175_ & new_n345_;
  assign new_n347_ = id1_1_ & ~new_n346_;
  assign new_n348_ = ~id1_1_ & new_n346_;
  assign od1_241_ = new_n347_ | new_n348_;
  assign new_n350_ = new_n110_ & new_n264_;
  assign new_n351_ = new_n292_ & new_n350_;
  assign new_n352_ = ~new_n311_ & new_n351_;
  assign new_n353_ = ~new_n292_ & new_n350_;
  assign new_n354_ = new_n311_ & new_n353_;
  assign new_n355_ = new_n110_ & ~new_n264_;
  assign new_n356_ = new_n292_ & new_n355_;
  assign new_n357_ = new_n311_ & new_n356_;
  assign new_n358_ = ~new_n110_ & new_n264_;
  assign new_n359_ = new_n292_ & new_n358_;
  assign new_n360_ = new_n311_ & new_n359_;
  assign new_n361_ = ~new_n352_ & ~new_n354_;
  assign new_n362_ = ~new_n357_ & new_n361_;
  assign new_n363_ = ~new_n360_ & new_n362_;
  assign new_n364_ = ~new_n147_ & ~new_n363_;
  assign new_n365_ = new_n175_ & new_n364_;
  assign new_n366_ = new_n203_ & new_n365_;
  assign new_n367_ = ~new_n222_ & new_n366_;
  assign new_n368_ = ~new_n311_ & new_n367_;
  assign new_n369_ = id20_20_ & ~new_n368_;
  assign new_n370_ = ~id20_20_ & new_n368_;
  assign od20_222_ = new_n369_ | new_n370_;
  assign new_n372_ = ~new_n264_ & new_n367_;
  assign new_n373_ = id21_21_ & ~new_n372_;
  assign new_n374_ = ~id21_21_ & new_n372_;
  assign od21_221_ = new_n373_ | new_n374_;
  assign new_n376_ = ~new_n292_ & new_n367_;
  assign new_n377_ = id22_22_ & ~new_n376_;
  assign new_n378_ = ~id22_22_ & new_n376_;
  assign od22_220_ = new_n377_ | new_n378_;
  assign new_n380_ = ~new_n175_ & new_n334_;
  assign new_n381_ = id5_5_ & ~new_n380_;
  assign new_n382_ = ~id5_5_ & new_n380_;
  assign od5_237_ = new_n381_ | new_n382_;
  assign new_n384_ = ~new_n175_ & new_n315_;
  assign new_n385_ = id9_9_ & ~new_n384_;
  assign new_n386_ = ~id9_9_ & new_n384_;
  assign od9_233_ = new_n385_ | new_n386_;
  assign new_n388_ = ~new_n203_ & new_n345_;
  assign new_n389_ = id2_2_ & ~new_n388_;
  assign new_n390_ = ~id2_2_ & new_n388_;
  assign od2_240_ = new_n389_ | new_n390_;
  assign new_n392_ = ~new_n110_ & new_n367_;
  assign new_n393_ = id23_23_ & ~new_n392_;
  assign new_n394_ = ~id23_23_ & new_n392_;
  assign od23_219_ = new_n393_ | new_n394_;
  assign new_n396_ = new_n147_ & ~new_n363_;
  assign new_n397_ = ~new_n175_ & new_n396_;
  assign new_n398_ = ~new_n203_ & new_n397_;
  assign new_n399_ = new_n222_ & new_n398_;
  assign new_n400_ = ~new_n311_ & new_n399_;
  assign new_n401_ = id24_24_ & ~new_n400_;
  assign new_n402_ = ~id24_24_ & new_n400_;
  assign od24_218_ = new_n401_ | new_n402_;
  assign new_n404_ = ~new_n264_ & new_n399_;
  assign new_n405_ = id25_25_ & ~new_n404_;
  assign new_n406_ = ~id25_25_ & new_n404_;
  assign od25_217_ = new_n405_ | new_n406_;
  assign new_n408_ = ~new_n292_ & new_n399_;
  assign new_n409_ = id26_26_ & ~new_n408_;
  assign new_n410_ = ~id26_26_ & new_n408_;
  assign od26_216_ = new_n409_ | new_n410_;
  assign new_n412_ = ~new_n110_ & new_n399_;
  assign new_n413_ = id27_27_ & ~new_n412_;
  assign new_n414_ = ~id27_27_ & new_n412_;
  assign od27_215_ = new_n413_ | new_n414_;
  assign new_n416_ = ~new_n175_ & new_n364_;
  assign new_n417_ = new_n203_ & new_n416_;
  assign new_n418_ = new_n222_ & new_n417_;
  assign new_n419_ = ~new_n311_ & new_n418_;
  assign new_n420_ = id28_28_ & ~new_n419_;
  assign new_n421_ = ~id28_28_ & new_n419_;
  assign od28_214_ = new_n420_ | new_n421_;
  assign new_n423_ = ~new_n264_ & new_n418_;
  assign new_n424_ = id29_29_ & ~new_n423_;
  assign new_n425_ = ~id29_29_ & new_n423_;
  assign od29_213_ = new_n424_ | new_n425_;
  assign new_n427_ = ~new_n292_ & new_n418_;
  assign new_n428_ = id30_30_ & ~new_n427_;
  assign new_n429_ = ~id30_30_ & new_n427_;
  assign od30_212_ = new_n428_ | new_n429_;
  assign new_n431_ = ~new_n110_ & new_n418_;
  assign new_n432_ = id31_31_ & ~new_n431_;
  assign new_n433_ = ~id31_31_ & new_n431_;
  assign od31_211_ = new_n432_ | new_n433_;
  assign new_n435_ = ~new_n203_ & new_n334_;
  assign new_n436_ = id6_6_ & ~new_n435_;
  assign new_n437_ = ~id6_6_ & new_n435_;
  assign od6_236_ = new_n436_ | new_n437_;
  assign new_n439_ = ~new_n175_ & new_n327_;
  assign new_n440_ = id13_13_ & ~new_n439_;
  assign new_n441_ = ~id13_13_ & new_n439_;
  assign od13_229_ = new_n440_ | new_n441_;
  assign new_n443_ = ~new_n203_ & new_n327_;
  assign new_n444_ = id14_14_ & ~new_n443_;
  assign new_n445_ = ~id14_14_ & new_n443_;
  assign od14_228_ = new_n444_ | new_n445_;
  assign new_n447_ = ~new_n147_ & new_n327_;
  assign new_n448_ = id15_15_ & ~new_n447_;
  assign new_n449_ = ~id15_15_ & new_n447_;
  assign od15_227_ = new_n448_ | new_n449_;
  assign new_n451_ = new_n175_ & new_n396_;
  assign new_n452_ = ~new_n203_ & new_n451_;
  assign new_n453_ = ~new_n222_ & new_n452_;
  assign new_n454_ = ~new_n311_ & new_n453_;
  assign new_n455_ = id16_16_ & ~new_n454_;
  assign new_n456_ = ~id16_16_ & new_n454_;
  assign od16_226_ = new_n455_ | new_n456_;
  assign new_n458_ = ~new_n264_ & new_n453_;
  assign new_n459_ = id17_17_ & ~new_n458_;
  assign new_n460_ = ~id17_17_ & new_n458_;
  assign od17_225_ = new_n459_ | new_n460_;
  assign new_n462_ = ~new_n292_ & new_n453_;
  assign new_n463_ = id18_18_ & ~new_n462_;
  assign new_n464_ = ~id18_18_ & new_n462_;
  assign od18_224_ = new_n463_ | new_n464_;
  assign new_n466_ = ~new_n110_ & new_n453_;
  assign new_n467_ = id19_19_ & ~new_n466_;
  assign new_n468_ = ~id19_19_ & new_n466_;
  assign od19_223_ = new_n467_ | new_n468_;
  assign new_n470_ = ~new_n147_ & new_n345_;
  assign new_n471_ = id3_3_ & ~new_n470_;
  assign new_n472_ = ~id3_3_ & new_n470_;
  assign od3_239_ = new_n471_ | new_n472_;
  assign new_n474_ = ~new_n147_ & new_n334_;
  assign new_n475_ = id7_7_ & ~new_n474_;
  assign new_n476_ = ~id7_7_ & new_n474_;
  assign od7_235_ = new_n475_ | new_n476_;
  assign new_n478_ = ~new_n222_ & new_n345_;
  assign new_n479_ = id0_0_ & ~new_n478_;
  assign new_n480_ = ~id0_0_ & new_n478_;
  assign od0_242_ = new_n479_ | new_n480_;
endmodule

