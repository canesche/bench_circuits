// Benchmark "testing" written by ABC on Thu Oct  8 22:16:45 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A106  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A106;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ , \new_[350]_ ,
    \new_[351]_ , \new_[352]_ , \new_[353]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[405]_ ,
    \new_[406]_ , \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ ,
    \new_[411]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[436]_ , \new_[437]_ , \new_[438]_ , \new_[439]_ , \new_[440]_ ,
    \new_[441]_ , \new_[442]_ , \new_[443]_ , \new_[444]_ , \new_[445]_ ,
    \new_[446]_ , \new_[447]_ , \new_[448]_ , \new_[449]_ , \new_[450]_ ,
    \new_[451]_ , \new_[452]_ , \new_[453]_ , \new_[454]_ , \new_[455]_ ,
    \new_[456]_ , \new_[457]_ , \new_[458]_ , \new_[459]_ , \new_[460]_ ,
    \new_[461]_ , \new_[462]_ , \new_[463]_ , \new_[464]_ , \new_[465]_ ,
    \new_[466]_ , \new_[467]_ , \new_[468]_ , \new_[469]_ , \new_[470]_ ,
    \new_[471]_ , \new_[472]_ , \new_[473]_ , \new_[474]_ , \new_[475]_ ,
    \new_[476]_ , \new_[477]_ , \new_[478]_ , \new_[479]_ , \new_[480]_ ,
    \new_[481]_ , \new_[482]_ , \new_[483]_ , \new_[484]_ , \new_[485]_ ,
    \new_[486]_ , \new_[487]_ , \new_[488]_ , \new_[489]_ , \new_[490]_ ,
    \new_[491]_ , \new_[492]_ , \new_[493]_ , \new_[494]_ , \new_[495]_ ,
    \new_[496]_ , \new_[497]_ , \new_[498]_ , \new_[499]_ , \new_[500]_ ,
    \new_[501]_ , \new_[502]_ , \new_[503]_ , \new_[504]_ , \new_[505]_ ,
    \new_[506]_ , \new_[507]_ , \new_[508]_ , \new_[509]_ , \new_[510]_ ,
    \new_[511]_ , \new_[512]_ , \new_[513]_ , \new_[514]_ , \new_[515]_ ,
    \new_[516]_ , \new_[517]_ , \new_[518]_ , \new_[519]_ , \new_[520]_ ,
    \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[525]_ ,
    \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ , \new_[530]_ ,
    \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ , \new_[535]_ ,
    \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ , \new_[540]_ ,
    \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ , \new_[545]_ ,
    \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ , \new_[550]_ ,
    \new_[551]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[566]_ , \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ ,
    \new_[571]_ , \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ ,
    \new_[576]_ , \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ ,
    \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[584]_ , \new_[585]_ ,
    \new_[586]_ , \new_[587]_ , \new_[588]_ , \new_[589]_ , \new_[590]_ ,
    \new_[591]_ , \new_[592]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[598]_ , \new_[599]_ , \new_[600]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ ,
    \new_[611]_ , \new_[612]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[616]_ , \new_[617]_ , \new_[618]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[626]_ , \new_[627]_ , \new_[628]_ , \new_[629]_ , \new_[630]_ ,
    \new_[631]_ , \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ ,
    \new_[636]_ , \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ ,
    \new_[641]_ , \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ ,
    \new_[646]_ , \new_[647]_ , \new_[648]_ , \new_[649]_ , \new_[650]_ ,
    \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[655]_ ,
    \new_[656]_ , \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ ,
    \new_[661]_ , \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ ,
    \new_[666]_ , \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ ,
    \new_[671]_ , \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ ,
    \new_[676]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ ,
    \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ ,
    \new_[686]_ , \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ ,
    \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ ,
    \new_[696]_ , \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ ,
    \new_[701]_ , \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ ,
    \new_[706]_ , \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ ,
    \new_[711]_ , \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ ,
    \new_[716]_ , \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ ,
    \new_[726]_ , \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ ,
    \new_[731]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[736]_ , \new_[737]_ , \new_[738]_ , \new_[739]_ , \new_[740]_ ,
    \new_[741]_ , \new_[742]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ ,
    \new_[746]_ , \new_[747]_ , \new_[748]_ , \new_[749]_ , \new_[750]_ ,
    \new_[751]_ , \new_[752]_ , \new_[753]_ , \new_[754]_ , \new_[755]_ ,
    \new_[756]_ , \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ ,
    \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ ,
    \new_[766]_ , \new_[767]_ , \new_[768]_ , \new_[769]_ , \new_[770]_ ,
    \new_[771]_ , \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ ,
    \new_[776]_ , \new_[777]_ , \new_[778]_ , \new_[779]_ , \new_[780]_ ,
    \new_[781]_ , \new_[782]_ , \new_[783]_ , \new_[784]_ , \new_[785]_ ,
    \new_[786]_ , \new_[787]_ , \new_[788]_ , \new_[789]_ , \new_[790]_ ,
    \new_[791]_ , \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ ,
    \new_[796]_ , \new_[797]_ , \new_[798]_ , \new_[799]_ , \new_[800]_ ,
    \new_[801]_ , \new_[802]_ , \new_[803]_ , \new_[804]_ , \new_[805]_ ,
    \new_[806]_ , \new_[807]_ , \new_[808]_ , \new_[809]_ , \new_[810]_ ,
    \new_[811]_ , \new_[812]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ ,
    \new_[816]_ , \new_[817]_ , \new_[818]_ , \new_[819]_ , \new_[820]_ ,
    \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[824]_ , \new_[825]_ ,
    \new_[826]_ , \new_[827]_ , \new_[828]_ , \new_[829]_ , \new_[830]_ ,
    \new_[831]_ , \new_[832]_ , \new_[833]_ , \new_[834]_ , \new_[835]_ ,
    \new_[836]_ , \new_[837]_ , \new_[838]_ , \new_[839]_ , \new_[840]_ ,
    \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[845]_ ,
    \new_[846]_ , \new_[847]_ , \new_[848]_ , \new_[849]_ , \new_[850]_ ,
    \new_[851]_ , \new_[852]_ , \new_[853]_ , \new_[854]_ , \new_[855]_ ,
    \new_[856]_ , \new_[857]_ , \new_[858]_ , \new_[859]_ , \new_[860]_ ,
    \new_[861]_ , \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[865]_ ,
    \new_[866]_ , \new_[867]_ , \new_[868]_ , \new_[869]_ , \new_[870]_ ,
    \new_[871]_ , \new_[872]_ , \new_[873]_ , \new_[874]_ , \new_[875]_ ,
    \new_[876]_ , \new_[877]_ , \new_[878]_ , \new_[879]_ , \new_[880]_ ,
    \new_[881]_ , \new_[882]_ , \new_[883]_ , \new_[884]_ , \new_[885]_ ,
    \new_[886]_ , \new_[887]_ , \new_[888]_ , \new_[889]_ , \new_[890]_ ,
    \new_[891]_ , \new_[892]_ , \new_[893]_ , \new_[894]_ , \new_[895]_ ,
    \new_[896]_ , \new_[897]_ , \new_[898]_ , \new_[899]_ , \new_[900]_ ,
    \new_[901]_ , \new_[902]_ , \new_[903]_ , \new_[904]_ , \new_[905]_ ,
    \new_[906]_ , \new_[907]_ , \new_[908]_ , \new_[909]_ , \new_[910]_ ,
    \new_[911]_ , \new_[912]_ , \new_[913]_ , \new_[914]_ , \new_[915]_ ,
    \new_[916]_ , \new_[917]_ , \new_[918]_ , \new_[919]_ , \new_[920]_ ,
    \new_[921]_ , \new_[922]_ , \new_[923]_ , \new_[924]_ , \new_[925]_ ,
    \new_[926]_ , \new_[927]_ , \new_[928]_ , \new_[929]_ , \new_[930]_ ,
    \new_[931]_ , \new_[932]_ , \new_[933]_ , \new_[934]_ , \new_[935]_ ,
    \new_[936]_ , \new_[937]_ , \new_[938]_ , \new_[939]_ , \new_[940]_ ,
    \new_[941]_ , \new_[942]_ , \new_[943]_ , \new_[944]_ , \new_[945]_ ,
    \new_[946]_ , \new_[947]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ ,
    \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[955]_ ,
    \new_[956]_ , \new_[957]_ , \new_[958]_ , \new_[959]_ , \new_[960]_ ,
    \new_[961]_ , \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ ,
    \new_[966]_ , \new_[967]_ , \new_[968]_ , \new_[969]_ , \new_[970]_ ,
    \new_[971]_ , \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[975]_ ,
    \new_[976]_ , \new_[977]_ , \new_[978]_ , \new_[979]_ , \new_[980]_ ,
    \new_[981]_ , \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ ,
    \new_[986]_ , \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ ,
    \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ ,
    \new_[996]_ , \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ ,
    \new_[1001]_ , \new_[1002]_ , \new_[1003]_ , \new_[1004]_ ,
    \new_[1005]_ , \new_[1006]_ , \new_[1007]_ , \new_[1008]_ ,
    \new_[1009]_ , \new_[1010]_ , \new_[1011]_ , \new_[1012]_ ,
    \new_[1013]_ , \new_[1014]_ , \new_[1015]_ , \new_[1016]_ ,
    \new_[1017]_ , \new_[1018]_ , \new_[1019]_ , \new_[1020]_ ,
    \new_[1021]_ , \new_[1022]_ , \new_[1023]_ , \new_[1024]_ ,
    \new_[1025]_ , \new_[1026]_ , \new_[1027]_ , \new_[1028]_ ,
    \new_[1029]_ , \new_[1030]_ , \new_[1031]_ , \new_[1032]_ ,
    \new_[1033]_ , \new_[1034]_ , \new_[1035]_ , \new_[1036]_ ,
    \new_[1037]_ , \new_[1038]_ , \new_[1039]_ , \new_[1040]_ ,
    \new_[1041]_ , \new_[1042]_ , \new_[1043]_ , \new_[1044]_ ,
    \new_[1045]_ , \new_[1046]_ , \new_[1047]_ , \new_[1048]_ ,
    \new_[1049]_ , \new_[1050]_ , \new_[1051]_ , \new_[1052]_ ,
    \new_[1053]_ , \new_[1054]_ , \new_[1055]_ , \new_[1056]_ ,
    \new_[1057]_ , \new_[1058]_ , \new_[1059]_ , \new_[1060]_ ,
    \new_[1061]_ , \new_[1062]_ , \new_[1063]_ , \new_[1064]_ ,
    \new_[1065]_ , \new_[1066]_ , \new_[1067]_ , \new_[1068]_ ,
    \new_[1069]_ , \new_[1070]_ , \new_[1071]_ , \new_[1072]_ ,
    \new_[1073]_ , \new_[1074]_ , \new_[1075]_ , \new_[1076]_ ,
    \new_[1077]_ , \new_[1078]_ , \new_[1079]_ , \new_[1080]_ ,
    \new_[1081]_ , \new_[1082]_ , \new_[1083]_ , \new_[1084]_ ,
    \new_[1085]_ , \new_[1086]_ , \new_[1087]_ , \new_[1088]_ ,
    \new_[1089]_ , \new_[1090]_ , \new_[1091]_ , \new_[1092]_ ,
    \new_[1093]_ , \new_[1094]_ , \new_[1095]_ , \new_[1096]_ ,
    \new_[1097]_ , \new_[1098]_ , \new_[1099]_ , \new_[1100]_ ,
    \new_[1101]_ , \new_[1102]_ , \new_[1103]_ , \new_[1104]_ ,
    \new_[1105]_ , \new_[1106]_ , \new_[1107]_ , \new_[1108]_ ,
    \new_[1109]_ , \new_[1110]_ , \new_[1111]_ , \new_[1112]_ ,
    \new_[1113]_ , \new_[1114]_ , \new_[1115]_ , \new_[1116]_ ,
    \new_[1117]_ , \new_[1118]_ , \new_[1119]_ , \new_[1122]_ ,
    \new_[1125]_ , \new_[1126]_ , \new_[1129]_ , \new_[1132]_ ,
    \new_[1133]_ , \new_[1134]_ , \new_[1137]_ , \new_[1140]_ ,
    \new_[1141]_ , \new_[1144]_ , \new_[1148]_ , \new_[1149]_ ,
    \new_[1150]_ , \new_[1151]_ , \new_[1152]_ , \new_[1155]_ ,
    \new_[1158]_ , \new_[1159]_ , \new_[1162]_ , \new_[1165]_ ,
    \new_[1166]_ , \new_[1167]_ , \new_[1170]_ , \new_[1173]_ ,
    \new_[1174]_ , \new_[1177]_ , \new_[1181]_ , \new_[1182]_ ,
    \new_[1183]_ , \new_[1184]_ , \new_[1185]_ , \new_[1186]_ ,
    \new_[1189]_ , \new_[1192]_ , \new_[1193]_ , \new_[1196]_ ,
    \new_[1199]_ , \new_[1200]_ , \new_[1201]_ , \new_[1204]_ ,
    \new_[1207]_ , \new_[1208]_ , \new_[1211]_ , \new_[1215]_ ,
    \new_[1216]_ , \new_[1217]_ , \new_[1218]_ , \new_[1219]_ ,
    \new_[1222]_ , \new_[1225]_ , \new_[1226]_ , \new_[1229]_ ,
    \new_[1233]_ , \new_[1234]_ , \new_[1235]_ , \new_[1236]_ ,
    \new_[1239]_ , \new_[1242]_ , \new_[1243]_ , \new_[1246]_ ,
    \new_[1250]_ , \new_[1251]_ , \new_[1252]_ , \new_[1253]_ ,
    \new_[1254]_ , \new_[1255]_ , \new_[1256]_ , \new_[1259]_ ,
    \new_[1262]_ , \new_[1263]_ , \new_[1266]_ , \new_[1269]_ ,
    \new_[1270]_ , \new_[1271]_ , \new_[1274]_ , \new_[1277]_ ,
    \new_[1278]_ , \new_[1281]_ , \new_[1285]_ , \new_[1286]_ ,
    \new_[1287]_ , \new_[1288]_ , \new_[1289]_ , \new_[1292]_ ,
    \new_[1295]_ , \new_[1296]_ , \new_[1299]_ , \new_[1303]_ ,
    \new_[1304]_ , \new_[1305]_ , \new_[1306]_ , \new_[1309]_ ,
    \new_[1312]_ , \new_[1313]_ , \new_[1316]_ , \new_[1320]_ ,
    \new_[1321]_ , \new_[1322]_ , \new_[1323]_ , \new_[1324]_ ,
    \new_[1325]_ , \new_[1328]_ , \new_[1331]_ , \new_[1332]_ ,
    \new_[1335]_ , \new_[1338]_ , \new_[1339]_ , \new_[1340]_ ,
    \new_[1343]_ , \new_[1346]_ , \new_[1347]_ , \new_[1350]_ ,
    \new_[1354]_ , \new_[1355]_ , \new_[1356]_ , \new_[1357]_ ,
    \new_[1358]_ , \new_[1361]_ , \new_[1364]_ , \new_[1365]_ ,
    \new_[1368]_ , \new_[1372]_ , \new_[1373]_ , \new_[1374]_ ,
    \new_[1375]_ , \new_[1378]_ , \new_[1381]_ , \new_[1382]_ ,
    \new_[1385]_ , \new_[1389]_ , \new_[1390]_ , \new_[1391]_ ,
    \new_[1392]_ , \new_[1393]_ , \new_[1394]_ , \new_[1395]_ ,
    \new_[1396]_ , \new_[1399]_ , \new_[1402]_ , \new_[1403]_ ,
    \new_[1406]_ , \new_[1409]_ , \new_[1410]_ , \new_[1411]_ ,
    \new_[1414]_ , \new_[1417]_ , \new_[1418]_ , \new_[1421]_ ,
    \new_[1425]_ , \new_[1426]_ , \new_[1427]_ , \new_[1428]_ ,
    \new_[1429]_ , \new_[1432]_ , \new_[1435]_ , \new_[1436]_ ,
    \new_[1439]_ , \new_[1443]_ , \new_[1444]_ , \new_[1445]_ ,
    \new_[1446]_ , \new_[1449]_ , \new_[1452]_ , \new_[1453]_ ,
    \new_[1456]_ , \new_[1460]_ , \new_[1461]_ , \new_[1462]_ ,
    \new_[1463]_ , \new_[1464]_ , \new_[1465]_ , \new_[1468]_ ,
    \new_[1471]_ , \new_[1472]_ , \new_[1475]_ , \new_[1478]_ ,
    \new_[1479]_ , \new_[1480]_ , \new_[1483]_ , \new_[1486]_ ,
    \new_[1487]_ , \new_[1490]_ , \new_[1494]_ , \new_[1495]_ ,
    \new_[1496]_ , \new_[1497]_ , \new_[1498]_ , \new_[1501]_ ,
    \new_[1504]_ , \new_[1505]_ , \new_[1508]_ , \new_[1512]_ ,
    \new_[1513]_ , \new_[1514]_ , \new_[1515]_ , \new_[1518]_ ,
    \new_[1521]_ , \new_[1522]_ , \new_[1525]_ , \new_[1529]_ ,
    \new_[1530]_ , \new_[1531]_ , \new_[1532]_ , \new_[1533]_ ,
    \new_[1534]_ , \new_[1535]_ , \new_[1538]_ , \new_[1541]_ ,
    \new_[1542]_ , \new_[1545]_ , \new_[1548]_ , \new_[1549]_ ,
    \new_[1550]_ , \new_[1553]_ , \new_[1556]_ , \new_[1557]_ ,
    \new_[1560]_ , \new_[1564]_ , \new_[1565]_ , \new_[1566]_ ,
    \new_[1567]_ , \new_[1568]_ , \new_[1571]_ , \new_[1574]_ ,
    \new_[1575]_ , \new_[1578]_ , \new_[1582]_ , \new_[1583]_ ,
    \new_[1584]_ , \new_[1585]_ , \new_[1588]_ , \new_[1591]_ ,
    \new_[1592]_ , \new_[1595]_ , \new_[1599]_ , \new_[1600]_ ,
    \new_[1601]_ , \new_[1602]_ , \new_[1603]_ , \new_[1604]_ ,
    \new_[1607]_ , \new_[1610]_ , \new_[1611]_ , \new_[1614]_ ,
    \new_[1617]_ , \new_[1618]_ , \new_[1619]_ , \new_[1622]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1629]_ , \new_[1633]_ ,
    \new_[1634]_ , \new_[1635]_ , \new_[1636]_ , \new_[1637]_ ,
    \new_[1640]_ , \new_[1643]_ , \new_[1644]_ , \new_[1647]_ ,
    \new_[1651]_ , \new_[1652]_ , \new_[1653]_ , \new_[1654]_ ,
    \new_[1657]_ , \new_[1660]_ , \new_[1661]_ , \new_[1664]_ ,
    \new_[1668]_ , \new_[1669]_ , \new_[1670]_ , \new_[1671]_ ,
    \new_[1672]_ , \new_[1673]_ , \new_[1674]_ , \new_[1675]_ ,
    \new_[1676]_ , \new_[1679]_ , \new_[1682]_ , \new_[1683]_ ,
    \new_[1686]_ , \new_[1689]_ , \new_[1690]_ , \new_[1691]_ ,
    \new_[1694]_ , \new_[1697]_ , \new_[1698]_ , \new_[1701]_ ,
    \new_[1705]_ , \new_[1706]_ , \new_[1707]_ , \new_[1708]_ ,
    \new_[1709]_ , \new_[1712]_ , \new_[1715]_ , \new_[1716]_ ,
    \new_[1719]_ , \new_[1723]_ , \new_[1724]_ , \new_[1725]_ ,
    \new_[1726]_ , \new_[1729]_ , \new_[1732]_ , \new_[1733]_ ,
    \new_[1736]_ , \new_[1740]_ , \new_[1741]_ , \new_[1742]_ ,
    \new_[1743]_ , \new_[1744]_ , \new_[1745]_ , \new_[1748]_ ,
    \new_[1751]_ , \new_[1752]_ , \new_[1755]_ , \new_[1758]_ ,
    \new_[1759]_ , \new_[1760]_ , \new_[1763]_ , \new_[1766]_ ,
    \new_[1767]_ , \new_[1770]_ , \new_[1774]_ , \new_[1775]_ ,
    \new_[1776]_ , \new_[1777]_ , \new_[1778]_ , \new_[1781]_ ,
    \new_[1784]_ , \new_[1785]_ , \new_[1788]_ , \new_[1792]_ ,
    \new_[1793]_ , \new_[1794]_ , \new_[1795]_ , \new_[1798]_ ,
    \new_[1801]_ , \new_[1802]_ , \new_[1805]_ , \new_[1809]_ ,
    \new_[1810]_ , \new_[1811]_ , \new_[1812]_ , \new_[1813]_ ,
    \new_[1814]_ , \new_[1815]_ , \new_[1818]_ , \new_[1821]_ ,
    \new_[1822]_ , \new_[1825]_ , \new_[1828]_ , \new_[1829]_ ,
    \new_[1830]_ , \new_[1833]_ , \new_[1836]_ , \new_[1837]_ ,
    \new_[1840]_ , \new_[1844]_ , \new_[1845]_ , \new_[1846]_ ,
    \new_[1847]_ , \new_[1848]_ , \new_[1851]_ , \new_[1854]_ ,
    \new_[1855]_ , \new_[1858]_ , \new_[1862]_ , \new_[1863]_ ,
    \new_[1864]_ , \new_[1865]_ , \new_[1868]_ , \new_[1871]_ ,
    \new_[1872]_ , \new_[1875]_ , \new_[1879]_ , \new_[1880]_ ,
    \new_[1881]_ , \new_[1882]_ , \new_[1883]_ , \new_[1884]_ ,
    \new_[1887]_ , \new_[1890]_ , \new_[1891]_ , \new_[1894]_ ,
    \new_[1897]_ , \new_[1898]_ , \new_[1899]_ , \new_[1902]_ ,
    \new_[1905]_ , \new_[1906]_ , \new_[1909]_ , \new_[1913]_ ,
    \new_[1914]_ , \new_[1915]_ , \new_[1916]_ , \new_[1917]_ ,
    \new_[1920]_ , \new_[1923]_ , \new_[1924]_ , \new_[1927]_ ,
    \new_[1931]_ , \new_[1932]_ , \new_[1933]_ , \new_[1934]_ ,
    \new_[1937]_ , \new_[1940]_ , \new_[1941]_ , \new_[1944]_ ,
    \new_[1948]_ , \new_[1949]_ , \new_[1950]_ , \new_[1951]_ ,
    \new_[1952]_ , \new_[1953]_ , \new_[1954]_ , \new_[1955]_ ,
    \new_[1958]_ , \new_[1961]_ , \new_[1962]_ , \new_[1965]_ ,
    \new_[1968]_ , \new_[1969]_ , \new_[1970]_ , \new_[1973]_ ,
    \new_[1976]_ , \new_[1977]_ , \new_[1980]_ , \new_[1984]_ ,
    \new_[1985]_ , \new_[1986]_ , \new_[1987]_ , \new_[1988]_ ,
    \new_[1991]_ , \new_[1994]_ , \new_[1995]_ , \new_[1998]_ ,
    \new_[2002]_ , \new_[2003]_ , \new_[2004]_ , \new_[2005]_ ,
    \new_[2008]_ , \new_[2011]_ , \new_[2012]_ , \new_[2015]_ ,
    \new_[2019]_ , \new_[2020]_ , \new_[2021]_ , \new_[2022]_ ,
    \new_[2023]_ , \new_[2024]_ , \new_[2027]_ , \new_[2030]_ ,
    \new_[2031]_ , \new_[2034]_ , \new_[2037]_ , \new_[2038]_ ,
    \new_[2039]_ , \new_[2042]_ , \new_[2045]_ , \new_[2046]_ ,
    \new_[2049]_ , \new_[2053]_ , \new_[2054]_ , \new_[2055]_ ,
    \new_[2056]_ , \new_[2057]_ , \new_[2060]_ , \new_[2063]_ ,
    \new_[2064]_ , \new_[2067]_ , \new_[2071]_ , \new_[2072]_ ,
    \new_[2073]_ , \new_[2074]_ , \new_[2077]_ , \new_[2080]_ ,
    \new_[2081]_ , \new_[2084]_ , \new_[2088]_ , \new_[2089]_ ,
    \new_[2090]_ , \new_[2091]_ , \new_[2092]_ , \new_[2093]_ ,
    \new_[2094]_ , \new_[2097]_ , \new_[2100]_ , \new_[2101]_ ,
    \new_[2104]_ , \new_[2107]_ , \new_[2108]_ , \new_[2109]_ ,
    \new_[2112]_ , \new_[2115]_ , \new_[2116]_ , \new_[2119]_ ,
    \new_[2123]_ , \new_[2124]_ , \new_[2125]_ , \new_[2126]_ ,
    \new_[2127]_ , \new_[2130]_ , \new_[2133]_ , \new_[2134]_ ,
    \new_[2137]_ , \new_[2141]_ , \new_[2142]_ , \new_[2143]_ ,
    \new_[2144]_ , \new_[2147]_ , \new_[2150]_ , \new_[2151]_ ,
    \new_[2154]_ , \new_[2158]_ , \new_[2159]_ , \new_[2160]_ ,
    \new_[2161]_ , \new_[2162]_ , \new_[2163]_ , \new_[2166]_ ,
    \new_[2169]_ , \new_[2170]_ , \new_[2173]_ , \new_[2176]_ ,
    \new_[2177]_ , \new_[2178]_ , \new_[2181]_ , \new_[2184]_ ,
    \new_[2185]_ , \new_[2188]_ , \new_[2192]_ , \new_[2193]_ ,
    \new_[2194]_ , \new_[2195]_ , \new_[2196]_ , \new_[2199]_ ,
    \new_[2202]_ , \new_[2203]_ , \new_[2206]_ , \new_[2210]_ ,
    \new_[2211]_ , \new_[2212]_ , \new_[2213]_ , \new_[2216]_ ,
    \new_[2219]_ , \new_[2220]_ , \new_[2223]_ , \new_[2227]_ ,
    \new_[2228]_ , \new_[2229]_ , \new_[2230]_ , \new_[2231]_ ,
    \new_[2232]_ , \new_[2233]_ , \new_[2234]_ , \new_[2235]_ ,
    \new_[2236]_ , \new_[2239]_ , \new_[2242]_ , \new_[2243]_ ,
    \new_[2246]_ , \new_[2249]_ , \new_[2250]_ , \new_[2251]_ ,
    \new_[2254]_ , \new_[2257]_ , \new_[2258]_ , \new_[2261]_ ,
    \new_[2265]_ , \new_[2266]_ , \new_[2267]_ , \new_[2268]_ ,
    \new_[2269]_ , \new_[2272]_ , \new_[2275]_ , \new_[2276]_ ,
    \new_[2279]_ , \new_[2283]_ , \new_[2284]_ , \new_[2285]_ ,
    \new_[2286]_ , \new_[2289]_ , \new_[2292]_ , \new_[2293]_ ,
    \new_[2296]_ , \new_[2300]_ , \new_[2301]_ , \new_[2302]_ ,
    \new_[2303]_ , \new_[2304]_ , \new_[2305]_ , \new_[2308]_ ,
    \new_[2311]_ , \new_[2312]_ , \new_[2315]_ , \new_[2318]_ ,
    \new_[2319]_ , \new_[2320]_ , \new_[2323]_ , \new_[2326]_ ,
    \new_[2327]_ , \new_[2330]_ , \new_[2334]_ , \new_[2335]_ ,
    \new_[2336]_ , \new_[2337]_ , \new_[2338]_ , \new_[2341]_ ,
    \new_[2344]_ , \new_[2345]_ , \new_[2348]_ , \new_[2352]_ ,
    \new_[2353]_ , \new_[2354]_ , \new_[2355]_ , \new_[2358]_ ,
    \new_[2361]_ , \new_[2362]_ , \new_[2365]_ , \new_[2369]_ ,
    \new_[2370]_ , \new_[2371]_ , \new_[2372]_ , \new_[2373]_ ,
    \new_[2374]_ , \new_[2375]_ , \new_[2378]_ , \new_[2381]_ ,
    \new_[2382]_ , \new_[2385]_ , \new_[2388]_ , \new_[2389]_ ,
    \new_[2390]_ , \new_[2393]_ , \new_[2396]_ , \new_[2397]_ ,
    \new_[2400]_ , \new_[2404]_ , \new_[2405]_ , \new_[2406]_ ,
    \new_[2407]_ , \new_[2408]_ , \new_[2411]_ , \new_[2414]_ ,
    \new_[2415]_ , \new_[2418]_ , \new_[2422]_ , \new_[2423]_ ,
    \new_[2424]_ , \new_[2425]_ , \new_[2428]_ , \new_[2431]_ ,
    \new_[2432]_ , \new_[2435]_ , \new_[2439]_ , \new_[2440]_ ,
    \new_[2441]_ , \new_[2442]_ , \new_[2443]_ , \new_[2444]_ ,
    \new_[2447]_ , \new_[2450]_ , \new_[2451]_ , \new_[2454]_ ,
    \new_[2457]_ , \new_[2458]_ , \new_[2459]_ , \new_[2462]_ ,
    \new_[2465]_ , \new_[2466]_ , \new_[2469]_ , \new_[2473]_ ,
    \new_[2474]_ , \new_[2475]_ , \new_[2476]_ , \new_[2477]_ ,
    \new_[2480]_ , \new_[2483]_ , \new_[2484]_ , \new_[2487]_ ,
    \new_[2491]_ , \new_[2492]_ , \new_[2493]_ , \new_[2494]_ ,
    \new_[2497]_ , \new_[2500]_ , \new_[2501]_ , \new_[2504]_ ,
    \new_[2508]_ , \new_[2509]_ , \new_[2510]_ , \new_[2511]_ ,
    \new_[2512]_ , \new_[2513]_ , \new_[2514]_ , \new_[2515]_ ,
    \new_[2518]_ , \new_[2521]_ , \new_[2522]_ , \new_[2525]_ ,
    \new_[2528]_ , \new_[2529]_ , \new_[2530]_ , \new_[2533]_ ,
    \new_[2536]_ , \new_[2537]_ , \new_[2540]_ , \new_[2544]_ ,
    \new_[2545]_ , \new_[2546]_ , \new_[2547]_ , \new_[2548]_ ,
    \new_[2551]_ , \new_[2554]_ , \new_[2555]_ , \new_[2558]_ ,
    \new_[2562]_ , \new_[2563]_ , \new_[2564]_ , \new_[2565]_ ,
    \new_[2568]_ , \new_[2571]_ , \new_[2572]_ , \new_[2575]_ ,
    \new_[2579]_ , \new_[2580]_ , \new_[2581]_ , \new_[2582]_ ,
    \new_[2583]_ , \new_[2584]_ , \new_[2587]_ , \new_[2590]_ ,
    \new_[2591]_ , \new_[2594]_ , \new_[2597]_ , \new_[2598]_ ,
    \new_[2599]_ , \new_[2602]_ , \new_[2605]_ , \new_[2606]_ ,
    \new_[2609]_ , \new_[2613]_ , \new_[2614]_ , \new_[2615]_ ,
    \new_[2616]_ , \new_[2617]_ , \new_[2620]_ , \new_[2623]_ ,
    \new_[2624]_ , \new_[2627]_ , \new_[2631]_ , \new_[2632]_ ,
    \new_[2633]_ , \new_[2634]_ , \new_[2637]_ , \new_[2640]_ ,
    \new_[2641]_ , \new_[2644]_ , \new_[2648]_ , \new_[2649]_ ,
    \new_[2650]_ , \new_[2651]_ , \new_[2652]_ , \new_[2653]_ ,
    \new_[2654]_ , \new_[2657]_ , \new_[2660]_ , \new_[2661]_ ,
    \new_[2664]_ , \new_[2667]_ , \new_[2668]_ , \new_[2669]_ ,
    \new_[2672]_ , \new_[2675]_ , \new_[2676]_ , \new_[2679]_ ,
    \new_[2683]_ , \new_[2684]_ , \new_[2685]_ , \new_[2686]_ ,
    \new_[2687]_ , \new_[2690]_ , \new_[2693]_ , \new_[2694]_ ,
    \new_[2697]_ , \new_[2701]_ , \new_[2702]_ , \new_[2703]_ ,
    \new_[2704]_ , \new_[2707]_ , \new_[2710]_ , \new_[2711]_ ,
    \new_[2714]_ , \new_[2718]_ , \new_[2719]_ , \new_[2720]_ ,
    \new_[2721]_ , \new_[2722]_ , \new_[2723]_ , \new_[2726]_ ,
    \new_[2729]_ , \new_[2730]_ , \new_[2733]_ , \new_[2736]_ ,
    \new_[2737]_ , \new_[2738]_ , \new_[2741]_ , \new_[2744]_ ,
    \new_[2745]_ , \new_[2748]_ , \new_[2752]_ , \new_[2753]_ ,
    \new_[2754]_ , \new_[2755]_ , \new_[2756]_ , \new_[2759]_ ,
    \new_[2762]_ , \new_[2763]_ , \new_[2766]_ , \new_[2770]_ ,
    \new_[2771]_ , \new_[2772]_ , \new_[2773]_ , \new_[2776]_ ,
    \new_[2779]_ , \new_[2780]_ , \new_[2783]_ , \new_[2787]_ ,
    \new_[2788]_ , \new_[2789]_ , \new_[2790]_ , \new_[2791]_ ,
    \new_[2792]_ , \new_[2793]_ , \new_[2794]_ , \new_[2795]_ ,
    \new_[2798]_ , \new_[2801]_ , \new_[2802]_ , \new_[2805]_ ,
    \new_[2808]_ , \new_[2809]_ , \new_[2810]_ , \new_[2813]_ ,
    \new_[2816]_ , \new_[2817]_ , \new_[2820]_ , \new_[2824]_ ,
    \new_[2825]_ , \new_[2826]_ , \new_[2827]_ , \new_[2828]_ ,
    \new_[2831]_ , \new_[2834]_ , \new_[2835]_ , \new_[2838]_ ,
    \new_[2842]_ , \new_[2843]_ , \new_[2844]_ , \new_[2845]_ ,
    \new_[2848]_ , \new_[2851]_ , \new_[2852]_ , \new_[2855]_ ,
    \new_[2859]_ , \new_[2860]_ , \new_[2861]_ , \new_[2862]_ ,
    \new_[2863]_ , \new_[2864]_ , \new_[2867]_ , \new_[2870]_ ,
    \new_[2871]_ , \new_[2874]_ , \new_[2877]_ , \new_[2878]_ ,
    \new_[2879]_ , \new_[2882]_ , \new_[2885]_ , \new_[2886]_ ,
    \new_[2889]_ , \new_[2893]_ , \new_[2894]_ , \new_[2895]_ ,
    \new_[2896]_ , \new_[2897]_ , \new_[2900]_ , \new_[2903]_ ,
    \new_[2904]_ , \new_[2907]_ , \new_[2911]_ , \new_[2912]_ ,
    \new_[2913]_ , \new_[2914]_ , \new_[2917]_ , \new_[2920]_ ,
    \new_[2921]_ , \new_[2924]_ , \new_[2928]_ , \new_[2929]_ ,
    \new_[2930]_ , \new_[2931]_ , \new_[2932]_ , \new_[2933]_ ,
    \new_[2934]_ , \new_[2937]_ , \new_[2940]_ , \new_[2941]_ ,
    \new_[2944]_ , \new_[2947]_ , \new_[2948]_ , \new_[2949]_ ,
    \new_[2952]_ , \new_[2955]_ , \new_[2956]_ , \new_[2959]_ ,
    \new_[2963]_ , \new_[2964]_ , \new_[2965]_ , \new_[2966]_ ,
    \new_[2967]_ , \new_[2970]_ , \new_[2973]_ , \new_[2974]_ ,
    \new_[2977]_ , \new_[2981]_ , \new_[2982]_ , \new_[2983]_ ,
    \new_[2984]_ , \new_[2987]_ , \new_[2990]_ , \new_[2991]_ ,
    \new_[2994]_ , \new_[2998]_ , \new_[2999]_ , \new_[3000]_ ,
    \new_[3001]_ , \new_[3002]_ , \new_[3003]_ , \new_[3006]_ ,
    \new_[3009]_ , \new_[3010]_ , \new_[3013]_ , \new_[3016]_ ,
    \new_[3017]_ , \new_[3018]_ , \new_[3021]_ , \new_[3024]_ ,
    \new_[3025]_ , \new_[3028]_ , \new_[3032]_ , \new_[3033]_ ,
    \new_[3034]_ , \new_[3035]_ , \new_[3036]_ , \new_[3039]_ ,
    \new_[3042]_ , \new_[3043]_ , \new_[3046]_ , \new_[3050]_ ,
    \new_[3051]_ , \new_[3052]_ , \new_[3053]_ , \new_[3056]_ ,
    \new_[3059]_ , \new_[3060]_ , \new_[3063]_ , \new_[3067]_ ,
    \new_[3068]_ , \new_[3069]_ , \new_[3070]_ , \new_[3071]_ ,
    \new_[3072]_ , \new_[3073]_ , \new_[3074]_ , \new_[3077]_ ,
    \new_[3080]_ , \new_[3081]_ , \new_[3084]_ , \new_[3087]_ ,
    \new_[3088]_ , \new_[3089]_ , \new_[3092]_ , \new_[3095]_ ,
    \new_[3096]_ , \new_[3099]_ , \new_[3103]_ , \new_[3104]_ ,
    \new_[3105]_ , \new_[3106]_ , \new_[3107]_ , \new_[3110]_ ,
    \new_[3113]_ , \new_[3114]_ , \new_[3117]_ , \new_[3121]_ ,
    \new_[3122]_ , \new_[3123]_ , \new_[3124]_ , \new_[3127]_ ,
    \new_[3130]_ , \new_[3131]_ , \new_[3134]_ , \new_[3138]_ ,
    \new_[3139]_ , \new_[3140]_ , \new_[3141]_ , \new_[3142]_ ,
    \new_[3143]_ , \new_[3146]_ , \new_[3149]_ , \new_[3150]_ ,
    \new_[3153]_ , \new_[3156]_ , \new_[3157]_ , \new_[3158]_ ,
    \new_[3161]_ , \new_[3164]_ , \new_[3165]_ , \new_[3168]_ ,
    \new_[3172]_ , \new_[3173]_ , \new_[3174]_ , \new_[3175]_ ,
    \new_[3176]_ , \new_[3179]_ , \new_[3182]_ , \new_[3183]_ ,
    \new_[3186]_ , \new_[3190]_ , \new_[3191]_ , \new_[3192]_ ,
    \new_[3193]_ , \new_[3196]_ , \new_[3199]_ , \new_[3200]_ ,
    \new_[3203]_ , \new_[3207]_ , \new_[3208]_ , \new_[3209]_ ,
    \new_[3210]_ , \new_[3211]_ , \new_[3212]_ , \new_[3213]_ ,
    \new_[3216]_ , \new_[3219]_ , \new_[3220]_ , \new_[3223]_ ,
    \new_[3226]_ , \new_[3227]_ , \new_[3228]_ , \new_[3231]_ ,
    \new_[3234]_ , \new_[3235]_ , \new_[3238]_ , \new_[3242]_ ,
    \new_[3243]_ , \new_[3244]_ , \new_[3245]_ , \new_[3246]_ ,
    \new_[3249]_ , \new_[3252]_ , \new_[3253]_ , \new_[3256]_ ,
    \new_[3260]_ , \new_[3261]_ , \new_[3262]_ , \new_[3263]_ ,
    \new_[3266]_ , \new_[3269]_ , \new_[3270]_ , \new_[3273]_ ,
    \new_[3277]_ , \new_[3278]_ , \new_[3279]_ , \new_[3280]_ ,
    \new_[3281]_ , \new_[3282]_ , \new_[3285]_ , \new_[3288]_ ,
    \new_[3289]_ , \new_[3292]_ , \new_[3295]_ , \new_[3296]_ ,
    \new_[3297]_ , \new_[3300]_ , \new_[3303]_ , \new_[3304]_ ,
    \new_[3307]_ , \new_[3311]_ , \new_[3312]_ , \new_[3313]_ ,
    \new_[3314]_ , \new_[3315]_ , \new_[3318]_ , \new_[3321]_ ,
    \new_[3322]_ , \new_[3325]_ , \new_[3329]_ , \new_[3330]_ ,
    \new_[3331]_ , \new_[3332]_ , \new_[3335]_ , \new_[3338]_ ,
    \new_[3339]_ , \new_[3342]_ , \new_[3346]_ , \new_[3347]_ ,
    \new_[3348]_ , \new_[3349]_ , \new_[3350]_ , \new_[3351]_ ,
    \new_[3352]_ , \new_[3353]_ , \new_[3354]_ , \new_[3355]_ ,
    \new_[3358]_ , \new_[3361]_ , \new_[3364]_ , \new_[3367]_ ,
    \new_[3370]_ , \new_[3373]_ , \new_[3377]_ , \new_[3378]_ ,
    \new_[3382]_ , \new_[3383]_ , \new_[3387]_ , \new_[3388]_ ,
    \new_[3392]_ , \new_[3393]_ , \new_[3397]_ , \new_[3398]_ ,
    \new_[3402]_ , \new_[3403]_ , \new_[3407]_ , \new_[3408]_ ,
    \new_[3412]_ , \new_[3413]_ , \new_[3417]_ , \new_[3418]_ ,
    \new_[3422]_ , \new_[3423]_ , \new_[3427]_ , \new_[3428]_ ,
    \new_[3432]_ , \new_[3433]_ , \new_[3437]_ , \new_[3438]_ ,
    \new_[3442]_ , \new_[3443]_ , \new_[3447]_ , \new_[3448]_ ,
    \new_[3452]_ , \new_[3453]_ , \new_[3457]_ , \new_[3458]_ ,
    \new_[3462]_ , \new_[3463]_ , \new_[3467]_ , \new_[3468]_ ,
    \new_[3472]_ , \new_[3473]_ , \new_[3477]_ , \new_[3478]_ ,
    \new_[3482]_ , \new_[3483]_ , \new_[3487]_ , \new_[3488]_ ,
    \new_[3492]_ , \new_[3493]_ , \new_[3496]_ , \new_[3499]_ ,
    \new_[3500]_ , \new_[3503]_ , \new_[3506]_ , \new_[3507]_ ,
    \new_[3510]_ , \new_[3513]_ , \new_[3514]_ , \new_[3517]_ ,
    \new_[3520]_ , \new_[3521]_ , \new_[3524]_ , \new_[3527]_ ,
    \new_[3528]_ , \new_[3531]_ , \new_[3534]_ , \new_[3535]_ ,
    \new_[3538]_ , \new_[3541]_ , \new_[3542]_ , \new_[3545]_ ,
    \new_[3548]_ , \new_[3549]_ , \new_[3552]_ , \new_[3555]_ ,
    \new_[3556]_ , \new_[3559]_ , \new_[3562]_ , \new_[3563]_ ,
    \new_[3566]_ , \new_[3569]_ , \new_[3570]_ , \new_[3573]_ ,
    \new_[3576]_ , \new_[3577]_ , \new_[3580]_ , \new_[3583]_ ,
    \new_[3584]_ , \new_[3587]_ , \new_[3590]_ , \new_[3591]_ ,
    \new_[3594]_ , \new_[3597]_ , \new_[3598]_ , \new_[3601]_ ,
    \new_[3604]_ , \new_[3605]_ , \new_[3608]_ , \new_[3611]_ ,
    \new_[3612]_ , \new_[3615]_ , \new_[3618]_ , \new_[3619]_ ,
    \new_[3622]_ , \new_[3625]_ , \new_[3626]_ , \new_[3629]_ ,
    \new_[3632]_ , \new_[3633]_ , \new_[3636]_ , \new_[3639]_ ,
    \new_[3640]_ , \new_[3643]_ , \new_[3646]_ , \new_[3647]_ ,
    \new_[3650]_ , \new_[3653]_ , \new_[3654]_ , \new_[3657]_ ,
    \new_[3660]_ , \new_[3661]_ , \new_[3664]_ , \new_[3667]_ ,
    \new_[3668]_ , \new_[3671]_ , \new_[3674]_ , \new_[3675]_ ,
    \new_[3678]_ , \new_[3681]_ , \new_[3682]_ , \new_[3685]_ ,
    \new_[3688]_ , \new_[3689]_ , \new_[3692]_ , \new_[3695]_ ,
    \new_[3696]_ , \new_[3699]_ , \new_[3702]_ , \new_[3703]_ ,
    \new_[3706]_ , \new_[3709]_ , \new_[3710]_ , \new_[3713]_ ,
    \new_[3716]_ , \new_[3717]_ , \new_[3720]_ , \new_[3723]_ ,
    \new_[3724]_ , \new_[3727]_ , \new_[3730]_ , \new_[3731]_ ,
    \new_[3734]_ , \new_[3737]_ , \new_[3738]_ , \new_[3741]_ ,
    \new_[3744]_ , \new_[3745]_ , \new_[3748]_ , \new_[3751]_ ,
    \new_[3752]_ , \new_[3755]_ , \new_[3758]_ , \new_[3759]_ ,
    \new_[3762]_ , \new_[3765]_ , \new_[3766]_ , \new_[3769]_ ,
    \new_[3772]_ , \new_[3773]_ , \new_[3776]_ , \new_[3779]_ ,
    \new_[3780]_ , \new_[3783]_ , \new_[3786]_ , \new_[3787]_ ,
    \new_[3790]_ , \new_[3793]_ , \new_[3794]_ , \new_[3797]_ ,
    \new_[3800]_ , \new_[3801]_ , \new_[3804]_ , \new_[3807]_ ,
    \new_[3808]_ , \new_[3811]_ , \new_[3814]_ , \new_[3815]_ ,
    \new_[3818]_ , \new_[3821]_ , \new_[3822]_ , \new_[3825]_ ,
    \new_[3828]_ , \new_[3829]_ , \new_[3832]_ , \new_[3835]_ ,
    \new_[3836]_ , \new_[3839]_ , \new_[3842]_ , \new_[3843]_ ,
    \new_[3846]_ , \new_[3849]_ , \new_[3850]_ , \new_[3853]_ ,
    \new_[3856]_ , \new_[3857]_ , \new_[3860]_ , \new_[3863]_ ,
    \new_[3864]_ , \new_[3867]_ , \new_[3870]_ , \new_[3871]_ ,
    \new_[3874]_ , \new_[3877]_ , \new_[3878]_ , \new_[3881]_ ,
    \new_[3884]_ , \new_[3885]_ , \new_[3888]_ , \new_[3891]_ ,
    \new_[3892]_ , \new_[3895]_ , \new_[3898]_ , \new_[3899]_ ,
    \new_[3902]_ , \new_[3905]_ , \new_[3906]_ , \new_[3909]_ ,
    \new_[3912]_ , \new_[3913]_ , \new_[3916]_ , \new_[3919]_ ,
    \new_[3920]_ , \new_[3923]_ , \new_[3926]_ , \new_[3927]_ ,
    \new_[3930]_ , \new_[3933]_ , \new_[3934]_ , \new_[3937]_ ,
    \new_[3940]_ , \new_[3941]_ , \new_[3944]_ , \new_[3947]_ ,
    \new_[3948]_ , \new_[3951]_ , \new_[3954]_ , \new_[3955]_ ,
    \new_[3958]_ , \new_[3961]_ , \new_[3962]_ , \new_[3965]_ ,
    \new_[3968]_ , \new_[3969]_ , \new_[3972]_ , \new_[3975]_ ,
    \new_[3976]_ , \new_[3979]_ , \new_[3982]_ , \new_[3983]_ ,
    \new_[3986]_ , \new_[3989]_ , \new_[3990]_ , \new_[3993]_ ,
    \new_[3996]_ , \new_[3997]_ , \new_[4000]_ , \new_[4003]_ ,
    \new_[4004]_ , \new_[4007]_ , \new_[4011]_ , \new_[4012]_ ,
    \new_[4013]_ , \new_[4016]_ , \new_[4019]_ , \new_[4020]_ ,
    \new_[4023]_ , \new_[4027]_ , \new_[4028]_ , \new_[4029]_ ,
    \new_[4032]_ , \new_[4035]_ , \new_[4036]_ , \new_[4039]_ ,
    \new_[4043]_ , \new_[4044]_ , \new_[4045]_ , \new_[4048]_ ,
    \new_[4051]_ , \new_[4052]_ , \new_[4055]_ , \new_[4059]_ ,
    \new_[4060]_ , \new_[4061]_ , \new_[4064]_ , \new_[4067]_ ,
    \new_[4068]_ , \new_[4071]_ , \new_[4075]_ , \new_[4076]_ ,
    \new_[4077]_ , \new_[4080]_ , \new_[4083]_ , \new_[4084]_ ,
    \new_[4087]_ , \new_[4091]_ , \new_[4092]_ , \new_[4093]_ ,
    \new_[4096]_ , \new_[4099]_ , \new_[4100]_ , \new_[4103]_ ,
    \new_[4107]_ , \new_[4108]_ , \new_[4109]_ , \new_[4112]_ ,
    \new_[4115]_ , \new_[4116]_ , \new_[4119]_ , \new_[4123]_ ,
    \new_[4124]_ , \new_[4125]_ , \new_[4128]_ , \new_[4131]_ ,
    \new_[4132]_ , \new_[4135]_ , \new_[4139]_ , \new_[4140]_ ,
    \new_[4141]_ , \new_[4144]_ , \new_[4147]_ , \new_[4148]_ ,
    \new_[4151]_ , \new_[4155]_ , \new_[4156]_ , \new_[4157]_ ,
    \new_[4160]_ , \new_[4163]_ , \new_[4164]_ , \new_[4167]_ ,
    \new_[4171]_ , \new_[4172]_ , \new_[4173]_ , \new_[4176]_ ,
    \new_[4179]_ , \new_[4180]_ , \new_[4183]_ , \new_[4187]_ ,
    \new_[4188]_ , \new_[4189]_ , \new_[4192]_ , \new_[4195]_ ,
    \new_[4196]_ , \new_[4199]_ , \new_[4203]_ , \new_[4204]_ ,
    \new_[4205]_ , \new_[4208]_ , \new_[4211]_ , \new_[4212]_ ,
    \new_[4215]_ , \new_[4219]_ , \new_[4220]_ , \new_[4221]_ ,
    \new_[4224]_ , \new_[4227]_ , \new_[4228]_ , \new_[4231]_ ,
    \new_[4235]_ , \new_[4236]_ , \new_[4237]_ , \new_[4240]_ ,
    \new_[4243]_ , \new_[4244]_ , \new_[4247]_ , \new_[4251]_ ,
    \new_[4252]_ , \new_[4253]_ , \new_[4256]_ , \new_[4259]_ ,
    \new_[4260]_ , \new_[4263]_ , \new_[4267]_ , \new_[4268]_ ,
    \new_[4269]_ , \new_[4272]_ , \new_[4275]_ , \new_[4276]_ ,
    \new_[4279]_ , \new_[4283]_ , \new_[4284]_ , \new_[4285]_ ,
    \new_[4288]_ , \new_[4291]_ , \new_[4292]_ , \new_[4295]_ ,
    \new_[4299]_ , \new_[4300]_ , \new_[4301]_ , \new_[4304]_ ,
    \new_[4307]_ , \new_[4308]_ , \new_[4311]_ , \new_[4315]_ ,
    \new_[4316]_ , \new_[4317]_ , \new_[4320]_ , \new_[4323]_ ,
    \new_[4324]_ , \new_[4327]_ , \new_[4331]_ , \new_[4332]_ ,
    \new_[4333]_ , \new_[4336]_ , \new_[4339]_ , \new_[4340]_ ,
    \new_[4343]_ , \new_[4347]_ , \new_[4348]_ , \new_[4349]_ ,
    \new_[4352]_ , \new_[4355]_ , \new_[4356]_ , \new_[4359]_ ,
    \new_[4363]_ , \new_[4364]_ , \new_[4365]_ , \new_[4368]_ ,
    \new_[4371]_ , \new_[4372]_ , \new_[4375]_ , \new_[4379]_ ,
    \new_[4380]_ , \new_[4381]_ , \new_[4384]_ , \new_[4387]_ ,
    \new_[4388]_ , \new_[4391]_ , \new_[4395]_ , \new_[4396]_ ,
    \new_[4397]_ , \new_[4400]_ , \new_[4403]_ , \new_[4404]_ ,
    \new_[4407]_ , \new_[4411]_ , \new_[4412]_ , \new_[4413]_ ,
    \new_[4416]_ , \new_[4419]_ , \new_[4420]_ , \new_[4423]_ ,
    \new_[4427]_ , \new_[4428]_ , \new_[4429]_ , \new_[4432]_ ,
    \new_[4435]_ , \new_[4436]_ , \new_[4439]_ , \new_[4443]_ ,
    \new_[4444]_ , \new_[4445]_ , \new_[4448]_ , \new_[4451]_ ,
    \new_[4452]_ , \new_[4455]_ , \new_[4459]_ , \new_[4460]_ ,
    \new_[4461]_ , \new_[4464]_ , \new_[4467]_ , \new_[4468]_ ,
    \new_[4471]_ , \new_[4475]_ , \new_[4476]_ , \new_[4477]_ ,
    \new_[4480]_ , \new_[4483]_ , \new_[4484]_ , \new_[4487]_ ,
    \new_[4491]_ , \new_[4492]_ , \new_[4493]_ , \new_[4496]_ ,
    \new_[4499]_ , \new_[4500]_ , \new_[4503]_ , \new_[4507]_ ,
    \new_[4508]_ , \new_[4509]_ , \new_[4512]_ , \new_[4515]_ ,
    \new_[4516]_ , \new_[4519]_ , \new_[4523]_ , \new_[4524]_ ,
    \new_[4525]_ , \new_[4528]_ , \new_[4531]_ , \new_[4532]_ ,
    \new_[4535]_ , \new_[4539]_ , \new_[4540]_ , \new_[4541]_ ,
    \new_[4544]_ , \new_[4547]_ , \new_[4548]_ , \new_[4551]_ ,
    \new_[4555]_ , \new_[4556]_ , \new_[4557]_ , \new_[4560]_ ,
    \new_[4563]_ , \new_[4564]_ , \new_[4567]_ , \new_[4571]_ ,
    \new_[4572]_ , \new_[4573]_ , \new_[4576]_ , \new_[4579]_ ,
    \new_[4580]_ , \new_[4583]_ , \new_[4587]_ , \new_[4588]_ ,
    \new_[4589]_ , \new_[4592]_ , \new_[4595]_ , \new_[4596]_ ,
    \new_[4599]_ , \new_[4603]_ , \new_[4604]_ , \new_[4605]_ ,
    \new_[4608]_ , \new_[4611]_ , \new_[4612]_ , \new_[4615]_ ,
    \new_[4619]_ , \new_[4620]_ , \new_[4621]_ , \new_[4624]_ ,
    \new_[4627]_ , \new_[4628]_ , \new_[4631]_ , \new_[4635]_ ,
    \new_[4636]_ , \new_[4637]_ , \new_[4640]_ , \new_[4643]_ ,
    \new_[4644]_ , \new_[4647]_ , \new_[4651]_ , \new_[4652]_ ,
    \new_[4653]_ , \new_[4656]_ , \new_[4659]_ , \new_[4660]_ ,
    \new_[4663]_ , \new_[4667]_ , \new_[4668]_ , \new_[4669]_ ,
    \new_[4672]_ , \new_[4675]_ , \new_[4676]_ , \new_[4679]_ ,
    \new_[4683]_ , \new_[4684]_ , \new_[4685]_ , \new_[4688]_ ,
    \new_[4691]_ , \new_[4692]_ , \new_[4695]_ , \new_[4699]_ ,
    \new_[4700]_ , \new_[4701]_ , \new_[4704]_ , \new_[4707]_ ,
    \new_[4708]_ , \new_[4711]_ , \new_[4715]_ , \new_[4716]_ ,
    \new_[4717]_ , \new_[4720]_ , \new_[4723]_ , \new_[4724]_ ,
    \new_[4727]_ , \new_[4731]_ , \new_[4732]_ , \new_[4733]_ ,
    \new_[4736]_ , \new_[4739]_ , \new_[4740]_ , \new_[4743]_ ,
    \new_[4747]_ , \new_[4748]_ , \new_[4749]_ , \new_[4752]_ ,
    \new_[4755]_ , \new_[4756]_ , \new_[4759]_ , \new_[4763]_ ,
    \new_[4764]_ , \new_[4765]_ , \new_[4768]_ , \new_[4771]_ ,
    \new_[4772]_ , \new_[4775]_ , \new_[4779]_ , \new_[4780]_ ,
    \new_[4781]_ , \new_[4784]_ , \new_[4787]_ , \new_[4788]_ ,
    \new_[4791]_ , \new_[4795]_ , \new_[4796]_ , \new_[4797]_ ,
    \new_[4800]_ , \new_[4803]_ , \new_[4804]_ , \new_[4807]_ ,
    \new_[4811]_ , \new_[4812]_ , \new_[4813]_ , \new_[4816]_ ,
    \new_[4819]_ , \new_[4820]_ , \new_[4823]_ , \new_[4827]_ ,
    \new_[4828]_ , \new_[4829]_ , \new_[4832]_ , \new_[4835]_ ,
    \new_[4836]_ , \new_[4839]_ , \new_[4843]_ , \new_[4844]_ ,
    \new_[4845]_ , \new_[4848]_ , \new_[4851]_ , \new_[4852]_ ,
    \new_[4855]_ , \new_[4859]_ , \new_[4860]_ , \new_[4861]_ ,
    \new_[4864]_ , \new_[4867]_ , \new_[4868]_ , \new_[4871]_ ,
    \new_[4875]_ , \new_[4876]_ , \new_[4877]_ , \new_[4880]_ ,
    \new_[4883]_ , \new_[4884]_ , \new_[4887]_ , \new_[4891]_ ,
    \new_[4892]_ , \new_[4893]_ , \new_[4896]_ , \new_[4899]_ ,
    \new_[4900]_ , \new_[4903]_ , \new_[4907]_ , \new_[4908]_ ,
    \new_[4909]_ , \new_[4912]_ , \new_[4915]_ , \new_[4916]_ ,
    \new_[4919]_ , \new_[4923]_ , \new_[4924]_ , \new_[4925]_ ,
    \new_[4928]_ , \new_[4931]_ , \new_[4932]_ , \new_[4935]_ ,
    \new_[4939]_ , \new_[4940]_ , \new_[4941]_ , \new_[4944]_ ,
    \new_[4947]_ , \new_[4948]_ , \new_[4951]_ , \new_[4955]_ ,
    \new_[4956]_ , \new_[4957]_ , \new_[4960]_ , \new_[4963]_ ,
    \new_[4964]_ , \new_[4967]_ , \new_[4971]_ , \new_[4972]_ ,
    \new_[4973]_ , \new_[4976]_ , \new_[4979]_ , \new_[4980]_ ,
    \new_[4983]_ , \new_[4987]_ , \new_[4988]_ , \new_[4989]_ ,
    \new_[4992]_ , \new_[4996]_ , \new_[4997]_ , \new_[4998]_ ,
    \new_[5001]_ , \new_[5005]_ , \new_[5006]_ , \new_[5007]_ ,
    \new_[5010]_ , \new_[5014]_ , \new_[5015]_ , \new_[5016]_ ,
    \new_[5019]_ , \new_[5023]_ , \new_[5024]_ , \new_[5025]_ ,
    \new_[5028]_ , \new_[5032]_ , \new_[5033]_ , \new_[5034]_ ,
    \new_[5037]_ , \new_[5041]_ , \new_[5042]_ , \new_[5043]_ ,
    \new_[5046]_ , \new_[5050]_ , \new_[5051]_ , \new_[5052]_ ,
    \new_[5055]_ , \new_[5059]_ , \new_[5060]_ , \new_[5061]_ ,
    \new_[5064]_ , \new_[5068]_ , \new_[5069]_ , \new_[5070]_ ,
    \new_[5073]_ , \new_[5077]_ , \new_[5078]_ , \new_[5079]_ ,
    \new_[5082]_ , \new_[5086]_ , \new_[5087]_ , \new_[5088]_ ,
    \new_[5091]_ , \new_[5095]_ , \new_[5096]_ , \new_[5097]_ ,
    \new_[5100]_ , \new_[5104]_ , \new_[5105]_ , \new_[5106]_ ,
    \new_[5109]_ , \new_[5113]_ , \new_[5114]_ , \new_[5115]_ ,
    \new_[5118]_ , \new_[5122]_ , \new_[5123]_ , \new_[5124]_ ,
    \new_[5127]_ , \new_[5131]_ , \new_[5132]_ , \new_[5133]_ ,
    \new_[5136]_ , \new_[5140]_ , \new_[5141]_ , \new_[5142]_ ,
    \new_[5145]_ , \new_[5149]_ , \new_[5150]_ , \new_[5151]_ ,
    \new_[5154]_ , \new_[5158]_ , \new_[5159]_ , \new_[5160]_ ,
    \new_[5163]_ , \new_[5167]_ , \new_[5168]_ , \new_[5169]_ ,
    \new_[5172]_ , \new_[5176]_ , \new_[5177]_ , \new_[5178]_ ,
    \new_[5181]_ , \new_[5185]_ , \new_[5186]_ , \new_[5187]_ ,
    \new_[5190]_ , \new_[5194]_ , \new_[5195]_ , \new_[5196]_ ,
    \new_[5199]_ , \new_[5203]_ , \new_[5204]_ , \new_[5205]_ ,
    \new_[5208]_ , \new_[5212]_ , \new_[5213]_ , \new_[5214]_ ,
    \new_[5217]_ , \new_[5221]_ , \new_[5222]_ , \new_[5223]_ ,
    \new_[5226]_ , \new_[5230]_ , \new_[5231]_ , \new_[5232]_ ,
    \new_[5235]_ , \new_[5239]_ , \new_[5240]_ , \new_[5241]_ ,
    \new_[5244]_ , \new_[5248]_ , \new_[5249]_ , \new_[5250]_ ,
    \new_[5253]_ , \new_[5257]_ , \new_[5258]_ , \new_[5259]_ ,
    \new_[5262]_ , \new_[5266]_ , \new_[5267]_ , \new_[5268]_ ,
    \new_[5271]_ , \new_[5275]_ , \new_[5276]_ , \new_[5277]_ ,
    \new_[5280]_ , \new_[5284]_ , \new_[5285]_ , \new_[5286]_ ,
    \new_[5289]_ , \new_[5293]_ , \new_[5294]_ , \new_[5295]_ ,
    \new_[5298]_ , \new_[5302]_ , \new_[5303]_ , \new_[5304]_ ,
    \new_[5307]_ , \new_[5311]_ , \new_[5312]_ , \new_[5313]_ ,
    \new_[5316]_ , \new_[5320]_ , \new_[5321]_ , \new_[5322]_ ,
    \new_[5325]_ , \new_[5329]_ , \new_[5330]_ , \new_[5331]_ ,
    \new_[5334]_ , \new_[5338]_ , \new_[5339]_ , \new_[5340]_ ,
    \new_[5343]_ , \new_[5347]_ , \new_[5348]_ , \new_[5349]_ ,
    \new_[5352]_ , \new_[5356]_ , \new_[5357]_ , \new_[5358]_ ,
    \new_[5361]_ , \new_[5365]_ , \new_[5366]_ , \new_[5367]_ ,
    \new_[5370]_ , \new_[5374]_ , \new_[5375]_ , \new_[5376]_ ,
    \new_[5379]_ , \new_[5383]_ , \new_[5384]_ , \new_[5385]_ ,
    \new_[5388]_ , \new_[5392]_ , \new_[5393]_ , \new_[5394]_ ,
    \new_[5397]_ , \new_[5401]_ , \new_[5402]_ , \new_[5403]_ ,
    \new_[5406]_ , \new_[5410]_ , \new_[5411]_ , \new_[5412]_ ,
    \new_[5415]_ , \new_[5419]_ , \new_[5420]_ , \new_[5421]_ ,
    \new_[5424]_ , \new_[5428]_ , \new_[5429]_ , \new_[5430]_ ,
    \new_[5433]_ , \new_[5437]_ , \new_[5438]_ , \new_[5439]_ ,
    \new_[5442]_ , \new_[5446]_ , \new_[5447]_ , \new_[5448]_ ,
    \new_[5451]_ , \new_[5455]_ , \new_[5456]_ , \new_[5457]_ ,
    \new_[5460]_ , \new_[5464]_ , \new_[5465]_ , \new_[5466]_ ,
    \new_[5469]_ , \new_[5473]_ , \new_[5474]_ , \new_[5475]_ ,
    \new_[5478]_ , \new_[5482]_ , \new_[5483]_ , \new_[5484]_ ,
    \new_[5487]_ , \new_[5491]_ , \new_[5492]_ , \new_[5493]_ ,
    \new_[5496]_ , \new_[5500]_ , \new_[5501]_ , \new_[5502]_ ,
    \new_[5505]_ , \new_[5509]_ , \new_[5510]_ , \new_[5511]_ ,
    \new_[5514]_ , \new_[5518]_ , \new_[5519]_ , \new_[5520]_ ,
    \new_[5523]_ , \new_[5527]_ , \new_[5528]_ , \new_[5529]_ ,
    \new_[5532]_ , \new_[5536]_ , \new_[5537]_ , \new_[5538]_ ,
    \new_[5541]_ , \new_[5545]_ , \new_[5546]_ , \new_[5547]_ ,
    \new_[5550]_ , \new_[5554]_ , \new_[5555]_ , \new_[5556]_ ,
    \new_[5559]_ , \new_[5563]_ , \new_[5564]_ , \new_[5565]_ ,
    \new_[5568]_ , \new_[5572]_ , \new_[5573]_ , \new_[5574]_ ,
    \new_[5577]_ , \new_[5581]_ , \new_[5582]_ , \new_[5583]_ ,
    \new_[5586]_ , \new_[5590]_ , \new_[5591]_ , \new_[5592]_ ,
    \new_[5595]_ , \new_[5599]_ , \new_[5600]_ , \new_[5601]_ ,
    \new_[5604]_ , \new_[5608]_ , \new_[5609]_ , \new_[5610]_ ,
    \new_[5613]_ , \new_[5617]_ , \new_[5618]_ , \new_[5619]_ ,
    \new_[5622]_ , \new_[5626]_ , \new_[5627]_ , \new_[5628]_ ,
    \new_[5631]_ , \new_[5635]_ , \new_[5636]_ , \new_[5637]_ ,
    \new_[5640]_ , \new_[5644]_ , \new_[5645]_ , \new_[5646]_ ,
    \new_[5649]_ , \new_[5653]_ , \new_[5654]_ , \new_[5655]_ ,
    \new_[5658]_ , \new_[5662]_ , \new_[5663]_ , \new_[5664]_ ,
    \new_[5667]_ , \new_[5671]_ , \new_[5672]_ , \new_[5673]_ ,
    \new_[5676]_ , \new_[5680]_ , \new_[5681]_ , \new_[5682]_ ,
    \new_[5685]_ , \new_[5689]_ , \new_[5690]_ , \new_[5691]_ ,
    \new_[5694]_ , \new_[5698]_ , \new_[5699]_ , \new_[5700]_ ,
    \new_[5703]_ , \new_[5707]_ , \new_[5708]_ , \new_[5709]_ ,
    \new_[5712]_ , \new_[5716]_ , \new_[5717]_ , \new_[5718]_ ,
    \new_[5721]_ , \new_[5725]_ , \new_[5726]_ , \new_[5727]_ ,
    \new_[5730]_ , \new_[5734]_ , \new_[5735]_ , \new_[5736]_ ,
    \new_[5739]_ , \new_[5743]_ , \new_[5744]_ , \new_[5745]_ ,
    \new_[5748]_ , \new_[5752]_ , \new_[5753]_ , \new_[5754]_ ,
    \new_[5757]_ , \new_[5761]_ , \new_[5762]_ , \new_[5763]_ ,
    \new_[5766]_ , \new_[5770]_ , \new_[5771]_ , \new_[5772]_ ,
    \new_[5775]_ , \new_[5779]_ , \new_[5780]_ , \new_[5781]_ ,
    \new_[5784]_ , \new_[5788]_ , \new_[5789]_ , \new_[5790]_ ,
    \new_[5793]_ , \new_[5797]_ , \new_[5798]_ , \new_[5799]_ ,
    \new_[5802]_ , \new_[5806]_ , \new_[5807]_ , \new_[5808]_ ,
    \new_[5811]_ , \new_[5815]_ , \new_[5816]_ , \new_[5817]_ ,
    \new_[5820]_ , \new_[5824]_ , \new_[5825]_ , \new_[5826]_ ,
    \new_[5829]_ , \new_[5833]_ , \new_[5834]_ , \new_[5835]_ ,
    \new_[5838]_ , \new_[5842]_ , \new_[5843]_ , \new_[5844]_ ,
    \new_[5847]_ , \new_[5851]_ , \new_[5852]_ , \new_[5853]_ ,
    \new_[5856]_ , \new_[5860]_ , \new_[5861]_ , \new_[5862]_ ,
    \new_[5865]_ , \new_[5869]_ , \new_[5870]_ , \new_[5871]_ ,
    \new_[5874]_ , \new_[5878]_ , \new_[5879]_ , \new_[5880]_ ,
    \new_[5883]_ , \new_[5887]_ , \new_[5888]_ , \new_[5889]_ ,
    \new_[5892]_ , \new_[5896]_ , \new_[5897]_ , \new_[5898]_ ,
    \new_[5901]_ , \new_[5905]_ , \new_[5906]_ , \new_[5907]_ ,
    \new_[5910]_ , \new_[5914]_ , \new_[5915]_ , \new_[5916]_ ,
    \new_[5919]_ , \new_[5923]_ , \new_[5924]_ , \new_[5925]_ ,
    \new_[5928]_ , \new_[5932]_ , \new_[5933]_ , \new_[5934]_ ,
    \new_[5937]_ , \new_[5941]_ , \new_[5942]_ , \new_[5943]_ ,
    \new_[5946]_ , \new_[5950]_ , \new_[5951]_ , \new_[5952]_ ,
    \new_[5955]_ , \new_[5959]_ , \new_[5960]_ , \new_[5961]_ ,
    \new_[5964]_ , \new_[5968]_ , \new_[5969]_ , \new_[5970]_ ,
    \new_[5973]_ , \new_[5977]_ , \new_[5978]_ , \new_[5979]_ ,
    \new_[5982]_ , \new_[5986]_ , \new_[5987]_ , \new_[5988]_ ,
    \new_[5991]_ , \new_[5995]_ , \new_[5996]_ , \new_[5997]_ ,
    \new_[6000]_ , \new_[6004]_ , \new_[6005]_ , \new_[6006]_ ,
    \new_[6009]_ , \new_[6013]_ , \new_[6014]_ , \new_[6015]_ ,
    \new_[6018]_ , \new_[6022]_ , \new_[6023]_ , \new_[6024]_ ,
    \new_[6027]_ , \new_[6031]_ , \new_[6032]_ , \new_[6033]_ ,
    \new_[6036]_ , \new_[6040]_ , \new_[6041]_ , \new_[6042]_ ,
    \new_[6045]_ , \new_[6049]_ , \new_[6050]_ , \new_[6051]_ ,
    \new_[6054]_ , \new_[6058]_ , \new_[6059]_ , \new_[6060]_ ,
    \new_[6063]_ , \new_[6067]_ , \new_[6068]_ , \new_[6069]_ ,
    \new_[6072]_ , \new_[6076]_ , \new_[6077]_ , \new_[6078]_ ,
    \new_[6081]_ , \new_[6085]_ , \new_[6086]_ , \new_[6087]_ ,
    \new_[6090]_ , \new_[6094]_ , \new_[6095]_ , \new_[6096]_ ,
    \new_[6099]_ , \new_[6103]_ , \new_[6104]_ , \new_[6105]_ ,
    \new_[6108]_ , \new_[6112]_ , \new_[6113]_ , \new_[6114]_ ,
    \new_[6117]_ , \new_[6121]_ , \new_[6122]_ , \new_[6123]_ ,
    \new_[6126]_ , \new_[6130]_ , \new_[6131]_ , \new_[6132]_ ,
    \new_[6135]_ , \new_[6139]_ , \new_[6140]_ , \new_[6141]_ ,
    \new_[6144]_ , \new_[6148]_ , \new_[6149]_ , \new_[6150]_ ,
    \new_[6153]_ , \new_[6157]_ , \new_[6158]_ , \new_[6159]_ ,
    \new_[6162]_ , \new_[6166]_ , \new_[6167]_ , \new_[6168]_ ,
    \new_[6171]_ , \new_[6175]_ , \new_[6176]_ , \new_[6177]_ ,
    \new_[6180]_ , \new_[6184]_ , \new_[6185]_ , \new_[6186]_ ,
    \new_[6189]_ , \new_[6193]_ , \new_[6194]_ , \new_[6195]_ ,
    \new_[6198]_ , \new_[6202]_ , \new_[6203]_ , \new_[6204]_ ,
    \new_[6207]_ , \new_[6211]_ , \new_[6212]_ , \new_[6213]_ ,
    \new_[6216]_ , \new_[6220]_ , \new_[6221]_ , \new_[6222]_ ,
    \new_[6225]_ , \new_[6229]_ , \new_[6230]_ , \new_[6231]_ ,
    \new_[6234]_ , \new_[6238]_ , \new_[6239]_ , \new_[6240]_ ,
    \new_[6243]_ , \new_[6247]_ , \new_[6248]_ , \new_[6249]_ ,
    \new_[6252]_ , \new_[6256]_ , \new_[6257]_ , \new_[6258]_ ,
    \new_[6261]_ , \new_[6265]_ , \new_[6266]_ , \new_[6267]_ ,
    \new_[6270]_ , \new_[6274]_ , \new_[6275]_ , \new_[6276]_ ,
    \new_[6279]_ , \new_[6283]_ , \new_[6284]_ , \new_[6285]_ ,
    \new_[6288]_ , \new_[6292]_ , \new_[6293]_ , \new_[6294]_ ,
    \new_[6297]_ , \new_[6301]_ , \new_[6302]_ , \new_[6303]_ ,
    \new_[6306]_ , \new_[6310]_ , \new_[6311]_ , \new_[6312]_ ,
    \new_[6315]_ , \new_[6319]_ , \new_[6320]_ , \new_[6321]_ ,
    \new_[6324]_ , \new_[6328]_ , \new_[6329]_ , \new_[6330]_ ,
    \new_[6333]_ , \new_[6337]_ , \new_[6338]_ , \new_[6339]_ ,
    \new_[6342]_ , \new_[6346]_ , \new_[6347]_ , \new_[6348]_ ,
    \new_[6351]_ , \new_[6355]_ , \new_[6356]_ , \new_[6357]_ ,
    \new_[6360]_ , \new_[6364]_ , \new_[6365]_ , \new_[6366]_ ,
    \new_[6369]_ , \new_[6373]_ , \new_[6374]_ , \new_[6375]_ ,
    \new_[6378]_ , \new_[6382]_ , \new_[6383]_ , \new_[6384]_ ,
    \new_[6387]_ , \new_[6391]_ , \new_[6392]_ , \new_[6393]_ ,
    \new_[6396]_ , \new_[6400]_ , \new_[6401]_ , \new_[6402]_ ,
    \new_[6405]_ , \new_[6409]_ , \new_[6410]_ , \new_[6411]_ ,
    \new_[6414]_ , \new_[6418]_ , \new_[6419]_ , \new_[6420]_ ,
    \new_[6423]_ , \new_[6427]_ , \new_[6428]_ , \new_[6429]_ ,
    \new_[6432]_ , \new_[6436]_ , \new_[6437]_ , \new_[6438]_ ,
    \new_[6441]_ , \new_[6445]_ , \new_[6446]_ , \new_[6447]_ ,
    \new_[6450]_ , \new_[6454]_ , \new_[6455]_ , \new_[6456]_ ,
    \new_[6459]_ , \new_[6463]_ , \new_[6464]_ , \new_[6465]_ ,
    \new_[6468]_ , \new_[6472]_ , \new_[6473]_ , \new_[6474]_ ,
    \new_[6477]_ , \new_[6481]_ , \new_[6482]_ , \new_[6483]_ ,
    \new_[6486]_ , \new_[6490]_ , \new_[6491]_ , \new_[6492]_ ,
    \new_[6495]_ , \new_[6499]_ , \new_[6500]_ , \new_[6501]_ ,
    \new_[6504]_ , \new_[6508]_ , \new_[6509]_ , \new_[6510]_ ,
    \new_[6513]_ , \new_[6517]_ , \new_[6518]_ , \new_[6519]_ ,
    \new_[6522]_ , \new_[6526]_ , \new_[6527]_ , \new_[6528]_ ,
    \new_[6531]_ , \new_[6535]_ , \new_[6536]_ , \new_[6537]_ ,
    \new_[6540]_ , \new_[6544]_ , \new_[6545]_ , \new_[6546]_ ,
    \new_[6549]_ , \new_[6553]_ , \new_[6554]_ , \new_[6555]_ ,
    \new_[6558]_ , \new_[6562]_ , \new_[6563]_ , \new_[6564]_ ,
    \new_[6567]_ , \new_[6571]_ , \new_[6572]_ , \new_[6573]_ ,
    \new_[6576]_ , \new_[6580]_ , \new_[6581]_ , \new_[6582]_ ,
    \new_[6585]_ , \new_[6589]_ , \new_[6590]_ , \new_[6591]_ ,
    \new_[6594]_ , \new_[6598]_ , \new_[6599]_ , \new_[6600]_ ,
    \new_[6603]_ , \new_[6607]_ , \new_[6608]_ , \new_[6609]_ ,
    \new_[6612]_ , \new_[6616]_ , \new_[6617]_ , \new_[6618]_ ,
    \new_[6621]_ , \new_[6625]_ , \new_[6626]_ , \new_[6627]_ ,
    \new_[6630]_ , \new_[6634]_ , \new_[6635]_ , \new_[6636]_ ,
    \new_[6639]_ , \new_[6643]_ , \new_[6644]_ , \new_[6645]_ ,
    \new_[6648]_ , \new_[6652]_ , \new_[6653]_ , \new_[6654]_ ,
    \new_[6657]_ , \new_[6661]_ , \new_[6662]_ , \new_[6663]_ ,
    \new_[6666]_ , \new_[6670]_ , \new_[6671]_ , \new_[6672]_ ,
    \new_[6675]_ , \new_[6679]_ , \new_[6680]_ , \new_[6681]_ ,
    \new_[6684]_ , \new_[6688]_ , \new_[6689]_ , \new_[6690]_ ,
    \new_[6693]_ , \new_[6697]_ , \new_[6698]_ , \new_[6699]_ ,
    \new_[6702]_ , \new_[6706]_ , \new_[6707]_ , \new_[6708]_ ,
    \new_[6711]_ , \new_[6715]_ , \new_[6716]_ , \new_[6717]_ ,
    \new_[6720]_ , \new_[6724]_ , \new_[6725]_ , \new_[6726]_ ,
    \new_[6729]_ , \new_[6733]_ , \new_[6734]_ , \new_[6735]_ ,
    \new_[6738]_ , \new_[6742]_ , \new_[6743]_ , \new_[6744]_ ,
    \new_[6747]_ , \new_[6751]_ , \new_[6752]_ , \new_[6753]_ ,
    \new_[6756]_ , \new_[6760]_ , \new_[6761]_ , \new_[6762]_ ,
    \new_[6765]_ , \new_[6769]_ , \new_[6770]_ , \new_[6771]_ ,
    \new_[6774]_ , \new_[6778]_ , \new_[6779]_ , \new_[6780]_ ,
    \new_[6783]_ , \new_[6787]_ , \new_[6788]_ , \new_[6789]_ ,
    \new_[6792]_ , \new_[6796]_ , \new_[6797]_ , \new_[6798]_ ,
    \new_[6801]_ , \new_[6805]_ , \new_[6806]_ , \new_[6807]_ ,
    \new_[6810]_ , \new_[6814]_ , \new_[6815]_ , \new_[6816]_ ,
    \new_[6819]_ , \new_[6823]_ , \new_[6824]_ , \new_[6825]_ ,
    \new_[6828]_ , \new_[6832]_ , \new_[6833]_ , \new_[6834]_ ,
    \new_[6837]_ , \new_[6841]_ , \new_[6842]_ , \new_[6843]_ ,
    \new_[6846]_ , \new_[6850]_ , \new_[6851]_ , \new_[6852]_ ,
    \new_[6855]_ , \new_[6859]_ , \new_[6860]_ , \new_[6861]_ ,
    \new_[6864]_ , \new_[6868]_ , \new_[6869]_ , \new_[6870]_ ,
    \new_[6873]_ , \new_[6877]_ , \new_[6878]_ , \new_[6879]_ ,
    \new_[6882]_ , \new_[6886]_ , \new_[6887]_ , \new_[6888]_ ,
    \new_[6891]_ , \new_[6895]_ , \new_[6896]_ , \new_[6897]_ ,
    \new_[6900]_ , \new_[6904]_ , \new_[6905]_ , \new_[6906]_ ,
    \new_[6909]_ , \new_[6913]_ , \new_[6914]_ , \new_[6915]_ ,
    \new_[6918]_ , \new_[6922]_ , \new_[6923]_ , \new_[6924]_ ,
    \new_[6927]_ , \new_[6931]_ , \new_[6932]_ , \new_[6933]_ ,
    \new_[6936]_ , \new_[6940]_ , \new_[6941]_ , \new_[6942]_ ,
    \new_[6945]_ , \new_[6949]_ , \new_[6950]_ , \new_[6951]_ ,
    \new_[6954]_ , \new_[6958]_ , \new_[6959]_ , \new_[6960]_ ,
    \new_[6963]_ , \new_[6967]_ , \new_[6968]_ , \new_[6969]_ ,
    \new_[6972]_ , \new_[6976]_ , \new_[6977]_ , \new_[6978]_ ,
    \new_[6981]_ , \new_[6985]_ , \new_[6986]_ , \new_[6987]_ ,
    \new_[6990]_ , \new_[6994]_ , \new_[6995]_ , \new_[6996]_ ,
    \new_[6999]_ , \new_[7003]_ , \new_[7004]_ , \new_[7005]_ ,
    \new_[7008]_ , \new_[7012]_ , \new_[7013]_ , \new_[7014]_ ,
    \new_[7017]_ , \new_[7021]_ , \new_[7022]_ , \new_[7023]_ ,
    \new_[7026]_ , \new_[7030]_ , \new_[7031]_ , \new_[7032]_ ,
    \new_[7035]_ , \new_[7039]_ , \new_[7040]_ , \new_[7041]_ ,
    \new_[7044]_ , \new_[7048]_ , \new_[7049]_ , \new_[7050]_ ,
    \new_[7053]_ , \new_[7057]_ , \new_[7058]_ , \new_[7059]_ ,
    \new_[7062]_ , \new_[7066]_ , \new_[7067]_ , \new_[7068]_ ,
    \new_[7071]_ , \new_[7075]_ , \new_[7076]_ , \new_[7077]_ ,
    \new_[7080]_ , \new_[7084]_ , \new_[7085]_ , \new_[7086]_ ,
    \new_[7089]_ , \new_[7093]_ , \new_[7094]_ , \new_[7095]_ ,
    \new_[7098]_ , \new_[7102]_ , \new_[7103]_ , \new_[7104]_ ,
    \new_[7107]_ , \new_[7111]_ , \new_[7112]_ , \new_[7113]_ ,
    \new_[7116]_ , \new_[7120]_ , \new_[7121]_ , \new_[7122]_ ,
    \new_[7125]_ , \new_[7129]_ , \new_[7130]_ , \new_[7131]_ ,
    \new_[7134]_ , \new_[7138]_ , \new_[7139]_ , \new_[7140]_ ,
    \new_[7143]_ , \new_[7147]_ , \new_[7148]_ , \new_[7149]_ ,
    \new_[7152]_ , \new_[7156]_ , \new_[7157]_ , \new_[7158]_ ,
    \new_[7161]_ , \new_[7165]_ , \new_[7166]_ , \new_[7167]_ ,
    \new_[7170]_ , \new_[7174]_ , \new_[7175]_ , \new_[7176]_ ,
    \new_[7179]_ , \new_[7183]_ , \new_[7184]_ , \new_[7185]_ ,
    \new_[7188]_ , \new_[7192]_ , \new_[7193]_ , \new_[7194]_ ,
    \new_[7197]_ , \new_[7201]_ , \new_[7202]_ , \new_[7203]_ ,
    \new_[7206]_ , \new_[7210]_ , \new_[7211]_ , \new_[7212]_ ,
    \new_[7215]_ , \new_[7219]_ , \new_[7220]_ , \new_[7221]_ ,
    \new_[7224]_ , \new_[7228]_ , \new_[7229]_ , \new_[7230]_ ,
    \new_[7233]_ , \new_[7237]_ , \new_[7238]_ , \new_[7239]_ ,
    \new_[7242]_ , \new_[7246]_ , \new_[7247]_ , \new_[7248]_ ,
    \new_[7251]_ , \new_[7255]_ , \new_[7256]_ , \new_[7257]_ ,
    \new_[7260]_ , \new_[7264]_ , \new_[7265]_ , \new_[7266]_ ,
    \new_[7269]_ , \new_[7273]_ , \new_[7274]_ , \new_[7275]_ ,
    \new_[7278]_ , \new_[7282]_ , \new_[7283]_ , \new_[7284]_ ,
    \new_[7287]_ , \new_[7291]_ , \new_[7292]_ , \new_[7293]_ ,
    \new_[7296]_ , \new_[7300]_ , \new_[7301]_ , \new_[7302]_ ,
    \new_[7305]_ , \new_[7309]_ , \new_[7310]_ , \new_[7311]_ ,
    \new_[7314]_ , \new_[7318]_ , \new_[7319]_ , \new_[7320]_ ,
    \new_[7323]_ , \new_[7327]_ , \new_[7328]_ , \new_[7329]_ ,
    \new_[7332]_ , \new_[7336]_ , \new_[7337]_ , \new_[7338]_ ,
    \new_[7341]_ , \new_[7345]_ , \new_[7346]_ , \new_[7347]_ ,
    \new_[7350]_ , \new_[7354]_ , \new_[7355]_ , \new_[7356]_ ,
    \new_[7359]_ , \new_[7363]_ , \new_[7364]_ , \new_[7365]_ ,
    \new_[7368]_ , \new_[7372]_ , \new_[7373]_ , \new_[7374]_ ,
    \new_[7377]_ , \new_[7381]_ , \new_[7382]_ , \new_[7383]_ ,
    \new_[7386]_ , \new_[7390]_ , \new_[7391]_ , \new_[7392]_ ,
    \new_[7395]_ , \new_[7399]_ , \new_[7400]_ , \new_[7401]_ ,
    \new_[7404]_ , \new_[7408]_ , \new_[7409]_ , \new_[7410]_ ,
    \new_[7413]_ , \new_[7417]_ , \new_[7418]_ , \new_[7419]_ ,
    \new_[7422]_ , \new_[7426]_ , \new_[7427]_ , \new_[7428]_ ,
    \new_[7431]_ , \new_[7435]_ , \new_[7436]_ , \new_[7437]_ ,
    \new_[7440]_ , \new_[7444]_ , \new_[7445]_ , \new_[7446]_ ,
    \new_[7449]_ , \new_[7453]_ , \new_[7454]_ , \new_[7455]_ ,
    \new_[7458]_ , \new_[7462]_ , \new_[7463]_ , \new_[7464]_ ,
    \new_[7467]_ , \new_[7471]_ , \new_[7472]_ , \new_[7473]_ ,
    \new_[7476]_ , \new_[7480]_ , \new_[7481]_ , \new_[7482]_ ,
    \new_[7485]_ , \new_[7489]_ , \new_[7490]_ , \new_[7491]_ ,
    \new_[7494]_ , \new_[7498]_ , \new_[7499]_ , \new_[7500]_ ,
    \new_[7503]_ , \new_[7507]_ , \new_[7508]_ , \new_[7509]_ ,
    \new_[7512]_ , \new_[7516]_ , \new_[7517]_ , \new_[7518]_ ,
    \new_[7521]_ , \new_[7525]_ , \new_[7526]_ , \new_[7527]_ ,
    \new_[7530]_ , \new_[7534]_ , \new_[7535]_ , \new_[7536]_ ,
    \new_[7539]_ , \new_[7543]_ , \new_[7544]_ , \new_[7545]_ ,
    \new_[7548]_ , \new_[7552]_ , \new_[7553]_ , \new_[7554]_ ,
    \new_[7557]_ , \new_[7561]_ , \new_[7562]_ , \new_[7563]_ ,
    \new_[7566]_ , \new_[7570]_ , \new_[7571]_ , \new_[7572]_ ,
    \new_[7575]_ , \new_[7579]_ , \new_[7580]_ , \new_[7581]_ ,
    \new_[7584]_ , \new_[7588]_ , \new_[7589]_ , \new_[7590]_ ,
    \new_[7593]_ , \new_[7597]_ , \new_[7598]_ , \new_[7599]_ ,
    \new_[7602]_ , \new_[7606]_ , \new_[7607]_ , \new_[7608]_ ,
    \new_[7611]_ , \new_[7615]_ , \new_[7616]_ , \new_[7617]_ ,
    \new_[7620]_ , \new_[7624]_ , \new_[7625]_ , \new_[7626]_ ,
    \new_[7629]_ , \new_[7633]_ , \new_[7634]_ , \new_[7635]_ ,
    \new_[7638]_ , \new_[7642]_ , \new_[7643]_ , \new_[7644]_ ,
    \new_[7647]_ , \new_[7651]_ , \new_[7652]_ , \new_[7653]_ ,
    \new_[7656]_ , \new_[7660]_ , \new_[7661]_ , \new_[7662]_ ,
    \new_[7665]_ , \new_[7669]_ , \new_[7670]_ , \new_[7671]_ ,
    \new_[7674]_ , \new_[7678]_ , \new_[7679]_ , \new_[7680]_ ,
    \new_[7683]_ , \new_[7687]_ , \new_[7688]_ , \new_[7689]_ ,
    \new_[7692]_ , \new_[7696]_ , \new_[7697]_ , \new_[7698]_ ,
    \new_[7701]_ , \new_[7705]_ , \new_[7706]_ , \new_[7707]_ ,
    \new_[7710]_ , \new_[7714]_ , \new_[7715]_ , \new_[7716]_ ,
    \new_[7719]_ , \new_[7723]_ , \new_[7724]_ , \new_[7725]_ ,
    \new_[7728]_ , \new_[7732]_ , \new_[7733]_ , \new_[7734]_ ,
    \new_[7737]_ , \new_[7741]_ , \new_[7742]_ , \new_[7743]_ ,
    \new_[7746]_ , \new_[7750]_ , \new_[7751]_ , \new_[7752]_ ,
    \new_[7755]_ , \new_[7759]_ , \new_[7760]_ , \new_[7761]_ ,
    \new_[7764]_ , \new_[7768]_ , \new_[7769]_ , \new_[7770]_ ,
    \new_[7773]_ , \new_[7777]_ , \new_[7778]_ , \new_[7779]_ ,
    \new_[7782]_ , \new_[7786]_ , \new_[7787]_ , \new_[7788]_ ,
    \new_[7791]_ , \new_[7795]_ , \new_[7796]_ , \new_[7797]_ ,
    \new_[7800]_ , \new_[7804]_ , \new_[7805]_ , \new_[7806]_ ,
    \new_[7809]_ , \new_[7813]_ , \new_[7814]_ , \new_[7815]_ ,
    \new_[7818]_ , \new_[7822]_ , \new_[7823]_ , \new_[7824]_ ,
    \new_[7827]_ , \new_[7831]_ , \new_[7832]_ , \new_[7833]_ ,
    \new_[7836]_ , \new_[7840]_ , \new_[7841]_ , \new_[7842]_ ,
    \new_[7845]_ , \new_[7849]_ , \new_[7850]_ , \new_[7851]_ ,
    \new_[7854]_ , \new_[7858]_ , \new_[7859]_ , \new_[7860]_ ,
    \new_[7863]_ , \new_[7867]_ , \new_[7868]_ , \new_[7869]_ ,
    \new_[7872]_ , \new_[7876]_ , \new_[7877]_ , \new_[7878]_ ,
    \new_[7881]_ , \new_[7885]_ , \new_[7886]_ , \new_[7887]_ ,
    \new_[7890]_ , \new_[7894]_ , \new_[7895]_ , \new_[7896]_ ,
    \new_[7899]_ , \new_[7903]_ , \new_[7904]_ , \new_[7905]_ ,
    \new_[7908]_ , \new_[7912]_ , \new_[7913]_ , \new_[7914]_ ,
    \new_[7917]_ , \new_[7921]_ , \new_[7922]_ , \new_[7923]_ ,
    \new_[7926]_ , \new_[7930]_ , \new_[7931]_ , \new_[7932]_ ,
    \new_[7935]_ , \new_[7939]_ , \new_[7940]_ , \new_[7941]_ ,
    \new_[7944]_ , \new_[7948]_ , \new_[7949]_ , \new_[7950]_ ,
    \new_[7953]_ , \new_[7957]_ , \new_[7958]_ , \new_[7959]_ ,
    \new_[7962]_ , \new_[7966]_ , \new_[7967]_ , \new_[7968]_ ,
    \new_[7971]_ , \new_[7975]_ , \new_[7976]_ , \new_[7977]_ ,
    \new_[7980]_ , \new_[7984]_ , \new_[7985]_ , \new_[7986]_ ,
    \new_[7989]_ , \new_[7993]_ , \new_[7994]_ , \new_[7995]_ ,
    \new_[7998]_ , \new_[8002]_ , \new_[8003]_ , \new_[8004]_ ,
    \new_[8007]_ , \new_[8011]_ , \new_[8012]_ , \new_[8013]_ ,
    \new_[8016]_ , \new_[8020]_ , \new_[8021]_ , \new_[8022]_ ,
    \new_[8025]_ , \new_[8029]_ , \new_[8030]_ , \new_[8031]_ ,
    \new_[8034]_ , \new_[8038]_ , \new_[8039]_ , \new_[8040]_ ,
    \new_[8043]_ , \new_[8047]_ , \new_[8048]_ , \new_[8049]_ ,
    \new_[8052]_ , \new_[8056]_ , \new_[8057]_ , \new_[8058]_ ,
    \new_[8061]_ , \new_[8065]_ , \new_[8066]_ , \new_[8067]_ ,
    \new_[8070]_ , \new_[8074]_ , \new_[8075]_ , \new_[8076]_ ,
    \new_[8079]_ , \new_[8083]_ , \new_[8084]_ , \new_[8085]_ ,
    \new_[8088]_ , \new_[8092]_ , \new_[8093]_ , \new_[8094]_ ,
    \new_[8097]_ , \new_[8101]_ , \new_[8102]_ , \new_[8103]_ ,
    \new_[8106]_ , \new_[8110]_ , \new_[8111]_ , \new_[8112]_ ,
    \new_[8115]_ , \new_[8119]_ , \new_[8120]_ , \new_[8121]_ ,
    \new_[8124]_ , \new_[8128]_ , \new_[8129]_ , \new_[8130]_ ,
    \new_[8134]_ , \new_[8135]_ , \new_[8139]_ , \new_[8140]_ ,
    \new_[8141]_ , \new_[8144]_ , \new_[8148]_ , \new_[8149]_ ,
    \new_[8150]_ , \new_[8154]_ , \new_[8155]_ , \new_[8159]_ ,
    \new_[8160]_ , \new_[8161]_ , \new_[8164]_ , \new_[8168]_ ,
    \new_[8169]_ , \new_[8170]_ , \new_[8174]_ , \new_[8175]_ ,
    \new_[8179]_ , \new_[8180]_ , \new_[8181]_ , \new_[8184]_ ,
    \new_[8188]_ , \new_[8189]_ , \new_[8190]_ , \new_[8194]_ ,
    \new_[8195]_ , \new_[8199]_ , \new_[8200]_ , \new_[8201]_ ,
    \new_[8204]_ , \new_[8208]_ , \new_[8209]_ , \new_[8210]_ ,
    \new_[8214]_ , \new_[8215]_ , \new_[8219]_ , \new_[8220]_ ,
    \new_[8221]_ , \new_[8224]_ , \new_[8228]_ , \new_[8229]_ ,
    \new_[8230]_ , \new_[8234]_ , \new_[8235]_ , \new_[8239]_ ,
    \new_[8240]_ , \new_[8241]_ , \new_[8244]_ , \new_[8248]_ ,
    \new_[8249]_ , \new_[8250]_ , \new_[8254]_ , \new_[8255]_ ,
    \new_[8259]_ , \new_[8260]_ , \new_[8261]_ , \new_[8264]_ ,
    \new_[8268]_ , \new_[8269]_ , \new_[8270]_ , \new_[8274]_ ,
    \new_[8275]_ , \new_[8279]_ , \new_[8280]_ , \new_[8281]_ ,
    \new_[8284]_ , \new_[8288]_ , \new_[8289]_ , \new_[8290]_ ,
    \new_[8294]_ , \new_[8295]_ , \new_[8299]_ , \new_[8300]_ ,
    \new_[8301]_ , \new_[8304]_ , \new_[8308]_ , \new_[8309]_ ,
    \new_[8310]_ , \new_[8314]_ , \new_[8315]_ , \new_[8319]_ ,
    \new_[8320]_ , \new_[8321]_ , \new_[8324]_ , \new_[8328]_ ,
    \new_[8329]_ , \new_[8330]_ , \new_[8334]_ , \new_[8335]_ ,
    \new_[8339]_ , \new_[8340]_ , \new_[8341]_ , \new_[8344]_ ,
    \new_[8348]_ , \new_[8349]_ , \new_[8350]_ , \new_[8354]_ ,
    \new_[8355]_ , \new_[8359]_ , \new_[8360]_ , \new_[8361]_ ,
    \new_[8364]_ , \new_[8368]_ , \new_[8369]_ , \new_[8370]_ ,
    \new_[8374]_ , \new_[8375]_ , \new_[8379]_ , \new_[8380]_ ,
    \new_[8381]_ , \new_[8384]_ , \new_[8388]_ , \new_[8389]_ ,
    \new_[8390]_ , \new_[8394]_ , \new_[8395]_ , \new_[8399]_ ,
    \new_[8400]_ , \new_[8401]_ , \new_[8404]_ , \new_[8408]_ ,
    \new_[8409]_ , \new_[8410]_ , \new_[8414]_ , \new_[8415]_ ,
    \new_[8419]_ , \new_[8420]_ , \new_[8421]_ , \new_[8424]_ ,
    \new_[8428]_ , \new_[8429]_ , \new_[8430]_ , \new_[8434]_ ,
    \new_[8435]_ , \new_[8439]_ , \new_[8440]_ , \new_[8441]_ ,
    \new_[8444]_ , \new_[8448]_ , \new_[8449]_ , \new_[8450]_ ,
    \new_[8454]_ , \new_[8455]_ , \new_[8459]_ , \new_[8460]_ ,
    \new_[8461]_ , \new_[8464]_ , \new_[8468]_ , \new_[8469]_ ,
    \new_[8470]_ , \new_[8474]_ , \new_[8475]_ , \new_[8479]_ ,
    \new_[8480]_ , \new_[8481]_ , \new_[8484]_ , \new_[8488]_ ,
    \new_[8489]_ , \new_[8490]_ , \new_[8494]_ , \new_[8495]_ ,
    \new_[8499]_ , \new_[8500]_ , \new_[8501]_ , \new_[8504]_ ,
    \new_[8508]_ , \new_[8509]_ , \new_[8510]_ , \new_[8514]_ ,
    \new_[8515]_ , \new_[8519]_ , \new_[8520]_ , \new_[8521]_ ,
    \new_[8524]_ , \new_[8528]_ , \new_[8529]_ , \new_[8530]_ ,
    \new_[8534]_ , \new_[8535]_ , \new_[8539]_ , \new_[8540]_ ,
    \new_[8541]_ , \new_[8544]_ , \new_[8548]_ , \new_[8549]_ ,
    \new_[8550]_ , \new_[8554]_ , \new_[8555]_ , \new_[8559]_ ,
    \new_[8560]_ , \new_[8561]_ , \new_[8564]_ , \new_[8568]_ ,
    \new_[8569]_ , \new_[8570]_ , \new_[8574]_ , \new_[8575]_ ,
    \new_[8579]_ , \new_[8580]_ , \new_[8581]_ , \new_[8584]_ ,
    \new_[8588]_ , \new_[8589]_ , \new_[8590]_ , \new_[8594]_ ,
    \new_[8595]_ , \new_[8599]_ , \new_[8600]_ , \new_[8601]_ ,
    \new_[8604]_ , \new_[8608]_ , \new_[8609]_ , \new_[8610]_ ,
    \new_[8614]_ , \new_[8615]_ , \new_[8619]_ , \new_[8620]_ ,
    \new_[8621]_ , \new_[8624]_ , \new_[8628]_ , \new_[8629]_ ,
    \new_[8630]_ , \new_[8634]_ , \new_[8635]_ , \new_[8639]_ ,
    \new_[8640]_ , \new_[8641]_ , \new_[8644]_ , \new_[8648]_ ,
    \new_[8649]_ , \new_[8650]_ , \new_[8654]_ , \new_[8655]_ ,
    \new_[8659]_ , \new_[8660]_ , \new_[8661]_ , \new_[8664]_ ,
    \new_[8668]_ , \new_[8669]_ , \new_[8670]_ , \new_[8674]_ ,
    \new_[8675]_ , \new_[8679]_ , \new_[8680]_ , \new_[8681]_ ,
    \new_[8684]_ , \new_[8688]_ , \new_[8689]_ , \new_[8690]_ ,
    \new_[8694]_ , \new_[8695]_ , \new_[8699]_ , \new_[8700]_ ,
    \new_[8701]_ , \new_[8704]_ , \new_[8708]_ , \new_[8709]_ ,
    \new_[8710]_ , \new_[8714]_ , \new_[8715]_ , \new_[8719]_ ,
    \new_[8720]_ , \new_[8721]_ , \new_[8724]_ , \new_[8728]_ ,
    \new_[8729]_ , \new_[8730]_ , \new_[8734]_ , \new_[8735]_ ,
    \new_[8739]_ , \new_[8740]_ , \new_[8741]_ , \new_[8744]_ ,
    \new_[8748]_ , \new_[8749]_ , \new_[8750]_ , \new_[8754]_ ,
    \new_[8755]_ , \new_[8759]_ , \new_[8760]_ , \new_[8761]_ ,
    \new_[8764]_ , \new_[8768]_ , \new_[8769]_ , \new_[8770]_ ,
    \new_[8774]_ , \new_[8775]_ , \new_[8779]_ , \new_[8780]_ ,
    \new_[8781]_ , \new_[8784]_ , \new_[8788]_ , \new_[8789]_ ,
    \new_[8790]_ , \new_[8794]_ , \new_[8795]_ , \new_[8799]_ ,
    \new_[8800]_ , \new_[8801]_ , \new_[8804]_ , \new_[8808]_ ,
    \new_[8809]_ , \new_[8810]_ , \new_[8814]_ , \new_[8815]_ ,
    \new_[8819]_ , \new_[8820]_ , \new_[8821]_ , \new_[8824]_ ,
    \new_[8828]_ , \new_[8829]_ , \new_[8830]_ , \new_[8834]_ ,
    \new_[8835]_ , \new_[8839]_ , \new_[8840]_ , \new_[8841]_ ,
    \new_[8844]_ , \new_[8848]_ , \new_[8849]_ , \new_[8850]_ ,
    \new_[8854]_ , \new_[8855]_ , \new_[8859]_ , \new_[8860]_ ,
    \new_[8861]_ , \new_[8864]_ , \new_[8868]_ , \new_[8869]_ ,
    \new_[8870]_ , \new_[8874]_ , \new_[8875]_ , \new_[8879]_ ,
    \new_[8880]_ , \new_[8881]_ , \new_[8884]_ , \new_[8888]_ ,
    \new_[8889]_ , \new_[8890]_ , \new_[8894]_ , \new_[8895]_ ,
    \new_[8899]_ , \new_[8900]_ , \new_[8901]_ , \new_[8904]_ ,
    \new_[8908]_ , \new_[8909]_ , \new_[8910]_ , \new_[8914]_ ,
    \new_[8915]_ , \new_[8919]_ , \new_[8920]_ , \new_[8921]_ ,
    \new_[8924]_ , \new_[8928]_ , \new_[8929]_ , \new_[8930]_ ,
    \new_[8934]_ , \new_[8935]_ , \new_[8939]_ , \new_[8940]_ ,
    \new_[8941]_ , \new_[8944]_ , \new_[8948]_ , \new_[8949]_ ,
    \new_[8950]_ , \new_[8954]_ , \new_[8955]_ , \new_[8959]_ ,
    \new_[8960]_ , \new_[8961]_ , \new_[8964]_ , \new_[8968]_ ,
    \new_[8969]_ , \new_[8970]_ , \new_[8974]_ , \new_[8975]_ ,
    \new_[8979]_ , \new_[8980]_ , \new_[8981]_ , \new_[8984]_ ,
    \new_[8988]_ , \new_[8989]_ , \new_[8990]_ , \new_[8994]_ ,
    \new_[8995]_ , \new_[8999]_ , \new_[9000]_ , \new_[9001]_ ,
    \new_[9004]_ , \new_[9008]_ , \new_[9009]_ , \new_[9010]_ ,
    \new_[9014]_ , \new_[9015]_ , \new_[9019]_ , \new_[9020]_ ,
    \new_[9021]_ , \new_[9024]_ , \new_[9028]_ , \new_[9029]_ ,
    \new_[9030]_ , \new_[9034]_ , \new_[9035]_ , \new_[9039]_ ,
    \new_[9040]_ , \new_[9041]_ , \new_[9044]_ , \new_[9048]_ ,
    \new_[9049]_ , \new_[9050]_ , \new_[9054]_ , \new_[9055]_ ,
    \new_[9059]_ , \new_[9060]_ , \new_[9061]_ , \new_[9064]_ ,
    \new_[9068]_ , \new_[9069]_ , \new_[9070]_ , \new_[9074]_ ,
    \new_[9075]_ , \new_[9079]_ , \new_[9080]_ , \new_[9081]_ ,
    \new_[9084]_ , \new_[9088]_ , \new_[9089]_ , \new_[9090]_ ,
    \new_[9094]_ , \new_[9095]_ , \new_[9099]_ , \new_[9100]_ ,
    \new_[9101]_ , \new_[9104]_ , \new_[9108]_ , \new_[9109]_ ,
    \new_[9110]_ , \new_[9114]_ , \new_[9115]_ , \new_[9119]_ ,
    \new_[9120]_ , \new_[9121]_ , \new_[9124]_ , \new_[9128]_ ,
    \new_[9129]_ , \new_[9130]_ , \new_[9134]_ , \new_[9135]_ ,
    \new_[9139]_ , \new_[9140]_ , \new_[9141]_ , \new_[9144]_ ,
    \new_[9148]_ , \new_[9149]_ , \new_[9150]_ , \new_[9154]_ ,
    \new_[9155]_ , \new_[9159]_ , \new_[9160]_ , \new_[9161]_ ,
    \new_[9164]_ , \new_[9168]_ , \new_[9169]_ , \new_[9170]_ ,
    \new_[9174]_ , \new_[9175]_ , \new_[9179]_ , \new_[9180]_ ,
    \new_[9181]_ , \new_[9184]_ , \new_[9188]_ , \new_[9189]_ ,
    \new_[9190]_ , \new_[9194]_ , \new_[9195]_ , \new_[9199]_ ,
    \new_[9200]_ , \new_[9201]_ , \new_[9204]_ , \new_[9208]_ ,
    \new_[9209]_ , \new_[9210]_ , \new_[9214]_ , \new_[9215]_ ,
    \new_[9219]_ , \new_[9220]_ , \new_[9221]_ , \new_[9224]_ ,
    \new_[9228]_ , \new_[9229]_ , \new_[9230]_ , \new_[9234]_ ,
    \new_[9235]_ , \new_[9239]_ , \new_[9240]_ , \new_[9241]_ ,
    \new_[9244]_ , \new_[9248]_ , \new_[9249]_ , \new_[9250]_ ,
    \new_[9254]_ , \new_[9255]_ , \new_[9259]_ , \new_[9260]_ ,
    \new_[9261]_ , \new_[9264]_ , \new_[9268]_ , \new_[9269]_ ,
    \new_[9270]_ , \new_[9274]_ , \new_[9275]_ , \new_[9279]_ ,
    \new_[9280]_ , \new_[9281]_ , \new_[9284]_ , \new_[9288]_ ,
    \new_[9289]_ , \new_[9290]_ , \new_[9294]_ , \new_[9295]_ ,
    \new_[9299]_ , \new_[9300]_ , \new_[9301]_ , \new_[9304]_ ,
    \new_[9308]_ , \new_[9309]_ , \new_[9310]_ , \new_[9314]_ ,
    \new_[9315]_ , \new_[9319]_ , \new_[9320]_ , \new_[9321]_ ,
    \new_[9324]_ , \new_[9328]_ , \new_[9329]_ , \new_[9330]_ ,
    \new_[9334]_ , \new_[9335]_ , \new_[9339]_ , \new_[9340]_ ,
    \new_[9341]_ , \new_[9344]_ , \new_[9348]_ , \new_[9349]_ ,
    \new_[9350]_ , \new_[9354]_ , \new_[9355]_ , \new_[9359]_ ,
    \new_[9360]_ , \new_[9361]_ , \new_[9364]_ , \new_[9368]_ ,
    \new_[9369]_ , \new_[9370]_ , \new_[9374]_ , \new_[9375]_ ,
    \new_[9379]_ , \new_[9380]_ , \new_[9381]_ , \new_[9384]_ ,
    \new_[9388]_ , \new_[9389]_ , \new_[9390]_ , \new_[9394]_ ,
    \new_[9395]_ , \new_[9399]_ , \new_[9400]_ , \new_[9401]_ ,
    \new_[9404]_ , \new_[9408]_ , \new_[9409]_ , \new_[9410]_ ,
    \new_[9414]_ , \new_[9415]_ , \new_[9419]_ , \new_[9420]_ ,
    \new_[9421]_ , \new_[9424]_ , \new_[9428]_ , \new_[9429]_ ,
    \new_[9430]_ , \new_[9434]_ , \new_[9435]_ , \new_[9439]_ ,
    \new_[9440]_ , \new_[9441]_ , \new_[9444]_ , \new_[9448]_ ,
    \new_[9449]_ , \new_[9450]_ , \new_[9454]_ , \new_[9455]_ ,
    \new_[9459]_ , \new_[9460]_ , \new_[9461]_ , \new_[9464]_ ,
    \new_[9468]_ , \new_[9469]_ , \new_[9470]_ , \new_[9474]_ ,
    \new_[9475]_ , \new_[9479]_ , \new_[9480]_ , \new_[9481]_ ,
    \new_[9484]_ , \new_[9488]_ , \new_[9489]_ , \new_[9490]_ ,
    \new_[9494]_ , \new_[9495]_ , \new_[9499]_ , \new_[9500]_ ,
    \new_[9501]_ , \new_[9504]_ , \new_[9508]_ , \new_[9509]_ ,
    \new_[9510]_ , \new_[9514]_ , \new_[9515]_ , \new_[9519]_ ,
    \new_[9520]_ , \new_[9521]_ , \new_[9524]_ , \new_[9528]_ ,
    \new_[9529]_ , \new_[9530]_ , \new_[9534]_ , \new_[9535]_ ,
    \new_[9539]_ , \new_[9540]_ , \new_[9541]_ , \new_[9544]_ ,
    \new_[9548]_ , \new_[9549]_ , \new_[9550]_ , \new_[9554]_ ,
    \new_[9555]_ , \new_[9559]_ , \new_[9560]_ , \new_[9561]_ ,
    \new_[9564]_ , \new_[9568]_ , \new_[9569]_ , \new_[9570]_ ,
    \new_[9574]_ , \new_[9575]_ , \new_[9579]_ , \new_[9580]_ ,
    \new_[9581]_ , \new_[9584]_ , \new_[9588]_ , \new_[9589]_ ,
    \new_[9590]_ , \new_[9594]_ , \new_[9595]_ , \new_[9599]_ ,
    \new_[9600]_ , \new_[9601]_ , \new_[9604]_ , \new_[9608]_ ,
    \new_[9609]_ , \new_[9610]_ , \new_[9614]_ , \new_[9615]_ ,
    \new_[9619]_ , \new_[9620]_ , \new_[9621]_ , \new_[9624]_ ,
    \new_[9628]_ , \new_[9629]_ , \new_[9630]_ , \new_[9634]_ ,
    \new_[9635]_ , \new_[9639]_ , \new_[9640]_ , \new_[9641]_ ,
    \new_[9644]_ , \new_[9648]_ , \new_[9649]_ , \new_[9650]_ ,
    \new_[9654]_ , \new_[9655]_ , \new_[9659]_ , \new_[9660]_ ,
    \new_[9661]_ , \new_[9664]_ , \new_[9668]_ , \new_[9669]_ ,
    \new_[9670]_ , \new_[9674]_ , \new_[9675]_ , \new_[9679]_ ,
    \new_[9680]_ , \new_[9681]_ , \new_[9684]_ , \new_[9688]_ ,
    \new_[9689]_ , \new_[9690]_ , \new_[9694]_ , \new_[9695]_ ,
    \new_[9699]_ , \new_[9700]_ , \new_[9701]_ , \new_[9704]_ ,
    \new_[9708]_ , \new_[9709]_ , \new_[9710]_ , \new_[9714]_ ,
    \new_[9715]_ , \new_[9719]_ , \new_[9720]_ , \new_[9721]_ ,
    \new_[9724]_ , \new_[9728]_ , \new_[9729]_ , \new_[9730]_ ,
    \new_[9734]_ , \new_[9735]_ , \new_[9739]_ , \new_[9740]_ ,
    \new_[9741]_ , \new_[9744]_ , \new_[9748]_ , \new_[9749]_ ,
    \new_[9750]_ , \new_[9754]_ , \new_[9755]_ , \new_[9759]_ ,
    \new_[9760]_ , \new_[9761]_ , \new_[9764]_ , \new_[9768]_ ,
    \new_[9769]_ , \new_[9770]_ , \new_[9774]_ , \new_[9775]_ ,
    \new_[9779]_ , \new_[9780]_ , \new_[9781]_ , \new_[9784]_ ,
    \new_[9788]_ , \new_[9789]_ , \new_[9790]_ , \new_[9794]_ ,
    \new_[9795]_ , \new_[9799]_ , \new_[9800]_ , \new_[9801]_ ,
    \new_[9804]_ , \new_[9808]_ , \new_[9809]_ , \new_[9810]_ ,
    \new_[9814]_ , \new_[9815]_ , \new_[9819]_ , \new_[9820]_ ,
    \new_[9821]_ , \new_[9824]_ , \new_[9828]_ , \new_[9829]_ ,
    \new_[9830]_ , \new_[9834]_ , \new_[9835]_ , \new_[9839]_ ,
    \new_[9840]_ , \new_[9841]_ , \new_[9844]_ , \new_[9848]_ ,
    \new_[9849]_ , \new_[9850]_ , \new_[9854]_ , \new_[9855]_ ,
    \new_[9859]_ , \new_[9860]_ , \new_[9861]_ , \new_[9864]_ ,
    \new_[9868]_ , \new_[9869]_ , \new_[9870]_ , \new_[9874]_ ,
    \new_[9875]_ , \new_[9879]_ , \new_[9880]_ , \new_[9881]_ ,
    \new_[9884]_ , \new_[9888]_ , \new_[9889]_ , \new_[9890]_ ,
    \new_[9894]_ , \new_[9895]_ , \new_[9899]_ , \new_[9900]_ ,
    \new_[9901]_ , \new_[9904]_ , \new_[9908]_ , \new_[9909]_ ,
    \new_[9910]_ , \new_[9914]_ , \new_[9915]_ , \new_[9919]_ ,
    \new_[9920]_ , \new_[9921]_ , \new_[9924]_ , \new_[9928]_ ,
    \new_[9929]_ , \new_[9930]_ , \new_[9934]_ , \new_[9935]_ ,
    \new_[9939]_ , \new_[9940]_ , \new_[9941]_ , \new_[9944]_ ,
    \new_[9948]_ , \new_[9949]_ , \new_[9950]_ , \new_[9954]_ ,
    \new_[9955]_ , \new_[9959]_ , \new_[9960]_ , \new_[9961]_ ,
    \new_[9964]_ , \new_[9968]_ , \new_[9969]_ , \new_[9970]_ ,
    \new_[9974]_ , \new_[9975]_ , \new_[9979]_ , \new_[9980]_ ,
    \new_[9981]_ , \new_[9984]_ , \new_[9988]_ , \new_[9989]_ ,
    \new_[9990]_ , \new_[9994]_ , \new_[9995]_ , \new_[9999]_ ,
    \new_[10000]_ , \new_[10001]_ , \new_[10004]_ , \new_[10008]_ ,
    \new_[10009]_ , \new_[10010]_ , \new_[10014]_ , \new_[10015]_ ,
    \new_[10019]_ , \new_[10020]_ , \new_[10021]_ , \new_[10024]_ ,
    \new_[10028]_ , \new_[10029]_ , \new_[10030]_ , \new_[10034]_ ,
    \new_[10035]_ , \new_[10039]_ , \new_[10040]_ , \new_[10041]_ ,
    \new_[10044]_ , \new_[10048]_ , \new_[10049]_ , \new_[10050]_ ,
    \new_[10054]_ , \new_[10055]_ , \new_[10059]_ , \new_[10060]_ ,
    \new_[10061]_ , \new_[10064]_ , \new_[10068]_ , \new_[10069]_ ,
    \new_[10070]_ , \new_[10074]_ , \new_[10075]_ , \new_[10079]_ ,
    \new_[10080]_ , \new_[10081]_ , \new_[10084]_ , \new_[10088]_ ,
    \new_[10089]_ , \new_[10090]_ , \new_[10094]_ , \new_[10095]_ ,
    \new_[10099]_ , \new_[10100]_ , \new_[10101]_ , \new_[10104]_ ,
    \new_[10108]_ , \new_[10109]_ , \new_[10110]_ , \new_[10114]_ ,
    \new_[10115]_ , \new_[10119]_ , \new_[10120]_ , \new_[10121]_ ,
    \new_[10124]_ , \new_[10128]_ , \new_[10129]_ , \new_[10130]_ ,
    \new_[10134]_ , \new_[10135]_ , \new_[10139]_ , \new_[10140]_ ,
    \new_[10141]_ , \new_[10144]_ , \new_[10148]_ , \new_[10149]_ ,
    \new_[10150]_ , \new_[10154]_ , \new_[10155]_ , \new_[10159]_ ,
    \new_[10160]_ , \new_[10161]_ , \new_[10164]_ , \new_[10168]_ ,
    \new_[10169]_ , \new_[10170]_ , \new_[10174]_ , \new_[10175]_ ,
    \new_[10179]_ , \new_[10180]_ , \new_[10181]_ , \new_[10184]_ ,
    \new_[10188]_ , \new_[10189]_ , \new_[10190]_ , \new_[10194]_ ,
    \new_[10195]_ , \new_[10199]_ , \new_[10200]_ , \new_[10201]_ ,
    \new_[10204]_ , \new_[10208]_ , \new_[10209]_ , \new_[10210]_ ,
    \new_[10214]_ , \new_[10215]_ , \new_[10219]_ , \new_[10220]_ ,
    \new_[10221]_ , \new_[10224]_ , \new_[10228]_ , \new_[10229]_ ,
    \new_[10230]_ , \new_[10234]_ , \new_[10235]_ , \new_[10239]_ ,
    \new_[10240]_ , \new_[10241]_ , \new_[10244]_ , \new_[10248]_ ,
    \new_[10249]_ , \new_[10250]_ , \new_[10254]_ , \new_[10255]_ ,
    \new_[10259]_ , \new_[10260]_ , \new_[10261]_ , \new_[10264]_ ,
    \new_[10268]_ , \new_[10269]_ , \new_[10270]_ , \new_[10274]_ ,
    \new_[10275]_ , \new_[10279]_ , \new_[10280]_ , \new_[10281]_ ,
    \new_[10284]_ , \new_[10288]_ , \new_[10289]_ , \new_[10290]_ ,
    \new_[10294]_ , \new_[10295]_ , \new_[10299]_ , \new_[10300]_ ,
    \new_[10301]_ , \new_[10304]_ , \new_[10308]_ , \new_[10309]_ ,
    \new_[10310]_ , \new_[10314]_ , \new_[10315]_ , \new_[10319]_ ,
    \new_[10320]_ , \new_[10321]_ , \new_[10324]_ , \new_[10328]_ ,
    \new_[10329]_ , \new_[10330]_ , \new_[10334]_ , \new_[10335]_ ,
    \new_[10339]_ , \new_[10340]_ , \new_[10341]_ , \new_[10344]_ ,
    \new_[10348]_ , \new_[10349]_ , \new_[10350]_ , \new_[10354]_ ,
    \new_[10355]_ , \new_[10359]_ , \new_[10360]_ , \new_[10361]_ ,
    \new_[10364]_ , \new_[10368]_ , \new_[10369]_ , \new_[10370]_ ,
    \new_[10374]_ , \new_[10375]_ , \new_[10379]_ , \new_[10380]_ ,
    \new_[10381]_ , \new_[10384]_ , \new_[10388]_ , \new_[10389]_ ,
    \new_[10390]_ , \new_[10394]_ , \new_[10395]_ , \new_[10399]_ ,
    \new_[10400]_ , \new_[10401]_ , \new_[10404]_ , \new_[10408]_ ,
    \new_[10409]_ , \new_[10410]_ , \new_[10414]_ , \new_[10415]_ ,
    \new_[10419]_ , \new_[10420]_ , \new_[10421]_ , \new_[10424]_ ,
    \new_[10428]_ , \new_[10429]_ , \new_[10430]_ , \new_[10434]_ ,
    \new_[10435]_ , \new_[10439]_ , \new_[10440]_ , \new_[10441]_ ,
    \new_[10444]_ , \new_[10448]_ , \new_[10449]_ , \new_[10450]_ ,
    \new_[10454]_ , \new_[10455]_ , \new_[10459]_ , \new_[10460]_ ,
    \new_[10461]_ , \new_[10464]_ , \new_[10468]_ , \new_[10469]_ ,
    \new_[10470]_ , \new_[10474]_ , \new_[10475]_ , \new_[10479]_ ,
    \new_[10480]_ , \new_[10481]_ , \new_[10484]_ , \new_[10488]_ ,
    \new_[10489]_ , \new_[10490]_ , \new_[10494]_ , \new_[10495]_ ,
    \new_[10499]_ , \new_[10500]_ , \new_[10501]_ , \new_[10504]_ ,
    \new_[10508]_ , \new_[10509]_ , \new_[10510]_ , \new_[10514]_ ,
    \new_[10515]_ , \new_[10519]_ , \new_[10520]_ , \new_[10521]_ ,
    \new_[10524]_ , \new_[10528]_ , \new_[10529]_ , \new_[10530]_ ,
    \new_[10534]_ , \new_[10535]_ , \new_[10539]_ , \new_[10540]_ ,
    \new_[10541]_ , \new_[10544]_ , \new_[10548]_ , \new_[10549]_ ,
    \new_[10550]_ , \new_[10554]_ , \new_[10555]_ , \new_[10559]_ ,
    \new_[10560]_ , \new_[10561]_ , \new_[10564]_ , \new_[10568]_ ,
    \new_[10569]_ , \new_[10570]_ , \new_[10574]_ , \new_[10575]_ ,
    \new_[10579]_ , \new_[10580]_ , \new_[10581]_ , \new_[10584]_ ,
    \new_[10588]_ , \new_[10589]_ , \new_[10590]_ , \new_[10594]_ ,
    \new_[10595]_ , \new_[10599]_ , \new_[10600]_ , \new_[10601]_ ,
    \new_[10604]_ , \new_[10608]_ , \new_[10609]_ , \new_[10610]_ ,
    \new_[10614]_ , \new_[10615]_ , \new_[10619]_ , \new_[10620]_ ,
    \new_[10621]_ , \new_[10624]_ , \new_[10628]_ , \new_[10629]_ ,
    \new_[10630]_ , \new_[10634]_ , \new_[10635]_ , \new_[10639]_ ,
    \new_[10640]_ , \new_[10641]_ , \new_[10644]_ , \new_[10648]_ ,
    \new_[10649]_ , \new_[10650]_ , \new_[10654]_ , \new_[10655]_ ,
    \new_[10659]_ , \new_[10660]_ , \new_[10661]_ , \new_[10664]_ ,
    \new_[10668]_ , \new_[10669]_ , \new_[10670]_ , \new_[10674]_ ,
    \new_[10675]_ , \new_[10679]_ , \new_[10680]_ , \new_[10681]_ ,
    \new_[10684]_ , \new_[10688]_ , \new_[10689]_ , \new_[10690]_ ,
    \new_[10694]_ , \new_[10695]_ , \new_[10699]_ , \new_[10700]_ ,
    \new_[10701]_ , \new_[10704]_ , \new_[10708]_ , \new_[10709]_ ,
    \new_[10710]_ , \new_[10714]_ , \new_[10715]_ , \new_[10719]_ ,
    \new_[10720]_ , \new_[10721]_ , \new_[10724]_ , \new_[10728]_ ,
    \new_[10729]_ , \new_[10730]_ , \new_[10734]_ , \new_[10735]_ ,
    \new_[10739]_ , \new_[10740]_ , \new_[10741]_ , \new_[10744]_ ,
    \new_[10748]_ , \new_[10749]_ , \new_[10750]_ , \new_[10754]_ ,
    \new_[10755]_ , \new_[10759]_ , \new_[10760]_ , \new_[10761]_ ,
    \new_[10764]_ , \new_[10768]_ , \new_[10769]_ , \new_[10770]_ ,
    \new_[10774]_ , \new_[10775]_ , \new_[10779]_ , \new_[10780]_ ,
    \new_[10781]_ , \new_[10784]_ , \new_[10788]_ , \new_[10789]_ ,
    \new_[10790]_ , \new_[10794]_ , \new_[10795]_ , \new_[10799]_ ,
    \new_[10800]_ , \new_[10801]_ , \new_[10804]_ , \new_[10808]_ ,
    \new_[10809]_ , \new_[10810]_ , \new_[10814]_ , \new_[10815]_ ,
    \new_[10819]_ , \new_[10820]_ , \new_[10821]_ , \new_[10824]_ ,
    \new_[10828]_ , \new_[10829]_ , \new_[10830]_ , \new_[10834]_ ,
    \new_[10835]_ , \new_[10839]_ , \new_[10840]_ , \new_[10841]_ ,
    \new_[10844]_ , \new_[10848]_ , \new_[10849]_ , \new_[10850]_ ,
    \new_[10854]_ , \new_[10855]_ , \new_[10859]_ , \new_[10860]_ ,
    \new_[10861]_ , \new_[10864]_ , \new_[10868]_ , \new_[10869]_ ,
    \new_[10870]_ , \new_[10874]_ , \new_[10875]_ , \new_[10879]_ ,
    \new_[10880]_ , \new_[10881]_ , \new_[10884]_ , \new_[10888]_ ,
    \new_[10889]_ , \new_[10890]_ , \new_[10894]_ , \new_[10895]_ ,
    \new_[10899]_ , \new_[10900]_ , \new_[10901]_ , \new_[10904]_ ,
    \new_[10908]_ , \new_[10909]_ , \new_[10910]_ , \new_[10914]_ ,
    \new_[10915]_ , \new_[10919]_ , \new_[10920]_ , \new_[10921]_ ,
    \new_[10924]_ , \new_[10928]_ , \new_[10929]_ , \new_[10930]_ ,
    \new_[10934]_ , \new_[10935]_ , \new_[10939]_ , \new_[10940]_ ,
    \new_[10941]_ , \new_[10944]_ , \new_[10948]_ , \new_[10949]_ ,
    \new_[10950]_ , \new_[10954]_ , \new_[10955]_ , \new_[10959]_ ,
    \new_[10960]_ , \new_[10961]_ , \new_[10964]_ , \new_[10968]_ ,
    \new_[10969]_ , \new_[10970]_ , \new_[10974]_ , \new_[10975]_ ,
    \new_[10979]_ , \new_[10980]_ , \new_[10981]_ , \new_[10984]_ ,
    \new_[10988]_ , \new_[10989]_ , \new_[10990]_ , \new_[10994]_ ,
    \new_[10995]_ , \new_[10999]_ , \new_[11000]_ , \new_[11001]_ ,
    \new_[11004]_ , \new_[11008]_ , \new_[11009]_ , \new_[11010]_ ,
    \new_[11014]_ , \new_[11015]_ , \new_[11019]_ , \new_[11020]_ ,
    \new_[11021]_ , \new_[11024]_ , \new_[11028]_ , \new_[11029]_ ,
    \new_[11030]_ , \new_[11034]_ , \new_[11035]_ , \new_[11039]_ ,
    \new_[11040]_ , \new_[11041]_ , \new_[11044]_ , \new_[11048]_ ,
    \new_[11049]_ , \new_[11050]_ , \new_[11054]_ , \new_[11055]_ ,
    \new_[11059]_ , \new_[11060]_ , \new_[11061]_ , \new_[11064]_ ,
    \new_[11068]_ , \new_[11069]_ , \new_[11070]_ , \new_[11074]_ ,
    \new_[11075]_ , \new_[11079]_ , \new_[11080]_ , \new_[11081]_ ,
    \new_[11084]_ , \new_[11088]_ , \new_[11089]_ , \new_[11090]_ ,
    \new_[11094]_ , \new_[11095]_ , \new_[11099]_ , \new_[11100]_ ,
    \new_[11101]_ , \new_[11104]_ , \new_[11108]_ , \new_[11109]_ ,
    \new_[11110]_ , \new_[11114]_ , \new_[11115]_ , \new_[11119]_ ,
    \new_[11120]_ , \new_[11121]_ , \new_[11124]_ , \new_[11128]_ ,
    \new_[11129]_ , \new_[11130]_ , \new_[11134]_ , \new_[11135]_ ,
    \new_[11139]_ , \new_[11140]_ , \new_[11141]_ , \new_[11144]_ ,
    \new_[11148]_ , \new_[11149]_ , \new_[11150]_ , \new_[11154]_ ,
    \new_[11155]_ , \new_[11159]_ , \new_[11160]_ , \new_[11161]_ ,
    \new_[11164]_ , \new_[11168]_ , \new_[11169]_ , \new_[11170]_ ,
    \new_[11174]_ , \new_[11175]_ , \new_[11179]_ , \new_[11180]_ ,
    \new_[11181]_ , \new_[11184]_ , \new_[11188]_ , \new_[11189]_ ,
    \new_[11190]_ , \new_[11194]_ , \new_[11195]_ , \new_[11199]_ ,
    \new_[11200]_ , \new_[11201]_ , \new_[11204]_ , \new_[11208]_ ,
    \new_[11209]_ , \new_[11210]_ , \new_[11214]_ , \new_[11215]_ ,
    \new_[11219]_ , \new_[11220]_ , \new_[11221]_ , \new_[11224]_ ,
    \new_[11228]_ , \new_[11229]_ , \new_[11230]_ , \new_[11234]_ ,
    \new_[11235]_ , \new_[11239]_ , \new_[11240]_ , \new_[11241]_ ,
    \new_[11244]_ , \new_[11248]_ , \new_[11249]_ , \new_[11250]_ ,
    \new_[11254]_ , \new_[11255]_ , \new_[11259]_ , \new_[11260]_ ,
    \new_[11261]_ , \new_[11264]_ , \new_[11268]_ , \new_[11269]_ ,
    \new_[11270]_ , \new_[11274]_ , \new_[11275]_ , \new_[11279]_ ,
    \new_[11280]_ , \new_[11281]_ , \new_[11284]_ , \new_[11288]_ ,
    \new_[11289]_ , \new_[11290]_ , \new_[11294]_ , \new_[11295]_ ,
    \new_[11299]_ , \new_[11300]_ , \new_[11301]_ , \new_[11304]_ ,
    \new_[11308]_ , \new_[11309]_ , \new_[11310]_ , \new_[11314]_ ,
    \new_[11315]_ , \new_[11319]_ , \new_[11320]_ , \new_[11321]_ ,
    \new_[11324]_ , \new_[11328]_ , \new_[11329]_ , \new_[11330]_ ,
    \new_[11334]_ , \new_[11335]_ , \new_[11339]_ , \new_[11340]_ ,
    \new_[11341]_ , \new_[11344]_ , \new_[11348]_ , \new_[11349]_ ,
    \new_[11350]_ , \new_[11354]_ , \new_[11355]_ , \new_[11359]_ ,
    \new_[11360]_ , \new_[11361]_ , \new_[11364]_ , \new_[11368]_ ,
    \new_[11369]_ , \new_[11370]_ , \new_[11374]_ , \new_[11375]_ ,
    \new_[11379]_ , \new_[11380]_ , \new_[11381]_ , \new_[11384]_ ,
    \new_[11388]_ , \new_[11389]_ , \new_[11390]_ , \new_[11394]_ ,
    \new_[11395]_ , \new_[11399]_ , \new_[11400]_ , \new_[11401]_ ,
    \new_[11404]_ , \new_[11408]_ , \new_[11409]_ , \new_[11410]_ ,
    \new_[11414]_ , \new_[11415]_ , \new_[11419]_ , \new_[11420]_ ,
    \new_[11421]_ , \new_[11424]_ , \new_[11428]_ , \new_[11429]_ ,
    \new_[11430]_ , \new_[11434]_ , \new_[11435]_ , \new_[11439]_ ,
    \new_[11440]_ , \new_[11441]_ , \new_[11444]_ , \new_[11448]_ ,
    \new_[11449]_ , \new_[11450]_ , \new_[11454]_ , \new_[11455]_ ,
    \new_[11459]_ , \new_[11460]_ , \new_[11461]_ , \new_[11464]_ ,
    \new_[11468]_ , \new_[11469]_ , \new_[11470]_ , \new_[11474]_ ,
    \new_[11475]_ , \new_[11479]_ , \new_[11480]_ , \new_[11481]_ ,
    \new_[11484]_ , \new_[11488]_ , \new_[11489]_ , \new_[11490]_ ,
    \new_[11494]_ , \new_[11495]_ , \new_[11499]_ , \new_[11500]_ ,
    \new_[11501]_ , \new_[11504]_ , \new_[11508]_ , \new_[11509]_ ,
    \new_[11510]_ , \new_[11514]_ , \new_[11515]_ , \new_[11519]_ ,
    \new_[11520]_ , \new_[11521]_ , \new_[11524]_ , \new_[11528]_ ,
    \new_[11529]_ , \new_[11530]_ , \new_[11534]_ , \new_[11535]_ ,
    \new_[11539]_ , \new_[11540]_ , \new_[11541]_ , \new_[11544]_ ,
    \new_[11548]_ , \new_[11549]_ , \new_[11550]_ , \new_[11554]_ ,
    \new_[11555]_ , \new_[11559]_ , \new_[11560]_ , \new_[11561]_ ,
    \new_[11564]_ , \new_[11568]_ , \new_[11569]_ , \new_[11570]_ ,
    \new_[11574]_ , \new_[11575]_ , \new_[11579]_ , \new_[11580]_ ,
    \new_[11581]_ , \new_[11584]_ , \new_[11588]_ , \new_[11589]_ ,
    \new_[11590]_ , \new_[11594]_ , \new_[11595]_ , \new_[11599]_ ,
    \new_[11600]_ , \new_[11601]_ , \new_[11604]_ , \new_[11608]_ ,
    \new_[11609]_ , \new_[11610]_ , \new_[11614]_ , \new_[11615]_ ,
    \new_[11619]_ , \new_[11620]_ , \new_[11621]_ , \new_[11624]_ ,
    \new_[11628]_ , \new_[11629]_ , \new_[11630]_ , \new_[11634]_ ,
    \new_[11635]_ , \new_[11639]_ , \new_[11640]_ , \new_[11641]_ ,
    \new_[11644]_ , \new_[11648]_ , \new_[11649]_ , \new_[11650]_ ,
    \new_[11654]_ , \new_[11655]_ , \new_[11659]_ , \new_[11660]_ ,
    \new_[11661]_ , \new_[11664]_ , \new_[11668]_ , \new_[11669]_ ,
    \new_[11670]_ , \new_[11674]_ , \new_[11675]_ , \new_[11679]_ ,
    \new_[11680]_ , \new_[11681]_ , \new_[11684]_ , \new_[11688]_ ,
    \new_[11689]_ , \new_[11690]_ , \new_[11694]_ , \new_[11695]_ ,
    \new_[11699]_ , \new_[11700]_ , \new_[11701]_ , \new_[11704]_ ,
    \new_[11708]_ , \new_[11709]_ , \new_[11710]_ , \new_[11714]_ ,
    \new_[11715]_ , \new_[11719]_ , \new_[11720]_ , \new_[11721]_ ,
    \new_[11724]_ , \new_[11728]_ , \new_[11729]_ , \new_[11730]_ ,
    \new_[11734]_ , \new_[11735]_ , \new_[11739]_ , \new_[11740]_ ,
    \new_[11741]_ , \new_[11744]_ , \new_[11748]_ , \new_[11749]_ ,
    \new_[11750]_ , \new_[11754]_ , \new_[11755]_ , \new_[11759]_ ,
    \new_[11760]_ , \new_[11761]_ , \new_[11764]_ , \new_[11768]_ ,
    \new_[11769]_ , \new_[11770]_ , \new_[11774]_ , \new_[11775]_ ,
    \new_[11779]_ , \new_[11780]_ , \new_[11781]_ , \new_[11784]_ ,
    \new_[11788]_ , \new_[11789]_ , \new_[11790]_ , \new_[11794]_ ,
    \new_[11795]_ , \new_[11799]_ , \new_[11800]_ , \new_[11801]_ ,
    \new_[11804]_ , \new_[11808]_ , \new_[11809]_ , \new_[11810]_ ,
    \new_[11814]_ , \new_[11815]_ , \new_[11819]_ , \new_[11820]_ ,
    \new_[11821]_ , \new_[11824]_ , \new_[11828]_ , \new_[11829]_ ,
    \new_[11830]_ , \new_[11834]_ , \new_[11835]_ , \new_[11839]_ ,
    \new_[11840]_ , \new_[11841]_ , \new_[11844]_ , \new_[11848]_ ,
    \new_[11849]_ , \new_[11850]_ , \new_[11854]_ , \new_[11855]_ ,
    \new_[11859]_ , \new_[11860]_ , \new_[11861]_ , \new_[11864]_ ,
    \new_[11868]_ , \new_[11869]_ , \new_[11870]_ , \new_[11874]_ ,
    \new_[11875]_ , \new_[11879]_ , \new_[11880]_ , \new_[11881]_ ,
    \new_[11884]_ , \new_[11888]_ , \new_[11889]_ , \new_[11890]_ ,
    \new_[11894]_ , \new_[11895]_ , \new_[11899]_ , \new_[11900]_ ,
    \new_[11901]_ , \new_[11904]_ , \new_[11908]_ , \new_[11909]_ ,
    \new_[11910]_ , \new_[11914]_ , \new_[11915]_ , \new_[11919]_ ,
    \new_[11920]_ , \new_[11921]_ , \new_[11924]_ , \new_[11928]_ ,
    \new_[11929]_ , \new_[11930]_ , \new_[11934]_ , \new_[11935]_ ,
    \new_[11939]_ , \new_[11940]_ , \new_[11941]_ , \new_[11944]_ ,
    \new_[11948]_ , \new_[11949]_ , \new_[11950]_ , \new_[11954]_ ,
    \new_[11955]_ , \new_[11959]_ , \new_[11960]_ , \new_[11961]_ ,
    \new_[11964]_ , \new_[11968]_ , \new_[11969]_ , \new_[11970]_ ,
    \new_[11974]_ , \new_[11975]_ , \new_[11979]_ , \new_[11980]_ ,
    \new_[11981]_ , \new_[11984]_ , \new_[11988]_ , \new_[11989]_ ,
    \new_[11990]_ , \new_[11994]_ , \new_[11995]_ , \new_[11999]_ ,
    \new_[12000]_ , \new_[12001]_ , \new_[12004]_ , \new_[12008]_ ,
    \new_[12009]_ , \new_[12010]_ , \new_[12014]_ , \new_[12015]_ ,
    \new_[12019]_ , \new_[12020]_ , \new_[12021]_ , \new_[12024]_ ,
    \new_[12028]_ , \new_[12029]_ , \new_[12030]_ , \new_[12034]_ ,
    \new_[12035]_ , \new_[12039]_ , \new_[12040]_ , \new_[12041]_ ,
    \new_[12044]_ , \new_[12048]_ , \new_[12049]_ , \new_[12050]_ ,
    \new_[12054]_ , \new_[12055]_ , \new_[12059]_ , \new_[12060]_ ,
    \new_[12061]_ , \new_[12064]_ , \new_[12068]_ , \new_[12069]_ ,
    \new_[12070]_ , \new_[12074]_ , \new_[12075]_ , \new_[12079]_ ,
    \new_[12080]_ , \new_[12081]_ , \new_[12084]_ , \new_[12088]_ ,
    \new_[12089]_ , \new_[12090]_ , \new_[12094]_ , \new_[12095]_ ,
    \new_[12099]_ , \new_[12100]_ , \new_[12101]_ , \new_[12104]_ ,
    \new_[12108]_ , \new_[12109]_ , \new_[12110]_ , \new_[12114]_ ,
    \new_[12115]_ , \new_[12119]_ , \new_[12120]_ , \new_[12121]_ ,
    \new_[12124]_ , \new_[12128]_ , \new_[12129]_ , \new_[12130]_ ,
    \new_[12134]_ , \new_[12135]_ , \new_[12139]_ , \new_[12140]_ ,
    \new_[12141]_ , \new_[12144]_ , \new_[12148]_ , \new_[12149]_ ,
    \new_[12150]_ , \new_[12154]_ , \new_[12155]_ , \new_[12159]_ ,
    \new_[12160]_ , \new_[12161]_ , \new_[12164]_ , \new_[12168]_ ,
    \new_[12169]_ , \new_[12170]_ , \new_[12174]_ , \new_[12175]_ ,
    \new_[12179]_ , \new_[12180]_ , \new_[12181]_ , \new_[12184]_ ,
    \new_[12188]_ , \new_[12189]_ , \new_[12190]_ , \new_[12194]_ ,
    \new_[12195]_ , \new_[12199]_ , \new_[12200]_ , \new_[12201]_ ,
    \new_[12204]_ , \new_[12208]_ , \new_[12209]_ , \new_[12210]_ ,
    \new_[12214]_ , \new_[12215]_ , \new_[12219]_ , \new_[12220]_ ,
    \new_[12221]_ , \new_[12225]_ , \new_[12226]_ , \new_[12230]_ ,
    \new_[12231]_ , \new_[12232]_ , \new_[12236]_ , \new_[12237]_ ,
    \new_[12241]_ , \new_[12242]_ , \new_[12243]_ , \new_[12247]_ ,
    \new_[12248]_ , \new_[12252]_ , \new_[12253]_ , \new_[12254]_ ,
    \new_[12258]_ , \new_[12259]_ , \new_[12263]_ , \new_[12264]_ ,
    \new_[12265]_ , \new_[12269]_ , \new_[12270]_ , \new_[12274]_ ,
    \new_[12275]_ , \new_[12276]_ , \new_[12280]_ , \new_[12281]_ ,
    \new_[12285]_ , \new_[12286]_ , \new_[12287]_ , \new_[12291]_ ,
    \new_[12292]_ , \new_[12296]_ , \new_[12297]_ , \new_[12298]_ ,
    \new_[12302]_ , \new_[12303]_ , \new_[12307]_ , \new_[12308]_ ,
    \new_[12309]_ , \new_[12313]_ , \new_[12314]_ , \new_[12318]_ ,
    \new_[12319]_ , \new_[12320]_ , \new_[12324]_ , \new_[12325]_ ,
    \new_[12329]_ , \new_[12330]_ , \new_[12331]_ , \new_[12335]_ ,
    \new_[12336]_ , \new_[12340]_ , \new_[12341]_ , \new_[12342]_ ,
    \new_[12346]_ , \new_[12347]_ , \new_[12351]_ , \new_[12352]_ ,
    \new_[12353]_ , \new_[12357]_ , \new_[12358]_ , \new_[12362]_ ,
    \new_[12363]_ , \new_[12364]_ , \new_[12368]_ , \new_[12369]_ ,
    \new_[12373]_ , \new_[12374]_ , \new_[12375]_ , \new_[12379]_ ,
    \new_[12380]_ , \new_[12384]_ , \new_[12385]_ , \new_[12386]_ ,
    \new_[12390]_ , \new_[12391]_ , \new_[12395]_ , \new_[12396]_ ,
    \new_[12397]_ , \new_[12401]_ , \new_[12402]_ , \new_[12406]_ ,
    \new_[12407]_ , \new_[12408]_ , \new_[12412]_ , \new_[12413]_ ,
    \new_[12417]_ , \new_[12418]_ , \new_[12419]_ , \new_[12423]_ ,
    \new_[12424]_ , \new_[12428]_ , \new_[12429]_ , \new_[12430]_ ,
    \new_[12434]_ , \new_[12435]_ , \new_[12439]_ , \new_[12440]_ ,
    \new_[12441]_ , \new_[12445]_ , \new_[12446]_ , \new_[12450]_ ,
    \new_[12451]_ , \new_[12452]_ , \new_[12456]_ , \new_[12457]_ ,
    \new_[12461]_ , \new_[12462]_ , \new_[12463]_ , \new_[12467]_ ,
    \new_[12468]_ , \new_[12472]_ , \new_[12473]_ , \new_[12474]_ ,
    \new_[12478]_ , \new_[12479]_ , \new_[12483]_ , \new_[12484]_ ,
    \new_[12485]_ , \new_[12489]_ , \new_[12490]_ , \new_[12494]_ ,
    \new_[12495]_ , \new_[12496]_ , \new_[12500]_ , \new_[12501]_ ,
    \new_[12505]_ , \new_[12506]_ , \new_[12507]_ , \new_[12511]_ ,
    \new_[12512]_ , \new_[12516]_ , \new_[12517]_ , \new_[12518]_ ,
    \new_[12522]_ , \new_[12523]_ , \new_[12527]_ , \new_[12528]_ ,
    \new_[12529]_ , \new_[12533]_ , \new_[12534]_ , \new_[12538]_ ,
    \new_[12539]_ , \new_[12540]_ , \new_[12544]_ , \new_[12545]_ ,
    \new_[12549]_ , \new_[12550]_ , \new_[12551]_ , \new_[12555]_ ,
    \new_[12556]_ , \new_[12560]_ , \new_[12561]_ , \new_[12562]_ ,
    \new_[12566]_ , \new_[12567]_ , \new_[12571]_ , \new_[12572]_ ,
    \new_[12573]_ , \new_[12577]_ , \new_[12578]_ , \new_[12582]_ ,
    \new_[12583]_ , \new_[12584]_ , \new_[12588]_ , \new_[12589]_ ,
    \new_[12593]_ , \new_[12594]_ , \new_[12595]_ , \new_[12599]_ ,
    \new_[12600]_ , \new_[12604]_ , \new_[12605]_ , \new_[12606]_ ,
    \new_[12610]_ , \new_[12611]_ , \new_[12615]_ , \new_[12616]_ ,
    \new_[12617]_ , \new_[12621]_ , \new_[12622]_ , \new_[12626]_ ,
    \new_[12627]_ , \new_[12628]_ , \new_[12632]_ , \new_[12633]_ ,
    \new_[12637]_ , \new_[12638]_ , \new_[12639]_ , \new_[12643]_ ,
    \new_[12644]_ , \new_[12648]_ , \new_[12649]_ , \new_[12650]_ ,
    \new_[12654]_ , \new_[12655]_ , \new_[12659]_ , \new_[12660]_ ,
    \new_[12661]_ , \new_[12665]_ , \new_[12666]_ , \new_[12670]_ ,
    \new_[12671]_ , \new_[12672]_ , \new_[12676]_ , \new_[12677]_ ,
    \new_[12681]_ , \new_[12682]_ , \new_[12683]_ , \new_[12687]_ ,
    \new_[12688]_ , \new_[12692]_ , \new_[12693]_ , \new_[12694]_ ,
    \new_[12698]_ , \new_[12699]_ , \new_[12703]_ , \new_[12704]_ ,
    \new_[12705]_ , \new_[12709]_ , \new_[12710]_ , \new_[12714]_ ,
    \new_[12715]_ , \new_[12716]_ , \new_[12720]_ , \new_[12721]_ ,
    \new_[12725]_ , \new_[12726]_ , \new_[12727]_ , \new_[12731]_ ,
    \new_[12732]_ , \new_[12736]_ , \new_[12737]_ , \new_[12738]_ ,
    \new_[12742]_ , \new_[12743]_ , \new_[12747]_ , \new_[12748]_ ,
    \new_[12749]_ , \new_[12753]_ , \new_[12754]_ , \new_[12758]_ ,
    \new_[12759]_ , \new_[12760]_ , \new_[12764]_ , \new_[12765]_ ,
    \new_[12769]_ , \new_[12770]_ , \new_[12771]_ , \new_[12775]_ ,
    \new_[12776]_ , \new_[12780]_ , \new_[12781]_ , \new_[12782]_ ,
    \new_[12786]_ , \new_[12787]_ , \new_[12791]_ , \new_[12792]_ ,
    \new_[12793]_ , \new_[12797]_ , \new_[12798]_ , \new_[12802]_ ,
    \new_[12803]_ , \new_[12804]_ , \new_[12808]_ , \new_[12809]_ ,
    \new_[12813]_ , \new_[12814]_ , \new_[12815]_ , \new_[12819]_ ,
    \new_[12820]_ , \new_[12824]_ , \new_[12825]_ , \new_[12826]_ ,
    \new_[12830]_ , \new_[12831]_ , \new_[12835]_ , \new_[12836]_ ,
    \new_[12837]_ , \new_[12841]_ , \new_[12842]_ , \new_[12846]_ ,
    \new_[12847]_ , \new_[12848]_ , \new_[12852]_ , \new_[12853]_ ,
    \new_[12857]_ , \new_[12858]_ , \new_[12859]_ , \new_[12863]_ ,
    \new_[12864]_ , \new_[12868]_ , \new_[12869]_ , \new_[12870]_ ,
    \new_[12874]_ , \new_[12875]_ , \new_[12879]_ , \new_[12880]_ ,
    \new_[12881]_ , \new_[12885]_ , \new_[12886]_ , \new_[12890]_ ,
    \new_[12891]_ , \new_[12892]_ , \new_[12896]_ , \new_[12897]_ ,
    \new_[12901]_ , \new_[12902]_ , \new_[12903]_ , \new_[12907]_ ,
    \new_[12908]_ , \new_[12912]_ , \new_[12913]_ , \new_[12914]_ ,
    \new_[12918]_ , \new_[12919]_ , \new_[12923]_ , \new_[12924]_ ,
    \new_[12925]_ , \new_[12929]_ , \new_[12930]_ , \new_[12934]_ ,
    \new_[12935]_ , \new_[12936]_ , \new_[12940]_ , \new_[12941]_ ,
    \new_[12945]_ , \new_[12946]_ , \new_[12947]_ , \new_[12951]_ ,
    \new_[12952]_ , \new_[12956]_ , \new_[12957]_ , \new_[12958]_ ,
    \new_[12962]_ , \new_[12963]_ , \new_[12967]_ , \new_[12968]_ ,
    \new_[12969]_ , \new_[12973]_ , \new_[12974]_ , \new_[12978]_ ,
    \new_[12979]_ , \new_[12980]_ , \new_[12984]_ , \new_[12985]_ ,
    \new_[12989]_ , \new_[12990]_ , \new_[12991]_ , \new_[12995]_ ,
    \new_[12996]_ , \new_[13000]_ , \new_[13001]_ , \new_[13002]_ ,
    \new_[13006]_ , \new_[13007]_ , \new_[13011]_ , \new_[13012]_ ,
    \new_[13013]_ , \new_[13017]_ , \new_[13018]_ , \new_[13022]_ ,
    \new_[13023]_ , \new_[13024]_ , \new_[13028]_ , \new_[13029]_ ,
    \new_[13033]_ , \new_[13034]_ , \new_[13035]_ , \new_[13039]_ ,
    \new_[13040]_ , \new_[13044]_ , \new_[13045]_ , \new_[13046]_ ,
    \new_[13050]_ , \new_[13051]_ , \new_[13055]_ , \new_[13056]_ ,
    \new_[13057]_ , \new_[13061]_ , \new_[13062]_ , \new_[13066]_ ,
    \new_[13067]_ , \new_[13068]_ , \new_[13072]_ , \new_[13073]_ ,
    \new_[13077]_ , \new_[13078]_ , \new_[13079]_ , \new_[13083]_ ,
    \new_[13084]_ , \new_[13088]_ , \new_[13089]_ , \new_[13090]_ ,
    \new_[13094]_ , \new_[13095]_ , \new_[13099]_ , \new_[13100]_ ,
    \new_[13101]_ , \new_[13105]_ , \new_[13106]_ , \new_[13110]_ ,
    \new_[13111]_ , \new_[13112]_ , \new_[13116]_ , \new_[13117]_ ,
    \new_[13121]_ , \new_[13122]_ , \new_[13123]_ , \new_[13127]_ ,
    \new_[13128]_ , \new_[13132]_ , \new_[13133]_ , \new_[13134]_ ,
    \new_[13138]_ , \new_[13139]_ , \new_[13143]_ , \new_[13144]_ ,
    \new_[13145]_ , \new_[13149]_ , \new_[13150]_ , \new_[13154]_ ,
    \new_[13155]_ , \new_[13156]_ , \new_[13160]_ , \new_[13161]_ ,
    \new_[13165]_ , \new_[13166]_ , \new_[13167]_ , \new_[13171]_ ,
    \new_[13172]_ , \new_[13176]_ , \new_[13177]_ , \new_[13178]_ ,
    \new_[13182]_ , \new_[13183]_ , \new_[13187]_ , \new_[13188]_ ,
    \new_[13189]_ , \new_[13193]_ , \new_[13194]_ , \new_[13198]_ ,
    \new_[13199]_ , \new_[13200]_ , \new_[13204]_ , \new_[13205]_ ,
    \new_[13209]_ , \new_[13210]_ , \new_[13211]_ , \new_[13215]_ ,
    \new_[13216]_ , \new_[13220]_ , \new_[13221]_ , \new_[13222]_ ,
    \new_[13226]_ , \new_[13227]_ , \new_[13231]_ , \new_[13232]_ ,
    \new_[13233]_ , \new_[13237]_ , \new_[13238]_ , \new_[13242]_ ,
    \new_[13243]_ , \new_[13244]_ , \new_[13248]_ , \new_[13249]_ ,
    \new_[13253]_ , \new_[13254]_ , \new_[13255]_ , \new_[13259]_ ,
    \new_[13260]_ , \new_[13264]_ , \new_[13265]_ , \new_[13266]_ ,
    \new_[13270]_ , \new_[13271]_ , \new_[13275]_ , \new_[13276]_ ,
    \new_[13277]_ , \new_[13281]_ , \new_[13282]_ , \new_[13286]_ ,
    \new_[13287]_ , \new_[13288]_ , \new_[13292]_ , \new_[13293]_ ,
    \new_[13297]_ , \new_[13298]_ , \new_[13299]_ , \new_[13303]_ ,
    \new_[13304]_ , \new_[13308]_ , \new_[13309]_ , \new_[13310]_ ,
    \new_[13314]_ , \new_[13315]_ , \new_[13319]_ , \new_[13320]_ ,
    \new_[13321]_ , \new_[13325]_ , \new_[13326]_ , \new_[13330]_ ,
    \new_[13331]_ , \new_[13332]_ , \new_[13336]_ , \new_[13337]_ ,
    \new_[13341]_ , \new_[13342]_ , \new_[13343]_ , \new_[13347]_ ,
    \new_[13348]_ , \new_[13352]_ , \new_[13353]_ , \new_[13354]_ ,
    \new_[13358]_ , \new_[13359]_ , \new_[13363]_ , \new_[13364]_ ,
    \new_[13365]_ , \new_[13369]_ , \new_[13370]_ , \new_[13374]_ ,
    \new_[13375]_ , \new_[13376]_ , \new_[13380]_ , \new_[13381]_ ,
    \new_[13385]_ , \new_[13386]_ , \new_[13387]_ , \new_[13391]_ ,
    \new_[13392]_ , \new_[13396]_ , \new_[13397]_ , \new_[13398]_ ,
    \new_[13402]_ , \new_[13403]_ , \new_[13407]_ , \new_[13408]_ ,
    \new_[13409]_ , \new_[13413]_ , \new_[13414]_ , \new_[13418]_ ,
    \new_[13419]_ , \new_[13420]_ , \new_[13424]_ , \new_[13425]_ ,
    \new_[13429]_ , \new_[13430]_ , \new_[13431]_ , \new_[13435]_ ,
    \new_[13436]_ , \new_[13440]_ , \new_[13441]_ , \new_[13442]_ ,
    \new_[13446]_ , \new_[13447]_ , \new_[13451]_ , \new_[13452]_ ,
    \new_[13453]_ , \new_[13457]_ , \new_[13458]_ , \new_[13462]_ ,
    \new_[13463]_ , \new_[13464]_ , \new_[13468]_ , \new_[13469]_ ,
    \new_[13473]_ , \new_[13474]_ , \new_[13475]_ , \new_[13479]_ ,
    \new_[13480]_ , \new_[13484]_ , \new_[13485]_ , \new_[13486]_ ,
    \new_[13490]_ , \new_[13491]_ , \new_[13495]_ , \new_[13496]_ ,
    \new_[13497]_ , \new_[13501]_ , \new_[13502]_ , \new_[13506]_ ,
    \new_[13507]_ , \new_[13508]_ , \new_[13512]_ , \new_[13513]_ ,
    \new_[13517]_ , \new_[13518]_ , \new_[13519]_ , \new_[13523]_ ,
    \new_[13524]_ , \new_[13528]_ , \new_[13529]_ , \new_[13530]_ ,
    \new_[13534]_ , \new_[13535]_ , \new_[13539]_ , \new_[13540]_ ,
    \new_[13541]_ , \new_[13545]_ , \new_[13546]_ , \new_[13550]_ ,
    \new_[13551]_ , \new_[13552]_ , \new_[13556]_ , \new_[13557]_ ,
    \new_[13561]_ , \new_[13562]_ , \new_[13563]_ , \new_[13567]_ ,
    \new_[13568]_ , \new_[13572]_ , \new_[13573]_ , \new_[13574]_ ,
    \new_[13578]_ , \new_[13579]_ , \new_[13583]_ , \new_[13584]_ ,
    \new_[13585]_ , \new_[13589]_ , \new_[13590]_ , \new_[13594]_ ,
    \new_[13595]_ , \new_[13596]_ , \new_[13600]_ , \new_[13601]_ ,
    \new_[13605]_ , \new_[13606]_ , \new_[13607]_ , \new_[13611]_ ,
    \new_[13612]_ , \new_[13616]_ , \new_[13617]_ , \new_[13618]_ ,
    \new_[13622]_ , \new_[13623]_ , \new_[13627]_ , \new_[13628]_ ,
    \new_[13629]_ , \new_[13633]_ , \new_[13634]_ , \new_[13638]_ ,
    \new_[13639]_ , \new_[13640]_ , \new_[13644]_ , \new_[13645]_ ,
    \new_[13649]_ , \new_[13650]_ , \new_[13651]_ , \new_[13655]_ ,
    \new_[13656]_ , \new_[13660]_ , \new_[13661]_ , \new_[13662]_ ,
    \new_[13666]_ , \new_[13667]_ , \new_[13671]_ , \new_[13672]_ ,
    \new_[13673]_ , \new_[13677]_ , \new_[13678]_ , \new_[13682]_ ,
    \new_[13683]_ , \new_[13684]_ , \new_[13688]_ , \new_[13689]_ ,
    \new_[13693]_ , \new_[13694]_ , \new_[13695]_ , \new_[13699]_ ,
    \new_[13700]_ , \new_[13704]_ , \new_[13705]_ , \new_[13706]_ ,
    \new_[13710]_ , \new_[13711]_ , \new_[13715]_ , \new_[13716]_ ,
    \new_[13717]_ , \new_[13721]_ , \new_[13722]_ , \new_[13726]_ ,
    \new_[13727]_ , \new_[13728]_ , \new_[13732]_ , \new_[13733]_ ,
    \new_[13737]_ , \new_[13738]_ , \new_[13739]_ , \new_[13743]_ ,
    \new_[13744]_ , \new_[13748]_ , \new_[13749]_ , \new_[13750]_ ,
    \new_[13754]_ , \new_[13755]_ , \new_[13759]_ , \new_[13760]_ ,
    \new_[13761]_ , \new_[13765]_ , \new_[13766]_ , \new_[13770]_ ,
    \new_[13771]_ , \new_[13772]_ , \new_[13776]_ , \new_[13777]_ ,
    \new_[13781]_ , \new_[13782]_ , \new_[13783]_ , \new_[13787]_ ,
    \new_[13788]_ , \new_[13792]_ , \new_[13793]_ , \new_[13794]_ ,
    \new_[13798]_ , \new_[13799]_ , \new_[13803]_ , \new_[13804]_ ,
    \new_[13805]_ , \new_[13809]_ , \new_[13810]_ , \new_[13814]_ ,
    \new_[13815]_ , \new_[13816]_ , \new_[13820]_ , \new_[13821]_ ,
    \new_[13825]_ , \new_[13826]_ , \new_[13827]_ , \new_[13831]_ ,
    \new_[13832]_ , \new_[13836]_ , \new_[13837]_ , \new_[13838]_ ,
    \new_[13842]_ , \new_[13843]_ , \new_[13847]_ , \new_[13848]_ ,
    \new_[13849]_ , \new_[13853]_ , \new_[13854]_ , \new_[13858]_ ,
    \new_[13859]_ , \new_[13860]_ , \new_[13864]_ , \new_[13865]_ ,
    \new_[13869]_ , \new_[13870]_ , \new_[13871]_ , \new_[13875]_ ,
    \new_[13876]_ , \new_[13880]_ , \new_[13881]_ , \new_[13882]_ ,
    \new_[13886]_ , \new_[13887]_ , \new_[13891]_ , \new_[13892]_ ,
    \new_[13893]_ , \new_[13897]_ , \new_[13898]_ , \new_[13902]_ ,
    \new_[13903]_ , \new_[13904]_ , \new_[13908]_ , \new_[13909]_ ,
    \new_[13913]_ , \new_[13914]_ , \new_[13915]_ , \new_[13919]_ ,
    \new_[13920]_ , \new_[13924]_ , \new_[13925]_ , \new_[13926]_ ,
    \new_[13930]_ , \new_[13931]_ , \new_[13935]_ , \new_[13936]_ ,
    \new_[13937]_ , \new_[13941]_ , \new_[13942]_ , \new_[13946]_ ,
    \new_[13947]_ , \new_[13948]_ , \new_[13952]_ , \new_[13953]_ ,
    \new_[13957]_ , \new_[13958]_ , \new_[13959]_ , \new_[13963]_ ,
    \new_[13964]_ , \new_[13968]_ , \new_[13969]_ , \new_[13970]_ ,
    \new_[13974]_ , \new_[13975]_ , \new_[13979]_ , \new_[13980]_ ,
    \new_[13981]_ , \new_[13985]_ , \new_[13986]_ , \new_[13990]_ ,
    \new_[13991]_ , \new_[13992]_ , \new_[13996]_ , \new_[13997]_ ,
    \new_[14001]_ , \new_[14002]_ , \new_[14003]_ , \new_[14007]_ ,
    \new_[14008]_ , \new_[14012]_ , \new_[14013]_ , \new_[14014]_ ,
    \new_[14018]_ , \new_[14019]_ , \new_[14023]_ , \new_[14024]_ ,
    \new_[14025]_ , \new_[14029]_ , \new_[14030]_ , \new_[14034]_ ,
    \new_[14035]_ , \new_[14036]_ , \new_[14040]_ , \new_[14041]_ ,
    \new_[14045]_ , \new_[14046]_ , \new_[14047]_ , \new_[14051]_ ,
    \new_[14052]_ , \new_[14056]_ , \new_[14057]_ , \new_[14058]_ ,
    \new_[14062]_ , \new_[14063]_ , \new_[14067]_ , \new_[14068]_ ,
    \new_[14069]_ , \new_[14073]_ , \new_[14074]_ , \new_[14078]_ ,
    \new_[14079]_ , \new_[14080]_ , \new_[14084]_ , \new_[14085]_ ,
    \new_[14089]_ , \new_[14090]_ , \new_[14091]_ , \new_[14095]_ ,
    \new_[14096]_ , \new_[14100]_ , \new_[14101]_ , \new_[14102]_ ,
    \new_[14106]_ , \new_[14107]_ , \new_[14111]_ , \new_[14112]_ ,
    \new_[14113]_ , \new_[14117]_ , \new_[14118]_ , \new_[14122]_ ,
    \new_[14123]_ , \new_[14124]_ , \new_[14128]_ , \new_[14129]_ ,
    \new_[14133]_ , \new_[14134]_ , \new_[14135]_ , \new_[14139]_ ,
    \new_[14140]_ , \new_[14144]_ , \new_[14145]_ , \new_[14146]_ ,
    \new_[14150]_ , \new_[14151]_ , \new_[14155]_ , \new_[14156]_ ,
    \new_[14157]_ , \new_[14161]_ , \new_[14162]_ , \new_[14166]_ ,
    \new_[14167]_ , \new_[14168]_ , \new_[14172]_ , \new_[14173]_ ,
    \new_[14177]_ , \new_[14178]_ , \new_[14179]_ , \new_[14183]_ ,
    \new_[14184]_ , \new_[14188]_ , \new_[14189]_ , \new_[14190]_ ,
    \new_[14194]_ , \new_[14195]_ , \new_[14199]_ , \new_[14200]_ ,
    \new_[14201]_ , \new_[14205]_ , \new_[14206]_ , \new_[14210]_ ,
    \new_[14211]_ , \new_[14212]_ , \new_[14216]_ , \new_[14217]_ ,
    \new_[14221]_ , \new_[14222]_ , \new_[14223]_ , \new_[14227]_ ,
    \new_[14228]_ , \new_[14232]_ , \new_[14233]_ , \new_[14234]_ ,
    \new_[14238]_ , \new_[14239]_ , \new_[14243]_ , \new_[14244]_ ,
    \new_[14245]_ , \new_[14249]_ , \new_[14250]_ , \new_[14254]_ ,
    \new_[14255]_ , \new_[14256]_ , \new_[14260]_ , \new_[14261]_ ,
    \new_[14265]_ , \new_[14266]_ , \new_[14267]_ , \new_[14271]_ ,
    \new_[14272]_ , \new_[14276]_ , \new_[14277]_ , \new_[14278]_ ,
    \new_[14282]_ , \new_[14283]_ , \new_[14287]_ , \new_[14288]_ ,
    \new_[14289]_ , \new_[14293]_ , \new_[14294]_ , \new_[14298]_ ,
    \new_[14299]_ , \new_[14300]_ , \new_[14304]_ , \new_[14305]_ ,
    \new_[14309]_ , \new_[14310]_ , \new_[14311]_ , \new_[14315]_ ,
    \new_[14316]_ , \new_[14320]_ , \new_[14321]_ , \new_[14322]_ ,
    \new_[14326]_ , \new_[14327]_ , \new_[14331]_ , \new_[14332]_ ,
    \new_[14333]_ , \new_[14337]_ , \new_[14338]_ , \new_[14342]_ ,
    \new_[14343]_ , \new_[14344]_ , \new_[14348]_ , \new_[14349]_ ,
    \new_[14353]_ , \new_[14354]_ , \new_[14355]_ , \new_[14359]_ ,
    \new_[14360]_ , \new_[14364]_ , \new_[14365]_ , \new_[14366]_ ,
    \new_[14370]_ , \new_[14371]_ , \new_[14375]_ , \new_[14376]_ ,
    \new_[14377]_ , \new_[14381]_ , \new_[14382]_ , \new_[14386]_ ,
    \new_[14387]_ , \new_[14388]_ , \new_[14392]_ , \new_[14393]_ ,
    \new_[14397]_ , \new_[14398]_ , \new_[14399]_ , \new_[14403]_ ,
    \new_[14404]_ , \new_[14408]_ , \new_[14409]_ , \new_[14410]_ ,
    \new_[14414]_ , \new_[14415]_ , \new_[14419]_ , \new_[14420]_ ,
    \new_[14421]_ , \new_[14425]_ , \new_[14426]_ , \new_[14430]_ ,
    \new_[14431]_ , \new_[14432]_ , \new_[14436]_ , \new_[14437]_ ,
    \new_[14441]_ , \new_[14442]_ , \new_[14443]_ , \new_[14447]_ ,
    \new_[14448]_ , \new_[14452]_ , \new_[14453]_ , \new_[14454]_ ,
    \new_[14458]_ , \new_[14459]_ , \new_[14463]_ , \new_[14464]_ ,
    \new_[14465]_ , \new_[14469]_ , \new_[14470]_ , \new_[14474]_ ,
    \new_[14475]_ , \new_[14476]_ , \new_[14480]_ , \new_[14481]_ ,
    \new_[14485]_ , \new_[14486]_ , \new_[14487]_ , \new_[14491]_ ,
    \new_[14492]_ , \new_[14496]_ , \new_[14497]_ , \new_[14498]_ ,
    \new_[14502]_ , \new_[14503]_ , \new_[14507]_ , \new_[14508]_ ,
    \new_[14509]_ , \new_[14513]_ , \new_[14514]_ , \new_[14518]_ ,
    \new_[14519]_ , \new_[14520]_ , \new_[14524]_ , \new_[14525]_ ,
    \new_[14529]_ , \new_[14530]_ , \new_[14531]_ , \new_[14535]_ ,
    \new_[14536]_ , \new_[14540]_ , \new_[14541]_ , \new_[14542]_ ,
    \new_[14546]_ , \new_[14547]_ , \new_[14551]_ , \new_[14552]_ ,
    \new_[14553]_ , \new_[14557]_ , \new_[14558]_ , \new_[14562]_ ,
    \new_[14563]_ , \new_[14564]_ , \new_[14568]_ , \new_[14569]_ ,
    \new_[14573]_ , \new_[14574]_ , \new_[14575]_ , \new_[14579]_ ,
    \new_[14580]_ , \new_[14584]_ , \new_[14585]_ , \new_[14586]_ ,
    \new_[14590]_ , \new_[14591]_ , \new_[14595]_ , \new_[14596]_ ,
    \new_[14597]_ , \new_[14601]_ , \new_[14602]_ , \new_[14606]_ ,
    \new_[14607]_ , \new_[14608]_ , \new_[14612]_ , \new_[14613]_ ,
    \new_[14617]_ , \new_[14618]_ , \new_[14619]_ , \new_[14623]_ ,
    \new_[14624]_ , \new_[14628]_ , \new_[14629]_ , \new_[14630]_ ,
    \new_[14634]_ , \new_[14635]_ , \new_[14639]_ , \new_[14640]_ ,
    \new_[14641]_ , \new_[14645]_ , \new_[14646]_ , \new_[14650]_ ,
    \new_[14651]_ , \new_[14652]_ , \new_[14656]_ , \new_[14657]_ ,
    \new_[14661]_ , \new_[14662]_ , \new_[14663]_ , \new_[14667]_ ,
    \new_[14668]_ , \new_[14672]_ , \new_[14673]_ , \new_[14674]_ ,
    \new_[14678]_ , \new_[14679]_ , \new_[14683]_ , \new_[14684]_ ,
    \new_[14685]_ , \new_[14689]_ , \new_[14690]_ , \new_[14694]_ ,
    \new_[14695]_ , \new_[14696]_ , \new_[14700]_ , \new_[14701]_ ,
    \new_[14705]_ , \new_[14706]_ , \new_[14707]_ , \new_[14711]_ ,
    \new_[14712]_ , \new_[14716]_ , \new_[14717]_ , \new_[14718]_ ,
    \new_[14722]_ , \new_[14723]_ , \new_[14727]_ , \new_[14728]_ ,
    \new_[14729]_ , \new_[14733]_ , \new_[14734]_ , \new_[14738]_ ,
    \new_[14739]_ , \new_[14740]_ , \new_[14744]_ , \new_[14745]_ ,
    \new_[14749]_ , \new_[14750]_ , \new_[14751]_ , \new_[14755]_ ,
    \new_[14756]_ , \new_[14760]_ , \new_[14761]_ , \new_[14762]_ ,
    \new_[14766]_ , \new_[14767]_ , \new_[14771]_ , \new_[14772]_ ,
    \new_[14773]_ , \new_[14777]_ , \new_[14778]_ , \new_[14782]_ ,
    \new_[14783]_ , \new_[14784]_ , \new_[14788]_ , \new_[14789]_ ,
    \new_[14793]_ , \new_[14794]_ , \new_[14795]_ , \new_[14799]_ ,
    \new_[14800]_ , \new_[14804]_ , \new_[14805]_ , \new_[14806]_ ,
    \new_[14810]_ , \new_[14811]_ , \new_[14815]_ , \new_[14816]_ ,
    \new_[14817]_ , \new_[14821]_ , \new_[14822]_ , \new_[14826]_ ,
    \new_[14827]_ , \new_[14828]_ , \new_[14832]_ , \new_[14833]_ ,
    \new_[14837]_ , \new_[14838]_ , \new_[14839]_ , \new_[14843]_ ,
    \new_[14844]_ , \new_[14848]_ , \new_[14849]_ , \new_[14850]_ ,
    \new_[14854]_ , \new_[14855]_ , \new_[14859]_ , \new_[14860]_ ,
    \new_[14861]_ , \new_[14865]_ , \new_[14866]_ , \new_[14870]_ ,
    \new_[14871]_ , \new_[14872]_ , \new_[14876]_ , \new_[14877]_ ,
    \new_[14881]_ , \new_[14882]_ , \new_[14883]_ , \new_[14887]_ ,
    \new_[14888]_ , \new_[14892]_ , \new_[14893]_ , \new_[14894]_ ,
    \new_[14898]_ , \new_[14899]_ , \new_[14903]_ , \new_[14904]_ ,
    \new_[14905]_ , \new_[14909]_ , \new_[14910]_ , \new_[14914]_ ,
    \new_[14915]_ , \new_[14916]_ , \new_[14920]_ , \new_[14921]_ ,
    \new_[14925]_ , \new_[14926]_ , \new_[14927]_ , \new_[14931]_ ,
    \new_[14932]_ , \new_[14936]_ , \new_[14937]_ , \new_[14938]_ ,
    \new_[14942]_ , \new_[14943]_ , \new_[14947]_ , \new_[14948]_ ,
    \new_[14949]_ , \new_[14953]_ , \new_[14954]_ , \new_[14958]_ ,
    \new_[14959]_ , \new_[14960]_ , \new_[14964]_ , \new_[14965]_ ,
    \new_[14969]_ , \new_[14970]_ , \new_[14971]_ , \new_[14975]_ ,
    \new_[14976]_ , \new_[14980]_ , \new_[14981]_ , \new_[14982]_ ,
    \new_[14986]_ , \new_[14987]_ , \new_[14991]_ , \new_[14992]_ ,
    \new_[14993]_ , \new_[14997]_ , \new_[14998]_ , \new_[15002]_ ,
    \new_[15003]_ , \new_[15004]_ , \new_[15008]_ , \new_[15009]_ ,
    \new_[15013]_ , \new_[15014]_ , \new_[15015]_ , \new_[15019]_ ,
    \new_[15020]_ , \new_[15024]_ , \new_[15025]_ , \new_[15026]_ ,
    \new_[15030]_ , \new_[15031]_ , \new_[15035]_ , \new_[15036]_ ,
    \new_[15037]_ , \new_[15041]_ , \new_[15042]_ , \new_[15046]_ ,
    \new_[15047]_ , \new_[15048]_ , \new_[15052]_ , \new_[15053]_ ,
    \new_[15057]_ , \new_[15058]_ , \new_[15059]_ , \new_[15063]_ ,
    \new_[15064]_ , \new_[15068]_ , \new_[15069]_ , \new_[15070]_ ,
    \new_[15074]_ , \new_[15075]_ , \new_[15079]_ , \new_[15080]_ ,
    \new_[15081]_ , \new_[15085]_ , \new_[15086]_ , \new_[15090]_ ,
    \new_[15091]_ , \new_[15092]_ , \new_[15096]_ , \new_[15097]_ ,
    \new_[15101]_ , \new_[15102]_ , \new_[15103]_ , \new_[15107]_ ,
    \new_[15108]_ , \new_[15112]_ , \new_[15113]_ , \new_[15114]_ ,
    \new_[15118]_ , \new_[15119]_ , \new_[15123]_ , \new_[15124]_ ,
    \new_[15125]_ , \new_[15129]_ , \new_[15130]_ , \new_[15134]_ ,
    \new_[15135]_ , \new_[15136]_ , \new_[15140]_ , \new_[15141]_ ,
    \new_[15145]_ , \new_[15146]_ , \new_[15147]_ , \new_[15151]_ ,
    \new_[15152]_ , \new_[15156]_ , \new_[15157]_ , \new_[15158]_ ,
    \new_[15162]_ , \new_[15163]_ , \new_[15167]_ , \new_[15168]_ ,
    \new_[15169]_ , \new_[15173]_ , \new_[15174]_ , \new_[15178]_ ,
    \new_[15179]_ , \new_[15180]_ , \new_[15184]_ , \new_[15185]_ ,
    \new_[15189]_ , \new_[15190]_ , \new_[15191]_ , \new_[15195]_ ,
    \new_[15196]_ , \new_[15200]_ , \new_[15201]_ , \new_[15202]_ ,
    \new_[15206]_ , \new_[15207]_ , \new_[15211]_ , \new_[15212]_ ,
    \new_[15213]_ , \new_[15217]_ , \new_[15218]_ , \new_[15222]_ ,
    \new_[15223]_ , \new_[15224]_ , \new_[15228]_ , \new_[15229]_ ,
    \new_[15233]_ , \new_[15234]_ , \new_[15235]_ , \new_[15239]_ ,
    \new_[15240]_ , \new_[15244]_ , \new_[15245]_ , \new_[15246]_ ,
    \new_[15250]_ , \new_[15251]_ , \new_[15255]_ , \new_[15256]_ ,
    \new_[15257]_ , \new_[15261]_ , \new_[15262]_ , \new_[15266]_ ,
    \new_[15267]_ , \new_[15268]_ , \new_[15272]_ , \new_[15273]_ ,
    \new_[15277]_ , \new_[15278]_ , \new_[15279]_ , \new_[15283]_ ,
    \new_[15284]_ , \new_[15288]_ , \new_[15289]_ , \new_[15290]_ ,
    \new_[15294]_ , \new_[15295]_ , \new_[15299]_ , \new_[15300]_ ,
    \new_[15301]_ , \new_[15305]_ , \new_[15306]_ , \new_[15310]_ ,
    \new_[15311]_ , \new_[15312]_ , \new_[15316]_ , \new_[15317]_ ,
    \new_[15321]_ , \new_[15322]_ , \new_[15323]_ , \new_[15327]_ ,
    \new_[15328]_ , \new_[15332]_ , \new_[15333]_ , \new_[15334]_ ,
    \new_[15338]_ , \new_[15339]_ , \new_[15343]_ , \new_[15344]_ ,
    \new_[15345]_ , \new_[15349]_ , \new_[15350]_ , \new_[15354]_ ,
    \new_[15355]_ , \new_[15356]_ , \new_[15360]_ , \new_[15361]_ ,
    \new_[15365]_ , \new_[15366]_ , \new_[15367]_ , \new_[15371]_ ,
    \new_[15372]_ , \new_[15376]_ , \new_[15377]_ , \new_[15378]_ ,
    \new_[15382]_ , \new_[15383]_ , \new_[15387]_ , \new_[15388]_ ,
    \new_[15389]_ , \new_[15393]_ , \new_[15394]_ , \new_[15398]_ ,
    \new_[15399]_ , \new_[15400]_ , \new_[15404]_ , \new_[15405]_ ,
    \new_[15409]_ , \new_[15410]_ , \new_[15411]_ , \new_[15415]_ ,
    \new_[15416]_ , \new_[15420]_ , \new_[15421]_ , \new_[15422]_ ,
    \new_[15426]_ , \new_[15427]_ , \new_[15431]_ , \new_[15432]_ ,
    \new_[15433]_ , \new_[15437]_ , \new_[15438]_ , \new_[15442]_ ,
    \new_[15443]_ , \new_[15444]_ , \new_[15448]_ , \new_[15449]_ ,
    \new_[15453]_ , \new_[15454]_ , \new_[15455]_ , \new_[15459]_ ,
    \new_[15460]_ , \new_[15464]_ , \new_[15465]_ , \new_[15466]_ ,
    \new_[15470]_ , \new_[15471]_ , \new_[15475]_ , \new_[15476]_ ,
    \new_[15477]_ , \new_[15481]_ , \new_[15482]_ , \new_[15486]_ ,
    \new_[15487]_ , \new_[15488]_ , \new_[15492]_ , \new_[15493]_ ,
    \new_[15497]_ , \new_[15498]_ , \new_[15499]_ , \new_[15503]_ ,
    \new_[15504]_ , \new_[15508]_ , \new_[15509]_ , \new_[15510]_ ,
    \new_[15514]_ , \new_[15515]_ , \new_[15519]_ , \new_[15520]_ ,
    \new_[15521]_ , \new_[15525]_ , \new_[15526]_ , \new_[15530]_ ,
    \new_[15531]_ , \new_[15532]_ , \new_[15536]_ , \new_[15537]_ ,
    \new_[15541]_ , \new_[15542]_ , \new_[15543]_ , \new_[15547]_ ,
    \new_[15548]_ , \new_[15552]_ , \new_[15553]_ , \new_[15554]_ ,
    \new_[15558]_ , \new_[15559]_ , \new_[15563]_ , \new_[15564]_ ,
    \new_[15565]_ , \new_[15569]_ , \new_[15570]_ , \new_[15574]_ ,
    \new_[15575]_ , \new_[15576]_ , \new_[15580]_ , \new_[15581]_ ,
    \new_[15585]_ , \new_[15586]_ , \new_[15587]_ , \new_[15591]_ ,
    \new_[15592]_ , \new_[15596]_ , \new_[15597]_ , \new_[15598]_ ,
    \new_[15602]_ , \new_[15603]_ , \new_[15607]_ , \new_[15608]_ ,
    \new_[15609]_ , \new_[15613]_ , \new_[15614]_ , \new_[15618]_ ,
    \new_[15619]_ , \new_[15620]_ , \new_[15624]_ , \new_[15625]_ ,
    \new_[15629]_ , \new_[15630]_ , \new_[15631]_ , \new_[15635]_ ,
    \new_[15636]_ , \new_[15640]_ , \new_[15641]_ , \new_[15642]_ ,
    \new_[15646]_ , \new_[15647]_ , \new_[15651]_ , \new_[15652]_ ,
    \new_[15653]_ , \new_[15657]_ , \new_[15658]_ , \new_[15662]_ ,
    \new_[15663]_ , \new_[15664]_ , \new_[15668]_ , \new_[15669]_ ,
    \new_[15673]_ , \new_[15674]_ , \new_[15675]_ , \new_[15679]_ ,
    \new_[15680]_ , \new_[15684]_ , \new_[15685]_ , \new_[15686]_ ,
    \new_[15690]_ , \new_[15691]_ , \new_[15695]_ , \new_[15696]_ ,
    \new_[15697]_ , \new_[15701]_ , \new_[15702]_ , \new_[15706]_ ,
    \new_[15707]_ , \new_[15708]_ , \new_[15712]_ , \new_[15713]_ ,
    \new_[15717]_ , \new_[15718]_ , \new_[15719]_ , \new_[15723]_ ,
    \new_[15724]_ , \new_[15728]_ , \new_[15729]_ , \new_[15730]_ ,
    \new_[15734]_ , \new_[15735]_ , \new_[15739]_ , \new_[15740]_ ,
    \new_[15741]_ , \new_[15745]_ , \new_[15746]_ , \new_[15750]_ ,
    \new_[15751]_ , \new_[15752]_ , \new_[15756]_ , \new_[15757]_ ,
    \new_[15761]_ , \new_[15762]_ , \new_[15763]_ , \new_[15767]_ ,
    \new_[15768]_ , \new_[15772]_ , \new_[15773]_ , \new_[15774]_ ,
    \new_[15778]_ , \new_[15779]_ , \new_[15783]_ , \new_[15784]_ ,
    \new_[15785]_ , \new_[15789]_ , \new_[15790]_ , \new_[15794]_ ,
    \new_[15795]_ , \new_[15796]_ , \new_[15800]_ , \new_[15801]_ ,
    \new_[15805]_ , \new_[15806]_ , \new_[15807]_ , \new_[15811]_ ,
    \new_[15812]_ , \new_[15816]_ , \new_[15817]_ , \new_[15818]_ ,
    \new_[15822]_ , \new_[15823]_ , \new_[15827]_ , \new_[15828]_ ,
    \new_[15829]_ , \new_[15833]_ , \new_[15834]_ , \new_[15838]_ ,
    \new_[15839]_ , \new_[15840]_ , \new_[15844]_ , \new_[15845]_ ,
    \new_[15849]_ , \new_[15850]_ , \new_[15851]_ , \new_[15855]_ ,
    \new_[15856]_ , \new_[15860]_ , \new_[15861]_ , \new_[15862]_ ,
    \new_[15866]_ , \new_[15867]_ , \new_[15871]_ , \new_[15872]_ ,
    \new_[15873]_ , \new_[15877]_ , \new_[15878]_ , \new_[15882]_ ,
    \new_[15883]_ , \new_[15884]_ , \new_[15888]_ , \new_[15889]_ ,
    \new_[15893]_ , \new_[15894]_ , \new_[15895]_ , \new_[15899]_ ,
    \new_[15900]_ , \new_[15904]_ , \new_[15905]_ , \new_[15906]_ ,
    \new_[15910]_ , \new_[15911]_ , \new_[15915]_ , \new_[15916]_ ,
    \new_[15917]_ , \new_[15921]_ , \new_[15922]_ , \new_[15926]_ ,
    \new_[15927]_ , \new_[15928]_ , \new_[15932]_ , \new_[15933]_ ,
    \new_[15937]_ , \new_[15938]_ , \new_[15939]_ , \new_[15943]_ ,
    \new_[15944]_ , \new_[15948]_ , \new_[15949]_ , \new_[15950]_ ,
    \new_[15954]_ , \new_[15955]_ , \new_[15959]_ , \new_[15960]_ ,
    \new_[15961]_ , \new_[15965]_ , \new_[15966]_ , \new_[15970]_ ,
    \new_[15971]_ , \new_[15972]_ , \new_[15976]_ , \new_[15977]_ ,
    \new_[15981]_ , \new_[15982]_ , \new_[15983]_ , \new_[15987]_ ,
    \new_[15988]_ , \new_[15992]_ , \new_[15993]_ , \new_[15994]_ ,
    \new_[15998]_ , \new_[15999]_ , \new_[16003]_ , \new_[16004]_ ,
    \new_[16005]_ , \new_[16009]_ , \new_[16010]_ , \new_[16014]_ ,
    \new_[16015]_ , \new_[16016]_ , \new_[16020]_ , \new_[16021]_ ,
    \new_[16025]_ , \new_[16026]_ , \new_[16027]_ , \new_[16031]_ ,
    \new_[16032]_ , \new_[16036]_ , \new_[16037]_ , \new_[16038]_ ,
    \new_[16042]_ , \new_[16043]_ , \new_[16047]_ , \new_[16048]_ ,
    \new_[16049]_ , \new_[16053]_ , \new_[16054]_ , \new_[16058]_ ,
    \new_[16059]_ , \new_[16060]_ , \new_[16064]_ , \new_[16065]_ ,
    \new_[16069]_ , \new_[16070]_ , \new_[16071]_ , \new_[16075]_ ,
    \new_[16076]_ , \new_[16080]_ , \new_[16081]_ , \new_[16082]_ ,
    \new_[16086]_ , \new_[16087]_ , \new_[16091]_ , \new_[16092]_ ,
    \new_[16093]_ , \new_[16097]_ , \new_[16098]_ , \new_[16102]_ ,
    \new_[16103]_ , \new_[16104]_ , \new_[16108]_ , \new_[16109]_ ,
    \new_[16113]_ , \new_[16114]_ , \new_[16115]_ , \new_[16119]_ ,
    \new_[16120]_ , \new_[16124]_ , \new_[16125]_ , \new_[16126]_ ,
    \new_[16130]_ , \new_[16131]_ , \new_[16135]_ , \new_[16136]_ ,
    \new_[16137]_ , \new_[16141]_ , \new_[16142]_ , \new_[16146]_ ,
    \new_[16147]_ , \new_[16148]_ , \new_[16152]_ , \new_[16153]_ ,
    \new_[16157]_ , \new_[16158]_ , \new_[16159]_ , \new_[16163]_ ,
    \new_[16164]_ , \new_[16168]_ , \new_[16169]_ , \new_[16170]_ ,
    \new_[16174]_ , \new_[16175]_ , \new_[16179]_ , \new_[16180]_ ,
    \new_[16181]_ , \new_[16185]_ , \new_[16186]_ , \new_[16190]_ ,
    \new_[16191]_ , \new_[16192]_ , \new_[16196]_ , \new_[16197]_ ,
    \new_[16201]_ , \new_[16202]_ , \new_[16203]_ , \new_[16207]_ ,
    \new_[16208]_ , \new_[16212]_ , \new_[16213]_ , \new_[16214]_ ,
    \new_[16218]_ , \new_[16219]_ , \new_[16223]_ , \new_[16224]_ ,
    \new_[16225]_ , \new_[16229]_ , \new_[16230]_ , \new_[16234]_ ,
    \new_[16235]_ , \new_[16236]_ , \new_[16240]_ , \new_[16241]_ ,
    \new_[16245]_ , \new_[16246]_ , \new_[16247]_ , \new_[16251]_ ,
    \new_[16252]_ , \new_[16256]_ , \new_[16257]_ , \new_[16258]_ ,
    \new_[16262]_ , \new_[16263]_ , \new_[16267]_ , \new_[16268]_ ,
    \new_[16269]_ , \new_[16273]_ , \new_[16274]_ , \new_[16278]_ ,
    \new_[16279]_ , \new_[16280]_ , \new_[16284]_ , \new_[16285]_ ,
    \new_[16289]_ , \new_[16290]_ , \new_[16291]_ , \new_[16295]_ ,
    \new_[16296]_ , \new_[16300]_ , \new_[16301]_ , \new_[16302]_ ,
    \new_[16306]_ , \new_[16307]_ , \new_[16311]_ , \new_[16312]_ ,
    \new_[16313]_ , \new_[16317]_ , \new_[16318]_ , \new_[16322]_ ,
    \new_[16323]_ , \new_[16324]_ , \new_[16328]_ , \new_[16329]_ ,
    \new_[16333]_ , \new_[16334]_ , \new_[16335]_ , \new_[16339]_ ,
    \new_[16340]_ , \new_[16344]_ , \new_[16345]_ , \new_[16346]_ ,
    \new_[16350]_ , \new_[16351]_ , \new_[16355]_ , \new_[16356]_ ,
    \new_[16357]_ , \new_[16361]_ , \new_[16362]_ , \new_[16366]_ ,
    \new_[16367]_ , \new_[16368]_ , \new_[16372]_ , \new_[16373]_ ,
    \new_[16377]_ , \new_[16378]_ , \new_[16379]_ , \new_[16383]_ ,
    \new_[16384]_ , \new_[16388]_ , \new_[16389]_ , \new_[16390]_ ,
    \new_[16394]_ , \new_[16395]_ , \new_[16399]_ , \new_[16400]_ ,
    \new_[16401]_ , \new_[16405]_ , \new_[16406]_ , \new_[16410]_ ,
    \new_[16411]_ , \new_[16412]_ , \new_[16416]_ , \new_[16417]_ ,
    \new_[16421]_ , \new_[16422]_ , \new_[16423]_ , \new_[16427]_ ,
    \new_[16428]_ , \new_[16432]_ , \new_[16433]_ , \new_[16434]_ ,
    \new_[16438]_ , \new_[16439]_ , \new_[16443]_ , \new_[16444]_ ,
    \new_[16445]_ , \new_[16449]_ , \new_[16450]_ , \new_[16454]_ ,
    \new_[16455]_ , \new_[16456]_ , \new_[16460]_ , \new_[16461]_ ,
    \new_[16465]_ , \new_[16466]_ , \new_[16467]_ , \new_[16471]_ ,
    \new_[16472]_ , \new_[16476]_ , \new_[16477]_ , \new_[16478]_ ,
    \new_[16482]_ , \new_[16483]_ , \new_[16487]_ , \new_[16488]_ ,
    \new_[16489]_ , \new_[16493]_ , \new_[16494]_ , \new_[16498]_ ,
    \new_[16499]_ , \new_[16500]_ , \new_[16504]_ , \new_[16505]_ ,
    \new_[16509]_ , \new_[16510]_ , \new_[16511]_ , \new_[16515]_ ,
    \new_[16516]_ , \new_[16520]_ , \new_[16521]_ , \new_[16522]_ ,
    \new_[16526]_ , \new_[16527]_ , \new_[16531]_ , \new_[16532]_ ,
    \new_[16533]_ , \new_[16537]_ , \new_[16538]_ , \new_[16542]_ ,
    \new_[16543]_ , \new_[16544]_ , \new_[16548]_ , \new_[16549]_ ,
    \new_[16553]_ , \new_[16554]_ , \new_[16555]_ , \new_[16559]_ ,
    \new_[16560]_ , \new_[16564]_ , \new_[16565]_ , \new_[16566]_ ,
    \new_[16570]_ , \new_[16571]_ , \new_[16575]_ , \new_[16576]_ ,
    \new_[16577]_ , \new_[16581]_ , \new_[16582]_ , \new_[16586]_ ,
    \new_[16587]_ , \new_[16588]_ , \new_[16592]_ , \new_[16593]_ ,
    \new_[16597]_ , \new_[16598]_ , \new_[16599]_ , \new_[16603]_ ,
    \new_[16604]_ , \new_[16608]_ , \new_[16609]_ , \new_[16610]_ ,
    \new_[16614]_ , \new_[16615]_ , \new_[16619]_ , \new_[16620]_ ,
    \new_[16621]_ , \new_[16625]_ , \new_[16626]_ , \new_[16630]_ ,
    \new_[16631]_ , \new_[16632]_ , \new_[16636]_ , \new_[16637]_ ,
    \new_[16641]_ , \new_[16642]_ , \new_[16643]_ , \new_[16647]_ ,
    \new_[16648]_ , \new_[16652]_ , \new_[16653]_ , \new_[16654]_ ,
    \new_[16658]_ , \new_[16659]_ , \new_[16663]_ , \new_[16664]_ ,
    \new_[16665]_ , \new_[16669]_ , \new_[16670]_ , \new_[16674]_ ,
    \new_[16675]_ , \new_[16676]_ , \new_[16680]_ , \new_[16681]_ ,
    \new_[16685]_ , \new_[16686]_ , \new_[16687]_ , \new_[16691]_ ,
    \new_[16692]_ , \new_[16696]_ , \new_[16697]_ , \new_[16698]_ ,
    \new_[16702]_ , \new_[16703]_ , \new_[16707]_ , \new_[16708]_ ,
    \new_[16709]_ , \new_[16713]_ , \new_[16714]_ , \new_[16718]_ ,
    \new_[16719]_ , \new_[16720]_ , \new_[16724]_ , \new_[16725]_ ,
    \new_[16729]_ , \new_[16730]_ , \new_[16731]_ , \new_[16735]_ ,
    \new_[16736]_ , \new_[16740]_ , \new_[16741]_ , \new_[16742]_ ,
    \new_[16746]_ , \new_[16747]_ , \new_[16751]_ , \new_[16752]_ ,
    \new_[16753]_ , \new_[16757]_ , \new_[16758]_ , \new_[16762]_ ,
    \new_[16763]_ , \new_[16764]_ , \new_[16768]_ , \new_[16769]_ ,
    \new_[16773]_ , \new_[16774]_ , \new_[16775]_ , \new_[16779]_ ,
    \new_[16780]_ , \new_[16784]_ , \new_[16785]_ , \new_[16786]_ ,
    \new_[16790]_ , \new_[16791]_ , \new_[16795]_ , \new_[16796]_ ,
    \new_[16797]_ , \new_[16801]_ , \new_[16802]_ , \new_[16806]_ ,
    \new_[16807]_ , \new_[16808]_ , \new_[16812]_ , \new_[16813]_ ,
    \new_[16817]_ , \new_[16818]_ , \new_[16819]_ , \new_[16823]_ ,
    \new_[16824]_ , \new_[16828]_ , \new_[16829]_ , \new_[16830]_ ,
    \new_[16834]_ , \new_[16835]_ , \new_[16839]_ , \new_[16840]_ ,
    \new_[16841]_ , \new_[16845]_ , \new_[16846]_ , \new_[16850]_ ,
    \new_[16851]_ , \new_[16852]_ , \new_[16856]_ , \new_[16857]_ ,
    \new_[16861]_ , \new_[16862]_ , \new_[16863]_ , \new_[16867]_ ,
    \new_[16868]_ , \new_[16872]_ , \new_[16873]_ , \new_[16874]_ ,
    \new_[16878]_ , \new_[16879]_ , \new_[16883]_ , \new_[16884]_ ,
    \new_[16885]_ , \new_[16889]_ , \new_[16890]_ , \new_[16894]_ ,
    \new_[16895]_ , \new_[16896]_ , \new_[16900]_ , \new_[16901]_ ,
    \new_[16905]_ , \new_[16906]_ , \new_[16907]_ , \new_[16911]_ ,
    \new_[16912]_ , \new_[16916]_ , \new_[16917]_ , \new_[16918]_ ,
    \new_[16922]_ , \new_[16923]_ , \new_[16927]_ , \new_[16928]_ ,
    \new_[16929]_ , \new_[16933]_ , \new_[16934]_ , \new_[16938]_ ,
    \new_[16939]_ , \new_[16940]_ , \new_[16944]_ , \new_[16945]_ ,
    \new_[16949]_ , \new_[16950]_ , \new_[16951]_ , \new_[16955]_ ,
    \new_[16956]_ , \new_[16960]_ , \new_[16961]_ , \new_[16962]_ ,
    \new_[16966]_ , \new_[16967]_ , \new_[16971]_ , \new_[16972]_ ,
    \new_[16973]_ , \new_[16977]_ , \new_[16978]_ , \new_[16982]_ ,
    \new_[16983]_ , \new_[16984]_ , \new_[16988]_ , \new_[16989]_ ,
    \new_[16993]_ , \new_[16994]_ , \new_[16995]_ , \new_[16999]_ ,
    \new_[17000]_ , \new_[17004]_ , \new_[17005]_ , \new_[17006]_ ,
    \new_[17010]_ , \new_[17011]_ , \new_[17015]_ , \new_[17016]_ ,
    \new_[17017]_ , \new_[17021]_ , \new_[17022]_ , \new_[17026]_ ,
    \new_[17027]_ , \new_[17028]_ , \new_[17032]_ , \new_[17033]_ ,
    \new_[17037]_ , \new_[17038]_ , \new_[17039]_ , \new_[17043]_ ,
    \new_[17044]_ , \new_[17048]_ , \new_[17049]_ , \new_[17050]_ ,
    \new_[17054]_ , \new_[17055]_ , \new_[17059]_ , \new_[17060]_ ,
    \new_[17061]_ , \new_[17065]_ , \new_[17066]_ , \new_[17070]_ ,
    \new_[17071]_ , \new_[17072]_ , \new_[17076]_ , \new_[17077]_ ,
    \new_[17081]_ , \new_[17082]_ , \new_[17083]_ , \new_[17087]_ ,
    \new_[17088]_ , \new_[17092]_ , \new_[17093]_ , \new_[17094]_ ,
    \new_[17098]_ , \new_[17099]_ , \new_[17103]_ , \new_[17104]_ ,
    \new_[17105]_ , \new_[17109]_ , \new_[17110]_ , \new_[17114]_ ,
    \new_[17115]_ , \new_[17116]_ , \new_[17120]_ , \new_[17121]_ ,
    \new_[17125]_ , \new_[17126]_ , \new_[17127]_ , \new_[17131]_ ,
    \new_[17132]_ , \new_[17136]_ , \new_[17137]_ , \new_[17138]_ ,
    \new_[17142]_ , \new_[17143]_ , \new_[17147]_ , \new_[17148]_ ,
    \new_[17149]_ , \new_[17153]_ , \new_[17154]_ , \new_[17158]_ ,
    \new_[17159]_ , \new_[17160]_ , \new_[17164]_ , \new_[17165]_ ,
    \new_[17169]_ , \new_[17170]_ , \new_[17171]_ , \new_[17175]_ ,
    \new_[17176]_ , \new_[17180]_ , \new_[17181]_ , \new_[17182]_ ,
    \new_[17186]_ , \new_[17187]_ , \new_[17191]_ , \new_[17192]_ ,
    \new_[17193]_ , \new_[17197]_ , \new_[17198]_ , \new_[17202]_ ,
    \new_[17203]_ , \new_[17204]_ , \new_[17208]_ , \new_[17209]_ ,
    \new_[17213]_ , \new_[17214]_ , \new_[17215]_ , \new_[17219]_ ,
    \new_[17220]_ , \new_[17224]_ , \new_[17225]_ , \new_[17226]_ ,
    \new_[17230]_ , \new_[17231]_ , \new_[17235]_ , \new_[17236]_ ,
    \new_[17237]_ , \new_[17241]_ , \new_[17242]_ , \new_[17246]_ ,
    \new_[17247]_ , \new_[17248]_ , \new_[17252]_ , \new_[17253]_ ,
    \new_[17257]_ , \new_[17258]_ , \new_[17259]_ , \new_[17263]_ ,
    \new_[17264]_ , \new_[17268]_ , \new_[17269]_ , \new_[17270]_ ,
    \new_[17274]_ , \new_[17275]_ , \new_[17279]_ , \new_[17280]_ ,
    \new_[17281]_ , \new_[17285]_ , \new_[17286]_ , \new_[17290]_ ,
    \new_[17291]_ , \new_[17292]_ , \new_[17296]_ , \new_[17297]_ ,
    \new_[17301]_ , \new_[17302]_ , \new_[17303]_ , \new_[17307]_ ,
    \new_[17308]_ , \new_[17312]_ , \new_[17313]_ , \new_[17314]_ ,
    \new_[17318]_ , \new_[17319]_ , \new_[17323]_ , \new_[17324]_ ,
    \new_[17325]_ , \new_[17329]_ , \new_[17330]_ , \new_[17334]_ ,
    \new_[17335]_ , \new_[17336]_ , \new_[17340]_ , \new_[17341]_ ,
    \new_[17345]_ , \new_[17346]_ , \new_[17347]_ , \new_[17351]_ ,
    \new_[17352]_ , \new_[17356]_ , \new_[17357]_ , \new_[17358]_ ,
    \new_[17362]_ , \new_[17363]_ , \new_[17367]_ , \new_[17368]_ ,
    \new_[17369]_ , \new_[17373]_ , \new_[17374]_ , \new_[17378]_ ,
    \new_[17379]_ , \new_[17380]_ , \new_[17384]_ , \new_[17385]_ ,
    \new_[17389]_ , \new_[17390]_ , \new_[17391]_ , \new_[17395]_ ,
    \new_[17396]_ , \new_[17400]_ , \new_[17401]_ , \new_[17402]_ ,
    \new_[17406]_ , \new_[17407]_ , \new_[17411]_ , \new_[17412]_ ,
    \new_[17413]_ , \new_[17417]_ , \new_[17418]_ , \new_[17422]_ ,
    \new_[17423]_ , \new_[17424]_ , \new_[17428]_ , \new_[17429]_ ,
    \new_[17433]_ , \new_[17434]_ , \new_[17435]_ , \new_[17439]_ ,
    \new_[17440]_ , \new_[17444]_ , \new_[17445]_ , \new_[17446]_ ,
    \new_[17450]_ , \new_[17451]_ , \new_[17455]_ , \new_[17456]_ ,
    \new_[17457]_ , \new_[17461]_ , \new_[17462]_ , \new_[17466]_ ,
    \new_[17467]_ , \new_[17468]_ , \new_[17472]_ , \new_[17473]_ ,
    \new_[17477]_ , \new_[17478]_ , \new_[17479]_ , \new_[17483]_ ,
    \new_[17484]_ , \new_[17488]_ , \new_[17489]_ , \new_[17490]_ ,
    \new_[17494]_ , \new_[17495]_ , \new_[17499]_ , \new_[17500]_ ,
    \new_[17501]_ , \new_[17505]_ , \new_[17506]_ , \new_[17510]_ ,
    \new_[17511]_ , \new_[17512]_ , \new_[17516]_ , \new_[17517]_ ,
    \new_[17521]_ , \new_[17522]_ , \new_[17523]_ , \new_[17527]_ ,
    \new_[17528]_ , \new_[17532]_ , \new_[17533]_ , \new_[17534]_ ,
    \new_[17538]_ , \new_[17539]_ , \new_[17543]_ , \new_[17544]_ ,
    \new_[17545]_ , \new_[17549]_ , \new_[17550]_ , \new_[17554]_ ,
    \new_[17555]_ , \new_[17556]_ , \new_[17560]_ , \new_[17561]_ ,
    \new_[17565]_ , \new_[17566]_ , \new_[17567]_ , \new_[17571]_ ,
    \new_[17572]_ , \new_[17576]_ , \new_[17577]_ , \new_[17578]_ ,
    \new_[17582]_ , \new_[17583]_ , \new_[17587]_ , \new_[17588]_ ,
    \new_[17589]_ , \new_[17593]_ , \new_[17594]_ , \new_[17598]_ ,
    \new_[17599]_ , \new_[17600]_ , \new_[17604]_ , \new_[17605]_ ,
    \new_[17609]_ , \new_[17610]_ , \new_[17611]_ , \new_[17615]_ ,
    \new_[17616]_ , \new_[17620]_ , \new_[17621]_ , \new_[17622]_ ,
    \new_[17626]_ , \new_[17627]_ , \new_[17631]_ , \new_[17632]_ ,
    \new_[17633]_ , \new_[17637]_ , \new_[17638]_ , \new_[17642]_ ,
    \new_[17643]_ , \new_[17644]_ , \new_[17648]_ , \new_[17649]_ ,
    \new_[17653]_ , \new_[17654]_ , \new_[17655]_ , \new_[17659]_ ,
    \new_[17660]_ , \new_[17664]_ , \new_[17665]_ , \new_[17666]_ ,
    \new_[17670]_ , \new_[17671]_ , \new_[17675]_ , \new_[17676]_ ,
    \new_[17677]_ , \new_[17681]_ , \new_[17682]_ , \new_[17686]_ ,
    \new_[17687]_ , \new_[17688]_ , \new_[17692]_ , \new_[17693]_ ,
    \new_[17697]_ , \new_[17698]_ , \new_[17699]_ , \new_[17703]_ ,
    \new_[17704]_ , \new_[17708]_ , \new_[17709]_ , \new_[17710]_ ,
    \new_[17714]_ , \new_[17715]_ , \new_[17719]_ , \new_[17720]_ ,
    \new_[17721]_ , \new_[17725]_ , \new_[17726]_ , \new_[17730]_ ,
    \new_[17731]_ , \new_[17732]_ , \new_[17736]_ , \new_[17737]_ ,
    \new_[17741]_ , \new_[17742]_ , \new_[17743]_ , \new_[17747]_ ,
    \new_[17748]_ , \new_[17752]_ , \new_[17753]_ , \new_[17754]_ ,
    \new_[17758]_ , \new_[17759]_ , \new_[17763]_ , \new_[17764]_ ,
    \new_[17765]_ , \new_[17769]_ , \new_[17770]_ , \new_[17774]_ ,
    \new_[17775]_ , \new_[17776]_ , \new_[17780]_ , \new_[17781]_ ,
    \new_[17785]_ , \new_[17786]_ , \new_[17787]_ , \new_[17791]_ ,
    \new_[17792]_ , \new_[17796]_ , \new_[17797]_ , \new_[17798]_ ,
    \new_[17802]_ , \new_[17803]_ , \new_[17807]_ , \new_[17808]_ ,
    \new_[17809]_ , \new_[17813]_ , \new_[17814]_ , \new_[17818]_ ,
    \new_[17819]_ , \new_[17820]_ , \new_[17824]_ , \new_[17825]_ ,
    \new_[17829]_ , \new_[17830]_ , \new_[17831]_ , \new_[17835]_ ,
    \new_[17836]_ , \new_[17840]_ , \new_[17841]_ , \new_[17842]_ ,
    \new_[17846]_ , \new_[17847]_ , \new_[17851]_ , \new_[17852]_ ,
    \new_[17853]_ , \new_[17857]_ , \new_[17858]_ , \new_[17862]_ ,
    \new_[17863]_ , \new_[17864]_ , \new_[17868]_ , \new_[17869]_ ,
    \new_[17873]_ , \new_[17874]_ , \new_[17875]_ , \new_[17879]_ ,
    \new_[17880]_ , \new_[17884]_ , \new_[17885]_ , \new_[17886]_ ,
    \new_[17890]_ , \new_[17891]_ , \new_[17895]_ , \new_[17896]_ ,
    \new_[17897]_ , \new_[17901]_ , \new_[17902]_ , \new_[17906]_ ,
    \new_[17907]_ , \new_[17908]_ , \new_[17912]_ , \new_[17913]_ ,
    \new_[17917]_ , \new_[17918]_ , \new_[17919]_ , \new_[17923]_ ,
    \new_[17924]_ , \new_[17928]_ , \new_[17929]_ , \new_[17930]_ ,
    \new_[17934]_ , \new_[17935]_ , \new_[17939]_ , \new_[17940]_ ,
    \new_[17941]_ , \new_[17945]_ , \new_[17946]_ , \new_[17950]_ ,
    \new_[17951]_ , \new_[17952]_ , \new_[17956]_ , \new_[17957]_ ,
    \new_[17961]_ , \new_[17962]_ , \new_[17963]_ , \new_[17967]_ ,
    \new_[17968]_ , \new_[17972]_ , \new_[17973]_ , \new_[17974]_ ,
    \new_[17978]_ , \new_[17979]_ , \new_[17983]_ , \new_[17984]_ ,
    \new_[17985]_ , \new_[17989]_ , \new_[17990]_ , \new_[17994]_ ,
    \new_[17995]_ , \new_[17996]_ , \new_[18000]_ , \new_[18001]_ ,
    \new_[18005]_ , \new_[18006]_ , \new_[18007]_ , \new_[18011]_ ,
    \new_[18012]_ , \new_[18016]_ , \new_[18017]_ , \new_[18018]_ ,
    \new_[18022]_ , \new_[18023]_ , \new_[18027]_ , \new_[18028]_ ,
    \new_[18029]_ , \new_[18033]_ , \new_[18034]_ , \new_[18038]_ ,
    \new_[18039]_ , \new_[18040]_ , \new_[18044]_ , \new_[18045]_ ,
    \new_[18049]_ , \new_[18050]_ , \new_[18051]_ , \new_[18055]_ ,
    \new_[18056]_ , \new_[18060]_ , \new_[18061]_ , \new_[18062]_ ,
    \new_[18066]_ , \new_[18067]_ , \new_[18071]_ , \new_[18072]_ ,
    \new_[18073]_ , \new_[18077]_ , \new_[18078]_ , \new_[18082]_ ,
    \new_[18083]_ , \new_[18084]_ , \new_[18088]_ , \new_[18089]_ ,
    \new_[18093]_ , \new_[18094]_ , \new_[18095]_ , \new_[18099]_ ,
    \new_[18100]_ , \new_[18104]_ , \new_[18105]_ , \new_[18106]_ ,
    \new_[18110]_ , \new_[18111]_ , \new_[18115]_ , \new_[18116]_ ,
    \new_[18117]_ , \new_[18121]_ , \new_[18122]_ , \new_[18126]_ ,
    \new_[18127]_ , \new_[18128]_ , \new_[18132]_ , \new_[18133]_ ,
    \new_[18137]_ , \new_[18138]_ , \new_[18139]_ , \new_[18143]_ ,
    \new_[18144]_ , \new_[18148]_ , \new_[18149]_ , \new_[18150]_ ,
    \new_[18154]_ , \new_[18155]_ , \new_[18159]_ , \new_[18160]_ ,
    \new_[18161]_ , \new_[18165]_ , \new_[18166]_ , \new_[18170]_ ,
    \new_[18171]_ , \new_[18172]_ , \new_[18176]_ , \new_[18177]_ ,
    \new_[18181]_ , \new_[18182]_ , \new_[18183]_ , \new_[18187]_ ,
    \new_[18188]_ , \new_[18192]_ , \new_[18193]_ , \new_[18194]_ ,
    \new_[18198]_ , \new_[18199]_ , \new_[18203]_ , \new_[18204]_ ,
    \new_[18205]_ , \new_[18209]_ , \new_[18210]_ , \new_[18214]_ ,
    \new_[18215]_ , \new_[18216]_ , \new_[18220]_ , \new_[18221]_ ,
    \new_[18225]_ , \new_[18226]_ , \new_[18227]_ , \new_[18231]_ ,
    \new_[18232]_ , \new_[18236]_ , \new_[18237]_ , \new_[18238]_ ,
    \new_[18242]_ , \new_[18243]_ , \new_[18247]_ , \new_[18248]_ ,
    \new_[18249]_ , \new_[18253]_ , \new_[18254]_ , \new_[18258]_ ,
    \new_[18259]_ , \new_[18260]_ , \new_[18264]_ , \new_[18265]_ ,
    \new_[18269]_ , \new_[18270]_ , \new_[18271]_ , \new_[18275]_ ,
    \new_[18276]_ , \new_[18280]_ , \new_[18281]_ , \new_[18282]_ ,
    \new_[18286]_ , \new_[18287]_ , \new_[18291]_ , \new_[18292]_ ,
    \new_[18293]_ , \new_[18297]_ , \new_[18298]_ , \new_[18302]_ ,
    \new_[18303]_ , \new_[18304]_ , \new_[18308]_ , \new_[18309]_ ,
    \new_[18313]_ , \new_[18314]_ , \new_[18315]_ , \new_[18319]_ ,
    \new_[18320]_ , \new_[18324]_ , \new_[18325]_ , \new_[18326]_ ,
    \new_[18330]_ , \new_[18331]_ , \new_[18335]_ , \new_[18336]_ ,
    \new_[18337]_ , \new_[18341]_ , \new_[18342]_ , \new_[18346]_ ,
    \new_[18347]_ , \new_[18348]_ , \new_[18352]_ , \new_[18353]_ ,
    \new_[18357]_ , \new_[18358]_ , \new_[18359]_ , \new_[18363]_ ,
    \new_[18364]_ , \new_[18368]_ , \new_[18369]_ , \new_[18370]_ ,
    \new_[18374]_ , \new_[18375]_ , \new_[18379]_ , \new_[18380]_ ,
    \new_[18381]_ , \new_[18385]_ , \new_[18386]_ , \new_[18390]_ ,
    \new_[18391]_ , \new_[18392]_ , \new_[18396]_ , \new_[18397]_ ,
    \new_[18401]_ , \new_[18402]_ , \new_[18403]_ , \new_[18407]_ ,
    \new_[18408]_ , \new_[18412]_ , \new_[18413]_ , \new_[18414]_ ,
    \new_[18418]_ , \new_[18419]_ , \new_[18423]_ , \new_[18424]_ ,
    \new_[18425]_ , \new_[18429]_ , \new_[18430]_ , \new_[18434]_ ,
    \new_[18435]_ , \new_[18436]_ , \new_[18440]_ , \new_[18441]_ ,
    \new_[18445]_ , \new_[18446]_ , \new_[18447]_ , \new_[18451]_ ,
    \new_[18452]_ , \new_[18456]_ , \new_[18457]_ , \new_[18458]_ ,
    \new_[18462]_ , \new_[18463]_ , \new_[18467]_ , \new_[18468]_ ,
    \new_[18469]_ , \new_[18473]_ , \new_[18474]_ , \new_[18478]_ ,
    \new_[18479]_ , \new_[18480]_ , \new_[18484]_ , \new_[18485]_ ,
    \new_[18489]_ , \new_[18490]_ , \new_[18491]_ , \new_[18495]_ ,
    \new_[18496]_ , \new_[18500]_ , \new_[18501]_ , \new_[18502]_ ,
    \new_[18506]_ , \new_[18507]_ , \new_[18511]_ , \new_[18512]_ ,
    \new_[18513]_ , \new_[18517]_ , \new_[18518]_ , \new_[18522]_ ,
    \new_[18523]_ , \new_[18524]_ , \new_[18528]_ , \new_[18529]_ ,
    \new_[18533]_ , \new_[18534]_ , \new_[18535]_ , \new_[18539]_ ,
    \new_[18540]_ , \new_[18544]_ , \new_[18545]_ , \new_[18546]_ ,
    \new_[18550]_ , \new_[18551]_ , \new_[18555]_ , \new_[18556]_ ,
    \new_[18557]_ , \new_[18561]_ , \new_[18562]_ , \new_[18566]_ ,
    \new_[18567]_ , \new_[18568]_ , \new_[18572]_ , \new_[18573]_ ,
    \new_[18577]_ , \new_[18578]_ , \new_[18579]_ , \new_[18583]_ ,
    \new_[18584]_ , \new_[18588]_ , \new_[18589]_ , \new_[18590]_ ,
    \new_[18594]_ , \new_[18595]_ , \new_[18599]_ , \new_[18600]_ ,
    \new_[18601]_ , \new_[18605]_ , \new_[18606]_ , \new_[18610]_ ,
    \new_[18611]_ , \new_[18612]_ , \new_[18616]_ , \new_[18617]_ ,
    \new_[18621]_ , \new_[18622]_ , \new_[18623]_ , \new_[18627]_ ,
    \new_[18628]_ , \new_[18632]_ , \new_[18633]_ , \new_[18634]_ ,
    \new_[18638]_ , \new_[18639]_ , \new_[18643]_ , \new_[18644]_ ,
    \new_[18645]_ , \new_[18649]_ , \new_[18650]_ , \new_[18654]_ ,
    \new_[18655]_ , \new_[18656]_ , \new_[18660]_ , \new_[18661]_ ,
    \new_[18665]_ , \new_[18666]_ , \new_[18667]_ , \new_[18671]_ ,
    \new_[18672]_ , \new_[18676]_ , \new_[18677]_ , \new_[18678]_ ,
    \new_[18682]_ , \new_[18683]_ , \new_[18687]_ , \new_[18688]_ ,
    \new_[18689]_ , \new_[18693]_ , \new_[18694]_ , \new_[18698]_ ,
    \new_[18699]_ , \new_[18700]_ , \new_[18704]_ , \new_[18705]_ ,
    \new_[18709]_ , \new_[18710]_ , \new_[18711]_ , \new_[18715]_ ,
    \new_[18716]_ , \new_[18720]_ , \new_[18721]_ , \new_[18722]_ ,
    \new_[18726]_ , \new_[18727]_ , \new_[18731]_ , \new_[18732]_ ,
    \new_[18733]_ , \new_[18737]_ , \new_[18738]_ , \new_[18742]_ ,
    \new_[18743]_ , \new_[18744]_ , \new_[18748]_ , \new_[18749]_ ,
    \new_[18753]_ , \new_[18754]_ , \new_[18755]_ , \new_[18759]_ ,
    \new_[18760]_ , \new_[18764]_ , \new_[18765]_ , \new_[18766]_ ,
    \new_[18770]_ , \new_[18771]_ , \new_[18775]_ , \new_[18776]_ ,
    \new_[18777]_ , \new_[18781]_ , \new_[18782]_ , \new_[18786]_ ,
    \new_[18787]_ , \new_[18788]_ , \new_[18792]_ , \new_[18793]_ ,
    \new_[18797]_ , \new_[18798]_ , \new_[18799]_ , \new_[18803]_ ,
    \new_[18804]_ , \new_[18808]_ , \new_[18809]_ , \new_[18810]_ ,
    \new_[18814]_ , \new_[18815]_ , \new_[18819]_ , \new_[18820]_ ,
    \new_[18821]_ , \new_[18825]_ , \new_[18826]_ , \new_[18830]_ ,
    \new_[18831]_ , \new_[18832]_ , \new_[18836]_ , \new_[18837]_ ,
    \new_[18841]_ , \new_[18842]_ , \new_[18843]_ , \new_[18847]_ ,
    \new_[18848]_ , \new_[18852]_ , \new_[18853]_ , \new_[18854]_ ,
    \new_[18858]_ , \new_[18859]_ , \new_[18863]_ , \new_[18864]_ ,
    \new_[18865]_ , \new_[18869]_ , \new_[18870]_ , \new_[18874]_ ,
    \new_[18875]_ , \new_[18876]_ , \new_[18880]_ , \new_[18881]_ ,
    \new_[18885]_ , \new_[18886]_ , \new_[18887]_ , \new_[18891]_ ,
    \new_[18892]_ , \new_[18896]_ , \new_[18897]_ , \new_[18898]_ ,
    \new_[18902]_ , \new_[18903]_ , \new_[18907]_ , \new_[18908]_ ,
    \new_[18909]_ , \new_[18913]_ , \new_[18914]_ , \new_[18918]_ ,
    \new_[18919]_ , \new_[18920]_ , \new_[18924]_ , \new_[18925]_ ,
    \new_[18929]_ , \new_[18930]_ , \new_[18931]_ , \new_[18935]_ ,
    \new_[18936]_ , \new_[18940]_ , \new_[18941]_ , \new_[18942]_ ,
    \new_[18946]_ , \new_[18947]_ , \new_[18951]_ , \new_[18952]_ ,
    \new_[18953]_ , \new_[18957]_ , \new_[18958]_ , \new_[18962]_ ,
    \new_[18963]_ , \new_[18964]_ , \new_[18968]_ , \new_[18969]_ ,
    \new_[18973]_ , \new_[18974]_ , \new_[18975]_ , \new_[18979]_ ,
    \new_[18980]_ , \new_[18984]_ , \new_[18985]_ , \new_[18986]_ ,
    \new_[18990]_ , \new_[18991]_ , \new_[18995]_ , \new_[18996]_ ,
    \new_[18997]_ , \new_[19001]_ , \new_[19002]_ , \new_[19006]_ ,
    \new_[19007]_ , \new_[19008]_ , \new_[19012]_ , \new_[19013]_ ,
    \new_[19017]_ , \new_[19018]_ , \new_[19019]_ , \new_[19023]_ ,
    \new_[19024]_ , \new_[19028]_ , \new_[19029]_ , \new_[19030]_ ,
    \new_[19034]_ , \new_[19035]_ , \new_[19038]_ , \new_[19041]_ ,
    \new_[19042]_ , \new_[19043]_ , \new_[19047]_ , \new_[19048]_ ,
    \new_[19052]_ , \new_[19053]_ , \new_[19054]_ , \new_[19058]_ ,
    \new_[19059]_ , \new_[19062]_ , \new_[19065]_ , \new_[19066]_ ,
    \new_[19067]_ , \new_[19071]_ , \new_[19072]_ , \new_[19076]_ ,
    \new_[19077]_ , \new_[19078]_ , \new_[19082]_ , \new_[19083]_ ,
    \new_[19086]_ , \new_[19089]_ , \new_[19090]_ , \new_[19091]_ ,
    \new_[19095]_ , \new_[19096]_ , \new_[19100]_ , \new_[19101]_ ,
    \new_[19102]_ , \new_[19106]_ , \new_[19107]_ , \new_[19110]_ ,
    \new_[19113]_ , \new_[19114]_ , \new_[19115]_ , \new_[19119]_ ,
    \new_[19120]_ , \new_[19124]_ , \new_[19125]_ , \new_[19126]_ ,
    \new_[19130]_ , \new_[19131]_ , \new_[19134]_ , \new_[19137]_ ,
    \new_[19138]_ , \new_[19139]_ , \new_[19143]_ , \new_[19144]_ ,
    \new_[19148]_ , \new_[19149]_ , \new_[19150]_ , \new_[19154]_ ,
    \new_[19155]_ , \new_[19158]_ , \new_[19161]_ , \new_[19162]_ ,
    \new_[19163]_ , \new_[19167]_ , \new_[19168]_ , \new_[19172]_ ,
    \new_[19173]_ , \new_[19174]_ , \new_[19178]_ , \new_[19179]_ ,
    \new_[19182]_ , \new_[19185]_ , \new_[19186]_ , \new_[19187]_ ,
    \new_[19191]_ , \new_[19192]_ , \new_[19196]_ , \new_[19197]_ ,
    \new_[19198]_ , \new_[19202]_ , \new_[19203]_ , \new_[19206]_ ,
    \new_[19209]_ , \new_[19210]_ , \new_[19211]_ , \new_[19215]_ ,
    \new_[19216]_ , \new_[19220]_ , \new_[19221]_ , \new_[19222]_ ,
    \new_[19226]_ , \new_[19227]_ , \new_[19230]_ , \new_[19233]_ ,
    \new_[19234]_ , \new_[19235]_ , \new_[19239]_ , \new_[19240]_ ,
    \new_[19244]_ , \new_[19245]_ , \new_[19246]_ , \new_[19250]_ ,
    \new_[19251]_ , \new_[19254]_ , \new_[19257]_ , \new_[19258]_ ,
    \new_[19259]_ , \new_[19263]_ , \new_[19264]_ , \new_[19268]_ ,
    \new_[19269]_ , \new_[19270]_ , \new_[19274]_ , \new_[19275]_ ,
    \new_[19278]_ , \new_[19281]_ , \new_[19282]_ , \new_[19283]_ ,
    \new_[19287]_ , \new_[19288]_ , \new_[19292]_ , \new_[19293]_ ,
    \new_[19294]_ , \new_[19298]_ , \new_[19299]_ , \new_[19302]_ ,
    \new_[19305]_ , \new_[19306]_ , \new_[19307]_ , \new_[19311]_ ,
    \new_[19312]_ , \new_[19316]_ , \new_[19317]_ , \new_[19318]_ ,
    \new_[19322]_ , \new_[19323]_ , \new_[19326]_ , \new_[19329]_ ,
    \new_[19330]_ , \new_[19331]_ , \new_[19335]_ , \new_[19336]_ ,
    \new_[19340]_ , \new_[19341]_ , \new_[19342]_ , \new_[19346]_ ,
    \new_[19347]_ , \new_[19350]_ , \new_[19353]_ , \new_[19354]_ ,
    \new_[19355]_ , \new_[19359]_ , \new_[19360]_ , \new_[19364]_ ,
    \new_[19365]_ , \new_[19366]_ , \new_[19370]_ , \new_[19371]_ ,
    \new_[19374]_ , \new_[19377]_ , \new_[19378]_ , \new_[19379]_ ,
    \new_[19383]_ , \new_[19384]_ , \new_[19388]_ , \new_[19389]_ ,
    \new_[19390]_ , \new_[19394]_ , \new_[19395]_ , \new_[19398]_ ,
    \new_[19401]_ , \new_[19402]_ , \new_[19403]_ , \new_[19407]_ ,
    \new_[19408]_ , \new_[19412]_ , \new_[19413]_ , \new_[19414]_ ,
    \new_[19418]_ , \new_[19419]_ , \new_[19422]_ , \new_[19425]_ ,
    \new_[19426]_ , \new_[19427]_ , \new_[19431]_ , \new_[19432]_ ,
    \new_[19436]_ , \new_[19437]_ , \new_[19438]_ , \new_[19442]_ ,
    \new_[19443]_ , \new_[19446]_ , \new_[19449]_ , \new_[19450]_ ,
    \new_[19451]_ , \new_[19455]_ , \new_[19456]_ , \new_[19460]_ ,
    \new_[19461]_ , \new_[19462]_ , \new_[19466]_ , \new_[19467]_ ,
    \new_[19470]_ , \new_[19473]_ , \new_[19474]_ , \new_[19475]_ ,
    \new_[19479]_ , \new_[19480]_ , \new_[19484]_ , \new_[19485]_ ,
    \new_[19486]_ , \new_[19490]_ , \new_[19491]_ , \new_[19494]_ ,
    \new_[19497]_ , \new_[19498]_ , \new_[19499]_ , \new_[19503]_ ,
    \new_[19504]_ , \new_[19508]_ , \new_[19509]_ , \new_[19510]_ ,
    \new_[19514]_ , \new_[19515]_ , \new_[19518]_ , \new_[19521]_ ,
    \new_[19522]_ , \new_[19523]_ , \new_[19527]_ , \new_[19528]_ ,
    \new_[19532]_ , \new_[19533]_ , \new_[19534]_ , \new_[19538]_ ,
    \new_[19539]_ , \new_[19542]_ , \new_[19545]_ , \new_[19546]_ ,
    \new_[19547]_ , \new_[19551]_ , \new_[19552]_ , \new_[19556]_ ,
    \new_[19557]_ , \new_[19558]_ , \new_[19562]_ , \new_[19563]_ ,
    \new_[19566]_ , \new_[19569]_ , \new_[19570]_ , \new_[19571]_ ,
    \new_[19575]_ , \new_[19576]_ , \new_[19580]_ , \new_[19581]_ ,
    \new_[19582]_ , \new_[19586]_ , \new_[19587]_ , \new_[19590]_ ,
    \new_[19593]_ , \new_[19594]_ , \new_[19595]_ , \new_[19599]_ ,
    \new_[19600]_ , \new_[19604]_ , \new_[19605]_ , \new_[19606]_ ,
    \new_[19610]_ , \new_[19611]_ , \new_[19614]_ , \new_[19617]_ ,
    \new_[19618]_ , \new_[19619]_ , \new_[19623]_ , \new_[19624]_ ,
    \new_[19628]_ , \new_[19629]_ , \new_[19630]_ , \new_[19634]_ ,
    \new_[19635]_ , \new_[19638]_ , \new_[19641]_ , \new_[19642]_ ,
    \new_[19643]_ , \new_[19647]_ , \new_[19648]_ , \new_[19652]_ ,
    \new_[19653]_ , \new_[19654]_ , \new_[19658]_ , \new_[19659]_ ,
    \new_[19662]_ , \new_[19665]_ , \new_[19666]_ , \new_[19667]_ ,
    \new_[19671]_ , \new_[19672]_ , \new_[19676]_ , \new_[19677]_ ,
    \new_[19678]_ , \new_[19682]_ , \new_[19683]_ , \new_[19686]_ ,
    \new_[19689]_ , \new_[19690]_ , \new_[19691]_ , \new_[19695]_ ,
    \new_[19696]_ , \new_[19700]_ , \new_[19701]_ , \new_[19702]_ ,
    \new_[19706]_ , \new_[19707]_ , \new_[19710]_ , \new_[19713]_ ,
    \new_[19714]_ , \new_[19715]_ , \new_[19719]_ , \new_[19720]_ ,
    \new_[19724]_ , \new_[19725]_ , \new_[19726]_ , \new_[19730]_ ,
    \new_[19731]_ , \new_[19734]_ , \new_[19737]_ , \new_[19738]_ ,
    \new_[19739]_ , \new_[19743]_ , \new_[19744]_ , \new_[19748]_ ,
    \new_[19749]_ , \new_[19750]_ , \new_[19754]_ , \new_[19755]_ ,
    \new_[19758]_ , \new_[19761]_ , \new_[19762]_ , \new_[19763]_ ,
    \new_[19767]_ , \new_[19768]_ , \new_[19772]_ , \new_[19773]_ ,
    \new_[19774]_ , \new_[19778]_ , \new_[19779]_ , \new_[19782]_ ,
    \new_[19785]_ , \new_[19786]_ , \new_[19787]_ , \new_[19791]_ ,
    \new_[19792]_ , \new_[19796]_ , \new_[19797]_ , \new_[19798]_ ,
    \new_[19802]_ , \new_[19803]_ , \new_[19806]_ , \new_[19809]_ ,
    \new_[19810]_ , \new_[19811]_ , \new_[19815]_ , \new_[19816]_ ,
    \new_[19820]_ , \new_[19821]_ , \new_[19822]_ , \new_[19826]_ ,
    \new_[19827]_ , \new_[19830]_ , \new_[19833]_ , \new_[19834]_ ,
    \new_[19835]_ , \new_[19839]_ , \new_[19840]_ , \new_[19844]_ ,
    \new_[19845]_ , \new_[19846]_ , \new_[19850]_ , \new_[19851]_ ,
    \new_[19854]_ , \new_[19857]_ , \new_[19858]_ , \new_[19859]_ ,
    \new_[19863]_ , \new_[19864]_ , \new_[19868]_ , \new_[19869]_ ,
    \new_[19870]_ , \new_[19874]_ , \new_[19875]_ , \new_[19878]_ ,
    \new_[19881]_ , \new_[19882]_ , \new_[19883]_ , \new_[19887]_ ,
    \new_[19888]_ , \new_[19892]_ , \new_[19893]_ , \new_[19894]_ ,
    \new_[19898]_ , \new_[19899]_ , \new_[19902]_ , \new_[19905]_ ,
    \new_[19906]_ , \new_[19907]_ , \new_[19911]_ , \new_[19912]_ ,
    \new_[19916]_ , \new_[19917]_ , \new_[19918]_ , \new_[19922]_ ,
    \new_[19923]_ , \new_[19926]_ , \new_[19929]_ , \new_[19930]_ ,
    \new_[19931]_ , \new_[19935]_ , \new_[19936]_ , \new_[19940]_ ,
    \new_[19941]_ , \new_[19942]_ , \new_[19946]_ , \new_[19947]_ ,
    \new_[19950]_ , \new_[19953]_ , \new_[19954]_ , \new_[19955]_ ,
    \new_[19959]_ , \new_[19960]_ , \new_[19964]_ , \new_[19965]_ ,
    \new_[19966]_ , \new_[19970]_ , \new_[19971]_ , \new_[19974]_ ,
    \new_[19977]_ , \new_[19978]_ , \new_[19979]_ , \new_[19983]_ ,
    \new_[19984]_ , \new_[19988]_ , \new_[19989]_ , \new_[19990]_ ,
    \new_[19994]_ , \new_[19995]_ , \new_[19998]_ , \new_[20001]_ ,
    \new_[20002]_ , \new_[20003]_ , \new_[20007]_ , \new_[20008]_ ,
    \new_[20012]_ , \new_[20013]_ , \new_[20014]_ , \new_[20018]_ ,
    \new_[20019]_ , \new_[20022]_ , \new_[20025]_ , \new_[20026]_ ,
    \new_[20027]_ , \new_[20031]_ , \new_[20032]_ , \new_[20036]_ ,
    \new_[20037]_ , \new_[20038]_ , \new_[20042]_ , \new_[20043]_ ,
    \new_[20046]_ , \new_[20049]_ , \new_[20050]_ , \new_[20051]_ ,
    \new_[20055]_ , \new_[20056]_ , \new_[20060]_ , \new_[20061]_ ,
    \new_[20062]_ , \new_[20066]_ , \new_[20067]_ , \new_[20070]_ ,
    \new_[20073]_ , \new_[20074]_ , \new_[20075]_ , \new_[20079]_ ,
    \new_[20080]_ , \new_[20084]_ , \new_[20085]_ , \new_[20086]_ ,
    \new_[20090]_ , \new_[20091]_ , \new_[20094]_ , \new_[20097]_ ,
    \new_[20098]_ , \new_[20099]_ , \new_[20103]_ , \new_[20104]_ ,
    \new_[20108]_ , \new_[20109]_ , \new_[20110]_ , \new_[20114]_ ,
    \new_[20115]_ , \new_[20118]_ , \new_[20121]_ , \new_[20122]_ ,
    \new_[20123]_ , \new_[20127]_ , \new_[20128]_ , \new_[20132]_ ,
    \new_[20133]_ , \new_[20134]_ , \new_[20138]_ , \new_[20139]_ ,
    \new_[20142]_ , \new_[20145]_ , \new_[20146]_ , \new_[20147]_ ,
    \new_[20151]_ , \new_[20152]_ , \new_[20156]_ , \new_[20157]_ ,
    \new_[20158]_ , \new_[20162]_ , \new_[20163]_ , \new_[20166]_ ,
    \new_[20169]_ , \new_[20170]_ , \new_[20171]_ , \new_[20175]_ ,
    \new_[20176]_ , \new_[20180]_ , \new_[20181]_ , \new_[20182]_ ,
    \new_[20186]_ , \new_[20187]_ , \new_[20190]_ , \new_[20193]_ ,
    \new_[20194]_ , \new_[20195]_ , \new_[20199]_ , \new_[20200]_ ,
    \new_[20204]_ , \new_[20205]_ , \new_[20206]_ , \new_[20210]_ ,
    \new_[20211]_ , \new_[20214]_ , \new_[20217]_ , \new_[20218]_ ,
    \new_[20219]_ , \new_[20223]_ , \new_[20224]_ , \new_[20228]_ ,
    \new_[20229]_ , \new_[20230]_ , \new_[20234]_ , \new_[20235]_ ,
    \new_[20238]_ , \new_[20241]_ , \new_[20242]_ , \new_[20243]_ ,
    \new_[20247]_ , \new_[20248]_ , \new_[20252]_ , \new_[20253]_ ,
    \new_[20254]_ , \new_[20258]_ , \new_[20259]_ , \new_[20262]_ ,
    \new_[20265]_ , \new_[20266]_ , \new_[20267]_ , \new_[20271]_ ,
    \new_[20272]_ , \new_[20276]_ , \new_[20277]_ , \new_[20278]_ ,
    \new_[20282]_ , \new_[20283]_ , \new_[20286]_ , \new_[20289]_ ,
    \new_[20290]_ , \new_[20291]_ , \new_[20295]_ , \new_[20296]_ ,
    \new_[20300]_ , \new_[20301]_ , \new_[20302]_ , \new_[20306]_ ,
    \new_[20307]_ , \new_[20310]_ , \new_[20313]_ , \new_[20314]_ ,
    \new_[20315]_ , \new_[20319]_ , \new_[20320]_ , \new_[20324]_ ,
    \new_[20325]_ , \new_[20326]_ , \new_[20330]_ , \new_[20331]_ ,
    \new_[20334]_ , \new_[20337]_ , \new_[20338]_ , \new_[20339]_ ,
    \new_[20343]_ , \new_[20344]_ , \new_[20348]_ , \new_[20349]_ ,
    \new_[20350]_ , \new_[20354]_ , \new_[20355]_ , \new_[20358]_ ,
    \new_[20361]_ , \new_[20362]_ , \new_[20363]_ , \new_[20367]_ ,
    \new_[20368]_ , \new_[20372]_ , \new_[20373]_ , \new_[20374]_ ,
    \new_[20378]_ , \new_[20379]_ , \new_[20382]_ , \new_[20385]_ ,
    \new_[20386]_ , \new_[20387]_ , \new_[20391]_ , \new_[20392]_ ,
    \new_[20396]_ , \new_[20397]_ , \new_[20398]_ , \new_[20402]_ ,
    \new_[20403]_ , \new_[20406]_ , \new_[20409]_ , \new_[20410]_ ,
    \new_[20411]_ , \new_[20415]_ , \new_[20416]_ , \new_[20420]_ ,
    \new_[20421]_ , \new_[20422]_ , \new_[20426]_ , \new_[20427]_ ,
    \new_[20430]_ , \new_[20433]_ , \new_[20434]_ , \new_[20435]_ ,
    \new_[20439]_ , \new_[20440]_ , \new_[20444]_ , \new_[20445]_ ,
    \new_[20446]_ , \new_[20450]_ , \new_[20451]_ , \new_[20454]_ ,
    \new_[20457]_ , \new_[20458]_ , \new_[20459]_ , \new_[20463]_ ,
    \new_[20464]_ , \new_[20468]_ , \new_[20469]_ , \new_[20470]_ ,
    \new_[20474]_ , \new_[20475]_ , \new_[20478]_ , \new_[20481]_ ,
    \new_[20482]_ , \new_[20483]_ , \new_[20487]_ , \new_[20488]_ ,
    \new_[20492]_ , \new_[20493]_ , \new_[20494]_ , \new_[20498]_ ,
    \new_[20499]_ , \new_[20502]_ , \new_[20505]_ , \new_[20506]_ ,
    \new_[20507]_ , \new_[20511]_ , \new_[20512]_ , \new_[20516]_ ,
    \new_[20517]_ , \new_[20518]_ , \new_[20522]_ , \new_[20523]_ ,
    \new_[20526]_ , \new_[20529]_ , \new_[20530]_ , \new_[20531]_ ,
    \new_[20535]_ , \new_[20536]_ , \new_[20540]_ , \new_[20541]_ ,
    \new_[20542]_ , \new_[20546]_ , \new_[20547]_ , \new_[20550]_ ,
    \new_[20553]_ , \new_[20554]_ , \new_[20555]_ , \new_[20559]_ ,
    \new_[20560]_ , \new_[20564]_ , \new_[20565]_ , \new_[20566]_ ,
    \new_[20570]_ , \new_[20571]_ , \new_[20574]_ , \new_[20577]_ ,
    \new_[20578]_ , \new_[20579]_ , \new_[20583]_ , \new_[20584]_ ,
    \new_[20588]_ , \new_[20589]_ , \new_[20590]_ , \new_[20594]_ ,
    \new_[20595]_ , \new_[20598]_ , \new_[20601]_ , \new_[20602]_ ,
    \new_[20603]_ , \new_[20607]_ , \new_[20608]_ , \new_[20612]_ ,
    \new_[20613]_ , \new_[20614]_ , \new_[20618]_ , \new_[20619]_ ,
    \new_[20622]_ , \new_[20625]_ , \new_[20626]_ , \new_[20627]_ ,
    \new_[20631]_ , \new_[20632]_ , \new_[20636]_ , \new_[20637]_ ,
    \new_[20638]_ , \new_[20642]_ , \new_[20643]_ , \new_[20646]_ ,
    \new_[20649]_ , \new_[20650]_ , \new_[20651]_ , \new_[20655]_ ,
    \new_[20656]_ , \new_[20660]_ , \new_[20661]_ , \new_[20662]_ ,
    \new_[20666]_ , \new_[20667]_ , \new_[20670]_ , \new_[20673]_ ,
    \new_[20674]_ , \new_[20675]_ , \new_[20679]_ , \new_[20680]_ ,
    \new_[20684]_ , \new_[20685]_ , \new_[20686]_ , \new_[20690]_ ,
    \new_[20691]_ , \new_[20694]_ , \new_[20697]_ , \new_[20698]_ ,
    \new_[20699]_ , \new_[20703]_ , \new_[20704]_ , \new_[20708]_ ,
    \new_[20709]_ , \new_[20710]_ , \new_[20714]_ , \new_[20715]_ ,
    \new_[20718]_ , \new_[20721]_ , \new_[20722]_ , \new_[20723]_ ,
    \new_[20727]_ , \new_[20728]_ , \new_[20732]_ , \new_[20733]_ ,
    \new_[20734]_ , \new_[20738]_ , \new_[20739]_ , \new_[20742]_ ,
    \new_[20745]_ , \new_[20746]_ , \new_[20747]_ , \new_[20751]_ ,
    \new_[20752]_ , \new_[20756]_ , \new_[20757]_ , \new_[20758]_ ,
    \new_[20762]_ , \new_[20763]_ , \new_[20766]_ , \new_[20769]_ ,
    \new_[20770]_ , \new_[20771]_ , \new_[20775]_ , \new_[20776]_ ,
    \new_[20780]_ , \new_[20781]_ , \new_[20782]_ , \new_[20786]_ ,
    \new_[20787]_ , \new_[20790]_ , \new_[20793]_ , \new_[20794]_ ,
    \new_[20795]_ , \new_[20799]_ , \new_[20800]_ , \new_[20804]_ ,
    \new_[20805]_ , \new_[20806]_ , \new_[20810]_ , \new_[20811]_ ,
    \new_[20814]_ , \new_[20817]_ , \new_[20818]_ , \new_[20819]_ ,
    \new_[20823]_ , \new_[20824]_ , \new_[20828]_ , \new_[20829]_ ,
    \new_[20830]_ , \new_[20834]_ , \new_[20835]_ , \new_[20838]_ ,
    \new_[20841]_ , \new_[20842]_ , \new_[20843]_ , \new_[20847]_ ,
    \new_[20848]_ , \new_[20852]_ , \new_[20853]_ , \new_[20854]_ ,
    \new_[20858]_ , \new_[20859]_ , \new_[20862]_ , \new_[20865]_ ,
    \new_[20866]_ , \new_[20867]_ , \new_[20871]_ , \new_[20872]_ ,
    \new_[20876]_ , \new_[20877]_ , \new_[20878]_ , \new_[20882]_ ,
    \new_[20883]_ , \new_[20886]_ , \new_[20889]_ , \new_[20890]_ ,
    \new_[20891]_ , \new_[20895]_ , \new_[20896]_ , \new_[20900]_ ,
    \new_[20901]_ , \new_[20902]_ , \new_[20906]_ , \new_[20907]_ ,
    \new_[20910]_ , \new_[20913]_ , \new_[20914]_ , \new_[20915]_ ,
    \new_[20919]_ , \new_[20920]_ , \new_[20924]_ , \new_[20925]_ ,
    \new_[20926]_ , \new_[20930]_ , \new_[20931]_ , \new_[20934]_ ,
    \new_[20937]_ , \new_[20938]_ , \new_[20939]_ , \new_[20943]_ ,
    \new_[20944]_ , \new_[20948]_ , \new_[20949]_ , \new_[20950]_ ,
    \new_[20954]_ , \new_[20955]_ , \new_[20958]_ , \new_[20961]_ ,
    \new_[20962]_ , \new_[20963]_ , \new_[20967]_ , \new_[20968]_ ,
    \new_[20972]_ , \new_[20973]_ , \new_[20974]_ , \new_[20978]_ ,
    \new_[20979]_ , \new_[20982]_ , \new_[20985]_ , \new_[20986]_ ,
    \new_[20987]_ , \new_[20991]_ , \new_[20992]_ , \new_[20996]_ ,
    \new_[20997]_ , \new_[20998]_ , \new_[21002]_ , \new_[21003]_ ,
    \new_[21006]_ , \new_[21009]_ , \new_[21010]_ , \new_[21011]_ ,
    \new_[21015]_ , \new_[21016]_ , \new_[21020]_ , \new_[21021]_ ,
    \new_[21022]_ , \new_[21026]_ , \new_[21027]_ , \new_[21030]_ ,
    \new_[21033]_ , \new_[21034]_ , \new_[21035]_ , \new_[21039]_ ,
    \new_[21040]_ , \new_[21044]_ , \new_[21045]_ , \new_[21046]_ ,
    \new_[21050]_ , \new_[21051]_ , \new_[21054]_ , \new_[21057]_ ,
    \new_[21058]_ , \new_[21059]_ , \new_[21063]_ , \new_[21064]_ ,
    \new_[21068]_ , \new_[21069]_ , \new_[21070]_ , \new_[21074]_ ,
    \new_[21075]_ , \new_[21078]_ , \new_[21081]_ , \new_[21082]_ ,
    \new_[21083]_ , \new_[21087]_ , \new_[21088]_ , \new_[21092]_ ,
    \new_[21093]_ , \new_[21094]_ , \new_[21098]_ , \new_[21099]_ ,
    \new_[21102]_ , \new_[21105]_ , \new_[21106]_ , \new_[21107]_ ,
    \new_[21111]_ , \new_[21112]_ , \new_[21116]_ , \new_[21117]_ ,
    \new_[21118]_ , \new_[21122]_ , \new_[21123]_ , \new_[21126]_ ,
    \new_[21129]_ , \new_[21130]_ , \new_[21131]_ , \new_[21135]_ ,
    \new_[21136]_ , \new_[21140]_ , \new_[21141]_ , \new_[21142]_ ,
    \new_[21146]_ , \new_[21147]_ , \new_[21150]_ , \new_[21153]_ ,
    \new_[21154]_ , \new_[21155]_ , \new_[21159]_ , \new_[21160]_ ,
    \new_[21164]_ , \new_[21165]_ , \new_[21166]_ , \new_[21170]_ ,
    \new_[21171]_ , \new_[21174]_ , \new_[21177]_ , \new_[21178]_ ,
    \new_[21179]_ , \new_[21183]_ , \new_[21184]_ , \new_[21188]_ ,
    \new_[21189]_ , \new_[21190]_ , \new_[21194]_ , \new_[21195]_ ,
    \new_[21198]_ , \new_[21201]_ , \new_[21202]_ , \new_[21203]_ ,
    \new_[21207]_ , \new_[21208]_ , \new_[21212]_ , \new_[21213]_ ,
    \new_[21214]_ , \new_[21218]_ , \new_[21219]_ , \new_[21222]_ ,
    \new_[21225]_ , \new_[21226]_ , \new_[21227]_ , \new_[21231]_ ,
    \new_[21232]_ , \new_[21236]_ , \new_[21237]_ , \new_[21238]_ ,
    \new_[21242]_ , \new_[21243]_ , \new_[21246]_ , \new_[21249]_ ,
    \new_[21250]_ , \new_[21251]_ , \new_[21255]_ , \new_[21256]_ ,
    \new_[21260]_ , \new_[21261]_ , \new_[21262]_ , \new_[21266]_ ,
    \new_[21267]_ , \new_[21270]_ , \new_[21273]_ , \new_[21274]_ ,
    \new_[21275]_ , \new_[21279]_ , \new_[21280]_ , \new_[21284]_ ,
    \new_[21285]_ , \new_[21286]_ , \new_[21290]_ , \new_[21291]_ ,
    \new_[21294]_ , \new_[21297]_ , \new_[21298]_ , \new_[21299]_ ,
    \new_[21303]_ , \new_[21304]_ , \new_[21308]_ , \new_[21309]_ ,
    \new_[21310]_ , \new_[21314]_ , \new_[21315]_ , \new_[21318]_ ,
    \new_[21321]_ , \new_[21322]_ , \new_[21323]_ , \new_[21327]_ ,
    \new_[21328]_ , \new_[21332]_ , \new_[21333]_ , \new_[21334]_ ,
    \new_[21338]_ , \new_[21339]_ , \new_[21342]_ , \new_[21345]_ ,
    \new_[21346]_ , \new_[21347]_ , \new_[21351]_ , \new_[21352]_ ,
    \new_[21356]_ , \new_[21357]_ , \new_[21358]_ , \new_[21362]_ ,
    \new_[21363]_ , \new_[21366]_ , \new_[21369]_ , \new_[21370]_ ,
    \new_[21371]_ , \new_[21375]_ , \new_[21376]_ , \new_[21380]_ ,
    \new_[21381]_ , \new_[21382]_ , \new_[21386]_ , \new_[21387]_ ,
    \new_[21390]_ , \new_[21393]_ , \new_[21394]_ , \new_[21395]_ ,
    \new_[21399]_ , \new_[21400]_ , \new_[21404]_ , \new_[21405]_ ,
    \new_[21406]_ , \new_[21410]_ , \new_[21411]_ , \new_[21414]_ ,
    \new_[21417]_ , \new_[21418]_ , \new_[21419]_ , \new_[21423]_ ,
    \new_[21424]_ , \new_[21428]_ , \new_[21429]_ , \new_[21430]_ ,
    \new_[21434]_ , \new_[21435]_ , \new_[21438]_ , \new_[21441]_ ,
    \new_[21442]_ , \new_[21443]_ , \new_[21447]_ , \new_[21448]_ ,
    \new_[21452]_ , \new_[21453]_ , \new_[21454]_ , \new_[21458]_ ,
    \new_[21459]_ , \new_[21462]_ , \new_[21465]_ , \new_[21466]_ ,
    \new_[21467]_ , \new_[21471]_ , \new_[21472]_ , \new_[21476]_ ,
    \new_[21477]_ , \new_[21478]_ , \new_[21482]_ , \new_[21483]_ ,
    \new_[21486]_ , \new_[21489]_ , \new_[21490]_ , \new_[21491]_ ,
    \new_[21495]_ , \new_[21496]_ , \new_[21500]_ , \new_[21501]_ ,
    \new_[21502]_ , \new_[21506]_ , \new_[21507]_ , \new_[21510]_ ,
    \new_[21513]_ , \new_[21514]_ , \new_[21515]_ , \new_[21519]_ ,
    \new_[21520]_ , \new_[21524]_ , \new_[21525]_ , \new_[21526]_ ,
    \new_[21530]_ , \new_[21531]_ , \new_[21534]_ , \new_[21537]_ ,
    \new_[21538]_ , \new_[21539]_ , \new_[21543]_ , \new_[21544]_ ,
    \new_[21548]_ , \new_[21549]_ , \new_[21550]_ , \new_[21554]_ ,
    \new_[21555]_ , \new_[21558]_ , \new_[21561]_ , \new_[21562]_ ,
    \new_[21563]_ , \new_[21567]_ , \new_[21568]_ , \new_[21572]_ ,
    \new_[21573]_ , \new_[21574]_ , \new_[21578]_ , \new_[21579]_ ,
    \new_[21582]_ , \new_[21585]_ , \new_[21586]_ , \new_[21587]_ ,
    \new_[21591]_ , \new_[21592]_ , \new_[21596]_ , \new_[21597]_ ,
    \new_[21598]_ , \new_[21602]_ , \new_[21603]_ , \new_[21606]_ ,
    \new_[21609]_ , \new_[21610]_ , \new_[21611]_ , \new_[21615]_ ,
    \new_[21616]_ , \new_[21620]_ , \new_[21621]_ , \new_[21622]_ ,
    \new_[21626]_ , \new_[21627]_ , \new_[21630]_ , \new_[21633]_ ,
    \new_[21634]_ , \new_[21635]_ , \new_[21639]_ , \new_[21640]_ ,
    \new_[21644]_ , \new_[21645]_ , \new_[21646]_ , \new_[21650]_ ,
    \new_[21651]_ , \new_[21654]_ , \new_[21657]_ , \new_[21658]_ ,
    \new_[21659]_ , \new_[21663]_ , \new_[21664]_ , \new_[21668]_ ,
    \new_[21669]_ , \new_[21670]_ , \new_[21674]_ , \new_[21675]_ ,
    \new_[21678]_ , \new_[21681]_ , \new_[21682]_ , \new_[21683]_ ,
    \new_[21687]_ , \new_[21688]_ , \new_[21692]_ , \new_[21693]_ ,
    \new_[21694]_ , \new_[21698]_ , \new_[21699]_ , \new_[21702]_ ,
    \new_[21705]_ , \new_[21706]_ , \new_[21707]_ , \new_[21711]_ ,
    \new_[21712]_ , \new_[21716]_ , \new_[21717]_ , \new_[21718]_ ,
    \new_[21722]_ , \new_[21723]_ , \new_[21726]_ , \new_[21729]_ ,
    \new_[21730]_ , \new_[21731]_ , \new_[21735]_ , \new_[21736]_ ,
    \new_[21740]_ , \new_[21741]_ , \new_[21742]_ , \new_[21746]_ ,
    \new_[21747]_ , \new_[21750]_ , \new_[21753]_ , \new_[21754]_ ,
    \new_[21755]_ , \new_[21759]_ , \new_[21760]_ , \new_[21764]_ ,
    \new_[21765]_ , \new_[21766]_ , \new_[21770]_ , \new_[21771]_ ,
    \new_[21774]_ , \new_[21777]_ , \new_[21778]_ , \new_[21779]_ ,
    \new_[21783]_ , \new_[21784]_ , \new_[21788]_ , \new_[21789]_ ,
    \new_[21790]_ , \new_[21794]_ , \new_[21795]_ , \new_[21798]_ ,
    \new_[21801]_ , \new_[21802]_ , \new_[21803]_ , \new_[21807]_ ,
    \new_[21808]_ , \new_[21812]_ , \new_[21813]_ , \new_[21814]_ ,
    \new_[21818]_ , \new_[21819]_ , \new_[21822]_ , \new_[21825]_ ,
    \new_[21826]_ , \new_[21827]_ , \new_[21831]_ , \new_[21832]_ ,
    \new_[21836]_ , \new_[21837]_ , \new_[21838]_ , \new_[21842]_ ,
    \new_[21843]_ , \new_[21846]_ , \new_[21849]_ , \new_[21850]_ ,
    \new_[21851]_ , \new_[21855]_ , \new_[21856]_ , \new_[21860]_ ,
    \new_[21861]_ , \new_[21862]_ , \new_[21866]_ , \new_[21867]_ ,
    \new_[21870]_ , \new_[21873]_ , \new_[21874]_ , \new_[21875]_ ,
    \new_[21879]_ , \new_[21880]_ , \new_[21884]_ , \new_[21885]_ ,
    \new_[21886]_ , \new_[21890]_ , \new_[21891]_ , \new_[21894]_ ,
    \new_[21897]_ , \new_[21898]_ , \new_[21899]_ , \new_[21903]_ ,
    \new_[21904]_ , \new_[21908]_ , \new_[21909]_ , \new_[21910]_ ,
    \new_[21914]_ , \new_[21915]_ , \new_[21918]_ , \new_[21921]_ ,
    \new_[21922]_ , \new_[21923]_ , \new_[21927]_ , \new_[21928]_ ,
    \new_[21932]_ , \new_[21933]_ , \new_[21934]_ , \new_[21938]_ ,
    \new_[21939]_ , \new_[21942]_ , \new_[21945]_ , \new_[21946]_ ,
    \new_[21947]_ , \new_[21951]_ , \new_[21952]_ , \new_[21956]_ ,
    \new_[21957]_ , \new_[21958]_ , \new_[21962]_ , \new_[21963]_ ,
    \new_[21966]_ , \new_[21969]_ , \new_[21970]_ , \new_[21971]_ ,
    \new_[21975]_ , \new_[21976]_ , \new_[21980]_ , \new_[21981]_ ,
    \new_[21982]_ , \new_[21986]_ , \new_[21987]_ , \new_[21990]_ ,
    \new_[21993]_ , \new_[21994]_ , \new_[21995]_ , \new_[21999]_ ,
    \new_[22000]_ , \new_[22004]_ , \new_[22005]_ , \new_[22006]_ ,
    \new_[22010]_ , \new_[22011]_ , \new_[22014]_ , \new_[22017]_ ,
    \new_[22018]_ , \new_[22019]_ , \new_[22023]_ , \new_[22024]_ ,
    \new_[22028]_ , \new_[22029]_ , \new_[22030]_ , \new_[22034]_ ,
    \new_[22035]_ , \new_[22038]_ , \new_[22041]_ , \new_[22042]_ ,
    \new_[22043]_ , \new_[22047]_ , \new_[22048]_ , \new_[22052]_ ,
    \new_[22053]_ , \new_[22054]_ , \new_[22058]_ , \new_[22059]_ ,
    \new_[22062]_ , \new_[22065]_ , \new_[22066]_ , \new_[22067]_ ,
    \new_[22071]_ , \new_[22072]_ , \new_[22076]_ , \new_[22077]_ ,
    \new_[22078]_ , \new_[22082]_ , \new_[22083]_ , \new_[22086]_ ,
    \new_[22089]_ , \new_[22090]_ , \new_[22091]_ , \new_[22095]_ ,
    \new_[22096]_ , \new_[22100]_ , \new_[22101]_ , \new_[22102]_ ,
    \new_[22106]_ , \new_[22107]_ , \new_[22110]_ , \new_[22113]_ ,
    \new_[22114]_ , \new_[22115]_ , \new_[22119]_ , \new_[22120]_ ,
    \new_[22124]_ , \new_[22125]_ , \new_[22126]_ , \new_[22130]_ ,
    \new_[22131]_ , \new_[22134]_ , \new_[22137]_ , \new_[22138]_ ,
    \new_[22139]_ , \new_[22143]_ , \new_[22144]_ , \new_[22148]_ ,
    \new_[22149]_ , \new_[22150]_ , \new_[22154]_ , \new_[22155]_ ,
    \new_[22158]_ , \new_[22161]_ , \new_[22162]_ , \new_[22163]_ ,
    \new_[22167]_ , \new_[22168]_ , \new_[22172]_ , \new_[22173]_ ,
    \new_[22174]_ , \new_[22178]_ , \new_[22179]_ , \new_[22182]_ ,
    \new_[22185]_ , \new_[22186]_ , \new_[22187]_ , \new_[22191]_ ,
    \new_[22192]_ , \new_[22196]_ , \new_[22197]_ , \new_[22198]_ ,
    \new_[22202]_ , \new_[22203]_ , \new_[22206]_ , \new_[22209]_ ,
    \new_[22210]_ , \new_[22211]_ , \new_[22215]_ , \new_[22216]_ ,
    \new_[22220]_ , \new_[22221]_ , \new_[22222]_ , \new_[22226]_ ,
    \new_[22227]_ , \new_[22230]_ , \new_[22233]_ , \new_[22234]_ ,
    \new_[22235]_ , \new_[22239]_ , \new_[22240]_ , \new_[22244]_ ,
    \new_[22245]_ , \new_[22246]_ , \new_[22250]_ , \new_[22251]_ ,
    \new_[22254]_ , \new_[22257]_ , \new_[22258]_ , \new_[22259]_ ,
    \new_[22263]_ , \new_[22264]_ , \new_[22268]_ , \new_[22269]_ ,
    \new_[22270]_ , \new_[22274]_ , \new_[22275]_ , \new_[22278]_ ,
    \new_[22281]_ , \new_[22282]_ , \new_[22283]_ , \new_[22287]_ ,
    \new_[22288]_ , \new_[22292]_ , \new_[22293]_ , \new_[22294]_ ,
    \new_[22298]_ , \new_[22299]_ , \new_[22302]_ , \new_[22305]_ ,
    \new_[22306]_ , \new_[22307]_ , \new_[22311]_ , \new_[22312]_ ,
    \new_[22316]_ , \new_[22317]_ , \new_[22318]_ , \new_[22322]_ ,
    \new_[22323]_ , \new_[22326]_ , \new_[22329]_ , \new_[22330]_ ,
    \new_[22331]_ , \new_[22335]_ , \new_[22336]_ , \new_[22340]_ ,
    \new_[22341]_ , \new_[22342]_ , \new_[22346]_ , \new_[22347]_ ,
    \new_[22350]_ , \new_[22353]_ , \new_[22354]_ , \new_[22355]_ ,
    \new_[22359]_ , \new_[22360]_ , \new_[22364]_ , \new_[22365]_ ,
    \new_[22366]_ , \new_[22370]_ , \new_[22371]_ , \new_[22374]_ ,
    \new_[22377]_ , \new_[22378]_ , \new_[22379]_ , \new_[22383]_ ,
    \new_[22384]_ , \new_[22388]_ , \new_[22389]_ , \new_[22390]_ ,
    \new_[22394]_ , \new_[22395]_ , \new_[22398]_ , \new_[22401]_ ,
    \new_[22402]_ , \new_[22403]_ , \new_[22407]_ , \new_[22408]_ ,
    \new_[22412]_ , \new_[22413]_ , \new_[22414]_ , \new_[22418]_ ,
    \new_[22419]_ , \new_[22422]_ , \new_[22425]_ , \new_[22426]_ ,
    \new_[22427]_ , \new_[22431]_ , \new_[22432]_ , \new_[22436]_ ,
    \new_[22437]_ , \new_[22438]_ , \new_[22442]_ , \new_[22443]_ ,
    \new_[22446]_ , \new_[22449]_ , \new_[22450]_ , \new_[22451]_ ,
    \new_[22455]_ , \new_[22456]_ , \new_[22460]_ , \new_[22461]_ ,
    \new_[22462]_ , \new_[22466]_ , \new_[22467]_ , \new_[22470]_ ,
    \new_[22473]_ , \new_[22474]_ , \new_[22475]_ , \new_[22479]_ ,
    \new_[22480]_ , \new_[22484]_ , \new_[22485]_ , \new_[22486]_ ,
    \new_[22490]_ , \new_[22491]_ , \new_[22494]_ , \new_[22497]_ ,
    \new_[22498]_ , \new_[22499]_ , \new_[22503]_ , \new_[22504]_ ,
    \new_[22508]_ , \new_[22509]_ , \new_[22510]_ , \new_[22514]_ ,
    \new_[22515]_ , \new_[22518]_ , \new_[22521]_ , \new_[22522]_ ,
    \new_[22523]_ , \new_[22527]_ , \new_[22528]_ , \new_[22532]_ ,
    \new_[22533]_ , \new_[22534]_ , \new_[22538]_ , \new_[22539]_ ,
    \new_[22542]_ , \new_[22545]_ , \new_[22546]_ , \new_[22547]_ ,
    \new_[22551]_ , \new_[22552]_ , \new_[22556]_ , \new_[22557]_ ,
    \new_[22558]_ , \new_[22562]_ , \new_[22563]_ , \new_[22566]_ ,
    \new_[22569]_ , \new_[22570]_ , \new_[22571]_ , \new_[22575]_ ,
    \new_[22576]_ , \new_[22580]_ , \new_[22581]_ , \new_[22582]_ ,
    \new_[22586]_ , \new_[22587]_ , \new_[22590]_ , \new_[22593]_ ,
    \new_[22594]_ , \new_[22595]_ , \new_[22599]_ , \new_[22600]_ ,
    \new_[22604]_ , \new_[22605]_ , \new_[22606]_ , \new_[22610]_ ,
    \new_[22611]_ , \new_[22614]_ , \new_[22617]_ , \new_[22618]_ ,
    \new_[22619]_ , \new_[22623]_ , \new_[22624]_ , \new_[22628]_ ,
    \new_[22629]_ , \new_[22630]_ , \new_[22634]_ , \new_[22635]_ ,
    \new_[22638]_ , \new_[22641]_ , \new_[22642]_ , \new_[22643]_ ,
    \new_[22647]_ , \new_[22648]_ , \new_[22652]_ , \new_[22653]_ ,
    \new_[22654]_ , \new_[22658]_ , \new_[22659]_ , \new_[22662]_ ,
    \new_[22665]_ , \new_[22666]_ , \new_[22667]_ , \new_[22671]_ ,
    \new_[22672]_ , \new_[22676]_ , \new_[22677]_ , \new_[22678]_ ,
    \new_[22682]_ , \new_[22683]_ , \new_[22686]_ , \new_[22689]_ ,
    \new_[22690]_ , \new_[22691]_ , \new_[22695]_ , \new_[22696]_ ,
    \new_[22700]_ , \new_[22701]_ , \new_[22702]_ , \new_[22706]_ ,
    \new_[22707]_ , \new_[22710]_ , \new_[22713]_ , \new_[22714]_ ,
    \new_[22715]_ , \new_[22719]_ , \new_[22720]_ , \new_[22724]_ ,
    \new_[22725]_ , \new_[22726]_ , \new_[22730]_ , \new_[22731]_ ,
    \new_[22734]_ , \new_[22737]_ , \new_[22738]_ , \new_[22739]_ ,
    \new_[22743]_ , \new_[22744]_ , \new_[22748]_ , \new_[22749]_ ,
    \new_[22750]_ , \new_[22754]_ , \new_[22755]_ , \new_[22758]_ ,
    \new_[22761]_ , \new_[22762]_ , \new_[22763]_ , \new_[22767]_ ,
    \new_[22768]_ , \new_[22772]_ , \new_[22773]_ , \new_[22774]_ ,
    \new_[22778]_ , \new_[22779]_ , \new_[22782]_ , \new_[22785]_ ,
    \new_[22786]_ , \new_[22787]_ , \new_[22791]_ , \new_[22792]_ ,
    \new_[22796]_ , \new_[22797]_ , \new_[22798]_ , \new_[22802]_ ,
    \new_[22803]_ , \new_[22806]_ , \new_[22809]_ , \new_[22810]_ ,
    \new_[22811]_ , \new_[22815]_ , \new_[22816]_ , \new_[22820]_ ,
    \new_[22821]_ , \new_[22822]_ , \new_[22826]_ , \new_[22827]_ ,
    \new_[22830]_ , \new_[22833]_ , \new_[22834]_ , \new_[22835]_ ,
    \new_[22839]_ , \new_[22840]_ , \new_[22844]_ , \new_[22845]_ ,
    \new_[22846]_ , \new_[22850]_ , \new_[22851]_ , \new_[22854]_ ,
    \new_[22857]_ , \new_[22858]_ , \new_[22859]_ , \new_[22863]_ ,
    \new_[22864]_ , \new_[22868]_ , \new_[22869]_ , \new_[22870]_ ,
    \new_[22874]_ , \new_[22875]_ , \new_[22878]_ , \new_[22881]_ ,
    \new_[22882]_ , \new_[22883]_ , \new_[22887]_ , \new_[22888]_ ,
    \new_[22892]_ , \new_[22893]_ , \new_[22894]_ , \new_[22898]_ ,
    \new_[22899]_ , \new_[22902]_ , \new_[22905]_ , \new_[22906]_ ,
    \new_[22907]_ , \new_[22911]_ , \new_[22912]_ , \new_[22916]_ ,
    \new_[22917]_ , \new_[22918]_ , \new_[22922]_ , \new_[22923]_ ,
    \new_[22926]_ , \new_[22929]_ , \new_[22930]_ , \new_[22931]_ ,
    \new_[22935]_ , \new_[22936]_ , \new_[22940]_ , \new_[22941]_ ,
    \new_[22942]_ , \new_[22946]_ , \new_[22947]_ , \new_[22950]_ ,
    \new_[22953]_ , \new_[22954]_ , \new_[22955]_ , \new_[22959]_ ,
    \new_[22960]_ , \new_[22964]_ , \new_[22965]_ , \new_[22966]_ ,
    \new_[22970]_ , \new_[22971]_ , \new_[22974]_ , \new_[22977]_ ,
    \new_[22978]_ , \new_[22979]_ , \new_[22983]_ , \new_[22984]_ ,
    \new_[22988]_ , \new_[22989]_ , \new_[22990]_ , \new_[22994]_ ,
    \new_[22995]_ , \new_[22998]_ , \new_[23001]_ , \new_[23002]_ ,
    \new_[23003]_ , \new_[23007]_ , \new_[23008]_ , \new_[23012]_ ,
    \new_[23013]_ , \new_[23014]_ , \new_[23018]_ , \new_[23019]_ ,
    \new_[23022]_ , \new_[23025]_ , \new_[23026]_ , \new_[23027]_ ,
    \new_[23031]_ , \new_[23032]_ , \new_[23036]_ , \new_[23037]_ ,
    \new_[23038]_ , \new_[23042]_ , \new_[23043]_ , \new_[23046]_ ,
    \new_[23049]_ , \new_[23050]_ , \new_[23051]_ , \new_[23055]_ ,
    \new_[23056]_ , \new_[23060]_ , \new_[23061]_ , \new_[23062]_ ,
    \new_[23066]_ , \new_[23067]_ , \new_[23070]_ , \new_[23073]_ ,
    \new_[23074]_ , \new_[23075]_ , \new_[23079]_ , \new_[23080]_ ,
    \new_[23084]_ , \new_[23085]_ , \new_[23086]_ , \new_[23090]_ ,
    \new_[23091]_ , \new_[23094]_ , \new_[23097]_ , \new_[23098]_ ,
    \new_[23099]_ , \new_[23103]_ , \new_[23104]_ , \new_[23108]_ ,
    \new_[23109]_ , \new_[23110]_ , \new_[23114]_ , \new_[23115]_ ,
    \new_[23118]_ , \new_[23121]_ , \new_[23122]_ , \new_[23123]_ ,
    \new_[23127]_ , \new_[23128]_ , \new_[23132]_ , \new_[23133]_ ,
    \new_[23134]_ , \new_[23138]_ , \new_[23139]_ , \new_[23142]_ ,
    \new_[23145]_ , \new_[23146]_ , \new_[23147]_ , \new_[23151]_ ,
    \new_[23152]_ , \new_[23156]_ , \new_[23157]_ , \new_[23158]_ ,
    \new_[23162]_ , \new_[23163]_ , \new_[23166]_ , \new_[23169]_ ,
    \new_[23170]_ , \new_[23171]_ , \new_[23175]_ , \new_[23176]_ ,
    \new_[23180]_ , \new_[23181]_ , \new_[23182]_ , \new_[23186]_ ,
    \new_[23187]_ , \new_[23190]_ , \new_[23193]_ , \new_[23194]_ ,
    \new_[23195]_ , \new_[23199]_ , \new_[23200]_ , \new_[23204]_ ,
    \new_[23205]_ , \new_[23206]_ , \new_[23210]_ , \new_[23211]_ ,
    \new_[23214]_ , \new_[23217]_ , \new_[23218]_ , \new_[23219]_ ,
    \new_[23223]_ , \new_[23224]_ , \new_[23228]_ , \new_[23229]_ ,
    \new_[23230]_ , \new_[23234]_ , \new_[23235]_ , \new_[23238]_ ,
    \new_[23241]_ , \new_[23242]_ , \new_[23243]_ , \new_[23247]_ ,
    \new_[23248]_ , \new_[23251]_ , \new_[23254]_ , \new_[23255]_ ,
    \new_[23256]_ , \new_[23260]_ , \new_[23261]_ , \new_[23264]_ ,
    \new_[23267]_ , \new_[23268]_ , \new_[23269]_ , \new_[23273]_ ,
    \new_[23274]_ , \new_[23277]_ , \new_[23280]_ , \new_[23281]_ ,
    \new_[23282]_ , \new_[23286]_ , \new_[23287]_ , \new_[23290]_ ,
    \new_[23293]_ , \new_[23294]_ , \new_[23295]_ , \new_[23299]_ ,
    \new_[23300]_ , \new_[23303]_ , \new_[23306]_ , \new_[23307]_ ,
    \new_[23308]_ , \new_[23312]_ , \new_[23313]_ , \new_[23316]_ ,
    \new_[23319]_ , \new_[23320]_ , \new_[23321]_ , \new_[23325]_ ,
    \new_[23326]_ , \new_[23329]_ , \new_[23332]_ , \new_[23333]_ ,
    \new_[23334]_ , \new_[23338]_ , \new_[23339]_ , \new_[23342]_ ,
    \new_[23345]_ , \new_[23346]_ , \new_[23347]_ , \new_[23351]_ ,
    \new_[23352]_ , \new_[23355]_ , \new_[23358]_ , \new_[23359]_ ,
    \new_[23360]_ , \new_[23364]_ , \new_[23365]_ , \new_[23368]_ ,
    \new_[23371]_ , \new_[23372]_ , \new_[23373]_ , \new_[23377]_ ,
    \new_[23378]_ , \new_[23381]_ , \new_[23384]_ , \new_[23385]_ ,
    \new_[23386]_ , \new_[23390]_ , \new_[23391]_ , \new_[23394]_ ,
    \new_[23397]_ , \new_[23398]_ , \new_[23399]_ , \new_[23403]_ ,
    \new_[23404]_ , \new_[23407]_ , \new_[23410]_ , \new_[23411]_ ,
    \new_[23412]_ , \new_[23416]_ , \new_[23417]_ , \new_[23420]_ ,
    \new_[23423]_ , \new_[23424]_ , \new_[23425]_ , \new_[23429]_ ,
    \new_[23430]_ , \new_[23433]_ , \new_[23436]_ , \new_[23437]_ ,
    \new_[23438]_ , \new_[23442]_ , \new_[23443]_ , \new_[23446]_ ,
    \new_[23449]_ , \new_[23450]_ , \new_[23451]_ , \new_[23455]_ ,
    \new_[23456]_ , \new_[23459]_ , \new_[23462]_ , \new_[23463]_ ,
    \new_[23464]_ , \new_[23468]_ , \new_[23469]_ , \new_[23472]_ ,
    \new_[23475]_ , \new_[23476]_ , \new_[23477]_ , \new_[23481]_ ,
    \new_[23482]_ , \new_[23485]_ , \new_[23488]_ , \new_[23489]_ ,
    \new_[23490]_ , \new_[23494]_ , \new_[23495]_ , \new_[23498]_ ,
    \new_[23501]_ , \new_[23502]_ , \new_[23503]_ , \new_[23507]_ ,
    \new_[23508]_ , \new_[23511]_ , \new_[23514]_ , \new_[23515]_ ,
    \new_[23516]_ , \new_[23520]_ , \new_[23521]_ , \new_[23524]_ ,
    \new_[23527]_ , \new_[23528]_ , \new_[23529]_ , \new_[23533]_ ,
    \new_[23534]_ , \new_[23537]_ , \new_[23540]_ , \new_[23541]_ ,
    \new_[23542]_ , \new_[23546]_ , \new_[23547]_ , \new_[23550]_ ,
    \new_[23553]_ , \new_[23554]_ , \new_[23555]_ , \new_[23559]_ ,
    \new_[23560]_ , \new_[23563]_ , \new_[23566]_ , \new_[23567]_ ,
    \new_[23568]_ , \new_[23572]_ , \new_[23573]_ , \new_[23576]_ ,
    \new_[23579]_ , \new_[23580]_ , \new_[23581]_ , \new_[23585]_ ,
    \new_[23586]_ , \new_[23589]_ , \new_[23592]_ , \new_[23593]_ ,
    \new_[23594]_ , \new_[23598]_ , \new_[23599]_ , \new_[23602]_ ,
    \new_[23605]_ , \new_[23606]_ , \new_[23607]_ , \new_[23611]_ ,
    \new_[23612]_ , \new_[23615]_ , \new_[23618]_ , \new_[23619]_ ,
    \new_[23620]_ , \new_[23624]_ , \new_[23625]_ , \new_[23628]_ ,
    \new_[23631]_ , \new_[23632]_ , \new_[23633]_ , \new_[23637]_ ,
    \new_[23638]_ , \new_[23641]_ , \new_[23644]_ , \new_[23645]_ ,
    \new_[23646]_ , \new_[23650]_ , \new_[23651]_ , \new_[23654]_ ,
    \new_[23657]_ , \new_[23658]_ , \new_[23659]_ , \new_[23663]_ ,
    \new_[23664]_ , \new_[23667]_ , \new_[23670]_ , \new_[23671]_ ,
    \new_[23672]_ , \new_[23676]_ , \new_[23677]_ , \new_[23680]_ ,
    \new_[23683]_ , \new_[23684]_ , \new_[23685]_ , \new_[23689]_ ,
    \new_[23690]_ , \new_[23693]_ , \new_[23696]_ , \new_[23697]_ ,
    \new_[23698]_ , \new_[23702]_ , \new_[23703]_ , \new_[23706]_ ,
    \new_[23709]_ , \new_[23710]_ , \new_[23711]_ , \new_[23715]_ ,
    \new_[23716]_ , \new_[23719]_ , \new_[23722]_ , \new_[23723]_ ,
    \new_[23724]_ , \new_[23728]_ , \new_[23729]_ , \new_[23732]_ ,
    \new_[23735]_ , \new_[23736]_ , \new_[23737]_ , \new_[23741]_ ,
    \new_[23742]_ , \new_[23745]_ , \new_[23748]_ , \new_[23749]_ ,
    \new_[23750]_ , \new_[23754]_ , \new_[23755]_ , \new_[23758]_ ,
    \new_[23761]_ , \new_[23762]_ , \new_[23763]_ , \new_[23767]_ ,
    \new_[23768]_ , \new_[23771]_ , \new_[23774]_ , \new_[23775]_ ,
    \new_[23776]_ , \new_[23780]_ , \new_[23781]_ , \new_[23784]_ ,
    \new_[23787]_ , \new_[23788]_ , \new_[23789]_ , \new_[23793]_ ,
    \new_[23794]_ , \new_[23797]_ , \new_[23800]_ , \new_[23801]_ ,
    \new_[23802]_ , \new_[23806]_ , \new_[23807]_ , \new_[23810]_ ,
    \new_[23813]_ , \new_[23814]_ , \new_[23815]_ , \new_[23819]_ ,
    \new_[23820]_ , \new_[23823]_ , \new_[23826]_ , \new_[23827]_ ,
    \new_[23828]_ , \new_[23832]_ , \new_[23833]_ , \new_[23836]_ ,
    \new_[23839]_ , \new_[23840]_ , \new_[23841]_ , \new_[23845]_ ,
    \new_[23846]_ , \new_[23849]_ , \new_[23852]_ , \new_[23853]_ ,
    \new_[23854]_ , \new_[23858]_ , \new_[23859]_ , \new_[23862]_ ,
    \new_[23865]_ , \new_[23866]_ , \new_[23867]_ , \new_[23871]_ ,
    \new_[23872]_ , \new_[23875]_ , \new_[23878]_ , \new_[23879]_ ,
    \new_[23880]_ , \new_[23884]_ , \new_[23885]_ , \new_[23888]_ ,
    \new_[23891]_ , \new_[23892]_ , \new_[23893]_ , \new_[23897]_ ,
    \new_[23898]_ , \new_[23901]_ , \new_[23904]_ , \new_[23905]_ ,
    \new_[23906]_ , \new_[23910]_ , \new_[23911]_ , \new_[23914]_ ,
    \new_[23917]_ , \new_[23918]_ , \new_[23919]_ , \new_[23923]_ ,
    \new_[23924]_ , \new_[23927]_ , \new_[23930]_ , \new_[23931]_ ,
    \new_[23932]_ , \new_[23936]_ , \new_[23937]_ , \new_[23940]_ ,
    \new_[23943]_ , \new_[23944]_ , \new_[23945]_ , \new_[23949]_ ,
    \new_[23950]_ , \new_[23953]_ , \new_[23956]_ , \new_[23957]_ ,
    \new_[23958]_ , \new_[23962]_ , \new_[23963]_ , \new_[23966]_ ,
    \new_[23969]_ , \new_[23970]_ , \new_[23971]_ , \new_[23975]_ ,
    \new_[23976]_ , \new_[23979]_ , \new_[23982]_ , \new_[23983]_ ,
    \new_[23984]_ , \new_[23988]_ , \new_[23989]_ , \new_[23992]_ ,
    \new_[23995]_ , \new_[23996]_ , \new_[23997]_ , \new_[24001]_ ,
    \new_[24002]_ , \new_[24005]_ , \new_[24008]_ , \new_[24009]_ ,
    \new_[24010]_ , \new_[24014]_ , \new_[24015]_ , \new_[24018]_ ,
    \new_[24021]_ , \new_[24022]_ , \new_[24023]_ , \new_[24027]_ ,
    \new_[24028]_ , \new_[24031]_ , \new_[24034]_ , \new_[24035]_ ,
    \new_[24036]_ , \new_[24040]_ , \new_[24041]_ , \new_[24044]_ ,
    \new_[24047]_ , \new_[24048]_ , \new_[24049]_ , \new_[24053]_ ,
    \new_[24054]_ , \new_[24057]_ , \new_[24060]_ , \new_[24061]_ ,
    \new_[24062]_ , \new_[24066]_ , \new_[24067]_ , \new_[24070]_ ,
    \new_[24073]_ , \new_[24074]_ , \new_[24075]_ , \new_[24079]_ ,
    \new_[24080]_ , \new_[24083]_ , \new_[24086]_ , \new_[24087]_ ,
    \new_[24088]_ , \new_[24092]_ , \new_[24093]_ , \new_[24096]_ ,
    \new_[24099]_ , \new_[24100]_ , \new_[24101]_ , \new_[24105]_ ,
    \new_[24106]_ , \new_[24109]_ , \new_[24112]_ , \new_[24113]_ ,
    \new_[24114]_ , \new_[24118]_ , \new_[24119]_ , \new_[24122]_ ,
    \new_[24125]_ , \new_[24126]_ , \new_[24127]_ , \new_[24131]_ ,
    \new_[24132]_ , \new_[24135]_ , \new_[24138]_ , \new_[24139]_ ,
    \new_[24140]_ , \new_[24144]_ , \new_[24145]_ , \new_[24148]_ ,
    \new_[24151]_ , \new_[24152]_ , \new_[24153]_ , \new_[24157]_ ,
    \new_[24158]_ , \new_[24161]_ , \new_[24164]_ , \new_[24165]_ ,
    \new_[24166]_ , \new_[24170]_ , \new_[24171]_ , \new_[24174]_ ,
    \new_[24177]_ , \new_[24178]_ , \new_[24179]_ , \new_[24183]_ ,
    \new_[24184]_ , \new_[24187]_ , \new_[24190]_ , \new_[24191]_ ,
    \new_[24192]_ , \new_[24196]_ , \new_[24197]_ , \new_[24200]_ ,
    \new_[24203]_ , \new_[24204]_ , \new_[24205]_ , \new_[24209]_ ,
    \new_[24210]_ , \new_[24213]_ , \new_[24216]_ , \new_[24217]_ ,
    \new_[24218]_ , \new_[24222]_ , \new_[24223]_ , \new_[24226]_ ,
    \new_[24229]_ , \new_[24230]_ , \new_[24231]_ , \new_[24235]_ ,
    \new_[24236]_ , \new_[24239]_ , \new_[24242]_ , \new_[24243]_ ,
    \new_[24244]_ , \new_[24248]_ , \new_[24249]_ , \new_[24252]_ ,
    \new_[24255]_ , \new_[24256]_ , \new_[24257]_ , \new_[24261]_ ,
    \new_[24262]_ , \new_[24265]_ , \new_[24268]_ , \new_[24269]_ ,
    \new_[24270]_ , \new_[24274]_ , \new_[24275]_ , \new_[24278]_ ,
    \new_[24281]_ , \new_[24282]_ , \new_[24283]_ , \new_[24287]_ ,
    \new_[24288]_ , \new_[24291]_ , \new_[24294]_ , \new_[24295]_ ,
    \new_[24296]_ , \new_[24300]_ , \new_[24301]_ , \new_[24304]_ ,
    \new_[24307]_ , \new_[24308]_ , \new_[24309]_ , \new_[24313]_ ,
    \new_[24314]_ , \new_[24317]_ , \new_[24320]_ , \new_[24321]_ ,
    \new_[24322]_ , \new_[24326]_ , \new_[24327]_ , \new_[24330]_ ,
    \new_[24333]_ , \new_[24334]_ , \new_[24335]_ , \new_[24339]_ ,
    \new_[24340]_ , \new_[24343]_ , \new_[24346]_ , \new_[24347]_ ,
    \new_[24348]_ , \new_[24352]_ , \new_[24353]_ , \new_[24356]_ ,
    \new_[24359]_ , \new_[24360]_ , \new_[24361]_ , \new_[24365]_ ,
    \new_[24366]_ , \new_[24369]_ , \new_[24372]_ , \new_[24373]_ ,
    \new_[24374]_ , \new_[24378]_ , \new_[24379]_ , \new_[24382]_ ,
    \new_[24385]_ , \new_[24386]_ , \new_[24387]_ , \new_[24391]_ ,
    \new_[24392]_ , \new_[24395]_ , \new_[24398]_ , \new_[24399]_ ,
    \new_[24400]_ , \new_[24404]_ , \new_[24405]_ , \new_[24408]_ ,
    \new_[24411]_ , \new_[24412]_ , \new_[24413]_ , \new_[24417]_ ,
    \new_[24418]_ , \new_[24421]_ , \new_[24424]_ , \new_[24425]_ ,
    \new_[24426]_ , \new_[24430]_ , \new_[24431]_ , \new_[24434]_ ,
    \new_[24437]_ , \new_[24438]_ , \new_[24439]_ , \new_[24443]_ ,
    \new_[24444]_ , \new_[24447]_ , \new_[24450]_ , \new_[24451]_ ,
    \new_[24452]_ , \new_[24456]_ , \new_[24457]_ , \new_[24460]_ ,
    \new_[24463]_ , \new_[24464]_ , \new_[24465]_ , \new_[24469]_ ,
    \new_[24470]_ , \new_[24473]_ , \new_[24476]_ , \new_[24477]_ ,
    \new_[24478]_ , \new_[24482]_ , \new_[24483]_ , \new_[24486]_ ,
    \new_[24489]_ , \new_[24490]_ , \new_[24491]_ , \new_[24495]_ ,
    \new_[24496]_ , \new_[24499]_ , \new_[24502]_ , \new_[24503]_ ,
    \new_[24504]_ , \new_[24508]_ , \new_[24509]_ , \new_[24512]_ ,
    \new_[24515]_ , \new_[24516]_ , \new_[24517]_ , \new_[24521]_ ,
    \new_[24522]_ , \new_[24525]_ , \new_[24528]_ , \new_[24529]_ ,
    \new_[24530]_ , \new_[24534]_ , \new_[24535]_ , \new_[24538]_ ,
    \new_[24541]_ , \new_[24542]_ , \new_[24543]_ , \new_[24547]_ ,
    \new_[24548]_ , \new_[24551]_ , \new_[24554]_ , \new_[24555]_ ,
    \new_[24556]_ , \new_[24560]_ , \new_[24561]_ , \new_[24564]_ ,
    \new_[24567]_ , \new_[24568]_ , \new_[24569]_ , \new_[24573]_ ,
    \new_[24574]_ , \new_[24577]_ , \new_[24580]_ , \new_[24581]_ ,
    \new_[24582]_ , \new_[24586]_ , \new_[24587]_ , \new_[24590]_ ,
    \new_[24593]_ , \new_[24594]_ , \new_[24595]_ , \new_[24599]_ ,
    \new_[24600]_ , \new_[24603]_ , \new_[24606]_ , \new_[24607]_ ,
    \new_[24608]_ , \new_[24612]_ , \new_[24613]_ , \new_[24616]_ ,
    \new_[24619]_ , \new_[24620]_ , \new_[24621]_ , \new_[24625]_ ,
    \new_[24626]_ , \new_[24629]_ , \new_[24632]_ , \new_[24633]_ ,
    \new_[24634]_ , \new_[24638]_ , \new_[24639]_ , \new_[24642]_ ,
    \new_[24645]_ , \new_[24646]_ , \new_[24647]_ , \new_[24651]_ ,
    \new_[24652]_ , \new_[24655]_ , \new_[24658]_ , \new_[24659]_ ,
    \new_[24660]_ , \new_[24664]_ , \new_[24665]_ , \new_[24668]_ ,
    \new_[24671]_ , \new_[24672]_ , \new_[24673]_ , \new_[24677]_ ,
    \new_[24678]_ , \new_[24681]_ , \new_[24684]_ , \new_[24685]_ ,
    \new_[24686]_ , \new_[24690]_ , \new_[24691]_ , \new_[24694]_ ,
    \new_[24697]_ , \new_[24698]_ , \new_[24699]_ , \new_[24703]_ ,
    \new_[24704]_ , \new_[24707]_ , \new_[24710]_ , \new_[24711]_ ,
    \new_[24712]_ , \new_[24716]_ , \new_[24717]_ , \new_[24720]_ ,
    \new_[24723]_ , \new_[24724]_ , \new_[24725]_ , \new_[24729]_ ,
    \new_[24730]_ , \new_[24733]_ , \new_[24736]_ , \new_[24737]_ ,
    \new_[24738]_ , \new_[24742]_ , \new_[24743]_ , \new_[24746]_ ,
    \new_[24749]_ , \new_[24750]_ , \new_[24751]_ , \new_[24755]_ ,
    \new_[24756]_ , \new_[24759]_ , \new_[24762]_ , \new_[24763]_ ,
    \new_[24764]_ , \new_[24768]_ , \new_[24769]_ , \new_[24772]_ ,
    \new_[24775]_ , \new_[24776]_ , \new_[24777]_ , \new_[24781]_ ,
    \new_[24782]_ , \new_[24785]_ , \new_[24788]_ , \new_[24789]_ ,
    \new_[24790]_ , \new_[24794]_ , \new_[24795]_ , \new_[24798]_ ,
    \new_[24801]_ , \new_[24802]_ , \new_[24803]_ , \new_[24807]_ ,
    \new_[24808]_ , \new_[24811]_ , \new_[24814]_ , \new_[24815]_ ,
    \new_[24816]_ , \new_[24820]_ , \new_[24821]_ , \new_[24824]_ ,
    \new_[24827]_ , \new_[24828]_ , \new_[24829]_ , \new_[24833]_ ,
    \new_[24834]_ , \new_[24837]_ , \new_[24840]_ , \new_[24841]_ ,
    \new_[24842]_ , \new_[24846]_ , \new_[24847]_ , \new_[24850]_ ,
    \new_[24853]_ , \new_[24854]_ , \new_[24855]_ , \new_[24859]_ ,
    \new_[24860]_ , \new_[24863]_ , \new_[24866]_ , \new_[24867]_ ,
    \new_[24868]_ , \new_[24872]_ , \new_[24873]_ , \new_[24876]_ ,
    \new_[24879]_ , \new_[24880]_ , \new_[24881]_ , \new_[24885]_ ,
    \new_[24886]_ , \new_[24889]_ , \new_[24892]_ , \new_[24893]_ ,
    \new_[24894]_ , \new_[24898]_ , \new_[24899]_ , \new_[24902]_ ,
    \new_[24905]_ , \new_[24906]_ , \new_[24907]_ , \new_[24911]_ ,
    \new_[24912]_ , \new_[24915]_ , \new_[24918]_ , \new_[24919]_ ,
    \new_[24920]_ , \new_[24924]_ , \new_[24925]_ , \new_[24928]_ ,
    \new_[24931]_ , \new_[24932]_ , \new_[24933]_ , \new_[24937]_ ,
    \new_[24938]_ , \new_[24941]_ , \new_[24944]_ , \new_[24945]_ ,
    \new_[24946]_ , \new_[24950]_ , \new_[24951]_ , \new_[24954]_ ,
    \new_[24957]_ , \new_[24958]_ , \new_[24959]_ , \new_[24963]_ ,
    \new_[24964]_ , \new_[24967]_ , \new_[24970]_ , \new_[24971]_ ,
    \new_[24972]_ , \new_[24976]_ , \new_[24977]_ , \new_[24980]_ ,
    \new_[24983]_ , \new_[24984]_ , \new_[24985]_ , \new_[24989]_ ,
    \new_[24990]_ , \new_[24993]_ , \new_[24996]_ , \new_[24997]_ ,
    \new_[24998]_ , \new_[25002]_ , \new_[25003]_ , \new_[25006]_ ,
    \new_[25009]_ , \new_[25010]_ , \new_[25011]_ , \new_[25015]_ ,
    \new_[25016]_ , \new_[25019]_ , \new_[25022]_ , \new_[25023]_ ,
    \new_[25024]_ , \new_[25028]_ , \new_[25029]_ , \new_[25032]_ ,
    \new_[25035]_ , \new_[25036]_ , \new_[25037]_ , \new_[25041]_ ,
    \new_[25042]_ , \new_[25045]_ , \new_[25048]_ , \new_[25049]_ ,
    \new_[25050]_ , \new_[25054]_ , \new_[25055]_ , \new_[25058]_ ,
    \new_[25061]_ , \new_[25062]_ , \new_[25063]_ , \new_[25067]_ ,
    \new_[25068]_ , \new_[25071]_ , \new_[25074]_ , \new_[25075]_ ,
    \new_[25076]_ , \new_[25080]_ , \new_[25081]_ , \new_[25084]_ ,
    \new_[25087]_ , \new_[25088]_ , \new_[25089]_ , \new_[25093]_ ,
    \new_[25094]_ , \new_[25097]_ , \new_[25100]_ , \new_[25101]_ ,
    \new_[25102]_ , \new_[25106]_ , \new_[25107]_ , \new_[25110]_ ,
    \new_[25113]_ , \new_[25114]_ , \new_[25115]_ , \new_[25119]_ ,
    \new_[25120]_ , \new_[25123]_ , \new_[25126]_ , \new_[25127]_ ,
    \new_[25128]_ , \new_[25132]_ , \new_[25133]_ , \new_[25136]_ ,
    \new_[25139]_ , \new_[25140]_ , \new_[25141]_ , \new_[25145]_ ,
    \new_[25146]_ , \new_[25149]_ , \new_[25152]_ , \new_[25153]_ ,
    \new_[25154]_ , \new_[25158]_ , \new_[25159]_ , \new_[25162]_ ,
    \new_[25165]_ , \new_[25166]_ , \new_[25167]_ , \new_[25171]_ ,
    \new_[25172]_ , \new_[25175]_ , \new_[25178]_ , \new_[25179]_ ,
    \new_[25180]_ , \new_[25184]_ , \new_[25185]_ , \new_[25188]_ ,
    \new_[25191]_ , \new_[25192]_ , \new_[25193]_ , \new_[25197]_ ,
    \new_[25198]_ , \new_[25201]_ , \new_[25204]_ , \new_[25205]_ ,
    \new_[25206]_ , \new_[25210]_ , \new_[25211]_ , \new_[25214]_ ,
    \new_[25217]_ , \new_[25218]_ , \new_[25219]_ , \new_[25223]_ ,
    \new_[25224]_ , \new_[25227]_ , \new_[25230]_ , \new_[25231]_ ,
    \new_[25232]_ , \new_[25236]_ , \new_[25237]_ , \new_[25240]_ ,
    \new_[25243]_ , \new_[25244]_ , \new_[25245]_ , \new_[25249]_ ,
    \new_[25250]_ , \new_[25253]_ , \new_[25256]_ , \new_[25257]_ ,
    \new_[25258]_ , \new_[25262]_ , \new_[25263]_ , \new_[25266]_ ,
    \new_[25269]_ , \new_[25270]_ , \new_[25271]_ , \new_[25275]_ ,
    \new_[25276]_ , \new_[25279]_ , \new_[25282]_ , \new_[25283]_ ,
    \new_[25284]_ , \new_[25288]_ , \new_[25289]_ , \new_[25292]_ ,
    \new_[25295]_ , \new_[25296]_ , \new_[25297]_ , \new_[25301]_ ,
    \new_[25302]_ , \new_[25305]_ , \new_[25308]_ , \new_[25309]_ ,
    \new_[25310]_ , \new_[25314]_ , \new_[25315]_ , \new_[25318]_ ,
    \new_[25321]_ , \new_[25322]_ , \new_[25323]_ , \new_[25327]_ ,
    \new_[25328]_ , \new_[25331]_ , \new_[25334]_ , \new_[25335]_ ,
    \new_[25336]_ , \new_[25340]_ , \new_[25341]_ , \new_[25344]_ ,
    \new_[25347]_ , \new_[25348]_ , \new_[25349]_ , \new_[25353]_ ,
    \new_[25354]_ , \new_[25357]_ , \new_[25360]_ , \new_[25361]_ ,
    \new_[25362]_ , \new_[25366]_ , \new_[25367]_ , \new_[25370]_ ,
    \new_[25373]_ , \new_[25374]_ , \new_[25375]_ , \new_[25379]_ ,
    \new_[25380]_ , \new_[25383]_ , \new_[25386]_ , \new_[25387]_ ,
    \new_[25388]_ , \new_[25392]_ , \new_[25393]_ , \new_[25396]_ ,
    \new_[25399]_ , \new_[25400]_ , \new_[25401]_ , \new_[25405]_ ,
    \new_[25406]_ , \new_[25409]_ , \new_[25412]_ , \new_[25413]_ ,
    \new_[25414]_ , \new_[25418]_ , \new_[25419]_ , \new_[25422]_ ,
    \new_[25425]_ , \new_[25426]_ , \new_[25427]_ , \new_[25431]_ ,
    \new_[25432]_ , \new_[25435]_ , \new_[25438]_ , \new_[25439]_ ,
    \new_[25440]_ , \new_[25444]_ , \new_[25445]_ , \new_[25448]_ ,
    \new_[25451]_ , \new_[25452]_ , \new_[25453]_ , \new_[25457]_ ,
    \new_[25458]_ , \new_[25461]_ , \new_[25464]_ , \new_[25465]_ ,
    \new_[25466]_ , \new_[25470]_ , \new_[25471]_ , \new_[25474]_ ,
    \new_[25477]_ , \new_[25478]_ , \new_[25479]_ , \new_[25483]_ ,
    \new_[25484]_ , \new_[25487]_ , \new_[25490]_ , \new_[25491]_ ,
    \new_[25492]_ , \new_[25496]_ , \new_[25497]_ , \new_[25500]_ ,
    \new_[25503]_ , \new_[25504]_ , \new_[25505]_ , \new_[25509]_ ,
    \new_[25510]_ , \new_[25513]_ , \new_[25516]_ , \new_[25517]_ ,
    \new_[25518]_ , \new_[25522]_ , \new_[25523]_ , \new_[25526]_ ,
    \new_[25529]_ , \new_[25530]_ , \new_[25531]_ , \new_[25535]_ ,
    \new_[25536]_ , \new_[25539]_ , \new_[25542]_ , \new_[25543]_ ,
    \new_[25544]_ , \new_[25548]_ , \new_[25549]_ , \new_[25552]_ ,
    \new_[25555]_ , \new_[25556]_ , \new_[25557]_ , \new_[25561]_ ,
    \new_[25562]_ , \new_[25565]_ , \new_[25568]_ , \new_[25569]_ ,
    \new_[25570]_ , \new_[25574]_ , \new_[25575]_ , \new_[25578]_ ,
    \new_[25581]_ , \new_[25582]_ , \new_[25583]_ , \new_[25587]_ ,
    \new_[25588]_ , \new_[25591]_ , \new_[25594]_ , \new_[25595]_ ,
    \new_[25596]_ , \new_[25600]_ , \new_[25601]_ , \new_[25604]_ ,
    \new_[25607]_ , \new_[25608]_ , \new_[25609]_ , \new_[25613]_ ,
    \new_[25614]_ , \new_[25617]_ , \new_[25620]_ , \new_[25621]_ ,
    \new_[25622]_ , \new_[25626]_ , \new_[25627]_ , \new_[25630]_ ,
    \new_[25633]_ , \new_[25634]_ , \new_[25635]_ , \new_[25639]_ ,
    \new_[25640]_ , \new_[25643]_ , \new_[25646]_ , \new_[25647]_ ,
    \new_[25648]_ , \new_[25652]_ , \new_[25653]_ , \new_[25656]_ ,
    \new_[25659]_ , \new_[25660]_ , \new_[25661]_ , \new_[25665]_ ,
    \new_[25666]_ , \new_[25669]_ , \new_[25672]_ , \new_[25673]_ ,
    \new_[25674]_ , \new_[25678]_ , \new_[25679]_ , \new_[25682]_ ,
    \new_[25685]_ , \new_[25686]_ , \new_[25687]_ , \new_[25691]_ ,
    \new_[25692]_ , \new_[25695]_ , \new_[25698]_ , \new_[25699]_ ,
    \new_[25700]_ , \new_[25704]_ , \new_[25705]_ , \new_[25708]_ ,
    \new_[25711]_ , \new_[25712]_ , \new_[25713]_ , \new_[25717]_ ,
    \new_[25718]_ , \new_[25721]_ , \new_[25724]_ , \new_[25725]_ ,
    \new_[25726]_ , \new_[25730]_ , \new_[25731]_ , \new_[25734]_ ,
    \new_[25737]_ , \new_[25738]_ , \new_[25739]_ , \new_[25743]_ ,
    \new_[25744]_ , \new_[25747]_ , \new_[25750]_ , \new_[25751]_ ,
    \new_[25752]_ , \new_[25756]_ , \new_[25757]_ , \new_[25760]_ ,
    \new_[25763]_ , \new_[25764]_ , \new_[25765]_ , \new_[25769]_ ,
    \new_[25770]_ , \new_[25773]_ , \new_[25776]_ , \new_[25777]_ ,
    \new_[25778]_ , \new_[25782]_ , \new_[25783]_ , \new_[25786]_ ,
    \new_[25789]_ , \new_[25790]_ , \new_[25791]_ , \new_[25795]_ ,
    \new_[25796]_ , \new_[25799]_ , \new_[25802]_ , \new_[25803]_ ,
    \new_[25804]_ , \new_[25808]_ , \new_[25809]_ , \new_[25812]_ ,
    \new_[25815]_ , \new_[25816]_ , \new_[25817]_ , \new_[25821]_ ,
    \new_[25822]_ , \new_[25825]_ , \new_[25828]_ , \new_[25829]_ ,
    \new_[25830]_ , \new_[25834]_ , \new_[25835]_ , \new_[25838]_ ,
    \new_[25841]_ , \new_[25842]_ , \new_[25843]_ , \new_[25847]_ ,
    \new_[25848]_ , \new_[25851]_ , \new_[25854]_ , \new_[25855]_ ,
    \new_[25856]_ , \new_[25860]_ , \new_[25861]_ , \new_[25864]_ ,
    \new_[25867]_ , \new_[25868]_ , \new_[25869]_ , \new_[25873]_ ,
    \new_[25874]_ , \new_[25877]_ , \new_[25880]_ , \new_[25881]_ ,
    \new_[25882]_ , \new_[25886]_ , \new_[25887]_ , \new_[25890]_ ,
    \new_[25893]_ , \new_[25894]_ , \new_[25895]_ , \new_[25899]_ ,
    \new_[25900]_ , \new_[25903]_ , \new_[25906]_ , \new_[25907]_ ,
    \new_[25908]_ , \new_[25912]_ , \new_[25913]_ , \new_[25916]_ ,
    \new_[25919]_ , \new_[25920]_ , \new_[25921]_ , \new_[25925]_ ,
    \new_[25926]_ , \new_[25929]_ , \new_[25932]_ , \new_[25933]_ ,
    \new_[25934]_ , \new_[25938]_ , \new_[25939]_ , \new_[25942]_ ,
    \new_[25945]_ , \new_[25946]_ , \new_[25947]_ , \new_[25951]_ ,
    \new_[25952]_ , \new_[25955]_ , \new_[25958]_ , \new_[25959]_ ,
    \new_[25960]_ , \new_[25964]_ , \new_[25965]_ , \new_[25968]_ ,
    \new_[25971]_ , \new_[25972]_ , \new_[25973]_ , \new_[25977]_ ,
    \new_[25978]_ , \new_[25981]_ , \new_[25984]_ , \new_[25985]_ ,
    \new_[25986]_ , \new_[25990]_ , \new_[25991]_ , \new_[25994]_ ,
    \new_[25997]_ , \new_[25998]_ , \new_[25999]_ , \new_[26003]_ ,
    \new_[26004]_ , \new_[26007]_ , \new_[26010]_ , \new_[26011]_ ,
    \new_[26012]_ , \new_[26016]_ , \new_[26017]_ , \new_[26020]_ ,
    \new_[26023]_ , \new_[26024]_ , \new_[26025]_ , \new_[26029]_ ,
    \new_[26030]_ , \new_[26033]_ , \new_[26036]_ , \new_[26037]_ ,
    \new_[26038]_ , \new_[26042]_ , \new_[26043]_ , \new_[26046]_ ,
    \new_[26049]_ , \new_[26050]_ , \new_[26051]_ , \new_[26055]_ ,
    \new_[26056]_ , \new_[26059]_ , \new_[26062]_ , \new_[26063]_ ,
    \new_[26064]_ , \new_[26068]_ , \new_[26069]_ , \new_[26072]_ ,
    \new_[26075]_ , \new_[26076]_ , \new_[26077]_ , \new_[26081]_ ,
    \new_[26082]_ , \new_[26085]_ , \new_[26088]_ , \new_[26089]_ ,
    \new_[26090]_ , \new_[26094]_ , \new_[26095]_ , \new_[26098]_ ,
    \new_[26101]_ , \new_[26102]_ , \new_[26103]_ , \new_[26107]_ ,
    \new_[26108]_ , \new_[26111]_ , \new_[26114]_ , \new_[26115]_ ,
    \new_[26116]_ , \new_[26120]_ , \new_[26121]_ , \new_[26124]_ ,
    \new_[26127]_ , \new_[26128]_ , \new_[26129]_ , \new_[26133]_ ,
    \new_[26134]_ , \new_[26137]_ , \new_[26140]_ , \new_[26141]_ ,
    \new_[26142]_ , \new_[26146]_ , \new_[26147]_ , \new_[26150]_ ,
    \new_[26153]_ , \new_[26154]_ , \new_[26155]_ , \new_[26159]_ ,
    \new_[26160]_ , \new_[26163]_ , \new_[26166]_ , \new_[26167]_ ,
    \new_[26168]_ , \new_[26172]_ , \new_[26173]_ , \new_[26176]_ ,
    \new_[26179]_ , \new_[26180]_ , \new_[26181]_ , \new_[26185]_ ,
    \new_[26186]_ , \new_[26189]_ , \new_[26192]_ , \new_[26193]_ ,
    \new_[26194]_ , \new_[26198]_ , \new_[26199]_ , \new_[26202]_ ,
    \new_[26205]_ , \new_[26206]_ , \new_[26207]_ , \new_[26211]_ ,
    \new_[26212]_ , \new_[26215]_ , \new_[26218]_ , \new_[26219]_ ,
    \new_[26220]_ , \new_[26223]_ , \new_[26226]_ , \new_[26227]_ ,
    \new_[26230]_ , \new_[26233]_ , \new_[26234]_ , \new_[26235]_ ,
    \new_[26239]_ , \new_[26240]_ , \new_[26243]_ , \new_[26246]_ ,
    \new_[26247]_ , \new_[26248]_ , \new_[26251]_ , \new_[26254]_ ,
    \new_[26255]_ , \new_[26258]_ , \new_[26261]_ , \new_[26262]_ ,
    \new_[26263]_ , \new_[26267]_ , \new_[26268]_ , \new_[26271]_ ,
    \new_[26274]_ , \new_[26275]_ , \new_[26276]_ , \new_[26279]_ ,
    \new_[26282]_ , \new_[26283]_ , \new_[26286]_ , \new_[26289]_ ,
    \new_[26290]_ , \new_[26291]_ , \new_[26295]_ , \new_[26296]_ ,
    \new_[26299]_ , \new_[26302]_ , \new_[26303]_ , \new_[26304]_ ,
    \new_[26307]_ , \new_[26310]_ , \new_[26311]_ , \new_[26314]_ ,
    \new_[26317]_ , \new_[26318]_ , \new_[26319]_ , \new_[26323]_ ,
    \new_[26324]_ , \new_[26327]_ , \new_[26330]_ , \new_[26331]_ ,
    \new_[26332]_ , \new_[26335]_ , \new_[26338]_ , \new_[26339]_ ,
    \new_[26342]_ , \new_[26345]_ , \new_[26346]_ , \new_[26347]_ ,
    \new_[26351]_ , \new_[26352]_ , \new_[26355]_ , \new_[26358]_ ,
    \new_[26359]_ , \new_[26360]_ , \new_[26363]_ , \new_[26366]_ ,
    \new_[26367]_ , \new_[26370]_ , \new_[26373]_ , \new_[26374]_ ,
    \new_[26375]_ , \new_[26379]_ , \new_[26380]_ , \new_[26383]_ ,
    \new_[26386]_ , \new_[26387]_ , \new_[26388]_ , \new_[26391]_ ,
    \new_[26394]_ , \new_[26395]_ , \new_[26398]_ , \new_[26401]_ ,
    \new_[26402]_ , \new_[26403]_ , \new_[26407]_ , \new_[26408]_ ,
    \new_[26411]_ , \new_[26414]_ , \new_[26415]_ , \new_[26416]_ ,
    \new_[26419]_ , \new_[26422]_ , \new_[26423]_ , \new_[26426]_ ,
    \new_[26429]_ , \new_[26430]_ , \new_[26431]_ , \new_[26435]_ ,
    \new_[26436]_ , \new_[26439]_ , \new_[26442]_ , \new_[26443]_ ,
    \new_[26444]_ , \new_[26447]_ , \new_[26450]_ , \new_[26451]_ ,
    \new_[26454]_ , \new_[26457]_ , \new_[26458]_ , \new_[26459]_ ,
    \new_[26463]_ , \new_[26464]_ , \new_[26467]_ , \new_[26470]_ ,
    \new_[26471]_ , \new_[26472]_ , \new_[26475]_ , \new_[26478]_ ,
    \new_[26479]_ , \new_[26482]_ , \new_[26485]_ , \new_[26486]_ ,
    \new_[26487]_ , \new_[26491]_ , \new_[26492]_ , \new_[26495]_ ,
    \new_[26498]_ , \new_[26499]_ , \new_[26500]_ , \new_[26503]_ ,
    \new_[26506]_ , \new_[26507]_ , \new_[26510]_ , \new_[26513]_ ,
    \new_[26514]_ , \new_[26515]_ , \new_[26519]_ , \new_[26520]_ ,
    \new_[26523]_ , \new_[26526]_ , \new_[26527]_ , \new_[26528]_ ,
    \new_[26531]_ , \new_[26534]_ , \new_[26535]_ , \new_[26538]_ ,
    \new_[26541]_ , \new_[26542]_ , \new_[26543]_ , \new_[26547]_ ,
    \new_[26548]_ , \new_[26551]_ , \new_[26554]_ , \new_[26555]_ ,
    \new_[26556]_ , \new_[26559]_ , \new_[26562]_ , \new_[26563]_ ,
    \new_[26566]_ , \new_[26569]_ , \new_[26570]_ , \new_[26571]_ ,
    \new_[26575]_ , \new_[26576]_ , \new_[26579]_ , \new_[26582]_ ,
    \new_[26583]_ , \new_[26584]_ , \new_[26587]_ , \new_[26590]_ ,
    \new_[26591]_ , \new_[26594]_ , \new_[26597]_ , \new_[26598]_ ,
    \new_[26599]_ , \new_[26603]_ , \new_[26604]_ , \new_[26607]_ ,
    \new_[26610]_ , \new_[26611]_ , \new_[26612]_ , \new_[26615]_ ,
    \new_[26618]_ , \new_[26619]_ , \new_[26622]_ , \new_[26625]_ ,
    \new_[26626]_ , \new_[26627]_ , \new_[26631]_ , \new_[26632]_ ,
    \new_[26635]_ , \new_[26638]_ , \new_[26639]_ , \new_[26640]_ ,
    \new_[26643]_ , \new_[26646]_ , \new_[26647]_ , \new_[26650]_ ,
    \new_[26653]_ , \new_[26654]_ , \new_[26655]_ , \new_[26659]_ ,
    \new_[26660]_ , \new_[26663]_ , \new_[26666]_ , \new_[26667]_ ,
    \new_[26668]_ , \new_[26671]_ , \new_[26674]_ , \new_[26675]_ ,
    \new_[26678]_ , \new_[26681]_ , \new_[26682]_ , \new_[26683]_ ,
    \new_[26687]_ , \new_[26688]_ , \new_[26691]_ , \new_[26694]_ ,
    \new_[26695]_ , \new_[26696]_ , \new_[26699]_ , \new_[26702]_ ,
    \new_[26703]_ , \new_[26706]_ , \new_[26709]_ , \new_[26710]_ ,
    \new_[26711]_ , \new_[26715]_ , \new_[26716]_ , \new_[26719]_ ,
    \new_[26722]_ , \new_[26723]_ , \new_[26724]_ , \new_[26727]_ ,
    \new_[26730]_ , \new_[26731]_ , \new_[26734]_ , \new_[26737]_ ,
    \new_[26738]_ , \new_[26739]_ , \new_[26743]_ , \new_[26744]_ ,
    \new_[26747]_ , \new_[26750]_ , \new_[26751]_ , \new_[26752]_ ,
    \new_[26755]_ , \new_[26758]_ , \new_[26759]_ , \new_[26762]_ ,
    \new_[26765]_ , \new_[26766]_ , \new_[26767]_ , \new_[26771]_ ,
    \new_[26772]_ , \new_[26775]_ , \new_[26778]_ , \new_[26779]_ ,
    \new_[26780]_ , \new_[26783]_ , \new_[26786]_ , \new_[26787]_ ,
    \new_[26790]_ , \new_[26793]_ , \new_[26794]_ , \new_[26795]_ ,
    \new_[26799]_ , \new_[26800]_ , \new_[26803]_ , \new_[26806]_ ,
    \new_[26807]_ , \new_[26808]_ , \new_[26811]_ , \new_[26814]_ ,
    \new_[26815]_ , \new_[26818]_ , \new_[26821]_ , \new_[26822]_ ,
    \new_[26823]_ , \new_[26827]_ , \new_[26828]_ , \new_[26831]_ ,
    \new_[26834]_ , \new_[26835]_ , \new_[26836]_ , \new_[26839]_ ,
    \new_[26842]_ , \new_[26843]_ , \new_[26846]_ , \new_[26849]_ ,
    \new_[26850]_ , \new_[26851]_ , \new_[26855]_ , \new_[26856]_ ,
    \new_[26859]_ , \new_[26862]_ , \new_[26863]_ , \new_[26864]_ ,
    \new_[26867]_ , \new_[26870]_ , \new_[26871]_ , \new_[26874]_ ,
    \new_[26877]_ , \new_[26878]_ , \new_[26879]_ , \new_[26883]_ ,
    \new_[26884]_ , \new_[26887]_ , \new_[26890]_ , \new_[26891]_ ,
    \new_[26892]_ , \new_[26895]_ , \new_[26898]_ , \new_[26899]_ ,
    \new_[26902]_ , \new_[26905]_ , \new_[26906]_ , \new_[26907]_ ,
    \new_[26911]_ , \new_[26912]_ , \new_[26915]_ , \new_[26918]_ ,
    \new_[26919]_ , \new_[26920]_ , \new_[26923]_ , \new_[26926]_ ,
    \new_[26927]_ , \new_[26930]_ , \new_[26933]_ , \new_[26934]_ ,
    \new_[26935]_ , \new_[26939]_ , \new_[26940]_ , \new_[26943]_ ,
    \new_[26946]_ , \new_[26947]_ , \new_[26948]_ , \new_[26951]_ ,
    \new_[26954]_ , \new_[26955]_ , \new_[26958]_ , \new_[26961]_ ,
    \new_[26962]_ , \new_[26963]_ , \new_[26967]_ , \new_[26968]_ ,
    \new_[26971]_ , \new_[26974]_ , \new_[26975]_ , \new_[26976]_ ,
    \new_[26979]_ , \new_[26982]_ , \new_[26983]_ , \new_[26986]_ ,
    \new_[26989]_ , \new_[26990]_ , \new_[26991]_ ;
  assign A106 = \new_[3355]_  | \new_[2236]_ ;
  assign \new_[1]_  = \new_[26991]_  & \new_[26976]_ ;
  assign \new_[2]_  = \new_[26963]_  & \new_[26948]_ ;
  assign \new_[3]_  = \new_[26935]_  & \new_[26920]_ ;
  assign \new_[4]_  = \new_[26907]_  & \new_[26892]_ ;
  assign \new_[5]_  = \new_[26879]_  & \new_[26864]_ ;
  assign \new_[6]_  = \new_[26851]_  & \new_[26836]_ ;
  assign \new_[7]_  = \new_[26823]_  & \new_[26808]_ ;
  assign \new_[8]_  = \new_[26795]_  & \new_[26780]_ ;
  assign \new_[9]_  = \new_[26767]_  & \new_[26752]_ ;
  assign \new_[10]_  = \new_[26739]_  & \new_[26724]_ ;
  assign \new_[11]_  = \new_[26711]_  & \new_[26696]_ ;
  assign \new_[12]_  = \new_[26683]_  & \new_[26668]_ ;
  assign \new_[13]_  = \new_[26655]_  & \new_[26640]_ ;
  assign \new_[14]_  = \new_[26627]_  & \new_[26612]_ ;
  assign \new_[15]_  = \new_[26599]_  & \new_[26584]_ ;
  assign \new_[16]_  = \new_[26571]_  & \new_[26556]_ ;
  assign \new_[17]_  = \new_[26543]_  & \new_[26528]_ ;
  assign \new_[18]_  = \new_[26515]_  & \new_[26500]_ ;
  assign \new_[19]_  = \new_[26487]_  & \new_[26472]_ ;
  assign \new_[20]_  = \new_[26459]_  & \new_[26444]_ ;
  assign \new_[21]_  = \new_[26431]_  & \new_[26416]_ ;
  assign \new_[22]_  = \new_[26403]_  & \new_[26388]_ ;
  assign \new_[23]_  = \new_[26375]_  & \new_[26360]_ ;
  assign \new_[24]_  = \new_[26347]_  & \new_[26332]_ ;
  assign \new_[25]_  = \new_[26319]_  & \new_[26304]_ ;
  assign \new_[26]_  = \new_[26291]_  & \new_[26276]_ ;
  assign \new_[27]_  = \new_[26263]_  & \new_[26248]_ ;
  assign \new_[28]_  = \new_[26235]_  & \new_[26220]_ ;
  assign \new_[29]_  = \new_[26207]_  & \new_[26194]_ ;
  assign \new_[30]_  = \new_[26181]_  & \new_[26168]_ ;
  assign \new_[31]_  = \new_[26155]_  & \new_[26142]_ ;
  assign \new_[32]_  = \new_[26129]_  & \new_[26116]_ ;
  assign \new_[33]_  = \new_[26103]_  & \new_[26090]_ ;
  assign \new_[34]_  = \new_[26077]_  & \new_[26064]_ ;
  assign \new_[35]_  = \new_[26051]_  & \new_[26038]_ ;
  assign \new_[36]_  = \new_[26025]_  & \new_[26012]_ ;
  assign \new_[37]_  = \new_[25999]_  & \new_[25986]_ ;
  assign \new_[38]_  = \new_[25973]_  & \new_[25960]_ ;
  assign \new_[39]_  = \new_[25947]_  & \new_[25934]_ ;
  assign \new_[40]_  = \new_[25921]_  & \new_[25908]_ ;
  assign \new_[41]_  = \new_[25895]_  & \new_[25882]_ ;
  assign \new_[42]_  = \new_[25869]_  & \new_[25856]_ ;
  assign \new_[43]_  = \new_[25843]_  & \new_[25830]_ ;
  assign \new_[44]_  = \new_[25817]_  & \new_[25804]_ ;
  assign \new_[45]_  = \new_[25791]_  & \new_[25778]_ ;
  assign \new_[46]_  = \new_[25765]_  & \new_[25752]_ ;
  assign \new_[47]_  = \new_[25739]_  & \new_[25726]_ ;
  assign \new_[48]_  = \new_[25713]_  & \new_[25700]_ ;
  assign \new_[49]_  = \new_[25687]_  & \new_[25674]_ ;
  assign \new_[50]_  = \new_[25661]_  & \new_[25648]_ ;
  assign \new_[51]_  = \new_[25635]_  & \new_[25622]_ ;
  assign \new_[52]_  = \new_[25609]_  & \new_[25596]_ ;
  assign \new_[53]_  = \new_[25583]_  & \new_[25570]_ ;
  assign \new_[54]_  = \new_[25557]_  & \new_[25544]_ ;
  assign \new_[55]_  = \new_[25531]_  & \new_[25518]_ ;
  assign \new_[56]_  = \new_[25505]_  & \new_[25492]_ ;
  assign \new_[57]_  = \new_[25479]_  & \new_[25466]_ ;
  assign \new_[58]_  = \new_[25453]_  & \new_[25440]_ ;
  assign \new_[59]_  = \new_[25427]_  & \new_[25414]_ ;
  assign \new_[60]_  = \new_[25401]_  & \new_[25388]_ ;
  assign \new_[61]_  = \new_[25375]_  & \new_[25362]_ ;
  assign \new_[62]_  = \new_[25349]_  & \new_[25336]_ ;
  assign \new_[63]_  = \new_[25323]_  & \new_[25310]_ ;
  assign \new_[64]_  = \new_[25297]_  & \new_[25284]_ ;
  assign \new_[65]_  = \new_[25271]_  & \new_[25258]_ ;
  assign \new_[66]_  = \new_[25245]_  & \new_[25232]_ ;
  assign \new_[67]_  = \new_[25219]_  & \new_[25206]_ ;
  assign \new_[68]_  = \new_[25193]_  & \new_[25180]_ ;
  assign \new_[69]_  = \new_[25167]_  & \new_[25154]_ ;
  assign \new_[70]_  = \new_[25141]_  & \new_[25128]_ ;
  assign \new_[71]_  = \new_[25115]_  & \new_[25102]_ ;
  assign \new_[72]_  = \new_[25089]_  & \new_[25076]_ ;
  assign \new_[73]_  = \new_[25063]_  & \new_[25050]_ ;
  assign \new_[74]_  = \new_[25037]_  & \new_[25024]_ ;
  assign \new_[75]_  = \new_[25011]_  & \new_[24998]_ ;
  assign \new_[76]_  = \new_[24985]_  & \new_[24972]_ ;
  assign \new_[77]_  = \new_[24959]_  & \new_[24946]_ ;
  assign \new_[78]_  = \new_[24933]_  & \new_[24920]_ ;
  assign \new_[79]_  = \new_[24907]_  & \new_[24894]_ ;
  assign \new_[80]_  = \new_[24881]_  & \new_[24868]_ ;
  assign \new_[81]_  = \new_[24855]_  & \new_[24842]_ ;
  assign \new_[82]_  = \new_[24829]_  & \new_[24816]_ ;
  assign \new_[83]_  = \new_[24803]_  & \new_[24790]_ ;
  assign \new_[84]_  = \new_[24777]_  & \new_[24764]_ ;
  assign \new_[85]_  = \new_[24751]_  & \new_[24738]_ ;
  assign \new_[86]_  = \new_[24725]_  & \new_[24712]_ ;
  assign \new_[87]_  = \new_[24699]_  & \new_[24686]_ ;
  assign \new_[88]_  = \new_[24673]_  & \new_[24660]_ ;
  assign \new_[89]_  = \new_[24647]_  & \new_[24634]_ ;
  assign \new_[90]_  = \new_[24621]_  & \new_[24608]_ ;
  assign \new_[91]_  = \new_[24595]_  & \new_[24582]_ ;
  assign \new_[92]_  = \new_[24569]_  & \new_[24556]_ ;
  assign \new_[93]_  = \new_[24543]_  & \new_[24530]_ ;
  assign \new_[94]_  = \new_[24517]_  & \new_[24504]_ ;
  assign \new_[95]_  = \new_[24491]_  & \new_[24478]_ ;
  assign \new_[96]_  = \new_[24465]_  & \new_[24452]_ ;
  assign \new_[97]_  = \new_[24439]_  & \new_[24426]_ ;
  assign \new_[98]_  = \new_[24413]_  & \new_[24400]_ ;
  assign \new_[99]_  = \new_[24387]_  & \new_[24374]_ ;
  assign \new_[100]_  = \new_[24361]_  & \new_[24348]_ ;
  assign \new_[101]_  = \new_[24335]_  & \new_[24322]_ ;
  assign \new_[102]_  = \new_[24309]_  & \new_[24296]_ ;
  assign \new_[103]_  = \new_[24283]_  & \new_[24270]_ ;
  assign \new_[104]_  = \new_[24257]_  & \new_[24244]_ ;
  assign \new_[105]_  = \new_[24231]_  & \new_[24218]_ ;
  assign \new_[106]_  = \new_[24205]_  & \new_[24192]_ ;
  assign \new_[107]_  = \new_[24179]_  & \new_[24166]_ ;
  assign \new_[108]_  = \new_[24153]_  & \new_[24140]_ ;
  assign \new_[109]_  = \new_[24127]_  & \new_[24114]_ ;
  assign \new_[110]_  = \new_[24101]_  & \new_[24088]_ ;
  assign \new_[111]_  = \new_[24075]_  & \new_[24062]_ ;
  assign \new_[112]_  = \new_[24049]_  & \new_[24036]_ ;
  assign \new_[113]_  = \new_[24023]_  & \new_[24010]_ ;
  assign \new_[114]_  = \new_[23997]_  & \new_[23984]_ ;
  assign \new_[115]_  = \new_[23971]_  & \new_[23958]_ ;
  assign \new_[116]_  = \new_[23945]_  & \new_[23932]_ ;
  assign \new_[117]_  = \new_[23919]_  & \new_[23906]_ ;
  assign \new_[118]_  = \new_[23893]_  & \new_[23880]_ ;
  assign \new_[119]_  = \new_[23867]_  & \new_[23854]_ ;
  assign \new_[120]_  = \new_[23841]_  & \new_[23828]_ ;
  assign \new_[121]_  = \new_[23815]_  & \new_[23802]_ ;
  assign \new_[122]_  = \new_[23789]_  & \new_[23776]_ ;
  assign \new_[123]_  = \new_[23763]_  & \new_[23750]_ ;
  assign \new_[124]_  = \new_[23737]_  & \new_[23724]_ ;
  assign \new_[125]_  = \new_[23711]_  & \new_[23698]_ ;
  assign \new_[126]_  = \new_[23685]_  & \new_[23672]_ ;
  assign \new_[127]_  = \new_[23659]_  & \new_[23646]_ ;
  assign \new_[128]_  = \new_[23633]_  & \new_[23620]_ ;
  assign \new_[129]_  = \new_[23607]_  & \new_[23594]_ ;
  assign \new_[130]_  = \new_[23581]_  & \new_[23568]_ ;
  assign \new_[131]_  = \new_[23555]_  & \new_[23542]_ ;
  assign \new_[132]_  = \new_[23529]_  & \new_[23516]_ ;
  assign \new_[133]_  = \new_[23503]_  & \new_[23490]_ ;
  assign \new_[134]_  = \new_[23477]_  & \new_[23464]_ ;
  assign \new_[135]_  = \new_[23451]_  & \new_[23438]_ ;
  assign \new_[136]_  = \new_[23425]_  & \new_[23412]_ ;
  assign \new_[137]_  = \new_[23399]_  & \new_[23386]_ ;
  assign \new_[138]_  = \new_[23373]_  & \new_[23360]_ ;
  assign \new_[139]_  = \new_[23347]_  & \new_[23334]_ ;
  assign \new_[140]_  = \new_[23321]_  & \new_[23308]_ ;
  assign \new_[141]_  = \new_[23295]_  & \new_[23282]_ ;
  assign \new_[142]_  = \new_[23269]_  & \new_[23256]_ ;
  assign \new_[143]_  = \new_[23243]_  & \new_[23230]_ ;
  assign \new_[144]_  = \new_[23219]_  & \new_[23206]_ ;
  assign \new_[145]_  = \new_[23195]_  & \new_[23182]_ ;
  assign \new_[146]_  = \new_[23171]_  & \new_[23158]_ ;
  assign \new_[147]_  = \new_[23147]_  & \new_[23134]_ ;
  assign \new_[148]_  = \new_[23123]_  & \new_[23110]_ ;
  assign \new_[149]_  = \new_[23099]_  & \new_[23086]_ ;
  assign \new_[150]_  = \new_[23075]_  & \new_[23062]_ ;
  assign \new_[151]_  = \new_[23051]_  & \new_[23038]_ ;
  assign \new_[152]_  = \new_[23027]_  & \new_[23014]_ ;
  assign \new_[153]_  = \new_[23003]_  & \new_[22990]_ ;
  assign \new_[154]_  = \new_[22979]_  & \new_[22966]_ ;
  assign \new_[155]_  = \new_[22955]_  & \new_[22942]_ ;
  assign \new_[156]_  = \new_[22931]_  & \new_[22918]_ ;
  assign \new_[157]_  = \new_[22907]_  & \new_[22894]_ ;
  assign \new_[158]_  = \new_[22883]_  & \new_[22870]_ ;
  assign \new_[159]_  = \new_[22859]_  & \new_[22846]_ ;
  assign \new_[160]_  = \new_[22835]_  & \new_[22822]_ ;
  assign \new_[161]_  = \new_[22811]_  & \new_[22798]_ ;
  assign \new_[162]_  = \new_[22787]_  & \new_[22774]_ ;
  assign \new_[163]_  = \new_[22763]_  & \new_[22750]_ ;
  assign \new_[164]_  = \new_[22739]_  & \new_[22726]_ ;
  assign \new_[165]_  = \new_[22715]_  & \new_[22702]_ ;
  assign \new_[166]_  = \new_[22691]_  & \new_[22678]_ ;
  assign \new_[167]_  = \new_[22667]_  & \new_[22654]_ ;
  assign \new_[168]_  = \new_[22643]_  & \new_[22630]_ ;
  assign \new_[169]_  = \new_[22619]_  & \new_[22606]_ ;
  assign \new_[170]_  = \new_[22595]_  & \new_[22582]_ ;
  assign \new_[171]_  = \new_[22571]_  & \new_[22558]_ ;
  assign \new_[172]_  = \new_[22547]_  & \new_[22534]_ ;
  assign \new_[173]_  = \new_[22523]_  & \new_[22510]_ ;
  assign \new_[174]_  = \new_[22499]_  & \new_[22486]_ ;
  assign \new_[175]_  = \new_[22475]_  & \new_[22462]_ ;
  assign \new_[176]_  = \new_[22451]_  & \new_[22438]_ ;
  assign \new_[177]_  = \new_[22427]_  & \new_[22414]_ ;
  assign \new_[178]_  = \new_[22403]_  & \new_[22390]_ ;
  assign \new_[179]_  = \new_[22379]_  & \new_[22366]_ ;
  assign \new_[180]_  = \new_[22355]_  & \new_[22342]_ ;
  assign \new_[181]_  = \new_[22331]_  & \new_[22318]_ ;
  assign \new_[182]_  = \new_[22307]_  & \new_[22294]_ ;
  assign \new_[183]_  = \new_[22283]_  & \new_[22270]_ ;
  assign \new_[184]_  = \new_[22259]_  & \new_[22246]_ ;
  assign \new_[185]_  = \new_[22235]_  & \new_[22222]_ ;
  assign \new_[186]_  = \new_[22211]_  & \new_[22198]_ ;
  assign \new_[187]_  = \new_[22187]_  & \new_[22174]_ ;
  assign \new_[188]_  = \new_[22163]_  & \new_[22150]_ ;
  assign \new_[189]_  = \new_[22139]_  & \new_[22126]_ ;
  assign \new_[190]_  = \new_[22115]_  & \new_[22102]_ ;
  assign \new_[191]_  = \new_[22091]_  & \new_[22078]_ ;
  assign \new_[192]_  = \new_[22067]_  & \new_[22054]_ ;
  assign \new_[193]_  = \new_[22043]_  & \new_[22030]_ ;
  assign \new_[194]_  = \new_[22019]_  & \new_[22006]_ ;
  assign \new_[195]_  = \new_[21995]_  & \new_[21982]_ ;
  assign \new_[196]_  = \new_[21971]_  & \new_[21958]_ ;
  assign \new_[197]_  = \new_[21947]_  & \new_[21934]_ ;
  assign \new_[198]_  = \new_[21923]_  & \new_[21910]_ ;
  assign \new_[199]_  = \new_[21899]_  & \new_[21886]_ ;
  assign \new_[200]_  = \new_[21875]_  & \new_[21862]_ ;
  assign \new_[201]_  = \new_[21851]_  & \new_[21838]_ ;
  assign \new_[202]_  = \new_[21827]_  & \new_[21814]_ ;
  assign \new_[203]_  = \new_[21803]_  & \new_[21790]_ ;
  assign \new_[204]_  = \new_[21779]_  & \new_[21766]_ ;
  assign \new_[205]_  = \new_[21755]_  & \new_[21742]_ ;
  assign \new_[206]_  = \new_[21731]_  & \new_[21718]_ ;
  assign \new_[207]_  = \new_[21707]_  & \new_[21694]_ ;
  assign \new_[208]_  = \new_[21683]_  & \new_[21670]_ ;
  assign \new_[209]_  = \new_[21659]_  & \new_[21646]_ ;
  assign \new_[210]_  = \new_[21635]_  & \new_[21622]_ ;
  assign \new_[211]_  = \new_[21611]_  & \new_[21598]_ ;
  assign \new_[212]_  = \new_[21587]_  & \new_[21574]_ ;
  assign \new_[213]_  = \new_[21563]_  & \new_[21550]_ ;
  assign \new_[214]_  = \new_[21539]_  & \new_[21526]_ ;
  assign \new_[215]_  = \new_[21515]_  & \new_[21502]_ ;
  assign \new_[216]_  = \new_[21491]_  & \new_[21478]_ ;
  assign \new_[217]_  = \new_[21467]_  & \new_[21454]_ ;
  assign \new_[218]_  = \new_[21443]_  & \new_[21430]_ ;
  assign \new_[219]_  = \new_[21419]_  & \new_[21406]_ ;
  assign \new_[220]_  = \new_[21395]_  & \new_[21382]_ ;
  assign \new_[221]_  = \new_[21371]_  & \new_[21358]_ ;
  assign \new_[222]_  = \new_[21347]_  & \new_[21334]_ ;
  assign \new_[223]_  = \new_[21323]_  & \new_[21310]_ ;
  assign \new_[224]_  = \new_[21299]_  & \new_[21286]_ ;
  assign \new_[225]_  = \new_[21275]_  & \new_[21262]_ ;
  assign \new_[226]_  = \new_[21251]_  & \new_[21238]_ ;
  assign \new_[227]_  = \new_[21227]_  & \new_[21214]_ ;
  assign \new_[228]_  = \new_[21203]_  & \new_[21190]_ ;
  assign \new_[229]_  = \new_[21179]_  & \new_[21166]_ ;
  assign \new_[230]_  = \new_[21155]_  & \new_[21142]_ ;
  assign \new_[231]_  = \new_[21131]_  & \new_[21118]_ ;
  assign \new_[232]_  = \new_[21107]_  & \new_[21094]_ ;
  assign \new_[233]_  = \new_[21083]_  & \new_[21070]_ ;
  assign \new_[234]_  = \new_[21059]_  & \new_[21046]_ ;
  assign \new_[235]_  = \new_[21035]_  & \new_[21022]_ ;
  assign \new_[236]_  = \new_[21011]_  & \new_[20998]_ ;
  assign \new_[237]_  = \new_[20987]_  & \new_[20974]_ ;
  assign \new_[238]_  = \new_[20963]_  & \new_[20950]_ ;
  assign \new_[239]_  = \new_[20939]_  & \new_[20926]_ ;
  assign \new_[240]_  = \new_[20915]_  & \new_[20902]_ ;
  assign \new_[241]_  = \new_[20891]_  & \new_[20878]_ ;
  assign \new_[242]_  = \new_[20867]_  & \new_[20854]_ ;
  assign \new_[243]_  = \new_[20843]_  & \new_[20830]_ ;
  assign \new_[244]_  = \new_[20819]_  & \new_[20806]_ ;
  assign \new_[245]_  = \new_[20795]_  & \new_[20782]_ ;
  assign \new_[246]_  = \new_[20771]_  & \new_[20758]_ ;
  assign \new_[247]_  = \new_[20747]_  & \new_[20734]_ ;
  assign \new_[248]_  = \new_[20723]_  & \new_[20710]_ ;
  assign \new_[249]_  = \new_[20699]_  & \new_[20686]_ ;
  assign \new_[250]_  = \new_[20675]_  & \new_[20662]_ ;
  assign \new_[251]_  = \new_[20651]_  & \new_[20638]_ ;
  assign \new_[252]_  = \new_[20627]_  & \new_[20614]_ ;
  assign \new_[253]_  = \new_[20603]_  & \new_[20590]_ ;
  assign \new_[254]_  = \new_[20579]_  & \new_[20566]_ ;
  assign \new_[255]_  = \new_[20555]_  & \new_[20542]_ ;
  assign \new_[256]_  = \new_[20531]_  & \new_[20518]_ ;
  assign \new_[257]_  = \new_[20507]_  & \new_[20494]_ ;
  assign \new_[258]_  = \new_[20483]_  & \new_[20470]_ ;
  assign \new_[259]_  = \new_[20459]_  & \new_[20446]_ ;
  assign \new_[260]_  = \new_[20435]_  & \new_[20422]_ ;
  assign \new_[261]_  = \new_[20411]_  & \new_[20398]_ ;
  assign \new_[262]_  = \new_[20387]_  & \new_[20374]_ ;
  assign \new_[263]_  = \new_[20363]_  & \new_[20350]_ ;
  assign \new_[264]_  = \new_[20339]_  & \new_[20326]_ ;
  assign \new_[265]_  = \new_[20315]_  & \new_[20302]_ ;
  assign \new_[266]_  = \new_[20291]_  & \new_[20278]_ ;
  assign \new_[267]_  = \new_[20267]_  & \new_[20254]_ ;
  assign \new_[268]_  = \new_[20243]_  & \new_[20230]_ ;
  assign \new_[269]_  = \new_[20219]_  & \new_[20206]_ ;
  assign \new_[270]_  = \new_[20195]_  & \new_[20182]_ ;
  assign \new_[271]_  = \new_[20171]_  & \new_[20158]_ ;
  assign \new_[272]_  = \new_[20147]_  & \new_[20134]_ ;
  assign \new_[273]_  = \new_[20123]_  & \new_[20110]_ ;
  assign \new_[274]_  = \new_[20099]_  & \new_[20086]_ ;
  assign \new_[275]_  = \new_[20075]_  & \new_[20062]_ ;
  assign \new_[276]_  = \new_[20051]_  & \new_[20038]_ ;
  assign \new_[277]_  = \new_[20027]_  & \new_[20014]_ ;
  assign \new_[278]_  = \new_[20003]_  & \new_[19990]_ ;
  assign \new_[279]_  = \new_[19979]_  & \new_[19966]_ ;
  assign \new_[280]_  = \new_[19955]_  & \new_[19942]_ ;
  assign \new_[281]_  = \new_[19931]_  & \new_[19918]_ ;
  assign \new_[282]_  = \new_[19907]_  & \new_[19894]_ ;
  assign \new_[283]_  = \new_[19883]_  & \new_[19870]_ ;
  assign \new_[284]_  = \new_[19859]_  & \new_[19846]_ ;
  assign \new_[285]_  = \new_[19835]_  & \new_[19822]_ ;
  assign \new_[286]_  = \new_[19811]_  & \new_[19798]_ ;
  assign \new_[287]_  = \new_[19787]_  & \new_[19774]_ ;
  assign \new_[288]_  = \new_[19763]_  & \new_[19750]_ ;
  assign \new_[289]_  = \new_[19739]_  & \new_[19726]_ ;
  assign \new_[290]_  = \new_[19715]_  & \new_[19702]_ ;
  assign \new_[291]_  = \new_[19691]_  & \new_[19678]_ ;
  assign \new_[292]_  = \new_[19667]_  & \new_[19654]_ ;
  assign \new_[293]_  = \new_[19643]_  & \new_[19630]_ ;
  assign \new_[294]_  = \new_[19619]_  & \new_[19606]_ ;
  assign \new_[295]_  = \new_[19595]_  & \new_[19582]_ ;
  assign \new_[296]_  = \new_[19571]_  & \new_[19558]_ ;
  assign \new_[297]_  = \new_[19547]_  & \new_[19534]_ ;
  assign \new_[298]_  = \new_[19523]_  & \new_[19510]_ ;
  assign \new_[299]_  = \new_[19499]_  & \new_[19486]_ ;
  assign \new_[300]_  = \new_[19475]_  & \new_[19462]_ ;
  assign \new_[301]_  = \new_[19451]_  & \new_[19438]_ ;
  assign \new_[302]_  = \new_[19427]_  & \new_[19414]_ ;
  assign \new_[303]_  = \new_[19403]_  & \new_[19390]_ ;
  assign \new_[304]_  = \new_[19379]_  & \new_[19366]_ ;
  assign \new_[305]_  = \new_[19355]_  & \new_[19342]_ ;
  assign \new_[306]_  = \new_[19331]_  & \new_[19318]_ ;
  assign \new_[307]_  = \new_[19307]_  & \new_[19294]_ ;
  assign \new_[308]_  = \new_[19283]_  & \new_[19270]_ ;
  assign \new_[309]_  = \new_[19259]_  & \new_[19246]_ ;
  assign \new_[310]_  = \new_[19235]_  & \new_[19222]_ ;
  assign \new_[311]_  = \new_[19211]_  & \new_[19198]_ ;
  assign \new_[312]_  = \new_[19187]_  & \new_[19174]_ ;
  assign \new_[313]_  = \new_[19163]_  & \new_[19150]_ ;
  assign \new_[314]_  = \new_[19139]_  & \new_[19126]_ ;
  assign \new_[315]_  = \new_[19115]_  & \new_[19102]_ ;
  assign \new_[316]_  = \new_[19091]_  & \new_[19078]_ ;
  assign \new_[317]_  = \new_[19067]_  & \new_[19054]_ ;
  assign \new_[318]_  = \new_[19043]_  & \new_[19030]_ ;
  assign \new_[319]_  = \new_[19019]_  & \new_[19008]_ ;
  assign \new_[320]_  = \new_[18997]_  & \new_[18986]_ ;
  assign \new_[321]_  = \new_[18975]_  & \new_[18964]_ ;
  assign \new_[322]_  = \new_[18953]_  & \new_[18942]_ ;
  assign \new_[323]_  = \new_[18931]_  & \new_[18920]_ ;
  assign \new_[324]_  = \new_[18909]_  & \new_[18898]_ ;
  assign \new_[325]_  = \new_[18887]_  & \new_[18876]_ ;
  assign \new_[326]_  = \new_[18865]_  & \new_[18854]_ ;
  assign \new_[327]_  = \new_[18843]_  & \new_[18832]_ ;
  assign \new_[328]_  = \new_[18821]_  & \new_[18810]_ ;
  assign \new_[329]_  = \new_[18799]_  & \new_[18788]_ ;
  assign \new_[330]_  = \new_[18777]_  & \new_[18766]_ ;
  assign \new_[331]_  = \new_[18755]_  & \new_[18744]_ ;
  assign \new_[332]_  = \new_[18733]_  & \new_[18722]_ ;
  assign \new_[333]_  = \new_[18711]_  & \new_[18700]_ ;
  assign \new_[334]_  = \new_[18689]_  & \new_[18678]_ ;
  assign \new_[335]_  = \new_[18667]_  & \new_[18656]_ ;
  assign \new_[336]_  = \new_[18645]_  & \new_[18634]_ ;
  assign \new_[337]_  = \new_[18623]_  & \new_[18612]_ ;
  assign \new_[338]_  = \new_[18601]_  & \new_[18590]_ ;
  assign \new_[339]_  = \new_[18579]_  & \new_[18568]_ ;
  assign \new_[340]_  = \new_[18557]_  & \new_[18546]_ ;
  assign \new_[341]_  = \new_[18535]_  & \new_[18524]_ ;
  assign \new_[342]_  = \new_[18513]_  & \new_[18502]_ ;
  assign \new_[343]_  = \new_[18491]_  & \new_[18480]_ ;
  assign \new_[344]_  = \new_[18469]_  & \new_[18458]_ ;
  assign \new_[345]_  = \new_[18447]_  & \new_[18436]_ ;
  assign \new_[346]_  = \new_[18425]_  & \new_[18414]_ ;
  assign \new_[347]_  = \new_[18403]_  & \new_[18392]_ ;
  assign \new_[348]_  = \new_[18381]_  & \new_[18370]_ ;
  assign \new_[349]_  = \new_[18359]_  & \new_[18348]_ ;
  assign \new_[350]_  = \new_[18337]_  & \new_[18326]_ ;
  assign \new_[351]_  = \new_[18315]_  & \new_[18304]_ ;
  assign \new_[352]_  = \new_[18293]_  & \new_[18282]_ ;
  assign \new_[353]_  = \new_[18271]_  & \new_[18260]_ ;
  assign \new_[354]_  = \new_[18249]_  & \new_[18238]_ ;
  assign \new_[355]_  = \new_[18227]_  & \new_[18216]_ ;
  assign \new_[356]_  = \new_[18205]_  & \new_[18194]_ ;
  assign \new_[357]_  = \new_[18183]_  & \new_[18172]_ ;
  assign \new_[358]_  = \new_[18161]_  & \new_[18150]_ ;
  assign \new_[359]_  = \new_[18139]_  & \new_[18128]_ ;
  assign \new_[360]_  = \new_[18117]_  & \new_[18106]_ ;
  assign \new_[361]_  = \new_[18095]_  & \new_[18084]_ ;
  assign \new_[362]_  = \new_[18073]_  & \new_[18062]_ ;
  assign \new_[363]_  = \new_[18051]_  & \new_[18040]_ ;
  assign \new_[364]_  = \new_[18029]_  & \new_[18018]_ ;
  assign \new_[365]_  = \new_[18007]_  & \new_[17996]_ ;
  assign \new_[366]_  = \new_[17985]_  & \new_[17974]_ ;
  assign \new_[367]_  = \new_[17963]_  & \new_[17952]_ ;
  assign \new_[368]_  = \new_[17941]_  & \new_[17930]_ ;
  assign \new_[369]_  = \new_[17919]_  & \new_[17908]_ ;
  assign \new_[370]_  = \new_[17897]_  & \new_[17886]_ ;
  assign \new_[371]_  = \new_[17875]_  & \new_[17864]_ ;
  assign \new_[372]_  = \new_[17853]_  & \new_[17842]_ ;
  assign \new_[373]_  = \new_[17831]_  & \new_[17820]_ ;
  assign \new_[374]_  = \new_[17809]_  & \new_[17798]_ ;
  assign \new_[375]_  = \new_[17787]_  & \new_[17776]_ ;
  assign \new_[376]_  = \new_[17765]_  & \new_[17754]_ ;
  assign \new_[377]_  = \new_[17743]_  & \new_[17732]_ ;
  assign \new_[378]_  = \new_[17721]_  & \new_[17710]_ ;
  assign \new_[379]_  = \new_[17699]_  & \new_[17688]_ ;
  assign \new_[380]_  = \new_[17677]_  & \new_[17666]_ ;
  assign \new_[381]_  = \new_[17655]_  & \new_[17644]_ ;
  assign \new_[382]_  = \new_[17633]_  & \new_[17622]_ ;
  assign \new_[383]_  = \new_[17611]_  & \new_[17600]_ ;
  assign \new_[384]_  = \new_[17589]_  & \new_[17578]_ ;
  assign \new_[385]_  = \new_[17567]_  & \new_[17556]_ ;
  assign \new_[386]_  = \new_[17545]_  & \new_[17534]_ ;
  assign \new_[387]_  = \new_[17523]_  & \new_[17512]_ ;
  assign \new_[388]_  = \new_[17501]_  & \new_[17490]_ ;
  assign \new_[389]_  = \new_[17479]_  & \new_[17468]_ ;
  assign \new_[390]_  = \new_[17457]_  & \new_[17446]_ ;
  assign \new_[391]_  = \new_[17435]_  & \new_[17424]_ ;
  assign \new_[392]_  = \new_[17413]_  & \new_[17402]_ ;
  assign \new_[393]_  = \new_[17391]_  & \new_[17380]_ ;
  assign \new_[394]_  = \new_[17369]_  & \new_[17358]_ ;
  assign \new_[395]_  = \new_[17347]_  & \new_[17336]_ ;
  assign \new_[396]_  = \new_[17325]_  & \new_[17314]_ ;
  assign \new_[397]_  = \new_[17303]_  & \new_[17292]_ ;
  assign \new_[398]_  = \new_[17281]_  & \new_[17270]_ ;
  assign \new_[399]_  = \new_[17259]_  & \new_[17248]_ ;
  assign \new_[400]_  = \new_[17237]_  & \new_[17226]_ ;
  assign \new_[401]_  = \new_[17215]_  & \new_[17204]_ ;
  assign \new_[402]_  = \new_[17193]_  & \new_[17182]_ ;
  assign \new_[403]_  = \new_[17171]_  & \new_[17160]_ ;
  assign \new_[404]_  = \new_[17149]_  & \new_[17138]_ ;
  assign \new_[405]_  = \new_[17127]_  & \new_[17116]_ ;
  assign \new_[406]_  = \new_[17105]_  & \new_[17094]_ ;
  assign \new_[407]_  = \new_[17083]_  & \new_[17072]_ ;
  assign \new_[408]_  = \new_[17061]_  & \new_[17050]_ ;
  assign \new_[409]_  = \new_[17039]_  & \new_[17028]_ ;
  assign \new_[410]_  = \new_[17017]_  & \new_[17006]_ ;
  assign \new_[411]_  = \new_[16995]_  & \new_[16984]_ ;
  assign \new_[412]_  = \new_[16973]_  & \new_[16962]_ ;
  assign \new_[413]_  = \new_[16951]_  & \new_[16940]_ ;
  assign \new_[414]_  = \new_[16929]_  & \new_[16918]_ ;
  assign \new_[415]_  = \new_[16907]_  & \new_[16896]_ ;
  assign \new_[416]_  = \new_[16885]_  & \new_[16874]_ ;
  assign \new_[417]_  = \new_[16863]_  & \new_[16852]_ ;
  assign \new_[418]_  = \new_[16841]_  & \new_[16830]_ ;
  assign \new_[419]_  = \new_[16819]_  & \new_[16808]_ ;
  assign \new_[420]_  = \new_[16797]_  & \new_[16786]_ ;
  assign \new_[421]_  = \new_[16775]_  & \new_[16764]_ ;
  assign \new_[422]_  = \new_[16753]_  & \new_[16742]_ ;
  assign \new_[423]_  = \new_[16731]_  & \new_[16720]_ ;
  assign \new_[424]_  = \new_[16709]_  & \new_[16698]_ ;
  assign \new_[425]_  = \new_[16687]_  & \new_[16676]_ ;
  assign \new_[426]_  = \new_[16665]_  & \new_[16654]_ ;
  assign \new_[427]_  = \new_[16643]_  & \new_[16632]_ ;
  assign \new_[428]_  = \new_[16621]_  & \new_[16610]_ ;
  assign \new_[429]_  = \new_[16599]_  & \new_[16588]_ ;
  assign \new_[430]_  = \new_[16577]_  & \new_[16566]_ ;
  assign \new_[431]_  = \new_[16555]_  & \new_[16544]_ ;
  assign \new_[432]_  = \new_[16533]_  & \new_[16522]_ ;
  assign \new_[433]_  = \new_[16511]_  & \new_[16500]_ ;
  assign \new_[434]_  = \new_[16489]_  & \new_[16478]_ ;
  assign \new_[435]_  = \new_[16467]_  & \new_[16456]_ ;
  assign \new_[436]_  = \new_[16445]_  & \new_[16434]_ ;
  assign \new_[437]_  = \new_[16423]_  & \new_[16412]_ ;
  assign \new_[438]_  = \new_[16401]_  & \new_[16390]_ ;
  assign \new_[439]_  = \new_[16379]_  & \new_[16368]_ ;
  assign \new_[440]_  = \new_[16357]_  & \new_[16346]_ ;
  assign \new_[441]_  = \new_[16335]_  & \new_[16324]_ ;
  assign \new_[442]_  = \new_[16313]_  & \new_[16302]_ ;
  assign \new_[443]_  = \new_[16291]_  & \new_[16280]_ ;
  assign \new_[444]_  = \new_[16269]_  & \new_[16258]_ ;
  assign \new_[445]_  = \new_[16247]_  & \new_[16236]_ ;
  assign \new_[446]_  = \new_[16225]_  & \new_[16214]_ ;
  assign \new_[447]_  = \new_[16203]_  & \new_[16192]_ ;
  assign \new_[448]_  = \new_[16181]_  & \new_[16170]_ ;
  assign \new_[449]_  = \new_[16159]_  & \new_[16148]_ ;
  assign \new_[450]_  = \new_[16137]_  & \new_[16126]_ ;
  assign \new_[451]_  = \new_[16115]_  & \new_[16104]_ ;
  assign \new_[452]_  = \new_[16093]_  & \new_[16082]_ ;
  assign \new_[453]_  = \new_[16071]_  & \new_[16060]_ ;
  assign \new_[454]_  = \new_[16049]_  & \new_[16038]_ ;
  assign \new_[455]_  = \new_[16027]_  & \new_[16016]_ ;
  assign \new_[456]_  = \new_[16005]_  & \new_[15994]_ ;
  assign \new_[457]_  = \new_[15983]_  & \new_[15972]_ ;
  assign \new_[458]_  = \new_[15961]_  & \new_[15950]_ ;
  assign \new_[459]_  = \new_[15939]_  & \new_[15928]_ ;
  assign \new_[460]_  = \new_[15917]_  & \new_[15906]_ ;
  assign \new_[461]_  = \new_[15895]_  & \new_[15884]_ ;
  assign \new_[462]_  = \new_[15873]_  & \new_[15862]_ ;
  assign \new_[463]_  = \new_[15851]_  & \new_[15840]_ ;
  assign \new_[464]_  = \new_[15829]_  & \new_[15818]_ ;
  assign \new_[465]_  = \new_[15807]_  & \new_[15796]_ ;
  assign \new_[466]_  = \new_[15785]_  & \new_[15774]_ ;
  assign \new_[467]_  = \new_[15763]_  & \new_[15752]_ ;
  assign \new_[468]_  = \new_[15741]_  & \new_[15730]_ ;
  assign \new_[469]_  = \new_[15719]_  & \new_[15708]_ ;
  assign \new_[470]_  = \new_[15697]_  & \new_[15686]_ ;
  assign \new_[471]_  = \new_[15675]_  & \new_[15664]_ ;
  assign \new_[472]_  = \new_[15653]_  & \new_[15642]_ ;
  assign \new_[473]_  = \new_[15631]_  & \new_[15620]_ ;
  assign \new_[474]_  = \new_[15609]_  & \new_[15598]_ ;
  assign \new_[475]_  = \new_[15587]_  & \new_[15576]_ ;
  assign \new_[476]_  = \new_[15565]_  & \new_[15554]_ ;
  assign \new_[477]_  = \new_[15543]_  & \new_[15532]_ ;
  assign \new_[478]_  = \new_[15521]_  & \new_[15510]_ ;
  assign \new_[479]_  = \new_[15499]_  & \new_[15488]_ ;
  assign \new_[480]_  = \new_[15477]_  & \new_[15466]_ ;
  assign \new_[481]_  = \new_[15455]_  & \new_[15444]_ ;
  assign \new_[482]_  = \new_[15433]_  & \new_[15422]_ ;
  assign \new_[483]_  = \new_[15411]_  & \new_[15400]_ ;
  assign \new_[484]_  = \new_[15389]_  & \new_[15378]_ ;
  assign \new_[485]_  = \new_[15367]_  & \new_[15356]_ ;
  assign \new_[486]_  = \new_[15345]_  & \new_[15334]_ ;
  assign \new_[487]_  = \new_[15323]_  & \new_[15312]_ ;
  assign \new_[488]_  = \new_[15301]_  & \new_[15290]_ ;
  assign \new_[489]_  = \new_[15279]_  & \new_[15268]_ ;
  assign \new_[490]_  = \new_[15257]_  & \new_[15246]_ ;
  assign \new_[491]_  = \new_[15235]_  & \new_[15224]_ ;
  assign \new_[492]_  = \new_[15213]_  & \new_[15202]_ ;
  assign \new_[493]_  = \new_[15191]_  & \new_[15180]_ ;
  assign \new_[494]_  = \new_[15169]_  & \new_[15158]_ ;
  assign \new_[495]_  = \new_[15147]_  & \new_[15136]_ ;
  assign \new_[496]_  = \new_[15125]_  & \new_[15114]_ ;
  assign \new_[497]_  = \new_[15103]_  & \new_[15092]_ ;
  assign \new_[498]_  = \new_[15081]_  & \new_[15070]_ ;
  assign \new_[499]_  = \new_[15059]_  & \new_[15048]_ ;
  assign \new_[500]_  = \new_[15037]_  & \new_[15026]_ ;
  assign \new_[501]_  = \new_[15015]_  & \new_[15004]_ ;
  assign \new_[502]_  = \new_[14993]_  & \new_[14982]_ ;
  assign \new_[503]_  = \new_[14971]_  & \new_[14960]_ ;
  assign \new_[504]_  = \new_[14949]_  & \new_[14938]_ ;
  assign \new_[505]_  = \new_[14927]_  & \new_[14916]_ ;
  assign \new_[506]_  = \new_[14905]_  & \new_[14894]_ ;
  assign \new_[507]_  = \new_[14883]_  & \new_[14872]_ ;
  assign \new_[508]_  = \new_[14861]_  & \new_[14850]_ ;
  assign \new_[509]_  = \new_[14839]_  & \new_[14828]_ ;
  assign \new_[510]_  = \new_[14817]_  & \new_[14806]_ ;
  assign \new_[511]_  = \new_[14795]_  & \new_[14784]_ ;
  assign \new_[512]_  = \new_[14773]_  & \new_[14762]_ ;
  assign \new_[513]_  = \new_[14751]_  & \new_[14740]_ ;
  assign \new_[514]_  = \new_[14729]_  & \new_[14718]_ ;
  assign \new_[515]_  = \new_[14707]_  & \new_[14696]_ ;
  assign \new_[516]_  = \new_[14685]_  & \new_[14674]_ ;
  assign \new_[517]_  = \new_[14663]_  & \new_[14652]_ ;
  assign \new_[518]_  = \new_[14641]_  & \new_[14630]_ ;
  assign \new_[519]_  = \new_[14619]_  & \new_[14608]_ ;
  assign \new_[520]_  = \new_[14597]_  & \new_[14586]_ ;
  assign \new_[521]_  = \new_[14575]_  & \new_[14564]_ ;
  assign \new_[522]_  = \new_[14553]_  & \new_[14542]_ ;
  assign \new_[523]_  = \new_[14531]_  & \new_[14520]_ ;
  assign \new_[524]_  = \new_[14509]_  & \new_[14498]_ ;
  assign \new_[525]_  = \new_[14487]_  & \new_[14476]_ ;
  assign \new_[526]_  = \new_[14465]_  & \new_[14454]_ ;
  assign \new_[527]_  = \new_[14443]_  & \new_[14432]_ ;
  assign \new_[528]_  = \new_[14421]_  & \new_[14410]_ ;
  assign \new_[529]_  = \new_[14399]_  & \new_[14388]_ ;
  assign \new_[530]_  = \new_[14377]_  & \new_[14366]_ ;
  assign \new_[531]_  = \new_[14355]_  & \new_[14344]_ ;
  assign \new_[532]_  = \new_[14333]_  & \new_[14322]_ ;
  assign \new_[533]_  = \new_[14311]_  & \new_[14300]_ ;
  assign \new_[534]_  = \new_[14289]_  & \new_[14278]_ ;
  assign \new_[535]_  = \new_[14267]_  & \new_[14256]_ ;
  assign \new_[536]_  = \new_[14245]_  & \new_[14234]_ ;
  assign \new_[537]_  = \new_[14223]_  & \new_[14212]_ ;
  assign \new_[538]_  = \new_[14201]_  & \new_[14190]_ ;
  assign \new_[539]_  = \new_[14179]_  & \new_[14168]_ ;
  assign \new_[540]_  = \new_[14157]_  & \new_[14146]_ ;
  assign \new_[541]_  = \new_[14135]_  & \new_[14124]_ ;
  assign \new_[542]_  = \new_[14113]_  & \new_[14102]_ ;
  assign \new_[543]_  = \new_[14091]_  & \new_[14080]_ ;
  assign \new_[544]_  = \new_[14069]_  & \new_[14058]_ ;
  assign \new_[545]_  = \new_[14047]_  & \new_[14036]_ ;
  assign \new_[546]_  = \new_[14025]_  & \new_[14014]_ ;
  assign \new_[547]_  = \new_[14003]_  & \new_[13992]_ ;
  assign \new_[548]_  = \new_[13981]_  & \new_[13970]_ ;
  assign \new_[549]_  = \new_[13959]_  & \new_[13948]_ ;
  assign \new_[550]_  = \new_[13937]_  & \new_[13926]_ ;
  assign \new_[551]_  = \new_[13915]_  & \new_[13904]_ ;
  assign \new_[552]_  = \new_[13893]_  & \new_[13882]_ ;
  assign \new_[553]_  = \new_[13871]_  & \new_[13860]_ ;
  assign \new_[554]_  = \new_[13849]_  & \new_[13838]_ ;
  assign \new_[555]_  = \new_[13827]_  & \new_[13816]_ ;
  assign \new_[556]_  = \new_[13805]_  & \new_[13794]_ ;
  assign \new_[557]_  = \new_[13783]_  & \new_[13772]_ ;
  assign \new_[558]_  = \new_[13761]_  & \new_[13750]_ ;
  assign \new_[559]_  = \new_[13739]_  & \new_[13728]_ ;
  assign \new_[560]_  = \new_[13717]_  & \new_[13706]_ ;
  assign \new_[561]_  = \new_[13695]_  & \new_[13684]_ ;
  assign \new_[562]_  = \new_[13673]_  & \new_[13662]_ ;
  assign \new_[563]_  = \new_[13651]_  & \new_[13640]_ ;
  assign \new_[564]_  = \new_[13629]_  & \new_[13618]_ ;
  assign \new_[565]_  = \new_[13607]_  & \new_[13596]_ ;
  assign \new_[566]_  = \new_[13585]_  & \new_[13574]_ ;
  assign \new_[567]_  = \new_[13563]_  & \new_[13552]_ ;
  assign \new_[568]_  = \new_[13541]_  & \new_[13530]_ ;
  assign \new_[569]_  = \new_[13519]_  & \new_[13508]_ ;
  assign \new_[570]_  = \new_[13497]_  & \new_[13486]_ ;
  assign \new_[571]_  = \new_[13475]_  & \new_[13464]_ ;
  assign \new_[572]_  = \new_[13453]_  & \new_[13442]_ ;
  assign \new_[573]_  = \new_[13431]_  & \new_[13420]_ ;
  assign \new_[574]_  = \new_[13409]_  & \new_[13398]_ ;
  assign \new_[575]_  = \new_[13387]_  & \new_[13376]_ ;
  assign \new_[576]_  = \new_[13365]_  & \new_[13354]_ ;
  assign \new_[577]_  = \new_[13343]_  & \new_[13332]_ ;
  assign \new_[578]_  = \new_[13321]_  & \new_[13310]_ ;
  assign \new_[579]_  = \new_[13299]_  & \new_[13288]_ ;
  assign \new_[580]_  = \new_[13277]_  & \new_[13266]_ ;
  assign \new_[581]_  = \new_[13255]_  & \new_[13244]_ ;
  assign \new_[582]_  = \new_[13233]_  & \new_[13222]_ ;
  assign \new_[583]_  = \new_[13211]_  & \new_[13200]_ ;
  assign \new_[584]_  = \new_[13189]_  & \new_[13178]_ ;
  assign \new_[585]_  = \new_[13167]_  & \new_[13156]_ ;
  assign \new_[586]_  = \new_[13145]_  & \new_[13134]_ ;
  assign \new_[587]_  = \new_[13123]_  & \new_[13112]_ ;
  assign \new_[588]_  = \new_[13101]_  & \new_[13090]_ ;
  assign \new_[589]_  = \new_[13079]_  & \new_[13068]_ ;
  assign \new_[590]_  = \new_[13057]_  & \new_[13046]_ ;
  assign \new_[591]_  = \new_[13035]_  & \new_[13024]_ ;
  assign \new_[592]_  = \new_[13013]_  & \new_[13002]_ ;
  assign \new_[593]_  = \new_[12991]_  & \new_[12980]_ ;
  assign \new_[594]_  = \new_[12969]_  & \new_[12958]_ ;
  assign \new_[595]_  = \new_[12947]_  & \new_[12936]_ ;
  assign \new_[596]_  = \new_[12925]_  & \new_[12914]_ ;
  assign \new_[597]_  = \new_[12903]_  & \new_[12892]_ ;
  assign \new_[598]_  = \new_[12881]_  & \new_[12870]_ ;
  assign \new_[599]_  = \new_[12859]_  & \new_[12848]_ ;
  assign \new_[600]_  = \new_[12837]_  & \new_[12826]_ ;
  assign \new_[601]_  = \new_[12815]_  & \new_[12804]_ ;
  assign \new_[602]_  = \new_[12793]_  & \new_[12782]_ ;
  assign \new_[603]_  = \new_[12771]_  & \new_[12760]_ ;
  assign \new_[604]_  = \new_[12749]_  & \new_[12738]_ ;
  assign \new_[605]_  = \new_[12727]_  & \new_[12716]_ ;
  assign \new_[606]_  = \new_[12705]_  & \new_[12694]_ ;
  assign \new_[607]_  = \new_[12683]_  & \new_[12672]_ ;
  assign \new_[608]_  = \new_[12661]_  & \new_[12650]_ ;
  assign \new_[609]_  = \new_[12639]_  & \new_[12628]_ ;
  assign \new_[610]_  = \new_[12617]_  & \new_[12606]_ ;
  assign \new_[611]_  = \new_[12595]_  & \new_[12584]_ ;
  assign \new_[612]_  = \new_[12573]_  & \new_[12562]_ ;
  assign \new_[613]_  = \new_[12551]_  & \new_[12540]_ ;
  assign \new_[614]_  = \new_[12529]_  & \new_[12518]_ ;
  assign \new_[615]_  = \new_[12507]_  & \new_[12496]_ ;
  assign \new_[616]_  = \new_[12485]_  & \new_[12474]_ ;
  assign \new_[617]_  = \new_[12463]_  & \new_[12452]_ ;
  assign \new_[618]_  = \new_[12441]_  & \new_[12430]_ ;
  assign \new_[619]_  = \new_[12419]_  & \new_[12408]_ ;
  assign \new_[620]_  = \new_[12397]_  & \new_[12386]_ ;
  assign \new_[621]_  = \new_[12375]_  & \new_[12364]_ ;
  assign \new_[622]_  = \new_[12353]_  & \new_[12342]_ ;
  assign \new_[623]_  = \new_[12331]_  & \new_[12320]_ ;
  assign \new_[624]_  = \new_[12309]_  & \new_[12298]_ ;
  assign \new_[625]_  = \new_[12287]_  & \new_[12276]_ ;
  assign \new_[626]_  = \new_[12265]_  & \new_[12254]_ ;
  assign \new_[627]_  = \new_[12243]_  & \new_[12232]_ ;
  assign \new_[628]_  = \new_[12221]_  & \new_[12210]_ ;
  assign \new_[629]_  = \new_[12201]_  & \new_[12190]_ ;
  assign \new_[630]_  = \new_[12181]_  & \new_[12170]_ ;
  assign \new_[631]_  = \new_[12161]_  & \new_[12150]_ ;
  assign \new_[632]_  = \new_[12141]_  & \new_[12130]_ ;
  assign \new_[633]_  = \new_[12121]_  & \new_[12110]_ ;
  assign \new_[634]_  = \new_[12101]_  & \new_[12090]_ ;
  assign \new_[635]_  = \new_[12081]_  & \new_[12070]_ ;
  assign \new_[636]_  = \new_[12061]_  & \new_[12050]_ ;
  assign \new_[637]_  = \new_[12041]_  & \new_[12030]_ ;
  assign \new_[638]_  = \new_[12021]_  & \new_[12010]_ ;
  assign \new_[639]_  = \new_[12001]_  & \new_[11990]_ ;
  assign \new_[640]_  = \new_[11981]_  & \new_[11970]_ ;
  assign \new_[641]_  = \new_[11961]_  & \new_[11950]_ ;
  assign \new_[642]_  = \new_[11941]_  & \new_[11930]_ ;
  assign \new_[643]_  = \new_[11921]_  & \new_[11910]_ ;
  assign \new_[644]_  = \new_[11901]_  & \new_[11890]_ ;
  assign \new_[645]_  = \new_[11881]_  & \new_[11870]_ ;
  assign \new_[646]_  = \new_[11861]_  & \new_[11850]_ ;
  assign \new_[647]_  = \new_[11841]_  & \new_[11830]_ ;
  assign \new_[648]_  = \new_[11821]_  & \new_[11810]_ ;
  assign \new_[649]_  = \new_[11801]_  & \new_[11790]_ ;
  assign \new_[650]_  = \new_[11781]_  & \new_[11770]_ ;
  assign \new_[651]_  = \new_[11761]_  & \new_[11750]_ ;
  assign \new_[652]_  = \new_[11741]_  & \new_[11730]_ ;
  assign \new_[653]_  = \new_[11721]_  & \new_[11710]_ ;
  assign \new_[654]_  = \new_[11701]_  & \new_[11690]_ ;
  assign \new_[655]_  = \new_[11681]_  & \new_[11670]_ ;
  assign \new_[656]_  = \new_[11661]_  & \new_[11650]_ ;
  assign \new_[657]_  = \new_[11641]_  & \new_[11630]_ ;
  assign \new_[658]_  = \new_[11621]_  & \new_[11610]_ ;
  assign \new_[659]_  = \new_[11601]_  & \new_[11590]_ ;
  assign \new_[660]_  = \new_[11581]_  & \new_[11570]_ ;
  assign \new_[661]_  = \new_[11561]_  & \new_[11550]_ ;
  assign \new_[662]_  = \new_[11541]_  & \new_[11530]_ ;
  assign \new_[663]_  = \new_[11521]_  & \new_[11510]_ ;
  assign \new_[664]_  = \new_[11501]_  & \new_[11490]_ ;
  assign \new_[665]_  = \new_[11481]_  & \new_[11470]_ ;
  assign \new_[666]_  = \new_[11461]_  & \new_[11450]_ ;
  assign \new_[667]_  = \new_[11441]_  & \new_[11430]_ ;
  assign \new_[668]_  = \new_[11421]_  & \new_[11410]_ ;
  assign \new_[669]_  = \new_[11401]_  & \new_[11390]_ ;
  assign \new_[670]_  = \new_[11381]_  & \new_[11370]_ ;
  assign \new_[671]_  = \new_[11361]_  & \new_[11350]_ ;
  assign \new_[672]_  = \new_[11341]_  & \new_[11330]_ ;
  assign \new_[673]_  = \new_[11321]_  & \new_[11310]_ ;
  assign \new_[674]_  = \new_[11301]_  & \new_[11290]_ ;
  assign \new_[675]_  = \new_[11281]_  & \new_[11270]_ ;
  assign \new_[676]_  = \new_[11261]_  & \new_[11250]_ ;
  assign \new_[677]_  = \new_[11241]_  & \new_[11230]_ ;
  assign \new_[678]_  = \new_[11221]_  & \new_[11210]_ ;
  assign \new_[679]_  = \new_[11201]_  & \new_[11190]_ ;
  assign \new_[680]_  = \new_[11181]_  & \new_[11170]_ ;
  assign \new_[681]_  = \new_[11161]_  & \new_[11150]_ ;
  assign \new_[682]_  = \new_[11141]_  & \new_[11130]_ ;
  assign \new_[683]_  = \new_[11121]_  & \new_[11110]_ ;
  assign \new_[684]_  = \new_[11101]_  & \new_[11090]_ ;
  assign \new_[685]_  = \new_[11081]_  & \new_[11070]_ ;
  assign \new_[686]_  = \new_[11061]_  & \new_[11050]_ ;
  assign \new_[687]_  = \new_[11041]_  & \new_[11030]_ ;
  assign \new_[688]_  = \new_[11021]_  & \new_[11010]_ ;
  assign \new_[689]_  = \new_[11001]_  & \new_[10990]_ ;
  assign \new_[690]_  = \new_[10981]_  & \new_[10970]_ ;
  assign \new_[691]_  = \new_[10961]_  & \new_[10950]_ ;
  assign \new_[692]_  = \new_[10941]_  & \new_[10930]_ ;
  assign \new_[693]_  = \new_[10921]_  & \new_[10910]_ ;
  assign \new_[694]_  = \new_[10901]_  & \new_[10890]_ ;
  assign \new_[695]_  = \new_[10881]_  & \new_[10870]_ ;
  assign \new_[696]_  = \new_[10861]_  & \new_[10850]_ ;
  assign \new_[697]_  = \new_[10841]_  & \new_[10830]_ ;
  assign \new_[698]_  = \new_[10821]_  & \new_[10810]_ ;
  assign \new_[699]_  = \new_[10801]_  & \new_[10790]_ ;
  assign \new_[700]_  = \new_[10781]_  & \new_[10770]_ ;
  assign \new_[701]_  = \new_[10761]_  & \new_[10750]_ ;
  assign \new_[702]_  = \new_[10741]_  & \new_[10730]_ ;
  assign \new_[703]_  = \new_[10721]_  & \new_[10710]_ ;
  assign \new_[704]_  = \new_[10701]_  & \new_[10690]_ ;
  assign \new_[705]_  = \new_[10681]_  & \new_[10670]_ ;
  assign \new_[706]_  = \new_[10661]_  & \new_[10650]_ ;
  assign \new_[707]_  = \new_[10641]_  & \new_[10630]_ ;
  assign \new_[708]_  = \new_[10621]_  & \new_[10610]_ ;
  assign \new_[709]_  = \new_[10601]_  & \new_[10590]_ ;
  assign \new_[710]_  = \new_[10581]_  & \new_[10570]_ ;
  assign \new_[711]_  = \new_[10561]_  & \new_[10550]_ ;
  assign \new_[712]_  = \new_[10541]_  & \new_[10530]_ ;
  assign \new_[713]_  = \new_[10521]_  & \new_[10510]_ ;
  assign \new_[714]_  = \new_[10501]_  & \new_[10490]_ ;
  assign \new_[715]_  = \new_[10481]_  & \new_[10470]_ ;
  assign \new_[716]_  = \new_[10461]_  & \new_[10450]_ ;
  assign \new_[717]_  = \new_[10441]_  & \new_[10430]_ ;
  assign \new_[718]_  = \new_[10421]_  & \new_[10410]_ ;
  assign \new_[719]_  = \new_[10401]_  & \new_[10390]_ ;
  assign \new_[720]_  = \new_[10381]_  & \new_[10370]_ ;
  assign \new_[721]_  = \new_[10361]_  & \new_[10350]_ ;
  assign \new_[722]_  = \new_[10341]_  & \new_[10330]_ ;
  assign \new_[723]_  = \new_[10321]_  & \new_[10310]_ ;
  assign \new_[724]_  = \new_[10301]_  & \new_[10290]_ ;
  assign \new_[725]_  = \new_[10281]_  & \new_[10270]_ ;
  assign \new_[726]_  = \new_[10261]_  & \new_[10250]_ ;
  assign \new_[727]_  = \new_[10241]_  & \new_[10230]_ ;
  assign \new_[728]_  = \new_[10221]_  & \new_[10210]_ ;
  assign \new_[729]_  = \new_[10201]_  & \new_[10190]_ ;
  assign \new_[730]_  = \new_[10181]_  & \new_[10170]_ ;
  assign \new_[731]_  = \new_[10161]_  & \new_[10150]_ ;
  assign \new_[732]_  = \new_[10141]_  & \new_[10130]_ ;
  assign \new_[733]_  = \new_[10121]_  & \new_[10110]_ ;
  assign \new_[734]_  = \new_[10101]_  & \new_[10090]_ ;
  assign \new_[735]_  = \new_[10081]_  & \new_[10070]_ ;
  assign \new_[736]_  = \new_[10061]_  & \new_[10050]_ ;
  assign \new_[737]_  = \new_[10041]_  & \new_[10030]_ ;
  assign \new_[738]_  = \new_[10021]_  & \new_[10010]_ ;
  assign \new_[739]_  = \new_[10001]_  & \new_[9990]_ ;
  assign \new_[740]_  = \new_[9981]_  & \new_[9970]_ ;
  assign \new_[741]_  = \new_[9961]_  & \new_[9950]_ ;
  assign \new_[742]_  = \new_[9941]_  & \new_[9930]_ ;
  assign \new_[743]_  = \new_[9921]_  & \new_[9910]_ ;
  assign \new_[744]_  = \new_[9901]_  & \new_[9890]_ ;
  assign \new_[745]_  = \new_[9881]_  & \new_[9870]_ ;
  assign \new_[746]_  = \new_[9861]_  & \new_[9850]_ ;
  assign \new_[747]_  = \new_[9841]_  & \new_[9830]_ ;
  assign \new_[748]_  = \new_[9821]_  & \new_[9810]_ ;
  assign \new_[749]_  = \new_[9801]_  & \new_[9790]_ ;
  assign \new_[750]_  = \new_[9781]_  & \new_[9770]_ ;
  assign \new_[751]_  = \new_[9761]_  & \new_[9750]_ ;
  assign \new_[752]_  = \new_[9741]_  & \new_[9730]_ ;
  assign \new_[753]_  = \new_[9721]_  & \new_[9710]_ ;
  assign \new_[754]_  = \new_[9701]_  & \new_[9690]_ ;
  assign \new_[755]_  = \new_[9681]_  & \new_[9670]_ ;
  assign \new_[756]_  = \new_[9661]_  & \new_[9650]_ ;
  assign \new_[757]_  = \new_[9641]_  & \new_[9630]_ ;
  assign \new_[758]_  = \new_[9621]_  & \new_[9610]_ ;
  assign \new_[759]_  = \new_[9601]_  & \new_[9590]_ ;
  assign \new_[760]_  = \new_[9581]_  & \new_[9570]_ ;
  assign \new_[761]_  = \new_[9561]_  & \new_[9550]_ ;
  assign \new_[762]_  = \new_[9541]_  & \new_[9530]_ ;
  assign \new_[763]_  = \new_[9521]_  & \new_[9510]_ ;
  assign \new_[764]_  = \new_[9501]_  & \new_[9490]_ ;
  assign \new_[765]_  = \new_[9481]_  & \new_[9470]_ ;
  assign \new_[766]_  = \new_[9461]_  & \new_[9450]_ ;
  assign \new_[767]_  = \new_[9441]_  & \new_[9430]_ ;
  assign \new_[768]_  = \new_[9421]_  & \new_[9410]_ ;
  assign \new_[769]_  = \new_[9401]_  & \new_[9390]_ ;
  assign \new_[770]_  = \new_[9381]_  & \new_[9370]_ ;
  assign \new_[771]_  = \new_[9361]_  & \new_[9350]_ ;
  assign \new_[772]_  = \new_[9341]_  & \new_[9330]_ ;
  assign \new_[773]_  = \new_[9321]_  & \new_[9310]_ ;
  assign \new_[774]_  = \new_[9301]_  & \new_[9290]_ ;
  assign \new_[775]_  = \new_[9281]_  & \new_[9270]_ ;
  assign \new_[776]_  = \new_[9261]_  & \new_[9250]_ ;
  assign \new_[777]_  = \new_[9241]_  & \new_[9230]_ ;
  assign \new_[778]_  = \new_[9221]_  & \new_[9210]_ ;
  assign \new_[779]_  = \new_[9201]_  & \new_[9190]_ ;
  assign \new_[780]_  = \new_[9181]_  & \new_[9170]_ ;
  assign \new_[781]_  = \new_[9161]_  & \new_[9150]_ ;
  assign \new_[782]_  = \new_[9141]_  & \new_[9130]_ ;
  assign \new_[783]_  = \new_[9121]_  & \new_[9110]_ ;
  assign \new_[784]_  = \new_[9101]_  & \new_[9090]_ ;
  assign \new_[785]_  = \new_[9081]_  & \new_[9070]_ ;
  assign \new_[786]_  = \new_[9061]_  & \new_[9050]_ ;
  assign \new_[787]_  = \new_[9041]_  & \new_[9030]_ ;
  assign \new_[788]_  = \new_[9021]_  & \new_[9010]_ ;
  assign \new_[789]_  = \new_[9001]_  & \new_[8990]_ ;
  assign \new_[790]_  = \new_[8981]_  & \new_[8970]_ ;
  assign \new_[791]_  = \new_[8961]_  & \new_[8950]_ ;
  assign \new_[792]_  = \new_[8941]_  & \new_[8930]_ ;
  assign \new_[793]_  = \new_[8921]_  & \new_[8910]_ ;
  assign \new_[794]_  = \new_[8901]_  & \new_[8890]_ ;
  assign \new_[795]_  = \new_[8881]_  & \new_[8870]_ ;
  assign \new_[796]_  = \new_[8861]_  & \new_[8850]_ ;
  assign \new_[797]_  = \new_[8841]_  & \new_[8830]_ ;
  assign \new_[798]_  = \new_[8821]_  & \new_[8810]_ ;
  assign \new_[799]_  = \new_[8801]_  & \new_[8790]_ ;
  assign \new_[800]_  = \new_[8781]_  & \new_[8770]_ ;
  assign \new_[801]_  = \new_[8761]_  & \new_[8750]_ ;
  assign \new_[802]_  = \new_[8741]_  & \new_[8730]_ ;
  assign \new_[803]_  = \new_[8721]_  & \new_[8710]_ ;
  assign \new_[804]_  = \new_[8701]_  & \new_[8690]_ ;
  assign \new_[805]_  = \new_[8681]_  & \new_[8670]_ ;
  assign \new_[806]_  = \new_[8661]_  & \new_[8650]_ ;
  assign \new_[807]_  = \new_[8641]_  & \new_[8630]_ ;
  assign \new_[808]_  = \new_[8621]_  & \new_[8610]_ ;
  assign \new_[809]_  = \new_[8601]_  & \new_[8590]_ ;
  assign \new_[810]_  = \new_[8581]_  & \new_[8570]_ ;
  assign \new_[811]_  = \new_[8561]_  & \new_[8550]_ ;
  assign \new_[812]_  = \new_[8541]_  & \new_[8530]_ ;
  assign \new_[813]_  = \new_[8521]_  & \new_[8510]_ ;
  assign \new_[814]_  = \new_[8501]_  & \new_[8490]_ ;
  assign \new_[815]_  = \new_[8481]_  & \new_[8470]_ ;
  assign \new_[816]_  = \new_[8461]_  & \new_[8450]_ ;
  assign \new_[817]_  = \new_[8441]_  & \new_[8430]_ ;
  assign \new_[818]_  = \new_[8421]_  & \new_[8410]_ ;
  assign \new_[819]_  = \new_[8401]_  & \new_[8390]_ ;
  assign \new_[820]_  = \new_[8381]_  & \new_[8370]_ ;
  assign \new_[821]_  = \new_[8361]_  & \new_[8350]_ ;
  assign \new_[822]_  = \new_[8341]_  & \new_[8330]_ ;
  assign \new_[823]_  = \new_[8321]_  & \new_[8310]_ ;
  assign \new_[824]_  = \new_[8301]_  & \new_[8290]_ ;
  assign \new_[825]_  = \new_[8281]_  & \new_[8270]_ ;
  assign \new_[826]_  = \new_[8261]_  & \new_[8250]_ ;
  assign \new_[827]_  = \new_[8241]_  & \new_[8230]_ ;
  assign \new_[828]_  = \new_[8221]_  & \new_[8210]_ ;
  assign \new_[829]_  = \new_[8201]_  & \new_[8190]_ ;
  assign \new_[830]_  = \new_[8181]_  & \new_[8170]_ ;
  assign \new_[831]_  = \new_[8161]_  & \new_[8150]_ ;
  assign \new_[832]_  = \new_[8141]_  & \new_[8130]_ ;
  assign \new_[833]_  = \new_[8121]_  & \new_[8112]_ ;
  assign \new_[834]_  = \new_[8103]_  & \new_[8094]_ ;
  assign \new_[835]_  = \new_[8085]_  & \new_[8076]_ ;
  assign \new_[836]_  = \new_[8067]_  & \new_[8058]_ ;
  assign \new_[837]_  = \new_[8049]_  & \new_[8040]_ ;
  assign \new_[838]_  = \new_[8031]_  & \new_[8022]_ ;
  assign \new_[839]_  = \new_[8013]_  & \new_[8004]_ ;
  assign \new_[840]_  = \new_[7995]_  & \new_[7986]_ ;
  assign \new_[841]_  = \new_[7977]_  & \new_[7968]_ ;
  assign \new_[842]_  = \new_[7959]_  & \new_[7950]_ ;
  assign \new_[843]_  = \new_[7941]_  & \new_[7932]_ ;
  assign \new_[844]_  = \new_[7923]_  & \new_[7914]_ ;
  assign \new_[845]_  = \new_[7905]_  & \new_[7896]_ ;
  assign \new_[846]_  = \new_[7887]_  & \new_[7878]_ ;
  assign \new_[847]_  = \new_[7869]_  & \new_[7860]_ ;
  assign \new_[848]_  = \new_[7851]_  & \new_[7842]_ ;
  assign \new_[849]_  = \new_[7833]_  & \new_[7824]_ ;
  assign \new_[850]_  = \new_[7815]_  & \new_[7806]_ ;
  assign \new_[851]_  = \new_[7797]_  & \new_[7788]_ ;
  assign \new_[852]_  = \new_[7779]_  & \new_[7770]_ ;
  assign \new_[853]_  = \new_[7761]_  & \new_[7752]_ ;
  assign \new_[854]_  = \new_[7743]_  & \new_[7734]_ ;
  assign \new_[855]_  = \new_[7725]_  & \new_[7716]_ ;
  assign \new_[856]_  = \new_[7707]_  & \new_[7698]_ ;
  assign \new_[857]_  = \new_[7689]_  & \new_[7680]_ ;
  assign \new_[858]_  = \new_[7671]_  & \new_[7662]_ ;
  assign \new_[859]_  = \new_[7653]_  & \new_[7644]_ ;
  assign \new_[860]_  = \new_[7635]_  & \new_[7626]_ ;
  assign \new_[861]_  = \new_[7617]_  & \new_[7608]_ ;
  assign \new_[862]_  = \new_[7599]_  & \new_[7590]_ ;
  assign \new_[863]_  = \new_[7581]_  & \new_[7572]_ ;
  assign \new_[864]_  = \new_[7563]_  & \new_[7554]_ ;
  assign \new_[865]_  = \new_[7545]_  & \new_[7536]_ ;
  assign \new_[866]_  = \new_[7527]_  & \new_[7518]_ ;
  assign \new_[867]_  = \new_[7509]_  & \new_[7500]_ ;
  assign \new_[868]_  = \new_[7491]_  & \new_[7482]_ ;
  assign \new_[869]_  = \new_[7473]_  & \new_[7464]_ ;
  assign \new_[870]_  = \new_[7455]_  & \new_[7446]_ ;
  assign \new_[871]_  = \new_[7437]_  & \new_[7428]_ ;
  assign \new_[872]_  = \new_[7419]_  & \new_[7410]_ ;
  assign \new_[873]_  = \new_[7401]_  & \new_[7392]_ ;
  assign \new_[874]_  = \new_[7383]_  & \new_[7374]_ ;
  assign \new_[875]_  = \new_[7365]_  & \new_[7356]_ ;
  assign \new_[876]_  = \new_[7347]_  & \new_[7338]_ ;
  assign \new_[877]_  = \new_[7329]_  & \new_[7320]_ ;
  assign \new_[878]_  = \new_[7311]_  & \new_[7302]_ ;
  assign \new_[879]_  = \new_[7293]_  & \new_[7284]_ ;
  assign \new_[880]_  = \new_[7275]_  & \new_[7266]_ ;
  assign \new_[881]_  = \new_[7257]_  & \new_[7248]_ ;
  assign \new_[882]_  = \new_[7239]_  & \new_[7230]_ ;
  assign \new_[883]_  = \new_[7221]_  & \new_[7212]_ ;
  assign \new_[884]_  = \new_[7203]_  & \new_[7194]_ ;
  assign \new_[885]_  = \new_[7185]_  & \new_[7176]_ ;
  assign \new_[886]_  = \new_[7167]_  & \new_[7158]_ ;
  assign \new_[887]_  = \new_[7149]_  & \new_[7140]_ ;
  assign \new_[888]_  = \new_[7131]_  & \new_[7122]_ ;
  assign \new_[889]_  = \new_[7113]_  & \new_[7104]_ ;
  assign \new_[890]_  = \new_[7095]_  & \new_[7086]_ ;
  assign \new_[891]_  = \new_[7077]_  & \new_[7068]_ ;
  assign \new_[892]_  = \new_[7059]_  & \new_[7050]_ ;
  assign \new_[893]_  = \new_[7041]_  & \new_[7032]_ ;
  assign \new_[894]_  = \new_[7023]_  & \new_[7014]_ ;
  assign \new_[895]_  = \new_[7005]_  & \new_[6996]_ ;
  assign \new_[896]_  = \new_[6987]_  & \new_[6978]_ ;
  assign \new_[897]_  = \new_[6969]_  & \new_[6960]_ ;
  assign \new_[898]_  = \new_[6951]_  & \new_[6942]_ ;
  assign \new_[899]_  = \new_[6933]_  & \new_[6924]_ ;
  assign \new_[900]_  = \new_[6915]_  & \new_[6906]_ ;
  assign \new_[901]_  = \new_[6897]_  & \new_[6888]_ ;
  assign \new_[902]_  = \new_[6879]_  & \new_[6870]_ ;
  assign \new_[903]_  = \new_[6861]_  & \new_[6852]_ ;
  assign \new_[904]_  = \new_[6843]_  & \new_[6834]_ ;
  assign \new_[905]_  = \new_[6825]_  & \new_[6816]_ ;
  assign \new_[906]_  = \new_[6807]_  & \new_[6798]_ ;
  assign \new_[907]_  = \new_[6789]_  & \new_[6780]_ ;
  assign \new_[908]_  = \new_[6771]_  & \new_[6762]_ ;
  assign \new_[909]_  = \new_[6753]_  & \new_[6744]_ ;
  assign \new_[910]_  = \new_[6735]_  & \new_[6726]_ ;
  assign \new_[911]_  = \new_[6717]_  & \new_[6708]_ ;
  assign \new_[912]_  = \new_[6699]_  & \new_[6690]_ ;
  assign \new_[913]_  = \new_[6681]_  & \new_[6672]_ ;
  assign \new_[914]_  = \new_[6663]_  & \new_[6654]_ ;
  assign \new_[915]_  = \new_[6645]_  & \new_[6636]_ ;
  assign \new_[916]_  = \new_[6627]_  & \new_[6618]_ ;
  assign \new_[917]_  = \new_[6609]_  & \new_[6600]_ ;
  assign \new_[918]_  = \new_[6591]_  & \new_[6582]_ ;
  assign \new_[919]_  = \new_[6573]_  & \new_[6564]_ ;
  assign \new_[920]_  = \new_[6555]_  & \new_[6546]_ ;
  assign \new_[921]_  = \new_[6537]_  & \new_[6528]_ ;
  assign \new_[922]_  = \new_[6519]_  & \new_[6510]_ ;
  assign \new_[923]_  = \new_[6501]_  & \new_[6492]_ ;
  assign \new_[924]_  = \new_[6483]_  & \new_[6474]_ ;
  assign \new_[925]_  = \new_[6465]_  & \new_[6456]_ ;
  assign \new_[926]_  = \new_[6447]_  & \new_[6438]_ ;
  assign \new_[927]_  = \new_[6429]_  & \new_[6420]_ ;
  assign \new_[928]_  = \new_[6411]_  & \new_[6402]_ ;
  assign \new_[929]_  = \new_[6393]_  & \new_[6384]_ ;
  assign \new_[930]_  = \new_[6375]_  & \new_[6366]_ ;
  assign \new_[931]_  = \new_[6357]_  & \new_[6348]_ ;
  assign \new_[932]_  = \new_[6339]_  & \new_[6330]_ ;
  assign \new_[933]_  = \new_[6321]_  & \new_[6312]_ ;
  assign \new_[934]_  = \new_[6303]_  & \new_[6294]_ ;
  assign \new_[935]_  = \new_[6285]_  & \new_[6276]_ ;
  assign \new_[936]_  = \new_[6267]_  & \new_[6258]_ ;
  assign \new_[937]_  = \new_[6249]_  & \new_[6240]_ ;
  assign \new_[938]_  = \new_[6231]_  & \new_[6222]_ ;
  assign \new_[939]_  = \new_[6213]_  & \new_[6204]_ ;
  assign \new_[940]_  = \new_[6195]_  & \new_[6186]_ ;
  assign \new_[941]_  = \new_[6177]_  & \new_[6168]_ ;
  assign \new_[942]_  = \new_[6159]_  & \new_[6150]_ ;
  assign \new_[943]_  = \new_[6141]_  & \new_[6132]_ ;
  assign \new_[944]_  = \new_[6123]_  & \new_[6114]_ ;
  assign \new_[945]_  = \new_[6105]_  & \new_[6096]_ ;
  assign \new_[946]_  = \new_[6087]_  & \new_[6078]_ ;
  assign \new_[947]_  = \new_[6069]_  & \new_[6060]_ ;
  assign \new_[948]_  = \new_[6051]_  & \new_[6042]_ ;
  assign \new_[949]_  = \new_[6033]_  & \new_[6024]_ ;
  assign \new_[950]_  = \new_[6015]_  & \new_[6006]_ ;
  assign \new_[951]_  = \new_[5997]_  & \new_[5988]_ ;
  assign \new_[952]_  = \new_[5979]_  & \new_[5970]_ ;
  assign \new_[953]_  = \new_[5961]_  & \new_[5952]_ ;
  assign \new_[954]_  = \new_[5943]_  & \new_[5934]_ ;
  assign \new_[955]_  = \new_[5925]_  & \new_[5916]_ ;
  assign \new_[956]_  = \new_[5907]_  & \new_[5898]_ ;
  assign \new_[957]_  = \new_[5889]_  & \new_[5880]_ ;
  assign \new_[958]_  = \new_[5871]_  & \new_[5862]_ ;
  assign \new_[959]_  = \new_[5853]_  & \new_[5844]_ ;
  assign \new_[960]_  = \new_[5835]_  & \new_[5826]_ ;
  assign \new_[961]_  = \new_[5817]_  & \new_[5808]_ ;
  assign \new_[962]_  = \new_[5799]_  & \new_[5790]_ ;
  assign \new_[963]_  = \new_[5781]_  & \new_[5772]_ ;
  assign \new_[964]_  = \new_[5763]_  & \new_[5754]_ ;
  assign \new_[965]_  = \new_[5745]_  & \new_[5736]_ ;
  assign \new_[966]_  = \new_[5727]_  & \new_[5718]_ ;
  assign \new_[967]_  = \new_[5709]_  & \new_[5700]_ ;
  assign \new_[968]_  = \new_[5691]_  & \new_[5682]_ ;
  assign \new_[969]_  = \new_[5673]_  & \new_[5664]_ ;
  assign \new_[970]_  = \new_[5655]_  & \new_[5646]_ ;
  assign \new_[971]_  = \new_[5637]_  & \new_[5628]_ ;
  assign \new_[972]_  = \new_[5619]_  & \new_[5610]_ ;
  assign \new_[973]_  = \new_[5601]_  & \new_[5592]_ ;
  assign \new_[974]_  = \new_[5583]_  & \new_[5574]_ ;
  assign \new_[975]_  = \new_[5565]_  & \new_[5556]_ ;
  assign \new_[976]_  = \new_[5547]_  & \new_[5538]_ ;
  assign \new_[977]_  = \new_[5529]_  & \new_[5520]_ ;
  assign \new_[978]_  = \new_[5511]_  & \new_[5502]_ ;
  assign \new_[979]_  = \new_[5493]_  & \new_[5484]_ ;
  assign \new_[980]_  = \new_[5475]_  & \new_[5466]_ ;
  assign \new_[981]_  = \new_[5457]_  & \new_[5448]_ ;
  assign \new_[982]_  = \new_[5439]_  & \new_[5430]_ ;
  assign \new_[983]_  = \new_[5421]_  & \new_[5412]_ ;
  assign \new_[984]_  = \new_[5403]_  & \new_[5394]_ ;
  assign \new_[985]_  = \new_[5385]_  & \new_[5376]_ ;
  assign \new_[986]_  = \new_[5367]_  & \new_[5358]_ ;
  assign \new_[987]_  = \new_[5349]_  & \new_[5340]_ ;
  assign \new_[988]_  = \new_[5331]_  & \new_[5322]_ ;
  assign \new_[989]_  = \new_[5313]_  & \new_[5304]_ ;
  assign \new_[990]_  = \new_[5295]_  & \new_[5286]_ ;
  assign \new_[991]_  = \new_[5277]_  & \new_[5268]_ ;
  assign \new_[992]_  = \new_[5259]_  & \new_[5250]_ ;
  assign \new_[993]_  = \new_[5241]_  & \new_[5232]_ ;
  assign \new_[994]_  = \new_[5223]_  & \new_[5214]_ ;
  assign \new_[995]_  = \new_[5205]_  & \new_[5196]_ ;
  assign \new_[996]_  = \new_[5187]_  & \new_[5178]_ ;
  assign \new_[997]_  = \new_[5169]_  & \new_[5160]_ ;
  assign \new_[998]_  = \new_[5151]_  & \new_[5142]_ ;
  assign \new_[999]_  = \new_[5133]_  & \new_[5124]_ ;
  assign \new_[1000]_  = \new_[5115]_  & \new_[5106]_ ;
  assign \new_[1001]_  = \new_[5097]_  & \new_[5088]_ ;
  assign \new_[1002]_  = \new_[5079]_  & \new_[5070]_ ;
  assign \new_[1003]_  = \new_[5061]_  & \new_[5052]_ ;
  assign \new_[1004]_  = \new_[5043]_  & \new_[5034]_ ;
  assign \new_[1005]_  = \new_[5025]_  & \new_[5016]_ ;
  assign \new_[1006]_  = \new_[5007]_  & \new_[4998]_ ;
  assign \new_[1007]_  = \new_[4989]_  & \new_[4980]_ ;
  assign \new_[1008]_  = \new_[4973]_  & \new_[4964]_ ;
  assign \new_[1009]_  = \new_[4957]_  & \new_[4948]_ ;
  assign \new_[1010]_  = \new_[4941]_  & \new_[4932]_ ;
  assign \new_[1011]_  = \new_[4925]_  & \new_[4916]_ ;
  assign \new_[1012]_  = \new_[4909]_  & \new_[4900]_ ;
  assign \new_[1013]_  = \new_[4893]_  & \new_[4884]_ ;
  assign \new_[1014]_  = \new_[4877]_  & \new_[4868]_ ;
  assign \new_[1015]_  = \new_[4861]_  & \new_[4852]_ ;
  assign \new_[1016]_  = \new_[4845]_  & \new_[4836]_ ;
  assign \new_[1017]_  = \new_[4829]_  & \new_[4820]_ ;
  assign \new_[1018]_  = \new_[4813]_  & \new_[4804]_ ;
  assign \new_[1019]_  = \new_[4797]_  & \new_[4788]_ ;
  assign \new_[1020]_  = \new_[4781]_  & \new_[4772]_ ;
  assign \new_[1021]_  = \new_[4765]_  & \new_[4756]_ ;
  assign \new_[1022]_  = \new_[4749]_  & \new_[4740]_ ;
  assign \new_[1023]_  = \new_[4733]_  & \new_[4724]_ ;
  assign \new_[1024]_  = \new_[4717]_  & \new_[4708]_ ;
  assign \new_[1025]_  = \new_[4701]_  & \new_[4692]_ ;
  assign \new_[1026]_  = \new_[4685]_  & \new_[4676]_ ;
  assign \new_[1027]_  = \new_[4669]_  & \new_[4660]_ ;
  assign \new_[1028]_  = \new_[4653]_  & \new_[4644]_ ;
  assign \new_[1029]_  = \new_[4637]_  & \new_[4628]_ ;
  assign \new_[1030]_  = \new_[4621]_  & \new_[4612]_ ;
  assign \new_[1031]_  = \new_[4605]_  & \new_[4596]_ ;
  assign \new_[1032]_  = \new_[4589]_  & \new_[4580]_ ;
  assign \new_[1033]_  = \new_[4573]_  & \new_[4564]_ ;
  assign \new_[1034]_  = \new_[4557]_  & \new_[4548]_ ;
  assign \new_[1035]_  = \new_[4541]_  & \new_[4532]_ ;
  assign \new_[1036]_  = \new_[4525]_  & \new_[4516]_ ;
  assign \new_[1037]_  = \new_[4509]_  & \new_[4500]_ ;
  assign \new_[1038]_  = \new_[4493]_  & \new_[4484]_ ;
  assign \new_[1039]_  = \new_[4477]_  & \new_[4468]_ ;
  assign \new_[1040]_  = \new_[4461]_  & \new_[4452]_ ;
  assign \new_[1041]_  = \new_[4445]_  & \new_[4436]_ ;
  assign \new_[1042]_  = \new_[4429]_  & \new_[4420]_ ;
  assign \new_[1043]_  = \new_[4413]_  & \new_[4404]_ ;
  assign \new_[1044]_  = \new_[4397]_  & \new_[4388]_ ;
  assign \new_[1045]_  = \new_[4381]_  & \new_[4372]_ ;
  assign \new_[1046]_  = \new_[4365]_  & \new_[4356]_ ;
  assign \new_[1047]_  = \new_[4349]_  & \new_[4340]_ ;
  assign \new_[1048]_  = \new_[4333]_  & \new_[4324]_ ;
  assign \new_[1049]_  = \new_[4317]_  & \new_[4308]_ ;
  assign \new_[1050]_  = \new_[4301]_  & \new_[4292]_ ;
  assign \new_[1051]_  = \new_[4285]_  & \new_[4276]_ ;
  assign \new_[1052]_  = \new_[4269]_  & \new_[4260]_ ;
  assign \new_[1053]_  = \new_[4253]_  & \new_[4244]_ ;
  assign \new_[1054]_  = \new_[4237]_  & \new_[4228]_ ;
  assign \new_[1055]_  = \new_[4221]_  & \new_[4212]_ ;
  assign \new_[1056]_  = \new_[4205]_  & \new_[4196]_ ;
  assign \new_[1057]_  = \new_[4189]_  & \new_[4180]_ ;
  assign \new_[1058]_  = \new_[4173]_  & \new_[4164]_ ;
  assign \new_[1059]_  = \new_[4157]_  & \new_[4148]_ ;
  assign \new_[1060]_  = \new_[4141]_  & \new_[4132]_ ;
  assign \new_[1061]_  = \new_[4125]_  & \new_[4116]_ ;
  assign \new_[1062]_  = \new_[4109]_  & \new_[4100]_ ;
  assign \new_[1063]_  = \new_[4093]_  & \new_[4084]_ ;
  assign \new_[1064]_  = \new_[4077]_  & \new_[4068]_ ;
  assign \new_[1065]_  = \new_[4061]_  & \new_[4052]_ ;
  assign \new_[1066]_  = \new_[4045]_  & \new_[4036]_ ;
  assign \new_[1067]_  = \new_[4029]_  & \new_[4020]_ ;
  assign \new_[1068]_  = \new_[4013]_  & \new_[4004]_ ;
  assign \new_[1069]_  = \new_[3997]_  & \new_[3990]_ ;
  assign \new_[1070]_  = \new_[3983]_  & \new_[3976]_ ;
  assign \new_[1071]_  = \new_[3969]_  & \new_[3962]_ ;
  assign \new_[1072]_  = \new_[3955]_  & \new_[3948]_ ;
  assign \new_[1073]_  = \new_[3941]_  & \new_[3934]_ ;
  assign \new_[1074]_  = \new_[3927]_  & \new_[3920]_ ;
  assign \new_[1075]_  = \new_[3913]_  & \new_[3906]_ ;
  assign \new_[1076]_  = \new_[3899]_  & \new_[3892]_ ;
  assign \new_[1077]_  = \new_[3885]_  & \new_[3878]_ ;
  assign \new_[1078]_  = \new_[3871]_  & \new_[3864]_ ;
  assign \new_[1079]_  = \new_[3857]_  & \new_[3850]_ ;
  assign \new_[1080]_  = \new_[3843]_  & \new_[3836]_ ;
  assign \new_[1081]_  = \new_[3829]_  & \new_[3822]_ ;
  assign \new_[1082]_  = \new_[3815]_  & \new_[3808]_ ;
  assign \new_[1083]_  = \new_[3801]_  & \new_[3794]_ ;
  assign \new_[1084]_  = \new_[3787]_  & \new_[3780]_ ;
  assign \new_[1085]_  = \new_[3773]_  & \new_[3766]_ ;
  assign \new_[1086]_  = \new_[3759]_  & \new_[3752]_ ;
  assign \new_[1087]_  = \new_[3745]_  & \new_[3738]_ ;
  assign \new_[1088]_  = \new_[3731]_  & \new_[3724]_ ;
  assign \new_[1089]_  = \new_[3717]_  & \new_[3710]_ ;
  assign \new_[1090]_  = \new_[3703]_  & \new_[3696]_ ;
  assign \new_[1091]_  = \new_[3689]_  & \new_[3682]_ ;
  assign \new_[1092]_  = \new_[3675]_  & \new_[3668]_ ;
  assign \new_[1093]_  = \new_[3661]_  & \new_[3654]_ ;
  assign \new_[1094]_  = \new_[3647]_  & \new_[3640]_ ;
  assign \new_[1095]_  = \new_[3633]_  & \new_[3626]_ ;
  assign \new_[1096]_  = \new_[3619]_  & \new_[3612]_ ;
  assign \new_[1097]_  = \new_[3605]_  & \new_[3598]_ ;
  assign \new_[1098]_  = \new_[3591]_  & \new_[3584]_ ;
  assign \new_[1099]_  = \new_[3577]_  & \new_[3570]_ ;
  assign \new_[1100]_  = \new_[3563]_  & \new_[3556]_ ;
  assign \new_[1101]_  = \new_[3549]_  & \new_[3542]_ ;
  assign \new_[1102]_  = \new_[3535]_  & \new_[3528]_ ;
  assign \new_[1103]_  = \new_[3521]_  & \new_[3514]_ ;
  assign \new_[1104]_  = \new_[3507]_  & \new_[3500]_ ;
  assign \new_[1105]_  = \new_[3493]_  & \new_[3488]_ ;
  assign \new_[1106]_  = \new_[3483]_  & \new_[3478]_ ;
  assign \new_[1107]_  = \new_[3473]_  & \new_[3468]_ ;
  assign \new_[1108]_  = \new_[3463]_  & \new_[3458]_ ;
  assign \new_[1109]_  = \new_[3453]_  & \new_[3448]_ ;
  assign \new_[1110]_  = \new_[3443]_  & \new_[3438]_ ;
  assign \new_[1111]_  = \new_[3433]_  & \new_[3428]_ ;
  assign \new_[1112]_  = \new_[3423]_  & \new_[3418]_ ;
  assign \new_[1113]_  = \new_[3413]_  & \new_[3408]_ ;
  assign \new_[1114]_  = \new_[3403]_  & \new_[3398]_ ;
  assign \new_[1115]_  = \new_[3393]_  & \new_[3388]_ ;
  assign \new_[1116]_  = \new_[3383]_  & \new_[3378]_ ;
  assign \new_[1117]_  = \new_[3373]_  & \new_[3370]_ ;
  assign \new_[1118]_  = \new_[3367]_  & \new_[3364]_ ;
  assign \new_[1119]_  = \new_[3361]_  & \new_[3358]_ ;
  assign \new_[1122]_  = \new_[1118]_  | \new_[1119]_ ;
  assign \new_[1125]_  = \new_[1116]_  | \new_[1117]_ ;
  assign \new_[1126]_  = \new_[1125]_  | \new_[1122]_ ;
  assign \new_[1129]_  = \new_[1114]_  | \new_[1115]_ ;
  assign \new_[1132]_  = \new_[1112]_  | \new_[1113]_ ;
  assign \new_[1133]_  = \new_[1132]_  | \new_[1129]_ ;
  assign \new_[1134]_  = \new_[1133]_  | \new_[1126]_ ;
  assign \new_[1137]_  = \new_[1110]_  | \new_[1111]_ ;
  assign \new_[1140]_  = \new_[1108]_  | \new_[1109]_ ;
  assign \new_[1141]_  = \new_[1140]_  | \new_[1137]_ ;
  assign \new_[1144]_  = \new_[1106]_  | \new_[1107]_ ;
  assign \new_[1148]_  = \new_[1103]_  | \new_[1104]_ ;
  assign \new_[1149]_  = \new_[1105]_  | \new_[1148]_ ;
  assign \new_[1150]_  = \new_[1149]_  | \new_[1144]_ ;
  assign \new_[1151]_  = \new_[1150]_  | \new_[1141]_ ;
  assign \new_[1152]_  = \new_[1151]_  | \new_[1134]_ ;
  assign \new_[1155]_  = \new_[1101]_  | \new_[1102]_ ;
  assign \new_[1158]_  = \new_[1099]_  | \new_[1100]_ ;
  assign \new_[1159]_  = \new_[1158]_  | \new_[1155]_ ;
  assign \new_[1162]_  = \new_[1097]_  | \new_[1098]_ ;
  assign \new_[1165]_  = \new_[1095]_  | \new_[1096]_ ;
  assign \new_[1166]_  = \new_[1165]_  | \new_[1162]_ ;
  assign \new_[1167]_  = \new_[1166]_  | \new_[1159]_ ;
  assign \new_[1170]_  = \new_[1093]_  | \new_[1094]_ ;
  assign \new_[1173]_  = \new_[1091]_  | \new_[1092]_ ;
  assign \new_[1174]_  = \new_[1173]_  | \new_[1170]_ ;
  assign \new_[1177]_  = \new_[1089]_  | \new_[1090]_ ;
  assign \new_[1181]_  = \new_[1086]_  | \new_[1087]_ ;
  assign \new_[1182]_  = \new_[1088]_  | \new_[1181]_ ;
  assign \new_[1183]_  = \new_[1182]_  | \new_[1177]_ ;
  assign \new_[1184]_  = \new_[1183]_  | \new_[1174]_ ;
  assign \new_[1185]_  = \new_[1184]_  | \new_[1167]_ ;
  assign \new_[1186]_  = \new_[1185]_  | \new_[1152]_ ;
  assign \new_[1189]_  = \new_[1084]_  | \new_[1085]_ ;
  assign \new_[1192]_  = \new_[1082]_  | \new_[1083]_ ;
  assign \new_[1193]_  = \new_[1192]_  | \new_[1189]_ ;
  assign \new_[1196]_  = \new_[1080]_  | \new_[1081]_ ;
  assign \new_[1199]_  = \new_[1078]_  | \new_[1079]_ ;
  assign \new_[1200]_  = \new_[1199]_  | \new_[1196]_ ;
  assign \new_[1201]_  = \new_[1200]_  | \new_[1193]_ ;
  assign \new_[1204]_  = \new_[1076]_  | \new_[1077]_ ;
  assign \new_[1207]_  = \new_[1074]_  | \new_[1075]_ ;
  assign \new_[1208]_  = \new_[1207]_  | \new_[1204]_ ;
  assign \new_[1211]_  = \new_[1072]_  | \new_[1073]_ ;
  assign \new_[1215]_  = \new_[1069]_  | \new_[1070]_ ;
  assign \new_[1216]_  = \new_[1071]_  | \new_[1215]_ ;
  assign \new_[1217]_  = \new_[1216]_  | \new_[1211]_ ;
  assign \new_[1218]_  = \new_[1217]_  | \new_[1208]_ ;
  assign \new_[1219]_  = \new_[1218]_  | \new_[1201]_ ;
  assign \new_[1222]_  = \new_[1067]_  | \new_[1068]_ ;
  assign \new_[1225]_  = \new_[1065]_  | \new_[1066]_ ;
  assign \new_[1226]_  = \new_[1225]_  | \new_[1222]_ ;
  assign \new_[1229]_  = \new_[1063]_  | \new_[1064]_ ;
  assign \new_[1233]_  = \new_[1060]_  | \new_[1061]_ ;
  assign \new_[1234]_  = \new_[1062]_  | \new_[1233]_ ;
  assign \new_[1235]_  = \new_[1234]_  | \new_[1229]_ ;
  assign \new_[1236]_  = \new_[1235]_  | \new_[1226]_ ;
  assign \new_[1239]_  = \new_[1058]_  | \new_[1059]_ ;
  assign \new_[1242]_  = \new_[1056]_  | \new_[1057]_ ;
  assign \new_[1243]_  = \new_[1242]_  | \new_[1239]_ ;
  assign \new_[1246]_  = \new_[1054]_  | \new_[1055]_ ;
  assign \new_[1250]_  = \new_[1051]_  | \new_[1052]_ ;
  assign \new_[1251]_  = \new_[1053]_  | \new_[1250]_ ;
  assign \new_[1252]_  = \new_[1251]_  | \new_[1246]_ ;
  assign \new_[1253]_  = \new_[1252]_  | \new_[1243]_ ;
  assign \new_[1254]_  = \new_[1253]_  | \new_[1236]_ ;
  assign \new_[1255]_  = \new_[1254]_  | \new_[1219]_ ;
  assign \new_[1256]_  = \new_[1255]_  | \new_[1186]_ ;
  assign \new_[1259]_  = \new_[1049]_  | \new_[1050]_ ;
  assign \new_[1262]_  = \new_[1047]_  | \new_[1048]_ ;
  assign \new_[1263]_  = \new_[1262]_  | \new_[1259]_ ;
  assign \new_[1266]_  = \new_[1045]_  | \new_[1046]_ ;
  assign \new_[1269]_  = \new_[1043]_  | \new_[1044]_ ;
  assign \new_[1270]_  = \new_[1269]_  | \new_[1266]_ ;
  assign \new_[1271]_  = \new_[1270]_  | \new_[1263]_ ;
  assign \new_[1274]_  = \new_[1041]_  | \new_[1042]_ ;
  assign \new_[1277]_  = \new_[1039]_  | \new_[1040]_ ;
  assign \new_[1278]_  = \new_[1277]_  | \new_[1274]_ ;
  assign \new_[1281]_  = \new_[1037]_  | \new_[1038]_ ;
  assign \new_[1285]_  = \new_[1034]_  | \new_[1035]_ ;
  assign \new_[1286]_  = \new_[1036]_  | \new_[1285]_ ;
  assign \new_[1287]_  = \new_[1286]_  | \new_[1281]_ ;
  assign \new_[1288]_  = \new_[1287]_  | \new_[1278]_ ;
  assign \new_[1289]_  = \new_[1288]_  | \new_[1271]_ ;
  assign \new_[1292]_  = \new_[1032]_  | \new_[1033]_ ;
  assign \new_[1295]_  = \new_[1030]_  | \new_[1031]_ ;
  assign \new_[1296]_  = \new_[1295]_  | \new_[1292]_ ;
  assign \new_[1299]_  = \new_[1028]_  | \new_[1029]_ ;
  assign \new_[1303]_  = \new_[1025]_  | \new_[1026]_ ;
  assign \new_[1304]_  = \new_[1027]_  | \new_[1303]_ ;
  assign \new_[1305]_  = \new_[1304]_  | \new_[1299]_ ;
  assign \new_[1306]_  = \new_[1305]_  | \new_[1296]_ ;
  assign \new_[1309]_  = \new_[1023]_  | \new_[1024]_ ;
  assign \new_[1312]_  = \new_[1021]_  | \new_[1022]_ ;
  assign \new_[1313]_  = \new_[1312]_  | \new_[1309]_ ;
  assign \new_[1316]_  = \new_[1019]_  | \new_[1020]_ ;
  assign \new_[1320]_  = \new_[1016]_  | \new_[1017]_ ;
  assign \new_[1321]_  = \new_[1018]_  | \new_[1320]_ ;
  assign \new_[1322]_  = \new_[1321]_  | \new_[1316]_ ;
  assign \new_[1323]_  = \new_[1322]_  | \new_[1313]_ ;
  assign \new_[1324]_  = \new_[1323]_  | \new_[1306]_ ;
  assign \new_[1325]_  = \new_[1324]_  | \new_[1289]_ ;
  assign \new_[1328]_  = \new_[1014]_  | \new_[1015]_ ;
  assign \new_[1331]_  = \new_[1012]_  | \new_[1013]_ ;
  assign \new_[1332]_  = \new_[1331]_  | \new_[1328]_ ;
  assign \new_[1335]_  = \new_[1010]_  | \new_[1011]_ ;
  assign \new_[1338]_  = \new_[1008]_  | \new_[1009]_ ;
  assign \new_[1339]_  = \new_[1338]_  | \new_[1335]_ ;
  assign \new_[1340]_  = \new_[1339]_  | \new_[1332]_ ;
  assign \new_[1343]_  = \new_[1006]_  | \new_[1007]_ ;
  assign \new_[1346]_  = \new_[1004]_  | \new_[1005]_ ;
  assign \new_[1347]_  = \new_[1346]_  | \new_[1343]_ ;
  assign \new_[1350]_  = \new_[1002]_  | \new_[1003]_ ;
  assign \new_[1354]_  = \new_[999]_  | \new_[1000]_ ;
  assign \new_[1355]_  = \new_[1001]_  | \new_[1354]_ ;
  assign \new_[1356]_  = \new_[1355]_  | \new_[1350]_ ;
  assign \new_[1357]_  = \new_[1356]_  | \new_[1347]_ ;
  assign \new_[1358]_  = \new_[1357]_  | \new_[1340]_ ;
  assign \new_[1361]_  = \new_[997]_  | \new_[998]_ ;
  assign \new_[1364]_  = \new_[995]_  | \new_[996]_ ;
  assign \new_[1365]_  = \new_[1364]_  | \new_[1361]_ ;
  assign \new_[1368]_  = \new_[993]_  | \new_[994]_ ;
  assign \new_[1372]_  = \new_[990]_  | \new_[991]_ ;
  assign \new_[1373]_  = \new_[992]_  | \new_[1372]_ ;
  assign \new_[1374]_  = \new_[1373]_  | \new_[1368]_ ;
  assign \new_[1375]_  = \new_[1374]_  | \new_[1365]_ ;
  assign \new_[1378]_  = \new_[988]_  | \new_[989]_ ;
  assign \new_[1381]_  = \new_[986]_  | \new_[987]_ ;
  assign \new_[1382]_  = \new_[1381]_  | \new_[1378]_ ;
  assign \new_[1385]_  = \new_[984]_  | \new_[985]_ ;
  assign \new_[1389]_  = \new_[981]_  | \new_[982]_ ;
  assign \new_[1390]_  = \new_[983]_  | \new_[1389]_ ;
  assign \new_[1391]_  = \new_[1390]_  | \new_[1385]_ ;
  assign \new_[1392]_  = \new_[1391]_  | \new_[1382]_ ;
  assign \new_[1393]_  = \new_[1392]_  | \new_[1375]_ ;
  assign \new_[1394]_  = \new_[1393]_  | \new_[1358]_ ;
  assign \new_[1395]_  = \new_[1394]_  | \new_[1325]_ ;
  assign \new_[1396]_  = \new_[1395]_  | \new_[1256]_ ;
  assign \new_[1399]_  = \new_[979]_  | \new_[980]_ ;
  assign \new_[1402]_  = \new_[977]_  | \new_[978]_ ;
  assign \new_[1403]_  = \new_[1402]_  | \new_[1399]_ ;
  assign \new_[1406]_  = \new_[975]_  | \new_[976]_ ;
  assign \new_[1409]_  = \new_[973]_  | \new_[974]_ ;
  assign \new_[1410]_  = \new_[1409]_  | \new_[1406]_ ;
  assign \new_[1411]_  = \new_[1410]_  | \new_[1403]_ ;
  assign \new_[1414]_  = \new_[971]_  | \new_[972]_ ;
  assign \new_[1417]_  = \new_[969]_  | \new_[970]_ ;
  assign \new_[1418]_  = \new_[1417]_  | \new_[1414]_ ;
  assign \new_[1421]_  = \new_[967]_  | \new_[968]_ ;
  assign \new_[1425]_  = \new_[964]_  | \new_[965]_ ;
  assign \new_[1426]_  = \new_[966]_  | \new_[1425]_ ;
  assign \new_[1427]_  = \new_[1426]_  | \new_[1421]_ ;
  assign \new_[1428]_  = \new_[1427]_  | \new_[1418]_ ;
  assign \new_[1429]_  = \new_[1428]_  | \new_[1411]_ ;
  assign \new_[1432]_  = \new_[962]_  | \new_[963]_ ;
  assign \new_[1435]_  = \new_[960]_  | \new_[961]_ ;
  assign \new_[1436]_  = \new_[1435]_  | \new_[1432]_ ;
  assign \new_[1439]_  = \new_[958]_  | \new_[959]_ ;
  assign \new_[1443]_  = \new_[955]_  | \new_[956]_ ;
  assign \new_[1444]_  = \new_[957]_  | \new_[1443]_ ;
  assign \new_[1445]_  = \new_[1444]_  | \new_[1439]_ ;
  assign \new_[1446]_  = \new_[1445]_  | \new_[1436]_ ;
  assign \new_[1449]_  = \new_[953]_  | \new_[954]_ ;
  assign \new_[1452]_  = \new_[951]_  | \new_[952]_ ;
  assign \new_[1453]_  = \new_[1452]_  | \new_[1449]_ ;
  assign \new_[1456]_  = \new_[949]_  | \new_[950]_ ;
  assign \new_[1460]_  = \new_[946]_  | \new_[947]_ ;
  assign \new_[1461]_  = \new_[948]_  | \new_[1460]_ ;
  assign \new_[1462]_  = \new_[1461]_  | \new_[1456]_ ;
  assign \new_[1463]_  = \new_[1462]_  | \new_[1453]_ ;
  assign \new_[1464]_  = \new_[1463]_  | \new_[1446]_ ;
  assign \new_[1465]_  = \new_[1464]_  | \new_[1429]_ ;
  assign \new_[1468]_  = \new_[944]_  | \new_[945]_ ;
  assign \new_[1471]_  = \new_[942]_  | \new_[943]_ ;
  assign \new_[1472]_  = \new_[1471]_  | \new_[1468]_ ;
  assign \new_[1475]_  = \new_[940]_  | \new_[941]_ ;
  assign \new_[1478]_  = \new_[938]_  | \new_[939]_ ;
  assign \new_[1479]_  = \new_[1478]_  | \new_[1475]_ ;
  assign \new_[1480]_  = \new_[1479]_  | \new_[1472]_ ;
  assign \new_[1483]_  = \new_[936]_  | \new_[937]_ ;
  assign \new_[1486]_  = \new_[934]_  | \new_[935]_ ;
  assign \new_[1487]_  = \new_[1486]_  | \new_[1483]_ ;
  assign \new_[1490]_  = \new_[932]_  | \new_[933]_ ;
  assign \new_[1494]_  = \new_[929]_  | \new_[930]_ ;
  assign \new_[1495]_  = \new_[931]_  | \new_[1494]_ ;
  assign \new_[1496]_  = \new_[1495]_  | \new_[1490]_ ;
  assign \new_[1497]_  = \new_[1496]_  | \new_[1487]_ ;
  assign \new_[1498]_  = \new_[1497]_  | \new_[1480]_ ;
  assign \new_[1501]_  = \new_[927]_  | \new_[928]_ ;
  assign \new_[1504]_  = \new_[925]_  | \new_[926]_ ;
  assign \new_[1505]_  = \new_[1504]_  | \new_[1501]_ ;
  assign \new_[1508]_  = \new_[923]_  | \new_[924]_ ;
  assign \new_[1512]_  = \new_[920]_  | \new_[921]_ ;
  assign \new_[1513]_  = \new_[922]_  | \new_[1512]_ ;
  assign \new_[1514]_  = \new_[1513]_  | \new_[1508]_ ;
  assign \new_[1515]_  = \new_[1514]_  | \new_[1505]_ ;
  assign \new_[1518]_  = \new_[918]_  | \new_[919]_ ;
  assign \new_[1521]_  = \new_[916]_  | \new_[917]_ ;
  assign \new_[1522]_  = \new_[1521]_  | \new_[1518]_ ;
  assign \new_[1525]_  = \new_[914]_  | \new_[915]_ ;
  assign \new_[1529]_  = \new_[911]_  | \new_[912]_ ;
  assign \new_[1530]_  = \new_[913]_  | \new_[1529]_ ;
  assign \new_[1531]_  = \new_[1530]_  | \new_[1525]_ ;
  assign \new_[1532]_  = \new_[1531]_  | \new_[1522]_ ;
  assign \new_[1533]_  = \new_[1532]_  | \new_[1515]_ ;
  assign \new_[1534]_  = \new_[1533]_  | \new_[1498]_ ;
  assign \new_[1535]_  = \new_[1534]_  | \new_[1465]_ ;
  assign \new_[1538]_  = \new_[909]_  | \new_[910]_ ;
  assign \new_[1541]_  = \new_[907]_  | \new_[908]_ ;
  assign \new_[1542]_  = \new_[1541]_  | \new_[1538]_ ;
  assign \new_[1545]_  = \new_[905]_  | \new_[906]_ ;
  assign \new_[1548]_  = \new_[903]_  | \new_[904]_ ;
  assign \new_[1549]_  = \new_[1548]_  | \new_[1545]_ ;
  assign \new_[1550]_  = \new_[1549]_  | \new_[1542]_ ;
  assign \new_[1553]_  = \new_[901]_  | \new_[902]_ ;
  assign \new_[1556]_  = \new_[899]_  | \new_[900]_ ;
  assign \new_[1557]_  = \new_[1556]_  | \new_[1553]_ ;
  assign \new_[1560]_  = \new_[897]_  | \new_[898]_ ;
  assign \new_[1564]_  = \new_[894]_  | \new_[895]_ ;
  assign \new_[1565]_  = \new_[896]_  | \new_[1564]_ ;
  assign \new_[1566]_  = \new_[1565]_  | \new_[1560]_ ;
  assign \new_[1567]_  = \new_[1566]_  | \new_[1557]_ ;
  assign \new_[1568]_  = \new_[1567]_  | \new_[1550]_ ;
  assign \new_[1571]_  = \new_[892]_  | \new_[893]_ ;
  assign \new_[1574]_  = \new_[890]_  | \new_[891]_ ;
  assign \new_[1575]_  = \new_[1574]_  | \new_[1571]_ ;
  assign \new_[1578]_  = \new_[888]_  | \new_[889]_ ;
  assign \new_[1582]_  = \new_[885]_  | \new_[886]_ ;
  assign \new_[1583]_  = \new_[887]_  | \new_[1582]_ ;
  assign \new_[1584]_  = \new_[1583]_  | \new_[1578]_ ;
  assign \new_[1585]_  = \new_[1584]_  | \new_[1575]_ ;
  assign \new_[1588]_  = \new_[883]_  | \new_[884]_ ;
  assign \new_[1591]_  = \new_[881]_  | \new_[882]_ ;
  assign \new_[1592]_  = \new_[1591]_  | \new_[1588]_ ;
  assign \new_[1595]_  = \new_[879]_  | \new_[880]_ ;
  assign \new_[1599]_  = \new_[876]_  | \new_[877]_ ;
  assign \new_[1600]_  = \new_[878]_  | \new_[1599]_ ;
  assign \new_[1601]_  = \new_[1600]_  | \new_[1595]_ ;
  assign \new_[1602]_  = \new_[1601]_  | \new_[1592]_ ;
  assign \new_[1603]_  = \new_[1602]_  | \new_[1585]_ ;
  assign \new_[1604]_  = \new_[1603]_  | \new_[1568]_ ;
  assign \new_[1607]_  = \new_[874]_  | \new_[875]_ ;
  assign \new_[1610]_  = \new_[872]_  | \new_[873]_ ;
  assign \new_[1611]_  = \new_[1610]_  | \new_[1607]_ ;
  assign \new_[1614]_  = \new_[870]_  | \new_[871]_ ;
  assign \new_[1617]_  = \new_[868]_  | \new_[869]_ ;
  assign \new_[1618]_  = \new_[1617]_  | \new_[1614]_ ;
  assign \new_[1619]_  = \new_[1618]_  | \new_[1611]_ ;
  assign \new_[1622]_  = \new_[866]_  | \new_[867]_ ;
  assign \new_[1625]_  = \new_[864]_  | \new_[865]_ ;
  assign \new_[1626]_  = \new_[1625]_  | \new_[1622]_ ;
  assign \new_[1629]_  = \new_[862]_  | \new_[863]_ ;
  assign \new_[1633]_  = \new_[859]_  | \new_[860]_ ;
  assign \new_[1634]_  = \new_[861]_  | \new_[1633]_ ;
  assign \new_[1635]_  = \new_[1634]_  | \new_[1629]_ ;
  assign \new_[1636]_  = \new_[1635]_  | \new_[1626]_ ;
  assign \new_[1637]_  = \new_[1636]_  | \new_[1619]_ ;
  assign \new_[1640]_  = \new_[857]_  | \new_[858]_ ;
  assign \new_[1643]_  = \new_[855]_  | \new_[856]_ ;
  assign \new_[1644]_  = \new_[1643]_  | \new_[1640]_ ;
  assign \new_[1647]_  = \new_[853]_  | \new_[854]_ ;
  assign \new_[1651]_  = \new_[850]_  | \new_[851]_ ;
  assign \new_[1652]_  = \new_[852]_  | \new_[1651]_ ;
  assign \new_[1653]_  = \new_[1652]_  | \new_[1647]_ ;
  assign \new_[1654]_  = \new_[1653]_  | \new_[1644]_ ;
  assign \new_[1657]_  = \new_[848]_  | \new_[849]_ ;
  assign \new_[1660]_  = \new_[846]_  | \new_[847]_ ;
  assign \new_[1661]_  = \new_[1660]_  | \new_[1657]_ ;
  assign \new_[1664]_  = \new_[844]_  | \new_[845]_ ;
  assign \new_[1668]_  = \new_[841]_  | \new_[842]_ ;
  assign \new_[1669]_  = \new_[843]_  | \new_[1668]_ ;
  assign \new_[1670]_  = \new_[1669]_  | \new_[1664]_ ;
  assign \new_[1671]_  = \new_[1670]_  | \new_[1661]_ ;
  assign \new_[1672]_  = \new_[1671]_  | \new_[1654]_ ;
  assign \new_[1673]_  = \new_[1672]_  | \new_[1637]_ ;
  assign \new_[1674]_  = \new_[1673]_  | \new_[1604]_ ;
  assign \new_[1675]_  = \new_[1674]_  | \new_[1535]_ ;
  assign \new_[1676]_  = \new_[1675]_  | \new_[1396]_ ;
  assign \new_[1679]_  = \new_[839]_  | \new_[840]_ ;
  assign \new_[1682]_  = \new_[837]_  | \new_[838]_ ;
  assign \new_[1683]_  = \new_[1682]_  | \new_[1679]_ ;
  assign \new_[1686]_  = \new_[835]_  | \new_[836]_ ;
  assign \new_[1689]_  = \new_[833]_  | \new_[834]_ ;
  assign \new_[1690]_  = \new_[1689]_  | \new_[1686]_ ;
  assign \new_[1691]_  = \new_[1690]_  | \new_[1683]_ ;
  assign \new_[1694]_  = \new_[831]_  | \new_[832]_ ;
  assign \new_[1697]_  = \new_[829]_  | \new_[830]_ ;
  assign \new_[1698]_  = \new_[1697]_  | \new_[1694]_ ;
  assign \new_[1701]_  = \new_[827]_  | \new_[828]_ ;
  assign \new_[1705]_  = \new_[824]_  | \new_[825]_ ;
  assign \new_[1706]_  = \new_[826]_  | \new_[1705]_ ;
  assign \new_[1707]_  = \new_[1706]_  | \new_[1701]_ ;
  assign \new_[1708]_  = \new_[1707]_  | \new_[1698]_ ;
  assign \new_[1709]_  = \new_[1708]_  | \new_[1691]_ ;
  assign \new_[1712]_  = \new_[822]_  | \new_[823]_ ;
  assign \new_[1715]_  = \new_[820]_  | \new_[821]_ ;
  assign \new_[1716]_  = \new_[1715]_  | \new_[1712]_ ;
  assign \new_[1719]_  = \new_[818]_  | \new_[819]_ ;
  assign \new_[1723]_  = \new_[815]_  | \new_[816]_ ;
  assign \new_[1724]_  = \new_[817]_  | \new_[1723]_ ;
  assign \new_[1725]_  = \new_[1724]_  | \new_[1719]_ ;
  assign \new_[1726]_  = \new_[1725]_  | \new_[1716]_ ;
  assign \new_[1729]_  = \new_[813]_  | \new_[814]_ ;
  assign \new_[1732]_  = \new_[811]_  | \new_[812]_ ;
  assign \new_[1733]_  = \new_[1732]_  | \new_[1729]_ ;
  assign \new_[1736]_  = \new_[809]_  | \new_[810]_ ;
  assign \new_[1740]_  = \new_[806]_  | \new_[807]_ ;
  assign \new_[1741]_  = \new_[808]_  | \new_[1740]_ ;
  assign \new_[1742]_  = \new_[1741]_  | \new_[1736]_ ;
  assign \new_[1743]_  = \new_[1742]_  | \new_[1733]_ ;
  assign \new_[1744]_  = \new_[1743]_  | \new_[1726]_ ;
  assign \new_[1745]_  = \new_[1744]_  | \new_[1709]_ ;
  assign \new_[1748]_  = \new_[804]_  | \new_[805]_ ;
  assign \new_[1751]_  = \new_[802]_  | \new_[803]_ ;
  assign \new_[1752]_  = \new_[1751]_  | \new_[1748]_ ;
  assign \new_[1755]_  = \new_[800]_  | \new_[801]_ ;
  assign \new_[1758]_  = \new_[798]_  | \new_[799]_ ;
  assign \new_[1759]_  = \new_[1758]_  | \new_[1755]_ ;
  assign \new_[1760]_  = \new_[1759]_  | \new_[1752]_ ;
  assign \new_[1763]_  = \new_[796]_  | \new_[797]_ ;
  assign \new_[1766]_  = \new_[794]_  | \new_[795]_ ;
  assign \new_[1767]_  = \new_[1766]_  | \new_[1763]_ ;
  assign \new_[1770]_  = \new_[792]_  | \new_[793]_ ;
  assign \new_[1774]_  = \new_[789]_  | \new_[790]_ ;
  assign \new_[1775]_  = \new_[791]_  | \new_[1774]_ ;
  assign \new_[1776]_  = \new_[1775]_  | \new_[1770]_ ;
  assign \new_[1777]_  = \new_[1776]_  | \new_[1767]_ ;
  assign \new_[1778]_  = \new_[1777]_  | \new_[1760]_ ;
  assign \new_[1781]_  = \new_[787]_  | \new_[788]_ ;
  assign \new_[1784]_  = \new_[785]_  | \new_[786]_ ;
  assign \new_[1785]_  = \new_[1784]_  | \new_[1781]_ ;
  assign \new_[1788]_  = \new_[783]_  | \new_[784]_ ;
  assign \new_[1792]_  = \new_[780]_  | \new_[781]_ ;
  assign \new_[1793]_  = \new_[782]_  | \new_[1792]_ ;
  assign \new_[1794]_  = \new_[1793]_  | \new_[1788]_ ;
  assign \new_[1795]_  = \new_[1794]_  | \new_[1785]_ ;
  assign \new_[1798]_  = \new_[778]_  | \new_[779]_ ;
  assign \new_[1801]_  = \new_[776]_  | \new_[777]_ ;
  assign \new_[1802]_  = \new_[1801]_  | \new_[1798]_ ;
  assign \new_[1805]_  = \new_[774]_  | \new_[775]_ ;
  assign \new_[1809]_  = \new_[771]_  | \new_[772]_ ;
  assign \new_[1810]_  = \new_[773]_  | \new_[1809]_ ;
  assign \new_[1811]_  = \new_[1810]_  | \new_[1805]_ ;
  assign \new_[1812]_  = \new_[1811]_  | \new_[1802]_ ;
  assign \new_[1813]_  = \new_[1812]_  | \new_[1795]_ ;
  assign \new_[1814]_  = \new_[1813]_  | \new_[1778]_ ;
  assign \new_[1815]_  = \new_[1814]_  | \new_[1745]_ ;
  assign \new_[1818]_  = \new_[769]_  | \new_[770]_ ;
  assign \new_[1821]_  = \new_[767]_  | \new_[768]_ ;
  assign \new_[1822]_  = \new_[1821]_  | \new_[1818]_ ;
  assign \new_[1825]_  = \new_[765]_  | \new_[766]_ ;
  assign \new_[1828]_  = \new_[763]_  | \new_[764]_ ;
  assign \new_[1829]_  = \new_[1828]_  | \new_[1825]_ ;
  assign \new_[1830]_  = \new_[1829]_  | \new_[1822]_ ;
  assign \new_[1833]_  = \new_[761]_  | \new_[762]_ ;
  assign \new_[1836]_  = \new_[759]_  | \new_[760]_ ;
  assign \new_[1837]_  = \new_[1836]_  | \new_[1833]_ ;
  assign \new_[1840]_  = \new_[757]_  | \new_[758]_ ;
  assign \new_[1844]_  = \new_[754]_  | \new_[755]_ ;
  assign \new_[1845]_  = \new_[756]_  | \new_[1844]_ ;
  assign \new_[1846]_  = \new_[1845]_  | \new_[1840]_ ;
  assign \new_[1847]_  = \new_[1846]_  | \new_[1837]_ ;
  assign \new_[1848]_  = \new_[1847]_  | \new_[1830]_ ;
  assign \new_[1851]_  = \new_[752]_  | \new_[753]_ ;
  assign \new_[1854]_  = \new_[750]_  | \new_[751]_ ;
  assign \new_[1855]_  = \new_[1854]_  | \new_[1851]_ ;
  assign \new_[1858]_  = \new_[748]_  | \new_[749]_ ;
  assign \new_[1862]_  = \new_[745]_  | \new_[746]_ ;
  assign \new_[1863]_  = \new_[747]_  | \new_[1862]_ ;
  assign \new_[1864]_  = \new_[1863]_  | \new_[1858]_ ;
  assign \new_[1865]_  = \new_[1864]_  | \new_[1855]_ ;
  assign \new_[1868]_  = \new_[743]_  | \new_[744]_ ;
  assign \new_[1871]_  = \new_[741]_  | \new_[742]_ ;
  assign \new_[1872]_  = \new_[1871]_  | \new_[1868]_ ;
  assign \new_[1875]_  = \new_[739]_  | \new_[740]_ ;
  assign \new_[1879]_  = \new_[736]_  | \new_[737]_ ;
  assign \new_[1880]_  = \new_[738]_  | \new_[1879]_ ;
  assign \new_[1881]_  = \new_[1880]_  | \new_[1875]_ ;
  assign \new_[1882]_  = \new_[1881]_  | \new_[1872]_ ;
  assign \new_[1883]_  = \new_[1882]_  | \new_[1865]_ ;
  assign \new_[1884]_  = \new_[1883]_  | \new_[1848]_ ;
  assign \new_[1887]_  = \new_[734]_  | \new_[735]_ ;
  assign \new_[1890]_  = \new_[732]_  | \new_[733]_ ;
  assign \new_[1891]_  = \new_[1890]_  | \new_[1887]_ ;
  assign \new_[1894]_  = \new_[730]_  | \new_[731]_ ;
  assign \new_[1897]_  = \new_[728]_  | \new_[729]_ ;
  assign \new_[1898]_  = \new_[1897]_  | \new_[1894]_ ;
  assign \new_[1899]_  = \new_[1898]_  | \new_[1891]_ ;
  assign \new_[1902]_  = \new_[726]_  | \new_[727]_ ;
  assign \new_[1905]_  = \new_[724]_  | \new_[725]_ ;
  assign \new_[1906]_  = \new_[1905]_  | \new_[1902]_ ;
  assign \new_[1909]_  = \new_[722]_  | \new_[723]_ ;
  assign \new_[1913]_  = \new_[719]_  | \new_[720]_ ;
  assign \new_[1914]_  = \new_[721]_  | \new_[1913]_ ;
  assign \new_[1915]_  = \new_[1914]_  | \new_[1909]_ ;
  assign \new_[1916]_  = \new_[1915]_  | \new_[1906]_ ;
  assign \new_[1917]_  = \new_[1916]_  | \new_[1899]_ ;
  assign \new_[1920]_  = \new_[717]_  | \new_[718]_ ;
  assign \new_[1923]_  = \new_[715]_  | \new_[716]_ ;
  assign \new_[1924]_  = \new_[1923]_  | \new_[1920]_ ;
  assign \new_[1927]_  = \new_[713]_  | \new_[714]_ ;
  assign \new_[1931]_  = \new_[710]_  | \new_[711]_ ;
  assign \new_[1932]_  = \new_[712]_  | \new_[1931]_ ;
  assign \new_[1933]_  = \new_[1932]_  | \new_[1927]_ ;
  assign \new_[1934]_  = \new_[1933]_  | \new_[1924]_ ;
  assign \new_[1937]_  = \new_[708]_  | \new_[709]_ ;
  assign \new_[1940]_  = \new_[706]_  | \new_[707]_ ;
  assign \new_[1941]_  = \new_[1940]_  | \new_[1937]_ ;
  assign \new_[1944]_  = \new_[704]_  | \new_[705]_ ;
  assign \new_[1948]_  = \new_[701]_  | \new_[702]_ ;
  assign \new_[1949]_  = \new_[703]_  | \new_[1948]_ ;
  assign \new_[1950]_  = \new_[1949]_  | \new_[1944]_ ;
  assign \new_[1951]_  = \new_[1950]_  | \new_[1941]_ ;
  assign \new_[1952]_  = \new_[1951]_  | \new_[1934]_ ;
  assign \new_[1953]_  = \new_[1952]_  | \new_[1917]_ ;
  assign \new_[1954]_  = \new_[1953]_  | \new_[1884]_ ;
  assign \new_[1955]_  = \new_[1954]_  | \new_[1815]_ ;
  assign \new_[1958]_  = \new_[699]_  | \new_[700]_ ;
  assign \new_[1961]_  = \new_[697]_  | \new_[698]_ ;
  assign \new_[1962]_  = \new_[1961]_  | \new_[1958]_ ;
  assign \new_[1965]_  = \new_[695]_  | \new_[696]_ ;
  assign \new_[1968]_  = \new_[693]_  | \new_[694]_ ;
  assign \new_[1969]_  = \new_[1968]_  | \new_[1965]_ ;
  assign \new_[1970]_  = \new_[1969]_  | \new_[1962]_ ;
  assign \new_[1973]_  = \new_[691]_  | \new_[692]_ ;
  assign \new_[1976]_  = \new_[689]_  | \new_[690]_ ;
  assign \new_[1977]_  = \new_[1976]_  | \new_[1973]_ ;
  assign \new_[1980]_  = \new_[687]_  | \new_[688]_ ;
  assign \new_[1984]_  = \new_[684]_  | \new_[685]_ ;
  assign \new_[1985]_  = \new_[686]_  | \new_[1984]_ ;
  assign \new_[1986]_  = \new_[1985]_  | \new_[1980]_ ;
  assign \new_[1987]_  = \new_[1986]_  | \new_[1977]_ ;
  assign \new_[1988]_  = \new_[1987]_  | \new_[1970]_ ;
  assign \new_[1991]_  = \new_[682]_  | \new_[683]_ ;
  assign \new_[1994]_  = \new_[680]_  | \new_[681]_ ;
  assign \new_[1995]_  = \new_[1994]_  | \new_[1991]_ ;
  assign \new_[1998]_  = \new_[678]_  | \new_[679]_ ;
  assign \new_[2002]_  = \new_[675]_  | \new_[676]_ ;
  assign \new_[2003]_  = \new_[677]_  | \new_[2002]_ ;
  assign \new_[2004]_  = \new_[2003]_  | \new_[1998]_ ;
  assign \new_[2005]_  = \new_[2004]_  | \new_[1995]_ ;
  assign \new_[2008]_  = \new_[673]_  | \new_[674]_ ;
  assign \new_[2011]_  = \new_[671]_  | \new_[672]_ ;
  assign \new_[2012]_  = \new_[2011]_  | \new_[2008]_ ;
  assign \new_[2015]_  = \new_[669]_  | \new_[670]_ ;
  assign \new_[2019]_  = \new_[666]_  | \new_[667]_ ;
  assign \new_[2020]_  = \new_[668]_  | \new_[2019]_ ;
  assign \new_[2021]_  = \new_[2020]_  | \new_[2015]_ ;
  assign \new_[2022]_  = \new_[2021]_  | \new_[2012]_ ;
  assign \new_[2023]_  = \new_[2022]_  | \new_[2005]_ ;
  assign \new_[2024]_  = \new_[2023]_  | \new_[1988]_ ;
  assign \new_[2027]_  = \new_[664]_  | \new_[665]_ ;
  assign \new_[2030]_  = \new_[662]_  | \new_[663]_ ;
  assign \new_[2031]_  = \new_[2030]_  | \new_[2027]_ ;
  assign \new_[2034]_  = \new_[660]_  | \new_[661]_ ;
  assign \new_[2037]_  = \new_[658]_  | \new_[659]_ ;
  assign \new_[2038]_  = \new_[2037]_  | \new_[2034]_ ;
  assign \new_[2039]_  = \new_[2038]_  | \new_[2031]_ ;
  assign \new_[2042]_  = \new_[656]_  | \new_[657]_ ;
  assign \new_[2045]_  = \new_[654]_  | \new_[655]_ ;
  assign \new_[2046]_  = \new_[2045]_  | \new_[2042]_ ;
  assign \new_[2049]_  = \new_[652]_  | \new_[653]_ ;
  assign \new_[2053]_  = \new_[649]_  | \new_[650]_ ;
  assign \new_[2054]_  = \new_[651]_  | \new_[2053]_ ;
  assign \new_[2055]_  = \new_[2054]_  | \new_[2049]_ ;
  assign \new_[2056]_  = \new_[2055]_  | \new_[2046]_ ;
  assign \new_[2057]_  = \new_[2056]_  | \new_[2039]_ ;
  assign \new_[2060]_  = \new_[647]_  | \new_[648]_ ;
  assign \new_[2063]_  = \new_[645]_  | \new_[646]_ ;
  assign \new_[2064]_  = \new_[2063]_  | \new_[2060]_ ;
  assign \new_[2067]_  = \new_[643]_  | \new_[644]_ ;
  assign \new_[2071]_  = \new_[640]_  | \new_[641]_ ;
  assign \new_[2072]_  = \new_[642]_  | \new_[2071]_ ;
  assign \new_[2073]_  = \new_[2072]_  | \new_[2067]_ ;
  assign \new_[2074]_  = \new_[2073]_  | \new_[2064]_ ;
  assign \new_[2077]_  = \new_[638]_  | \new_[639]_ ;
  assign \new_[2080]_  = \new_[636]_  | \new_[637]_ ;
  assign \new_[2081]_  = \new_[2080]_  | \new_[2077]_ ;
  assign \new_[2084]_  = \new_[634]_  | \new_[635]_ ;
  assign \new_[2088]_  = \new_[631]_  | \new_[632]_ ;
  assign \new_[2089]_  = \new_[633]_  | \new_[2088]_ ;
  assign \new_[2090]_  = \new_[2089]_  | \new_[2084]_ ;
  assign \new_[2091]_  = \new_[2090]_  | \new_[2081]_ ;
  assign \new_[2092]_  = \new_[2091]_  | \new_[2074]_ ;
  assign \new_[2093]_  = \new_[2092]_  | \new_[2057]_ ;
  assign \new_[2094]_  = \new_[2093]_  | \new_[2024]_ ;
  assign \new_[2097]_  = \new_[629]_  | \new_[630]_ ;
  assign \new_[2100]_  = \new_[627]_  | \new_[628]_ ;
  assign \new_[2101]_  = \new_[2100]_  | \new_[2097]_ ;
  assign \new_[2104]_  = \new_[625]_  | \new_[626]_ ;
  assign \new_[2107]_  = \new_[623]_  | \new_[624]_ ;
  assign \new_[2108]_  = \new_[2107]_  | \new_[2104]_ ;
  assign \new_[2109]_  = \new_[2108]_  | \new_[2101]_ ;
  assign \new_[2112]_  = \new_[621]_  | \new_[622]_ ;
  assign \new_[2115]_  = \new_[619]_  | \new_[620]_ ;
  assign \new_[2116]_  = \new_[2115]_  | \new_[2112]_ ;
  assign \new_[2119]_  = \new_[617]_  | \new_[618]_ ;
  assign \new_[2123]_  = \new_[614]_  | \new_[615]_ ;
  assign \new_[2124]_  = \new_[616]_  | \new_[2123]_ ;
  assign \new_[2125]_  = \new_[2124]_  | \new_[2119]_ ;
  assign \new_[2126]_  = \new_[2125]_  | \new_[2116]_ ;
  assign \new_[2127]_  = \new_[2126]_  | \new_[2109]_ ;
  assign \new_[2130]_  = \new_[612]_  | \new_[613]_ ;
  assign \new_[2133]_  = \new_[610]_  | \new_[611]_ ;
  assign \new_[2134]_  = \new_[2133]_  | \new_[2130]_ ;
  assign \new_[2137]_  = \new_[608]_  | \new_[609]_ ;
  assign \new_[2141]_  = \new_[605]_  | \new_[606]_ ;
  assign \new_[2142]_  = \new_[607]_  | \new_[2141]_ ;
  assign \new_[2143]_  = \new_[2142]_  | \new_[2137]_ ;
  assign \new_[2144]_  = \new_[2143]_  | \new_[2134]_ ;
  assign \new_[2147]_  = \new_[603]_  | \new_[604]_ ;
  assign \new_[2150]_  = \new_[601]_  | \new_[602]_ ;
  assign \new_[2151]_  = \new_[2150]_  | \new_[2147]_ ;
  assign \new_[2154]_  = \new_[599]_  | \new_[600]_ ;
  assign \new_[2158]_  = \new_[596]_  | \new_[597]_ ;
  assign \new_[2159]_  = \new_[598]_  | \new_[2158]_ ;
  assign \new_[2160]_  = \new_[2159]_  | \new_[2154]_ ;
  assign \new_[2161]_  = \new_[2160]_  | \new_[2151]_ ;
  assign \new_[2162]_  = \new_[2161]_  | \new_[2144]_ ;
  assign \new_[2163]_  = \new_[2162]_  | \new_[2127]_ ;
  assign \new_[2166]_  = \new_[594]_  | \new_[595]_ ;
  assign \new_[2169]_  = \new_[592]_  | \new_[593]_ ;
  assign \new_[2170]_  = \new_[2169]_  | \new_[2166]_ ;
  assign \new_[2173]_  = \new_[590]_  | \new_[591]_ ;
  assign \new_[2176]_  = \new_[588]_  | \new_[589]_ ;
  assign \new_[2177]_  = \new_[2176]_  | \new_[2173]_ ;
  assign \new_[2178]_  = \new_[2177]_  | \new_[2170]_ ;
  assign \new_[2181]_  = \new_[586]_  | \new_[587]_ ;
  assign \new_[2184]_  = \new_[584]_  | \new_[585]_ ;
  assign \new_[2185]_  = \new_[2184]_  | \new_[2181]_ ;
  assign \new_[2188]_  = \new_[582]_  | \new_[583]_ ;
  assign \new_[2192]_  = \new_[579]_  | \new_[580]_ ;
  assign \new_[2193]_  = \new_[581]_  | \new_[2192]_ ;
  assign \new_[2194]_  = \new_[2193]_  | \new_[2188]_ ;
  assign \new_[2195]_  = \new_[2194]_  | \new_[2185]_ ;
  assign \new_[2196]_  = \new_[2195]_  | \new_[2178]_ ;
  assign \new_[2199]_  = \new_[577]_  | \new_[578]_ ;
  assign \new_[2202]_  = \new_[575]_  | \new_[576]_ ;
  assign \new_[2203]_  = \new_[2202]_  | \new_[2199]_ ;
  assign \new_[2206]_  = \new_[573]_  | \new_[574]_ ;
  assign \new_[2210]_  = \new_[570]_  | \new_[571]_ ;
  assign \new_[2211]_  = \new_[572]_  | \new_[2210]_ ;
  assign \new_[2212]_  = \new_[2211]_  | \new_[2206]_ ;
  assign \new_[2213]_  = \new_[2212]_  | \new_[2203]_ ;
  assign \new_[2216]_  = \new_[568]_  | \new_[569]_ ;
  assign \new_[2219]_  = \new_[566]_  | \new_[567]_ ;
  assign \new_[2220]_  = \new_[2219]_  | \new_[2216]_ ;
  assign \new_[2223]_  = \new_[564]_  | \new_[565]_ ;
  assign \new_[2227]_  = \new_[561]_  | \new_[562]_ ;
  assign \new_[2228]_  = \new_[563]_  | \new_[2227]_ ;
  assign \new_[2229]_  = \new_[2228]_  | \new_[2223]_ ;
  assign \new_[2230]_  = \new_[2229]_  | \new_[2220]_ ;
  assign \new_[2231]_  = \new_[2230]_  | \new_[2213]_ ;
  assign \new_[2232]_  = \new_[2231]_  | \new_[2196]_ ;
  assign \new_[2233]_  = \new_[2232]_  | \new_[2163]_ ;
  assign \new_[2234]_  = \new_[2233]_  | \new_[2094]_ ;
  assign \new_[2235]_  = \new_[2234]_  | \new_[1955]_ ;
  assign \new_[2236]_  = \new_[2235]_  | \new_[1676]_ ;
  assign \new_[2239]_  = \new_[559]_  | \new_[560]_ ;
  assign \new_[2242]_  = \new_[557]_  | \new_[558]_ ;
  assign \new_[2243]_  = \new_[2242]_  | \new_[2239]_ ;
  assign \new_[2246]_  = \new_[555]_  | \new_[556]_ ;
  assign \new_[2249]_  = \new_[553]_  | \new_[554]_ ;
  assign \new_[2250]_  = \new_[2249]_  | \new_[2246]_ ;
  assign \new_[2251]_  = \new_[2250]_  | \new_[2243]_ ;
  assign \new_[2254]_  = \new_[551]_  | \new_[552]_ ;
  assign \new_[2257]_  = \new_[549]_  | \new_[550]_ ;
  assign \new_[2258]_  = \new_[2257]_  | \new_[2254]_ ;
  assign \new_[2261]_  = \new_[547]_  | \new_[548]_ ;
  assign \new_[2265]_  = \new_[544]_  | \new_[545]_ ;
  assign \new_[2266]_  = \new_[546]_  | \new_[2265]_ ;
  assign \new_[2267]_  = \new_[2266]_  | \new_[2261]_ ;
  assign \new_[2268]_  = \new_[2267]_  | \new_[2258]_ ;
  assign \new_[2269]_  = \new_[2268]_  | \new_[2251]_ ;
  assign \new_[2272]_  = \new_[542]_  | \new_[543]_ ;
  assign \new_[2275]_  = \new_[540]_  | \new_[541]_ ;
  assign \new_[2276]_  = \new_[2275]_  | \new_[2272]_ ;
  assign \new_[2279]_  = \new_[538]_  | \new_[539]_ ;
  assign \new_[2283]_  = \new_[535]_  | \new_[536]_ ;
  assign \new_[2284]_  = \new_[537]_  | \new_[2283]_ ;
  assign \new_[2285]_  = \new_[2284]_  | \new_[2279]_ ;
  assign \new_[2286]_  = \new_[2285]_  | \new_[2276]_ ;
  assign \new_[2289]_  = \new_[533]_  | \new_[534]_ ;
  assign \new_[2292]_  = \new_[531]_  | \new_[532]_ ;
  assign \new_[2293]_  = \new_[2292]_  | \new_[2289]_ ;
  assign \new_[2296]_  = \new_[529]_  | \new_[530]_ ;
  assign \new_[2300]_  = \new_[526]_  | \new_[527]_ ;
  assign \new_[2301]_  = \new_[528]_  | \new_[2300]_ ;
  assign \new_[2302]_  = \new_[2301]_  | \new_[2296]_ ;
  assign \new_[2303]_  = \new_[2302]_  | \new_[2293]_ ;
  assign \new_[2304]_  = \new_[2303]_  | \new_[2286]_ ;
  assign \new_[2305]_  = \new_[2304]_  | \new_[2269]_ ;
  assign \new_[2308]_  = \new_[524]_  | \new_[525]_ ;
  assign \new_[2311]_  = \new_[522]_  | \new_[523]_ ;
  assign \new_[2312]_  = \new_[2311]_  | \new_[2308]_ ;
  assign \new_[2315]_  = \new_[520]_  | \new_[521]_ ;
  assign \new_[2318]_  = \new_[518]_  | \new_[519]_ ;
  assign \new_[2319]_  = \new_[2318]_  | \new_[2315]_ ;
  assign \new_[2320]_  = \new_[2319]_  | \new_[2312]_ ;
  assign \new_[2323]_  = \new_[516]_  | \new_[517]_ ;
  assign \new_[2326]_  = \new_[514]_  | \new_[515]_ ;
  assign \new_[2327]_  = \new_[2326]_  | \new_[2323]_ ;
  assign \new_[2330]_  = \new_[512]_  | \new_[513]_ ;
  assign \new_[2334]_  = \new_[509]_  | \new_[510]_ ;
  assign \new_[2335]_  = \new_[511]_  | \new_[2334]_ ;
  assign \new_[2336]_  = \new_[2335]_  | \new_[2330]_ ;
  assign \new_[2337]_  = \new_[2336]_  | \new_[2327]_ ;
  assign \new_[2338]_  = \new_[2337]_  | \new_[2320]_ ;
  assign \new_[2341]_  = \new_[507]_  | \new_[508]_ ;
  assign \new_[2344]_  = \new_[505]_  | \new_[506]_ ;
  assign \new_[2345]_  = \new_[2344]_  | \new_[2341]_ ;
  assign \new_[2348]_  = \new_[503]_  | \new_[504]_ ;
  assign \new_[2352]_  = \new_[500]_  | \new_[501]_ ;
  assign \new_[2353]_  = \new_[502]_  | \new_[2352]_ ;
  assign \new_[2354]_  = \new_[2353]_  | \new_[2348]_ ;
  assign \new_[2355]_  = \new_[2354]_  | \new_[2345]_ ;
  assign \new_[2358]_  = \new_[498]_  | \new_[499]_ ;
  assign \new_[2361]_  = \new_[496]_  | \new_[497]_ ;
  assign \new_[2362]_  = \new_[2361]_  | \new_[2358]_ ;
  assign \new_[2365]_  = \new_[494]_  | \new_[495]_ ;
  assign \new_[2369]_  = \new_[491]_  | \new_[492]_ ;
  assign \new_[2370]_  = \new_[493]_  | \new_[2369]_ ;
  assign \new_[2371]_  = \new_[2370]_  | \new_[2365]_ ;
  assign \new_[2372]_  = \new_[2371]_  | \new_[2362]_ ;
  assign \new_[2373]_  = \new_[2372]_  | \new_[2355]_ ;
  assign \new_[2374]_  = \new_[2373]_  | \new_[2338]_ ;
  assign \new_[2375]_  = \new_[2374]_  | \new_[2305]_ ;
  assign \new_[2378]_  = \new_[489]_  | \new_[490]_ ;
  assign \new_[2381]_  = \new_[487]_  | \new_[488]_ ;
  assign \new_[2382]_  = \new_[2381]_  | \new_[2378]_ ;
  assign \new_[2385]_  = \new_[485]_  | \new_[486]_ ;
  assign \new_[2388]_  = \new_[483]_  | \new_[484]_ ;
  assign \new_[2389]_  = \new_[2388]_  | \new_[2385]_ ;
  assign \new_[2390]_  = \new_[2389]_  | \new_[2382]_ ;
  assign \new_[2393]_  = \new_[481]_  | \new_[482]_ ;
  assign \new_[2396]_  = \new_[479]_  | \new_[480]_ ;
  assign \new_[2397]_  = \new_[2396]_  | \new_[2393]_ ;
  assign \new_[2400]_  = \new_[477]_  | \new_[478]_ ;
  assign \new_[2404]_  = \new_[474]_  | \new_[475]_ ;
  assign \new_[2405]_  = \new_[476]_  | \new_[2404]_ ;
  assign \new_[2406]_  = \new_[2405]_  | \new_[2400]_ ;
  assign \new_[2407]_  = \new_[2406]_  | \new_[2397]_ ;
  assign \new_[2408]_  = \new_[2407]_  | \new_[2390]_ ;
  assign \new_[2411]_  = \new_[472]_  | \new_[473]_ ;
  assign \new_[2414]_  = \new_[470]_  | \new_[471]_ ;
  assign \new_[2415]_  = \new_[2414]_  | \new_[2411]_ ;
  assign \new_[2418]_  = \new_[468]_  | \new_[469]_ ;
  assign \new_[2422]_  = \new_[465]_  | \new_[466]_ ;
  assign \new_[2423]_  = \new_[467]_  | \new_[2422]_ ;
  assign \new_[2424]_  = \new_[2423]_  | \new_[2418]_ ;
  assign \new_[2425]_  = \new_[2424]_  | \new_[2415]_ ;
  assign \new_[2428]_  = \new_[463]_  | \new_[464]_ ;
  assign \new_[2431]_  = \new_[461]_  | \new_[462]_ ;
  assign \new_[2432]_  = \new_[2431]_  | \new_[2428]_ ;
  assign \new_[2435]_  = \new_[459]_  | \new_[460]_ ;
  assign \new_[2439]_  = \new_[456]_  | \new_[457]_ ;
  assign \new_[2440]_  = \new_[458]_  | \new_[2439]_ ;
  assign \new_[2441]_  = \new_[2440]_  | \new_[2435]_ ;
  assign \new_[2442]_  = \new_[2441]_  | \new_[2432]_ ;
  assign \new_[2443]_  = \new_[2442]_  | \new_[2425]_ ;
  assign \new_[2444]_  = \new_[2443]_  | \new_[2408]_ ;
  assign \new_[2447]_  = \new_[454]_  | \new_[455]_ ;
  assign \new_[2450]_  = \new_[452]_  | \new_[453]_ ;
  assign \new_[2451]_  = \new_[2450]_  | \new_[2447]_ ;
  assign \new_[2454]_  = \new_[450]_  | \new_[451]_ ;
  assign \new_[2457]_  = \new_[448]_  | \new_[449]_ ;
  assign \new_[2458]_  = \new_[2457]_  | \new_[2454]_ ;
  assign \new_[2459]_  = \new_[2458]_  | \new_[2451]_ ;
  assign \new_[2462]_  = \new_[446]_  | \new_[447]_ ;
  assign \new_[2465]_  = \new_[444]_  | \new_[445]_ ;
  assign \new_[2466]_  = \new_[2465]_  | \new_[2462]_ ;
  assign \new_[2469]_  = \new_[442]_  | \new_[443]_ ;
  assign \new_[2473]_  = \new_[439]_  | \new_[440]_ ;
  assign \new_[2474]_  = \new_[441]_  | \new_[2473]_ ;
  assign \new_[2475]_  = \new_[2474]_  | \new_[2469]_ ;
  assign \new_[2476]_  = \new_[2475]_  | \new_[2466]_ ;
  assign \new_[2477]_  = \new_[2476]_  | \new_[2459]_ ;
  assign \new_[2480]_  = \new_[437]_  | \new_[438]_ ;
  assign \new_[2483]_  = \new_[435]_  | \new_[436]_ ;
  assign \new_[2484]_  = \new_[2483]_  | \new_[2480]_ ;
  assign \new_[2487]_  = \new_[433]_  | \new_[434]_ ;
  assign \new_[2491]_  = \new_[430]_  | \new_[431]_ ;
  assign \new_[2492]_  = \new_[432]_  | \new_[2491]_ ;
  assign \new_[2493]_  = \new_[2492]_  | \new_[2487]_ ;
  assign \new_[2494]_  = \new_[2493]_  | \new_[2484]_ ;
  assign \new_[2497]_  = \new_[428]_  | \new_[429]_ ;
  assign \new_[2500]_  = \new_[426]_  | \new_[427]_ ;
  assign \new_[2501]_  = \new_[2500]_  | \new_[2497]_ ;
  assign \new_[2504]_  = \new_[424]_  | \new_[425]_ ;
  assign \new_[2508]_  = \new_[421]_  | \new_[422]_ ;
  assign \new_[2509]_  = \new_[423]_  | \new_[2508]_ ;
  assign \new_[2510]_  = \new_[2509]_  | \new_[2504]_ ;
  assign \new_[2511]_  = \new_[2510]_  | \new_[2501]_ ;
  assign \new_[2512]_  = \new_[2511]_  | \new_[2494]_ ;
  assign \new_[2513]_  = \new_[2512]_  | \new_[2477]_ ;
  assign \new_[2514]_  = \new_[2513]_  | \new_[2444]_ ;
  assign \new_[2515]_  = \new_[2514]_  | \new_[2375]_ ;
  assign \new_[2518]_  = \new_[419]_  | \new_[420]_ ;
  assign \new_[2521]_  = \new_[417]_  | \new_[418]_ ;
  assign \new_[2522]_  = \new_[2521]_  | \new_[2518]_ ;
  assign \new_[2525]_  = \new_[415]_  | \new_[416]_ ;
  assign \new_[2528]_  = \new_[413]_  | \new_[414]_ ;
  assign \new_[2529]_  = \new_[2528]_  | \new_[2525]_ ;
  assign \new_[2530]_  = \new_[2529]_  | \new_[2522]_ ;
  assign \new_[2533]_  = \new_[411]_  | \new_[412]_ ;
  assign \new_[2536]_  = \new_[409]_  | \new_[410]_ ;
  assign \new_[2537]_  = \new_[2536]_  | \new_[2533]_ ;
  assign \new_[2540]_  = \new_[407]_  | \new_[408]_ ;
  assign \new_[2544]_  = \new_[404]_  | \new_[405]_ ;
  assign \new_[2545]_  = \new_[406]_  | \new_[2544]_ ;
  assign \new_[2546]_  = \new_[2545]_  | \new_[2540]_ ;
  assign \new_[2547]_  = \new_[2546]_  | \new_[2537]_ ;
  assign \new_[2548]_  = \new_[2547]_  | \new_[2530]_ ;
  assign \new_[2551]_  = \new_[402]_  | \new_[403]_ ;
  assign \new_[2554]_  = \new_[400]_  | \new_[401]_ ;
  assign \new_[2555]_  = \new_[2554]_  | \new_[2551]_ ;
  assign \new_[2558]_  = \new_[398]_  | \new_[399]_ ;
  assign \new_[2562]_  = \new_[395]_  | \new_[396]_ ;
  assign \new_[2563]_  = \new_[397]_  | \new_[2562]_ ;
  assign \new_[2564]_  = \new_[2563]_  | \new_[2558]_ ;
  assign \new_[2565]_  = \new_[2564]_  | \new_[2555]_ ;
  assign \new_[2568]_  = \new_[393]_  | \new_[394]_ ;
  assign \new_[2571]_  = \new_[391]_  | \new_[392]_ ;
  assign \new_[2572]_  = \new_[2571]_  | \new_[2568]_ ;
  assign \new_[2575]_  = \new_[389]_  | \new_[390]_ ;
  assign \new_[2579]_  = \new_[386]_  | \new_[387]_ ;
  assign \new_[2580]_  = \new_[388]_  | \new_[2579]_ ;
  assign \new_[2581]_  = \new_[2580]_  | \new_[2575]_ ;
  assign \new_[2582]_  = \new_[2581]_  | \new_[2572]_ ;
  assign \new_[2583]_  = \new_[2582]_  | \new_[2565]_ ;
  assign \new_[2584]_  = \new_[2583]_  | \new_[2548]_ ;
  assign \new_[2587]_  = \new_[384]_  | \new_[385]_ ;
  assign \new_[2590]_  = \new_[382]_  | \new_[383]_ ;
  assign \new_[2591]_  = \new_[2590]_  | \new_[2587]_ ;
  assign \new_[2594]_  = \new_[380]_  | \new_[381]_ ;
  assign \new_[2597]_  = \new_[378]_  | \new_[379]_ ;
  assign \new_[2598]_  = \new_[2597]_  | \new_[2594]_ ;
  assign \new_[2599]_  = \new_[2598]_  | \new_[2591]_ ;
  assign \new_[2602]_  = \new_[376]_  | \new_[377]_ ;
  assign \new_[2605]_  = \new_[374]_  | \new_[375]_ ;
  assign \new_[2606]_  = \new_[2605]_  | \new_[2602]_ ;
  assign \new_[2609]_  = \new_[372]_  | \new_[373]_ ;
  assign \new_[2613]_  = \new_[369]_  | \new_[370]_ ;
  assign \new_[2614]_  = \new_[371]_  | \new_[2613]_ ;
  assign \new_[2615]_  = \new_[2614]_  | \new_[2609]_ ;
  assign \new_[2616]_  = \new_[2615]_  | \new_[2606]_ ;
  assign \new_[2617]_  = \new_[2616]_  | \new_[2599]_ ;
  assign \new_[2620]_  = \new_[367]_  | \new_[368]_ ;
  assign \new_[2623]_  = \new_[365]_  | \new_[366]_ ;
  assign \new_[2624]_  = \new_[2623]_  | \new_[2620]_ ;
  assign \new_[2627]_  = \new_[363]_  | \new_[364]_ ;
  assign \new_[2631]_  = \new_[360]_  | \new_[361]_ ;
  assign \new_[2632]_  = \new_[362]_  | \new_[2631]_ ;
  assign \new_[2633]_  = \new_[2632]_  | \new_[2627]_ ;
  assign \new_[2634]_  = \new_[2633]_  | \new_[2624]_ ;
  assign \new_[2637]_  = \new_[358]_  | \new_[359]_ ;
  assign \new_[2640]_  = \new_[356]_  | \new_[357]_ ;
  assign \new_[2641]_  = \new_[2640]_  | \new_[2637]_ ;
  assign \new_[2644]_  = \new_[354]_  | \new_[355]_ ;
  assign \new_[2648]_  = \new_[351]_  | \new_[352]_ ;
  assign \new_[2649]_  = \new_[353]_  | \new_[2648]_ ;
  assign \new_[2650]_  = \new_[2649]_  | \new_[2644]_ ;
  assign \new_[2651]_  = \new_[2650]_  | \new_[2641]_ ;
  assign \new_[2652]_  = \new_[2651]_  | \new_[2634]_ ;
  assign \new_[2653]_  = \new_[2652]_  | \new_[2617]_ ;
  assign \new_[2654]_  = \new_[2653]_  | \new_[2584]_ ;
  assign \new_[2657]_  = \new_[349]_  | \new_[350]_ ;
  assign \new_[2660]_  = \new_[347]_  | \new_[348]_ ;
  assign \new_[2661]_  = \new_[2660]_  | \new_[2657]_ ;
  assign \new_[2664]_  = \new_[345]_  | \new_[346]_ ;
  assign \new_[2667]_  = \new_[343]_  | \new_[344]_ ;
  assign \new_[2668]_  = \new_[2667]_  | \new_[2664]_ ;
  assign \new_[2669]_  = \new_[2668]_  | \new_[2661]_ ;
  assign \new_[2672]_  = \new_[341]_  | \new_[342]_ ;
  assign \new_[2675]_  = \new_[339]_  | \new_[340]_ ;
  assign \new_[2676]_  = \new_[2675]_  | \new_[2672]_ ;
  assign \new_[2679]_  = \new_[337]_  | \new_[338]_ ;
  assign \new_[2683]_  = \new_[334]_  | \new_[335]_ ;
  assign \new_[2684]_  = \new_[336]_  | \new_[2683]_ ;
  assign \new_[2685]_  = \new_[2684]_  | \new_[2679]_ ;
  assign \new_[2686]_  = \new_[2685]_  | \new_[2676]_ ;
  assign \new_[2687]_  = \new_[2686]_  | \new_[2669]_ ;
  assign \new_[2690]_  = \new_[332]_  | \new_[333]_ ;
  assign \new_[2693]_  = \new_[330]_  | \new_[331]_ ;
  assign \new_[2694]_  = \new_[2693]_  | \new_[2690]_ ;
  assign \new_[2697]_  = \new_[328]_  | \new_[329]_ ;
  assign \new_[2701]_  = \new_[325]_  | \new_[326]_ ;
  assign \new_[2702]_  = \new_[327]_  | \new_[2701]_ ;
  assign \new_[2703]_  = \new_[2702]_  | \new_[2697]_ ;
  assign \new_[2704]_  = \new_[2703]_  | \new_[2694]_ ;
  assign \new_[2707]_  = \new_[323]_  | \new_[324]_ ;
  assign \new_[2710]_  = \new_[321]_  | \new_[322]_ ;
  assign \new_[2711]_  = \new_[2710]_  | \new_[2707]_ ;
  assign \new_[2714]_  = \new_[319]_  | \new_[320]_ ;
  assign \new_[2718]_  = \new_[316]_  | \new_[317]_ ;
  assign \new_[2719]_  = \new_[318]_  | \new_[2718]_ ;
  assign \new_[2720]_  = \new_[2719]_  | \new_[2714]_ ;
  assign \new_[2721]_  = \new_[2720]_  | \new_[2711]_ ;
  assign \new_[2722]_  = \new_[2721]_  | \new_[2704]_ ;
  assign \new_[2723]_  = \new_[2722]_  | \new_[2687]_ ;
  assign \new_[2726]_  = \new_[314]_  | \new_[315]_ ;
  assign \new_[2729]_  = \new_[312]_  | \new_[313]_ ;
  assign \new_[2730]_  = \new_[2729]_  | \new_[2726]_ ;
  assign \new_[2733]_  = \new_[310]_  | \new_[311]_ ;
  assign \new_[2736]_  = \new_[308]_  | \new_[309]_ ;
  assign \new_[2737]_  = \new_[2736]_  | \new_[2733]_ ;
  assign \new_[2738]_  = \new_[2737]_  | \new_[2730]_ ;
  assign \new_[2741]_  = \new_[306]_  | \new_[307]_ ;
  assign \new_[2744]_  = \new_[304]_  | \new_[305]_ ;
  assign \new_[2745]_  = \new_[2744]_  | \new_[2741]_ ;
  assign \new_[2748]_  = \new_[302]_  | \new_[303]_ ;
  assign \new_[2752]_  = \new_[299]_  | \new_[300]_ ;
  assign \new_[2753]_  = \new_[301]_  | \new_[2752]_ ;
  assign \new_[2754]_  = \new_[2753]_  | \new_[2748]_ ;
  assign \new_[2755]_  = \new_[2754]_  | \new_[2745]_ ;
  assign \new_[2756]_  = \new_[2755]_  | \new_[2738]_ ;
  assign \new_[2759]_  = \new_[297]_  | \new_[298]_ ;
  assign \new_[2762]_  = \new_[295]_  | \new_[296]_ ;
  assign \new_[2763]_  = \new_[2762]_  | \new_[2759]_ ;
  assign \new_[2766]_  = \new_[293]_  | \new_[294]_ ;
  assign \new_[2770]_  = \new_[290]_  | \new_[291]_ ;
  assign \new_[2771]_  = \new_[292]_  | \new_[2770]_ ;
  assign \new_[2772]_  = \new_[2771]_  | \new_[2766]_ ;
  assign \new_[2773]_  = \new_[2772]_  | \new_[2763]_ ;
  assign \new_[2776]_  = \new_[288]_  | \new_[289]_ ;
  assign \new_[2779]_  = \new_[286]_  | \new_[287]_ ;
  assign \new_[2780]_  = \new_[2779]_  | \new_[2776]_ ;
  assign \new_[2783]_  = \new_[284]_  | \new_[285]_ ;
  assign \new_[2787]_  = \new_[281]_  | \new_[282]_ ;
  assign \new_[2788]_  = \new_[283]_  | \new_[2787]_ ;
  assign \new_[2789]_  = \new_[2788]_  | \new_[2783]_ ;
  assign \new_[2790]_  = \new_[2789]_  | \new_[2780]_ ;
  assign \new_[2791]_  = \new_[2790]_  | \new_[2773]_ ;
  assign \new_[2792]_  = \new_[2791]_  | \new_[2756]_ ;
  assign \new_[2793]_  = \new_[2792]_  | \new_[2723]_ ;
  assign \new_[2794]_  = \new_[2793]_  | \new_[2654]_ ;
  assign \new_[2795]_  = \new_[2794]_  | \new_[2515]_ ;
  assign \new_[2798]_  = \new_[279]_  | \new_[280]_ ;
  assign \new_[2801]_  = \new_[277]_  | \new_[278]_ ;
  assign \new_[2802]_  = \new_[2801]_  | \new_[2798]_ ;
  assign \new_[2805]_  = \new_[275]_  | \new_[276]_ ;
  assign \new_[2808]_  = \new_[273]_  | \new_[274]_ ;
  assign \new_[2809]_  = \new_[2808]_  | \new_[2805]_ ;
  assign \new_[2810]_  = \new_[2809]_  | \new_[2802]_ ;
  assign \new_[2813]_  = \new_[271]_  | \new_[272]_ ;
  assign \new_[2816]_  = \new_[269]_  | \new_[270]_ ;
  assign \new_[2817]_  = \new_[2816]_  | \new_[2813]_ ;
  assign \new_[2820]_  = \new_[267]_  | \new_[268]_ ;
  assign \new_[2824]_  = \new_[264]_  | \new_[265]_ ;
  assign \new_[2825]_  = \new_[266]_  | \new_[2824]_ ;
  assign \new_[2826]_  = \new_[2825]_  | \new_[2820]_ ;
  assign \new_[2827]_  = \new_[2826]_  | \new_[2817]_ ;
  assign \new_[2828]_  = \new_[2827]_  | \new_[2810]_ ;
  assign \new_[2831]_  = \new_[262]_  | \new_[263]_ ;
  assign \new_[2834]_  = \new_[260]_  | \new_[261]_ ;
  assign \new_[2835]_  = \new_[2834]_  | \new_[2831]_ ;
  assign \new_[2838]_  = \new_[258]_  | \new_[259]_ ;
  assign \new_[2842]_  = \new_[255]_  | \new_[256]_ ;
  assign \new_[2843]_  = \new_[257]_  | \new_[2842]_ ;
  assign \new_[2844]_  = \new_[2843]_  | \new_[2838]_ ;
  assign \new_[2845]_  = \new_[2844]_  | \new_[2835]_ ;
  assign \new_[2848]_  = \new_[253]_  | \new_[254]_ ;
  assign \new_[2851]_  = \new_[251]_  | \new_[252]_ ;
  assign \new_[2852]_  = \new_[2851]_  | \new_[2848]_ ;
  assign \new_[2855]_  = \new_[249]_  | \new_[250]_ ;
  assign \new_[2859]_  = \new_[246]_  | \new_[247]_ ;
  assign \new_[2860]_  = \new_[248]_  | \new_[2859]_ ;
  assign \new_[2861]_  = \new_[2860]_  | \new_[2855]_ ;
  assign \new_[2862]_  = \new_[2861]_  | \new_[2852]_ ;
  assign \new_[2863]_  = \new_[2862]_  | \new_[2845]_ ;
  assign \new_[2864]_  = \new_[2863]_  | \new_[2828]_ ;
  assign \new_[2867]_  = \new_[244]_  | \new_[245]_ ;
  assign \new_[2870]_  = \new_[242]_  | \new_[243]_ ;
  assign \new_[2871]_  = \new_[2870]_  | \new_[2867]_ ;
  assign \new_[2874]_  = \new_[240]_  | \new_[241]_ ;
  assign \new_[2877]_  = \new_[238]_  | \new_[239]_ ;
  assign \new_[2878]_  = \new_[2877]_  | \new_[2874]_ ;
  assign \new_[2879]_  = \new_[2878]_  | \new_[2871]_ ;
  assign \new_[2882]_  = \new_[236]_  | \new_[237]_ ;
  assign \new_[2885]_  = \new_[234]_  | \new_[235]_ ;
  assign \new_[2886]_  = \new_[2885]_  | \new_[2882]_ ;
  assign \new_[2889]_  = \new_[232]_  | \new_[233]_ ;
  assign \new_[2893]_  = \new_[229]_  | \new_[230]_ ;
  assign \new_[2894]_  = \new_[231]_  | \new_[2893]_ ;
  assign \new_[2895]_  = \new_[2894]_  | \new_[2889]_ ;
  assign \new_[2896]_  = \new_[2895]_  | \new_[2886]_ ;
  assign \new_[2897]_  = \new_[2896]_  | \new_[2879]_ ;
  assign \new_[2900]_  = \new_[227]_  | \new_[228]_ ;
  assign \new_[2903]_  = \new_[225]_  | \new_[226]_ ;
  assign \new_[2904]_  = \new_[2903]_  | \new_[2900]_ ;
  assign \new_[2907]_  = \new_[223]_  | \new_[224]_ ;
  assign \new_[2911]_  = \new_[220]_  | \new_[221]_ ;
  assign \new_[2912]_  = \new_[222]_  | \new_[2911]_ ;
  assign \new_[2913]_  = \new_[2912]_  | \new_[2907]_ ;
  assign \new_[2914]_  = \new_[2913]_  | \new_[2904]_ ;
  assign \new_[2917]_  = \new_[218]_  | \new_[219]_ ;
  assign \new_[2920]_  = \new_[216]_  | \new_[217]_ ;
  assign \new_[2921]_  = \new_[2920]_  | \new_[2917]_ ;
  assign \new_[2924]_  = \new_[214]_  | \new_[215]_ ;
  assign \new_[2928]_  = \new_[211]_  | \new_[212]_ ;
  assign \new_[2929]_  = \new_[213]_  | \new_[2928]_ ;
  assign \new_[2930]_  = \new_[2929]_  | \new_[2924]_ ;
  assign \new_[2931]_  = \new_[2930]_  | \new_[2921]_ ;
  assign \new_[2932]_  = \new_[2931]_  | \new_[2914]_ ;
  assign \new_[2933]_  = \new_[2932]_  | \new_[2897]_ ;
  assign \new_[2934]_  = \new_[2933]_  | \new_[2864]_ ;
  assign \new_[2937]_  = \new_[209]_  | \new_[210]_ ;
  assign \new_[2940]_  = \new_[207]_  | \new_[208]_ ;
  assign \new_[2941]_  = \new_[2940]_  | \new_[2937]_ ;
  assign \new_[2944]_  = \new_[205]_  | \new_[206]_ ;
  assign \new_[2947]_  = \new_[203]_  | \new_[204]_ ;
  assign \new_[2948]_  = \new_[2947]_  | \new_[2944]_ ;
  assign \new_[2949]_  = \new_[2948]_  | \new_[2941]_ ;
  assign \new_[2952]_  = \new_[201]_  | \new_[202]_ ;
  assign \new_[2955]_  = \new_[199]_  | \new_[200]_ ;
  assign \new_[2956]_  = \new_[2955]_  | \new_[2952]_ ;
  assign \new_[2959]_  = \new_[197]_  | \new_[198]_ ;
  assign \new_[2963]_  = \new_[194]_  | \new_[195]_ ;
  assign \new_[2964]_  = \new_[196]_  | \new_[2963]_ ;
  assign \new_[2965]_  = \new_[2964]_  | \new_[2959]_ ;
  assign \new_[2966]_  = \new_[2965]_  | \new_[2956]_ ;
  assign \new_[2967]_  = \new_[2966]_  | \new_[2949]_ ;
  assign \new_[2970]_  = \new_[192]_  | \new_[193]_ ;
  assign \new_[2973]_  = \new_[190]_  | \new_[191]_ ;
  assign \new_[2974]_  = \new_[2973]_  | \new_[2970]_ ;
  assign \new_[2977]_  = \new_[188]_  | \new_[189]_ ;
  assign \new_[2981]_  = \new_[185]_  | \new_[186]_ ;
  assign \new_[2982]_  = \new_[187]_  | \new_[2981]_ ;
  assign \new_[2983]_  = \new_[2982]_  | \new_[2977]_ ;
  assign \new_[2984]_  = \new_[2983]_  | \new_[2974]_ ;
  assign \new_[2987]_  = \new_[183]_  | \new_[184]_ ;
  assign \new_[2990]_  = \new_[181]_  | \new_[182]_ ;
  assign \new_[2991]_  = \new_[2990]_  | \new_[2987]_ ;
  assign \new_[2994]_  = \new_[179]_  | \new_[180]_ ;
  assign \new_[2998]_  = \new_[176]_  | \new_[177]_ ;
  assign \new_[2999]_  = \new_[178]_  | \new_[2998]_ ;
  assign \new_[3000]_  = \new_[2999]_  | \new_[2994]_ ;
  assign \new_[3001]_  = \new_[3000]_  | \new_[2991]_ ;
  assign \new_[3002]_  = \new_[3001]_  | \new_[2984]_ ;
  assign \new_[3003]_  = \new_[3002]_  | \new_[2967]_ ;
  assign \new_[3006]_  = \new_[174]_  | \new_[175]_ ;
  assign \new_[3009]_  = \new_[172]_  | \new_[173]_ ;
  assign \new_[3010]_  = \new_[3009]_  | \new_[3006]_ ;
  assign \new_[3013]_  = \new_[170]_  | \new_[171]_ ;
  assign \new_[3016]_  = \new_[168]_  | \new_[169]_ ;
  assign \new_[3017]_  = \new_[3016]_  | \new_[3013]_ ;
  assign \new_[3018]_  = \new_[3017]_  | \new_[3010]_ ;
  assign \new_[3021]_  = \new_[166]_  | \new_[167]_ ;
  assign \new_[3024]_  = \new_[164]_  | \new_[165]_ ;
  assign \new_[3025]_  = \new_[3024]_  | \new_[3021]_ ;
  assign \new_[3028]_  = \new_[162]_  | \new_[163]_ ;
  assign \new_[3032]_  = \new_[159]_  | \new_[160]_ ;
  assign \new_[3033]_  = \new_[161]_  | \new_[3032]_ ;
  assign \new_[3034]_  = \new_[3033]_  | \new_[3028]_ ;
  assign \new_[3035]_  = \new_[3034]_  | \new_[3025]_ ;
  assign \new_[3036]_  = \new_[3035]_  | \new_[3018]_ ;
  assign \new_[3039]_  = \new_[157]_  | \new_[158]_ ;
  assign \new_[3042]_  = \new_[155]_  | \new_[156]_ ;
  assign \new_[3043]_  = \new_[3042]_  | \new_[3039]_ ;
  assign \new_[3046]_  = \new_[153]_  | \new_[154]_ ;
  assign \new_[3050]_  = \new_[150]_  | \new_[151]_ ;
  assign \new_[3051]_  = \new_[152]_  | \new_[3050]_ ;
  assign \new_[3052]_  = \new_[3051]_  | \new_[3046]_ ;
  assign \new_[3053]_  = \new_[3052]_  | \new_[3043]_ ;
  assign \new_[3056]_  = \new_[148]_  | \new_[149]_ ;
  assign \new_[3059]_  = \new_[146]_  | \new_[147]_ ;
  assign \new_[3060]_  = \new_[3059]_  | \new_[3056]_ ;
  assign \new_[3063]_  = \new_[144]_  | \new_[145]_ ;
  assign \new_[3067]_  = \new_[141]_  | \new_[142]_ ;
  assign \new_[3068]_  = \new_[143]_  | \new_[3067]_ ;
  assign \new_[3069]_  = \new_[3068]_  | \new_[3063]_ ;
  assign \new_[3070]_  = \new_[3069]_  | \new_[3060]_ ;
  assign \new_[3071]_  = \new_[3070]_  | \new_[3053]_ ;
  assign \new_[3072]_  = \new_[3071]_  | \new_[3036]_ ;
  assign \new_[3073]_  = \new_[3072]_  | \new_[3003]_ ;
  assign \new_[3074]_  = \new_[3073]_  | \new_[2934]_ ;
  assign \new_[3077]_  = \new_[139]_  | \new_[140]_ ;
  assign \new_[3080]_  = \new_[137]_  | \new_[138]_ ;
  assign \new_[3081]_  = \new_[3080]_  | \new_[3077]_ ;
  assign \new_[3084]_  = \new_[135]_  | \new_[136]_ ;
  assign \new_[3087]_  = \new_[133]_  | \new_[134]_ ;
  assign \new_[3088]_  = \new_[3087]_  | \new_[3084]_ ;
  assign \new_[3089]_  = \new_[3088]_  | \new_[3081]_ ;
  assign \new_[3092]_  = \new_[131]_  | \new_[132]_ ;
  assign \new_[3095]_  = \new_[129]_  | \new_[130]_ ;
  assign \new_[3096]_  = \new_[3095]_  | \new_[3092]_ ;
  assign \new_[3099]_  = \new_[127]_  | \new_[128]_ ;
  assign \new_[3103]_  = \new_[124]_  | \new_[125]_ ;
  assign \new_[3104]_  = \new_[126]_  | \new_[3103]_ ;
  assign \new_[3105]_  = \new_[3104]_  | \new_[3099]_ ;
  assign \new_[3106]_  = \new_[3105]_  | \new_[3096]_ ;
  assign \new_[3107]_  = \new_[3106]_  | \new_[3089]_ ;
  assign \new_[3110]_  = \new_[122]_  | \new_[123]_ ;
  assign \new_[3113]_  = \new_[120]_  | \new_[121]_ ;
  assign \new_[3114]_  = \new_[3113]_  | \new_[3110]_ ;
  assign \new_[3117]_  = \new_[118]_  | \new_[119]_ ;
  assign \new_[3121]_  = \new_[115]_  | \new_[116]_ ;
  assign \new_[3122]_  = \new_[117]_  | \new_[3121]_ ;
  assign \new_[3123]_  = \new_[3122]_  | \new_[3117]_ ;
  assign \new_[3124]_  = \new_[3123]_  | \new_[3114]_ ;
  assign \new_[3127]_  = \new_[113]_  | \new_[114]_ ;
  assign \new_[3130]_  = \new_[111]_  | \new_[112]_ ;
  assign \new_[3131]_  = \new_[3130]_  | \new_[3127]_ ;
  assign \new_[3134]_  = \new_[109]_  | \new_[110]_ ;
  assign \new_[3138]_  = \new_[106]_  | \new_[107]_ ;
  assign \new_[3139]_  = \new_[108]_  | \new_[3138]_ ;
  assign \new_[3140]_  = \new_[3139]_  | \new_[3134]_ ;
  assign \new_[3141]_  = \new_[3140]_  | \new_[3131]_ ;
  assign \new_[3142]_  = \new_[3141]_  | \new_[3124]_ ;
  assign \new_[3143]_  = \new_[3142]_  | \new_[3107]_ ;
  assign \new_[3146]_  = \new_[104]_  | \new_[105]_ ;
  assign \new_[3149]_  = \new_[102]_  | \new_[103]_ ;
  assign \new_[3150]_  = \new_[3149]_  | \new_[3146]_ ;
  assign \new_[3153]_  = \new_[100]_  | \new_[101]_ ;
  assign \new_[3156]_  = \new_[98]_  | \new_[99]_ ;
  assign \new_[3157]_  = \new_[3156]_  | \new_[3153]_ ;
  assign \new_[3158]_  = \new_[3157]_  | \new_[3150]_ ;
  assign \new_[3161]_  = \new_[96]_  | \new_[97]_ ;
  assign \new_[3164]_  = \new_[94]_  | \new_[95]_ ;
  assign \new_[3165]_  = \new_[3164]_  | \new_[3161]_ ;
  assign \new_[3168]_  = \new_[92]_  | \new_[93]_ ;
  assign \new_[3172]_  = \new_[89]_  | \new_[90]_ ;
  assign \new_[3173]_  = \new_[91]_  | \new_[3172]_ ;
  assign \new_[3174]_  = \new_[3173]_  | \new_[3168]_ ;
  assign \new_[3175]_  = \new_[3174]_  | \new_[3165]_ ;
  assign \new_[3176]_  = \new_[3175]_  | \new_[3158]_ ;
  assign \new_[3179]_  = \new_[87]_  | \new_[88]_ ;
  assign \new_[3182]_  = \new_[85]_  | \new_[86]_ ;
  assign \new_[3183]_  = \new_[3182]_  | \new_[3179]_ ;
  assign \new_[3186]_  = \new_[83]_  | \new_[84]_ ;
  assign \new_[3190]_  = \new_[80]_  | \new_[81]_ ;
  assign \new_[3191]_  = \new_[82]_  | \new_[3190]_ ;
  assign \new_[3192]_  = \new_[3191]_  | \new_[3186]_ ;
  assign \new_[3193]_  = \new_[3192]_  | \new_[3183]_ ;
  assign \new_[3196]_  = \new_[78]_  | \new_[79]_ ;
  assign \new_[3199]_  = \new_[76]_  | \new_[77]_ ;
  assign \new_[3200]_  = \new_[3199]_  | \new_[3196]_ ;
  assign \new_[3203]_  = \new_[74]_  | \new_[75]_ ;
  assign \new_[3207]_  = \new_[71]_  | \new_[72]_ ;
  assign \new_[3208]_  = \new_[73]_  | \new_[3207]_ ;
  assign \new_[3209]_  = \new_[3208]_  | \new_[3203]_ ;
  assign \new_[3210]_  = \new_[3209]_  | \new_[3200]_ ;
  assign \new_[3211]_  = \new_[3210]_  | \new_[3193]_ ;
  assign \new_[3212]_  = \new_[3211]_  | \new_[3176]_ ;
  assign \new_[3213]_  = \new_[3212]_  | \new_[3143]_ ;
  assign \new_[3216]_  = \new_[69]_  | \new_[70]_ ;
  assign \new_[3219]_  = \new_[67]_  | \new_[68]_ ;
  assign \new_[3220]_  = \new_[3219]_  | \new_[3216]_ ;
  assign \new_[3223]_  = \new_[65]_  | \new_[66]_ ;
  assign \new_[3226]_  = \new_[63]_  | \new_[64]_ ;
  assign \new_[3227]_  = \new_[3226]_  | \new_[3223]_ ;
  assign \new_[3228]_  = \new_[3227]_  | \new_[3220]_ ;
  assign \new_[3231]_  = \new_[61]_  | \new_[62]_ ;
  assign \new_[3234]_  = \new_[59]_  | \new_[60]_ ;
  assign \new_[3235]_  = \new_[3234]_  | \new_[3231]_ ;
  assign \new_[3238]_  = \new_[57]_  | \new_[58]_ ;
  assign \new_[3242]_  = \new_[54]_  | \new_[55]_ ;
  assign \new_[3243]_  = \new_[56]_  | \new_[3242]_ ;
  assign \new_[3244]_  = \new_[3243]_  | \new_[3238]_ ;
  assign \new_[3245]_  = \new_[3244]_  | \new_[3235]_ ;
  assign \new_[3246]_  = \new_[3245]_  | \new_[3228]_ ;
  assign \new_[3249]_  = \new_[52]_  | \new_[53]_ ;
  assign \new_[3252]_  = \new_[50]_  | \new_[51]_ ;
  assign \new_[3253]_  = \new_[3252]_  | \new_[3249]_ ;
  assign \new_[3256]_  = \new_[48]_  | \new_[49]_ ;
  assign \new_[3260]_  = \new_[45]_  | \new_[46]_ ;
  assign \new_[3261]_  = \new_[47]_  | \new_[3260]_ ;
  assign \new_[3262]_  = \new_[3261]_  | \new_[3256]_ ;
  assign \new_[3263]_  = \new_[3262]_  | \new_[3253]_ ;
  assign \new_[3266]_  = \new_[43]_  | \new_[44]_ ;
  assign \new_[3269]_  = \new_[41]_  | \new_[42]_ ;
  assign \new_[3270]_  = \new_[3269]_  | \new_[3266]_ ;
  assign \new_[3273]_  = \new_[39]_  | \new_[40]_ ;
  assign \new_[3277]_  = \new_[36]_  | \new_[37]_ ;
  assign \new_[3278]_  = \new_[38]_  | \new_[3277]_ ;
  assign \new_[3279]_  = \new_[3278]_  | \new_[3273]_ ;
  assign \new_[3280]_  = \new_[3279]_  | \new_[3270]_ ;
  assign \new_[3281]_  = \new_[3280]_  | \new_[3263]_ ;
  assign \new_[3282]_  = \new_[3281]_  | \new_[3246]_ ;
  assign \new_[3285]_  = \new_[34]_  | \new_[35]_ ;
  assign \new_[3288]_  = \new_[32]_  | \new_[33]_ ;
  assign \new_[3289]_  = \new_[3288]_  | \new_[3285]_ ;
  assign \new_[3292]_  = \new_[30]_  | \new_[31]_ ;
  assign \new_[3295]_  = \new_[28]_  | \new_[29]_ ;
  assign \new_[3296]_  = \new_[3295]_  | \new_[3292]_ ;
  assign \new_[3297]_  = \new_[3296]_  | \new_[3289]_ ;
  assign \new_[3300]_  = \new_[26]_  | \new_[27]_ ;
  assign \new_[3303]_  = \new_[24]_  | \new_[25]_ ;
  assign \new_[3304]_  = \new_[3303]_  | \new_[3300]_ ;
  assign \new_[3307]_  = \new_[22]_  | \new_[23]_ ;
  assign \new_[3311]_  = \new_[19]_  | \new_[20]_ ;
  assign \new_[3312]_  = \new_[21]_  | \new_[3311]_ ;
  assign \new_[3313]_  = \new_[3312]_  | \new_[3307]_ ;
  assign \new_[3314]_  = \new_[3313]_  | \new_[3304]_ ;
  assign \new_[3315]_  = \new_[3314]_  | \new_[3297]_ ;
  assign \new_[3318]_  = \new_[17]_  | \new_[18]_ ;
  assign \new_[3321]_  = \new_[15]_  | \new_[16]_ ;
  assign \new_[3322]_  = \new_[3321]_  | \new_[3318]_ ;
  assign \new_[3325]_  = \new_[13]_  | \new_[14]_ ;
  assign \new_[3329]_  = \new_[10]_  | \new_[11]_ ;
  assign \new_[3330]_  = \new_[12]_  | \new_[3329]_ ;
  assign \new_[3331]_  = \new_[3330]_  | \new_[3325]_ ;
  assign \new_[3332]_  = \new_[3331]_  | \new_[3322]_ ;
  assign \new_[3335]_  = \new_[8]_  | \new_[9]_ ;
  assign \new_[3338]_  = \new_[6]_  | \new_[7]_ ;
  assign \new_[3339]_  = \new_[3338]_  | \new_[3335]_ ;
  assign \new_[3342]_  = \new_[4]_  | \new_[5]_ ;
  assign \new_[3346]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[3347]_  = \new_[3]_  | \new_[3346]_ ;
  assign \new_[3348]_  = \new_[3347]_  | \new_[3342]_ ;
  assign \new_[3349]_  = \new_[3348]_  | \new_[3339]_ ;
  assign \new_[3350]_  = \new_[3349]_  | \new_[3332]_ ;
  assign \new_[3351]_  = \new_[3350]_  | \new_[3315]_ ;
  assign \new_[3352]_  = \new_[3351]_  | \new_[3282]_ ;
  assign \new_[3353]_  = \new_[3352]_  | \new_[3213]_ ;
  assign \new_[3354]_  = \new_[3353]_  | \new_[3074]_ ;
  assign \new_[3355]_  = \new_[3354]_  | \new_[2795]_ ;
  assign \new_[3358]_  = A200 & ~A199;
  assign \new_[3361]_  = A233 & ~A232;
  assign \new_[3364]_  = A166 & A168;
  assign \new_[3367]_  = A233 & ~A232;
  assign \new_[3370]_  = A167 & A168;
  assign \new_[3373]_  = A233 & ~A232;
  assign \new_[3377]_  = A232 & A200;
  assign \new_[3378]_  = ~A199 & \new_[3377]_ ;
  assign \new_[3382]_  = A235 & A234;
  assign \new_[3383]_  = ~A233 & \new_[3382]_ ;
  assign \new_[3387]_  = A232 & A200;
  assign \new_[3388]_  = ~A199 & \new_[3387]_ ;
  assign \new_[3392]_  = A236 & A234;
  assign \new_[3393]_  = ~A233 & \new_[3392]_ ;
  assign \new_[3397]_  = A201 & ~A200;
  assign \new_[3398]_  = A199 & \new_[3397]_ ;
  assign \new_[3402]_  = A233 & ~A232;
  assign \new_[3403]_  = A202 & \new_[3402]_ ;
  assign \new_[3407]_  = A201 & ~A200;
  assign \new_[3408]_  = A199 & \new_[3407]_ ;
  assign \new_[3412]_  = A233 & ~A232;
  assign \new_[3413]_  = A203 & \new_[3412]_ ;
  assign \new_[3417]_  = A232 & A166;
  assign \new_[3418]_  = A168 & \new_[3417]_ ;
  assign \new_[3422]_  = A235 & A234;
  assign \new_[3423]_  = ~A233 & \new_[3422]_ ;
  assign \new_[3427]_  = A232 & A166;
  assign \new_[3428]_  = A168 & \new_[3427]_ ;
  assign \new_[3432]_  = A236 & A234;
  assign \new_[3433]_  = ~A233 & \new_[3432]_ ;
  assign \new_[3437]_  = A232 & A167;
  assign \new_[3438]_  = A168 & \new_[3437]_ ;
  assign \new_[3442]_  = A235 & A234;
  assign \new_[3443]_  = ~A233 & \new_[3442]_ ;
  assign \new_[3447]_  = A232 & A167;
  assign \new_[3448]_  = A168 & \new_[3447]_ ;
  assign \new_[3452]_  = A236 & A234;
  assign \new_[3453]_  = ~A233 & \new_[3452]_ ;
  assign \new_[3457]_  = A167 & A169;
  assign \new_[3458]_  = ~A170 & \new_[3457]_ ;
  assign \new_[3462]_  = A233 & ~A232;
  assign \new_[3463]_  = A166 & \new_[3462]_ ;
  assign \new_[3467]_  = ~A167 & A169;
  assign \new_[3468]_  = ~A170 & \new_[3467]_ ;
  assign \new_[3472]_  = A233 & ~A232;
  assign \new_[3473]_  = ~A166 & \new_[3472]_ ;
  assign \new_[3477]_  = A167 & ~A169;
  assign \new_[3478]_  = A170 & \new_[3477]_ ;
  assign \new_[3482]_  = A233 & ~A232;
  assign \new_[3483]_  = ~A166 & \new_[3482]_ ;
  assign \new_[3487]_  = ~A167 & ~A169;
  assign \new_[3488]_  = A170 & \new_[3487]_ ;
  assign \new_[3492]_  = A233 & ~A232;
  assign \new_[3493]_  = A166 & \new_[3492]_ ;
  assign \new_[3496]_  = ~A200 & A199;
  assign \new_[3499]_  = A202 & A201;
  assign \new_[3500]_  = \new_[3499]_  & \new_[3496]_ ;
  assign \new_[3503]_  = ~A233 & A232;
  assign \new_[3506]_  = A235 & A234;
  assign \new_[3507]_  = \new_[3506]_  & \new_[3503]_ ;
  assign \new_[3510]_  = ~A200 & A199;
  assign \new_[3513]_  = A202 & A201;
  assign \new_[3514]_  = \new_[3513]_  & \new_[3510]_ ;
  assign \new_[3517]_  = ~A233 & A232;
  assign \new_[3520]_  = A236 & A234;
  assign \new_[3521]_  = \new_[3520]_  & \new_[3517]_ ;
  assign \new_[3524]_  = ~A200 & A199;
  assign \new_[3527]_  = A203 & A201;
  assign \new_[3528]_  = \new_[3527]_  & \new_[3524]_ ;
  assign \new_[3531]_  = ~A233 & A232;
  assign \new_[3534]_  = A235 & A234;
  assign \new_[3535]_  = \new_[3534]_  & \new_[3531]_ ;
  assign \new_[3538]_  = ~A200 & A199;
  assign \new_[3541]_  = A203 & A201;
  assign \new_[3542]_  = \new_[3541]_  & \new_[3538]_ ;
  assign \new_[3545]_  = ~A233 & A232;
  assign \new_[3548]_  = A236 & A234;
  assign \new_[3549]_  = \new_[3548]_  & \new_[3545]_ ;
  assign \new_[3552]_  = A166 & A168;
  assign \new_[3555]_  = A200 & A199;
  assign \new_[3556]_  = \new_[3555]_  & \new_[3552]_ ;
  assign \new_[3559]_  = A266 & A265;
  assign \new_[3562]_  = A299 & ~A298;
  assign \new_[3563]_  = \new_[3562]_  & \new_[3559]_ ;
  assign \new_[3566]_  = A166 & A168;
  assign \new_[3569]_  = A200 & A199;
  assign \new_[3570]_  = \new_[3569]_  & \new_[3566]_ ;
  assign \new_[3573]_  = ~A267 & ~A266;
  assign \new_[3576]_  = A299 & ~A298;
  assign \new_[3577]_  = \new_[3576]_  & \new_[3573]_ ;
  assign \new_[3580]_  = A166 & A168;
  assign \new_[3583]_  = A200 & A199;
  assign \new_[3584]_  = \new_[3583]_  & \new_[3580]_ ;
  assign \new_[3587]_  = ~A266 & ~A265;
  assign \new_[3590]_  = A299 & ~A298;
  assign \new_[3591]_  = \new_[3590]_  & \new_[3587]_ ;
  assign \new_[3594]_  = A166 & A168;
  assign \new_[3597]_  = A200 & ~A199;
  assign \new_[3598]_  = \new_[3597]_  & \new_[3594]_ ;
  assign \new_[3601]_  = A266 & ~A265;
  assign \new_[3604]_  = ~A300 & A298;
  assign \new_[3605]_  = \new_[3604]_  & \new_[3601]_ ;
  assign \new_[3608]_  = A166 & A168;
  assign \new_[3611]_  = A200 & ~A199;
  assign \new_[3612]_  = \new_[3611]_  & \new_[3608]_ ;
  assign \new_[3615]_  = A266 & ~A265;
  assign \new_[3618]_  = A299 & A298;
  assign \new_[3619]_  = \new_[3618]_  & \new_[3615]_ ;
  assign \new_[3622]_  = A166 & A168;
  assign \new_[3625]_  = A200 & ~A199;
  assign \new_[3626]_  = \new_[3625]_  & \new_[3622]_ ;
  assign \new_[3629]_  = A266 & ~A265;
  assign \new_[3632]_  = ~A299 & ~A298;
  assign \new_[3633]_  = \new_[3632]_  & \new_[3629]_ ;
  assign \new_[3636]_  = A166 & A168;
  assign \new_[3639]_  = ~A201 & ~A200;
  assign \new_[3640]_  = \new_[3639]_  & \new_[3636]_ ;
  assign \new_[3643]_  = A266 & A265;
  assign \new_[3646]_  = A299 & ~A298;
  assign \new_[3647]_  = \new_[3646]_  & \new_[3643]_ ;
  assign \new_[3650]_  = A166 & A168;
  assign \new_[3653]_  = ~A201 & ~A200;
  assign \new_[3654]_  = \new_[3653]_  & \new_[3650]_ ;
  assign \new_[3657]_  = ~A267 & ~A266;
  assign \new_[3660]_  = A299 & ~A298;
  assign \new_[3661]_  = \new_[3660]_  & \new_[3657]_ ;
  assign \new_[3664]_  = A166 & A168;
  assign \new_[3667]_  = ~A201 & ~A200;
  assign \new_[3668]_  = \new_[3667]_  & \new_[3664]_ ;
  assign \new_[3671]_  = ~A266 & ~A265;
  assign \new_[3674]_  = A299 & ~A298;
  assign \new_[3675]_  = \new_[3674]_  & \new_[3671]_ ;
  assign \new_[3678]_  = A166 & A168;
  assign \new_[3681]_  = ~A200 & ~A199;
  assign \new_[3682]_  = \new_[3681]_  & \new_[3678]_ ;
  assign \new_[3685]_  = A266 & A265;
  assign \new_[3688]_  = A299 & ~A298;
  assign \new_[3689]_  = \new_[3688]_  & \new_[3685]_ ;
  assign \new_[3692]_  = A166 & A168;
  assign \new_[3695]_  = ~A200 & ~A199;
  assign \new_[3696]_  = \new_[3695]_  & \new_[3692]_ ;
  assign \new_[3699]_  = ~A267 & ~A266;
  assign \new_[3702]_  = A299 & ~A298;
  assign \new_[3703]_  = \new_[3702]_  & \new_[3699]_ ;
  assign \new_[3706]_  = A166 & A168;
  assign \new_[3709]_  = ~A200 & ~A199;
  assign \new_[3710]_  = \new_[3709]_  & \new_[3706]_ ;
  assign \new_[3713]_  = ~A266 & ~A265;
  assign \new_[3716]_  = A299 & ~A298;
  assign \new_[3717]_  = \new_[3716]_  & \new_[3713]_ ;
  assign \new_[3720]_  = A167 & A168;
  assign \new_[3723]_  = A200 & A199;
  assign \new_[3724]_  = \new_[3723]_  & \new_[3720]_ ;
  assign \new_[3727]_  = A266 & A265;
  assign \new_[3730]_  = A299 & ~A298;
  assign \new_[3731]_  = \new_[3730]_  & \new_[3727]_ ;
  assign \new_[3734]_  = A167 & A168;
  assign \new_[3737]_  = A200 & A199;
  assign \new_[3738]_  = \new_[3737]_  & \new_[3734]_ ;
  assign \new_[3741]_  = ~A267 & ~A266;
  assign \new_[3744]_  = A299 & ~A298;
  assign \new_[3745]_  = \new_[3744]_  & \new_[3741]_ ;
  assign \new_[3748]_  = A167 & A168;
  assign \new_[3751]_  = A200 & A199;
  assign \new_[3752]_  = \new_[3751]_  & \new_[3748]_ ;
  assign \new_[3755]_  = ~A266 & ~A265;
  assign \new_[3758]_  = A299 & ~A298;
  assign \new_[3759]_  = \new_[3758]_  & \new_[3755]_ ;
  assign \new_[3762]_  = A167 & A168;
  assign \new_[3765]_  = A200 & ~A199;
  assign \new_[3766]_  = \new_[3765]_  & \new_[3762]_ ;
  assign \new_[3769]_  = A266 & ~A265;
  assign \new_[3772]_  = ~A300 & A298;
  assign \new_[3773]_  = \new_[3772]_  & \new_[3769]_ ;
  assign \new_[3776]_  = A167 & A168;
  assign \new_[3779]_  = A200 & ~A199;
  assign \new_[3780]_  = \new_[3779]_  & \new_[3776]_ ;
  assign \new_[3783]_  = A266 & ~A265;
  assign \new_[3786]_  = A299 & A298;
  assign \new_[3787]_  = \new_[3786]_  & \new_[3783]_ ;
  assign \new_[3790]_  = A167 & A168;
  assign \new_[3793]_  = A200 & ~A199;
  assign \new_[3794]_  = \new_[3793]_  & \new_[3790]_ ;
  assign \new_[3797]_  = A266 & ~A265;
  assign \new_[3800]_  = ~A299 & ~A298;
  assign \new_[3801]_  = \new_[3800]_  & \new_[3797]_ ;
  assign \new_[3804]_  = A167 & A168;
  assign \new_[3807]_  = ~A201 & ~A200;
  assign \new_[3808]_  = \new_[3807]_  & \new_[3804]_ ;
  assign \new_[3811]_  = A266 & A265;
  assign \new_[3814]_  = A299 & ~A298;
  assign \new_[3815]_  = \new_[3814]_  & \new_[3811]_ ;
  assign \new_[3818]_  = A167 & A168;
  assign \new_[3821]_  = ~A201 & ~A200;
  assign \new_[3822]_  = \new_[3821]_  & \new_[3818]_ ;
  assign \new_[3825]_  = ~A267 & ~A266;
  assign \new_[3828]_  = A299 & ~A298;
  assign \new_[3829]_  = \new_[3828]_  & \new_[3825]_ ;
  assign \new_[3832]_  = A167 & A168;
  assign \new_[3835]_  = ~A201 & ~A200;
  assign \new_[3836]_  = \new_[3835]_  & \new_[3832]_ ;
  assign \new_[3839]_  = ~A266 & ~A265;
  assign \new_[3842]_  = A299 & ~A298;
  assign \new_[3843]_  = \new_[3842]_  & \new_[3839]_ ;
  assign \new_[3846]_  = A167 & A168;
  assign \new_[3849]_  = ~A200 & ~A199;
  assign \new_[3850]_  = \new_[3849]_  & \new_[3846]_ ;
  assign \new_[3853]_  = A266 & A265;
  assign \new_[3856]_  = A299 & ~A298;
  assign \new_[3857]_  = \new_[3856]_  & \new_[3853]_ ;
  assign \new_[3860]_  = A167 & A168;
  assign \new_[3863]_  = ~A200 & ~A199;
  assign \new_[3864]_  = \new_[3863]_  & \new_[3860]_ ;
  assign \new_[3867]_  = ~A267 & ~A266;
  assign \new_[3870]_  = A299 & ~A298;
  assign \new_[3871]_  = \new_[3870]_  & \new_[3867]_ ;
  assign \new_[3874]_  = A167 & A168;
  assign \new_[3877]_  = ~A200 & ~A199;
  assign \new_[3878]_  = \new_[3877]_  & \new_[3874]_ ;
  assign \new_[3881]_  = ~A266 & ~A265;
  assign \new_[3884]_  = A299 & ~A298;
  assign \new_[3885]_  = \new_[3884]_  & \new_[3881]_ ;
  assign \new_[3888]_  = A169 & ~A170;
  assign \new_[3891]_  = A166 & A167;
  assign \new_[3892]_  = \new_[3891]_  & \new_[3888]_ ;
  assign \new_[3895]_  = ~A233 & A232;
  assign \new_[3898]_  = A235 & A234;
  assign \new_[3899]_  = \new_[3898]_  & \new_[3895]_ ;
  assign \new_[3902]_  = A169 & ~A170;
  assign \new_[3905]_  = A166 & A167;
  assign \new_[3906]_  = \new_[3905]_  & \new_[3902]_ ;
  assign \new_[3909]_  = ~A233 & A232;
  assign \new_[3912]_  = A236 & A234;
  assign \new_[3913]_  = \new_[3912]_  & \new_[3909]_ ;
  assign \new_[3916]_  = A169 & ~A170;
  assign \new_[3919]_  = ~A166 & ~A167;
  assign \new_[3920]_  = \new_[3919]_  & \new_[3916]_ ;
  assign \new_[3923]_  = ~A233 & A232;
  assign \new_[3926]_  = A235 & A234;
  assign \new_[3927]_  = \new_[3926]_  & \new_[3923]_ ;
  assign \new_[3930]_  = A169 & ~A170;
  assign \new_[3933]_  = ~A166 & ~A167;
  assign \new_[3934]_  = \new_[3933]_  & \new_[3930]_ ;
  assign \new_[3937]_  = ~A233 & A232;
  assign \new_[3940]_  = A236 & A234;
  assign \new_[3941]_  = \new_[3940]_  & \new_[3937]_ ;
  assign \new_[3944]_  = ~A169 & A170;
  assign \new_[3947]_  = ~A166 & A167;
  assign \new_[3948]_  = \new_[3947]_  & \new_[3944]_ ;
  assign \new_[3951]_  = ~A233 & A232;
  assign \new_[3954]_  = A235 & A234;
  assign \new_[3955]_  = \new_[3954]_  & \new_[3951]_ ;
  assign \new_[3958]_  = ~A169 & A170;
  assign \new_[3961]_  = ~A166 & A167;
  assign \new_[3962]_  = \new_[3961]_  & \new_[3958]_ ;
  assign \new_[3965]_  = ~A233 & A232;
  assign \new_[3968]_  = A236 & A234;
  assign \new_[3969]_  = \new_[3968]_  & \new_[3965]_ ;
  assign \new_[3972]_  = ~A169 & A170;
  assign \new_[3975]_  = A166 & ~A167;
  assign \new_[3976]_  = \new_[3975]_  & \new_[3972]_ ;
  assign \new_[3979]_  = ~A233 & A232;
  assign \new_[3982]_  = A235 & A234;
  assign \new_[3983]_  = \new_[3982]_  & \new_[3979]_ ;
  assign \new_[3986]_  = ~A169 & A170;
  assign \new_[3989]_  = A166 & ~A167;
  assign \new_[3990]_  = \new_[3989]_  & \new_[3986]_ ;
  assign \new_[3993]_  = ~A233 & A232;
  assign \new_[3996]_  = A236 & A234;
  assign \new_[3997]_  = \new_[3996]_  & \new_[3993]_ ;
  assign \new_[4000]_  = A166 & A168;
  assign \new_[4003]_  = A200 & A199;
  assign \new_[4004]_  = \new_[4003]_  & \new_[4000]_ ;
  assign \new_[4007]_  = ~A268 & ~A266;
  assign \new_[4011]_  = A299 & ~A298;
  assign \new_[4012]_  = ~A269 & \new_[4011]_ ;
  assign \new_[4013]_  = \new_[4012]_  & \new_[4007]_ ;
  assign \new_[4016]_  = A166 & A168;
  assign \new_[4019]_  = A200 & ~A199;
  assign \new_[4020]_  = \new_[4019]_  & \new_[4016]_ ;
  assign \new_[4023]_  = A266 & ~A265;
  assign \new_[4027]_  = ~A302 & ~A301;
  assign \new_[4028]_  = A298 & \new_[4027]_ ;
  assign \new_[4029]_  = \new_[4028]_  & \new_[4023]_ ;
  assign \new_[4032]_  = A166 & A168;
  assign \new_[4035]_  = ~A202 & ~A200;
  assign \new_[4036]_  = \new_[4035]_  & \new_[4032]_ ;
  assign \new_[4039]_  = A265 & ~A203;
  assign \new_[4043]_  = A299 & ~A298;
  assign \new_[4044]_  = A266 & \new_[4043]_ ;
  assign \new_[4045]_  = \new_[4044]_  & \new_[4039]_ ;
  assign \new_[4048]_  = A166 & A168;
  assign \new_[4051]_  = ~A202 & ~A200;
  assign \new_[4052]_  = \new_[4051]_  & \new_[4048]_ ;
  assign \new_[4055]_  = ~A266 & ~A203;
  assign \new_[4059]_  = A299 & ~A298;
  assign \new_[4060]_  = ~A267 & \new_[4059]_ ;
  assign \new_[4061]_  = \new_[4060]_  & \new_[4055]_ ;
  assign \new_[4064]_  = A166 & A168;
  assign \new_[4067]_  = ~A202 & ~A200;
  assign \new_[4068]_  = \new_[4067]_  & \new_[4064]_ ;
  assign \new_[4071]_  = ~A265 & ~A203;
  assign \new_[4075]_  = A299 & ~A298;
  assign \new_[4076]_  = ~A266 & \new_[4075]_ ;
  assign \new_[4077]_  = \new_[4076]_  & \new_[4071]_ ;
  assign \new_[4080]_  = A166 & A168;
  assign \new_[4083]_  = ~A201 & ~A200;
  assign \new_[4084]_  = \new_[4083]_  & \new_[4080]_ ;
  assign \new_[4087]_  = ~A268 & ~A266;
  assign \new_[4091]_  = A299 & ~A298;
  assign \new_[4092]_  = ~A269 & \new_[4091]_ ;
  assign \new_[4093]_  = \new_[4092]_  & \new_[4087]_ ;
  assign \new_[4096]_  = A166 & A168;
  assign \new_[4099]_  = ~A200 & ~A199;
  assign \new_[4100]_  = \new_[4099]_  & \new_[4096]_ ;
  assign \new_[4103]_  = ~A268 & ~A266;
  assign \new_[4107]_  = A299 & ~A298;
  assign \new_[4108]_  = ~A269 & \new_[4107]_ ;
  assign \new_[4109]_  = \new_[4108]_  & \new_[4103]_ ;
  assign \new_[4112]_  = A167 & A168;
  assign \new_[4115]_  = A200 & A199;
  assign \new_[4116]_  = \new_[4115]_  & \new_[4112]_ ;
  assign \new_[4119]_  = ~A268 & ~A266;
  assign \new_[4123]_  = A299 & ~A298;
  assign \new_[4124]_  = ~A269 & \new_[4123]_ ;
  assign \new_[4125]_  = \new_[4124]_  & \new_[4119]_ ;
  assign \new_[4128]_  = A167 & A168;
  assign \new_[4131]_  = A200 & ~A199;
  assign \new_[4132]_  = \new_[4131]_  & \new_[4128]_ ;
  assign \new_[4135]_  = A266 & ~A265;
  assign \new_[4139]_  = ~A302 & ~A301;
  assign \new_[4140]_  = A298 & \new_[4139]_ ;
  assign \new_[4141]_  = \new_[4140]_  & \new_[4135]_ ;
  assign \new_[4144]_  = A167 & A168;
  assign \new_[4147]_  = ~A202 & ~A200;
  assign \new_[4148]_  = \new_[4147]_  & \new_[4144]_ ;
  assign \new_[4151]_  = A265 & ~A203;
  assign \new_[4155]_  = A299 & ~A298;
  assign \new_[4156]_  = A266 & \new_[4155]_ ;
  assign \new_[4157]_  = \new_[4156]_  & \new_[4151]_ ;
  assign \new_[4160]_  = A167 & A168;
  assign \new_[4163]_  = ~A202 & ~A200;
  assign \new_[4164]_  = \new_[4163]_  & \new_[4160]_ ;
  assign \new_[4167]_  = ~A266 & ~A203;
  assign \new_[4171]_  = A299 & ~A298;
  assign \new_[4172]_  = ~A267 & \new_[4171]_ ;
  assign \new_[4173]_  = \new_[4172]_  & \new_[4167]_ ;
  assign \new_[4176]_  = A167 & A168;
  assign \new_[4179]_  = ~A202 & ~A200;
  assign \new_[4180]_  = \new_[4179]_  & \new_[4176]_ ;
  assign \new_[4183]_  = ~A265 & ~A203;
  assign \new_[4187]_  = A299 & ~A298;
  assign \new_[4188]_  = ~A266 & \new_[4187]_ ;
  assign \new_[4189]_  = \new_[4188]_  & \new_[4183]_ ;
  assign \new_[4192]_  = A167 & A168;
  assign \new_[4195]_  = ~A201 & ~A200;
  assign \new_[4196]_  = \new_[4195]_  & \new_[4192]_ ;
  assign \new_[4199]_  = ~A268 & ~A266;
  assign \new_[4203]_  = A299 & ~A298;
  assign \new_[4204]_  = ~A269 & \new_[4203]_ ;
  assign \new_[4205]_  = \new_[4204]_  & \new_[4199]_ ;
  assign \new_[4208]_  = A167 & A168;
  assign \new_[4211]_  = ~A200 & ~A199;
  assign \new_[4212]_  = \new_[4211]_  & \new_[4208]_ ;
  assign \new_[4215]_  = ~A268 & ~A266;
  assign \new_[4219]_  = A299 & ~A298;
  assign \new_[4220]_  = ~A269 & \new_[4219]_ ;
  assign \new_[4221]_  = \new_[4220]_  & \new_[4215]_ ;
  assign \new_[4224]_  = ~A167 & A170;
  assign \new_[4227]_  = A199 & ~A166;
  assign \new_[4228]_  = \new_[4227]_  & \new_[4224]_ ;
  assign \new_[4231]_  = ~A265 & A200;
  assign \new_[4235]_  = ~A300 & A298;
  assign \new_[4236]_  = A266 & \new_[4235]_ ;
  assign \new_[4237]_  = \new_[4236]_  & \new_[4231]_ ;
  assign \new_[4240]_  = ~A167 & A170;
  assign \new_[4243]_  = A199 & ~A166;
  assign \new_[4244]_  = \new_[4243]_  & \new_[4240]_ ;
  assign \new_[4247]_  = ~A265 & A200;
  assign \new_[4251]_  = A299 & A298;
  assign \new_[4252]_  = A266 & \new_[4251]_ ;
  assign \new_[4253]_  = \new_[4252]_  & \new_[4247]_ ;
  assign \new_[4256]_  = ~A167 & A170;
  assign \new_[4259]_  = A199 & ~A166;
  assign \new_[4260]_  = \new_[4259]_  & \new_[4256]_ ;
  assign \new_[4263]_  = ~A265 & A200;
  assign \new_[4267]_  = ~A299 & ~A298;
  assign \new_[4268]_  = A266 & \new_[4267]_ ;
  assign \new_[4269]_  = \new_[4268]_  & \new_[4263]_ ;
  assign \new_[4272]_  = ~A167 & A170;
  assign \new_[4275]_  = ~A199 & ~A166;
  assign \new_[4276]_  = \new_[4275]_  & \new_[4272]_ ;
  assign \new_[4279]_  = A265 & A200;
  assign \new_[4283]_  = A299 & ~A298;
  assign \new_[4284]_  = A266 & \new_[4283]_ ;
  assign \new_[4285]_  = \new_[4284]_  & \new_[4279]_ ;
  assign \new_[4288]_  = ~A167 & A170;
  assign \new_[4291]_  = ~A199 & ~A166;
  assign \new_[4292]_  = \new_[4291]_  & \new_[4288]_ ;
  assign \new_[4295]_  = ~A266 & A200;
  assign \new_[4299]_  = A299 & ~A298;
  assign \new_[4300]_  = ~A267 & \new_[4299]_ ;
  assign \new_[4301]_  = \new_[4300]_  & \new_[4295]_ ;
  assign \new_[4304]_  = ~A167 & A170;
  assign \new_[4307]_  = ~A199 & ~A166;
  assign \new_[4308]_  = \new_[4307]_  & \new_[4304]_ ;
  assign \new_[4311]_  = ~A265 & A200;
  assign \new_[4315]_  = A299 & ~A298;
  assign \new_[4316]_  = ~A266 & \new_[4315]_ ;
  assign \new_[4317]_  = \new_[4316]_  & \new_[4311]_ ;
  assign \new_[4320]_  = ~A167 & A170;
  assign \new_[4323]_  = ~A200 & ~A166;
  assign \new_[4324]_  = \new_[4323]_  & \new_[4320]_ ;
  assign \new_[4327]_  = ~A265 & ~A201;
  assign \new_[4331]_  = ~A300 & A298;
  assign \new_[4332]_  = A266 & \new_[4331]_ ;
  assign \new_[4333]_  = \new_[4332]_  & \new_[4327]_ ;
  assign \new_[4336]_  = ~A167 & A170;
  assign \new_[4339]_  = ~A200 & ~A166;
  assign \new_[4340]_  = \new_[4339]_  & \new_[4336]_ ;
  assign \new_[4343]_  = ~A265 & ~A201;
  assign \new_[4347]_  = A299 & A298;
  assign \new_[4348]_  = A266 & \new_[4347]_ ;
  assign \new_[4349]_  = \new_[4348]_  & \new_[4343]_ ;
  assign \new_[4352]_  = ~A167 & A170;
  assign \new_[4355]_  = ~A200 & ~A166;
  assign \new_[4356]_  = \new_[4355]_  & \new_[4352]_ ;
  assign \new_[4359]_  = ~A265 & ~A201;
  assign \new_[4363]_  = ~A299 & ~A298;
  assign \new_[4364]_  = A266 & \new_[4363]_ ;
  assign \new_[4365]_  = \new_[4364]_  & \new_[4359]_ ;
  assign \new_[4368]_  = ~A167 & A170;
  assign \new_[4371]_  = ~A199 & ~A166;
  assign \new_[4372]_  = \new_[4371]_  & \new_[4368]_ ;
  assign \new_[4375]_  = ~A265 & ~A200;
  assign \new_[4379]_  = ~A300 & A298;
  assign \new_[4380]_  = A266 & \new_[4379]_ ;
  assign \new_[4381]_  = \new_[4380]_  & \new_[4375]_ ;
  assign \new_[4384]_  = ~A167 & A170;
  assign \new_[4387]_  = ~A199 & ~A166;
  assign \new_[4388]_  = \new_[4387]_  & \new_[4384]_ ;
  assign \new_[4391]_  = ~A265 & ~A200;
  assign \new_[4395]_  = A299 & A298;
  assign \new_[4396]_  = A266 & \new_[4395]_ ;
  assign \new_[4397]_  = \new_[4396]_  & \new_[4391]_ ;
  assign \new_[4400]_  = ~A167 & A170;
  assign \new_[4403]_  = ~A199 & ~A166;
  assign \new_[4404]_  = \new_[4403]_  & \new_[4400]_ ;
  assign \new_[4407]_  = ~A265 & ~A200;
  assign \new_[4411]_  = ~A299 & ~A298;
  assign \new_[4412]_  = A266 & \new_[4411]_ ;
  assign \new_[4413]_  = \new_[4412]_  & \new_[4407]_ ;
  assign \new_[4416]_  = A169 & A170;
  assign \new_[4419]_  = A199 & ~A168;
  assign \new_[4420]_  = \new_[4419]_  & \new_[4416]_ ;
  assign \new_[4423]_  = ~A265 & A200;
  assign \new_[4427]_  = ~A300 & A298;
  assign \new_[4428]_  = A266 & \new_[4427]_ ;
  assign \new_[4429]_  = \new_[4428]_  & \new_[4423]_ ;
  assign \new_[4432]_  = A169 & A170;
  assign \new_[4435]_  = A199 & ~A168;
  assign \new_[4436]_  = \new_[4435]_  & \new_[4432]_ ;
  assign \new_[4439]_  = ~A265 & A200;
  assign \new_[4443]_  = A299 & A298;
  assign \new_[4444]_  = A266 & \new_[4443]_ ;
  assign \new_[4445]_  = \new_[4444]_  & \new_[4439]_ ;
  assign \new_[4448]_  = A169 & A170;
  assign \new_[4451]_  = A199 & ~A168;
  assign \new_[4452]_  = \new_[4451]_  & \new_[4448]_ ;
  assign \new_[4455]_  = ~A265 & A200;
  assign \new_[4459]_  = ~A299 & ~A298;
  assign \new_[4460]_  = A266 & \new_[4459]_ ;
  assign \new_[4461]_  = \new_[4460]_  & \new_[4455]_ ;
  assign \new_[4464]_  = A169 & A170;
  assign \new_[4467]_  = ~A199 & ~A168;
  assign \new_[4468]_  = \new_[4467]_  & \new_[4464]_ ;
  assign \new_[4471]_  = A265 & A200;
  assign \new_[4475]_  = A299 & ~A298;
  assign \new_[4476]_  = A266 & \new_[4475]_ ;
  assign \new_[4477]_  = \new_[4476]_  & \new_[4471]_ ;
  assign \new_[4480]_  = A169 & A170;
  assign \new_[4483]_  = ~A199 & ~A168;
  assign \new_[4484]_  = \new_[4483]_  & \new_[4480]_ ;
  assign \new_[4487]_  = ~A266 & A200;
  assign \new_[4491]_  = A299 & ~A298;
  assign \new_[4492]_  = ~A267 & \new_[4491]_ ;
  assign \new_[4493]_  = \new_[4492]_  & \new_[4487]_ ;
  assign \new_[4496]_  = A169 & A170;
  assign \new_[4499]_  = ~A199 & ~A168;
  assign \new_[4500]_  = \new_[4499]_  & \new_[4496]_ ;
  assign \new_[4503]_  = ~A265 & A200;
  assign \new_[4507]_  = A299 & ~A298;
  assign \new_[4508]_  = ~A266 & \new_[4507]_ ;
  assign \new_[4509]_  = \new_[4508]_  & \new_[4503]_ ;
  assign \new_[4512]_  = A169 & A170;
  assign \new_[4515]_  = ~A200 & ~A168;
  assign \new_[4516]_  = \new_[4515]_  & \new_[4512]_ ;
  assign \new_[4519]_  = ~A265 & ~A201;
  assign \new_[4523]_  = ~A300 & A298;
  assign \new_[4524]_  = A266 & \new_[4523]_ ;
  assign \new_[4525]_  = \new_[4524]_  & \new_[4519]_ ;
  assign \new_[4528]_  = A169 & A170;
  assign \new_[4531]_  = ~A200 & ~A168;
  assign \new_[4532]_  = \new_[4531]_  & \new_[4528]_ ;
  assign \new_[4535]_  = ~A265 & ~A201;
  assign \new_[4539]_  = A299 & A298;
  assign \new_[4540]_  = A266 & \new_[4539]_ ;
  assign \new_[4541]_  = \new_[4540]_  & \new_[4535]_ ;
  assign \new_[4544]_  = A169 & A170;
  assign \new_[4547]_  = ~A200 & ~A168;
  assign \new_[4548]_  = \new_[4547]_  & \new_[4544]_ ;
  assign \new_[4551]_  = ~A265 & ~A201;
  assign \new_[4555]_  = ~A299 & ~A298;
  assign \new_[4556]_  = A266 & \new_[4555]_ ;
  assign \new_[4557]_  = \new_[4556]_  & \new_[4551]_ ;
  assign \new_[4560]_  = A169 & A170;
  assign \new_[4563]_  = ~A199 & ~A168;
  assign \new_[4564]_  = \new_[4563]_  & \new_[4560]_ ;
  assign \new_[4567]_  = ~A265 & ~A200;
  assign \new_[4571]_  = ~A300 & A298;
  assign \new_[4572]_  = A266 & \new_[4571]_ ;
  assign \new_[4573]_  = \new_[4572]_  & \new_[4567]_ ;
  assign \new_[4576]_  = A169 & A170;
  assign \new_[4579]_  = ~A199 & ~A168;
  assign \new_[4580]_  = \new_[4579]_  & \new_[4576]_ ;
  assign \new_[4583]_  = ~A265 & ~A200;
  assign \new_[4587]_  = A299 & A298;
  assign \new_[4588]_  = A266 & \new_[4587]_ ;
  assign \new_[4589]_  = \new_[4588]_  & \new_[4583]_ ;
  assign \new_[4592]_  = A169 & A170;
  assign \new_[4595]_  = ~A199 & ~A168;
  assign \new_[4596]_  = \new_[4595]_  & \new_[4592]_ ;
  assign \new_[4599]_  = ~A265 & ~A200;
  assign \new_[4603]_  = ~A299 & ~A298;
  assign \new_[4604]_  = A266 & \new_[4603]_ ;
  assign \new_[4605]_  = \new_[4604]_  & \new_[4599]_ ;
  assign \new_[4608]_  = ~A167 & ~A169;
  assign \new_[4611]_  = A199 & ~A166;
  assign \new_[4612]_  = \new_[4611]_  & \new_[4608]_ ;
  assign \new_[4615]_  = ~A265 & A200;
  assign \new_[4619]_  = ~A300 & A298;
  assign \new_[4620]_  = A266 & \new_[4619]_ ;
  assign \new_[4621]_  = \new_[4620]_  & \new_[4615]_ ;
  assign \new_[4624]_  = ~A167 & ~A169;
  assign \new_[4627]_  = A199 & ~A166;
  assign \new_[4628]_  = \new_[4627]_  & \new_[4624]_ ;
  assign \new_[4631]_  = ~A265 & A200;
  assign \new_[4635]_  = A299 & A298;
  assign \new_[4636]_  = A266 & \new_[4635]_ ;
  assign \new_[4637]_  = \new_[4636]_  & \new_[4631]_ ;
  assign \new_[4640]_  = ~A167 & ~A169;
  assign \new_[4643]_  = A199 & ~A166;
  assign \new_[4644]_  = \new_[4643]_  & \new_[4640]_ ;
  assign \new_[4647]_  = ~A265 & A200;
  assign \new_[4651]_  = ~A299 & ~A298;
  assign \new_[4652]_  = A266 & \new_[4651]_ ;
  assign \new_[4653]_  = \new_[4652]_  & \new_[4647]_ ;
  assign \new_[4656]_  = ~A167 & ~A169;
  assign \new_[4659]_  = ~A199 & ~A166;
  assign \new_[4660]_  = \new_[4659]_  & \new_[4656]_ ;
  assign \new_[4663]_  = A265 & A200;
  assign \new_[4667]_  = A299 & ~A298;
  assign \new_[4668]_  = A266 & \new_[4667]_ ;
  assign \new_[4669]_  = \new_[4668]_  & \new_[4663]_ ;
  assign \new_[4672]_  = ~A167 & ~A169;
  assign \new_[4675]_  = ~A199 & ~A166;
  assign \new_[4676]_  = \new_[4675]_  & \new_[4672]_ ;
  assign \new_[4679]_  = ~A266 & A200;
  assign \new_[4683]_  = A299 & ~A298;
  assign \new_[4684]_  = ~A267 & \new_[4683]_ ;
  assign \new_[4685]_  = \new_[4684]_  & \new_[4679]_ ;
  assign \new_[4688]_  = ~A167 & ~A169;
  assign \new_[4691]_  = ~A199 & ~A166;
  assign \new_[4692]_  = \new_[4691]_  & \new_[4688]_ ;
  assign \new_[4695]_  = ~A265 & A200;
  assign \new_[4699]_  = A299 & ~A298;
  assign \new_[4700]_  = ~A266 & \new_[4699]_ ;
  assign \new_[4701]_  = \new_[4700]_  & \new_[4695]_ ;
  assign \new_[4704]_  = ~A167 & ~A169;
  assign \new_[4707]_  = ~A200 & ~A166;
  assign \new_[4708]_  = \new_[4707]_  & \new_[4704]_ ;
  assign \new_[4711]_  = ~A265 & ~A201;
  assign \new_[4715]_  = ~A300 & A298;
  assign \new_[4716]_  = A266 & \new_[4715]_ ;
  assign \new_[4717]_  = \new_[4716]_  & \new_[4711]_ ;
  assign \new_[4720]_  = ~A167 & ~A169;
  assign \new_[4723]_  = ~A200 & ~A166;
  assign \new_[4724]_  = \new_[4723]_  & \new_[4720]_ ;
  assign \new_[4727]_  = ~A265 & ~A201;
  assign \new_[4731]_  = A299 & A298;
  assign \new_[4732]_  = A266 & \new_[4731]_ ;
  assign \new_[4733]_  = \new_[4732]_  & \new_[4727]_ ;
  assign \new_[4736]_  = ~A167 & ~A169;
  assign \new_[4739]_  = ~A200 & ~A166;
  assign \new_[4740]_  = \new_[4739]_  & \new_[4736]_ ;
  assign \new_[4743]_  = ~A265 & ~A201;
  assign \new_[4747]_  = ~A299 & ~A298;
  assign \new_[4748]_  = A266 & \new_[4747]_ ;
  assign \new_[4749]_  = \new_[4748]_  & \new_[4743]_ ;
  assign \new_[4752]_  = ~A167 & ~A169;
  assign \new_[4755]_  = ~A199 & ~A166;
  assign \new_[4756]_  = \new_[4755]_  & \new_[4752]_ ;
  assign \new_[4759]_  = ~A265 & ~A200;
  assign \new_[4763]_  = ~A300 & A298;
  assign \new_[4764]_  = A266 & \new_[4763]_ ;
  assign \new_[4765]_  = \new_[4764]_  & \new_[4759]_ ;
  assign \new_[4768]_  = ~A167 & ~A169;
  assign \new_[4771]_  = ~A199 & ~A166;
  assign \new_[4772]_  = \new_[4771]_  & \new_[4768]_ ;
  assign \new_[4775]_  = ~A265 & ~A200;
  assign \new_[4779]_  = A299 & A298;
  assign \new_[4780]_  = A266 & \new_[4779]_ ;
  assign \new_[4781]_  = \new_[4780]_  & \new_[4775]_ ;
  assign \new_[4784]_  = ~A167 & ~A169;
  assign \new_[4787]_  = ~A199 & ~A166;
  assign \new_[4788]_  = \new_[4787]_  & \new_[4784]_ ;
  assign \new_[4791]_  = ~A265 & ~A200;
  assign \new_[4795]_  = ~A299 & ~A298;
  assign \new_[4796]_  = A266 & \new_[4795]_ ;
  assign \new_[4797]_  = \new_[4796]_  & \new_[4791]_ ;
  assign \new_[4800]_  = ~A169 & ~A170;
  assign \new_[4803]_  = A199 & ~A168;
  assign \new_[4804]_  = \new_[4803]_  & \new_[4800]_ ;
  assign \new_[4807]_  = ~A265 & A200;
  assign \new_[4811]_  = ~A300 & A298;
  assign \new_[4812]_  = A266 & \new_[4811]_ ;
  assign \new_[4813]_  = \new_[4812]_  & \new_[4807]_ ;
  assign \new_[4816]_  = ~A169 & ~A170;
  assign \new_[4819]_  = A199 & ~A168;
  assign \new_[4820]_  = \new_[4819]_  & \new_[4816]_ ;
  assign \new_[4823]_  = ~A265 & A200;
  assign \new_[4827]_  = A299 & A298;
  assign \new_[4828]_  = A266 & \new_[4827]_ ;
  assign \new_[4829]_  = \new_[4828]_  & \new_[4823]_ ;
  assign \new_[4832]_  = ~A169 & ~A170;
  assign \new_[4835]_  = A199 & ~A168;
  assign \new_[4836]_  = \new_[4835]_  & \new_[4832]_ ;
  assign \new_[4839]_  = ~A265 & A200;
  assign \new_[4843]_  = ~A299 & ~A298;
  assign \new_[4844]_  = A266 & \new_[4843]_ ;
  assign \new_[4845]_  = \new_[4844]_  & \new_[4839]_ ;
  assign \new_[4848]_  = ~A169 & ~A170;
  assign \new_[4851]_  = ~A199 & ~A168;
  assign \new_[4852]_  = \new_[4851]_  & \new_[4848]_ ;
  assign \new_[4855]_  = A265 & A200;
  assign \new_[4859]_  = A299 & ~A298;
  assign \new_[4860]_  = A266 & \new_[4859]_ ;
  assign \new_[4861]_  = \new_[4860]_  & \new_[4855]_ ;
  assign \new_[4864]_  = ~A169 & ~A170;
  assign \new_[4867]_  = ~A199 & ~A168;
  assign \new_[4868]_  = \new_[4867]_  & \new_[4864]_ ;
  assign \new_[4871]_  = ~A266 & A200;
  assign \new_[4875]_  = A299 & ~A298;
  assign \new_[4876]_  = ~A267 & \new_[4875]_ ;
  assign \new_[4877]_  = \new_[4876]_  & \new_[4871]_ ;
  assign \new_[4880]_  = ~A169 & ~A170;
  assign \new_[4883]_  = ~A199 & ~A168;
  assign \new_[4884]_  = \new_[4883]_  & \new_[4880]_ ;
  assign \new_[4887]_  = ~A265 & A200;
  assign \new_[4891]_  = A299 & ~A298;
  assign \new_[4892]_  = ~A266 & \new_[4891]_ ;
  assign \new_[4893]_  = \new_[4892]_  & \new_[4887]_ ;
  assign \new_[4896]_  = ~A169 & ~A170;
  assign \new_[4899]_  = ~A200 & ~A168;
  assign \new_[4900]_  = \new_[4899]_  & \new_[4896]_ ;
  assign \new_[4903]_  = ~A265 & ~A201;
  assign \new_[4907]_  = ~A300 & A298;
  assign \new_[4908]_  = A266 & \new_[4907]_ ;
  assign \new_[4909]_  = \new_[4908]_  & \new_[4903]_ ;
  assign \new_[4912]_  = ~A169 & ~A170;
  assign \new_[4915]_  = ~A200 & ~A168;
  assign \new_[4916]_  = \new_[4915]_  & \new_[4912]_ ;
  assign \new_[4919]_  = ~A265 & ~A201;
  assign \new_[4923]_  = A299 & A298;
  assign \new_[4924]_  = A266 & \new_[4923]_ ;
  assign \new_[4925]_  = \new_[4924]_  & \new_[4919]_ ;
  assign \new_[4928]_  = ~A169 & ~A170;
  assign \new_[4931]_  = ~A200 & ~A168;
  assign \new_[4932]_  = \new_[4931]_  & \new_[4928]_ ;
  assign \new_[4935]_  = ~A265 & ~A201;
  assign \new_[4939]_  = ~A299 & ~A298;
  assign \new_[4940]_  = A266 & \new_[4939]_ ;
  assign \new_[4941]_  = \new_[4940]_  & \new_[4935]_ ;
  assign \new_[4944]_  = ~A169 & ~A170;
  assign \new_[4947]_  = ~A199 & ~A168;
  assign \new_[4948]_  = \new_[4947]_  & \new_[4944]_ ;
  assign \new_[4951]_  = ~A265 & ~A200;
  assign \new_[4955]_  = ~A300 & A298;
  assign \new_[4956]_  = A266 & \new_[4955]_ ;
  assign \new_[4957]_  = \new_[4956]_  & \new_[4951]_ ;
  assign \new_[4960]_  = ~A169 & ~A170;
  assign \new_[4963]_  = ~A199 & ~A168;
  assign \new_[4964]_  = \new_[4963]_  & \new_[4960]_ ;
  assign \new_[4967]_  = ~A265 & ~A200;
  assign \new_[4971]_  = A299 & A298;
  assign \new_[4972]_  = A266 & \new_[4971]_ ;
  assign \new_[4973]_  = \new_[4972]_  & \new_[4967]_ ;
  assign \new_[4976]_  = ~A169 & ~A170;
  assign \new_[4979]_  = ~A199 & ~A168;
  assign \new_[4980]_  = \new_[4979]_  & \new_[4976]_ ;
  assign \new_[4983]_  = ~A265 & ~A200;
  assign \new_[4987]_  = ~A299 & ~A298;
  assign \new_[4988]_  = A266 & \new_[4987]_ ;
  assign \new_[4989]_  = \new_[4988]_  & \new_[4983]_ ;
  assign \new_[4992]_  = A166 & A168;
  assign \new_[4996]_  = A265 & A200;
  assign \new_[4997]_  = A199 & \new_[4996]_ ;
  assign \new_[4998]_  = \new_[4997]_  & \new_[4992]_ ;
  assign \new_[5001]_  = A298 & A266;
  assign \new_[5005]_  = A301 & A300;
  assign \new_[5006]_  = ~A299 & \new_[5005]_ ;
  assign \new_[5007]_  = \new_[5006]_  & \new_[5001]_ ;
  assign \new_[5010]_  = A166 & A168;
  assign \new_[5014]_  = A265 & A200;
  assign \new_[5015]_  = A199 & \new_[5014]_ ;
  assign \new_[5016]_  = \new_[5015]_  & \new_[5010]_ ;
  assign \new_[5019]_  = A298 & A266;
  assign \new_[5023]_  = A302 & A300;
  assign \new_[5024]_  = ~A299 & \new_[5023]_ ;
  assign \new_[5025]_  = \new_[5024]_  & \new_[5019]_ ;
  assign \new_[5028]_  = A166 & A168;
  assign \new_[5032]_  = ~A266 & A200;
  assign \new_[5033]_  = A199 & \new_[5032]_ ;
  assign \new_[5034]_  = \new_[5033]_  & \new_[5028]_ ;
  assign \new_[5037]_  = A298 & ~A267;
  assign \new_[5041]_  = A301 & A300;
  assign \new_[5042]_  = ~A299 & \new_[5041]_ ;
  assign \new_[5043]_  = \new_[5042]_  & \new_[5037]_ ;
  assign \new_[5046]_  = A166 & A168;
  assign \new_[5050]_  = ~A266 & A200;
  assign \new_[5051]_  = A199 & \new_[5050]_ ;
  assign \new_[5052]_  = \new_[5051]_  & \new_[5046]_ ;
  assign \new_[5055]_  = A298 & ~A267;
  assign \new_[5059]_  = A302 & A300;
  assign \new_[5060]_  = ~A299 & \new_[5059]_ ;
  assign \new_[5061]_  = \new_[5060]_  & \new_[5055]_ ;
  assign \new_[5064]_  = A166 & A168;
  assign \new_[5068]_  = ~A265 & A200;
  assign \new_[5069]_  = A199 & \new_[5068]_ ;
  assign \new_[5070]_  = \new_[5069]_  & \new_[5064]_ ;
  assign \new_[5073]_  = A298 & ~A266;
  assign \new_[5077]_  = A301 & A300;
  assign \new_[5078]_  = ~A299 & \new_[5077]_ ;
  assign \new_[5079]_  = \new_[5078]_  & \new_[5073]_ ;
  assign \new_[5082]_  = A166 & A168;
  assign \new_[5086]_  = ~A265 & A200;
  assign \new_[5087]_  = A199 & \new_[5086]_ ;
  assign \new_[5088]_  = \new_[5087]_  & \new_[5082]_ ;
  assign \new_[5091]_  = A298 & ~A266;
  assign \new_[5095]_  = A302 & A300;
  assign \new_[5096]_  = ~A299 & \new_[5095]_ ;
  assign \new_[5097]_  = \new_[5096]_  & \new_[5091]_ ;
  assign \new_[5100]_  = A166 & A168;
  assign \new_[5104]_  = A265 & A200;
  assign \new_[5105]_  = ~A199 & \new_[5104]_ ;
  assign \new_[5106]_  = \new_[5105]_  & \new_[5100]_ ;
  assign \new_[5109]_  = A267 & ~A266;
  assign \new_[5113]_  = ~A300 & A298;
  assign \new_[5114]_  = A268 & \new_[5113]_ ;
  assign \new_[5115]_  = \new_[5114]_  & \new_[5109]_ ;
  assign \new_[5118]_  = A166 & A168;
  assign \new_[5122]_  = A265 & A200;
  assign \new_[5123]_  = ~A199 & \new_[5122]_ ;
  assign \new_[5124]_  = \new_[5123]_  & \new_[5118]_ ;
  assign \new_[5127]_  = A267 & ~A266;
  assign \new_[5131]_  = A299 & A298;
  assign \new_[5132]_  = A268 & \new_[5131]_ ;
  assign \new_[5133]_  = \new_[5132]_  & \new_[5127]_ ;
  assign \new_[5136]_  = A166 & A168;
  assign \new_[5140]_  = A265 & A200;
  assign \new_[5141]_  = ~A199 & \new_[5140]_ ;
  assign \new_[5142]_  = \new_[5141]_  & \new_[5136]_ ;
  assign \new_[5145]_  = A267 & ~A266;
  assign \new_[5149]_  = ~A299 & ~A298;
  assign \new_[5150]_  = A268 & \new_[5149]_ ;
  assign \new_[5151]_  = \new_[5150]_  & \new_[5145]_ ;
  assign \new_[5154]_  = A166 & A168;
  assign \new_[5158]_  = A265 & A200;
  assign \new_[5159]_  = ~A199 & \new_[5158]_ ;
  assign \new_[5160]_  = \new_[5159]_  & \new_[5154]_ ;
  assign \new_[5163]_  = A267 & ~A266;
  assign \new_[5167]_  = ~A300 & A298;
  assign \new_[5168]_  = A269 & \new_[5167]_ ;
  assign \new_[5169]_  = \new_[5168]_  & \new_[5163]_ ;
  assign \new_[5172]_  = A166 & A168;
  assign \new_[5176]_  = A265 & A200;
  assign \new_[5177]_  = ~A199 & \new_[5176]_ ;
  assign \new_[5178]_  = \new_[5177]_  & \new_[5172]_ ;
  assign \new_[5181]_  = A267 & ~A266;
  assign \new_[5185]_  = A299 & A298;
  assign \new_[5186]_  = A269 & \new_[5185]_ ;
  assign \new_[5187]_  = \new_[5186]_  & \new_[5181]_ ;
  assign \new_[5190]_  = A166 & A168;
  assign \new_[5194]_  = A265 & A200;
  assign \new_[5195]_  = ~A199 & \new_[5194]_ ;
  assign \new_[5196]_  = \new_[5195]_  & \new_[5190]_ ;
  assign \new_[5199]_  = A267 & ~A266;
  assign \new_[5203]_  = ~A299 & ~A298;
  assign \new_[5204]_  = A269 & \new_[5203]_ ;
  assign \new_[5205]_  = \new_[5204]_  & \new_[5199]_ ;
  assign \new_[5208]_  = A166 & A168;
  assign \new_[5212]_  = ~A203 & ~A202;
  assign \new_[5213]_  = ~A200 & \new_[5212]_ ;
  assign \new_[5214]_  = \new_[5213]_  & \new_[5208]_ ;
  assign \new_[5217]_  = ~A268 & ~A266;
  assign \new_[5221]_  = A299 & ~A298;
  assign \new_[5222]_  = ~A269 & \new_[5221]_ ;
  assign \new_[5223]_  = \new_[5222]_  & \new_[5217]_ ;
  assign \new_[5226]_  = A166 & A168;
  assign \new_[5230]_  = A265 & ~A201;
  assign \new_[5231]_  = ~A200 & \new_[5230]_ ;
  assign \new_[5232]_  = \new_[5231]_  & \new_[5226]_ ;
  assign \new_[5235]_  = A298 & A266;
  assign \new_[5239]_  = A301 & A300;
  assign \new_[5240]_  = ~A299 & \new_[5239]_ ;
  assign \new_[5241]_  = \new_[5240]_  & \new_[5235]_ ;
  assign \new_[5244]_  = A166 & A168;
  assign \new_[5248]_  = A265 & ~A201;
  assign \new_[5249]_  = ~A200 & \new_[5248]_ ;
  assign \new_[5250]_  = \new_[5249]_  & \new_[5244]_ ;
  assign \new_[5253]_  = A298 & A266;
  assign \new_[5257]_  = A302 & A300;
  assign \new_[5258]_  = ~A299 & \new_[5257]_ ;
  assign \new_[5259]_  = \new_[5258]_  & \new_[5253]_ ;
  assign \new_[5262]_  = A166 & A168;
  assign \new_[5266]_  = ~A266 & ~A201;
  assign \new_[5267]_  = ~A200 & \new_[5266]_ ;
  assign \new_[5268]_  = \new_[5267]_  & \new_[5262]_ ;
  assign \new_[5271]_  = A298 & ~A267;
  assign \new_[5275]_  = A301 & A300;
  assign \new_[5276]_  = ~A299 & \new_[5275]_ ;
  assign \new_[5277]_  = \new_[5276]_  & \new_[5271]_ ;
  assign \new_[5280]_  = A166 & A168;
  assign \new_[5284]_  = ~A266 & ~A201;
  assign \new_[5285]_  = ~A200 & \new_[5284]_ ;
  assign \new_[5286]_  = \new_[5285]_  & \new_[5280]_ ;
  assign \new_[5289]_  = A298 & ~A267;
  assign \new_[5293]_  = A302 & A300;
  assign \new_[5294]_  = ~A299 & \new_[5293]_ ;
  assign \new_[5295]_  = \new_[5294]_  & \new_[5289]_ ;
  assign \new_[5298]_  = A166 & A168;
  assign \new_[5302]_  = ~A265 & ~A201;
  assign \new_[5303]_  = ~A200 & \new_[5302]_ ;
  assign \new_[5304]_  = \new_[5303]_  & \new_[5298]_ ;
  assign \new_[5307]_  = A298 & ~A266;
  assign \new_[5311]_  = A301 & A300;
  assign \new_[5312]_  = ~A299 & \new_[5311]_ ;
  assign \new_[5313]_  = \new_[5312]_  & \new_[5307]_ ;
  assign \new_[5316]_  = A166 & A168;
  assign \new_[5320]_  = ~A265 & ~A201;
  assign \new_[5321]_  = ~A200 & \new_[5320]_ ;
  assign \new_[5322]_  = \new_[5321]_  & \new_[5316]_ ;
  assign \new_[5325]_  = A298 & ~A266;
  assign \new_[5329]_  = A302 & A300;
  assign \new_[5330]_  = ~A299 & \new_[5329]_ ;
  assign \new_[5331]_  = \new_[5330]_  & \new_[5325]_ ;
  assign \new_[5334]_  = A166 & A168;
  assign \new_[5338]_  = A201 & ~A200;
  assign \new_[5339]_  = A199 & \new_[5338]_ ;
  assign \new_[5340]_  = \new_[5339]_  & \new_[5334]_ ;
  assign \new_[5343]_  = ~A265 & A202;
  assign \new_[5347]_  = ~A300 & A298;
  assign \new_[5348]_  = A266 & \new_[5347]_ ;
  assign \new_[5349]_  = \new_[5348]_  & \new_[5343]_ ;
  assign \new_[5352]_  = A166 & A168;
  assign \new_[5356]_  = A201 & ~A200;
  assign \new_[5357]_  = A199 & \new_[5356]_ ;
  assign \new_[5358]_  = \new_[5357]_  & \new_[5352]_ ;
  assign \new_[5361]_  = ~A265 & A202;
  assign \new_[5365]_  = A299 & A298;
  assign \new_[5366]_  = A266 & \new_[5365]_ ;
  assign \new_[5367]_  = \new_[5366]_  & \new_[5361]_ ;
  assign \new_[5370]_  = A166 & A168;
  assign \new_[5374]_  = A201 & ~A200;
  assign \new_[5375]_  = A199 & \new_[5374]_ ;
  assign \new_[5376]_  = \new_[5375]_  & \new_[5370]_ ;
  assign \new_[5379]_  = ~A265 & A202;
  assign \new_[5383]_  = ~A299 & ~A298;
  assign \new_[5384]_  = A266 & \new_[5383]_ ;
  assign \new_[5385]_  = \new_[5384]_  & \new_[5379]_ ;
  assign \new_[5388]_  = A166 & A168;
  assign \new_[5392]_  = A201 & ~A200;
  assign \new_[5393]_  = A199 & \new_[5392]_ ;
  assign \new_[5394]_  = \new_[5393]_  & \new_[5388]_ ;
  assign \new_[5397]_  = ~A265 & A203;
  assign \new_[5401]_  = ~A300 & A298;
  assign \new_[5402]_  = A266 & \new_[5401]_ ;
  assign \new_[5403]_  = \new_[5402]_  & \new_[5397]_ ;
  assign \new_[5406]_  = A166 & A168;
  assign \new_[5410]_  = A201 & ~A200;
  assign \new_[5411]_  = A199 & \new_[5410]_ ;
  assign \new_[5412]_  = \new_[5411]_  & \new_[5406]_ ;
  assign \new_[5415]_  = ~A265 & A203;
  assign \new_[5419]_  = A299 & A298;
  assign \new_[5420]_  = A266 & \new_[5419]_ ;
  assign \new_[5421]_  = \new_[5420]_  & \new_[5415]_ ;
  assign \new_[5424]_  = A166 & A168;
  assign \new_[5428]_  = A201 & ~A200;
  assign \new_[5429]_  = A199 & \new_[5428]_ ;
  assign \new_[5430]_  = \new_[5429]_  & \new_[5424]_ ;
  assign \new_[5433]_  = ~A265 & A203;
  assign \new_[5437]_  = ~A299 & ~A298;
  assign \new_[5438]_  = A266 & \new_[5437]_ ;
  assign \new_[5439]_  = \new_[5438]_  & \new_[5433]_ ;
  assign \new_[5442]_  = A166 & A168;
  assign \new_[5446]_  = A265 & ~A200;
  assign \new_[5447]_  = ~A199 & \new_[5446]_ ;
  assign \new_[5448]_  = \new_[5447]_  & \new_[5442]_ ;
  assign \new_[5451]_  = A298 & A266;
  assign \new_[5455]_  = A301 & A300;
  assign \new_[5456]_  = ~A299 & \new_[5455]_ ;
  assign \new_[5457]_  = \new_[5456]_  & \new_[5451]_ ;
  assign \new_[5460]_  = A166 & A168;
  assign \new_[5464]_  = A265 & ~A200;
  assign \new_[5465]_  = ~A199 & \new_[5464]_ ;
  assign \new_[5466]_  = \new_[5465]_  & \new_[5460]_ ;
  assign \new_[5469]_  = A298 & A266;
  assign \new_[5473]_  = A302 & A300;
  assign \new_[5474]_  = ~A299 & \new_[5473]_ ;
  assign \new_[5475]_  = \new_[5474]_  & \new_[5469]_ ;
  assign \new_[5478]_  = A166 & A168;
  assign \new_[5482]_  = ~A266 & ~A200;
  assign \new_[5483]_  = ~A199 & \new_[5482]_ ;
  assign \new_[5484]_  = \new_[5483]_  & \new_[5478]_ ;
  assign \new_[5487]_  = A298 & ~A267;
  assign \new_[5491]_  = A301 & A300;
  assign \new_[5492]_  = ~A299 & \new_[5491]_ ;
  assign \new_[5493]_  = \new_[5492]_  & \new_[5487]_ ;
  assign \new_[5496]_  = A166 & A168;
  assign \new_[5500]_  = ~A266 & ~A200;
  assign \new_[5501]_  = ~A199 & \new_[5500]_ ;
  assign \new_[5502]_  = \new_[5501]_  & \new_[5496]_ ;
  assign \new_[5505]_  = A298 & ~A267;
  assign \new_[5509]_  = A302 & A300;
  assign \new_[5510]_  = ~A299 & \new_[5509]_ ;
  assign \new_[5511]_  = \new_[5510]_  & \new_[5505]_ ;
  assign \new_[5514]_  = A166 & A168;
  assign \new_[5518]_  = ~A265 & ~A200;
  assign \new_[5519]_  = ~A199 & \new_[5518]_ ;
  assign \new_[5520]_  = \new_[5519]_  & \new_[5514]_ ;
  assign \new_[5523]_  = A298 & ~A266;
  assign \new_[5527]_  = A301 & A300;
  assign \new_[5528]_  = ~A299 & \new_[5527]_ ;
  assign \new_[5529]_  = \new_[5528]_  & \new_[5523]_ ;
  assign \new_[5532]_  = A166 & A168;
  assign \new_[5536]_  = ~A265 & ~A200;
  assign \new_[5537]_  = ~A199 & \new_[5536]_ ;
  assign \new_[5538]_  = \new_[5537]_  & \new_[5532]_ ;
  assign \new_[5541]_  = A298 & ~A266;
  assign \new_[5545]_  = A302 & A300;
  assign \new_[5546]_  = ~A299 & \new_[5545]_ ;
  assign \new_[5547]_  = \new_[5546]_  & \new_[5541]_ ;
  assign \new_[5550]_  = A167 & A168;
  assign \new_[5554]_  = A265 & A200;
  assign \new_[5555]_  = A199 & \new_[5554]_ ;
  assign \new_[5556]_  = \new_[5555]_  & \new_[5550]_ ;
  assign \new_[5559]_  = A298 & A266;
  assign \new_[5563]_  = A301 & A300;
  assign \new_[5564]_  = ~A299 & \new_[5563]_ ;
  assign \new_[5565]_  = \new_[5564]_  & \new_[5559]_ ;
  assign \new_[5568]_  = A167 & A168;
  assign \new_[5572]_  = A265 & A200;
  assign \new_[5573]_  = A199 & \new_[5572]_ ;
  assign \new_[5574]_  = \new_[5573]_  & \new_[5568]_ ;
  assign \new_[5577]_  = A298 & A266;
  assign \new_[5581]_  = A302 & A300;
  assign \new_[5582]_  = ~A299 & \new_[5581]_ ;
  assign \new_[5583]_  = \new_[5582]_  & \new_[5577]_ ;
  assign \new_[5586]_  = A167 & A168;
  assign \new_[5590]_  = ~A266 & A200;
  assign \new_[5591]_  = A199 & \new_[5590]_ ;
  assign \new_[5592]_  = \new_[5591]_  & \new_[5586]_ ;
  assign \new_[5595]_  = A298 & ~A267;
  assign \new_[5599]_  = A301 & A300;
  assign \new_[5600]_  = ~A299 & \new_[5599]_ ;
  assign \new_[5601]_  = \new_[5600]_  & \new_[5595]_ ;
  assign \new_[5604]_  = A167 & A168;
  assign \new_[5608]_  = ~A266 & A200;
  assign \new_[5609]_  = A199 & \new_[5608]_ ;
  assign \new_[5610]_  = \new_[5609]_  & \new_[5604]_ ;
  assign \new_[5613]_  = A298 & ~A267;
  assign \new_[5617]_  = A302 & A300;
  assign \new_[5618]_  = ~A299 & \new_[5617]_ ;
  assign \new_[5619]_  = \new_[5618]_  & \new_[5613]_ ;
  assign \new_[5622]_  = A167 & A168;
  assign \new_[5626]_  = ~A265 & A200;
  assign \new_[5627]_  = A199 & \new_[5626]_ ;
  assign \new_[5628]_  = \new_[5627]_  & \new_[5622]_ ;
  assign \new_[5631]_  = A298 & ~A266;
  assign \new_[5635]_  = A301 & A300;
  assign \new_[5636]_  = ~A299 & \new_[5635]_ ;
  assign \new_[5637]_  = \new_[5636]_  & \new_[5631]_ ;
  assign \new_[5640]_  = A167 & A168;
  assign \new_[5644]_  = ~A265 & A200;
  assign \new_[5645]_  = A199 & \new_[5644]_ ;
  assign \new_[5646]_  = \new_[5645]_  & \new_[5640]_ ;
  assign \new_[5649]_  = A298 & ~A266;
  assign \new_[5653]_  = A302 & A300;
  assign \new_[5654]_  = ~A299 & \new_[5653]_ ;
  assign \new_[5655]_  = \new_[5654]_  & \new_[5649]_ ;
  assign \new_[5658]_  = A167 & A168;
  assign \new_[5662]_  = A265 & A200;
  assign \new_[5663]_  = ~A199 & \new_[5662]_ ;
  assign \new_[5664]_  = \new_[5663]_  & \new_[5658]_ ;
  assign \new_[5667]_  = A267 & ~A266;
  assign \new_[5671]_  = ~A300 & A298;
  assign \new_[5672]_  = A268 & \new_[5671]_ ;
  assign \new_[5673]_  = \new_[5672]_  & \new_[5667]_ ;
  assign \new_[5676]_  = A167 & A168;
  assign \new_[5680]_  = A265 & A200;
  assign \new_[5681]_  = ~A199 & \new_[5680]_ ;
  assign \new_[5682]_  = \new_[5681]_  & \new_[5676]_ ;
  assign \new_[5685]_  = A267 & ~A266;
  assign \new_[5689]_  = A299 & A298;
  assign \new_[5690]_  = A268 & \new_[5689]_ ;
  assign \new_[5691]_  = \new_[5690]_  & \new_[5685]_ ;
  assign \new_[5694]_  = A167 & A168;
  assign \new_[5698]_  = A265 & A200;
  assign \new_[5699]_  = ~A199 & \new_[5698]_ ;
  assign \new_[5700]_  = \new_[5699]_  & \new_[5694]_ ;
  assign \new_[5703]_  = A267 & ~A266;
  assign \new_[5707]_  = ~A299 & ~A298;
  assign \new_[5708]_  = A268 & \new_[5707]_ ;
  assign \new_[5709]_  = \new_[5708]_  & \new_[5703]_ ;
  assign \new_[5712]_  = A167 & A168;
  assign \new_[5716]_  = A265 & A200;
  assign \new_[5717]_  = ~A199 & \new_[5716]_ ;
  assign \new_[5718]_  = \new_[5717]_  & \new_[5712]_ ;
  assign \new_[5721]_  = A267 & ~A266;
  assign \new_[5725]_  = ~A300 & A298;
  assign \new_[5726]_  = A269 & \new_[5725]_ ;
  assign \new_[5727]_  = \new_[5726]_  & \new_[5721]_ ;
  assign \new_[5730]_  = A167 & A168;
  assign \new_[5734]_  = A265 & A200;
  assign \new_[5735]_  = ~A199 & \new_[5734]_ ;
  assign \new_[5736]_  = \new_[5735]_  & \new_[5730]_ ;
  assign \new_[5739]_  = A267 & ~A266;
  assign \new_[5743]_  = A299 & A298;
  assign \new_[5744]_  = A269 & \new_[5743]_ ;
  assign \new_[5745]_  = \new_[5744]_  & \new_[5739]_ ;
  assign \new_[5748]_  = A167 & A168;
  assign \new_[5752]_  = A265 & A200;
  assign \new_[5753]_  = ~A199 & \new_[5752]_ ;
  assign \new_[5754]_  = \new_[5753]_  & \new_[5748]_ ;
  assign \new_[5757]_  = A267 & ~A266;
  assign \new_[5761]_  = ~A299 & ~A298;
  assign \new_[5762]_  = A269 & \new_[5761]_ ;
  assign \new_[5763]_  = \new_[5762]_  & \new_[5757]_ ;
  assign \new_[5766]_  = A167 & A168;
  assign \new_[5770]_  = ~A203 & ~A202;
  assign \new_[5771]_  = ~A200 & \new_[5770]_ ;
  assign \new_[5772]_  = \new_[5771]_  & \new_[5766]_ ;
  assign \new_[5775]_  = ~A268 & ~A266;
  assign \new_[5779]_  = A299 & ~A298;
  assign \new_[5780]_  = ~A269 & \new_[5779]_ ;
  assign \new_[5781]_  = \new_[5780]_  & \new_[5775]_ ;
  assign \new_[5784]_  = A167 & A168;
  assign \new_[5788]_  = A265 & ~A201;
  assign \new_[5789]_  = ~A200 & \new_[5788]_ ;
  assign \new_[5790]_  = \new_[5789]_  & \new_[5784]_ ;
  assign \new_[5793]_  = A298 & A266;
  assign \new_[5797]_  = A301 & A300;
  assign \new_[5798]_  = ~A299 & \new_[5797]_ ;
  assign \new_[5799]_  = \new_[5798]_  & \new_[5793]_ ;
  assign \new_[5802]_  = A167 & A168;
  assign \new_[5806]_  = A265 & ~A201;
  assign \new_[5807]_  = ~A200 & \new_[5806]_ ;
  assign \new_[5808]_  = \new_[5807]_  & \new_[5802]_ ;
  assign \new_[5811]_  = A298 & A266;
  assign \new_[5815]_  = A302 & A300;
  assign \new_[5816]_  = ~A299 & \new_[5815]_ ;
  assign \new_[5817]_  = \new_[5816]_  & \new_[5811]_ ;
  assign \new_[5820]_  = A167 & A168;
  assign \new_[5824]_  = ~A266 & ~A201;
  assign \new_[5825]_  = ~A200 & \new_[5824]_ ;
  assign \new_[5826]_  = \new_[5825]_  & \new_[5820]_ ;
  assign \new_[5829]_  = A298 & ~A267;
  assign \new_[5833]_  = A301 & A300;
  assign \new_[5834]_  = ~A299 & \new_[5833]_ ;
  assign \new_[5835]_  = \new_[5834]_  & \new_[5829]_ ;
  assign \new_[5838]_  = A167 & A168;
  assign \new_[5842]_  = ~A266 & ~A201;
  assign \new_[5843]_  = ~A200 & \new_[5842]_ ;
  assign \new_[5844]_  = \new_[5843]_  & \new_[5838]_ ;
  assign \new_[5847]_  = A298 & ~A267;
  assign \new_[5851]_  = A302 & A300;
  assign \new_[5852]_  = ~A299 & \new_[5851]_ ;
  assign \new_[5853]_  = \new_[5852]_  & \new_[5847]_ ;
  assign \new_[5856]_  = A167 & A168;
  assign \new_[5860]_  = ~A265 & ~A201;
  assign \new_[5861]_  = ~A200 & \new_[5860]_ ;
  assign \new_[5862]_  = \new_[5861]_  & \new_[5856]_ ;
  assign \new_[5865]_  = A298 & ~A266;
  assign \new_[5869]_  = A301 & A300;
  assign \new_[5870]_  = ~A299 & \new_[5869]_ ;
  assign \new_[5871]_  = \new_[5870]_  & \new_[5865]_ ;
  assign \new_[5874]_  = A167 & A168;
  assign \new_[5878]_  = ~A265 & ~A201;
  assign \new_[5879]_  = ~A200 & \new_[5878]_ ;
  assign \new_[5880]_  = \new_[5879]_  & \new_[5874]_ ;
  assign \new_[5883]_  = A298 & ~A266;
  assign \new_[5887]_  = A302 & A300;
  assign \new_[5888]_  = ~A299 & \new_[5887]_ ;
  assign \new_[5889]_  = \new_[5888]_  & \new_[5883]_ ;
  assign \new_[5892]_  = A167 & A168;
  assign \new_[5896]_  = A201 & ~A200;
  assign \new_[5897]_  = A199 & \new_[5896]_ ;
  assign \new_[5898]_  = \new_[5897]_  & \new_[5892]_ ;
  assign \new_[5901]_  = ~A265 & A202;
  assign \new_[5905]_  = ~A300 & A298;
  assign \new_[5906]_  = A266 & \new_[5905]_ ;
  assign \new_[5907]_  = \new_[5906]_  & \new_[5901]_ ;
  assign \new_[5910]_  = A167 & A168;
  assign \new_[5914]_  = A201 & ~A200;
  assign \new_[5915]_  = A199 & \new_[5914]_ ;
  assign \new_[5916]_  = \new_[5915]_  & \new_[5910]_ ;
  assign \new_[5919]_  = ~A265 & A202;
  assign \new_[5923]_  = A299 & A298;
  assign \new_[5924]_  = A266 & \new_[5923]_ ;
  assign \new_[5925]_  = \new_[5924]_  & \new_[5919]_ ;
  assign \new_[5928]_  = A167 & A168;
  assign \new_[5932]_  = A201 & ~A200;
  assign \new_[5933]_  = A199 & \new_[5932]_ ;
  assign \new_[5934]_  = \new_[5933]_  & \new_[5928]_ ;
  assign \new_[5937]_  = ~A265 & A202;
  assign \new_[5941]_  = ~A299 & ~A298;
  assign \new_[5942]_  = A266 & \new_[5941]_ ;
  assign \new_[5943]_  = \new_[5942]_  & \new_[5937]_ ;
  assign \new_[5946]_  = A167 & A168;
  assign \new_[5950]_  = A201 & ~A200;
  assign \new_[5951]_  = A199 & \new_[5950]_ ;
  assign \new_[5952]_  = \new_[5951]_  & \new_[5946]_ ;
  assign \new_[5955]_  = ~A265 & A203;
  assign \new_[5959]_  = ~A300 & A298;
  assign \new_[5960]_  = A266 & \new_[5959]_ ;
  assign \new_[5961]_  = \new_[5960]_  & \new_[5955]_ ;
  assign \new_[5964]_  = A167 & A168;
  assign \new_[5968]_  = A201 & ~A200;
  assign \new_[5969]_  = A199 & \new_[5968]_ ;
  assign \new_[5970]_  = \new_[5969]_  & \new_[5964]_ ;
  assign \new_[5973]_  = ~A265 & A203;
  assign \new_[5977]_  = A299 & A298;
  assign \new_[5978]_  = A266 & \new_[5977]_ ;
  assign \new_[5979]_  = \new_[5978]_  & \new_[5973]_ ;
  assign \new_[5982]_  = A167 & A168;
  assign \new_[5986]_  = A201 & ~A200;
  assign \new_[5987]_  = A199 & \new_[5986]_ ;
  assign \new_[5988]_  = \new_[5987]_  & \new_[5982]_ ;
  assign \new_[5991]_  = ~A265 & A203;
  assign \new_[5995]_  = ~A299 & ~A298;
  assign \new_[5996]_  = A266 & \new_[5995]_ ;
  assign \new_[5997]_  = \new_[5996]_  & \new_[5991]_ ;
  assign \new_[6000]_  = A167 & A168;
  assign \new_[6004]_  = A265 & ~A200;
  assign \new_[6005]_  = ~A199 & \new_[6004]_ ;
  assign \new_[6006]_  = \new_[6005]_  & \new_[6000]_ ;
  assign \new_[6009]_  = A298 & A266;
  assign \new_[6013]_  = A301 & A300;
  assign \new_[6014]_  = ~A299 & \new_[6013]_ ;
  assign \new_[6015]_  = \new_[6014]_  & \new_[6009]_ ;
  assign \new_[6018]_  = A167 & A168;
  assign \new_[6022]_  = A265 & ~A200;
  assign \new_[6023]_  = ~A199 & \new_[6022]_ ;
  assign \new_[6024]_  = \new_[6023]_  & \new_[6018]_ ;
  assign \new_[6027]_  = A298 & A266;
  assign \new_[6031]_  = A302 & A300;
  assign \new_[6032]_  = ~A299 & \new_[6031]_ ;
  assign \new_[6033]_  = \new_[6032]_  & \new_[6027]_ ;
  assign \new_[6036]_  = A167 & A168;
  assign \new_[6040]_  = ~A266 & ~A200;
  assign \new_[6041]_  = ~A199 & \new_[6040]_ ;
  assign \new_[6042]_  = \new_[6041]_  & \new_[6036]_ ;
  assign \new_[6045]_  = A298 & ~A267;
  assign \new_[6049]_  = A301 & A300;
  assign \new_[6050]_  = ~A299 & \new_[6049]_ ;
  assign \new_[6051]_  = \new_[6050]_  & \new_[6045]_ ;
  assign \new_[6054]_  = A167 & A168;
  assign \new_[6058]_  = ~A266 & ~A200;
  assign \new_[6059]_  = ~A199 & \new_[6058]_ ;
  assign \new_[6060]_  = \new_[6059]_  & \new_[6054]_ ;
  assign \new_[6063]_  = A298 & ~A267;
  assign \new_[6067]_  = A302 & A300;
  assign \new_[6068]_  = ~A299 & \new_[6067]_ ;
  assign \new_[6069]_  = \new_[6068]_  & \new_[6063]_ ;
  assign \new_[6072]_  = A167 & A168;
  assign \new_[6076]_  = ~A265 & ~A200;
  assign \new_[6077]_  = ~A199 & \new_[6076]_ ;
  assign \new_[6078]_  = \new_[6077]_  & \new_[6072]_ ;
  assign \new_[6081]_  = A298 & ~A266;
  assign \new_[6085]_  = A301 & A300;
  assign \new_[6086]_  = ~A299 & \new_[6085]_ ;
  assign \new_[6087]_  = \new_[6086]_  & \new_[6081]_ ;
  assign \new_[6090]_  = A167 & A168;
  assign \new_[6094]_  = ~A265 & ~A200;
  assign \new_[6095]_  = ~A199 & \new_[6094]_ ;
  assign \new_[6096]_  = \new_[6095]_  & \new_[6090]_ ;
  assign \new_[6099]_  = A298 & ~A266;
  assign \new_[6103]_  = A302 & A300;
  assign \new_[6104]_  = ~A299 & \new_[6103]_ ;
  assign \new_[6105]_  = \new_[6104]_  & \new_[6099]_ ;
  assign \new_[6108]_  = ~A167 & A170;
  assign \new_[6112]_  = A200 & A199;
  assign \new_[6113]_  = ~A166 & \new_[6112]_ ;
  assign \new_[6114]_  = \new_[6113]_  & \new_[6108]_ ;
  assign \new_[6117]_  = A266 & ~A265;
  assign \new_[6121]_  = ~A302 & ~A301;
  assign \new_[6122]_  = A298 & \new_[6121]_ ;
  assign \new_[6123]_  = \new_[6122]_  & \new_[6117]_ ;
  assign \new_[6126]_  = ~A167 & A170;
  assign \new_[6130]_  = A200 & ~A199;
  assign \new_[6131]_  = ~A166 & \new_[6130]_ ;
  assign \new_[6132]_  = \new_[6131]_  & \new_[6126]_ ;
  assign \new_[6135]_  = ~A268 & ~A266;
  assign \new_[6139]_  = A299 & ~A298;
  assign \new_[6140]_  = ~A269 & \new_[6139]_ ;
  assign \new_[6141]_  = \new_[6140]_  & \new_[6135]_ ;
  assign \new_[6144]_  = ~A167 & A170;
  assign \new_[6148]_  = ~A202 & ~A200;
  assign \new_[6149]_  = ~A166 & \new_[6148]_ ;
  assign \new_[6150]_  = \new_[6149]_  & \new_[6144]_ ;
  assign \new_[6153]_  = ~A265 & ~A203;
  assign \new_[6157]_  = ~A300 & A298;
  assign \new_[6158]_  = A266 & \new_[6157]_ ;
  assign \new_[6159]_  = \new_[6158]_  & \new_[6153]_ ;
  assign \new_[6162]_  = ~A167 & A170;
  assign \new_[6166]_  = ~A202 & ~A200;
  assign \new_[6167]_  = ~A166 & \new_[6166]_ ;
  assign \new_[6168]_  = \new_[6167]_  & \new_[6162]_ ;
  assign \new_[6171]_  = ~A265 & ~A203;
  assign \new_[6175]_  = A299 & A298;
  assign \new_[6176]_  = A266 & \new_[6175]_ ;
  assign \new_[6177]_  = \new_[6176]_  & \new_[6171]_ ;
  assign \new_[6180]_  = ~A167 & A170;
  assign \new_[6184]_  = ~A202 & ~A200;
  assign \new_[6185]_  = ~A166 & \new_[6184]_ ;
  assign \new_[6186]_  = \new_[6185]_  & \new_[6180]_ ;
  assign \new_[6189]_  = ~A265 & ~A203;
  assign \new_[6193]_  = ~A299 & ~A298;
  assign \new_[6194]_  = A266 & \new_[6193]_ ;
  assign \new_[6195]_  = \new_[6194]_  & \new_[6189]_ ;
  assign \new_[6198]_  = ~A167 & A170;
  assign \new_[6202]_  = ~A201 & ~A200;
  assign \new_[6203]_  = ~A166 & \new_[6202]_ ;
  assign \new_[6204]_  = \new_[6203]_  & \new_[6198]_ ;
  assign \new_[6207]_  = A266 & ~A265;
  assign \new_[6211]_  = ~A302 & ~A301;
  assign \new_[6212]_  = A298 & \new_[6211]_ ;
  assign \new_[6213]_  = \new_[6212]_  & \new_[6207]_ ;
  assign \new_[6216]_  = ~A167 & A170;
  assign \new_[6220]_  = ~A200 & ~A199;
  assign \new_[6221]_  = ~A166 & \new_[6220]_ ;
  assign \new_[6222]_  = \new_[6221]_  & \new_[6216]_ ;
  assign \new_[6225]_  = A266 & ~A265;
  assign \new_[6229]_  = ~A302 & ~A301;
  assign \new_[6230]_  = A298 & \new_[6229]_ ;
  assign \new_[6231]_  = \new_[6230]_  & \new_[6225]_ ;
  assign \new_[6234]_  = ~A168 & A169;
  assign \new_[6238]_  = A199 & ~A166;
  assign \new_[6239]_  = A167 & \new_[6238]_ ;
  assign \new_[6240]_  = \new_[6239]_  & \new_[6234]_ ;
  assign \new_[6243]_  = ~A265 & A200;
  assign \new_[6247]_  = ~A300 & A298;
  assign \new_[6248]_  = A266 & \new_[6247]_ ;
  assign \new_[6249]_  = \new_[6248]_  & \new_[6243]_ ;
  assign \new_[6252]_  = ~A168 & A169;
  assign \new_[6256]_  = A199 & ~A166;
  assign \new_[6257]_  = A167 & \new_[6256]_ ;
  assign \new_[6258]_  = \new_[6257]_  & \new_[6252]_ ;
  assign \new_[6261]_  = ~A265 & A200;
  assign \new_[6265]_  = A299 & A298;
  assign \new_[6266]_  = A266 & \new_[6265]_ ;
  assign \new_[6267]_  = \new_[6266]_  & \new_[6261]_ ;
  assign \new_[6270]_  = ~A168 & A169;
  assign \new_[6274]_  = A199 & ~A166;
  assign \new_[6275]_  = A167 & \new_[6274]_ ;
  assign \new_[6276]_  = \new_[6275]_  & \new_[6270]_ ;
  assign \new_[6279]_  = ~A265 & A200;
  assign \new_[6283]_  = ~A299 & ~A298;
  assign \new_[6284]_  = A266 & \new_[6283]_ ;
  assign \new_[6285]_  = \new_[6284]_  & \new_[6279]_ ;
  assign \new_[6288]_  = ~A168 & A169;
  assign \new_[6292]_  = ~A199 & ~A166;
  assign \new_[6293]_  = A167 & \new_[6292]_ ;
  assign \new_[6294]_  = \new_[6293]_  & \new_[6288]_ ;
  assign \new_[6297]_  = A265 & A200;
  assign \new_[6301]_  = A299 & ~A298;
  assign \new_[6302]_  = A266 & \new_[6301]_ ;
  assign \new_[6303]_  = \new_[6302]_  & \new_[6297]_ ;
  assign \new_[6306]_  = ~A168 & A169;
  assign \new_[6310]_  = ~A199 & ~A166;
  assign \new_[6311]_  = A167 & \new_[6310]_ ;
  assign \new_[6312]_  = \new_[6311]_  & \new_[6306]_ ;
  assign \new_[6315]_  = ~A266 & A200;
  assign \new_[6319]_  = A299 & ~A298;
  assign \new_[6320]_  = ~A267 & \new_[6319]_ ;
  assign \new_[6321]_  = \new_[6320]_  & \new_[6315]_ ;
  assign \new_[6324]_  = ~A168 & A169;
  assign \new_[6328]_  = ~A199 & ~A166;
  assign \new_[6329]_  = A167 & \new_[6328]_ ;
  assign \new_[6330]_  = \new_[6329]_  & \new_[6324]_ ;
  assign \new_[6333]_  = ~A265 & A200;
  assign \new_[6337]_  = A299 & ~A298;
  assign \new_[6338]_  = ~A266 & \new_[6337]_ ;
  assign \new_[6339]_  = \new_[6338]_  & \new_[6333]_ ;
  assign \new_[6342]_  = ~A168 & A169;
  assign \new_[6346]_  = ~A200 & ~A166;
  assign \new_[6347]_  = A167 & \new_[6346]_ ;
  assign \new_[6348]_  = \new_[6347]_  & \new_[6342]_ ;
  assign \new_[6351]_  = ~A265 & ~A201;
  assign \new_[6355]_  = ~A300 & A298;
  assign \new_[6356]_  = A266 & \new_[6355]_ ;
  assign \new_[6357]_  = \new_[6356]_  & \new_[6351]_ ;
  assign \new_[6360]_  = ~A168 & A169;
  assign \new_[6364]_  = ~A200 & ~A166;
  assign \new_[6365]_  = A167 & \new_[6364]_ ;
  assign \new_[6366]_  = \new_[6365]_  & \new_[6360]_ ;
  assign \new_[6369]_  = ~A265 & ~A201;
  assign \new_[6373]_  = A299 & A298;
  assign \new_[6374]_  = A266 & \new_[6373]_ ;
  assign \new_[6375]_  = \new_[6374]_  & \new_[6369]_ ;
  assign \new_[6378]_  = ~A168 & A169;
  assign \new_[6382]_  = ~A200 & ~A166;
  assign \new_[6383]_  = A167 & \new_[6382]_ ;
  assign \new_[6384]_  = \new_[6383]_  & \new_[6378]_ ;
  assign \new_[6387]_  = ~A265 & ~A201;
  assign \new_[6391]_  = ~A299 & ~A298;
  assign \new_[6392]_  = A266 & \new_[6391]_ ;
  assign \new_[6393]_  = \new_[6392]_  & \new_[6387]_ ;
  assign \new_[6396]_  = ~A168 & A169;
  assign \new_[6400]_  = ~A199 & ~A166;
  assign \new_[6401]_  = A167 & \new_[6400]_ ;
  assign \new_[6402]_  = \new_[6401]_  & \new_[6396]_ ;
  assign \new_[6405]_  = ~A265 & ~A200;
  assign \new_[6409]_  = ~A300 & A298;
  assign \new_[6410]_  = A266 & \new_[6409]_ ;
  assign \new_[6411]_  = \new_[6410]_  & \new_[6405]_ ;
  assign \new_[6414]_  = ~A168 & A169;
  assign \new_[6418]_  = ~A199 & ~A166;
  assign \new_[6419]_  = A167 & \new_[6418]_ ;
  assign \new_[6420]_  = \new_[6419]_  & \new_[6414]_ ;
  assign \new_[6423]_  = ~A265 & ~A200;
  assign \new_[6427]_  = A299 & A298;
  assign \new_[6428]_  = A266 & \new_[6427]_ ;
  assign \new_[6429]_  = \new_[6428]_  & \new_[6423]_ ;
  assign \new_[6432]_  = ~A168 & A169;
  assign \new_[6436]_  = ~A199 & ~A166;
  assign \new_[6437]_  = A167 & \new_[6436]_ ;
  assign \new_[6438]_  = \new_[6437]_  & \new_[6432]_ ;
  assign \new_[6441]_  = ~A265 & ~A200;
  assign \new_[6445]_  = ~A299 & ~A298;
  assign \new_[6446]_  = A266 & \new_[6445]_ ;
  assign \new_[6447]_  = \new_[6446]_  & \new_[6441]_ ;
  assign \new_[6450]_  = ~A168 & A169;
  assign \new_[6454]_  = A199 & A166;
  assign \new_[6455]_  = ~A167 & \new_[6454]_ ;
  assign \new_[6456]_  = \new_[6455]_  & \new_[6450]_ ;
  assign \new_[6459]_  = ~A265 & A200;
  assign \new_[6463]_  = ~A300 & A298;
  assign \new_[6464]_  = A266 & \new_[6463]_ ;
  assign \new_[6465]_  = \new_[6464]_  & \new_[6459]_ ;
  assign \new_[6468]_  = ~A168 & A169;
  assign \new_[6472]_  = A199 & A166;
  assign \new_[6473]_  = ~A167 & \new_[6472]_ ;
  assign \new_[6474]_  = \new_[6473]_  & \new_[6468]_ ;
  assign \new_[6477]_  = ~A265 & A200;
  assign \new_[6481]_  = A299 & A298;
  assign \new_[6482]_  = A266 & \new_[6481]_ ;
  assign \new_[6483]_  = \new_[6482]_  & \new_[6477]_ ;
  assign \new_[6486]_  = ~A168 & A169;
  assign \new_[6490]_  = A199 & A166;
  assign \new_[6491]_  = ~A167 & \new_[6490]_ ;
  assign \new_[6492]_  = \new_[6491]_  & \new_[6486]_ ;
  assign \new_[6495]_  = ~A265 & A200;
  assign \new_[6499]_  = ~A299 & ~A298;
  assign \new_[6500]_  = A266 & \new_[6499]_ ;
  assign \new_[6501]_  = \new_[6500]_  & \new_[6495]_ ;
  assign \new_[6504]_  = ~A168 & A169;
  assign \new_[6508]_  = ~A199 & A166;
  assign \new_[6509]_  = ~A167 & \new_[6508]_ ;
  assign \new_[6510]_  = \new_[6509]_  & \new_[6504]_ ;
  assign \new_[6513]_  = A265 & A200;
  assign \new_[6517]_  = A299 & ~A298;
  assign \new_[6518]_  = A266 & \new_[6517]_ ;
  assign \new_[6519]_  = \new_[6518]_  & \new_[6513]_ ;
  assign \new_[6522]_  = ~A168 & A169;
  assign \new_[6526]_  = ~A199 & A166;
  assign \new_[6527]_  = ~A167 & \new_[6526]_ ;
  assign \new_[6528]_  = \new_[6527]_  & \new_[6522]_ ;
  assign \new_[6531]_  = ~A266 & A200;
  assign \new_[6535]_  = A299 & ~A298;
  assign \new_[6536]_  = ~A267 & \new_[6535]_ ;
  assign \new_[6537]_  = \new_[6536]_  & \new_[6531]_ ;
  assign \new_[6540]_  = ~A168 & A169;
  assign \new_[6544]_  = ~A199 & A166;
  assign \new_[6545]_  = ~A167 & \new_[6544]_ ;
  assign \new_[6546]_  = \new_[6545]_  & \new_[6540]_ ;
  assign \new_[6549]_  = ~A265 & A200;
  assign \new_[6553]_  = A299 & ~A298;
  assign \new_[6554]_  = ~A266 & \new_[6553]_ ;
  assign \new_[6555]_  = \new_[6554]_  & \new_[6549]_ ;
  assign \new_[6558]_  = ~A168 & A169;
  assign \new_[6562]_  = ~A200 & A166;
  assign \new_[6563]_  = ~A167 & \new_[6562]_ ;
  assign \new_[6564]_  = \new_[6563]_  & \new_[6558]_ ;
  assign \new_[6567]_  = ~A265 & ~A201;
  assign \new_[6571]_  = ~A300 & A298;
  assign \new_[6572]_  = A266 & \new_[6571]_ ;
  assign \new_[6573]_  = \new_[6572]_  & \new_[6567]_ ;
  assign \new_[6576]_  = ~A168 & A169;
  assign \new_[6580]_  = ~A200 & A166;
  assign \new_[6581]_  = ~A167 & \new_[6580]_ ;
  assign \new_[6582]_  = \new_[6581]_  & \new_[6576]_ ;
  assign \new_[6585]_  = ~A265 & ~A201;
  assign \new_[6589]_  = A299 & A298;
  assign \new_[6590]_  = A266 & \new_[6589]_ ;
  assign \new_[6591]_  = \new_[6590]_  & \new_[6585]_ ;
  assign \new_[6594]_  = ~A168 & A169;
  assign \new_[6598]_  = ~A200 & A166;
  assign \new_[6599]_  = ~A167 & \new_[6598]_ ;
  assign \new_[6600]_  = \new_[6599]_  & \new_[6594]_ ;
  assign \new_[6603]_  = ~A265 & ~A201;
  assign \new_[6607]_  = ~A299 & ~A298;
  assign \new_[6608]_  = A266 & \new_[6607]_ ;
  assign \new_[6609]_  = \new_[6608]_  & \new_[6603]_ ;
  assign \new_[6612]_  = ~A168 & A169;
  assign \new_[6616]_  = ~A199 & A166;
  assign \new_[6617]_  = ~A167 & \new_[6616]_ ;
  assign \new_[6618]_  = \new_[6617]_  & \new_[6612]_ ;
  assign \new_[6621]_  = ~A265 & ~A200;
  assign \new_[6625]_  = ~A300 & A298;
  assign \new_[6626]_  = A266 & \new_[6625]_ ;
  assign \new_[6627]_  = \new_[6626]_  & \new_[6621]_ ;
  assign \new_[6630]_  = ~A168 & A169;
  assign \new_[6634]_  = ~A199 & A166;
  assign \new_[6635]_  = ~A167 & \new_[6634]_ ;
  assign \new_[6636]_  = \new_[6635]_  & \new_[6630]_ ;
  assign \new_[6639]_  = ~A265 & ~A200;
  assign \new_[6643]_  = A299 & A298;
  assign \new_[6644]_  = A266 & \new_[6643]_ ;
  assign \new_[6645]_  = \new_[6644]_  & \new_[6639]_ ;
  assign \new_[6648]_  = ~A168 & A169;
  assign \new_[6652]_  = ~A199 & A166;
  assign \new_[6653]_  = ~A167 & \new_[6652]_ ;
  assign \new_[6654]_  = \new_[6653]_  & \new_[6648]_ ;
  assign \new_[6657]_  = ~A265 & ~A200;
  assign \new_[6661]_  = ~A299 & ~A298;
  assign \new_[6662]_  = A266 & \new_[6661]_ ;
  assign \new_[6663]_  = \new_[6662]_  & \new_[6657]_ ;
  assign \new_[6666]_  = A169 & A170;
  assign \new_[6670]_  = A200 & A199;
  assign \new_[6671]_  = ~A168 & \new_[6670]_ ;
  assign \new_[6672]_  = \new_[6671]_  & \new_[6666]_ ;
  assign \new_[6675]_  = A266 & ~A265;
  assign \new_[6679]_  = ~A302 & ~A301;
  assign \new_[6680]_  = A298 & \new_[6679]_ ;
  assign \new_[6681]_  = \new_[6680]_  & \new_[6675]_ ;
  assign \new_[6684]_  = A169 & A170;
  assign \new_[6688]_  = A200 & ~A199;
  assign \new_[6689]_  = ~A168 & \new_[6688]_ ;
  assign \new_[6690]_  = \new_[6689]_  & \new_[6684]_ ;
  assign \new_[6693]_  = ~A268 & ~A266;
  assign \new_[6697]_  = A299 & ~A298;
  assign \new_[6698]_  = ~A269 & \new_[6697]_ ;
  assign \new_[6699]_  = \new_[6698]_  & \new_[6693]_ ;
  assign \new_[6702]_  = A169 & A170;
  assign \new_[6706]_  = ~A202 & ~A200;
  assign \new_[6707]_  = ~A168 & \new_[6706]_ ;
  assign \new_[6708]_  = \new_[6707]_  & \new_[6702]_ ;
  assign \new_[6711]_  = ~A265 & ~A203;
  assign \new_[6715]_  = ~A300 & A298;
  assign \new_[6716]_  = A266 & \new_[6715]_ ;
  assign \new_[6717]_  = \new_[6716]_  & \new_[6711]_ ;
  assign \new_[6720]_  = A169 & A170;
  assign \new_[6724]_  = ~A202 & ~A200;
  assign \new_[6725]_  = ~A168 & \new_[6724]_ ;
  assign \new_[6726]_  = \new_[6725]_  & \new_[6720]_ ;
  assign \new_[6729]_  = ~A265 & ~A203;
  assign \new_[6733]_  = A299 & A298;
  assign \new_[6734]_  = A266 & \new_[6733]_ ;
  assign \new_[6735]_  = \new_[6734]_  & \new_[6729]_ ;
  assign \new_[6738]_  = A169 & A170;
  assign \new_[6742]_  = ~A202 & ~A200;
  assign \new_[6743]_  = ~A168 & \new_[6742]_ ;
  assign \new_[6744]_  = \new_[6743]_  & \new_[6738]_ ;
  assign \new_[6747]_  = ~A265 & ~A203;
  assign \new_[6751]_  = ~A299 & ~A298;
  assign \new_[6752]_  = A266 & \new_[6751]_ ;
  assign \new_[6753]_  = \new_[6752]_  & \new_[6747]_ ;
  assign \new_[6756]_  = A169 & A170;
  assign \new_[6760]_  = ~A201 & ~A200;
  assign \new_[6761]_  = ~A168 & \new_[6760]_ ;
  assign \new_[6762]_  = \new_[6761]_  & \new_[6756]_ ;
  assign \new_[6765]_  = A266 & ~A265;
  assign \new_[6769]_  = ~A302 & ~A301;
  assign \new_[6770]_  = A298 & \new_[6769]_ ;
  assign \new_[6771]_  = \new_[6770]_  & \new_[6765]_ ;
  assign \new_[6774]_  = A169 & A170;
  assign \new_[6778]_  = ~A200 & ~A199;
  assign \new_[6779]_  = ~A168 & \new_[6778]_ ;
  assign \new_[6780]_  = \new_[6779]_  & \new_[6774]_ ;
  assign \new_[6783]_  = A266 & ~A265;
  assign \new_[6787]_  = ~A302 & ~A301;
  assign \new_[6788]_  = A298 & \new_[6787]_ ;
  assign \new_[6789]_  = \new_[6788]_  & \new_[6783]_ ;
  assign \new_[6792]_  = A169 & ~A170;
  assign \new_[6796]_  = A199 & A166;
  assign \new_[6797]_  = A167 & \new_[6796]_ ;
  assign \new_[6798]_  = \new_[6797]_  & \new_[6792]_ ;
  assign \new_[6801]_  = A265 & A200;
  assign \new_[6805]_  = A299 & ~A298;
  assign \new_[6806]_  = A266 & \new_[6805]_ ;
  assign \new_[6807]_  = \new_[6806]_  & \new_[6801]_ ;
  assign \new_[6810]_  = A169 & ~A170;
  assign \new_[6814]_  = A199 & A166;
  assign \new_[6815]_  = A167 & \new_[6814]_ ;
  assign \new_[6816]_  = \new_[6815]_  & \new_[6810]_ ;
  assign \new_[6819]_  = ~A266 & A200;
  assign \new_[6823]_  = A299 & ~A298;
  assign \new_[6824]_  = ~A267 & \new_[6823]_ ;
  assign \new_[6825]_  = \new_[6824]_  & \new_[6819]_ ;
  assign \new_[6828]_  = A169 & ~A170;
  assign \new_[6832]_  = A199 & A166;
  assign \new_[6833]_  = A167 & \new_[6832]_ ;
  assign \new_[6834]_  = \new_[6833]_  & \new_[6828]_ ;
  assign \new_[6837]_  = ~A265 & A200;
  assign \new_[6841]_  = A299 & ~A298;
  assign \new_[6842]_  = ~A266 & \new_[6841]_ ;
  assign \new_[6843]_  = \new_[6842]_  & \new_[6837]_ ;
  assign \new_[6846]_  = A169 & ~A170;
  assign \new_[6850]_  = ~A199 & A166;
  assign \new_[6851]_  = A167 & \new_[6850]_ ;
  assign \new_[6852]_  = \new_[6851]_  & \new_[6846]_ ;
  assign \new_[6855]_  = ~A265 & A200;
  assign \new_[6859]_  = ~A300 & A298;
  assign \new_[6860]_  = A266 & \new_[6859]_ ;
  assign \new_[6861]_  = \new_[6860]_  & \new_[6855]_ ;
  assign \new_[6864]_  = A169 & ~A170;
  assign \new_[6868]_  = ~A199 & A166;
  assign \new_[6869]_  = A167 & \new_[6868]_ ;
  assign \new_[6870]_  = \new_[6869]_  & \new_[6864]_ ;
  assign \new_[6873]_  = ~A265 & A200;
  assign \new_[6877]_  = A299 & A298;
  assign \new_[6878]_  = A266 & \new_[6877]_ ;
  assign \new_[6879]_  = \new_[6878]_  & \new_[6873]_ ;
  assign \new_[6882]_  = A169 & ~A170;
  assign \new_[6886]_  = ~A199 & A166;
  assign \new_[6887]_  = A167 & \new_[6886]_ ;
  assign \new_[6888]_  = \new_[6887]_  & \new_[6882]_ ;
  assign \new_[6891]_  = ~A265 & A200;
  assign \new_[6895]_  = ~A299 & ~A298;
  assign \new_[6896]_  = A266 & \new_[6895]_ ;
  assign \new_[6897]_  = \new_[6896]_  & \new_[6891]_ ;
  assign \new_[6900]_  = A169 & ~A170;
  assign \new_[6904]_  = ~A200 & A166;
  assign \new_[6905]_  = A167 & \new_[6904]_ ;
  assign \new_[6906]_  = \new_[6905]_  & \new_[6900]_ ;
  assign \new_[6909]_  = A265 & ~A201;
  assign \new_[6913]_  = A299 & ~A298;
  assign \new_[6914]_  = A266 & \new_[6913]_ ;
  assign \new_[6915]_  = \new_[6914]_  & \new_[6909]_ ;
  assign \new_[6918]_  = A169 & ~A170;
  assign \new_[6922]_  = ~A200 & A166;
  assign \new_[6923]_  = A167 & \new_[6922]_ ;
  assign \new_[6924]_  = \new_[6923]_  & \new_[6918]_ ;
  assign \new_[6927]_  = ~A266 & ~A201;
  assign \new_[6931]_  = A299 & ~A298;
  assign \new_[6932]_  = ~A267 & \new_[6931]_ ;
  assign \new_[6933]_  = \new_[6932]_  & \new_[6927]_ ;
  assign \new_[6936]_  = A169 & ~A170;
  assign \new_[6940]_  = ~A200 & A166;
  assign \new_[6941]_  = A167 & \new_[6940]_ ;
  assign \new_[6942]_  = \new_[6941]_  & \new_[6936]_ ;
  assign \new_[6945]_  = ~A265 & ~A201;
  assign \new_[6949]_  = A299 & ~A298;
  assign \new_[6950]_  = ~A266 & \new_[6949]_ ;
  assign \new_[6951]_  = \new_[6950]_  & \new_[6945]_ ;
  assign \new_[6954]_  = A169 & ~A170;
  assign \new_[6958]_  = ~A199 & A166;
  assign \new_[6959]_  = A167 & \new_[6958]_ ;
  assign \new_[6960]_  = \new_[6959]_  & \new_[6954]_ ;
  assign \new_[6963]_  = A265 & ~A200;
  assign \new_[6967]_  = A299 & ~A298;
  assign \new_[6968]_  = A266 & \new_[6967]_ ;
  assign \new_[6969]_  = \new_[6968]_  & \new_[6963]_ ;
  assign \new_[6972]_  = A169 & ~A170;
  assign \new_[6976]_  = ~A199 & A166;
  assign \new_[6977]_  = A167 & \new_[6976]_ ;
  assign \new_[6978]_  = \new_[6977]_  & \new_[6972]_ ;
  assign \new_[6981]_  = ~A266 & ~A200;
  assign \new_[6985]_  = A299 & ~A298;
  assign \new_[6986]_  = ~A267 & \new_[6985]_ ;
  assign \new_[6987]_  = \new_[6986]_  & \new_[6981]_ ;
  assign \new_[6990]_  = A169 & ~A170;
  assign \new_[6994]_  = ~A199 & A166;
  assign \new_[6995]_  = A167 & \new_[6994]_ ;
  assign \new_[6996]_  = \new_[6995]_  & \new_[6990]_ ;
  assign \new_[6999]_  = ~A265 & ~A200;
  assign \new_[7003]_  = A299 & ~A298;
  assign \new_[7004]_  = ~A266 & \new_[7003]_ ;
  assign \new_[7005]_  = \new_[7004]_  & \new_[6999]_ ;
  assign \new_[7008]_  = A169 & ~A170;
  assign \new_[7012]_  = A199 & ~A166;
  assign \new_[7013]_  = ~A167 & \new_[7012]_ ;
  assign \new_[7014]_  = \new_[7013]_  & \new_[7008]_ ;
  assign \new_[7017]_  = A265 & A200;
  assign \new_[7021]_  = A299 & ~A298;
  assign \new_[7022]_  = A266 & \new_[7021]_ ;
  assign \new_[7023]_  = \new_[7022]_  & \new_[7017]_ ;
  assign \new_[7026]_  = A169 & ~A170;
  assign \new_[7030]_  = A199 & ~A166;
  assign \new_[7031]_  = ~A167 & \new_[7030]_ ;
  assign \new_[7032]_  = \new_[7031]_  & \new_[7026]_ ;
  assign \new_[7035]_  = ~A266 & A200;
  assign \new_[7039]_  = A299 & ~A298;
  assign \new_[7040]_  = ~A267 & \new_[7039]_ ;
  assign \new_[7041]_  = \new_[7040]_  & \new_[7035]_ ;
  assign \new_[7044]_  = A169 & ~A170;
  assign \new_[7048]_  = A199 & ~A166;
  assign \new_[7049]_  = ~A167 & \new_[7048]_ ;
  assign \new_[7050]_  = \new_[7049]_  & \new_[7044]_ ;
  assign \new_[7053]_  = ~A265 & A200;
  assign \new_[7057]_  = A299 & ~A298;
  assign \new_[7058]_  = ~A266 & \new_[7057]_ ;
  assign \new_[7059]_  = \new_[7058]_  & \new_[7053]_ ;
  assign \new_[7062]_  = A169 & ~A170;
  assign \new_[7066]_  = ~A199 & ~A166;
  assign \new_[7067]_  = ~A167 & \new_[7066]_ ;
  assign \new_[7068]_  = \new_[7067]_  & \new_[7062]_ ;
  assign \new_[7071]_  = ~A265 & A200;
  assign \new_[7075]_  = ~A300 & A298;
  assign \new_[7076]_  = A266 & \new_[7075]_ ;
  assign \new_[7077]_  = \new_[7076]_  & \new_[7071]_ ;
  assign \new_[7080]_  = A169 & ~A170;
  assign \new_[7084]_  = ~A199 & ~A166;
  assign \new_[7085]_  = ~A167 & \new_[7084]_ ;
  assign \new_[7086]_  = \new_[7085]_  & \new_[7080]_ ;
  assign \new_[7089]_  = ~A265 & A200;
  assign \new_[7093]_  = A299 & A298;
  assign \new_[7094]_  = A266 & \new_[7093]_ ;
  assign \new_[7095]_  = \new_[7094]_  & \new_[7089]_ ;
  assign \new_[7098]_  = A169 & ~A170;
  assign \new_[7102]_  = ~A199 & ~A166;
  assign \new_[7103]_  = ~A167 & \new_[7102]_ ;
  assign \new_[7104]_  = \new_[7103]_  & \new_[7098]_ ;
  assign \new_[7107]_  = ~A265 & A200;
  assign \new_[7111]_  = ~A299 & ~A298;
  assign \new_[7112]_  = A266 & \new_[7111]_ ;
  assign \new_[7113]_  = \new_[7112]_  & \new_[7107]_ ;
  assign \new_[7116]_  = A169 & ~A170;
  assign \new_[7120]_  = ~A200 & ~A166;
  assign \new_[7121]_  = ~A167 & \new_[7120]_ ;
  assign \new_[7122]_  = \new_[7121]_  & \new_[7116]_ ;
  assign \new_[7125]_  = A265 & ~A201;
  assign \new_[7129]_  = A299 & ~A298;
  assign \new_[7130]_  = A266 & \new_[7129]_ ;
  assign \new_[7131]_  = \new_[7130]_  & \new_[7125]_ ;
  assign \new_[7134]_  = A169 & ~A170;
  assign \new_[7138]_  = ~A200 & ~A166;
  assign \new_[7139]_  = ~A167 & \new_[7138]_ ;
  assign \new_[7140]_  = \new_[7139]_  & \new_[7134]_ ;
  assign \new_[7143]_  = ~A266 & ~A201;
  assign \new_[7147]_  = A299 & ~A298;
  assign \new_[7148]_  = ~A267 & \new_[7147]_ ;
  assign \new_[7149]_  = \new_[7148]_  & \new_[7143]_ ;
  assign \new_[7152]_  = A169 & ~A170;
  assign \new_[7156]_  = ~A200 & ~A166;
  assign \new_[7157]_  = ~A167 & \new_[7156]_ ;
  assign \new_[7158]_  = \new_[7157]_  & \new_[7152]_ ;
  assign \new_[7161]_  = ~A265 & ~A201;
  assign \new_[7165]_  = A299 & ~A298;
  assign \new_[7166]_  = ~A266 & \new_[7165]_ ;
  assign \new_[7167]_  = \new_[7166]_  & \new_[7161]_ ;
  assign \new_[7170]_  = A169 & ~A170;
  assign \new_[7174]_  = ~A199 & ~A166;
  assign \new_[7175]_  = ~A167 & \new_[7174]_ ;
  assign \new_[7176]_  = \new_[7175]_  & \new_[7170]_ ;
  assign \new_[7179]_  = A265 & ~A200;
  assign \new_[7183]_  = A299 & ~A298;
  assign \new_[7184]_  = A266 & \new_[7183]_ ;
  assign \new_[7185]_  = \new_[7184]_  & \new_[7179]_ ;
  assign \new_[7188]_  = A169 & ~A170;
  assign \new_[7192]_  = ~A199 & ~A166;
  assign \new_[7193]_  = ~A167 & \new_[7192]_ ;
  assign \new_[7194]_  = \new_[7193]_  & \new_[7188]_ ;
  assign \new_[7197]_  = ~A266 & ~A200;
  assign \new_[7201]_  = A299 & ~A298;
  assign \new_[7202]_  = ~A267 & \new_[7201]_ ;
  assign \new_[7203]_  = \new_[7202]_  & \new_[7197]_ ;
  assign \new_[7206]_  = A169 & ~A170;
  assign \new_[7210]_  = ~A199 & ~A166;
  assign \new_[7211]_  = ~A167 & \new_[7210]_ ;
  assign \new_[7212]_  = \new_[7211]_  & \new_[7206]_ ;
  assign \new_[7215]_  = ~A265 & ~A200;
  assign \new_[7219]_  = A299 & ~A298;
  assign \new_[7220]_  = ~A266 & \new_[7219]_ ;
  assign \new_[7221]_  = \new_[7220]_  & \new_[7215]_ ;
  assign \new_[7224]_  = ~A167 & ~A169;
  assign \new_[7228]_  = A200 & A199;
  assign \new_[7229]_  = ~A166 & \new_[7228]_ ;
  assign \new_[7230]_  = \new_[7229]_  & \new_[7224]_ ;
  assign \new_[7233]_  = A266 & ~A265;
  assign \new_[7237]_  = ~A302 & ~A301;
  assign \new_[7238]_  = A298 & \new_[7237]_ ;
  assign \new_[7239]_  = \new_[7238]_  & \new_[7233]_ ;
  assign \new_[7242]_  = ~A167 & ~A169;
  assign \new_[7246]_  = A200 & ~A199;
  assign \new_[7247]_  = ~A166 & \new_[7246]_ ;
  assign \new_[7248]_  = \new_[7247]_  & \new_[7242]_ ;
  assign \new_[7251]_  = ~A268 & ~A266;
  assign \new_[7255]_  = A299 & ~A298;
  assign \new_[7256]_  = ~A269 & \new_[7255]_ ;
  assign \new_[7257]_  = \new_[7256]_  & \new_[7251]_ ;
  assign \new_[7260]_  = ~A167 & ~A169;
  assign \new_[7264]_  = ~A202 & ~A200;
  assign \new_[7265]_  = ~A166 & \new_[7264]_ ;
  assign \new_[7266]_  = \new_[7265]_  & \new_[7260]_ ;
  assign \new_[7269]_  = ~A265 & ~A203;
  assign \new_[7273]_  = ~A300 & A298;
  assign \new_[7274]_  = A266 & \new_[7273]_ ;
  assign \new_[7275]_  = \new_[7274]_  & \new_[7269]_ ;
  assign \new_[7278]_  = ~A167 & ~A169;
  assign \new_[7282]_  = ~A202 & ~A200;
  assign \new_[7283]_  = ~A166 & \new_[7282]_ ;
  assign \new_[7284]_  = \new_[7283]_  & \new_[7278]_ ;
  assign \new_[7287]_  = ~A265 & ~A203;
  assign \new_[7291]_  = A299 & A298;
  assign \new_[7292]_  = A266 & \new_[7291]_ ;
  assign \new_[7293]_  = \new_[7292]_  & \new_[7287]_ ;
  assign \new_[7296]_  = ~A167 & ~A169;
  assign \new_[7300]_  = ~A202 & ~A200;
  assign \new_[7301]_  = ~A166 & \new_[7300]_ ;
  assign \new_[7302]_  = \new_[7301]_  & \new_[7296]_ ;
  assign \new_[7305]_  = ~A265 & ~A203;
  assign \new_[7309]_  = ~A299 & ~A298;
  assign \new_[7310]_  = A266 & \new_[7309]_ ;
  assign \new_[7311]_  = \new_[7310]_  & \new_[7305]_ ;
  assign \new_[7314]_  = ~A167 & ~A169;
  assign \new_[7318]_  = ~A201 & ~A200;
  assign \new_[7319]_  = ~A166 & \new_[7318]_ ;
  assign \new_[7320]_  = \new_[7319]_  & \new_[7314]_ ;
  assign \new_[7323]_  = A266 & ~A265;
  assign \new_[7327]_  = ~A302 & ~A301;
  assign \new_[7328]_  = A298 & \new_[7327]_ ;
  assign \new_[7329]_  = \new_[7328]_  & \new_[7323]_ ;
  assign \new_[7332]_  = ~A167 & ~A169;
  assign \new_[7336]_  = ~A200 & ~A199;
  assign \new_[7337]_  = ~A166 & \new_[7336]_ ;
  assign \new_[7338]_  = \new_[7337]_  & \new_[7332]_ ;
  assign \new_[7341]_  = A266 & ~A265;
  assign \new_[7345]_  = ~A302 & ~A301;
  assign \new_[7346]_  = A298 & \new_[7345]_ ;
  assign \new_[7347]_  = \new_[7346]_  & \new_[7341]_ ;
  assign \new_[7350]_  = ~A168 & ~A169;
  assign \new_[7354]_  = A199 & A166;
  assign \new_[7355]_  = A167 & \new_[7354]_ ;
  assign \new_[7356]_  = \new_[7355]_  & \new_[7350]_ ;
  assign \new_[7359]_  = ~A265 & A200;
  assign \new_[7363]_  = ~A300 & A298;
  assign \new_[7364]_  = A266 & \new_[7363]_ ;
  assign \new_[7365]_  = \new_[7364]_  & \new_[7359]_ ;
  assign \new_[7368]_  = ~A168 & ~A169;
  assign \new_[7372]_  = A199 & A166;
  assign \new_[7373]_  = A167 & \new_[7372]_ ;
  assign \new_[7374]_  = \new_[7373]_  & \new_[7368]_ ;
  assign \new_[7377]_  = ~A265 & A200;
  assign \new_[7381]_  = A299 & A298;
  assign \new_[7382]_  = A266 & \new_[7381]_ ;
  assign \new_[7383]_  = \new_[7382]_  & \new_[7377]_ ;
  assign \new_[7386]_  = ~A168 & ~A169;
  assign \new_[7390]_  = A199 & A166;
  assign \new_[7391]_  = A167 & \new_[7390]_ ;
  assign \new_[7392]_  = \new_[7391]_  & \new_[7386]_ ;
  assign \new_[7395]_  = ~A265 & A200;
  assign \new_[7399]_  = ~A299 & ~A298;
  assign \new_[7400]_  = A266 & \new_[7399]_ ;
  assign \new_[7401]_  = \new_[7400]_  & \new_[7395]_ ;
  assign \new_[7404]_  = ~A168 & ~A169;
  assign \new_[7408]_  = ~A199 & A166;
  assign \new_[7409]_  = A167 & \new_[7408]_ ;
  assign \new_[7410]_  = \new_[7409]_  & \new_[7404]_ ;
  assign \new_[7413]_  = A265 & A200;
  assign \new_[7417]_  = A299 & ~A298;
  assign \new_[7418]_  = A266 & \new_[7417]_ ;
  assign \new_[7419]_  = \new_[7418]_  & \new_[7413]_ ;
  assign \new_[7422]_  = ~A168 & ~A169;
  assign \new_[7426]_  = ~A199 & A166;
  assign \new_[7427]_  = A167 & \new_[7426]_ ;
  assign \new_[7428]_  = \new_[7427]_  & \new_[7422]_ ;
  assign \new_[7431]_  = ~A266 & A200;
  assign \new_[7435]_  = A299 & ~A298;
  assign \new_[7436]_  = ~A267 & \new_[7435]_ ;
  assign \new_[7437]_  = \new_[7436]_  & \new_[7431]_ ;
  assign \new_[7440]_  = ~A168 & ~A169;
  assign \new_[7444]_  = ~A199 & A166;
  assign \new_[7445]_  = A167 & \new_[7444]_ ;
  assign \new_[7446]_  = \new_[7445]_  & \new_[7440]_ ;
  assign \new_[7449]_  = ~A265 & A200;
  assign \new_[7453]_  = A299 & ~A298;
  assign \new_[7454]_  = ~A266 & \new_[7453]_ ;
  assign \new_[7455]_  = \new_[7454]_  & \new_[7449]_ ;
  assign \new_[7458]_  = ~A168 & ~A169;
  assign \new_[7462]_  = ~A200 & A166;
  assign \new_[7463]_  = A167 & \new_[7462]_ ;
  assign \new_[7464]_  = \new_[7463]_  & \new_[7458]_ ;
  assign \new_[7467]_  = ~A265 & ~A201;
  assign \new_[7471]_  = ~A300 & A298;
  assign \new_[7472]_  = A266 & \new_[7471]_ ;
  assign \new_[7473]_  = \new_[7472]_  & \new_[7467]_ ;
  assign \new_[7476]_  = ~A168 & ~A169;
  assign \new_[7480]_  = ~A200 & A166;
  assign \new_[7481]_  = A167 & \new_[7480]_ ;
  assign \new_[7482]_  = \new_[7481]_  & \new_[7476]_ ;
  assign \new_[7485]_  = ~A265 & ~A201;
  assign \new_[7489]_  = A299 & A298;
  assign \new_[7490]_  = A266 & \new_[7489]_ ;
  assign \new_[7491]_  = \new_[7490]_  & \new_[7485]_ ;
  assign \new_[7494]_  = ~A168 & ~A169;
  assign \new_[7498]_  = ~A200 & A166;
  assign \new_[7499]_  = A167 & \new_[7498]_ ;
  assign \new_[7500]_  = \new_[7499]_  & \new_[7494]_ ;
  assign \new_[7503]_  = ~A265 & ~A201;
  assign \new_[7507]_  = ~A299 & ~A298;
  assign \new_[7508]_  = A266 & \new_[7507]_ ;
  assign \new_[7509]_  = \new_[7508]_  & \new_[7503]_ ;
  assign \new_[7512]_  = ~A168 & ~A169;
  assign \new_[7516]_  = ~A199 & A166;
  assign \new_[7517]_  = A167 & \new_[7516]_ ;
  assign \new_[7518]_  = \new_[7517]_  & \new_[7512]_ ;
  assign \new_[7521]_  = ~A265 & ~A200;
  assign \new_[7525]_  = ~A300 & A298;
  assign \new_[7526]_  = A266 & \new_[7525]_ ;
  assign \new_[7527]_  = \new_[7526]_  & \new_[7521]_ ;
  assign \new_[7530]_  = ~A168 & ~A169;
  assign \new_[7534]_  = ~A199 & A166;
  assign \new_[7535]_  = A167 & \new_[7534]_ ;
  assign \new_[7536]_  = \new_[7535]_  & \new_[7530]_ ;
  assign \new_[7539]_  = ~A265 & ~A200;
  assign \new_[7543]_  = A299 & A298;
  assign \new_[7544]_  = A266 & \new_[7543]_ ;
  assign \new_[7545]_  = \new_[7544]_  & \new_[7539]_ ;
  assign \new_[7548]_  = ~A168 & ~A169;
  assign \new_[7552]_  = ~A199 & A166;
  assign \new_[7553]_  = A167 & \new_[7552]_ ;
  assign \new_[7554]_  = \new_[7553]_  & \new_[7548]_ ;
  assign \new_[7557]_  = ~A265 & ~A200;
  assign \new_[7561]_  = ~A299 & ~A298;
  assign \new_[7562]_  = A266 & \new_[7561]_ ;
  assign \new_[7563]_  = \new_[7562]_  & \new_[7557]_ ;
  assign \new_[7566]_  = ~A169 & A170;
  assign \new_[7570]_  = A199 & ~A166;
  assign \new_[7571]_  = A167 & \new_[7570]_ ;
  assign \new_[7572]_  = \new_[7571]_  & \new_[7566]_ ;
  assign \new_[7575]_  = A265 & A200;
  assign \new_[7579]_  = A299 & ~A298;
  assign \new_[7580]_  = A266 & \new_[7579]_ ;
  assign \new_[7581]_  = \new_[7580]_  & \new_[7575]_ ;
  assign \new_[7584]_  = ~A169 & A170;
  assign \new_[7588]_  = A199 & ~A166;
  assign \new_[7589]_  = A167 & \new_[7588]_ ;
  assign \new_[7590]_  = \new_[7589]_  & \new_[7584]_ ;
  assign \new_[7593]_  = ~A266 & A200;
  assign \new_[7597]_  = A299 & ~A298;
  assign \new_[7598]_  = ~A267 & \new_[7597]_ ;
  assign \new_[7599]_  = \new_[7598]_  & \new_[7593]_ ;
  assign \new_[7602]_  = ~A169 & A170;
  assign \new_[7606]_  = A199 & ~A166;
  assign \new_[7607]_  = A167 & \new_[7606]_ ;
  assign \new_[7608]_  = \new_[7607]_  & \new_[7602]_ ;
  assign \new_[7611]_  = ~A265 & A200;
  assign \new_[7615]_  = A299 & ~A298;
  assign \new_[7616]_  = ~A266 & \new_[7615]_ ;
  assign \new_[7617]_  = \new_[7616]_  & \new_[7611]_ ;
  assign \new_[7620]_  = ~A169 & A170;
  assign \new_[7624]_  = ~A199 & ~A166;
  assign \new_[7625]_  = A167 & \new_[7624]_ ;
  assign \new_[7626]_  = \new_[7625]_  & \new_[7620]_ ;
  assign \new_[7629]_  = ~A265 & A200;
  assign \new_[7633]_  = ~A300 & A298;
  assign \new_[7634]_  = A266 & \new_[7633]_ ;
  assign \new_[7635]_  = \new_[7634]_  & \new_[7629]_ ;
  assign \new_[7638]_  = ~A169 & A170;
  assign \new_[7642]_  = ~A199 & ~A166;
  assign \new_[7643]_  = A167 & \new_[7642]_ ;
  assign \new_[7644]_  = \new_[7643]_  & \new_[7638]_ ;
  assign \new_[7647]_  = ~A265 & A200;
  assign \new_[7651]_  = A299 & A298;
  assign \new_[7652]_  = A266 & \new_[7651]_ ;
  assign \new_[7653]_  = \new_[7652]_  & \new_[7647]_ ;
  assign \new_[7656]_  = ~A169 & A170;
  assign \new_[7660]_  = ~A199 & ~A166;
  assign \new_[7661]_  = A167 & \new_[7660]_ ;
  assign \new_[7662]_  = \new_[7661]_  & \new_[7656]_ ;
  assign \new_[7665]_  = ~A265 & A200;
  assign \new_[7669]_  = ~A299 & ~A298;
  assign \new_[7670]_  = A266 & \new_[7669]_ ;
  assign \new_[7671]_  = \new_[7670]_  & \new_[7665]_ ;
  assign \new_[7674]_  = ~A169 & A170;
  assign \new_[7678]_  = ~A200 & ~A166;
  assign \new_[7679]_  = A167 & \new_[7678]_ ;
  assign \new_[7680]_  = \new_[7679]_  & \new_[7674]_ ;
  assign \new_[7683]_  = A265 & ~A201;
  assign \new_[7687]_  = A299 & ~A298;
  assign \new_[7688]_  = A266 & \new_[7687]_ ;
  assign \new_[7689]_  = \new_[7688]_  & \new_[7683]_ ;
  assign \new_[7692]_  = ~A169 & A170;
  assign \new_[7696]_  = ~A200 & ~A166;
  assign \new_[7697]_  = A167 & \new_[7696]_ ;
  assign \new_[7698]_  = \new_[7697]_  & \new_[7692]_ ;
  assign \new_[7701]_  = ~A266 & ~A201;
  assign \new_[7705]_  = A299 & ~A298;
  assign \new_[7706]_  = ~A267 & \new_[7705]_ ;
  assign \new_[7707]_  = \new_[7706]_  & \new_[7701]_ ;
  assign \new_[7710]_  = ~A169 & A170;
  assign \new_[7714]_  = ~A200 & ~A166;
  assign \new_[7715]_  = A167 & \new_[7714]_ ;
  assign \new_[7716]_  = \new_[7715]_  & \new_[7710]_ ;
  assign \new_[7719]_  = ~A265 & ~A201;
  assign \new_[7723]_  = A299 & ~A298;
  assign \new_[7724]_  = ~A266 & \new_[7723]_ ;
  assign \new_[7725]_  = \new_[7724]_  & \new_[7719]_ ;
  assign \new_[7728]_  = ~A169 & A170;
  assign \new_[7732]_  = ~A199 & ~A166;
  assign \new_[7733]_  = A167 & \new_[7732]_ ;
  assign \new_[7734]_  = \new_[7733]_  & \new_[7728]_ ;
  assign \new_[7737]_  = A265 & ~A200;
  assign \new_[7741]_  = A299 & ~A298;
  assign \new_[7742]_  = A266 & \new_[7741]_ ;
  assign \new_[7743]_  = \new_[7742]_  & \new_[7737]_ ;
  assign \new_[7746]_  = ~A169 & A170;
  assign \new_[7750]_  = ~A199 & ~A166;
  assign \new_[7751]_  = A167 & \new_[7750]_ ;
  assign \new_[7752]_  = \new_[7751]_  & \new_[7746]_ ;
  assign \new_[7755]_  = ~A266 & ~A200;
  assign \new_[7759]_  = A299 & ~A298;
  assign \new_[7760]_  = ~A267 & \new_[7759]_ ;
  assign \new_[7761]_  = \new_[7760]_  & \new_[7755]_ ;
  assign \new_[7764]_  = ~A169 & A170;
  assign \new_[7768]_  = ~A199 & ~A166;
  assign \new_[7769]_  = A167 & \new_[7768]_ ;
  assign \new_[7770]_  = \new_[7769]_  & \new_[7764]_ ;
  assign \new_[7773]_  = ~A265 & ~A200;
  assign \new_[7777]_  = A299 & ~A298;
  assign \new_[7778]_  = ~A266 & \new_[7777]_ ;
  assign \new_[7779]_  = \new_[7778]_  & \new_[7773]_ ;
  assign \new_[7782]_  = ~A169 & A170;
  assign \new_[7786]_  = A199 & A166;
  assign \new_[7787]_  = ~A167 & \new_[7786]_ ;
  assign \new_[7788]_  = \new_[7787]_  & \new_[7782]_ ;
  assign \new_[7791]_  = A265 & A200;
  assign \new_[7795]_  = A299 & ~A298;
  assign \new_[7796]_  = A266 & \new_[7795]_ ;
  assign \new_[7797]_  = \new_[7796]_  & \new_[7791]_ ;
  assign \new_[7800]_  = ~A169 & A170;
  assign \new_[7804]_  = A199 & A166;
  assign \new_[7805]_  = ~A167 & \new_[7804]_ ;
  assign \new_[7806]_  = \new_[7805]_  & \new_[7800]_ ;
  assign \new_[7809]_  = ~A266 & A200;
  assign \new_[7813]_  = A299 & ~A298;
  assign \new_[7814]_  = ~A267 & \new_[7813]_ ;
  assign \new_[7815]_  = \new_[7814]_  & \new_[7809]_ ;
  assign \new_[7818]_  = ~A169 & A170;
  assign \new_[7822]_  = A199 & A166;
  assign \new_[7823]_  = ~A167 & \new_[7822]_ ;
  assign \new_[7824]_  = \new_[7823]_  & \new_[7818]_ ;
  assign \new_[7827]_  = ~A265 & A200;
  assign \new_[7831]_  = A299 & ~A298;
  assign \new_[7832]_  = ~A266 & \new_[7831]_ ;
  assign \new_[7833]_  = \new_[7832]_  & \new_[7827]_ ;
  assign \new_[7836]_  = ~A169 & A170;
  assign \new_[7840]_  = ~A199 & A166;
  assign \new_[7841]_  = ~A167 & \new_[7840]_ ;
  assign \new_[7842]_  = \new_[7841]_  & \new_[7836]_ ;
  assign \new_[7845]_  = ~A265 & A200;
  assign \new_[7849]_  = ~A300 & A298;
  assign \new_[7850]_  = A266 & \new_[7849]_ ;
  assign \new_[7851]_  = \new_[7850]_  & \new_[7845]_ ;
  assign \new_[7854]_  = ~A169 & A170;
  assign \new_[7858]_  = ~A199 & A166;
  assign \new_[7859]_  = ~A167 & \new_[7858]_ ;
  assign \new_[7860]_  = \new_[7859]_  & \new_[7854]_ ;
  assign \new_[7863]_  = ~A265 & A200;
  assign \new_[7867]_  = A299 & A298;
  assign \new_[7868]_  = A266 & \new_[7867]_ ;
  assign \new_[7869]_  = \new_[7868]_  & \new_[7863]_ ;
  assign \new_[7872]_  = ~A169 & A170;
  assign \new_[7876]_  = ~A199 & A166;
  assign \new_[7877]_  = ~A167 & \new_[7876]_ ;
  assign \new_[7878]_  = \new_[7877]_  & \new_[7872]_ ;
  assign \new_[7881]_  = ~A265 & A200;
  assign \new_[7885]_  = ~A299 & ~A298;
  assign \new_[7886]_  = A266 & \new_[7885]_ ;
  assign \new_[7887]_  = \new_[7886]_  & \new_[7881]_ ;
  assign \new_[7890]_  = ~A169 & A170;
  assign \new_[7894]_  = ~A200 & A166;
  assign \new_[7895]_  = ~A167 & \new_[7894]_ ;
  assign \new_[7896]_  = \new_[7895]_  & \new_[7890]_ ;
  assign \new_[7899]_  = A265 & ~A201;
  assign \new_[7903]_  = A299 & ~A298;
  assign \new_[7904]_  = A266 & \new_[7903]_ ;
  assign \new_[7905]_  = \new_[7904]_  & \new_[7899]_ ;
  assign \new_[7908]_  = ~A169 & A170;
  assign \new_[7912]_  = ~A200 & A166;
  assign \new_[7913]_  = ~A167 & \new_[7912]_ ;
  assign \new_[7914]_  = \new_[7913]_  & \new_[7908]_ ;
  assign \new_[7917]_  = ~A266 & ~A201;
  assign \new_[7921]_  = A299 & ~A298;
  assign \new_[7922]_  = ~A267 & \new_[7921]_ ;
  assign \new_[7923]_  = \new_[7922]_  & \new_[7917]_ ;
  assign \new_[7926]_  = ~A169 & A170;
  assign \new_[7930]_  = ~A200 & A166;
  assign \new_[7931]_  = ~A167 & \new_[7930]_ ;
  assign \new_[7932]_  = \new_[7931]_  & \new_[7926]_ ;
  assign \new_[7935]_  = ~A265 & ~A201;
  assign \new_[7939]_  = A299 & ~A298;
  assign \new_[7940]_  = ~A266 & \new_[7939]_ ;
  assign \new_[7941]_  = \new_[7940]_  & \new_[7935]_ ;
  assign \new_[7944]_  = ~A169 & A170;
  assign \new_[7948]_  = ~A199 & A166;
  assign \new_[7949]_  = ~A167 & \new_[7948]_ ;
  assign \new_[7950]_  = \new_[7949]_  & \new_[7944]_ ;
  assign \new_[7953]_  = A265 & ~A200;
  assign \new_[7957]_  = A299 & ~A298;
  assign \new_[7958]_  = A266 & \new_[7957]_ ;
  assign \new_[7959]_  = \new_[7958]_  & \new_[7953]_ ;
  assign \new_[7962]_  = ~A169 & A170;
  assign \new_[7966]_  = ~A199 & A166;
  assign \new_[7967]_  = ~A167 & \new_[7966]_ ;
  assign \new_[7968]_  = \new_[7967]_  & \new_[7962]_ ;
  assign \new_[7971]_  = ~A266 & ~A200;
  assign \new_[7975]_  = A299 & ~A298;
  assign \new_[7976]_  = ~A267 & \new_[7975]_ ;
  assign \new_[7977]_  = \new_[7976]_  & \new_[7971]_ ;
  assign \new_[7980]_  = ~A169 & A170;
  assign \new_[7984]_  = ~A199 & A166;
  assign \new_[7985]_  = ~A167 & \new_[7984]_ ;
  assign \new_[7986]_  = \new_[7985]_  & \new_[7980]_ ;
  assign \new_[7989]_  = ~A265 & ~A200;
  assign \new_[7993]_  = A299 & ~A298;
  assign \new_[7994]_  = ~A266 & \new_[7993]_ ;
  assign \new_[7995]_  = \new_[7994]_  & \new_[7989]_ ;
  assign \new_[7998]_  = ~A169 & ~A170;
  assign \new_[8002]_  = A200 & A199;
  assign \new_[8003]_  = ~A168 & \new_[8002]_ ;
  assign \new_[8004]_  = \new_[8003]_  & \new_[7998]_ ;
  assign \new_[8007]_  = A266 & ~A265;
  assign \new_[8011]_  = ~A302 & ~A301;
  assign \new_[8012]_  = A298 & \new_[8011]_ ;
  assign \new_[8013]_  = \new_[8012]_  & \new_[8007]_ ;
  assign \new_[8016]_  = ~A169 & ~A170;
  assign \new_[8020]_  = A200 & ~A199;
  assign \new_[8021]_  = ~A168 & \new_[8020]_ ;
  assign \new_[8022]_  = \new_[8021]_  & \new_[8016]_ ;
  assign \new_[8025]_  = ~A268 & ~A266;
  assign \new_[8029]_  = A299 & ~A298;
  assign \new_[8030]_  = ~A269 & \new_[8029]_ ;
  assign \new_[8031]_  = \new_[8030]_  & \new_[8025]_ ;
  assign \new_[8034]_  = ~A169 & ~A170;
  assign \new_[8038]_  = ~A202 & ~A200;
  assign \new_[8039]_  = ~A168 & \new_[8038]_ ;
  assign \new_[8040]_  = \new_[8039]_  & \new_[8034]_ ;
  assign \new_[8043]_  = ~A265 & ~A203;
  assign \new_[8047]_  = ~A300 & A298;
  assign \new_[8048]_  = A266 & \new_[8047]_ ;
  assign \new_[8049]_  = \new_[8048]_  & \new_[8043]_ ;
  assign \new_[8052]_  = ~A169 & ~A170;
  assign \new_[8056]_  = ~A202 & ~A200;
  assign \new_[8057]_  = ~A168 & \new_[8056]_ ;
  assign \new_[8058]_  = \new_[8057]_  & \new_[8052]_ ;
  assign \new_[8061]_  = ~A265 & ~A203;
  assign \new_[8065]_  = A299 & A298;
  assign \new_[8066]_  = A266 & \new_[8065]_ ;
  assign \new_[8067]_  = \new_[8066]_  & \new_[8061]_ ;
  assign \new_[8070]_  = ~A169 & ~A170;
  assign \new_[8074]_  = ~A202 & ~A200;
  assign \new_[8075]_  = ~A168 & \new_[8074]_ ;
  assign \new_[8076]_  = \new_[8075]_  & \new_[8070]_ ;
  assign \new_[8079]_  = ~A265 & ~A203;
  assign \new_[8083]_  = ~A299 & ~A298;
  assign \new_[8084]_  = A266 & \new_[8083]_ ;
  assign \new_[8085]_  = \new_[8084]_  & \new_[8079]_ ;
  assign \new_[8088]_  = ~A169 & ~A170;
  assign \new_[8092]_  = ~A201 & ~A200;
  assign \new_[8093]_  = ~A168 & \new_[8092]_ ;
  assign \new_[8094]_  = \new_[8093]_  & \new_[8088]_ ;
  assign \new_[8097]_  = A266 & ~A265;
  assign \new_[8101]_  = ~A302 & ~A301;
  assign \new_[8102]_  = A298 & \new_[8101]_ ;
  assign \new_[8103]_  = \new_[8102]_  & \new_[8097]_ ;
  assign \new_[8106]_  = ~A169 & ~A170;
  assign \new_[8110]_  = ~A200 & ~A199;
  assign \new_[8111]_  = ~A168 & \new_[8110]_ ;
  assign \new_[8112]_  = \new_[8111]_  & \new_[8106]_ ;
  assign \new_[8115]_  = A266 & ~A265;
  assign \new_[8119]_  = ~A302 & ~A301;
  assign \new_[8120]_  = A298 & \new_[8119]_ ;
  assign \new_[8121]_  = \new_[8120]_  & \new_[8115]_ ;
  assign \new_[8124]_  = A166 & A168;
  assign \new_[8128]_  = ~A266 & A200;
  assign \new_[8129]_  = A199 & \new_[8128]_ ;
  assign \new_[8130]_  = \new_[8129]_  & \new_[8124]_ ;
  assign \new_[8134]_  = A298 & ~A269;
  assign \new_[8135]_  = ~A268 & \new_[8134]_ ;
  assign \new_[8139]_  = A301 & A300;
  assign \new_[8140]_  = ~A299 & \new_[8139]_ ;
  assign \new_[8141]_  = \new_[8140]_  & \new_[8135]_ ;
  assign \new_[8144]_  = A166 & A168;
  assign \new_[8148]_  = ~A266 & A200;
  assign \new_[8149]_  = A199 & \new_[8148]_ ;
  assign \new_[8150]_  = \new_[8149]_  & \new_[8144]_ ;
  assign \new_[8154]_  = A298 & ~A269;
  assign \new_[8155]_  = ~A268 & \new_[8154]_ ;
  assign \new_[8159]_  = A302 & A300;
  assign \new_[8160]_  = ~A299 & \new_[8159]_ ;
  assign \new_[8161]_  = \new_[8160]_  & \new_[8155]_ ;
  assign \new_[8164]_  = A166 & A168;
  assign \new_[8168]_  = A265 & A200;
  assign \new_[8169]_  = ~A199 & \new_[8168]_ ;
  assign \new_[8170]_  = \new_[8169]_  & \new_[8164]_ ;
  assign \new_[8174]_  = A268 & A267;
  assign \new_[8175]_  = ~A266 & \new_[8174]_ ;
  assign \new_[8179]_  = ~A302 & ~A301;
  assign \new_[8180]_  = A298 & \new_[8179]_ ;
  assign \new_[8181]_  = \new_[8180]_  & \new_[8175]_ ;
  assign \new_[8184]_  = A166 & A168;
  assign \new_[8188]_  = A265 & A200;
  assign \new_[8189]_  = ~A199 & \new_[8188]_ ;
  assign \new_[8190]_  = \new_[8189]_  & \new_[8184]_ ;
  assign \new_[8194]_  = A269 & A267;
  assign \new_[8195]_  = ~A266 & \new_[8194]_ ;
  assign \new_[8199]_  = ~A302 & ~A301;
  assign \new_[8200]_  = A298 & \new_[8199]_ ;
  assign \new_[8201]_  = \new_[8200]_  & \new_[8195]_ ;
  assign \new_[8204]_  = A166 & A168;
  assign \new_[8208]_  = ~A203 & ~A202;
  assign \new_[8209]_  = ~A200 & \new_[8208]_ ;
  assign \new_[8210]_  = \new_[8209]_  & \new_[8204]_ ;
  assign \new_[8214]_  = A298 & A266;
  assign \new_[8215]_  = A265 & \new_[8214]_ ;
  assign \new_[8219]_  = A301 & A300;
  assign \new_[8220]_  = ~A299 & \new_[8219]_ ;
  assign \new_[8221]_  = \new_[8220]_  & \new_[8215]_ ;
  assign \new_[8224]_  = A166 & A168;
  assign \new_[8228]_  = ~A203 & ~A202;
  assign \new_[8229]_  = ~A200 & \new_[8228]_ ;
  assign \new_[8230]_  = \new_[8229]_  & \new_[8224]_ ;
  assign \new_[8234]_  = A298 & A266;
  assign \new_[8235]_  = A265 & \new_[8234]_ ;
  assign \new_[8239]_  = A302 & A300;
  assign \new_[8240]_  = ~A299 & \new_[8239]_ ;
  assign \new_[8241]_  = \new_[8240]_  & \new_[8235]_ ;
  assign \new_[8244]_  = A166 & A168;
  assign \new_[8248]_  = ~A203 & ~A202;
  assign \new_[8249]_  = ~A200 & \new_[8248]_ ;
  assign \new_[8250]_  = \new_[8249]_  & \new_[8244]_ ;
  assign \new_[8254]_  = A298 & ~A267;
  assign \new_[8255]_  = ~A266 & \new_[8254]_ ;
  assign \new_[8259]_  = A301 & A300;
  assign \new_[8260]_  = ~A299 & \new_[8259]_ ;
  assign \new_[8261]_  = \new_[8260]_  & \new_[8255]_ ;
  assign \new_[8264]_  = A166 & A168;
  assign \new_[8268]_  = ~A203 & ~A202;
  assign \new_[8269]_  = ~A200 & \new_[8268]_ ;
  assign \new_[8270]_  = \new_[8269]_  & \new_[8264]_ ;
  assign \new_[8274]_  = A298 & ~A267;
  assign \new_[8275]_  = ~A266 & \new_[8274]_ ;
  assign \new_[8279]_  = A302 & A300;
  assign \new_[8280]_  = ~A299 & \new_[8279]_ ;
  assign \new_[8281]_  = \new_[8280]_  & \new_[8275]_ ;
  assign \new_[8284]_  = A166 & A168;
  assign \new_[8288]_  = ~A203 & ~A202;
  assign \new_[8289]_  = ~A200 & \new_[8288]_ ;
  assign \new_[8290]_  = \new_[8289]_  & \new_[8284]_ ;
  assign \new_[8294]_  = A298 & ~A266;
  assign \new_[8295]_  = ~A265 & \new_[8294]_ ;
  assign \new_[8299]_  = A301 & A300;
  assign \new_[8300]_  = ~A299 & \new_[8299]_ ;
  assign \new_[8301]_  = \new_[8300]_  & \new_[8295]_ ;
  assign \new_[8304]_  = A166 & A168;
  assign \new_[8308]_  = ~A203 & ~A202;
  assign \new_[8309]_  = ~A200 & \new_[8308]_ ;
  assign \new_[8310]_  = \new_[8309]_  & \new_[8304]_ ;
  assign \new_[8314]_  = A298 & ~A266;
  assign \new_[8315]_  = ~A265 & \new_[8314]_ ;
  assign \new_[8319]_  = A302 & A300;
  assign \new_[8320]_  = ~A299 & \new_[8319]_ ;
  assign \new_[8321]_  = \new_[8320]_  & \new_[8315]_ ;
  assign \new_[8324]_  = A166 & A168;
  assign \new_[8328]_  = ~A266 & ~A201;
  assign \new_[8329]_  = ~A200 & \new_[8328]_ ;
  assign \new_[8330]_  = \new_[8329]_  & \new_[8324]_ ;
  assign \new_[8334]_  = A298 & ~A269;
  assign \new_[8335]_  = ~A268 & \new_[8334]_ ;
  assign \new_[8339]_  = A301 & A300;
  assign \new_[8340]_  = ~A299 & \new_[8339]_ ;
  assign \new_[8341]_  = \new_[8340]_  & \new_[8335]_ ;
  assign \new_[8344]_  = A166 & A168;
  assign \new_[8348]_  = ~A266 & ~A201;
  assign \new_[8349]_  = ~A200 & \new_[8348]_ ;
  assign \new_[8350]_  = \new_[8349]_  & \new_[8344]_ ;
  assign \new_[8354]_  = A298 & ~A269;
  assign \new_[8355]_  = ~A268 & \new_[8354]_ ;
  assign \new_[8359]_  = A302 & A300;
  assign \new_[8360]_  = ~A299 & \new_[8359]_ ;
  assign \new_[8361]_  = \new_[8360]_  & \new_[8355]_ ;
  assign \new_[8364]_  = A166 & A168;
  assign \new_[8368]_  = A201 & ~A200;
  assign \new_[8369]_  = A199 & \new_[8368]_ ;
  assign \new_[8370]_  = \new_[8369]_  & \new_[8364]_ ;
  assign \new_[8374]_  = A266 & ~A265;
  assign \new_[8375]_  = A202 & \new_[8374]_ ;
  assign \new_[8379]_  = ~A302 & ~A301;
  assign \new_[8380]_  = A298 & \new_[8379]_ ;
  assign \new_[8381]_  = \new_[8380]_  & \new_[8375]_ ;
  assign \new_[8384]_  = A166 & A168;
  assign \new_[8388]_  = A201 & ~A200;
  assign \new_[8389]_  = A199 & \new_[8388]_ ;
  assign \new_[8390]_  = \new_[8389]_  & \new_[8384]_ ;
  assign \new_[8394]_  = A266 & ~A265;
  assign \new_[8395]_  = A203 & \new_[8394]_ ;
  assign \new_[8399]_  = ~A302 & ~A301;
  assign \new_[8400]_  = A298 & \new_[8399]_ ;
  assign \new_[8401]_  = \new_[8400]_  & \new_[8395]_ ;
  assign \new_[8404]_  = A166 & A168;
  assign \new_[8408]_  = ~A266 & ~A200;
  assign \new_[8409]_  = ~A199 & \new_[8408]_ ;
  assign \new_[8410]_  = \new_[8409]_  & \new_[8404]_ ;
  assign \new_[8414]_  = A298 & ~A269;
  assign \new_[8415]_  = ~A268 & \new_[8414]_ ;
  assign \new_[8419]_  = A301 & A300;
  assign \new_[8420]_  = ~A299 & \new_[8419]_ ;
  assign \new_[8421]_  = \new_[8420]_  & \new_[8415]_ ;
  assign \new_[8424]_  = A166 & A168;
  assign \new_[8428]_  = ~A266 & ~A200;
  assign \new_[8429]_  = ~A199 & \new_[8428]_ ;
  assign \new_[8430]_  = \new_[8429]_  & \new_[8424]_ ;
  assign \new_[8434]_  = A298 & ~A269;
  assign \new_[8435]_  = ~A268 & \new_[8434]_ ;
  assign \new_[8439]_  = A302 & A300;
  assign \new_[8440]_  = ~A299 & \new_[8439]_ ;
  assign \new_[8441]_  = \new_[8440]_  & \new_[8435]_ ;
  assign \new_[8444]_  = A167 & A168;
  assign \new_[8448]_  = ~A266 & A200;
  assign \new_[8449]_  = A199 & \new_[8448]_ ;
  assign \new_[8450]_  = \new_[8449]_  & \new_[8444]_ ;
  assign \new_[8454]_  = A298 & ~A269;
  assign \new_[8455]_  = ~A268 & \new_[8454]_ ;
  assign \new_[8459]_  = A301 & A300;
  assign \new_[8460]_  = ~A299 & \new_[8459]_ ;
  assign \new_[8461]_  = \new_[8460]_  & \new_[8455]_ ;
  assign \new_[8464]_  = A167 & A168;
  assign \new_[8468]_  = ~A266 & A200;
  assign \new_[8469]_  = A199 & \new_[8468]_ ;
  assign \new_[8470]_  = \new_[8469]_  & \new_[8464]_ ;
  assign \new_[8474]_  = A298 & ~A269;
  assign \new_[8475]_  = ~A268 & \new_[8474]_ ;
  assign \new_[8479]_  = A302 & A300;
  assign \new_[8480]_  = ~A299 & \new_[8479]_ ;
  assign \new_[8481]_  = \new_[8480]_  & \new_[8475]_ ;
  assign \new_[8484]_  = A167 & A168;
  assign \new_[8488]_  = A265 & A200;
  assign \new_[8489]_  = ~A199 & \new_[8488]_ ;
  assign \new_[8490]_  = \new_[8489]_  & \new_[8484]_ ;
  assign \new_[8494]_  = A268 & A267;
  assign \new_[8495]_  = ~A266 & \new_[8494]_ ;
  assign \new_[8499]_  = ~A302 & ~A301;
  assign \new_[8500]_  = A298 & \new_[8499]_ ;
  assign \new_[8501]_  = \new_[8500]_  & \new_[8495]_ ;
  assign \new_[8504]_  = A167 & A168;
  assign \new_[8508]_  = A265 & A200;
  assign \new_[8509]_  = ~A199 & \new_[8508]_ ;
  assign \new_[8510]_  = \new_[8509]_  & \new_[8504]_ ;
  assign \new_[8514]_  = A269 & A267;
  assign \new_[8515]_  = ~A266 & \new_[8514]_ ;
  assign \new_[8519]_  = ~A302 & ~A301;
  assign \new_[8520]_  = A298 & \new_[8519]_ ;
  assign \new_[8521]_  = \new_[8520]_  & \new_[8515]_ ;
  assign \new_[8524]_  = A167 & A168;
  assign \new_[8528]_  = ~A203 & ~A202;
  assign \new_[8529]_  = ~A200 & \new_[8528]_ ;
  assign \new_[8530]_  = \new_[8529]_  & \new_[8524]_ ;
  assign \new_[8534]_  = A298 & A266;
  assign \new_[8535]_  = A265 & \new_[8534]_ ;
  assign \new_[8539]_  = A301 & A300;
  assign \new_[8540]_  = ~A299 & \new_[8539]_ ;
  assign \new_[8541]_  = \new_[8540]_  & \new_[8535]_ ;
  assign \new_[8544]_  = A167 & A168;
  assign \new_[8548]_  = ~A203 & ~A202;
  assign \new_[8549]_  = ~A200 & \new_[8548]_ ;
  assign \new_[8550]_  = \new_[8549]_  & \new_[8544]_ ;
  assign \new_[8554]_  = A298 & A266;
  assign \new_[8555]_  = A265 & \new_[8554]_ ;
  assign \new_[8559]_  = A302 & A300;
  assign \new_[8560]_  = ~A299 & \new_[8559]_ ;
  assign \new_[8561]_  = \new_[8560]_  & \new_[8555]_ ;
  assign \new_[8564]_  = A167 & A168;
  assign \new_[8568]_  = ~A203 & ~A202;
  assign \new_[8569]_  = ~A200 & \new_[8568]_ ;
  assign \new_[8570]_  = \new_[8569]_  & \new_[8564]_ ;
  assign \new_[8574]_  = A298 & ~A267;
  assign \new_[8575]_  = ~A266 & \new_[8574]_ ;
  assign \new_[8579]_  = A301 & A300;
  assign \new_[8580]_  = ~A299 & \new_[8579]_ ;
  assign \new_[8581]_  = \new_[8580]_  & \new_[8575]_ ;
  assign \new_[8584]_  = A167 & A168;
  assign \new_[8588]_  = ~A203 & ~A202;
  assign \new_[8589]_  = ~A200 & \new_[8588]_ ;
  assign \new_[8590]_  = \new_[8589]_  & \new_[8584]_ ;
  assign \new_[8594]_  = A298 & ~A267;
  assign \new_[8595]_  = ~A266 & \new_[8594]_ ;
  assign \new_[8599]_  = A302 & A300;
  assign \new_[8600]_  = ~A299 & \new_[8599]_ ;
  assign \new_[8601]_  = \new_[8600]_  & \new_[8595]_ ;
  assign \new_[8604]_  = A167 & A168;
  assign \new_[8608]_  = ~A203 & ~A202;
  assign \new_[8609]_  = ~A200 & \new_[8608]_ ;
  assign \new_[8610]_  = \new_[8609]_  & \new_[8604]_ ;
  assign \new_[8614]_  = A298 & ~A266;
  assign \new_[8615]_  = ~A265 & \new_[8614]_ ;
  assign \new_[8619]_  = A301 & A300;
  assign \new_[8620]_  = ~A299 & \new_[8619]_ ;
  assign \new_[8621]_  = \new_[8620]_  & \new_[8615]_ ;
  assign \new_[8624]_  = A167 & A168;
  assign \new_[8628]_  = ~A203 & ~A202;
  assign \new_[8629]_  = ~A200 & \new_[8628]_ ;
  assign \new_[8630]_  = \new_[8629]_  & \new_[8624]_ ;
  assign \new_[8634]_  = A298 & ~A266;
  assign \new_[8635]_  = ~A265 & \new_[8634]_ ;
  assign \new_[8639]_  = A302 & A300;
  assign \new_[8640]_  = ~A299 & \new_[8639]_ ;
  assign \new_[8641]_  = \new_[8640]_  & \new_[8635]_ ;
  assign \new_[8644]_  = A167 & A168;
  assign \new_[8648]_  = ~A266 & ~A201;
  assign \new_[8649]_  = ~A200 & \new_[8648]_ ;
  assign \new_[8650]_  = \new_[8649]_  & \new_[8644]_ ;
  assign \new_[8654]_  = A298 & ~A269;
  assign \new_[8655]_  = ~A268 & \new_[8654]_ ;
  assign \new_[8659]_  = A301 & A300;
  assign \new_[8660]_  = ~A299 & \new_[8659]_ ;
  assign \new_[8661]_  = \new_[8660]_  & \new_[8655]_ ;
  assign \new_[8664]_  = A167 & A168;
  assign \new_[8668]_  = ~A266 & ~A201;
  assign \new_[8669]_  = ~A200 & \new_[8668]_ ;
  assign \new_[8670]_  = \new_[8669]_  & \new_[8664]_ ;
  assign \new_[8674]_  = A298 & ~A269;
  assign \new_[8675]_  = ~A268 & \new_[8674]_ ;
  assign \new_[8679]_  = A302 & A300;
  assign \new_[8680]_  = ~A299 & \new_[8679]_ ;
  assign \new_[8681]_  = \new_[8680]_  & \new_[8675]_ ;
  assign \new_[8684]_  = A167 & A168;
  assign \new_[8688]_  = A201 & ~A200;
  assign \new_[8689]_  = A199 & \new_[8688]_ ;
  assign \new_[8690]_  = \new_[8689]_  & \new_[8684]_ ;
  assign \new_[8694]_  = A266 & ~A265;
  assign \new_[8695]_  = A202 & \new_[8694]_ ;
  assign \new_[8699]_  = ~A302 & ~A301;
  assign \new_[8700]_  = A298 & \new_[8699]_ ;
  assign \new_[8701]_  = \new_[8700]_  & \new_[8695]_ ;
  assign \new_[8704]_  = A167 & A168;
  assign \new_[8708]_  = A201 & ~A200;
  assign \new_[8709]_  = A199 & \new_[8708]_ ;
  assign \new_[8710]_  = \new_[8709]_  & \new_[8704]_ ;
  assign \new_[8714]_  = A266 & ~A265;
  assign \new_[8715]_  = A203 & \new_[8714]_ ;
  assign \new_[8719]_  = ~A302 & ~A301;
  assign \new_[8720]_  = A298 & \new_[8719]_ ;
  assign \new_[8721]_  = \new_[8720]_  & \new_[8715]_ ;
  assign \new_[8724]_  = A167 & A168;
  assign \new_[8728]_  = ~A266 & ~A200;
  assign \new_[8729]_  = ~A199 & \new_[8728]_ ;
  assign \new_[8730]_  = \new_[8729]_  & \new_[8724]_ ;
  assign \new_[8734]_  = A298 & ~A269;
  assign \new_[8735]_  = ~A268 & \new_[8734]_ ;
  assign \new_[8739]_  = A301 & A300;
  assign \new_[8740]_  = ~A299 & \new_[8739]_ ;
  assign \new_[8741]_  = \new_[8740]_  & \new_[8735]_ ;
  assign \new_[8744]_  = A167 & A168;
  assign \new_[8748]_  = ~A266 & ~A200;
  assign \new_[8749]_  = ~A199 & \new_[8748]_ ;
  assign \new_[8750]_  = \new_[8749]_  & \new_[8744]_ ;
  assign \new_[8754]_  = A298 & ~A269;
  assign \new_[8755]_  = ~A268 & \new_[8754]_ ;
  assign \new_[8759]_  = A302 & A300;
  assign \new_[8760]_  = ~A299 & \new_[8759]_ ;
  assign \new_[8761]_  = \new_[8760]_  & \new_[8755]_ ;
  assign \new_[8764]_  = ~A167 & A170;
  assign \new_[8768]_  = A200 & A199;
  assign \new_[8769]_  = ~A166 & \new_[8768]_ ;
  assign \new_[8770]_  = \new_[8769]_  & \new_[8764]_ ;
  assign \new_[8774]_  = A267 & ~A266;
  assign \new_[8775]_  = A265 & \new_[8774]_ ;
  assign \new_[8779]_  = ~A300 & A298;
  assign \new_[8780]_  = A268 & \new_[8779]_ ;
  assign \new_[8781]_  = \new_[8780]_  & \new_[8775]_ ;
  assign \new_[8784]_  = ~A167 & A170;
  assign \new_[8788]_  = A200 & A199;
  assign \new_[8789]_  = ~A166 & \new_[8788]_ ;
  assign \new_[8790]_  = \new_[8789]_  & \new_[8784]_ ;
  assign \new_[8794]_  = A267 & ~A266;
  assign \new_[8795]_  = A265 & \new_[8794]_ ;
  assign \new_[8799]_  = A299 & A298;
  assign \new_[8800]_  = A268 & \new_[8799]_ ;
  assign \new_[8801]_  = \new_[8800]_  & \new_[8795]_ ;
  assign \new_[8804]_  = ~A167 & A170;
  assign \new_[8808]_  = A200 & A199;
  assign \new_[8809]_  = ~A166 & \new_[8808]_ ;
  assign \new_[8810]_  = \new_[8809]_  & \new_[8804]_ ;
  assign \new_[8814]_  = A267 & ~A266;
  assign \new_[8815]_  = A265 & \new_[8814]_ ;
  assign \new_[8819]_  = ~A299 & ~A298;
  assign \new_[8820]_  = A268 & \new_[8819]_ ;
  assign \new_[8821]_  = \new_[8820]_  & \new_[8815]_ ;
  assign \new_[8824]_  = ~A167 & A170;
  assign \new_[8828]_  = A200 & A199;
  assign \new_[8829]_  = ~A166 & \new_[8828]_ ;
  assign \new_[8830]_  = \new_[8829]_  & \new_[8824]_ ;
  assign \new_[8834]_  = A267 & ~A266;
  assign \new_[8835]_  = A265 & \new_[8834]_ ;
  assign \new_[8839]_  = ~A300 & A298;
  assign \new_[8840]_  = A269 & \new_[8839]_ ;
  assign \new_[8841]_  = \new_[8840]_  & \new_[8835]_ ;
  assign \new_[8844]_  = ~A167 & A170;
  assign \new_[8848]_  = A200 & A199;
  assign \new_[8849]_  = ~A166 & \new_[8848]_ ;
  assign \new_[8850]_  = \new_[8849]_  & \new_[8844]_ ;
  assign \new_[8854]_  = A267 & ~A266;
  assign \new_[8855]_  = A265 & \new_[8854]_ ;
  assign \new_[8859]_  = A299 & A298;
  assign \new_[8860]_  = A269 & \new_[8859]_ ;
  assign \new_[8861]_  = \new_[8860]_  & \new_[8855]_ ;
  assign \new_[8864]_  = ~A167 & A170;
  assign \new_[8868]_  = A200 & A199;
  assign \new_[8869]_  = ~A166 & \new_[8868]_ ;
  assign \new_[8870]_  = \new_[8869]_  & \new_[8864]_ ;
  assign \new_[8874]_  = A267 & ~A266;
  assign \new_[8875]_  = A265 & \new_[8874]_ ;
  assign \new_[8879]_  = ~A299 & ~A298;
  assign \new_[8880]_  = A269 & \new_[8879]_ ;
  assign \new_[8881]_  = \new_[8880]_  & \new_[8875]_ ;
  assign \new_[8884]_  = ~A167 & A170;
  assign \new_[8888]_  = A200 & ~A199;
  assign \new_[8889]_  = ~A166 & \new_[8888]_ ;
  assign \new_[8890]_  = \new_[8889]_  & \new_[8884]_ ;
  assign \new_[8894]_  = A298 & A266;
  assign \new_[8895]_  = A265 & \new_[8894]_ ;
  assign \new_[8899]_  = A301 & A300;
  assign \new_[8900]_  = ~A299 & \new_[8899]_ ;
  assign \new_[8901]_  = \new_[8900]_  & \new_[8895]_ ;
  assign \new_[8904]_  = ~A167 & A170;
  assign \new_[8908]_  = A200 & ~A199;
  assign \new_[8909]_  = ~A166 & \new_[8908]_ ;
  assign \new_[8910]_  = \new_[8909]_  & \new_[8904]_ ;
  assign \new_[8914]_  = A298 & A266;
  assign \new_[8915]_  = A265 & \new_[8914]_ ;
  assign \new_[8919]_  = A302 & A300;
  assign \new_[8920]_  = ~A299 & \new_[8919]_ ;
  assign \new_[8921]_  = \new_[8920]_  & \new_[8915]_ ;
  assign \new_[8924]_  = ~A167 & A170;
  assign \new_[8928]_  = A200 & ~A199;
  assign \new_[8929]_  = ~A166 & \new_[8928]_ ;
  assign \new_[8930]_  = \new_[8929]_  & \new_[8924]_ ;
  assign \new_[8934]_  = A298 & ~A267;
  assign \new_[8935]_  = ~A266 & \new_[8934]_ ;
  assign \new_[8939]_  = A301 & A300;
  assign \new_[8940]_  = ~A299 & \new_[8939]_ ;
  assign \new_[8941]_  = \new_[8940]_  & \new_[8935]_ ;
  assign \new_[8944]_  = ~A167 & A170;
  assign \new_[8948]_  = A200 & ~A199;
  assign \new_[8949]_  = ~A166 & \new_[8948]_ ;
  assign \new_[8950]_  = \new_[8949]_  & \new_[8944]_ ;
  assign \new_[8954]_  = A298 & ~A267;
  assign \new_[8955]_  = ~A266 & \new_[8954]_ ;
  assign \new_[8959]_  = A302 & A300;
  assign \new_[8960]_  = ~A299 & \new_[8959]_ ;
  assign \new_[8961]_  = \new_[8960]_  & \new_[8955]_ ;
  assign \new_[8964]_  = ~A167 & A170;
  assign \new_[8968]_  = A200 & ~A199;
  assign \new_[8969]_  = ~A166 & \new_[8968]_ ;
  assign \new_[8970]_  = \new_[8969]_  & \new_[8964]_ ;
  assign \new_[8974]_  = A298 & ~A266;
  assign \new_[8975]_  = ~A265 & \new_[8974]_ ;
  assign \new_[8979]_  = A301 & A300;
  assign \new_[8980]_  = ~A299 & \new_[8979]_ ;
  assign \new_[8981]_  = \new_[8980]_  & \new_[8975]_ ;
  assign \new_[8984]_  = ~A167 & A170;
  assign \new_[8988]_  = A200 & ~A199;
  assign \new_[8989]_  = ~A166 & \new_[8988]_ ;
  assign \new_[8990]_  = \new_[8989]_  & \new_[8984]_ ;
  assign \new_[8994]_  = A298 & ~A266;
  assign \new_[8995]_  = ~A265 & \new_[8994]_ ;
  assign \new_[8999]_  = A302 & A300;
  assign \new_[9000]_  = ~A299 & \new_[8999]_ ;
  assign \new_[9001]_  = \new_[9000]_  & \new_[8995]_ ;
  assign \new_[9004]_  = ~A167 & A170;
  assign \new_[9008]_  = ~A202 & ~A200;
  assign \new_[9009]_  = ~A166 & \new_[9008]_ ;
  assign \new_[9010]_  = \new_[9009]_  & \new_[9004]_ ;
  assign \new_[9014]_  = A266 & ~A265;
  assign \new_[9015]_  = ~A203 & \new_[9014]_ ;
  assign \new_[9019]_  = ~A302 & ~A301;
  assign \new_[9020]_  = A298 & \new_[9019]_ ;
  assign \new_[9021]_  = \new_[9020]_  & \new_[9015]_ ;
  assign \new_[9024]_  = ~A167 & A170;
  assign \new_[9028]_  = ~A201 & ~A200;
  assign \new_[9029]_  = ~A166 & \new_[9028]_ ;
  assign \new_[9030]_  = \new_[9029]_  & \new_[9024]_ ;
  assign \new_[9034]_  = A267 & ~A266;
  assign \new_[9035]_  = A265 & \new_[9034]_ ;
  assign \new_[9039]_  = ~A300 & A298;
  assign \new_[9040]_  = A268 & \new_[9039]_ ;
  assign \new_[9041]_  = \new_[9040]_  & \new_[9035]_ ;
  assign \new_[9044]_  = ~A167 & A170;
  assign \new_[9048]_  = ~A201 & ~A200;
  assign \new_[9049]_  = ~A166 & \new_[9048]_ ;
  assign \new_[9050]_  = \new_[9049]_  & \new_[9044]_ ;
  assign \new_[9054]_  = A267 & ~A266;
  assign \new_[9055]_  = A265 & \new_[9054]_ ;
  assign \new_[9059]_  = A299 & A298;
  assign \new_[9060]_  = A268 & \new_[9059]_ ;
  assign \new_[9061]_  = \new_[9060]_  & \new_[9055]_ ;
  assign \new_[9064]_  = ~A167 & A170;
  assign \new_[9068]_  = ~A201 & ~A200;
  assign \new_[9069]_  = ~A166 & \new_[9068]_ ;
  assign \new_[9070]_  = \new_[9069]_  & \new_[9064]_ ;
  assign \new_[9074]_  = A267 & ~A266;
  assign \new_[9075]_  = A265 & \new_[9074]_ ;
  assign \new_[9079]_  = ~A299 & ~A298;
  assign \new_[9080]_  = A268 & \new_[9079]_ ;
  assign \new_[9081]_  = \new_[9080]_  & \new_[9075]_ ;
  assign \new_[9084]_  = ~A167 & A170;
  assign \new_[9088]_  = ~A201 & ~A200;
  assign \new_[9089]_  = ~A166 & \new_[9088]_ ;
  assign \new_[9090]_  = \new_[9089]_  & \new_[9084]_ ;
  assign \new_[9094]_  = A267 & ~A266;
  assign \new_[9095]_  = A265 & \new_[9094]_ ;
  assign \new_[9099]_  = ~A300 & A298;
  assign \new_[9100]_  = A269 & \new_[9099]_ ;
  assign \new_[9101]_  = \new_[9100]_  & \new_[9095]_ ;
  assign \new_[9104]_  = ~A167 & A170;
  assign \new_[9108]_  = ~A201 & ~A200;
  assign \new_[9109]_  = ~A166 & \new_[9108]_ ;
  assign \new_[9110]_  = \new_[9109]_  & \new_[9104]_ ;
  assign \new_[9114]_  = A267 & ~A266;
  assign \new_[9115]_  = A265 & \new_[9114]_ ;
  assign \new_[9119]_  = A299 & A298;
  assign \new_[9120]_  = A269 & \new_[9119]_ ;
  assign \new_[9121]_  = \new_[9120]_  & \new_[9115]_ ;
  assign \new_[9124]_  = ~A167 & A170;
  assign \new_[9128]_  = ~A201 & ~A200;
  assign \new_[9129]_  = ~A166 & \new_[9128]_ ;
  assign \new_[9130]_  = \new_[9129]_  & \new_[9124]_ ;
  assign \new_[9134]_  = A267 & ~A266;
  assign \new_[9135]_  = A265 & \new_[9134]_ ;
  assign \new_[9139]_  = ~A299 & ~A298;
  assign \new_[9140]_  = A269 & \new_[9139]_ ;
  assign \new_[9141]_  = \new_[9140]_  & \new_[9135]_ ;
  assign \new_[9144]_  = ~A167 & A170;
  assign \new_[9148]_  = ~A200 & A199;
  assign \new_[9149]_  = ~A166 & \new_[9148]_ ;
  assign \new_[9150]_  = \new_[9149]_  & \new_[9144]_ ;
  assign \new_[9154]_  = A265 & A202;
  assign \new_[9155]_  = A201 & \new_[9154]_ ;
  assign \new_[9159]_  = A299 & ~A298;
  assign \new_[9160]_  = A266 & \new_[9159]_ ;
  assign \new_[9161]_  = \new_[9160]_  & \new_[9155]_ ;
  assign \new_[9164]_  = ~A167 & A170;
  assign \new_[9168]_  = ~A200 & A199;
  assign \new_[9169]_  = ~A166 & \new_[9168]_ ;
  assign \new_[9170]_  = \new_[9169]_  & \new_[9164]_ ;
  assign \new_[9174]_  = ~A266 & A202;
  assign \new_[9175]_  = A201 & \new_[9174]_ ;
  assign \new_[9179]_  = A299 & ~A298;
  assign \new_[9180]_  = ~A267 & \new_[9179]_ ;
  assign \new_[9181]_  = \new_[9180]_  & \new_[9175]_ ;
  assign \new_[9184]_  = ~A167 & A170;
  assign \new_[9188]_  = ~A200 & A199;
  assign \new_[9189]_  = ~A166 & \new_[9188]_ ;
  assign \new_[9190]_  = \new_[9189]_  & \new_[9184]_ ;
  assign \new_[9194]_  = ~A265 & A202;
  assign \new_[9195]_  = A201 & \new_[9194]_ ;
  assign \new_[9199]_  = A299 & ~A298;
  assign \new_[9200]_  = ~A266 & \new_[9199]_ ;
  assign \new_[9201]_  = \new_[9200]_  & \new_[9195]_ ;
  assign \new_[9204]_  = ~A167 & A170;
  assign \new_[9208]_  = ~A200 & A199;
  assign \new_[9209]_  = ~A166 & \new_[9208]_ ;
  assign \new_[9210]_  = \new_[9209]_  & \new_[9204]_ ;
  assign \new_[9214]_  = A265 & A203;
  assign \new_[9215]_  = A201 & \new_[9214]_ ;
  assign \new_[9219]_  = A299 & ~A298;
  assign \new_[9220]_  = A266 & \new_[9219]_ ;
  assign \new_[9221]_  = \new_[9220]_  & \new_[9215]_ ;
  assign \new_[9224]_  = ~A167 & A170;
  assign \new_[9228]_  = ~A200 & A199;
  assign \new_[9229]_  = ~A166 & \new_[9228]_ ;
  assign \new_[9230]_  = \new_[9229]_  & \new_[9224]_ ;
  assign \new_[9234]_  = ~A266 & A203;
  assign \new_[9235]_  = A201 & \new_[9234]_ ;
  assign \new_[9239]_  = A299 & ~A298;
  assign \new_[9240]_  = ~A267 & \new_[9239]_ ;
  assign \new_[9241]_  = \new_[9240]_  & \new_[9235]_ ;
  assign \new_[9244]_  = ~A167 & A170;
  assign \new_[9248]_  = ~A200 & A199;
  assign \new_[9249]_  = ~A166 & \new_[9248]_ ;
  assign \new_[9250]_  = \new_[9249]_  & \new_[9244]_ ;
  assign \new_[9254]_  = ~A265 & A203;
  assign \new_[9255]_  = A201 & \new_[9254]_ ;
  assign \new_[9259]_  = A299 & ~A298;
  assign \new_[9260]_  = ~A266 & \new_[9259]_ ;
  assign \new_[9261]_  = \new_[9260]_  & \new_[9255]_ ;
  assign \new_[9264]_  = ~A167 & A170;
  assign \new_[9268]_  = ~A200 & ~A199;
  assign \new_[9269]_  = ~A166 & \new_[9268]_ ;
  assign \new_[9270]_  = \new_[9269]_  & \new_[9264]_ ;
  assign \new_[9274]_  = A267 & ~A266;
  assign \new_[9275]_  = A265 & \new_[9274]_ ;
  assign \new_[9279]_  = ~A300 & A298;
  assign \new_[9280]_  = A268 & \new_[9279]_ ;
  assign \new_[9281]_  = \new_[9280]_  & \new_[9275]_ ;
  assign \new_[9284]_  = ~A167 & A170;
  assign \new_[9288]_  = ~A200 & ~A199;
  assign \new_[9289]_  = ~A166 & \new_[9288]_ ;
  assign \new_[9290]_  = \new_[9289]_  & \new_[9284]_ ;
  assign \new_[9294]_  = A267 & ~A266;
  assign \new_[9295]_  = A265 & \new_[9294]_ ;
  assign \new_[9299]_  = A299 & A298;
  assign \new_[9300]_  = A268 & \new_[9299]_ ;
  assign \new_[9301]_  = \new_[9300]_  & \new_[9295]_ ;
  assign \new_[9304]_  = ~A167 & A170;
  assign \new_[9308]_  = ~A200 & ~A199;
  assign \new_[9309]_  = ~A166 & \new_[9308]_ ;
  assign \new_[9310]_  = \new_[9309]_  & \new_[9304]_ ;
  assign \new_[9314]_  = A267 & ~A266;
  assign \new_[9315]_  = A265 & \new_[9314]_ ;
  assign \new_[9319]_  = ~A299 & ~A298;
  assign \new_[9320]_  = A268 & \new_[9319]_ ;
  assign \new_[9321]_  = \new_[9320]_  & \new_[9315]_ ;
  assign \new_[9324]_  = ~A167 & A170;
  assign \new_[9328]_  = ~A200 & ~A199;
  assign \new_[9329]_  = ~A166 & \new_[9328]_ ;
  assign \new_[9330]_  = \new_[9329]_  & \new_[9324]_ ;
  assign \new_[9334]_  = A267 & ~A266;
  assign \new_[9335]_  = A265 & \new_[9334]_ ;
  assign \new_[9339]_  = ~A300 & A298;
  assign \new_[9340]_  = A269 & \new_[9339]_ ;
  assign \new_[9341]_  = \new_[9340]_  & \new_[9335]_ ;
  assign \new_[9344]_  = ~A167 & A170;
  assign \new_[9348]_  = ~A200 & ~A199;
  assign \new_[9349]_  = ~A166 & \new_[9348]_ ;
  assign \new_[9350]_  = \new_[9349]_  & \new_[9344]_ ;
  assign \new_[9354]_  = A267 & ~A266;
  assign \new_[9355]_  = A265 & \new_[9354]_ ;
  assign \new_[9359]_  = A299 & A298;
  assign \new_[9360]_  = A269 & \new_[9359]_ ;
  assign \new_[9361]_  = \new_[9360]_  & \new_[9355]_ ;
  assign \new_[9364]_  = ~A167 & A170;
  assign \new_[9368]_  = ~A200 & ~A199;
  assign \new_[9369]_  = ~A166 & \new_[9368]_ ;
  assign \new_[9370]_  = \new_[9369]_  & \new_[9364]_ ;
  assign \new_[9374]_  = A267 & ~A266;
  assign \new_[9375]_  = A265 & \new_[9374]_ ;
  assign \new_[9379]_  = ~A299 & ~A298;
  assign \new_[9380]_  = A269 & \new_[9379]_ ;
  assign \new_[9381]_  = \new_[9380]_  & \new_[9375]_ ;
  assign \new_[9384]_  = ~A168 & A169;
  assign \new_[9388]_  = A199 & ~A166;
  assign \new_[9389]_  = A167 & \new_[9388]_ ;
  assign \new_[9390]_  = \new_[9389]_  & \new_[9384]_ ;
  assign \new_[9394]_  = A266 & ~A265;
  assign \new_[9395]_  = A200 & \new_[9394]_ ;
  assign \new_[9399]_  = ~A302 & ~A301;
  assign \new_[9400]_  = A298 & \new_[9399]_ ;
  assign \new_[9401]_  = \new_[9400]_  & \new_[9395]_ ;
  assign \new_[9404]_  = ~A168 & A169;
  assign \new_[9408]_  = ~A199 & ~A166;
  assign \new_[9409]_  = A167 & \new_[9408]_ ;
  assign \new_[9410]_  = \new_[9409]_  & \new_[9404]_ ;
  assign \new_[9414]_  = ~A268 & ~A266;
  assign \new_[9415]_  = A200 & \new_[9414]_ ;
  assign \new_[9419]_  = A299 & ~A298;
  assign \new_[9420]_  = ~A269 & \new_[9419]_ ;
  assign \new_[9421]_  = \new_[9420]_  & \new_[9415]_ ;
  assign \new_[9424]_  = ~A168 & A169;
  assign \new_[9428]_  = ~A200 & ~A166;
  assign \new_[9429]_  = A167 & \new_[9428]_ ;
  assign \new_[9430]_  = \new_[9429]_  & \new_[9424]_ ;
  assign \new_[9434]_  = ~A265 & ~A203;
  assign \new_[9435]_  = ~A202 & \new_[9434]_ ;
  assign \new_[9439]_  = ~A300 & A298;
  assign \new_[9440]_  = A266 & \new_[9439]_ ;
  assign \new_[9441]_  = \new_[9440]_  & \new_[9435]_ ;
  assign \new_[9444]_  = ~A168 & A169;
  assign \new_[9448]_  = ~A200 & ~A166;
  assign \new_[9449]_  = A167 & \new_[9448]_ ;
  assign \new_[9450]_  = \new_[9449]_  & \new_[9444]_ ;
  assign \new_[9454]_  = ~A265 & ~A203;
  assign \new_[9455]_  = ~A202 & \new_[9454]_ ;
  assign \new_[9459]_  = A299 & A298;
  assign \new_[9460]_  = A266 & \new_[9459]_ ;
  assign \new_[9461]_  = \new_[9460]_  & \new_[9455]_ ;
  assign \new_[9464]_  = ~A168 & A169;
  assign \new_[9468]_  = ~A200 & ~A166;
  assign \new_[9469]_  = A167 & \new_[9468]_ ;
  assign \new_[9470]_  = \new_[9469]_  & \new_[9464]_ ;
  assign \new_[9474]_  = ~A265 & ~A203;
  assign \new_[9475]_  = ~A202 & \new_[9474]_ ;
  assign \new_[9479]_  = ~A299 & ~A298;
  assign \new_[9480]_  = A266 & \new_[9479]_ ;
  assign \new_[9481]_  = \new_[9480]_  & \new_[9475]_ ;
  assign \new_[9484]_  = ~A168 & A169;
  assign \new_[9488]_  = ~A200 & ~A166;
  assign \new_[9489]_  = A167 & \new_[9488]_ ;
  assign \new_[9490]_  = \new_[9489]_  & \new_[9484]_ ;
  assign \new_[9494]_  = A266 & ~A265;
  assign \new_[9495]_  = ~A201 & \new_[9494]_ ;
  assign \new_[9499]_  = ~A302 & ~A301;
  assign \new_[9500]_  = A298 & \new_[9499]_ ;
  assign \new_[9501]_  = \new_[9500]_  & \new_[9495]_ ;
  assign \new_[9504]_  = ~A168 & A169;
  assign \new_[9508]_  = ~A199 & ~A166;
  assign \new_[9509]_  = A167 & \new_[9508]_ ;
  assign \new_[9510]_  = \new_[9509]_  & \new_[9504]_ ;
  assign \new_[9514]_  = A266 & ~A265;
  assign \new_[9515]_  = ~A200 & \new_[9514]_ ;
  assign \new_[9519]_  = ~A302 & ~A301;
  assign \new_[9520]_  = A298 & \new_[9519]_ ;
  assign \new_[9521]_  = \new_[9520]_  & \new_[9515]_ ;
  assign \new_[9524]_  = ~A168 & A169;
  assign \new_[9528]_  = A199 & A166;
  assign \new_[9529]_  = ~A167 & \new_[9528]_ ;
  assign \new_[9530]_  = \new_[9529]_  & \new_[9524]_ ;
  assign \new_[9534]_  = A266 & ~A265;
  assign \new_[9535]_  = A200 & \new_[9534]_ ;
  assign \new_[9539]_  = ~A302 & ~A301;
  assign \new_[9540]_  = A298 & \new_[9539]_ ;
  assign \new_[9541]_  = \new_[9540]_  & \new_[9535]_ ;
  assign \new_[9544]_  = ~A168 & A169;
  assign \new_[9548]_  = ~A199 & A166;
  assign \new_[9549]_  = ~A167 & \new_[9548]_ ;
  assign \new_[9550]_  = \new_[9549]_  & \new_[9544]_ ;
  assign \new_[9554]_  = ~A268 & ~A266;
  assign \new_[9555]_  = A200 & \new_[9554]_ ;
  assign \new_[9559]_  = A299 & ~A298;
  assign \new_[9560]_  = ~A269 & \new_[9559]_ ;
  assign \new_[9561]_  = \new_[9560]_  & \new_[9555]_ ;
  assign \new_[9564]_  = ~A168 & A169;
  assign \new_[9568]_  = ~A200 & A166;
  assign \new_[9569]_  = ~A167 & \new_[9568]_ ;
  assign \new_[9570]_  = \new_[9569]_  & \new_[9564]_ ;
  assign \new_[9574]_  = ~A265 & ~A203;
  assign \new_[9575]_  = ~A202 & \new_[9574]_ ;
  assign \new_[9579]_  = ~A300 & A298;
  assign \new_[9580]_  = A266 & \new_[9579]_ ;
  assign \new_[9581]_  = \new_[9580]_  & \new_[9575]_ ;
  assign \new_[9584]_  = ~A168 & A169;
  assign \new_[9588]_  = ~A200 & A166;
  assign \new_[9589]_  = ~A167 & \new_[9588]_ ;
  assign \new_[9590]_  = \new_[9589]_  & \new_[9584]_ ;
  assign \new_[9594]_  = ~A265 & ~A203;
  assign \new_[9595]_  = ~A202 & \new_[9594]_ ;
  assign \new_[9599]_  = A299 & A298;
  assign \new_[9600]_  = A266 & \new_[9599]_ ;
  assign \new_[9601]_  = \new_[9600]_  & \new_[9595]_ ;
  assign \new_[9604]_  = ~A168 & A169;
  assign \new_[9608]_  = ~A200 & A166;
  assign \new_[9609]_  = ~A167 & \new_[9608]_ ;
  assign \new_[9610]_  = \new_[9609]_  & \new_[9604]_ ;
  assign \new_[9614]_  = ~A265 & ~A203;
  assign \new_[9615]_  = ~A202 & \new_[9614]_ ;
  assign \new_[9619]_  = ~A299 & ~A298;
  assign \new_[9620]_  = A266 & \new_[9619]_ ;
  assign \new_[9621]_  = \new_[9620]_  & \new_[9615]_ ;
  assign \new_[9624]_  = ~A168 & A169;
  assign \new_[9628]_  = ~A200 & A166;
  assign \new_[9629]_  = ~A167 & \new_[9628]_ ;
  assign \new_[9630]_  = \new_[9629]_  & \new_[9624]_ ;
  assign \new_[9634]_  = A266 & ~A265;
  assign \new_[9635]_  = ~A201 & \new_[9634]_ ;
  assign \new_[9639]_  = ~A302 & ~A301;
  assign \new_[9640]_  = A298 & \new_[9639]_ ;
  assign \new_[9641]_  = \new_[9640]_  & \new_[9635]_ ;
  assign \new_[9644]_  = ~A168 & A169;
  assign \new_[9648]_  = ~A199 & A166;
  assign \new_[9649]_  = ~A167 & \new_[9648]_ ;
  assign \new_[9650]_  = \new_[9649]_  & \new_[9644]_ ;
  assign \new_[9654]_  = A266 & ~A265;
  assign \new_[9655]_  = ~A200 & \new_[9654]_ ;
  assign \new_[9659]_  = ~A302 & ~A301;
  assign \new_[9660]_  = A298 & \new_[9659]_ ;
  assign \new_[9661]_  = \new_[9660]_  & \new_[9655]_ ;
  assign \new_[9664]_  = A169 & A170;
  assign \new_[9668]_  = A200 & A199;
  assign \new_[9669]_  = ~A168 & \new_[9668]_ ;
  assign \new_[9670]_  = \new_[9669]_  & \new_[9664]_ ;
  assign \new_[9674]_  = A267 & ~A266;
  assign \new_[9675]_  = A265 & \new_[9674]_ ;
  assign \new_[9679]_  = ~A300 & A298;
  assign \new_[9680]_  = A268 & \new_[9679]_ ;
  assign \new_[9681]_  = \new_[9680]_  & \new_[9675]_ ;
  assign \new_[9684]_  = A169 & A170;
  assign \new_[9688]_  = A200 & A199;
  assign \new_[9689]_  = ~A168 & \new_[9688]_ ;
  assign \new_[9690]_  = \new_[9689]_  & \new_[9684]_ ;
  assign \new_[9694]_  = A267 & ~A266;
  assign \new_[9695]_  = A265 & \new_[9694]_ ;
  assign \new_[9699]_  = A299 & A298;
  assign \new_[9700]_  = A268 & \new_[9699]_ ;
  assign \new_[9701]_  = \new_[9700]_  & \new_[9695]_ ;
  assign \new_[9704]_  = A169 & A170;
  assign \new_[9708]_  = A200 & A199;
  assign \new_[9709]_  = ~A168 & \new_[9708]_ ;
  assign \new_[9710]_  = \new_[9709]_  & \new_[9704]_ ;
  assign \new_[9714]_  = A267 & ~A266;
  assign \new_[9715]_  = A265 & \new_[9714]_ ;
  assign \new_[9719]_  = ~A299 & ~A298;
  assign \new_[9720]_  = A268 & \new_[9719]_ ;
  assign \new_[9721]_  = \new_[9720]_  & \new_[9715]_ ;
  assign \new_[9724]_  = A169 & A170;
  assign \new_[9728]_  = A200 & A199;
  assign \new_[9729]_  = ~A168 & \new_[9728]_ ;
  assign \new_[9730]_  = \new_[9729]_  & \new_[9724]_ ;
  assign \new_[9734]_  = A267 & ~A266;
  assign \new_[9735]_  = A265 & \new_[9734]_ ;
  assign \new_[9739]_  = ~A300 & A298;
  assign \new_[9740]_  = A269 & \new_[9739]_ ;
  assign \new_[9741]_  = \new_[9740]_  & \new_[9735]_ ;
  assign \new_[9744]_  = A169 & A170;
  assign \new_[9748]_  = A200 & A199;
  assign \new_[9749]_  = ~A168 & \new_[9748]_ ;
  assign \new_[9750]_  = \new_[9749]_  & \new_[9744]_ ;
  assign \new_[9754]_  = A267 & ~A266;
  assign \new_[9755]_  = A265 & \new_[9754]_ ;
  assign \new_[9759]_  = A299 & A298;
  assign \new_[9760]_  = A269 & \new_[9759]_ ;
  assign \new_[9761]_  = \new_[9760]_  & \new_[9755]_ ;
  assign \new_[9764]_  = A169 & A170;
  assign \new_[9768]_  = A200 & A199;
  assign \new_[9769]_  = ~A168 & \new_[9768]_ ;
  assign \new_[9770]_  = \new_[9769]_  & \new_[9764]_ ;
  assign \new_[9774]_  = A267 & ~A266;
  assign \new_[9775]_  = A265 & \new_[9774]_ ;
  assign \new_[9779]_  = ~A299 & ~A298;
  assign \new_[9780]_  = A269 & \new_[9779]_ ;
  assign \new_[9781]_  = \new_[9780]_  & \new_[9775]_ ;
  assign \new_[9784]_  = A169 & A170;
  assign \new_[9788]_  = A200 & ~A199;
  assign \new_[9789]_  = ~A168 & \new_[9788]_ ;
  assign \new_[9790]_  = \new_[9789]_  & \new_[9784]_ ;
  assign \new_[9794]_  = A298 & A266;
  assign \new_[9795]_  = A265 & \new_[9794]_ ;
  assign \new_[9799]_  = A301 & A300;
  assign \new_[9800]_  = ~A299 & \new_[9799]_ ;
  assign \new_[9801]_  = \new_[9800]_  & \new_[9795]_ ;
  assign \new_[9804]_  = A169 & A170;
  assign \new_[9808]_  = A200 & ~A199;
  assign \new_[9809]_  = ~A168 & \new_[9808]_ ;
  assign \new_[9810]_  = \new_[9809]_  & \new_[9804]_ ;
  assign \new_[9814]_  = A298 & A266;
  assign \new_[9815]_  = A265 & \new_[9814]_ ;
  assign \new_[9819]_  = A302 & A300;
  assign \new_[9820]_  = ~A299 & \new_[9819]_ ;
  assign \new_[9821]_  = \new_[9820]_  & \new_[9815]_ ;
  assign \new_[9824]_  = A169 & A170;
  assign \new_[9828]_  = A200 & ~A199;
  assign \new_[9829]_  = ~A168 & \new_[9828]_ ;
  assign \new_[9830]_  = \new_[9829]_  & \new_[9824]_ ;
  assign \new_[9834]_  = A298 & ~A267;
  assign \new_[9835]_  = ~A266 & \new_[9834]_ ;
  assign \new_[9839]_  = A301 & A300;
  assign \new_[9840]_  = ~A299 & \new_[9839]_ ;
  assign \new_[9841]_  = \new_[9840]_  & \new_[9835]_ ;
  assign \new_[9844]_  = A169 & A170;
  assign \new_[9848]_  = A200 & ~A199;
  assign \new_[9849]_  = ~A168 & \new_[9848]_ ;
  assign \new_[9850]_  = \new_[9849]_  & \new_[9844]_ ;
  assign \new_[9854]_  = A298 & ~A267;
  assign \new_[9855]_  = ~A266 & \new_[9854]_ ;
  assign \new_[9859]_  = A302 & A300;
  assign \new_[9860]_  = ~A299 & \new_[9859]_ ;
  assign \new_[9861]_  = \new_[9860]_  & \new_[9855]_ ;
  assign \new_[9864]_  = A169 & A170;
  assign \new_[9868]_  = A200 & ~A199;
  assign \new_[9869]_  = ~A168 & \new_[9868]_ ;
  assign \new_[9870]_  = \new_[9869]_  & \new_[9864]_ ;
  assign \new_[9874]_  = A298 & ~A266;
  assign \new_[9875]_  = ~A265 & \new_[9874]_ ;
  assign \new_[9879]_  = A301 & A300;
  assign \new_[9880]_  = ~A299 & \new_[9879]_ ;
  assign \new_[9881]_  = \new_[9880]_  & \new_[9875]_ ;
  assign \new_[9884]_  = A169 & A170;
  assign \new_[9888]_  = A200 & ~A199;
  assign \new_[9889]_  = ~A168 & \new_[9888]_ ;
  assign \new_[9890]_  = \new_[9889]_  & \new_[9884]_ ;
  assign \new_[9894]_  = A298 & ~A266;
  assign \new_[9895]_  = ~A265 & \new_[9894]_ ;
  assign \new_[9899]_  = A302 & A300;
  assign \new_[9900]_  = ~A299 & \new_[9899]_ ;
  assign \new_[9901]_  = \new_[9900]_  & \new_[9895]_ ;
  assign \new_[9904]_  = A169 & A170;
  assign \new_[9908]_  = ~A202 & ~A200;
  assign \new_[9909]_  = ~A168 & \new_[9908]_ ;
  assign \new_[9910]_  = \new_[9909]_  & \new_[9904]_ ;
  assign \new_[9914]_  = A266 & ~A265;
  assign \new_[9915]_  = ~A203 & \new_[9914]_ ;
  assign \new_[9919]_  = ~A302 & ~A301;
  assign \new_[9920]_  = A298 & \new_[9919]_ ;
  assign \new_[9921]_  = \new_[9920]_  & \new_[9915]_ ;
  assign \new_[9924]_  = A169 & A170;
  assign \new_[9928]_  = ~A201 & ~A200;
  assign \new_[9929]_  = ~A168 & \new_[9928]_ ;
  assign \new_[9930]_  = \new_[9929]_  & \new_[9924]_ ;
  assign \new_[9934]_  = A267 & ~A266;
  assign \new_[9935]_  = A265 & \new_[9934]_ ;
  assign \new_[9939]_  = ~A300 & A298;
  assign \new_[9940]_  = A268 & \new_[9939]_ ;
  assign \new_[9941]_  = \new_[9940]_  & \new_[9935]_ ;
  assign \new_[9944]_  = A169 & A170;
  assign \new_[9948]_  = ~A201 & ~A200;
  assign \new_[9949]_  = ~A168 & \new_[9948]_ ;
  assign \new_[9950]_  = \new_[9949]_  & \new_[9944]_ ;
  assign \new_[9954]_  = A267 & ~A266;
  assign \new_[9955]_  = A265 & \new_[9954]_ ;
  assign \new_[9959]_  = A299 & A298;
  assign \new_[9960]_  = A268 & \new_[9959]_ ;
  assign \new_[9961]_  = \new_[9960]_  & \new_[9955]_ ;
  assign \new_[9964]_  = A169 & A170;
  assign \new_[9968]_  = ~A201 & ~A200;
  assign \new_[9969]_  = ~A168 & \new_[9968]_ ;
  assign \new_[9970]_  = \new_[9969]_  & \new_[9964]_ ;
  assign \new_[9974]_  = A267 & ~A266;
  assign \new_[9975]_  = A265 & \new_[9974]_ ;
  assign \new_[9979]_  = ~A299 & ~A298;
  assign \new_[9980]_  = A268 & \new_[9979]_ ;
  assign \new_[9981]_  = \new_[9980]_  & \new_[9975]_ ;
  assign \new_[9984]_  = A169 & A170;
  assign \new_[9988]_  = ~A201 & ~A200;
  assign \new_[9989]_  = ~A168 & \new_[9988]_ ;
  assign \new_[9990]_  = \new_[9989]_  & \new_[9984]_ ;
  assign \new_[9994]_  = A267 & ~A266;
  assign \new_[9995]_  = A265 & \new_[9994]_ ;
  assign \new_[9999]_  = ~A300 & A298;
  assign \new_[10000]_  = A269 & \new_[9999]_ ;
  assign \new_[10001]_  = \new_[10000]_  & \new_[9995]_ ;
  assign \new_[10004]_  = A169 & A170;
  assign \new_[10008]_  = ~A201 & ~A200;
  assign \new_[10009]_  = ~A168 & \new_[10008]_ ;
  assign \new_[10010]_  = \new_[10009]_  & \new_[10004]_ ;
  assign \new_[10014]_  = A267 & ~A266;
  assign \new_[10015]_  = A265 & \new_[10014]_ ;
  assign \new_[10019]_  = A299 & A298;
  assign \new_[10020]_  = A269 & \new_[10019]_ ;
  assign \new_[10021]_  = \new_[10020]_  & \new_[10015]_ ;
  assign \new_[10024]_  = A169 & A170;
  assign \new_[10028]_  = ~A201 & ~A200;
  assign \new_[10029]_  = ~A168 & \new_[10028]_ ;
  assign \new_[10030]_  = \new_[10029]_  & \new_[10024]_ ;
  assign \new_[10034]_  = A267 & ~A266;
  assign \new_[10035]_  = A265 & \new_[10034]_ ;
  assign \new_[10039]_  = ~A299 & ~A298;
  assign \new_[10040]_  = A269 & \new_[10039]_ ;
  assign \new_[10041]_  = \new_[10040]_  & \new_[10035]_ ;
  assign \new_[10044]_  = A169 & A170;
  assign \new_[10048]_  = ~A200 & A199;
  assign \new_[10049]_  = ~A168 & \new_[10048]_ ;
  assign \new_[10050]_  = \new_[10049]_  & \new_[10044]_ ;
  assign \new_[10054]_  = A265 & A202;
  assign \new_[10055]_  = A201 & \new_[10054]_ ;
  assign \new_[10059]_  = A299 & ~A298;
  assign \new_[10060]_  = A266 & \new_[10059]_ ;
  assign \new_[10061]_  = \new_[10060]_  & \new_[10055]_ ;
  assign \new_[10064]_  = A169 & A170;
  assign \new_[10068]_  = ~A200 & A199;
  assign \new_[10069]_  = ~A168 & \new_[10068]_ ;
  assign \new_[10070]_  = \new_[10069]_  & \new_[10064]_ ;
  assign \new_[10074]_  = ~A266 & A202;
  assign \new_[10075]_  = A201 & \new_[10074]_ ;
  assign \new_[10079]_  = A299 & ~A298;
  assign \new_[10080]_  = ~A267 & \new_[10079]_ ;
  assign \new_[10081]_  = \new_[10080]_  & \new_[10075]_ ;
  assign \new_[10084]_  = A169 & A170;
  assign \new_[10088]_  = ~A200 & A199;
  assign \new_[10089]_  = ~A168 & \new_[10088]_ ;
  assign \new_[10090]_  = \new_[10089]_  & \new_[10084]_ ;
  assign \new_[10094]_  = ~A265 & A202;
  assign \new_[10095]_  = A201 & \new_[10094]_ ;
  assign \new_[10099]_  = A299 & ~A298;
  assign \new_[10100]_  = ~A266 & \new_[10099]_ ;
  assign \new_[10101]_  = \new_[10100]_  & \new_[10095]_ ;
  assign \new_[10104]_  = A169 & A170;
  assign \new_[10108]_  = ~A200 & A199;
  assign \new_[10109]_  = ~A168 & \new_[10108]_ ;
  assign \new_[10110]_  = \new_[10109]_  & \new_[10104]_ ;
  assign \new_[10114]_  = A265 & A203;
  assign \new_[10115]_  = A201 & \new_[10114]_ ;
  assign \new_[10119]_  = A299 & ~A298;
  assign \new_[10120]_  = A266 & \new_[10119]_ ;
  assign \new_[10121]_  = \new_[10120]_  & \new_[10115]_ ;
  assign \new_[10124]_  = A169 & A170;
  assign \new_[10128]_  = ~A200 & A199;
  assign \new_[10129]_  = ~A168 & \new_[10128]_ ;
  assign \new_[10130]_  = \new_[10129]_  & \new_[10124]_ ;
  assign \new_[10134]_  = ~A266 & A203;
  assign \new_[10135]_  = A201 & \new_[10134]_ ;
  assign \new_[10139]_  = A299 & ~A298;
  assign \new_[10140]_  = ~A267 & \new_[10139]_ ;
  assign \new_[10141]_  = \new_[10140]_  & \new_[10135]_ ;
  assign \new_[10144]_  = A169 & A170;
  assign \new_[10148]_  = ~A200 & A199;
  assign \new_[10149]_  = ~A168 & \new_[10148]_ ;
  assign \new_[10150]_  = \new_[10149]_  & \new_[10144]_ ;
  assign \new_[10154]_  = ~A265 & A203;
  assign \new_[10155]_  = A201 & \new_[10154]_ ;
  assign \new_[10159]_  = A299 & ~A298;
  assign \new_[10160]_  = ~A266 & \new_[10159]_ ;
  assign \new_[10161]_  = \new_[10160]_  & \new_[10155]_ ;
  assign \new_[10164]_  = A169 & A170;
  assign \new_[10168]_  = ~A200 & ~A199;
  assign \new_[10169]_  = ~A168 & \new_[10168]_ ;
  assign \new_[10170]_  = \new_[10169]_  & \new_[10164]_ ;
  assign \new_[10174]_  = A267 & ~A266;
  assign \new_[10175]_  = A265 & \new_[10174]_ ;
  assign \new_[10179]_  = ~A300 & A298;
  assign \new_[10180]_  = A268 & \new_[10179]_ ;
  assign \new_[10181]_  = \new_[10180]_  & \new_[10175]_ ;
  assign \new_[10184]_  = A169 & A170;
  assign \new_[10188]_  = ~A200 & ~A199;
  assign \new_[10189]_  = ~A168 & \new_[10188]_ ;
  assign \new_[10190]_  = \new_[10189]_  & \new_[10184]_ ;
  assign \new_[10194]_  = A267 & ~A266;
  assign \new_[10195]_  = A265 & \new_[10194]_ ;
  assign \new_[10199]_  = A299 & A298;
  assign \new_[10200]_  = A268 & \new_[10199]_ ;
  assign \new_[10201]_  = \new_[10200]_  & \new_[10195]_ ;
  assign \new_[10204]_  = A169 & A170;
  assign \new_[10208]_  = ~A200 & ~A199;
  assign \new_[10209]_  = ~A168 & \new_[10208]_ ;
  assign \new_[10210]_  = \new_[10209]_  & \new_[10204]_ ;
  assign \new_[10214]_  = A267 & ~A266;
  assign \new_[10215]_  = A265 & \new_[10214]_ ;
  assign \new_[10219]_  = ~A299 & ~A298;
  assign \new_[10220]_  = A268 & \new_[10219]_ ;
  assign \new_[10221]_  = \new_[10220]_  & \new_[10215]_ ;
  assign \new_[10224]_  = A169 & A170;
  assign \new_[10228]_  = ~A200 & ~A199;
  assign \new_[10229]_  = ~A168 & \new_[10228]_ ;
  assign \new_[10230]_  = \new_[10229]_  & \new_[10224]_ ;
  assign \new_[10234]_  = A267 & ~A266;
  assign \new_[10235]_  = A265 & \new_[10234]_ ;
  assign \new_[10239]_  = ~A300 & A298;
  assign \new_[10240]_  = A269 & \new_[10239]_ ;
  assign \new_[10241]_  = \new_[10240]_  & \new_[10235]_ ;
  assign \new_[10244]_  = A169 & A170;
  assign \new_[10248]_  = ~A200 & ~A199;
  assign \new_[10249]_  = ~A168 & \new_[10248]_ ;
  assign \new_[10250]_  = \new_[10249]_  & \new_[10244]_ ;
  assign \new_[10254]_  = A267 & ~A266;
  assign \new_[10255]_  = A265 & \new_[10254]_ ;
  assign \new_[10259]_  = A299 & A298;
  assign \new_[10260]_  = A269 & \new_[10259]_ ;
  assign \new_[10261]_  = \new_[10260]_  & \new_[10255]_ ;
  assign \new_[10264]_  = A169 & A170;
  assign \new_[10268]_  = ~A200 & ~A199;
  assign \new_[10269]_  = ~A168 & \new_[10268]_ ;
  assign \new_[10270]_  = \new_[10269]_  & \new_[10264]_ ;
  assign \new_[10274]_  = A267 & ~A266;
  assign \new_[10275]_  = A265 & \new_[10274]_ ;
  assign \new_[10279]_  = ~A299 & ~A298;
  assign \new_[10280]_  = A269 & \new_[10279]_ ;
  assign \new_[10281]_  = \new_[10280]_  & \new_[10275]_ ;
  assign \new_[10284]_  = A169 & ~A170;
  assign \new_[10288]_  = A199 & A166;
  assign \new_[10289]_  = A167 & \new_[10288]_ ;
  assign \new_[10290]_  = \new_[10289]_  & \new_[10284]_ ;
  assign \new_[10294]_  = ~A268 & ~A266;
  assign \new_[10295]_  = A200 & \new_[10294]_ ;
  assign \new_[10299]_  = A299 & ~A298;
  assign \new_[10300]_  = ~A269 & \new_[10299]_ ;
  assign \new_[10301]_  = \new_[10300]_  & \new_[10295]_ ;
  assign \new_[10304]_  = A169 & ~A170;
  assign \new_[10308]_  = ~A199 & A166;
  assign \new_[10309]_  = A167 & \new_[10308]_ ;
  assign \new_[10310]_  = \new_[10309]_  & \new_[10304]_ ;
  assign \new_[10314]_  = A266 & ~A265;
  assign \new_[10315]_  = A200 & \new_[10314]_ ;
  assign \new_[10319]_  = ~A302 & ~A301;
  assign \new_[10320]_  = A298 & \new_[10319]_ ;
  assign \new_[10321]_  = \new_[10320]_  & \new_[10315]_ ;
  assign \new_[10324]_  = A169 & ~A170;
  assign \new_[10328]_  = ~A200 & A166;
  assign \new_[10329]_  = A167 & \new_[10328]_ ;
  assign \new_[10330]_  = \new_[10329]_  & \new_[10324]_ ;
  assign \new_[10334]_  = A265 & ~A203;
  assign \new_[10335]_  = ~A202 & \new_[10334]_ ;
  assign \new_[10339]_  = A299 & ~A298;
  assign \new_[10340]_  = A266 & \new_[10339]_ ;
  assign \new_[10341]_  = \new_[10340]_  & \new_[10335]_ ;
  assign \new_[10344]_  = A169 & ~A170;
  assign \new_[10348]_  = ~A200 & A166;
  assign \new_[10349]_  = A167 & \new_[10348]_ ;
  assign \new_[10350]_  = \new_[10349]_  & \new_[10344]_ ;
  assign \new_[10354]_  = ~A266 & ~A203;
  assign \new_[10355]_  = ~A202 & \new_[10354]_ ;
  assign \new_[10359]_  = A299 & ~A298;
  assign \new_[10360]_  = ~A267 & \new_[10359]_ ;
  assign \new_[10361]_  = \new_[10360]_  & \new_[10355]_ ;
  assign \new_[10364]_  = A169 & ~A170;
  assign \new_[10368]_  = ~A200 & A166;
  assign \new_[10369]_  = A167 & \new_[10368]_ ;
  assign \new_[10370]_  = \new_[10369]_  & \new_[10364]_ ;
  assign \new_[10374]_  = ~A265 & ~A203;
  assign \new_[10375]_  = ~A202 & \new_[10374]_ ;
  assign \new_[10379]_  = A299 & ~A298;
  assign \new_[10380]_  = ~A266 & \new_[10379]_ ;
  assign \new_[10381]_  = \new_[10380]_  & \new_[10375]_ ;
  assign \new_[10384]_  = A169 & ~A170;
  assign \new_[10388]_  = ~A200 & A166;
  assign \new_[10389]_  = A167 & \new_[10388]_ ;
  assign \new_[10390]_  = \new_[10389]_  & \new_[10384]_ ;
  assign \new_[10394]_  = ~A268 & ~A266;
  assign \new_[10395]_  = ~A201 & \new_[10394]_ ;
  assign \new_[10399]_  = A299 & ~A298;
  assign \new_[10400]_  = ~A269 & \new_[10399]_ ;
  assign \new_[10401]_  = \new_[10400]_  & \new_[10395]_ ;
  assign \new_[10404]_  = A169 & ~A170;
  assign \new_[10408]_  = ~A199 & A166;
  assign \new_[10409]_  = A167 & \new_[10408]_ ;
  assign \new_[10410]_  = \new_[10409]_  & \new_[10404]_ ;
  assign \new_[10414]_  = ~A268 & ~A266;
  assign \new_[10415]_  = ~A200 & \new_[10414]_ ;
  assign \new_[10419]_  = A299 & ~A298;
  assign \new_[10420]_  = ~A269 & \new_[10419]_ ;
  assign \new_[10421]_  = \new_[10420]_  & \new_[10415]_ ;
  assign \new_[10424]_  = A169 & ~A170;
  assign \new_[10428]_  = A199 & ~A166;
  assign \new_[10429]_  = ~A167 & \new_[10428]_ ;
  assign \new_[10430]_  = \new_[10429]_  & \new_[10424]_ ;
  assign \new_[10434]_  = ~A268 & ~A266;
  assign \new_[10435]_  = A200 & \new_[10434]_ ;
  assign \new_[10439]_  = A299 & ~A298;
  assign \new_[10440]_  = ~A269 & \new_[10439]_ ;
  assign \new_[10441]_  = \new_[10440]_  & \new_[10435]_ ;
  assign \new_[10444]_  = A169 & ~A170;
  assign \new_[10448]_  = ~A199 & ~A166;
  assign \new_[10449]_  = ~A167 & \new_[10448]_ ;
  assign \new_[10450]_  = \new_[10449]_  & \new_[10444]_ ;
  assign \new_[10454]_  = A266 & ~A265;
  assign \new_[10455]_  = A200 & \new_[10454]_ ;
  assign \new_[10459]_  = ~A302 & ~A301;
  assign \new_[10460]_  = A298 & \new_[10459]_ ;
  assign \new_[10461]_  = \new_[10460]_  & \new_[10455]_ ;
  assign \new_[10464]_  = A169 & ~A170;
  assign \new_[10468]_  = ~A200 & ~A166;
  assign \new_[10469]_  = ~A167 & \new_[10468]_ ;
  assign \new_[10470]_  = \new_[10469]_  & \new_[10464]_ ;
  assign \new_[10474]_  = A265 & ~A203;
  assign \new_[10475]_  = ~A202 & \new_[10474]_ ;
  assign \new_[10479]_  = A299 & ~A298;
  assign \new_[10480]_  = A266 & \new_[10479]_ ;
  assign \new_[10481]_  = \new_[10480]_  & \new_[10475]_ ;
  assign \new_[10484]_  = A169 & ~A170;
  assign \new_[10488]_  = ~A200 & ~A166;
  assign \new_[10489]_  = ~A167 & \new_[10488]_ ;
  assign \new_[10490]_  = \new_[10489]_  & \new_[10484]_ ;
  assign \new_[10494]_  = ~A266 & ~A203;
  assign \new_[10495]_  = ~A202 & \new_[10494]_ ;
  assign \new_[10499]_  = A299 & ~A298;
  assign \new_[10500]_  = ~A267 & \new_[10499]_ ;
  assign \new_[10501]_  = \new_[10500]_  & \new_[10495]_ ;
  assign \new_[10504]_  = A169 & ~A170;
  assign \new_[10508]_  = ~A200 & ~A166;
  assign \new_[10509]_  = ~A167 & \new_[10508]_ ;
  assign \new_[10510]_  = \new_[10509]_  & \new_[10504]_ ;
  assign \new_[10514]_  = ~A265 & ~A203;
  assign \new_[10515]_  = ~A202 & \new_[10514]_ ;
  assign \new_[10519]_  = A299 & ~A298;
  assign \new_[10520]_  = ~A266 & \new_[10519]_ ;
  assign \new_[10521]_  = \new_[10520]_  & \new_[10515]_ ;
  assign \new_[10524]_  = A169 & ~A170;
  assign \new_[10528]_  = ~A200 & ~A166;
  assign \new_[10529]_  = ~A167 & \new_[10528]_ ;
  assign \new_[10530]_  = \new_[10529]_  & \new_[10524]_ ;
  assign \new_[10534]_  = ~A268 & ~A266;
  assign \new_[10535]_  = ~A201 & \new_[10534]_ ;
  assign \new_[10539]_  = A299 & ~A298;
  assign \new_[10540]_  = ~A269 & \new_[10539]_ ;
  assign \new_[10541]_  = \new_[10540]_  & \new_[10535]_ ;
  assign \new_[10544]_  = A169 & ~A170;
  assign \new_[10548]_  = ~A199 & ~A166;
  assign \new_[10549]_  = ~A167 & \new_[10548]_ ;
  assign \new_[10550]_  = \new_[10549]_  & \new_[10544]_ ;
  assign \new_[10554]_  = ~A268 & ~A266;
  assign \new_[10555]_  = ~A200 & \new_[10554]_ ;
  assign \new_[10559]_  = A299 & ~A298;
  assign \new_[10560]_  = ~A269 & \new_[10559]_ ;
  assign \new_[10561]_  = \new_[10560]_  & \new_[10555]_ ;
  assign \new_[10564]_  = ~A167 & ~A169;
  assign \new_[10568]_  = A200 & A199;
  assign \new_[10569]_  = ~A166 & \new_[10568]_ ;
  assign \new_[10570]_  = \new_[10569]_  & \new_[10564]_ ;
  assign \new_[10574]_  = A267 & ~A266;
  assign \new_[10575]_  = A265 & \new_[10574]_ ;
  assign \new_[10579]_  = ~A300 & A298;
  assign \new_[10580]_  = A268 & \new_[10579]_ ;
  assign \new_[10581]_  = \new_[10580]_  & \new_[10575]_ ;
  assign \new_[10584]_  = ~A167 & ~A169;
  assign \new_[10588]_  = A200 & A199;
  assign \new_[10589]_  = ~A166 & \new_[10588]_ ;
  assign \new_[10590]_  = \new_[10589]_  & \new_[10584]_ ;
  assign \new_[10594]_  = A267 & ~A266;
  assign \new_[10595]_  = A265 & \new_[10594]_ ;
  assign \new_[10599]_  = A299 & A298;
  assign \new_[10600]_  = A268 & \new_[10599]_ ;
  assign \new_[10601]_  = \new_[10600]_  & \new_[10595]_ ;
  assign \new_[10604]_  = ~A167 & ~A169;
  assign \new_[10608]_  = A200 & A199;
  assign \new_[10609]_  = ~A166 & \new_[10608]_ ;
  assign \new_[10610]_  = \new_[10609]_  & \new_[10604]_ ;
  assign \new_[10614]_  = A267 & ~A266;
  assign \new_[10615]_  = A265 & \new_[10614]_ ;
  assign \new_[10619]_  = ~A299 & ~A298;
  assign \new_[10620]_  = A268 & \new_[10619]_ ;
  assign \new_[10621]_  = \new_[10620]_  & \new_[10615]_ ;
  assign \new_[10624]_  = ~A167 & ~A169;
  assign \new_[10628]_  = A200 & A199;
  assign \new_[10629]_  = ~A166 & \new_[10628]_ ;
  assign \new_[10630]_  = \new_[10629]_  & \new_[10624]_ ;
  assign \new_[10634]_  = A267 & ~A266;
  assign \new_[10635]_  = A265 & \new_[10634]_ ;
  assign \new_[10639]_  = ~A300 & A298;
  assign \new_[10640]_  = A269 & \new_[10639]_ ;
  assign \new_[10641]_  = \new_[10640]_  & \new_[10635]_ ;
  assign \new_[10644]_  = ~A167 & ~A169;
  assign \new_[10648]_  = A200 & A199;
  assign \new_[10649]_  = ~A166 & \new_[10648]_ ;
  assign \new_[10650]_  = \new_[10649]_  & \new_[10644]_ ;
  assign \new_[10654]_  = A267 & ~A266;
  assign \new_[10655]_  = A265 & \new_[10654]_ ;
  assign \new_[10659]_  = A299 & A298;
  assign \new_[10660]_  = A269 & \new_[10659]_ ;
  assign \new_[10661]_  = \new_[10660]_  & \new_[10655]_ ;
  assign \new_[10664]_  = ~A167 & ~A169;
  assign \new_[10668]_  = A200 & A199;
  assign \new_[10669]_  = ~A166 & \new_[10668]_ ;
  assign \new_[10670]_  = \new_[10669]_  & \new_[10664]_ ;
  assign \new_[10674]_  = A267 & ~A266;
  assign \new_[10675]_  = A265 & \new_[10674]_ ;
  assign \new_[10679]_  = ~A299 & ~A298;
  assign \new_[10680]_  = A269 & \new_[10679]_ ;
  assign \new_[10681]_  = \new_[10680]_  & \new_[10675]_ ;
  assign \new_[10684]_  = ~A167 & ~A169;
  assign \new_[10688]_  = A200 & ~A199;
  assign \new_[10689]_  = ~A166 & \new_[10688]_ ;
  assign \new_[10690]_  = \new_[10689]_  & \new_[10684]_ ;
  assign \new_[10694]_  = A298 & A266;
  assign \new_[10695]_  = A265 & \new_[10694]_ ;
  assign \new_[10699]_  = A301 & A300;
  assign \new_[10700]_  = ~A299 & \new_[10699]_ ;
  assign \new_[10701]_  = \new_[10700]_  & \new_[10695]_ ;
  assign \new_[10704]_  = ~A167 & ~A169;
  assign \new_[10708]_  = A200 & ~A199;
  assign \new_[10709]_  = ~A166 & \new_[10708]_ ;
  assign \new_[10710]_  = \new_[10709]_  & \new_[10704]_ ;
  assign \new_[10714]_  = A298 & A266;
  assign \new_[10715]_  = A265 & \new_[10714]_ ;
  assign \new_[10719]_  = A302 & A300;
  assign \new_[10720]_  = ~A299 & \new_[10719]_ ;
  assign \new_[10721]_  = \new_[10720]_  & \new_[10715]_ ;
  assign \new_[10724]_  = ~A167 & ~A169;
  assign \new_[10728]_  = A200 & ~A199;
  assign \new_[10729]_  = ~A166 & \new_[10728]_ ;
  assign \new_[10730]_  = \new_[10729]_  & \new_[10724]_ ;
  assign \new_[10734]_  = A298 & ~A267;
  assign \new_[10735]_  = ~A266 & \new_[10734]_ ;
  assign \new_[10739]_  = A301 & A300;
  assign \new_[10740]_  = ~A299 & \new_[10739]_ ;
  assign \new_[10741]_  = \new_[10740]_  & \new_[10735]_ ;
  assign \new_[10744]_  = ~A167 & ~A169;
  assign \new_[10748]_  = A200 & ~A199;
  assign \new_[10749]_  = ~A166 & \new_[10748]_ ;
  assign \new_[10750]_  = \new_[10749]_  & \new_[10744]_ ;
  assign \new_[10754]_  = A298 & ~A267;
  assign \new_[10755]_  = ~A266 & \new_[10754]_ ;
  assign \new_[10759]_  = A302 & A300;
  assign \new_[10760]_  = ~A299 & \new_[10759]_ ;
  assign \new_[10761]_  = \new_[10760]_  & \new_[10755]_ ;
  assign \new_[10764]_  = ~A167 & ~A169;
  assign \new_[10768]_  = A200 & ~A199;
  assign \new_[10769]_  = ~A166 & \new_[10768]_ ;
  assign \new_[10770]_  = \new_[10769]_  & \new_[10764]_ ;
  assign \new_[10774]_  = A298 & ~A266;
  assign \new_[10775]_  = ~A265 & \new_[10774]_ ;
  assign \new_[10779]_  = A301 & A300;
  assign \new_[10780]_  = ~A299 & \new_[10779]_ ;
  assign \new_[10781]_  = \new_[10780]_  & \new_[10775]_ ;
  assign \new_[10784]_  = ~A167 & ~A169;
  assign \new_[10788]_  = A200 & ~A199;
  assign \new_[10789]_  = ~A166 & \new_[10788]_ ;
  assign \new_[10790]_  = \new_[10789]_  & \new_[10784]_ ;
  assign \new_[10794]_  = A298 & ~A266;
  assign \new_[10795]_  = ~A265 & \new_[10794]_ ;
  assign \new_[10799]_  = A302 & A300;
  assign \new_[10800]_  = ~A299 & \new_[10799]_ ;
  assign \new_[10801]_  = \new_[10800]_  & \new_[10795]_ ;
  assign \new_[10804]_  = ~A167 & ~A169;
  assign \new_[10808]_  = ~A202 & ~A200;
  assign \new_[10809]_  = ~A166 & \new_[10808]_ ;
  assign \new_[10810]_  = \new_[10809]_  & \new_[10804]_ ;
  assign \new_[10814]_  = A266 & ~A265;
  assign \new_[10815]_  = ~A203 & \new_[10814]_ ;
  assign \new_[10819]_  = ~A302 & ~A301;
  assign \new_[10820]_  = A298 & \new_[10819]_ ;
  assign \new_[10821]_  = \new_[10820]_  & \new_[10815]_ ;
  assign \new_[10824]_  = ~A167 & ~A169;
  assign \new_[10828]_  = ~A201 & ~A200;
  assign \new_[10829]_  = ~A166 & \new_[10828]_ ;
  assign \new_[10830]_  = \new_[10829]_  & \new_[10824]_ ;
  assign \new_[10834]_  = A267 & ~A266;
  assign \new_[10835]_  = A265 & \new_[10834]_ ;
  assign \new_[10839]_  = ~A300 & A298;
  assign \new_[10840]_  = A268 & \new_[10839]_ ;
  assign \new_[10841]_  = \new_[10840]_  & \new_[10835]_ ;
  assign \new_[10844]_  = ~A167 & ~A169;
  assign \new_[10848]_  = ~A201 & ~A200;
  assign \new_[10849]_  = ~A166 & \new_[10848]_ ;
  assign \new_[10850]_  = \new_[10849]_  & \new_[10844]_ ;
  assign \new_[10854]_  = A267 & ~A266;
  assign \new_[10855]_  = A265 & \new_[10854]_ ;
  assign \new_[10859]_  = A299 & A298;
  assign \new_[10860]_  = A268 & \new_[10859]_ ;
  assign \new_[10861]_  = \new_[10860]_  & \new_[10855]_ ;
  assign \new_[10864]_  = ~A167 & ~A169;
  assign \new_[10868]_  = ~A201 & ~A200;
  assign \new_[10869]_  = ~A166 & \new_[10868]_ ;
  assign \new_[10870]_  = \new_[10869]_  & \new_[10864]_ ;
  assign \new_[10874]_  = A267 & ~A266;
  assign \new_[10875]_  = A265 & \new_[10874]_ ;
  assign \new_[10879]_  = ~A299 & ~A298;
  assign \new_[10880]_  = A268 & \new_[10879]_ ;
  assign \new_[10881]_  = \new_[10880]_  & \new_[10875]_ ;
  assign \new_[10884]_  = ~A167 & ~A169;
  assign \new_[10888]_  = ~A201 & ~A200;
  assign \new_[10889]_  = ~A166 & \new_[10888]_ ;
  assign \new_[10890]_  = \new_[10889]_  & \new_[10884]_ ;
  assign \new_[10894]_  = A267 & ~A266;
  assign \new_[10895]_  = A265 & \new_[10894]_ ;
  assign \new_[10899]_  = ~A300 & A298;
  assign \new_[10900]_  = A269 & \new_[10899]_ ;
  assign \new_[10901]_  = \new_[10900]_  & \new_[10895]_ ;
  assign \new_[10904]_  = ~A167 & ~A169;
  assign \new_[10908]_  = ~A201 & ~A200;
  assign \new_[10909]_  = ~A166 & \new_[10908]_ ;
  assign \new_[10910]_  = \new_[10909]_  & \new_[10904]_ ;
  assign \new_[10914]_  = A267 & ~A266;
  assign \new_[10915]_  = A265 & \new_[10914]_ ;
  assign \new_[10919]_  = A299 & A298;
  assign \new_[10920]_  = A269 & \new_[10919]_ ;
  assign \new_[10921]_  = \new_[10920]_  & \new_[10915]_ ;
  assign \new_[10924]_  = ~A167 & ~A169;
  assign \new_[10928]_  = ~A201 & ~A200;
  assign \new_[10929]_  = ~A166 & \new_[10928]_ ;
  assign \new_[10930]_  = \new_[10929]_  & \new_[10924]_ ;
  assign \new_[10934]_  = A267 & ~A266;
  assign \new_[10935]_  = A265 & \new_[10934]_ ;
  assign \new_[10939]_  = ~A299 & ~A298;
  assign \new_[10940]_  = A269 & \new_[10939]_ ;
  assign \new_[10941]_  = \new_[10940]_  & \new_[10935]_ ;
  assign \new_[10944]_  = ~A167 & ~A169;
  assign \new_[10948]_  = ~A200 & A199;
  assign \new_[10949]_  = ~A166 & \new_[10948]_ ;
  assign \new_[10950]_  = \new_[10949]_  & \new_[10944]_ ;
  assign \new_[10954]_  = A265 & A202;
  assign \new_[10955]_  = A201 & \new_[10954]_ ;
  assign \new_[10959]_  = A299 & ~A298;
  assign \new_[10960]_  = A266 & \new_[10959]_ ;
  assign \new_[10961]_  = \new_[10960]_  & \new_[10955]_ ;
  assign \new_[10964]_  = ~A167 & ~A169;
  assign \new_[10968]_  = ~A200 & A199;
  assign \new_[10969]_  = ~A166 & \new_[10968]_ ;
  assign \new_[10970]_  = \new_[10969]_  & \new_[10964]_ ;
  assign \new_[10974]_  = ~A266 & A202;
  assign \new_[10975]_  = A201 & \new_[10974]_ ;
  assign \new_[10979]_  = A299 & ~A298;
  assign \new_[10980]_  = ~A267 & \new_[10979]_ ;
  assign \new_[10981]_  = \new_[10980]_  & \new_[10975]_ ;
  assign \new_[10984]_  = ~A167 & ~A169;
  assign \new_[10988]_  = ~A200 & A199;
  assign \new_[10989]_  = ~A166 & \new_[10988]_ ;
  assign \new_[10990]_  = \new_[10989]_  & \new_[10984]_ ;
  assign \new_[10994]_  = ~A265 & A202;
  assign \new_[10995]_  = A201 & \new_[10994]_ ;
  assign \new_[10999]_  = A299 & ~A298;
  assign \new_[11000]_  = ~A266 & \new_[10999]_ ;
  assign \new_[11001]_  = \new_[11000]_  & \new_[10995]_ ;
  assign \new_[11004]_  = ~A167 & ~A169;
  assign \new_[11008]_  = ~A200 & A199;
  assign \new_[11009]_  = ~A166 & \new_[11008]_ ;
  assign \new_[11010]_  = \new_[11009]_  & \new_[11004]_ ;
  assign \new_[11014]_  = A265 & A203;
  assign \new_[11015]_  = A201 & \new_[11014]_ ;
  assign \new_[11019]_  = A299 & ~A298;
  assign \new_[11020]_  = A266 & \new_[11019]_ ;
  assign \new_[11021]_  = \new_[11020]_  & \new_[11015]_ ;
  assign \new_[11024]_  = ~A167 & ~A169;
  assign \new_[11028]_  = ~A200 & A199;
  assign \new_[11029]_  = ~A166 & \new_[11028]_ ;
  assign \new_[11030]_  = \new_[11029]_  & \new_[11024]_ ;
  assign \new_[11034]_  = ~A266 & A203;
  assign \new_[11035]_  = A201 & \new_[11034]_ ;
  assign \new_[11039]_  = A299 & ~A298;
  assign \new_[11040]_  = ~A267 & \new_[11039]_ ;
  assign \new_[11041]_  = \new_[11040]_  & \new_[11035]_ ;
  assign \new_[11044]_  = ~A167 & ~A169;
  assign \new_[11048]_  = ~A200 & A199;
  assign \new_[11049]_  = ~A166 & \new_[11048]_ ;
  assign \new_[11050]_  = \new_[11049]_  & \new_[11044]_ ;
  assign \new_[11054]_  = ~A265 & A203;
  assign \new_[11055]_  = A201 & \new_[11054]_ ;
  assign \new_[11059]_  = A299 & ~A298;
  assign \new_[11060]_  = ~A266 & \new_[11059]_ ;
  assign \new_[11061]_  = \new_[11060]_  & \new_[11055]_ ;
  assign \new_[11064]_  = ~A167 & ~A169;
  assign \new_[11068]_  = ~A200 & ~A199;
  assign \new_[11069]_  = ~A166 & \new_[11068]_ ;
  assign \new_[11070]_  = \new_[11069]_  & \new_[11064]_ ;
  assign \new_[11074]_  = A267 & ~A266;
  assign \new_[11075]_  = A265 & \new_[11074]_ ;
  assign \new_[11079]_  = ~A300 & A298;
  assign \new_[11080]_  = A268 & \new_[11079]_ ;
  assign \new_[11081]_  = \new_[11080]_  & \new_[11075]_ ;
  assign \new_[11084]_  = ~A167 & ~A169;
  assign \new_[11088]_  = ~A200 & ~A199;
  assign \new_[11089]_  = ~A166 & \new_[11088]_ ;
  assign \new_[11090]_  = \new_[11089]_  & \new_[11084]_ ;
  assign \new_[11094]_  = A267 & ~A266;
  assign \new_[11095]_  = A265 & \new_[11094]_ ;
  assign \new_[11099]_  = A299 & A298;
  assign \new_[11100]_  = A268 & \new_[11099]_ ;
  assign \new_[11101]_  = \new_[11100]_  & \new_[11095]_ ;
  assign \new_[11104]_  = ~A167 & ~A169;
  assign \new_[11108]_  = ~A200 & ~A199;
  assign \new_[11109]_  = ~A166 & \new_[11108]_ ;
  assign \new_[11110]_  = \new_[11109]_  & \new_[11104]_ ;
  assign \new_[11114]_  = A267 & ~A266;
  assign \new_[11115]_  = A265 & \new_[11114]_ ;
  assign \new_[11119]_  = ~A299 & ~A298;
  assign \new_[11120]_  = A268 & \new_[11119]_ ;
  assign \new_[11121]_  = \new_[11120]_  & \new_[11115]_ ;
  assign \new_[11124]_  = ~A167 & ~A169;
  assign \new_[11128]_  = ~A200 & ~A199;
  assign \new_[11129]_  = ~A166 & \new_[11128]_ ;
  assign \new_[11130]_  = \new_[11129]_  & \new_[11124]_ ;
  assign \new_[11134]_  = A267 & ~A266;
  assign \new_[11135]_  = A265 & \new_[11134]_ ;
  assign \new_[11139]_  = ~A300 & A298;
  assign \new_[11140]_  = A269 & \new_[11139]_ ;
  assign \new_[11141]_  = \new_[11140]_  & \new_[11135]_ ;
  assign \new_[11144]_  = ~A167 & ~A169;
  assign \new_[11148]_  = ~A200 & ~A199;
  assign \new_[11149]_  = ~A166 & \new_[11148]_ ;
  assign \new_[11150]_  = \new_[11149]_  & \new_[11144]_ ;
  assign \new_[11154]_  = A267 & ~A266;
  assign \new_[11155]_  = A265 & \new_[11154]_ ;
  assign \new_[11159]_  = A299 & A298;
  assign \new_[11160]_  = A269 & \new_[11159]_ ;
  assign \new_[11161]_  = \new_[11160]_  & \new_[11155]_ ;
  assign \new_[11164]_  = ~A167 & ~A169;
  assign \new_[11168]_  = ~A200 & ~A199;
  assign \new_[11169]_  = ~A166 & \new_[11168]_ ;
  assign \new_[11170]_  = \new_[11169]_  & \new_[11164]_ ;
  assign \new_[11174]_  = A267 & ~A266;
  assign \new_[11175]_  = A265 & \new_[11174]_ ;
  assign \new_[11179]_  = ~A299 & ~A298;
  assign \new_[11180]_  = A269 & \new_[11179]_ ;
  assign \new_[11181]_  = \new_[11180]_  & \new_[11175]_ ;
  assign \new_[11184]_  = ~A168 & ~A169;
  assign \new_[11188]_  = A199 & A166;
  assign \new_[11189]_  = A167 & \new_[11188]_ ;
  assign \new_[11190]_  = \new_[11189]_  & \new_[11184]_ ;
  assign \new_[11194]_  = A266 & ~A265;
  assign \new_[11195]_  = A200 & \new_[11194]_ ;
  assign \new_[11199]_  = ~A302 & ~A301;
  assign \new_[11200]_  = A298 & \new_[11199]_ ;
  assign \new_[11201]_  = \new_[11200]_  & \new_[11195]_ ;
  assign \new_[11204]_  = ~A168 & ~A169;
  assign \new_[11208]_  = ~A199 & A166;
  assign \new_[11209]_  = A167 & \new_[11208]_ ;
  assign \new_[11210]_  = \new_[11209]_  & \new_[11204]_ ;
  assign \new_[11214]_  = ~A268 & ~A266;
  assign \new_[11215]_  = A200 & \new_[11214]_ ;
  assign \new_[11219]_  = A299 & ~A298;
  assign \new_[11220]_  = ~A269 & \new_[11219]_ ;
  assign \new_[11221]_  = \new_[11220]_  & \new_[11215]_ ;
  assign \new_[11224]_  = ~A168 & ~A169;
  assign \new_[11228]_  = ~A200 & A166;
  assign \new_[11229]_  = A167 & \new_[11228]_ ;
  assign \new_[11230]_  = \new_[11229]_  & \new_[11224]_ ;
  assign \new_[11234]_  = ~A265 & ~A203;
  assign \new_[11235]_  = ~A202 & \new_[11234]_ ;
  assign \new_[11239]_  = ~A300 & A298;
  assign \new_[11240]_  = A266 & \new_[11239]_ ;
  assign \new_[11241]_  = \new_[11240]_  & \new_[11235]_ ;
  assign \new_[11244]_  = ~A168 & ~A169;
  assign \new_[11248]_  = ~A200 & A166;
  assign \new_[11249]_  = A167 & \new_[11248]_ ;
  assign \new_[11250]_  = \new_[11249]_  & \new_[11244]_ ;
  assign \new_[11254]_  = ~A265 & ~A203;
  assign \new_[11255]_  = ~A202 & \new_[11254]_ ;
  assign \new_[11259]_  = A299 & A298;
  assign \new_[11260]_  = A266 & \new_[11259]_ ;
  assign \new_[11261]_  = \new_[11260]_  & \new_[11255]_ ;
  assign \new_[11264]_  = ~A168 & ~A169;
  assign \new_[11268]_  = ~A200 & A166;
  assign \new_[11269]_  = A167 & \new_[11268]_ ;
  assign \new_[11270]_  = \new_[11269]_  & \new_[11264]_ ;
  assign \new_[11274]_  = ~A265 & ~A203;
  assign \new_[11275]_  = ~A202 & \new_[11274]_ ;
  assign \new_[11279]_  = ~A299 & ~A298;
  assign \new_[11280]_  = A266 & \new_[11279]_ ;
  assign \new_[11281]_  = \new_[11280]_  & \new_[11275]_ ;
  assign \new_[11284]_  = ~A168 & ~A169;
  assign \new_[11288]_  = ~A200 & A166;
  assign \new_[11289]_  = A167 & \new_[11288]_ ;
  assign \new_[11290]_  = \new_[11289]_  & \new_[11284]_ ;
  assign \new_[11294]_  = A266 & ~A265;
  assign \new_[11295]_  = ~A201 & \new_[11294]_ ;
  assign \new_[11299]_  = ~A302 & ~A301;
  assign \new_[11300]_  = A298 & \new_[11299]_ ;
  assign \new_[11301]_  = \new_[11300]_  & \new_[11295]_ ;
  assign \new_[11304]_  = ~A168 & ~A169;
  assign \new_[11308]_  = ~A199 & A166;
  assign \new_[11309]_  = A167 & \new_[11308]_ ;
  assign \new_[11310]_  = \new_[11309]_  & \new_[11304]_ ;
  assign \new_[11314]_  = A266 & ~A265;
  assign \new_[11315]_  = ~A200 & \new_[11314]_ ;
  assign \new_[11319]_  = ~A302 & ~A301;
  assign \new_[11320]_  = A298 & \new_[11319]_ ;
  assign \new_[11321]_  = \new_[11320]_  & \new_[11315]_ ;
  assign \new_[11324]_  = ~A169 & A170;
  assign \new_[11328]_  = A199 & ~A166;
  assign \new_[11329]_  = A167 & \new_[11328]_ ;
  assign \new_[11330]_  = \new_[11329]_  & \new_[11324]_ ;
  assign \new_[11334]_  = ~A268 & ~A266;
  assign \new_[11335]_  = A200 & \new_[11334]_ ;
  assign \new_[11339]_  = A299 & ~A298;
  assign \new_[11340]_  = ~A269 & \new_[11339]_ ;
  assign \new_[11341]_  = \new_[11340]_  & \new_[11335]_ ;
  assign \new_[11344]_  = ~A169 & A170;
  assign \new_[11348]_  = ~A199 & ~A166;
  assign \new_[11349]_  = A167 & \new_[11348]_ ;
  assign \new_[11350]_  = \new_[11349]_  & \new_[11344]_ ;
  assign \new_[11354]_  = A266 & ~A265;
  assign \new_[11355]_  = A200 & \new_[11354]_ ;
  assign \new_[11359]_  = ~A302 & ~A301;
  assign \new_[11360]_  = A298 & \new_[11359]_ ;
  assign \new_[11361]_  = \new_[11360]_  & \new_[11355]_ ;
  assign \new_[11364]_  = ~A169 & A170;
  assign \new_[11368]_  = ~A200 & ~A166;
  assign \new_[11369]_  = A167 & \new_[11368]_ ;
  assign \new_[11370]_  = \new_[11369]_  & \new_[11364]_ ;
  assign \new_[11374]_  = A265 & ~A203;
  assign \new_[11375]_  = ~A202 & \new_[11374]_ ;
  assign \new_[11379]_  = A299 & ~A298;
  assign \new_[11380]_  = A266 & \new_[11379]_ ;
  assign \new_[11381]_  = \new_[11380]_  & \new_[11375]_ ;
  assign \new_[11384]_  = ~A169 & A170;
  assign \new_[11388]_  = ~A200 & ~A166;
  assign \new_[11389]_  = A167 & \new_[11388]_ ;
  assign \new_[11390]_  = \new_[11389]_  & \new_[11384]_ ;
  assign \new_[11394]_  = ~A266 & ~A203;
  assign \new_[11395]_  = ~A202 & \new_[11394]_ ;
  assign \new_[11399]_  = A299 & ~A298;
  assign \new_[11400]_  = ~A267 & \new_[11399]_ ;
  assign \new_[11401]_  = \new_[11400]_  & \new_[11395]_ ;
  assign \new_[11404]_  = ~A169 & A170;
  assign \new_[11408]_  = ~A200 & ~A166;
  assign \new_[11409]_  = A167 & \new_[11408]_ ;
  assign \new_[11410]_  = \new_[11409]_  & \new_[11404]_ ;
  assign \new_[11414]_  = ~A265 & ~A203;
  assign \new_[11415]_  = ~A202 & \new_[11414]_ ;
  assign \new_[11419]_  = A299 & ~A298;
  assign \new_[11420]_  = ~A266 & \new_[11419]_ ;
  assign \new_[11421]_  = \new_[11420]_  & \new_[11415]_ ;
  assign \new_[11424]_  = ~A169 & A170;
  assign \new_[11428]_  = ~A200 & ~A166;
  assign \new_[11429]_  = A167 & \new_[11428]_ ;
  assign \new_[11430]_  = \new_[11429]_  & \new_[11424]_ ;
  assign \new_[11434]_  = ~A268 & ~A266;
  assign \new_[11435]_  = ~A201 & \new_[11434]_ ;
  assign \new_[11439]_  = A299 & ~A298;
  assign \new_[11440]_  = ~A269 & \new_[11439]_ ;
  assign \new_[11441]_  = \new_[11440]_  & \new_[11435]_ ;
  assign \new_[11444]_  = ~A169 & A170;
  assign \new_[11448]_  = ~A199 & ~A166;
  assign \new_[11449]_  = A167 & \new_[11448]_ ;
  assign \new_[11450]_  = \new_[11449]_  & \new_[11444]_ ;
  assign \new_[11454]_  = ~A268 & ~A266;
  assign \new_[11455]_  = ~A200 & \new_[11454]_ ;
  assign \new_[11459]_  = A299 & ~A298;
  assign \new_[11460]_  = ~A269 & \new_[11459]_ ;
  assign \new_[11461]_  = \new_[11460]_  & \new_[11455]_ ;
  assign \new_[11464]_  = ~A169 & A170;
  assign \new_[11468]_  = A199 & A166;
  assign \new_[11469]_  = ~A167 & \new_[11468]_ ;
  assign \new_[11470]_  = \new_[11469]_  & \new_[11464]_ ;
  assign \new_[11474]_  = ~A268 & ~A266;
  assign \new_[11475]_  = A200 & \new_[11474]_ ;
  assign \new_[11479]_  = A299 & ~A298;
  assign \new_[11480]_  = ~A269 & \new_[11479]_ ;
  assign \new_[11481]_  = \new_[11480]_  & \new_[11475]_ ;
  assign \new_[11484]_  = ~A169 & A170;
  assign \new_[11488]_  = ~A199 & A166;
  assign \new_[11489]_  = ~A167 & \new_[11488]_ ;
  assign \new_[11490]_  = \new_[11489]_  & \new_[11484]_ ;
  assign \new_[11494]_  = A266 & ~A265;
  assign \new_[11495]_  = A200 & \new_[11494]_ ;
  assign \new_[11499]_  = ~A302 & ~A301;
  assign \new_[11500]_  = A298 & \new_[11499]_ ;
  assign \new_[11501]_  = \new_[11500]_  & \new_[11495]_ ;
  assign \new_[11504]_  = ~A169 & A170;
  assign \new_[11508]_  = ~A200 & A166;
  assign \new_[11509]_  = ~A167 & \new_[11508]_ ;
  assign \new_[11510]_  = \new_[11509]_  & \new_[11504]_ ;
  assign \new_[11514]_  = A265 & ~A203;
  assign \new_[11515]_  = ~A202 & \new_[11514]_ ;
  assign \new_[11519]_  = A299 & ~A298;
  assign \new_[11520]_  = A266 & \new_[11519]_ ;
  assign \new_[11521]_  = \new_[11520]_  & \new_[11515]_ ;
  assign \new_[11524]_  = ~A169 & A170;
  assign \new_[11528]_  = ~A200 & A166;
  assign \new_[11529]_  = ~A167 & \new_[11528]_ ;
  assign \new_[11530]_  = \new_[11529]_  & \new_[11524]_ ;
  assign \new_[11534]_  = ~A266 & ~A203;
  assign \new_[11535]_  = ~A202 & \new_[11534]_ ;
  assign \new_[11539]_  = A299 & ~A298;
  assign \new_[11540]_  = ~A267 & \new_[11539]_ ;
  assign \new_[11541]_  = \new_[11540]_  & \new_[11535]_ ;
  assign \new_[11544]_  = ~A169 & A170;
  assign \new_[11548]_  = ~A200 & A166;
  assign \new_[11549]_  = ~A167 & \new_[11548]_ ;
  assign \new_[11550]_  = \new_[11549]_  & \new_[11544]_ ;
  assign \new_[11554]_  = ~A265 & ~A203;
  assign \new_[11555]_  = ~A202 & \new_[11554]_ ;
  assign \new_[11559]_  = A299 & ~A298;
  assign \new_[11560]_  = ~A266 & \new_[11559]_ ;
  assign \new_[11561]_  = \new_[11560]_  & \new_[11555]_ ;
  assign \new_[11564]_  = ~A169 & A170;
  assign \new_[11568]_  = ~A200 & A166;
  assign \new_[11569]_  = ~A167 & \new_[11568]_ ;
  assign \new_[11570]_  = \new_[11569]_  & \new_[11564]_ ;
  assign \new_[11574]_  = ~A268 & ~A266;
  assign \new_[11575]_  = ~A201 & \new_[11574]_ ;
  assign \new_[11579]_  = A299 & ~A298;
  assign \new_[11580]_  = ~A269 & \new_[11579]_ ;
  assign \new_[11581]_  = \new_[11580]_  & \new_[11575]_ ;
  assign \new_[11584]_  = ~A169 & A170;
  assign \new_[11588]_  = ~A199 & A166;
  assign \new_[11589]_  = ~A167 & \new_[11588]_ ;
  assign \new_[11590]_  = \new_[11589]_  & \new_[11584]_ ;
  assign \new_[11594]_  = ~A268 & ~A266;
  assign \new_[11595]_  = ~A200 & \new_[11594]_ ;
  assign \new_[11599]_  = A299 & ~A298;
  assign \new_[11600]_  = ~A269 & \new_[11599]_ ;
  assign \new_[11601]_  = \new_[11600]_  & \new_[11595]_ ;
  assign \new_[11604]_  = ~A169 & ~A170;
  assign \new_[11608]_  = A200 & A199;
  assign \new_[11609]_  = ~A168 & \new_[11608]_ ;
  assign \new_[11610]_  = \new_[11609]_  & \new_[11604]_ ;
  assign \new_[11614]_  = A267 & ~A266;
  assign \new_[11615]_  = A265 & \new_[11614]_ ;
  assign \new_[11619]_  = ~A300 & A298;
  assign \new_[11620]_  = A268 & \new_[11619]_ ;
  assign \new_[11621]_  = \new_[11620]_  & \new_[11615]_ ;
  assign \new_[11624]_  = ~A169 & ~A170;
  assign \new_[11628]_  = A200 & A199;
  assign \new_[11629]_  = ~A168 & \new_[11628]_ ;
  assign \new_[11630]_  = \new_[11629]_  & \new_[11624]_ ;
  assign \new_[11634]_  = A267 & ~A266;
  assign \new_[11635]_  = A265 & \new_[11634]_ ;
  assign \new_[11639]_  = A299 & A298;
  assign \new_[11640]_  = A268 & \new_[11639]_ ;
  assign \new_[11641]_  = \new_[11640]_  & \new_[11635]_ ;
  assign \new_[11644]_  = ~A169 & ~A170;
  assign \new_[11648]_  = A200 & A199;
  assign \new_[11649]_  = ~A168 & \new_[11648]_ ;
  assign \new_[11650]_  = \new_[11649]_  & \new_[11644]_ ;
  assign \new_[11654]_  = A267 & ~A266;
  assign \new_[11655]_  = A265 & \new_[11654]_ ;
  assign \new_[11659]_  = ~A299 & ~A298;
  assign \new_[11660]_  = A268 & \new_[11659]_ ;
  assign \new_[11661]_  = \new_[11660]_  & \new_[11655]_ ;
  assign \new_[11664]_  = ~A169 & ~A170;
  assign \new_[11668]_  = A200 & A199;
  assign \new_[11669]_  = ~A168 & \new_[11668]_ ;
  assign \new_[11670]_  = \new_[11669]_  & \new_[11664]_ ;
  assign \new_[11674]_  = A267 & ~A266;
  assign \new_[11675]_  = A265 & \new_[11674]_ ;
  assign \new_[11679]_  = ~A300 & A298;
  assign \new_[11680]_  = A269 & \new_[11679]_ ;
  assign \new_[11681]_  = \new_[11680]_  & \new_[11675]_ ;
  assign \new_[11684]_  = ~A169 & ~A170;
  assign \new_[11688]_  = A200 & A199;
  assign \new_[11689]_  = ~A168 & \new_[11688]_ ;
  assign \new_[11690]_  = \new_[11689]_  & \new_[11684]_ ;
  assign \new_[11694]_  = A267 & ~A266;
  assign \new_[11695]_  = A265 & \new_[11694]_ ;
  assign \new_[11699]_  = A299 & A298;
  assign \new_[11700]_  = A269 & \new_[11699]_ ;
  assign \new_[11701]_  = \new_[11700]_  & \new_[11695]_ ;
  assign \new_[11704]_  = ~A169 & ~A170;
  assign \new_[11708]_  = A200 & A199;
  assign \new_[11709]_  = ~A168 & \new_[11708]_ ;
  assign \new_[11710]_  = \new_[11709]_  & \new_[11704]_ ;
  assign \new_[11714]_  = A267 & ~A266;
  assign \new_[11715]_  = A265 & \new_[11714]_ ;
  assign \new_[11719]_  = ~A299 & ~A298;
  assign \new_[11720]_  = A269 & \new_[11719]_ ;
  assign \new_[11721]_  = \new_[11720]_  & \new_[11715]_ ;
  assign \new_[11724]_  = ~A169 & ~A170;
  assign \new_[11728]_  = A200 & ~A199;
  assign \new_[11729]_  = ~A168 & \new_[11728]_ ;
  assign \new_[11730]_  = \new_[11729]_  & \new_[11724]_ ;
  assign \new_[11734]_  = A298 & A266;
  assign \new_[11735]_  = A265 & \new_[11734]_ ;
  assign \new_[11739]_  = A301 & A300;
  assign \new_[11740]_  = ~A299 & \new_[11739]_ ;
  assign \new_[11741]_  = \new_[11740]_  & \new_[11735]_ ;
  assign \new_[11744]_  = ~A169 & ~A170;
  assign \new_[11748]_  = A200 & ~A199;
  assign \new_[11749]_  = ~A168 & \new_[11748]_ ;
  assign \new_[11750]_  = \new_[11749]_  & \new_[11744]_ ;
  assign \new_[11754]_  = A298 & A266;
  assign \new_[11755]_  = A265 & \new_[11754]_ ;
  assign \new_[11759]_  = A302 & A300;
  assign \new_[11760]_  = ~A299 & \new_[11759]_ ;
  assign \new_[11761]_  = \new_[11760]_  & \new_[11755]_ ;
  assign \new_[11764]_  = ~A169 & ~A170;
  assign \new_[11768]_  = A200 & ~A199;
  assign \new_[11769]_  = ~A168 & \new_[11768]_ ;
  assign \new_[11770]_  = \new_[11769]_  & \new_[11764]_ ;
  assign \new_[11774]_  = A298 & ~A267;
  assign \new_[11775]_  = ~A266 & \new_[11774]_ ;
  assign \new_[11779]_  = A301 & A300;
  assign \new_[11780]_  = ~A299 & \new_[11779]_ ;
  assign \new_[11781]_  = \new_[11780]_  & \new_[11775]_ ;
  assign \new_[11784]_  = ~A169 & ~A170;
  assign \new_[11788]_  = A200 & ~A199;
  assign \new_[11789]_  = ~A168 & \new_[11788]_ ;
  assign \new_[11790]_  = \new_[11789]_  & \new_[11784]_ ;
  assign \new_[11794]_  = A298 & ~A267;
  assign \new_[11795]_  = ~A266 & \new_[11794]_ ;
  assign \new_[11799]_  = A302 & A300;
  assign \new_[11800]_  = ~A299 & \new_[11799]_ ;
  assign \new_[11801]_  = \new_[11800]_  & \new_[11795]_ ;
  assign \new_[11804]_  = ~A169 & ~A170;
  assign \new_[11808]_  = A200 & ~A199;
  assign \new_[11809]_  = ~A168 & \new_[11808]_ ;
  assign \new_[11810]_  = \new_[11809]_  & \new_[11804]_ ;
  assign \new_[11814]_  = A298 & ~A266;
  assign \new_[11815]_  = ~A265 & \new_[11814]_ ;
  assign \new_[11819]_  = A301 & A300;
  assign \new_[11820]_  = ~A299 & \new_[11819]_ ;
  assign \new_[11821]_  = \new_[11820]_  & \new_[11815]_ ;
  assign \new_[11824]_  = ~A169 & ~A170;
  assign \new_[11828]_  = A200 & ~A199;
  assign \new_[11829]_  = ~A168 & \new_[11828]_ ;
  assign \new_[11830]_  = \new_[11829]_  & \new_[11824]_ ;
  assign \new_[11834]_  = A298 & ~A266;
  assign \new_[11835]_  = ~A265 & \new_[11834]_ ;
  assign \new_[11839]_  = A302 & A300;
  assign \new_[11840]_  = ~A299 & \new_[11839]_ ;
  assign \new_[11841]_  = \new_[11840]_  & \new_[11835]_ ;
  assign \new_[11844]_  = ~A169 & ~A170;
  assign \new_[11848]_  = ~A202 & ~A200;
  assign \new_[11849]_  = ~A168 & \new_[11848]_ ;
  assign \new_[11850]_  = \new_[11849]_  & \new_[11844]_ ;
  assign \new_[11854]_  = A266 & ~A265;
  assign \new_[11855]_  = ~A203 & \new_[11854]_ ;
  assign \new_[11859]_  = ~A302 & ~A301;
  assign \new_[11860]_  = A298 & \new_[11859]_ ;
  assign \new_[11861]_  = \new_[11860]_  & \new_[11855]_ ;
  assign \new_[11864]_  = ~A169 & ~A170;
  assign \new_[11868]_  = ~A201 & ~A200;
  assign \new_[11869]_  = ~A168 & \new_[11868]_ ;
  assign \new_[11870]_  = \new_[11869]_  & \new_[11864]_ ;
  assign \new_[11874]_  = A267 & ~A266;
  assign \new_[11875]_  = A265 & \new_[11874]_ ;
  assign \new_[11879]_  = ~A300 & A298;
  assign \new_[11880]_  = A268 & \new_[11879]_ ;
  assign \new_[11881]_  = \new_[11880]_  & \new_[11875]_ ;
  assign \new_[11884]_  = ~A169 & ~A170;
  assign \new_[11888]_  = ~A201 & ~A200;
  assign \new_[11889]_  = ~A168 & \new_[11888]_ ;
  assign \new_[11890]_  = \new_[11889]_  & \new_[11884]_ ;
  assign \new_[11894]_  = A267 & ~A266;
  assign \new_[11895]_  = A265 & \new_[11894]_ ;
  assign \new_[11899]_  = A299 & A298;
  assign \new_[11900]_  = A268 & \new_[11899]_ ;
  assign \new_[11901]_  = \new_[11900]_  & \new_[11895]_ ;
  assign \new_[11904]_  = ~A169 & ~A170;
  assign \new_[11908]_  = ~A201 & ~A200;
  assign \new_[11909]_  = ~A168 & \new_[11908]_ ;
  assign \new_[11910]_  = \new_[11909]_  & \new_[11904]_ ;
  assign \new_[11914]_  = A267 & ~A266;
  assign \new_[11915]_  = A265 & \new_[11914]_ ;
  assign \new_[11919]_  = ~A299 & ~A298;
  assign \new_[11920]_  = A268 & \new_[11919]_ ;
  assign \new_[11921]_  = \new_[11920]_  & \new_[11915]_ ;
  assign \new_[11924]_  = ~A169 & ~A170;
  assign \new_[11928]_  = ~A201 & ~A200;
  assign \new_[11929]_  = ~A168 & \new_[11928]_ ;
  assign \new_[11930]_  = \new_[11929]_  & \new_[11924]_ ;
  assign \new_[11934]_  = A267 & ~A266;
  assign \new_[11935]_  = A265 & \new_[11934]_ ;
  assign \new_[11939]_  = ~A300 & A298;
  assign \new_[11940]_  = A269 & \new_[11939]_ ;
  assign \new_[11941]_  = \new_[11940]_  & \new_[11935]_ ;
  assign \new_[11944]_  = ~A169 & ~A170;
  assign \new_[11948]_  = ~A201 & ~A200;
  assign \new_[11949]_  = ~A168 & \new_[11948]_ ;
  assign \new_[11950]_  = \new_[11949]_  & \new_[11944]_ ;
  assign \new_[11954]_  = A267 & ~A266;
  assign \new_[11955]_  = A265 & \new_[11954]_ ;
  assign \new_[11959]_  = A299 & A298;
  assign \new_[11960]_  = A269 & \new_[11959]_ ;
  assign \new_[11961]_  = \new_[11960]_  & \new_[11955]_ ;
  assign \new_[11964]_  = ~A169 & ~A170;
  assign \new_[11968]_  = ~A201 & ~A200;
  assign \new_[11969]_  = ~A168 & \new_[11968]_ ;
  assign \new_[11970]_  = \new_[11969]_  & \new_[11964]_ ;
  assign \new_[11974]_  = A267 & ~A266;
  assign \new_[11975]_  = A265 & \new_[11974]_ ;
  assign \new_[11979]_  = ~A299 & ~A298;
  assign \new_[11980]_  = A269 & \new_[11979]_ ;
  assign \new_[11981]_  = \new_[11980]_  & \new_[11975]_ ;
  assign \new_[11984]_  = ~A169 & ~A170;
  assign \new_[11988]_  = ~A200 & A199;
  assign \new_[11989]_  = ~A168 & \new_[11988]_ ;
  assign \new_[11990]_  = \new_[11989]_  & \new_[11984]_ ;
  assign \new_[11994]_  = A265 & A202;
  assign \new_[11995]_  = A201 & \new_[11994]_ ;
  assign \new_[11999]_  = A299 & ~A298;
  assign \new_[12000]_  = A266 & \new_[11999]_ ;
  assign \new_[12001]_  = \new_[12000]_  & \new_[11995]_ ;
  assign \new_[12004]_  = ~A169 & ~A170;
  assign \new_[12008]_  = ~A200 & A199;
  assign \new_[12009]_  = ~A168 & \new_[12008]_ ;
  assign \new_[12010]_  = \new_[12009]_  & \new_[12004]_ ;
  assign \new_[12014]_  = ~A266 & A202;
  assign \new_[12015]_  = A201 & \new_[12014]_ ;
  assign \new_[12019]_  = A299 & ~A298;
  assign \new_[12020]_  = ~A267 & \new_[12019]_ ;
  assign \new_[12021]_  = \new_[12020]_  & \new_[12015]_ ;
  assign \new_[12024]_  = ~A169 & ~A170;
  assign \new_[12028]_  = ~A200 & A199;
  assign \new_[12029]_  = ~A168 & \new_[12028]_ ;
  assign \new_[12030]_  = \new_[12029]_  & \new_[12024]_ ;
  assign \new_[12034]_  = ~A265 & A202;
  assign \new_[12035]_  = A201 & \new_[12034]_ ;
  assign \new_[12039]_  = A299 & ~A298;
  assign \new_[12040]_  = ~A266 & \new_[12039]_ ;
  assign \new_[12041]_  = \new_[12040]_  & \new_[12035]_ ;
  assign \new_[12044]_  = ~A169 & ~A170;
  assign \new_[12048]_  = ~A200 & A199;
  assign \new_[12049]_  = ~A168 & \new_[12048]_ ;
  assign \new_[12050]_  = \new_[12049]_  & \new_[12044]_ ;
  assign \new_[12054]_  = A265 & A203;
  assign \new_[12055]_  = A201 & \new_[12054]_ ;
  assign \new_[12059]_  = A299 & ~A298;
  assign \new_[12060]_  = A266 & \new_[12059]_ ;
  assign \new_[12061]_  = \new_[12060]_  & \new_[12055]_ ;
  assign \new_[12064]_  = ~A169 & ~A170;
  assign \new_[12068]_  = ~A200 & A199;
  assign \new_[12069]_  = ~A168 & \new_[12068]_ ;
  assign \new_[12070]_  = \new_[12069]_  & \new_[12064]_ ;
  assign \new_[12074]_  = ~A266 & A203;
  assign \new_[12075]_  = A201 & \new_[12074]_ ;
  assign \new_[12079]_  = A299 & ~A298;
  assign \new_[12080]_  = ~A267 & \new_[12079]_ ;
  assign \new_[12081]_  = \new_[12080]_  & \new_[12075]_ ;
  assign \new_[12084]_  = ~A169 & ~A170;
  assign \new_[12088]_  = ~A200 & A199;
  assign \new_[12089]_  = ~A168 & \new_[12088]_ ;
  assign \new_[12090]_  = \new_[12089]_  & \new_[12084]_ ;
  assign \new_[12094]_  = ~A265 & A203;
  assign \new_[12095]_  = A201 & \new_[12094]_ ;
  assign \new_[12099]_  = A299 & ~A298;
  assign \new_[12100]_  = ~A266 & \new_[12099]_ ;
  assign \new_[12101]_  = \new_[12100]_  & \new_[12095]_ ;
  assign \new_[12104]_  = ~A169 & ~A170;
  assign \new_[12108]_  = ~A200 & ~A199;
  assign \new_[12109]_  = ~A168 & \new_[12108]_ ;
  assign \new_[12110]_  = \new_[12109]_  & \new_[12104]_ ;
  assign \new_[12114]_  = A267 & ~A266;
  assign \new_[12115]_  = A265 & \new_[12114]_ ;
  assign \new_[12119]_  = ~A300 & A298;
  assign \new_[12120]_  = A268 & \new_[12119]_ ;
  assign \new_[12121]_  = \new_[12120]_  & \new_[12115]_ ;
  assign \new_[12124]_  = ~A169 & ~A170;
  assign \new_[12128]_  = ~A200 & ~A199;
  assign \new_[12129]_  = ~A168 & \new_[12128]_ ;
  assign \new_[12130]_  = \new_[12129]_  & \new_[12124]_ ;
  assign \new_[12134]_  = A267 & ~A266;
  assign \new_[12135]_  = A265 & \new_[12134]_ ;
  assign \new_[12139]_  = A299 & A298;
  assign \new_[12140]_  = A268 & \new_[12139]_ ;
  assign \new_[12141]_  = \new_[12140]_  & \new_[12135]_ ;
  assign \new_[12144]_  = ~A169 & ~A170;
  assign \new_[12148]_  = ~A200 & ~A199;
  assign \new_[12149]_  = ~A168 & \new_[12148]_ ;
  assign \new_[12150]_  = \new_[12149]_  & \new_[12144]_ ;
  assign \new_[12154]_  = A267 & ~A266;
  assign \new_[12155]_  = A265 & \new_[12154]_ ;
  assign \new_[12159]_  = ~A299 & ~A298;
  assign \new_[12160]_  = A268 & \new_[12159]_ ;
  assign \new_[12161]_  = \new_[12160]_  & \new_[12155]_ ;
  assign \new_[12164]_  = ~A169 & ~A170;
  assign \new_[12168]_  = ~A200 & ~A199;
  assign \new_[12169]_  = ~A168 & \new_[12168]_ ;
  assign \new_[12170]_  = \new_[12169]_  & \new_[12164]_ ;
  assign \new_[12174]_  = A267 & ~A266;
  assign \new_[12175]_  = A265 & \new_[12174]_ ;
  assign \new_[12179]_  = ~A300 & A298;
  assign \new_[12180]_  = A269 & \new_[12179]_ ;
  assign \new_[12181]_  = \new_[12180]_  & \new_[12175]_ ;
  assign \new_[12184]_  = ~A169 & ~A170;
  assign \new_[12188]_  = ~A200 & ~A199;
  assign \new_[12189]_  = ~A168 & \new_[12188]_ ;
  assign \new_[12190]_  = \new_[12189]_  & \new_[12184]_ ;
  assign \new_[12194]_  = A267 & ~A266;
  assign \new_[12195]_  = A265 & \new_[12194]_ ;
  assign \new_[12199]_  = A299 & A298;
  assign \new_[12200]_  = A269 & \new_[12199]_ ;
  assign \new_[12201]_  = \new_[12200]_  & \new_[12195]_ ;
  assign \new_[12204]_  = ~A169 & ~A170;
  assign \new_[12208]_  = ~A200 & ~A199;
  assign \new_[12209]_  = ~A168 & \new_[12208]_ ;
  assign \new_[12210]_  = \new_[12209]_  & \new_[12204]_ ;
  assign \new_[12214]_  = A267 & ~A266;
  assign \new_[12215]_  = A265 & \new_[12214]_ ;
  assign \new_[12219]_  = ~A299 & ~A298;
  assign \new_[12220]_  = A269 & \new_[12219]_ ;
  assign \new_[12221]_  = \new_[12220]_  & \new_[12215]_ ;
  assign \new_[12225]_  = ~A200 & A166;
  assign \new_[12226]_  = A168 & \new_[12225]_ ;
  assign \new_[12230]_  = ~A266 & ~A203;
  assign \new_[12231]_  = ~A202 & \new_[12230]_ ;
  assign \new_[12232]_  = \new_[12231]_  & \new_[12226]_ ;
  assign \new_[12236]_  = A298 & ~A269;
  assign \new_[12237]_  = ~A268 & \new_[12236]_ ;
  assign \new_[12241]_  = A301 & A300;
  assign \new_[12242]_  = ~A299 & \new_[12241]_ ;
  assign \new_[12243]_  = \new_[12242]_  & \new_[12237]_ ;
  assign \new_[12247]_  = ~A200 & A166;
  assign \new_[12248]_  = A168 & \new_[12247]_ ;
  assign \new_[12252]_  = ~A266 & ~A203;
  assign \new_[12253]_  = ~A202 & \new_[12252]_ ;
  assign \new_[12254]_  = \new_[12253]_  & \new_[12248]_ ;
  assign \new_[12258]_  = A298 & ~A269;
  assign \new_[12259]_  = ~A268 & \new_[12258]_ ;
  assign \new_[12263]_  = A302 & A300;
  assign \new_[12264]_  = ~A299 & \new_[12263]_ ;
  assign \new_[12265]_  = \new_[12264]_  & \new_[12259]_ ;
  assign \new_[12269]_  = A199 & A166;
  assign \new_[12270]_  = A168 & \new_[12269]_ ;
  assign \new_[12274]_  = A202 & A201;
  assign \new_[12275]_  = ~A200 & \new_[12274]_ ;
  assign \new_[12276]_  = \new_[12275]_  & \new_[12270]_ ;
  assign \new_[12280]_  = A267 & ~A266;
  assign \new_[12281]_  = A265 & \new_[12280]_ ;
  assign \new_[12285]_  = ~A300 & A298;
  assign \new_[12286]_  = A268 & \new_[12285]_ ;
  assign \new_[12287]_  = \new_[12286]_  & \new_[12281]_ ;
  assign \new_[12291]_  = A199 & A166;
  assign \new_[12292]_  = A168 & \new_[12291]_ ;
  assign \new_[12296]_  = A202 & A201;
  assign \new_[12297]_  = ~A200 & \new_[12296]_ ;
  assign \new_[12298]_  = \new_[12297]_  & \new_[12292]_ ;
  assign \new_[12302]_  = A267 & ~A266;
  assign \new_[12303]_  = A265 & \new_[12302]_ ;
  assign \new_[12307]_  = A299 & A298;
  assign \new_[12308]_  = A268 & \new_[12307]_ ;
  assign \new_[12309]_  = \new_[12308]_  & \new_[12303]_ ;
  assign \new_[12313]_  = A199 & A166;
  assign \new_[12314]_  = A168 & \new_[12313]_ ;
  assign \new_[12318]_  = A202 & A201;
  assign \new_[12319]_  = ~A200 & \new_[12318]_ ;
  assign \new_[12320]_  = \new_[12319]_  & \new_[12314]_ ;
  assign \new_[12324]_  = A267 & ~A266;
  assign \new_[12325]_  = A265 & \new_[12324]_ ;
  assign \new_[12329]_  = ~A299 & ~A298;
  assign \new_[12330]_  = A268 & \new_[12329]_ ;
  assign \new_[12331]_  = \new_[12330]_  & \new_[12325]_ ;
  assign \new_[12335]_  = A199 & A166;
  assign \new_[12336]_  = A168 & \new_[12335]_ ;
  assign \new_[12340]_  = A202 & A201;
  assign \new_[12341]_  = ~A200 & \new_[12340]_ ;
  assign \new_[12342]_  = \new_[12341]_  & \new_[12336]_ ;
  assign \new_[12346]_  = A267 & ~A266;
  assign \new_[12347]_  = A265 & \new_[12346]_ ;
  assign \new_[12351]_  = ~A300 & A298;
  assign \new_[12352]_  = A269 & \new_[12351]_ ;
  assign \new_[12353]_  = \new_[12352]_  & \new_[12347]_ ;
  assign \new_[12357]_  = A199 & A166;
  assign \new_[12358]_  = A168 & \new_[12357]_ ;
  assign \new_[12362]_  = A202 & A201;
  assign \new_[12363]_  = ~A200 & \new_[12362]_ ;
  assign \new_[12364]_  = \new_[12363]_  & \new_[12358]_ ;
  assign \new_[12368]_  = A267 & ~A266;
  assign \new_[12369]_  = A265 & \new_[12368]_ ;
  assign \new_[12373]_  = A299 & A298;
  assign \new_[12374]_  = A269 & \new_[12373]_ ;
  assign \new_[12375]_  = \new_[12374]_  & \new_[12369]_ ;
  assign \new_[12379]_  = A199 & A166;
  assign \new_[12380]_  = A168 & \new_[12379]_ ;
  assign \new_[12384]_  = A202 & A201;
  assign \new_[12385]_  = ~A200 & \new_[12384]_ ;
  assign \new_[12386]_  = \new_[12385]_  & \new_[12380]_ ;
  assign \new_[12390]_  = A267 & ~A266;
  assign \new_[12391]_  = A265 & \new_[12390]_ ;
  assign \new_[12395]_  = ~A299 & ~A298;
  assign \new_[12396]_  = A269 & \new_[12395]_ ;
  assign \new_[12397]_  = \new_[12396]_  & \new_[12391]_ ;
  assign \new_[12401]_  = A199 & A166;
  assign \new_[12402]_  = A168 & \new_[12401]_ ;
  assign \new_[12406]_  = A203 & A201;
  assign \new_[12407]_  = ~A200 & \new_[12406]_ ;
  assign \new_[12408]_  = \new_[12407]_  & \new_[12402]_ ;
  assign \new_[12412]_  = A267 & ~A266;
  assign \new_[12413]_  = A265 & \new_[12412]_ ;
  assign \new_[12417]_  = ~A300 & A298;
  assign \new_[12418]_  = A268 & \new_[12417]_ ;
  assign \new_[12419]_  = \new_[12418]_  & \new_[12413]_ ;
  assign \new_[12423]_  = A199 & A166;
  assign \new_[12424]_  = A168 & \new_[12423]_ ;
  assign \new_[12428]_  = A203 & A201;
  assign \new_[12429]_  = ~A200 & \new_[12428]_ ;
  assign \new_[12430]_  = \new_[12429]_  & \new_[12424]_ ;
  assign \new_[12434]_  = A267 & ~A266;
  assign \new_[12435]_  = A265 & \new_[12434]_ ;
  assign \new_[12439]_  = A299 & A298;
  assign \new_[12440]_  = A268 & \new_[12439]_ ;
  assign \new_[12441]_  = \new_[12440]_  & \new_[12435]_ ;
  assign \new_[12445]_  = A199 & A166;
  assign \new_[12446]_  = A168 & \new_[12445]_ ;
  assign \new_[12450]_  = A203 & A201;
  assign \new_[12451]_  = ~A200 & \new_[12450]_ ;
  assign \new_[12452]_  = \new_[12451]_  & \new_[12446]_ ;
  assign \new_[12456]_  = A267 & ~A266;
  assign \new_[12457]_  = A265 & \new_[12456]_ ;
  assign \new_[12461]_  = ~A299 & ~A298;
  assign \new_[12462]_  = A268 & \new_[12461]_ ;
  assign \new_[12463]_  = \new_[12462]_  & \new_[12457]_ ;
  assign \new_[12467]_  = A199 & A166;
  assign \new_[12468]_  = A168 & \new_[12467]_ ;
  assign \new_[12472]_  = A203 & A201;
  assign \new_[12473]_  = ~A200 & \new_[12472]_ ;
  assign \new_[12474]_  = \new_[12473]_  & \new_[12468]_ ;
  assign \new_[12478]_  = A267 & ~A266;
  assign \new_[12479]_  = A265 & \new_[12478]_ ;
  assign \new_[12483]_  = ~A300 & A298;
  assign \new_[12484]_  = A269 & \new_[12483]_ ;
  assign \new_[12485]_  = \new_[12484]_  & \new_[12479]_ ;
  assign \new_[12489]_  = A199 & A166;
  assign \new_[12490]_  = A168 & \new_[12489]_ ;
  assign \new_[12494]_  = A203 & A201;
  assign \new_[12495]_  = ~A200 & \new_[12494]_ ;
  assign \new_[12496]_  = \new_[12495]_  & \new_[12490]_ ;
  assign \new_[12500]_  = A267 & ~A266;
  assign \new_[12501]_  = A265 & \new_[12500]_ ;
  assign \new_[12505]_  = A299 & A298;
  assign \new_[12506]_  = A269 & \new_[12505]_ ;
  assign \new_[12507]_  = \new_[12506]_  & \new_[12501]_ ;
  assign \new_[12511]_  = A199 & A166;
  assign \new_[12512]_  = A168 & \new_[12511]_ ;
  assign \new_[12516]_  = A203 & A201;
  assign \new_[12517]_  = ~A200 & \new_[12516]_ ;
  assign \new_[12518]_  = \new_[12517]_  & \new_[12512]_ ;
  assign \new_[12522]_  = A267 & ~A266;
  assign \new_[12523]_  = A265 & \new_[12522]_ ;
  assign \new_[12527]_  = ~A299 & ~A298;
  assign \new_[12528]_  = A269 & \new_[12527]_ ;
  assign \new_[12529]_  = \new_[12528]_  & \new_[12523]_ ;
  assign \new_[12533]_  = ~A200 & A167;
  assign \new_[12534]_  = A168 & \new_[12533]_ ;
  assign \new_[12538]_  = ~A266 & ~A203;
  assign \new_[12539]_  = ~A202 & \new_[12538]_ ;
  assign \new_[12540]_  = \new_[12539]_  & \new_[12534]_ ;
  assign \new_[12544]_  = A298 & ~A269;
  assign \new_[12545]_  = ~A268 & \new_[12544]_ ;
  assign \new_[12549]_  = A301 & A300;
  assign \new_[12550]_  = ~A299 & \new_[12549]_ ;
  assign \new_[12551]_  = \new_[12550]_  & \new_[12545]_ ;
  assign \new_[12555]_  = ~A200 & A167;
  assign \new_[12556]_  = A168 & \new_[12555]_ ;
  assign \new_[12560]_  = ~A266 & ~A203;
  assign \new_[12561]_  = ~A202 & \new_[12560]_ ;
  assign \new_[12562]_  = \new_[12561]_  & \new_[12556]_ ;
  assign \new_[12566]_  = A298 & ~A269;
  assign \new_[12567]_  = ~A268 & \new_[12566]_ ;
  assign \new_[12571]_  = A302 & A300;
  assign \new_[12572]_  = ~A299 & \new_[12571]_ ;
  assign \new_[12573]_  = \new_[12572]_  & \new_[12567]_ ;
  assign \new_[12577]_  = A199 & A167;
  assign \new_[12578]_  = A168 & \new_[12577]_ ;
  assign \new_[12582]_  = A202 & A201;
  assign \new_[12583]_  = ~A200 & \new_[12582]_ ;
  assign \new_[12584]_  = \new_[12583]_  & \new_[12578]_ ;
  assign \new_[12588]_  = A267 & ~A266;
  assign \new_[12589]_  = A265 & \new_[12588]_ ;
  assign \new_[12593]_  = ~A300 & A298;
  assign \new_[12594]_  = A268 & \new_[12593]_ ;
  assign \new_[12595]_  = \new_[12594]_  & \new_[12589]_ ;
  assign \new_[12599]_  = A199 & A167;
  assign \new_[12600]_  = A168 & \new_[12599]_ ;
  assign \new_[12604]_  = A202 & A201;
  assign \new_[12605]_  = ~A200 & \new_[12604]_ ;
  assign \new_[12606]_  = \new_[12605]_  & \new_[12600]_ ;
  assign \new_[12610]_  = A267 & ~A266;
  assign \new_[12611]_  = A265 & \new_[12610]_ ;
  assign \new_[12615]_  = A299 & A298;
  assign \new_[12616]_  = A268 & \new_[12615]_ ;
  assign \new_[12617]_  = \new_[12616]_  & \new_[12611]_ ;
  assign \new_[12621]_  = A199 & A167;
  assign \new_[12622]_  = A168 & \new_[12621]_ ;
  assign \new_[12626]_  = A202 & A201;
  assign \new_[12627]_  = ~A200 & \new_[12626]_ ;
  assign \new_[12628]_  = \new_[12627]_  & \new_[12622]_ ;
  assign \new_[12632]_  = A267 & ~A266;
  assign \new_[12633]_  = A265 & \new_[12632]_ ;
  assign \new_[12637]_  = ~A299 & ~A298;
  assign \new_[12638]_  = A268 & \new_[12637]_ ;
  assign \new_[12639]_  = \new_[12638]_  & \new_[12633]_ ;
  assign \new_[12643]_  = A199 & A167;
  assign \new_[12644]_  = A168 & \new_[12643]_ ;
  assign \new_[12648]_  = A202 & A201;
  assign \new_[12649]_  = ~A200 & \new_[12648]_ ;
  assign \new_[12650]_  = \new_[12649]_  & \new_[12644]_ ;
  assign \new_[12654]_  = A267 & ~A266;
  assign \new_[12655]_  = A265 & \new_[12654]_ ;
  assign \new_[12659]_  = ~A300 & A298;
  assign \new_[12660]_  = A269 & \new_[12659]_ ;
  assign \new_[12661]_  = \new_[12660]_  & \new_[12655]_ ;
  assign \new_[12665]_  = A199 & A167;
  assign \new_[12666]_  = A168 & \new_[12665]_ ;
  assign \new_[12670]_  = A202 & A201;
  assign \new_[12671]_  = ~A200 & \new_[12670]_ ;
  assign \new_[12672]_  = \new_[12671]_  & \new_[12666]_ ;
  assign \new_[12676]_  = A267 & ~A266;
  assign \new_[12677]_  = A265 & \new_[12676]_ ;
  assign \new_[12681]_  = A299 & A298;
  assign \new_[12682]_  = A269 & \new_[12681]_ ;
  assign \new_[12683]_  = \new_[12682]_  & \new_[12677]_ ;
  assign \new_[12687]_  = A199 & A167;
  assign \new_[12688]_  = A168 & \new_[12687]_ ;
  assign \new_[12692]_  = A202 & A201;
  assign \new_[12693]_  = ~A200 & \new_[12692]_ ;
  assign \new_[12694]_  = \new_[12693]_  & \new_[12688]_ ;
  assign \new_[12698]_  = A267 & ~A266;
  assign \new_[12699]_  = A265 & \new_[12698]_ ;
  assign \new_[12703]_  = ~A299 & ~A298;
  assign \new_[12704]_  = A269 & \new_[12703]_ ;
  assign \new_[12705]_  = \new_[12704]_  & \new_[12699]_ ;
  assign \new_[12709]_  = A199 & A167;
  assign \new_[12710]_  = A168 & \new_[12709]_ ;
  assign \new_[12714]_  = A203 & A201;
  assign \new_[12715]_  = ~A200 & \new_[12714]_ ;
  assign \new_[12716]_  = \new_[12715]_  & \new_[12710]_ ;
  assign \new_[12720]_  = A267 & ~A266;
  assign \new_[12721]_  = A265 & \new_[12720]_ ;
  assign \new_[12725]_  = ~A300 & A298;
  assign \new_[12726]_  = A268 & \new_[12725]_ ;
  assign \new_[12727]_  = \new_[12726]_  & \new_[12721]_ ;
  assign \new_[12731]_  = A199 & A167;
  assign \new_[12732]_  = A168 & \new_[12731]_ ;
  assign \new_[12736]_  = A203 & A201;
  assign \new_[12737]_  = ~A200 & \new_[12736]_ ;
  assign \new_[12738]_  = \new_[12737]_  & \new_[12732]_ ;
  assign \new_[12742]_  = A267 & ~A266;
  assign \new_[12743]_  = A265 & \new_[12742]_ ;
  assign \new_[12747]_  = A299 & A298;
  assign \new_[12748]_  = A268 & \new_[12747]_ ;
  assign \new_[12749]_  = \new_[12748]_  & \new_[12743]_ ;
  assign \new_[12753]_  = A199 & A167;
  assign \new_[12754]_  = A168 & \new_[12753]_ ;
  assign \new_[12758]_  = A203 & A201;
  assign \new_[12759]_  = ~A200 & \new_[12758]_ ;
  assign \new_[12760]_  = \new_[12759]_  & \new_[12754]_ ;
  assign \new_[12764]_  = A267 & ~A266;
  assign \new_[12765]_  = A265 & \new_[12764]_ ;
  assign \new_[12769]_  = ~A299 & ~A298;
  assign \new_[12770]_  = A268 & \new_[12769]_ ;
  assign \new_[12771]_  = \new_[12770]_  & \new_[12765]_ ;
  assign \new_[12775]_  = A199 & A167;
  assign \new_[12776]_  = A168 & \new_[12775]_ ;
  assign \new_[12780]_  = A203 & A201;
  assign \new_[12781]_  = ~A200 & \new_[12780]_ ;
  assign \new_[12782]_  = \new_[12781]_  & \new_[12776]_ ;
  assign \new_[12786]_  = A267 & ~A266;
  assign \new_[12787]_  = A265 & \new_[12786]_ ;
  assign \new_[12791]_  = ~A300 & A298;
  assign \new_[12792]_  = A269 & \new_[12791]_ ;
  assign \new_[12793]_  = \new_[12792]_  & \new_[12787]_ ;
  assign \new_[12797]_  = A199 & A167;
  assign \new_[12798]_  = A168 & \new_[12797]_ ;
  assign \new_[12802]_  = A203 & A201;
  assign \new_[12803]_  = ~A200 & \new_[12802]_ ;
  assign \new_[12804]_  = \new_[12803]_  & \new_[12798]_ ;
  assign \new_[12808]_  = A267 & ~A266;
  assign \new_[12809]_  = A265 & \new_[12808]_ ;
  assign \new_[12813]_  = A299 & A298;
  assign \new_[12814]_  = A269 & \new_[12813]_ ;
  assign \new_[12815]_  = \new_[12814]_  & \new_[12809]_ ;
  assign \new_[12819]_  = A199 & A167;
  assign \new_[12820]_  = A168 & \new_[12819]_ ;
  assign \new_[12824]_  = A203 & A201;
  assign \new_[12825]_  = ~A200 & \new_[12824]_ ;
  assign \new_[12826]_  = \new_[12825]_  & \new_[12820]_ ;
  assign \new_[12830]_  = A267 & ~A266;
  assign \new_[12831]_  = A265 & \new_[12830]_ ;
  assign \new_[12835]_  = ~A299 & ~A298;
  assign \new_[12836]_  = A269 & \new_[12835]_ ;
  assign \new_[12837]_  = \new_[12836]_  & \new_[12831]_ ;
  assign \new_[12841]_  = ~A166 & ~A167;
  assign \new_[12842]_  = A170 & \new_[12841]_ ;
  assign \new_[12846]_  = A265 & A200;
  assign \new_[12847]_  = A199 & \new_[12846]_ ;
  assign \new_[12848]_  = \new_[12847]_  & \new_[12842]_ ;
  assign \new_[12852]_  = A268 & A267;
  assign \new_[12853]_  = ~A266 & \new_[12852]_ ;
  assign \new_[12857]_  = ~A302 & ~A301;
  assign \new_[12858]_  = A298 & \new_[12857]_ ;
  assign \new_[12859]_  = \new_[12858]_  & \new_[12853]_ ;
  assign \new_[12863]_  = ~A166 & ~A167;
  assign \new_[12864]_  = A170 & \new_[12863]_ ;
  assign \new_[12868]_  = A265 & A200;
  assign \new_[12869]_  = A199 & \new_[12868]_ ;
  assign \new_[12870]_  = \new_[12869]_  & \new_[12864]_ ;
  assign \new_[12874]_  = A269 & A267;
  assign \new_[12875]_  = ~A266 & \new_[12874]_ ;
  assign \new_[12879]_  = ~A302 & ~A301;
  assign \new_[12880]_  = A298 & \new_[12879]_ ;
  assign \new_[12881]_  = \new_[12880]_  & \new_[12875]_ ;
  assign \new_[12885]_  = ~A166 & ~A167;
  assign \new_[12886]_  = A170 & \new_[12885]_ ;
  assign \new_[12890]_  = ~A266 & A200;
  assign \new_[12891]_  = ~A199 & \new_[12890]_ ;
  assign \new_[12892]_  = \new_[12891]_  & \new_[12886]_ ;
  assign \new_[12896]_  = A298 & ~A269;
  assign \new_[12897]_  = ~A268 & \new_[12896]_ ;
  assign \new_[12901]_  = A301 & A300;
  assign \new_[12902]_  = ~A299 & \new_[12901]_ ;
  assign \new_[12903]_  = \new_[12902]_  & \new_[12897]_ ;
  assign \new_[12907]_  = ~A166 & ~A167;
  assign \new_[12908]_  = A170 & \new_[12907]_ ;
  assign \new_[12912]_  = ~A266 & A200;
  assign \new_[12913]_  = ~A199 & \new_[12912]_ ;
  assign \new_[12914]_  = \new_[12913]_  & \new_[12908]_ ;
  assign \new_[12918]_  = A298 & ~A269;
  assign \new_[12919]_  = ~A268 & \new_[12918]_ ;
  assign \new_[12923]_  = A302 & A300;
  assign \new_[12924]_  = ~A299 & \new_[12923]_ ;
  assign \new_[12925]_  = \new_[12924]_  & \new_[12919]_ ;
  assign \new_[12929]_  = ~A166 & ~A167;
  assign \new_[12930]_  = A170 & \new_[12929]_ ;
  assign \new_[12934]_  = ~A203 & ~A202;
  assign \new_[12935]_  = ~A200 & \new_[12934]_ ;
  assign \new_[12936]_  = \new_[12935]_  & \new_[12930]_ ;
  assign \new_[12940]_  = A267 & ~A266;
  assign \new_[12941]_  = A265 & \new_[12940]_ ;
  assign \new_[12945]_  = ~A300 & A298;
  assign \new_[12946]_  = A268 & \new_[12945]_ ;
  assign \new_[12947]_  = \new_[12946]_  & \new_[12941]_ ;
  assign \new_[12951]_  = ~A166 & ~A167;
  assign \new_[12952]_  = A170 & \new_[12951]_ ;
  assign \new_[12956]_  = ~A203 & ~A202;
  assign \new_[12957]_  = ~A200 & \new_[12956]_ ;
  assign \new_[12958]_  = \new_[12957]_  & \new_[12952]_ ;
  assign \new_[12962]_  = A267 & ~A266;
  assign \new_[12963]_  = A265 & \new_[12962]_ ;
  assign \new_[12967]_  = A299 & A298;
  assign \new_[12968]_  = A268 & \new_[12967]_ ;
  assign \new_[12969]_  = \new_[12968]_  & \new_[12963]_ ;
  assign \new_[12973]_  = ~A166 & ~A167;
  assign \new_[12974]_  = A170 & \new_[12973]_ ;
  assign \new_[12978]_  = ~A203 & ~A202;
  assign \new_[12979]_  = ~A200 & \new_[12978]_ ;
  assign \new_[12980]_  = \new_[12979]_  & \new_[12974]_ ;
  assign \new_[12984]_  = A267 & ~A266;
  assign \new_[12985]_  = A265 & \new_[12984]_ ;
  assign \new_[12989]_  = ~A299 & ~A298;
  assign \new_[12990]_  = A268 & \new_[12989]_ ;
  assign \new_[12991]_  = \new_[12990]_  & \new_[12985]_ ;
  assign \new_[12995]_  = ~A166 & ~A167;
  assign \new_[12996]_  = A170 & \new_[12995]_ ;
  assign \new_[13000]_  = ~A203 & ~A202;
  assign \new_[13001]_  = ~A200 & \new_[13000]_ ;
  assign \new_[13002]_  = \new_[13001]_  & \new_[12996]_ ;
  assign \new_[13006]_  = A267 & ~A266;
  assign \new_[13007]_  = A265 & \new_[13006]_ ;
  assign \new_[13011]_  = ~A300 & A298;
  assign \new_[13012]_  = A269 & \new_[13011]_ ;
  assign \new_[13013]_  = \new_[13012]_  & \new_[13007]_ ;
  assign \new_[13017]_  = ~A166 & ~A167;
  assign \new_[13018]_  = A170 & \new_[13017]_ ;
  assign \new_[13022]_  = ~A203 & ~A202;
  assign \new_[13023]_  = ~A200 & \new_[13022]_ ;
  assign \new_[13024]_  = \new_[13023]_  & \new_[13018]_ ;
  assign \new_[13028]_  = A267 & ~A266;
  assign \new_[13029]_  = A265 & \new_[13028]_ ;
  assign \new_[13033]_  = A299 & A298;
  assign \new_[13034]_  = A269 & \new_[13033]_ ;
  assign \new_[13035]_  = \new_[13034]_  & \new_[13029]_ ;
  assign \new_[13039]_  = ~A166 & ~A167;
  assign \new_[13040]_  = A170 & \new_[13039]_ ;
  assign \new_[13044]_  = ~A203 & ~A202;
  assign \new_[13045]_  = ~A200 & \new_[13044]_ ;
  assign \new_[13046]_  = \new_[13045]_  & \new_[13040]_ ;
  assign \new_[13050]_  = A267 & ~A266;
  assign \new_[13051]_  = A265 & \new_[13050]_ ;
  assign \new_[13055]_  = ~A299 & ~A298;
  assign \new_[13056]_  = A269 & \new_[13055]_ ;
  assign \new_[13057]_  = \new_[13056]_  & \new_[13051]_ ;
  assign \new_[13061]_  = ~A166 & ~A167;
  assign \new_[13062]_  = A170 & \new_[13061]_ ;
  assign \new_[13066]_  = A265 & ~A201;
  assign \new_[13067]_  = ~A200 & \new_[13066]_ ;
  assign \new_[13068]_  = \new_[13067]_  & \new_[13062]_ ;
  assign \new_[13072]_  = A268 & A267;
  assign \new_[13073]_  = ~A266 & \new_[13072]_ ;
  assign \new_[13077]_  = ~A302 & ~A301;
  assign \new_[13078]_  = A298 & \new_[13077]_ ;
  assign \new_[13079]_  = \new_[13078]_  & \new_[13073]_ ;
  assign \new_[13083]_  = ~A166 & ~A167;
  assign \new_[13084]_  = A170 & \new_[13083]_ ;
  assign \new_[13088]_  = A265 & ~A201;
  assign \new_[13089]_  = ~A200 & \new_[13088]_ ;
  assign \new_[13090]_  = \new_[13089]_  & \new_[13084]_ ;
  assign \new_[13094]_  = A269 & A267;
  assign \new_[13095]_  = ~A266 & \new_[13094]_ ;
  assign \new_[13099]_  = ~A302 & ~A301;
  assign \new_[13100]_  = A298 & \new_[13099]_ ;
  assign \new_[13101]_  = \new_[13100]_  & \new_[13095]_ ;
  assign \new_[13105]_  = ~A166 & ~A167;
  assign \new_[13106]_  = A170 & \new_[13105]_ ;
  assign \new_[13110]_  = A201 & ~A200;
  assign \new_[13111]_  = A199 & \new_[13110]_ ;
  assign \new_[13112]_  = \new_[13111]_  & \new_[13106]_ ;
  assign \new_[13116]_  = ~A268 & ~A266;
  assign \new_[13117]_  = A202 & \new_[13116]_ ;
  assign \new_[13121]_  = A299 & ~A298;
  assign \new_[13122]_  = ~A269 & \new_[13121]_ ;
  assign \new_[13123]_  = \new_[13122]_  & \new_[13117]_ ;
  assign \new_[13127]_  = ~A166 & ~A167;
  assign \new_[13128]_  = A170 & \new_[13127]_ ;
  assign \new_[13132]_  = A201 & ~A200;
  assign \new_[13133]_  = A199 & \new_[13132]_ ;
  assign \new_[13134]_  = \new_[13133]_  & \new_[13128]_ ;
  assign \new_[13138]_  = ~A268 & ~A266;
  assign \new_[13139]_  = A203 & \new_[13138]_ ;
  assign \new_[13143]_  = A299 & ~A298;
  assign \new_[13144]_  = ~A269 & \new_[13143]_ ;
  assign \new_[13145]_  = \new_[13144]_  & \new_[13139]_ ;
  assign \new_[13149]_  = ~A166 & ~A167;
  assign \new_[13150]_  = A170 & \new_[13149]_ ;
  assign \new_[13154]_  = A265 & ~A200;
  assign \new_[13155]_  = ~A199 & \new_[13154]_ ;
  assign \new_[13156]_  = \new_[13155]_  & \new_[13150]_ ;
  assign \new_[13160]_  = A268 & A267;
  assign \new_[13161]_  = ~A266 & \new_[13160]_ ;
  assign \new_[13165]_  = ~A302 & ~A301;
  assign \new_[13166]_  = A298 & \new_[13165]_ ;
  assign \new_[13167]_  = \new_[13166]_  & \new_[13161]_ ;
  assign \new_[13171]_  = ~A166 & ~A167;
  assign \new_[13172]_  = A170 & \new_[13171]_ ;
  assign \new_[13176]_  = A265 & ~A200;
  assign \new_[13177]_  = ~A199 & \new_[13176]_ ;
  assign \new_[13178]_  = \new_[13177]_  & \new_[13172]_ ;
  assign \new_[13182]_  = A269 & A267;
  assign \new_[13183]_  = ~A266 & \new_[13182]_ ;
  assign \new_[13187]_  = ~A302 & ~A301;
  assign \new_[13188]_  = A298 & \new_[13187]_ ;
  assign \new_[13189]_  = \new_[13188]_  & \new_[13183]_ ;
  assign \new_[13193]_  = A167 & ~A168;
  assign \new_[13194]_  = A169 & \new_[13193]_ ;
  assign \new_[13198]_  = A200 & A199;
  assign \new_[13199]_  = ~A166 & \new_[13198]_ ;
  assign \new_[13200]_  = \new_[13199]_  & \new_[13194]_ ;
  assign \new_[13204]_  = A267 & ~A266;
  assign \new_[13205]_  = A265 & \new_[13204]_ ;
  assign \new_[13209]_  = ~A300 & A298;
  assign \new_[13210]_  = A268 & \new_[13209]_ ;
  assign \new_[13211]_  = \new_[13210]_  & \new_[13205]_ ;
  assign \new_[13215]_  = A167 & ~A168;
  assign \new_[13216]_  = A169 & \new_[13215]_ ;
  assign \new_[13220]_  = A200 & A199;
  assign \new_[13221]_  = ~A166 & \new_[13220]_ ;
  assign \new_[13222]_  = \new_[13221]_  & \new_[13216]_ ;
  assign \new_[13226]_  = A267 & ~A266;
  assign \new_[13227]_  = A265 & \new_[13226]_ ;
  assign \new_[13231]_  = A299 & A298;
  assign \new_[13232]_  = A268 & \new_[13231]_ ;
  assign \new_[13233]_  = \new_[13232]_  & \new_[13227]_ ;
  assign \new_[13237]_  = A167 & ~A168;
  assign \new_[13238]_  = A169 & \new_[13237]_ ;
  assign \new_[13242]_  = A200 & A199;
  assign \new_[13243]_  = ~A166 & \new_[13242]_ ;
  assign \new_[13244]_  = \new_[13243]_  & \new_[13238]_ ;
  assign \new_[13248]_  = A267 & ~A266;
  assign \new_[13249]_  = A265 & \new_[13248]_ ;
  assign \new_[13253]_  = ~A299 & ~A298;
  assign \new_[13254]_  = A268 & \new_[13253]_ ;
  assign \new_[13255]_  = \new_[13254]_  & \new_[13249]_ ;
  assign \new_[13259]_  = A167 & ~A168;
  assign \new_[13260]_  = A169 & \new_[13259]_ ;
  assign \new_[13264]_  = A200 & A199;
  assign \new_[13265]_  = ~A166 & \new_[13264]_ ;
  assign \new_[13266]_  = \new_[13265]_  & \new_[13260]_ ;
  assign \new_[13270]_  = A267 & ~A266;
  assign \new_[13271]_  = A265 & \new_[13270]_ ;
  assign \new_[13275]_  = ~A300 & A298;
  assign \new_[13276]_  = A269 & \new_[13275]_ ;
  assign \new_[13277]_  = \new_[13276]_  & \new_[13271]_ ;
  assign \new_[13281]_  = A167 & ~A168;
  assign \new_[13282]_  = A169 & \new_[13281]_ ;
  assign \new_[13286]_  = A200 & A199;
  assign \new_[13287]_  = ~A166 & \new_[13286]_ ;
  assign \new_[13288]_  = \new_[13287]_  & \new_[13282]_ ;
  assign \new_[13292]_  = A267 & ~A266;
  assign \new_[13293]_  = A265 & \new_[13292]_ ;
  assign \new_[13297]_  = A299 & A298;
  assign \new_[13298]_  = A269 & \new_[13297]_ ;
  assign \new_[13299]_  = \new_[13298]_  & \new_[13293]_ ;
  assign \new_[13303]_  = A167 & ~A168;
  assign \new_[13304]_  = A169 & \new_[13303]_ ;
  assign \new_[13308]_  = A200 & A199;
  assign \new_[13309]_  = ~A166 & \new_[13308]_ ;
  assign \new_[13310]_  = \new_[13309]_  & \new_[13304]_ ;
  assign \new_[13314]_  = A267 & ~A266;
  assign \new_[13315]_  = A265 & \new_[13314]_ ;
  assign \new_[13319]_  = ~A299 & ~A298;
  assign \new_[13320]_  = A269 & \new_[13319]_ ;
  assign \new_[13321]_  = \new_[13320]_  & \new_[13315]_ ;
  assign \new_[13325]_  = A167 & ~A168;
  assign \new_[13326]_  = A169 & \new_[13325]_ ;
  assign \new_[13330]_  = A200 & ~A199;
  assign \new_[13331]_  = ~A166 & \new_[13330]_ ;
  assign \new_[13332]_  = \new_[13331]_  & \new_[13326]_ ;
  assign \new_[13336]_  = A298 & A266;
  assign \new_[13337]_  = A265 & \new_[13336]_ ;
  assign \new_[13341]_  = A301 & A300;
  assign \new_[13342]_  = ~A299 & \new_[13341]_ ;
  assign \new_[13343]_  = \new_[13342]_  & \new_[13337]_ ;
  assign \new_[13347]_  = A167 & ~A168;
  assign \new_[13348]_  = A169 & \new_[13347]_ ;
  assign \new_[13352]_  = A200 & ~A199;
  assign \new_[13353]_  = ~A166 & \new_[13352]_ ;
  assign \new_[13354]_  = \new_[13353]_  & \new_[13348]_ ;
  assign \new_[13358]_  = A298 & A266;
  assign \new_[13359]_  = A265 & \new_[13358]_ ;
  assign \new_[13363]_  = A302 & A300;
  assign \new_[13364]_  = ~A299 & \new_[13363]_ ;
  assign \new_[13365]_  = \new_[13364]_  & \new_[13359]_ ;
  assign \new_[13369]_  = A167 & ~A168;
  assign \new_[13370]_  = A169 & \new_[13369]_ ;
  assign \new_[13374]_  = A200 & ~A199;
  assign \new_[13375]_  = ~A166 & \new_[13374]_ ;
  assign \new_[13376]_  = \new_[13375]_  & \new_[13370]_ ;
  assign \new_[13380]_  = A298 & ~A267;
  assign \new_[13381]_  = ~A266 & \new_[13380]_ ;
  assign \new_[13385]_  = A301 & A300;
  assign \new_[13386]_  = ~A299 & \new_[13385]_ ;
  assign \new_[13387]_  = \new_[13386]_  & \new_[13381]_ ;
  assign \new_[13391]_  = A167 & ~A168;
  assign \new_[13392]_  = A169 & \new_[13391]_ ;
  assign \new_[13396]_  = A200 & ~A199;
  assign \new_[13397]_  = ~A166 & \new_[13396]_ ;
  assign \new_[13398]_  = \new_[13397]_  & \new_[13392]_ ;
  assign \new_[13402]_  = A298 & ~A267;
  assign \new_[13403]_  = ~A266 & \new_[13402]_ ;
  assign \new_[13407]_  = A302 & A300;
  assign \new_[13408]_  = ~A299 & \new_[13407]_ ;
  assign \new_[13409]_  = \new_[13408]_  & \new_[13403]_ ;
  assign \new_[13413]_  = A167 & ~A168;
  assign \new_[13414]_  = A169 & \new_[13413]_ ;
  assign \new_[13418]_  = A200 & ~A199;
  assign \new_[13419]_  = ~A166 & \new_[13418]_ ;
  assign \new_[13420]_  = \new_[13419]_  & \new_[13414]_ ;
  assign \new_[13424]_  = A298 & ~A266;
  assign \new_[13425]_  = ~A265 & \new_[13424]_ ;
  assign \new_[13429]_  = A301 & A300;
  assign \new_[13430]_  = ~A299 & \new_[13429]_ ;
  assign \new_[13431]_  = \new_[13430]_  & \new_[13425]_ ;
  assign \new_[13435]_  = A167 & ~A168;
  assign \new_[13436]_  = A169 & \new_[13435]_ ;
  assign \new_[13440]_  = A200 & ~A199;
  assign \new_[13441]_  = ~A166 & \new_[13440]_ ;
  assign \new_[13442]_  = \new_[13441]_  & \new_[13436]_ ;
  assign \new_[13446]_  = A298 & ~A266;
  assign \new_[13447]_  = ~A265 & \new_[13446]_ ;
  assign \new_[13451]_  = A302 & A300;
  assign \new_[13452]_  = ~A299 & \new_[13451]_ ;
  assign \new_[13453]_  = \new_[13452]_  & \new_[13447]_ ;
  assign \new_[13457]_  = A167 & ~A168;
  assign \new_[13458]_  = A169 & \new_[13457]_ ;
  assign \new_[13462]_  = ~A202 & ~A200;
  assign \new_[13463]_  = ~A166 & \new_[13462]_ ;
  assign \new_[13464]_  = \new_[13463]_  & \new_[13458]_ ;
  assign \new_[13468]_  = A266 & ~A265;
  assign \new_[13469]_  = ~A203 & \new_[13468]_ ;
  assign \new_[13473]_  = ~A302 & ~A301;
  assign \new_[13474]_  = A298 & \new_[13473]_ ;
  assign \new_[13475]_  = \new_[13474]_  & \new_[13469]_ ;
  assign \new_[13479]_  = A167 & ~A168;
  assign \new_[13480]_  = A169 & \new_[13479]_ ;
  assign \new_[13484]_  = ~A201 & ~A200;
  assign \new_[13485]_  = ~A166 & \new_[13484]_ ;
  assign \new_[13486]_  = \new_[13485]_  & \new_[13480]_ ;
  assign \new_[13490]_  = A267 & ~A266;
  assign \new_[13491]_  = A265 & \new_[13490]_ ;
  assign \new_[13495]_  = ~A300 & A298;
  assign \new_[13496]_  = A268 & \new_[13495]_ ;
  assign \new_[13497]_  = \new_[13496]_  & \new_[13491]_ ;
  assign \new_[13501]_  = A167 & ~A168;
  assign \new_[13502]_  = A169 & \new_[13501]_ ;
  assign \new_[13506]_  = ~A201 & ~A200;
  assign \new_[13507]_  = ~A166 & \new_[13506]_ ;
  assign \new_[13508]_  = \new_[13507]_  & \new_[13502]_ ;
  assign \new_[13512]_  = A267 & ~A266;
  assign \new_[13513]_  = A265 & \new_[13512]_ ;
  assign \new_[13517]_  = A299 & A298;
  assign \new_[13518]_  = A268 & \new_[13517]_ ;
  assign \new_[13519]_  = \new_[13518]_  & \new_[13513]_ ;
  assign \new_[13523]_  = A167 & ~A168;
  assign \new_[13524]_  = A169 & \new_[13523]_ ;
  assign \new_[13528]_  = ~A201 & ~A200;
  assign \new_[13529]_  = ~A166 & \new_[13528]_ ;
  assign \new_[13530]_  = \new_[13529]_  & \new_[13524]_ ;
  assign \new_[13534]_  = A267 & ~A266;
  assign \new_[13535]_  = A265 & \new_[13534]_ ;
  assign \new_[13539]_  = ~A299 & ~A298;
  assign \new_[13540]_  = A268 & \new_[13539]_ ;
  assign \new_[13541]_  = \new_[13540]_  & \new_[13535]_ ;
  assign \new_[13545]_  = A167 & ~A168;
  assign \new_[13546]_  = A169 & \new_[13545]_ ;
  assign \new_[13550]_  = ~A201 & ~A200;
  assign \new_[13551]_  = ~A166 & \new_[13550]_ ;
  assign \new_[13552]_  = \new_[13551]_  & \new_[13546]_ ;
  assign \new_[13556]_  = A267 & ~A266;
  assign \new_[13557]_  = A265 & \new_[13556]_ ;
  assign \new_[13561]_  = ~A300 & A298;
  assign \new_[13562]_  = A269 & \new_[13561]_ ;
  assign \new_[13563]_  = \new_[13562]_  & \new_[13557]_ ;
  assign \new_[13567]_  = A167 & ~A168;
  assign \new_[13568]_  = A169 & \new_[13567]_ ;
  assign \new_[13572]_  = ~A201 & ~A200;
  assign \new_[13573]_  = ~A166 & \new_[13572]_ ;
  assign \new_[13574]_  = \new_[13573]_  & \new_[13568]_ ;
  assign \new_[13578]_  = A267 & ~A266;
  assign \new_[13579]_  = A265 & \new_[13578]_ ;
  assign \new_[13583]_  = A299 & A298;
  assign \new_[13584]_  = A269 & \new_[13583]_ ;
  assign \new_[13585]_  = \new_[13584]_  & \new_[13579]_ ;
  assign \new_[13589]_  = A167 & ~A168;
  assign \new_[13590]_  = A169 & \new_[13589]_ ;
  assign \new_[13594]_  = ~A201 & ~A200;
  assign \new_[13595]_  = ~A166 & \new_[13594]_ ;
  assign \new_[13596]_  = \new_[13595]_  & \new_[13590]_ ;
  assign \new_[13600]_  = A267 & ~A266;
  assign \new_[13601]_  = A265 & \new_[13600]_ ;
  assign \new_[13605]_  = ~A299 & ~A298;
  assign \new_[13606]_  = A269 & \new_[13605]_ ;
  assign \new_[13607]_  = \new_[13606]_  & \new_[13601]_ ;
  assign \new_[13611]_  = A167 & ~A168;
  assign \new_[13612]_  = A169 & \new_[13611]_ ;
  assign \new_[13616]_  = ~A200 & A199;
  assign \new_[13617]_  = ~A166 & \new_[13616]_ ;
  assign \new_[13618]_  = \new_[13617]_  & \new_[13612]_ ;
  assign \new_[13622]_  = A265 & A202;
  assign \new_[13623]_  = A201 & \new_[13622]_ ;
  assign \new_[13627]_  = A299 & ~A298;
  assign \new_[13628]_  = A266 & \new_[13627]_ ;
  assign \new_[13629]_  = \new_[13628]_  & \new_[13623]_ ;
  assign \new_[13633]_  = A167 & ~A168;
  assign \new_[13634]_  = A169 & \new_[13633]_ ;
  assign \new_[13638]_  = ~A200 & A199;
  assign \new_[13639]_  = ~A166 & \new_[13638]_ ;
  assign \new_[13640]_  = \new_[13639]_  & \new_[13634]_ ;
  assign \new_[13644]_  = ~A266 & A202;
  assign \new_[13645]_  = A201 & \new_[13644]_ ;
  assign \new_[13649]_  = A299 & ~A298;
  assign \new_[13650]_  = ~A267 & \new_[13649]_ ;
  assign \new_[13651]_  = \new_[13650]_  & \new_[13645]_ ;
  assign \new_[13655]_  = A167 & ~A168;
  assign \new_[13656]_  = A169 & \new_[13655]_ ;
  assign \new_[13660]_  = ~A200 & A199;
  assign \new_[13661]_  = ~A166 & \new_[13660]_ ;
  assign \new_[13662]_  = \new_[13661]_  & \new_[13656]_ ;
  assign \new_[13666]_  = ~A265 & A202;
  assign \new_[13667]_  = A201 & \new_[13666]_ ;
  assign \new_[13671]_  = A299 & ~A298;
  assign \new_[13672]_  = ~A266 & \new_[13671]_ ;
  assign \new_[13673]_  = \new_[13672]_  & \new_[13667]_ ;
  assign \new_[13677]_  = A167 & ~A168;
  assign \new_[13678]_  = A169 & \new_[13677]_ ;
  assign \new_[13682]_  = ~A200 & A199;
  assign \new_[13683]_  = ~A166 & \new_[13682]_ ;
  assign \new_[13684]_  = \new_[13683]_  & \new_[13678]_ ;
  assign \new_[13688]_  = A265 & A203;
  assign \new_[13689]_  = A201 & \new_[13688]_ ;
  assign \new_[13693]_  = A299 & ~A298;
  assign \new_[13694]_  = A266 & \new_[13693]_ ;
  assign \new_[13695]_  = \new_[13694]_  & \new_[13689]_ ;
  assign \new_[13699]_  = A167 & ~A168;
  assign \new_[13700]_  = A169 & \new_[13699]_ ;
  assign \new_[13704]_  = ~A200 & A199;
  assign \new_[13705]_  = ~A166 & \new_[13704]_ ;
  assign \new_[13706]_  = \new_[13705]_  & \new_[13700]_ ;
  assign \new_[13710]_  = ~A266 & A203;
  assign \new_[13711]_  = A201 & \new_[13710]_ ;
  assign \new_[13715]_  = A299 & ~A298;
  assign \new_[13716]_  = ~A267 & \new_[13715]_ ;
  assign \new_[13717]_  = \new_[13716]_  & \new_[13711]_ ;
  assign \new_[13721]_  = A167 & ~A168;
  assign \new_[13722]_  = A169 & \new_[13721]_ ;
  assign \new_[13726]_  = ~A200 & A199;
  assign \new_[13727]_  = ~A166 & \new_[13726]_ ;
  assign \new_[13728]_  = \new_[13727]_  & \new_[13722]_ ;
  assign \new_[13732]_  = ~A265 & A203;
  assign \new_[13733]_  = A201 & \new_[13732]_ ;
  assign \new_[13737]_  = A299 & ~A298;
  assign \new_[13738]_  = ~A266 & \new_[13737]_ ;
  assign \new_[13739]_  = \new_[13738]_  & \new_[13733]_ ;
  assign \new_[13743]_  = A167 & ~A168;
  assign \new_[13744]_  = A169 & \new_[13743]_ ;
  assign \new_[13748]_  = ~A200 & ~A199;
  assign \new_[13749]_  = ~A166 & \new_[13748]_ ;
  assign \new_[13750]_  = \new_[13749]_  & \new_[13744]_ ;
  assign \new_[13754]_  = A267 & ~A266;
  assign \new_[13755]_  = A265 & \new_[13754]_ ;
  assign \new_[13759]_  = ~A300 & A298;
  assign \new_[13760]_  = A268 & \new_[13759]_ ;
  assign \new_[13761]_  = \new_[13760]_  & \new_[13755]_ ;
  assign \new_[13765]_  = A167 & ~A168;
  assign \new_[13766]_  = A169 & \new_[13765]_ ;
  assign \new_[13770]_  = ~A200 & ~A199;
  assign \new_[13771]_  = ~A166 & \new_[13770]_ ;
  assign \new_[13772]_  = \new_[13771]_  & \new_[13766]_ ;
  assign \new_[13776]_  = A267 & ~A266;
  assign \new_[13777]_  = A265 & \new_[13776]_ ;
  assign \new_[13781]_  = A299 & A298;
  assign \new_[13782]_  = A268 & \new_[13781]_ ;
  assign \new_[13783]_  = \new_[13782]_  & \new_[13777]_ ;
  assign \new_[13787]_  = A167 & ~A168;
  assign \new_[13788]_  = A169 & \new_[13787]_ ;
  assign \new_[13792]_  = ~A200 & ~A199;
  assign \new_[13793]_  = ~A166 & \new_[13792]_ ;
  assign \new_[13794]_  = \new_[13793]_  & \new_[13788]_ ;
  assign \new_[13798]_  = A267 & ~A266;
  assign \new_[13799]_  = A265 & \new_[13798]_ ;
  assign \new_[13803]_  = ~A299 & ~A298;
  assign \new_[13804]_  = A268 & \new_[13803]_ ;
  assign \new_[13805]_  = \new_[13804]_  & \new_[13799]_ ;
  assign \new_[13809]_  = A167 & ~A168;
  assign \new_[13810]_  = A169 & \new_[13809]_ ;
  assign \new_[13814]_  = ~A200 & ~A199;
  assign \new_[13815]_  = ~A166 & \new_[13814]_ ;
  assign \new_[13816]_  = \new_[13815]_  & \new_[13810]_ ;
  assign \new_[13820]_  = A267 & ~A266;
  assign \new_[13821]_  = A265 & \new_[13820]_ ;
  assign \new_[13825]_  = ~A300 & A298;
  assign \new_[13826]_  = A269 & \new_[13825]_ ;
  assign \new_[13827]_  = \new_[13826]_  & \new_[13821]_ ;
  assign \new_[13831]_  = A167 & ~A168;
  assign \new_[13832]_  = A169 & \new_[13831]_ ;
  assign \new_[13836]_  = ~A200 & ~A199;
  assign \new_[13837]_  = ~A166 & \new_[13836]_ ;
  assign \new_[13838]_  = \new_[13837]_  & \new_[13832]_ ;
  assign \new_[13842]_  = A267 & ~A266;
  assign \new_[13843]_  = A265 & \new_[13842]_ ;
  assign \new_[13847]_  = A299 & A298;
  assign \new_[13848]_  = A269 & \new_[13847]_ ;
  assign \new_[13849]_  = \new_[13848]_  & \new_[13843]_ ;
  assign \new_[13853]_  = A167 & ~A168;
  assign \new_[13854]_  = A169 & \new_[13853]_ ;
  assign \new_[13858]_  = ~A200 & ~A199;
  assign \new_[13859]_  = ~A166 & \new_[13858]_ ;
  assign \new_[13860]_  = \new_[13859]_  & \new_[13854]_ ;
  assign \new_[13864]_  = A267 & ~A266;
  assign \new_[13865]_  = A265 & \new_[13864]_ ;
  assign \new_[13869]_  = ~A299 & ~A298;
  assign \new_[13870]_  = A269 & \new_[13869]_ ;
  assign \new_[13871]_  = \new_[13870]_  & \new_[13865]_ ;
  assign \new_[13875]_  = ~A167 & ~A168;
  assign \new_[13876]_  = A169 & \new_[13875]_ ;
  assign \new_[13880]_  = A200 & A199;
  assign \new_[13881]_  = A166 & \new_[13880]_ ;
  assign \new_[13882]_  = \new_[13881]_  & \new_[13876]_ ;
  assign \new_[13886]_  = A267 & ~A266;
  assign \new_[13887]_  = A265 & \new_[13886]_ ;
  assign \new_[13891]_  = ~A300 & A298;
  assign \new_[13892]_  = A268 & \new_[13891]_ ;
  assign \new_[13893]_  = \new_[13892]_  & \new_[13887]_ ;
  assign \new_[13897]_  = ~A167 & ~A168;
  assign \new_[13898]_  = A169 & \new_[13897]_ ;
  assign \new_[13902]_  = A200 & A199;
  assign \new_[13903]_  = A166 & \new_[13902]_ ;
  assign \new_[13904]_  = \new_[13903]_  & \new_[13898]_ ;
  assign \new_[13908]_  = A267 & ~A266;
  assign \new_[13909]_  = A265 & \new_[13908]_ ;
  assign \new_[13913]_  = A299 & A298;
  assign \new_[13914]_  = A268 & \new_[13913]_ ;
  assign \new_[13915]_  = \new_[13914]_  & \new_[13909]_ ;
  assign \new_[13919]_  = ~A167 & ~A168;
  assign \new_[13920]_  = A169 & \new_[13919]_ ;
  assign \new_[13924]_  = A200 & A199;
  assign \new_[13925]_  = A166 & \new_[13924]_ ;
  assign \new_[13926]_  = \new_[13925]_  & \new_[13920]_ ;
  assign \new_[13930]_  = A267 & ~A266;
  assign \new_[13931]_  = A265 & \new_[13930]_ ;
  assign \new_[13935]_  = ~A299 & ~A298;
  assign \new_[13936]_  = A268 & \new_[13935]_ ;
  assign \new_[13937]_  = \new_[13936]_  & \new_[13931]_ ;
  assign \new_[13941]_  = ~A167 & ~A168;
  assign \new_[13942]_  = A169 & \new_[13941]_ ;
  assign \new_[13946]_  = A200 & A199;
  assign \new_[13947]_  = A166 & \new_[13946]_ ;
  assign \new_[13948]_  = \new_[13947]_  & \new_[13942]_ ;
  assign \new_[13952]_  = A267 & ~A266;
  assign \new_[13953]_  = A265 & \new_[13952]_ ;
  assign \new_[13957]_  = ~A300 & A298;
  assign \new_[13958]_  = A269 & \new_[13957]_ ;
  assign \new_[13959]_  = \new_[13958]_  & \new_[13953]_ ;
  assign \new_[13963]_  = ~A167 & ~A168;
  assign \new_[13964]_  = A169 & \new_[13963]_ ;
  assign \new_[13968]_  = A200 & A199;
  assign \new_[13969]_  = A166 & \new_[13968]_ ;
  assign \new_[13970]_  = \new_[13969]_  & \new_[13964]_ ;
  assign \new_[13974]_  = A267 & ~A266;
  assign \new_[13975]_  = A265 & \new_[13974]_ ;
  assign \new_[13979]_  = A299 & A298;
  assign \new_[13980]_  = A269 & \new_[13979]_ ;
  assign \new_[13981]_  = \new_[13980]_  & \new_[13975]_ ;
  assign \new_[13985]_  = ~A167 & ~A168;
  assign \new_[13986]_  = A169 & \new_[13985]_ ;
  assign \new_[13990]_  = A200 & A199;
  assign \new_[13991]_  = A166 & \new_[13990]_ ;
  assign \new_[13992]_  = \new_[13991]_  & \new_[13986]_ ;
  assign \new_[13996]_  = A267 & ~A266;
  assign \new_[13997]_  = A265 & \new_[13996]_ ;
  assign \new_[14001]_  = ~A299 & ~A298;
  assign \new_[14002]_  = A269 & \new_[14001]_ ;
  assign \new_[14003]_  = \new_[14002]_  & \new_[13997]_ ;
  assign \new_[14007]_  = ~A167 & ~A168;
  assign \new_[14008]_  = A169 & \new_[14007]_ ;
  assign \new_[14012]_  = A200 & ~A199;
  assign \new_[14013]_  = A166 & \new_[14012]_ ;
  assign \new_[14014]_  = \new_[14013]_  & \new_[14008]_ ;
  assign \new_[14018]_  = A298 & A266;
  assign \new_[14019]_  = A265 & \new_[14018]_ ;
  assign \new_[14023]_  = A301 & A300;
  assign \new_[14024]_  = ~A299 & \new_[14023]_ ;
  assign \new_[14025]_  = \new_[14024]_  & \new_[14019]_ ;
  assign \new_[14029]_  = ~A167 & ~A168;
  assign \new_[14030]_  = A169 & \new_[14029]_ ;
  assign \new_[14034]_  = A200 & ~A199;
  assign \new_[14035]_  = A166 & \new_[14034]_ ;
  assign \new_[14036]_  = \new_[14035]_  & \new_[14030]_ ;
  assign \new_[14040]_  = A298 & A266;
  assign \new_[14041]_  = A265 & \new_[14040]_ ;
  assign \new_[14045]_  = A302 & A300;
  assign \new_[14046]_  = ~A299 & \new_[14045]_ ;
  assign \new_[14047]_  = \new_[14046]_  & \new_[14041]_ ;
  assign \new_[14051]_  = ~A167 & ~A168;
  assign \new_[14052]_  = A169 & \new_[14051]_ ;
  assign \new_[14056]_  = A200 & ~A199;
  assign \new_[14057]_  = A166 & \new_[14056]_ ;
  assign \new_[14058]_  = \new_[14057]_  & \new_[14052]_ ;
  assign \new_[14062]_  = A298 & ~A267;
  assign \new_[14063]_  = ~A266 & \new_[14062]_ ;
  assign \new_[14067]_  = A301 & A300;
  assign \new_[14068]_  = ~A299 & \new_[14067]_ ;
  assign \new_[14069]_  = \new_[14068]_  & \new_[14063]_ ;
  assign \new_[14073]_  = ~A167 & ~A168;
  assign \new_[14074]_  = A169 & \new_[14073]_ ;
  assign \new_[14078]_  = A200 & ~A199;
  assign \new_[14079]_  = A166 & \new_[14078]_ ;
  assign \new_[14080]_  = \new_[14079]_  & \new_[14074]_ ;
  assign \new_[14084]_  = A298 & ~A267;
  assign \new_[14085]_  = ~A266 & \new_[14084]_ ;
  assign \new_[14089]_  = A302 & A300;
  assign \new_[14090]_  = ~A299 & \new_[14089]_ ;
  assign \new_[14091]_  = \new_[14090]_  & \new_[14085]_ ;
  assign \new_[14095]_  = ~A167 & ~A168;
  assign \new_[14096]_  = A169 & \new_[14095]_ ;
  assign \new_[14100]_  = A200 & ~A199;
  assign \new_[14101]_  = A166 & \new_[14100]_ ;
  assign \new_[14102]_  = \new_[14101]_  & \new_[14096]_ ;
  assign \new_[14106]_  = A298 & ~A266;
  assign \new_[14107]_  = ~A265 & \new_[14106]_ ;
  assign \new_[14111]_  = A301 & A300;
  assign \new_[14112]_  = ~A299 & \new_[14111]_ ;
  assign \new_[14113]_  = \new_[14112]_  & \new_[14107]_ ;
  assign \new_[14117]_  = ~A167 & ~A168;
  assign \new_[14118]_  = A169 & \new_[14117]_ ;
  assign \new_[14122]_  = A200 & ~A199;
  assign \new_[14123]_  = A166 & \new_[14122]_ ;
  assign \new_[14124]_  = \new_[14123]_  & \new_[14118]_ ;
  assign \new_[14128]_  = A298 & ~A266;
  assign \new_[14129]_  = ~A265 & \new_[14128]_ ;
  assign \new_[14133]_  = A302 & A300;
  assign \new_[14134]_  = ~A299 & \new_[14133]_ ;
  assign \new_[14135]_  = \new_[14134]_  & \new_[14129]_ ;
  assign \new_[14139]_  = ~A167 & ~A168;
  assign \new_[14140]_  = A169 & \new_[14139]_ ;
  assign \new_[14144]_  = ~A202 & ~A200;
  assign \new_[14145]_  = A166 & \new_[14144]_ ;
  assign \new_[14146]_  = \new_[14145]_  & \new_[14140]_ ;
  assign \new_[14150]_  = A266 & ~A265;
  assign \new_[14151]_  = ~A203 & \new_[14150]_ ;
  assign \new_[14155]_  = ~A302 & ~A301;
  assign \new_[14156]_  = A298 & \new_[14155]_ ;
  assign \new_[14157]_  = \new_[14156]_  & \new_[14151]_ ;
  assign \new_[14161]_  = ~A167 & ~A168;
  assign \new_[14162]_  = A169 & \new_[14161]_ ;
  assign \new_[14166]_  = ~A201 & ~A200;
  assign \new_[14167]_  = A166 & \new_[14166]_ ;
  assign \new_[14168]_  = \new_[14167]_  & \new_[14162]_ ;
  assign \new_[14172]_  = A267 & ~A266;
  assign \new_[14173]_  = A265 & \new_[14172]_ ;
  assign \new_[14177]_  = ~A300 & A298;
  assign \new_[14178]_  = A268 & \new_[14177]_ ;
  assign \new_[14179]_  = \new_[14178]_  & \new_[14173]_ ;
  assign \new_[14183]_  = ~A167 & ~A168;
  assign \new_[14184]_  = A169 & \new_[14183]_ ;
  assign \new_[14188]_  = ~A201 & ~A200;
  assign \new_[14189]_  = A166 & \new_[14188]_ ;
  assign \new_[14190]_  = \new_[14189]_  & \new_[14184]_ ;
  assign \new_[14194]_  = A267 & ~A266;
  assign \new_[14195]_  = A265 & \new_[14194]_ ;
  assign \new_[14199]_  = A299 & A298;
  assign \new_[14200]_  = A268 & \new_[14199]_ ;
  assign \new_[14201]_  = \new_[14200]_  & \new_[14195]_ ;
  assign \new_[14205]_  = ~A167 & ~A168;
  assign \new_[14206]_  = A169 & \new_[14205]_ ;
  assign \new_[14210]_  = ~A201 & ~A200;
  assign \new_[14211]_  = A166 & \new_[14210]_ ;
  assign \new_[14212]_  = \new_[14211]_  & \new_[14206]_ ;
  assign \new_[14216]_  = A267 & ~A266;
  assign \new_[14217]_  = A265 & \new_[14216]_ ;
  assign \new_[14221]_  = ~A299 & ~A298;
  assign \new_[14222]_  = A268 & \new_[14221]_ ;
  assign \new_[14223]_  = \new_[14222]_  & \new_[14217]_ ;
  assign \new_[14227]_  = ~A167 & ~A168;
  assign \new_[14228]_  = A169 & \new_[14227]_ ;
  assign \new_[14232]_  = ~A201 & ~A200;
  assign \new_[14233]_  = A166 & \new_[14232]_ ;
  assign \new_[14234]_  = \new_[14233]_  & \new_[14228]_ ;
  assign \new_[14238]_  = A267 & ~A266;
  assign \new_[14239]_  = A265 & \new_[14238]_ ;
  assign \new_[14243]_  = ~A300 & A298;
  assign \new_[14244]_  = A269 & \new_[14243]_ ;
  assign \new_[14245]_  = \new_[14244]_  & \new_[14239]_ ;
  assign \new_[14249]_  = ~A167 & ~A168;
  assign \new_[14250]_  = A169 & \new_[14249]_ ;
  assign \new_[14254]_  = ~A201 & ~A200;
  assign \new_[14255]_  = A166 & \new_[14254]_ ;
  assign \new_[14256]_  = \new_[14255]_  & \new_[14250]_ ;
  assign \new_[14260]_  = A267 & ~A266;
  assign \new_[14261]_  = A265 & \new_[14260]_ ;
  assign \new_[14265]_  = A299 & A298;
  assign \new_[14266]_  = A269 & \new_[14265]_ ;
  assign \new_[14267]_  = \new_[14266]_  & \new_[14261]_ ;
  assign \new_[14271]_  = ~A167 & ~A168;
  assign \new_[14272]_  = A169 & \new_[14271]_ ;
  assign \new_[14276]_  = ~A201 & ~A200;
  assign \new_[14277]_  = A166 & \new_[14276]_ ;
  assign \new_[14278]_  = \new_[14277]_  & \new_[14272]_ ;
  assign \new_[14282]_  = A267 & ~A266;
  assign \new_[14283]_  = A265 & \new_[14282]_ ;
  assign \new_[14287]_  = ~A299 & ~A298;
  assign \new_[14288]_  = A269 & \new_[14287]_ ;
  assign \new_[14289]_  = \new_[14288]_  & \new_[14283]_ ;
  assign \new_[14293]_  = ~A167 & ~A168;
  assign \new_[14294]_  = A169 & \new_[14293]_ ;
  assign \new_[14298]_  = ~A200 & A199;
  assign \new_[14299]_  = A166 & \new_[14298]_ ;
  assign \new_[14300]_  = \new_[14299]_  & \new_[14294]_ ;
  assign \new_[14304]_  = A265 & A202;
  assign \new_[14305]_  = A201 & \new_[14304]_ ;
  assign \new_[14309]_  = A299 & ~A298;
  assign \new_[14310]_  = A266 & \new_[14309]_ ;
  assign \new_[14311]_  = \new_[14310]_  & \new_[14305]_ ;
  assign \new_[14315]_  = ~A167 & ~A168;
  assign \new_[14316]_  = A169 & \new_[14315]_ ;
  assign \new_[14320]_  = ~A200 & A199;
  assign \new_[14321]_  = A166 & \new_[14320]_ ;
  assign \new_[14322]_  = \new_[14321]_  & \new_[14316]_ ;
  assign \new_[14326]_  = ~A266 & A202;
  assign \new_[14327]_  = A201 & \new_[14326]_ ;
  assign \new_[14331]_  = A299 & ~A298;
  assign \new_[14332]_  = ~A267 & \new_[14331]_ ;
  assign \new_[14333]_  = \new_[14332]_  & \new_[14327]_ ;
  assign \new_[14337]_  = ~A167 & ~A168;
  assign \new_[14338]_  = A169 & \new_[14337]_ ;
  assign \new_[14342]_  = ~A200 & A199;
  assign \new_[14343]_  = A166 & \new_[14342]_ ;
  assign \new_[14344]_  = \new_[14343]_  & \new_[14338]_ ;
  assign \new_[14348]_  = ~A265 & A202;
  assign \new_[14349]_  = A201 & \new_[14348]_ ;
  assign \new_[14353]_  = A299 & ~A298;
  assign \new_[14354]_  = ~A266 & \new_[14353]_ ;
  assign \new_[14355]_  = \new_[14354]_  & \new_[14349]_ ;
  assign \new_[14359]_  = ~A167 & ~A168;
  assign \new_[14360]_  = A169 & \new_[14359]_ ;
  assign \new_[14364]_  = ~A200 & A199;
  assign \new_[14365]_  = A166 & \new_[14364]_ ;
  assign \new_[14366]_  = \new_[14365]_  & \new_[14360]_ ;
  assign \new_[14370]_  = A265 & A203;
  assign \new_[14371]_  = A201 & \new_[14370]_ ;
  assign \new_[14375]_  = A299 & ~A298;
  assign \new_[14376]_  = A266 & \new_[14375]_ ;
  assign \new_[14377]_  = \new_[14376]_  & \new_[14371]_ ;
  assign \new_[14381]_  = ~A167 & ~A168;
  assign \new_[14382]_  = A169 & \new_[14381]_ ;
  assign \new_[14386]_  = ~A200 & A199;
  assign \new_[14387]_  = A166 & \new_[14386]_ ;
  assign \new_[14388]_  = \new_[14387]_  & \new_[14382]_ ;
  assign \new_[14392]_  = ~A266 & A203;
  assign \new_[14393]_  = A201 & \new_[14392]_ ;
  assign \new_[14397]_  = A299 & ~A298;
  assign \new_[14398]_  = ~A267 & \new_[14397]_ ;
  assign \new_[14399]_  = \new_[14398]_  & \new_[14393]_ ;
  assign \new_[14403]_  = ~A167 & ~A168;
  assign \new_[14404]_  = A169 & \new_[14403]_ ;
  assign \new_[14408]_  = ~A200 & A199;
  assign \new_[14409]_  = A166 & \new_[14408]_ ;
  assign \new_[14410]_  = \new_[14409]_  & \new_[14404]_ ;
  assign \new_[14414]_  = ~A265 & A203;
  assign \new_[14415]_  = A201 & \new_[14414]_ ;
  assign \new_[14419]_  = A299 & ~A298;
  assign \new_[14420]_  = ~A266 & \new_[14419]_ ;
  assign \new_[14421]_  = \new_[14420]_  & \new_[14415]_ ;
  assign \new_[14425]_  = ~A167 & ~A168;
  assign \new_[14426]_  = A169 & \new_[14425]_ ;
  assign \new_[14430]_  = ~A200 & ~A199;
  assign \new_[14431]_  = A166 & \new_[14430]_ ;
  assign \new_[14432]_  = \new_[14431]_  & \new_[14426]_ ;
  assign \new_[14436]_  = A267 & ~A266;
  assign \new_[14437]_  = A265 & \new_[14436]_ ;
  assign \new_[14441]_  = ~A300 & A298;
  assign \new_[14442]_  = A268 & \new_[14441]_ ;
  assign \new_[14443]_  = \new_[14442]_  & \new_[14437]_ ;
  assign \new_[14447]_  = ~A167 & ~A168;
  assign \new_[14448]_  = A169 & \new_[14447]_ ;
  assign \new_[14452]_  = ~A200 & ~A199;
  assign \new_[14453]_  = A166 & \new_[14452]_ ;
  assign \new_[14454]_  = \new_[14453]_  & \new_[14448]_ ;
  assign \new_[14458]_  = A267 & ~A266;
  assign \new_[14459]_  = A265 & \new_[14458]_ ;
  assign \new_[14463]_  = A299 & A298;
  assign \new_[14464]_  = A268 & \new_[14463]_ ;
  assign \new_[14465]_  = \new_[14464]_  & \new_[14459]_ ;
  assign \new_[14469]_  = ~A167 & ~A168;
  assign \new_[14470]_  = A169 & \new_[14469]_ ;
  assign \new_[14474]_  = ~A200 & ~A199;
  assign \new_[14475]_  = A166 & \new_[14474]_ ;
  assign \new_[14476]_  = \new_[14475]_  & \new_[14470]_ ;
  assign \new_[14480]_  = A267 & ~A266;
  assign \new_[14481]_  = A265 & \new_[14480]_ ;
  assign \new_[14485]_  = ~A299 & ~A298;
  assign \new_[14486]_  = A268 & \new_[14485]_ ;
  assign \new_[14487]_  = \new_[14486]_  & \new_[14481]_ ;
  assign \new_[14491]_  = ~A167 & ~A168;
  assign \new_[14492]_  = A169 & \new_[14491]_ ;
  assign \new_[14496]_  = ~A200 & ~A199;
  assign \new_[14497]_  = A166 & \new_[14496]_ ;
  assign \new_[14498]_  = \new_[14497]_  & \new_[14492]_ ;
  assign \new_[14502]_  = A267 & ~A266;
  assign \new_[14503]_  = A265 & \new_[14502]_ ;
  assign \new_[14507]_  = ~A300 & A298;
  assign \new_[14508]_  = A269 & \new_[14507]_ ;
  assign \new_[14509]_  = \new_[14508]_  & \new_[14503]_ ;
  assign \new_[14513]_  = ~A167 & ~A168;
  assign \new_[14514]_  = A169 & \new_[14513]_ ;
  assign \new_[14518]_  = ~A200 & ~A199;
  assign \new_[14519]_  = A166 & \new_[14518]_ ;
  assign \new_[14520]_  = \new_[14519]_  & \new_[14514]_ ;
  assign \new_[14524]_  = A267 & ~A266;
  assign \new_[14525]_  = A265 & \new_[14524]_ ;
  assign \new_[14529]_  = A299 & A298;
  assign \new_[14530]_  = A269 & \new_[14529]_ ;
  assign \new_[14531]_  = \new_[14530]_  & \new_[14525]_ ;
  assign \new_[14535]_  = ~A167 & ~A168;
  assign \new_[14536]_  = A169 & \new_[14535]_ ;
  assign \new_[14540]_  = ~A200 & ~A199;
  assign \new_[14541]_  = A166 & \new_[14540]_ ;
  assign \new_[14542]_  = \new_[14541]_  & \new_[14536]_ ;
  assign \new_[14546]_  = A267 & ~A266;
  assign \new_[14547]_  = A265 & \new_[14546]_ ;
  assign \new_[14551]_  = ~A299 & ~A298;
  assign \new_[14552]_  = A269 & \new_[14551]_ ;
  assign \new_[14553]_  = \new_[14552]_  & \new_[14547]_ ;
  assign \new_[14557]_  = ~A168 & A169;
  assign \new_[14558]_  = A170 & \new_[14557]_ ;
  assign \new_[14562]_  = A265 & A200;
  assign \new_[14563]_  = A199 & \new_[14562]_ ;
  assign \new_[14564]_  = \new_[14563]_  & \new_[14558]_ ;
  assign \new_[14568]_  = A268 & A267;
  assign \new_[14569]_  = ~A266 & \new_[14568]_ ;
  assign \new_[14573]_  = ~A302 & ~A301;
  assign \new_[14574]_  = A298 & \new_[14573]_ ;
  assign \new_[14575]_  = \new_[14574]_  & \new_[14569]_ ;
  assign \new_[14579]_  = ~A168 & A169;
  assign \new_[14580]_  = A170 & \new_[14579]_ ;
  assign \new_[14584]_  = A265 & A200;
  assign \new_[14585]_  = A199 & \new_[14584]_ ;
  assign \new_[14586]_  = \new_[14585]_  & \new_[14580]_ ;
  assign \new_[14590]_  = A269 & A267;
  assign \new_[14591]_  = ~A266 & \new_[14590]_ ;
  assign \new_[14595]_  = ~A302 & ~A301;
  assign \new_[14596]_  = A298 & \new_[14595]_ ;
  assign \new_[14597]_  = \new_[14596]_  & \new_[14591]_ ;
  assign \new_[14601]_  = ~A168 & A169;
  assign \new_[14602]_  = A170 & \new_[14601]_ ;
  assign \new_[14606]_  = ~A266 & A200;
  assign \new_[14607]_  = ~A199 & \new_[14606]_ ;
  assign \new_[14608]_  = \new_[14607]_  & \new_[14602]_ ;
  assign \new_[14612]_  = A298 & ~A269;
  assign \new_[14613]_  = ~A268 & \new_[14612]_ ;
  assign \new_[14617]_  = A301 & A300;
  assign \new_[14618]_  = ~A299 & \new_[14617]_ ;
  assign \new_[14619]_  = \new_[14618]_  & \new_[14613]_ ;
  assign \new_[14623]_  = ~A168 & A169;
  assign \new_[14624]_  = A170 & \new_[14623]_ ;
  assign \new_[14628]_  = ~A266 & A200;
  assign \new_[14629]_  = ~A199 & \new_[14628]_ ;
  assign \new_[14630]_  = \new_[14629]_  & \new_[14624]_ ;
  assign \new_[14634]_  = A298 & ~A269;
  assign \new_[14635]_  = ~A268 & \new_[14634]_ ;
  assign \new_[14639]_  = A302 & A300;
  assign \new_[14640]_  = ~A299 & \new_[14639]_ ;
  assign \new_[14641]_  = \new_[14640]_  & \new_[14635]_ ;
  assign \new_[14645]_  = ~A168 & A169;
  assign \new_[14646]_  = A170 & \new_[14645]_ ;
  assign \new_[14650]_  = ~A203 & ~A202;
  assign \new_[14651]_  = ~A200 & \new_[14650]_ ;
  assign \new_[14652]_  = \new_[14651]_  & \new_[14646]_ ;
  assign \new_[14656]_  = A267 & ~A266;
  assign \new_[14657]_  = A265 & \new_[14656]_ ;
  assign \new_[14661]_  = ~A300 & A298;
  assign \new_[14662]_  = A268 & \new_[14661]_ ;
  assign \new_[14663]_  = \new_[14662]_  & \new_[14657]_ ;
  assign \new_[14667]_  = ~A168 & A169;
  assign \new_[14668]_  = A170 & \new_[14667]_ ;
  assign \new_[14672]_  = ~A203 & ~A202;
  assign \new_[14673]_  = ~A200 & \new_[14672]_ ;
  assign \new_[14674]_  = \new_[14673]_  & \new_[14668]_ ;
  assign \new_[14678]_  = A267 & ~A266;
  assign \new_[14679]_  = A265 & \new_[14678]_ ;
  assign \new_[14683]_  = A299 & A298;
  assign \new_[14684]_  = A268 & \new_[14683]_ ;
  assign \new_[14685]_  = \new_[14684]_  & \new_[14679]_ ;
  assign \new_[14689]_  = ~A168 & A169;
  assign \new_[14690]_  = A170 & \new_[14689]_ ;
  assign \new_[14694]_  = ~A203 & ~A202;
  assign \new_[14695]_  = ~A200 & \new_[14694]_ ;
  assign \new_[14696]_  = \new_[14695]_  & \new_[14690]_ ;
  assign \new_[14700]_  = A267 & ~A266;
  assign \new_[14701]_  = A265 & \new_[14700]_ ;
  assign \new_[14705]_  = ~A299 & ~A298;
  assign \new_[14706]_  = A268 & \new_[14705]_ ;
  assign \new_[14707]_  = \new_[14706]_  & \new_[14701]_ ;
  assign \new_[14711]_  = ~A168 & A169;
  assign \new_[14712]_  = A170 & \new_[14711]_ ;
  assign \new_[14716]_  = ~A203 & ~A202;
  assign \new_[14717]_  = ~A200 & \new_[14716]_ ;
  assign \new_[14718]_  = \new_[14717]_  & \new_[14712]_ ;
  assign \new_[14722]_  = A267 & ~A266;
  assign \new_[14723]_  = A265 & \new_[14722]_ ;
  assign \new_[14727]_  = ~A300 & A298;
  assign \new_[14728]_  = A269 & \new_[14727]_ ;
  assign \new_[14729]_  = \new_[14728]_  & \new_[14723]_ ;
  assign \new_[14733]_  = ~A168 & A169;
  assign \new_[14734]_  = A170 & \new_[14733]_ ;
  assign \new_[14738]_  = ~A203 & ~A202;
  assign \new_[14739]_  = ~A200 & \new_[14738]_ ;
  assign \new_[14740]_  = \new_[14739]_  & \new_[14734]_ ;
  assign \new_[14744]_  = A267 & ~A266;
  assign \new_[14745]_  = A265 & \new_[14744]_ ;
  assign \new_[14749]_  = A299 & A298;
  assign \new_[14750]_  = A269 & \new_[14749]_ ;
  assign \new_[14751]_  = \new_[14750]_  & \new_[14745]_ ;
  assign \new_[14755]_  = ~A168 & A169;
  assign \new_[14756]_  = A170 & \new_[14755]_ ;
  assign \new_[14760]_  = ~A203 & ~A202;
  assign \new_[14761]_  = ~A200 & \new_[14760]_ ;
  assign \new_[14762]_  = \new_[14761]_  & \new_[14756]_ ;
  assign \new_[14766]_  = A267 & ~A266;
  assign \new_[14767]_  = A265 & \new_[14766]_ ;
  assign \new_[14771]_  = ~A299 & ~A298;
  assign \new_[14772]_  = A269 & \new_[14771]_ ;
  assign \new_[14773]_  = \new_[14772]_  & \new_[14767]_ ;
  assign \new_[14777]_  = ~A168 & A169;
  assign \new_[14778]_  = A170 & \new_[14777]_ ;
  assign \new_[14782]_  = A265 & ~A201;
  assign \new_[14783]_  = ~A200 & \new_[14782]_ ;
  assign \new_[14784]_  = \new_[14783]_  & \new_[14778]_ ;
  assign \new_[14788]_  = A268 & A267;
  assign \new_[14789]_  = ~A266 & \new_[14788]_ ;
  assign \new_[14793]_  = ~A302 & ~A301;
  assign \new_[14794]_  = A298 & \new_[14793]_ ;
  assign \new_[14795]_  = \new_[14794]_  & \new_[14789]_ ;
  assign \new_[14799]_  = ~A168 & A169;
  assign \new_[14800]_  = A170 & \new_[14799]_ ;
  assign \new_[14804]_  = A265 & ~A201;
  assign \new_[14805]_  = ~A200 & \new_[14804]_ ;
  assign \new_[14806]_  = \new_[14805]_  & \new_[14800]_ ;
  assign \new_[14810]_  = A269 & A267;
  assign \new_[14811]_  = ~A266 & \new_[14810]_ ;
  assign \new_[14815]_  = ~A302 & ~A301;
  assign \new_[14816]_  = A298 & \new_[14815]_ ;
  assign \new_[14817]_  = \new_[14816]_  & \new_[14811]_ ;
  assign \new_[14821]_  = ~A168 & A169;
  assign \new_[14822]_  = A170 & \new_[14821]_ ;
  assign \new_[14826]_  = A201 & ~A200;
  assign \new_[14827]_  = A199 & \new_[14826]_ ;
  assign \new_[14828]_  = \new_[14827]_  & \new_[14822]_ ;
  assign \new_[14832]_  = ~A268 & ~A266;
  assign \new_[14833]_  = A202 & \new_[14832]_ ;
  assign \new_[14837]_  = A299 & ~A298;
  assign \new_[14838]_  = ~A269 & \new_[14837]_ ;
  assign \new_[14839]_  = \new_[14838]_  & \new_[14833]_ ;
  assign \new_[14843]_  = ~A168 & A169;
  assign \new_[14844]_  = A170 & \new_[14843]_ ;
  assign \new_[14848]_  = A201 & ~A200;
  assign \new_[14849]_  = A199 & \new_[14848]_ ;
  assign \new_[14850]_  = \new_[14849]_  & \new_[14844]_ ;
  assign \new_[14854]_  = ~A268 & ~A266;
  assign \new_[14855]_  = A203 & \new_[14854]_ ;
  assign \new_[14859]_  = A299 & ~A298;
  assign \new_[14860]_  = ~A269 & \new_[14859]_ ;
  assign \new_[14861]_  = \new_[14860]_  & \new_[14855]_ ;
  assign \new_[14865]_  = ~A168 & A169;
  assign \new_[14866]_  = A170 & \new_[14865]_ ;
  assign \new_[14870]_  = A265 & ~A200;
  assign \new_[14871]_  = ~A199 & \new_[14870]_ ;
  assign \new_[14872]_  = \new_[14871]_  & \new_[14866]_ ;
  assign \new_[14876]_  = A268 & A267;
  assign \new_[14877]_  = ~A266 & \new_[14876]_ ;
  assign \new_[14881]_  = ~A302 & ~A301;
  assign \new_[14882]_  = A298 & \new_[14881]_ ;
  assign \new_[14883]_  = \new_[14882]_  & \new_[14877]_ ;
  assign \new_[14887]_  = ~A168 & A169;
  assign \new_[14888]_  = A170 & \new_[14887]_ ;
  assign \new_[14892]_  = A265 & ~A200;
  assign \new_[14893]_  = ~A199 & \new_[14892]_ ;
  assign \new_[14894]_  = \new_[14893]_  & \new_[14888]_ ;
  assign \new_[14898]_  = A269 & A267;
  assign \new_[14899]_  = ~A266 & \new_[14898]_ ;
  assign \new_[14903]_  = ~A302 & ~A301;
  assign \new_[14904]_  = A298 & \new_[14903]_ ;
  assign \new_[14905]_  = \new_[14904]_  & \new_[14899]_ ;
  assign \new_[14909]_  = A167 & A169;
  assign \new_[14910]_  = ~A170 & \new_[14909]_ ;
  assign \new_[14914]_  = A200 & A199;
  assign \new_[14915]_  = A166 & \new_[14914]_ ;
  assign \new_[14916]_  = \new_[14915]_  & \new_[14910]_ ;
  assign \new_[14920]_  = A298 & A266;
  assign \new_[14921]_  = A265 & \new_[14920]_ ;
  assign \new_[14925]_  = A301 & A300;
  assign \new_[14926]_  = ~A299 & \new_[14925]_ ;
  assign \new_[14927]_  = \new_[14926]_  & \new_[14921]_ ;
  assign \new_[14931]_  = A167 & A169;
  assign \new_[14932]_  = ~A170 & \new_[14931]_ ;
  assign \new_[14936]_  = A200 & A199;
  assign \new_[14937]_  = A166 & \new_[14936]_ ;
  assign \new_[14938]_  = \new_[14937]_  & \new_[14932]_ ;
  assign \new_[14942]_  = A298 & A266;
  assign \new_[14943]_  = A265 & \new_[14942]_ ;
  assign \new_[14947]_  = A302 & A300;
  assign \new_[14948]_  = ~A299 & \new_[14947]_ ;
  assign \new_[14949]_  = \new_[14948]_  & \new_[14943]_ ;
  assign \new_[14953]_  = A167 & A169;
  assign \new_[14954]_  = ~A170 & \new_[14953]_ ;
  assign \new_[14958]_  = A200 & A199;
  assign \new_[14959]_  = A166 & \new_[14958]_ ;
  assign \new_[14960]_  = \new_[14959]_  & \new_[14954]_ ;
  assign \new_[14964]_  = A298 & ~A267;
  assign \new_[14965]_  = ~A266 & \new_[14964]_ ;
  assign \new_[14969]_  = A301 & A300;
  assign \new_[14970]_  = ~A299 & \new_[14969]_ ;
  assign \new_[14971]_  = \new_[14970]_  & \new_[14965]_ ;
  assign \new_[14975]_  = A167 & A169;
  assign \new_[14976]_  = ~A170 & \new_[14975]_ ;
  assign \new_[14980]_  = A200 & A199;
  assign \new_[14981]_  = A166 & \new_[14980]_ ;
  assign \new_[14982]_  = \new_[14981]_  & \new_[14976]_ ;
  assign \new_[14986]_  = A298 & ~A267;
  assign \new_[14987]_  = ~A266 & \new_[14986]_ ;
  assign \new_[14991]_  = A302 & A300;
  assign \new_[14992]_  = ~A299 & \new_[14991]_ ;
  assign \new_[14993]_  = \new_[14992]_  & \new_[14987]_ ;
  assign \new_[14997]_  = A167 & A169;
  assign \new_[14998]_  = ~A170 & \new_[14997]_ ;
  assign \new_[15002]_  = A200 & A199;
  assign \new_[15003]_  = A166 & \new_[15002]_ ;
  assign \new_[15004]_  = \new_[15003]_  & \new_[14998]_ ;
  assign \new_[15008]_  = A298 & ~A266;
  assign \new_[15009]_  = ~A265 & \new_[15008]_ ;
  assign \new_[15013]_  = A301 & A300;
  assign \new_[15014]_  = ~A299 & \new_[15013]_ ;
  assign \new_[15015]_  = \new_[15014]_  & \new_[15009]_ ;
  assign \new_[15019]_  = A167 & A169;
  assign \new_[15020]_  = ~A170 & \new_[15019]_ ;
  assign \new_[15024]_  = A200 & A199;
  assign \new_[15025]_  = A166 & \new_[15024]_ ;
  assign \new_[15026]_  = \new_[15025]_  & \new_[15020]_ ;
  assign \new_[15030]_  = A298 & ~A266;
  assign \new_[15031]_  = ~A265 & \new_[15030]_ ;
  assign \new_[15035]_  = A302 & A300;
  assign \new_[15036]_  = ~A299 & \new_[15035]_ ;
  assign \new_[15037]_  = \new_[15036]_  & \new_[15031]_ ;
  assign \new_[15041]_  = A167 & A169;
  assign \new_[15042]_  = ~A170 & \new_[15041]_ ;
  assign \new_[15046]_  = A200 & ~A199;
  assign \new_[15047]_  = A166 & \new_[15046]_ ;
  assign \new_[15048]_  = \new_[15047]_  & \new_[15042]_ ;
  assign \new_[15052]_  = A267 & ~A266;
  assign \new_[15053]_  = A265 & \new_[15052]_ ;
  assign \new_[15057]_  = ~A300 & A298;
  assign \new_[15058]_  = A268 & \new_[15057]_ ;
  assign \new_[15059]_  = \new_[15058]_  & \new_[15053]_ ;
  assign \new_[15063]_  = A167 & A169;
  assign \new_[15064]_  = ~A170 & \new_[15063]_ ;
  assign \new_[15068]_  = A200 & ~A199;
  assign \new_[15069]_  = A166 & \new_[15068]_ ;
  assign \new_[15070]_  = \new_[15069]_  & \new_[15064]_ ;
  assign \new_[15074]_  = A267 & ~A266;
  assign \new_[15075]_  = A265 & \new_[15074]_ ;
  assign \new_[15079]_  = A299 & A298;
  assign \new_[15080]_  = A268 & \new_[15079]_ ;
  assign \new_[15081]_  = \new_[15080]_  & \new_[15075]_ ;
  assign \new_[15085]_  = A167 & A169;
  assign \new_[15086]_  = ~A170 & \new_[15085]_ ;
  assign \new_[15090]_  = A200 & ~A199;
  assign \new_[15091]_  = A166 & \new_[15090]_ ;
  assign \new_[15092]_  = \new_[15091]_  & \new_[15086]_ ;
  assign \new_[15096]_  = A267 & ~A266;
  assign \new_[15097]_  = A265 & \new_[15096]_ ;
  assign \new_[15101]_  = ~A299 & ~A298;
  assign \new_[15102]_  = A268 & \new_[15101]_ ;
  assign \new_[15103]_  = \new_[15102]_  & \new_[15097]_ ;
  assign \new_[15107]_  = A167 & A169;
  assign \new_[15108]_  = ~A170 & \new_[15107]_ ;
  assign \new_[15112]_  = A200 & ~A199;
  assign \new_[15113]_  = A166 & \new_[15112]_ ;
  assign \new_[15114]_  = \new_[15113]_  & \new_[15108]_ ;
  assign \new_[15118]_  = A267 & ~A266;
  assign \new_[15119]_  = A265 & \new_[15118]_ ;
  assign \new_[15123]_  = ~A300 & A298;
  assign \new_[15124]_  = A269 & \new_[15123]_ ;
  assign \new_[15125]_  = \new_[15124]_  & \new_[15119]_ ;
  assign \new_[15129]_  = A167 & A169;
  assign \new_[15130]_  = ~A170 & \new_[15129]_ ;
  assign \new_[15134]_  = A200 & ~A199;
  assign \new_[15135]_  = A166 & \new_[15134]_ ;
  assign \new_[15136]_  = \new_[15135]_  & \new_[15130]_ ;
  assign \new_[15140]_  = A267 & ~A266;
  assign \new_[15141]_  = A265 & \new_[15140]_ ;
  assign \new_[15145]_  = A299 & A298;
  assign \new_[15146]_  = A269 & \new_[15145]_ ;
  assign \new_[15147]_  = \new_[15146]_  & \new_[15141]_ ;
  assign \new_[15151]_  = A167 & A169;
  assign \new_[15152]_  = ~A170 & \new_[15151]_ ;
  assign \new_[15156]_  = A200 & ~A199;
  assign \new_[15157]_  = A166 & \new_[15156]_ ;
  assign \new_[15158]_  = \new_[15157]_  & \new_[15152]_ ;
  assign \new_[15162]_  = A267 & ~A266;
  assign \new_[15163]_  = A265 & \new_[15162]_ ;
  assign \new_[15167]_  = ~A299 & ~A298;
  assign \new_[15168]_  = A269 & \new_[15167]_ ;
  assign \new_[15169]_  = \new_[15168]_  & \new_[15163]_ ;
  assign \new_[15173]_  = A167 & A169;
  assign \new_[15174]_  = ~A170 & \new_[15173]_ ;
  assign \new_[15178]_  = ~A202 & ~A200;
  assign \new_[15179]_  = A166 & \new_[15178]_ ;
  assign \new_[15180]_  = \new_[15179]_  & \new_[15174]_ ;
  assign \new_[15184]_  = ~A268 & ~A266;
  assign \new_[15185]_  = ~A203 & \new_[15184]_ ;
  assign \new_[15189]_  = A299 & ~A298;
  assign \new_[15190]_  = ~A269 & \new_[15189]_ ;
  assign \new_[15191]_  = \new_[15190]_  & \new_[15185]_ ;
  assign \new_[15195]_  = A167 & A169;
  assign \new_[15196]_  = ~A170 & \new_[15195]_ ;
  assign \new_[15200]_  = ~A201 & ~A200;
  assign \new_[15201]_  = A166 & \new_[15200]_ ;
  assign \new_[15202]_  = \new_[15201]_  & \new_[15196]_ ;
  assign \new_[15206]_  = A298 & A266;
  assign \new_[15207]_  = A265 & \new_[15206]_ ;
  assign \new_[15211]_  = A301 & A300;
  assign \new_[15212]_  = ~A299 & \new_[15211]_ ;
  assign \new_[15213]_  = \new_[15212]_  & \new_[15207]_ ;
  assign \new_[15217]_  = A167 & A169;
  assign \new_[15218]_  = ~A170 & \new_[15217]_ ;
  assign \new_[15222]_  = ~A201 & ~A200;
  assign \new_[15223]_  = A166 & \new_[15222]_ ;
  assign \new_[15224]_  = \new_[15223]_  & \new_[15218]_ ;
  assign \new_[15228]_  = A298 & A266;
  assign \new_[15229]_  = A265 & \new_[15228]_ ;
  assign \new_[15233]_  = A302 & A300;
  assign \new_[15234]_  = ~A299 & \new_[15233]_ ;
  assign \new_[15235]_  = \new_[15234]_  & \new_[15229]_ ;
  assign \new_[15239]_  = A167 & A169;
  assign \new_[15240]_  = ~A170 & \new_[15239]_ ;
  assign \new_[15244]_  = ~A201 & ~A200;
  assign \new_[15245]_  = A166 & \new_[15244]_ ;
  assign \new_[15246]_  = \new_[15245]_  & \new_[15240]_ ;
  assign \new_[15250]_  = A298 & ~A267;
  assign \new_[15251]_  = ~A266 & \new_[15250]_ ;
  assign \new_[15255]_  = A301 & A300;
  assign \new_[15256]_  = ~A299 & \new_[15255]_ ;
  assign \new_[15257]_  = \new_[15256]_  & \new_[15251]_ ;
  assign \new_[15261]_  = A167 & A169;
  assign \new_[15262]_  = ~A170 & \new_[15261]_ ;
  assign \new_[15266]_  = ~A201 & ~A200;
  assign \new_[15267]_  = A166 & \new_[15266]_ ;
  assign \new_[15268]_  = \new_[15267]_  & \new_[15262]_ ;
  assign \new_[15272]_  = A298 & ~A267;
  assign \new_[15273]_  = ~A266 & \new_[15272]_ ;
  assign \new_[15277]_  = A302 & A300;
  assign \new_[15278]_  = ~A299 & \new_[15277]_ ;
  assign \new_[15279]_  = \new_[15278]_  & \new_[15273]_ ;
  assign \new_[15283]_  = A167 & A169;
  assign \new_[15284]_  = ~A170 & \new_[15283]_ ;
  assign \new_[15288]_  = ~A201 & ~A200;
  assign \new_[15289]_  = A166 & \new_[15288]_ ;
  assign \new_[15290]_  = \new_[15289]_  & \new_[15284]_ ;
  assign \new_[15294]_  = A298 & ~A266;
  assign \new_[15295]_  = ~A265 & \new_[15294]_ ;
  assign \new_[15299]_  = A301 & A300;
  assign \new_[15300]_  = ~A299 & \new_[15299]_ ;
  assign \new_[15301]_  = \new_[15300]_  & \new_[15295]_ ;
  assign \new_[15305]_  = A167 & A169;
  assign \new_[15306]_  = ~A170 & \new_[15305]_ ;
  assign \new_[15310]_  = ~A201 & ~A200;
  assign \new_[15311]_  = A166 & \new_[15310]_ ;
  assign \new_[15312]_  = \new_[15311]_  & \new_[15306]_ ;
  assign \new_[15316]_  = A298 & ~A266;
  assign \new_[15317]_  = ~A265 & \new_[15316]_ ;
  assign \new_[15321]_  = A302 & A300;
  assign \new_[15322]_  = ~A299 & \new_[15321]_ ;
  assign \new_[15323]_  = \new_[15322]_  & \new_[15317]_ ;
  assign \new_[15327]_  = A167 & A169;
  assign \new_[15328]_  = ~A170 & \new_[15327]_ ;
  assign \new_[15332]_  = ~A200 & A199;
  assign \new_[15333]_  = A166 & \new_[15332]_ ;
  assign \new_[15334]_  = \new_[15333]_  & \new_[15328]_ ;
  assign \new_[15338]_  = ~A265 & A202;
  assign \new_[15339]_  = A201 & \new_[15338]_ ;
  assign \new_[15343]_  = ~A300 & A298;
  assign \new_[15344]_  = A266 & \new_[15343]_ ;
  assign \new_[15345]_  = \new_[15344]_  & \new_[15339]_ ;
  assign \new_[15349]_  = A167 & A169;
  assign \new_[15350]_  = ~A170 & \new_[15349]_ ;
  assign \new_[15354]_  = ~A200 & A199;
  assign \new_[15355]_  = A166 & \new_[15354]_ ;
  assign \new_[15356]_  = \new_[15355]_  & \new_[15350]_ ;
  assign \new_[15360]_  = ~A265 & A202;
  assign \new_[15361]_  = A201 & \new_[15360]_ ;
  assign \new_[15365]_  = A299 & A298;
  assign \new_[15366]_  = A266 & \new_[15365]_ ;
  assign \new_[15367]_  = \new_[15366]_  & \new_[15361]_ ;
  assign \new_[15371]_  = A167 & A169;
  assign \new_[15372]_  = ~A170 & \new_[15371]_ ;
  assign \new_[15376]_  = ~A200 & A199;
  assign \new_[15377]_  = A166 & \new_[15376]_ ;
  assign \new_[15378]_  = \new_[15377]_  & \new_[15372]_ ;
  assign \new_[15382]_  = ~A265 & A202;
  assign \new_[15383]_  = A201 & \new_[15382]_ ;
  assign \new_[15387]_  = ~A299 & ~A298;
  assign \new_[15388]_  = A266 & \new_[15387]_ ;
  assign \new_[15389]_  = \new_[15388]_  & \new_[15383]_ ;
  assign \new_[15393]_  = A167 & A169;
  assign \new_[15394]_  = ~A170 & \new_[15393]_ ;
  assign \new_[15398]_  = ~A200 & A199;
  assign \new_[15399]_  = A166 & \new_[15398]_ ;
  assign \new_[15400]_  = \new_[15399]_  & \new_[15394]_ ;
  assign \new_[15404]_  = ~A265 & A203;
  assign \new_[15405]_  = A201 & \new_[15404]_ ;
  assign \new_[15409]_  = ~A300 & A298;
  assign \new_[15410]_  = A266 & \new_[15409]_ ;
  assign \new_[15411]_  = \new_[15410]_  & \new_[15405]_ ;
  assign \new_[15415]_  = A167 & A169;
  assign \new_[15416]_  = ~A170 & \new_[15415]_ ;
  assign \new_[15420]_  = ~A200 & A199;
  assign \new_[15421]_  = A166 & \new_[15420]_ ;
  assign \new_[15422]_  = \new_[15421]_  & \new_[15416]_ ;
  assign \new_[15426]_  = ~A265 & A203;
  assign \new_[15427]_  = A201 & \new_[15426]_ ;
  assign \new_[15431]_  = A299 & A298;
  assign \new_[15432]_  = A266 & \new_[15431]_ ;
  assign \new_[15433]_  = \new_[15432]_  & \new_[15427]_ ;
  assign \new_[15437]_  = A167 & A169;
  assign \new_[15438]_  = ~A170 & \new_[15437]_ ;
  assign \new_[15442]_  = ~A200 & A199;
  assign \new_[15443]_  = A166 & \new_[15442]_ ;
  assign \new_[15444]_  = \new_[15443]_  & \new_[15438]_ ;
  assign \new_[15448]_  = ~A265 & A203;
  assign \new_[15449]_  = A201 & \new_[15448]_ ;
  assign \new_[15453]_  = ~A299 & ~A298;
  assign \new_[15454]_  = A266 & \new_[15453]_ ;
  assign \new_[15455]_  = \new_[15454]_  & \new_[15449]_ ;
  assign \new_[15459]_  = A167 & A169;
  assign \new_[15460]_  = ~A170 & \new_[15459]_ ;
  assign \new_[15464]_  = ~A200 & ~A199;
  assign \new_[15465]_  = A166 & \new_[15464]_ ;
  assign \new_[15466]_  = \new_[15465]_  & \new_[15460]_ ;
  assign \new_[15470]_  = A298 & A266;
  assign \new_[15471]_  = A265 & \new_[15470]_ ;
  assign \new_[15475]_  = A301 & A300;
  assign \new_[15476]_  = ~A299 & \new_[15475]_ ;
  assign \new_[15477]_  = \new_[15476]_  & \new_[15471]_ ;
  assign \new_[15481]_  = A167 & A169;
  assign \new_[15482]_  = ~A170 & \new_[15481]_ ;
  assign \new_[15486]_  = ~A200 & ~A199;
  assign \new_[15487]_  = A166 & \new_[15486]_ ;
  assign \new_[15488]_  = \new_[15487]_  & \new_[15482]_ ;
  assign \new_[15492]_  = A298 & A266;
  assign \new_[15493]_  = A265 & \new_[15492]_ ;
  assign \new_[15497]_  = A302 & A300;
  assign \new_[15498]_  = ~A299 & \new_[15497]_ ;
  assign \new_[15499]_  = \new_[15498]_  & \new_[15493]_ ;
  assign \new_[15503]_  = A167 & A169;
  assign \new_[15504]_  = ~A170 & \new_[15503]_ ;
  assign \new_[15508]_  = ~A200 & ~A199;
  assign \new_[15509]_  = A166 & \new_[15508]_ ;
  assign \new_[15510]_  = \new_[15509]_  & \new_[15504]_ ;
  assign \new_[15514]_  = A298 & ~A267;
  assign \new_[15515]_  = ~A266 & \new_[15514]_ ;
  assign \new_[15519]_  = A301 & A300;
  assign \new_[15520]_  = ~A299 & \new_[15519]_ ;
  assign \new_[15521]_  = \new_[15520]_  & \new_[15515]_ ;
  assign \new_[15525]_  = A167 & A169;
  assign \new_[15526]_  = ~A170 & \new_[15525]_ ;
  assign \new_[15530]_  = ~A200 & ~A199;
  assign \new_[15531]_  = A166 & \new_[15530]_ ;
  assign \new_[15532]_  = \new_[15531]_  & \new_[15526]_ ;
  assign \new_[15536]_  = A298 & ~A267;
  assign \new_[15537]_  = ~A266 & \new_[15536]_ ;
  assign \new_[15541]_  = A302 & A300;
  assign \new_[15542]_  = ~A299 & \new_[15541]_ ;
  assign \new_[15543]_  = \new_[15542]_  & \new_[15537]_ ;
  assign \new_[15547]_  = A167 & A169;
  assign \new_[15548]_  = ~A170 & \new_[15547]_ ;
  assign \new_[15552]_  = ~A200 & ~A199;
  assign \new_[15553]_  = A166 & \new_[15552]_ ;
  assign \new_[15554]_  = \new_[15553]_  & \new_[15548]_ ;
  assign \new_[15558]_  = A298 & ~A266;
  assign \new_[15559]_  = ~A265 & \new_[15558]_ ;
  assign \new_[15563]_  = A301 & A300;
  assign \new_[15564]_  = ~A299 & \new_[15563]_ ;
  assign \new_[15565]_  = \new_[15564]_  & \new_[15559]_ ;
  assign \new_[15569]_  = A167 & A169;
  assign \new_[15570]_  = ~A170 & \new_[15569]_ ;
  assign \new_[15574]_  = ~A200 & ~A199;
  assign \new_[15575]_  = A166 & \new_[15574]_ ;
  assign \new_[15576]_  = \new_[15575]_  & \new_[15570]_ ;
  assign \new_[15580]_  = A298 & ~A266;
  assign \new_[15581]_  = ~A265 & \new_[15580]_ ;
  assign \new_[15585]_  = A302 & A300;
  assign \new_[15586]_  = ~A299 & \new_[15585]_ ;
  assign \new_[15587]_  = \new_[15586]_  & \new_[15581]_ ;
  assign \new_[15591]_  = ~A167 & A169;
  assign \new_[15592]_  = ~A170 & \new_[15591]_ ;
  assign \new_[15596]_  = A200 & A199;
  assign \new_[15597]_  = ~A166 & \new_[15596]_ ;
  assign \new_[15598]_  = \new_[15597]_  & \new_[15592]_ ;
  assign \new_[15602]_  = A298 & A266;
  assign \new_[15603]_  = A265 & \new_[15602]_ ;
  assign \new_[15607]_  = A301 & A300;
  assign \new_[15608]_  = ~A299 & \new_[15607]_ ;
  assign \new_[15609]_  = \new_[15608]_  & \new_[15603]_ ;
  assign \new_[15613]_  = ~A167 & A169;
  assign \new_[15614]_  = ~A170 & \new_[15613]_ ;
  assign \new_[15618]_  = A200 & A199;
  assign \new_[15619]_  = ~A166 & \new_[15618]_ ;
  assign \new_[15620]_  = \new_[15619]_  & \new_[15614]_ ;
  assign \new_[15624]_  = A298 & A266;
  assign \new_[15625]_  = A265 & \new_[15624]_ ;
  assign \new_[15629]_  = A302 & A300;
  assign \new_[15630]_  = ~A299 & \new_[15629]_ ;
  assign \new_[15631]_  = \new_[15630]_  & \new_[15625]_ ;
  assign \new_[15635]_  = ~A167 & A169;
  assign \new_[15636]_  = ~A170 & \new_[15635]_ ;
  assign \new_[15640]_  = A200 & A199;
  assign \new_[15641]_  = ~A166 & \new_[15640]_ ;
  assign \new_[15642]_  = \new_[15641]_  & \new_[15636]_ ;
  assign \new_[15646]_  = A298 & ~A267;
  assign \new_[15647]_  = ~A266 & \new_[15646]_ ;
  assign \new_[15651]_  = A301 & A300;
  assign \new_[15652]_  = ~A299 & \new_[15651]_ ;
  assign \new_[15653]_  = \new_[15652]_  & \new_[15647]_ ;
  assign \new_[15657]_  = ~A167 & A169;
  assign \new_[15658]_  = ~A170 & \new_[15657]_ ;
  assign \new_[15662]_  = A200 & A199;
  assign \new_[15663]_  = ~A166 & \new_[15662]_ ;
  assign \new_[15664]_  = \new_[15663]_  & \new_[15658]_ ;
  assign \new_[15668]_  = A298 & ~A267;
  assign \new_[15669]_  = ~A266 & \new_[15668]_ ;
  assign \new_[15673]_  = A302 & A300;
  assign \new_[15674]_  = ~A299 & \new_[15673]_ ;
  assign \new_[15675]_  = \new_[15674]_  & \new_[15669]_ ;
  assign \new_[15679]_  = ~A167 & A169;
  assign \new_[15680]_  = ~A170 & \new_[15679]_ ;
  assign \new_[15684]_  = A200 & A199;
  assign \new_[15685]_  = ~A166 & \new_[15684]_ ;
  assign \new_[15686]_  = \new_[15685]_  & \new_[15680]_ ;
  assign \new_[15690]_  = A298 & ~A266;
  assign \new_[15691]_  = ~A265 & \new_[15690]_ ;
  assign \new_[15695]_  = A301 & A300;
  assign \new_[15696]_  = ~A299 & \new_[15695]_ ;
  assign \new_[15697]_  = \new_[15696]_  & \new_[15691]_ ;
  assign \new_[15701]_  = ~A167 & A169;
  assign \new_[15702]_  = ~A170 & \new_[15701]_ ;
  assign \new_[15706]_  = A200 & A199;
  assign \new_[15707]_  = ~A166 & \new_[15706]_ ;
  assign \new_[15708]_  = \new_[15707]_  & \new_[15702]_ ;
  assign \new_[15712]_  = A298 & ~A266;
  assign \new_[15713]_  = ~A265 & \new_[15712]_ ;
  assign \new_[15717]_  = A302 & A300;
  assign \new_[15718]_  = ~A299 & \new_[15717]_ ;
  assign \new_[15719]_  = \new_[15718]_  & \new_[15713]_ ;
  assign \new_[15723]_  = ~A167 & A169;
  assign \new_[15724]_  = ~A170 & \new_[15723]_ ;
  assign \new_[15728]_  = A200 & ~A199;
  assign \new_[15729]_  = ~A166 & \new_[15728]_ ;
  assign \new_[15730]_  = \new_[15729]_  & \new_[15724]_ ;
  assign \new_[15734]_  = A267 & ~A266;
  assign \new_[15735]_  = A265 & \new_[15734]_ ;
  assign \new_[15739]_  = ~A300 & A298;
  assign \new_[15740]_  = A268 & \new_[15739]_ ;
  assign \new_[15741]_  = \new_[15740]_  & \new_[15735]_ ;
  assign \new_[15745]_  = ~A167 & A169;
  assign \new_[15746]_  = ~A170 & \new_[15745]_ ;
  assign \new_[15750]_  = A200 & ~A199;
  assign \new_[15751]_  = ~A166 & \new_[15750]_ ;
  assign \new_[15752]_  = \new_[15751]_  & \new_[15746]_ ;
  assign \new_[15756]_  = A267 & ~A266;
  assign \new_[15757]_  = A265 & \new_[15756]_ ;
  assign \new_[15761]_  = A299 & A298;
  assign \new_[15762]_  = A268 & \new_[15761]_ ;
  assign \new_[15763]_  = \new_[15762]_  & \new_[15757]_ ;
  assign \new_[15767]_  = ~A167 & A169;
  assign \new_[15768]_  = ~A170 & \new_[15767]_ ;
  assign \new_[15772]_  = A200 & ~A199;
  assign \new_[15773]_  = ~A166 & \new_[15772]_ ;
  assign \new_[15774]_  = \new_[15773]_  & \new_[15768]_ ;
  assign \new_[15778]_  = A267 & ~A266;
  assign \new_[15779]_  = A265 & \new_[15778]_ ;
  assign \new_[15783]_  = ~A299 & ~A298;
  assign \new_[15784]_  = A268 & \new_[15783]_ ;
  assign \new_[15785]_  = \new_[15784]_  & \new_[15779]_ ;
  assign \new_[15789]_  = ~A167 & A169;
  assign \new_[15790]_  = ~A170 & \new_[15789]_ ;
  assign \new_[15794]_  = A200 & ~A199;
  assign \new_[15795]_  = ~A166 & \new_[15794]_ ;
  assign \new_[15796]_  = \new_[15795]_  & \new_[15790]_ ;
  assign \new_[15800]_  = A267 & ~A266;
  assign \new_[15801]_  = A265 & \new_[15800]_ ;
  assign \new_[15805]_  = ~A300 & A298;
  assign \new_[15806]_  = A269 & \new_[15805]_ ;
  assign \new_[15807]_  = \new_[15806]_  & \new_[15801]_ ;
  assign \new_[15811]_  = ~A167 & A169;
  assign \new_[15812]_  = ~A170 & \new_[15811]_ ;
  assign \new_[15816]_  = A200 & ~A199;
  assign \new_[15817]_  = ~A166 & \new_[15816]_ ;
  assign \new_[15818]_  = \new_[15817]_  & \new_[15812]_ ;
  assign \new_[15822]_  = A267 & ~A266;
  assign \new_[15823]_  = A265 & \new_[15822]_ ;
  assign \new_[15827]_  = A299 & A298;
  assign \new_[15828]_  = A269 & \new_[15827]_ ;
  assign \new_[15829]_  = \new_[15828]_  & \new_[15823]_ ;
  assign \new_[15833]_  = ~A167 & A169;
  assign \new_[15834]_  = ~A170 & \new_[15833]_ ;
  assign \new_[15838]_  = A200 & ~A199;
  assign \new_[15839]_  = ~A166 & \new_[15838]_ ;
  assign \new_[15840]_  = \new_[15839]_  & \new_[15834]_ ;
  assign \new_[15844]_  = A267 & ~A266;
  assign \new_[15845]_  = A265 & \new_[15844]_ ;
  assign \new_[15849]_  = ~A299 & ~A298;
  assign \new_[15850]_  = A269 & \new_[15849]_ ;
  assign \new_[15851]_  = \new_[15850]_  & \new_[15845]_ ;
  assign \new_[15855]_  = ~A167 & A169;
  assign \new_[15856]_  = ~A170 & \new_[15855]_ ;
  assign \new_[15860]_  = ~A202 & ~A200;
  assign \new_[15861]_  = ~A166 & \new_[15860]_ ;
  assign \new_[15862]_  = \new_[15861]_  & \new_[15856]_ ;
  assign \new_[15866]_  = ~A268 & ~A266;
  assign \new_[15867]_  = ~A203 & \new_[15866]_ ;
  assign \new_[15871]_  = A299 & ~A298;
  assign \new_[15872]_  = ~A269 & \new_[15871]_ ;
  assign \new_[15873]_  = \new_[15872]_  & \new_[15867]_ ;
  assign \new_[15877]_  = ~A167 & A169;
  assign \new_[15878]_  = ~A170 & \new_[15877]_ ;
  assign \new_[15882]_  = ~A201 & ~A200;
  assign \new_[15883]_  = ~A166 & \new_[15882]_ ;
  assign \new_[15884]_  = \new_[15883]_  & \new_[15878]_ ;
  assign \new_[15888]_  = A298 & A266;
  assign \new_[15889]_  = A265 & \new_[15888]_ ;
  assign \new_[15893]_  = A301 & A300;
  assign \new_[15894]_  = ~A299 & \new_[15893]_ ;
  assign \new_[15895]_  = \new_[15894]_  & \new_[15889]_ ;
  assign \new_[15899]_  = ~A167 & A169;
  assign \new_[15900]_  = ~A170 & \new_[15899]_ ;
  assign \new_[15904]_  = ~A201 & ~A200;
  assign \new_[15905]_  = ~A166 & \new_[15904]_ ;
  assign \new_[15906]_  = \new_[15905]_  & \new_[15900]_ ;
  assign \new_[15910]_  = A298 & A266;
  assign \new_[15911]_  = A265 & \new_[15910]_ ;
  assign \new_[15915]_  = A302 & A300;
  assign \new_[15916]_  = ~A299 & \new_[15915]_ ;
  assign \new_[15917]_  = \new_[15916]_  & \new_[15911]_ ;
  assign \new_[15921]_  = ~A167 & A169;
  assign \new_[15922]_  = ~A170 & \new_[15921]_ ;
  assign \new_[15926]_  = ~A201 & ~A200;
  assign \new_[15927]_  = ~A166 & \new_[15926]_ ;
  assign \new_[15928]_  = \new_[15927]_  & \new_[15922]_ ;
  assign \new_[15932]_  = A298 & ~A267;
  assign \new_[15933]_  = ~A266 & \new_[15932]_ ;
  assign \new_[15937]_  = A301 & A300;
  assign \new_[15938]_  = ~A299 & \new_[15937]_ ;
  assign \new_[15939]_  = \new_[15938]_  & \new_[15933]_ ;
  assign \new_[15943]_  = ~A167 & A169;
  assign \new_[15944]_  = ~A170 & \new_[15943]_ ;
  assign \new_[15948]_  = ~A201 & ~A200;
  assign \new_[15949]_  = ~A166 & \new_[15948]_ ;
  assign \new_[15950]_  = \new_[15949]_  & \new_[15944]_ ;
  assign \new_[15954]_  = A298 & ~A267;
  assign \new_[15955]_  = ~A266 & \new_[15954]_ ;
  assign \new_[15959]_  = A302 & A300;
  assign \new_[15960]_  = ~A299 & \new_[15959]_ ;
  assign \new_[15961]_  = \new_[15960]_  & \new_[15955]_ ;
  assign \new_[15965]_  = ~A167 & A169;
  assign \new_[15966]_  = ~A170 & \new_[15965]_ ;
  assign \new_[15970]_  = ~A201 & ~A200;
  assign \new_[15971]_  = ~A166 & \new_[15970]_ ;
  assign \new_[15972]_  = \new_[15971]_  & \new_[15966]_ ;
  assign \new_[15976]_  = A298 & ~A266;
  assign \new_[15977]_  = ~A265 & \new_[15976]_ ;
  assign \new_[15981]_  = A301 & A300;
  assign \new_[15982]_  = ~A299 & \new_[15981]_ ;
  assign \new_[15983]_  = \new_[15982]_  & \new_[15977]_ ;
  assign \new_[15987]_  = ~A167 & A169;
  assign \new_[15988]_  = ~A170 & \new_[15987]_ ;
  assign \new_[15992]_  = ~A201 & ~A200;
  assign \new_[15993]_  = ~A166 & \new_[15992]_ ;
  assign \new_[15994]_  = \new_[15993]_  & \new_[15988]_ ;
  assign \new_[15998]_  = A298 & ~A266;
  assign \new_[15999]_  = ~A265 & \new_[15998]_ ;
  assign \new_[16003]_  = A302 & A300;
  assign \new_[16004]_  = ~A299 & \new_[16003]_ ;
  assign \new_[16005]_  = \new_[16004]_  & \new_[15999]_ ;
  assign \new_[16009]_  = ~A167 & A169;
  assign \new_[16010]_  = ~A170 & \new_[16009]_ ;
  assign \new_[16014]_  = ~A200 & A199;
  assign \new_[16015]_  = ~A166 & \new_[16014]_ ;
  assign \new_[16016]_  = \new_[16015]_  & \new_[16010]_ ;
  assign \new_[16020]_  = ~A265 & A202;
  assign \new_[16021]_  = A201 & \new_[16020]_ ;
  assign \new_[16025]_  = ~A300 & A298;
  assign \new_[16026]_  = A266 & \new_[16025]_ ;
  assign \new_[16027]_  = \new_[16026]_  & \new_[16021]_ ;
  assign \new_[16031]_  = ~A167 & A169;
  assign \new_[16032]_  = ~A170 & \new_[16031]_ ;
  assign \new_[16036]_  = ~A200 & A199;
  assign \new_[16037]_  = ~A166 & \new_[16036]_ ;
  assign \new_[16038]_  = \new_[16037]_  & \new_[16032]_ ;
  assign \new_[16042]_  = ~A265 & A202;
  assign \new_[16043]_  = A201 & \new_[16042]_ ;
  assign \new_[16047]_  = A299 & A298;
  assign \new_[16048]_  = A266 & \new_[16047]_ ;
  assign \new_[16049]_  = \new_[16048]_  & \new_[16043]_ ;
  assign \new_[16053]_  = ~A167 & A169;
  assign \new_[16054]_  = ~A170 & \new_[16053]_ ;
  assign \new_[16058]_  = ~A200 & A199;
  assign \new_[16059]_  = ~A166 & \new_[16058]_ ;
  assign \new_[16060]_  = \new_[16059]_  & \new_[16054]_ ;
  assign \new_[16064]_  = ~A265 & A202;
  assign \new_[16065]_  = A201 & \new_[16064]_ ;
  assign \new_[16069]_  = ~A299 & ~A298;
  assign \new_[16070]_  = A266 & \new_[16069]_ ;
  assign \new_[16071]_  = \new_[16070]_  & \new_[16065]_ ;
  assign \new_[16075]_  = ~A167 & A169;
  assign \new_[16076]_  = ~A170 & \new_[16075]_ ;
  assign \new_[16080]_  = ~A200 & A199;
  assign \new_[16081]_  = ~A166 & \new_[16080]_ ;
  assign \new_[16082]_  = \new_[16081]_  & \new_[16076]_ ;
  assign \new_[16086]_  = ~A265 & A203;
  assign \new_[16087]_  = A201 & \new_[16086]_ ;
  assign \new_[16091]_  = ~A300 & A298;
  assign \new_[16092]_  = A266 & \new_[16091]_ ;
  assign \new_[16093]_  = \new_[16092]_  & \new_[16087]_ ;
  assign \new_[16097]_  = ~A167 & A169;
  assign \new_[16098]_  = ~A170 & \new_[16097]_ ;
  assign \new_[16102]_  = ~A200 & A199;
  assign \new_[16103]_  = ~A166 & \new_[16102]_ ;
  assign \new_[16104]_  = \new_[16103]_  & \new_[16098]_ ;
  assign \new_[16108]_  = ~A265 & A203;
  assign \new_[16109]_  = A201 & \new_[16108]_ ;
  assign \new_[16113]_  = A299 & A298;
  assign \new_[16114]_  = A266 & \new_[16113]_ ;
  assign \new_[16115]_  = \new_[16114]_  & \new_[16109]_ ;
  assign \new_[16119]_  = ~A167 & A169;
  assign \new_[16120]_  = ~A170 & \new_[16119]_ ;
  assign \new_[16124]_  = ~A200 & A199;
  assign \new_[16125]_  = ~A166 & \new_[16124]_ ;
  assign \new_[16126]_  = \new_[16125]_  & \new_[16120]_ ;
  assign \new_[16130]_  = ~A265 & A203;
  assign \new_[16131]_  = A201 & \new_[16130]_ ;
  assign \new_[16135]_  = ~A299 & ~A298;
  assign \new_[16136]_  = A266 & \new_[16135]_ ;
  assign \new_[16137]_  = \new_[16136]_  & \new_[16131]_ ;
  assign \new_[16141]_  = ~A167 & A169;
  assign \new_[16142]_  = ~A170 & \new_[16141]_ ;
  assign \new_[16146]_  = ~A200 & ~A199;
  assign \new_[16147]_  = ~A166 & \new_[16146]_ ;
  assign \new_[16148]_  = \new_[16147]_  & \new_[16142]_ ;
  assign \new_[16152]_  = A298 & A266;
  assign \new_[16153]_  = A265 & \new_[16152]_ ;
  assign \new_[16157]_  = A301 & A300;
  assign \new_[16158]_  = ~A299 & \new_[16157]_ ;
  assign \new_[16159]_  = \new_[16158]_  & \new_[16153]_ ;
  assign \new_[16163]_  = ~A167 & A169;
  assign \new_[16164]_  = ~A170 & \new_[16163]_ ;
  assign \new_[16168]_  = ~A200 & ~A199;
  assign \new_[16169]_  = ~A166 & \new_[16168]_ ;
  assign \new_[16170]_  = \new_[16169]_  & \new_[16164]_ ;
  assign \new_[16174]_  = A298 & A266;
  assign \new_[16175]_  = A265 & \new_[16174]_ ;
  assign \new_[16179]_  = A302 & A300;
  assign \new_[16180]_  = ~A299 & \new_[16179]_ ;
  assign \new_[16181]_  = \new_[16180]_  & \new_[16175]_ ;
  assign \new_[16185]_  = ~A167 & A169;
  assign \new_[16186]_  = ~A170 & \new_[16185]_ ;
  assign \new_[16190]_  = ~A200 & ~A199;
  assign \new_[16191]_  = ~A166 & \new_[16190]_ ;
  assign \new_[16192]_  = \new_[16191]_  & \new_[16186]_ ;
  assign \new_[16196]_  = A298 & ~A267;
  assign \new_[16197]_  = ~A266 & \new_[16196]_ ;
  assign \new_[16201]_  = A301 & A300;
  assign \new_[16202]_  = ~A299 & \new_[16201]_ ;
  assign \new_[16203]_  = \new_[16202]_  & \new_[16197]_ ;
  assign \new_[16207]_  = ~A167 & A169;
  assign \new_[16208]_  = ~A170 & \new_[16207]_ ;
  assign \new_[16212]_  = ~A200 & ~A199;
  assign \new_[16213]_  = ~A166 & \new_[16212]_ ;
  assign \new_[16214]_  = \new_[16213]_  & \new_[16208]_ ;
  assign \new_[16218]_  = A298 & ~A267;
  assign \new_[16219]_  = ~A266 & \new_[16218]_ ;
  assign \new_[16223]_  = A302 & A300;
  assign \new_[16224]_  = ~A299 & \new_[16223]_ ;
  assign \new_[16225]_  = \new_[16224]_  & \new_[16219]_ ;
  assign \new_[16229]_  = ~A167 & A169;
  assign \new_[16230]_  = ~A170 & \new_[16229]_ ;
  assign \new_[16234]_  = ~A200 & ~A199;
  assign \new_[16235]_  = ~A166 & \new_[16234]_ ;
  assign \new_[16236]_  = \new_[16235]_  & \new_[16230]_ ;
  assign \new_[16240]_  = A298 & ~A266;
  assign \new_[16241]_  = ~A265 & \new_[16240]_ ;
  assign \new_[16245]_  = A301 & A300;
  assign \new_[16246]_  = ~A299 & \new_[16245]_ ;
  assign \new_[16247]_  = \new_[16246]_  & \new_[16241]_ ;
  assign \new_[16251]_  = ~A167 & A169;
  assign \new_[16252]_  = ~A170 & \new_[16251]_ ;
  assign \new_[16256]_  = ~A200 & ~A199;
  assign \new_[16257]_  = ~A166 & \new_[16256]_ ;
  assign \new_[16258]_  = \new_[16257]_  & \new_[16252]_ ;
  assign \new_[16262]_  = A298 & ~A266;
  assign \new_[16263]_  = ~A265 & \new_[16262]_ ;
  assign \new_[16267]_  = A302 & A300;
  assign \new_[16268]_  = ~A299 & \new_[16267]_ ;
  assign \new_[16269]_  = \new_[16268]_  & \new_[16263]_ ;
  assign \new_[16273]_  = ~A166 & ~A167;
  assign \new_[16274]_  = ~A169 & \new_[16273]_ ;
  assign \new_[16278]_  = A265 & A200;
  assign \new_[16279]_  = A199 & \new_[16278]_ ;
  assign \new_[16280]_  = \new_[16279]_  & \new_[16274]_ ;
  assign \new_[16284]_  = A268 & A267;
  assign \new_[16285]_  = ~A266 & \new_[16284]_ ;
  assign \new_[16289]_  = ~A302 & ~A301;
  assign \new_[16290]_  = A298 & \new_[16289]_ ;
  assign \new_[16291]_  = \new_[16290]_  & \new_[16285]_ ;
  assign \new_[16295]_  = ~A166 & ~A167;
  assign \new_[16296]_  = ~A169 & \new_[16295]_ ;
  assign \new_[16300]_  = A265 & A200;
  assign \new_[16301]_  = A199 & \new_[16300]_ ;
  assign \new_[16302]_  = \new_[16301]_  & \new_[16296]_ ;
  assign \new_[16306]_  = A269 & A267;
  assign \new_[16307]_  = ~A266 & \new_[16306]_ ;
  assign \new_[16311]_  = ~A302 & ~A301;
  assign \new_[16312]_  = A298 & \new_[16311]_ ;
  assign \new_[16313]_  = \new_[16312]_  & \new_[16307]_ ;
  assign \new_[16317]_  = ~A166 & ~A167;
  assign \new_[16318]_  = ~A169 & \new_[16317]_ ;
  assign \new_[16322]_  = ~A266 & A200;
  assign \new_[16323]_  = ~A199 & \new_[16322]_ ;
  assign \new_[16324]_  = \new_[16323]_  & \new_[16318]_ ;
  assign \new_[16328]_  = A298 & ~A269;
  assign \new_[16329]_  = ~A268 & \new_[16328]_ ;
  assign \new_[16333]_  = A301 & A300;
  assign \new_[16334]_  = ~A299 & \new_[16333]_ ;
  assign \new_[16335]_  = \new_[16334]_  & \new_[16329]_ ;
  assign \new_[16339]_  = ~A166 & ~A167;
  assign \new_[16340]_  = ~A169 & \new_[16339]_ ;
  assign \new_[16344]_  = ~A266 & A200;
  assign \new_[16345]_  = ~A199 & \new_[16344]_ ;
  assign \new_[16346]_  = \new_[16345]_  & \new_[16340]_ ;
  assign \new_[16350]_  = A298 & ~A269;
  assign \new_[16351]_  = ~A268 & \new_[16350]_ ;
  assign \new_[16355]_  = A302 & A300;
  assign \new_[16356]_  = ~A299 & \new_[16355]_ ;
  assign \new_[16357]_  = \new_[16356]_  & \new_[16351]_ ;
  assign \new_[16361]_  = ~A166 & ~A167;
  assign \new_[16362]_  = ~A169 & \new_[16361]_ ;
  assign \new_[16366]_  = ~A203 & ~A202;
  assign \new_[16367]_  = ~A200 & \new_[16366]_ ;
  assign \new_[16368]_  = \new_[16367]_  & \new_[16362]_ ;
  assign \new_[16372]_  = A267 & ~A266;
  assign \new_[16373]_  = A265 & \new_[16372]_ ;
  assign \new_[16377]_  = ~A300 & A298;
  assign \new_[16378]_  = A268 & \new_[16377]_ ;
  assign \new_[16379]_  = \new_[16378]_  & \new_[16373]_ ;
  assign \new_[16383]_  = ~A166 & ~A167;
  assign \new_[16384]_  = ~A169 & \new_[16383]_ ;
  assign \new_[16388]_  = ~A203 & ~A202;
  assign \new_[16389]_  = ~A200 & \new_[16388]_ ;
  assign \new_[16390]_  = \new_[16389]_  & \new_[16384]_ ;
  assign \new_[16394]_  = A267 & ~A266;
  assign \new_[16395]_  = A265 & \new_[16394]_ ;
  assign \new_[16399]_  = A299 & A298;
  assign \new_[16400]_  = A268 & \new_[16399]_ ;
  assign \new_[16401]_  = \new_[16400]_  & \new_[16395]_ ;
  assign \new_[16405]_  = ~A166 & ~A167;
  assign \new_[16406]_  = ~A169 & \new_[16405]_ ;
  assign \new_[16410]_  = ~A203 & ~A202;
  assign \new_[16411]_  = ~A200 & \new_[16410]_ ;
  assign \new_[16412]_  = \new_[16411]_  & \new_[16406]_ ;
  assign \new_[16416]_  = A267 & ~A266;
  assign \new_[16417]_  = A265 & \new_[16416]_ ;
  assign \new_[16421]_  = ~A299 & ~A298;
  assign \new_[16422]_  = A268 & \new_[16421]_ ;
  assign \new_[16423]_  = \new_[16422]_  & \new_[16417]_ ;
  assign \new_[16427]_  = ~A166 & ~A167;
  assign \new_[16428]_  = ~A169 & \new_[16427]_ ;
  assign \new_[16432]_  = ~A203 & ~A202;
  assign \new_[16433]_  = ~A200 & \new_[16432]_ ;
  assign \new_[16434]_  = \new_[16433]_  & \new_[16428]_ ;
  assign \new_[16438]_  = A267 & ~A266;
  assign \new_[16439]_  = A265 & \new_[16438]_ ;
  assign \new_[16443]_  = ~A300 & A298;
  assign \new_[16444]_  = A269 & \new_[16443]_ ;
  assign \new_[16445]_  = \new_[16444]_  & \new_[16439]_ ;
  assign \new_[16449]_  = ~A166 & ~A167;
  assign \new_[16450]_  = ~A169 & \new_[16449]_ ;
  assign \new_[16454]_  = ~A203 & ~A202;
  assign \new_[16455]_  = ~A200 & \new_[16454]_ ;
  assign \new_[16456]_  = \new_[16455]_  & \new_[16450]_ ;
  assign \new_[16460]_  = A267 & ~A266;
  assign \new_[16461]_  = A265 & \new_[16460]_ ;
  assign \new_[16465]_  = A299 & A298;
  assign \new_[16466]_  = A269 & \new_[16465]_ ;
  assign \new_[16467]_  = \new_[16466]_  & \new_[16461]_ ;
  assign \new_[16471]_  = ~A166 & ~A167;
  assign \new_[16472]_  = ~A169 & \new_[16471]_ ;
  assign \new_[16476]_  = ~A203 & ~A202;
  assign \new_[16477]_  = ~A200 & \new_[16476]_ ;
  assign \new_[16478]_  = \new_[16477]_  & \new_[16472]_ ;
  assign \new_[16482]_  = A267 & ~A266;
  assign \new_[16483]_  = A265 & \new_[16482]_ ;
  assign \new_[16487]_  = ~A299 & ~A298;
  assign \new_[16488]_  = A269 & \new_[16487]_ ;
  assign \new_[16489]_  = \new_[16488]_  & \new_[16483]_ ;
  assign \new_[16493]_  = ~A166 & ~A167;
  assign \new_[16494]_  = ~A169 & \new_[16493]_ ;
  assign \new_[16498]_  = A265 & ~A201;
  assign \new_[16499]_  = ~A200 & \new_[16498]_ ;
  assign \new_[16500]_  = \new_[16499]_  & \new_[16494]_ ;
  assign \new_[16504]_  = A268 & A267;
  assign \new_[16505]_  = ~A266 & \new_[16504]_ ;
  assign \new_[16509]_  = ~A302 & ~A301;
  assign \new_[16510]_  = A298 & \new_[16509]_ ;
  assign \new_[16511]_  = \new_[16510]_  & \new_[16505]_ ;
  assign \new_[16515]_  = ~A166 & ~A167;
  assign \new_[16516]_  = ~A169 & \new_[16515]_ ;
  assign \new_[16520]_  = A265 & ~A201;
  assign \new_[16521]_  = ~A200 & \new_[16520]_ ;
  assign \new_[16522]_  = \new_[16521]_  & \new_[16516]_ ;
  assign \new_[16526]_  = A269 & A267;
  assign \new_[16527]_  = ~A266 & \new_[16526]_ ;
  assign \new_[16531]_  = ~A302 & ~A301;
  assign \new_[16532]_  = A298 & \new_[16531]_ ;
  assign \new_[16533]_  = \new_[16532]_  & \new_[16527]_ ;
  assign \new_[16537]_  = ~A166 & ~A167;
  assign \new_[16538]_  = ~A169 & \new_[16537]_ ;
  assign \new_[16542]_  = A201 & ~A200;
  assign \new_[16543]_  = A199 & \new_[16542]_ ;
  assign \new_[16544]_  = \new_[16543]_  & \new_[16538]_ ;
  assign \new_[16548]_  = ~A268 & ~A266;
  assign \new_[16549]_  = A202 & \new_[16548]_ ;
  assign \new_[16553]_  = A299 & ~A298;
  assign \new_[16554]_  = ~A269 & \new_[16553]_ ;
  assign \new_[16555]_  = \new_[16554]_  & \new_[16549]_ ;
  assign \new_[16559]_  = ~A166 & ~A167;
  assign \new_[16560]_  = ~A169 & \new_[16559]_ ;
  assign \new_[16564]_  = A201 & ~A200;
  assign \new_[16565]_  = A199 & \new_[16564]_ ;
  assign \new_[16566]_  = \new_[16565]_  & \new_[16560]_ ;
  assign \new_[16570]_  = ~A268 & ~A266;
  assign \new_[16571]_  = A203 & \new_[16570]_ ;
  assign \new_[16575]_  = A299 & ~A298;
  assign \new_[16576]_  = ~A269 & \new_[16575]_ ;
  assign \new_[16577]_  = \new_[16576]_  & \new_[16571]_ ;
  assign \new_[16581]_  = ~A166 & ~A167;
  assign \new_[16582]_  = ~A169 & \new_[16581]_ ;
  assign \new_[16586]_  = A265 & ~A200;
  assign \new_[16587]_  = ~A199 & \new_[16586]_ ;
  assign \new_[16588]_  = \new_[16587]_  & \new_[16582]_ ;
  assign \new_[16592]_  = A268 & A267;
  assign \new_[16593]_  = ~A266 & \new_[16592]_ ;
  assign \new_[16597]_  = ~A302 & ~A301;
  assign \new_[16598]_  = A298 & \new_[16597]_ ;
  assign \new_[16599]_  = \new_[16598]_  & \new_[16593]_ ;
  assign \new_[16603]_  = ~A166 & ~A167;
  assign \new_[16604]_  = ~A169 & \new_[16603]_ ;
  assign \new_[16608]_  = A265 & ~A200;
  assign \new_[16609]_  = ~A199 & \new_[16608]_ ;
  assign \new_[16610]_  = \new_[16609]_  & \new_[16604]_ ;
  assign \new_[16614]_  = A269 & A267;
  assign \new_[16615]_  = ~A266 & \new_[16614]_ ;
  assign \new_[16619]_  = ~A302 & ~A301;
  assign \new_[16620]_  = A298 & \new_[16619]_ ;
  assign \new_[16621]_  = \new_[16620]_  & \new_[16615]_ ;
  assign \new_[16625]_  = A167 & ~A168;
  assign \new_[16626]_  = ~A169 & \new_[16625]_ ;
  assign \new_[16630]_  = A200 & A199;
  assign \new_[16631]_  = A166 & \new_[16630]_ ;
  assign \new_[16632]_  = \new_[16631]_  & \new_[16626]_ ;
  assign \new_[16636]_  = A267 & ~A266;
  assign \new_[16637]_  = A265 & \new_[16636]_ ;
  assign \new_[16641]_  = ~A300 & A298;
  assign \new_[16642]_  = A268 & \new_[16641]_ ;
  assign \new_[16643]_  = \new_[16642]_  & \new_[16637]_ ;
  assign \new_[16647]_  = A167 & ~A168;
  assign \new_[16648]_  = ~A169 & \new_[16647]_ ;
  assign \new_[16652]_  = A200 & A199;
  assign \new_[16653]_  = A166 & \new_[16652]_ ;
  assign \new_[16654]_  = \new_[16653]_  & \new_[16648]_ ;
  assign \new_[16658]_  = A267 & ~A266;
  assign \new_[16659]_  = A265 & \new_[16658]_ ;
  assign \new_[16663]_  = A299 & A298;
  assign \new_[16664]_  = A268 & \new_[16663]_ ;
  assign \new_[16665]_  = \new_[16664]_  & \new_[16659]_ ;
  assign \new_[16669]_  = A167 & ~A168;
  assign \new_[16670]_  = ~A169 & \new_[16669]_ ;
  assign \new_[16674]_  = A200 & A199;
  assign \new_[16675]_  = A166 & \new_[16674]_ ;
  assign \new_[16676]_  = \new_[16675]_  & \new_[16670]_ ;
  assign \new_[16680]_  = A267 & ~A266;
  assign \new_[16681]_  = A265 & \new_[16680]_ ;
  assign \new_[16685]_  = ~A299 & ~A298;
  assign \new_[16686]_  = A268 & \new_[16685]_ ;
  assign \new_[16687]_  = \new_[16686]_  & \new_[16681]_ ;
  assign \new_[16691]_  = A167 & ~A168;
  assign \new_[16692]_  = ~A169 & \new_[16691]_ ;
  assign \new_[16696]_  = A200 & A199;
  assign \new_[16697]_  = A166 & \new_[16696]_ ;
  assign \new_[16698]_  = \new_[16697]_  & \new_[16692]_ ;
  assign \new_[16702]_  = A267 & ~A266;
  assign \new_[16703]_  = A265 & \new_[16702]_ ;
  assign \new_[16707]_  = ~A300 & A298;
  assign \new_[16708]_  = A269 & \new_[16707]_ ;
  assign \new_[16709]_  = \new_[16708]_  & \new_[16703]_ ;
  assign \new_[16713]_  = A167 & ~A168;
  assign \new_[16714]_  = ~A169 & \new_[16713]_ ;
  assign \new_[16718]_  = A200 & A199;
  assign \new_[16719]_  = A166 & \new_[16718]_ ;
  assign \new_[16720]_  = \new_[16719]_  & \new_[16714]_ ;
  assign \new_[16724]_  = A267 & ~A266;
  assign \new_[16725]_  = A265 & \new_[16724]_ ;
  assign \new_[16729]_  = A299 & A298;
  assign \new_[16730]_  = A269 & \new_[16729]_ ;
  assign \new_[16731]_  = \new_[16730]_  & \new_[16725]_ ;
  assign \new_[16735]_  = A167 & ~A168;
  assign \new_[16736]_  = ~A169 & \new_[16735]_ ;
  assign \new_[16740]_  = A200 & A199;
  assign \new_[16741]_  = A166 & \new_[16740]_ ;
  assign \new_[16742]_  = \new_[16741]_  & \new_[16736]_ ;
  assign \new_[16746]_  = A267 & ~A266;
  assign \new_[16747]_  = A265 & \new_[16746]_ ;
  assign \new_[16751]_  = ~A299 & ~A298;
  assign \new_[16752]_  = A269 & \new_[16751]_ ;
  assign \new_[16753]_  = \new_[16752]_  & \new_[16747]_ ;
  assign \new_[16757]_  = A167 & ~A168;
  assign \new_[16758]_  = ~A169 & \new_[16757]_ ;
  assign \new_[16762]_  = A200 & ~A199;
  assign \new_[16763]_  = A166 & \new_[16762]_ ;
  assign \new_[16764]_  = \new_[16763]_  & \new_[16758]_ ;
  assign \new_[16768]_  = A298 & A266;
  assign \new_[16769]_  = A265 & \new_[16768]_ ;
  assign \new_[16773]_  = A301 & A300;
  assign \new_[16774]_  = ~A299 & \new_[16773]_ ;
  assign \new_[16775]_  = \new_[16774]_  & \new_[16769]_ ;
  assign \new_[16779]_  = A167 & ~A168;
  assign \new_[16780]_  = ~A169 & \new_[16779]_ ;
  assign \new_[16784]_  = A200 & ~A199;
  assign \new_[16785]_  = A166 & \new_[16784]_ ;
  assign \new_[16786]_  = \new_[16785]_  & \new_[16780]_ ;
  assign \new_[16790]_  = A298 & A266;
  assign \new_[16791]_  = A265 & \new_[16790]_ ;
  assign \new_[16795]_  = A302 & A300;
  assign \new_[16796]_  = ~A299 & \new_[16795]_ ;
  assign \new_[16797]_  = \new_[16796]_  & \new_[16791]_ ;
  assign \new_[16801]_  = A167 & ~A168;
  assign \new_[16802]_  = ~A169 & \new_[16801]_ ;
  assign \new_[16806]_  = A200 & ~A199;
  assign \new_[16807]_  = A166 & \new_[16806]_ ;
  assign \new_[16808]_  = \new_[16807]_  & \new_[16802]_ ;
  assign \new_[16812]_  = A298 & ~A267;
  assign \new_[16813]_  = ~A266 & \new_[16812]_ ;
  assign \new_[16817]_  = A301 & A300;
  assign \new_[16818]_  = ~A299 & \new_[16817]_ ;
  assign \new_[16819]_  = \new_[16818]_  & \new_[16813]_ ;
  assign \new_[16823]_  = A167 & ~A168;
  assign \new_[16824]_  = ~A169 & \new_[16823]_ ;
  assign \new_[16828]_  = A200 & ~A199;
  assign \new_[16829]_  = A166 & \new_[16828]_ ;
  assign \new_[16830]_  = \new_[16829]_  & \new_[16824]_ ;
  assign \new_[16834]_  = A298 & ~A267;
  assign \new_[16835]_  = ~A266 & \new_[16834]_ ;
  assign \new_[16839]_  = A302 & A300;
  assign \new_[16840]_  = ~A299 & \new_[16839]_ ;
  assign \new_[16841]_  = \new_[16840]_  & \new_[16835]_ ;
  assign \new_[16845]_  = A167 & ~A168;
  assign \new_[16846]_  = ~A169 & \new_[16845]_ ;
  assign \new_[16850]_  = A200 & ~A199;
  assign \new_[16851]_  = A166 & \new_[16850]_ ;
  assign \new_[16852]_  = \new_[16851]_  & \new_[16846]_ ;
  assign \new_[16856]_  = A298 & ~A266;
  assign \new_[16857]_  = ~A265 & \new_[16856]_ ;
  assign \new_[16861]_  = A301 & A300;
  assign \new_[16862]_  = ~A299 & \new_[16861]_ ;
  assign \new_[16863]_  = \new_[16862]_  & \new_[16857]_ ;
  assign \new_[16867]_  = A167 & ~A168;
  assign \new_[16868]_  = ~A169 & \new_[16867]_ ;
  assign \new_[16872]_  = A200 & ~A199;
  assign \new_[16873]_  = A166 & \new_[16872]_ ;
  assign \new_[16874]_  = \new_[16873]_  & \new_[16868]_ ;
  assign \new_[16878]_  = A298 & ~A266;
  assign \new_[16879]_  = ~A265 & \new_[16878]_ ;
  assign \new_[16883]_  = A302 & A300;
  assign \new_[16884]_  = ~A299 & \new_[16883]_ ;
  assign \new_[16885]_  = \new_[16884]_  & \new_[16879]_ ;
  assign \new_[16889]_  = A167 & ~A168;
  assign \new_[16890]_  = ~A169 & \new_[16889]_ ;
  assign \new_[16894]_  = ~A202 & ~A200;
  assign \new_[16895]_  = A166 & \new_[16894]_ ;
  assign \new_[16896]_  = \new_[16895]_  & \new_[16890]_ ;
  assign \new_[16900]_  = A266 & ~A265;
  assign \new_[16901]_  = ~A203 & \new_[16900]_ ;
  assign \new_[16905]_  = ~A302 & ~A301;
  assign \new_[16906]_  = A298 & \new_[16905]_ ;
  assign \new_[16907]_  = \new_[16906]_  & \new_[16901]_ ;
  assign \new_[16911]_  = A167 & ~A168;
  assign \new_[16912]_  = ~A169 & \new_[16911]_ ;
  assign \new_[16916]_  = ~A201 & ~A200;
  assign \new_[16917]_  = A166 & \new_[16916]_ ;
  assign \new_[16918]_  = \new_[16917]_  & \new_[16912]_ ;
  assign \new_[16922]_  = A267 & ~A266;
  assign \new_[16923]_  = A265 & \new_[16922]_ ;
  assign \new_[16927]_  = ~A300 & A298;
  assign \new_[16928]_  = A268 & \new_[16927]_ ;
  assign \new_[16929]_  = \new_[16928]_  & \new_[16923]_ ;
  assign \new_[16933]_  = A167 & ~A168;
  assign \new_[16934]_  = ~A169 & \new_[16933]_ ;
  assign \new_[16938]_  = ~A201 & ~A200;
  assign \new_[16939]_  = A166 & \new_[16938]_ ;
  assign \new_[16940]_  = \new_[16939]_  & \new_[16934]_ ;
  assign \new_[16944]_  = A267 & ~A266;
  assign \new_[16945]_  = A265 & \new_[16944]_ ;
  assign \new_[16949]_  = A299 & A298;
  assign \new_[16950]_  = A268 & \new_[16949]_ ;
  assign \new_[16951]_  = \new_[16950]_  & \new_[16945]_ ;
  assign \new_[16955]_  = A167 & ~A168;
  assign \new_[16956]_  = ~A169 & \new_[16955]_ ;
  assign \new_[16960]_  = ~A201 & ~A200;
  assign \new_[16961]_  = A166 & \new_[16960]_ ;
  assign \new_[16962]_  = \new_[16961]_  & \new_[16956]_ ;
  assign \new_[16966]_  = A267 & ~A266;
  assign \new_[16967]_  = A265 & \new_[16966]_ ;
  assign \new_[16971]_  = ~A299 & ~A298;
  assign \new_[16972]_  = A268 & \new_[16971]_ ;
  assign \new_[16973]_  = \new_[16972]_  & \new_[16967]_ ;
  assign \new_[16977]_  = A167 & ~A168;
  assign \new_[16978]_  = ~A169 & \new_[16977]_ ;
  assign \new_[16982]_  = ~A201 & ~A200;
  assign \new_[16983]_  = A166 & \new_[16982]_ ;
  assign \new_[16984]_  = \new_[16983]_  & \new_[16978]_ ;
  assign \new_[16988]_  = A267 & ~A266;
  assign \new_[16989]_  = A265 & \new_[16988]_ ;
  assign \new_[16993]_  = ~A300 & A298;
  assign \new_[16994]_  = A269 & \new_[16993]_ ;
  assign \new_[16995]_  = \new_[16994]_  & \new_[16989]_ ;
  assign \new_[16999]_  = A167 & ~A168;
  assign \new_[17000]_  = ~A169 & \new_[16999]_ ;
  assign \new_[17004]_  = ~A201 & ~A200;
  assign \new_[17005]_  = A166 & \new_[17004]_ ;
  assign \new_[17006]_  = \new_[17005]_  & \new_[17000]_ ;
  assign \new_[17010]_  = A267 & ~A266;
  assign \new_[17011]_  = A265 & \new_[17010]_ ;
  assign \new_[17015]_  = A299 & A298;
  assign \new_[17016]_  = A269 & \new_[17015]_ ;
  assign \new_[17017]_  = \new_[17016]_  & \new_[17011]_ ;
  assign \new_[17021]_  = A167 & ~A168;
  assign \new_[17022]_  = ~A169 & \new_[17021]_ ;
  assign \new_[17026]_  = ~A201 & ~A200;
  assign \new_[17027]_  = A166 & \new_[17026]_ ;
  assign \new_[17028]_  = \new_[17027]_  & \new_[17022]_ ;
  assign \new_[17032]_  = A267 & ~A266;
  assign \new_[17033]_  = A265 & \new_[17032]_ ;
  assign \new_[17037]_  = ~A299 & ~A298;
  assign \new_[17038]_  = A269 & \new_[17037]_ ;
  assign \new_[17039]_  = \new_[17038]_  & \new_[17033]_ ;
  assign \new_[17043]_  = A167 & ~A168;
  assign \new_[17044]_  = ~A169 & \new_[17043]_ ;
  assign \new_[17048]_  = ~A200 & A199;
  assign \new_[17049]_  = A166 & \new_[17048]_ ;
  assign \new_[17050]_  = \new_[17049]_  & \new_[17044]_ ;
  assign \new_[17054]_  = A265 & A202;
  assign \new_[17055]_  = A201 & \new_[17054]_ ;
  assign \new_[17059]_  = A299 & ~A298;
  assign \new_[17060]_  = A266 & \new_[17059]_ ;
  assign \new_[17061]_  = \new_[17060]_  & \new_[17055]_ ;
  assign \new_[17065]_  = A167 & ~A168;
  assign \new_[17066]_  = ~A169 & \new_[17065]_ ;
  assign \new_[17070]_  = ~A200 & A199;
  assign \new_[17071]_  = A166 & \new_[17070]_ ;
  assign \new_[17072]_  = \new_[17071]_  & \new_[17066]_ ;
  assign \new_[17076]_  = ~A266 & A202;
  assign \new_[17077]_  = A201 & \new_[17076]_ ;
  assign \new_[17081]_  = A299 & ~A298;
  assign \new_[17082]_  = ~A267 & \new_[17081]_ ;
  assign \new_[17083]_  = \new_[17082]_  & \new_[17077]_ ;
  assign \new_[17087]_  = A167 & ~A168;
  assign \new_[17088]_  = ~A169 & \new_[17087]_ ;
  assign \new_[17092]_  = ~A200 & A199;
  assign \new_[17093]_  = A166 & \new_[17092]_ ;
  assign \new_[17094]_  = \new_[17093]_  & \new_[17088]_ ;
  assign \new_[17098]_  = ~A265 & A202;
  assign \new_[17099]_  = A201 & \new_[17098]_ ;
  assign \new_[17103]_  = A299 & ~A298;
  assign \new_[17104]_  = ~A266 & \new_[17103]_ ;
  assign \new_[17105]_  = \new_[17104]_  & \new_[17099]_ ;
  assign \new_[17109]_  = A167 & ~A168;
  assign \new_[17110]_  = ~A169 & \new_[17109]_ ;
  assign \new_[17114]_  = ~A200 & A199;
  assign \new_[17115]_  = A166 & \new_[17114]_ ;
  assign \new_[17116]_  = \new_[17115]_  & \new_[17110]_ ;
  assign \new_[17120]_  = A265 & A203;
  assign \new_[17121]_  = A201 & \new_[17120]_ ;
  assign \new_[17125]_  = A299 & ~A298;
  assign \new_[17126]_  = A266 & \new_[17125]_ ;
  assign \new_[17127]_  = \new_[17126]_  & \new_[17121]_ ;
  assign \new_[17131]_  = A167 & ~A168;
  assign \new_[17132]_  = ~A169 & \new_[17131]_ ;
  assign \new_[17136]_  = ~A200 & A199;
  assign \new_[17137]_  = A166 & \new_[17136]_ ;
  assign \new_[17138]_  = \new_[17137]_  & \new_[17132]_ ;
  assign \new_[17142]_  = ~A266 & A203;
  assign \new_[17143]_  = A201 & \new_[17142]_ ;
  assign \new_[17147]_  = A299 & ~A298;
  assign \new_[17148]_  = ~A267 & \new_[17147]_ ;
  assign \new_[17149]_  = \new_[17148]_  & \new_[17143]_ ;
  assign \new_[17153]_  = A167 & ~A168;
  assign \new_[17154]_  = ~A169 & \new_[17153]_ ;
  assign \new_[17158]_  = ~A200 & A199;
  assign \new_[17159]_  = A166 & \new_[17158]_ ;
  assign \new_[17160]_  = \new_[17159]_  & \new_[17154]_ ;
  assign \new_[17164]_  = ~A265 & A203;
  assign \new_[17165]_  = A201 & \new_[17164]_ ;
  assign \new_[17169]_  = A299 & ~A298;
  assign \new_[17170]_  = ~A266 & \new_[17169]_ ;
  assign \new_[17171]_  = \new_[17170]_  & \new_[17165]_ ;
  assign \new_[17175]_  = A167 & ~A168;
  assign \new_[17176]_  = ~A169 & \new_[17175]_ ;
  assign \new_[17180]_  = ~A200 & ~A199;
  assign \new_[17181]_  = A166 & \new_[17180]_ ;
  assign \new_[17182]_  = \new_[17181]_  & \new_[17176]_ ;
  assign \new_[17186]_  = A267 & ~A266;
  assign \new_[17187]_  = A265 & \new_[17186]_ ;
  assign \new_[17191]_  = ~A300 & A298;
  assign \new_[17192]_  = A268 & \new_[17191]_ ;
  assign \new_[17193]_  = \new_[17192]_  & \new_[17187]_ ;
  assign \new_[17197]_  = A167 & ~A168;
  assign \new_[17198]_  = ~A169 & \new_[17197]_ ;
  assign \new_[17202]_  = ~A200 & ~A199;
  assign \new_[17203]_  = A166 & \new_[17202]_ ;
  assign \new_[17204]_  = \new_[17203]_  & \new_[17198]_ ;
  assign \new_[17208]_  = A267 & ~A266;
  assign \new_[17209]_  = A265 & \new_[17208]_ ;
  assign \new_[17213]_  = A299 & A298;
  assign \new_[17214]_  = A268 & \new_[17213]_ ;
  assign \new_[17215]_  = \new_[17214]_  & \new_[17209]_ ;
  assign \new_[17219]_  = A167 & ~A168;
  assign \new_[17220]_  = ~A169 & \new_[17219]_ ;
  assign \new_[17224]_  = ~A200 & ~A199;
  assign \new_[17225]_  = A166 & \new_[17224]_ ;
  assign \new_[17226]_  = \new_[17225]_  & \new_[17220]_ ;
  assign \new_[17230]_  = A267 & ~A266;
  assign \new_[17231]_  = A265 & \new_[17230]_ ;
  assign \new_[17235]_  = ~A299 & ~A298;
  assign \new_[17236]_  = A268 & \new_[17235]_ ;
  assign \new_[17237]_  = \new_[17236]_  & \new_[17231]_ ;
  assign \new_[17241]_  = A167 & ~A168;
  assign \new_[17242]_  = ~A169 & \new_[17241]_ ;
  assign \new_[17246]_  = ~A200 & ~A199;
  assign \new_[17247]_  = A166 & \new_[17246]_ ;
  assign \new_[17248]_  = \new_[17247]_  & \new_[17242]_ ;
  assign \new_[17252]_  = A267 & ~A266;
  assign \new_[17253]_  = A265 & \new_[17252]_ ;
  assign \new_[17257]_  = ~A300 & A298;
  assign \new_[17258]_  = A269 & \new_[17257]_ ;
  assign \new_[17259]_  = \new_[17258]_  & \new_[17253]_ ;
  assign \new_[17263]_  = A167 & ~A168;
  assign \new_[17264]_  = ~A169 & \new_[17263]_ ;
  assign \new_[17268]_  = ~A200 & ~A199;
  assign \new_[17269]_  = A166 & \new_[17268]_ ;
  assign \new_[17270]_  = \new_[17269]_  & \new_[17264]_ ;
  assign \new_[17274]_  = A267 & ~A266;
  assign \new_[17275]_  = A265 & \new_[17274]_ ;
  assign \new_[17279]_  = A299 & A298;
  assign \new_[17280]_  = A269 & \new_[17279]_ ;
  assign \new_[17281]_  = \new_[17280]_  & \new_[17275]_ ;
  assign \new_[17285]_  = A167 & ~A168;
  assign \new_[17286]_  = ~A169 & \new_[17285]_ ;
  assign \new_[17290]_  = ~A200 & ~A199;
  assign \new_[17291]_  = A166 & \new_[17290]_ ;
  assign \new_[17292]_  = \new_[17291]_  & \new_[17286]_ ;
  assign \new_[17296]_  = A267 & ~A266;
  assign \new_[17297]_  = A265 & \new_[17296]_ ;
  assign \new_[17301]_  = ~A299 & ~A298;
  assign \new_[17302]_  = A269 & \new_[17301]_ ;
  assign \new_[17303]_  = \new_[17302]_  & \new_[17297]_ ;
  assign \new_[17307]_  = A167 & ~A169;
  assign \new_[17308]_  = A170 & \new_[17307]_ ;
  assign \new_[17312]_  = A200 & A199;
  assign \new_[17313]_  = ~A166 & \new_[17312]_ ;
  assign \new_[17314]_  = \new_[17313]_  & \new_[17308]_ ;
  assign \new_[17318]_  = A298 & A266;
  assign \new_[17319]_  = A265 & \new_[17318]_ ;
  assign \new_[17323]_  = A301 & A300;
  assign \new_[17324]_  = ~A299 & \new_[17323]_ ;
  assign \new_[17325]_  = \new_[17324]_  & \new_[17319]_ ;
  assign \new_[17329]_  = A167 & ~A169;
  assign \new_[17330]_  = A170 & \new_[17329]_ ;
  assign \new_[17334]_  = A200 & A199;
  assign \new_[17335]_  = ~A166 & \new_[17334]_ ;
  assign \new_[17336]_  = \new_[17335]_  & \new_[17330]_ ;
  assign \new_[17340]_  = A298 & A266;
  assign \new_[17341]_  = A265 & \new_[17340]_ ;
  assign \new_[17345]_  = A302 & A300;
  assign \new_[17346]_  = ~A299 & \new_[17345]_ ;
  assign \new_[17347]_  = \new_[17346]_  & \new_[17341]_ ;
  assign \new_[17351]_  = A167 & ~A169;
  assign \new_[17352]_  = A170 & \new_[17351]_ ;
  assign \new_[17356]_  = A200 & A199;
  assign \new_[17357]_  = ~A166 & \new_[17356]_ ;
  assign \new_[17358]_  = \new_[17357]_  & \new_[17352]_ ;
  assign \new_[17362]_  = A298 & ~A267;
  assign \new_[17363]_  = ~A266 & \new_[17362]_ ;
  assign \new_[17367]_  = A301 & A300;
  assign \new_[17368]_  = ~A299 & \new_[17367]_ ;
  assign \new_[17369]_  = \new_[17368]_  & \new_[17363]_ ;
  assign \new_[17373]_  = A167 & ~A169;
  assign \new_[17374]_  = A170 & \new_[17373]_ ;
  assign \new_[17378]_  = A200 & A199;
  assign \new_[17379]_  = ~A166 & \new_[17378]_ ;
  assign \new_[17380]_  = \new_[17379]_  & \new_[17374]_ ;
  assign \new_[17384]_  = A298 & ~A267;
  assign \new_[17385]_  = ~A266 & \new_[17384]_ ;
  assign \new_[17389]_  = A302 & A300;
  assign \new_[17390]_  = ~A299 & \new_[17389]_ ;
  assign \new_[17391]_  = \new_[17390]_  & \new_[17385]_ ;
  assign \new_[17395]_  = A167 & ~A169;
  assign \new_[17396]_  = A170 & \new_[17395]_ ;
  assign \new_[17400]_  = A200 & A199;
  assign \new_[17401]_  = ~A166 & \new_[17400]_ ;
  assign \new_[17402]_  = \new_[17401]_  & \new_[17396]_ ;
  assign \new_[17406]_  = A298 & ~A266;
  assign \new_[17407]_  = ~A265 & \new_[17406]_ ;
  assign \new_[17411]_  = A301 & A300;
  assign \new_[17412]_  = ~A299 & \new_[17411]_ ;
  assign \new_[17413]_  = \new_[17412]_  & \new_[17407]_ ;
  assign \new_[17417]_  = A167 & ~A169;
  assign \new_[17418]_  = A170 & \new_[17417]_ ;
  assign \new_[17422]_  = A200 & A199;
  assign \new_[17423]_  = ~A166 & \new_[17422]_ ;
  assign \new_[17424]_  = \new_[17423]_  & \new_[17418]_ ;
  assign \new_[17428]_  = A298 & ~A266;
  assign \new_[17429]_  = ~A265 & \new_[17428]_ ;
  assign \new_[17433]_  = A302 & A300;
  assign \new_[17434]_  = ~A299 & \new_[17433]_ ;
  assign \new_[17435]_  = \new_[17434]_  & \new_[17429]_ ;
  assign \new_[17439]_  = A167 & ~A169;
  assign \new_[17440]_  = A170 & \new_[17439]_ ;
  assign \new_[17444]_  = A200 & ~A199;
  assign \new_[17445]_  = ~A166 & \new_[17444]_ ;
  assign \new_[17446]_  = \new_[17445]_  & \new_[17440]_ ;
  assign \new_[17450]_  = A267 & ~A266;
  assign \new_[17451]_  = A265 & \new_[17450]_ ;
  assign \new_[17455]_  = ~A300 & A298;
  assign \new_[17456]_  = A268 & \new_[17455]_ ;
  assign \new_[17457]_  = \new_[17456]_  & \new_[17451]_ ;
  assign \new_[17461]_  = A167 & ~A169;
  assign \new_[17462]_  = A170 & \new_[17461]_ ;
  assign \new_[17466]_  = A200 & ~A199;
  assign \new_[17467]_  = ~A166 & \new_[17466]_ ;
  assign \new_[17468]_  = \new_[17467]_  & \new_[17462]_ ;
  assign \new_[17472]_  = A267 & ~A266;
  assign \new_[17473]_  = A265 & \new_[17472]_ ;
  assign \new_[17477]_  = A299 & A298;
  assign \new_[17478]_  = A268 & \new_[17477]_ ;
  assign \new_[17479]_  = \new_[17478]_  & \new_[17473]_ ;
  assign \new_[17483]_  = A167 & ~A169;
  assign \new_[17484]_  = A170 & \new_[17483]_ ;
  assign \new_[17488]_  = A200 & ~A199;
  assign \new_[17489]_  = ~A166 & \new_[17488]_ ;
  assign \new_[17490]_  = \new_[17489]_  & \new_[17484]_ ;
  assign \new_[17494]_  = A267 & ~A266;
  assign \new_[17495]_  = A265 & \new_[17494]_ ;
  assign \new_[17499]_  = ~A299 & ~A298;
  assign \new_[17500]_  = A268 & \new_[17499]_ ;
  assign \new_[17501]_  = \new_[17500]_  & \new_[17495]_ ;
  assign \new_[17505]_  = A167 & ~A169;
  assign \new_[17506]_  = A170 & \new_[17505]_ ;
  assign \new_[17510]_  = A200 & ~A199;
  assign \new_[17511]_  = ~A166 & \new_[17510]_ ;
  assign \new_[17512]_  = \new_[17511]_  & \new_[17506]_ ;
  assign \new_[17516]_  = A267 & ~A266;
  assign \new_[17517]_  = A265 & \new_[17516]_ ;
  assign \new_[17521]_  = ~A300 & A298;
  assign \new_[17522]_  = A269 & \new_[17521]_ ;
  assign \new_[17523]_  = \new_[17522]_  & \new_[17517]_ ;
  assign \new_[17527]_  = A167 & ~A169;
  assign \new_[17528]_  = A170 & \new_[17527]_ ;
  assign \new_[17532]_  = A200 & ~A199;
  assign \new_[17533]_  = ~A166 & \new_[17532]_ ;
  assign \new_[17534]_  = \new_[17533]_  & \new_[17528]_ ;
  assign \new_[17538]_  = A267 & ~A266;
  assign \new_[17539]_  = A265 & \new_[17538]_ ;
  assign \new_[17543]_  = A299 & A298;
  assign \new_[17544]_  = A269 & \new_[17543]_ ;
  assign \new_[17545]_  = \new_[17544]_  & \new_[17539]_ ;
  assign \new_[17549]_  = A167 & ~A169;
  assign \new_[17550]_  = A170 & \new_[17549]_ ;
  assign \new_[17554]_  = A200 & ~A199;
  assign \new_[17555]_  = ~A166 & \new_[17554]_ ;
  assign \new_[17556]_  = \new_[17555]_  & \new_[17550]_ ;
  assign \new_[17560]_  = A267 & ~A266;
  assign \new_[17561]_  = A265 & \new_[17560]_ ;
  assign \new_[17565]_  = ~A299 & ~A298;
  assign \new_[17566]_  = A269 & \new_[17565]_ ;
  assign \new_[17567]_  = \new_[17566]_  & \new_[17561]_ ;
  assign \new_[17571]_  = A167 & ~A169;
  assign \new_[17572]_  = A170 & \new_[17571]_ ;
  assign \new_[17576]_  = ~A202 & ~A200;
  assign \new_[17577]_  = ~A166 & \new_[17576]_ ;
  assign \new_[17578]_  = \new_[17577]_  & \new_[17572]_ ;
  assign \new_[17582]_  = ~A268 & ~A266;
  assign \new_[17583]_  = ~A203 & \new_[17582]_ ;
  assign \new_[17587]_  = A299 & ~A298;
  assign \new_[17588]_  = ~A269 & \new_[17587]_ ;
  assign \new_[17589]_  = \new_[17588]_  & \new_[17583]_ ;
  assign \new_[17593]_  = A167 & ~A169;
  assign \new_[17594]_  = A170 & \new_[17593]_ ;
  assign \new_[17598]_  = ~A201 & ~A200;
  assign \new_[17599]_  = ~A166 & \new_[17598]_ ;
  assign \new_[17600]_  = \new_[17599]_  & \new_[17594]_ ;
  assign \new_[17604]_  = A298 & A266;
  assign \new_[17605]_  = A265 & \new_[17604]_ ;
  assign \new_[17609]_  = A301 & A300;
  assign \new_[17610]_  = ~A299 & \new_[17609]_ ;
  assign \new_[17611]_  = \new_[17610]_  & \new_[17605]_ ;
  assign \new_[17615]_  = A167 & ~A169;
  assign \new_[17616]_  = A170 & \new_[17615]_ ;
  assign \new_[17620]_  = ~A201 & ~A200;
  assign \new_[17621]_  = ~A166 & \new_[17620]_ ;
  assign \new_[17622]_  = \new_[17621]_  & \new_[17616]_ ;
  assign \new_[17626]_  = A298 & A266;
  assign \new_[17627]_  = A265 & \new_[17626]_ ;
  assign \new_[17631]_  = A302 & A300;
  assign \new_[17632]_  = ~A299 & \new_[17631]_ ;
  assign \new_[17633]_  = \new_[17632]_  & \new_[17627]_ ;
  assign \new_[17637]_  = A167 & ~A169;
  assign \new_[17638]_  = A170 & \new_[17637]_ ;
  assign \new_[17642]_  = ~A201 & ~A200;
  assign \new_[17643]_  = ~A166 & \new_[17642]_ ;
  assign \new_[17644]_  = \new_[17643]_  & \new_[17638]_ ;
  assign \new_[17648]_  = A298 & ~A267;
  assign \new_[17649]_  = ~A266 & \new_[17648]_ ;
  assign \new_[17653]_  = A301 & A300;
  assign \new_[17654]_  = ~A299 & \new_[17653]_ ;
  assign \new_[17655]_  = \new_[17654]_  & \new_[17649]_ ;
  assign \new_[17659]_  = A167 & ~A169;
  assign \new_[17660]_  = A170 & \new_[17659]_ ;
  assign \new_[17664]_  = ~A201 & ~A200;
  assign \new_[17665]_  = ~A166 & \new_[17664]_ ;
  assign \new_[17666]_  = \new_[17665]_  & \new_[17660]_ ;
  assign \new_[17670]_  = A298 & ~A267;
  assign \new_[17671]_  = ~A266 & \new_[17670]_ ;
  assign \new_[17675]_  = A302 & A300;
  assign \new_[17676]_  = ~A299 & \new_[17675]_ ;
  assign \new_[17677]_  = \new_[17676]_  & \new_[17671]_ ;
  assign \new_[17681]_  = A167 & ~A169;
  assign \new_[17682]_  = A170 & \new_[17681]_ ;
  assign \new_[17686]_  = ~A201 & ~A200;
  assign \new_[17687]_  = ~A166 & \new_[17686]_ ;
  assign \new_[17688]_  = \new_[17687]_  & \new_[17682]_ ;
  assign \new_[17692]_  = A298 & ~A266;
  assign \new_[17693]_  = ~A265 & \new_[17692]_ ;
  assign \new_[17697]_  = A301 & A300;
  assign \new_[17698]_  = ~A299 & \new_[17697]_ ;
  assign \new_[17699]_  = \new_[17698]_  & \new_[17693]_ ;
  assign \new_[17703]_  = A167 & ~A169;
  assign \new_[17704]_  = A170 & \new_[17703]_ ;
  assign \new_[17708]_  = ~A201 & ~A200;
  assign \new_[17709]_  = ~A166 & \new_[17708]_ ;
  assign \new_[17710]_  = \new_[17709]_  & \new_[17704]_ ;
  assign \new_[17714]_  = A298 & ~A266;
  assign \new_[17715]_  = ~A265 & \new_[17714]_ ;
  assign \new_[17719]_  = A302 & A300;
  assign \new_[17720]_  = ~A299 & \new_[17719]_ ;
  assign \new_[17721]_  = \new_[17720]_  & \new_[17715]_ ;
  assign \new_[17725]_  = A167 & ~A169;
  assign \new_[17726]_  = A170 & \new_[17725]_ ;
  assign \new_[17730]_  = ~A200 & A199;
  assign \new_[17731]_  = ~A166 & \new_[17730]_ ;
  assign \new_[17732]_  = \new_[17731]_  & \new_[17726]_ ;
  assign \new_[17736]_  = ~A265 & A202;
  assign \new_[17737]_  = A201 & \new_[17736]_ ;
  assign \new_[17741]_  = ~A300 & A298;
  assign \new_[17742]_  = A266 & \new_[17741]_ ;
  assign \new_[17743]_  = \new_[17742]_  & \new_[17737]_ ;
  assign \new_[17747]_  = A167 & ~A169;
  assign \new_[17748]_  = A170 & \new_[17747]_ ;
  assign \new_[17752]_  = ~A200 & A199;
  assign \new_[17753]_  = ~A166 & \new_[17752]_ ;
  assign \new_[17754]_  = \new_[17753]_  & \new_[17748]_ ;
  assign \new_[17758]_  = ~A265 & A202;
  assign \new_[17759]_  = A201 & \new_[17758]_ ;
  assign \new_[17763]_  = A299 & A298;
  assign \new_[17764]_  = A266 & \new_[17763]_ ;
  assign \new_[17765]_  = \new_[17764]_  & \new_[17759]_ ;
  assign \new_[17769]_  = A167 & ~A169;
  assign \new_[17770]_  = A170 & \new_[17769]_ ;
  assign \new_[17774]_  = ~A200 & A199;
  assign \new_[17775]_  = ~A166 & \new_[17774]_ ;
  assign \new_[17776]_  = \new_[17775]_  & \new_[17770]_ ;
  assign \new_[17780]_  = ~A265 & A202;
  assign \new_[17781]_  = A201 & \new_[17780]_ ;
  assign \new_[17785]_  = ~A299 & ~A298;
  assign \new_[17786]_  = A266 & \new_[17785]_ ;
  assign \new_[17787]_  = \new_[17786]_  & \new_[17781]_ ;
  assign \new_[17791]_  = A167 & ~A169;
  assign \new_[17792]_  = A170 & \new_[17791]_ ;
  assign \new_[17796]_  = ~A200 & A199;
  assign \new_[17797]_  = ~A166 & \new_[17796]_ ;
  assign \new_[17798]_  = \new_[17797]_  & \new_[17792]_ ;
  assign \new_[17802]_  = ~A265 & A203;
  assign \new_[17803]_  = A201 & \new_[17802]_ ;
  assign \new_[17807]_  = ~A300 & A298;
  assign \new_[17808]_  = A266 & \new_[17807]_ ;
  assign \new_[17809]_  = \new_[17808]_  & \new_[17803]_ ;
  assign \new_[17813]_  = A167 & ~A169;
  assign \new_[17814]_  = A170 & \new_[17813]_ ;
  assign \new_[17818]_  = ~A200 & A199;
  assign \new_[17819]_  = ~A166 & \new_[17818]_ ;
  assign \new_[17820]_  = \new_[17819]_  & \new_[17814]_ ;
  assign \new_[17824]_  = ~A265 & A203;
  assign \new_[17825]_  = A201 & \new_[17824]_ ;
  assign \new_[17829]_  = A299 & A298;
  assign \new_[17830]_  = A266 & \new_[17829]_ ;
  assign \new_[17831]_  = \new_[17830]_  & \new_[17825]_ ;
  assign \new_[17835]_  = A167 & ~A169;
  assign \new_[17836]_  = A170 & \new_[17835]_ ;
  assign \new_[17840]_  = ~A200 & A199;
  assign \new_[17841]_  = ~A166 & \new_[17840]_ ;
  assign \new_[17842]_  = \new_[17841]_  & \new_[17836]_ ;
  assign \new_[17846]_  = ~A265 & A203;
  assign \new_[17847]_  = A201 & \new_[17846]_ ;
  assign \new_[17851]_  = ~A299 & ~A298;
  assign \new_[17852]_  = A266 & \new_[17851]_ ;
  assign \new_[17853]_  = \new_[17852]_  & \new_[17847]_ ;
  assign \new_[17857]_  = A167 & ~A169;
  assign \new_[17858]_  = A170 & \new_[17857]_ ;
  assign \new_[17862]_  = ~A200 & ~A199;
  assign \new_[17863]_  = ~A166 & \new_[17862]_ ;
  assign \new_[17864]_  = \new_[17863]_  & \new_[17858]_ ;
  assign \new_[17868]_  = A298 & A266;
  assign \new_[17869]_  = A265 & \new_[17868]_ ;
  assign \new_[17873]_  = A301 & A300;
  assign \new_[17874]_  = ~A299 & \new_[17873]_ ;
  assign \new_[17875]_  = \new_[17874]_  & \new_[17869]_ ;
  assign \new_[17879]_  = A167 & ~A169;
  assign \new_[17880]_  = A170 & \new_[17879]_ ;
  assign \new_[17884]_  = ~A200 & ~A199;
  assign \new_[17885]_  = ~A166 & \new_[17884]_ ;
  assign \new_[17886]_  = \new_[17885]_  & \new_[17880]_ ;
  assign \new_[17890]_  = A298 & A266;
  assign \new_[17891]_  = A265 & \new_[17890]_ ;
  assign \new_[17895]_  = A302 & A300;
  assign \new_[17896]_  = ~A299 & \new_[17895]_ ;
  assign \new_[17897]_  = \new_[17896]_  & \new_[17891]_ ;
  assign \new_[17901]_  = A167 & ~A169;
  assign \new_[17902]_  = A170 & \new_[17901]_ ;
  assign \new_[17906]_  = ~A200 & ~A199;
  assign \new_[17907]_  = ~A166 & \new_[17906]_ ;
  assign \new_[17908]_  = \new_[17907]_  & \new_[17902]_ ;
  assign \new_[17912]_  = A298 & ~A267;
  assign \new_[17913]_  = ~A266 & \new_[17912]_ ;
  assign \new_[17917]_  = A301 & A300;
  assign \new_[17918]_  = ~A299 & \new_[17917]_ ;
  assign \new_[17919]_  = \new_[17918]_  & \new_[17913]_ ;
  assign \new_[17923]_  = A167 & ~A169;
  assign \new_[17924]_  = A170 & \new_[17923]_ ;
  assign \new_[17928]_  = ~A200 & ~A199;
  assign \new_[17929]_  = ~A166 & \new_[17928]_ ;
  assign \new_[17930]_  = \new_[17929]_  & \new_[17924]_ ;
  assign \new_[17934]_  = A298 & ~A267;
  assign \new_[17935]_  = ~A266 & \new_[17934]_ ;
  assign \new_[17939]_  = A302 & A300;
  assign \new_[17940]_  = ~A299 & \new_[17939]_ ;
  assign \new_[17941]_  = \new_[17940]_  & \new_[17935]_ ;
  assign \new_[17945]_  = A167 & ~A169;
  assign \new_[17946]_  = A170 & \new_[17945]_ ;
  assign \new_[17950]_  = ~A200 & ~A199;
  assign \new_[17951]_  = ~A166 & \new_[17950]_ ;
  assign \new_[17952]_  = \new_[17951]_  & \new_[17946]_ ;
  assign \new_[17956]_  = A298 & ~A266;
  assign \new_[17957]_  = ~A265 & \new_[17956]_ ;
  assign \new_[17961]_  = A301 & A300;
  assign \new_[17962]_  = ~A299 & \new_[17961]_ ;
  assign \new_[17963]_  = \new_[17962]_  & \new_[17957]_ ;
  assign \new_[17967]_  = A167 & ~A169;
  assign \new_[17968]_  = A170 & \new_[17967]_ ;
  assign \new_[17972]_  = ~A200 & ~A199;
  assign \new_[17973]_  = ~A166 & \new_[17972]_ ;
  assign \new_[17974]_  = \new_[17973]_  & \new_[17968]_ ;
  assign \new_[17978]_  = A298 & ~A266;
  assign \new_[17979]_  = ~A265 & \new_[17978]_ ;
  assign \new_[17983]_  = A302 & A300;
  assign \new_[17984]_  = ~A299 & \new_[17983]_ ;
  assign \new_[17985]_  = \new_[17984]_  & \new_[17979]_ ;
  assign \new_[17989]_  = ~A167 & ~A169;
  assign \new_[17990]_  = A170 & \new_[17989]_ ;
  assign \new_[17994]_  = A200 & A199;
  assign \new_[17995]_  = A166 & \new_[17994]_ ;
  assign \new_[17996]_  = \new_[17995]_  & \new_[17990]_ ;
  assign \new_[18000]_  = A298 & A266;
  assign \new_[18001]_  = A265 & \new_[18000]_ ;
  assign \new_[18005]_  = A301 & A300;
  assign \new_[18006]_  = ~A299 & \new_[18005]_ ;
  assign \new_[18007]_  = \new_[18006]_  & \new_[18001]_ ;
  assign \new_[18011]_  = ~A167 & ~A169;
  assign \new_[18012]_  = A170 & \new_[18011]_ ;
  assign \new_[18016]_  = A200 & A199;
  assign \new_[18017]_  = A166 & \new_[18016]_ ;
  assign \new_[18018]_  = \new_[18017]_  & \new_[18012]_ ;
  assign \new_[18022]_  = A298 & A266;
  assign \new_[18023]_  = A265 & \new_[18022]_ ;
  assign \new_[18027]_  = A302 & A300;
  assign \new_[18028]_  = ~A299 & \new_[18027]_ ;
  assign \new_[18029]_  = \new_[18028]_  & \new_[18023]_ ;
  assign \new_[18033]_  = ~A167 & ~A169;
  assign \new_[18034]_  = A170 & \new_[18033]_ ;
  assign \new_[18038]_  = A200 & A199;
  assign \new_[18039]_  = A166 & \new_[18038]_ ;
  assign \new_[18040]_  = \new_[18039]_  & \new_[18034]_ ;
  assign \new_[18044]_  = A298 & ~A267;
  assign \new_[18045]_  = ~A266 & \new_[18044]_ ;
  assign \new_[18049]_  = A301 & A300;
  assign \new_[18050]_  = ~A299 & \new_[18049]_ ;
  assign \new_[18051]_  = \new_[18050]_  & \new_[18045]_ ;
  assign \new_[18055]_  = ~A167 & ~A169;
  assign \new_[18056]_  = A170 & \new_[18055]_ ;
  assign \new_[18060]_  = A200 & A199;
  assign \new_[18061]_  = A166 & \new_[18060]_ ;
  assign \new_[18062]_  = \new_[18061]_  & \new_[18056]_ ;
  assign \new_[18066]_  = A298 & ~A267;
  assign \new_[18067]_  = ~A266 & \new_[18066]_ ;
  assign \new_[18071]_  = A302 & A300;
  assign \new_[18072]_  = ~A299 & \new_[18071]_ ;
  assign \new_[18073]_  = \new_[18072]_  & \new_[18067]_ ;
  assign \new_[18077]_  = ~A167 & ~A169;
  assign \new_[18078]_  = A170 & \new_[18077]_ ;
  assign \new_[18082]_  = A200 & A199;
  assign \new_[18083]_  = A166 & \new_[18082]_ ;
  assign \new_[18084]_  = \new_[18083]_  & \new_[18078]_ ;
  assign \new_[18088]_  = A298 & ~A266;
  assign \new_[18089]_  = ~A265 & \new_[18088]_ ;
  assign \new_[18093]_  = A301 & A300;
  assign \new_[18094]_  = ~A299 & \new_[18093]_ ;
  assign \new_[18095]_  = \new_[18094]_  & \new_[18089]_ ;
  assign \new_[18099]_  = ~A167 & ~A169;
  assign \new_[18100]_  = A170 & \new_[18099]_ ;
  assign \new_[18104]_  = A200 & A199;
  assign \new_[18105]_  = A166 & \new_[18104]_ ;
  assign \new_[18106]_  = \new_[18105]_  & \new_[18100]_ ;
  assign \new_[18110]_  = A298 & ~A266;
  assign \new_[18111]_  = ~A265 & \new_[18110]_ ;
  assign \new_[18115]_  = A302 & A300;
  assign \new_[18116]_  = ~A299 & \new_[18115]_ ;
  assign \new_[18117]_  = \new_[18116]_  & \new_[18111]_ ;
  assign \new_[18121]_  = ~A167 & ~A169;
  assign \new_[18122]_  = A170 & \new_[18121]_ ;
  assign \new_[18126]_  = A200 & ~A199;
  assign \new_[18127]_  = A166 & \new_[18126]_ ;
  assign \new_[18128]_  = \new_[18127]_  & \new_[18122]_ ;
  assign \new_[18132]_  = A267 & ~A266;
  assign \new_[18133]_  = A265 & \new_[18132]_ ;
  assign \new_[18137]_  = ~A300 & A298;
  assign \new_[18138]_  = A268 & \new_[18137]_ ;
  assign \new_[18139]_  = \new_[18138]_  & \new_[18133]_ ;
  assign \new_[18143]_  = ~A167 & ~A169;
  assign \new_[18144]_  = A170 & \new_[18143]_ ;
  assign \new_[18148]_  = A200 & ~A199;
  assign \new_[18149]_  = A166 & \new_[18148]_ ;
  assign \new_[18150]_  = \new_[18149]_  & \new_[18144]_ ;
  assign \new_[18154]_  = A267 & ~A266;
  assign \new_[18155]_  = A265 & \new_[18154]_ ;
  assign \new_[18159]_  = A299 & A298;
  assign \new_[18160]_  = A268 & \new_[18159]_ ;
  assign \new_[18161]_  = \new_[18160]_  & \new_[18155]_ ;
  assign \new_[18165]_  = ~A167 & ~A169;
  assign \new_[18166]_  = A170 & \new_[18165]_ ;
  assign \new_[18170]_  = A200 & ~A199;
  assign \new_[18171]_  = A166 & \new_[18170]_ ;
  assign \new_[18172]_  = \new_[18171]_  & \new_[18166]_ ;
  assign \new_[18176]_  = A267 & ~A266;
  assign \new_[18177]_  = A265 & \new_[18176]_ ;
  assign \new_[18181]_  = ~A299 & ~A298;
  assign \new_[18182]_  = A268 & \new_[18181]_ ;
  assign \new_[18183]_  = \new_[18182]_  & \new_[18177]_ ;
  assign \new_[18187]_  = ~A167 & ~A169;
  assign \new_[18188]_  = A170 & \new_[18187]_ ;
  assign \new_[18192]_  = A200 & ~A199;
  assign \new_[18193]_  = A166 & \new_[18192]_ ;
  assign \new_[18194]_  = \new_[18193]_  & \new_[18188]_ ;
  assign \new_[18198]_  = A267 & ~A266;
  assign \new_[18199]_  = A265 & \new_[18198]_ ;
  assign \new_[18203]_  = ~A300 & A298;
  assign \new_[18204]_  = A269 & \new_[18203]_ ;
  assign \new_[18205]_  = \new_[18204]_  & \new_[18199]_ ;
  assign \new_[18209]_  = ~A167 & ~A169;
  assign \new_[18210]_  = A170 & \new_[18209]_ ;
  assign \new_[18214]_  = A200 & ~A199;
  assign \new_[18215]_  = A166 & \new_[18214]_ ;
  assign \new_[18216]_  = \new_[18215]_  & \new_[18210]_ ;
  assign \new_[18220]_  = A267 & ~A266;
  assign \new_[18221]_  = A265 & \new_[18220]_ ;
  assign \new_[18225]_  = A299 & A298;
  assign \new_[18226]_  = A269 & \new_[18225]_ ;
  assign \new_[18227]_  = \new_[18226]_  & \new_[18221]_ ;
  assign \new_[18231]_  = ~A167 & ~A169;
  assign \new_[18232]_  = A170 & \new_[18231]_ ;
  assign \new_[18236]_  = A200 & ~A199;
  assign \new_[18237]_  = A166 & \new_[18236]_ ;
  assign \new_[18238]_  = \new_[18237]_  & \new_[18232]_ ;
  assign \new_[18242]_  = A267 & ~A266;
  assign \new_[18243]_  = A265 & \new_[18242]_ ;
  assign \new_[18247]_  = ~A299 & ~A298;
  assign \new_[18248]_  = A269 & \new_[18247]_ ;
  assign \new_[18249]_  = \new_[18248]_  & \new_[18243]_ ;
  assign \new_[18253]_  = ~A167 & ~A169;
  assign \new_[18254]_  = A170 & \new_[18253]_ ;
  assign \new_[18258]_  = ~A202 & ~A200;
  assign \new_[18259]_  = A166 & \new_[18258]_ ;
  assign \new_[18260]_  = \new_[18259]_  & \new_[18254]_ ;
  assign \new_[18264]_  = ~A268 & ~A266;
  assign \new_[18265]_  = ~A203 & \new_[18264]_ ;
  assign \new_[18269]_  = A299 & ~A298;
  assign \new_[18270]_  = ~A269 & \new_[18269]_ ;
  assign \new_[18271]_  = \new_[18270]_  & \new_[18265]_ ;
  assign \new_[18275]_  = ~A167 & ~A169;
  assign \new_[18276]_  = A170 & \new_[18275]_ ;
  assign \new_[18280]_  = ~A201 & ~A200;
  assign \new_[18281]_  = A166 & \new_[18280]_ ;
  assign \new_[18282]_  = \new_[18281]_  & \new_[18276]_ ;
  assign \new_[18286]_  = A298 & A266;
  assign \new_[18287]_  = A265 & \new_[18286]_ ;
  assign \new_[18291]_  = A301 & A300;
  assign \new_[18292]_  = ~A299 & \new_[18291]_ ;
  assign \new_[18293]_  = \new_[18292]_  & \new_[18287]_ ;
  assign \new_[18297]_  = ~A167 & ~A169;
  assign \new_[18298]_  = A170 & \new_[18297]_ ;
  assign \new_[18302]_  = ~A201 & ~A200;
  assign \new_[18303]_  = A166 & \new_[18302]_ ;
  assign \new_[18304]_  = \new_[18303]_  & \new_[18298]_ ;
  assign \new_[18308]_  = A298 & A266;
  assign \new_[18309]_  = A265 & \new_[18308]_ ;
  assign \new_[18313]_  = A302 & A300;
  assign \new_[18314]_  = ~A299 & \new_[18313]_ ;
  assign \new_[18315]_  = \new_[18314]_  & \new_[18309]_ ;
  assign \new_[18319]_  = ~A167 & ~A169;
  assign \new_[18320]_  = A170 & \new_[18319]_ ;
  assign \new_[18324]_  = ~A201 & ~A200;
  assign \new_[18325]_  = A166 & \new_[18324]_ ;
  assign \new_[18326]_  = \new_[18325]_  & \new_[18320]_ ;
  assign \new_[18330]_  = A298 & ~A267;
  assign \new_[18331]_  = ~A266 & \new_[18330]_ ;
  assign \new_[18335]_  = A301 & A300;
  assign \new_[18336]_  = ~A299 & \new_[18335]_ ;
  assign \new_[18337]_  = \new_[18336]_  & \new_[18331]_ ;
  assign \new_[18341]_  = ~A167 & ~A169;
  assign \new_[18342]_  = A170 & \new_[18341]_ ;
  assign \new_[18346]_  = ~A201 & ~A200;
  assign \new_[18347]_  = A166 & \new_[18346]_ ;
  assign \new_[18348]_  = \new_[18347]_  & \new_[18342]_ ;
  assign \new_[18352]_  = A298 & ~A267;
  assign \new_[18353]_  = ~A266 & \new_[18352]_ ;
  assign \new_[18357]_  = A302 & A300;
  assign \new_[18358]_  = ~A299 & \new_[18357]_ ;
  assign \new_[18359]_  = \new_[18358]_  & \new_[18353]_ ;
  assign \new_[18363]_  = ~A167 & ~A169;
  assign \new_[18364]_  = A170 & \new_[18363]_ ;
  assign \new_[18368]_  = ~A201 & ~A200;
  assign \new_[18369]_  = A166 & \new_[18368]_ ;
  assign \new_[18370]_  = \new_[18369]_  & \new_[18364]_ ;
  assign \new_[18374]_  = A298 & ~A266;
  assign \new_[18375]_  = ~A265 & \new_[18374]_ ;
  assign \new_[18379]_  = A301 & A300;
  assign \new_[18380]_  = ~A299 & \new_[18379]_ ;
  assign \new_[18381]_  = \new_[18380]_  & \new_[18375]_ ;
  assign \new_[18385]_  = ~A167 & ~A169;
  assign \new_[18386]_  = A170 & \new_[18385]_ ;
  assign \new_[18390]_  = ~A201 & ~A200;
  assign \new_[18391]_  = A166 & \new_[18390]_ ;
  assign \new_[18392]_  = \new_[18391]_  & \new_[18386]_ ;
  assign \new_[18396]_  = A298 & ~A266;
  assign \new_[18397]_  = ~A265 & \new_[18396]_ ;
  assign \new_[18401]_  = A302 & A300;
  assign \new_[18402]_  = ~A299 & \new_[18401]_ ;
  assign \new_[18403]_  = \new_[18402]_  & \new_[18397]_ ;
  assign \new_[18407]_  = ~A167 & ~A169;
  assign \new_[18408]_  = A170 & \new_[18407]_ ;
  assign \new_[18412]_  = ~A200 & A199;
  assign \new_[18413]_  = A166 & \new_[18412]_ ;
  assign \new_[18414]_  = \new_[18413]_  & \new_[18408]_ ;
  assign \new_[18418]_  = ~A265 & A202;
  assign \new_[18419]_  = A201 & \new_[18418]_ ;
  assign \new_[18423]_  = ~A300 & A298;
  assign \new_[18424]_  = A266 & \new_[18423]_ ;
  assign \new_[18425]_  = \new_[18424]_  & \new_[18419]_ ;
  assign \new_[18429]_  = ~A167 & ~A169;
  assign \new_[18430]_  = A170 & \new_[18429]_ ;
  assign \new_[18434]_  = ~A200 & A199;
  assign \new_[18435]_  = A166 & \new_[18434]_ ;
  assign \new_[18436]_  = \new_[18435]_  & \new_[18430]_ ;
  assign \new_[18440]_  = ~A265 & A202;
  assign \new_[18441]_  = A201 & \new_[18440]_ ;
  assign \new_[18445]_  = A299 & A298;
  assign \new_[18446]_  = A266 & \new_[18445]_ ;
  assign \new_[18447]_  = \new_[18446]_  & \new_[18441]_ ;
  assign \new_[18451]_  = ~A167 & ~A169;
  assign \new_[18452]_  = A170 & \new_[18451]_ ;
  assign \new_[18456]_  = ~A200 & A199;
  assign \new_[18457]_  = A166 & \new_[18456]_ ;
  assign \new_[18458]_  = \new_[18457]_  & \new_[18452]_ ;
  assign \new_[18462]_  = ~A265 & A202;
  assign \new_[18463]_  = A201 & \new_[18462]_ ;
  assign \new_[18467]_  = ~A299 & ~A298;
  assign \new_[18468]_  = A266 & \new_[18467]_ ;
  assign \new_[18469]_  = \new_[18468]_  & \new_[18463]_ ;
  assign \new_[18473]_  = ~A167 & ~A169;
  assign \new_[18474]_  = A170 & \new_[18473]_ ;
  assign \new_[18478]_  = ~A200 & A199;
  assign \new_[18479]_  = A166 & \new_[18478]_ ;
  assign \new_[18480]_  = \new_[18479]_  & \new_[18474]_ ;
  assign \new_[18484]_  = ~A265 & A203;
  assign \new_[18485]_  = A201 & \new_[18484]_ ;
  assign \new_[18489]_  = ~A300 & A298;
  assign \new_[18490]_  = A266 & \new_[18489]_ ;
  assign \new_[18491]_  = \new_[18490]_  & \new_[18485]_ ;
  assign \new_[18495]_  = ~A167 & ~A169;
  assign \new_[18496]_  = A170 & \new_[18495]_ ;
  assign \new_[18500]_  = ~A200 & A199;
  assign \new_[18501]_  = A166 & \new_[18500]_ ;
  assign \new_[18502]_  = \new_[18501]_  & \new_[18496]_ ;
  assign \new_[18506]_  = ~A265 & A203;
  assign \new_[18507]_  = A201 & \new_[18506]_ ;
  assign \new_[18511]_  = A299 & A298;
  assign \new_[18512]_  = A266 & \new_[18511]_ ;
  assign \new_[18513]_  = \new_[18512]_  & \new_[18507]_ ;
  assign \new_[18517]_  = ~A167 & ~A169;
  assign \new_[18518]_  = A170 & \new_[18517]_ ;
  assign \new_[18522]_  = ~A200 & A199;
  assign \new_[18523]_  = A166 & \new_[18522]_ ;
  assign \new_[18524]_  = \new_[18523]_  & \new_[18518]_ ;
  assign \new_[18528]_  = ~A265 & A203;
  assign \new_[18529]_  = A201 & \new_[18528]_ ;
  assign \new_[18533]_  = ~A299 & ~A298;
  assign \new_[18534]_  = A266 & \new_[18533]_ ;
  assign \new_[18535]_  = \new_[18534]_  & \new_[18529]_ ;
  assign \new_[18539]_  = ~A167 & ~A169;
  assign \new_[18540]_  = A170 & \new_[18539]_ ;
  assign \new_[18544]_  = ~A200 & ~A199;
  assign \new_[18545]_  = A166 & \new_[18544]_ ;
  assign \new_[18546]_  = \new_[18545]_  & \new_[18540]_ ;
  assign \new_[18550]_  = A298 & A266;
  assign \new_[18551]_  = A265 & \new_[18550]_ ;
  assign \new_[18555]_  = A301 & A300;
  assign \new_[18556]_  = ~A299 & \new_[18555]_ ;
  assign \new_[18557]_  = \new_[18556]_  & \new_[18551]_ ;
  assign \new_[18561]_  = ~A167 & ~A169;
  assign \new_[18562]_  = A170 & \new_[18561]_ ;
  assign \new_[18566]_  = ~A200 & ~A199;
  assign \new_[18567]_  = A166 & \new_[18566]_ ;
  assign \new_[18568]_  = \new_[18567]_  & \new_[18562]_ ;
  assign \new_[18572]_  = A298 & A266;
  assign \new_[18573]_  = A265 & \new_[18572]_ ;
  assign \new_[18577]_  = A302 & A300;
  assign \new_[18578]_  = ~A299 & \new_[18577]_ ;
  assign \new_[18579]_  = \new_[18578]_  & \new_[18573]_ ;
  assign \new_[18583]_  = ~A167 & ~A169;
  assign \new_[18584]_  = A170 & \new_[18583]_ ;
  assign \new_[18588]_  = ~A200 & ~A199;
  assign \new_[18589]_  = A166 & \new_[18588]_ ;
  assign \new_[18590]_  = \new_[18589]_  & \new_[18584]_ ;
  assign \new_[18594]_  = A298 & ~A267;
  assign \new_[18595]_  = ~A266 & \new_[18594]_ ;
  assign \new_[18599]_  = A301 & A300;
  assign \new_[18600]_  = ~A299 & \new_[18599]_ ;
  assign \new_[18601]_  = \new_[18600]_  & \new_[18595]_ ;
  assign \new_[18605]_  = ~A167 & ~A169;
  assign \new_[18606]_  = A170 & \new_[18605]_ ;
  assign \new_[18610]_  = ~A200 & ~A199;
  assign \new_[18611]_  = A166 & \new_[18610]_ ;
  assign \new_[18612]_  = \new_[18611]_  & \new_[18606]_ ;
  assign \new_[18616]_  = A298 & ~A267;
  assign \new_[18617]_  = ~A266 & \new_[18616]_ ;
  assign \new_[18621]_  = A302 & A300;
  assign \new_[18622]_  = ~A299 & \new_[18621]_ ;
  assign \new_[18623]_  = \new_[18622]_  & \new_[18617]_ ;
  assign \new_[18627]_  = ~A167 & ~A169;
  assign \new_[18628]_  = A170 & \new_[18627]_ ;
  assign \new_[18632]_  = ~A200 & ~A199;
  assign \new_[18633]_  = A166 & \new_[18632]_ ;
  assign \new_[18634]_  = \new_[18633]_  & \new_[18628]_ ;
  assign \new_[18638]_  = A298 & ~A266;
  assign \new_[18639]_  = ~A265 & \new_[18638]_ ;
  assign \new_[18643]_  = A301 & A300;
  assign \new_[18644]_  = ~A299 & \new_[18643]_ ;
  assign \new_[18645]_  = \new_[18644]_  & \new_[18639]_ ;
  assign \new_[18649]_  = ~A167 & ~A169;
  assign \new_[18650]_  = A170 & \new_[18649]_ ;
  assign \new_[18654]_  = ~A200 & ~A199;
  assign \new_[18655]_  = A166 & \new_[18654]_ ;
  assign \new_[18656]_  = \new_[18655]_  & \new_[18650]_ ;
  assign \new_[18660]_  = A298 & ~A266;
  assign \new_[18661]_  = ~A265 & \new_[18660]_ ;
  assign \new_[18665]_  = A302 & A300;
  assign \new_[18666]_  = ~A299 & \new_[18665]_ ;
  assign \new_[18667]_  = \new_[18666]_  & \new_[18661]_ ;
  assign \new_[18671]_  = ~A168 & ~A169;
  assign \new_[18672]_  = ~A170 & \new_[18671]_ ;
  assign \new_[18676]_  = A265 & A200;
  assign \new_[18677]_  = A199 & \new_[18676]_ ;
  assign \new_[18678]_  = \new_[18677]_  & \new_[18672]_ ;
  assign \new_[18682]_  = A268 & A267;
  assign \new_[18683]_  = ~A266 & \new_[18682]_ ;
  assign \new_[18687]_  = ~A302 & ~A301;
  assign \new_[18688]_  = A298 & \new_[18687]_ ;
  assign \new_[18689]_  = \new_[18688]_  & \new_[18683]_ ;
  assign \new_[18693]_  = ~A168 & ~A169;
  assign \new_[18694]_  = ~A170 & \new_[18693]_ ;
  assign \new_[18698]_  = A265 & A200;
  assign \new_[18699]_  = A199 & \new_[18698]_ ;
  assign \new_[18700]_  = \new_[18699]_  & \new_[18694]_ ;
  assign \new_[18704]_  = A269 & A267;
  assign \new_[18705]_  = ~A266 & \new_[18704]_ ;
  assign \new_[18709]_  = ~A302 & ~A301;
  assign \new_[18710]_  = A298 & \new_[18709]_ ;
  assign \new_[18711]_  = \new_[18710]_  & \new_[18705]_ ;
  assign \new_[18715]_  = ~A168 & ~A169;
  assign \new_[18716]_  = ~A170 & \new_[18715]_ ;
  assign \new_[18720]_  = ~A266 & A200;
  assign \new_[18721]_  = ~A199 & \new_[18720]_ ;
  assign \new_[18722]_  = \new_[18721]_  & \new_[18716]_ ;
  assign \new_[18726]_  = A298 & ~A269;
  assign \new_[18727]_  = ~A268 & \new_[18726]_ ;
  assign \new_[18731]_  = A301 & A300;
  assign \new_[18732]_  = ~A299 & \new_[18731]_ ;
  assign \new_[18733]_  = \new_[18732]_  & \new_[18727]_ ;
  assign \new_[18737]_  = ~A168 & ~A169;
  assign \new_[18738]_  = ~A170 & \new_[18737]_ ;
  assign \new_[18742]_  = ~A266 & A200;
  assign \new_[18743]_  = ~A199 & \new_[18742]_ ;
  assign \new_[18744]_  = \new_[18743]_  & \new_[18738]_ ;
  assign \new_[18748]_  = A298 & ~A269;
  assign \new_[18749]_  = ~A268 & \new_[18748]_ ;
  assign \new_[18753]_  = A302 & A300;
  assign \new_[18754]_  = ~A299 & \new_[18753]_ ;
  assign \new_[18755]_  = \new_[18754]_  & \new_[18749]_ ;
  assign \new_[18759]_  = ~A168 & ~A169;
  assign \new_[18760]_  = ~A170 & \new_[18759]_ ;
  assign \new_[18764]_  = ~A203 & ~A202;
  assign \new_[18765]_  = ~A200 & \new_[18764]_ ;
  assign \new_[18766]_  = \new_[18765]_  & \new_[18760]_ ;
  assign \new_[18770]_  = A267 & ~A266;
  assign \new_[18771]_  = A265 & \new_[18770]_ ;
  assign \new_[18775]_  = ~A300 & A298;
  assign \new_[18776]_  = A268 & \new_[18775]_ ;
  assign \new_[18777]_  = \new_[18776]_  & \new_[18771]_ ;
  assign \new_[18781]_  = ~A168 & ~A169;
  assign \new_[18782]_  = ~A170 & \new_[18781]_ ;
  assign \new_[18786]_  = ~A203 & ~A202;
  assign \new_[18787]_  = ~A200 & \new_[18786]_ ;
  assign \new_[18788]_  = \new_[18787]_  & \new_[18782]_ ;
  assign \new_[18792]_  = A267 & ~A266;
  assign \new_[18793]_  = A265 & \new_[18792]_ ;
  assign \new_[18797]_  = A299 & A298;
  assign \new_[18798]_  = A268 & \new_[18797]_ ;
  assign \new_[18799]_  = \new_[18798]_  & \new_[18793]_ ;
  assign \new_[18803]_  = ~A168 & ~A169;
  assign \new_[18804]_  = ~A170 & \new_[18803]_ ;
  assign \new_[18808]_  = ~A203 & ~A202;
  assign \new_[18809]_  = ~A200 & \new_[18808]_ ;
  assign \new_[18810]_  = \new_[18809]_  & \new_[18804]_ ;
  assign \new_[18814]_  = A267 & ~A266;
  assign \new_[18815]_  = A265 & \new_[18814]_ ;
  assign \new_[18819]_  = ~A299 & ~A298;
  assign \new_[18820]_  = A268 & \new_[18819]_ ;
  assign \new_[18821]_  = \new_[18820]_  & \new_[18815]_ ;
  assign \new_[18825]_  = ~A168 & ~A169;
  assign \new_[18826]_  = ~A170 & \new_[18825]_ ;
  assign \new_[18830]_  = ~A203 & ~A202;
  assign \new_[18831]_  = ~A200 & \new_[18830]_ ;
  assign \new_[18832]_  = \new_[18831]_  & \new_[18826]_ ;
  assign \new_[18836]_  = A267 & ~A266;
  assign \new_[18837]_  = A265 & \new_[18836]_ ;
  assign \new_[18841]_  = ~A300 & A298;
  assign \new_[18842]_  = A269 & \new_[18841]_ ;
  assign \new_[18843]_  = \new_[18842]_  & \new_[18837]_ ;
  assign \new_[18847]_  = ~A168 & ~A169;
  assign \new_[18848]_  = ~A170 & \new_[18847]_ ;
  assign \new_[18852]_  = ~A203 & ~A202;
  assign \new_[18853]_  = ~A200 & \new_[18852]_ ;
  assign \new_[18854]_  = \new_[18853]_  & \new_[18848]_ ;
  assign \new_[18858]_  = A267 & ~A266;
  assign \new_[18859]_  = A265 & \new_[18858]_ ;
  assign \new_[18863]_  = A299 & A298;
  assign \new_[18864]_  = A269 & \new_[18863]_ ;
  assign \new_[18865]_  = \new_[18864]_  & \new_[18859]_ ;
  assign \new_[18869]_  = ~A168 & ~A169;
  assign \new_[18870]_  = ~A170 & \new_[18869]_ ;
  assign \new_[18874]_  = ~A203 & ~A202;
  assign \new_[18875]_  = ~A200 & \new_[18874]_ ;
  assign \new_[18876]_  = \new_[18875]_  & \new_[18870]_ ;
  assign \new_[18880]_  = A267 & ~A266;
  assign \new_[18881]_  = A265 & \new_[18880]_ ;
  assign \new_[18885]_  = ~A299 & ~A298;
  assign \new_[18886]_  = A269 & \new_[18885]_ ;
  assign \new_[18887]_  = \new_[18886]_  & \new_[18881]_ ;
  assign \new_[18891]_  = ~A168 & ~A169;
  assign \new_[18892]_  = ~A170 & \new_[18891]_ ;
  assign \new_[18896]_  = A265 & ~A201;
  assign \new_[18897]_  = ~A200 & \new_[18896]_ ;
  assign \new_[18898]_  = \new_[18897]_  & \new_[18892]_ ;
  assign \new_[18902]_  = A268 & A267;
  assign \new_[18903]_  = ~A266 & \new_[18902]_ ;
  assign \new_[18907]_  = ~A302 & ~A301;
  assign \new_[18908]_  = A298 & \new_[18907]_ ;
  assign \new_[18909]_  = \new_[18908]_  & \new_[18903]_ ;
  assign \new_[18913]_  = ~A168 & ~A169;
  assign \new_[18914]_  = ~A170 & \new_[18913]_ ;
  assign \new_[18918]_  = A265 & ~A201;
  assign \new_[18919]_  = ~A200 & \new_[18918]_ ;
  assign \new_[18920]_  = \new_[18919]_  & \new_[18914]_ ;
  assign \new_[18924]_  = A269 & A267;
  assign \new_[18925]_  = ~A266 & \new_[18924]_ ;
  assign \new_[18929]_  = ~A302 & ~A301;
  assign \new_[18930]_  = A298 & \new_[18929]_ ;
  assign \new_[18931]_  = \new_[18930]_  & \new_[18925]_ ;
  assign \new_[18935]_  = ~A168 & ~A169;
  assign \new_[18936]_  = ~A170 & \new_[18935]_ ;
  assign \new_[18940]_  = A201 & ~A200;
  assign \new_[18941]_  = A199 & \new_[18940]_ ;
  assign \new_[18942]_  = \new_[18941]_  & \new_[18936]_ ;
  assign \new_[18946]_  = ~A268 & ~A266;
  assign \new_[18947]_  = A202 & \new_[18946]_ ;
  assign \new_[18951]_  = A299 & ~A298;
  assign \new_[18952]_  = ~A269 & \new_[18951]_ ;
  assign \new_[18953]_  = \new_[18952]_  & \new_[18947]_ ;
  assign \new_[18957]_  = ~A168 & ~A169;
  assign \new_[18958]_  = ~A170 & \new_[18957]_ ;
  assign \new_[18962]_  = A201 & ~A200;
  assign \new_[18963]_  = A199 & \new_[18962]_ ;
  assign \new_[18964]_  = \new_[18963]_  & \new_[18958]_ ;
  assign \new_[18968]_  = ~A268 & ~A266;
  assign \new_[18969]_  = A203 & \new_[18968]_ ;
  assign \new_[18973]_  = A299 & ~A298;
  assign \new_[18974]_  = ~A269 & \new_[18973]_ ;
  assign \new_[18975]_  = \new_[18974]_  & \new_[18969]_ ;
  assign \new_[18979]_  = ~A168 & ~A169;
  assign \new_[18980]_  = ~A170 & \new_[18979]_ ;
  assign \new_[18984]_  = A265 & ~A200;
  assign \new_[18985]_  = ~A199 & \new_[18984]_ ;
  assign \new_[18986]_  = \new_[18985]_  & \new_[18980]_ ;
  assign \new_[18990]_  = A268 & A267;
  assign \new_[18991]_  = ~A266 & \new_[18990]_ ;
  assign \new_[18995]_  = ~A302 & ~A301;
  assign \new_[18996]_  = A298 & \new_[18995]_ ;
  assign \new_[18997]_  = \new_[18996]_  & \new_[18991]_ ;
  assign \new_[19001]_  = ~A168 & ~A169;
  assign \new_[19002]_  = ~A170 & \new_[19001]_ ;
  assign \new_[19006]_  = A265 & ~A200;
  assign \new_[19007]_  = ~A199 & \new_[19006]_ ;
  assign \new_[19008]_  = \new_[19007]_  & \new_[19002]_ ;
  assign \new_[19012]_  = A269 & A267;
  assign \new_[19013]_  = ~A266 & \new_[19012]_ ;
  assign \new_[19017]_  = ~A302 & ~A301;
  assign \new_[19018]_  = A298 & \new_[19017]_ ;
  assign \new_[19019]_  = \new_[19018]_  & \new_[19013]_ ;
  assign \new_[19023]_  = A199 & A166;
  assign \new_[19024]_  = A168 & \new_[19023]_ ;
  assign \new_[19028]_  = A202 & A201;
  assign \new_[19029]_  = ~A200 & \new_[19028]_ ;
  assign \new_[19030]_  = \new_[19029]_  & \new_[19024]_ ;
  assign \new_[19034]_  = A267 & ~A266;
  assign \new_[19035]_  = A265 & \new_[19034]_ ;
  assign \new_[19038]_  = A298 & A268;
  assign \new_[19041]_  = ~A302 & ~A301;
  assign \new_[19042]_  = \new_[19041]_  & \new_[19038]_ ;
  assign \new_[19043]_  = \new_[19042]_  & \new_[19035]_ ;
  assign \new_[19047]_  = A199 & A166;
  assign \new_[19048]_  = A168 & \new_[19047]_ ;
  assign \new_[19052]_  = A202 & A201;
  assign \new_[19053]_  = ~A200 & \new_[19052]_ ;
  assign \new_[19054]_  = \new_[19053]_  & \new_[19048]_ ;
  assign \new_[19058]_  = A267 & ~A266;
  assign \new_[19059]_  = A265 & \new_[19058]_ ;
  assign \new_[19062]_  = A298 & A269;
  assign \new_[19065]_  = ~A302 & ~A301;
  assign \new_[19066]_  = \new_[19065]_  & \new_[19062]_ ;
  assign \new_[19067]_  = \new_[19066]_  & \new_[19059]_ ;
  assign \new_[19071]_  = A199 & A166;
  assign \new_[19072]_  = A168 & \new_[19071]_ ;
  assign \new_[19076]_  = A203 & A201;
  assign \new_[19077]_  = ~A200 & \new_[19076]_ ;
  assign \new_[19078]_  = \new_[19077]_  & \new_[19072]_ ;
  assign \new_[19082]_  = A267 & ~A266;
  assign \new_[19083]_  = A265 & \new_[19082]_ ;
  assign \new_[19086]_  = A298 & A268;
  assign \new_[19089]_  = ~A302 & ~A301;
  assign \new_[19090]_  = \new_[19089]_  & \new_[19086]_ ;
  assign \new_[19091]_  = \new_[19090]_  & \new_[19083]_ ;
  assign \new_[19095]_  = A199 & A166;
  assign \new_[19096]_  = A168 & \new_[19095]_ ;
  assign \new_[19100]_  = A203 & A201;
  assign \new_[19101]_  = ~A200 & \new_[19100]_ ;
  assign \new_[19102]_  = \new_[19101]_  & \new_[19096]_ ;
  assign \new_[19106]_  = A267 & ~A266;
  assign \new_[19107]_  = A265 & \new_[19106]_ ;
  assign \new_[19110]_  = A298 & A269;
  assign \new_[19113]_  = ~A302 & ~A301;
  assign \new_[19114]_  = \new_[19113]_  & \new_[19110]_ ;
  assign \new_[19115]_  = \new_[19114]_  & \new_[19107]_ ;
  assign \new_[19119]_  = A199 & A167;
  assign \new_[19120]_  = A168 & \new_[19119]_ ;
  assign \new_[19124]_  = A202 & A201;
  assign \new_[19125]_  = ~A200 & \new_[19124]_ ;
  assign \new_[19126]_  = \new_[19125]_  & \new_[19120]_ ;
  assign \new_[19130]_  = A267 & ~A266;
  assign \new_[19131]_  = A265 & \new_[19130]_ ;
  assign \new_[19134]_  = A298 & A268;
  assign \new_[19137]_  = ~A302 & ~A301;
  assign \new_[19138]_  = \new_[19137]_  & \new_[19134]_ ;
  assign \new_[19139]_  = \new_[19138]_  & \new_[19131]_ ;
  assign \new_[19143]_  = A199 & A167;
  assign \new_[19144]_  = A168 & \new_[19143]_ ;
  assign \new_[19148]_  = A202 & A201;
  assign \new_[19149]_  = ~A200 & \new_[19148]_ ;
  assign \new_[19150]_  = \new_[19149]_  & \new_[19144]_ ;
  assign \new_[19154]_  = A267 & ~A266;
  assign \new_[19155]_  = A265 & \new_[19154]_ ;
  assign \new_[19158]_  = A298 & A269;
  assign \new_[19161]_  = ~A302 & ~A301;
  assign \new_[19162]_  = \new_[19161]_  & \new_[19158]_ ;
  assign \new_[19163]_  = \new_[19162]_  & \new_[19155]_ ;
  assign \new_[19167]_  = A199 & A167;
  assign \new_[19168]_  = A168 & \new_[19167]_ ;
  assign \new_[19172]_  = A203 & A201;
  assign \new_[19173]_  = ~A200 & \new_[19172]_ ;
  assign \new_[19174]_  = \new_[19173]_  & \new_[19168]_ ;
  assign \new_[19178]_  = A267 & ~A266;
  assign \new_[19179]_  = A265 & \new_[19178]_ ;
  assign \new_[19182]_  = A298 & A268;
  assign \new_[19185]_  = ~A302 & ~A301;
  assign \new_[19186]_  = \new_[19185]_  & \new_[19182]_ ;
  assign \new_[19187]_  = \new_[19186]_  & \new_[19179]_ ;
  assign \new_[19191]_  = A199 & A167;
  assign \new_[19192]_  = A168 & \new_[19191]_ ;
  assign \new_[19196]_  = A203 & A201;
  assign \new_[19197]_  = ~A200 & \new_[19196]_ ;
  assign \new_[19198]_  = \new_[19197]_  & \new_[19192]_ ;
  assign \new_[19202]_  = A267 & ~A266;
  assign \new_[19203]_  = A265 & \new_[19202]_ ;
  assign \new_[19206]_  = A298 & A269;
  assign \new_[19209]_  = ~A302 & ~A301;
  assign \new_[19210]_  = \new_[19209]_  & \new_[19206]_ ;
  assign \new_[19211]_  = \new_[19210]_  & \new_[19203]_ ;
  assign \new_[19215]_  = ~A166 & ~A167;
  assign \new_[19216]_  = A170 & \new_[19215]_ ;
  assign \new_[19220]_  = ~A203 & ~A202;
  assign \new_[19221]_  = ~A200 & \new_[19220]_ ;
  assign \new_[19222]_  = \new_[19221]_  & \new_[19216]_ ;
  assign \new_[19226]_  = A267 & ~A266;
  assign \new_[19227]_  = A265 & \new_[19226]_ ;
  assign \new_[19230]_  = A298 & A268;
  assign \new_[19233]_  = ~A302 & ~A301;
  assign \new_[19234]_  = \new_[19233]_  & \new_[19230]_ ;
  assign \new_[19235]_  = \new_[19234]_  & \new_[19227]_ ;
  assign \new_[19239]_  = ~A166 & ~A167;
  assign \new_[19240]_  = A170 & \new_[19239]_ ;
  assign \new_[19244]_  = ~A203 & ~A202;
  assign \new_[19245]_  = ~A200 & \new_[19244]_ ;
  assign \new_[19246]_  = \new_[19245]_  & \new_[19240]_ ;
  assign \new_[19250]_  = A267 & ~A266;
  assign \new_[19251]_  = A265 & \new_[19250]_ ;
  assign \new_[19254]_  = A298 & A269;
  assign \new_[19257]_  = ~A302 & ~A301;
  assign \new_[19258]_  = \new_[19257]_  & \new_[19254]_ ;
  assign \new_[19259]_  = \new_[19258]_  & \new_[19251]_ ;
  assign \new_[19263]_  = ~A166 & ~A167;
  assign \new_[19264]_  = A170 & \new_[19263]_ ;
  assign \new_[19268]_  = A201 & ~A200;
  assign \new_[19269]_  = A199 & \new_[19268]_ ;
  assign \new_[19270]_  = \new_[19269]_  & \new_[19264]_ ;
  assign \new_[19274]_  = A266 & A265;
  assign \new_[19275]_  = A202 & \new_[19274]_ ;
  assign \new_[19278]_  = ~A299 & A298;
  assign \new_[19281]_  = A301 & A300;
  assign \new_[19282]_  = \new_[19281]_  & \new_[19278]_ ;
  assign \new_[19283]_  = \new_[19282]_  & \new_[19275]_ ;
  assign \new_[19287]_  = ~A166 & ~A167;
  assign \new_[19288]_  = A170 & \new_[19287]_ ;
  assign \new_[19292]_  = A201 & ~A200;
  assign \new_[19293]_  = A199 & \new_[19292]_ ;
  assign \new_[19294]_  = \new_[19293]_  & \new_[19288]_ ;
  assign \new_[19298]_  = A266 & A265;
  assign \new_[19299]_  = A202 & \new_[19298]_ ;
  assign \new_[19302]_  = ~A299 & A298;
  assign \new_[19305]_  = A302 & A300;
  assign \new_[19306]_  = \new_[19305]_  & \new_[19302]_ ;
  assign \new_[19307]_  = \new_[19306]_  & \new_[19299]_ ;
  assign \new_[19311]_  = ~A166 & ~A167;
  assign \new_[19312]_  = A170 & \new_[19311]_ ;
  assign \new_[19316]_  = A201 & ~A200;
  assign \new_[19317]_  = A199 & \new_[19316]_ ;
  assign \new_[19318]_  = \new_[19317]_  & \new_[19312]_ ;
  assign \new_[19322]_  = ~A267 & ~A266;
  assign \new_[19323]_  = A202 & \new_[19322]_ ;
  assign \new_[19326]_  = ~A299 & A298;
  assign \new_[19329]_  = A301 & A300;
  assign \new_[19330]_  = \new_[19329]_  & \new_[19326]_ ;
  assign \new_[19331]_  = \new_[19330]_  & \new_[19323]_ ;
  assign \new_[19335]_  = ~A166 & ~A167;
  assign \new_[19336]_  = A170 & \new_[19335]_ ;
  assign \new_[19340]_  = A201 & ~A200;
  assign \new_[19341]_  = A199 & \new_[19340]_ ;
  assign \new_[19342]_  = \new_[19341]_  & \new_[19336]_ ;
  assign \new_[19346]_  = ~A267 & ~A266;
  assign \new_[19347]_  = A202 & \new_[19346]_ ;
  assign \new_[19350]_  = ~A299 & A298;
  assign \new_[19353]_  = A302 & A300;
  assign \new_[19354]_  = \new_[19353]_  & \new_[19350]_ ;
  assign \new_[19355]_  = \new_[19354]_  & \new_[19347]_ ;
  assign \new_[19359]_  = ~A166 & ~A167;
  assign \new_[19360]_  = A170 & \new_[19359]_ ;
  assign \new_[19364]_  = A201 & ~A200;
  assign \new_[19365]_  = A199 & \new_[19364]_ ;
  assign \new_[19366]_  = \new_[19365]_  & \new_[19360]_ ;
  assign \new_[19370]_  = ~A266 & ~A265;
  assign \new_[19371]_  = A202 & \new_[19370]_ ;
  assign \new_[19374]_  = ~A299 & A298;
  assign \new_[19377]_  = A301 & A300;
  assign \new_[19378]_  = \new_[19377]_  & \new_[19374]_ ;
  assign \new_[19379]_  = \new_[19378]_  & \new_[19371]_ ;
  assign \new_[19383]_  = ~A166 & ~A167;
  assign \new_[19384]_  = A170 & \new_[19383]_ ;
  assign \new_[19388]_  = A201 & ~A200;
  assign \new_[19389]_  = A199 & \new_[19388]_ ;
  assign \new_[19390]_  = \new_[19389]_  & \new_[19384]_ ;
  assign \new_[19394]_  = ~A266 & ~A265;
  assign \new_[19395]_  = A202 & \new_[19394]_ ;
  assign \new_[19398]_  = ~A299 & A298;
  assign \new_[19401]_  = A302 & A300;
  assign \new_[19402]_  = \new_[19401]_  & \new_[19398]_ ;
  assign \new_[19403]_  = \new_[19402]_  & \new_[19395]_ ;
  assign \new_[19407]_  = ~A166 & ~A167;
  assign \new_[19408]_  = A170 & \new_[19407]_ ;
  assign \new_[19412]_  = A201 & ~A200;
  assign \new_[19413]_  = A199 & \new_[19412]_ ;
  assign \new_[19414]_  = \new_[19413]_  & \new_[19408]_ ;
  assign \new_[19418]_  = A266 & A265;
  assign \new_[19419]_  = A203 & \new_[19418]_ ;
  assign \new_[19422]_  = ~A299 & A298;
  assign \new_[19425]_  = A301 & A300;
  assign \new_[19426]_  = \new_[19425]_  & \new_[19422]_ ;
  assign \new_[19427]_  = \new_[19426]_  & \new_[19419]_ ;
  assign \new_[19431]_  = ~A166 & ~A167;
  assign \new_[19432]_  = A170 & \new_[19431]_ ;
  assign \new_[19436]_  = A201 & ~A200;
  assign \new_[19437]_  = A199 & \new_[19436]_ ;
  assign \new_[19438]_  = \new_[19437]_  & \new_[19432]_ ;
  assign \new_[19442]_  = A266 & A265;
  assign \new_[19443]_  = A203 & \new_[19442]_ ;
  assign \new_[19446]_  = ~A299 & A298;
  assign \new_[19449]_  = A302 & A300;
  assign \new_[19450]_  = \new_[19449]_  & \new_[19446]_ ;
  assign \new_[19451]_  = \new_[19450]_  & \new_[19443]_ ;
  assign \new_[19455]_  = ~A166 & ~A167;
  assign \new_[19456]_  = A170 & \new_[19455]_ ;
  assign \new_[19460]_  = A201 & ~A200;
  assign \new_[19461]_  = A199 & \new_[19460]_ ;
  assign \new_[19462]_  = \new_[19461]_  & \new_[19456]_ ;
  assign \new_[19466]_  = ~A267 & ~A266;
  assign \new_[19467]_  = A203 & \new_[19466]_ ;
  assign \new_[19470]_  = ~A299 & A298;
  assign \new_[19473]_  = A301 & A300;
  assign \new_[19474]_  = \new_[19473]_  & \new_[19470]_ ;
  assign \new_[19475]_  = \new_[19474]_  & \new_[19467]_ ;
  assign \new_[19479]_  = ~A166 & ~A167;
  assign \new_[19480]_  = A170 & \new_[19479]_ ;
  assign \new_[19484]_  = A201 & ~A200;
  assign \new_[19485]_  = A199 & \new_[19484]_ ;
  assign \new_[19486]_  = \new_[19485]_  & \new_[19480]_ ;
  assign \new_[19490]_  = ~A267 & ~A266;
  assign \new_[19491]_  = A203 & \new_[19490]_ ;
  assign \new_[19494]_  = ~A299 & A298;
  assign \new_[19497]_  = A302 & A300;
  assign \new_[19498]_  = \new_[19497]_  & \new_[19494]_ ;
  assign \new_[19499]_  = \new_[19498]_  & \new_[19491]_ ;
  assign \new_[19503]_  = ~A166 & ~A167;
  assign \new_[19504]_  = A170 & \new_[19503]_ ;
  assign \new_[19508]_  = A201 & ~A200;
  assign \new_[19509]_  = A199 & \new_[19508]_ ;
  assign \new_[19510]_  = \new_[19509]_  & \new_[19504]_ ;
  assign \new_[19514]_  = ~A266 & ~A265;
  assign \new_[19515]_  = A203 & \new_[19514]_ ;
  assign \new_[19518]_  = ~A299 & A298;
  assign \new_[19521]_  = A301 & A300;
  assign \new_[19522]_  = \new_[19521]_  & \new_[19518]_ ;
  assign \new_[19523]_  = \new_[19522]_  & \new_[19515]_ ;
  assign \new_[19527]_  = ~A166 & ~A167;
  assign \new_[19528]_  = A170 & \new_[19527]_ ;
  assign \new_[19532]_  = A201 & ~A200;
  assign \new_[19533]_  = A199 & \new_[19532]_ ;
  assign \new_[19534]_  = \new_[19533]_  & \new_[19528]_ ;
  assign \new_[19538]_  = ~A266 & ~A265;
  assign \new_[19539]_  = A203 & \new_[19538]_ ;
  assign \new_[19542]_  = ~A299 & A298;
  assign \new_[19545]_  = A302 & A300;
  assign \new_[19546]_  = \new_[19545]_  & \new_[19542]_ ;
  assign \new_[19547]_  = \new_[19546]_  & \new_[19539]_ ;
  assign \new_[19551]_  = A167 & ~A168;
  assign \new_[19552]_  = A169 & \new_[19551]_ ;
  assign \new_[19556]_  = A200 & A199;
  assign \new_[19557]_  = ~A166 & \new_[19556]_ ;
  assign \new_[19558]_  = \new_[19557]_  & \new_[19552]_ ;
  assign \new_[19562]_  = A267 & ~A266;
  assign \new_[19563]_  = A265 & \new_[19562]_ ;
  assign \new_[19566]_  = A298 & A268;
  assign \new_[19569]_  = ~A302 & ~A301;
  assign \new_[19570]_  = \new_[19569]_  & \new_[19566]_ ;
  assign \new_[19571]_  = \new_[19570]_  & \new_[19563]_ ;
  assign \new_[19575]_  = A167 & ~A168;
  assign \new_[19576]_  = A169 & \new_[19575]_ ;
  assign \new_[19580]_  = A200 & A199;
  assign \new_[19581]_  = ~A166 & \new_[19580]_ ;
  assign \new_[19582]_  = \new_[19581]_  & \new_[19576]_ ;
  assign \new_[19586]_  = A267 & ~A266;
  assign \new_[19587]_  = A265 & \new_[19586]_ ;
  assign \new_[19590]_  = A298 & A269;
  assign \new_[19593]_  = ~A302 & ~A301;
  assign \new_[19594]_  = \new_[19593]_  & \new_[19590]_ ;
  assign \new_[19595]_  = \new_[19594]_  & \new_[19587]_ ;
  assign \new_[19599]_  = A167 & ~A168;
  assign \new_[19600]_  = A169 & \new_[19599]_ ;
  assign \new_[19604]_  = A200 & ~A199;
  assign \new_[19605]_  = ~A166 & \new_[19604]_ ;
  assign \new_[19606]_  = \new_[19605]_  & \new_[19600]_ ;
  assign \new_[19610]_  = ~A269 & ~A268;
  assign \new_[19611]_  = ~A266 & \new_[19610]_ ;
  assign \new_[19614]_  = ~A299 & A298;
  assign \new_[19617]_  = A301 & A300;
  assign \new_[19618]_  = \new_[19617]_  & \new_[19614]_ ;
  assign \new_[19619]_  = \new_[19618]_  & \new_[19611]_ ;
  assign \new_[19623]_  = A167 & ~A168;
  assign \new_[19624]_  = A169 & \new_[19623]_ ;
  assign \new_[19628]_  = A200 & ~A199;
  assign \new_[19629]_  = ~A166 & \new_[19628]_ ;
  assign \new_[19630]_  = \new_[19629]_  & \new_[19624]_ ;
  assign \new_[19634]_  = ~A269 & ~A268;
  assign \new_[19635]_  = ~A266 & \new_[19634]_ ;
  assign \new_[19638]_  = ~A299 & A298;
  assign \new_[19641]_  = A302 & A300;
  assign \new_[19642]_  = \new_[19641]_  & \new_[19638]_ ;
  assign \new_[19643]_  = \new_[19642]_  & \new_[19635]_ ;
  assign \new_[19647]_  = A167 & ~A168;
  assign \new_[19648]_  = A169 & \new_[19647]_ ;
  assign \new_[19652]_  = ~A202 & ~A200;
  assign \new_[19653]_  = ~A166 & \new_[19652]_ ;
  assign \new_[19654]_  = \new_[19653]_  & \new_[19648]_ ;
  assign \new_[19658]_  = ~A266 & A265;
  assign \new_[19659]_  = ~A203 & \new_[19658]_ ;
  assign \new_[19662]_  = A268 & A267;
  assign \new_[19665]_  = ~A300 & A298;
  assign \new_[19666]_  = \new_[19665]_  & \new_[19662]_ ;
  assign \new_[19667]_  = \new_[19666]_  & \new_[19659]_ ;
  assign \new_[19671]_  = A167 & ~A168;
  assign \new_[19672]_  = A169 & \new_[19671]_ ;
  assign \new_[19676]_  = ~A202 & ~A200;
  assign \new_[19677]_  = ~A166 & \new_[19676]_ ;
  assign \new_[19678]_  = \new_[19677]_  & \new_[19672]_ ;
  assign \new_[19682]_  = ~A266 & A265;
  assign \new_[19683]_  = ~A203 & \new_[19682]_ ;
  assign \new_[19686]_  = A268 & A267;
  assign \new_[19689]_  = A299 & A298;
  assign \new_[19690]_  = \new_[19689]_  & \new_[19686]_ ;
  assign \new_[19691]_  = \new_[19690]_  & \new_[19683]_ ;
  assign \new_[19695]_  = A167 & ~A168;
  assign \new_[19696]_  = A169 & \new_[19695]_ ;
  assign \new_[19700]_  = ~A202 & ~A200;
  assign \new_[19701]_  = ~A166 & \new_[19700]_ ;
  assign \new_[19702]_  = \new_[19701]_  & \new_[19696]_ ;
  assign \new_[19706]_  = ~A266 & A265;
  assign \new_[19707]_  = ~A203 & \new_[19706]_ ;
  assign \new_[19710]_  = A268 & A267;
  assign \new_[19713]_  = ~A299 & ~A298;
  assign \new_[19714]_  = \new_[19713]_  & \new_[19710]_ ;
  assign \new_[19715]_  = \new_[19714]_  & \new_[19707]_ ;
  assign \new_[19719]_  = A167 & ~A168;
  assign \new_[19720]_  = A169 & \new_[19719]_ ;
  assign \new_[19724]_  = ~A202 & ~A200;
  assign \new_[19725]_  = ~A166 & \new_[19724]_ ;
  assign \new_[19726]_  = \new_[19725]_  & \new_[19720]_ ;
  assign \new_[19730]_  = ~A266 & A265;
  assign \new_[19731]_  = ~A203 & \new_[19730]_ ;
  assign \new_[19734]_  = A269 & A267;
  assign \new_[19737]_  = ~A300 & A298;
  assign \new_[19738]_  = \new_[19737]_  & \new_[19734]_ ;
  assign \new_[19739]_  = \new_[19738]_  & \new_[19731]_ ;
  assign \new_[19743]_  = A167 & ~A168;
  assign \new_[19744]_  = A169 & \new_[19743]_ ;
  assign \new_[19748]_  = ~A202 & ~A200;
  assign \new_[19749]_  = ~A166 & \new_[19748]_ ;
  assign \new_[19750]_  = \new_[19749]_  & \new_[19744]_ ;
  assign \new_[19754]_  = ~A266 & A265;
  assign \new_[19755]_  = ~A203 & \new_[19754]_ ;
  assign \new_[19758]_  = A269 & A267;
  assign \new_[19761]_  = A299 & A298;
  assign \new_[19762]_  = \new_[19761]_  & \new_[19758]_ ;
  assign \new_[19763]_  = \new_[19762]_  & \new_[19755]_ ;
  assign \new_[19767]_  = A167 & ~A168;
  assign \new_[19768]_  = A169 & \new_[19767]_ ;
  assign \new_[19772]_  = ~A202 & ~A200;
  assign \new_[19773]_  = ~A166 & \new_[19772]_ ;
  assign \new_[19774]_  = \new_[19773]_  & \new_[19768]_ ;
  assign \new_[19778]_  = ~A266 & A265;
  assign \new_[19779]_  = ~A203 & \new_[19778]_ ;
  assign \new_[19782]_  = A269 & A267;
  assign \new_[19785]_  = ~A299 & ~A298;
  assign \new_[19786]_  = \new_[19785]_  & \new_[19782]_ ;
  assign \new_[19787]_  = \new_[19786]_  & \new_[19779]_ ;
  assign \new_[19791]_  = A167 & ~A168;
  assign \new_[19792]_  = A169 & \new_[19791]_ ;
  assign \new_[19796]_  = ~A201 & ~A200;
  assign \new_[19797]_  = ~A166 & \new_[19796]_ ;
  assign \new_[19798]_  = \new_[19797]_  & \new_[19792]_ ;
  assign \new_[19802]_  = A267 & ~A266;
  assign \new_[19803]_  = A265 & \new_[19802]_ ;
  assign \new_[19806]_  = A298 & A268;
  assign \new_[19809]_  = ~A302 & ~A301;
  assign \new_[19810]_  = \new_[19809]_  & \new_[19806]_ ;
  assign \new_[19811]_  = \new_[19810]_  & \new_[19803]_ ;
  assign \new_[19815]_  = A167 & ~A168;
  assign \new_[19816]_  = A169 & \new_[19815]_ ;
  assign \new_[19820]_  = ~A201 & ~A200;
  assign \new_[19821]_  = ~A166 & \new_[19820]_ ;
  assign \new_[19822]_  = \new_[19821]_  & \new_[19816]_ ;
  assign \new_[19826]_  = A267 & ~A266;
  assign \new_[19827]_  = A265 & \new_[19826]_ ;
  assign \new_[19830]_  = A298 & A269;
  assign \new_[19833]_  = ~A302 & ~A301;
  assign \new_[19834]_  = \new_[19833]_  & \new_[19830]_ ;
  assign \new_[19835]_  = \new_[19834]_  & \new_[19827]_ ;
  assign \new_[19839]_  = A167 & ~A168;
  assign \new_[19840]_  = A169 & \new_[19839]_ ;
  assign \new_[19844]_  = ~A200 & A199;
  assign \new_[19845]_  = ~A166 & \new_[19844]_ ;
  assign \new_[19846]_  = \new_[19845]_  & \new_[19840]_ ;
  assign \new_[19850]_  = ~A266 & A202;
  assign \new_[19851]_  = A201 & \new_[19850]_ ;
  assign \new_[19854]_  = ~A269 & ~A268;
  assign \new_[19857]_  = A299 & ~A298;
  assign \new_[19858]_  = \new_[19857]_  & \new_[19854]_ ;
  assign \new_[19859]_  = \new_[19858]_  & \new_[19851]_ ;
  assign \new_[19863]_  = A167 & ~A168;
  assign \new_[19864]_  = A169 & \new_[19863]_ ;
  assign \new_[19868]_  = ~A200 & A199;
  assign \new_[19869]_  = ~A166 & \new_[19868]_ ;
  assign \new_[19870]_  = \new_[19869]_  & \new_[19864]_ ;
  assign \new_[19874]_  = ~A266 & A203;
  assign \new_[19875]_  = A201 & \new_[19874]_ ;
  assign \new_[19878]_  = ~A269 & ~A268;
  assign \new_[19881]_  = A299 & ~A298;
  assign \new_[19882]_  = \new_[19881]_  & \new_[19878]_ ;
  assign \new_[19883]_  = \new_[19882]_  & \new_[19875]_ ;
  assign \new_[19887]_  = A167 & ~A168;
  assign \new_[19888]_  = A169 & \new_[19887]_ ;
  assign \new_[19892]_  = ~A200 & ~A199;
  assign \new_[19893]_  = ~A166 & \new_[19892]_ ;
  assign \new_[19894]_  = \new_[19893]_  & \new_[19888]_ ;
  assign \new_[19898]_  = A267 & ~A266;
  assign \new_[19899]_  = A265 & \new_[19898]_ ;
  assign \new_[19902]_  = A298 & A268;
  assign \new_[19905]_  = ~A302 & ~A301;
  assign \new_[19906]_  = \new_[19905]_  & \new_[19902]_ ;
  assign \new_[19907]_  = \new_[19906]_  & \new_[19899]_ ;
  assign \new_[19911]_  = A167 & ~A168;
  assign \new_[19912]_  = A169 & \new_[19911]_ ;
  assign \new_[19916]_  = ~A200 & ~A199;
  assign \new_[19917]_  = ~A166 & \new_[19916]_ ;
  assign \new_[19918]_  = \new_[19917]_  & \new_[19912]_ ;
  assign \new_[19922]_  = A267 & ~A266;
  assign \new_[19923]_  = A265 & \new_[19922]_ ;
  assign \new_[19926]_  = A298 & A269;
  assign \new_[19929]_  = ~A302 & ~A301;
  assign \new_[19930]_  = \new_[19929]_  & \new_[19926]_ ;
  assign \new_[19931]_  = \new_[19930]_  & \new_[19923]_ ;
  assign \new_[19935]_  = ~A167 & ~A168;
  assign \new_[19936]_  = A169 & \new_[19935]_ ;
  assign \new_[19940]_  = A200 & A199;
  assign \new_[19941]_  = A166 & \new_[19940]_ ;
  assign \new_[19942]_  = \new_[19941]_  & \new_[19936]_ ;
  assign \new_[19946]_  = A267 & ~A266;
  assign \new_[19947]_  = A265 & \new_[19946]_ ;
  assign \new_[19950]_  = A298 & A268;
  assign \new_[19953]_  = ~A302 & ~A301;
  assign \new_[19954]_  = \new_[19953]_  & \new_[19950]_ ;
  assign \new_[19955]_  = \new_[19954]_  & \new_[19947]_ ;
  assign \new_[19959]_  = ~A167 & ~A168;
  assign \new_[19960]_  = A169 & \new_[19959]_ ;
  assign \new_[19964]_  = A200 & A199;
  assign \new_[19965]_  = A166 & \new_[19964]_ ;
  assign \new_[19966]_  = \new_[19965]_  & \new_[19960]_ ;
  assign \new_[19970]_  = A267 & ~A266;
  assign \new_[19971]_  = A265 & \new_[19970]_ ;
  assign \new_[19974]_  = A298 & A269;
  assign \new_[19977]_  = ~A302 & ~A301;
  assign \new_[19978]_  = \new_[19977]_  & \new_[19974]_ ;
  assign \new_[19979]_  = \new_[19978]_  & \new_[19971]_ ;
  assign \new_[19983]_  = ~A167 & ~A168;
  assign \new_[19984]_  = A169 & \new_[19983]_ ;
  assign \new_[19988]_  = A200 & ~A199;
  assign \new_[19989]_  = A166 & \new_[19988]_ ;
  assign \new_[19990]_  = \new_[19989]_  & \new_[19984]_ ;
  assign \new_[19994]_  = ~A269 & ~A268;
  assign \new_[19995]_  = ~A266 & \new_[19994]_ ;
  assign \new_[19998]_  = ~A299 & A298;
  assign \new_[20001]_  = A301 & A300;
  assign \new_[20002]_  = \new_[20001]_  & \new_[19998]_ ;
  assign \new_[20003]_  = \new_[20002]_  & \new_[19995]_ ;
  assign \new_[20007]_  = ~A167 & ~A168;
  assign \new_[20008]_  = A169 & \new_[20007]_ ;
  assign \new_[20012]_  = A200 & ~A199;
  assign \new_[20013]_  = A166 & \new_[20012]_ ;
  assign \new_[20014]_  = \new_[20013]_  & \new_[20008]_ ;
  assign \new_[20018]_  = ~A269 & ~A268;
  assign \new_[20019]_  = ~A266 & \new_[20018]_ ;
  assign \new_[20022]_  = ~A299 & A298;
  assign \new_[20025]_  = A302 & A300;
  assign \new_[20026]_  = \new_[20025]_  & \new_[20022]_ ;
  assign \new_[20027]_  = \new_[20026]_  & \new_[20019]_ ;
  assign \new_[20031]_  = ~A167 & ~A168;
  assign \new_[20032]_  = A169 & \new_[20031]_ ;
  assign \new_[20036]_  = ~A202 & ~A200;
  assign \new_[20037]_  = A166 & \new_[20036]_ ;
  assign \new_[20038]_  = \new_[20037]_  & \new_[20032]_ ;
  assign \new_[20042]_  = ~A266 & A265;
  assign \new_[20043]_  = ~A203 & \new_[20042]_ ;
  assign \new_[20046]_  = A268 & A267;
  assign \new_[20049]_  = ~A300 & A298;
  assign \new_[20050]_  = \new_[20049]_  & \new_[20046]_ ;
  assign \new_[20051]_  = \new_[20050]_  & \new_[20043]_ ;
  assign \new_[20055]_  = ~A167 & ~A168;
  assign \new_[20056]_  = A169 & \new_[20055]_ ;
  assign \new_[20060]_  = ~A202 & ~A200;
  assign \new_[20061]_  = A166 & \new_[20060]_ ;
  assign \new_[20062]_  = \new_[20061]_  & \new_[20056]_ ;
  assign \new_[20066]_  = ~A266 & A265;
  assign \new_[20067]_  = ~A203 & \new_[20066]_ ;
  assign \new_[20070]_  = A268 & A267;
  assign \new_[20073]_  = A299 & A298;
  assign \new_[20074]_  = \new_[20073]_  & \new_[20070]_ ;
  assign \new_[20075]_  = \new_[20074]_  & \new_[20067]_ ;
  assign \new_[20079]_  = ~A167 & ~A168;
  assign \new_[20080]_  = A169 & \new_[20079]_ ;
  assign \new_[20084]_  = ~A202 & ~A200;
  assign \new_[20085]_  = A166 & \new_[20084]_ ;
  assign \new_[20086]_  = \new_[20085]_  & \new_[20080]_ ;
  assign \new_[20090]_  = ~A266 & A265;
  assign \new_[20091]_  = ~A203 & \new_[20090]_ ;
  assign \new_[20094]_  = A268 & A267;
  assign \new_[20097]_  = ~A299 & ~A298;
  assign \new_[20098]_  = \new_[20097]_  & \new_[20094]_ ;
  assign \new_[20099]_  = \new_[20098]_  & \new_[20091]_ ;
  assign \new_[20103]_  = ~A167 & ~A168;
  assign \new_[20104]_  = A169 & \new_[20103]_ ;
  assign \new_[20108]_  = ~A202 & ~A200;
  assign \new_[20109]_  = A166 & \new_[20108]_ ;
  assign \new_[20110]_  = \new_[20109]_  & \new_[20104]_ ;
  assign \new_[20114]_  = ~A266 & A265;
  assign \new_[20115]_  = ~A203 & \new_[20114]_ ;
  assign \new_[20118]_  = A269 & A267;
  assign \new_[20121]_  = ~A300 & A298;
  assign \new_[20122]_  = \new_[20121]_  & \new_[20118]_ ;
  assign \new_[20123]_  = \new_[20122]_  & \new_[20115]_ ;
  assign \new_[20127]_  = ~A167 & ~A168;
  assign \new_[20128]_  = A169 & \new_[20127]_ ;
  assign \new_[20132]_  = ~A202 & ~A200;
  assign \new_[20133]_  = A166 & \new_[20132]_ ;
  assign \new_[20134]_  = \new_[20133]_  & \new_[20128]_ ;
  assign \new_[20138]_  = ~A266 & A265;
  assign \new_[20139]_  = ~A203 & \new_[20138]_ ;
  assign \new_[20142]_  = A269 & A267;
  assign \new_[20145]_  = A299 & A298;
  assign \new_[20146]_  = \new_[20145]_  & \new_[20142]_ ;
  assign \new_[20147]_  = \new_[20146]_  & \new_[20139]_ ;
  assign \new_[20151]_  = ~A167 & ~A168;
  assign \new_[20152]_  = A169 & \new_[20151]_ ;
  assign \new_[20156]_  = ~A202 & ~A200;
  assign \new_[20157]_  = A166 & \new_[20156]_ ;
  assign \new_[20158]_  = \new_[20157]_  & \new_[20152]_ ;
  assign \new_[20162]_  = ~A266 & A265;
  assign \new_[20163]_  = ~A203 & \new_[20162]_ ;
  assign \new_[20166]_  = A269 & A267;
  assign \new_[20169]_  = ~A299 & ~A298;
  assign \new_[20170]_  = \new_[20169]_  & \new_[20166]_ ;
  assign \new_[20171]_  = \new_[20170]_  & \new_[20163]_ ;
  assign \new_[20175]_  = ~A167 & ~A168;
  assign \new_[20176]_  = A169 & \new_[20175]_ ;
  assign \new_[20180]_  = ~A201 & ~A200;
  assign \new_[20181]_  = A166 & \new_[20180]_ ;
  assign \new_[20182]_  = \new_[20181]_  & \new_[20176]_ ;
  assign \new_[20186]_  = A267 & ~A266;
  assign \new_[20187]_  = A265 & \new_[20186]_ ;
  assign \new_[20190]_  = A298 & A268;
  assign \new_[20193]_  = ~A302 & ~A301;
  assign \new_[20194]_  = \new_[20193]_  & \new_[20190]_ ;
  assign \new_[20195]_  = \new_[20194]_  & \new_[20187]_ ;
  assign \new_[20199]_  = ~A167 & ~A168;
  assign \new_[20200]_  = A169 & \new_[20199]_ ;
  assign \new_[20204]_  = ~A201 & ~A200;
  assign \new_[20205]_  = A166 & \new_[20204]_ ;
  assign \new_[20206]_  = \new_[20205]_  & \new_[20200]_ ;
  assign \new_[20210]_  = A267 & ~A266;
  assign \new_[20211]_  = A265 & \new_[20210]_ ;
  assign \new_[20214]_  = A298 & A269;
  assign \new_[20217]_  = ~A302 & ~A301;
  assign \new_[20218]_  = \new_[20217]_  & \new_[20214]_ ;
  assign \new_[20219]_  = \new_[20218]_  & \new_[20211]_ ;
  assign \new_[20223]_  = ~A167 & ~A168;
  assign \new_[20224]_  = A169 & \new_[20223]_ ;
  assign \new_[20228]_  = ~A200 & A199;
  assign \new_[20229]_  = A166 & \new_[20228]_ ;
  assign \new_[20230]_  = \new_[20229]_  & \new_[20224]_ ;
  assign \new_[20234]_  = ~A266 & A202;
  assign \new_[20235]_  = A201 & \new_[20234]_ ;
  assign \new_[20238]_  = ~A269 & ~A268;
  assign \new_[20241]_  = A299 & ~A298;
  assign \new_[20242]_  = \new_[20241]_  & \new_[20238]_ ;
  assign \new_[20243]_  = \new_[20242]_  & \new_[20235]_ ;
  assign \new_[20247]_  = ~A167 & ~A168;
  assign \new_[20248]_  = A169 & \new_[20247]_ ;
  assign \new_[20252]_  = ~A200 & A199;
  assign \new_[20253]_  = A166 & \new_[20252]_ ;
  assign \new_[20254]_  = \new_[20253]_  & \new_[20248]_ ;
  assign \new_[20258]_  = ~A266 & A203;
  assign \new_[20259]_  = A201 & \new_[20258]_ ;
  assign \new_[20262]_  = ~A269 & ~A268;
  assign \new_[20265]_  = A299 & ~A298;
  assign \new_[20266]_  = \new_[20265]_  & \new_[20262]_ ;
  assign \new_[20267]_  = \new_[20266]_  & \new_[20259]_ ;
  assign \new_[20271]_  = ~A167 & ~A168;
  assign \new_[20272]_  = A169 & \new_[20271]_ ;
  assign \new_[20276]_  = ~A200 & ~A199;
  assign \new_[20277]_  = A166 & \new_[20276]_ ;
  assign \new_[20278]_  = \new_[20277]_  & \new_[20272]_ ;
  assign \new_[20282]_  = A267 & ~A266;
  assign \new_[20283]_  = A265 & \new_[20282]_ ;
  assign \new_[20286]_  = A298 & A268;
  assign \new_[20289]_  = ~A302 & ~A301;
  assign \new_[20290]_  = \new_[20289]_  & \new_[20286]_ ;
  assign \new_[20291]_  = \new_[20290]_  & \new_[20283]_ ;
  assign \new_[20295]_  = ~A167 & ~A168;
  assign \new_[20296]_  = A169 & \new_[20295]_ ;
  assign \new_[20300]_  = ~A200 & ~A199;
  assign \new_[20301]_  = A166 & \new_[20300]_ ;
  assign \new_[20302]_  = \new_[20301]_  & \new_[20296]_ ;
  assign \new_[20306]_  = A267 & ~A266;
  assign \new_[20307]_  = A265 & \new_[20306]_ ;
  assign \new_[20310]_  = A298 & A269;
  assign \new_[20313]_  = ~A302 & ~A301;
  assign \new_[20314]_  = \new_[20313]_  & \new_[20310]_ ;
  assign \new_[20315]_  = \new_[20314]_  & \new_[20307]_ ;
  assign \new_[20319]_  = ~A168 & A169;
  assign \new_[20320]_  = A170 & \new_[20319]_ ;
  assign \new_[20324]_  = ~A203 & ~A202;
  assign \new_[20325]_  = ~A200 & \new_[20324]_ ;
  assign \new_[20326]_  = \new_[20325]_  & \new_[20320]_ ;
  assign \new_[20330]_  = A267 & ~A266;
  assign \new_[20331]_  = A265 & \new_[20330]_ ;
  assign \new_[20334]_  = A298 & A268;
  assign \new_[20337]_  = ~A302 & ~A301;
  assign \new_[20338]_  = \new_[20337]_  & \new_[20334]_ ;
  assign \new_[20339]_  = \new_[20338]_  & \new_[20331]_ ;
  assign \new_[20343]_  = ~A168 & A169;
  assign \new_[20344]_  = A170 & \new_[20343]_ ;
  assign \new_[20348]_  = ~A203 & ~A202;
  assign \new_[20349]_  = ~A200 & \new_[20348]_ ;
  assign \new_[20350]_  = \new_[20349]_  & \new_[20344]_ ;
  assign \new_[20354]_  = A267 & ~A266;
  assign \new_[20355]_  = A265 & \new_[20354]_ ;
  assign \new_[20358]_  = A298 & A269;
  assign \new_[20361]_  = ~A302 & ~A301;
  assign \new_[20362]_  = \new_[20361]_  & \new_[20358]_ ;
  assign \new_[20363]_  = \new_[20362]_  & \new_[20355]_ ;
  assign \new_[20367]_  = ~A168 & A169;
  assign \new_[20368]_  = A170 & \new_[20367]_ ;
  assign \new_[20372]_  = A201 & ~A200;
  assign \new_[20373]_  = A199 & \new_[20372]_ ;
  assign \new_[20374]_  = \new_[20373]_  & \new_[20368]_ ;
  assign \new_[20378]_  = A266 & A265;
  assign \new_[20379]_  = A202 & \new_[20378]_ ;
  assign \new_[20382]_  = ~A299 & A298;
  assign \new_[20385]_  = A301 & A300;
  assign \new_[20386]_  = \new_[20385]_  & \new_[20382]_ ;
  assign \new_[20387]_  = \new_[20386]_  & \new_[20379]_ ;
  assign \new_[20391]_  = ~A168 & A169;
  assign \new_[20392]_  = A170 & \new_[20391]_ ;
  assign \new_[20396]_  = A201 & ~A200;
  assign \new_[20397]_  = A199 & \new_[20396]_ ;
  assign \new_[20398]_  = \new_[20397]_  & \new_[20392]_ ;
  assign \new_[20402]_  = A266 & A265;
  assign \new_[20403]_  = A202 & \new_[20402]_ ;
  assign \new_[20406]_  = ~A299 & A298;
  assign \new_[20409]_  = A302 & A300;
  assign \new_[20410]_  = \new_[20409]_  & \new_[20406]_ ;
  assign \new_[20411]_  = \new_[20410]_  & \new_[20403]_ ;
  assign \new_[20415]_  = ~A168 & A169;
  assign \new_[20416]_  = A170 & \new_[20415]_ ;
  assign \new_[20420]_  = A201 & ~A200;
  assign \new_[20421]_  = A199 & \new_[20420]_ ;
  assign \new_[20422]_  = \new_[20421]_  & \new_[20416]_ ;
  assign \new_[20426]_  = ~A267 & ~A266;
  assign \new_[20427]_  = A202 & \new_[20426]_ ;
  assign \new_[20430]_  = ~A299 & A298;
  assign \new_[20433]_  = A301 & A300;
  assign \new_[20434]_  = \new_[20433]_  & \new_[20430]_ ;
  assign \new_[20435]_  = \new_[20434]_  & \new_[20427]_ ;
  assign \new_[20439]_  = ~A168 & A169;
  assign \new_[20440]_  = A170 & \new_[20439]_ ;
  assign \new_[20444]_  = A201 & ~A200;
  assign \new_[20445]_  = A199 & \new_[20444]_ ;
  assign \new_[20446]_  = \new_[20445]_  & \new_[20440]_ ;
  assign \new_[20450]_  = ~A267 & ~A266;
  assign \new_[20451]_  = A202 & \new_[20450]_ ;
  assign \new_[20454]_  = ~A299 & A298;
  assign \new_[20457]_  = A302 & A300;
  assign \new_[20458]_  = \new_[20457]_  & \new_[20454]_ ;
  assign \new_[20459]_  = \new_[20458]_  & \new_[20451]_ ;
  assign \new_[20463]_  = ~A168 & A169;
  assign \new_[20464]_  = A170 & \new_[20463]_ ;
  assign \new_[20468]_  = A201 & ~A200;
  assign \new_[20469]_  = A199 & \new_[20468]_ ;
  assign \new_[20470]_  = \new_[20469]_  & \new_[20464]_ ;
  assign \new_[20474]_  = ~A266 & ~A265;
  assign \new_[20475]_  = A202 & \new_[20474]_ ;
  assign \new_[20478]_  = ~A299 & A298;
  assign \new_[20481]_  = A301 & A300;
  assign \new_[20482]_  = \new_[20481]_  & \new_[20478]_ ;
  assign \new_[20483]_  = \new_[20482]_  & \new_[20475]_ ;
  assign \new_[20487]_  = ~A168 & A169;
  assign \new_[20488]_  = A170 & \new_[20487]_ ;
  assign \new_[20492]_  = A201 & ~A200;
  assign \new_[20493]_  = A199 & \new_[20492]_ ;
  assign \new_[20494]_  = \new_[20493]_  & \new_[20488]_ ;
  assign \new_[20498]_  = ~A266 & ~A265;
  assign \new_[20499]_  = A202 & \new_[20498]_ ;
  assign \new_[20502]_  = ~A299 & A298;
  assign \new_[20505]_  = A302 & A300;
  assign \new_[20506]_  = \new_[20505]_  & \new_[20502]_ ;
  assign \new_[20507]_  = \new_[20506]_  & \new_[20499]_ ;
  assign \new_[20511]_  = ~A168 & A169;
  assign \new_[20512]_  = A170 & \new_[20511]_ ;
  assign \new_[20516]_  = A201 & ~A200;
  assign \new_[20517]_  = A199 & \new_[20516]_ ;
  assign \new_[20518]_  = \new_[20517]_  & \new_[20512]_ ;
  assign \new_[20522]_  = A266 & A265;
  assign \new_[20523]_  = A203 & \new_[20522]_ ;
  assign \new_[20526]_  = ~A299 & A298;
  assign \new_[20529]_  = A301 & A300;
  assign \new_[20530]_  = \new_[20529]_  & \new_[20526]_ ;
  assign \new_[20531]_  = \new_[20530]_  & \new_[20523]_ ;
  assign \new_[20535]_  = ~A168 & A169;
  assign \new_[20536]_  = A170 & \new_[20535]_ ;
  assign \new_[20540]_  = A201 & ~A200;
  assign \new_[20541]_  = A199 & \new_[20540]_ ;
  assign \new_[20542]_  = \new_[20541]_  & \new_[20536]_ ;
  assign \new_[20546]_  = A266 & A265;
  assign \new_[20547]_  = A203 & \new_[20546]_ ;
  assign \new_[20550]_  = ~A299 & A298;
  assign \new_[20553]_  = A302 & A300;
  assign \new_[20554]_  = \new_[20553]_  & \new_[20550]_ ;
  assign \new_[20555]_  = \new_[20554]_  & \new_[20547]_ ;
  assign \new_[20559]_  = ~A168 & A169;
  assign \new_[20560]_  = A170 & \new_[20559]_ ;
  assign \new_[20564]_  = A201 & ~A200;
  assign \new_[20565]_  = A199 & \new_[20564]_ ;
  assign \new_[20566]_  = \new_[20565]_  & \new_[20560]_ ;
  assign \new_[20570]_  = ~A267 & ~A266;
  assign \new_[20571]_  = A203 & \new_[20570]_ ;
  assign \new_[20574]_  = ~A299 & A298;
  assign \new_[20577]_  = A301 & A300;
  assign \new_[20578]_  = \new_[20577]_  & \new_[20574]_ ;
  assign \new_[20579]_  = \new_[20578]_  & \new_[20571]_ ;
  assign \new_[20583]_  = ~A168 & A169;
  assign \new_[20584]_  = A170 & \new_[20583]_ ;
  assign \new_[20588]_  = A201 & ~A200;
  assign \new_[20589]_  = A199 & \new_[20588]_ ;
  assign \new_[20590]_  = \new_[20589]_  & \new_[20584]_ ;
  assign \new_[20594]_  = ~A267 & ~A266;
  assign \new_[20595]_  = A203 & \new_[20594]_ ;
  assign \new_[20598]_  = ~A299 & A298;
  assign \new_[20601]_  = A302 & A300;
  assign \new_[20602]_  = \new_[20601]_  & \new_[20598]_ ;
  assign \new_[20603]_  = \new_[20602]_  & \new_[20595]_ ;
  assign \new_[20607]_  = ~A168 & A169;
  assign \new_[20608]_  = A170 & \new_[20607]_ ;
  assign \new_[20612]_  = A201 & ~A200;
  assign \new_[20613]_  = A199 & \new_[20612]_ ;
  assign \new_[20614]_  = \new_[20613]_  & \new_[20608]_ ;
  assign \new_[20618]_  = ~A266 & ~A265;
  assign \new_[20619]_  = A203 & \new_[20618]_ ;
  assign \new_[20622]_  = ~A299 & A298;
  assign \new_[20625]_  = A301 & A300;
  assign \new_[20626]_  = \new_[20625]_  & \new_[20622]_ ;
  assign \new_[20627]_  = \new_[20626]_  & \new_[20619]_ ;
  assign \new_[20631]_  = ~A168 & A169;
  assign \new_[20632]_  = A170 & \new_[20631]_ ;
  assign \new_[20636]_  = A201 & ~A200;
  assign \new_[20637]_  = A199 & \new_[20636]_ ;
  assign \new_[20638]_  = \new_[20637]_  & \new_[20632]_ ;
  assign \new_[20642]_  = ~A266 & ~A265;
  assign \new_[20643]_  = A203 & \new_[20642]_ ;
  assign \new_[20646]_  = ~A299 & A298;
  assign \new_[20649]_  = A302 & A300;
  assign \new_[20650]_  = \new_[20649]_  & \new_[20646]_ ;
  assign \new_[20651]_  = \new_[20650]_  & \new_[20643]_ ;
  assign \new_[20655]_  = A167 & A169;
  assign \new_[20656]_  = ~A170 & \new_[20655]_ ;
  assign \new_[20660]_  = A200 & A199;
  assign \new_[20661]_  = A166 & \new_[20660]_ ;
  assign \new_[20662]_  = \new_[20661]_  & \new_[20656]_ ;
  assign \new_[20666]_  = ~A269 & ~A268;
  assign \new_[20667]_  = ~A266 & \new_[20666]_ ;
  assign \new_[20670]_  = ~A299 & A298;
  assign \new_[20673]_  = A301 & A300;
  assign \new_[20674]_  = \new_[20673]_  & \new_[20670]_ ;
  assign \new_[20675]_  = \new_[20674]_  & \new_[20667]_ ;
  assign \new_[20679]_  = A167 & A169;
  assign \new_[20680]_  = ~A170 & \new_[20679]_ ;
  assign \new_[20684]_  = A200 & A199;
  assign \new_[20685]_  = A166 & \new_[20684]_ ;
  assign \new_[20686]_  = \new_[20685]_  & \new_[20680]_ ;
  assign \new_[20690]_  = ~A269 & ~A268;
  assign \new_[20691]_  = ~A266 & \new_[20690]_ ;
  assign \new_[20694]_  = ~A299 & A298;
  assign \new_[20697]_  = A302 & A300;
  assign \new_[20698]_  = \new_[20697]_  & \new_[20694]_ ;
  assign \new_[20699]_  = \new_[20698]_  & \new_[20691]_ ;
  assign \new_[20703]_  = A167 & A169;
  assign \new_[20704]_  = ~A170 & \new_[20703]_ ;
  assign \new_[20708]_  = A200 & ~A199;
  assign \new_[20709]_  = A166 & \new_[20708]_ ;
  assign \new_[20710]_  = \new_[20709]_  & \new_[20704]_ ;
  assign \new_[20714]_  = A267 & ~A266;
  assign \new_[20715]_  = A265 & \new_[20714]_ ;
  assign \new_[20718]_  = A298 & A268;
  assign \new_[20721]_  = ~A302 & ~A301;
  assign \new_[20722]_  = \new_[20721]_  & \new_[20718]_ ;
  assign \new_[20723]_  = \new_[20722]_  & \new_[20715]_ ;
  assign \new_[20727]_  = A167 & A169;
  assign \new_[20728]_  = ~A170 & \new_[20727]_ ;
  assign \new_[20732]_  = A200 & ~A199;
  assign \new_[20733]_  = A166 & \new_[20732]_ ;
  assign \new_[20734]_  = \new_[20733]_  & \new_[20728]_ ;
  assign \new_[20738]_  = A267 & ~A266;
  assign \new_[20739]_  = A265 & \new_[20738]_ ;
  assign \new_[20742]_  = A298 & A269;
  assign \new_[20745]_  = ~A302 & ~A301;
  assign \new_[20746]_  = \new_[20745]_  & \new_[20742]_ ;
  assign \new_[20747]_  = \new_[20746]_  & \new_[20739]_ ;
  assign \new_[20751]_  = A167 & A169;
  assign \new_[20752]_  = ~A170 & \new_[20751]_ ;
  assign \new_[20756]_  = ~A202 & ~A200;
  assign \new_[20757]_  = A166 & \new_[20756]_ ;
  assign \new_[20758]_  = \new_[20757]_  & \new_[20752]_ ;
  assign \new_[20762]_  = A266 & A265;
  assign \new_[20763]_  = ~A203 & \new_[20762]_ ;
  assign \new_[20766]_  = ~A299 & A298;
  assign \new_[20769]_  = A301 & A300;
  assign \new_[20770]_  = \new_[20769]_  & \new_[20766]_ ;
  assign \new_[20771]_  = \new_[20770]_  & \new_[20763]_ ;
  assign \new_[20775]_  = A167 & A169;
  assign \new_[20776]_  = ~A170 & \new_[20775]_ ;
  assign \new_[20780]_  = ~A202 & ~A200;
  assign \new_[20781]_  = A166 & \new_[20780]_ ;
  assign \new_[20782]_  = \new_[20781]_  & \new_[20776]_ ;
  assign \new_[20786]_  = A266 & A265;
  assign \new_[20787]_  = ~A203 & \new_[20786]_ ;
  assign \new_[20790]_  = ~A299 & A298;
  assign \new_[20793]_  = A302 & A300;
  assign \new_[20794]_  = \new_[20793]_  & \new_[20790]_ ;
  assign \new_[20795]_  = \new_[20794]_  & \new_[20787]_ ;
  assign \new_[20799]_  = A167 & A169;
  assign \new_[20800]_  = ~A170 & \new_[20799]_ ;
  assign \new_[20804]_  = ~A202 & ~A200;
  assign \new_[20805]_  = A166 & \new_[20804]_ ;
  assign \new_[20806]_  = \new_[20805]_  & \new_[20800]_ ;
  assign \new_[20810]_  = ~A267 & ~A266;
  assign \new_[20811]_  = ~A203 & \new_[20810]_ ;
  assign \new_[20814]_  = ~A299 & A298;
  assign \new_[20817]_  = A301 & A300;
  assign \new_[20818]_  = \new_[20817]_  & \new_[20814]_ ;
  assign \new_[20819]_  = \new_[20818]_  & \new_[20811]_ ;
  assign \new_[20823]_  = A167 & A169;
  assign \new_[20824]_  = ~A170 & \new_[20823]_ ;
  assign \new_[20828]_  = ~A202 & ~A200;
  assign \new_[20829]_  = A166 & \new_[20828]_ ;
  assign \new_[20830]_  = \new_[20829]_  & \new_[20824]_ ;
  assign \new_[20834]_  = ~A267 & ~A266;
  assign \new_[20835]_  = ~A203 & \new_[20834]_ ;
  assign \new_[20838]_  = ~A299 & A298;
  assign \new_[20841]_  = A302 & A300;
  assign \new_[20842]_  = \new_[20841]_  & \new_[20838]_ ;
  assign \new_[20843]_  = \new_[20842]_  & \new_[20835]_ ;
  assign \new_[20847]_  = A167 & A169;
  assign \new_[20848]_  = ~A170 & \new_[20847]_ ;
  assign \new_[20852]_  = ~A202 & ~A200;
  assign \new_[20853]_  = A166 & \new_[20852]_ ;
  assign \new_[20854]_  = \new_[20853]_  & \new_[20848]_ ;
  assign \new_[20858]_  = ~A266 & ~A265;
  assign \new_[20859]_  = ~A203 & \new_[20858]_ ;
  assign \new_[20862]_  = ~A299 & A298;
  assign \new_[20865]_  = A301 & A300;
  assign \new_[20866]_  = \new_[20865]_  & \new_[20862]_ ;
  assign \new_[20867]_  = \new_[20866]_  & \new_[20859]_ ;
  assign \new_[20871]_  = A167 & A169;
  assign \new_[20872]_  = ~A170 & \new_[20871]_ ;
  assign \new_[20876]_  = ~A202 & ~A200;
  assign \new_[20877]_  = A166 & \new_[20876]_ ;
  assign \new_[20878]_  = \new_[20877]_  & \new_[20872]_ ;
  assign \new_[20882]_  = ~A266 & ~A265;
  assign \new_[20883]_  = ~A203 & \new_[20882]_ ;
  assign \new_[20886]_  = ~A299 & A298;
  assign \new_[20889]_  = A302 & A300;
  assign \new_[20890]_  = \new_[20889]_  & \new_[20886]_ ;
  assign \new_[20891]_  = \new_[20890]_  & \new_[20883]_ ;
  assign \new_[20895]_  = A167 & A169;
  assign \new_[20896]_  = ~A170 & \new_[20895]_ ;
  assign \new_[20900]_  = ~A201 & ~A200;
  assign \new_[20901]_  = A166 & \new_[20900]_ ;
  assign \new_[20902]_  = \new_[20901]_  & \new_[20896]_ ;
  assign \new_[20906]_  = ~A269 & ~A268;
  assign \new_[20907]_  = ~A266 & \new_[20906]_ ;
  assign \new_[20910]_  = ~A299 & A298;
  assign \new_[20913]_  = A301 & A300;
  assign \new_[20914]_  = \new_[20913]_  & \new_[20910]_ ;
  assign \new_[20915]_  = \new_[20914]_  & \new_[20907]_ ;
  assign \new_[20919]_  = A167 & A169;
  assign \new_[20920]_  = ~A170 & \new_[20919]_ ;
  assign \new_[20924]_  = ~A201 & ~A200;
  assign \new_[20925]_  = A166 & \new_[20924]_ ;
  assign \new_[20926]_  = \new_[20925]_  & \new_[20920]_ ;
  assign \new_[20930]_  = ~A269 & ~A268;
  assign \new_[20931]_  = ~A266 & \new_[20930]_ ;
  assign \new_[20934]_  = ~A299 & A298;
  assign \new_[20937]_  = A302 & A300;
  assign \new_[20938]_  = \new_[20937]_  & \new_[20934]_ ;
  assign \new_[20939]_  = \new_[20938]_  & \new_[20931]_ ;
  assign \new_[20943]_  = A167 & A169;
  assign \new_[20944]_  = ~A170 & \new_[20943]_ ;
  assign \new_[20948]_  = ~A200 & A199;
  assign \new_[20949]_  = A166 & \new_[20948]_ ;
  assign \new_[20950]_  = \new_[20949]_  & \new_[20944]_ ;
  assign \new_[20954]_  = ~A265 & A202;
  assign \new_[20955]_  = A201 & \new_[20954]_ ;
  assign \new_[20958]_  = A298 & A266;
  assign \new_[20961]_  = ~A302 & ~A301;
  assign \new_[20962]_  = \new_[20961]_  & \new_[20958]_ ;
  assign \new_[20963]_  = \new_[20962]_  & \new_[20955]_ ;
  assign \new_[20967]_  = A167 & A169;
  assign \new_[20968]_  = ~A170 & \new_[20967]_ ;
  assign \new_[20972]_  = ~A200 & A199;
  assign \new_[20973]_  = A166 & \new_[20972]_ ;
  assign \new_[20974]_  = \new_[20973]_  & \new_[20968]_ ;
  assign \new_[20978]_  = ~A265 & A203;
  assign \new_[20979]_  = A201 & \new_[20978]_ ;
  assign \new_[20982]_  = A298 & A266;
  assign \new_[20985]_  = ~A302 & ~A301;
  assign \new_[20986]_  = \new_[20985]_  & \new_[20982]_ ;
  assign \new_[20987]_  = \new_[20986]_  & \new_[20979]_ ;
  assign \new_[20991]_  = A167 & A169;
  assign \new_[20992]_  = ~A170 & \new_[20991]_ ;
  assign \new_[20996]_  = ~A200 & ~A199;
  assign \new_[20997]_  = A166 & \new_[20996]_ ;
  assign \new_[20998]_  = \new_[20997]_  & \new_[20992]_ ;
  assign \new_[21002]_  = ~A269 & ~A268;
  assign \new_[21003]_  = ~A266 & \new_[21002]_ ;
  assign \new_[21006]_  = ~A299 & A298;
  assign \new_[21009]_  = A301 & A300;
  assign \new_[21010]_  = \new_[21009]_  & \new_[21006]_ ;
  assign \new_[21011]_  = \new_[21010]_  & \new_[21003]_ ;
  assign \new_[21015]_  = A167 & A169;
  assign \new_[21016]_  = ~A170 & \new_[21015]_ ;
  assign \new_[21020]_  = ~A200 & ~A199;
  assign \new_[21021]_  = A166 & \new_[21020]_ ;
  assign \new_[21022]_  = \new_[21021]_  & \new_[21016]_ ;
  assign \new_[21026]_  = ~A269 & ~A268;
  assign \new_[21027]_  = ~A266 & \new_[21026]_ ;
  assign \new_[21030]_  = ~A299 & A298;
  assign \new_[21033]_  = A302 & A300;
  assign \new_[21034]_  = \new_[21033]_  & \new_[21030]_ ;
  assign \new_[21035]_  = \new_[21034]_  & \new_[21027]_ ;
  assign \new_[21039]_  = ~A167 & A169;
  assign \new_[21040]_  = ~A170 & \new_[21039]_ ;
  assign \new_[21044]_  = A200 & A199;
  assign \new_[21045]_  = ~A166 & \new_[21044]_ ;
  assign \new_[21046]_  = \new_[21045]_  & \new_[21040]_ ;
  assign \new_[21050]_  = ~A269 & ~A268;
  assign \new_[21051]_  = ~A266 & \new_[21050]_ ;
  assign \new_[21054]_  = ~A299 & A298;
  assign \new_[21057]_  = A301 & A300;
  assign \new_[21058]_  = \new_[21057]_  & \new_[21054]_ ;
  assign \new_[21059]_  = \new_[21058]_  & \new_[21051]_ ;
  assign \new_[21063]_  = ~A167 & A169;
  assign \new_[21064]_  = ~A170 & \new_[21063]_ ;
  assign \new_[21068]_  = A200 & A199;
  assign \new_[21069]_  = ~A166 & \new_[21068]_ ;
  assign \new_[21070]_  = \new_[21069]_  & \new_[21064]_ ;
  assign \new_[21074]_  = ~A269 & ~A268;
  assign \new_[21075]_  = ~A266 & \new_[21074]_ ;
  assign \new_[21078]_  = ~A299 & A298;
  assign \new_[21081]_  = A302 & A300;
  assign \new_[21082]_  = \new_[21081]_  & \new_[21078]_ ;
  assign \new_[21083]_  = \new_[21082]_  & \new_[21075]_ ;
  assign \new_[21087]_  = ~A167 & A169;
  assign \new_[21088]_  = ~A170 & \new_[21087]_ ;
  assign \new_[21092]_  = A200 & ~A199;
  assign \new_[21093]_  = ~A166 & \new_[21092]_ ;
  assign \new_[21094]_  = \new_[21093]_  & \new_[21088]_ ;
  assign \new_[21098]_  = A267 & ~A266;
  assign \new_[21099]_  = A265 & \new_[21098]_ ;
  assign \new_[21102]_  = A298 & A268;
  assign \new_[21105]_  = ~A302 & ~A301;
  assign \new_[21106]_  = \new_[21105]_  & \new_[21102]_ ;
  assign \new_[21107]_  = \new_[21106]_  & \new_[21099]_ ;
  assign \new_[21111]_  = ~A167 & A169;
  assign \new_[21112]_  = ~A170 & \new_[21111]_ ;
  assign \new_[21116]_  = A200 & ~A199;
  assign \new_[21117]_  = ~A166 & \new_[21116]_ ;
  assign \new_[21118]_  = \new_[21117]_  & \new_[21112]_ ;
  assign \new_[21122]_  = A267 & ~A266;
  assign \new_[21123]_  = A265 & \new_[21122]_ ;
  assign \new_[21126]_  = A298 & A269;
  assign \new_[21129]_  = ~A302 & ~A301;
  assign \new_[21130]_  = \new_[21129]_  & \new_[21126]_ ;
  assign \new_[21131]_  = \new_[21130]_  & \new_[21123]_ ;
  assign \new_[21135]_  = ~A167 & A169;
  assign \new_[21136]_  = ~A170 & \new_[21135]_ ;
  assign \new_[21140]_  = ~A202 & ~A200;
  assign \new_[21141]_  = ~A166 & \new_[21140]_ ;
  assign \new_[21142]_  = \new_[21141]_  & \new_[21136]_ ;
  assign \new_[21146]_  = A266 & A265;
  assign \new_[21147]_  = ~A203 & \new_[21146]_ ;
  assign \new_[21150]_  = ~A299 & A298;
  assign \new_[21153]_  = A301 & A300;
  assign \new_[21154]_  = \new_[21153]_  & \new_[21150]_ ;
  assign \new_[21155]_  = \new_[21154]_  & \new_[21147]_ ;
  assign \new_[21159]_  = ~A167 & A169;
  assign \new_[21160]_  = ~A170 & \new_[21159]_ ;
  assign \new_[21164]_  = ~A202 & ~A200;
  assign \new_[21165]_  = ~A166 & \new_[21164]_ ;
  assign \new_[21166]_  = \new_[21165]_  & \new_[21160]_ ;
  assign \new_[21170]_  = A266 & A265;
  assign \new_[21171]_  = ~A203 & \new_[21170]_ ;
  assign \new_[21174]_  = ~A299 & A298;
  assign \new_[21177]_  = A302 & A300;
  assign \new_[21178]_  = \new_[21177]_  & \new_[21174]_ ;
  assign \new_[21179]_  = \new_[21178]_  & \new_[21171]_ ;
  assign \new_[21183]_  = ~A167 & A169;
  assign \new_[21184]_  = ~A170 & \new_[21183]_ ;
  assign \new_[21188]_  = ~A202 & ~A200;
  assign \new_[21189]_  = ~A166 & \new_[21188]_ ;
  assign \new_[21190]_  = \new_[21189]_  & \new_[21184]_ ;
  assign \new_[21194]_  = ~A267 & ~A266;
  assign \new_[21195]_  = ~A203 & \new_[21194]_ ;
  assign \new_[21198]_  = ~A299 & A298;
  assign \new_[21201]_  = A301 & A300;
  assign \new_[21202]_  = \new_[21201]_  & \new_[21198]_ ;
  assign \new_[21203]_  = \new_[21202]_  & \new_[21195]_ ;
  assign \new_[21207]_  = ~A167 & A169;
  assign \new_[21208]_  = ~A170 & \new_[21207]_ ;
  assign \new_[21212]_  = ~A202 & ~A200;
  assign \new_[21213]_  = ~A166 & \new_[21212]_ ;
  assign \new_[21214]_  = \new_[21213]_  & \new_[21208]_ ;
  assign \new_[21218]_  = ~A267 & ~A266;
  assign \new_[21219]_  = ~A203 & \new_[21218]_ ;
  assign \new_[21222]_  = ~A299 & A298;
  assign \new_[21225]_  = A302 & A300;
  assign \new_[21226]_  = \new_[21225]_  & \new_[21222]_ ;
  assign \new_[21227]_  = \new_[21226]_  & \new_[21219]_ ;
  assign \new_[21231]_  = ~A167 & A169;
  assign \new_[21232]_  = ~A170 & \new_[21231]_ ;
  assign \new_[21236]_  = ~A202 & ~A200;
  assign \new_[21237]_  = ~A166 & \new_[21236]_ ;
  assign \new_[21238]_  = \new_[21237]_  & \new_[21232]_ ;
  assign \new_[21242]_  = ~A266 & ~A265;
  assign \new_[21243]_  = ~A203 & \new_[21242]_ ;
  assign \new_[21246]_  = ~A299 & A298;
  assign \new_[21249]_  = A301 & A300;
  assign \new_[21250]_  = \new_[21249]_  & \new_[21246]_ ;
  assign \new_[21251]_  = \new_[21250]_  & \new_[21243]_ ;
  assign \new_[21255]_  = ~A167 & A169;
  assign \new_[21256]_  = ~A170 & \new_[21255]_ ;
  assign \new_[21260]_  = ~A202 & ~A200;
  assign \new_[21261]_  = ~A166 & \new_[21260]_ ;
  assign \new_[21262]_  = \new_[21261]_  & \new_[21256]_ ;
  assign \new_[21266]_  = ~A266 & ~A265;
  assign \new_[21267]_  = ~A203 & \new_[21266]_ ;
  assign \new_[21270]_  = ~A299 & A298;
  assign \new_[21273]_  = A302 & A300;
  assign \new_[21274]_  = \new_[21273]_  & \new_[21270]_ ;
  assign \new_[21275]_  = \new_[21274]_  & \new_[21267]_ ;
  assign \new_[21279]_  = ~A167 & A169;
  assign \new_[21280]_  = ~A170 & \new_[21279]_ ;
  assign \new_[21284]_  = ~A201 & ~A200;
  assign \new_[21285]_  = ~A166 & \new_[21284]_ ;
  assign \new_[21286]_  = \new_[21285]_  & \new_[21280]_ ;
  assign \new_[21290]_  = ~A269 & ~A268;
  assign \new_[21291]_  = ~A266 & \new_[21290]_ ;
  assign \new_[21294]_  = ~A299 & A298;
  assign \new_[21297]_  = A301 & A300;
  assign \new_[21298]_  = \new_[21297]_  & \new_[21294]_ ;
  assign \new_[21299]_  = \new_[21298]_  & \new_[21291]_ ;
  assign \new_[21303]_  = ~A167 & A169;
  assign \new_[21304]_  = ~A170 & \new_[21303]_ ;
  assign \new_[21308]_  = ~A201 & ~A200;
  assign \new_[21309]_  = ~A166 & \new_[21308]_ ;
  assign \new_[21310]_  = \new_[21309]_  & \new_[21304]_ ;
  assign \new_[21314]_  = ~A269 & ~A268;
  assign \new_[21315]_  = ~A266 & \new_[21314]_ ;
  assign \new_[21318]_  = ~A299 & A298;
  assign \new_[21321]_  = A302 & A300;
  assign \new_[21322]_  = \new_[21321]_  & \new_[21318]_ ;
  assign \new_[21323]_  = \new_[21322]_  & \new_[21315]_ ;
  assign \new_[21327]_  = ~A167 & A169;
  assign \new_[21328]_  = ~A170 & \new_[21327]_ ;
  assign \new_[21332]_  = ~A200 & A199;
  assign \new_[21333]_  = ~A166 & \new_[21332]_ ;
  assign \new_[21334]_  = \new_[21333]_  & \new_[21328]_ ;
  assign \new_[21338]_  = ~A265 & A202;
  assign \new_[21339]_  = A201 & \new_[21338]_ ;
  assign \new_[21342]_  = A298 & A266;
  assign \new_[21345]_  = ~A302 & ~A301;
  assign \new_[21346]_  = \new_[21345]_  & \new_[21342]_ ;
  assign \new_[21347]_  = \new_[21346]_  & \new_[21339]_ ;
  assign \new_[21351]_  = ~A167 & A169;
  assign \new_[21352]_  = ~A170 & \new_[21351]_ ;
  assign \new_[21356]_  = ~A200 & A199;
  assign \new_[21357]_  = ~A166 & \new_[21356]_ ;
  assign \new_[21358]_  = \new_[21357]_  & \new_[21352]_ ;
  assign \new_[21362]_  = ~A265 & A203;
  assign \new_[21363]_  = A201 & \new_[21362]_ ;
  assign \new_[21366]_  = A298 & A266;
  assign \new_[21369]_  = ~A302 & ~A301;
  assign \new_[21370]_  = \new_[21369]_  & \new_[21366]_ ;
  assign \new_[21371]_  = \new_[21370]_  & \new_[21363]_ ;
  assign \new_[21375]_  = ~A167 & A169;
  assign \new_[21376]_  = ~A170 & \new_[21375]_ ;
  assign \new_[21380]_  = ~A200 & ~A199;
  assign \new_[21381]_  = ~A166 & \new_[21380]_ ;
  assign \new_[21382]_  = \new_[21381]_  & \new_[21376]_ ;
  assign \new_[21386]_  = ~A269 & ~A268;
  assign \new_[21387]_  = ~A266 & \new_[21386]_ ;
  assign \new_[21390]_  = ~A299 & A298;
  assign \new_[21393]_  = A301 & A300;
  assign \new_[21394]_  = \new_[21393]_  & \new_[21390]_ ;
  assign \new_[21395]_  = \new_[21394]_  & \new_[21387]_ ;
  assign \new_[21399]_  = ~A167 & A169;
  assign \new_[21400]_  = ~A170 & \new_[21399]_ ;
  assign \new_[21404]_  = ~A200 & ~A199;
  assign \new_[21405]_  = ~A166 & \new_[21404]_ ;
  assign \new_[21406]_  = \new_[21405]_  & \new_[21400]_ ;
  assign \new_[21410]_  = ~A269 & ~A268;
  assign \new_[21411]_  = ~A266 & \new_[21410]_ ;
  assign \new_[21414]_  = ~A299 & A298;
  assign \new_[21417]_  = A302 & A300;
  assign \new_[21418]_  = \new_[21417]_  & \new_[21414]_ ;
  assign \new_[21419]_  = \new_[21418]_  & \new_[21411]_ ;
  assign \new_[21423]_  = ~A166 & ~A167;
  assign \new_[21424]_  = ~A169 & \new_[21423]_ ;
  assign \new_[21428]_  = ~A203 & ~A202;
  assign \new_[21429]_  = ~A200 & \new_[21428]_ ;
  assign \new_[21430]_  = \new_[21429]_  & \new_[21424]_ ;
  assign \new_[21434]_  = A267 & ~A266;
  assign \new_[21435]_  = A265 & \new_[21434]_ ;
  assign \new_[21438]_  = A298 & A268;
  assign \new_[21441]_  = ~A302 & ~A301;
  assign \new_[21442]_  = \new_[21441]_  & \new_[21438]_ ;
  assign \new_[21443]_  = \new_[21442]_  & \new_[21435]_ ;
  assign \new_[21447]_  = ~A166 & ~A167;
  assign \new_[21448]_  = ~A169 & \new_[21447]_ ;
  assign \new_[21452]_  = ~A203 & ~A202;
  assign \new_[21453]_  = ~A200 & \new_[21452]_ ;
  assign \new_[21454]_  = \new_[21453]_  & \new_[21448]_ ;
  assign \new_[21458]_  = A267 & ~A266;
  assign \new_[21459]_  = A265 & \new_[21458]_ ;
  assign \new_[21462]_  = A298 & A269;
  assign \new_[21465]_  = ~A302 & ~A301;
  assign \new_[21466]_  = \new_[21465]_  & \new_[21462]_ ;
  assign \new_[21467]_  = \new_[21466]_  & \new_[21459]_ ;
  assign \new_[21471]_  = ~A166 & ~A167;
  assign \new_[21472]_  = ~A169 & \new_[21471]_ ;
  assign \new_[21476]_  = A201 & ~A200;
  assign \new_[21477]_  = A199 & \new_[21476]_ ;
  assign \new_[21478]_  = \new_[21477]_  & \new_[21472]_ ;
  assign \new_[21482]_  = A266 & A265;
  assign \new_[21483]_  = A202 & \new_[21482]_ ;
  assign \new_[21486]_  = ~A299 & A298;
  assign \new_[21489]_  = A301 & A300;
  assign \new_[21490]_  = \new_[21489]_  & \new_[21486]_ ;
  assign \new_[21491]_  = \new_[21490]_  & \new_[21483]_ ;
  assign \new_[21495]_  = ~A166 & ~A167;
  assign \new_[21496]_  = ~A169 & \new_[21495]_ ;
  assign \new_[21500]_  = A201 & ~A200;
  assign \new_[21501]_  = A199 & \new_[21500]_ ;
  assign \new_[21502]_  = \new_[21501]_  & \new_[21496]_ ;
  assign \new_[21506]_  = A266 & A265;
  assign \new_[21507]_  = A202 & \new_[21506]_ ;
  assign \new_[21510]_  = ~A299 & A298;
  assign \new_[21513]_  = A302 & A300;
  assign \new_[21514]_  = \new_[21513]_  & \new_[21510]_ ;
  assign \new_[21515]_  = \new_[21514]_  & \new_[21507]_ ;
  assign \new_[21519]_  = ~A166 & ~A167;
  assign \new_[21520]_  = ~A169 & \new_[21519]_ ;
  assign \new_[21524]_  = A201 & ~A200;
  assign \new_[21525]_  = A199 & \new_[21524]_ ;
  assign \new_[21526]_  = \new_[21525]_  & \new_[21520]_ ;
  assign \new_[21530]_  = ~A267 & ~A266;
  assign \new_[21531]_  = A202 & \new_[21530]_ ;
  assign \new_[21534]_  = ~A299 & A298;
  assign \new_[21537]_  = A301 & A300;
  assign \new_[21538]_  = \new_[21537]_  & \new_[21534]_ ;
  assign \new_[21539]_  = \new_[21538]_  & \new_[21531]_ ;
  assign \new_[21543]_  = ~A166 & ~A167;
  assign \new_[21544]_  = ~A169 & \new_[21543]_ ;
  assign \new_[21548]_  = A201 & ~A200;
  assign \new_[21549]_  = A199 & \new_[21548]_ ;
  assign \new_[21550]_  = \new_[21549]_  & \new_[21544]_ ;
  assign \new_[21554]_  = ~A267 & ~A266;
  assign \new_[21555]_  = A202 & \new_[21554]_ ;
  assign \new_[21558]_  = ~A299 & A298;
  assign \new_[21561]_  = A302 & A300;
  assign \new_[21562]_  = \new_[21561]_  & \new_[21558]_ ;
  assign \new_[21563]_  = \new_[21562]_  & \new_[21555]_ ;
  assign \new_[21567]_  = ~A166 & ~A167;
  assign \new_[21568]_  = ~A169 & \new_[21567]_ ;
  assign \new_[21572]_  = A201 & ~A200;
  assign \new_[21573]_  = A199 & \new_[21572]_ ;
  assign \new_[21574]_  = \new_[21573]_  & \new_[21568]_ ;
  assign \new_[21578]_  = ~A266 & ~A265;
  assign \new_[21579]_  = A202 & \new_[21578]_ ;
  assign \new_[21582]_  = ~A299 & A298;
  assign \new_[21585]_  = A301 & A300;
  assign \new_[21586]_  = \new_[21585]_  & \new_[21582]_ ;
  assign \new_[21587]_  = \new_[21586]_  & \new_[21579]_ ;
  assign \new_[21591]_  = ~A166 & ~A167;
  assign \new_[21592]_  = ~A169 & \new_[21591]_ ;
  assign \new_[21596]_  = A201 & ~A200;
  assign \new_[21597]_  = A199 & \new_[21596]_ ;
  assign \new_[21598]_  = \new_[21597]_  & \new_[21592]_ ;
  assign \new_[21602]_  = ~A266 & ~A265;
  assign \new_[21603]_  = A202 & \new_[21602]_ ;
  assign \new_[21606]_  = ~A299 & A298;
  assign \new_[21609]_  = A302 & A300;
  assign \new_[21610]_  = \new_[21609]_  & \new_[21606]_ ;
  assign \new_[21611]_  = \new_[21610]_  & \new_[21603]_ ;
  assign \new_[21615]_  = ~A166 & ~A167;
  assign \new_[21616]_  = ~A169 & \new_[21615]_ ;
  assign \new_[21620]_  = A201 & ~A200;
  assign \new_[21621]_  = A199 & \new_[21620]_ ;
  assign \new_[21622]_  = \new_[21621]_  & \new_[21616]_ ;
  assign \new_[21626]_  = A266 & A265;
  assign \new_[21627]_  = A203 & \new_[21626]_ ;
  assign \new_[21630]_  = ~A299 & A298;
  assign \new_[21633]_  = A301 & A300;
  assign \new_[21634]_  = \new_[21633]_  & \new_[21630]_ ;
  assign \new_[21635]_  = \new_[21634]_  & \new_[21627]_ ;
  assign \new_[21639]_  = ~A166 & ~A167;
  assign \new_[21640]_  = ~A169 & \new_[21639]_ ;
  assign \new_[21644]_  = A201 & ~A200;
  assign \new_[21645]_  = A199 & \new_[21644]_ ;
  assign \new_[21646]_  = \new_[21645]_  & \new_[21640]_ ;
  assign \new_[21650]_  = A266 & A265;
  assign \new_[21651]_  = A203 & \new_[21650]_ ;
  assign \new_[21654]_  = ~A299 & A298;
  assign \new_[21657]_  = A302 & A300;
  assign \new_[21658]_  = \new_[21657]_  & \new_[21654]_ ;
  assign \new_[21659]_  = \new_[21658]_  & \new_[21651]_ ;
  assign \new_[21663]_  = ~A166 & ~A167;
  assign \new_[21664]_  = ~A169 & \new_[21663]_ ;
  assign \new_[21668]_  = A201 & ~A200;
  assign \new_[21669]_  = A199 & \new_[21668]_ ;
  assign \new_[21670]_  = \new_[21669]_  & \new_[21664]_ ;
  assign \new_[21674]_  = ~A267 & ~A266;
  assign \new_[21675]_  = A203 & \new_[21674]_ ;
  assign \new_[21678]_  = ~A299 & A298;
  assign \new_[21681]_  = A301 & A300;
  assign \new_[21682]_  = \new_[21681]_  & \new_[21678]_ ;
  assign \new_[21683]_  = \new_[21682]_  & \new_[21675]_ ;
  assign \new_[21687]_  = ~A166 & ~A167;
  assign \new_[21688]_  = ~A169 & \new_[21687]_ ;
  assign \new_[21692]_  = A201 & ~A200;
  assign \new_[21693]_  = A199 & \new_[21692]_ ;
  assign \new_[21694]_  = \new_[21693]_  & \new_[21688]_ ;
  assign \new_[21698]_  = ~A267 & ~A266;
  assign \new_[21699]_  = A203 & \new_[21698]_ ;
  assign \new_[21702]_  = ~A299 & A298;
  assign \new_[21705]_  = A302 & A300;
  assign \new_[21706]_  = \new_[21705]_  & \new_[21702]_ ;
  assign \new_[21707]_  = \new_[21706]_  & \new_[21699]_ ;
  assign \new_[21711]_  = ~A166 & ~A167;
  assign \new_[21712]_  = ~A169 & \new_[21711]_ ;
  assign \new_[21716]_  = A201 & ~A200;
  assign \new_[21717]_  = A199 & \new_[21716]_ ;
  assign \new_[21718]_  = \new_[21717]_  & \new_[21712]_ ;
  assign \new_[21722]_  = ~A266 & ~A265;
  assign \new_[21723]_  = A203 & \new_[21722]_ ;
  assign \new_[21726]_  = ~A299 & A298;
  assign \new_[21729]_  = A301 & A300;
  assign \new_[21730]_  = \new_[21729]_  & \new_[21726]_ ;
  assign \new_[21731]_  = \new_[21730]_  & \new_[21723]_ ;
  assign \new_[21735]_  = ~A166 & ~A167;
  assign \new_[21736]_  = ~A169 & \new_[21735]_ ;
  assign \new_[21740]_  = A201 & ~A200;
  assign \new_[21741]_  = A199 & \new_[21740]_ ;
  assign \new_[21742]_  = \new_[21741]_  & \new_[21736]_ ;
  assign \new_[21746]_  = ~A266 & ~A265;
  assign \new_[21747]_  = A203 & \new_[21746]_ ;
  assign \new_[21750]_  = ~A299 & A298;
  assign \new_[21753]_  = A302 & A300;
  assign \new_[21754]_  = \new_[21753]_  & \new_[21750]_ ;
  assign \new_[21755]_  = \new_[21754]_  & \new_[21747]_ ;
  assign \new_[21759]_  = A167 & ~A168;
  assign \new_[21760]_  = ~A169 & \new_[21759]_ ;
  assign \new_[21764]_  = A200 & A199;
  assign \new_[21765]_  = A166 & \new_[21764]_ ;
  assign \new_[21766]_  = \new_[21765]_  & \new_[21760]_ ;
  assign \new_[21770]_  = A267 & ~A266;
  assign \new_[21771]_  = A265 & \new_[21770]_ ;
  assign \new_[21774]_  = A298 & A268;
  assign \new_[21777]_  = ~A302 & ~A301;
  assign \new_[21778]_  = \new_[21777]_  & \new_[21774]_ ;
  assign \new_[21779]_  = \new_[21778]_  & \new_[21771]_ ;
  assign \new_[21783]_  = A167 & ~A168;
  assign \new_[21784]_  = ~A169 & \new_[21783]_ ;
  assign \new_[21788]_  = A200 & A199;
  assign \new_[21789]_  = A166 & \new_[21788]_ ;
  assign \new_[21790]_  = \new_[21789]_  & \new_[21784]_ ;
  assign \new_[21794]_  = A267 & ~A266;
  assign \new_[21795]_  = A265 & \new_[21794]_ ;
  assign \new_[21798]_  = A298 & A269;
  assign \new_[21801]_  = ~A302 & ~A301;
  assign \new_[21802]_  = \new_[21801]_  & \new_[21798]_ ;
  assign \new_[21803]_  = \new_[21802]_  & \new_[21795]_ ;
  assign \new_[21807]_  = A167 & ~A168;
  assign \new_[21808]_  = ~A169 & \new_[21807]_ ;
  assign \new_[21812]_  = A200 & ~A199;
  assign \new_[21813]_  = A166 & \new_[21812]_ ;
  assign \new_[21814]_  = \new_[21813]_  & \new_[21808]_ ;
  assign \new_[21818]_  = ~A269 & ~A268;
  assign \new_[21819]_  = ~A266 & \new_[21818]_ ;
  assign \new_[21822]_  = ~A299 & A298;
  assign \new_[21825]_  = A301 & A300;
  assign \new_[21826]_  = \new_[21825]_  & \new_[21822]_ ;
  assign \new_[21827]_  = \new_[21826]_  & \new_[21819]_ ;
  assign \new_[21831]_  = A167 & ~A168;
  assign \new_[21832]_  = ~A169 & \new_[21831]_ ;
  assign \new_[21836]_  = A200 & ~A199;
  assign \new_[21837]_  = A166 & \new_[21836]_ ;
  assign \new_[21838]_  = \new_[21837]_  & \new_[21832]_ ;
  assign \new_[21842]_  = ~A269 & ~A268;
  assign \new_[21843]_  = ~A266 & \new_[21842]_ ;
  assign \new_[21846]_  = ~A299 & A298;
  assign \new_[21849]_  = A302 & A300;
  assign \new_[21850]_  = \new_[21849]_  & \new_[21846]_ ;
  assign \new_[21851]_  = \new_[21850]_  & \new_[21843]_ ;
  assign \new_[21855]_  = A167 & ~A168;
  assign \new_[21856]_  = ~A169 & \new_[21855]_ ;
  assign \new_[21860]_  = ~A202 & ~A200;
  assign \new_[21861]_  = A166 & \new_[21860]_ ;
  assign \new_[21862]_  = \new_[21861]_  & \new_[21856]_ ;
  assign \new_[21866]_  = ~A266 & A265;
  assign \new_[21867]_  = ~A203 & \new_[21866]_ ;
  assign \new_[21870]_  = A268 & A267;
  assign \new_[21873]_  = ~A300 & A298;
  assign \new_[21874]_  = \new_[21873]_  & \new_[21870]_ ;
  assign \new_[21875]_  = \new_[21874]_  & \new_[21867]_ ;
  assign \new_[21879]_  = A167 & ~A168;
  assign \new_[21880]_  = ~A169 & \new_[21879]_ ;
  assign \new_[21884]_  = ~A202 & ~A200;
  assign \new_[21885]_  = A166 & \new_[21884]_ ;
  assign \new_[21886]_  = \new_[21885]_  & \new_[21880]_ ;
  assign \new_[21890]_  = ~A266 & A265;
  assign \new_[21891]_  = ~A203 & \new_[21890]_ ;
  assign \new_[21894]_  = A268 & A267;
  assign \new_[21897]_  = A299 & A298;
  assign \new_[21898]_  = \new_[21897]_  & \new_[21894]_ ;
  assign \new_[21899]_  = \new_[21898]_  & \new_[21891]_ ;
  assign \new_[21903]_  = A167 & ~A168;
  assign \new_[21904]_  = ~A169 & \new_[21903]_ ;
  assign \new_[21908]_  = ~A202 & ~A200;
  assign \new_[21909]_  = A166 & \new_[21908]_ ;
  assign \new_[21910]_  = \new_[21909]_  & \new_[21904]_ ;
  assign \new_[21914]_  = ~A266 & A265;
  assign \new_[21915]_  = ~A203 & \new_[21914]_ ;
  assign \new_[21918]_  = A268 & A267;
  assign \new_[21921]_  = ~A299 & ~A298;
  assign \new_[21922]_  = \new_[21921]_  & \new_[21918]_ ;
  assign \new_[21923]_  = \new_[21922]_  & \new_[21915]_ ;
  assign \new_[21927]_  = A167 & ~A168;
  assign \new_[21928]_  = ~A169 & \new_[21927]_ ;
  assign \new_[21932]_  = ~A202 & ~A200;
  assign \new_[21933]_  = A166 & \new_[21932]_ ;
  assign \new_[21934]_  = \new_[21933]_  & \new_[21928]_ ;
  assign \new_[21938]_  = ~A266 & A265;
  assign \new_[21939]_  = ~A203 & \new_[21938]_ ;
  assign \new_[21942]_  = A269 & A267;
  assign \new_[21945]_  = ~A300 & A298;
  assign \new_[21946]_  = \new_[21945]_  & \new_[21942]_ ;
  assign \new_[21947]_  = \new_[21946]_  & \new_[21939]_ ;
  assign \new_[21951]_  = A167 & ~A168;
  assign \new_[21952]_  = ~A169 & \new_[21951]_ ;
  assign \new_[21956]_  = ~A202 & ~A200;
  assign \new_[21957]_  = A166 & \new_[21956]_ ;
  assign \new_[21958]_  = \new_[21957]_  & \new_[21952]_ ;
  assign \new_[21962]_  = ~A266 & A265;
  assign \new_[21963]_  = ~A203 & \new_[21962]_ ;
  assign \new_[21966]_  = A269 & A267;
  assign \new_[21969]_  = A299 & A298;
  assign \new_[21970]_  = \new_[21969]_  & \new_[21966]_ ;
  assign \new_[21971]_  = \new_[21970]_  & \new_[21963]_ ;
  assign \new_[21975]_  = A167 & ~A168;
  assign \new_[21976]_  = ~A169 & \new_[21975]_ ;
  assign \new_[21980]_  = ~A202 & ~A200;
  assign \new_[21981]_  = A166 & \new_[21980]_ ;
  assign \new_[21982]_  = \new_[21981]_  & \new_[21976]_ ;
  assign \new_[21986]_  = ~A266 & A265;
  assign \new_[21987]_  = ~A203 & \new_[21986]_ ;
  assign \new_[21990]_  = A269 & A267;
  assign \new_[21993]_  = ~A299 & ~A298;
  assign \new_[21994]_  = \new_[21993]_  & \new_[21990]_ ;
  assign \new_[21995]_  = \new_[21994]_  & \new_[21987]_ ;
  assign \new_[21999]_  = A167 & ~A168;
  assign \new_[22000]_  = ~A169 & \new_[21999]_ ;
  assign \new_[22004]_  = ~A201 & ~A200;
  assign \new_[22005]_  = A166 & \new_[22004]_ ;
  assign \new_[22006]_  = \new_[22005]_  & \new_[22000]_ ;
  assign \new_[22010]_  = A267 & ~A266;
  assign \new_[22011]_  = A265 & \new_[22010]_ ;
  assign \new_[22014]_  = A298 & A268;
  assign \new_[22017]_  = ~A302 & ~A301;
  assign \new_[22018]_  = \new_[22017]_  & \new_[22014]_ ;
  assign \new_[22019]_  = \new_[22018]_  & \new_[22011]_ ;
  assign \new_[22023]_  = A167 & ~A168;
  assign \new_[22024]_  = ~A169 & \new_[22023]_ ;
  assign \new_[22028]_  = ~A201 & ~A200;
  assign \new_[22029]_  = A166 & \new_[22028]_ ;
  assign \new_[22030]_  = \new_[22029]_  & \new_[22024]_ ;
  assign \new_[22034]_  = A267 & ~A266;
  assign \new_[22035]_  = A265 & \new_[22034]_ ;
  assign \new_[22038]_  = A298 & A269;
  assign \new_[22041]_  = ~A302 & ~A301;
  assign \new_[22042]_  = \new_[22041]_  & \new_[22038]_ ;
  assign \new_[22043]_  = \new_[22042]_  & \new_[22035]_ ;
  assign \new_[22047]_  = A167 & ~A168;
  assign \new_[22048]_  = ~A169 & \new_[22047]_ ;
  assign \new_[22052]_  = ~A200 & A199;
  assign \new_[22053]_  = A166 & \new_[22052]_ ;
  assign \new_[22054]_  = \new_[22053]_  & \new_[22048]_ ;
  assign \new_[22058]_  = ~A266 & A202;
  assign \new_[22059]_  = A201 & \new_[22058]_ ;
  assign \new_[22062]_  = ~A269 & ~A268;
  assign \new_[22065]_  = A299 & ~A298;
  assign \new_[22066]_  = \new_[22065]_  & \new_[22062]_ ;
  assign \new_[22067]_  = \new_[22066]_  & \new_[22059]_ ;
  assign \new_[22071]_  = A167 & ~A168;
  assign \new_[22072]_  = ~A169 & \new_[22071]_ ;
  assign \new_[22076]_  = ~A200 & A199;
  assign \new_[22077]_  = A166 & \new_[22076]_ ;
  assign \new_[22078]_  = \new_[22077]_  & \new_[22072]_ ;
  assign \new_[22082]_  = ~A266 & A203;
  assign \new_[22083]_  = A201 & \new_[22082]_ ;
  assign \new_[22086]_  = ~A269 & ~A268;
  assign \new_[22089]_  = A299 & ~A298;
  assign \new_[22090]_  = \new_[22089]_  & \new_[22086]_ ;
  assign \new_[22091]_  = \new_[22090]_  & \new_[22083]_ ;
  assign \new_[22095]_  = A167 & ~A168;
  assign \new_[22096]_  = ~A169 & \new_[22095]_ ;
  assign \new_[22100]_  = ~A200 & ~A199;
  assign \new_[22101]_  = A166 & \new_[22100]_ ;
  assign \new_[22102]_  = \new_[22101]_  & \new_[22096]_ ;
  assign \new_[22106]_  = A267 & ~A266;
  assign \new_[22107]_  = A265 & \new_[22106]_ ;
  assign \new_[22110]_  = A298 & A268;
  assign \new_[22113]_  = ~A302 & ~A301;
  assign \new_[22114]_  = \new_[22113]_  & \new_[22110]_ ;
  assign \new_[22115]_  = \new_[22114]_  & \new_[22107]_ ;
  assign \new_[22119]_  = A167 & ~A168;
  assign \new_[22120]_  = ~A169 & \new_[22119]_ ;
  assign \new_[22124]_  = ~A200 & ~A199;
  assign \new_[22125]_  = A166 & \new_[22124]_ ;
  assign \new_[22126]_  = \new_[22125]_  & \new_[22120]_ ;
  assign \new_[22130]_  = A267 & ~A266;
  assign \new_[22131]_  = A265 & \new_[22130]_ ;
  assign \new_[22134]_  = A298 & A269;
  assign \new_[22137]_  = ~A302 & ~A301;
  assign \new_[22138]_  = \new_[22137]_  & \new_[22134]_ ;
  assign \new_[22139]_  = \new_[22138]_  & \new_[22131]_ ;
  assign \new_[22143]_  = A167 & ~A169;
  assign \new_[22144]_  = A170 & \new_[22143]_ ;
  assign \new_[22148]_  = A200 & A199;
  assign \new_[22149]_  = ~A166 & \new_[22148]_ ;
  assign \new_[22150]_  = \new_[22149]_  & \new_[22144]_ ;
  assign \new_[22154]_  = ~A269 & ~A268;
  assign \new_[22155]_  = ~A266 & \new_[22154]_ ;
  assign \new_[22158]_  = ~A299 & A298;
  assign \new_[22161]_  = A301 & A300;
  assign \new_[22162]_  = \new_[22161]_  & \new_[22158]_ ;
  assign \new_[22163]_  = \new_[22162]_  & \new_[22155]_ ;
  assign \new_[22167]_  = A167 & ~A169;
  assign \new_[22168]_  = A170 & \new_[22167]_ ;
  assign \new_[22172]_  = A200 & A199;
  assign \new_[22173]_  = ~A166 & \new_[22172]_ ;
  assign \new_[22174]_  = \new_[22173]_  & \new_[22168]_ ;
  assign \new_[22178]_  = ~A269 & ~A268;
  assign \new_[22179]_  = ~A266 & \new_[22178]_ ;
  assign \new_[22182]_  = ~A299 & A298;
  assign \new_[22185]_  = A302 & A300;
  assign \new_[22186]_  = \new_[22185]_  & \new_[22182]_ ;
  assign \new_[22187]_  = \new_[22186]_  & \new_[22179]_ ;
  assign \new_[22191]_  = A167 & ~A169;
  assign \new_[22192]_  = A170 & \new_[22191]_ ;
  assign \new_[22196]_  = A200 & ~A199;
  assign \new_[22197]_  = ~A166 & \new_[22196]_ ;
  assign \new_[22198]_  = \new_[22197]_  & \new_[22192]_ ;
  assign \new_[22202]_  = A267 & ~A266;
  assign \new_[22203]_  = A265 & \new_[22202]_ ;
  assign \new_[22206]_  = A298 & A268;
  assign \new_[22209]_  = ~A302 & ~A301;
  assign \new_[22210]_  = \new_[22209]_  & \new_[22206]_ ;
  assign \new_[22211]_  = \new_[22210]_  & \new_[22203]_ ;
  assign \new_[22215]_  = A167 & ~A169;
  assign \new_[22216]_  = A170 & \new_[22215]_ ;
  assign \new_[22220]_  = A200 & ~A199;
  assign \new_[22221]_  = ~A166 & \new_[22220]_ ;
  assign \new_[22222]_  = \new_[22221]_  & \new_[22216]_ ;
  assign \new_[22226]_  = A267 & ~A266;
  assign \new_[22227]_  = A265 & \new_[22226]_ ;
  assign \new_[22230]_  = A298 & A269;
  assign \new_[22233]_  = ~A302 & ~A301;
  assign \new_[22234]_  = \new_[22233]_  & \new_[22230]_ ;
  assign \new_[22235]_  = \new_[22234]_  & \new_[22227]_ ;
  assign \new_[22239]_  = A167 & ~A169;
  assign \new_[22240]_  = A170 & \new_[22239]_ ;
  assign \new_[22244]_  = ~A202 & ~A200;
  assign \new_[22245]_  = ~A166 & \new_[22244]_ ;
  assign \new_[22246]_  = \new_[22245]_  & \new_[22240]_ ;
  assign \new_[22250]_  = A266 & A265;
  assign \new_[22251]_  = ~A203 & \new_[22250]_ ;
  assign \new_[22254]_  = ~A299 & A298;
  assign \new_[22257]_  = A301 & A300;
  assign \new_[22258]_  = \new_[22257]_  & \new_[22254]_ ;
  assign \new_[22259]_  = \new_[22258]_  & \new_[22251]_ ;
  assign \new_[22263]_  = A167 & ~A169;
  assign \new_[22264]_  = A170 & \new_[22263]_ ;
  assign \new_[22268]_  = ~A202 & ~A200;
  assign \new_[22269]_  = ~A166 & \new_[22268]_ ;
  assign \new_[22270]_  = \new_[22269]_  & \new_[22264]_ ;
  assign \new_[22274]_  = A266 & A265;
  assign \new_[22275]_  = ~A203 & \new_[22274]_ ;
  assign \new_[22278]_  = ~A299 & A298;
  assign \new_[22281]_  = A302 & A300;
  assign \new_[22282]_  = \new_[22281]_  & \new_[22278]_ ;
  assign \new_[22283]_  = \new_[22282]_  & \new_[22275]_ ;
  assign \new_[22287]_  = A167 & ~A169;
  assign \new_[22288]_  = A170 & \new_[22287]_ ;
  assign \new_[22292]_  = ~A202 & ~A200;
  assign \new_[22293]_  = ~A166 & \new_[22292]_ ;
  assign \new_[22294]_  = \new_[22293]_  & \new_[22288]_ ;
  assign \new_[22298]_  = ~A267 & ~A266;
  assign \new_[22299]_  = ~A203 & \new_[22298]_ ;
  assign \new_[22302]_  = ~A299 & A298;
  assign \new_[22305]_  = A301 & A300;
  assign \new_[22306]_  = \new_[22305]_  & \new_[22302]_ ;
  assign \new_[22307]_  = \new_[22306]_  & \new_[22299]_ ;
  assign \new_[22311]_  = A167 & ~A169;
  assign \new_[22312]_  = A170 & \new_[22311]_ ;
  assign \new_[22316]_  = ~A202 & ~A200;
  assign \new_[22317]_  = ~A166 & \new_[22316]_ ;
  assign \new_[22318]_  = \new_[22317]_  & \new_[22312]_ ;
  assign \new_[22322]_  = ~A267 & ~A266;
  assign \new_[22323]_  = ~A203 & \new_[22322]_ ;
  assign \new_[22326]_  = ~A299 & A298;
  assign \new_[22329]_  = A302 & A300;
  assign \new_[22330]_  = \new_[22329]_  & \new_[22326]_ ;
  assign \new_[22331]_  = \new_[22330]_  & \new_[22323]_ ;
  assign \new_[22335]_  = A167 & ~A169;
  assign \new_[22336]_  = A170 & \new_[22335]_ ;
  assign \new_[22340]_  = ~A202 & ~A200;
  assign \new_[22341]_  = ~A166 & \new_[22340]_ ;
  assign \new_[22342]_  = \new_[22341]_  & \new_[22336]_ ;
  assign \new_[22346]_  = ~A266 & ~A265;
  assign \new_[22347]_  = ~A203 & \new_[22346]_ ;
  assign \new_[22350]_  = ~A299 & A298;
  assign \new_[22353]_  = A301 & A300;
  assign \new_[22354]_  = \new_[22353]_  & \new_[22350]_ ;
  assign \new_[22355]_  = \new_[22354]_  & \new_[22347]_ ;
  assign \new_[22359]_  = A167 & ~A169;
  assign \new_[22360]_  = A170 & \new_[22359]_ ;
  assign \new_[22364]_  = ~A202 & ~A200;
  assign \new_[22365]_  = ~A166 & \new_[22364]_ ;
  assign \new_[22366]_  = \new_[22365]_  & \new_[22360]_ ;
  assign \new_[22370]_  = ~A266 & ~A265;
  assign \new_[22371]_  = ~A203 & \new_[22370]_ ;
  assign \new_[22374]_  = ~A299 & A298;
  assign \new_[22377]_  = A302 & A300;
  assign \new_[22378]_  = \new_[22377]_  & \new_[22374]_ ;
  assign \new_[22379]_  = \new_[22378]_  & \new_[22371]_ ;
  assign \new_[22383]_  = A167 & ~A169;
  assign \new_[22384]_  = A170 & \new_[22383]_ ;
  assign \new_[22388]_  = ~A201 & ~A200;
  assign \new_[22389]_  = ~A166 & \new_[22388]_ ;
  assign \new_[22390]_  = \new_[22389]_  & \new_[22384]_ ;
  assign \new_[22394]_  = ~A269 & ~A268;
  assign \new_[22395]_  = ~A266 & \new_[22394]_ ;
  assign \new_[22398]_  = ~A299 & A298;
  assign \new_[22401]_  = A301 & A300;
  assign \new_[22402]_  = \new_[22401]_  & \new_[22398]_ ;
  assign \new_[22403]_  = \new_[22402]_  & \new_[22395]_ ;
  assign \new_[22407]_  = A167 & ~A169;
  assign \new_[22408]_  = A170 & \new_[22407]_ ;
  assign \new_[22412]_  = ~A201 & ~A200;
  assign \new_[22413]_  = ~A166 & \new_[22412]_ ;
  assign \new_[22414]_  = \new_[22413]_  & \new_[22408]_ ;
  assign \new_[22418]_  = ~A269 & ~A268;
  assign \new_[22419]_  = ~A266 & \new_[22418]_ ;
  assign \new_[22422]_  = ~A299 & A298;
  assign \new_[22425]_  = A302 & A300;
  assign \new_[22426]_  = \new_[22425]_  & \new_[22422]_ ;
  assign \new_[22427]_  = \new_[22426]_  & \new_[22419]_ ;
  assign \new_[22431]_  = A167 & ~A169;
  assign \new_[22432]_  = A170 & \new_[22431]_ ;
  assign \new_[22436]_  = ~A200 & A199;
  assign \new_[22437]_  = ~A166 & \new_[22436]_ ;
  assign \new_[22438]_  = \new_[22437]_  & \new_[22432]_ ;
  assign \new_[22442]_  = ~A265 & A202;
  assign \new_[22443]_  = A201 & \new_[22442]_ ;
  assign \new_[22446]_  = A298 & A266;
  assign \new_[22449]_  = ~A302 & ~A301;
  assign \new_[22450]_  = \new_[22449]_  & \new_[22446]_ ;
  assign \new_[22451]_  = \new_[22450]_  & \new_[22443]_ ;
  assign \new_[22455]_  = A167 & ~A169;
  assign \new_[22456]_  = A170 & \new_[22455]_ ;
  assign \new_[22460]_  = ~A200 & A199;
  assign \new_[22461]_  = ~A166 & \new_[22460]_ ;
  assign \new_[22462]_  = \new_[22461]_  & \new_[22456]_ ;
  assign \new_[22466]_  = ~A265 & A203;
  assign \new_[22467]_  = A201 & \new_[22466]_ ;
  assign \new_[22470]_  = A298 & A266;
  assign \new_[22473]_  = ~A302 & ~A301;
  assign \new_[22474]_  = \new_[22473]_  & \new_[22470]_ ;
  assign \new_[22475]_  = \new_[22474]_  & \new_[22467]_ ;
  assign \new_[22479]_  = A167 & ~A169;
  assign \new_[22480]_  = A170 & \new_[22479]_ ;
  assign \new_[22484]_  = ~A200 & ~A199;
  assign \new_[22485]_  = ~A166 & \new_[22484]_ ;
  assign \new_[22486]_  = \new_[22485]_  & \new_[22480]_ ;
  assign \new_[22490]_  = ~A269 & ~A268;
  assign \new_[22491]_  = ~A266 & \new_[22490]_ ;
  assign \new_[22494]_  = ~A299 & A298;
  assign \new_[22497]_  = A301 & A300;
  assign \new_[22498]_  = \new_[22497]_  & \new_[22494]_ ;
  assign \new_[22499]_  = \new_[22498]_  & \new_[22491]_ ;
  assign \new_[22503]_  = A167 & ~A169;
  assign \new_[22504]_  = A170 & \new_[22503]_ ;
  assign \new_[22508]_  = ~A200 & ~A199;
  assign \new_[22509]_  = ~A166 & \new_[22508]_ ;
  assign \new_[22510]_  = \new_[22509]_  & \new_[22504]_ ;
  assign \new_[22514]_  = ~A269 & ~A268;
  assign \new_[22515]_  = ~A266 & \new_[22514]_ ;
  assign \new_[22518]_  = ~A299 & A298;
  assign \new_[22521]_  = A302 & A300;
  assign \new_[22522]_  = \new_[22521]_  & \new_[22518]_ ;
  assign \new_[22523]_  = \new_[22522]_  & \new_[22515]_ ;
  assign \new_[22527]_  = ~A167 & ~A169;
  assign \new_[22528]_  = A170 & \new_[22527]_ ;
  assign \new_[22532]_  = A200 & A199;
  assign \new_[22533]_  = A166 & \new_[22532]_ ;
  assign \new_[22534]_  = \new_[22533]_  & \new_[22528]_ ;
  assign \new_[22538]_  = ~A269 & ~A268;
  assign \new_[22539]_  = ~A266 & \new_[22538]_ ;
  assign \new_[22542]_  = ~A299 & A298;
  assign \new_[22545]_  = A301 & A300;
  assign \new_[22546]_  = \new_[22545]_  & \new_[22542]_ ;
  assign \new_[22547]_  = \new_[22546]_  & \new_[22539]_ ;
  assign \new_[22551]_  = ~A167 & ~A169;
  assign \new_[22552]_  = A170 & \new_[22551]_ ;
  assign \new_[22556]_  = A200 & A199;
  assign \new_[22557]_  = A166 & \new_[22556]_ ;
  assign \new_[22558]_  = \new_[22557]_  & \new_[22552]_ ;
  assign \new_[22562]_  = ~A269 & ~A268;
  assign \new_[22563]_  = ~A266 & \new_[22562]_ ;
  assign \new_[22566]_  = ~A299 & A298;
  assign \new_[22569]_  = A302 & A300;
  assign \new_[22570]_  = \new_[22569]_  & \new_[22566]_ ;
  assign \new_[22571]_  = \new_[22570]_  & \new_[22563]_ ;
  assign \new_[22575]_  = ~A167 & ~A169;
  assign \new_[22576]_  = A170 & \new_[22575]_ ;
  assign \new_[22580]_  = A200 & ~A199;
  assign \new_[22581]_  = A166 & \new_[22580]_ ;
  assign \new_[22582]_  = \new_[22581]_  & \new_[22576]_ ;
  assign \new_[22586]_  = A267 & ~A266;
  assign \new_[22587]_  = A265 & \new_[22586]_ ;
  assign \new_[22590]_  = A298 & A268;
  assign \new_[22593]_  = ~A302 & ~A301;
  assign \new_[22594]_  = \new_[22593]_  & \new_[22590]_ ;
  assign \new_[22595]_  = \new_[22594]_  & \new_[22587]_ ;
  assign \new_[22599]_  = ~A167 & ~A169;
  assign \new_[22600]_  = A170 & \new_[22599]_ ;
  assign \new_[22604]_  = A200 & ~A199;
  assign \new_[22605]_  = A166 & \new_[22604]_ ;
  assign \new_[22606]_  = \new_[22605]_  & \new_[22600]_ ;
  assign \new_[22610]_  = A267 & ~A266;
  assign \new_[22611]_  = A265 & \new_[22610]_ ;
  assign \new_[22614]_  = A298 & A269;
  assign \new_[22617]_  = ~A302 & ~A301;
  assign \new_[22618]_  = \new_[22617]_  & \new_[22614]_ ;
  assign \new_[22619]_  = \new_[22618]_  & \new_[22611]_ ;
  assign \new_[22623]_  = ~A167 & ~A169;
  assign \new_[22624]_  = A170 & \new_[22623]_ ;
  assign \new_[22628]_  = ~A202 & ~A200;
  assign \new_[22629]_  = A166 & \new_[22628]_ ;
  assign \new_[22630]_  = \new_[22629]_  & \new_[22624]_ ;
  assign \new_[22634]_  = A266 & A265;
  assign \new_[22635]_  = ~A203 & \new_[22634]_ ;
  assign \new_[22638]_  = ~A299 & A298;
  assign \new_[22641]_  = A301 & A300;
  assign \new_[22642]_  = \new_[22641]_  & \new_[22638]_ ;
  assign \new_[22643]_  = \new_[22642]_  & \new_[22635]_ ;
  assign \new_[22647]_  = ~A167 & ~A169;
  assign \new_[22648]_  = A170 & \new_[22647]_ ;
  assign \new_[22652]_  = ~A202 & ~A200;
  assign \new_[22653]_  = A166 & \new_[22652]_ ;
  assign \new_[22654]_  = \new_[22653]_  & \new_[22648]_ ;
  assign \new_[22658]_  = A266 & A265;
  assign \new_[22659]_  = ~A203 & \new_[22658]_ ;
  assign \new_[22662]_  = ~A299 & A298;
  assign \new_[22665]_  = A302 & A300;
  assign \new_[22666]_  = \new_[22665]_  & \new_[22662]_ ;
  assign \new_[22667]_  = \new_[22666]_  & \new_[22659]_ ;
  assign \new_[22671]_  = ~A167 & ~A169;
  assign \new_[22672]_  = A170 & \new_[22671]_ ;
  assign \new_[22676]_  = ~A202 & ~A200;
  assign \new_[22677]_  = A166 & \new_[22676]_ ;
  assign \new_[22678]_  = \new_[22677]_  & \new_[22672]_ ;
  assign \new_[22682]_  = ~A267 & ~A266;
  assign \new_[22683]_  = ~A203 & \new_[22682]_ ;
  assign \new_[22686]_  = ~A299 & A298;
  assign \new_[22689]_  = A301 & A300;
  assign \new_[22690]_  = \new_[22689]_  & \new_[22686]_ ;
  assign \new_[22691]_  = \new_[22690]_  & \new_[22683]_ ;
  assign \new_[22695]_  = ~A167 & ~A169;
  assign \new_[22696]_  = A170 & \new_[22695]_ ;
  assign \new_[22700]_  = ~A202 & ~A200;
  assign \new_[22701]_  = A166 & \new_[22700]_ ;
  assign \new_[22702]_  = \new_[22701]_  & \new_[22696]_ ;
  assign \new_[22706]_  = ~A267 & ~A266;
  assign \new_[22707]_  = ~A203 & \new_[22706]_ ;
  assign \new_[22710]_  = ~A299 & A298;
  assign \new_[22713]_  = A302 & A300;
  assign \new_[22714]_  = \new_[22713]_  & \new_[22710]_ ;
  assign \new_[22715]_  = \new_[22714]_  & \new_[22707]_ ;
  assign \new_[22719]_  = ~A167 & ~A169;
  assign \new_[22720]_  = A170 & \new_[22719]_ ;
  assign \new_[22724]_  = ~A202 & ~A200;
  assign \new_[22725]_  = A166 & \new_[22724]_ ;
  assign \new_[22726]_  = \new_[22725]_  & \new_[22720]_ ;
  assign \new_[22730]_  = ~A266 & ~A265;
  assign \new_[22731]_  = ~A203 & \new_[22730]_ ;
  assign \new_[22734]_  = ~A299 & A298;
  assign \new_[22737]_  = A301 & A300;
  assign \new_[22738]_  = \new_[22737]_  & \new_[22734]_ ;
  assign \new_[22739]_  = \new_[22738]_  & \new_[22731]_ ;
  assign \new_[22743]_  = ~A167 & ~A169;
  assign \new_[22744]_  = A170 & \new_[22743]_ ;
  assign \new_[22748]_  = ~A202 & ~A200;
  assign \new_[22749]_  = A166 & \new_[22748]_ ;
  assign \new_[22750]_  = \new_[22749]_  & \new_[22744]_ ;
  assign \new_[22754]_  = ~A266 & ~A265;
  assign \new_[22755]_  = ~A203 & \new_[22754]_ ;
  assign \new_[22758]_  = ~A299 & A298;
  assign \new_[22761]_  = A302 & A300;
  assign \new_[22762]_  = \new_[22761]_  & \new_[22758]_ ;
  assign \new_[22763]_  = \new_[22762]_  & \new_[22755]_ ;
  assign \new_[22767]_  = ~A167 & ~A169;
  assign \new_[22768]_  = A170 & \new_[22767]_ ;
  assign \new_[22772]_  = ~A201 & ~A200;
  assign \new_[22773]_  = A166 & \new_[22772]_ ;
  assign \new_[22774]_  = \new_[22773]_  & \new_[22768]_ ;
  assign \new_[22778]_  = ~A269 & ~A268;
  assign \new_[22779]_  = ~A266 & \new_[22778]_ ;
  assign \new_[22782]_  = ~A299 & A298;
  assign \new_[22785]_  = A301 & A300;
  assign \new_[22786]_  = \new_[22785]_  & \new_[22782]_ ;
  assign \new_[22787]_  = \new_[22786]_  & \new_[22779]_ ;
  assign \new_[22791]_  = ~A167 & ~A169;
  assign \new_[22792]_  = A170 & \new_[22791]_ ;
  assign \new_[22796]_  = ~A201 & ~A200;
  assign \new_[22797]_  = A166 & \new_[22796]_ ;
  assign \new_[22798]_  = \new_[22797]_  & \new_[22792]_ ;
  assign \new_[22802]_  = ~A269 & ~A268;
  assign \new_[22803]_  = ~A266 & \new_[22802]_ ;
  assign \new_[22806]_  = ~A299 & A298;
  assign \new_[22809]_  = A302 & A300;
  assign \new_[22810]_  = \new_[22809]_  & \new_[22806]_ ;
  assign \new_[22811]_  = \new_[22810]_  & \new_[22803]_ ;
  assign \new_[22815]_  = ~A167 & ~A169;
  assign \new_[22816]_  = A170 & \new_[22815]_ ;
  assign \new_[22820]_  = ~A200 & A199;
  assign \new_[22821]_  = A166 & \new_[22820]_ ;
  assign \new_[22822]_  = \new_[22821]_  & \new_[22816]_ ;
  assign \new_[22826]_  = ~A265 & A202;
  assign \new_[22827]_  = A201 & \new_[22826]_ ;
  assign \new_[22830]_  = A298 & A266;
  assign \new_[22833]_  = ~A302 & ~A301;
  assign \new_[22834]_  = \new_[22833]_  & \new_[22830]_ ;
  assign \new_[22835]_  = \new_[22834]_  & \new_[22827]_ ;
  assign \new_[22839]_  = ~A167 & ~A169;
  assign \new_[22840]_  = A170 & \new_[22839]_ ;
  assign \new_[22844]_  = ~A200 & A199;
  assign \new_[22845]_  = A166 & \new_[22844]_ ;
  assign \new_[22846]_  = \new_[22845]_  & \new_[22840]_ ;
  assign \new_[22850]_  = ~A265 & A203;
  assign \new_[22851]_  = A201 & \new_[22850]_ ;
  assign \new_[22854]_  = A298 & A266;
  assign \new_[22857]_  = ~A302 & ~A301;
  assign \new_[22858]_  = \new_[22857]_  & \new_[22854]_ ;
  assign \new_[22859]_  = \new_[22858]_  & \new_[22851]_ ;
  assign \new_[22863]_  = ~A167 & ~A169;
  assign \new_[22864]_  = A170 & \new_[22863]_ ;
  assign \new_[22868]_  = ~A200 & ~A199;
  assign \new_[22869]_  = A166 & \new_[22868]_ ;
  assign \new_[22870]_  = \new_[22869]_  & \new_[22864]_ ;
  assign \new_[22874]_  = ~A269 & ~A268;
  assign \new_[22875]_  = ~A266 & \new_[22874]_ ;
  assign \new_[22878]_  = ~A299 & A298;
  assign \new_[22881]_  = A301 & A300;
  assign \new_[22882]_  = \new_[22881]_  & \new_[22878]_ ;
  assign \new_[22883]_  = \new_[22882]_  & \new_[22875]_ ;
  assign \new_[22887]_  = ~A167 & ~A169;
  assign \new_[22888]_  = A170 & \new_[22887]_ ;
  assign \new_[22892]_  = ~A200 & ~A199;
  assign \new_[22893]_  = A166 & \new_[22892]_ ;
  assign \new_[22894]_  = \new_[22893]_  & \new_[22888]_ ;
  assign \new_[22898]_  = ~A269 & ~A268;
  assign \new_[22899]_  = ~A266 & \new_[22898]_ ;
  assign \new_[22902]_  = ~A299 & A298;
  assign \new_[22905]_  = A302 & A300;
  assign \new_[22906]_  = \new_[22905]_  & \new_[22902]_ ;
  assign \new_[22907]_  = \new_[22906]_  & \new_[22899]_ ;
  assign \new_[22911]_  = ~A168 & ~A169;
  assign \new_[22912]_  = ~A170 & \new_[22911]_ ;
  assign \new_[22916]_  = ~A203 & ~A202;
  assign \new_[22917]_  = ~A200 & \new_[22916]_ ;
  assign \new_[22918]_  = \new_[22917]_  & \new_[22912]_ ;
  assign \new_[22922]_  = A267 & ~A266;
  assign \new_[22923]_  = A265 & \new_[22922]_ ;
  assign \new_[22926]_  = A298 & A268;
  assign \new_[22929]_  = ~A302 & ~A301;
  assign \new_[22930]_  = \new_[22929]_  & \new_[22926]_ ;
  assign \new_[22931]_  = \new_[22930]_  & \new_[22923]_ ;
  assign \new_[22935]_  = ~A168 & ~A169;
  assign \new_[22936]_  = ~A170 & \new_[22935]_ ;
  assign \new_[22940]_  = ~A203 & ~A202;
  assign \new_[22941]_  = ~A200 & \new_[22940]_ ;
  assign \new_[22942]_  = \new_[22941]_  & \new_[22936]_ ;
  assign \new_[22946]_  = A267 & ~A266;
  assign \new_[22947]_  = A265 & \new_[22946]_ ;
  assign \new_[22950]_  = A298 & A269;
  assign \new_[22953]_  = ~A302 & ~A301;
  assign \new_[22954]_  = \new_[22953]_  & \new_[22950]_ ;
  assign \new_[22955]_  = \new_[22954]_  & \new_[22947]_ ;
  assign \new_[22959]_  = ~A168 & ~A169;
  assign \new_[22960]_  = ~A170 & \new_[22959]_ ;
  assign \new_[22964]_  = A201 & ~A200;
  assign \new_[22965]_  = A199 & \new_[22964]_ ;
  assign \new_[22966]_  = \new_[22965]_  & \new_[22960]_ ;
  assign \new_[22970]_  = A266 & A265;
  assign \new_[22971]_  = A202 & \new_[22970]_ ;
  assign \new_[22974]_  = ~A299 & A298;
  assign \new_[22977]_  = A301 & A300;
  assign \new_[22978]_  = \new_[22977]_  & \new_[22974]_ ;
  assign \new_[22979]_  = \new_[22978]_  & \new_[22971]_ ;
  assign \new_[22983]_  = ~A168 & ~A169;
  assign \new_[22984]_  = ~A170 & \new_[22983]_ ;
  assign \new_[22988]_  = A201 & ~A200;
  assign \new_[22989]_  = A199 & \new_[22988]_ ;
  assign \new_[22990]_  = \new_[22989]_  & \new_[22984]_ ;
  assign \new_[22994]_  = A266 & A265;
  assign \new_[22995]_  = A202 & \new_[22994]_ ;
  assign \new_[22998]_  = ~A299 & A298;
  assign \new_[23001]_  = A302 & A300;
  assign \new_[23002]_  = \new_[23001]_  & \new_[22998]_ ;
  assign \new_[23003]_  = \new_[23002]_  & \new_[22995]_ ;
  assign \new_[23007]_  = ~A168 & ~A169;
  assign \new_[23008]_  = ~A170 & \new_[23007]_ ;
  assign \new_[23012]_  = A201 & ~A200;
  assign \new_[23013]_  = A199 & \new_[23012]_ ;
  assign \new_[23014]_  = \new_[23013]_  & \new_[23008]_ ;
  assign \new_[23018]_  = ~A267 & ~A266;
  assign \new_[23019]_  = A202 & \new_[23018]_ ;
  assign \new_[23022]_  = ~A299 & A298;
  assign \new_[23025]_  = A301 & A300;
  assign \new_[23026]_  = \new_[23025]_  & \new_[23022]_ ;
  assign \new_[23027]_  = \new_[23026]_  & \new_[23019]_ ;
  assign \new_[23031]_  = ~A168 & ~A169;
  assign \new_[23032]_  = ~A170 & \new_[23031]_ ;
  assign \new_[23036]_  = A201 & ~A200;
  assign \new_[23037]_  = A199 & \new_[23036]_ ;
  assign \new_[23038]_  = \new_[23037]_  & \new_[23032]_ ;
  assign \new_[23042]_  = ~A267 & ~A266;
  assign \new_[23043]_  = A202 & \new_[23042]_ ;
  assign \new_[23046]_  = ~A299 & A298;
  assign \new_[23049]_  = A302 & A300;
  assign \new_[23050]_  = \new_[23049]_  & \new_[23046]_ ;
  assign \new_[23051]_  = \new_[23050]_  & \new_[23043]_ ;
  assign \new_[23055]_  = ~A168 & ~A169;
  assign \new_[23056]_  = ~A170 & \new_[23055]_ ;
  assign \new_[23060]_  = A201 & ~A200;
  assign \new_[23061]_  = A199 & \new_[23060]_ ;
  assign \new_[23062]_  = \new_[23061]_  & \new_[23056]_ ;
  assign \new_[23066]_  = ~A266 & ~A265;
  assign \new_[23067]_  = A202 & \new_[23066]_ ;
  assign \new_[23070]_  = ~A299 & A298;
  assign \new_[23073]_  = A301 & A300;
  assign \new_[23074]_  = \new_[23073]_  & \new_[23070]_ ;
  assign \new_[23075]_  = \new_[23074]_  & \new_[23067]_ ;
  assign \new_[23079]_  = ~A168 & ~A169;
  assign \new_[23080]_  = ~A170 & \new_[23079]_ ;
  assign \new_[23084]_  = A201 & ~A200;
  assign \new_[23085]_  = A199 & \new_[23084]_ ;
  assign \new_[23086]_  = \new_[23085]_  & \new_[23080]_ ;
  assign \new_[23090]_  = ~A266 & ~A265;
  assign \new_[23091]_  = A202 & \new_[23090]_ ;
  assign \new_[23094]_  = ~A299 & A298;
  assign \new_[23097]_  = A302 & A300;
  assign \new_[23098]_  = \new_[23097]_  & \new_[23094]_ ;
  assign \new_[23099]_  = \new_[23098]_  & \new_[23091]_ ;
  assign \new_[23103]_  = ~A168 & ~A169;
  assign \new_[23104]_  = ~A170 & \new_[23103]_ ;
  assign \new_[23108]_  = A201 & ~A200;
  assign \new_[23109]_  = A199 & \new_[23108]_ ;
  assign \new_[23110]_  = \new_[23109]_  & \new_[23104]_ ;
  assign \new_[23114]_  = A266 & A265;
  assign \new_[23115]_  = A203 & \new_[23114]_ ;
  assign \new_[23118]_  = ~A299 & A298;
  assign \new_[23121]_  = A301 & A300;
  assign \new_[23122]_  = \new_[23121]_  & \new_[23118]_ ;
  assign \new_[23123]_  = \new_[23122]_  & \new_[23115]_ ;
  assign \new_[23127]_  = ~A168 & ~A169;
  assign \new_[23128]_  = ~A170 & \new_[23127]_ ;
  assign \new_[23132]_  = A201 & ~A200;
  assign \new_[23133]_  = A199 & \new_[23132]_ ;
  assign \new_[23134]_  = \new_[23133]_  & \new_[23128]_ ;
  assign \new_[23138]_  = A266 & A265;
  assign \new_[23139]_  = A203 & \new_[23138]_ ;
  assign \new_[23142]_  = ~A299 & A298;
  assign \new_[23145]_  = A302 & A300;
  assign \new_[23146]_  = \new_[23145]_  & \new_[23142]_ ;
  assign \new_[23147]_  = \new_[23146]_  & \new_[23139]_ ;
  assign \new_[23151]_  = ~A168 & ~A169;
  assign \new_[23152]_  = ~A170 & \new_[23151]_ ;
  assign \new_[23156]_  = A201 & ~A200;
  assign \new_[23157]_  = A199 & \new_[23156]_ ;
  assign \new_[23158]_  = \new_[23157]_  & \new_[23152]_ ;
  assign \new_[23162]_  = ~A267 & ~A266;
  assign \new_[23163]_  = A203 & \new_[23162]_ ;
  assign \new_[23166]_  = ~A299 & A298;
  assign \new_[23169]_  = A301 & A300;
  assign \new_[23170]_  = \new_[23169]_  & \new_[23166]_ ;
  assign \new_[23171]_  = \new_[23170]_  & \new_[23163]_ ;
  assign \new_[23175]_  = ~A168 & ~A169;
  assign \new_[23176]_  = ~A170 & \new_[23175]_ ;
  assign \new_[23180]_  = A201 & ~A200;
  assign \new_[23181]_  = A199 & \new_[23180]_ ;
  assign \new_[23182]_  = \new_[23181]_  & \new_[23176]_ ;
  assign \new_[23186]_  = ~A267 & ~A266;
  assign \new_[23187]_  = A203 & \new_[23186]_ ;
  assign \new_[23190]_  = ~A299 & A298;
  assign \new_[23193]_  = A302 & A300;
  assign \new_[23194]_  = \new_[23193]_  & \new_[23190]_ ;
  assign \new_[23195]_  = \new_[23194]_  & \new_[23187]_ ;
  assign \new_[23199]_  = ~A168 & ~A169;
  assign \new_[23200]_  = ~A170 & \new_[23199]_ ;
  assign \new_[23204]_  = A201 & ~A200;
  assign \new_[23205]_  = A199 & \new_[23204]_ ;
  assign \new_[23206]_  = \new_[23205]_  & \new_[23200]_ ;
  assign \new_[23210]_  = ~A266 & ~A265;
  assign \new_[23211]_  = A203 & \new_[23210]_ ;
  assign \new_[23214]_  = ~A299 & A298;
  assign \new_[23217]_  = A301 & A300;
  assign \new_[23218]_  = \new_[23217]_  & \new_[23214]_ ;
  assign \new_[23219]_  = \new_[23218]_  & \new_[23211]_ ;
  assign \new_[23223]_  = ~A168 & ~A169;
  assign \new_[23224]_  = ~A170 & \new_[23223]_ ;
  assign \new_[23228]_  = A201 & ~A200;
  assign \new_[23229]_  = A199 & \new_[23228]_ ;
  assign \new_[23230]_  = \new_[23229]_  & \new_[23224]_ ;
  assign \new_[23234]_  = ~A266 & ~A265;
  assign \new_[23235]_  = A203 & \new_[23234]_ ;
  assign \new_[23238]_  = ~A299 & A298;
  assign \new_[23241]_  = A302 & A300;
  assign \new_[23242]_  = \new_[23241]_  & \new_[23238]_ ;
  assign \new_[23243]_  = \new_[23242]_  & \new_[23235]_ ;
  assign \new_[23247]_  = ~A166 & ~A167;
  assign \new_[23248]_  = A170 & \new_[23247]_ ;
  assign \new_[23251]_  = ~A200 & A199;
  assign \new_[23254]_  = A202 & A201;
  assign \new_[23255]_  = \new_[23254]_  & \new_[23251]_ ;
  assign \new_[23256]_  = \new_[23255]_  & \new_[23248]_ ;
  assign \new_[23260]_  = ~A269 & ~A268;
  assign \new_[23261]_  = ~A266 & \new_[23260]_ ;
  assign \new_[23264]_  = ~A299 & A298;
  assign \new_[23267]_  = A301 & A300;
  assign \new_[23268]_  = \new_[23267]_  & \new_[23264]_ ;
  assign \new_[23269]_  = \new_[23268]_  & \new_[23261]_ ;
  assign \new_[23273]_  = ~A166 & ~A167;
  assign \new_[23274]_  = A170 & \new_[23273]_ ;
  assign \new_[23277]_  = ~A200 & A199;
  assign \new_[23280]_  = A202 & A201;
  assign \new_[23281]_  = \new_[23280]_  & \new_[23277]_ ;
  assign \new_[23282]_  = \new_[23281]_  & \new_[23274]_ ;
  assign \new_[23286]_  = ~A269 & ~A268;
  assign \new_[23287]_  = ~A266 & \new_[23286]_ ;
  assign \new_[23290]_  = ~A299 & A298;
  assign \new_[23293]_  = A302 & A300;
  assign \new_[23294]_  = \new_[23293]_  & \new_[23290]_ ;
  assign \new_[23295]_  = \new_[23294]_  & \new_[23287]_ ;
  assign \new_[23299]_  = ~A166 & ~A167;
  assign \new_[23300]_  = A170 & \new_[23299]_ ;
  assign \new_[23303]_  = ~A200 & A199;
  assign \new_[23306]_  = A203 & A201;
  assign \new_[23307]_  = \new_[23306]_  & \new_[23303]_ ;
  assign \new_[23308]_  = \new_[23307]_  & \new_[23300]_ ;
  assign \new_[23312]_  = ~A269 & ~A268;
  assign \new_[23313]_  = ~A266 & \new_[23312]_ ;
  assign \new_[23316]_  = ~A299 & A298;
  assign \new_[23319]_  = A301 & A300;
  assign \new_[23320]_  = \new_[23319]_  & \new_[23316]_ ;
  assign \new_[23321]_  = \new_[23320]_  & \new_[23313]_ ;
  assign \new_[23325]_  = ~A166 & ~A167;
  assign \new_[23326]_  = A170 & \new_[23325]_ ;
  assign \new_[23329]_  = ~A200 & A199;
  assign \new_[23332]_  = A203 & A201;
  assign \new_[23333]_  = \new_[23332]_  & \new_[23329]_ ;
  assign \new_[23334]_  = \new_[23333]_  & \new_[23326]_ ;
  assign \new_[23338]_  = ~A269 & ~A268;
  assign \new_[23339]_  = ~A266 & \new_[23338]_ ;
  assign \new_[23342]_  = ~A299 & A298;
  assign \new_[23345]_  = A302 & A300;
  assign \new_[23346]_  = \new_[23345]_  & \new_[23342]_ ;
  assign \new_[23347]_  = \new_[23346]_  & \new_[23339]_ ;
  assign \new_[23351]_  = A167 & ~A168;
  assign \new_[23352]_  = A169 & \new_[23351]_ ;
  assign \new_[23355]_  = ~A200 & ~A166;
  assign \new_[23358]_  = ~A203 & ~A202;
  assign \new_[23359]_  = \new_[23358]_  & \new_[23355]_ ;
  assign \new_[23360]_  = \new_[23359]_  & \new_[23352]_ ;
  assign \new_[23364]_  = A267 & ~A266;
  assign \new_[23365]_  = A265 & \new_[23364]_ ;
  assign \new_[23368]_  = A298 & A268;
  assign \new_[23371]_  = ~A302 & ~A301;
  assign \new_[23372]_  = \new_[23371]_  & \new_[23368]_ ;
  assign \new_[23373]_  = \new_[23372]_  & \new_[23365]_ ;
  assign \new_[23377]_  = A167 & ~A168;
  assign \new_[23378]_  = A169 & \new_[23377]_ ;
  assign \new_[23381]_  = ~A200 & ~A166;
  assign \new_[23384]_  = ~A203 & ~A202;
  assign \new_[23385]_  = \new_[23384]_  & \new_[23381]_ ;
  assign \new_[23386]_  = \new_[23385]_  & \new_[23378]_ ;
  assign \new_[23390]_  = A267 & ~A266;
  assign \new_[23391]_  = A265 & \new_[23390]_ ;
  assign \new_[23394]_  = A298 & A269;
  assign \new_[23397]_  = ~A302 & ~A301;
  assign \new_[23398]_  = \new_[23397]_  & \new_[23394]_ ;
  assign \new_[23399]_  = \new_[23398]_  & \new_[23391]_ ;
  assign \new_[23403]_  = A167 & ~A168;
  assign \new_[23404]_  = A169 & \new_[23403]_ ;
  assign \new_[23407]_  = A199 & ~A166;
  assign \new_[23410]_  = A201 & ~A200;
  assign \new_[23411]_  = \new_[23410]_  & \new_[23407]_ ;
  assign \new_[23412]_  = \new_[23411]_  & \new_[23404]_ ;
  assign \new_[23416]_  = A266 & A265;
  assign \new_[23417]_  = A202 & \new_[23416]_ ;
  assign \new_[23420]_  = ~A299 & A298;
  assign \new_[23423]_  = A301 & A300;
  assign \new_[23424]_  = \new_[23423]_  & \new_[23420]_ ;
  assign \new_[23425]_  = \new_[23424]_  & \new_[23417]_ ;
  assign \new_[23429]_  = A167 & ~A168;
  assign \new_[23430]_  = A169 & \new_[23429]_ ;
  assign \new_[23433]_  = A199 & ~A166;
  assign \new_[23436]_  = A201 & ~A200;
  assign \new_[23437]_  = \new_[23436]_  & \new_[23433]_ ;
  assign \new_[23438]_  = \new_[23437]_  & \new_[23430]_ ;
  assign \new_[23442]_  = A266 & A265;
  assign \new_[23443]_  = A202 & \new_[23442]_ ;
  assign \new_[23446]_  = ~A299 & A298;
  assign \new_[23449]_  = A302 & A300;
  assign \new_[23450]_  = \new_[23449]_  & \new_[23446]_ ;
  assign \new_[23451]_  = \new_[23450]_  & \new_[23443]_ ;
  assign \new_[23455]_  = A167 & ~A168;
  assign \new_[23456]_  = A169 & \new_[23455]_ ;
  assign \new_[23459]_  = A199 & ~A166;
  assign \new_[23462]_  = A201 & ~A200;
  assign \new_[23463]_  = \new_[23462]_  & \new_[23459]_ ;
  assign \new_[23464]_  = \new_[23463]_  & \new_[23456]_ ;
  assign \new_[23468]_  = ~A267 & ~A266;
  assign \new_[23469]_  = A202 & \new_[23468]_ ;
  assign \new_[23472]_  = ~A299 & A298;
  assign \new_[23475]_  = A301 & A300;
  assign \new_[23476]_  = \new_[23475]_  & \new_[23472]_ ;
  assign \new_[23477]_  = \new_[23476]_  & \new_[23469]_ ;
  assign \new_[23481]_  = A167 & ~A168;
  assign \new_[23482]_  = A169 & \new_[23481]_ ;
  assign \new_[23485]_  = A199 & ~A166;
  assign \new_[23488]_  = A201 & ~A200;
  assign \new_[23489]_  = \new_[23488]_  & \new_[23485]_ ;
  assign \new_[23490]_  = \new_[23489]_  & \new_[23482]_ ;
  assign \new_[23494]_  = ~A267 & ~A266;
  assign \new_[23495]_  = A202 & \new_[23494]_ ;
  assign \new_[23498]_  = ~A299 & A298;
  assign \new_[23501]_  = A302 & A300;
  assign \new_[23502]_  = \new_[23501]_  & \new_[23498]_ ;
  assign \new_[23503]_  = \new_[23502]_  & \new_[23495]_ ;
  assign \new_[23507]_  = A167 & ~A168;
  assign \new_[23508]_  = A169 & \new_[23507]_ ;
  assign \new_[23511]_  = A199 & ~A166;
  assign \new_[23514]_  = A201 & ~A200;
  assign \new_[23515]_  = \new_[23514]_  & \new_[23511]_ ;
  assign \new_[23516]_  = \new_[23515]_  & \new_[23508]_ ;
  assign \new_[23520]_  = ~A266 & ~A265;
  assign \new_[23521]_  = A202 & \new_[23520]_ ;
  assign \new_[23524]_  = ~A299 & A298;
  assign \new_[23527]_  = A301 & A300;
  assign \new_[23528]_  = \new_[23527]_  & \new_[23524]_ ;
  assign \new_[23529]_  = \new_[23528]_  & \new_[23521]_ ;
  assign \new_[23533]_  = A167 & ~A168;
  assign \new_[23534]_  = A169 & \new_[23533]_ ;
  assign \new_[23537]_  = A199 & ~A166;
  assign \new_[23540]_  = A201 & ~A200;
  assign \new_[23541]_  = \new_[23540]_  & \new_[23537]_ ;
  assign \new_[23542]_  = \new_[23541]_  & \new_[23534]_ ;
  assign \new_[23546]_  = ~A266 & ~A265;
  assign \new_[23547]_  = A202 & \new_[23546]_ ;
  assign \new_[23550]_  = ~A299 & A298;
  assign \new_[23553]_  = A302 & A300;
  assign \new_[23554]_  = \new_[23553]_  & \new_[23550]_ ;
  assign \new_[23555]_  = \new_[23554]_  & \new_[23547]_ ;
  assign \new_[23559]_  = A167 & ~A168;
  assign \new_[23560]_  = A169 & \new_[23559]_ ;
  assign \new_[23563]_  = A199 & ~A166;
  assign \new_[23566]_  = A201 & ~A200;
  assign \new_[23567]_  = \new_[23566]_  & \new_[23563]_ ;
  assign \new_[23568]_  = \new_[23567]_  & \new_[23560]_ ;
  assign \new_[23572]_  = A266 & A265;
  assign \new_[23573]_  = A203 & \new_[23572]_ ;
  assign \new_[23576]_  = ~A299 & A298;
  assign \new_[23579]_  = A301 & A300;
  assign \new_[23580]_  = \new_[23579]_  & \new_[23576]_ ;
  assign \new_[23581]_  = \new_[23580]_  & \new_[23573]_ ;
  assign \new_[23585]_  = A167 & ~A168;
  assign \new_[23586]_  = A169 & \new_[23585]_ ;
  assign \new_[23589]_  = A199 & ~A166;
  assign \new_[23592]_  = A201 & ~A200;
  assign \new_[23593]_  = \new_[23592]_  & \new_[23589]_ ;
  assign \new_[23594]_  = \new_[23593]_  & \new_[23586]_ ;
  assign \new_[23598]_  = A266 & A265;
  assign \new_[23599]_  = A203 & \new_[23598]_ ;
  assign \new_[23602]_  = ~A299 & A298;
  assign \new_[23605]_  = A302 & A300;
  assign \new_[23606]_  = \new_[23605]_  & \new_[23602]_ ;
  assign \new_[23607]_  = \new_[23606]_  & \new_[23599]_ ;
  assign \new_[23611]_  = A167 & ~A168;
  assign \new_[23612]_  = A169 & \new_[23611]_ ;
  assign \new_[23615]_  = A199 & ~A166;
  assign \new_[23618]_  = A201 & ~A200;
  assign \new_[23619]_  = \new_[23618]_  & \new_[23615]_ ;
  assign \new_[23620]_  = \new_[23619]_  & \new_[23612]_ ;
  assign \new_[23624]_  = ~A267 & ~A266;
  assign \new_[23625]_  = A203 & \new_[23624]_ ;
  assign \new_[23628]_  = ~A299 & A298;
  assign \new_[23631]_  = A301 & A300;
  assign \new_[23632]_  = \new_[23631]_  & \new_[23628]_ ;
  assign \new_[23633]_  = \new_[23632]_  & \new_[23625]_ ;
  assign \new_[23637]_  = A167 & ~A168;
  assign \new_[23638]_  = A169 & \new_[23637]_ ;
  assign \new_[23641]_  = A199 & ~A166;
  assign \new_[23644]_  = A201 & ~A200;
  assign \new_[23645]_  = \new_[23644]_  & \new_[23641]_ ;
  assign \new_[23646]_  = \new_[23645]_  & \new_[23638]_ ;
  assign \new_[23650]_  = ~A267 & ~A266;
  assign \new_[23651]_  = A203 & \new_[23650]_ ;
  assign \new_[23654]_  = ~A299 & A298;
  assign \new_[23657]_  = A302 & A300;
  assign \new_[23658]_  = \new_[23657]_  & \new_[23654]_ ;
  assign \new_[23659]_  = \new_[23658]_  & \new_[23651]_ ;
  assign \new_[23663]_  = A167 & ~A168;
  assign \new_[23664]_  = A169 & \new_[23663]_ ;
  assign \new_[23667]_  = A199 & ~A166;
  assign \new_[23670]_  = A201 & ~A200;
  assign \new_[23671]_  = \new_[23670]_  & \new_[23667]_ ;
  assign \new_[23672]_  = \new_[23671]_  & \new_[23664]_ ;
  assign \new_[23676]_  = ~A266 & ~A265;
  assign \new_[23677]_  = A203 & \new_[23676]_ ;
  assign \new_[23680]_  = ~A299 & A298;
  assign \new_[23683]_  = A301 & A300;
  assign \new_[23684]_  = \new_[23683]_  & \new_[23680]_ ;
  assign \new_[23685]_  = \new_[23684]_  & \new_[23677]_ ;
  assign \new_[23689]_  = A167 & ~A168;
  assign \new_[23690]_  = A169 & \new_[23689]_ ;
  assign \new_[23693]_  = A199 & ~A166;
  assign \new_[23696]_  = A201 & ~A200;
  assign \new_[23697]_  = \new_[23696]_  & \new_[23693]_ ;
  assign \new_[23698]_  = \new_[23697]_  & \new_[23690]_ ;
  assign \new_[23702]_  = ~A266 & ~A265;
  assign \new_[23703]_  = A203 & \new_[23702]_ ;
  assign \new_[23706]_  = ~A299 & A298;
  assign \new_[23709]_  = A302 & A300;
  assign \new_[23710]_  = \new_[23709]_  & \new_[23706]_ ;
  assign \new_[23711]_  = \new_[23710]_  & \new_[23703]_ ;
  assign \new_[23715]_  = ~A167 & ~A168;
  assign \new_[23716]_  = A169 & \new_[23715]_ ;
  assign \new_[23719]_  = ~A200 & A166;
  assign \new_[23722]_  = ~A203 & ~A202;
  assign \new_[23723]_  = \new_[23722]_  & \new_[23719]_ ;
  assign \new_[23724]_  = \new_[23723]_  & \new_[23716]_ ;
  assign \new_[23728]_  = A267 & ~A266;
  assign \new_[23729]_  = A265 & \new_[23728]_ ;
  assign \new_[23732]_  = A298 & A268;
  assign \new_[23735]_  = ~A302 & ~A301;
  assign \new_[23736]_  = \new_[23735]_  & \new_[23732]_ ;
  assign \new_[23737]_  = \new_[23736]_  & \new_[23729]_ ;
  assign \new_[23741]_  = ~A167 & ~A168;
  assign \new_[23742]_  = A169 & \new_[23741]_ ;
  assign \new_[23745]_  = ~A200 & A166;
  assign \new_[23748]_  = ~A203 & ~A202;
  assign \new_[23749]_  = \new_[23748]_  & \new_[23745]_ ;
  assign \new_[23750]_  = \new_[23749]_  & \new_[23742]_ ;
  assign \new_[23754]_  = A267 & ~A266;
  assign \new_[23755]_  = A265 & \new_[23754]_ ;
  assign \new_[23758]_  = A298 & A269;
  assign \new_[23761]_  = ~A302 & ~A301;
  assign \new_[23762]_  = \new_[23761]_  & \new_[23758]_ ;
  assign \new_[23763]_  = \new_[23762]_  & \new_[23755]_ ;
  assign \new_[23767]_  = ~A167 & ~A168;
  assign \new_[23768]_  = A169 & \new_[23767]_ ;
  assign \new_[23771]_  = A199 & A166;
  assign \new_[23774]_  = A201 & ~A200;
  assign \new_[23775]_  = \new_[23774]_  & \new_[23771]_ ;
  assign \new_[23776]_  = \new_[23775]_  & \new_[23768]_ ;
  assign \new_[23780]_  = A266 & A265;
  assign \new_[23781]_  = A202 & \new_[23780]_ ;
  assign \new_[23784]_  = ~A299 & A298;
  assign \new_[23787]_  = A301 & A300;
  assign \new_[23788]_  = \new_[23787]_  & \new_[23784]_ ;
  assign \new_[23789]_  = \new_[23788]_  & \new_[23781]_ ;
  assign \new_[23793]_  = ~A167 & ~A168;
  assign \new_[23794]_  = A169 & \new_[23793]_ ;
  assign \new_[23797]_  = A199 & A166;
  assign \new_[23800]_  = A201 & ~A200;
  assign \new_[23801]_  = \new_[23800]_  & \new_[23797]_ ;
  assign \new_[23802]_  = \new_[23801]_  & \new_[23794]_ ;
  assign \new_[23806]_  = A266 & A265;
  assign \new_[23807]_  = A202 & \new_[23806]_ ;
  assign \new_[23810]_  = ~A299 & A298;
  assign \new_[23813]_  = A302 & A300;
  assign \new_[23814]_  = \new_[23813]_  & \new_[23810]_ ;
  assign \new_[23815]_  = \new_[23814]_  & \new_[23807]_ ;
  assign \new_[23819]_  = ~A167 & ~A168;
  assign \new_[23820]_  = A169 & \new_[23819]_ ;
  assign \new_[23823]_  = A199 & A166;
  assign \new_[23826]_  = A201 & ~A200;
  assign \new_[23827]_  = \new_[23826]_  & \new_[23823]_ ;
  assign \new_[23828]_  = \new_[23827]_  & \new_[23820]_ ;
  assign \new_[23832]_  = ~A267 & ~A266;
  assign \new_[23833]_  = A202 & \new_[23832]_ ;
  assign \new_[23836]_  = ~A299 & A298;
  assign \new_[23839]_  = A301 & A300;
  assign \new_[23840]_  = \new_[23839]_  & \new_[23836]_ ;
  assign \new_[23841]_  = \new_[23840]_  & \new_[23833]_ ;
  assign \new_[23845]_  = ~A167 & ~A168;
  assign \new_[23846]_  = A169 & \new_[23845]_ ;
  assign \new_[23849]_  = A199 & A166;
  assign \new_[23852]_  = A201 & ~A200;
  assign \new_[23853]_  = \new_[23852]_  & \new_[23849]_ ;
  assign \new_[23854]_  = \new_[23853]_  & \new_[23846]_ ;
  assign \new_[23858]_  = ~A267 & ~A266;
  assign \new_[23859]_  = A202 & \new_[23858]_ ;
  assign \new_[23862]_  = ~A299 & A298;
  assign \new_[23865]_  = A302 & A300;
  assign \new_[23866]_  = \new_[23865]_  & \new_[23862]_ ;
  assign \new_[23867]_  = \new_[23866]_  & \new_[23859]_ ;
  assign \new_[23871]_  = ~A167 & ~A168;
  assign \new_[23872]_  = A169 & \new_[23871]_ ;
  assign \new_[23875]_  = A199 & A166;
  assign \new_[23878]_  = A201 & ~A200;
  assign \new_[23879]_  = \new_[23878]_  & \new_[23875]_ ;
  assign \new_[23880]_  = \new_[23879]_  & \new_[23872]_ ;
  assign \new_[23884]_  = ~A266 & ~A265;
  assign \new_[23885]_  = A202 & \new_[23884]_ ;
  assign \new_[23888]_  = ~A299 & A298;
  assign \new_[23891]_  = A301 & A300;
  assign \new_[23892]_  = \new_[23891]_  & \new_[23888]_ ;
  assign \new_[23893]_  = \new_[23892]_  & \new_[23885]_ ;
  assign \new_[23897]_  = ~A167 & ~A168;
  assign \new_[23898]_  = A169 & \new_[23897]_ ;
  assign \new_[23901]_  = A199 & A166;
  assign \new_[23904]_  = A201 & ~A200;
  assign \new_[23905]_  = \new_[23904]_  & \new_[23901]_ ;
  assign \new_[23906]_  = \new_[23905]_  & \new_[23898]_ ;
  assign \new_[23910]_  = ~A266 & ~A265;
  assign \new_[23911]_  = A202 & \new_[23910]_ ;
  assign \new_[23914]_  = ~A299 & A298;
  assign \new_[23917]_  = A302 & A300;
  assign \new_[23918]_  = \new_[23917]_  & \new_[23914]_ ;
  assign \new_[23919]_  = \new_[23918]_  & \new_[23911]_ ;
  assign \new_[23923]_  = ~A167 & ~A168;
  assign \new_[23924]_  = A169 & \new_[23923]_ ;
  assign \new_[23927]_  = A199 & A166;
  assign \new_[23930]_  = A201 & ~A200;
  assign \new_[23931]_  = \new_[23930]_  & \new_[23927]_ ;
  assign \new_[23932]_  = \new_[23931]_  & \new_[23924]_ ;
  assign \new_[23936]_  = A266 & A265;
  assign \new_[23937]_  = A203 & \new_[23936]_ ;
  assign \new_[23940]_  = ~A299 & A298;
  assign \new_[23943]_  = A301 & A300;
  assign \new_[23944]_  = \new_[23943]_  & \new_[23940]_ ;
  assign \new_[23945]_  = \new_[23944]_  & \new_[23937]_ ;
  assign \new_[23949]_  = ~A167 & ~A168;
  assign \new_[23950]_  = A169 & \new_[23949]_ ;
  assign \new_[23953]_  = A199 & A166;
  assign \new_[23956]_  = A201 & ~A200;
  assign \new_[23957]_  = \new_[23956]_  & \new_[23953]_ ;
  assign \new_[23958]_  = \new_[23957]_  & \new_[23950]_ ;
  assign \new_[23962]_  = A266 & A265;
  assign \new_[23963]_  = A203 & \new_[23962]_ ;
  assign \new_[23966]_  = ~A299 & A298;
  assign \new_[23969]_  = A302 & A300;
  assign \new_[23970]_  = \new_[23969]_  & \new_[23966]_ ;
  assign \new_[23971]_  = \new_[23970]_  & \new_[23963]_ ;
  assign \new_[23975]_  = ~A167 & ~A168;
  assign \new_[23976]_  = A169 & \new_[23975]_ ;
  assign \new_[23979]_  = A199 & A166;
  assign \new_[23982]_  = A201 & ~A200;
  assign \new_[23983]_  = \new_[23982]_  & \new_[23979]_ ;
  assign \new_[23984]_  = \new_[23983]_  & \new_[23976]_ ;
  assign \new_[23988]_  = ~A267 & ~A266;
  assign \new_[23989]_  = A203 & \new_[23988]_ ;
  assign \new_[23992]_  = ~A299 & A298;
  assign \new_[23995]_  = A301 & A300;
  assign \new_[23996]_  = \new_[23995]_  & \new_[23992]_ ;
  assign \new_[23997]_  = \new_[23996]_  & \new_[23989]_ ;
  assign \new_[24001]_  = ~A167 & ~A168;
  assign \new_[24002]_  = A169 & \new_[24001]_ ;
  assign \new_[24005]_  = A199 & A166;
  assign \new_[24008]_  = A201 & ~A200;
  assign \new_[24009]_  = \new_[24008]_  & \new_[24005]_ ;
  assign \new_[24010]_  = \new_[24009]_  & \new_[24002]_ ;
  assign \new_[24014]_  = ~A267 & ~A266;
  assign \new_[24015]_  = A203 & \new_[24014]_ ;
  assign \new_[24018]_  = ~A299 & A298;
  assign \new_[24021]_  = A302 & A300;
  assign \new_[24022]_  = \new_[24021]_  & \new_[24018]_ ;
  assign \new_[24023]_  = \new_[24022]_  & \new_[24015]_ ;
  assign \new_[24027]_  = ~A167 & ~A168;
  assign \new_[24028]_  = A169 & \new_[24027]_ ;
  assign \new_[24031]_  = A199 & A166;
  assign \new_[24034]_  = A201 & ~A200;
  assign \new_[24035]_  = \new_[24034]_  & \new_[24031]_ ;
  assign \new_[24036]_  = \new_[24035]_  & \new_[24028]_ ;
  assign \new_[24040]_  = ~A266 & ~A265;
  assign \new_[24041]_  = A203 & \new_[24040]_ ;
  assign \new_[24044]_  = ~A299 & A298;
  assign \new_[24047]_  = A301 & A300;
  assign \new_[24048]_  = \new_[24047]_  & \new_[24044]_ ;
  assign \new_[24049]_  = \new_[24048]_  & \new_[24041]_ ;
  assign \new_[24053]_  = ~A167 & ~A168;
  assign \new_[24054]_  = A169 & \new_[24053]_ ;
  assign \new_[24057]_  = A199 & A166;
  assign \new_[24060]_  = A201 & ~A200;
  assign \new_[24061]_  = \new_[24060]_  & \new_[24057]_ ;
  assign \new_[24062]_  = \new_[24061]_  & \new_[24054]_ ;
  assign \new_[24066]_  = ~A266 & ~A265;
  assign \new_[24067]_  = A203 & \new_[24066]_ ;
  assign \new_[24070]_  = ~A299 & A298;
  assign \new_[24073]_  = A302 & A300;
  assign \new_[24074]_  = \new_[24073]_  & \new_[24070]_ ;
  assign \new_[24075]_  = \new_[24074]_  & \new_[24067]_ ;
  assign \new_[24079]_  = ~A168 & A169;
  assign \new_[24080]_  = A170 & \new_[24079]_ ;
  assign \new_[24083]_  = ~A200 & A199;
  assign \new_[24086]_  = A202 & A201;
  assign \new_[24087]_  = \new_[24086]_  & \new_[24083]_ ;
  assign \new_[24088]_  = \new_[24087]_  & \new_[24080]_ ;
  assign \new_[24092]_  = ~A269 & ~A268;
  assign \new_[24093]_  = ~A266 & \new_[24092]_ ;
  assign \new_[24096]_  = ~A299 & A298;
  assign \new_[24099]_  = A301 & A300;
  assign \new_[24100]_  = \new_[24099]_  & \new_[24096]_ ;
  assign \new_[24101]_  = \new_[24100]_  & \new_[24093]_ ;
  assign \new_[24105]_  = ~A168 & A169;
  assign \new_[24106]_  = A170 & \new_[24105]_ ;
  assign \new_[24109]_  = ~A200 & A199;
  assign \new_[24112]_  = A202 & A201;
  assign \new_[24113]_  = \new_[24112]_  & \new_[24109]_ ;
  assign \new_[24114]_  = \new_[24113]_  & \new_[24106]_ ;
  assign \new_[24118]_  = ~A269 & ~A268;
  assign \new_[24119]_  = ~A266 & \new_[24118]_ ;
  assign \new_[24122]_  = ~A299 & A298;
  assign \new_[24125]_  = A302 & A300;
  assign \new_[24126]_  = \new_[24125]_  & \new_[24122]_ ;
  assign \new_[24127]_  = \new_[24126]_  & \new_[24119]_ ;
  assign \new_[24131]_  = ~A168 & A169;
  assign \new_[24132]_  = A170 & \new_[24131]_ ;
  assign \new_[24135]_  = ~A200 & A199;
  assign \new_[24138]_  = A203 & A201;
  assign \new_[24139]_  = \new_[24138]_  & \new_[24135]_ ;
  assign \new_[24140]_  = \new_[24139]_  & \new_[24132]_ ;
  assign \new_[24144]_  = ~A269 & ~A268;
  assign \new_[24145]_  = ~A266 & \new_[24144]_ ;
  assign \new_[24148]_  = ~A299 & A298;
  assign \new_[24151]_  = A301 & A300;
  assign \new_[24152]_  = \new_[24151]_  & \new_[24148]_ ;
  assign \new_[24153]_  = \new_[24152]_  & \new_[24145]_ ;
  assign \new_[24157]_  = ~A168 & A169;
  assign \new_[24158]_  = A170 & \new_[24157]_ ;
  assign \new_[24161]_  = ~A200 & A199;
  assign \new_[24164]_  = A203 & A201;
  assign \new_[24165]_  = \new_[24164]_  & \new_[24161]_ ;
  assign \new_[24166]_  = \new_[24165]_  & \new_[24158]_ ;
  assign \new_[24170]_  = ~A269 & ~A268;
  assign \new_[24171]_  = ~A266 & \new_[24170]_ ;
  assign \new_[24174]_  = ~A299 & A298;
  assign \new_[24177]_  = A302 & A300;
  assign \new_[24178]_  = \new_[24177]_  & \new_[24174]_ ;
  assign \new_[24179]_  = \new_[24178]_  & \new_[24171]_ ;
  assign \new_[24183]_  = A167 & A169;
  assign \new_[24184]_  = ~A170 & \new_[24183]_ ;
  assign \new_[24187]_  = ~A200 & A166;
  assign \new_[24190]_  = ~A203 & ~A202;
  assign \new_[24191]_  = \new_[24190]_  & \new_[24187]_ ;
  assign \new_[24192]_  = \new_[24191]_  & \new_[24184]_ ;
  assign \new_[24196]_  = ~A269 & ~A268;
  assign \new_[24197]_  = ~A266 & \new_[24196]_ ;
  assign \new_[24200]_  = ~A299 & A298;
  assign \new_[24203]_  = A301 & A300;
  assign \new_[24204]_  = \new_[24203]_  & \new_[24200]_ ;
  assign \new_[24205]_  = \new_[24204]_  & \new_[24197]_ ;
  assign \new_[24209]_  = A167 & A169;
  assign \new_[24210]_  = ~A170 & \new_[24209]_ ;
  assign \new_[24213]_  = ~A200 & A166;
  assign \new_[24216]_  = ~A203 & ~A202;
  assign \new_[24217]_  = \new_[24216]_  & \new_[24213]_ ;
  assign \new_[24218]_  = \new_[24217]_  & \new_[24210]_ ;
  assign \new_[24222]_  = ~A269 & ~A268;
  assign \new_[24223]_  = ~A266 & \new_[24222]_ ;
  assign \new_[24226]_  = ~A299 & A298;
  assign \new_[24229]_  = A302 & A300;
  assign \new_[24230]_  = \new_[24229]_  & \new_[24226]_ ;
  assign \new_[24231]_  = \new_[24230]_  & \new_[24223]_ ;
  assign \new_[24235]_  = A167 & A169;
  assign \new_[24236]_  = ~A170 & \new_[24235]_ ;
  assign \new_[24239]_  = A199 & A166;
  assign \new_[24242]_  = A201 & ~A200;
  assign \new_[24243]_  = \new_[24242]_  & \new_[24239]_ ;
  assign \new_[24244]_  = \new_[24243]_  & \new_[24236]_ ;
  assign \new_[24248]_  = ~A266 & A265;
  assign \new_[24249]_  = A202 & \new_[24248]_ ;
  assign \new_[24252]_  = A268 & A267;
  assign \new_[24255]_  = ~A300 & A298;
  assign \new_[24256]_  = \new_[24255]_  & \new_[24252]_ ;
  assign \new_[24257]_  = \new_[24256]_  & \new_[24249]_ ;
  assign \new_[24261]_  = A167 & A169;
  assign \new_[24262]_  = ~A170 & \new_[24261]_ ;
  assign \new_[24265]_  = A199 & A166;
  assign \new_[24268]_  = A201 & ~A200;
  assign \new_[24269]_  = \new_[24268]_  & \new_[24265]_ ;
  assign \new_[24270]_  = \new_[24269]_  & \new_[24262]_ ;
  assign \new_[24274]_  = ~A266 & A265;
  assign \new_[24275]_  = A202 & \new_[24274]_ ;
  assign \new_[24278]_  = A268 & A267;
  assign \new_[24281]_  = A299 & A298;
  assign \new_[24282]_  = \new_[24281]_  & \new_[24278]_ ;
  assign \new_[24283]_  = \new_[24282]_  & \new_[24275]_ ;
  assign \new_[24287]_  = A167 & A169;
  assign \new_[24288]_  = ~A170 & \new_[24287]_ ;
  assign \new_[24291]_  = A199 & A166;
  assign \new_[24294]_  = A201 & ~A200;
  assign \new_[24295]_  = \new_[24294]_  & \new_[24291]_ ;
  assign \new_[24296]_  = \new_[24295]_  & \new_[24288]_ ;
  assign \new_[24300]_  = ~A266 & A265;
  assign \new_[24301]_  = A202 & \new_[24300]_ ;
  assign \new_[24304]_  = A268 & A267;
  assign \new_[24307]_  = ~A299 & ~A298;
  assign \new_[24308]_  = \new_[24307]_  & \new_[24304]_ ;
  assign \new_[24309]_  = \new_[24308]_  & \new_[24301]_ ;
  assign \new_[24313]_  = A167 & A169;
  assign \new_[24314]_  = ~A170 & \new_[24313]_ ;
  assign \new_[24317]_  = A199 & A166;
  assign \new_[24320]_  = A201 & ~A200;
  assign \new_[24321]_  = \new_[24320]_  & \new_[24317]_ ;
  assign \new_[24322]_  = \new_[24321]_  & \new_[24314]_ ;
  assign \new_[24326]_  = ~A266 & A265;
  assign \new_[24327]_  = A202 & \new_[24326]_ ;
  assign \new_[24330]_  = A269 & A267;
  assign \new_[24333]_  = ~A300 & A298;
  assign \new_[24334]_  = \new_[24333]_  & \new_[24330]_ ;
  assign \new_[24335]_  = \new_[24334]_  & \new_[24327]_ ;
  assign \new_[24339]_  = A167 & A169;
  assign \new_[24340]_  = ~A170 & \new_[24339]_ ;
  assign \new_[24343]_  = A199 & A166;
  assign \new_[24346]_  = A201 & ~A200;
  assign \new_[24347]_  = \new_[24346]_  & \new_[24343]_ ;
  assign \new_[24348]_  = \new_[24347]_  & \new_[24340]_ ;
  assign \new_[24352]_  = ~A266 & A265;
  assign \new_[24353]_  = A202 & \new_[24352]_ ;
  assign \new_[24356]_  = A269 & A267;
  assign \new_[24359]_  = A299 & A298;
  assign \new_[24360]_  = \new_[24359]_  & \new_[24356]_ ;
  assign \new_[24361]_  = \new_[24360]_  & \new_[24353]_ ;
  assign \new_[24365]_  = A167 & A169;
  assign \new_[24366]_  = ~A170 & \new_[24365]_ ;
  assign \new_[24369]_  = A199 & A166;
  assign \new_[24372]_  = A201 & ~A200;
  assign \new_[24373]_  = \new_[24372]_  & \new_[24369]_ ;
  assign \new_[24374]_  = \new_[24373]_  & \new_[24366]_ ;
  assign \new_[24378]_  = ~A266 & A265;
  assign \new_[24379]_  = A202 & \new_[24378]_ ;
  assign \new_[24382]_  = A269 & A267;
  assign \new_[24385]_  = ~A299 & ~A298;
  assign \new_[24386]_  = \new_[24385]_  & \new_[24382]_ ;
  assign \new_[24387]_  = \new_[24386]_  & \new_[24379]_ ;
  assign \new_[24391]_  = A167 & A169;
  assign \new_[24392]_  = ~A170 & \new_[24391]_ ;
  assign \new_[24395]_  = A199 & A166;
  assign \new_[24398]_  = A201 & ~A200;
  assign \new_[24399]_  = \new_[24398]_  & \new_[24395]_ ;
  assign \new_[24400]_  = \new_[24399]_  & \new_[24392]_ ;
  assign \new_[24404]_  = ~A266 & A265;
  assign \new_[24405]_  = A203 & \new_[24404]_ ;
  assign \new_[24408]_  = A268 & A267;
  assign \new_[24411]_  = ~A300 & A298;
  assign \new_[24412]_  = \new_[24411]_  & \new_[24408]_ ;
  assign \new_[24413]_  = \new_[24412]_  & \new_[24405]_ ;
  assign \new_[24417]_  = A167 & A169;
  assign \new_[24418]_  = ~A170 & \new_[24417]_ ;
  assign \new_[24421]_  = A199 & A166;
  assign \new_[24424]_  = A201 & ~A200;
  assign \new_[24425]_  = \new_[24424]_  & \new_[24421]_ ;
  assign \new_[24426]_  = \new_[24425]_  & \new_[24418]_ ;
  assign \new_[24430]_  = ~A266 & A265;
  assign \new_[24431]_  = A203 & \new_[24430]_ ;
  assign \new_[24434]_  = A268 & A267;
  assign \new_[24437]_  = A299 & A298;
  assign \new_[24438]_  = \new_[24437]_  & \new_[24434]_ ;
  assign \new_[24439]_  = \new_[24438]_  & \new_[24431]_ ;
  assign \new_[24443]_  = A167 & A169;
  assign \new_[24444]_  = ~A170 & \new_[24443]_ ;
  assign \new_[24447]_  = A199 & A166;
  assign \new_[24450]_  = A201 & ~A200;
  assign \new_[24451]_  = \new_[24450]_  & \new_[24447]_ ;
  assign \new_[24452]_  = \new_[24451]_  & \new_[24444]_ ;
  assign \new_[24456]_  = ~A266 & A265;
  assign \new_[24457]_  = A203 & \new_[24456]_ ;
  assign \new_[24460]_  = A268 & A267;
  assign \new_[24463]_  = ~A299 & ~A298;
  assign \new_[24464]_  = \new_[24463]_  & \new_[24460]_ ;
  assign \new_[24465]_  = \new_[24464]_  & \new_[24457]_ ;
  assign \new_[24469]_  = A167 & A169;
  assign \new_[24470]_  = ~A170 & \new_[24469]_ ;
  assign \new_[24473]_  = A199 & A166;
  assign \new_[24476]_  = A201 & ~A200;
  assign \new_[24477]_  = \new_[24476]_  & \new_[24473]_ ;
  assign \new_[24478]_  = \new_[24477]_  & \new_[24470]_ ;
  assign \new_[24482]_  = ~A266 & A265;
  assign \new_[24483]_  = A203 & \new_[24482]_ ;
  assign \new_[24486]_  = A269 & A267;
  assign \new_[24489]_  = ~A300 & A298;
  assign \new_[24490]_  = \new_[24489]_  & \new_[24486]_ ;
  assign \new_[24491]_  = \new_[24490]_  & \new_[24483]_ ;
  assign \new_[24495]_  = A167 & A169;
  assign \new_[24496]_  = ~A170 & \new_[24495]_ ;
  assign \new_[24499]_  = A199 & A166;
  assign \new_[24502]_  = A201 & ~A200;
  assign \new_[24503]_  = \new_[24502]_  & \new_[24499]_ ;
  assign \new_[24504]_  = \new_[24503]_  & \new_[24496]_ ;
  assign \new_[24508]_  = ~A266 & A265;
  assign \new_[24509]_  = A203 & \new_[24508]_ ;
  assign \new_[24512]_  = A269 & A267;
  assign \new_[24515]_  = A299 & A298;
  assign \new_[24516]_  = \new_[24515]_  & \new_[24512]_ ;
  assign \new_[24517]_  = \new_[24516]_  & \new_[24509]_ ;
  assign \new_[24521]_  = A167 & A169;
  assign \new_[24522]_  = ~A170 & \new_[24521]_ ;
  assign \new_[24525]_  = A199 & A166;
  assign \new_[24528]_  = A201 & ~A200;
  assign \new_[24529]_  = \new_[24528]_  & \new_[24525]_ ;
  assign \new_[24530]_  = \new_[24529]_  & \new_[24522]_ ;
  assign \new_[24534]_  = ~A266 & A265;
  assign \new_[24535]_  = A203 & \new_[24534]_ ;
  assign \new_[24538]_  = A269 & A267;
  assign \new_[24541]_  = ~A299 & ~A298;
  assign \new_[24542]_  = \new_[24541]_  & \new_[24538]_ ;
  assign \new_[24543]_  = \new_[24542]_  & \new_[24535]_ ;
  assign \new_[24547]_  = ~A167 & A169;
  assign \new_[24548]_  = ~A170 & \new_[24547]_ ;
  assign \new_[24551]_  = ~A200 & ~A166;
  assign \new_[24554]_  = ~A203 & ~A202;
  assign \new_[24555]_  = \new_[24554]_  & \new_[24551]_ ;
  assign \new_[24556]_  = \new_[24555]_  & \new_[24548]_ ;
  assign \new_[24560]_  = ~A269 & ~A268;
  assign \new_[24561]_  = ~A266 & \new_[24560]_ ;
  assign \new_[24564]_  = ~A299 & A298;
  assign \new_[24567]_  = A301 & A300;
  assign \new_[24568]_  = \new_[24567]_  & \new_[24564]_ ;
  assign \new_[24569]_  = \new_[24568]_  & \new_[24561]_ ;
  assign \new_[24573]_  = ~A167 & A169;
  assign \new_[24574]_  = ~A170 & \new_[24573]_ ;
  assign \new_[24577]_  = ~A200 & ~A166;
  assign \new_[24580]_  = ~A203 & ~A202;
  assign \new_[24581]_  = \new_[24580]_  & \new_[24577]_ ;
  assign \new_[24582]_  = \new_[24581]_  & \new_[24574]_ ;
  assign \new_[24586]_  = ~A269 & ~A268;
  assign \new_[24587]_  = ~A266 & \new_[24586]_ ;
  assign \new_[24590]_  = ~A299 & A298;
  assign \new_[24593]_  = A302 & A300;
  assign \new_[24594]_  = \new_[24593]_  & \new_[24590]_ ;
  assign \new_[24595]_  = \new_[24594]_  & \new_[24587]_ ;
  assign \new_[24599]_  = ~A167 & A169;
  assign \new_[24600]_  = ~A170 & \new_[24599]_ ;
  assign \new_[24603]_  = A199 & ~A166;
  assign \new_[24606]_  = A201 & ~A200;
  assign \new_[24607]_  = \new_[24606]_  & \new_[24603]_ ;
  assign \new_[24608]_  = \new_[24607]_  & \new_[24600]_ ;
  assign \new_[24612]_  = ~A266 & A265;
  assign \new_[24613]_  = A202 & \new_[24612]_ ;
  assign \new_[24616]_  = A268 & A267;
  assign \new_[24619]_  = ~A300 & A298;
  assign \new_[24620]_  = \new_[24619]_  & \new_[24616]_ ;
  assign \new_[24621]_  = \new_[24620]_  & \new_[24613]_ ;
  assign \new_[24625]_  = ~A167 & A169;
  assign \new_[24626]_  = ~A170 & \new_[24625]_ ;
  assign \new_[24629]_  = A199 & ~A166;
  assign \new_[24632]_  = A201 & ~A200;
  assign \new_[24633]_  = \new_[24632]_  & \new_[24629]_ ;
  assign \new_[24634]_  = \new_[24633]_  & \new_[24626]_ ;
  assign \new_[24638]_  = ~A266 & A265;
  assign \new_[24639]_  = A202 & \new_[24638]_ ;
  assign \new_[24642]_  = A268 & A267;
  assign \new_[24645]_  = A299 & A298;
  assign \new_[24646]_  = \new_[24645]_  & \new_[24642]_ ;
  assign \new_[24647]_  = \new_[24646]_  & \new_[24639]_ ;
  assign \new_[24651]_  = ~A167 & A169;
  assign \new_[24652]_  = ~A170 & \new_[24651]_ ;
  assign \new_[24655]_  = A199 & ~A166;
  assign \new_[24658]_  = A201 & ~A200;
  assign \new_[24659]_  = \new_[24658]_  & \new_[24655]_ ;
  assign \new_[24660]_  = \new_[24659]_  & \new_[24652]_ ;
  assign \new_[24664]_  = ~A266 & A265;
  assign \new_[24665]_  = A202 & \new_[24664]_ ;
  assign \new_[24668]_  = A268 & A267;
  assign \new_[24671]_  = ~A299 & ~A298;
  assign \new_[24672]_  = \new_[24671]_  & \new_[24668]_ ;
  assign \new_[24673]_  = \new_[24672]_  & \new_[24665]_ ;
  assign \new_[24677]_  = ~A167 & A169;
  assign \new_[24678]_  = ~A170 & \new_[24677]_ ;
  assign \new_[24681]_  = A199 & ~A166;
  assign \new_[24684]_  = A201 & ~A200;
  assign \new_[24685]_  = \new_[24684]_  & \new_[24681]_ ;
  assign \new_[24686]_  = \new_[24685]_  & \new_[24678]_ ;
  assign \new_[24690]_  = ~A266 & A265;
  assign \new_[24691]_  = A202 & \new_[24690]_ ;
  assign \new_[24694]_  = A269 & A267;
  assign \new_[24697]_  = ~A300 & A298;
  assign \new_[24698]_  = \new_[24697]_  & \new_[24694]_ ;
  assign \new_[24699]_  = \new_[24698]_  & \new_[24691]_ ;
  assign \new_[24703]_  = ~A167 & A169;
  assign \new_[24704]_  = ~A170 & \new_[24703]_ ;
  assign \new_[24707]_  = A199 & ~A166;
  assign \new_[24710]_  = A201 & ~A200;
  assign \new_[24711]_  = \new_[24710]_  & \new_[24707]_ ;
  assign \new_[24712]_  = \new_[24711]_  & \new_[24704]_ ;
  assign \new_[24716]_  = ~A266 & A265;
  assign \new_[24717]_  = A202 & \new_[24716]_ ;
  assign \new_[24720]_  = A269 & A267;
  assign \new_[24723]_  = A299 & A298;
  assign \new_[24724]_  = \new_[24723]_  & \new_[24720]_ ;
  assign \new_[24725]_  = \new_[24724]_  & \new_[24717]_ ;
  assign \new_[24729]_  = ~A167 & A169;
  assign \new_[24730]_  = ~A170 & \new_[24729]_ ;
  assign \new_[24733]_  = A199 & ~A166;
  assign \new_[24736]_  = A201 & ~A200;
  assign \new_[24737]_  = \new_[24736]_  & \new_[24733]_ ;
  assign \new_[24738]_  = \new_[24737]_  & \new_[24730]_ ;
  assign \new_[24742]_  = ~A266 & A265;
  assign \new_[24743]_  = A202 & \new_[24742]_ ;
  assign \new_[24746]_  = A269 & A267;
  assign \new_[24749]_  = ~A299 & ~A298;
  assign \new_[24750]_  = \new_[24749]_  & \new_[24746]_ ;
  assign \new_[24751]_  = \new_[24750]_  & \new_[24743]_ ;
  assign \new_[24755]_  = ~A167 & A169;
  assign \new_[24756]_  = ~A170 & \new_[24755]_ ;
  assign \new_[24759]_  = A199 & ~A166;
  assign \new_[24762]_  = A201 & ~A200;
  assign \new_[24763]_  = \new_[24762]_  & \new_[24759]_ ;
  assign \new_[24764]_  = \new_[24763]_  & \new_[24756]_ ;
  assign \new_[24768]_  = ~A266 & A265;
  assign \new_[24769]_  = A203 & \new_[24768]_ ;
  assign \new_[24772]_  = A268 & A267;
  assign \new_[24775]_  = ~A300 & A298;
  assign \new_[24776]_  = \new_[24775]_  & \new_[24772]_ ;
  assign \new_[24777]_  = \new_[24776]_  & \new_[24769]_ ;
  assign \new_[24781]_  = ~A167 & A169;
  assign \new_[24782]_  = ~A170 & \new_[24781]_ ;
  assign \new_[24785]_  = A199 & ~A166;
  assign \new_[24788]_  = A201 & ~A200;
  assign \new_[24789]_  = \new_[24788]_  & \new_[24785]_ ;
  assign \new_[24790]_  = \new_[24789]_  & \new_[24782]_ ;
  assign \new_[24794]_  = ~A266 & A265;
  assign \new_[24795]_  = A203 & \new_[24794]_ ;
  assign \new_[24798]_  = A268 & A267;
  assign \new_[24801]_  = A299 & A298;
  assign \new_[24802]_  = \new_[24801]_  & \new_[24798]_ ;
  assign \new_[24803]_  = \new_[24802]_  & \new_[24795]_ ;
  assign \new_[24807]_  = ~A167 & A169;
  assign \new_[24808]_  = ~A170 & \new_[24807]_ ;
  assign \new_[24811]_  = A199 & ~A166;
  assign \new_[24814]_  = A201 & ~A200;
  assign \new_[24815]_  = \new_[24814]_  & \new_[24811]_ ;
  assign \new_[24816]_  = \new_[24815]_  & \new_[24808]_ ;
  assign \new_[24820]_  = ~A266 & A265;
  assign \new_[24821]_  = A203 & \new_[24820]_ ;
  assign \new_[24824]_  = A268 & A267;
  assign \new_[24827]_  = ~A299 & ~A298;
  assign \new_[24828]_  = \new_[24827]_  & \new_[24824]_ ;
  assign \new_[24829]_  = \new_[24828]_  & \new_[24821]_ ;
  assign \new_[24833]_  = ~A167 & A169;
  assign \new_[24834]_  = ~A170 & \new_[24833]_ ;
  assign \new_[24837]_  = A199 & ~A166;
  assign \new_[24840]_  = A201 & ~A200;
  assign \new_[24841]_  = \new_[24840]_  & \new_[24837]_ ;
  assign \new_[24842]_  = \new_[24841]_  & \new_[24834]_ ;
  assign \new_[24846]_  = ~A266 & A265;
  assign \new_[24847]_  = A203 & \new_[24846]_ ;
  assign \new_[24850]_  = A269 & A267;
  assign \new_[24853]_  = ~A300 & A298;
  assign \new_[24854]_  = \new_[24853]_  & \new_[24850]_ ;
  assign \new_[24855]_  = \new_[24854]_  & \new_[24847]_ ;
  assign \new_[24859]_  = ~A167 & A169;
  assign \new_[24860]_  = ~A170 & \new_[24859]_ ;
  assign \new_[24863]_  = A199 & ~A166;
  assign \new_[24866]_  = A201 & ~A200;
  assign \new_[24867]_  = \new_[24866]_  & \new_[24863]_ ;
  assign \new_[24868]_  = \new_[24867]_  & \new_[24860]_ ;
  assign \new_[24872]_  = ~A266 & A265;
  assign \new_[24873]_  = A203 & \new_[24872]_ ;
  assign \new_[24876]_  = A269 & A267;
  assign \new_[24879]_  = A299 & A298;
  assign \new_[24880]_  = \new_[24879]_  & \new_[24876]_ ;
  assign \new_[24881]_  = \new_[24880]_  & \new_[24873]_ ;
  assign \new_[24885]_  = ~A167 & A169;
  assign \new_[24886]_  = ~A170 & \new_[24885]_ ;
  assign \new_[24889]_  = A199 & ~A166;
  assign \new_[24892]_  = A201 & ~A200;
  assign \new_[24893]_  = \new_[24892]_  & \new_[24889]_ ;
  assign \new_[24894]_  = \new_[24893]_  & \new_[24886]_ ;
  assign \new_[24898]_  = ~A266 & A265;
  assign \new_[24899]_  = A203 & \new_[24898]_ ;
  assign \new_[24902]_  = A269 & A267;
  assign \new_[24905]_  = ~A299 & ~A298;
  assign \new_[24906]_  = \new_[24905]_  & \new_[24902]_ ;
  assign \new_[24907]_  = \new_[24906]_  & \new_[24899]_ ;
  assign \new_[24911]_  = ~A166 & ~A167;
  assign \new_[24912]_  = ~A169 & \new_[24911]_ ;
  assign \new_[24915]_  = ~A200 & A199;
  assign \new_[24918]_  = A202 & A201;
  assign \new_[24919]_  = \new_[24918]_  & \new_[24915]_ ;
  assign \new_[24920]_  = \new_[24919]_  & \new_[24912]_ ;
  assign \new_[24924]_  = ~A269 & ~A268;
  assign \new_[24925]_  = ~A266 & \new_[24924]_ ;
  assign \new_[24928]_  = ~A299 & A298;
  assign \new_[24931]_  = A301 & A300;
  assign \new_[24932]_  = \new_[24931]_  & \new_[24928]_ ;
  assign \new_[24933]_  = \new_[24932]_  & \new_[24925]_ ;
  assign \new_[24937]_  = ~A166 & ~A167;
  assign \new_[24938]_  = ~A169 & \new_[24937]_ ;
  assign \new_[24941]_  = ~A200 & A199;
  assign \new_[24944]_  = A202 & A201;
  assign \new_[24945]_  = \new_[24944]_  & \new_[24941]_ ;
  assign \new_[24946]_  = \new_[24945]_  & \new_[24938]_ ;
  assign \new_[24950]_  = ~A269 & ~A268;
  assign \new_[24951]_  = ~A266 & \new_[24950]_ ;
  assign \new_[24954]_  = ~A299 & A298;
  assign \new_[24957]_  = A302 & A300;
  assign \new_[24958]_  = \new_[24957]_  & \new_[24954]_ ;
  assign \new_[24959]_  = \new_[24958]_  & \new_[24951]_ ;
  assign \new_[24963]_  = ~A166 & ~A167;
  assign \new_[24964]_  = ~A169 & \new_[24963]_ ;
  assign \new_[24967]_  = ~A200 & A199;
  assign \new_[24970]_  = A203 & A201;
  assign \new_[24971]_  = \new_[24970]_  & \new_[24967]_ ;
  assign \new_[24972]_  = \new_[24971]_  & \new_[24964]_ ;
  assign \new_[24976]_  = ~A269 & ~A268;
  assign \new_[24977]_  = ~A266 & \new_[24976]_ ;
  assign \new_[24980]_  = ~A299 & A298;
  assign \new_[24983]_  = A301 & A300;
  assign \new_[24984]_  = \new_[24983]_  & \new_[24980]_ ;
  assign \new_[24985]_  = \new_[24984]_  & \new_[24977]_ ;
  assign \new_[24989]_  = ~A166 & ~A167;
  assign \new_[24990]_  = ~A169 & \new_[24989]_ ;
  assign \new_[24993]_  = ~A200 & A199;
  assign \new_[24996]_  = A203 & A201;
  assign \new_[24997]_  = \new_[24996]_  & \new_[24993]_ ;
  assign \new_[24998]_  = \new_[24997]_  & \new_[24990]_ ;
  assign \new_[25002]_  = ~A269 & ~A268;
  assign \new_[25003]_  = ~A266 & \new_[25002]_ ;
  assign \new_[25006]_  = ~A299 & A298;
  assign \new_[25009]_  = A302 & A300;
  assign \new_[25010]_  = \new_[25009]_  & \new_[25006]_ ;
  assign \new_[25011]_  = \new_[25010]_  & \new_[25003]_ ;
  assign \new_[25015]_  = A167 & ~A168;
  assign \new_[25016]_  = ~A169 & \new_[25015]_ ;
  assign \new_[25019]_  = ~A200 & A166;
  assign \new_[25022]_  = ~A203 & ~A202;
  assign \new_[25023]_  = \new_[25022]_  & \new_[25019]_ ;
  assign \new_[25024]_  = \new_[25023]_  & \new_[25016]_ ;
  assign \new_[25028]_  = A267 & ~A266;
  assign \new_[25029]_  = A265 & \new_[25028]_ ;
  assign \new_[25032]_  = A298 & A268;
  assign \new_[25035]_  = ~A302 & ~A301;
  assign \new_[25036]_  = \new_[25035]_  & \new_[25032]_ ;
  assign \new_[25037]_  = \new_[25036]_  & \new_[25029]_ ;
  assign \new_[25041]_  = A167 & ~A168;
  assign \new_[25042]_  = ~A169 & \new_[25041]_ ;
  assign \new_[25045]_  = ~A200 & A166;
  assign \new_[25048]_  = ~A203 & ~A202;
  assign \new_[25049]_  = \new_[25048]_  & \new_[25045]_ ;
  assign \new_[25050]_  = \new_[25049]_  & \new_[25042]_ ;
  assign \new_[25054]_  = A267 & ~A266;
  assign \new_[25055]_  = A265 & \new_[25054]_ ;
  assign \new_[25058]_  = A298 & A269;
  assign \new_[25061]_  = ~A302 & ~A301;
  assign \new_[25062]_  = \new_[25061]_  & \new_[25058]_ ;
  assign \new_[25063]_  = \new_[25062]_  & \new_[25055]_ ;
  assign \new_[25067]_  = A167 & ~A168;
  assign \new_[25068]_  = ~A169 & \new_[25067]_ ;
  assign \new_[25071]_  = A199 & A166;
  assign \new_[25074]_  = A201 & ~A200;
  assign \new_[25075]_  = \new_[25074]_  & \new_[25071]_ ;
  assign \new_[25076]_  = \new_[25075]_  & \new_[25068]_ ;
  assign \new_[25080]_  = A266 & A265;
  assign \new_[25081]_  = A202 & \new_[25080]_ ;
  assign \new_[25084]_  = ~A299 & A298;
  assign \new_[25087]_  = A301 & A300;
  assign \new_[25088]_  = \new_[25087]_  & \new_[25084]_ ;
  assign \new_[25089]_  = \new_[25088]_  & \new_[25081]_ ;
  assign \new_[25093]_  = A167 & ~A168;
  assign \new_[25094]_  = ~A169 & \new_[25093]_ ;
  assign \new_[25097]_  = A199 & A166;
  assign \new_[25100]_  = A201 & ~A200;
  assign \new_[25101]_  = \new_[25100]_  & \new_[25097]_ ;
  assign \new_[25102]_  = \new_[25101]_  & \new_[25094]_ ;
  assign \new_[25106]_  = A266 & A265;
  assign \new_[25107]_  = A202 & \new_[25106]_ ;
  assign \new_[25110]_  = ~A299 & A298;
  assign \new_[25113]_  = A302 & A300;
  assign \new_[25114]_  = \new_[25113]_  & \new_[25110]_ ;
  assign \new_[25115]_  = \new_[25114]_  & \new_[25107]_ ;
  assign \new_[25119]_  = A167 & ~A168;
  assign \new_[25120]_  = ~A169 & \new_[25119]_ ;
  assign \new_[25123]_  = A199 & A166;
  assign \new_[25126]_  = A201 & ~A200;
  assign \new_[25127]_  = \new_[25126]_  & \new_[25123]_ ;
  assign \new_[25128]_  = \new_[25127]_  & \new_[25120]_ ;
  assign \new_[25132]_  = ~A267 & ~A266;
  assign \new_[25133]_  = A202 & \new_[25132]_ ;
  assign \new_[25136]_  = ~A299 & A298;
  assign \new_[25139]_  = A301 & A300;
  assign \new_[25140]_  = \new_[25139]_  & \new_[25136]_ ;
  assign \new_[25141]_  = \new_[25140]_  & \new_[25133]_ ;
  assign \new_[25145]_  = A167 & ~A168;
  assign \new_[25146]_  = ~A169 & \new_[25145]_ ;
  assign \new_[25149]_  = A199 & A166;
  assign \new_[25152]_  = A201 & ~A200;
  assign \new_[25153]_  = \new_[25152]_  & \new_[25149]_ ;
  assign \new_[25154]_  = \new_[25153]_  & \new_[25146]_ ;
  assign \new_[25158]_  = ~A267 & ~A266;
  assign \new_[25159]_  = A202 & \new_[25158]_ ;
  assign \new_[25162]_  = ~A299 & A298;
  assign \new_[25165]_  = A302 & A300;
  assign \new_[25166]_  = \new_[25165]_  & \new_[25162]_ ;
  assign \new_[25167]_  = \new_[25166]_  & \new_[25159]_ ;
  assign \new_[25171]_  = A167 & ~A168;
  assign \new_[25172]_  = ~A169 & \new_[25171]_ ;
  assign \new_[25175]_  = A199 & A166;
  assign \new_[25178]_  = A201 & ~A200;
  assign \new_[25179]_  = \new_[25178]_  & \new_[25175]_ ;
  assign \new_[25180]_  = \new_[25179]_  & \new_[25172]_ ;
  assign \new_[25184]_  = ~A266 & ~A265;
  assign \new_[25185]_  = A202 & \new_[25184]_ ;
  assign \new_[25188]_  = ~A299 & A298;
  assign \new_[25191]_  = A301 & A300;
  assign \new_[25192]_  = \new_[25191]_  & \new_[25188]_ ;
  assign \new_[25193]_  = \new_[25192]_  & \new_[25185]_ ;
  assign \new_[25197]_  = A167 & ~A168;
  assign \new_[25198]_  = ~A169 & \new_[25197]_ ;
  assign \new_[25201]_  = A199 & A166;
  assign \new_[25204]_  = A201 & ~A200;
  assign \new_[25205]_  = \new_[25204]_  & \new_[25201]_ ;
  assign \new_[25206]_  = \new_[25205]_  & \new_[25198]_ ;
  assign \new_[25210]_  = ~A266 & ~A265;
  assign \new_[25211]_  = A202 & \new_[25210]_ ;
  assign \new_[25214]_  = ~A299 & A298;
  assign \new_[25217]_  = A302 & A300;
  assign \new_[25218]_  = \new_[25217]_  & \new_[25214]_ ;
  assign \new_[25219]_  = \new_[25218]_  & \new_[25211]_ ;
  assign \new_[25223]_  = A167 & ~A168;
  assign \new_[25224]_  = ~A169 & \new_[25223]_ ;
  assign \new_[25227]_  = A199 & A166;
  assign \new_[25230]_  = A201 & ~A200;
  assign \new_[25231]_  = \new_[25230]_  & \new_[25227]_ ;
  assign \new_[25232]_  = \new_[25231]_  & \new_[25224]_ ;
  assign \new_[25236]_  = A266 & A265;
  assign \new_[25237]_  = A203 & \new_[25236]_ ;
  assign \new_[25240]_  = ~A299 & A298;
  assign \new_[25243]_  = A301 & A300;
  assign \new_[25244]_  = \new_[25243]_  & \new_[25240]_ ;
  assign \new_[25245]_  = \new_[25244]_  & \new_[25237]_ ;
  assign \new_[25249]_  = A167 & ~A168;
  assign \new_[25250]_  = ~A169 & \new_[25249]_ ;
  assign \new_[25253]_  = A199 & A166;
  assign \new_[25256]_  = A201 & ~A200;
  assign \new_[25257]_  = \new_[25256]_  & \new_[25253]_ ;
  assign \new_[25258]_  = \new_[25257]_  & \new_[25250]_ ;
  assign \new_[25262]_  = A266 & A265;
  assign \new_[25263]_  = A203 & \new_[25262]_ ;
  assign \new_[25266]_  = ~A299 & A298;
  assign \new_[25269]_  = A302 & A300;
  assign \new_[25270]_  = \new_[25269]_  & \new_[25266]_ ;
  assign \new_[25271]_  = \new_[25270]_  & \new_[25263]_ ;
  assign \new_[25275]_  = A167 & ~A168;
  assign \new_[25276]_  = ~A169 & \new_[25275]_ ;
  assign \new_[25279]_  = A199 & A166;
  assign \new_[25282]_  = A201 & ~A200;
  assign \new_[25283]_  = \new_[25282]_  & \new_[25279]_ ;
  assign \new_[25284]_  = \new_[25283]_  & \new_[25276]_ ;
  assign \new_[25288]_  = ~A267 & ~A266;
  assign \new_[25289]_  = A203 & \new_[25288]_ ;
  assign \new_[25292]_  = ~A299 & A298;
  assign \new_[25295]_  = A301 & A300;
  assign \new_[25296]_  = \new_[25295]_  & \new_[25292]_ ;
  assign \new_[25297]_  = \new_[25296]_  & \new_[25289]_ ;
  assign \new_[25301]_  = A167 & ~A168;
  assign \new_[25302]_  = ~A169 & \new_[25301]_ ;
  assign \new_[25305]_  = A199 & A166;
  assign \new_[25308]_  = A201 & ~A200;
  assign \new_[25309]_  = \new_[25308]_  & \new_[25305]_ ;
  assign \new_[25310]_  = \new_[25309]_  & \new_[25302]_ ;
  assign \new_[25314]_  = ~A267 & ~A266;
  assign \new_[25315]_  = A203 & \new_[25314]_ ;
  assign \new_[25318]_  = ~A299 & A298;
  assign \new_[25321]_  = A302 & A300;
  assign \new_[25322]_  = \new_[25321]_  & \new_[25318]_ ;
  assign \new_[25323]_  = \new_[25322]_  & \new_[25315]_ ;
  assign \new_[25327]_  = A167 & ~A168;
  assign \new_[25328]_  = ~A169 & \new_[25327]_ ;
  assign \new_[25331]_  = A199 & A166;
  assign \new_[25334]_  = A201 & ~A200;
  assign \new_[25335]_  = \new_[25334]_  & \new_[25331]_ ;
  assign \new_[25336]_  = \new_[25335]_  & \new_[25328]_ ;
  assign \new_[25340]_  = ~A266 & ~A265;
  assign \new_[25341]_  = A203 & \new_[25340]_ ;
  assign \new_[25344]_  = ~A299 & A298;
  assign \new_[25347]_  = A301 & A300;
  assign \new_[25348]_  = \new_[25347]_  & \new_[25344]_ ;
  assign \new_[25349]_  = \new_[25348]_  & \new_[25341]_ ;
  assign \new_[25353]_  = A167 & ~A168;
  assign \new_[25354]_  = ~A169 & \new_[25353]_ ;
  assign \new_[25357]_  = A199 & A166;
  assign \new_[25360]_  = A201 & ~A200;
  assign \new_[25361]_  = \new_[25360]_  & \new_[25357]_ ;
  assign \new_[25362]_  = \new_[25361]_  & \new_[25354]_ ;
  assign \new_[25366]_  = ~A266 & ~A265;
  assign \new_[25367]_  = A203 & \new_[25366]_ ;
  assign \new_[25370]_  = ~A299 & A298;
  assign \new_[25373]_  = A302 & A300;
  assign \new_[25374]_  = \new_[25373]_  & \new_[25370]_ ;
  assign \new_[25375]_  = \new_[25374]_  & \new_[25367]_ ;
  assign \new_[25379]_  = A167 & ~A169;
  assign \new_[25380]_  = A170 & \new_[25379]_ ;
  assign \new_[25383]_  = ~A200 & ~A166;
  assign \new_[25386]_  = ~A203 & ~A202;
  assign \new_[25387]_  = \new_[25386]_  & \new_[25383]_ ;
  assign \new_[25388]_  = \new_[25387]_  & \new_[25380]_ ;
  assign \new_[25392]_  = ~A269 & ~A268;
  assign \new_[25393]_  = ~A266 & \new_[25392]_ ;
  assign \new_[25396]_  = ~A299 & A298;
  assign \new_[25399]_  = A301 & A300;
  assign \new_[25400]_  = \new_[25399]_  & \new_[25396]_ ;
  assign \new_[25401]_  = \new_[25400]_  & \new_[25393]_ ;
  assign \new_[25405]_  = A167 & ~A169;
  assign \new_[25406]_  = A170 & \new_[25405]_ ;
  assign \new_[25409]_  = ~A200 & ~A166;
  assign \new_[25412]_  = ~A203 & ~A202;
  assign \new_[25413]_  = \new_[25412]_  & \new_[25409]_ ;
  assign \new_[25414]_  = \new_[25413]_  & \new_[25406]_ ;
  assign \new_[25418]_  = ~A269 & ~A268;
  assign \new_[25419]_  = ~A266 & \new_[25418]_ ;
  assign \new_[25422]_  = ~A299 & A298;
  assign \new_[25425]_  = A302 & A300;
  assign \new_[25426]_  = \new_[25425]_  & \new_[25422]_ ;
  assign \new_[25427]_  = \new_[25426]_  & \new_[25419]_ ;
  assign \new_[25431]_  = A167 & ~A169;
  assign \new_[25432]_  = A170 & \new_[25431]_ ;
  assign \new_[25435]_  = A199 & ~A166;
  assign \new_[25438]_  = A201 & ~A200;
  assign \new_[25439]_  = \new_[25438]_  & \new_[25435]_ ;
  assign \new_[25440]_  = \new_[25439]_  & \new_[25432]_ ;
  assign \new_[25444]_  = ~A266 & A265;
  assign \new_[25445]_  = A202 & \new_[25444]_ ;
  assign \new_[25448]_  = A268 & A267;
  assign \new_[25451]_  = ~A300 & A298;
  assign \new_[25452]_  = \new_[25451]_  & \new_[25448]_ ;
  assign \new_[25453]_  = \new_[25452]_  & \new_[25445]_ ;
  assign \new_[25457]_  = A167 & ~A169;
  assign \new_[25458]_  = A170 & \new_[25457]_ ;
  assign \new_[25461]_  = A199 & ~A166;
  assign \new_[25464]_  = A201 & ~A200;
  assign \new_[25465]_  = \new_[25464]_  & \new_[25461]_ ;
  assign \new_[25466]_  = \new_[25465]_  & \new_[25458]_ ;
  assign \new_[25470]_  = ~A266 & A265;
  assign \new_[25471]_  = A202 & \new_[25470]_ ;
  assign \new_[25474]_  = A268 & A267;
  assign \new_[25477]_  = A299 & A298;
  assign \new_[25478]_  = \new_[25477]_  & \new_[25474]_ ;
  assign \new_[25479]_  = \new_[25478]_  & \new_[25471]_ ;
  assign \new_[25483]_  = A167 & ~A169;
  assign \new_[25484]_  = A170 & \new_[25483]_ ;
  assign \new_[25487]_  = A199 & ~A166;
  assign \new_[25490]_  = A201 & ~A200;
  assign \new_[25491]_  = \new_[25490]_  & \new_[25487]_ ;
  assign \new_[25492]_  = \new_[25491]_  & \new_[25484]_ ;
  assign \new_[25496]_  = ~A266 & A265;
  assign \new_[25497]_  = A202 & \new_[25496]_ ;
  assign \new_[25500]_  = A268 & A267;
  assign \new_[25503]_  = ~A299 & ~A298;
  assign \new_[25504]_  = \new_[25503]_  & \new_[25500]_ ;
  assign \new_[25505]_  = \new_[25504]_  & \new_[25497]_ ;
  assign \new_[25509]_  = A167 & ~A169;
  assign \new_[25510]_  = A170 & \new_[25509]_ ;
  assign \new_[25513]_  = A199 & ~A166;
  assign \new_[25516]_  = A201 & ~A200;
  assign \new_[25517]_  = \new_[25516]_  & \new_[25513]_ ;
  assign \new_[25518]_  = \new_[25517]_  & \new_[25510]_ ;
  assign \new_[25522]_  = ~A266 & A265;
  assign \new_[25523]_  = A202 & \new_[25522]_ ;
  assign \new_[25526]_  = A269 & A267;
  assign \new_[25529]_  = ~A300 & A298;
  assign \new_[25530]_  = \new_[25529]_  & \new_[25526]_ ;
  assign \new_[25531]_  = \new_[25530]_  & \new_[25523]_ ;
  assign \new_[25535]_  = A167 & ~A169;
  assign \new_[25536]_  = A170 & \new_[25535]_ ;
  assign \new_[25539]_  = A199 & ~A166;
  assign \new_[25542]_  = A201 & ~A200;
  assign \new_[25543]_  = \new_[25542]_  & \new_[25539]_ ;
  assign \new_[25544]_  = \new_[25543]_  & \new_[25536]_ ;
  assign \new_[25548]_  = ~A266 & A265;
  assign \new_[25549]_  = A202 & \new_[25548]_ ;
  assign \new_[25552]_  = A269 & A267;
  assign \new_[25555]_  = A299 & A298;
  assign \new_[25556]_  = \new_[25555]_  & \new_[25552]_ ;
  assign \new_[25557]_  = \new_[25556]_  & \new_[25549]_ ;
  assign \new_[25561]_  = A167 & ~A169;
  assign \new_[25562]_  = A170 & \new_[25561]_ ;
  assign \new_[25565]_  = A199 & ~A166;
  assign \new_[25568]_  = A201 & ~A200;
  assign \new_[25569]_  = \new_[25568]_  & \new_[25565]_ ;
  assign \new_[25570]_  = \new_[25569]_  & \new_[25562]_ ;
  assign \new_[25574]_  = ~A266 & A265;
  assign \new_[25575]_  = A202 & \new_[25574]_ ;
  assign \new_[25578]_  = A269 & A267;
  assign \new_[25581]_  = ~A299 & ~A298;
  assign \new_[25582]_  = \new_[25581]_  & \new_[25578]_ ;
  assign \new_[25583]_  = \new_[25582]_  & \new_[25575]_ ;
  assign \new_[25587]_  = A167 & ~A169;
  assign \new_[25588]_  = A170 & \new_[25587]_ ;
  assign \new_[25591]_  = A199 & ~A166;
  assign \new_[25594]_  = A201 & ~A200;
  assign \new_[25595]_  = \new_[25594]_  & \new_[25591]_ ;
  assign \new_[25596]_  = \new_[25595]_  & \new_[25588]_ ;
  assign \new_[25600]_  = ~A266 & A265;
  assign \new_[25601]_  = A203 & \new_[25600]_ ;
  assign \new_[25604]_  = A268 & A267;
  assign \new_[25607]_  = ~A300 & A298;
  assign \new_[25608]_  = \new_[25607]_  & \new_[25604]_ ;
  assign \new_[25609]_  = \new_[25608]_  & \new_[25601]_ ;
  assign \new_[25613]_  = A167 & ~A169;
  assign \new_[25614]_  = A170 & \new_[25613]_ ;
  assign \new_[25617]_  = A199 & ~A166;
  assign \new_[25620]_  = A201 & ~A200;
  assign \new_[25621]_  = \new_[25620]_  & \new_[25617]_ ;
  assign \new_[25622]_  = \new_[25621]_  & \new_[25614]_ ;
  assign \new_[25626]_  = ~A266 & A265;
  assign \new_[25627]_  = A203 & \new_[25626]_ ;
  assign \new_[25630]_  = A268 & A267;
  assign \new_[25633]_  = A299 & A298;
  assign \new_[25634]_  = \new_[25633]_  & \new_[25630]_ ;
  assign \new_[25635]_  = \new_[25634]_  & \new_[25627]_ ;
  assign \new_[25639]_  = A167 & ~A169;
  assign \new_[25640]_  = A170 & \new_[25639]_ ;
  assign \new_[25643]_  = A199 & ~A166;
  assign \new_[25646]_  = A201 & ~A200;
  assign \new_[25647]_  = \new_[25646]_  & \new_[25643]_ ;
  assign \new_[25648]_  = \new_[25647]_  & \new_[25640]_ ;
  assign \new_[25652]_  = ~A266 & A265;
  assign \new_[25653]_  = A203 & \new_[25652]_ ;
  assign \new_[25656]_  = A268 & A267;
  assign \new_[25659]_  = ~A299 & ~A298;
  assign \new_[25660]_  = \new_[25659]_  & \new_[25656]_ ;
  assign \new_[25661]_  = \new_[25660]_  & \new_[25653]_ ;
  assign \new_[25665]_  = A167 & ~A169;
  assign \new_[25666]_  = A170 & \new_[25665]_ ;
  assign \new_[25669]_  = A199 & ~A166;
  assign \new_[25672]_  = A201 & ~A200;
  assign \new_[25673]_  = \new_[25672]_  & \new_[25669]_ ;
  assign \new_[25674]_  = \new_[25673]_  & \new_[25666]_ ;
  assign \new_[25678]_  = ~A266 & A265;
  assign \new_[25679]_  = A203 & \new_[25678]_ ;
  assign \new_[25682]_  = A269 & A267;
  assign \new_[25685]_  = ~A300 & A298;
  assign \new_[25686]_  = \new_[25685]_  & \new_[25682]_ ;
  assign \new_[25687]_  = \new_[25686]_  & \new_[25679]_ ;
  assign \new_[25691]_  = A167 & ~A169;
  assign \new_[25692]_  = A170 & \new_[25691]_ ;
  assign \new_[25695]_  = A199 & ~A166;
  assign \new_[25698]_  = A201 & ~A200;
  assign \new_[25699]_  = \new_[25698]_  & \new_[25695]_ ;
  assign \new_[25700]_  = \new_[25699]_  & \new_[25692]_ ;
  assign \new_[25704]_  = ~A266 & A265;
  assign \new_[25705]_  = A203 & \new_[25704]_ ;
  assign \new_[25708]_  = A269 & A267;
  assign \new_[25711]_  = A299 & A298;
  assign \new_[25712]_  = \new_[25711]_  & \new_[25708]_ ;
  assign \new_[25713]_  = \new_[25712]_  & \new_[25705]_ ;
  assign \new_[25717]_  = A167 & ~A169;
  assign \new_[25718]_  = A170 & \new_[25717]_ ;
  assign \new_[25721]_  = A199 & ~A166;
  assign \new_[25724]_  = A201 & ~A200;
  assign \new_[25725]_  = \new_[25724]_  & \new_[25721]_ ;
  assign \new_[25726]_  = \new_[25725]_  & \new_[25718]_ ;
  assign \new_[25730]_  = ~A266 & A265;
  assign \new_[25731]_  = A203 & \new_[25730]_ ;
  assign \new_[25734]_  = A269 & A267;
  assign \new_[25737]_  = ~A299 & ~A298;
  assign \new_[25738]_  = \new_[25737]_  & \new_[25734]_ ;
  assign \new_[25739]_  = \new_[25738]_  & \new_[25731]_ ;
  assign \new_[25743]_  = ~A167 & ~A169;
  assign \new_[25744]_  = A170 & \new_[25743]_ ;
  assign \new_[25747]_  = ~A200 & A166;
  assign \new_[25750]_  = ~A203 & ~A202;
  assign \new_[25751]_  = \new_[25750]_  & \new_[25747]_ ;
  assign \new_[25752]_  = \new_[25751]_  & \new_[25744]_ ;
  assign \new_[25756]_  = ~A269 & ~A268;
  assign \new_[25757]_  = ~A266 & \new_[25756]_ ;
  assign \new_[25760]_  = ~A299 & A298;
  assign \new_[25763]_  = A301 & A300;
  assign \new_[25764]_  = \new_[25763]_  & \new_[25760]_ ;
  assign \new_[25765]_  = \new_[25764]_  & \new_[25757]_ ;
  assign \new_[25769]_  = ~A167 & ~A169;
  assign \new_[25770]_  = A170 & \new_[25769]_ ;
  assign \new_[25773]_  = ~A200 & A166;
  assign \new_[25776]_  = ~A203 & ~A202;
  assign \new_[25777]_  = \new_[25776]_  & \new_[25773]_ ;
  assign \new_[25778]_  = \new_[25777]_  & \new_[25770]_ ;
  assign \new_[25782]_  = ~A269 & ~A268;
  assign \new_[25783]_  = ~A266 & \new_[25782]_ ;
  assign \new_[25786]_  = ~A299 & A298;
  assign \new_[25789]_  = A302 & A300;
  assign \new_[25790]_  = \new_[25789]_  & \new_[25786]_ ;
  assign \new_[25791]_  = \new_[25790]_  & \new_[25783]_ ;
  assign \new_[25795]_  = ~A167 & ~A169;
  assign \new_[25796]_  = A170 & \new_[25795]_ ;
  assign \new_[25799]_  = A199 & A166;
  assign \new_[25802]_  = A201 & ~A200;
  assign \new_[25803]_  = \new_[25802]_  & \new_[25799]_ ;
  assign \new_[25804]_  = \new_[25803]_  & \new_[25796]_ ;
  assign \new_[25808]_  = ~A266 & A265;
  assign \new_[25809]_  = A202 & \new_[25808]_ ;
  assign \new_[25812]_  = A268 & A267;
  assign \new_[25815]_  = ~A300 & A298;
  assign \new_[25816]_  = \new_[25815]_  & \new_[25812]_ ;
  assign \new_[25817]_  = \new_[25816]_  & \new_[25809]_ ;
  assign \new_[25821]_  = ~A167 & ~A169;
  assign \new_[25822]_  = A170 & \new_[25821]_ ;
  assign \new_[25825]_  = A199 & A166;
  assign \new_[25828]_  = A201 & ~A200;
  assign \new_[25829]_  = \new_[25828]_  & \new_[25825]_ ;
  assign \new_[25830]_  = \new_[25829]_  & \new_[25822]_ ;
  assign \new_[25834]_  = ~A266 & A265;
  assign \new_[25835]_  = A202 & \new_[25834]_ ;
  assign \new_[25838]_  = A268 & A267;
  assign \new_[25841]_  = A299 & A298;
  assign \new_[25842]_  = \new_[25841]_  & \new_[25838]_ ;
  assign \new_[25843]_  = \new_[25842]_  & \new_[25835]_ ;
  assign \new_[25847]_  = ~A167 & ~A169;
  assign \new_[25848]_  = A170 & \new_[25847]_ ;
  assign \new_[25851]_  = A199 & A166;
  assign \new_[25854]_  = A201 & ~A200;
  assign \new_[25855]_  = \new_[25854]_  & \new_[25851]_ ;
  assign \new_[25856]_  = \new_[25855]_  & \new_[25848]_ ;
  assign \new_[25860]_  = ~A266 & A265;
  assign \new_[25861]_  = A202 & \new_[25860]_ ;
  assign \new_[25864]_  = A268 & A267;
  assign \new_[25867]_  = ~A299 & ~A298;
  assign \new_[25868]_  = \new_[25867]_  & \new_[25864]_ ;
  assign \new_[25869]_  = \new_[25868]_  & \new_[25861]_ ;
  assign \new_[25873]_  = ~A167 & ~A169;
  assign \new_[25874]_  = A170 & \new_[25873]_ ;
  assign \new_[25877]_  = A199 & A166;
  assign \new_[25880]_  = A201 & ~A200;
  assign \new_[25881]_  = \new_[25880]_  & \new_[25877]_ ;
  assign \new_[25882]_  = \new_[25881]_  & \new_[25874]_ ;
  assign \new_[25886]_  = ~A266 & A265;
  assign \new_[25887]_  = A202 & \new_[25886]_ ;
  assign \new_[25890]_  = A269 & A267;
  assign \new_[25893]_  = ~A300 & A298;
  assign \new_[25894]_  = \new_[25893]_  & \new_[25890]_ ;
  assign \new_[25895]_  = \new_[25894]_  & \new_[25887]_ ;
  assign \new_[25899]_  = ~A167 & ~A169;
  assign \new_[25900]_  = A170 & \new_[25899]_ ;
  assign \new_[25903]_  = A199 & A166;
  assign \new_[25906]_  = A201 & ~A200;
  assign \new_[25907]_  = \new_[25906]_  & \new_[25903]_ ;
  assign \new_[25908]_  = \new_[25907]_  & \new_[25900]_ ;
  assign \new_[25912]_  = ~A266 & A265;
  assign \new_[25913]_  = A202 & \new_[25912]_ ;
  assign \new_[25916]_  = A269 & A267;
  assign \new_[25919]_  = A299 & A298;
  assign \new_[25920]_  = \new_[25919]_  & \new_[25916]_ ;
  assign \new_[25921]_  = \new_[25920]_  & \new_[25913]_ ;
  assign \new_[25925]_  = ~A167 & ~A169;
  assign \new_[25926]_  = A170 & \new_[25925]_ ;
  assign \new_[25929]_  = A199 & A166;
  assign \new_[25932]_  = A201 & ~A200;
  assign \new_[25933]_  = \new_[25932]_  & \new_[25929]_ ;
  assign \new_[25934]_  = \new_[25933]_  & \new_[25926]_ ;
  assign \new_[25938]_  = ~A266 & A265;
  assign \new_[25939]_  = A202 & \new_[25938]_ ;
  assign \new_[25942]_  = A269 & A267;
  assign \new_[25945]_  = ~A299 & ~A298;
  assign \new_[25946]_  = \new_[25945]_  & \new_[25942]_ ;
  assign \new_[25947]_  = \new_[25946]_  & \new_[25939]_ ;
  assign \new_[25951]_  = ~A167 & ~A169;
  assign \new_[25952]_  = A170 & \new_[25951]_ ;
  assign \new_[25955]_  = A199 & A166;
  assign \new_[25958]_  = A201 & ~A200;
  assign \new_[25959]_  = \new_[25958]_  & \new_[25955]_ ;
  assign \new_[25960]_  = \new_[25959]_  & \new_[25952]_ ;
  assign \new_[25964]_  = ~A266 & A265;
  assign \new_[25965]_  = A203 & \new_[25964]_ ;
  assign \new_[25968]_  = A268 & A267;
  assign \new_[25971]_  = ~A300 & A298;
  assign \new_[25972]_  = \new_[25971]_  & \new_[25968]_ ;
  assign \new_[25973]_  = \new_[25972]_  & \new_[25965]_ ;
  assign \new_[25977]_  = ~A167 & ~A169;
  assign \new_[25978]_  = A170 & \new_[25977]_ ;
  assign \new_[25981]_  = A199 & A166;
  assign \new_[25984]_  = A201 & ~A200;
  assign \new_[25985]_  = \new_[25984]_  & \new_[25981]_ ;
  assign \new_[25986]_  = \new_[25985]_  & \new_[25978]_ ;
  assign \new_[25990]_  = ~A266 & A265;
  assign \new_[25991]_  = A203 & \new_[25990]_ ;
  assign \new_[25994]_  = A268 & A267;
  assign \new_[25997]_  = A299 & A298;
  assign \new_[25998]_  = \new_[25997]_  & \new_[25994]_ ;
  assign \new_[25999]_  = \new_[25998]_  & \new_[25991]_ ;
  assign \new_[26003]_  = ~A167 & ~A169;
  assign \new_[26004]_  = A170 & \new_[26003]_ ;
  assign \new_[26007]_  = A199 & A166;
  assign \new_[26010]_  = A201 & ~A200;
  assign \new_[26011]_  = \new_[26010]_  & \new_[26007]_ ;
  assign \new_[26012]_  = \new_[26011]_  & \new_[26004]_ ;
  assign \new_[26016]_  = ~A266 & A265;
  assign \new_[26017]_  = A203 & \new_[26016]_ ;
  assign \new_[26020]_  = A268 & A267;
  assign \new_[26023]_  = ~A299 & ~A298;
  assign \new_[26024]_  = \new_[26023]_  & \new_[26020]_ ;
  assign \new_[26025]_  = \new_[26024]_  & \new_[26017]_ ;
  assign \new_[26029]_  = ~A167 & ~A169;
  assign \new_[26030]_  = A170 & \new_[26029]_ ;
  assign \new_[26033]_  = A199 & A166;
  assign \new_[26036]_  = A201 & ~A200;
  assign \new_[26037]_  = \new_[26036]_  & \new_[26033]_ ;
  assign \new_[26038]_  = \new_[26037]_  & \new_[26030]_ ;
  assign \new_[26042]_  = ~A266 & A265;
  assign \new_[26043]_  = A203 & \new_[26042]_ ;
  assign \new_[26046]_  = A269 & A267;
  assign \new_[26049]_  = ~A300 & A298;
  assign \new_[26050]_  = \new_[26049]_  & \new_[26046]_ ;
  assign \new_[26051]_  = \new_[26050]_  & \new_[26043]_ ;
  assign \new_[26055]_  = ~A167 & ~A169;
  assign \new_[26056]_  = A170 & \new_[26055]_ ;
  assign \new_[26059]_  = A199 & A166;
  assign \new_[26062]_  = A201 & ~A200;
  assign \new_[26063]_  = \new_[26062]_  & \new_[26059]_ ;
  assign \new_[26064]_  = \new_[26063]_  & \new_[26056]_ ;
  assign \new_[26068]_  = ~A266 & A265;
  assign \new_[26069]_  = A203 & \new_[26068]_ ;
  assign \new_[26072]_  = A269 & A267;
  assign \new_[26075]_  = A299 & A298;
  assign \new_[26076]_  = \new_[26075]_  & \new_[26072]_ ;
  assign \new_[26077]_  = \new_[26076]_  & \new_[26069]_ ;
  assign \new_[26081]_  = ~A167 & ~A169;
  assign \new_[26082]_  = A170 & \new_[26081]_ ;
  assign \new_[26085]_  = A199 & A166;
  assign \new_[26088]_  = A201 & ~A200;
  assign \new_[26089]_  = \new_[26088]_  & \new_[26085]_ ;
  assign \new_[26090]_  = \new_[26089]_  & \new_[26082]_ ;
  assign \new_[26094]_  = ~A266 & A265;
  assign \new_[26095]_  = A203 & \new_[26094]_ ;
  assign \new_[26098]_  = A269 & A267;
  assign \new_[26101]_  = ~A299 & ~A298;
  assign \new_[26102]_  = \new_[26101]_  & \new_[26098]_ ;
  assign \new_[26103]_  = \new_[26102]_  & \new_[26095]_ ;
  assign \new_[26107]_  = ~A168 & ~A169;
  assign \new_[26108]_  = ~A170 & \new_[26107]_ ;
  assign \new_[26111]_  = ~A200 & A199;
  assign \new_[26114]_  = A202 & A201;
  assign \new_[26115]_  = \new_[26114]_  & \new_[26111]_ ;
  assign \new_[26116]_  = \new_[26115]_  & \new_[26108]_ ;
  assign \new_[26120]_  = ~A269 & ~A268;
  assign \new_[26121]_  = ~A266 & \new_[26120]_ ;
  assign \new_[26124]_  = ~A299 & A298;
  assign \new_[26127]_  = A301 & A300;
  assign \new_[26128]_  = \new_[26127]_  & \new_[26124]_ ;
  assign \new_[26129]_  = \new_[26128]_  & \new_[26121]_ ;
  assign \new_[26133]_  = ~A168 & ~A169;
  assign \new_[26134]_  = ~A170 & \new_[26133]_ ;
  assign \new_[26137]_  = ~A200 & A199;
  assign \new_[26140]_  = A202 & A201;
  assign \new_[26141]_  = \new_[26140]_  & \new_[26137]_ ;
  assign \new_[26142]_  = \new_[26141]_  & \new_[26134]_ ;
  assign \new_[26146]_  = ~A269 & ~A268;
  assign \new_[26147]_  = ~A266 & \new_[26146]_ ;
  assign \new_[26150]_  = ~A299 & A298;
  assign \new_[26153]_  = A302 & A300;
  assign \new_[26154]_  = \new_[26153]_  & \new_[26150]_ ;
  assign \new_[26155]_  = \new_[26154]_  & \new_[26147]_ ;
  assign \new_[26159]_  = ~A168 & ~A169;
  assign \new_[26160]_  = ~A170 & \new_[26159]_ ;
  assign \new_[26163]_  = ~A200 & A199;
  assign \new_[26166]_  = A203 & A201;
  assign \new_[26167]_  = \new_[26166]_  & \new_[26163]_ ;
  assign \new_[26168]_  = \new_[26167]_  & \new_[26160]_ ;
  assign \new_[26172]_  = ~A269 & ~A268;
  assign \new_[26173]_  = ~A266 & \new_[26172]_ ;
  assign \new_[26176]_  = ~A299 & A298;
  assign \new_[26179]_  = A301 & A300;
  assign \new_[26180]_  = \new_[26179]_  & \new_[26176]_ ;
  assign \new_[26181]_  = \new_[26180]_  & \new_[26173]_ ;
  assign \new_[26185]_  = ~A168 & ~A169;
  assign \new_[26186]_  = ~A170 & \new_[26185]_ ;
  assign \new_[26189]_  = ~A200 & A199;
  assign \new_[26192]_  = A203 & A201;
  assign \new_[26193]_  = \new_[26192]_  & \new_[26189]_ ;
  assign \new_[26194]_  = \new_[26193]_  & \new_[26186]_ ;
  assign \new_[26198]_  = ~A269 & ~A268;
  assign \new_[26199]_  = ~A266 & \new_[26198]_ ;
  assign \new_[26202]_  = ~A299 & A298;
  assign \new_[26205]_  = A302 & A300;
  assign \new_[26206]_  = \new_[26205]_  & \new_[26202]_ ;
  assign \new_[26207]_  = \new_[26206]_  & \new_[26199]_ ;
  assign \new_[26211]_  = A167 & ~A168;
  assign \new_[26212]_  = A169 & \new_[26211]_ ;
  assign \new_[26215]_  = A199 & ~A166;
  assign \new_[26218]_  = A201 & ~A200;
  assign \new_[26219]_  = \new_[26218]_  & \new_[26215]_ ;
  assign \new_[26220]_  = \new_[26219]_  & \new_[26212]_ ;
  assign \new_[26223]_  = ~A266 & A202;
  assign \new_[26226]_  = ~A269 & ~A268;
  assign \new_[26227]_  = \new_[26226]_  & \new_[26223]_ ;
  assign \new_[26230]_  = ~A299 & A298;
  assign \new_[26233]_  = A301 & A300;
  assign \new_[26234]_  = \new_[26233]_  & \new_[26230]_ ;
  assign \new_[26235]_  = \new_[26234]_  & \new_[26227]_ ;
  assign \new_[26239]_  = A167 & ~A168;
  assign \new_[26240]_  = A169 & \new_[26239]_ ;
  assign \new_[26243]_  = A199 & ~A166;
  assign \new_[26246]_  = A201 & ~A200;
  assign \new_[26247]_  = \new_[26246]_  & \new_[26243]_ ;
  assign \new_[26248]_  = \new_[26247]_  & \new_[26240]_ ;
  assign \new_[26251]_  = ~A266 & A202;
  assign \new_[26254]_  = ~A269 & ~A268;
  assign \new_[26255]_  = \new_[26254]_  & \new_[26251]_ ;
  assign \new_[26258]_  = ~A299 & A298;
  assign \new_[26261]_  = A302 & A300;
  assign \new_[26262]_  = \new_[26261]_  & \new_[26258]_ ;
  assign \new_[26263]_  = \new_[26262]_  & \new_[26255]_ ;
  assign \new_[26267]_  = A167 & ~A168;
  assign \new_[26268]_  = A169 & \new_[26267]_ ;
  assign \new_[26271]_  = A199 & ~A166;
  assign \new_[26274]_  = A201 & ~A200;
  assign \new_[26275]_  = \new_[26274]_  & \new_[26271]_ ;
  assign \new_[26276]_  = \new_[26275]_  & \new_[26268]_ ;
  assign \new_[26279]_  = ~A266 & A203;
  assign \new_[26282]_  = ~A269 & ~A268;
  assign \new_[26283]_  = \new_[26282]_  & \new_[26279]_ ;
  assign \new_[26286]_  = ~A299 & A298;
  assign \new_[26289]_  = A301 & A300;
  assign \new_[26290]_  = \new_[26289]_  & \new_[26286]_ ;
  assign \new_[26291]_  = \new_[26290]_  & \new_[26283]_ ;
  assign \new_[26295]_  = A167 & ~A168;
  assign \new_[26296]_  = A169 & \new_[26295]_ ;
  assign \new_[26299]_  = A199 & ~A166;
  assign \new_[26302]_  = A201 & ~A200;
  assign \new_[26303]_  = \new_[26302]_  & \new_[26299]_ ;
  assign \new_[26304]_  = \new_[26303]_  & \new_[26296]_ ;
  assign \new_[26307]_  = ~A266 & A203;
  assign \new_[26310]_  = ~A269 & ~A268;
  assign \new_[26311]_  = \new_[26310]_  & \new_[26307]_ ;
  assign \new_[26314]_  = ~A299 & A298;
  assign \new_[26317]_  = A302 & A300;
  assign \new_[26318]_  = \new_[26317]_  & \new_[26314]_ ;
  assign \new_[26319]_  = \new_[26318]_  & \new_[26311]_ ;
  assign \new_[26323]_  = ~A167 & ~A168;
  assign \new_[26324]_  = A169 & \new_[26323]_ ;
  assign \new_[26327]_  = A199 & A166;
  assign \new_[26330]_  = A201 & ~A200;
  assign \new_[26331]_  = \new_[26330]_  & \new_[26327]_ ;
  assign \new_[26332]_  = \new_[26331]_  & \new_[26324]_ ;
  assign \new_[26335]_  = ~A266 & A202;
  assign \new_[26338]_  = ~A269 & ~A268;
  assign \new_[26339]_  = \new_[26338]_  & \new_[26335]_ ;
  assign \new_[26342]_  = ~A299 & A298;
  assign \new_[26345]_  = A301 & A300;
  assign \new_[26346]_  = \new_[26345]_  & \new_[26342]_ ;
  assign \new_[26347]_  = \new_[26346]_  & \new_[26339]_ ;
  assign \new_[26351]_  = ~A167 & ~A168;
  assign \new_[26352]_  = A169 & \new_[26351]_ ;
  assign \new_[26355]_  = A199 & A166;
  assign \new_[26358]_  = A201 & ~A200;
  assign \new_[26359]_  = \new_[26358]_  & \new_[26355]_ ;
  assign \new_[26360]_  = \new_[26359]_  & \new_[26352]_ ;
  assign \new_[26363]_  = ~A266 & A202;
  assign \new_[26366]_  = ~A269 & ~A268;
  assign \new_[26367]_  = \new_[26366]_  & \new_[26363]_ ;
  assign \new_[26370]_  = ~A299 & A298;
  assign \new_[26373]_  = A302 & A300;
  assign \new_[26374]_  = \new_[26373]_  & \new_[26370]_ ;
  assign \new_[26375]_  = \new_[26374]_  & \new_[26367]_ ;
  assign \new_[26379]_  = ~A167 & ~A168;
  assign \new_[26380]_  = A169 & \new_[26379]_ ;
  assign \new_[26383]_  = A199 & A166;
  assign \new_[26386]_  = A201 & ~A200;
  assign \new_[26387]_  = \new_[26386]_  & \new_[26383]_ ;
  assign \new_[26388]_  = \new_[26387]_  & \new_[26380]_ ;
  assign \new_[26391]_  = ~A266 & A203;
  assign \new_[26394]_  = ~A269 & ~A268;
  assign \new_[26395]_  = \new_[26394]_  & \new_[26391]_ ;
  assign \new_[26398]_  = ~A299 & A298;
  assign \new_[26401]_  = A301 & A300;
  assign \new_[26402]_  = \new_[26401]_  & \new_[26398]_ ;
  assign \new_[26403]_  = \new_[26402]_  & \new_[26395]_ ;
  assign \new_[26407]_  = ~A167 & ~A168;
  assign \new_[26408]_  = A169 & \new_[26407]_ ;
  assign \new_[26411]_  = A199 & A166;
  assign \new_[26414]_  = A201 & ~A200;
  assign \new_[26415]_  = \new_[26414]_  & \new_[26411]_ ;
  assign \new_[26416]_  = \new_[26415]_  & \new_[26408]_ ;
  assign \new_[26419]_  = ~A266 & A203;
  assign \new_[26422]_  = ~A269 & ~A268;
  assign \new_[26423]_  = \new_[26422]_  & \new_[26419]_ ;
  assign \new_[26426]_  = ~A299 & A298;
  assign \new_[26429]_  = A302 & A300;
  assign \new_[26430]_  = \new_[26429]_  & \new_[26426]_ ;
  assign \new_[26431]_  = \new_[26430]_  & \new_[26423]_ ;
  assign \new_[26435]_  = A167 & A169;
  assign \new_[26436]_  = ~A170 & \new_[26435]_ ;
  assign \new_[26439]_  = A199 & A166;
  assign \new_[26442]_  = A201 & ~A200;
  assign \new_[26443]_  = \new_[26442]_  & \new_[26439]_ ;
  assign \new_[26444]_  = \new_[26443]_  & \new_[26436]_ ;
  assign \new_[26447]_  = A265 & A202;
  assign \new_[26450]_  = A267 & ~A266;
  assign \new_[26451]_  = \new_[26450]_  & \new_[26447]_ ;
  assign \new_[26454]_  = A298 & A268;
  assign \new_[26457]_  = ~A302 & ~A301;
  assign \new_[26458]_  = \new_[26457]_  & \new_[26454]_ ;
  assign \new_[26459]_  = \new_[26458]_  & \new_[26451]_ ;
  assign \new_[26463]_  = A167 & A169;
  assign \new_[26464]_  = ~A170 & \new_[26463]_ ;
  assign \new_[26467]_  = A199 & A166;
  assign \new_[26470]_  = A201 & ~A200;
  assign \new_[26471]_  = \new_[26470]_  & \new_[26467]_ ;
  assign \new_[26472]_  = \new_[26471]_  & \new_[26464]_ ;
  assign \new_[26475]_  = A265 & A202;
  assign \new_[26478]_  = A267 & ~A266;
  assign \new_[26479]_  = \new_[26478]_  & \new_[26475]_ ;
  assign \new_[26482]_  = A298 & A269;
  assign \new_[26485]_  = ~A302 & ~A301;
  assign \new_[26486]_  = \new_[26485]_  & \new_[26482]_ ;
  assign \new_[26487]_  = \new_[26486]_  & \new_[26479]_ ;
  assign \new_[26491]_  = A167 & A169;
  assign \new_[26492]_  = ~A170 & \new_[26491]_ ;
  assign \new_[26495]_  = A199 & A166;
  assign \new_[26498]_  = A201 & ~A200;
  assign \new_[26499]_  = \new_[26498]_  & \new_[26495]_ ;
  assign \new_[26500]_  = \new_[26499]_  & \new_[26492]_ ;
  assign \new_[26503]_  = A265 & A203;
  assign \new_[26506]_  = A267 & ~A266;
  assign \new_[26507]_  = \new_[26506]_  & \new_[26503]_ ;
  assign \new_[26510]_  = A298 & A268;
  assign \new_[26513]_  = ~A302 & ~A301;
  assign \new_[26514]_  = \new_[26513]_  & \new_[26510]_ ;
  assign \new_[26515]_  = \new_[26514]_  & \new_[26507]_ ;
  assign \new_[26519]_  = A167 & A169;
  assign \new_[26520]_  = ~A170 & \new_[26519]_ ;
  assign \new_[26523]_  = A199 & A166;
  assign \new_[26526]_  = A201 & ~A200;
  assign \new_[26527]_  = \new_[26526]_  & \new_[26523]_ ;
  assign \new_[26528]_  = \new_[26527]_  & \new_[26520]_ ;
  assign \new_[26531]_  = A265 & A203;
  assign \new_[26534]_  = A267 & ~A266;
  assign \new_[26535]_  = \new_[26534]_  & \new_[26531]_ ;
  assign \new_[26538]_  = A298 & A269;
  assign \new_[26541]_  = ~A302 & ~A301;
  assign \new_[26542]_  = \new_[26541]_  & \new_[26538]_ ;
  assign \new_[26543]_  = \new_[26542]_  & \new_[26535]_ ;
  assign \new_[26547]_  = ~A167 & A169;
  assign \new_[26548]_  = ~A170 & \new_[26547]_ ;
  assign \new_[26551]_  = A199 & ~A166;
  assign \new_[26554]_  = A201 & ~A200;
  assign \new_[26555]_  = \new_[26554]_  & \new_[26551]_ ;
  assign \new_[26556]_  = \new_[26555]_  & \new_[26548]_ ;
  assign \new_[26559]_  = A265 & A202;
  assign \new_[26562]_  = A267 & ~A266;
  assign \new_[26563]_  = \new_[26562]_  & \new_[26559]_ ;
  assign \new_[26566]_  = A298 & A268;
  assign \new_[26569]_  = ~A302 & ~A301;
  assign \new_[26570]_  = \new_[26569]_  & \new_[26566]_ ;
  assign \new_[26571]_  = \new_[26570]_  & \new_[26563]_ ;
  assign \new_[26575]_  = ~A167 & A169;
  assign \new_[26576]_  = ~A170 & \new_[26575]_ ;
  assign \new_[26579]_  = A199 & ~A166;
  assign \new_[26582]_  = A201 & ~A200;
  assign \new_[26583]_  = \new_[26582]_  & \new_[26579]_ ;
  assign \new_[26584]_  = \new_[26583]_  & \new_[26576]_ ;
  assign \new_[26587]_  = A265 & A202;
  assign \new_[26590]_  = A267 & ~A266;
  assign \new_[26591]_  = \new_[26590]_  & \new_[26587]_ ;
  assign \new_[26594]_  = A298 & A269;
  assign \new_[26597]_  = ~A302 & ~A301;
  assign \new_[26598]_  = \new_[26597]_  & \new_[26594]_ ;
  assign \new_[26599]_  = \new_[26598]_  & \new_[26591]_ ;
  assign \new_[26603]_  = ~A167 & A169;
  assign \new_[26604]_  = ~A170 & \new_[26603]_ ;
  assign \new_[26607]_  = A199 & ~A166;
  assign \new_[26610]_  = A201 & ~A200;
  assign \new_[26611]_  = \new_[26610]_  & \new_[26607]_ ;
  assign \new_[26612]_  = \new_[26611]_  & \new_[26604]_ ;
  assign \new_[26615]_  = A265 & A203;
  assign \new_[26618]_  = A267 & ~A266;
  assign \new_[26619]_  = \new_[26618]_  & \new_[26615]_ ;
  assign \new_[26622]_  = A298 & A268;
  assign \new_[26625]_  = ~A302 & ~A301;
  assign \new_[26626]_  = \new_[26625]_  & \new_[26622]_ ;
  assign \new_[26627]_  = \new_[26626]_  & \new_[26619]_ ;
  assign \new_[26631]_  = ~A167 & A169;
  assign \new_[26632]_  = ~A170 & \new_[26631]_ ;
  assign \new_[26635]_  = A199 & ~A166;
  assign \new_[26638]_  = A201 & ~A200;
  assign \new_[26639]_  = \new_[26638]_  & \new_[26635]_ ;
  assign \new_[26640]_  = \new_[26639]_  & \new_[26632]_ ;
  assign \new_[26643]_  = A265 & A203;
  assign \new_[26646]_  = A267 & ~A266;
  assign \new_[26647]_  = \new_[26646]_  & \new_[26643]_ ;
  assign \new_[26650]_  = A298 & A269;
  assign \new_[26653]_  = ~A302 & ~A301;
  assign \new_[26654]_  = \new_[26653]_  & \new_[26650]_ ;
  assign \new_[26655]_  = \new_[26654]_  & \new_[26647]_ ;
  assign \new_[26659]_  = A167 & ~A168;
  assign \new_[26660]_  = ~A169 & \new_[26659]_ ;
  assign \new_[26663]_  = A199 & A166;
  assign \new_[26666]_  = A201 & ~A200;
  assign \new_[26667]_  = \new_[26666]_  & \new_[26663]_ ;
  assign \new_[26668]_  = \new_[26667]_  & \new_[26660]_ ;
  assign \new_[26671]_  = ~A266 & A202;
  assign \new_[26674]_  = ~A269 & ~A268;
  assign \new_[26675]_  = \new_[26674]_  & \new_[26671]_ ;
  assign \new_[26678]_  = ~A299 & A298;
  assign \new_[26681]_  = A301 & A300;
  assign \new_[26682]_  = \new_[26681]_  & \new_[26678]_ ;
  assign \new_[26683]_  = \new_[26682]_  & \new_[26675]_ ;
  assign \new_[26687]_  = A167 & ~A168;
  assign \new_[26688]_  = ~A169 & \new_[26687]_ ;
  assign \new_[26691]_  = A199 & A166;
  assign \new_[26694]_  = A201 & ~A200;
  assign \new_[26695]_  = \new_[26694]_  & \new_[26691]_ ;
  assign \new_[26696]_  = \new_[26695]_  & \new_[26688]_ ;
  assign \new_[26699]_  = ~A266 & A202;
  assign \new_[26702]_  = ~A269 & ~A268;
  assign \new_[26703]_  = \new_[26702]_  & \new_[26699]_ ;
  assign \new_[26706]_  = ~A299 & A298;
  assign \new_[26709]_  = A302 & A300;
  assign \new_[26710]_  = \new_[26709]_  & \new_[26706]_ ;
  assign \new_[26711]_  = \new_[26710]_  & \new_[26703]_ ;
  assign \new_[26715]_  = A167 & ~A168;
  assign \new_[26716]_  = ~A169 & \new_[26715]_ ;
  assign \new_[26719]_  = A199 & A166;
  assign \new_[26722]_  = A201 & ~A200;
  assign \new_[26723]_  = \new_[26722]_  & \new_[26719]_ ;
  assign \new_[26724]_  = \new_[26723]_  & \new_[26716]_ ;
  assign \new_[26727]_  = ~A266 & A203;
  assign \new_[26730]_  = ~A269 & ~A268;
  assign \new_[26731]_  = \new_[26730]_  & \new_[26727]_ ;
  assign \new_[26734]_  = ~A299 & A298;
  assign \new_[26737]_  = A301 & A300;
  assign \new_[26738]_  = \new_[26737]_  & \new_[26734]_ ;
  assign \new_[26739]_  = \new_[26738]_  & \new_[26731]_ ;
  assign \new_[26743]_  = A167 & ~A168;
  assign \new_[26744]_  = ~A169 & \new_[26743]_ ;
  assign \new_[26747]_  = A199 & A166;
  assign \new_[26750]_  = A201 & ~A200;
  assign \new_[26751]_  = \new_[26750]_  & \new_[26747]_ ;
  assign \new_[26752]_  = \new_[26751]_  & \new_[26744]_ ;
  assign \new_[26755]_  = ~A266 & A203;
  assign \new_[26758]_  = ~A269 & ~A268;
  assign \new_[26759]_  = \new_[26758]_  & \new_[26755]_ ;
  assign \new_[26762]_  = ~A299 & A298;
  assign \new_[26765]_  = A302 & A300;
  assign \new_[26766]_  = \new_[26765]_  & \new_[26762]_ ;
  assign \new_[26767]_  = \new_[26766]_  & \new_[26759]_ ;
  assign \new_[26771]_  = A167 & ~A169;
  assign \new_[26772]_  = A170 & \new_[26771]_ ;
  assign \new_[26775]_  = A199 & ~A166;
  assign \new_[26778]_  = A201 & ~A200;
  assign \new_[26779]_  = \new_[26778]_  & \new_[26775]_ ;
  assign \new_[26780]_  = \new_[26779]_  & \new_[26772]_ ;
  assign \new_[26783]_  = A265 & A202;
  assign \new_[26786]_  = A267 & ~A266;
  assign \new_[26787]_  = \new_[26786]_  & \new_[26783]_ ;
  assign \new_[26790]_  = A298 & A268;
  assign \new_[26793]_  = ~A302 & ~A301;
  assign \new_[26794]_  = \new_[26793]_  & \new_[26790]_ ;
  assign \new_[26795]_  = \new_[26794]_  & \new_[26787]_ ;
  assign \new_[26799]_  = A167 & ~A169;
  assign \new_[26800]_  = A170 & \new_[26799]_ ;
  assign \new_[26803]_  = A199 & ~A166;
  assign \new_[26806]_  = A201 & ~A200;
  assign \new_[26807]_  = \new_[26806]_  & \new_[26803]_ ;
  assign \new_[26808]_  = \new_[26807]_  & \new_[26800]_ ;
  assign \new_[26811]_  = A265 & A202;
  assign \new_[26814]_  = A267 & ~A266;
  assign \new_[26815]_  = \new_[26814]_  & \new_[26811]_ ;
  assign \new_[26818]_  = A298 & A269;
  assign \new_[26821]_  = ~A302 & ~A301;
  assign \new_[26822]_  = \new_[26821]_  & \new_[26818]_ ;
  assign \new_[26823]_  = \new_[26822]_  & \new_[26815]_ ;
  assign \new_[26827]_  = A167 & ~A169;
  assign \new_[26828]_  = A170 & \new_[26827]_ ;
  assign \new_[26831]_  = A199 & ~A166;
  assign \new_[26834]_  = A201 & ~A200;
  assign \new_[26835]_  = \new_[26834]_  & \new_[26831]_ ;
  assign \new_[26836]_  = \new_[26835]_  & \new_[26828]_ ;
  assign \new_[26839]_  = A265 & A203;
  assign \new_[26842]_  = A267 & ~A266;
  assign \new_[26843]_  = \new_[26842]_  & \new_[26839]_ ;
  assign \new_[26846]_  = A298 & A268;
  assign \new_[26849]_  = ~A302 & ~A301;
  assign \new_[26850]_  = \new_[26849]_  & \new_[26846]_ ;
  assign \new_[26851]_  = \new_[26850]_  & \new_[26843]_ ;
  assign \new_[26855]_  = A167 & ~A169;
  assign \new_[26856]_  = A170 & \new_[26855]_ ;
  assign \new_[26859]_  = A199 & ~A166;
  assign \new_[26862]_  = A201 & ~A200;
  assign \new_[26863]_  = \new_[26862]_  & \new_[26859]_ ;
  assign \new_[26864]_  = \new_[26863]_  & \new_[26856]_ ;
  assign \new_[26867]_  = A265 & A203;
  assign \new_[26870]_  = A267 & ~A266;
  assign \new_[26871]_  = \new_[26870]_  & \new_[26867]_ ;
  assign \new_[26874]_  = A298 & A269;
  assign \new_[26877]_  = ~A302 & ~A301;
  assign \new_[26878]_  = \new_[26877]_  & \new_[26874]_ ;
  assign \new_[26879]_  = \new_[26878]_  & \new_[26871]_ ;
  assign \new_[26883]_  = ~A167 & ~A169;
  assign \new_[26884]_  = A170 & \new_[26883]_ ;
  assign \new_[26887]_  = A199 & A166;
  assign \new_[26890]_  = A201 & ~A200;
  assign \new_[26891]_  = \new_[26890]_  & \new_[26887]_ ;
  assign \new_[26892]_  = \new_[26891]_  & \new_[26884]_ ;
  assign \new_[26895]_  = A265 & A202;
  assign \new_[26898]_  = A267 & ~A266;
  assign \new_[26899]_  = \new_[26898]_  & \new_[26895]_ ;
  assign \new_[26902]_  = A298 & A268;
  assign \new_[26905]_  = ~A302 & ~A301;
  assign \new_[26906]_  = \new_[26905]_  & \new_[26902]_ ;
  assign \new_[26907]_  = \new_[26906]_  & \new_[26899]_ ;
  assign \new_[26911]_  = ~A167 & ~A169;
  assign \new_[26912]_  = A170 & \new_[26911]_ ;
  assign \new_[26915]_  = A199 & A166;
  assign \new_[26918]_  = A201 & ~A200;
  assign \new_[26919]_  = \new_[26918]_  & \new_[26915]_ ;
  assign \new_[26920]_  = \new_[26919]_  & \new_[26912]_ ;
  assign \new_[26923]_  = A265 & A202;
  assign \new_[26926]_  = A267 & ~A266;
  assign \new_[26927]_  = \new_[26926]_  & \new_[26923]_ ;
  assign \new_[26930]_  = A298 & A269;
  assign \new_[26933]_  = ~A302 & ~A301;
  assign \new_[26934]_  = \new_[26933]_  & \new_[26930]_ ;
  assign \new_[26935]_  = \new_[26934]_  & \new_[26927]_ ;
  assign \new_[26939]_  = ~A167 & ~A169;
  assign \new_[26940]_  = A170 & \new_[26939]_ ;
  assign \new_[26943]_  = A199 & A166;
  assign \new_[26946]_  = A201 & ~A200;
  assign \new_[26947]_  = \new_[26946]_  & \new_[26943]_ ;
  assign \new_[26948]_  = \new_[26947]_  & \new_[26940]_ ;
  assign \new_[26951]_  = A265 & A203;
  assign \new_[26954]_  = A267 & ~A266;
  assign \new_[26955]_  = \new_[26954]_  & \new_[26951]_ ;
  assign \new_[26958]_  = A298 & A268;
  assign \new_[26961]_  = ~A302 & ~A301;
  assign \new_[26962]_  = \new_[26961]_  & \new_[26958]_ ;
  assign \new_[26963]_  = \new_[26962]_  & \new_[26955]_ ;
  assign \new_[26967]_  = ~A167 & ~A169;
  assign \new_[26968]_  = A170 & \new_[26967]_ ;
  assign \new_[26971]_  = A199 & A166;
  assign \new_[26974]_  = A201 & ~A200;
  assign \new_[26975]_  = \new_[26974]_  & \new_[26971]_ ;
  assign \new_[26976]_  = \new_[26975]_  & \new_[26968]_ ;
  assign \new_[26979]_  = A265 & A203;
  assign \new_[26982]_  = A267 & ~A266;
  assign \new_[26983]_  = \new_[26982]_  & \new_[26979]_ ;
  assign \new_[26986]_  = A298 & A269;
  assign \new_[26989]_  = ~A302 & ~A301;
  assign \new_[26990]_  = \new_[26989]_  & \new_[26986]_ ;
  assign \new_[26991]_  = \new_[26990]_  & \new_[26983]_ ;
endmodule


