// Benchmark "spi" written by ABC on Thu Oct  8 22:04:26 2020

module spi ( clock, 
    wb_clk_i, wb_rst_i, wb_we_i, wb_stb_i, wb_cyc_i, miso_pad_i,
    \wb_adr_i[0] , \wb_adr_i[1] , \wb_adr_i[2] , \wb_adr_i[3] ,
    \wb_adr_i[4] , \wb_dat_i[0] , \wb_dat_i[1] , \wb_dat_i[2] ,
    \wb_dat_i[3] , \wb_dat_i[4] , \wb_dat_i[5] , \wb_dat_i[6] ,
    \wb_dat_i[7] , \wb_dat_i[8] , \wb_dat_i[9] , \wb_dat_i[10] ,
    \wb_dat_i[11] , \wb_dat_i[12] , \wb_dat_i[13] , \wb_dat_i[14] ,
    \wb_dat_i[15] , \wb_dat_i[16] , \wb_dat_i[17] , \wb_dat_i[18] ,
    \wb_dat_i[19] , \wb_dat_i[20] , \wb_dat_i[21] , \wb_dat_i[22] ,
    \wb_dat_i[23] , \wb_dat_i[24] , \wb_dat_i[25] , \wb_dat_i[26] ,
    \wb_dat_i[27] , \wb_dat_i[28] , \wb_dat_i[29] , \wb_dat_i[30] ,
    \wb_dat_i[31] , \wb_sel_i[0] , \wb_sel_i[1] , \wb_sel_i[2] ,
    \wb_sel_i[3] ,
    \wb_dat_o[0] , \wb_dat_o[1] , \wb_dat_o[2] , \wb_dat_o[3] ,
    \wb_dat_o[4] , \wb_dat_o[5] , \wb_dat_o[6] , \wb_dat_o[7] ,
    \wb_dat_o[8] , \wb_dat_o[9] , \wb_dat_o[10] , \wb_dat_o[11] ,
    \wb_dat_o[12] , \wb_dat_o[13] , \wb_dat_o[14] , \wb_dat_o[15] ,
    \wb_dat_o[16] , \wb_dat_o[17] , \wb_dat_o[18] , \wb_dat_o[19] ,
    \wb_dat_o[20] , \wb_dat_o[21] , \wb_dat_o[22] , \wb_dat_o[23] ,
    \wb_dat_o[24] , \wb_dat_o[25] , \wb_dat_o[26] , \wb_dat_o[27] ,
    \wb_dat_o[28] , \wb_dat_o[29] , \wb_dat_o[30] , \wb_dat_o[31] ,
    wb_ack_o, wb_err_o, wb_int_o, sclk_pad_o, mosi_pad_o, \ss_pad_o[0] ,
    \ss_pad_o[1] , \ss_pad_o[2] , \ss_pad_o[3] , \ss_pad_o[4] ,
    \ss_pad_o[5] , \ss_pad_o[6] , \ss_pad_o[7]   );
  input  clock;
  input  wb_clk_i, wb_rst_i, wb_we_i, wb_stb_i, wb_cyc_i, miso_pad_i,
    \wb_adr_i[0] , \wb_adr_i[1] , \wb_adr_i[2] , \wb_adr_i[3] ,
    \wb_adr_i[4] , \wb_dat_i[0] , \wb_dat_i[1] , \wb_dat_i[2] ,
    \wb_dat_i[3] , \wb_dat_i[4] , \wb_dat_i[5] , \wb_dat_i[6] ,
    \wb_dat_i[7] , \wb_dat_i[8] , \wb_dat_i[9] , \wb_dat_i[10] ,
    \wb_dat_i[11] , \wb_dat_i[12] , \wb_dat_i[13] , \wb_dat_i[14] ,
    \wb_dat_i[15] , \wb_dat_i[16] , \wb_dat_i[17] , \wb_dat_i[18] ,
    \wb_dat_i[19] , \wb_dat_i[20] , \wb_dat_i[21] , \wb_dat_i[22] ,
    \wb_dat_i[23] , \wb_dat_i[24] , \wb_dat_i[25] , \wb_dat_i[26] ,
    \wb_dat_i[27] , \wb_dat_i[28] , \wb_dat_i[29] , \wb_dat_i[30] ,
    \wb_dat_i[31] , \wb_sel_i[0] , \wb_sel_i[1] , \wb_sel_i[2] ,
    \wb_sel_i[3] ;
  output \wb_dat_o[0] , \wb_dat_o[1] , \wb_dat_o[2] , \wb_dat_o[3] ,
    \wb_dat_o[4] , \wb_dat_o[5] , \wb_dat_o[6] , \wb_dat_o[7] ,
    \wb_dat_o[8] , \wb_dat_o[9] , \wb_dat_o[10] , \wb_dat_o[11] ,
    \wb_dat_o[12] , \wb_dat_o[13] , \wb_dat_o[14] , \wb_dat_o[15] ,
    \wb_dat_o[16] , \wb_dat_o[17] , \wb_dat_o[18] , \wb_dat_o[19] ,
    \wb_dat_o[20] , \wb_dat_o[21] , \wb_dat_o[22] , \wb_dat_o[23] ,
    \wb_dat_o[24] , \wb_dat_o[25] , \wb_dat_o[26] , \wb_dat_o[27] ,
    \wb_dat_o[28] , \wb_dat_o[29] , \wb_dat_o[30] , \wb_dat_o[31] ,
    wb_ack_o, wb_err_o, wb_int_o, sclk_pad_o, mosi_pad_o, \ss_pad_o[0] ,
    \ss_pad_o[1] , \ss_pad_o[2] , \ss_pad_o[3] , \ss_pad_o[4] ,
    \ss_pad_o[5] , \ss_pad_o[6] , \ss_pad_o[7] ;
  reg \\shift_data_reg[39] , \\shift_data_reg[56] , \\shift_data_reg[63] ,
    \\shift_data_reg[32] , \\shift_data_reg[65] , \\shift_data_reg[66] ,
    \\shift_data_reg[68] , \\shift_data_reg[71] , \\shift_data_reg[74] ,
    \\shift_data_reg[75] , \\shift_data_reg[76] , \\shift_data_reg[85] ,
    \\shift_data_reg[86] , \\shift_data_reg[87] , \\shift_data_reg[91] ,
    \\shift_data_reg[93] , \\shift_data_reg[94] , \\shift_data_reg[95] ,
    \\shift_data_reg[0] , \\shift_data_reg[2] , \\shift_data_reg[4] ,
    \\shift_data_reg[7] , \\shift_data_reg[8] , \\shift_data_reg[14] ,
    \\shift_data_reg[15] , \\shift_data_reg[16] , \\shift_data_reg[17] ,
    \\shift_data_reg[18] , \\shift_data_reg[1] , \\shift_data_reg[20] ,
    \\shift_data_reg[23] , \\shift_data_reg[92] , \\shift_data_reg[89] ,
    \\shift_data_reg[64] , \\shift_data_reg[67] , \\shift_data_reg[69] ,
    \\shift_data_reg[70] , \\shift_data_reg[72] , \\shift_data_reg[73] ,
    \\shift_data_reg[77] , \\shift_data_reg[80] , \\shift_data_reg[83] ,
    \\shift_data_reg[84] , \\shift_data_reg[81] , \\shift_data_reg[88] ,
    \\shift_data_reg[82] , \\shift_data_reg[90] , \\shift_data_reg[79] ,
    \\shift_data_reg[78] , \\shift_data_reg[26] , \\shift_data_reg[27] ,
    \\shift_data_reg[24] , \\shift_data_reg[29] , \\shift_data_reg[28] ,
    \\shift_data_reg[30] , \\shift_data_reg[31] , \\shift_data_reg[10] ,
    \\shift_data_reg[3] , \\shift_data_reg[5] , \\shift_data_reg[25] ,
    \\shift_data_reg[6] , \\shift_data_reg[12] , \\shift_data_reg[13] ,
    \\shift_data_reg[11] , \\shift_data_reg[9] , \\shift_data_reg[19] ,
    \\shift_data_reg[21] , \\shift_data_reg[22] , \\shift_data_reg[53] ,
    \\shift_data_reg[54] , \\shift_data_reg[51] , \\shift_data_reg[33] ,
    \\shift_data_reg[34] , \\shift_data_reg[35] , \\shift_data_reg[36] ,
    \\shift_data_reg[43] , \\shift_data_reg[45] , \\shift_data_reg[46] ,
    \\shift_data_reg[47] , \\shift_data_reg[57] , \\shift_data_reg[58] ,
    \\shift_data_reg[59] , \\shift_data_reg[61] , \\shift_data_reg[62] ,
    \\shift_data_reg[104] , \\shift_data_reg[111] , \\shift_data_reg[112] ,
    \\shift_data_reg[119] , \\shift_data_reg[121] , \\shift_data_reg[97] ,
    \\shift_data_reg[123] , \\shift_data_reg[125] , \\shift_data_reg[126] ,
    \\shift_data_reg[122] , \\shift_data_reg[127] , \\shift_data_reg[124] ,
    \\shift_data_reg[98] , \\shift_data_reg[114] , \\shift_data_reg[60] ,
    \\shift_data_reg[48] , \\shift_data_reg[41] , \\shift_data_reg[40] ,
    \\shift_data_reg[120] , \\shift_data_reg[105] , \\shift_data_reg[113] ,
    \\shift_data_reg[108] , \\shift_data_reg[37] , \\shift_data_reg[38] ,
    \\shift_data_reg[116] , \\shift_data_reg[42] , \\shift_data_reg[49] ,
    \\shift_data_reg[50] , \\shift_data_reg[44] , \\shift_data_reg[52] ,
    \\shift_data_reg[55] , \\shift_data_reg[103] , \\shift_data_reg[100] ,
    \\shift_data_reg[106] , \\shift_data_reg[96] , \\shift_data_reg[99] ,
    \\shift_data_reg[118] , \\shift_data_reg[115] , \\shift_data_reg[101] ,
    \\shift_data_reg[102] , \\shift_data_reg[107] , \\shift_data_reg[109] ,
    \\shift_data_reg[110] , \\shift_data_reg[117] , shift_s_out_reg,
    clgen_clk_out_reg, \\shift_cnt_reg[7] , \\ctrl_reg[8] ,
    \\clgen_cnt_reg[15] , \\shift_cnt_reg[6] , wb_int_o_reg,
    \\wb_dat_o_reg[9] , shift_tip_reg, \\wb_dat_o_reg[11] , \\ctrl_reg[9] ,
    \\shift_cnt_reg[4] , \\shift_cnt_reg[5] , \\clgen_cnt_reg[11] ,
    \\shift_cnt_reg[3] , \\ctrl_reg[11] , \\ctrl_reg[10] ,
    clgen_pos_edge_reg, clgen_neg_edge_reg, \\clgen_cnt_reg[14] ,
    \\shift_cnt_reg[2] , \\clgen_cnt_reg[13] , \\ctrl_reg[0] ,
    \\ctrl_reg[12] , \\ctrl_reg[13] , \\divider_reg[11] ,
    \\clgen_cnt_reg[12] , \\divider_reg[4] , \\ctrl_reg[2] ,
    \\divider_reg[15] , \\ctrl_reg[7] , \\clgen_cnt_reg[10] ,
    \\divider_reg[8] , \\ctrl_reg[5] , \\clgen_cnt_reg[3] ,
    \\divider_reg[13] , \\clgen_cnt_reg[5] , \\clgen_cnt_reg[0] ,
    \\clgen_cnt_reg[2] , \\clgen_cnt_reg[7] , \\clgen_cnt_reg[6] ,
    \\clgen_cnt_reg[9] , \\clgen_cnt_reg[1] , \\ctrl_reg[1] ,
    \\divider_reg[12] , \\divider_reg[10] , \\divider_reg[1] ,
    \\divider_reg[2] , \\ctrl_reg[3] , \\ctrl_reg[4] , \\ctrl_reg[6] ,
    \\divider_reg[0] , \\divider_reg[14] , \\divider_reg[3] ,
    \\divider_reg[5] , \\divider_reg[6] , \\divider_reg[7] ,
    \\divider_reg[9] , \\clgen_cnt_reg[4] , \\shift_cnt_reg[1] ,
    \\wb_dat_o_reg[7] , \\wb_dat_o_reg[3] , \\shift_cnt_reg[0] ,
    \\clgen_cnt_reg[8] , \\ss_reg[5] , \\ss_reg[3] , \\ss_reg[1] ,
    \\ss_reg[7] , \\ss_reg[0] , \\ss_reg[2] , \\ss_reg[4] , \\ss_reg[6] ,
    \\wb_dat_o_reg[4] , \\wb_dat_o_reg[5] , \\wb_dat_o_reg[0] ,
    \\wb_dat_o_reg[1] , \\wb_dat_o_reg[6] , \\wb_dat_o_reg[2] ,
    \\wb_dat_o_reg[10] , \\wb_dat_o_reg[13] , \\wb_dat_o_reg[14] ,
    \\wb_dat_o_reg[12] , \\wb_dat_o_reg[8] , \\wb_dat_o_reg[15] ,
    \\wb_dat_o_reg[26] , \\wb_dat_o_reg[16] , \\wb_dat_o_reg[18] ,
    \\wb_dat_o_reg[17] , \\wb_dat_o_reg[19] , \\wb_dat_o_reg[22] ,
    \\wb_dat_o_reg[27] , \\wb_dat_o_reg[21] , \\wb_dat_o_reg[31] ,
    \\wb_dat_o_reg[28] , \\wb_dat_o_reg[24] , \\wb_dat_o_reg[23] ,
    \\wb_dat_o_reg[30] , \\wb_dat_o_reg[20] , \\wb_dat_o_reg[29] ,
    \\wb_dat_o_reg[25] , wb_ack_o_reg;
  wire \new_[321]_ , \new_[324]_ , \new_[325]_ , \new_[326]_ , \new_[327]_ ,
    \new_[328]_ , \new_[329]_ , \new_[330]_ , \new_[331]_ , \new_[332]_ ,
    \new_[333]_ , \new_[334]_ , \new_[335]_ , \new_[336]_ , \new_[337]_ ,
    \new_[338]_ , \new_[339]_ , \new_[340]_ , \new_[341]_ , \new_[342]_ ,
    \new_[343]_ , \new_[344]_ , \new_[345]_ , \new_[346]_ , \new_[347]_ ,
    \new_[348]_ , \new_[349]_ , \new_[350]_ , \new_[351]_ , \new_[352]_ ,
    \new_[353]_ , \new_[354]_ , \new_[355]_ , \new_[356]_ , \new_[357]_ ,
    \new_[358]_ , \new_[359]_ , \new_[360]_ , \new_[361]_ , \new_[362]_ ,
    \new_[363]_ , \new_[364]_ , \new_[365]_ , \new_[366]_ , \new_[367]_ ,
    \new_[368]_ , \new_[369]_ , \new_[370]_ , \new_[371]_ , \new_[372]_ ,
    \new_[373]_ , \new_[374]_ , \new_[375]_ , \new_[376]_ , \new_[377]_ ,
    \new_[378]_ , \new_[379]_ , \new_[380]_ , \new_[381]_ , \new_[382]_ ,
    \new_[383]_ , \new_[384]_ , \new_[385]_ , \new_[386]_ , \new_[387]_ ,
    \new_[388]_ , \new_[389]_ , \new_[390]_ , \new_[391]_ , \new_[392]_ ,
    \new_[393]_ , \new_[394]_ , \new_[424]_ , \new_[425]_ , \new_[426]_ ,
    \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ , \new_[431]_ ,
    \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ , \new_[436]_ ,
    \new_[437]_ , \new_[438]_ , \new_[439]_ , \new_[440]_ , \new_[441]_ ,
    \new_[442]_ , \new_[443]_ , \new_[444]_ , \new_[445]_ , \new_[446]_ ,
    \new_[447]_ , \new_[464]_ , \new_[465]_ , \new_[468]_ , \new_[474]_ ,
    \new_[482]_ , \new_[486]_ , \new_[488]_ , \new_[492]_ , \new_[493]_ ,
    \new_[494]_ , \new_[495]_ , \new_[496]_ , \new_[497]_ , \new_[498]_ ,
    \new_[499]_ , \new_[500]_ , \new_[501]_ , \new_[502]_ , \new_[503]_ ,
    \new_[504]_ , \new_[505]_ , \new_[506]_ , \new_[507]_ , \new_[508]_ ,
    \new_[509]_ , \new_[515]_ , \new_[517]_ , \new_[518]_ , \new_[519]_ ,
    \new_[520]_ , \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ ,
    \new_[525]_ , \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ ,
    \new_[530]_ , \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ ,
    \new_[535]_ , \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ ,
    \new_[540]_ , \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ ,
    \new_[545]_ , \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[557]_ ,
    \new_[558]_ , \new_[559]_ , \new_[560]_ , \new_[561]_ , \new_[562]_ ,
    \new_[578]_ , \new_[579]_ , \new_[580]_ , \new_[581]_ , \new_[582]_ ,
    \new_[583]_ , \new_[584]_ , \new_[585]_ , \new_[586]_ , \new_[587]_ ,
    \new_[588]_ , \new_[589]_ , \new_[590]_ , \new_[591]_ , \new_[592]_ ,
    \new_[593]_ , \new_[594]_ , \new_[595]_ , \new_[596]_ , \new_[597]_ ,
    \new_[598]_ , \new_[599]_ , \new_[600]_ , \new_[601]_ , \new_[602]_ ,
    \new_[603]_ , \new_[604]_ , \new_[605]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ , \new_[636]_ ,
    \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ , \new_[641]_ ,
    \new_[642]_ , \new_[643]_ , \new_[649]_ , \new_[650]_ , \new_[651]_ ,
    \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[655]_ , \new_[656]_ ,
    \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ , \new_[661]_ ,
    \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ , \new_[666]_ ,
    \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ , \new_[671]_ ,
    \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ , \new_[676]_ ,
    \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ , \new_[681]_ ,
    \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ , \new_[686]_ ,
    \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ , \new_[691]_ ,
    \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ , \new_[696]_ ,
    \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ , \new_[701]_ ,
    \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ , \new_[706]_ ,
    \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ , \new_[711]_ ,
    \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ , \new_[716]_ ,
    \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ , \new_[721]_ ,
    \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ , \new_[726]_ ,
    \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ , \new_[731]_ ,
    \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ , \new_[736]_ ,
    \new_[737]_ , \new_[738]_ , \new_[739]_ , \new_[740]_ , \new_[741]_ ,
    \new_[742]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ , \new_[746]_ ,
    \new_[747]_ , \new_[748]_ , \new_[749]_ , \new_[750]_ , \new_[751]_ ,
    \new_[752]_ , \new_[753]_ , \new_[754]_ , \new_[755]_ , \new_[756]_ ,
    \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ , \new_[761]_ ,
    \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ , \new_[766]_ ,
    \new_[767]_ , \new_[768]_ , \new_[769]_ , \new_[770]_ , \new_[771]_ ,
    \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ , \new_[776]_ ,
    \new_[777]_ , \new_[778]_ , \new_[779]_ , \new_[780]_ , \new_[781]_ ,
    \new_[782]_ , \new_[783]_ , \new_[784]_ , \new_[785]_ , \new_[786]_ ,
    \new_[787]_ , \new_[788]_ , \new_[789]_ , \new_[790]_ , \new_[791]_ ,
    \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ , \new_[796]_ ,
    \new_[797]_ , \new_[798]_ , \new_[799]_ , \new_[800]_ , \new_[801]_ ,
    \new_[802]_ , \new_[803]_ , \new_[804]_ , \new_[805]_ , \new_[806]_ ,
    \new_[807]_ , \new_[808]_ , \new_[809]_ , \new_[810]_ , \new_[811]_ ,
    \new_[812]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ , \new_[816]_ ,
    \new_[817]_ , \new_[818]_ , \new_[819]_ , \new_[820]_ , \new_[821]_ ,
    \new_[822]_ , \new_[823]_ , \new_[824]_ , \new_[825]_ , \new_[826]_ ,
    \new_[827]_ , \new_[828]_ , \new_[829]_ , \new_[830]_ , \new_[831]_ ,
    \new_[832]_ , \new_[833]_ , \new_[834]_ , \new_[835]_ , \new_[836]_ ,
    \new_[837]_ , \new_[838]_ , \new_[839]_ , \new_[840]_ , \new_[841]_ ,
    \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[845]_ , \new_[846]_ ,
    \new_[847]_ , \new_[848]_ , \new_[849]_ , \new_[850]_ , \new_[851]_ ,
    \new_[852]_ , \new_[853]_ , \new_[854]_ , \new_[855]_ , \new_[856]_ ,
    \new_[857]_ , \new_[858]_ , \new_[859]_ , \new_[860]_ , \new_[861]_ ,
    \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[865]_ , \new_[866]_ ,
    \new_[867]_ , \new_[868]_ , \new_[869]_ , \new_[870]_ , \new_[871]_ ,
    \new_[872]_ , \new_[873]_ , \new_[874]_ , \new_[875]_ , \new_[876]_ ,
    \new_[877]_ , \new_[878]_ , \new_[879]_ , \new_[880]_ , \new_[881]_ ,
    \new_[882]_ , \new_[883]_ , \new_[884]_ , \new_[885]_ , \new_[886]_ ,
    \new_[887]_ , \new_[888]_ , \new_[889]_ , \new_[890]_ , \new_[891]_ ,
    \new_[892]_ , \new_[893]_ , \new_[894]_ , \new_[895]_ , \new_[896]_ ,
    \new_[897]_ , \new_[898]_ , \new_[899]_ , \new_[900]_ , \new_[901]_ ,
    \new_[902]_ , \new_[903]_ , \new_[904]_ , \new_[905]_ , \new_[906]_ ,
    \new_[907]_ , \new_[908]_ , \new_[909]_ , \new_[910]_ , \new_[911]_ ,
    \new_[912]_ , \new_[913]_ , \new_[914]_ , \new_[915]_ , \new_[916]_ ,
    \new_[917]_ , \new_[918]_ , \new_[919]_ , \new_[920]_ , \new_[921]_ ,
    \new_[922]_ , \new_[923]_ , \new_[924]_ , \new_[925]_ , \new_[926]_ ,
    \new_[927]_ , \new_[928]_ , \new_[929]_ , \new_[930]_ , \new_[931]_ ,
    \new_[932]_ , \new_[933]_ , \new_[934]_ , \new_[935]_ , \new_[936]_ ,
    \new_[937]_ , \new_[938]_ , \new_[939]_ , \new_[940]_ , \new_[941]_ ,
    \new_[942]_ , \new_[943]_ , \new_[944]_ , \new_[945]_ , \new_[946]_ ,
    \new_[947]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ , \new_[951]_ ,
    \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[955]_ , \new_[956]_ ,
    \new_[957]_ , \new_[958]_ , \new_[959]_ , \new_[960]_ , \new_[961]_ ,
    \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ , \new_[966]_ ,
    \new_[967]_ , \new_[968]_ , \new_[969]_ , \new_[970]_ , \new_[971]_ ,
    \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[975]_ , \new_[976]_ ,
    \new_[977]_ , \new_[978]_ , \new_[979]_ , \new_[980]_ , \new_[981]_ ,
    \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ , \new_[986]_ ,
    \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ , \new_[991]_ ,
    \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ , \new_[996]_ ,
    \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ , \new_[1001]_ ,
    \new_[1002]_ , \new_[1003]_ , \new_[1004]_ , \new_[1005]_ ,
    \new_[1006]_ , \new_[1007]_ , \new_[1008]_ , \new_[1009]_ ,
    \new_[1010]_ , \new_[1011]_ , \new_[1012]_ , \new_[1013]_ ,
    \new_[1014]_ , \new_[1015]_ , \new_[1016]_ , \new_[1017]_ ,
    \new_[1018]_ , \new_[1019]_ , \new_[1020]_ , \new_[1021]_ ,
    \new_[1022]_ , \new_[1023]_ , \new_[1024]_ , \new_[1025]_ ,
    \new_[1026]_ , \new_[1027]_ , \new_[1028]_ , \new_[1029]_ ,
    \new_[1030]_ , \new_[1031]_ , \new_[1032]_ , \new_[1033]_ ,
    \new_[1034]_ , \new_[1035]_ , \new_[1036]_ , \new_[1037]_ ,
    \new_[1038]_ , \new_[1039]_ , \new_[1040]_ , \new_[1041]_ ,
    \new_[1042]_ , \new_[1043]_ , \new_[1044]_ , \new_[1045]_ ,
    \new_[1046]_ , \new_[1047]_ , \new_[1048]_ , \new_[1049]_ ,
    \new_[1050]_ , \new_[1051]_ , \new_[1052]_ , \new_[1053]_ ,
    \new_[1054]_ , \new_[1055]_ , \new_[1056]_ , \new_[1057]_ ,
    \new_[1058]_ , \new_[1059]_ , \new_[1060]_ , \new_[1061]_ ,
    \new_[1062]_ , \new_[1063]_ , \new_[1064]_ , \new_[1065]_ ,
    \new_[1066]_ , \new_[1067]_ , \new_[1068]_ , \new_[1069]_ ,
    \new_[1070]_ , \new_[1071]_ , \new_[1072]_ , \new_[1073]_ ,
    \new_[1074]_ , \new_[1075]_ , \new_[1076]_ , \new_[1077]_ ,
    \new_[1078]_ , \new_[1079]_ , \new_[1080]_ , \new_[1081]_ ,
    \new_[1082]_ , \new_[1083]_ , \new_[1084]_ , \new_[1085]_ ,
    \new_[1086]_ , \new_[1087]_ , \new_[1088]_ , \new_[1089]_ ,
    \new_[1090]_ , \new_[1091]_ , \new_[1092]_ , \new_[1093]_ ,
    \new_[1094]_ , \new_[1095]_ , \new_[1096]_ , \new_[1097]_ ,
    \new_[1098]_ , \new_[1099]_ , \new_[1100]_ , \new_[1101]_ ,
    \new_[1102]_ , \new_[1103]_ , \new_[1104]_ , \new_[1105]_ ,
    \new_[1106]_ , \new_[1107]_ , \new_[1108]_ , \new_[1109]_ ,
    \new_[1110]_ , \new_[1111]_ , \new_[1112]_ , \new_[1113]_ ,
    \new_[1114]_ , \new_[1115]_ , \new_[1116]_ , \new_[1117]_ ,
    \new_[1118]_ , \new_[1119]_ , \new_[1120]_ , \new_[1121]_ ,
    \new_[1122]_ , \new_[1123]_ , \new_[1124]_ , \new_[1125]_ ,
    \new_[1126]_ , \new_[1127]_ , \new_[1128]_ , \new_[1129]_ ,
    \new_[1130]_ , \new_[1131]_ , \new_[1132]_ , \new_[1133]_ ,
    \new_[1134]_ , \new_[1135]_ , \new_[1136]_ , \new_[1137]_ ,
    \new_[1138]_ , \new_[1139]_ , \new_[1140]_ , \new_[1141]_ ,
    \new_[1142]_ , \new_[1143]_ , \new_[1144]_ , \new_[1145]_ ,
    \new_[1146]_ , \new_[1147]_ , \new_[1148]_ , \new_[1149]_ ,
    \new_[1150]_ , \new_[1151]_ , \new_[1152]_ , \new_[1153]_ ,
    \new_[1154]_ , \new_[1155]_ , \new_[1156]_ , \new_[1157]_ ,
    \new_[1158]_ , \new_[1159]_ , \new_[1160]_ , \new_[1161]_ ,
    \new_[1162]_ , \new_[1163]_ , \new_[1164]_ , \new_[1165]_ ,
    \new_[1166]_ , \new_[1167]_ , \new_[1168]_ , \new_[1169]_ ,
    \new_[1170]_ , \new_[1171]_ , \new_[1172]_ , \new_[1173]_ ,
    \new_[1174]_ , \new_[1175]_ , \new_[1176]_ , \new_[1177]_ ,
    \new_[1178]_ , \new_[1179]_ , \new_[1180]_ , \new_[1181]_ ,
    \new_[1182]_ , \new_[1183]_ , \new_[1184]_ , \new_[1185]_ ,
    \new_[1186]_ , \new_[1187]_ , \new_[1188]_ , \new_[1190]_ ,
    \new_[1191]_ , \new_[1192]_ , \new_[1193]_ , \new_[1194]_ ,
    \new_[1195]_ , \new_[1196]_ , \new_[1197]_ , \new_[1198]_ ,
    \new_[1199]_ , \new_[1200]_ , \new_[1201]_ , \new_[1202]_ ,
    \new_[1203]_ , \new_[1204]_ , \new_[1205]_ , \new_[1206]_ ,
    \new_[1207]_ , \new_[1208]_ , \new_[1209]_ , \new_[1210]_ ,
    \new_[1211]_ , \new_[1212]_ , \new_[1213]_ , \new_[1214]_ ,
    \new_[1215]_ , \new_[1216]_ , \new_[1217]_ , \new_[1218]_ ,
    \new_[1219]_ , \new_[1220]_ , \new_[1221]_ , \new_[1222]_ ,
    \new_[1223]_ , \new_[1224]_ , \new_[1225]_ , \new_[1226]_ ,
    \new_[1227]_ , \new_[1228]_ , \new_[1229]_ , \new_[1230]_ ,
    \new_[1231]_ , \new_[1232]_ , \new_[1233]_ , \new_[1234]_ ,
    \new_[1235]_ , \new_[1236]_ , \new_[1237]_ , \new_[1238]_ ,
    \new_[1239]_ , \new_[1240]_ , \new_[1241]_ , \new_[1242]_ ,
    \new_[1243]_ , \new_[1244]_ , \new_[1245]_ , \new_[1246]_ ,
    \new_[1247]_ , \new_[1248]_ , \new_[1249]_ , \new_[1250]_ ,
    \new_[1251]_ , \new_[1252]_ , \new_[1253]_ , \new_[1254]_ ,
    \new_[1255]_ , \new_[1256]_ , \new_[1257]_ , \new_[1258]_ ,
    \new_[1259]_ , \new_[1260]_ , \new_[1261]_ , \new_[1262]_ ,
    \new_[1263]_ , \new_[1264]_ , \new_[1265]_ , \new_[1266]_ ,
    \new_[1267]_ , \new_[1268]_ , \new_[1269]_ , \new_[1270]_ ,
    \new_[1271]_ , \new_[1272]_ , \new_[1273]_ , \new_[1274]_ ,
    \new_[1275]_ , \new_[1276]_ , \new_[1277]_ , \new_[1278]_ ,
    \new_[1279]_ , \new_[1280]_ , \new_[1281]_ , \new_[1282]_ ,
    \new_[1283]_ , \new_[1284]_ , \new_[1285]_ , \new_[1286]_ ,
    \new_[1287]_ , \new_[1288]_ , \new_[1289]_ , \new_[1290]_ ,
    \new_[1291]_ , \new_[1292]_ , \new_[1293]_ , \new_[1294]_ ,
    \new_[1295]_ , \new_[1296]_ , \new_[1297]_ , \new_[1298]_ ,
    \new_[1299]_ , \new_[1300]_ , \new_[1301]_ , \new_[1302]_ ,
    \new_[1303]_ , \new_[1304]_ , \new_[1305]_ , \new_[1306]_ ,
    \new_[1307]_ , \new_[1308]_ , \new_[1309]_ , \new_[1310]_ ,
    \new_[1311]_ , \new_[1312]_ , \new_[1314]_ , \new_[1315]_ ,
    \new_[1316]_ , \new_[1317]_ , \new_[1318]_ , \new_[1319]_ ,
    \new_[1320]_ , \new_[1321]_ , \new_[1322]_ , \new_[1323]_ ,
    \new_[1324]_ , \new_[1325]_ , \new_[1326]_ , \new_[1327]_ ,
    \new_[1328]_ , \new_[1329]_ , \new_[1330]_ , \new_[1331]_ ,
    \new_[1332]_ , \new_[1333]_ , \new_[1334]_ , \new_[1335]_ ,
    \new_[1336]_ , \new_[1337]_ , \new_[1338]_ , \new_[1339]_ ,
    \new_[1340]_ , \new_[1341]_ , \new_[1342]_ , \new_[1343]_ ,
    \new_[1344]_ , \new_[1345]_ , \new_[1346]_ , \new_[1347]_ ,
    \new_[1348]_ , \new_[1349]_ , \new_[1350]_ , \new_[1351]_ ,
    \new_[1352]_ , \new_[1353]_ , \new_[1354]_ , \new_[1355]_ ,
    \new_[1356]_ , \new_[1357]_ , \new_[1358]_ , \new_[1359]_ ,
    \new_[1360]_ , \new_[1361]_ , \new_[1362]_ , \new_[1363]_ ,
    \new_[1364]_ , \new_[1365]_ , \new_[1366]_ , \new_[1367]_ ,
    \new_[1368]_ , \new_[1369]_ , \new_[1370]_ , \new_[1371]_ ,
    \new_[1372]_ , \new_[1373]_ , \new_[1374]_ , \new_[1375]_ ,
    \new_[1376]_ , \new_[1377]_ , \new_[1378]_ , \new_[1379]_ ,
    \new_[1380]_ , \new_[1381]_ , \new_[1382]_ , \new_[1383]_ ,
    \new_[1384]_ , \new_[1385]_ , \new_[1386]_ , \new_[1387]_ ,
    \new_[1388]_ , \new_[1389]_ , \new_[1390]_ , \new_[1391]_ ,
    \new_[1392]_ , \new_[1393]_ , \new_[1394]_ , \new_[1395]_ ,
    \new_[1396]_ , \new_[1397]_ , \new_[1398]_ , \new_[1399]_ ,
    \new_[1400]_ , \new_[1401]_ , \new_[1402]_ , \new_[1403]_ ,
    \new_[1404]_ , \new_[1405]_ , \new_[1406]_ , \new_[1407]_ ,
    \new_[1408]_ , \new_[1409]_ , \new_[1410]_ , \new_[1411]_ ,
    \new_[1412]_ , \new_[1413]_ , \new_[1414]_ , \new_[1415]_ ,
    \new_[1416]_ , \new_[1417]_ , \new_[1418]_ , \new_[1419]_ ,
    \new_[1420]_ , \new_[1421]_ , \new_[1422]_ , \new_[1423]_ ,
    \new_[1424]_ , \new_[1425]_ , \new_[1426]_ , \new_[1427]_ ,
    \new_[1428]_ , \new_[1429]_ , \new_[1430]_ , \new_[1431]_ ,
    \new_[1432]_ , \new_[1433]_ , \new_[1434]_ , \new_[1435]_ ,
    \new_[1436]_ , \new_[1437]_ , \new_[1438]_ , \new_[1439]_ ,
    \new_[1440]_ , \new_[1441]_ , \new_[1442]_ , \new_[1443]_ ,
    \new_[1444]_ , \new_[1445]_ , \new_[1446]_ , \new_[1447]_ ,
    \new_[1448]_ , \new_[1449]_ , \new_[1450]_ , \new_[1451]_ ,
    \new_[1452]_ , \new_[1453]_ , \new_[1454]_ , \new_[1455]_ ,
    \new_[1456]_ , \new_[1457]_ , \new_[1458]_ , \new_[1459]_ ,
    \new_[1460]_ , \new_[1461]_ , \new_[1462]_ , \new_[1463]_ ,
    \new_[1464]_ , \new_[1465]_ , \new_[1466]_ , \new_[1467]_ ,
    \new_[1468]_ , \new_[1469]_ , \new_[1470]_ , \new_[1471]_ ,
    \new_[1472]_ , \new_[1473]_ , \new_[1474]_ , \new_[1475]_ ,
    \new_[1476]_ , \new_[1477]_ , \new_[1478]_ , \new_[1479]_ ,
    \new_[1480]_ , \new_[1481]_ , \new_[1482]_ , \new_[1483]_ ,
    \new_[1484]_ , \new_[1485]_ , \new_[1486]_ , \new_[1487]_ ,
    \new_[1488]_ , \new_[1489]_ , \new_[1490]_ , \new_[1491]_ ,
    \new_[1492]_ , \new_[1493]_ , \new_[1494]_ , \new_[1495]_ ,
    \new_[1496]_ , \new_[1497]_ , \new_[1498]_ , \new_[1499]_ ,
    \new_[1500]_ , \new_[1501]_ , \new_[1502]_ , \new_[1503]_ ,
    \new_[1504]_ , \new_[1505]_ , \new_[1506]_ , \new_[1507]_ ,
    \new_[1508]_ , \new_[1509]_ , \new_[1510]_ , \new_[1511]_ ,
    \new_[1512]_ , \new_[1513]_ , \new_[1514]_ , \new_[1515]_ ,
    \new_[1516]_ , \new_[1517]_ , \new_[1518]_ , \new_[1519]_ ,
    \new_[1520]_ , \new_[1521]_ , \new_[1522]_ , \new_[1523]_ ,
    \new_[1524]_ , \new_[1525]_ , \new_[1526]_ , \new_[1527]_ ,
    \new_[1528]_ , \new_[1529]_ , \new_[1530]_ , \new_[1531]_ ,
    \new_[1532]_ , \new_[1533]_ , \new_[1534]_ , \new_[1535]_ ,
    \new_[1536]_ , \new_[1537]_ , \new_[1538]_ , \new_[1539]_ ,
    \new_[1540]_ , \new_[1541]_ , \new_[1542]_ , \new_[1543]_ ,
    \new_[1544]_ , \new_[1545]_ , \new_[1546]_ , \new_[1547]_ ,
    \new_[1548]_ , \new_[1549]_ , \new_[1550]_ , \new_[1551]_ ,
    \new_[1552]_ , \new_[1553]_ , \new_[1555]_ , \new_[1556]_ ,
    \new_[1557]_ , \new_[1558]_ , \new_[1559]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1562]_ , \new_[1563]_ , \new_[1564]_ ,
    \new_[1565]_ , \new_[1566]_ , \new_[1567]_ , \new_[1568]_ ,
    \new_[1569]_ , \new_[1570]_ , \new_[1571]_ , \new_[1572]_ ,
    \new_[1573]_ , \new_[1574]_ , \new_[1575]_ , \new_[1576]_ ,
    \new_[1577]_ , \new_[1578]_ , \new_[1579]_ , \new_[1580]_ ,
    \new_[1581]_ , \new_[1582]_ , \new_[1583]_ , \new_[1584]_ ,
    \new_[1585]_ , \new_[1586]_ , \new_[1587]_ , \new_[1588]_ ,
    \new_[1589]_ , \new_[1590]_ , \new_[1591]_ , \new_[1592]_ ,
    \new_[1593]_ , \new_[1595]_ , \new_[1596]_ , \new_[1597]_ ,
    \new_[1600]_ , \new_[1601]_ , \new_[1602]_ , \new_[1603]_ ,
    \new_[1604]_ , \new_[1605]_ , \new_[1606]_ , \new_[1607]_ ,
    \new_[1608]_ , \new_[1609]_ , \new_[1610]_ , \new_[1611]_ ,
    \new_[1613]_ , \new_[1614]_ , \new_[1615]_ , \new_[1617]_ ,
    \new_[1618]_ , \new_[1619]_ , \new_[1620]_ , \new_[1621]_ ,
    \new_[1622]_ , \new_[1623]_ , \new_[1624]_ , \new_[1625]_ ,
    \new_[1626]_ , \new_[1627]_ , \new_[1628]_ , \new_[1629]_ ,
    \new_[1630]_ , \new_[1631]_ , \new_[1632]_ , \new_[1633]_ ,
    \new_[1634]_ , \new_[1635]_ , \new_[1636]_ , \new_[1637]_ ,
    \new_[1638]_ , \new_[1639]_ , \new_[1640]_ , \new_[1641]_ ,
    \new_[1642]_ , \new_[1643]_ , \new_[1644]_ , \new_[1645]_ ,
    \new_[1646]_ , \new_[1647]_ , \new_[1648]_ , \new_[1649]_ ,
    \new_[1650]_ , \new_[1651]_ , \new_[1652]_ , \new_[1653]_ ,
    \new_[1654]_ , \new_[1655]_ , \new_[1656]_ , \new_[1657]_ ,
    \new_[1658]_ , \new_[1659]_ , \new_[1660]_ , \new_[1662]_ ,
    \new_[1663]_ , \new_[1664]_ , \new_[1665]_ , \new_[1667]_ ,
    \new_[1668]_ , \new_[1669]_ , \new_[1670]_ , \new_[1671]_ ,
    \new_[1672]_ , \new_[1674]_ , \new_[1675]_ , \new_[1676]_ ,
    \new_[1677]_ , \new_[1678]_ , \new_[1679]_ , \new_[1680]_ ,
    \new_[1681]_ , \new_[1682]_ , \new_[1683]_ , \new_[1684]_ ,
    \new_[1685]_ , \new_[1686]_ , \new_[1687]_ , \new_[1688]_ ,
    \new_[1689]_ , \new_[1690]_ , \new_[1691]_ , \new_[1692]_ ,
    \new_[1693]_ , \new_[1694]_ , \new_[1695]_ , \new_[1696]_ ,
    \new_[1697]_ , \new_[1699]_ , \new_[1700]_ , \new_[1701]_ ,
    \new_[1702]_ , \new_[1703]_ , \new_[1704]_ , \new_[1705]_ ,
    \new_[1706]_ , \new_[1708]_ , \new_[1709]_ , \new_[1710]_ ,
    \new_[1711]_ , \new_[1712]_ , \new_[1713]_ , \new_[1714]_ ,
    \new_[1715]_ , \new_[1716]_ , \new_[1717]_ , \new_[1718]_ ,
    \new_[1719]_ , \new_[1720]_ , \new_[1721]_ , \new_[1722]_ ,
    \new_[1723]_ , \new_[1724]_ , \new_[1725]_ , \new_[1726]_ ,
    \new_[1727]_ , \new_[1728]_ , \new_[1729]_ , \new_[1730]_ ,
    \new_[1731]_ , \new_[1732]_ , \new_[1733]_ , \new_[1734]_ ,
    \new_[1735]_ , \new_[1736]_ , \new_[1737]_ , \new_[1738]_ ,
    \new_[1739]_ , \new_[1740]_ , \new_[1741]_ , \new_[1742]_ ,
    \new_[1743]_ , \new_[1744]_ , \new_[1745]_ , \new_[1746]_ ,
    \new_[1747]_ , \new_[1748]_ , \new_[1749]_ , \new_[1750]_ ,
    \new_[1751]_ , \new_[1752]_ , \new_[1753]_ , \new_[1754]_ ,
    \new_[1755]_ , \new_[1756]_ , \new_[1757]_ , \new_[1758]_ ,
    \new_[1759]_ , \new_[1760]_ , \new_[1761]_ , \new_[1762]_ ,
    \new_[1763]_ , \new_[1764]_ , \new_[1765]_ , \new_[1766]_ ,
    \new_[1768]_ , \new_[1769]_ , \new_[1770]_ , \new_[1771]_ ,
    \new_[1772]_ , \new_[1773]_ , \new_[1774]_ , \new_[1775]_ ,
    \new_[1776]_ , \new_[1777]_ , \new_[1780]_ , \new_[1781]_ ,
    \new_[1782]_ , \new_[1785]_ , \new_[1787]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1791]_ , \new_[1792]_ ,
    \new_[1793]_ , \new_[1794]_ , \new_[1795]_ , \new_[1796]_ ,
    \new_[1797]_ , \new_[1798]_ , \new_[1799]_ , \new_[1800]_ ,
    \new_[1801]_ , \new_[1802]_ , \new_[1803]_ , \new_[1804]_ ,
    \new_[1805]_ , \new_[1806]_ , \new_[1807]_ , \new_[1808]_ ,
    \new_[1809]_ , \new_[1810]_ , \new_[1811]_ , \new_[1812]_ ,
    \new_[1813]_ , \new_[1814]_ , \new_[1815]_ , \new_[1816]_ ,
    \new_[1817]_ , \new_[1818]_ , \new_[1819]_ , \new_[1820]_ ,
    \new_[1821]_ , \new_[1822]_ , \new_[1823]_ , \new_[1824]_ ,
    \new_[1825]_ , \new_[1826]_ , \new_[1827]_ , \new_[1828]_ ,
    \new_[1830]_ , \new_[1831]_ , \new_[1832]_ , \new_[1833]_ ,
    \new_[1834]_ , \new_[1835]_ , \new_[1836]_ , \new_[1837]_ ,
    \new_[1838]_ , \new_[1839]_ , \new_[1840]_ , \new_[1841]_ ,
    \new_[1842]_ , \new_[1843]_ , \new_[1844]_ , \new_[1846]_ ,
    \new_[1847]_ , \new_[1848]_ , \new_[1849]_ , \new_[1850]_ ,
    \new_[1851]_ , \new_[1852]_ , \new_[1853]_ , \new_[1854]_ ,
    \new_[1855]_ , \new_[1856]_ , \new_[1857]_ , \new_[1858]_ ,
    \new_[1859]_ , \new_[1860]_ , \new_[1861]_ , \new_[1862]_ ,
    \new_[1863]_ , \new_[1864]_ , \new_[1865]_ , \new_[1866]_ ,
    \new_[1867]_ , \new_[1868]_ , \new_[1869]_ , \new_[1870]_ ,
    \new_[1871]_ , \new_[1872]_ , \new_[1873]_ , \new_[1874]_ ,
    \new_[1875]_ , \new_[1876]_ , \new_[1877]_ , \new_[1878]_ ,
    \new_[1879]_ , \new_[1880]_ , \new_[1881]_ , \new_[1882]_ ,
    \new_[1883]_ , \new_[1884]_ , \new_[1885]_ , \new_[1886]_ ,
    \new_[1887]_ , \new_[1888]_ , \new_[1889]_ , \new_[1891]_ ,
    \new_[1892]_ , \new_[1893]_ , \new_[1894]_ , \new_[1895]_ ,
    \new_[1896]_ , \new_[1897]_ , \new_[1898]_ , \new_[1899]_ ,
    \new_[1900]_ , \new_[1901]_ , \new_[1902]_ , \new_[1903]_ ,
    \new_[1904]_ , \new_[1905]_ , \new_[1906]_ , \new_[1907]_ ,
    \new_[1908]_ , \new_[1909]_ , \new_[1910]_ , \new_[1911]_ ,
    \new_[1912]_ , \new_[1913]_ , \new_[1914]_ , \new_[1915]_ ,
    \new_[1916]_ , \new_[1917]_ , \new_[1918]_ , \new_[1919]_ ,
    \new_[1920]_ , \new_[1921]_ , \new_[1922]_ , \new_[1923]_ ,
    \new_[1924]_ , \new_[1925]_ , \new_[1926]_ , \new_[1927]_ ,
    \new_[1928]_ , \new_[1929]_ , \new_[1930]_ , \new_[1931]_ ,
    \new_[1932]_ , \new_[1933]_ , \new_[1934]_ , \new_[1935]_ ,
    \new_[1936]_ , \new_[1937]_ , \new_[1938]_ , \new_[1939]_ ,
    \new_[1940]_ , \new_[1941]_ , \new_[1942]_ , \new_[1943]_ ,
    \new_[1944]_ , \new_[1945]_ , \new_[1946]_ , \new_[1947]_ ,
    \new_[1948]_ , \new_[1949]_ , \new_[1950]_ , \new_[1951]_ ,
    \new_[1954]_ , \new_[1955]_ , \new_[1956]_ , \new_[1957]_ ,
    \new_[1958]_ , \new_[1959]_ , \new_[1960]_ , \new_[1961]_ ,
    \new_[1962]_ , \new_[1963]_ , \new_[1964]_ , \new_[1965]_ ,
    \new_[1966]_ , \new_[1967]_ , \new_[1968]_ , \new_[1969]_ ,
    \new_[1970]_ , \new_[1971]_ , \new_[1972]_ , \new_[1973]_ ,
    \new_[1974]_ , \new_[1975]_ , \new_[1976]_ , \new_[1977]_ ,
    \new_[1978]_ , \new_[1979]_ , \new_[1980]_ , \new_[1981]_ ,
    \new_[1982]_ , \new_[1983]_ , \new_[1984]_ , \new_[1985]_ ,
    \new_[1986]_ , \new_[1987]_ , \new_[1988]_ , \new_[1989]_ ,
    \new_[1990]_ , \new_[1991]_ , \new_[1992]_ , \new_[1993]_ ,
    \new_[1994]_ , \new_[1995]_ , \new_[1996]_ , \new_[1997]_ ,
    \new_[1998]_ , \new_[1999]_ , \new_[2000]_ , \new_[2001]_ ,
    \new_[2002]_ , \new_[2003]_ , \new_[2004]_ , \new_[2005]_ ,
    \new_[2006]_ , \new_[2007]_ , \new_[2008]_ , \new_[2009]_ ,
    \new_[2010]_ , \new_[2011]_ , \new_[2012]_ , \new_[2013]_ ,
    \new_[2014]_ , \new_[2015]_ , \new_[2016]_ , \new_[2017]_ ,
    \new_[2018]_ , \new_[2019]_ , \new_[2020]_ , \new_[2021]_ ,
    \new_[2022]_ , \new_[2023]_ , \new_[2025]_ , \new_[2026]_ ,
    \new_[2027]_ , \new_[2029]_ , \new_[2032]_ , \new_[2033]_ ,
    \new_[2035]_ , \new_[2036]_ , \new_[2037]_ , \new_[2038]_ ,
    \new_[2039]_ , \new_[2040]_ , \new_[2041]_ , \new_[2042]_ ,
    \new_[2043]_ , \new_[2044]_ , \new_[2045]_ , \new_[2046]_ ,
    \new_[2047]_ , \new_[2048]_ , \new_[2049]_ , \new_[2050]_ ,
    \new_[2051]_ , \new_[2052]_ , \new_[2053]_ , \new_[2054]_ ,
    \new_[2055]_ , \new_[2056]_ , \new_[2057]_ , \new_[2058]_ ,
    \new_[2059]_ , \new_[2060]_ , \new_[2061]_ , \new_[2062]_ ,
    \new_[2063]_ , \new_[2064]_ , \new_[2065]_ , \new_[2066]_ ,
    \new_[2067]_ , \new_[2068]_ , \new_[2069]_ , \new_[2070]_ ,
    \new_[2071]_ , \new_[2072]_ , \new_[2073]_ , \new_[2074]_ ,
    \new_[2075]_ , \new_[2076]_ , \new_[2077]_ , \new_[2081]_ ,
    \new_[2082]_ , \new_[2083]_ , \new_[2084]_ , \new_[2085]_ ,
    \new_[2086]_ , \new_[2087]_ , \new_[2088]_ , \new_[2089]_ ,
    \new_[2090]_ , \new_[2091]_ , \new_[2092]_ , \new_[2093]_ ,
    \new_[2094]_ , \new_[2095]_ , \new_[2096]_ , \new_[2097]_ ,
    \new_[2098]_ , \new_[2099]_ , \new_[2100]_ , \new_[2101]_ ,
    \new_[2102]_ , \new_[2103]_ , \new_[2104]_ , \new_[2105]_ ,
    \new_[2106]_ , \new_[2107]_ , \new_[2108]_ , \new_[2109]_ ,
    \new_[2110]_ , \new_[2111]_ , \new_[2112]_ , \new_[2113]_ ,
    \new_[2114]_ , \new_[2115]_ , \new_[2116]_ , \new_[2117]_ ,
    \new_[2118]_ , \new_[2119]_ , \new_[2120]_ , \new_[2121]_ ,
    \new_[2122]_ , \new_[2123]_ , \new_[2124]_ , \new_[2125]_ ,
    \new_[2126]_ , \new_[2129]_ , \new_[2130]_ , \new_[2131]_ ,
    \new_[2133]_ , \new_[2135]_ , \new_[2136]_ , \new_[2137]_ ,
    \new_[2138]_ , \new_[2139]_ , \new_[2140]_ , \new_[2141]_ ,
    \new_[2148]_ , \new_[2149]_ , \new_[2150]_ , \new_[2151]_ ,
    \new_[2152]_ , \new_[2177]_ , \new_[2178]_ , \new_[2179]_ ,
    \new_[2180]_ , \new_[2181]_ , \new_[2182]_ , \new_[2183]_ ,
    \new_[2184]_ , \new_[2185]_ , \new_[2186]_ , \new_[2187]_ ,
    \new_[2188]_ , \new_[2189]_ , \new_[2190]_ , \new_[2191]_ ,
    \new_[2192]_ , \new_[2193]_ , \new_[2194]_ , \new_[2195]_ ,
    \new_[2196]_ , \new_[2197]_ , \new_[2198]_ , \new_[2199]_ ,
    \new_[2200]_ , \new_[2201]_ , \new_[2202]_ , \new_[2204]_ ,
    \new_[2205]_ , \new_[2209]_ , \new_[2210]_ , \new_[2214]_ ,
    \new_[2215]_ , \new_[2216]_ , \new_[2217]_ , \new_[2219]_ ,
    \new_[2222]_ , \new_[2223]_ , \new_[2225]_ , \new_[2226]_ ,
    \new_[2227]_ , \new_[2228]_ , \new_[2229]_ , \new_[2230]_ ,
    \new_[2231]_ , \new_[2232]_ , \new_[2233]_ , \new_[2234]_ ,
    \new_[2235]_ , \new_[2236]_ , \new_[2237]_ , \new_[2238]_ ,
    \new_[2239]_ , \new_[2240]_ , \new_[2241]_ , \new_[2242]_ ,
    \new_[2243]_ , \new_[2244]_ , \new_[2245]_ , \new_[2246]_ ,
    \new_[2247]_ , \new_[2249]_ , \new_[2250]_ , \new_[2251]_ ,
    \new_[2252]_ , \new_[2253]_ , \new_[2254]_ , \new_[2255]_ ,
    \new_[2256]_ , \new_[2257]_ , \new_[2258]_ , \new_[2259]_ ,
    \new_[2260]_ , \new_[2261]_ , \new_[2262]_ , \new_[2263]_ ,
    \new_[2264]_ , \new_[2265]_ , \new_[2266]_ , \new_[2267]_ ,
    \new_[2268]_ , \new_[2269]_ , \new_[2270]_ , \new_[2271]_ ,
    \new_[2272]_ , \new_[2273]_ , \new_[2274]_ , \new_[2275]_ ,
    \new_[2276]_ , \new_[2277]_ , \new_[2278]_ , \new_[2279]_ ,
    \new_[2280]_ , \new_[2281]_ , \new_[2282]_ , \new_[2283]_ ,
    \new_[2284]_ , \new_[2285]_ , \new_[2286]_ , \new_[2292]_ ,
    \new_[2293]_ , \new_[2294]_ , \new_[2295]_ , \new_[2296]_ ,
    \new_[2297]_ , \new_[2298]_ , \new_[2299]_ , \new_[2300]_ ,
    \new_[2301]_ , \new_[2302]_ , \new_[2303]_ , \new_[2304]_ ,
    \new_[2305]_ , \new_[2306]_ , \new_[2307]_ , \new_[2308]_ ,
    \new_[2309]_ , \new_[2318]_ , \new_[2319]_ , \new_[2320]_ ,
    \new_[2321]_ , \new_[2322]_ , \new_[2323]_ , \new_[2324]_ ,
    \new_[2325]_ , \new_[2326]_ , \new_[2327]_ , \new_[2328]_ ,
    \new_[2329]_ , \new_[2330]_ , \new_[2331]_ , \new_[2332]_ ,
    \new_[2333]_ , \new_[2334]_ , \new_[2335]_ , \new_[2336]_ ,
    \new_[2337]_ , \new_[2338]_ , \new_[2339]_ , \new_[2340]_ ,
    \new_[2341]_ , \new_[2342]_ , \new_[2343]_ , \new_[2344]_ ,
    \new_[2345]_ , \new_[2346]_ , \new_[2347]_ , \new_[2348]_ ,
    \new_[2349]_ , \new_[2350]_ , \new_[2351]_ , \new_[2352]_ ,
    \new_[2353]_ , \new_[2354]_ , \new_[2355]_ , \new_[2356]_ ,
    \new_[2357]_ , \new_[2358]_ , \new_[2359]_ , \new_[2360]_ ,
    \new_[2361]_ , \new_[2362]_ , \new_[2363]_ , \new_[2364]_ ,
    \new_[2365]_ , \new_[2366]_ , \new_[2367]_ , \new_[2368]_ ,
    \new_[2369]_ , \new_[2370]_ , \new_[2371]_ , \new_[2372]_ ,
    \new_[2373]_ , \new_[2374]_ , \new_[2375]_ , \new_[2376]_ ,
    \new_[2377]_ , \new_[2378]_ , \new_[2379]_ , \new_[2380]_ ,
    \new_[2381]_ , \new_[2383]_ , \new_[2384]_ , \new_[2385]_ ,
    \new_[2386]_ , \new_[2387]_ , \new_[2388]_ , \new_[2389]_ ,
    \new_[2395]_ , \new_[2396]_ , \new_[2397]_ , \new_[2398]_ ,
    \new_[2399]_ , \new_[2400]_ , \new_[2401]_ , \new_[2402]_ ,
    \new_[2403]_ , \new_[2404]_ , \new_[2405]_ , \new_[2406]_ ,
    \new_[2407]_ , \new_[2408]_ , \new_[2409]_ , \new_[2410]_ ,
    \new_[2411]_ , \new_[2412]_ , \new_[2413]_ , \new_[2414]_ ,
    \new_[2415]_ , \new_[2416]_ , \new_[2417]_ , \new_[2418]_ ,
    \new_[2419]_ , \new_[2420]_ , \new_[2421]_ , \new_[2422]_ ,
    \new_[2423]_ , \new_[2424]_ , \new_[2425]_ , \new_[2426]_ ,
    \new_[2427]_ , \new_[2428]_ , \new_[2429]_ , \new_[2430]_ ,
    \new_[2431]_ , \new_[2432]_ , \new_[2433]_ , \new_[2434]_ ,
    \new_[2435]_ , \new_[2436]_ , \new_[2437]_ , \new_[2438]_ ,
    \new_[2439]_ , \new_[2440]_ , \new_[2441]_ , \new_[2442]_ ,
    \new_[2443]_ , \new_[2444]_ , \new_[2445]_ , \new_[2446]_ ,
    \new_[2447]_ , \new_[2448]_ , \new_[2449]_ , \new_[2450]_ ,
    \new_[2451]_ , \new_[2452]_ , \new_[2453]_ , \new_[2454]_ ,
    \new_[2455]_ , \new_[2456]_ , \new_[2457]_ , \new_[2458]_ ,
    \new_[2459]_ , \new_[2460]_ , \new_[2461]_ , \new_[2462]_ ,
    \new_[2463]_ , \new_[2464]_ , \new_[2465]_ , \new_[2467]_ ,
    \new_[2468]_ , \new_[2469]_ , \new_[2470]_ , \new_[2471]_ ,
    \new_[2472]_ , \new_[2473]_ , \new_[2474]_ , \new_[2475]_ ,
    \new_[2476]_ , \new_[2477]_ , \new_[2478]_ , \new_[2479]_ ,
    \new_[2480]_ , \new_[2481]_ , \new_[2483]_ , \new_[2484]_ ,
    \new_[2487]_ , \new_[2488]_ , \new_[2489]_ , \new_[2491]_ ,
    \new_[2493]_ , \new_[2495]_ , \new_[2498]_ , \new_[2514]_ ,
    \new_[2515]_ , \new_[2516]_ , \new_[2519]_ , \new_[2520]_ ,
    \new_[2521]_ , \new_[2524]_ , \new_[2525]_ , \new_[2528]_ ,
    \new_[2529]_ , \new_[2530]_ , \new_[2531]_ , \new_[2532]_ ,
    \new_[2533]_ , \new_[2534]_ , \new_[2535]_ , \new_[2536]_ ,
    \new_[2537]_ , \new_[2538]_ , \new_[2539]_ , \new_[2540]_ ,
    \new_[2541]_ , \new_[2542]_ , \new_[2543]_ , \new_[2544]_ ,
    \new_[2545]_ , \new_[2546]_ , \new_[2547]_ , \new_[2548]_ ,
    \new_[2549]_ , \new_[2550]_ , \new_[2551]_ , \new_[2552]_ ,
    \new_[2553]_ , \new_[2554]_ , \new_[2555]_ , \new_[2556]_ ,
    \new_[2557]_ , \new_[2558]_ , \new_[2559]_ , \new_[2560]_ ,
    \new_[2561]_ , \new_[2562]_ , \new_[2563]_ , \new_[2564]_ ,
    \new_[2565]_ , \new_[2566]_ , \new_[2567]_ , \new_[2568]_ ,
    \new_[2569]_ , \new_[2570]_ , \new_[2571]_ , \new_[2572]_ ,
    \new_[2573]_ , \new_[2574]_ , \new_[2575]_ , \new_[2576]_ ,
    \new_[2577]_ , \new_[2578]_ , \new_[2579]_ , \new_[2580]_ ,
    \new_[2581]_ , \new_[2582]_ , \new_[2583]_ , \new_[2584]_ ,
    \new_[2585]_ , \new_[2586]_ , \new_[2587]_ , \new_[2588]_ ,
    \new_[2589]_ , \new_[2590]_ , \new_[2591]_ , \new_[2592]_ ,
    \new_[2593]_ , \new_[2594]_ , \new_[2595]_ , \new_[2596]_ ,
    \new_[2597]_ , \new_[2598]_ , \new_[2599]_ , \new_[2600]_ ,
    \new_[2601]_ , \new_[2602]_ , \new_[2612]_ , \new_[2617]_ ,
    \new_[2620]_ , \new_[2621]_ , \new_[2622]_ , \new_[2623]_ ,
    \new_[2624]_ , \new_[2625]_ , \new_[2626]_ , \new_[2627]_ ,
    \new_[2628]_ , \new_[2629]_ , \new_[2630]_ , \new_[2631]_ ,
    \new_[2632]_ , \new_[2633]_ , \new_[2634]_ , \new_[2635]_ ,
    \new_[2636]_ , \new_[2637]_ , \new_[2638]_ , \new_[2639]_ ,
    \new_[2640]_ , \new_[2641]_ , \new_[2642]_ , \new_[2643]_ ,
    \new_[2644]_ , \new_[2645]_ , \new_[2646]_ , \new_[2647]_ ,
    \new_[2648]_ , \new_[2649]_ , \new_[2650]_ , \new_[2651]_ ,
    \new_[2652]_ , \new_[2653]_ , \new_[2655]_ , \new_[2656]_ ,
    \new_[2657]_ , \new_[2658]_ , \new_[2659]_ , \new_[2660]_ ,
    \new_[2661]_ , \new_[2662]_ , \new_[2663]_ , \new_[2664]_ ,
    \new_[2665]_ , \new_[2666]_ , \new_[2667]_ , \new_[2668]_ ,
    \new_[2669]_ , \new_[2670]_ , \new_[2671]_ , \new_[2672]_ ,
    \new_[2673]_ , \new_[2674]_ , \new_[2675]_ , \new_[2676]_ ,
    \new_[2677]_ , \new_[2678]_ , \new_[2679]_ , \new_[2680]_ ,
    \new_[2681]_ , \new_[2682]_ , \new_[2683]_ , \new_[2684]_ ,
    \new_[2685]_ , \new_[2686]_ , \new_[2687]_ , \new_[2688]_ ,
    \new_[2689]_ , \new_[2690]_ , \new_[2691]_ , \new_[2692]_ ,
    \new_[2693]_ , \new_[2694]_ , \new_[2695]_ , \new_[2696]_ ,
    \new_[2697]_ , \new_[2698]_ , \new_[2699]_ , \new_[2700]_ ,
    \new_[2701]_ , \new_[2702]_ , \new_[2703]_ , \new_[2704]_ ,
    \new_[2705]_ , \new_[2706]_ , \new_[2707]_ , \new_[2708]_ ,
    \new_[2709]_ , \new_[2710]_ , \new_[2711]_ , \new_[2712]_ ,
    \new_[2713]_ , \new_[2714]_ , \new_[2715]_ , \new_[2716]_ ,
    \new_[2717]_ , \new_[2718]_ , \new_[2719]_ , \new_[2720]_ ,
    \new_[2721]_ , \new_[2722]_ , \new_[2723]_ , \new_[2724]_ ,
    \new_[2725]_ , \new_[2726]_ , \new_[2727]_ , \new_[2728]_ ,
    \new_[2729]_ , \new_[2730]_ , \new_[2731]_ , \new_[2732]_ ,
    \new_[2733]_ , \new_[2734]_ , \new_[2735]_ , \new_[2736]_ ,
    \new_[2737]_ , \new_[2738]_ , \new_[2739]_ , \new_[2740]_ ,
    \new_[2741]_ , \new_[2742]_ , \new_[2743]_ , \new_[2744]_ ,
    \new_[2745]_ , \new_[2746]_ , \new_[2747]_ , \new_[2748]_ ,
    \new_[2749]_ , \new_[2750]_ , \new_[2751]_ , \new_[2752]_ ,
    \new_[2753]_ , \new_[2754]_ , \new_[2755]_ , \new_[2756]_ ,
    \new_[2757]_ , \new_[2758]_ , \new_[2759]_ , \new_[2760]_ ,
    \new_[2761]_ , \new_[2762]_ , \new_[2763]_ , \new_[2764]_ ,
    \new_[2765]_ , \new_[2766]_ , \new_[2767]_ , \new_[2768]_ ,
    \new_[2770]_ , \new_[2771]_ , \new_[2772]_ , \new_[2773]_ ,
    \new_[2774]_ , \new_[2775]_ , \new_[2776]_ , \new_[2777]_ ,
    \new_[2778]_ , \new_[2779]_ , \new_[2780]_ , \new_[2781]_ ,
    \new_[2782]_ , \new_[2783]_ , \new_[2784]_ , \new_[2785]_ ,
    \new_[2786]_ , \new_[2787]_ , \new_[2788]_ , \new_[2789]_ ,
    \new_[2790]_ , \new_[2791]_ , \new_[2792]_ , \new_[2793]_ ,
    \new_[2794]_ , \new_[2795]_ , \new_[2796]_ , \new_[2797]_ ,
    \new_[2798]_ , \new_[2799]_ , \new_[2800]_ , \new_[2801]_ ,
    \new_[2802]_ , \new_[2803]_ , \new_[2804]_ , \new_[2805]_ ,
    \new_[2806]_ , \new_[2807]_ , \new_[2808]_ , \new_[2809]_ ,
    \new_[2810]_ , \new_[2811]_ , \new_[2812]_ , \new_[2813]_ ,
    \new_[2814]_ , \new_[2815]_ , \new_[2816]_ , \new_[2817]_ ,
    \new_[2818]_ , \new_[2819]_ , \new_[2820]_ , \new_[2821]_ ,
    \new_[2822]_ , \new_[2823]_ , \new_[2824]_ , \new_[2825]_ ,
    \new_[2826]_ , \new_[2827]_ , \new_[2828]_ , \new_[2829]_ ,
    \new_[2830]_ , \new_[2831]_ , \new_[2832]_ , \new_[2833]_ ,
    \new_[2834]_ , \new_[2835]_ , \new_[2836]_ , \new_[2837]_ ,
    \new_[2838]_ , \new_[2839]_ , \new_[2840]_ , \new_[2841]_ ,
    \new_[2842]_ , \new_[2843]_ , \new_[2844]_ , \new_[2845]_ ,
    \new_[2846]_ , \new_[2847]_ , \new_[2848]_ , \new_[2849]_ ,
    \new_[2850]_ , \new_[2851]_ , \new_[2852]_ , \new_[2853]_ ,
    \new_[2854]_ , \new_[2855]_ , \new_[2856]_ , \new_[2857]_ ,
    \new_[2858]_ , \new_[2859]_ , \new_[2860]_ , \new_[2861]_ ,
    \new_[2862]_ , \new_[2863]_ , \new_[2864]_ , \new_[2865]_ ,
    \new_[2866]_ , \new_[2867]_ , \new_[2868]_ , \new_[2869]_ ,
    \new_[2870]_ , \new_[2871]_ , \new_[2872]_ , \new_[2873]_ ,
    \new_[2874]_ , \new_[2875]_ , \new_[2876]_ , \new_[2877]_ ,
    \new_[2878]_ , \new_[2879]_ , \new_[2880]_ , \new_[2881]_ ,
    \new_[2882]_ , \new_[2883]_ , \new_[2884]_ , \new_[2885]_ ,
    \new_[2886]_ , \new_[2887]_ , \new_[2888]_ , \new_[2889]_ ,
    \new_[2890]_ , \new_[2891]_ , \new_[2892]_ , \new_[2893]_ ,
    \new_[2894]_ , \new_[2895]_ , \new_[2896]_ , \new_[2897]_ ,
    \new_[2898]_ , \new_[2899]_ , \new_[2900]_ , \new_[2901]_ ,
    \new_[2902]_ , \new_[2903]_ , \new_[2904]_ , \new_[2905]_ ,
    \new_[2906]_ , \new_[2907]_ , \new_[2908]_ , \new_[2909]_ ,
    \new_[2910]_ , \new_[2911]_ , \new_[2912]_ , \new_[2913]_ ,
    \new_[2914]_ , \new_[2915]_ , \new_[2916]_ , \new_[2917]_ ,
    \new_[2918]_ , \new_[2919]_ , \new_[2920]_ , \new_[2921]_ ,
    \new_[2923]_ , \new_[2924]_ , \new_[2925]_ , \new_[2926]_ ,
    \new_[2927]_ , \new_[2928]_ , \new_[2929]_ , \new_[2930]_ ,
    \new_[2931]_ , \new_[2932]_ , \new_[2933]_ , \new_[2934]_ ,
    \new_[2935]_ , \new_[2936]_ , \new_[2937]_ , \new_[2938]_ ,
    \new_[2939]_ , \new_[2940]_ , \new_[2941]_ , \new_[2942]_ ,
    \new_[2943]_ , \new_[2944]_ , \new_[2945]_ , \new_[2946]_ ,
    \new_[2947]_ , \new_[2948]_ , \new_[2949]_ , \new_[2950]_ ,
    \new_[2951]_ , \new_[2952]_ , \new_[2953]_ , \new_[2954]_ ,
    \new_[2955]_ , \new_[2956]_ , \new_[2957]_ , \new_[2958]_ ,
    \new_[2959]_ , \new_[2960]_ , \new_[2961]_ , \new_[2962]_ ,
    \new_[2963]_ , \new_[2964]_ , \new_[2965]_ , \new_[2966]_ ,
    \new_[2967]_ , \new_[2968]_ , \new_[2969]_ , \new_[2970]_ ,
    \new_[2971]_ , \new_[2972]_ , \new_[2973]_ , \new_[2974]_ ,
    \new_[2975]_ , \new_[2976]_ , \new_[2977]_ , \new_[2978]_ ,
    \new_[2979]_ , \new_[2980]_ , \new_[2981]_ , \new_[2982]_ ,
    \new_[2983]_ , \new_[2984]_ , \new_[2985]_ , \new_[2986]_ ,
    \new_[2987]_ , \new_[2988]_ , \new_[2989]_ , \new_[2990]_ ,
    \new_[2991]_ , \new_[2992]_ , \new_[2993]_ , \new_[2994]_ ,
    \new_[2995]_ , \new_[2996]_ , \new_[2997]_ , \new_[2998]_ ,
    \new_[2999]_ , \new_[3000]_ , \new_[3001]_ , \new_[3002]_ ,
    \new_[3003]_ , \new_[3004]_ , \new_[3005]_ , \new_[3006]_ ,
    \new_[3007]_ , \new_[3008]_ , \new_[3009]_ , \new_[3010]_ ,
    \new_[3011]_ , \new_[3012]_ , \new_[3013]_ , \new_[3014]_ ,
    \new_[3015]_ , \new_[3016]_ , \new_[3017]_ , \new_[3018]_ ,
    \new_[3019]_ , \new_[3020]_ , \new_[3021]_ , \new_[3022]_ ,
    \new_[3023]_ , \new_[3024]_ , \new_[3025]_ , \new_[3026]_ ,
    \new_[3027]_ , \new_[3028]_ , \new_[3029]_ , \new_[3030]_ ,
    \new_[3031]_ , \new_[3032]_ , \new_[3033]_ , \new_[3034]_ ,
    \new_[3035]_ , \new_[3036]_ , \new_[3037]_ , \new_[3038]_ ,
    \new_[3039]_ , \new_[3040]_ , \new_[3041]_ , \new_[3042]_ ,
    \new_[3043]_ , \new_[3044]_ , \new_[3045]_ , \new_[3046]_ ,
    \new_[3047]_ , \new_[3048]_ , \new_[3049]_ , \new_[3050]_ ,
    \new_[3051]_ , \new_[3052]_ , \new_[3053]_ , \new_[3054]_ ,
    \new_[3055]_ , \new_[3056]_ , \new_[3057]_ , \new_[3058]_ ,
    \new_[3059]_ , \new_[3060]_ , \new_[3061]_ , \new_[3062]_ ,
    \new_[3063]_ , \new_[3064]_ , \new_[3065]_ , \new_[3066]_ ,
    \new_[3067]_ , \new_[3068]_ , \new_[3069]_ , \new_[3070]_ ,
    \new_[3071]_ , \new_[3072]_ , \new_[3073]_ , \new_[3074]_ ,
    \new_[3075]_ , \new_[3076]_ , \new_[3077]_ , \new_[3078]_ ,
    \new_[3079]_ , \new_[3080]_ , \new_[3081]_ , \new_[3082]_ ,
    \new_[3083]_ , \new_[3084]_ , \new_[3085]_ , \new_[3086]_ ,
    \new_[3087]_ , \new_[3088]_ , \new_[3089]_ , \new_[3090]_ ,
    \new_[3091]_ , \new_[3092]_ , \new_[3093]_ , \new_[3094]_ ,
    \new_[3095]_ , \new_[3096]_ , \new_[3097]_ , \new_[3098]_ ,
    \new_[3099]_ , \new_[3100]_ , \new_[3101]_ , \new_[3102]_ ,
    \new_[3103]_ , \new_[3104]_ , \new_[3105]_ , \new_[3106]_ ,
    \new_[3107]_ , \new_[3108]_ , \new_[3109]_ , \new_[3110]_ ,
    \new_[3111]_ , \new_[3112]_ , \new_[3113]_ , \new_[3114]_ ,
    \new_[3115]_ , \new_[3116]_ , \new_[3117]_ , \new_[3118]_ ,
    \new_[3119]_ , \new_[3120]_ , \new_[3121]_ , \new_[3122]_ ,
    \new_[3123]_ , \new_[3124]_ , \new_[3125]_ , \new_[3127]_ ,
    \new_[3128]_ , \new_[3129]_ , \new_[3130]_ , \new_[3131]_ ,
    \new_[3132]_ , \new_[3133]_ , \new_[3134]_ , \new_[3135]_ ,
    \new_[3136]_ , \new_[3137]_ , \new_[3138]_ , \new_[3139]_ ,
    \new_[3140]_ , \new_[3141]_ , \new_[3142]_ , \new_[3143]_ ,
    \new_[3144]_ , \new_[3145]_ , \new_[3146]_ , \new_[3147]_ ,
    \new_[3148]_ , \new_[3149]_ , \new_[3150]_ , \new_[3151]_ ,
    \new_[3152]_ , \new_[3153]_ , \new_[3154]_ , \new_[3155]_ ,
    \new_[3156]_ , \new_[3157]_ , \new_[3158]_ , \new_[3159]_ ,
    \new_[3160]_ , \new_[3161]_ , \new_[3162]_ , \new_[3163]_ ,
    \new_[3164]_ , \new_[3165]_ , \new_[3166]_ , \new_[3167]_ ,
    \new_[3168]_ , \new_[3169]_ , \new_[3170]_ , \new_[3171]_ ,
    \new_[3172]_ , \new_[3173]_ , \new_[3174]_ , \new_[3175]_ ,
    \new_[3176]_ , \new_[3177]_ , \new_[3178]_ , \new_[3179]_ ,
    \new_[3180]_ , \new_[3181]_ , \new_[3182]_ , \new_[3183]_ ,
    \new_[3184]_ , \new_[3185]_ , \new_[3186]_ , \new_[3187]_ ,
    \new_[3188]_ , \new_[3189]_ , \new_[3190]_ , \new_[3191]_ ,
    \new_[3192]_ , \new_[3193]_ , \new_[3194]_ , \new_[3195]_ ,
    \new_[3196]_ , \new_[3197]_ , \new_[3198]_ , \new_[3199]_ ,
    \new_[3200]_ , \new_[3201]_ , \new_[3202]_ , \new_[3203]_ ,
    \new_[3204]_ , \new_[3205]_ , \new_[3206]_ , \new_[3207]_ ,
    \new_[3208]_ , \new_[3209]_ , \new_[3210]_ , \new_[3211]_ ,
    \new_[3212]_ , \new_[3213]_ , \new_[3214]_ , \new_[3215]_ ,
    \new_[3216]_ , \new_[3217]_ , \new_[3218]_ , \new_[3219]_ ,
    \new_[3220]_ , \new_[3221]_ , \new_[3222]_ , \new_[3223]_ ,
    \new_[3224]_ , \new_[3225]_ , \new_[3226]_ , \new_[3227]_ ,
    \new_[3228]_ , \new_[3229]_ , \new_[3230]_ , \new_[3231]_ ,
    \new_[3232]_ , \new_[3233]_ , \new_[3234]_ , \new_[3235]_ ,
    \new_[3236]_ , \new_[3237]_ , \new_[3238]_ , \new_[3239]_ ,
    \new_[3240]_ , \new_[3241]_ , \new_[3242]_ , \new_[3243]_ ,
    \new_[3244]_ , \new_[3245]_ , \new_[3246]_ , \new_[3247]_ ,
    \new_[3248]_ , \new_[3249]_ , \new_[3250]_ , \new_[3251]_ ,
    \new_[3252]_ , \new_[3253]_ , \new_[3254]_ , \new_[3255]_ ,
    \new_[3256]_ , \new_[3257]_ , \new_[3258]_ , \new_[3259]_ ,
    \new_[3260]_ , \new_[3261]_ , \new_[3262]_ , \new_[3263]_ ,
    \new_[3264]_ , \new_[3265]_ , \new_[3266]_ , \new_[3267]_ ,
    \new_[3268]_ , \new_[3269]_ , \new_[3270]_ , \new_[3271]_ ,
    \new_[3272]_ , \new_[3273]_ , \new_[3274]_ , \new_[3275]_ ,
    \new_[3276]_ , \new_[3277]_ , \new_[3278]_ , \new_[3279]_ ,
    \new_[3280]_ , \new_[3281]_ , \new_[3282]_ , \new_[3283]_ ,
    \new_[3284]_ , \new_[3285]_ , \new_[3286]_ , \new_[3287]_ ,
    \new_[3288]_ , \new_[3289]_ , \new_[3290]_ , \new_[3291]_ ,
    \new_[3292]_ , \new_[3293]_ , \new_[3294]_ , \new_[3295]_ ,
    \new_[3296]_ , \new_[3297]_ , \new_[3298]_ , \new_[3299]_ ,
    \new_[3300]_ , \new_[3301]_ , \new_[3303]_ , \new_[3304]_ ,
    \new_[3305]_ , \new_[3306]_ , \new_[3307]_ , \new_[3308]_ ,
    \new_[3309]_ , \new_[3310]_ , \new_[3311]_ , \new_[3312]_ ,
    \new_[3313]_ , \new_[3314]_ , \new_[3315]_ , \new_[3316]_ ,
    \new_[3317]_ , \new_[3318]_ , \new_[3319]_ , \new_[3320]_ ,
    \new_[3321]_ , \new_[3322]_ , \new_[3323]_ , \new_[3324]_ ,
    \new_[3325]_ , \new_[3326]_ , \new_[3327]_ , \new_[3328]_ ,
    \new_[3329]_ , \new_[3330]_ , \new_[3331]_ , \new_[3332]_ ,
    \new_[3333]_ , \new_[3334]_ , \new_[3335]_ , \new_[3336]_ ,
    \new_[3337]_ , \new_[3338]_ , \new_[3339]_ , \new_[3340]_ ,
    \new_[3341]_ , \new_[3342]_ , \new_[3343]_ , \new_[3344]_ ,
    \new_[3345]_ , \new_[3346]_ , \new_[3347]_ , \new_[3348]_ ,
    \new_[3349]_ , \new_[3350]_ , \new_[3351]_ , \new_[3352]_ ,
    \new_[3353]_ , \new_[3354]_ , \new_[3355]_ , \new_[3356]_ ,
    \new_[3357]_ , \new_[3358]_ , \new_[3359]_ , \new_[3360]_ ,
    \new_[3361]_ , \new_[3362]_ , \new_[3363]_ , \new_[3364]_ ,
    \new_[3365]_ , \new_[3366]_ , \new_[3367]_ , \new_[3368]_ ,
    \new_[3369]_ , \new_[3370]_ , \new_[3371]_ , \new_[3372]_ ,
    \new_[3373]_ , \new_[3374]_ , \new_[3375]_ , \new_[3376]_ ,
    \new_[3377]_ , \new_[3378]_ , \new_[3379]_ , \new_[3380]_ ,
    \new_[3381]_ , \new_[3382]_ , \new_[3383]_ , \new_[3384]_ ,
    \new_[3385]_ , \new_[3386]_ , \new_[3387]_ , \new_[3388]_ ,
    \new_[3389]_ , \new_[3390]_ , \new_[3391]_ , \new_[3392]_ ,
    \new_[3393]_ , \new_[3394]_ , \new_[3395]_ , \new_[3396]_ ,
    \new_[3397]_ , \new_[3398]_ , \new_[3399]_ , \new_[3400]_ ,
    \new_[3401]_ , \new_[3402]_ , \new_[3403]_ , \new_[3404]_ ,
    \new_[3405]_ , \new_[3406]_ , \new_[3407]_ , \new_[3408]_ ,
    \new_[3409]_ , \new_[3410]_ , \new_[3411]_ , \new_[3412]_ ,
    \new_[3413]_ , \new_[3414]_ , \new_[3415]_ , \new_[3416]_ ,
    \new_[3417]_ , \new_[3418]_ , \new_[3419]_ , \new_[3420]_ ,
    \new_[3421]_ , \new_[3422]_ , \new_[3423]_ , \new_[3424]_ ,
    \new_[3425]_ , \new_[3426]_ , \new_[3427]_ , \new_[3428]_ ,
    \new_[3429]_ , \new_[3430]_ , \new_[3431]_ , \new_[3432]_ ,
    \new_[3433]_ , \new_[3434]_ , \new_[3435]_ , \new_[3436]_ ,
    \new_[3437]_ , \new_[3438]_ , \new_[3439]_ , \new_[3440]_ ,
    \new_[3441]_ , \new_[3442]_ , \new_[3443]_ , \new_[3444]_ ,
    \new_[3445]_ , \new_[3446]_ , \new_[3447]_ , \new_[3448]_ ,
    \new_[3449]_ , \new_[3450]_ , \new_[3451]_ , \new_[3452]_ ,
    \new_[3453]_ , \new_[3454]_ , \new_[3455]_ , \new_[3456]_ ,
    \new_[3457]_ , \new_[3458]_ , \new_[3459]_ , \new_[3460]_ ,
    \new_[3461]_ , \new_[3462]_ , \new_[3464]_ , \new_[3465]_ ,
    \new_[3466]_ , \new_[3467]_ , \new_[3468]_ , \new_[3469]_ ,
    \new_[3470]_ , \new_[3471]_ , \new_[3472]_ , \new_[3473]_ ,
    \new_[3474]_ , \new_[3475]_ , \new_[3476]_ , \new_[3477]_ ,
    \new_[3478]_ , \new_[3479]_ , \new_[3480]_ , \new_[3481]_ ,
    \new_[3482]_ , \new_[3483]_ , \new_[3484]_ , \new_[3485]_ ,
    \new_[3486]_ , \new_[3487]_ , \new_[3488]_ , \new_[3489]_ ,
    \new_[3490]_ , \new_[3492]_ , \new_[3493]_ , \new_[3494]_ ,
    \new_[3495]_ , \new_[3496]_ , \new_[3497]_ , \new_[3499]_ ,
    \new_[3500]_ , \new_[3501]_ , \new_[3502]_ , \new_[3503]_ ,
    \new_[3504]_ , \new_[3505]_ , \new_[3506]_ , \new_[3507]_ ,
    \new_[3508]_ , \new_[3509]_ , \new_[3510]_ , \new_[3511]_ ,
    \new_[3512]_ , \new_[3513]_ , \new_[3514]_ , \new_[3515]_ ,
    \new_[3516]_ , \new_[3517]_ , \new_[3518]_ , \new_[3519]_ ,
    \new_[3520]_ , \new_[3521]_ , \new_[3522]_ , \new_[3523]_ ,
    \new_[3524]_ , \new_[3525]_ , \new_[3526]_ , \new_[3527]_ ,
    \new_[3528]_ , \new_[3529]_ , \new_[3530]_ , \new_[3531]_ ,
    \new_[3532]_ , \new_[3533]_ , \new_[3534]_ , \new_[3535]_ ,
    \new_[3536]_ , \new_[3537]_ , \new_[3538]_ , \new_[3539]_ ,
    \new_[3540]_ , \new_[3541]_ , \new_[3542]_ , \new_[3543]_ ,
    \new_[3544]_ , \new_[3545]_ , \new_[3546]_ , \new_[3547]_ ,
    \new_[3548]_ , \new_[3549]_ , \new_[3550]_ , n186, n191, n196, n201,
    n206, n211, n216, n221, n226, n231, n236, n241, n246, n251, n256, n261,
    n266, n271, n276, n281, n286, n291, n296, n301, n306, n311, n316, n321,
    n326, n331, n336, n341, n346, n351, n356, n361, n366, n371, n376, n381,
    n386, n391, n396, n401, n406, n411, n416, n421, n426, n431, n436, n441,
    n446, n451, n456, n461, n466, n471, n476, n481, n486, n491, n496, n501,
    n506, n511, n516, n521, n526, n531, n536, n541, n546, n551, n556, n561,
    n566, n571, n576, n581, n586, n591, n596, n601, n606, n611, n616, n621,
    n626, n631, n636, n641, n646, n651, n656, n661, n666, n671, n676, n681,
    n686, n691, n696, n701, n706, n711, n716, n721, n726, n731, n736, n741,
    n746, n751, n756, n761, n766, n771, n776, n781, n786, n791, n796, n801,
    n806, n811, n816, n821, n826, n831, n836, n841, n846, n851, n856, n861,
    n866, n871, n876, n881, n886, n891, n896, n901, n906, n911, n916, n921,
    n926, n931, n936, n941, n946, n951, n956, n961, n966, n971, n976, n981,
    n986, n991, n996, n1001, n1006, n1011, n1016, n1021, n1026, n1031,
    n1036, n1041, n1046, n1051, n1056, n1061, n1066, n1071, n1076, n1081,
    n1086, n1091, n1096, n1101, n1106, n1111, n1116, n1121, n1126, n1131,
    n1136, n1141, n1146, n1151, n1156, n1161, n1166, n1171, n1176, n1181,
    n1186, n1191, n1196, n1201, n1206, n1211, n1216, n1221, n1226, n1231,
    n1236, n1241, n1246, n1251, n1256, n1261, n1266, n1271, n1276, n1281,
    n1286, n1291, n1296, n1301, n1306, n1311, n1316, n1321, n1326;
  assign \new_[321]_  = 1'b0;
  assign wb_err_o = \new_[321]_ ;
  assign \new_[324]_  = \\shift_data_reg[39] ;
  assign \new_[325]_  = \\shift_data_reg[56] ;
  assign \new_[326]_  = \\shift_data_reg[63] ;
  assign \new_[327]_  = \\shift_data_reg[32] ;
  assign \new_[328]_  = \\shift_data_reg[65] ;
  assign \new_[329]_  = \\shift_data_reg[66] ;
  assign \new_[330]_  = \\shift_data_reg[68] ;
  assign \new_[331]_  = \\shift_data_reg[71] ;
  assign \new_[332]_  = \\shift_data_reg[74] ;
  assign \new_[333]_  = \\shift_data_reg[75] ;
  assign \new_[334]_  = \\shift_data_reg[76] ;
  assign \new_[335]_  = \\shift_data_reg[85] ;
  assign \new_[336]_  = \\shift_data_reg[86] ;
  assign \new_[337]_  = \\shift_data_reg[87] ;
  assign \new_[338]_  = \\shift_data_reg[91] ;
  assign \new_[339]_  = \\shift_data_reg[93] ;
  assign \new_[340]_  = \\shift_data_reg[94] ;
  assign \new_[341]_  = \\shift_data_reg[95] ;
  assign \new_[342]_  = \\shift_data_reg[0] ;
  assign \new_[343]_  = \\shift_data_reg[2] ;
  assign \new_[344]_  = \\shift_data_reg[4] ;
  assign \new_[345]_  = \\shift_data_reg[7] ;
  assign \new_[346]_  = \\shift_data_reg[8] ;
  assign \new_[347]_  = \\shift_data_reg[14] ;
  assign \new_[348]_  = \\shift_data_reg[15] ;
  assign \new_[349]_  = \\shift_data_reg[16] ;
  assign \new_[350]_  = \\shift_data_reg[17] ;
  assign \new_[351]_  = \\shift_data_reg[18] ;
  assign \new_[352]_  = \\shift_data_reg[1] ;
  assign \new_[353]_  = \\shift_data_reg[20] ;
  assign \new_[354]_  = \\shift_data_reg[23] ;
  assign \new_[355]_  = \\shift_data_reg[92] ;
  assign \new_[356]_  = \\shift_data_reg[89] ;
  assign \new_[357]_  = \\shift_data_reg[64] ;
  assign \new_[358]_  = \\shift_data_reg[67] ;
  assign \new_[359]_  = \\shift_data_reg[69] ;
  assign \new_[360]_  = \\shift_data_reg[70] ;
  assign \new_[361]_  = \\shift_data_reg[72] ;
  assign \new_[362]_  = \\shift_data_reg[73] ;
  assign \new_[363]_  = \\shift_data_reg[77] ;
  assign \new_[364]_  = \\shift_data_reg[80] ;
  assign \new_[365]_  = \\shift_data_reg[83] ;
  assign \new_[366]_  = \\shift_data_reg[84] ;
  assign \new_[367]_  = \\shift_data_reg[81] ;
  assign \new_[368]_  = \\shift_data_reg[88] ;
  assign \new_[369]_  = \\shift_data_reg[82] ;
  assign \new_[370]_  = \\shift_data_reg[90] ;
  assign \new_[371]_  = \\shift_data_reg[79] ;
  assign \new_[372]_  = \\shift_data_reg[78] ;
  assign \new_[373]_  = \\shift_data_reg[26] ;
  assign \new_[374]_  = \\shift_data_reg[27] ;
  assign \new_[375]_  = \\shift_data_reg[24] ;
  assign \new_[376]_  = \\shift_data_reg[29] ;
  assign \new_[377]_  = \\shift_data_reg[28] ;
  assign \new_[378]_  = \\shift_data_reg[30] ;
  assign \new_[379]_  = \\shift_data_reg[31] ;
  assign \new_[380]_  = \\shift_data_reg[10] ;
  assign \new_[381]_  = \\shift_data_reg[3] ;
  assign \new_[382]_  = \\shift_data_reg[5] ;
  assign \new_[383]_  = \\shift_data_reg[25] ;
  assign \new_[384]_  = \\shift_data_reg[6] ;
  assign \new_[385]_  = \\shift_data_reg[12] ;
  assign \new_[386]_  = \\shift_data_reg[13] ;
  assign \new_[387]_  = \\shift_data_reg[11] ;
  assign \new_[388]_  = \\shift_data_reg[9] ;
  assign \new_[389]_  = \\shift_data_reg[19] ;
  assign \new_[390]_  = \\shift_data_reg[21] ;
  assign \new_[391]_  = \\shift_data_reg[22] ;
  assign \new_[392]_  = \\shift_data_reg[53] ;
  assign \new_[393]_  = \\shift_data_reg[54] ;
  assign \new_[394]_  = \\shift_data_reg[51] ;
  assign n216 = ~\new_[521]_  | ~\new_[1992]_ ;
  assign n221 = ~\new_[522]_  | ~\new_[1976]_ ;
  assign n226 = ~\new_[523]_  | ~\new_[1979]_ ;
  assign n231 = ~\new_[525]_  | ~\new_[1980]_ ;
  assign n236 = ~\new_[526]_  | ~\new_[1981]_ ;
  assign n241 = ~\new_[529]_  | ~\new_[1990]_ ;
  assign n196 = ~\new_[2246]_  | ~\new_[548]_ ;
  assign n246 = ~\new_[530]_  | ~\new_[2001]_ ;
  assign n251 = ~\new_[531]_  | ~\new_[1991]_ ;
  assign n256 = ~\new_[533]_  | ~\new_[1995]_ ;
  assign n261 = ~\new_[534]_  | ~\new_[1997]_ ;
  assign n201 = ~\new_[545]_  | ~\new_[2238]_ ;
  assign n266 = ~\new_[535]_  | ~\new_[2000]_ ;
  assign n186 = ~\new_[546]_  | ~\new_[2239]_ ;
  assign n271 = ~\new_[536]_  | ~\new_[1998]_ ;
  assign n191 = ~\new_[547]_  | ~\new_[2243]_ ;
  assign n281 = ~\new_[515]_  | ~\new_[2332]_ ;
  assign n286 = ~\new_[517]_  | ~\new_[2339]_ ;
  assign n276 = ~\new_[518]_  | ~\new_[2338]_ ;
  assign n291 = ~\new_[2345]_  | ~\new_[527]_ ;
  assign n296 = ~\new_[532]_  | ~\new_[2348]_ ;
  assign n301 = ~\new_[2351]_  | ~\new_[537]_ ;
  assign n306 = ~\new_[538]_  | ~\new_[2341]_ ;
  assign n311 = ~\new_[539]_  | ~\new_[2337]_ ;
  assign n316 = ~\new_[2352]_  | ~\new_[540]_ ;
  assign n321 = ~\new_[2335]_  | ~\new_[541]_ ;
  assign n326 = ~\new_[542]_  | ~\new_[2236]_ ;
  assign n331 = ~\new_[2347]_  | ~\new_[543]_ ;
  assign n336 = ~\new_[544]_  | ~\new_[2344]_ ;
  assign \new_[424]_  = \\shift_data_reg[33] ;
  assign \new_[425]_  = \\shift_data_reg[34] ;
  assign \new_[426]_  = \\shift_data_reg[35] ;
  assign \new_[427]_  = \\shift_data_reg[36] ;
  assign \new_[428]_  = \\shift_data_reg[43] ;
  assign \new_[429]_  = \\shift_data_reg[45] ;
  assign \new_[430]_  = \\shift_data_reg[46] ;
  assign \new_[431]_  = \\shift_data_reg[47] ;
  assign \new_[432]_  = \\shift_data_reg[57] ;
  assign \new_[433]_  = \\shift_data_reg[58] ;
  assign \new_[434]_  = \\shift_data_reg[59] ;
  assign \new_[435]_  = \\shift_data_reg[61] ;
  assign \new_[436]_  = \\shift_data_reg[62] ;
  assign \new_[437]_  = \\shift_data_reg[104] ;
  assign \new_[438]_  = \\shift_data_reg[111] ;
  assign \new_[439]_  = \\shift_data_reg[112] ;
  assign \new_[440]_  = \\shift_data_reg[119] ;
  assign \new_[441]_  = \\shift_data_reg[121] ;
  assign \new_[442]_  = \\shift_data_reg[97] ;
  assign \new_[443]_  = \\shift_data_reg[123] ;
  assign \new_[444]_  = \\shift_data_reg[125] ;
  assign \new_[445]_  = \\shift_data_reg[126] ;
  assign \new_[446]_  = \\shift_data_reg[122] ;
  assign \new_[447]_  = \\shift_data_reg[127] ;
  assign n206 = ~\new_[519]_  | ~\new_[1972]_ ;
  assign n211 = ~\new_[520]_  | ~\new_[1982]_ ;
  assign n361 = ~\new_[584]_  | ~\new_[1974]_ ;
  assign n366 = ~\new_[1975]_  | ~\new_[586]_ ;
  assign n371 = ~\new_[587]_  | ~\new_[1977]_ ;
  assign n376 = ~\new_[588]_  | ~\new_[1978]_ ;
  assign n381 = ~\new_[589]_  | ~\new_[1999]_ ;
  assign n426 = ~\new_[590]_  | ~\new_[1983]_ ;
  assign n421 = ~\new_[591]_  | ~\new_[1984]_ ;
  assign n401 = ~\new_[593]_  | ~\new_[1986]_ ;
  assign n411 = ~\new_[1970]_  | ~\new_[594]_ ;
  assign n386 = ~\new_[592]_  | ~\new_[1985]_ ;
  assign n391 = ~\new_[595]_  | ~\new_[1988]_ ;
  assign n396 = ~\new_[596]_  | ~\new_[1989]_ ;
  assign n406 = ~\new_[597]_  | ~\new_[1987]_ ;
  assign n416 = ~\new_[598]_  | ~\new_[1994]_ ;
  assign \new_[464]_  = \\shift_data_reg[124] ;
  assign \new_[465]_  = \\shift_data_reg[98] ;
  assign n346 = ~\new_[1993]_  | ~\new_[634]_ ;
  assign n341 = ~\new_[635]_  | ~\new_[1996]_ ;
  assign \new_[468]_  = \\shift_data_reg[114] ;
  assign n481 = ~\new_[2461]_  | ~\new_[633]_ ;
  assign n436 = ~\new_[2340]_  | ~\new_[637]_ ;
  assign n451 = ~\new_[2463]_  | ~\new_[638]_ ;
  assign n431 = ~\new_[2462]_  | ~\new_[636]_ ;
  assign n446 = ~\new_[2464]_  | ~\new_[639]_ ;
  assign \new_[474]_  = \\shift_data_reg[60] ;
  assign n456 = ~\new_[2333]_  | ~\new_[578]_ ;
  assign n461 = ~\new_[2334]_  | ~\new_[579]_ ;
  assign n471 = ~\new_[2336]_  | ~\new_[580]_ ;
  assign n476 = ~\new_[2343]_  | ~\new_[581]_ ;
  assign n486 = ~\new_[2346]_  | ~\new_[585]_ ;
  assign n466 = ~\new_[2233]_  | ~\new_[3278]_ ;
  assign n501 = ~\new_[2349]_  | ~\new_[599]_ ;
  assign \new_[482]_  = \\shift_data_reg[48] ;
  assign n491 = ~\new_[2235]_  | ~\new_[3285]_ ;
  assign n506 = ~\new_[2350]_  | ~\new_[600]_ ;
  assign n496 = ~\new_[2342]_  | ~\new_[601]_ ;
  assign \new_[486]_  = \\shift_data_reg[41] ;
  assign n511 = ~\new_[2353]_  | ~\new_[602]_ ;
  assign \new_[488]_  = \\shift_data_reg[40] ;
  assign n516 = ~\new_[2354]_  | ~\new_[603]_ ;
  assign n521 = ~\new_[2234]_  | ~\new_[604]_ ;
  assign n441 = ~\new_[2355]_  | ~\new_[605]_ ;
  assign \new_[492]_  = \\shift_data_reg[120] ;
  assign \new_[493]_  = \\shift_data_reg[105] ;
  assign \new_[494]_  = \\shift_data_reg[113] ;
  assign \new_[495]_  = \\shift_data_reg[108] ;
  assign \new_[496]_  = \\shift_data_reg[37] ;
  assign \new_[497]_  = \\shift_data_reg[38] ;
  assign \new_[498]_  = \\shift_data_reg[116] ;
  assign \new_[499]_  = \\shift_data_reg[42] ;
  assign \new_[500]_  = \\shift_data_reg[49] ;
  assign \new_[501]_  = \\shift_data_reg[50] ;
  assign \new_[502]_  = \\shift_data_reg[44] ;
  assign \new_[503]_  = \\shift_data_reg[52] ;
  assign \new_[504]_  = \\shift_data_reg[55] ;
  assign \new_[505]_  = \\shift_data_reg[103] ;
  assign \new_[506]_  = \\shift_data_reg[100] ;
  assign \new_[507]_  = \\shift_data_reg[106] ;
  assign \new_[508]_  = \\shift_data_reg[96] ;
  assign \new_[509]_  = \\shift_data_reg[99] ;
  assign n536 = ~\new_[619]_  | ~\new_[2416]_ ;
  assign n531 = ~\new_[621]_  | ~\new_[2458]_ ;
  assign n526 = ~\new_[620]_  | ~\new_[2418]_ ;
  assign n351 = ~\new_[582]_  | ~\new_[1971]_ ;
  assign n356 = ~\new_[583]_  | ~\new_[1973]_ ;
  assign \new_[515]_  = ~\new_[677]_  | ~\new_[2624]_ ;
  assign n636 = ~\new_[641]_  | ~\new_[2072]_ ;
  assign \new_[517]_  = ~\new_[678]_  | ~\new_[2624]_ ;
  assign \new_[518]_  = ~\new_[676]_  | ~\new_[2624]_ ;
  assign \new_[519]_  = ~\new_[649]_  | ~\new_[2561]_ ;
  assign \new_[520]_  = ~\new_[650]_  | ~\new_[2588]_ ;
  assign \new_[521]_  = ~\new_[651]_  | ~\new_[2559]_ ;
  assign \new_[522]_  = ~\new_[652]_  | ~\new_[2588]_ ;
  assign \new_[523]_  = ~\new_[653]_  | ~\new_[2559]_ ;
  assign \new_[524]_  = \\shift_data_reg[118] ;
  assign \new_[525]_  = ~\new_[654]_  | ~\new_[2588]_ ;
  assign \new_[526]_  = ~\new_[655]_  | ~\new_[2561]_ ;
  assign \new_[527]_  = ~\new_[3312]_  | (~\new_[2229]_  & ~\new_[730]_ );
  assign \new_[528]_  = \\shift_data_reg[115] ;
  assign \new_[529]_  = ~\new_[656]_  | ~\new_[2561]_ ;
  assign \new_[530]_  = ~\new_[657]_  | ~\new_[2564]_ ;
  assign \new_[531]_  = ~\new_[658]_  | ~\new_[2564]_ ;
  assign \new_[532]_  = ~\new_[679]_  | ~\new_[2624]_ ;
  assign \new_[533]_  = ~\new_[659]_  | ~\new_[2561]_ ;
  assign \new_[534]_  = ~\new_[660]_  | ~\new_[2588]_ ;
  assign \new_[535]_  = ~\new_[661]_  | ~\new_[2561]_ ;
  assign \new_[536]_  = ~\new_[662]_  | ~\new_[2588]_ ;
  assign \new_[537]_  = ~\new_[3312]_  | (~\new_[2230]_  & ~\new_[731]_ );
  assign \new_[538]_  = ~\new_[680]_  | ~\new_[2624]_ ;
  assign \new_[539]_  = ~\new_[681]_  | ~\new_[2624]_ ;
  assign \new_[540]_  = ~\new_[2562]_  | (~\new_[2231]_  & ~\new_[732]_ );
  assign \new_[541]_  = ~\new_[3312]_  | (~\new_[2228]_  & ~\new_[733]_ );
  assign \new_[542]_  = ~\new_[682]_  | ~\new_[2624]_ ;
  assign \new_[543]_  = ~\new_[3312]_  | (~\new_[2232]_  & ~\new_[734]_ );
  assign \new_[544]_  = ~\new_[683]_  | ~\new_[2624]_ ;
  assign \new_[545]_  = ~\new_[2397]_  & (~\new_[727]_  | ~\new_[2181]_ );
  assign \new_[546]_  = ~\new_[2404]_  & (~\new_[728]_  | ~\new_[2181]_ );
  assign \new_[547]_  = ~\new_[2420]_  & (~\new_[729]_  | ~\new_[2181]_ );
  assign \new_[548]_  = ~\new_[2428]_  & (~\new_[3359]_  | ~\new_[2181]_ );
  assign n651 = ~\new_[684]_  | ~\new_[2046]_ ;
  assign n656 = ~\new_[685]_  | ~\new_[2075]_ ;
  assign n606 = ~\new_[686]_  | ~\new_[2052]_ ;
  assign n611 = ~\new_[687]_  | ~\new_[2057]_ ;
  assign n616 = ~\new_[688]_  | ~\new_[2058]_ ;
  assign n621 = ~\new_[689]_  | ~\new_[2065]_ ;
  assign n626 = ~\new_[690]_  | ~\new_[2070]_ ;
  assign n631 = ~\new_[640]_  | ~\new_[2069]_ ;
  assign \new_[557]_  = \\shift_data_reg[101] ;
  assign \new_[558]_  = \\shift_data_reg[102] ;
  assign \new_[559]_  = \\shift_data_reg[107] ;
  assign \new_[560]_  = \\shift_data_reg[109] ;
  assign \new_[561]_  = \\shift_data_reg[110] ;
  assign \new_[562]_  = \\shift_data_reg[117] ;
  assign n641 = ~\new_[642]_  | ~\new_[2074]_ ;
  assign n646 = ~\new_[643]_  | ~\new_[2062]_ ;
  assign n541 = ~\new_[663]_  | ~\new_[2398]_ ;
  assign n546 = ~\new_[664]_  | ~\new_[2399]_ ;
  assign n551 = ~\new_[665]_  | ~\new_[2400]_ ;
  assign n556 = ~\new_[666]_  | ~\new_[2401]_ ;
  assign n561 = ~\new_[669]_  | ~\new_[2408]_ ;
  assign n566 = ~\new_[667]_  | ~\new_[2410]_ ;
  assign n571 = ~\new_[668]_  | ~\new_[2411]_ ;
  assign n576 = ~\new_[670]_  | ~\new_[2412]_ ;
  assign n581 = ~\new_[671]_  | ~\new_[2421]_ ;
  assign n586 = ~\new_[672]_  | ~\new_[2422]_ ;
  assign n591 = ~\new_[673]_  | ~\new_[2424]_ ;
  assign n596 = ~\new_[674]_  | ~\new_[2426]_ ;
  assign n601 = ~\new_[675]_  | ~\new_[2427]_ ;
  assign \new_[578]_  = ~\new_[2560]_  | (~\new_[755]_  & ~\new_[2226]_ );
  assign \new_[579]_  = ~\new_[3312]_  | (~\new_[756]_  & ~\new_[2227]_ );
  assign \new_[580]_  = ~\new_[2560]_  | (~\new_[757]_  & ~\new_[2323]_ );
  assign \new_[581]_  = ~\new_[2617]_  | (~\new_[2326]_  & ~\new_[758]_ );
  assign \new_[582]_  = ~\new_[700]_  | ~\new_[2559]_ ;
  assign \new_[583]_  = ~\new_[701]_  | ~\new_[2588]_ ;
  assign \new_[584]_  = ~\new_[702]_  | ~\new_[2559]_ ;
  assign \new_[585]_  = ~\new_[2560]_  | (~\new_[760]_  & ~\new_[2324]_ );
  assign \new_[586]_  = ~\new_[703]_  | ~\new_[2559]_ ;
  assign \new_[587]_  = ~\new_[704]_  | ~\new_[2559]_ ;
  assign \new_[588]_  = ~\new_[705]_  | ~\new_[2559]_ ;
  assign \new_[589]_  = ~\new_[706]_  | ~\new_[2559]_ ;
  assign \new_[590]_  = ~\new_[707]_  | ~\new_[2564]_ ;
  assign \new_[591]_  = ~\new_[708]_  | ~\new_[2564]_ ;
  assign \new_[592]_  = ~\new_[709]_  | ~\new_[2564]_ ;
  assign \new_[593]_  = ~\new_[710]_  | ~\new_[2561]_ ;
  assign \new_[594]_  = ~\new_[711]_  | ~\new_[2561]_ ;
  assign \new_[595]_  = ~\new_[712]_  | ~\new_[2588]_ ;
  assign \new_[596]_  = ~\new_[713]_  | ~\new_[2588]_ ;
  assign \new_[597]_  = ~\new_[714]_  | ~\new_[2564]_ ;
  assign \new_[598]_  = ~\new_[715]_  | ~\new_[2561]_ ;
  assign \new_[599]_  = ~\new_[2560]_  | (~\new_[763]_  & ~\new_[2327]_ );
  assign \new_[600]_  = ~\new_[2617]_  | (~\new_[764]_  & ~\new_[2325]_ );
  assign \new_[601]_  = ~\new_[2560]_  | (~\new_[2328]_  & ~\new_[765]_ );
  assign \new_[602]_  = ~\new_[2617]_  | (~\new_[2322]_  & ~\new_[766]_ );
  assign \new_[603]_  = ~\new_[2617]_  | (~\new_[767]_  & ~\new_[2329]_ );
  assign \new_[604]_  = ~\new_[3312]_  | (~\new_[768]_  & ~\new_[2330]_ );
  assign \new_[605]_  = ~\new_[2560]_  | (~\new_[769]_  & ~\new_[2331]_ );
  assign n701 = ~\new_[695]_  | ~\new_[2053]_ ;
  assign n706 = ~\new_[696]_  | ~\new_[2059]_ ;
  assign n711 = ~\new_[697]_  | ~\new_[2056]_ ;
  assign n726 = ~\new_[698]_  | ~\new_[2068]_ ;
  assign n696 = ~\new_[699]_  | ~\new_[2066]_ ;
  assign n766 = ~\new_[735]_  | ~\new_[2049]_ ;
  assign n761 = ~\new_[3226]_  | ~\new_[2051]_ ;
  assign n771 = ~\new_[736]_  | ~\new_[2054]_ ;
  assign n671 = ~\new_[737]_  | ~\new_[2060]_ ;
  assign n776 = ~\new_[738]_  | ~\new_[2067]_ ;
  assign n666 = ~\new_[691]_  | ~\new_[2071]_ ;
  assign n781 = ~\new_[692]_  | ~\new_[2048]_ ;
  assign n661 = ~\new_[3210]_  | ~\new_[2073]_ ;
  assign \new_[619]_  = (~\new_[739]_  | ~\new_[2183]_ ) & (~\new_[3311]_  | ~\new_[394]_ );
  assign \new_[620]_  = (~\new_[740]_  | ~\new_[2097]_ ) & (~\new_[3306]_  | ~\new_[392]_ );
  assign \new_[621]_  = (~\new_[741]_  | ~\new_[2098]_ ) & (~\new_[2626]_  | ~\new_[393]_ );
  assign n716 = ~\new_[716]_  | ~\new_[2402]_ ;
  assign n721 = ~\new_[717]_  | ~\new_[2403]_ ;
  assign n691 = ~\new_[718]_  | ~\new_[2405]_ ;
  assign n686 = ~\new_[719]_  | ~\new_[2406]_ ;
  assign n731 = ~\new_[721]_  | ~\new_[2407]_ ;
  assign n746 = ~\new_[720]_  | ~\new_[2409]_ ;
  assign n681 = ~\new_[722]_  | ~\new_[2413]_ ;
  assign n736 = ~\new_[723]_  | ~\new_[2414]_ ;
  assign n741 = ~\new_[724]_  | ~\new_[2415]_ ;
  assign n751 = ~\new_[725]_  | ~\new_[2417]_ ;
  assign n676 = ~\new_[726]_  | ~\new_[2425]_ ;
  assign \new_[633]_  = ~\new_[2617]_  | (~\new_[2318]_  & ~\new_[750]_ );
  assign \new_[634]_  = ~\new_[693]_  | ~\new_[2564]_ ;
  assign \new_[635]_  = ~\new_[694]_  | ~\new_[2564]_ ;
  assign \new_[636]_  = ~\new_[2617]_  | (~\new_[2319]_  & ~\new_[751]_ );
  assign \new_[637]_  = ~\new_[2617]_  | (~\new_[752]_  & ~\new_[2320]_ );
  assign \new_[638]_  = ~\new_[2617]_  | (~\new_[2321]_  & ~\new_[753]_ );
  assign \new_[639]_  = ~\new_[2560]_  | (~\new_[2225]_  & ~\new_[754]_ );
  assign \new_[640]_  = ~\new_[3218]_  | (~\new_[802]_  & ~\new_[2529]_ );
  assign \new_[641]_  = ~\new_[3218]_  | (~\new_[804]_  & ~\new_[2549]_ );
  assign \new_[642]_  = ~\new_[2098]_  | (~\new_[805]_  & ~\new_[2532]_ );
  assign \new_[643]_  = ~\new_[3310]_  | (~\new_[806]_  & ~\new_[2550]_ );
  assign n801 = ~\new_[3238]_  | ~\new_[2050]_ ;
  assign n806 = ~\new_[759]_  | ~\new_[2055]_ ;
  assign n791 = ~\new_[3264]_  | ~\new_[2061]_ ;
  assign n786 = ~\new_[762]_  | ~\new_[2064]_ ;
  assign n821 = ~\new_[761]_  | ~\new_[2063]_ ;
  assign \new_[649]_  = ~\new_[2430]_  | (~\new_[783]_  & ~\new_[2360]_ );
  assign \new_[650]_  = ~\new_[2431]_  | (~\new_[784]_  & ~\new_[2360]_ );
  assign \new_[651]_  = ~\new_[2433]_  | (~\new_[785]_  & ~\new_[2360]_ );
  assign \new_[652]_  = ~\new_[2436]_  | (~\new_[786]_  & ~\new_[2360]_ );
  assign \new_[653]_  = ~\new_[2439]_  | (~\new_[787]_  & ~\new_[2360]_ );
  assign \new_[654]_  = ~\new_[2440]_  | (~\new_[788]_  & ~\new_[2360]_ );
  assign \new_[655]_  = ~\new_[2443]_  | (~\new_[789]_  & ~\new_[2360]_ );
  assign \new_[656]_  = ~\new_[2460]_  | (~\new_[790]_  & ~\new_[2360]_ );
  assign \new_[657]_  = ~\new_[2456]_  | (~\new_[791]_  & ~\new_[2360]_ );
  assign \new_[658]_  = ~\new_[2450]_  | (~\new_[792]_  & ~\new_[2360]_ );
  assign \new_[659]_  = ~\new_[2452]_  | (~\new_[793]_  & ~\new_[2360]_ );
  assign \new_[660]_  = ~\new_[2454]_  | (~\new_[794]_  & ~\new_[2360]_ );
  assign \new_[661]_  = ~\new_[2459]_  | (~\new_[795]_  & ~\new_[2360]_ );
  assign \new_[662]_  = ~\new_[2455]_  | (~\new_[796]_  & ~\new_[2360]_ );
  assign \new_[663]_  = (~\new_[770]_  | ~\new_[2182]_ ) & (~\new_[2625]_  | ~\new_[424]_ );
  assign \new_[664]_  = (~\new_[771]_  | ~\new_[2183]_ ) & (~\new_[2626]_  | ~\new_[425]_ );
  assign \new_[665]_  = (~\new_[772]_  | ~\new_[2182]_ ) & (~\new_[2558]_  | ~\new_[426]_ );
  assign \new_[666]_  = (~\new_[773]_  | ~\new_[3310]_ ) & (~\new_[2632]_  | ~\new_[427]_ );
  assign \new_[667]_  = (~\new_[775]_  | ~\new_[2183]_ ) & (~\new_[3308]_  | ~\new_[429]_ );
  assign \new_[668]_  = (~\new_[776]_  | ~\new_[2097]_ ) & (~\new_[2626]_  | ~\new_[430]_ );
  assign \new_[669]_  = (~\new_[774]_  | ~\new_[2180]_ ) & (~\new_[2558]_  | ~\new_[428]_ );
  assign \new_[670]_  = (~\new_[777]_  | ~\new_[2180]_ ) & (~\new_[2626]_  | ~\new_[431]_ );
  assign \new_[671]_  = (~\new_[778]_  | ~\new_[2098]_ ) & (~\new_[2632]_  | ~\new_[432]_ );
  assign \new_[672]_  = (~\new_[779]_  | ~\new_[2183]_ ) & (~\new_[2632]_  | ~\new_[433]_ );
  assign \new_[673]_  = (~\new_[780]_  | ~\new_[2098]_ ) & (~\new_[2626]_  | ~\new_[434]_ );
  assign \new_[674]_  = (~\new_[781]_  | ~\new_[2180]_ ) & (~\new_[2625]_  | ~\new_[435]_ );
  assign \new_[675]_  = (~\new_[782]_  | ~\new_[2097]_ ) & (~\new_[3311]_  | ~\new_[436]_ );
  assign \new_[676]_  = ~\new_[743]_  | (~\new_[2240]_  & ~\new_[3146]_ );
  assign \new_[677]_  = ~\new_[742]_  | (~\new_[2240]_  & ~\new_[3176]_ );
  assign \new_[678]_  = ~\new_[744]_  | (~\new_[2240]_  & ~\new_[3199]_ );
  assign \new_[679]_  = ~\new_[745]_  | (~\new_[2240]_  & ~\new_[3113]_ );
  assign \new_[680]_  = ~\new_[746]_  | (~\new_[2240]_  & ~\new_[3138]_ );
  assign \new_[681]_  = ~\new_[747]_  | (~\new_[2240]_  & ~\new_[3084]_ );
  assign \new_[682]_  = ~\new_[748]_  | (~\new_[2240]_  & ~\new_[3139]_ );
  assign \new_[683]_  = ~\new_[749]_  | (~\new_[2240]_  & ~\new_[3195]_ );
  assign \new_[684]_  = ~\new_[3496]_  | (~\new_[803]_  & ~\new_[2531]_ );
  assign \new_[685]_  = ~\new_[2098]_  | (~\new_[807]_  & ~\new_[2540]_ );
  assign \new_[686]_  = ~\new_[3218]_  | (~\new_[797]_  & ~\new_[2534]_ );
  assign \new_[687]_  = ~\new_[3218]_  | (~\new_[798]_  & ~\new_[2539]_ );
  assign \new_[688]_  = ~\new_[2181]_  | (~\new_[799]_  & ~\new_[2541]_ );
  assign \new_[689]_  = ~\new_[2180]_  | (~\new_[800]_  & ~\new_[2584]_ );
  assign \new_[690]_  = ~\new_[2180]_  | (~\new_[801]_  & ~\new_[2547]_ );
  assign \new_[691]_  = ~\new_[3218]_  | (~\new_[853]_  & ~\new_[2548]_ );
  assign \new_[692]_  = ~\new_[3218]_  | (~\new_[854]_  & ~\new_[2533]_ );
  assign \new_[693]_  = ~\new_[2423]_  | (~\new_[808]_  & ~\new_[2360]_ );
  assign \new_[694]_  = ~\new_[2453]_  | (~\new_[809]_  & ~\new_[2360]_ );
  assign \new_[695]_  = ~\new_[3496]_  | (~\new_[810]_  & ~\new_[2535]_ );
  assign \new_[696]_  = ~\new_[2181]_  | (~\new_[812]_  & ~\new_[2542]_ );
  assign \new_[697]_  = ~\new_[2180]_  | (~\new_[811]_  & ~\new_[2538]_ );
  assign \new_[698]_  = ~\new_[3310]_  | (~\new_[813]_  & ~\new_[2546]_ );
  assign \new_[699]_  = ~\new_[3310]_  | (~\new_[3344]_  & ~\new_[2551]_ );
  assign \new_[700]_  = ~\new_[2429]_  | (~\new_[828]_  & ~\new_[2360]_ );
  assign \new_[701]_  = ~\new_[2432]_  | (~\new_[829]_  & ~\new_[2360]_ );
  assign \new_[702]_  = ~\new_[2434]_  | (~\new_[830]_  & ~\new_[2360]_ );
  assign \new_[703]_  = ~\new_[2435]_  | (~\new_[831]_  & ~\new_[2360]_ );
  assign \new_[704]_  = ~\new_[2437]_  | (~\new_[832]_  & ~\new_[2360]_ );
  assign \new_[705]_  = ~\new_[2438]_  | (~\new_[833]_  & ~\new_[2360]_ );
  assign \new_[706]_  = ~\new_[2444]_  | (~\new_[834]_  & ~\new_[2360]_ );
  assign \new_[707]_  = ~\new_[2445]_  | (~\new_[835]_  & ~\new_[2360]_ );
  assign \new_[708]_  = ~\new_[2441]_  | (~\new_[836]_  & ~\new_[2360]_ );
  assign \new_[709]_  = ~\new_[2446]_  | (~\new_[837]_  & ~\new_[2360]_ );
  assign \new_[710]_  = ~\new_[2457]_  | (~\new_[838]_  & ~\new_[2360]_ );
  assign \new_[711]_  = ~\new_[2447]_  | (~\new_[839]_  & ~\new_[2360]_ );
  assign \new_[712]_  = ~\new_[2448]_  | (~\new_[840]_  & ~\new_[2360]_ );
  assign \new_[713]_  = ~\new_[2449]_  | (~\new_[841]_  & ~\new_[2360]_ );
  assign \new_[714]_  = ~\new_[2442]_  | (~\new_[842]_  & ~\new_[2360]_ );
  assign \new_[715]_  = ~\new_[2451]_  | (~\new_[843]_  & ~\new_[2360]_ );
  assign \new_[716]_  = (~\new_[814]_  | ~\new_[2183]_ ) & (~\new_[3306]_  | ~\new_[496]_ );
  assign \new_[717]_  = (~\new_[815]_  | ~\new_[2180]_ ) & (~\new_[2558]_  | ~\new_[497]_ );
  assign \new_[718]_  = (~\new_[816]_  | ~\new_[2182]_ ) & (~\new_[2625]_  | ~\new_[488]_ );
  assign \new_[719]_  = (~\new_[817]_  | ~\new_[2182]_ ) & (~\new_[3311]_  | ~\new_[486]_ );
  assign \new_[720]_  = (~\new_[819]_  | ~\new_[2183]_ ) & (~\new_[2632]_  | ~\new_[502]_ );
  assign \new_[721]_  = (~\new_[818]_  | ~\new_[2183]_ ) & (~\new_[2626]_  | ~\new_[499]_ );
  assign \new_[722]_  = (~\new_[820]_  | ~\new_[3310]_ ) & (~\new_[3306]_  | ~\new_[482]_ );
  assign \new_[723]_  = (~\new_[821]_  | ~\new_[3310]_ ) & (~\new_[2558]_  | ~\new_[500]_ );
  assign \new_[724]_  = (~\new_[822]_  | ~\new_[2098]_ ) & (~\new_[2626]_  | ~\new_[501]_ );
  assign \new_[725]_  = (~\new_[823]_  | ~\new_[2097]_ ) & (~\new_[2626]_  | ~\new_[503]_ );
  assign \new_[726]_  = (~\new_[824]_  | ~\new_[2183]_ ) & (~\new_[2625]_  | ~\new_[474]_ );
  assign \new_[727]_  = ~\new_[2479]_  | (~\new_[825]_  & ~\new_[3364]_ );
  assign \new_[728]_  = ~\new_[2480]_  | (~\new_[826]_  & ~\new_[3364]_ );
  assign \new_[729]_  = ~\new_[2481]_  | (~\new_[827]_  & ~\new_[3364]_ );
  assign \new_[730]_  = ~\new_[3292]_  & (~\new_[2103]_  | ~\new_[844]_ );
  assign \new_[731]_  = ~\new_[2374]_  & (~\new_[2104]_  | ~\new_[845]_ );
  assign \new_[732]_  = ~\new_[3292]_  & (~\new_[2091]_  | ~\new_[846]_ );
  assign \new_[733]_  = ~\new_[3292]_  & (~\new_[2089]_  | ~\new_[847]_ );
  assign \new_[734]_  = ~\new_[3292]_  & (~\new_[2101]_  | ~\new_[848]_ );
  assign \new_[735]_  = ~\new_[2181]_  | (~\new_[849]_  & ~\new_[2583]_ );
  assign \new_[736]_  = ~\new_[3218]_  | (~\new_[850]_  & ~\new_[2536]_ );
  assign \new_[737]_  = ~\new_[2181]_  | (~\new_[851]_  & ~\new_[2543]_ );
  assign \new_[738]_  = ~\new_[2180]_  | (~\new_[852]_  & ~\new_[2545]_ );
  assign \new_[739]_  = ~\new_[2092]_  | (~\new_[895]_  & ~\new_[2276]_ );
  assign \new_[740]_  = ~\new_[2093]_  | (~\new_[896]_  & ~\new_[2276]_ );
  assign \new_[741]_  = ~\new_[2087]_  | (~\new_[897]_  & ~\new_[2276]_ );
  assign \new_[742]_  = ~\new_[2242]_  | ~\new_[885]_  | ~\new_[2194]_ ;
  assign \new_[743]_  = ~\new_[2241]_  | ~\new_[886]_  | ~\new_[2197]_ ;
  assign \new_[744]_  = ~\new_[2241]_  | ~\new_[887]_  | ~\new_[2202]_ ;
  assign \new_[745]_  = ~\new_[2242]_  | ~\new_[890]_  | ~\new_[2195]_ ;
  assign \new_[746]_  = ~\new_[2242]_  | ~\new_[891]_  | ~\new_[2201]_ ;
  assign \new_[747]_  = ~\new_[2241]_  | ~\new_[892]_  | ~\new_[2196]_ ;
  assign \new_[748]_  = ~\new_[2241]_  | ~\new_[893]_  | ~\new_[2199]_ ;
  assign \new_[749]_  = ~\new_[2242]_  | ~\new_[894]_  | ~\new_[2198]_ ;
  assign \new_[750]_  = ~\new_[3292]_  & (~\new_[2177]_  | ~\new_[866]_ );
  assign \new_[751]_  = ~\new_[2374]_  & (~\new_[2082]_  | ~\new_[867]_ );
  assign \new_[752]_  = ~\new_[3292]_  & (~\new_[2083]_  | ~\new_[868]_ );
  assign \new_[753]_  = ~\new_[2374]_  & (~\new_[2084]_  | ~\new_[869]_ );
  assign \new_[754]_  = ~\new_[3292]_  & (~\new_[2187]_  | ~\new_[870]_ );
  assign \new_[755]_  = ~\new_[3292]_  & (~\new_[2085]_  | ~\new_[871]_ );
  assign \new_[756]_  = ~\new_[3292]_  & (~\new_[2086]_  | ~\new_[872]_ );
  assign \new_[757]_  = ~\new_[2374]_  & (~\new_[2090]_  | ~\new_[873]_ );
  assign \new_[758]_  = ~\new_[3292]_  & (~\new_[2184]_  | ~\new_[874]_ );
  assign \new_[759]_  = ~\new_[3496]_  | (~\new_[3423]_  & ~\new_[2537]_ );
  assign \new_[760]_  = ~\new_[3292]_  & (~\new_[2100]_  | ~\new_[875]_ );
  assign \new_[761]_  = ~\new_[3496]_  | (~\new_[888]_  & ~\new_[2544]_ );
  assign \new_[762]_  = ~\new_[2098]_  | (~\new_[889]_  & ~\new_[2530]_ );
  assign \new_[763]_  = ~\new_[2374]_  & (~\new_[2102]_  | ~\new_[877]_ );
  assign \new_[764]_  = ~\new_[3292]_  & (~\new_[2088]_  | ~\new_[3294]_ );
  assign \new_[765]_  = ~\new_[3292]_  & (~\new_[2178]_  | ~\new_[880]_ );
  assign \new_[766]_  = ~\new_[2374]_  & (~\new_[2099]_  | ~\new_[881]_ );
  assign \new_[767]_  = ~\new_[3292]_  & (~\new_[2186]_  | ~\new_[882]_ );
  assign \new_[768]_  = ~\new_[2374]_  & (~\new_[2105]_  | ~\new_[883]_ );
  assign \new_[769]_  = ~\new_[3292]_  & (~\new_[2188]_  | ~\new_[884]_ );
  assign \new_[770]_  = \new_[933]_  ? \new_[2249]_  : \new_[424]_ ;
  assign \new_[771]_  = \new_[934]_  ? \new_[2276]_  : \new_[425]_ ;
  assign \new_[772]_  = \new_[935]_  ? \new_[2276]_  : \new_[426]_ ;
  assign \new_[773]_  = \new_[936]_  ? \new_[2276]_  : \new_[427]_ ;
  assign \new_[774]_  = \new_[937]_  ? \new_[2249]_  : \new_[428]_ ;
  assign \new_[775]_  = \new_[938]_  ? \new_[2249]_  : \new_[429]_ ;
  assign \new_[776]_  = \new_[939]_  ? \new_[2249]_  : \new_[430]_ ;
  assign \new_[777]_  = \new_[940]_  ? \new_[2276]_  : \new_[431]_ ;
  assign \new_[778]_  = \new_[942]_  ? \new_[2249]_  : \new_[432]_ ;
  assign \new_[779]_  = \new_[943]_  ? \new_[2249]_  : \new_[433]_ ;
  assign \new_[780]_  = \new_[944]_  ? \new_[2282]_  : \new_[434]_ ;
  assign \new_[781]_  = \new_[945]_  ? \new_[2249]_  : \new_[435]_ ;
  assign \new_[782]_  = \new_[946]_  ? \new_[2249]_  : \new_[436]_ ;
  assign \new_[783]_  = ~\new_[2367]_  & ~\new_[855]_ ;
  assign \new_[784]_  = ~\new_[2266]_  & ~\new_[856]_ ;
  assign \new_[785]_  = ~\new_[2267]_  & ~\new_[857]_ ;
  assign \new_[786]_  = ~\new_[2268]_  & ~\new_[858]_ ;
  assign \new_[787]_  = ~\new_[2270]_  & ~\new_[859]_ ;
  assign \new_[788]_  = ~\new_[2370]_  & ~\new_[860]_ ;
  assign \new_[789]_  = ~\new_[2271]_  & ~\new_[861]_ ;
  assign \new_[790]_  = ~\new_[2471]_  & ~\new_[862]_ ;
  assign \new_[791]_  = ~\new_[2472]_  & ~\new_[863]_ ;
  assign \new_[792]_  = ~\new_[2473]_  & ~\new_[864]_ ;
  assign \new_[793]_  = ~\new_[2278]_  & ~\new_[876]_ ;
  assign \new_[794]_  = ~\new_[2469]_  & ~\new_[878]_ ;
  assign \new_[795]_  = ~\new_[2277]_  & ~\new_[879]_ ;
  assign \new_[796]_  = ~\new_[2525]_  & ~\new_[865]_ ;
  assign \new_[797]_  = ~\new_[898]_  & ~\new_[2281]_ ;
  assign \new_[798]_  = ~\new_[899]_  & ~\new_[2283]_ ;
  assign \new_[799]_  = ~\new_[900]_  & ~\new_[2283]_ ;
  assign \new_[800]_  = ~\new_[901]_  & ~\new_[3214]_ ;
  assign \new_[801]_  = ~\new_[902]_  & ~\new_[2281]_ ;
  assign \new_[802]_  = ~\new_[903]_  & ~\new_[2281]_ ;
  assign \new_[803]_  = ~\new_[907]_  & ~\new_[2283]_ ;
  assign \new_[804]_  = ~\new_[904]_  & ~\new_[2283]_ ;
  assign \new_[805]_  = ~\new_[905]_  & ~\new_[3214]_ ;
  assign \new_[806]_  = ~\new_[906]_  & ~\new_[3214]_ ;
  assign \new_[807]_  = ~\new_[908]_  & ~\new_[3214]_ ;
  assign \new_[808]_  = ~\new_[2275]_  & ~\new_[910]_ ;
  assign \new_[809]_  = ~\new_[2264]_  & ~\new_[909]_ ;
  assign \new_[810]_  = ~\new_[931]_  & ~\new_[2283]_ ;
  assign \new_[811]_  = ~\new_[3424]_  & ~\new_[929]_ ;
  assign \new_[812]_  = ~\new_[932]_  & ~\new_[2283]_ ;
  assign \new_[813]_  = ~\new_[930]_  & ~\new_[3424]_ ;
  assign \new_[814]_  = \new_[955]_  ? \new_[2276]_  : \new_[496]_ ;
  assign \new_[815]_  = \new_[956]_  ? \new_[2276]_  : \new_[497]_ ;
  assign \new_[816]_  = \new_[957]_  ? \new_[2249]_  : \new_[488]_ ;
  assign \new_[817]_  = \new_[958]_  ? \new_[2249]_  : \new_[486]_ ;
  assign \new_[818]_  = \new_[959]_  ? \new_[2249]_  : \new_[499]_ ;
  assign \new_[819]_  = \new_[960]_  ? \new_[2249]_  : \new_[502]_ ;
  assign \new_[820]_  = \new_[961]_  ? \new_[2249]_  : \new_[482]_ ;
  assign \new_[821]_  = \new_[962]_  ? \new_[2282]_  : \new_[500]_ ;
  assign \new_[822]_  = \new_[963]_  ? \new_[2249]_  : \new_[501]_ ;
  assign \new_[823]_  = \new_[964]_  ? \new_[2249]_  : \new_[503]_ ;
  assign \new_[824]_  = \new_[965]_  ? \new_[2276]_  : \new_[474]_ ;
  assign \new_[825]_  = ~\new_[2364]_  & ~\new_[911]_ ;
  assign \new_[826]_  = ~\new_[2365]_  & ~\new_[925]_ ;
  assign \new_[827]_  = ~\new_[2366]_  & ~\new_[912]_ ;
  assign \new_[828]_  = ~\new_[2265]_  & ~\new_[913]_ ;
  assign \new_[829]_  = ~\new_[2368]_  & ~\new_[926]_ ;
  assign \new_[830]_  = ~\new_[2475]_  & ~\new_[914]_ ;
  assign \new_[831]_  = ~\new_[2468]_  & ~\new_[3220]_ ;
  assign \new_[832]_  = ~\new_[2269]_  & ~\new_[915]_ ;
  assign \new_[833]_  = ~\new_[2369]_  & ~\new_[916]_ ;
  assign \new_[834]_  = ~\new_[2467]_  & ~\new_[927]_ ;
  assign \new_[835]_  = ~\new_[2272]_  & ~\new_[928]_ ;
  assign \new_[836]_  = ~\new_[2375]_  & ~\new_[917]_ ;
  assign \new_[837]_  = ~\new_[2273]_  & ~\new_[918]_ ;
  assign \new_[838]_  = ~\new_[2470]_  & ~\new_[919]_ ;
  assign \new_[839]_  = ~\new_[2376]_  & ~\new_[920]_ ;
  assign \new_[840]_  = ~\new_[2274]_  & ~\new_[921]_ ;
  assign \new_[841]_  = ~\new_[2477]_  & ~\new_[922]_ ;
  assign \new_[842]_  = ~\new_[2474]_  & ~\new_[923]_ ;
  assign \new_[843]_  = ~\new_[2476]_  & ~\new_[924]_ ;
  assign \new_[844]_  = ~\new_[973]_  | ~\new_[2372]_  | ~\new_[1084]_ ;
  assign \new_[845]_  = ~\new_[966]_  | ~\new_[2372]_  | ~\new_[1100]_ ;
  assign \new_[846]_  = ~\new_[980]_  | ~\new_[2372]_  | ~\new_[1162]_ ;
  assign \new_[847]_  = ~\new_[981]_  | ~\new_[2372]_  | ~\new_[1163]_ ;
  assign \new_[848]_  = ~\new_[982]_  | ~\new_[2372]_  | ~\new_[1164]_ ;
  assign \new_[849]_  = ~\new_[941]_  & ~\new_[3424]_ ;
  assign \new_[850]_  = ~\new_[947]_  & ~\new_[2281]_ ;
  assign \new_[851]_  = ~\new_[3424]_  & ~\new_[948]_ ;
  assign \new_[852]_  = ~\new_[949]_  & ~\new_[3214]_ ;
  assign \new_[853]_  = ~\new_[950]_  & ~\new_[3424]_ ;
  assign \new_[854]_  = ~\new_[3424]_  & ~\new_[951]_ ;
  assign \new_[855]_  = ~\new_[2600]_  & (~\new_[1157]_  | ~\new_[1011]_ );
  assign \new_[856]_  = ~\new_[2591]_  & (~\new_[999]_  | ~\new_[1110]_ );
  assign \new_[857]_  = ~\new_[3225]_  & (~\new_[1001]_  | ~\new_[1112]_ );
  assign \new_[858]_  = ~\new_[2578]_  & (~\new_[1014]_  | ~\new_[1137]_ );
  assign \new_[859]_  = ~\new_[2577]_  & (~\new_[1117]_  | ~\new_[1015]_ );
  assign \new_[860]_  = ~\new_[2591]_  & (~\new_[1138]_  | ~\new_[1017]_ );
  assign \new_[861]_  = ~\new_[3225]_  & (~\new_[1018]_  | ~\new_[1119]_ );
  assign \new_[862]_  = ~\new_[2600]_  & (~\new_[1021]_  | ~\new_[1197]_ );
  assign \new_[863]_  = ~\new_[2600]_  & (~\new_[1198]_  | ~\new_[1022]_ );
  assign \new_[864]_  = ~\new_[2600]_  & (~\new_[1023]_  | ~\new_[1125]_ );
  assign \new_[865]_  = ~\new_[2578]_  & (~\new_[1141]_  | ~\new_[1026]_ );
  assign \new_[866]_  = ~\new_[988]_  | ~\new_[3298]_  | ~\new_[1132]_ ;
  assign \new_[867]_  = ~\new_[989]_  | ~\new_[3298]_  | ~\new_[1133]_ ;
  assign \new_[868]_  = ~\new_[1002]_  | ~\new_[3298]_  | ~\new_[1147]_ ;
  assign \new_[869]_  = ~\new_[990]_  | ~\new_[3298]_  | ~\new_[1134]_ ;
  assign \new_[870]_  = ~\new_[1003]_  | ~\new_[3298]_  | ~\new_[1148]_ ;
  assign \new_[871]_  = ~\new_[1005]_  | ~\new_[3298]_  | ~\new_[1149]_ ;
  assign \new_[872]_  = ~\new_[3298]_  | ~\new_[1006]_  | ~\new_[1209]_ ;
  assign \new_[873]_  = ~\new_[3298]_  | ~\new_[1007]_  | ~\new_[1077]_ ;
  assign \new_[874]_  = ~\new_[1000]_  | ~\new_[3298]_  | ~\new_[1111]_ ;
  assign \new_[875]_  = ~\new_[3298]_  | ~\new_[1013]_  | ~\new_[1114]_ ;
  assign \new_[876]_  = ~\new_[2577]_  & (~\new_[993]_  | ~\new_[1107]_ );
  assign \new_[877]_  = ~\new_[3298]_  | ~\new_[1025]_  | ~\new_[1085]_ ;
  assign \new_[878]_  = ~\new_[2577]_  & (~\new_[994]_  | ~\new_[1108]_ );
  assign \new_[879]_  = ~\new_[2577]_  & (~\new_[1109]_  | ~\new_[995]_ );
  assign \new_[880]_  = ~\new_[991]_  | ~\new_[3298]_  | ~\new_[1135]_ ;
  assign \new_[881]_  = ~\new_[992]_  | ~\new_[3298]_  | ~\new_[1101]_ ;
  assign \new_[882]_  = ~\new_[997]_  | ~\new_[3298]_  | ~\new_[1103]_ ;
  assign \new_[883]_  = ~\new_[3298]_  | ~\new_[1034]_  | ~\new_[1106]_ ;
  assign \new_[884]_  = ~\new_[3298]_  | ~\new_[987]_  | ~\new_[1225]_ ;
  assign \new_[885]_  = ~\new_[2514]_  | ~\new_[1004]_  | ~\new_[1208]_ ;
  assign \new_[886]_  = ~\new_[2514]_  | ~\new_[1019]_  | ~\new_[1212]_ ;
  assign \new_[887]_  = ~\new_[2524]_  | ~\new_[1008]_  | ~\new_[1211]_ ;
  assign \new_[888]_  = ~\new_[3253]_  & ~\new_[3214]_ ;
  assign \new_[889]_  = ~\new_[3299]_  & ~\new_[3214]_ ;
  assign \new_[890]_  = ~\new_[2524]_  | ~\new_[1024]_  | ~\new_[1217]_ ;
  assign \new_[891]_  = ~\new_[2514]_  | ~\new_[996]_  | ~\new_[1207]_ ;
  assign \new_[892]_  = ~\new_[2514]_  | ~\new_[1032]_  | ~\new_[1131]_ ;
  assign \new_[893]_  = ~\new_[2524]_  | ~\new_[1033]_  | ~\new_[1218]_ ;
  assign \new_[894]_  = ~\new_[2524]_  | ~\new_[998]_  | ~\new_[1192]_ ;
  assign \new_[895]_  = ~\new_[967]_  | (~\new_[1294]_  & ~\new_[394]_ );
  assign \new_[896]_  = ~\new_[968]_  | (~\new_[1295]_  & ~\new_[392]_ );
  assign \new_[897]_  = ~\new_[969]_  | (~\new_[1296]_  & ~\new_[393]_ );
  assign \new_[898]_  = ~\new_[970]_  & (~\new_[1266]_  | ~\new_[437]_ );
  assign \new_[899]_  = ~\new_[971]_  & (~\new_[1159]_  | ~\new_[438]_ );
  assign \new_[900]_  = ~\new_[972]_  & (~\new_[1368]_  | ~\new_[439]_ );
  assign \new_[901]_  = ~\new_[974]_  & (~\new_[1370]_  | ~\new_[440]_ );
  assign \new_[902]_  = ~\new_[976]_  & (~\new_[1097]_  | ~\new_[441]_ );
  assign \new_[903]_  = ~\new_[975]_  & (~\new_[1242]_  | ~\new_[442]_ );
  assign \new_[904]_  = ~\new_[977]_  & (~\new_[1371]_  | ~\new_[443]_ );
  assign \new_[905]_  = ~\new_[978]_  & (~\new_[1372]_  | ~\new_[444]_ );
  assign \new_[906]_  = ~\new_[979]_  & (~\new_[1373]_  | ~\new_[445]_ );
  assign \new_[907]_  = (~\new_[1035]_  | ~\new_[1080]_ ) & (~\new_[1098]_  | ~\new_[446]_ );
  assign \new_[908]_  = (~\new_[1035]_  | ~\new_[1332]_ ) & (~\new_[1369]_  | ~\new_[447]_ );
  assign \new_[909]_  = ~\new_[2591]_  & (~\new_[1038]_  | ~\new_[1081]_ );
  assign \new_[910]_  = ~\new_[2600]_  & (~\new_[1036]_  | ~\new_[1037]_ );
  assign \new_[911]_  = ~\new_[2596]_  & (~\new_[1043]_  | ~\new_[1193]_ );
  assign \new_[912]_  = ~\new_[2596]_  & (~\new_[1044]_  | ~\new_[1153]_ );
  assign \new_[913]_  = ~\new_[2600]_  & (~\new_[1046]_  | ~\new_[1213]_ );
  assign \new_[914]_  = ~\new_[2591]_  & (~\new_[1047]_  | ~\new_[1113]_ );
  assign \new_[915]_  = ~\new_[2600]_  & (~\new_[1048]_  | ~\new_[1115]_ );
  assign \new_[916]_  = ~\new_[2577]_  & (~\new_[1049]_  | ~\new_[1116]_ );
  assign \new_[917]_  = ~\new_[2578]_  & (~\new_[1050]_  | ~\new_[1235]_ );
  assign \new_[918]_  = ~\new_[2591]_  & (~\new_[1051]_  | ~\new_[1161]_ );
  assign \new_[919]_  = ~\new_[2591]_  & (~\new_[1052]_  | ~\new_[1268]_ );
  assign \new_[920]_  = ~\new_[2591]_  & (~\new_[1269]_  | ~\new_[1053]_ );
  assign \new_[921]_  = ~\new_[3225]_  & (~\new_[1054]_  | ~\new_[1196]_ );
  assign \new_[922]_  = ~\new_[2577]_  & (~\new_[1055]_  | ~\new_[1270]_ );
  assign \new_[923]_  = ~\new_[2600]_  & (~\new_[1056]_  | ~\new_[1139]_ );
  assign \new_[924]_  = ~\new_[2578]_  & (~\new_[1057]_  | ~\new_[1104]_ );
  assign \new_[925]_  = ~\new_[2596]_  & (~\new_[1039]_  | ~\new_[1206]_ );
  assign \new_[926]_  = ~\new_[2577]_  & (~\new_[1040]_  | ~\new_[1064]_ );
  assign \new_[927]_  = ~\new_[2577]_  & (~\new_[1041]_  | ~\new_[1086]_ );
  assign \new_[928]_  = ~\new_[2591]_  & (~\new_[1042]_  | ~\new_[1087]_ );
  assign \new_[929]_  = ~\new_[985]_  & (~\new_[1129]_  | ~\new_[495]_ );
  assign \new_[930]_  = ~\new_[986]_  & (~\new_[1191]_  | ~\new_[498]_ );
  assign \new_[931]_  = ~\new_[983]_  & (~\new_[1128]_  | ~\new_[493]_ );
  assign \new_[932]_  = ~\new_[984]_  & (~\new_[1190]_  | ~\new_[494]_ );
  assign \new_[933]_  = ~\new_[1146]_  & (~\new_[1058]_  | ~\new_[1292]_ );
  assign \new_[934]_  = ~\new_[1150]_  & (~\new_[1058]_  | ~\new_[3232]_ );
  assign \new_[935]_  = ~\new_[1083]_  & (~\new_[1061]_  | ~\new_[1143]_ );
  assign \new_[936]_  = ~\new_[1151]_  & (~\new_[1058]_  | ~\new_[1247]_ );
  assign \new_[937]_  = ~\new_[1260]_  & (~\new_[1058]_  | ~\new_[1378]_ );
  assign \new_[938]_  = ~\new_[1261]_  & (~\new_[1058]_  | ~\new_[1379]_ );
  assign \new_[939]_  = ~\new_[1262]_  & (~\new_[1062]_  | ~\new_[1380]_ );
  assign \new_[940]_  = ~\new_[1152]_  & (~\new_[1062]_  | ~\new_[1293]_ );
  assign \new_[941]_  = ~\new_[1009]_  & (~\new_[1229]_  | ~\new_[506]_ );
  assign \new_[942]_  = ~\new_[1078]_  & (~\new_[1058]_  | ~\new_[1122]_ );
  assign \new_[943]_  = ~\new_[1093]_  & (~\new_[1062]_  | ~\new_[1165]_ );
  assign \new_[944]_  = ~\new_[1154]_  & (~\new_[1058]_  | ~\new_[1297]_ );
  assign \new_[945]_  = ~\new_[1155]_  & (~\new_[1062]_  | ~\new_[1298]_ );
  assign \new_[946]_  = ~\new_[1156]_  & (~\new_[1058]_  | ~\new_[1299]_ );
  assign \new_[947]_  = ~\new_[1012]_  & (~\new_[1254]_  | ~\new_[507]_ );
  assign \new_[948]_  = ~\new_[1020]_  & (~\new_[1325]_  | ~\new_[468]_ );
  assign \new_[949]_  = ~\new_[1027]_  & (~\new_[1241]_  | ~\new_[508]_ );
  assign \new_[950]_  = ~\new_[1028]_  & (~\new_[1175]_  | ~\new_[465]_ );
  assign \new_[951]_  = ~\new_[1029]_  & (~\new_[1224]_  | ~\new_[509]_ );
  assign \new_[952]_  = (~\new_[1067]_  | ~\new_[1126]_ ) & (~\new_[1181]_  | ~\new_[3305]_ );
  assign \new_[953]_  = (~\new_[3430]_  | ~\new_[1226]_ ) & (~\new_[1287]_  | ~\new_[560]_ );
  assign \new_[954]_  = (~\new_[3430]_  | ~\new_[1227]_ ) & (~\new_[1288]_  | ~\new_[561]_ );
  assign \new_[955]_  = (~\new_[1067]_  | ~\new_[1258]_ ) & (~\new_[1327]_  | ~\new_[3179]_ );
  assign \new_[956]_  = (~\new_[1067]_  | ~\new_[1136]_ ) & (~\new_[1194]_  | ~\new_[3128]_ );
  assign \new_[957]_  = (~\new_[1067]_  | ~\new_[1127]_ ) & (~\new_[1183]_  | ~\new_[3153]_ );
  assign \new_[958]_  = (~\new_[1067]_  | ~\new_[1210]_ ) & (~\new_[1259]_  | ~\new_[3194]_ );
  assign \new_[959]_  = (~\new_[1067]_  | ~\new_[1222]_ ) & (~\new_[1281]_  | ~\new_[3160]_ );
  assign \new_[960]_  = (~\new_[1067]_  | ~\new_[1219]_ ) & (~\new_[1275]_  | ~\new_[3200]_ );
  assign \new_[961]_  = (~\new_[1067]_  | ~\new_[1249]_ ) & (~\new_[1310]_  | ~\new_[3169]_ );
  assign \new_[962]_  = (~\new_[1067]_  | ~\new_[1263]_ ) & (~\new_[1328]_  | ~\new_[3144]_ );
  assign \new_[963]_  = (~\new_[1067]_  | ~\new_[1282]_ ) & (~\new_[1339]_  | ~\new_[3114]_ );
  assign \new_[964]_  = (~\new_[1067]_  | ~\new_[1276]_ ) & (~\new_[1336]_  | ~\new_[3185]_ );
  assign \new_[965]_  = (~\new_[1067]_  | ~\new_[1079]_ ) & (~\new_[1094]_  | ~\new_[3133]_ );
  assign \new_[966]_  = ~\new_[1063]_  | ~\new_[1142]_ ;
  assign \new_[967]_  = ~\new_[1060]_  | ~\new_[1294]_ ;
  assign \new_[968]_  = ~\new_[1060]_  | ~\new_[1295]_ ;
  assign \new_[969]_  = ~\new_[1060]_  | ~\new_[1296]_ ;
  assign \new_[970]_  = ~\new_[1059]_  & ~\new_[1266]_ ;
  assign \new_[971]_  = ~\new_[1061]_  & ~\new_[1159]_ ;
  assign \new_[972]_  = ~\new_[1061]_  & ~\new_[1368]_ ;
  assign \new_[973]_  = ~\new_[1063]_  | ~\new_[1144]_ ;
  assign \new_[974]_  = ~\new_[1059]_  & ~\new_[1370]_ ;
  assign \new_[975]_  = ~\new_[1061]_  & ~\new_[1242]_ ;
  assign \new_[976]_  = ~\new_[1059]_  & ~\new_[1097]_ ;
  assign \new_[977]_  = ~\new_[1061]_  & ~\new_[1371]_ ;
  assign \new_[978]_  = ~\new_[1061]_  & ~\new_[1372]_ ;
  assign \new_[979]_  = ~\new_[1059]_  & ~\new_[1373]_ ;
  assign \new_[980]_  = ~\new_[1063]_  | ~\new_[1243]_ ;
  assign \new_[981]_  = ~\new_[1063]_  | ~\new_[1244]_ ;
  assign \new_[982]_  = ~\new_[1063]_  | ~\new_[1245]_ ;
  assign \new_[983]_  = ~\new_[1068]_  & ~\new_[1128]_ ;
  assign \new_[984]_  = ~\new_[1069]_  & ~\new_[1190]_ ;
  assign \new_[985]_  = ~\new_[1068]_  & ~\new_[1129]_ ;
  assign \new_[986]_  = ~\new_[1069]_  & ~\new_[1191]_ ;
  assign \new_[987]_  = ~\new_[1065]_  | ~\new_[1312]_ ;
  assign \new_[988]_  = ~\new_[1075]_  | ~\new_[1255]_ ;
  assign \new_[989]_  = ~\new_[1075]_  | ~\new_[1280]_ ;
  assign \new_[990]_  = ~\new_[1075]_  | ~\new_[1274]_ ;
  assign \new_[991]_  = ~\new_[1075]_  | ~\new_[1273]_ ;
  assign \new_[992]_  = ~\new_[1075]_  | ~\new_[1203]_ ;
  assign \new_[993]_  = ~\new_[1071]_  | ~\new_[1238]_ ;
  assign \new_[994]_  = ~\new_[1071]_  | ~\new_[1239]_ ;
  assign \new_[995]_  = ~\new_[1076]_  | ~\new_[1240]_ ;
  assign \new_[996]_  = ~\new_[1070]_  | ~\new_[1308]_ ;
  assign \new_[997]_  = ~\new_[1065]_  | ~\new_[1204]_ ;
  assign \new_[998]_  = ~\new_[1070]_  | ~\new_[1335]_ ;
  assign \new_[999]_  = ~\new_[1071]_  | ~\new_[1246]_ ;
  assign \new_[1000]_  = ~\new_[1075]_  | ~\new_[1178]_ ;
  assign \new_[1001]_  = ~\new_[1076]_  | ~\new_[1248]_ ;
  assign \new_[1002]_  = ~\new_[1066]_  | ~\new_[1289]_ ;
  assign \new_[1003]_  = ~\new_[1075]_  | ~\new_[1290]_ ;
  assign \new_[1004]_  = ~\new_[1070]_  | ~\new_[1343]_ ;
  assign \new_[1005]_  = ~\new_[1066]_  | ~\new_[1291]_ ;
  assign \new_[1006]_  = ~\new_[1065]_  | ~\new_[1344]_ ;
  assign \new_[1007]_  = ~\new_[1065]_  | ~\new_[1099]_ ;
  assign \new_[1008]_  = ~\new_[1070]_  | ~\new_[1346]_ ;
  assign \new_[1009]_  = ~\new_[1069]_  & ~\new_[1229]_ ;
  assign \new_[1010]_  = ~\new_[1068]_  & ~\new_[1250]_ ;
  assign \new_[1011]_  = ~\new_[1076]_  | ~\new_[1230]_ ;
  assign \new_[1012]_  = ~\new_[1068]_  & ~\new_[1254]_ ;
  assign \new_[1013]_  = ~\new_[1066]_  | ~\new_[1232]_ ;
  assign \new_[1014]_  = ~\new_[1071]_  | ~\new_[1220]_ ;
  assign \new_[1015]_  = ~\new_[1076]_  | ~\new_[1123]_ ;
  assign \new_[1016]_  = ~\new_[1066]_  | ~\new_[1177]_ ;
  assign \new_[1017]_  = ~\new_[1076]_  | ~\new_[1223]_ ;
  assign \new_[1018]_  = ~\new_[1076]_  | ~\new_[1124]_ ;
  assign \new_[1019]_  = ~\new_[1070]_  | ~\new_[1347]_ ;
  assign \new_[1020]_  = ~\new_[1068]_  & ~\new_[1325]_ ;
  assign \new_[1021]_  = ~\new_[1071]_  | ~\new_[1285]_ ;
  assign \new_[1022]_  = ~\new_[1076]_  | ~\new_[1286]_ ;
  assign \new_[1023]_  = ~\new_[1071]_  | ~\new_[1185]_ ;
  assign \new_[1024]_  = ~\new_[1070]_  | ~\new_[1307]_ ;
  assign \new_[1025]_  = ~\new_[1065]_  | ~\new_[1145]_ ;
  assign \new_[1026]_  = ~\new_[1076]_  | ~\new_[1221]_ ;
  assign \new_[1027]_  = ~\new_[1069]_  & ~\new_[1241]_ ;
  assign \new_[1028]_  = ~\new_[1069]_  & ~\new_[1175]_ ;
  assign \new_[1029]_  = ~\new_[1068]_  & ~\new_[1224]_ ;
  assign \new_[1030]_  = ~\new_[1068]_  & ~\new_[1095]_ ;
  assign \new_[1031]_  = ~\new_[1066]_  | ~\new_[1180]_ ;
  assign \new_[1032]_  = ~\new_[1070]_  | ~\new_[1202]_ ;
  assign \new_[1033]_  = ~\new_[1070]_  | ~\new_[1309]_ ;
  assign \new_[1034]_  = ~\new_[1065]_  | ~\new_[1205]_ ;
  assign \new_[1035]_  = ~\new_[1062]_ ;
  assign \new_[1036]_  = ~\new_[1082]_  | ~\new_[356]_ ;
  assign \new_[1037]_  = ~\new_[1089]_  | ~\new_[1102]_ ;
  assign \new_[1038]_  = ~\new_[1088]_  | ~\new_[1105]_ ;
  assign \new_[1039]_  = ~\new_[3428]_  | ~\new_[1377]_ ;
  assign \new_[1040]_  = ~\new_[1088]_  | ~\new_[1121]_ ;
  assign \new_[1041]_  = ~\new_[1088]_  | ~\new_[1214]_ ;
  assign \new_[1042]_  = ~\new_[1088]_  | ~\new_[1215]_ ;
  assign \new_[1043]_  = ~\new_[3428]_  | ~\new_[1256]_ ;
  assign \new_[1044]_  = ~\new_[3428]_  | ~\new_[1228]_ ;
  assign \new_[1045]_  = ~\new_[3428]_  | ~\new_[1277]_ ;
  assign \new_[1046]_  = ~\new_[1088]_  | ~\new_[1300]_ ;
  assign \new_[1047]_  = ~\new_[1088]_  | ~\new_[1166]_ ;
  assign \new_[1048]_  = ~\new_[1088]_  | ~\new_[1167]_ ;
  assign \new_[1049]_  = ~\new_[1088]_  | ~\new_[1168]_ ;
  assign \new_[1050]_  = ~\new_[1088]_  | ~\new_[1311]_ ;
  assign \new_[1051]_  = ~\new_[1088]_  | ~\new_[1303]_ ;
  assign \new_[1052]_  = ~\new_[1088]_  | ~\new_[1304]_ ;
  assign \new_[1053]_  = ~\new_[1089]_  | ~\new_[1305]_ ;
  assign \new_[1054]_  = ~\new_[1088]_  | ~\new_[1284]_ ;
  assign \new_[1055]_  = ~\new_[1088]_  | ~\new_[1306]_ ;
  assign \new_[1056]_  = ~\new_[1088]_  | ~\new_[1216]_ ;
  assign \new_[1057]_  = ~\new_[1088]_  | ~\new_[1140]_ ;
  assign \new_[1058]_  = ~\new_[1072]_ ;
  assign \new_[1059]_  = ~\new_[1072]_ ;
  assign \new_[1060]_  = ~\new_[1073]_ ;
  assign \new_[1061]_  = ~\new_[1073]_ ;
  assign \new_[1062]_  = ~\new_[1074]_ ;
  assign \new_[1063]_  = ~\new_[1074]_ ;
  assign \new_[1064]_  = ~\new_[1096]_  | ~\new_[358]_ ;
  assign \new_[1065]_  = ~\new_[3428]_ ;
  assign \new_[1066]_  = ~\new_[3428]_ ;
  assign \new_[1067]_  = ~\new_[1089]_ ;
  assign \new_[1068]_  = ~\new_[1090]_ ;
  assign \new_[1069]_  = ~\new_[1090]_ ;
  assign \new_[1070]_  = ~\new_[1091]_ ;
  assign \new_[1071]_  = ~\new_[1091]_ ;
  assign \new_[1072]_  = ~\new_[1092]_ ;
  assign \new_[1073]_  = ~\new_[1092]_ ;
  assign \new_[1074]_  = ~\new_[1092]_ ;
  assign \new_[1075]_  = \new_[1092]_ ;
  assign \new_[1076]_  = ~\new_[1092]_ ;
  assign \new_[1077]_  = \new_[1099]_  | \new_[381]_ ;
  assign \new_[1078]_  = ~\new_[1122]_  & ~\new_[432]_ ;
  assign \new_[1079]_  = ~\new_[1094]_ ;
  assign \new_[1080]_  = ~\new_[1098]_ ;
  assign \new_[1081]_  = ~\new_[1130]_  | ~\new_[355]_ ;
  assign \new_[1082]_  = ~\new_[1102]_ ;
  assign \new_[1083]_  = ~\new_[1143]_  & ~\new_[426]_ ;
  assign \new_[1084]_  = \new_[1144]_  | \new_[345]_ ;
  assign \new_[1085]_  = \new_[1145]_  | \new_[387]_ ;
  assign \new_[1086]_  = ~\new_[1158]_  | ~\new_[363]_ ;
  assign \new_[1087]_  = ~\new_[1160]_  | ~\new_[372]_ ;
  assign \new_[1088]_  = \new_[3429]_ ;
  assign \new_[1089]_  = \new_[3429]_ ;
  assign \new_[1090]_  = \new_[3429]_ ;
  assign \new_[1091]_  = ~\new_[3429]_ ;
  assign \new_[1092]_  = ~\new_[3429]_ ;
  assign \new_[1093]_  = ~\new_[1165]_  & ~\new_[433]_ ;
  assign \new_[1094]_  = ~\new_[1424]_  | ~\new_[1699]_  | ~\new_[1188]_ ;
  assign \new_[1095]_  = ~\new_[3276]_  | ~\new_[3406]_  | ~\new_[1188]_ ;
  assign \new_[1096]_  = ~\new_[1121]_ ;
  assign \new_[1097]_  = ~\new_[1186]_  | ~\new_[1381]_ ;
  assign \new_[1098]_  = ~\new_[1187]_  | ~\new_[1381]_ ;
  assign \new_[1099]_  = ~\new_[1182]_  & ~\new_[1699]_ ;
  assign \new_[1100]_  = ~\new_[1201]_  | ~\new_[3152]_ ;
  assign \new_[1101]_  = \new_[1203]_  | \new_[389]_ ;
  assign \new_[1102]_  = \new_[1199]_  & \new_[1768]_ ;
  assign \new_[1103]_  = \new_[1204]_  | \new_[390]_ ;
  assign \new_[1104]_  = ~\new_[1200]_  | ~\new_[370]_ ;
  assign \new_[1105]_  = ~\new_[1130]_ ;
  assign \new_[1106]_  = \new_[1205]_  | \new_[391]_ ;
  assign \new_[1107]_  = ~\new_[1172]_  | ~\new_[338]_ ;
  assign \new_[1108]_  = ~\new_[1173]_  | ~\new_[339]_ ;
  assign \new_[1109]_  = ~\new_[1174]_  | ~\new_[340]_ ;
  assign \new_[1110]_  = ~\new_[1176]_  | ~\new_[329]_ ;
  assign \new_[1111]_  = \new_[1178]_  | \new_[382]_ ;
  assign \new_[1112]_  = ~\new_[1179]_  | ~\new_[330]_ ;
  assign \new_[1113]_  = ~\new_[1231]_  | ~\new_[359]_ ;
  assign \new_[1114]_  = \new_[1232]_  | \new_[384]_ ;
  assign \new_[1115]_  = ~\new_[1233]_  | ~\new_[361]_ ;
  assign \new_[1116]_  = ~\new_[1234]_  | ~\new_[362]_ ;
  assign \new_[1117]_  = ~\new_[1169]_  | ~\new_[332]_ ;
  assign \new_[1118]_  = \new_[1177]_  | \new_[380]_ ;
  assign \new_[1119]_  = ~\new_[1170]_  | ~\new_[334]_ ;
  assign \new_[1120]_  = \new_[1180]_  | \new_[385]_ ;
  assign \new_[1121]_  = ~\new_[1184]_  & ~\new_[1699]_ ;
  assign \new_[1122]_  = \new_[1186]_  & \new_[3273]_ ;
  assign \new_[1123]_  = ~\new_[1169]_ ;
  assign \new_[1124]_  = ~\new_[1170]_ ;
  assign \new_[1125]_  = ~\new_[1251]_  | ~\new_[337]_ ;
  assign \new_[1126]_  = ~\new_[1181]_ ;
  assign \new_[1127]_  = ~\new_[1183]_ ;
  assign \new_[1128]_  = ~\new_[1418]_  | ~\new_[1768]_  | ~\new_[1331]_ ;
  assign \new_[1129]_  = ~\new_[1324]_  | ~\new_[3406]_  | ~\new_[1331]_ ;
  assign \new_[1130]_  = ~\new_[1426]_  | ~\new_[1699]_  | ~\new_[3205]_ ;
  assign \new_[1131]_  = ~\new_[1253]_  | ~\new_[349]_ ;
  assign \new_[1132]_  = \new_[1255]_  | \new_[383]_ ;
  assign \new_[1133]_  = \new_[1280]_  | \new_[373]_ ;
  assign \new_[1134]_  = \new_[1274]_  | \new_[377]_ ;
  assign \new_[1135]_  = \new_[1273]_  | \new_[386]_ ;
  assign \new_[1136]_  = ~\new_[1194]_ ;
  assign \new_[1137]_  = ~\new_[1278]_  | ~\new_[331]_ ;
  assign \new_[1138]_  = ~\new_[1283]_  | ~\new_[333]_ ;
  assign \new_[1139]_  = ~\new_[1271]_  | ~\new_[368]_ ;
  assign \new_[1140]_  = ~\new_[1200]_ ;
  assign \new_[1141]_  = ~\new_[1279]_  | ~\new_[341]_ ;
  assign \new_[1142]_  = ~\new_[1201]_ ;
  assign \new_[1143]_  = ~\new_[1257]_  & ~\new_[1699]_ ;
  assign \new_[1144]_  = ~\new_[1267]_  & ~\new_[1699]_ ;
  assign \new_[1145]_  = ~\new_[1272]_  & ~\new_[1699]_ ;
  assign \new_[1146]_  = ~\new_[1292]_  & ~\new_[424]_ ;
  assign \new_[1147]_  = \new_[1289]_  | \new_[374]_ ;
  assign \new_[1148]_  = \new_[1290]_  | \new_[376]_ ;
  assign \new_[1149]_  = \new_[1291]_  | \new_[378]_ ;
  assign \new_[1150]_  = ~\new_[3232]_  & ~\new_[425]_ ;
  assign \new_[1151]_  = ~\new_[1247]_  & ~\new_[427]_ ;
  assign \new_[1152]_  = ~\new_[1293]_  & ~\new_[431]_ ;
  assign \new_[1153]_  = ~\new_[3270]_  | ~\new_[325]_ ;
  assign \new_[1154]_  = ~\new_[1297]_  & ~\new_[434]_ ;
  assign \new_[1155]_  = ~\new_[1298]_  & ~\new_[435]_ ;
  assign \new_[1156]_  = ~\new_[1299]_  & ~\new_[436]_ ;
  assign \new_[1157]_  = ~\new_[1301]_  | ~\new_[328]_ ;
  assign \new_[1158]_  = ~\new_[1214]_ ;
  assign \new_[1159]_  = ~\new_[1520]_  | ~\new_[1402]_  | ~\new_[1324]_ ;
  assign \new_[1160]_  = ~\new_[1215]_ ;
  assign \new_[1161]_  = ~\new_[1236]_  | ~\new_[364]_ ;
  assign \new_[1162]_  = \new_[1243]_  | \new_[350]_ ;
  assign \new_[1163]_  = \new_[1244]_  | \new_[351]_ ;
  assign \new_[1164]_  = \new_[1245]_  | \new_[353]_ ;
  assign \new_[1165]_  = ~\new_[1252]_  & ~\new_[1388]_ ;
  assign \new_[1166]_  = ~\new_[1231]_ ;
  assign \new_[1167]_  = ~\new_[1233]_ ;
  assign \new_[1168]_  = ~\new_[1234]_ ;
  assign \new_[1169]_  = ~\new_[1318]_  | ~\new_[1391]_ ;
  assign \new_[1170]_  = ~\new_[1319]_  | ~\new_[1391]_ ;
  assign \new_[1171]_  = ~\new_[1237]_ ;
  assign \new_[1172]_  = ~\new_[1238]_ ;
  assign \new_[1173]_  = ~\new_[1239]_ ;
  assign \new_[1174]_  = ~\new_[1240]_ ;
  assign \new_[1175]_  = ~\new_[1322]_  | ~\new_[1420]_ ;
  assign \new_[1176]_  = ~\new_[1246]_ ;
  assign \new_[1177]_  = \new_[1318]_  & \new_[1382]_ ;
  assign \new_[1178]_  = \new_[1320]_  & \new_[1405]_ ;
  assign \new_[1179]_  = ~\new_[1248]_ ;
  assign \new_[1180]_  = \new_[1319]_  & \new_[1382]_ ;
  assign \new_[1181]_  = \new_[1321]_  | \new_[3233]_ ;
  assign \new_[1182]_  = ~\new_[1316]_  | ~\new_[1424]_ ;
  assign \new_[1183]_  = ~\new_[1366]_  | ~\new_[1424]_  | ~\new_[1442]_ ;
  assign \new_[1184]_  = ~\new_[1316]_  | ~\new_[3276]_ ;
  assign \new_[1185]_  = ~\new_[1251]_ ;
  assign \new_[1186]_  = ~\new_[1699]_  & ~\new_[1315]_ ;
  assign \new_[1187]_  = ~\new_[1252]_ ;
  assign \new_[1188]_  = ~\new_[1315]_  & ~\new_[1478]_ ;
  assign mosi_pad_o = shift_s_out_reg;
  assign \new_[1190]_  = ~\new_[1470]_  | ~\new_[1768]_  | ~\new_[1367]_ ;
  assign \new_[1191]_  = ~\new_[1458]_  | ~\new_[3406]_  | ~\new_[1367]_ ;
  assign \new_[1192]_  = \new_[1335]_  | \new_[3195]_ ;
  assign \new_[1193]_  = ~\new_[1326]_  | ~\new_[327]_ ;
  assign \new_[1194]_  = ~\new_[1448]_  | ~\new_[1699]_  | ~\new_[1376]_ ;
  assign \new_[1195]_  = ~\new_[1337]_  | ~\new_[326]_ ;
  assign \new_[1196]_  = ~\new_[1340]_  | ~\new_[365]_ ;
  assign \new_[1197]_  = ~\new_[1341]_  | ~\new_[335]_ ;
  assign \new_[1198]_  = ~\new_[1342]_  | ~\new_[336]_ ;
  assign \new_[1199]_  = \new_[1443]_  & \new_[3205]_ ;
  assign \new_[1200]_  = ~\new_[1352]_  | ~\new_[1522]_  | ~\new_[1443]_ ;
  assign \new_[1201]_  = ~\new_[1353]_  | ~\new_[1699]_  | ~\new_[1473]_ ;
  assign \new_[1202]_  = ~\new_[1253]_ ;
  assign \new_[1203]_  = \new_[1333]_  & \new_[1520]_ ;
  assign \new_[1204]_  = ~\new_[1334]_  & ~\new_[1479]_ ;
  assign \new_[1205]_  = ~\new_[1334]_  & ~\new_[1519]_ ;
  assign \new_[1206]_  = ~\new_[1345]_  | ~\new_[324]_ ;
  assign \new_[1207]_  = \new_[1308]_  | \new_[3138]_ ;
  assign \new_[1208]_  = \new_[1343]_  | \new_[3176]_ ;
  assign \new_[1209]_  = \new_[1344]_  | \new_[379]_ ;
  assign \new_[1210]_  = ~\new_[1259]_ ;
  assign \new_[1211]_  = \new_[1346]_  | \new_[3199]_ ;
  assign \new_[1212]_  = \new_[1347]_  | \new_[3146]_ ;
  assign \new_[1213]_  = ~\new_[1348]_  | ~\new_[357]_ ;
  assign \new_[1214]_  = \new_[1302]_  & \new_[1465]_ ;
  assign \new_[1215]_  = \new_[1466]_  & \new_[1302]_ ;
  assign \new_[1216]_  = ~\new_[1271]_ ;
  assign \new_[1217]_  = \new_[1307]_  | \new_[3113]_ ;
  assign \new_[1218]_  = \new_[1309]_  | \new_[3139]_ ;
  assign \new_[1219]_  = ~\new_[1275]_ ;
  assign \new_[1220]_  = ~\new_[1278]_ ;
  assign \new_[1221]_  = ~\new_[1279]_ ;
  assign \new_[1222]_  = ~\new_[1281]_ ;
  assign \new_[1223]_  = ~\new_[1283]_ ;
  assign \new_[1224]_  = ~\new_[1520]_  | ~\new_[1389]_  | ~\new_[1478]_  | ~\new_[3315]_ ;
  assign \new_[1225]_  = \new_[1312]_  | \new_[375]_ ;
  assign \new_[1226]_  = ~\new_[1287]_ ;
  assign \new_[1227]_  = ~\new_[1288]_ ;
  assign \new_[1228]_  = ~\new_[3270]_ ;
  assign \new_[1229]_  = ~\new_[1323]_  | ~\new_[1420]_ ;
  assign \new_[1230]_  = ~\new_[1301]_ ;
  assign \new_[1231]_  = ~\new_[1320]_  | ~\new_[1390]_ ;
  assign \new_[1232]_  = \new_[1317]_  & \new_[1405]_ ;
  assign \new_[1233]_  = ~\new_[1366]_  | ~\new_[1419]_  | ~\new_[1459]_ ;
  assign \new_[1234]_  = ~\new_[1314]_  | ~\new_[1391]_ ;
  assign \new_[1235]_  = ~\new_[1357]_  | ~\new_[371]_ ;
  assign \new_[1236]_  = ~\new_[1303]_ ;
  assign \new_[1237]_  = \new_[1359]_  | \new_[3258]_ ;
  assign \new_[1238]_  = ~\new_[1361]_  & ~\new_[1432]_ ;
  assign \new_[1239]_  = ~\new_[1362]_  & ~\new_[1432]_ ;
  assign \new_[1240]_  = ~\new_[1363]_  & ~\new_[1432]_ ;
  assign \new_[1241]_  = \new_[1365]_  | \new_[1385]_ ;
  assign \new_[1242]_  = \new_[1360]_  | \new_[1409]_ ;
  assign \new_[1243]_  = \new_[1421]_  & \new_[1356]_ ;
  assign \new_[1244]_  = \new_[1422]_  & \new_[1356]_ ;
  assign \new_[1245]_  = \new_[1423]_  & \new_[1356]_ ;
  assign \new_[1246]_  = ~\new_[3237]_  & ~\new_[1432]_ ;
  assign \new_[1247]_  = ~\new_[1364]_  & ~\new_[3233]_ ;
  assign \new_[1248]_  = ~\new_[1364]_  & ~\new_[1432]_ ;
  assign \new_[1249]_  = ~\new_[1310]_ ;
  assign \new_[1250]_  = ~\new_[3315]_  | ~\new_[3276]_  | ~\new_[1434]_ ;
  assign \new_[1251]_  = ~\new_[1401]_  | ~\new_[3276]_  | ~\new_[1453]_ ;
  assign \new_[1252]_  = ~\new_[3271]_  | ~\new_[1699]_  | ~\new_[3412]_ ;
  assign \new_[1253]_  = ~\new_[3401]_  | ~\new_[1417]_  | ~\new_[3542]_ ;
  assign \new_[1254]_  = ~\new_[1418]_  | ~\new_[1522]_  | ~\new_[1402]_ ;
  assign \new_[1255]_  = ~\new_[1374]_  & ~\new_[1399]_ ;
  assign \new_[1256]_  = ~\new_[1326]_ ;
  assign \new_[1257]_  = ~\new_[1435]_  | ~\new_[1376]_ ;
  assign \new_[1258]_  = ~\new_[1327]_ ;
  assign \new_[1259]_  = ~\new_[1442]_  | ~\new_[1481]_  | ~\new_[1768]_  | ~\new_[1386]_ ;
  assign \new_[1260]_  = ~\new_[1378]_  & ~\new_[428]_ ;
  assign \new_[1261]_  = ~\new_[1379]_  & ~\new_[429]_ ;
  assign \new_[1262]_  = ~\new_[1380]_  & ~\new_[430]_ ;
  assign \new_[1263]_  = ~\new_[1328]_ ;
  assign \new_[1264]_  = ~\new_[1329]_ ;
  assign \new_[1265]_  = ~\new_[1330]_ ;
  assign \new_[1266]_  = ~\new_[1402]_  | ~\new_[1366]_ ;
  assign \new_[1267]_  = ~\new_[1458]_  | ~\new_[1353]_ ;
  assign \new_[1268]_  = ~\new_[1349]_  | ~\new_[367]_ ;
  assign \new_[1269]_  = ~\new_[1350]_  | ~\new_[369]_ ;
  assign \new_[1270]_  = ~\new_[1351]_  | ~\new_[366]_ ;
  assign \new_[1271]_  = ~\new_[1425]_  | ~\new_[1352]_ ;
  assign \new_[1272]_  = ~\new_[1353]_  | ~\new_[1451]_ ;
  assign \new_[1273]_  = ~\new_[1354]_  & ~\new_[1461]_ ;
  assign \new_[1274]_  = ~\new_[1375]_  & ~\new_[1400]_ ;
  assign \new_[1275]_  = ~\new_[1442]_  | ~\new_[3401]_  | ~\new_[1472]_  | ~\new_[1386]_ ;
  assign \new_[1276]_  = ~\new_[1336]_ ;
  assign \new_[1277]_  = ~\new_[1337]_ ;
  assign \new_[1278]_  = ~\new_[1520]_  | ~\new_[1427]_  | ~\new_[1390]_ ;
  assign \new_[1279]_  = ~\new_[1520]_  | ~\new_[1352]_  | ~\new_[1426]_ ;
  assign \new_[1280]_  = ~\new_[1338]_ ;
  assign \new_[1281]_  = ~\new_[1442]_  | ~\new_[1482]_  | ~\new_[3412]_  | ~\new_[1386]_ ;
  assign \new_[1282]_  = ~\new_[1339]_ ;
  assign \new_[1283]_  = ~\new_[1428]_  | ~\new_[1520]_  | ~\new_[1478]_  | ~\new_[1391]_ ;
  assign \new_[1284]_  = ~\new_[1340]_ ;
  assign \new_[1285]_  = ~\new_[1341]_ ;
  assign \new_[1286]_  = ~\new_[1342]_ ;
  assign \new_[1287]_  = \new_[1414]_  | \new_[1355]_ ;
  assign \new_[1288]_  = \new_[1415]_  | \new_[1355]_ ;
  assign \new_[1289]_  = ~\new_[1361]_  & ~\new_[1392]_ ;
  assign \new_[1290]_  = ~\new_[1362]_  & ~\new_[1392]_ ;
  assign \new_[1291]_  = ~\new_[1363]_  & ~\new_[1392]_ ;
  assign \new_[1292]_  = ~\new_[1360]_  & ~\new_[3233]_ ;
  assign \new_[1293]_  = ~\new_[1383]_  & ~\new_[1365]_ ;
  assign \new_[1294]_  = ~\new_[1359]_  & ~\new_[1387]_ ;
  assign \new_[1295]_  = ~\new_[3256]_  & ~\new_[1387]_ ;
  assign \new_[1296]_  = ~\new_[3247]_  & ~\new_[1387]_ ;
  assign \new_[1297]_  = ~\new_[1361]_  & ~\new_[3233]_ ;
  assign \new_[1298]_  = ~\new_[1362]_  & ~\new_[3233]_ ;
  assign \new_[1299]_  = ~\new_[1363]_  & ~\new_[3233]_ ;
  assign \new_[1300]_  = ~\new_[1348]_ ;
  assign \new_[1301]_  = \new_[1360]_  | \new_[1432]_ ;
  assign \new_[1302]_  = \new_[1428]_  & \new_[1391]_ ;
  assign \new_[1303]_  = ~\new_[1398]_  & ~\new_[1385]_ ;
  assign \new_[1304]_  = ~\new_[1349]_ ;
  assign \new_[1305]_  = ~\new_[1350]_ ;
  assign \new_[1306]_  = ~\new_[1351]_ ;
  assign \new_[1307]_  = ~\new_[1437]_  & ~\new_[1384]_ ;
  assign \new_[1308]_  = ~\new_[1384]_  & ~\new_[1456]_ ;
  assign \new_[1309]_  = ~\new_[1457]_  & ~\new_[1384]_ ;
  assign \new_[1310]_  = ~\new_[1455]_  | ~\new_[1424]_  | ~\new_[1429]_ ;
  assign \new_[1311]_  = ~\new_[1357]_ ;
  assign \new_[1312]_  = ~\new_[1358]_ ;
  assign n826 = ~\new_[1504]_  | (~\new_[1517]_  & ~\new_[1416]_ );
  assign \new_[1314]_  = ~\new_[1395]_  & ~\new_[1699]_ ;
  assign \new_[1315]_  = ~\new_[1593]_  | ~\new_[3272]_ ;
  assign \new_[1316]_  = ~\new_[1472]_  & ~\new_[1394]_ ;
  assign \new_[1317]_  = ~\new_[1394]_  & ~\new_[1768]_ ;
  assign \new_[1318]_  = ~\new_[1396]_  & ~\new_[1593]_ ;
  assign \new_[1319]_  = ~\new_[1397]_  & ~\new_[1478]_ ;
  assign \new_[1320]_  = ~\new_[1393]_  & ~\new_[1699]_ ;
  assign \new_[1321]_  = ~\new_[1467]_  | ~\new_[1401]_ ;
  assign \new_[1322]_  = ~\new_[3237]_ ;
  assign \new_[1323]_  = ~\new_[1364]_ ;
  assign \new_[1324]_  = ~\new_[3208]_  & ~\new_[1478]_ ;
  assign \new_[1325]_  = ~\new_[1470]_  | ~\new_[1522]_  | ~\new_[1404]_ ;
  assign \new_[1326]_  = ~\new_[3401]_  | ~\new_[1435]_  | ~\new_[3313]_ ;
  assign \new_[1327]_  = ~\new_[1448]_  | ~\new_[1486]_  | ~\new_[3313]_ ;
  assign \new_[1328]_  = ~\new_[1429]_  | ~\new_[1481]_  | ~\new_[1768]_  | ~\new_[1408]_ ;
  assign \new_[1329]_  = ~\new_[1465]_  | ~\new_[1403]_ ;
  assign \new_[1330]_  = ~\new_[1466]_  | ~\new_[1403]_ ;
  assign \new_[1331]_  = \new_[1593]_  & \new_[1402]_ ;
  assign \new_[1332]_  = ~\new_[1369]_ ;
  assign \new_[1333]_  = \new_[1417]_  & \new_[3542]_ ;
  assign \new_[1334]_  = ~\new_[3542]_  | ~\new_[1430]_ ;
  assign \new_[1335]_  = \new_[3542]_  & \new_[1401]_ ;
  assign \new_[1336]_  = ~\new_[1429]_  | ~\new_[3401]_  | ~\new_[1472]_  | ~\new_[1408]_ ;
  assign \new_[1337]_  = ~\new_[1520]_  | ~\new_[3271]_  | ~\new_[1405]_ ;
  assign \new_[1338]_  = ~\new_[1431]_  | ~\new_[1482]_  | ~\new_[3412]_  | ~\new_[1412]_ ;
  assign \new_[1339]_  = ~\new_[1429]_  | ~\new_[1482]_  | ~\new_[3412]_  | ~\new_[1408]_ ;
  assign \new_[1340]_  = ~\new_[1453]_  | ~\new_[1520]_  | ~\new_[1478]_  | ~\new_[1411]_ ;
  assign \new_[1341]_  = ~\new_[1453]_  | ~\new_[1476]_  | ~\new_[1593]_  | ~\new_[1411]_ ;
  assign \new_[1342]_  = ~\new_[1453]_  | ~\new_[1477]_  | ~\new_[1699]_  | ~\new_[1411]_ ;
  assign \new_[1343]_  = ~\new_[1454]_  & ~\new_[1384]_ ;
  assign \new_[1344]_  = ~\new_[1383]_  & ~\new_[1398]_ ;
  assign \new_[1345]_  = ~\new_[1377]_ ;
  assign \new_[1346]_  = ~\new_[1446]_  & ~\new_[1384]_ ;
  assign \new_[1347]_  = ~\new_[1384]_  & ~\new_[1450]_ ;
  assign \new_[1348]_  = ~\new_[3401]_  | ~\new_[1381]_  | ~\new_[1427]_ ;
  assign \new_[1349]_  = ~\new_[1421]_  | ~\new_[1411]_ ;
  assign \new_[1350]_  = ~\new_[1422]_  | ~\new_[1411]_ ;
  assign \new_[1351]_  = ~\new_[1423]_  | ~\new_[1411]_ ;
  assign \new_[1352]_  = ~\new_[3206]_ ;
  assign \new_[1353]_  = ~\new_[1406]_  & ~\new_[1593]_ ;
  assign \new_[1354]_  = \new_[1699]_  | \new_[1406]_ ;
  assign \new_[1355]_  = ~\new_[3276]_  | ~\new_[3209]_ ;
  assign \new_[1356]_  = ~\new_[3276]_  & ~\new_[3209]_ ;
  assign \new_[1357]_  = ~\new_[1460]_  | ~\new_[3276]_  | ~\new_[1428]_ ;
  assign \new_[1358]_  = ~\new_[1431]_  | ~\new_[1424]_  | ~\new_[1425]_ ;
  assign \new_[1359]_  = ~\new_[1520]_  | ~\new_[1478]_  | ~\new_[1429]_ ;
  assign \new_[1360]_  = ~\new_[1481]_  | ~\new_[1768]_  | ~\new_[3315]_ ;
  assign \new_[1361]_  = ~\new_[1520]_  | ~\new_[1478]_  | ~\new_[1431]_ ;
  assign \new_[1362]_  = ~\new_[1431]_  | ~\new_[1593]_  | ~\new_[1476]_ ;
  assign \new_[1363]_  = ~\new_[1477]_  | ~\new_[1699]_  | ~\new_[1431]_ ;
  assign \new_[1364]_  = ~\new_[3315]_  | ~\new_[1472]_  | ~\new_[3401]_ ;
  assign \new_[1365]_  = ~\new_[3234]_  | ~\new_[3209]_ ;
  assign \new_[1366]_  = \new_[1418]_  & \new_[3401]_ ;
  assign \new_[1367]_  = \new_[1593]_  & \new_[1404]_ ;
  assign \new_[1368]_  = ~\new_[1404]_  | ~\new_[1455]_ ;
  assign \new_[1369]_  = ~\new_[1404]_  | ~\new_[1460]_ ;
  assign \new_[1370]_  = ~\new_[1520]_  | ~\new_[1404]_  | ~\new_[1458]_ ;
  assign \new_[1371]_  = ~\new_[1520]_  | ~\new_[1404]_  | ~\new_[1451]_ ;
  assign \new_[1372]_  = ~\new_[1473]_  | ~\new_[1404]_  | ~\new_[1486]_ ;
  assign \new_[1373]_  = ~\new_[1473]_  | ~\new_[1404]_  | ~\new_[1522]_ ;
  assign \new_[1374]_  = ~\new_[1768]_  | ~\new_[1412]_ ;
  assign \new_[1375]_  = ~\new_[1472]_  | ~\new_[1412]_ ;
  assign \new_[1376]_  = \new_[3313]_  & \new_[3412]_ ;
  assign \new_[1377]_  = \new_[3313]_  & \new_[1434]_ ;
  assign \new_[1378]_  = ~\new_[1413]_  & ~\new_[1407]_ ;
  assign \new_[1379]_  = ~\new_[1414]_  & ~\new_[1407]_ ;
  assign \new_[1380]_  = ~\new_[1415]_  & ~\new_[1407]_ ;
  assign \new_[1381]_  = ~\new_[1424]_  & ~\new_[1472]_ ;
  assign \new_[1382]_  = \new_[3277]_  & \new_[1459]_ ;
  assign \new_[1383]_  = ~\new_[1424]_  | ~\new_[1460]_ ;
  assign \new_[1384]_  = \new_[1406]_ ;
  assign \new_[1385]_  = ~\new_[3276]_  | ~\new_[1455]_ ;
  assign \new_[1386]_  = ~\new_[1407]_ ;
  assign \new_[1387]_  = ~\new_[1408]_ ;
  assign \new_[1388]_  = ~\new_[3273]_ ;
  assign \new_[1389]_  = ~\new_[1409]_ ;
  assign \new_[1390]_  = ~\new_[1478]_  & ~\new_[1424]_ ;
  assign \new_[1391]_  = ~\new_[1410]_ ;
  assign \new_[1392]_  = ~\new_[1412]_ ;
  assign \new_[1393]_  = ~\new_[1427]_  | ~\new_[1593]_ ;
  assign \new_[1394]_  = ~\new_[3412]_  | ~\new_[1427]_ ;
  assign \new_[1395]_  = ~\new_[1428]_  | ~\new_[1481]_ ;
  assign \new_[1396]_  = ~\new_[1428]_  | ~\new_[1482]_ ;
  assign \new_[1397]_  = ~\new_[1428]_  | ~\new_[3401]_ ;
  assign \new_[1398]_  = ~\new_[3235]_  | ~\new_[3208]_ ;
  assign \new_[1399]_  = ~\new_[1431]_  | ~\new_[1481]_ ;
  assign \new_[1400]_  = ~\new_[1431]_  | ~\new_[3401]_ ;
  assign \new_[1401]_  = \new_[1430]_  & \new_[1520]_ ;
  assign \new_[1402]_  = \new_[3543]_  & \new_[1420]_ ;
  assign \new_[1403]_  = \new_[3315]_  & \new_[1420]_ ;
  assign \new_[1404]_  = ~\new_[3209]_  & ~\new_[1433]_ ;
  assign \new_[1405]_  = ~\new_[3276]_  & ~\new_[1478]_ ;
  assign \new_[1406]_  = ~\new_[1436]_  | ~\new_[3549]_ ;
  assign \new_[1407]_  = ~\new_[3277]_  | ~\new_[3209]_ ;
  assign \new_[1408]_  = ~\new_[3276]_  & ~\new_[1459]_ ;
  assign \new_[1409]_  = ~\new_[1420]_ ;
  assign \new_[1410]_  = ~\new_[3207]_ ;
  assign \new_[1411]_  = ~\new_[3277]_  & ~\new_[3209]_ ;
  assign \new_[1412]_  = ~\new_[3545]_ ;
  assign \new_[1413]_  = ~\new_[1520]_  | ~\new_[1478]_  | ~\new_[1442]_ ;
  assign \new_[1414]_  = ~\new_[1476]_  | ~\new_[1593]_  | ~\new_[1442]_ ;
  assign \new_[1415]_  = ~\new_[1477]_  | ~\new_[1699]_  | ~\new_[1442]_ ;
  assign \new_[1416]_  = \new_[1444]_  ? \new_[1513]_  : \new_[1445]_ ;
  assign \new_[1417]_  = ~\new_[3209]_  & ~\new_[1472]_ ;
  assign \new_[1418]_  = ~\new_[3208]_  & ~\new_[1472]_ ;
  assign \new_[1419]_  = ~\new_[1432]_ ;
  assign \new_[1420]_  = ~\new_[1433]_ ;
  assign \new_[1421]_  = ~\new_[1439]_  & ~\new_[1699]_ ;
  assign \new_[1422]_  = ~\new_[1440]_  & ~\new_[1593]_ ;
  assign \new_[1423]_  = ~\new_[1441]_  & ~\new_[1478]_ ;
  assign \new_[1424]_  = ~\new_[3276]_ ;
  assign \new_[1425]_  = \new_[1443]_  & \new_[3401]_ ;
  assign \new_[1426]_  = ~\new_[3234]_  & ~\new_[1478]_ ;
  assign \new_[1427]_  = ~\new_[3548]_  & ~\new_[3314]_ ;
  assign \new_[1428]_  = \new_[1436]_ ;
  assign \new_[1429]_  = ~\new_[3235]_  & ~\new_[3209]_ ;
  assign \new_[1430]_  = ~\new_[3209]_  & ~\new_[1478]_ ;
  assign \new_[1431]_  = ~\new_[3532]_  & ~\new_[1467]_ ;
  assign \new_[1432]_  = ~\new_[3550]_  | ~\new_[3235]_ ;
  assign \new_[1433]_  = ~\new_[1447]_  | ~\new_[3538]_ ;
  assign \new_[1434]_  = \new_[1448]_  & \new_[1520]_ ;
  assign \new_[1435]_  = ~\new_[3235]_  & ~\new_[1472]_ ;
  assign \new_[1436]_  = ~\new_[3548]_  & ~\new_[3208]_ ;
  assign \new_[1437]_  = ~\new_[1451]_  | ~\new_[3401]_ ;
  assign \new_[1438]_  = ~\new_[1447]_ ;
  assign \new_[1439]_  = ~\new_[1453]_  | ~\new_[1481]_ ;
  assign \new_[1440]_  = ~\new_[1453]_  | ~\new_[1482]_ ;
  assign \new_[1441]_  = ~\new_[1453]_  | ~\new_[3401]_ ;
  assign \new_[1442]_  = ~\new_[1449]_ ;
  assign \new_[1443]_  = ~\new_[3234]_  & ~\new_[1472]_ ;
  assign \new_[1444]_  = \new_[1471]_  ? \new_[1592]_  : \new_[1463]_ ;
  assign \new_[1445]_  = \new_[1462]_  ? \new_[1592]_  : \new_[1464]_ ;
  assign \new_[1446]_  = ~\new_[1458]_  | ~\new_[3401]_ ;
  assign \new_[1447]_  = ~\new_[3546]_ ;
  assign \new_[1448]_  = ~\new_[3235]_  & ~\new_[1478]_ ;
  assign \new_[1449]_  = ~\new_[1452]_ ;
  assign \new_[1450]_  = ~\new_[1455]_ ;
  assign \new_[1451]_  = ~\new_[1467]_  & ~\new_[1472]_ ;
  assign \new_[1452]_  = ~\new_[3537]_  & ~\new_[1467]_ ;
  assign \new_[1453]_  = \new_[3537]_  & \new_[1467]_ ;
  assign \new_[1454]_  = ~\new_[1522]_  | ~\new_[1470]_ ;
  assign \new_[1455]_  = \new_[3401]_  & \new_[1470]_ ;
  assign \new_[1456]_  = ~\new_[1460]_ ;
  assign \new_[1457]_  = ~\new_[1486]_  | ~\new_[1470]_ ;
  assign \new_[1458]_  = ~\new_[3543]_  & ~\new_[3274]_ ;
  assign \new_[1459]_  = ~\new_[1467]_ ;
  assign \new_[1460]_  = \new_[1473]_  & \new_[1520]_ ;
  assign \new_[1461]_  = ~\new_[1593]_  | ~\new_[1473]_ ;
  assign \new_[1462]_  = ~\new_[1487]_  & (~\new_[1485]_  | ~\new_[1711]_ );
  assign \new_[1463]_  = ~\new_[1474]_  & (~\new_[1483]_  | ~\new_[1711]_ );
  assign \new_[1464]_  = ~\new_[1475]_  & (~\new_[1484]_  | ~\new_[1711]_ );
  assign \new_[1465]_  = \new_[1593]_  & \new_[1476]_ ;
  assign \new_[1466]_  = \new_[1699]_  & \new_[1477]_ ;
  assign \new_[1467]_  = ~\new_[3543]_ ;
  assign \new_[1468]_  = ~\new_[3445]_  | (~\new_[1497]_  & ~\new_[1489]_ );
  assign \new_[1469]_  = ~\new_[3520]_  | (~\new_[1488]_  & ~\new_[1496]_ );
  assign \new_[1470]_  = ~\new_[3543]_  & ~\new_[1472]_ ;
  assign \new_[1471]_  = \new_[1507]_  ? \new_[1711]_  : \new_[1515]_ ;
  assign \new_[1472]_  = ~\new_[3274]_ ;
  assign \new_[1473]_  = ~\new_[1467]_  & ~\new_[3274]_ ;
  assign \new_[1474]_  = ~\new_[1711]_  & (~\new_[1586]_  | ~\new_[1509]_ );
  assign \new_[1475]_  = ~\new_[1711]_  & (~\new_[1585]_  | ~\new_[1510]_ );
  assign \new_[1476]_  = ~\new_[3406]_  & ~\new_[3274]_ ;
  assign \new_[1477]_  = ~\new_[3274]_  & ~\new_[1674]_ ;
  assign \new_[1478]_  = ~\new_[1472]_ ;
  assign \new_[1479]_  = ~\new_[1486]_ ;
  assign \new_[1480]_  = \new_[3328]_  ? \new_[1514]_  : \new_[1785]_ ;
  assign \new_[1481]_  = ~\new_[1472]_  & ~\new_[3412]_ ;
  assign \new_[1482]_  = ~\new_[1768]_  & ~\new_[1472]_ ;
  assign \new_[1483]_  = ~\new_[1508]_  | (~\new_[1608]_  & ~\new_[1671]_ );
  assign \new_[1484]_  = ~\new_[1511]_  | (~\new_[1606]_  & ~\new_[1671]_ );
  assign \new_[1485]_  = ~\new_[1512]_  | (~\new_[1607]_  & ~\new_[1671]_ );
  assign \new_[1486]_  = ~\new_[1699]_  & ~\new_[3412]_ ;
  assign \new_[1487]_  = ~\new_[1516]_  & ~\new_[1711]_ ;
  assign \new_[1488]_  = ~\new_[1521]_  & (~\new_[1524]_  | ~\new_[1558]_ );
  assign \new_[1489]_  = ~\new_[3522]_  & (~\new_[1527]_  | ~\new_[1561]_ );
  assign \new_[1490]_  = ~\new_[3353]_  & (~\new_[1529]_  | ~\new_[1563]_ );
  assign \new_[1491]_  = ~\new_[3522]_  & (~\new_[1530]_  | ~\new_[1564]_ );
  assign \new_[1492]_  = ~\new_[3353]_  & (~\new_[1535]_  | ~\new_[1569]_ );
  assign \new_[1493]_  = ~\new_[1521]_  & (~\new_[1539]_  | ~\new_[1570]_ );
  assign \new_[1494]_  = ~\new_[1521]_  & (~\new_[1544]_  | ~\new_[1576]_ );
  assign \new_[1495]_  = ~\new_[3353]_  & (~\new_[1547]_  | ~\new_[1579]_ );
  assign \new_[1496]_  = ~\new_[3440]_  & (~\new_[1525]_  | ~\new_[1559]_ );
  assign \new_[1497]_  = ~\new_[3357]_  & (~\new_[1526]_  | ~\new_[1560]_ );
  assign \new_[1498]_  = ~\new_[3440]_  & (~\new_[1528]_  | ~\new_[1562]_ );
  assign \new_[1499]_  = ~\new_[3518]_  & (~\new_[1531]_  | ~\new_[1565]_ );
  assign \new_[1500]_  = ~\new_[3440]_  & (~\new_[1533]_  | ~\new_[1567]_ );
  assign \new_[1501]_  = ~\new_[3440]_  & (~\new_[1534]_  | ~\new_[1568]_ );
  assign \new_[1502]_  = ~\new_[3275]_  & (~\new_[1538]_  | ~\new_[1548]_ );
  assign \new_[1503]_  = ~\new_[3357]_  & (~\new_[1540]_  | ~\new_[1571]_ );
  assign \new_[1504]_  = ~\new_[1517]_  | ~mosi_pad_o;
  assign \new_[1505]_  = ~\new_[3440]_  & (~\new_[1545]_  | ~\new_[1577]_ );
  assign \new_[1506]_  = ~\new_[3357]_  & (~\new_[1546]_  | ~\new_[1578]_ );
  assign \new_[1507]_  = ~\new_[1588]_  & ~\new_[1518]_ ;
  assign \new_[1508]_  = ~\new_[1549]_  & (~\new_[1772]_  | ~\new_[1670]_ );
  assign \new_[1509]_  = ~\new_[1550]_  & (~\new_[1704]_  | ~\new_[1670]_ );
  assign \new_[1510]_  = ~\new_[1551]_  & (~\new_[1771]_  | ~\new_[1670]_ );
  assign \new_[1511]_  = ~\new_[1552]_  & (~\new_[1776]_  | ~\new_[1670]_ );
  assign \new_[1512]_  = ~\new_[1553]_  & (~\new_[1777]_  | ~\new_[1670]_ );
  assign \new_[1513]_  = (~\new_[1582]_  | ~\new_[2622]_ ) & (~\new_[2150]_  | ~\new_[2585]_ );
  assign \new_[1514]_  = ~\new_[1865]_  | ~\new_[1584]_  | ~\new_[1587]_ ;
  assign \new_[1515]_  = ~\new_[1555]_  & (~\new_[1664]_  | ~\new_[1670]_ );
  assign \new_[1516]_  = ~\new_[1556]_  & (~\new_[1663]_  | ~\new_[1670]_ );
  assign \new_[1517]_  = ~\new_[3145]_  & (~\new_[1591]_  | ~\new_[2223]_ );
  assign \new_[1518]_  = ~\new_[1589]_  | (~\new_[1601]_  & ~\new_[1788]_ );
  assign \new_[1519]_  = ~\new_[1522]_ ;
  assign \new_[1520]_  = \new_[1768]_  & \new_[3410]_ ;
  assign \new_[1521]_  = ~\new_[3518]_ ;
  assign \new_[1522]_  = ~\new_[1768]_  & ~\new_[1593]_ ;
  assign \new_[1523]_  = ~\new_[3411]_  | ~\new_[1622]_ ;
  assign \new_[1524]_  = ~\new_[3410]_  | ~\new_[1624]_ ;
  assign \new_[1525]_  = ~\new_[1677]_  | ~\new_[3411]_ ;
  assign \new_[1526]_  = ~\new_[3414]_  | ~\new_[1626]_ ;
  assign \new_[1527]_  = ~\new_[3410]_  | ~\new_[1679]_ ;
  assign \new_[1528]_  = ~\new_[3414]_  | ~\new_[1680]_ ;
  assign \new_[1529]_  = ~\new_[3410]_  | ~\new_[1630]_ ;
  assign \new_[1530]_  = ~\new_[3414]_  | ~\new_[1682]_ ;
  assign \new_[1531]_  = ~\new_[3411]_  | ~\new_[1633]_ ;
  assign \new_[1532]_  = ~\new_[3410]_  | ~\new_[1683]_ ;
  assign \new_[1533]_  = ~\new_[3414]_  | ~\new_[1640]_ ;
  assign \new_[1534]_  = ~\new_[3414]_  | ~\new_[1684]_ ;
  assign \new_[1535]_  = ~\new_[3411]_  | ~\new_[1643]_ ;
  assign \new_[1536]_  = ~\new_[3411]_  | ~\new_[1645]_ ;
  assign \new_[1537]_  = ~\new_[3414]_  | ~\new_[1614]_ ;
  assign \new_[1538]_  = ~\new_[3414]_  | ~\new_[1595]_ ;
  assign \new_[1539]_  = ~\new_[3414]_  | ~\new_[1649]_ ;
  assign \new_[1540]_  = ~\new_[3414]_  | ~\new_[1648]_ ;
  assign \new_[1541]_  = ~\new_[3414]_  | ~\new_[1646]_ ;
  assign \new_[1542]_  = ~\new_[3414]_  | ~\new_[1653]_ ;
  assign \new_[1543]_  = ~\new_[3414]_  | ~\new_[1655]_ ;
  assign \new_[1544]_  = ~\new_[3414]_  | ~\new_[1610]_ ;
  assign \new_[1545]_  = ~\new_[3411]_  | ~\new_[1609]_ ;
  assign \new_[1546]_  = ~\new_[3414]_  | ~\new_[1613]_ ;
  assign \new_[1547]_  = ~\new_[3410]_  | ~\new_[1660]_ ;
  assign \new_[1548]_  = ~\new_[1674]_  | ~\new_[1596]_ ;
  assign \new_[1549]_  = ~\new_[1602]_  & ~\new_[1788]_ ;
  assign \new_[1550]_  = ~\new_[1600]_  & ~\new_[1788]_ ;
  assign \new_[1551]_  = ~\new_[1603]_  & ~\new_[1788]_ ;
  assign \new_[1552]_  = ~\new_[1604]_  & ~\new_[1788]_ ;
  assign \new_[1553]_  = ~\new_[1605]_  & ~\new_[1788]_ ;
  assign sclk_pad_o = clgen_clk_out_reg;
  assign \new_[1555]_  = (~\new_[1696]_  & ~\new_[1788]_ ) | (~\new_[1702]_  & ~\new_[1671]_ );
  assign \new_[1556]_  = (~\new_[1697]_  & ~\new_[1788]_ ) | (~\new_[1706]_  & ~\new_[1671]_ );
  assign \new_[1557]_  = ~\new_[1617]_  | ~\new_[1623]_ ;
  assign \new_[1558]_  = ~\new_[1674]_  | ~\new_[1625]_ ;
  assign \new_[1559]_  = ~\new_[1617]_  | ~\new_[1678]_ ;
  assign \new_[1560]_  = ~\new_[3472]_  | ~\new_[1627]_ ;
  assign \new_[1561]_  = ~\new_[1618]_  | ~\new_[1628]_ ;
  assign \new_[1562]_  = ~\new_[1617]_  | ~\new_[1681]_ ;
  assign \new_[1563]_  = ~\new_[1674]_  | ~\new_[1631]_ ;
  assign \new_[1564]_  = ~\new_[1618]_  | ~\new_[1632]_ ;
  assign \new_[1565]_  = ~\new_[1674]_  | ~\new_[1634]_ ;
  assign \new_[1566]_  = ~\new_[1618]_  | ~\new_[1637]_ ;
  assign \new_[1567]_  = ~\new_[1619]_  | ~\new_[1641]_ ;
  assign \new_[1568]_  = ~\new_[1619]_  | ~\new_[1642]_ ;
  assign \new_[1569]_  = ~\new_[1674]_  | ~\new_[1644]_ ;
  assign \new_[1570]_  = ~\new_[1674]_  | ~\new_[1650]_ ;
  assign \new_[1571]_  = ~\new_[1674]_  | ~\new_[1651]_ ;
  assign \new_[1572]_  = ~\new_[1674]_  | ~\new_[1652]_ ;
  assign \new_[1573]_  = ~\new_[3472]_  | ~\new_[1654]_ ;
  assign \new_[1574]_  = ~\new_[1674]_  | ~\new_[1615]_ ;
  assign \new_[1575]_  = ~\new_[3472]_  | ~\new_[1611]_ ;
  assign \new_[1576]_  = ~\new_[1674]_  | ~\new_[1656]_ ;
  assign \new_[1577]_  = ~\new_[1617]_  | ~\new_[1657]_ ;
  assign \new_[1578]_  = ~\new_[3472]_  | ~\new_[1659]_ ;
  assign \new_[1579]_  = ~\new_[1621]_  | ~\new_[1618]_ ;
  assign \new_[1580]_  = \\shift_cnt_reg[7] ;
  assign \new_[1581]_  = ~\\ctrl_reg[8] ;
  assign \new_[1582]_  = \new_[2950]_  ^ \new_[1700]_ ;
  assign \new_[1583]_  = \\clgen_cnt_reg[15] ;
  assign \new_[1584]_  = ~\new_[1864]_  | ~\new_[1667]_ ;
  assign \new_[1585]_  = \new_[1705]_  | \new_[1671]_ ;
  assign \new_[1586]_  = \new_[1701]_  | \new_[1671]_ ;
  assign \new_[1587]_  = ~\new_[1864]_  | ~\new_[1857]_  | ~\new_[1757]_ ;
  assign \new_[1588]_  = ~\new_[1703]_  & ~\new_[1671]_ ;
  assign \new_[1589]_  = ~\new_[1770]_  | ~\new_[1670]_ ;
  assign \new_[1590]_  = ~\new_[1674]_  | ~\new_[1687]_ ;
  assign \new_[1591]_  = \new_[1789]_  ? \new_[1712]_  : \new_[1713]_ ;
  assign \new_[1592]_  = (~\new_[1769]_  | ~\new_[2622]_ ) & (~\new_[2262]_  | ~\new_[2585]_ );
  assign \new_[1593]_  = ~\new_[1620]_ ;
  assign n831 = sclk_pad_o ^ \new_[1766]_ ;
  assign \new_[1595]_  = ~\new_[1736]_  | ~\new_[1695]_ ;
  assign \new_[1596]_  = ~\new_[1737]_  | ~\new_[3368]_ ;
  assign \new_[1597]_  = \\shift_cnt_reg[6] ;
  assign wb_int_o = wb_int_o_reg;
  assign \wb_dat_o[9]  = \\wb_dat_o_reg[9] ;
  assign \new_[1600]_  = (~\new_[1775]_  | ~\new_[1881]_ ) & (~\new_[1833]_  | ~\new_[1966]_ );
  assign \new_[1601]_  = (~\new_[1774]_  | ~\new_[1966]_ ) & (~\new_[1834]_  | ~\new_[2044]_ );
  assign \new_[1602]_  = (~\new_[1836]_  | ~\new_[1966]_ ) & (~\new_[1885]_  | ~\new_[2044]_ );
  assign \new_[1603]_  = (~\new_[1773]_  | ~\new_[1881]_ ) & (~\new_[1884]_  | ~\new_[1966]_ );
  assign \new_[1604]_  = (~\new_[1835]_  | ~\new_[1881]_ ) & (~\new_[1886]_  | ~\new_[1966]_ );
  assign \new_[1605]_  = (~\new_[1837]_  | ~\new_[1881]_ ) & (~\new_[1887]_  | ~\new_[1966]_ );
  assign \new_[1606]_  = ~\new_[1710]_  & (~\new_[1846]_  | ~\new_[1780]_ );
  assign \new_[1607]_  = ~\new_[1708]_  & (~\new_[1846]_  | ~\new_[1782]_ );
  assign \new_[1608]_  = ~\new_[1709]_  & (~\new_[1846]_  | ~\new_[1781]_ );
  assign \new_[1609]_  = ~\new_[1824]_  | (~\new_[1831]_  & ~\new_[3186]_ );
  assign \new_[1610]_  = ~\new_[1752]_  | ~\new_[1764]_ ;
  assign \new_[1611]_  = ~\new_[1751]_  | ~\new_[1823]_ ;
  assign n836 = (~\new_[1787]_  & ~\new_[3145]_ ) | (~\new_[2557]_  & ~\new_[1658]_ );
  assign \new_[1613]_  = ~\new_[1753]_  | ~\new_[1826]_ ;
  assign \new_[1614]_  = ~\new_[1750]_  | ~\new_[1822]_ ;
  assign \new_[1615]_  = ~\new_[1749]_  | ~\new_[1763]_ ;
  assign n841 = (~\new_[1830]_  & ~\new_[2635]_ ) | (~\new_[2930]_  & ~\new_[2574]_ );
  assign \new_[1617]_  = ~\new_[3473]_ ;
  assign \new_[1618]_  = ~\new_[3473]_ ;
  assign \new_[1619]_  = ~\new_[3473]_ ;
  assign \new_[1620]_  = ~\new_[1674]_ ;
  assign \new_[1621]_  = ~\new_[1714]_  | (~\new_[1874]_  & ~\new_[3153]_ );
  assign \new_[1622]_  = ~\new_[1796]_  | (~\new_[3373]_  & ~\new_[3197]_ );
  assign \new_[1623]_  = ~\new_[1797]_  | (~\new_[1831]_  & ~\new_[3142]_ );
  assign \new_[1624]_  = ~\new_[1715]_  | ~\new_[1756]_ ;
  assign \new_[1625]_  = ~\new_[1716]_  | ~\new_[1798]_ ;
  assign \new_[1626]_  = ~\new_[1717]_  | ~\new_[1801]_ ;
  assign \new_[1627]_  = ~\new_[1718]_  | ~\new_[1802]_ ;
  assign \new_[1628]_  = ~\new_[1719]_  | (~\new_[1874]_  & ~\new_[3180]_ );
  assign \new_[1629]_  = ~\new_[1748]_  | (~\new_[1874]_  & ~\new_[3187]_ );
  assign \new_[1630]_  = ~\new_[1720]_  | (~\new_[1959]_  & ~\new_[3192]_ );
  assign \new_[1631]_  = ~\new_[1721]_  | (~\new_[1872]_  & ~\new_[3118]_ );
  assign \new_[1632]_  = ~\new_[1722]_  | (~\new_[1874]_  & ~\new_[3181]_ );
  assign \new_[1633]_  = ~\new_[1723]_  | (~\new_[1872]_  & ~\new_[3178]_ );
  assign \new_[1634]_  = ~\new_[1724]_  | (~\new_[1867]_  & ~\new_[3182]_ );
  assign \new_[1635]_  = ~\new_[1725]_  | ~\new_[1807]_ ;
  assign \new_[1636]_  = ~\new_[1726]_  | ~\new_[1808]_ ;
  assign \new_[1637]_  = ~\new_[1727]_  | (~\new_[1874]_  & ~\new_[3161]_ );
  assign \new_[1638]_  = ~\new_[1810]_  | (~\new_[3373]_  & ~\new_[3157]_ );
  assign \new_[1639]_  = ~\new_[1811]_  | (~\new_[1831]_  & ~\new_[3154]_ );
  assign \new_[1640]_  = ~\new_[1728]_  | (~\new_[1873]_  & ~\new_[3162]_ );
  assign \new_[1641]_  = ~\new_[1729]_  | (~\new_[1959]_  & ~\new_[3147]_ );
  assign \new_[1642]_  = ~\new_[1730]_  | (~\new_[1874]_  & ~\new_[3174]_ );
  assign \new_[1643]_  = ~\new_[1731]_  | (~\new_[1867]_  & ~\new_[3163]_ );
  assign \new_[1644]_  = ~\new_[1732]_  | (~\new_[1961]_  & ~\new_[3115]_ );
  assign \new_[1645]_  = ~\new_[1733]_  | (~\new_[1961]_  & ~\new_[3131]_ );
  assign \new_[1646]_  = ~\new_[1744]_  | ~\new_[1761]_ ;
  assign \new_[1647]_  = ~\new_[1741]_  | ~\new_[1813]_ ;
  assign \new_[1648]_  = ~\new_[1734]_  | ~\new_[1759]_ ;
  assign \new_[1649]_  = ~\new_[1738]_  | ~\new_[1755]_ ;
  assign \new_[1650]_  = ~\new_[1740]_  | ~\new_[1814]_ ;
  assign \new_[1651]_  = ~\new_[1742]_  | ~\new_[1760]_ ;
  assign \new_[1652]_  = ~\new_[1745]_  | ~\new_[1816]_ ;
  assign \new_[1653]_  = ~\new_[1746]_  | ~\new_[1819]_ ;
  assign \new_[1654]_  = ~\new_[1747]_  | ~\new_[1820]_ ;
  assign \new_[1655]_  = ~\new_[1735]_  | ~\new_[1762]_ ;
  assign \new_[1656]_  = ~\new_[1739]_  | ~\new_[1765]_ ;
  assign \new_[1657]_  = ~\new_[1825]_  | (~\new_[3406]_  & ~\new_[3191]_ );
  assign \new_[1658]_  = shift_tip_reg;
  assign \new_[1659]_  = ~\new_[1754]_  | ~\new_[1827]_ ;
  assign \new_[1660]_  = ~\new_[1828]_  | (~\new_[3373]_  & ~\new_[3183]_ );
  assign \wb_dat_o[11]  = \\wb_dat_o_reg[11] ;
  assign \new_[1662]_  = \\ctrl_reg[9] ;
  assign \new_[1663]_  = \new_[1894]_  ? \new_[2003]_  : \new_[1893]_ ;
  assign \new_[1664]_  = \new_[1906]_  ? \new_[2003]_  : \new_[1900]_ ;
  assign \new_[1665]_  = \\shift_cnt_reg[4] ;
  assign n846 = ~\new_[2302]_  | (~\new_[1852]_  & ~\new_[2519]_ );
  assign \new_[1667]_  = ~\new_[2037]_  | (~\new_[3417]_  & ~\new_[2036]_ );
  assign \new_[1668]_  = ~\new_[1951]_  & (~\new_[1857]_  | ~\new_[2033]_ );
  assign \new_[1669]_  = (~\new_[1858]_  | ~\new_[1857]_ ) & (~\new_[2140]_  | ~\new_[2131]_ );
  assign \new_[1670]_  = \new_[1788]_  & \new_[1966]_ ;
  assign \new_[1671]_  = ~\new_[1788]_  | ~\new_[2044]_ ;
  assign \new_[1672]_  = ~\new_[1790]_  | ~\new_[2590]_ ;
  assign n851 = (~\new_[2623]_  & ~\new_[3095]_  & ~\new_[1658]_ ) | (~\new_[3145]_  & ~\new_[2821]_  & ~\new_[1965]_ );
  assign \new_[1674]_  = \new_[3474]_ ;
  assign \new_[1675]_  = ~\new_[1791]_  | (~\new_[1873]_  & ~\new_[3128]_ );
  assign \new_[1676]_  = ~\new_[1792]_  | (~\new_[2041]_  & ~\new_[3166]_ );
  assign \new_[1677]_  = ~\new_[1793]_  | ~\new_[1799]_ ;
  assign \new_[1678]_  = ~\new_[1800]_  | (~\new_[1869]_  & ~\new_[3117]_ );
  assign \new_[1679]_  = ~\new_[1803]_  | (~\new_[1870]_  & ~\new_[3134]_ );
  assign \new_[1680]_  = ~\new_[1804]_  | (~\new_[1876]_  & ~\new_[3167]_ );
  assign \new_[1681]_  = ~\new_[1805]_  | (~\new_[1869]_  & ~\new_[3155]_ );
  assign \new_[1682]_  = ~\new_[1806]_  | (~\new_[1870]_  & ~\new_[3125]_ );
  assign \new_[1683]_  = ~\new_[1809]_  | (~\new_[1870]_  & ~\new_[3198]_ );
  assign \new_[1684]_  = ~\new_[1812]_  | (~\new_[1870]_  & ~\new_[3123]_ );
  assign \new_[1685]_  = ~\new_[1794]_  | (~\new_[1873]_  & ~\new_[3156]_ );
  assign \new_[1686]_  = ~\new_[1795]_  | (~\new_[1959]_  & ~\new_[3164]_ );
  assign \new_[1687]_  = ~\new_[1863]_  | (~\new_[1867]_  & ~\new_[3168]_ );
  assign \new_[1688]_  = ~\new_[1817]_  | (~\new_[1876]_  & ~\new_[3195]_ );
  assign \new_[1689]_  = ~\new_[1818]_  | (~\new_[1869]_  & ~\new_[3132]_ );
  assign \new_[1690]_  = \\shift_cnt_reg[5] ;
  assign \new_[1691]_  = ~\new_[1821]_  | (~\new_[1870]_  & ~\new_[3184]_ );
  assign \new_[1692]_  = \\clgen_cnt_reg[11] ;
  assign \new_[1693]_  = \\shift_cnt_reg[3] ;
  assign \new_[1694]_  = \\ctrl_reg[11] ;
  assign \new_[1695]_  = ~\new_[3406]_  | ~\new_[384]_ ;
  assign \new_[1696]_  = (~\new_[1882]_  | ~\new_[1966]_ ) & (~\new_[1883]_  | ~\new_[1881]_ );
  assign \new_[1697]_  = (~\new_[1889]_  | ~\new_[1966]_ ) & (~\new_[1888]_  | ~\new_[1881]_ );
  assign n856 = ~\new_[1832]_  | (~\new_[3171]_  & ~wb_ack_o);
  assign \new_[1699]_  = ~\new_[1768]_ ;
  assign \new_[1700]_  = ~\new_[1839]_  & ~\new_[2813]_ ;
  assign \new_[1701]_  = ~\new_[1840]_  & (~\new_[2002]_  | ~\new_[1912]_ );
  assign \new_[1702]_  = ~\new_[1844]_  & (~\new_[2003]_  | ~\new_[2012]_ );
  assign \new_[1703]_  = ~\new_[1843]_  & (~\new_[2002]_  | ~\new_[1909]_ );
  assign \new_[1704]_  = \new_[1847]_  ? \new_[2002]_  : \new_[1848]_ ;
  assign \new_[1705]_  = ~\new_[1841]_  & (~\new_[2002]_  | ~\new_[1913]_ );
  assign \new_[1706]_  = ~\new_[1842]_  & (~\new_[3381]_  | ~\new_[1898]_ );
  assign n861 = ~\new_[2698]_  | ~\new_[2780]_  | ~\new_[1838]_  | ~\new_[2773]_ ;
  assign \new_[1708]_  = ~\new_[1846]_  & ~\new_[1850]_ ;
  assign \new_[1709]_  = ~\new_[2003]_  & ~\new_[1851]_ ;
  assign \new_[1710]_  = ~\new_[2003]_  & ~\new_[1849]_ ;
  assign \new_[1711]_  = ~\new_[1855]_  & (~\new_[2378]_  | ~\new_[2106]_ );
  assign \new_[1712]_  = \\ctrl_reg[10] ;
  assign \new_[1713]_  = ~\new_[1790]_ ;
  assign \new_[1714]_  = ~\new_[1875]_  | ~\new_[486]_ ;
  assign \new_[1715]_  = ~\new_[1874]_  | ~\new_[443]_ ;
  assign \new_[1716]_  = ~\new_[1872]_  | ~\new_[441]_ ;
  assign \new_[1717]_  = ~\new_[1871]_  | ~\new_[440]_ ;
  assign \new_[1718]_  = ~\new_[1872]_  | ~\new_[562]_ ;
  assign \new_[1719]_  = ~\new_[494]_  | ~\new_[1867]_ ;
  assign \new_[1720]_  = ~\new_[3402]_  | ~\new_[559]_ ;
  assign \new_[1721]_  = ~\new_[1875]_  | ~\new_[493]_ ;
  assign \new_[1722]_  = ~\new_[1867]_  | ~\new_[442]_ ;
  assign \new_[1723]_  = ~\new_[1875]_  | ~\new_[505]_ ;
  assign \new_[1724]_  = ~\new_[1877]_  | ~\new_[557]_ ;
  assign \new_[1725]_  = ~\new_[1871]_  | ~\new_[337]_ ;
  assign \new_[1726]_  = ~\new_[1872]_  | ~\new_[335]_ ;
  assign \new_[1727]_  = ~\new_[1875]_  | ~\new_[367]_ ;
  assign \new_[1728]_  = ~\new_[1875]_  | ~\new_[341]_ ;
  assign \new_[1729]_  = ~\new_[1867]_  | ~\new_[339]_ ;
  assign \new_[1730]_  = ~\new_[1875]_  | ~\new_[359]_ ;
  assign \new_[1731]_  = ~\new_[1875]_  | ~\new_[358]_ ;
  assign \new_[1732]_  = ~\new_[1877]_  | ~\new_[328]_ ;
  assign \new_[1733]_  = ~\new_[1877]_  | ~\new_[333]_ ;
  assign \new_[1734]_  = ~\new_[1868]_  | ~\new_[348]_ ;
  assign \new_[1735]_  = ~\new_[1868]_  | ~\new_[504]_ ;
  assign \new_[1736]_  = ~\new_[1868]_  | ~\new_[345]_ ;
  assign \new_[1737]_  = ~\new_[1868]_  | ~\new_[382]_ ;
  assign \new_[1738]_  = ~\new_[1874]_  | ~\new_[381]_ ;
  assign \new_[1739]_  = ~\new_[1868]_  | ~\new_[432]_ ;
  assign \new_[1740]_  = ~\new_[1872]_  | ~\new_[352]_ ;
  assign \new_[1741]_  = ~\new_[1871]_  | ~\new_[387]_ ;
  assign \new_[1742]_  = ~\new_[1868]_  | ~\new_[386]_ ;
  assign \new_[1743]_  = ~\new_[1872]_  | ~\new_[388]_ ;
  assign \new_[1744]_  = ~\new_[1874]_  | ~\new_[389]_ ;
  assign \new_[1745]_  = ~\new_[1871]_  | ~\new_[350]_ ;
  assign \new_[1746]_  = ~\new_[1868]_  | ~\new_[379]_ ;
  assign \new_[1747]_  = ~\new_[1874]_  | ~\new_[376]_ ;
  assign \new_[1748]_  = ~\new_[1875]_  | ~\new_[383]_ ;
  assign \new_[1749]_  = ~\new_[1868]_  | ~\new_[392]_ ;
  assign \new_[1750]_  = ~\new_[1871]_  | ~\new_[394]_ ;
  assign \new_[1751]_  = ~\new_[1872]_  | ~\new_[500]_ ;
  assign \new_[1752]_  = ~\new_[1868]_  | ~\new_[434]_ ;
  assign \new_[1753]_  = ~\new_[1868]_  | ~\new_[431]_ ;
  assign \new_[1754]_  = ~\new_[1874]_  | ~\new_[429]_ ;
  assign \new_[1755]_  = ~\new_[1878]_  | ~\new_[343]_ ;
  assign \new_[1756]_  = ~\new_[1878]_  | ~\new_[446]_ ;
  assign \new_[1757]_  = ~\new_[3529]_ ;
  assign \new_[1758]_  = \new_[1866]_  | \new_[1694]_ ;
  assign \new_[1759]_  = ~\new_[1870]_  | ~\new_[347]_ ;
  assign \new_[1760]_  = ~\new_[1876]_  | ~\new_[385]_ ;
  assign \new_[1761]_  = ~\new_[1878]_  | ~\new_[351]_ ;
  assign \new_[1762]_  = ~\new_[1870]_  | ~\new_[393]_ ;
  assign \new_[1763]_  = ~\new_[1876]_  | ~\new_[503]_ ;
  assign \new_[1764]_  = ~\new_[1878]_  | ~\new_[433]_ ;
  assign \new_[1765]_  = ~\new_[1878]_  | ~\new_[325]_ ;
  assign \new_[1766]_  = ~\new_[1879]_  & ~\new_[2662]_ ;
  assign n866 = \new_[1880]_  | \new_[2761]_ ;
  assign \new_[1768]_  = ~\new_[3406]_ ;
  assign \new_[1769]_  = \new_[2732]_  ^ \new_[1968]_ ;
  assign \new_[1770]_  = \new_[1899]_  ? \new_[2025]_  : \new_[1903]_ ;
  assign \new_[1771]_  = \new_[1895]_  ? \new_[2002]_  : \new_[1902]_ ;
  assign \new_[1772]_  = \new_[1897]_  ? \new_[2002]_  : \new_[1910]_ ;
  assign \new_[1773]_  = \new_[2015]_  ? \new_[3381]_  : \new_[2019]_ ;
  assign \new_[1774]_  = \new_[2022]_  ? \new_[2003]_  : \new_[2013]_ ;
  assign \new_[1775]_  = \new_[2007]_  ? \new_[3381]_  : \new_[2020]_ ;
  assign \new_[1776]_  = \new_[1905]_  ? \new_[2025]_  : \new_[1904]_ ;
  assign \new_[1777]_  = \new_[1901]_  ? \new_[2002]_  : \new_[1896]_ ;
  assign n871 = ~\new_[2707]_  | ~\new_[2839]_  | ~\new_[1853]_  | ~\new_[2764]_ ;
  assign n876 = (~\new_[2574]_  & ~\new_[3072]_ ) | (~\new_[2279]_  & ~\new_[3331]_ );
  assign \new_[1780]_  = \new_[342]_  ? \new_[2498]_  : \new_[352]_ ;
  assign \new_[1781]_  = \new_[357]_  ? \new_[2498]_  : \new_[328]_ ;
  assign \new_[1782]_  = \new_[327]_  ? \new_[2498]_  : \new_[424]_ ;
  assign n891 = ~\new_[2299]_  | (~\new_[2021]_  & ~\new_[2519]_ );
  assign n881 = ~\new_[2359]_  | ~\new_[1920]_ ;
  assign \new_[1785]_  = ~\new_[3328]_ ;
  assign n896 = ~\new_[2358]_  | (~\new_[2027]_  & ~\new_[3145]_ );
  assign \new_[1787]_  = (~\new_[2035]_  | ~\new_[1789]_ ) & (~\new_[1580]_  | ~\new_[3137]_ );
  assign \new_[1788]_  = ~\new_[2215]_  & (~\new_[2081]_  | ~\new_[1694]_ );
  assign \new_[1789]_  = clgen_pos_edge_reg;
  assign \new_[1790]_  = ~clgen_neg_edge_reg;
  assign \new_[1791]_  = ~\new_[1960]_  | ~\new_[324]_ ;
  assign \new_[1792]_  = ~\new_[1960]_  | ~\new_[496]_ ;
  assign \new_[1793]_  = ~\new_[1959]_  | ~\new_[447]_ ;
  assign \new_[1794]_  = ~\new_[1960]_  | ~\new_[371]_ ;
  assign \new_[1795]_  = ~\new_[1960]_  | ~\new_[363]_ ;
  assign \new_[1796]_  = ~\new_[1956]_  | ~\new_[425]_ ;
  assign \new_[1797]_  = ~\new_[1954]_  | ~\new_[327]_ ;
  assign \new_[1798]_  = ~\new_[1955]_  | ~\new_[492]_ ;
  assign \new_[1799]_  = ~\new_[1954]_  | ~\new_[445]_ ;
  assign \new_[1800]_  = ~\new_[1954]_  | ~\new_[464]_ ;
  assign \new_[1801]_  = ~\new_[1955]_  | ~\new_[524]_ ;
  assign \new_[1802]_  = ~\new_[1962]_  | ~\new_[498]_ ;
  assign \new_[1803]_  = ~\new_[1954]_  | ~\new_[468]_ ;
  assign \new_[1804]_  = ~\new_[1956]_  | ~\new_[561]_ ;
  assign \new_[1805]_  = ~\new_[1954]_  | ~\new_[495]_ ;
  assign \new_[1806]_  = ~\new_[1958]_  | ~\new_[465]_ ;
  assign \new_[1807]_  = ~\new_[1955]_  | ~\new_[336]_ ;
  assign \new_[1808]_  = ~\new_[1962]_  | ~\new_[366]_ ;
  assign \new_[1809]_  = ~\new_[1958]_  | ~\new_[369]_ ;
  assign \new_[1810]_  = ~\new_[1962]_  | ~\new_[370]_ ;
  assign \new_[1811]_  = ~\new_[1954]_  | ~\new_[368]_ ;
  assign \new_[1812]_  = ~\new_[1958]_  | ~\new_[360]_ ;
  assign \new_[1813]_  = ~\new_[1955]_  | ~\new_[380]_ ;
  assign \new_[1814]_  = ~\new_[1955]_  | ~\new_[342]_ ;
  assign \new_[1815]_  = ~\new_[1962]_  | ~\new_[346]_ ;
  assign \new_[1816]_  = ~\new_[1955]_  | ~\new_[349]_ ;
  assign \new_[1817]_  = ~\new_[1956]_  | ~\new_[391]_ ;
  assign \new_[1818]_  = ~\new_[1954]_  | ~\new_[353]_ ;
  assign \new_[1819]_  = ~\new_[1962]_  | ~\new_[378]_ ;
  assign \new_[1820]_  = ~\new_[1956]_  | ~\new_[377]_ ;
  assign \new_[1821]_  = ~\new_[1958]_  | ~\new_[373]_ ;
  assign \new_[1822]_  = ~\new_[1955]_  | ~\new_[501]_ ;
  assign \new_[1823]_  = ~\new_[1962]_  | ~\new_[482]_ ;
  assign \new_[1824]_  = ~\new_[1962]_  | ~\new_[436]_ ;
  assign \new_[1825]_  = ~\new_[1954]_  | ~\new_[474]_ ;
  assign \new_[1826]_  = ~\new_[1962]_  | ~\new_[430]_ ;
  assign \new_[1827]_  = ~\new_[1956]_  | ~\new_[502]_ ;
  assign \new_[1828]_  = ~\new_[1958]_  | ~\new_[499]_ ;
  assign n886 = (~\new_[2623]_  & ~\new_[3175]_  & ~\new_[1658]_ ) | (~\new_[3145]_  & ~\new_[2816]_  & ~\new_[2151]_ );
  assign \new_[1830]_  = ~\new_[2761]_  & (~\new_[3158]_  | ~\new_[2045]_ );
  assign \new_[1831]_  = ~\new_[1867]_ ;
  assign \new_[1832]_  = ~\new_[1658]_  | ~\new_[1967]_  | ~\new_[3159]_ ;
  assign \new_[1833]_  = \new_[2114]_  ? \new_[3381]_  : \new_[2011]_ ;
  assign \new_[1834]_  = \new_[2010]_  ? \new_[3381]_  : \new_[2113]_ ;
  assign \new_[1835]_  = \new_[2018]_  ? \new_[3381]_  : \new_[2017]_ ;
  assign \new_[1836]_  = \new_[2014]_  ? \new_[3381]_  : \new_[2016]_ ;
  assign \new_[1837]_  = \new_[2008]_  ? \new_[3381]_  : \new_[2009]_ ;
  assign \new_[1838]_  = (~\new_[2832]_  | ~\new_[1950]_ ) & (~\new_[2768]_  | ~\new_[2590]_ );
  assign \new_[1839]_  = ~\new_[2190]_  | (~\new_[2006]_  & ~\new_[2850]_ );
  assign \new_[1840]_  = ~\new_[2025]_  & ~\new_[1911]_ ;
  assign \new_[1841]_  = ~\new_[2025]_  & ~\new_[1915]_ ;
  assign \new_[1842]_  = ~\new_[3381]_  & ~\new_[1914]_ ;
  assign \new_[1843]_  = ~\new_[2025]_  & ~\new_[1908]_ ;
  assign \new_[1844]_  = ~\new_[3381]_  & ~\new_[1907]_ ;
  assign n901 = (~\new_[2574]_  & ~\new_[3052]_ ) | (~\new_[2279]_  & ~\new_[2585]_ );
  assign \new_[1846]_  = ~\new_[2023]_ ;
  assign \new_[1847]_  = \new_[337]_  ? \new_[2362]_  : \new_[336]_ ;
  assign \new_[1848]_  = \new_[335]_  ? \new_[2362]_  : \new_[366]_ ;
  assign \new_[1849]_  = (~\new_[2362]_  | ~\new_[343]_ ) & (~\new_[2498]_  | ~\new_[381]_ );
  assign \new_[1850]_  = (~\new_[2362]_  | ~\new_[425]_ ) & (~\new_[2498]_  | ~\new_[426]_ );
  assign \new_[1851]_  = (~\new_[2362]_  | ~\new_[329]_ ) & (~\new_[2498]_  | ~\new_[358]_ );
  assign \new_[1852]_  = \new_[1583]_  ^ \new_[2125]_ ;
  assign \new_[1853]_  = (~\new_[2832]_  | ~\new_[1891]_ ) & (~\new_[2622]_  | ~\new_[2768]_ );
  assign \new_[1854]_  = \\clgen_cnt_reg[14] ;
  assign \new_[1855]_  = ~\new_[2077]_  | (~\new_[2380]_  & ~\new_[2622]_ );
  assign \new_[1856]_  = \\shift_cnt_reg[2] ;
  assign \new_[1857]_  = ~\new_[1924]_ ;
  assign \new_[1858]_  = ~\new_[1925]_ ;
  assign \new_[1859]_  = \\clgen_cnt_reg[13] ;
  assign \new_[1860]_  = \\ctrl_reg[0] ;
  assign \new_[1861]_  = ~\\ctrl_reg[12] ;
  assign \new_[1862]_  = ~\\ctrl_reg[13] ;
  assign \new_[1863]_  = ~\new_[2038]_  | ~\new_[362]_ ;
  assign \new_[1864]_  = ~\new_[2042]_  | ~\new_[3175]_ ;
  assign \new_[1865]_  = ~\new_[2043]_  | ~\new_[1926]_ ;
  assign \new_[1866]_  = (~\new_[2150]_  | ~\new_[3331]_ ) & (~\new_[2590]_  | ~\new_[1597]_ );
  assign \new_[1867]_  = ~\new_[1957]_ ;
  assign \new_[1868]_  = ~\new_[1958]_ ;
  assign \new_[1869]_  = ~\new_[1961]_ ;
  assign \new_[1870]_  = ~\new_[1960]_ ;
  assign \new_[1871]_  = ~\new_[1963]_ ;
  assign \new_[1872]_  = ~\new_[1963]_ ;
  assign \new_[1873]_  = ~\new_[1963]_ ;
  assign \new_[1874]_  = ~\new_[1963]_ ;
  assign \new_[1875]_  = ~\new_[1964]_ ;
  assign \new_[1876]_  = \new_[1964]_ ;
  assign \new_[1877]_  = ~\new_[3373]_ ;
  assign \new_[1878]_  = \new_[3373]_ ;
  assign \new_[1879]_  = ~\new_[2047]_  | ~\new_[1658]_ ;
  assign \new_[1880]_  = \new_[2045]_  & \new_[1658]_ ;
  assign \new_[1881]_  = ~\new_[1966]_ ;
  assign \new_[1882]_  = \new_[2108]_  ? \new_[3381]_  : \new_[2119]_ ;
  assign \new_[1883]_  = \new_[2112]_  ? \new_[3381]_  : \new_[2192]_ ;
  assign \new_[1884]_  = \new_[2116]_  ? \new_[3381]_  : \new_[2121]_ ;
  assign \new_[1885]_  = \new_[2111]_  ? \new_[3381]_  : \new_[2120]_ ;
  assign \new_[1886]_  = \new_[2115]_  ? \new_[3381]_  : \new_[2117]_ ;
  assign \new_[1887]_  = \new_[2123]_  ? \new_[3381]_  : \new_[2122]_ ;
  assign \new_[1888]_  = \new_[2118]_  ? \new_[3381]_  : \new_[2110]_ ;
  assign \new_[1889]_  = \new_[2107]_  ? \new_[3381]_  : \new_[2130]_ ;
  assign n906 = ~\new_[2005]_  | (~\new_[2574]_  & ~\new_[3034]_ );
  assign \new_[1891]_  = \\divider_reg[11] ;
  assign \new_[1892]_  = \\clgen_cnt_reg[12] ;
  assign \new_[1893]_  = \new_[392]_  ? \new_[2204]_  : \new_[503]_ ;
  assign \new_[1894]_  = \new_[504]_  ? \new_[2204]_  : \new_[393]_ ;
  assign \new_[1895]_  = \new_[354]_  ? \new_[2362]_  : \new_[391]_ ;
  assign \new_[1896]_  = \new_[496]_  ? \new_[2204]_  : \new_[427]_ ;
  assign \new_[1897]_  = \new_[331]_  ? \new_[2204]_  : \new_[360]_ ;
  assign \new_[1898]_  = \new_[500]_  ? \new_[2204]_  : \new_[482]_ ;
  assign \new_[1899]_  = \new_[440]_  ? \new_[2204]_  : \new_[524]_ ;
  assign \new_[1900]_  = \new_[557]_  ? \new_[2204]_  : \new_[506]_ ;
  assign \new_[1901]_  = \new_[324]_  ? \new_[2204]_  : \new_[497]_ ;
  assign \new_[1902]_  = \new_[390]_  ? \new_[2204]_  : \new_[353]_ ;
  assign \new_[1903]_  = \new_[498]_  ? \new_[2498]_  : \new_[562]_ ;
  assign \new_[1904]_  = \new_[344]_  ? \new_[2498]_  : \new_[382]_ ;
  assign \new_[1905]_  = \new_[384]_  ? \new_[2498]_  : \new_[345]_ ;
  assign \new_[1906]_  = \new_[558]_  ? \new_[2498]_  : \new_[505]_ ;
  assign \new_[1907]_  = (~\new_[2204]_  | ~\new_[465]_ ) & (~\new_[2498]_  | ~\new_[509]_ );
  assign \new_[1908]_  = (~\new_[2362]_  | ~\new_[468]_ ) & (~\new_[2498]_  | ~\new_[528]_ );
  assign \new_[1909]_  = \new_[439]_  ? \new_[2498]_  : \new_[494]_ ;
  assign \new_[1910]_  = \new_[330]_  ? \new_[2498]_  : \new_[359]_ ;
  assign \new_[1911]_  = (~\new_[2362]_  | ~\new_[369]_ ) & (~\new_[2498]_  | ~\new_[365]_ );
  assign \new_[1912]_  = \new_[364]_  ? \new_[2498]_  : \new_[367]_ ;
  assign \new_[1913]_  = \new_[349]_  ? \new_[2498]_  : \new_[350]_ ;
  assign \new_[1914]_  = (~\new_[2204]_  | ~\new_[501]_ ) & (~\new_[2498]_  | ~\new_[394]_ );
  assign \new_[1915]_  = (~\new_[2362]_  | ~\new_[351]_ ) & (~\new_[2498]_  | ~\new_[389]_ );
  assign \new_[1916]_  = \\divider_reg[4] ;
  assign \new_[1917]_  = \\ctrl_reg[2] ;
  assign \new_[1918]_  = \\divider_reg[15] ;
  assign \new_[1919]_  = ~\\ctrl_reg[7] ;
  assign \new_[1920]_  = ~\new_[2129]_  | ~\new_[1658]_ ;
  assign \new_[1921]_  = ~\new_[3331]_  | ~\new_[3137]_ ;
  assign \new_[1922]_  = \\clgen_cnt_reg[10] ;
  assign \new_[1923]_  = \\divider_reg[8] ;
  assign \new_[1924]_  = ~\new_[3528]_  | ~\new_[2140]_ ;
  assign \new_[1925]_  = ~\new_[2141]_  & (~\new_[2308]_  | ~\new_[3526]_ );
  assign \new_[1926]_  = \\ctrl_reg[5] ;
  assign \new_[1927]_  = \\clgen_cnt_reg[3] ;
  assign \new_[1928]_  = \\divider_reg[13] ;
  assign \new_[1929]_  = \\clgen_cnt_reg[5] ;
  assign \new_[1930]_  = \\clgen_cnt_reg[0] ;
  assign \new_[1931]_  = \\clgen_cnt_reg[2] ;
  assign \new_[1932]_  = \\clgen_cnt_reg[7] ;
  assign \new_[1933]_  = \\clgen_cnt_reg[6] ;
  assign \new_[1934]_  = \\clgen_cnt_reg[9] ;
  assign \new_[1935]_  = \\clgen_cnt_reg[1] ;
  assign \new_[1936]_  = \\ctrl_reg[1] ;
  assign \new_[1937]_  = \\divider_reg[12] ;
  assign \new_[1938]_  = \\divider_reg[10] ;
  assign \new_[1939]_  = \\divider_reg[1] ;
  assign \new_[1940]_  = \\divider_reg[2] ;
  assign \new_[1941]_  = \\ctrl_reg[3] ;
  assign \new_[1942]_  = \\ctrl_reg[4] ;
  assign \new_[1943]_  = \\ctrl_reg[6] ;
  assign \new_[1944]_  = \\divider_reg[0] ;
  assign \new_[1945]_  = \\divider_reg[14] ;
  assign \new_[1946]_  = \\divider_reg[3] ;
  assign \new_[1947]_  = \\divider_reg[5] ;
  assign \new_[1948]_  = \\divider_reg[6] ;
  assign \new_[1949]_  = \\divider_reg[7] ;
  assign \new_[1950]_  = \\divider_reg[9] ;
  assign \new_[1951]_  = ~\new_[2037]_ ;
  assign n916 = ~\new_[2149]_  & ~\new_[3145]_ ;
  assign n911 = ~\new_[2653]_  | ~\new_[2148]_ ;
  assign \new_[1954]_  = ~\new_[2038]_ ;
  assign \new_[1955]_  = ~\new_[2038]_ ;
  assign \new_[1956]_  = ~\new_[2038]_ ;
  assign \new_[1957]_  = ~\new_[2039]_ ;
  assign \new_[1958]_  = ~\new_[2039]_ ;
  assign \new_[1959]_  = ~\new_[2040]_ ;
  assign \new_[1960]_  = ~\new_[2040]_ ;
  assign \new_[1961]_  = ~\new_[2040]_ ;
  assign \new_[1962]_  = ~\new_[2041]_ ;
  assign \new_[1963]_  = ~\new_[2041]_ ;
  assign \new_[1964]_  = ~\new_[3403]_ ;
  assign \new_[1965]_  = ~\new_[2150]_  & ~\new_[3137]_ ;
  assign \new_[1966]_  = ~\new_[2044]_ ;
  assign \new_[1967]_  = ~\new_[2045]_ ;
  assign \new_[1968]_  = ~\new_[2191]_  | ~\new_[2675]_  | ~\new_[2373]_ ;
  assign \new_[1969]_  = \new_[2286]_  | \new_[2152]_ ;
  assign \new_[1970]_  = ~\new_[2094]_  | ~\new_[369]_ ;
  assign \new_[1971]_  = ~\new_[2094]_  | ~\new_[357]_ ;
  assign \new_[1972]_  = ~\new_[2094]_  | ~\new_[328]_ ;
  assign \new_[1973]_  = ~\new_[2094]_  | ~\new_[358]_ ;
  assign \new_[1974]_  = ~\new_[2096]_  | ~\new_[359]_ ;
  assign \new_[1975]_  = ~\new_[2094]_  | ~\new_[360]_ ;
  assign \new_[1976]_  = ~\new_[2094]_  | ~\new_[331]_ ;
  assign \new_[1977]_  = ~\new_[2094]_  | ~\new_[361]_ ;
  assign \new_[1978]_  = ~\new_[2095]_  | ~\new_[362]_ ;
  assign \new_[1979]_  = ~\new_[2095]_  | ~\new_[332]_ ;
  assign \new_[1980]_  = ~\new_[2095]_  | ~\new_[333]_ ;
  assign \new_[1981]_  = ~\new_[2095]_  | ~\new_[334]_ ;
  assign \new_[1982]_  = ~\new_[2095]_  | ~\new_[329]_ ;
  assign \new_[1983]_  = ~\new_[2095]_  | ~\new_[372]_ ;
  assign \new_[1984]_  = ~\new_[2095]_  | ~\new_[371]_ ;
  assign \new_[1985]_  = ~\new_[2244]_  | ~\new_[364]_ ;
  assign \new_[1986]_  = ~\new_[2096]_  | ~\new_[367]_ ;
  assign \new_[1987]_  = ~\new_[2096]_  | ~\new_[368]_ ;
  assign \new_[1988]_  = ~\new_[2096]_  | ~\new_[365]_ ;
  assign \new_[1989]_  = ~\new_[2244]_  | ~\new_[366]_ ;
  assign \new_[1990]_  = ~\new_[2096]_  | ~\new_[335]_ ;
  assign \new_[1991]_  = ~\new_[2244]_  | ~\new_[337]_ ;
  assign \new_[1992]_  = ~\new_[2244]_  | ~\new_[330]_ ;
  assign \new_[1993]_  = ~\new_[2244]_  | ~\new_[356]_ ;
  assign \new_[1994]_  = ~\new_[2244]_  | ~\new_[370]_ ;
  assign \new_[1995]_  = ~\new_[2095]_  | ~\new_[338]_ ;
  assign \new_[1996]_  = ~\new_[2244]_  | ~\new_[355]_ ;
  assign \new_[1997]_  = ~\new_[2244]_  | ~\new_[339]_ ;
  assign \new_[1998]_  = ~\new_[2094]_  | ~\new_[341]_ ;
  assign \new_[1999]_  = ~\new_[2096]_  | ~\new_[363]_ ;
  assign \new_[2000]_  = ~\new_[2096]_  | ~\new_[340]_ ;
  assign \new_[2001]_  = ~\new_[2096]_  | ~\new_[336]_ ;
  assign \new_[2002]_  = ~\new_[2023]_ ;
  assign \new_[2003]_  = ~\new_[2023]_ ;
  assign \new_[2004]_  = \\clgen_cnt_reg[4] ;
  assign \new_[2005]_  = ~\new_[2193]_  | ~\new_[1712]_ ;
  assign \new_[2006]_  = \new_[2200]_  & \new_[2675]_ ;
  assign \new_[2007]_  = \new_[338]_  ? \new_[2362]_  : \new_[370]_ ;
  assign \new_[2008]_  = \new_[428]_  ? \new_[2362]_  : \new_[499]_ ;
  assign \new_[2009]_  = \new_[486]_  ? \new_[2362]_  : \new_[488]_ ;
  assign \new_[2010]_  = \new_[446]_  ? \new_[2498]_  : \new_[443]_ ;
  assign \new_[2011]_  = \new_[355]_  ? \new_[2498]_  : \new_[339]_ ;
  assign \new_[2012]_  = \new_[508]_  ? \new_[2498]_  : \new_[442]_ ;
  assign \new_[2013]_  = \new_[464]_  ? \new_[2498]_  : \new_[444]_ ;
  assign \new_[2014]_  = \new_[372]_  ? \new_[2498]_  : \new_[371]_ ;
  assign \new_[2015]_  = \new_[373]_  ? \new_[2498]_  : \new_[374]_ ;
  assign \new_[2016]_  = \new_[334]_  ? \new_[2498]_  : \new_[363]_ ;
  assign \new_[2017]_  = \new_[346]_  ? \new_[2498]_  : \new_[388]_ ;
  assign \new_[2018]_  = \new_[380]_  ? \new_[2498]_  : \new_[387]_ ;
  assign \new_[2019]_  = \new_[375]_  ? \new_[2498]_  : \new_[383]_ ;
  assign \new_[2020]_  = \new_[368]_  ? \new_[2498]_  : \new_[356]_ ;
  assign \new_[2021]_  = ~\new_[2205]_  & (~\new_[2491]_  | ~\new_[1692]_ );
  assign \new_[2022]_  = \new_[445]_  ? \new_[2498]_  : \new_[447]_ ;
  assign \new_[2023]_  = ~\new_[3381]_ ;
  assign n921 = ~\new_[2301]_  | (~\new_[2292]_  & ~\new_[2519]_ );
  assign \new_[2025]_  = \new_[3381]_ ;
  assign \new_[2026]_  = ~\new_[3526]_  | ~\new_[2396]_  | ~\new_[2309]_ ;
  assign \new_[2027]_  = ~\new_[2214]_  | (~\new_[3061]_  & ~\new_[1789]_ );
  assign n931 = ~\new_[2300]_  | (~\new_[2293]_  & ~\new_[2519]_ );
  assign \new_[2029]_  = \\shift_cnt_reg[1] ;
  assign \wb_dat_o[7]  = \\wb_dat_o_reg[7] ;
  assign \wb_dat_o[3]  = \\wb_dat_o_reg[3] ;
  assign \new_[2032]_  = \\shift_cnt_reg[0] ;
  assign \new_[2033]_  = \new_[3511]_  & \new_[3526]_ ;
  assign n926 = (~\new_[2623]_  & ~\new_[3140]_  & ~\new_[1658]_ ) | (~\new_[3145]_  & ~\new_[2644]_  & ~\new_[2387]_ );
  assign \new_[2035]_  = ~\new_[2216]_  | (~\new_[2384]_  & ~\new_[1580]_ );
  assign \new_[2036]_  = ~\new_[2140]_ ;
  assign \new_[2037]_  = ~\new_[2219]_  | ~\new_[1942]_ ;
  assign \new_[2038]_  = ~\new_[3374]_ ;
  assign \new_[2039]_  = ~\new_[3374]_ ;
  assign \new_[2040]_  = \new_[3374]_ ;
  assign \new_[2041]_  = ~\new_[3374]_ ;
  assign \new_[2042]_  = ~\new_[2652]_  | ~\new_[2217]_ ;
  assign \new_[2043]_  = \new_[2652]_  & \new_[2217]_ ;
  assign \new_[2044]_  = ~\new_[2388]_  & (~\new_[2263]_  | ~\new_[2622]_ );
  assign \new_[2045]_  = \new_[2223]_  | \new_[3137]_ ;
  assign \new_[2046]_  = ~\new_[2222]_  | ~\new_[446]_ ;
  assign \new_[2047]_  = \new_[2223]_  | sclk_pad_o;
  assign \new_[2048]_  = ~\new_[2222]_  | ~\new_[509]_ ;
  assign \new_[2049]_  = ~\new_[2222]_  | ~\new_[506]_ ;
  assign \new_[2050]_  = ~\new_[2222]_  | ~\new_[558]_ ;
  assign \new_[2051]_  = ~\new_[2222]_  | ~\new_[505]_ ;
  assign \new_[2052]_  = ~\new_[2222]_  | ~\new_[437]_ ;
  assign \new_[2053]_  = ~\new_[2222]_  | ~\new_[493]_ ;
  assign \new_[2054]_  = ~\new_[2222]_  | ~\new_[507]_ ;
  assign \new_[2055]_  = ~\new_[2222]_  | ~\new_[559]_ ;
  assign \new_[2056]_  = ~\new_[2222]_  | ~\new_[495]_ ;
  assign \new_[2057]_  = ~\new_[2222]_  | ~\new_[438]_ ;
  assign \new_[2058]_  = ~\new_[2222]_  | ~\new_[439]_ ;
  assign \new_[2059]_  = ~\new_[2222]_  | ~\new_[494]_ ;
  assign \new_[2060]_  = ~\new_[2222]_  | ~\new_[468]_ ;
  assign \new_[2061]_  = ~\new_[2222]_  | ~\new_[528]_ ;
  assign \new_[2062]_  = ~\new_[2222]_  | ~\new_[445]_ ;
  assign \new_[2063]_  = ~\new_[2222]_  | ~\new_[562]_ ;
  assign \new_[2064]_  = ~\new_[2222]_  | ~\new_[524]_ ;
  assign \new_[2065]_  = ~\new_[2222]_  | ~\new_[440]_ ;
  assign \new_[2066]_  = ~\new_[2222]_  | ~\new_[492]_ ;
  assign \new_[2067]_  = ~\new_[2222]_  | ~\new_[508]_ ;
  assign \new_[2068]_  = ~\new_[2222]_  | ~\new_[498]_ ;
  assign \new_[2069]_  = ~\new_[2222]_  | ~\new_[442]_ ;
  assign \new_[2070]_  = ~\new_[2222]_  | ~\new_[441]_ ;
  assign \new_[2071]_  = ~\new_[2222]_  | ~\new_[465]_ ;
  assign \new_[2072]_  = ~\new_[2222]_  | ~\new_[443]_ ;
  assign \new_[2073]_  = ~\new_[2222]_  | ~\new_[464]_ ;
  assign \new_[2074]_  = ~\new_[2222]_  | ~\new_[444]_ ;
  assign \new_[2075]_  = ~\new_[2222]_  | ~\new_[447]_ ;
  assign \new_[2076]_  = \\clgen_cnt_reg[8] ;
  assign \new_[2077]_  = ~\new_[2622]_  | ~\new_[2189]_  | ~\new_[2587]_ ;
  assign n936 = ~\new_[2185]_  | (~\new_[2740]_  & ~\new_[2574]_ );
  assign n946 = (~\new_[2574]_  & ~\new_[3031]_ ) | (~\new_[2279]_  & ~\new_[1862]_ );
  assign n941 = (~\new_[2574]_  & ~\new_[3060]_ ) | (~\new_[2279]_  & ~\new_[1861]_ );
  assign \new_[2081]_  = \new_[2640]_  ^ \new_[2280]_ ;
  assign \new_[2082]_  = ~\new_[2282]_  | ~\new_[373]_ ;
  assign \new_[2083]_  = ~\new_[2282]_  | ~\new_[374]_ ;
  assign \new_[2084]_  = ~\new_[2282]_  | ~\new_[377]_ ;
  assign \new_[2085]_  = ~\new_[2282]_  | ~\new_[378]_ ;
  assign \new_[2086]_  = ~\new_[2282]_  | ~\new_[379]_ ;
  assign \new_[2087]_  = ~\new_[2276]_  | ~\new_[393]_ ;
  assign \new_[2088]_  = ~\new_[2282]_  | ~\new_[388]_ ;
  assign \new_[2089]_  = ~\new_[2282]_  | ~\new_[351]_ ;
  assign \new_[2090]_  = ~\new_[2282]_  | ~\new_[381]_ ;
  assign \new_[2091]_  = ~\new_[2282]_  | ~\new_[350]_ ;
  assign \new_[2092]_  = ~\new_[2276]_  | ~\new_[394]_ ;
  assign \new_[2093]_  = ~\new_[2276]_  | ~\new_[392]_ ;
  assign \new_[2094]_  = ~\new_[2179]_ ;
  assign \new_[2095]_  = ~\new_[2179]_ ;
  assign \new_[2096]_  = ~\new_[2179]_ ;
  assign \new_[2097]_  = ~\new_[3500]_ ;
  assign \new_[2098]_  = ~\new_[3500]_ ;
  assign \new_[2099]_  = ~\new_[2282]_  | ~\new_[389]_ ;
  assign \new_[2100]_  = ~\new_[2282]_  | ~\new_[384]_ ;
  assign \new_[2101]_  = ~\new_[2282]_  | ~\new_[353]_ ;
  assign \new_[2102]_  = ~\new_[2282]_  | ~\new_[387]_ ;
  assign \new_[2103]_  = ~\new_[2282]_  | ~\new_[345]_ ;
  assign \new_[2104]_  = ~\new_[2282]_  | ~\new_[347]_ ;
  assign \new_[2105]_  = ~\new_[2282]_  | ~\new_[391]_ ;
  assign \new_[2106]_  = ~\new_[2189]_ ;
  assign \new_[2107]_  = \new_[326]_  ? \new_[2204]_  : \new_[436]_ ;
  assign \new_[2108]_  = \new_[438]_  ? \new_[2362]_  : \new_[561]_ ;
  assign \new_[2109]_  = ~\\ss_reg[5] ;
  assign \new_[2110]_  = \new_[432]_  ? \new_[2362]_  : \new_[325]_ ;
  assign \new_[2111]_  = \new_[333]_  ? \new_[2204]_  : \new_[332]_ ;
  assign \new_[2112]_  = \new_[559]_  ? \new_[2362]_  : \new_[507]_ ;
  assign \new_[2113]_  = \new_[441]_  ? \new_[2204]_  : \new_[492]_ ;
  assign \new_[2114]_  = \new_[341]_  ? \new_[2204]_  : \new_[340]_ ;
  assign \new_[2115]_  = \new_[348]_  ? \new_[2362]_  : \new_[347]_ ;
  assign \new_[2116]_  = \new_[379]_  ? \new_[2204]_  : \new_[378]_ ;
  assign \new_[2117]_  = \new_[386]_  ? \new_[2362]_  : \new_[385]_ ;
  assign \new_[2118]_  = \new_[434]_  ? \new_[2204]_  : \new_[433]_ ;
  assign \new_[2119]_  = \new_[495]_  ? \new_[2498]_  : \new_[560]_ ;
  assign \new_[2120]_  = \new_[361]_  ? \new_[2498]_  : \new_[362]_ ;
  assign \new_[2121]_  = \new_[377]_  ? \new_[2498]_  : \new_[376]_ ;
  assign \new_[2122]_  = \new_[502]_  ? \new_[2498]_  : \new_[429]_ ;
  assign \new_[2123]_  = \new_[430]_  ? \new_[2498]_  : \new_[431]_ ;
  assign \new_[2124]_  = ~\\ss_reg[3] ;
  assign \new_[2125]_  = \new_[1859]_  | \new_[1854]_  | \new_[2285]_  | \new_[1892]_ ;
  assign \new_[2126]_  = ~\\ss_reg[1] ;
  assign n1021 = ~\new_[2296]_  | (~\new_[2495]_  & ~\new_[2519]_ );
  assign n956 = \new_[2379]_  ? \new_[2519]_  : \new_[1937]_ ;
  assign \new_[2129]_  = ~\new_[2642]_  & (~\new_[2380]_  | ~\new_[1789]_ );
  assign \new_[2130]_  = \new_[435]_  ? \new_[2362]_  : \new_[474]_ ;
  assign \new_[2131]_  = ~\new_[2210]_ ;
  assign n996 = ~\new_[2305]_  | (~\new_[2748]_  & ~\new_[2519]_ );
  assign \new_[2133]_  = ~\new_[2643]_  | (~\new_[2385]_  & ~\new_[3436]_ );
  assign n981 = \new_[2383]_  ? \new_[2519]_  : \new_[1938]_ ;
  assign \new_[2135]_  = ~\\ss_reg[7] ;
  assign \new_[2136]_  = ~\\ss_reg[0] ;
  assign \new_[2137]_  = ~\\ss_reg[2] ;
  assign \new_[2138]_  = ~\\ss_reg[4] ;
  assign \new_[2139]_  = ~\\ss_reg[6] ;
  assign \new_[2140]_  = ~\new_[2307]_  | ~\new_[3190]_ ;
  assign \new_[2141]_  = ~\new_[3408]_ ;
  assign n1006 = ~\new_[2294]_  | (~\new_[2687]_  & ~\new_[2519]_ );
  assign n1026 = ~\new_[2295]_  | (~\new_[2744]_  & ~\new_[2519]_ );
  assign n1011 = ~\new_[2298]_  | (~\new_[2519]_  & ~\new_[1930]_ );
  assign n1031 = ~\new_[2297]_  | (~\new_[2660]_  & ~\new_[2519]_ );
  assign n1016 = ~\new_[2304]_  | (~\new_[2785]_  & ~\new_[2519]_ );
  assign n1036 = ~\new_[2303]_  | (~\new_[2914]_  & ~\new_[2519]_ );
  assign \new_[2148]_  = (~\new_[2737]_  | ~\new_[2419]_ ) & (~\new_[2690]_  | ~sclk_pad_o);
  assign \new_[2149]_  = (~\new_[2419]_  | ~sclk_pad_o) & (~\new_[2690]_  | ~\new_[3121]_ );
  assign \new_[2150]_  = \new_[1597]_  ^ \new_[2357]_ ;
  assign \new_[2151]_  = ~\new_[2262]_  & ~\new_[3137]_ ;
  assign \new_[2152]_  = \new_[2262]_  & \new_[3331]_ ;
  assign n961 = ~\new_[2245]_  | (~\new_[2680]_  & ~\new_[3102]_ );
  assign n1051 = ~\new_[2253]_  | (~\new_[2680]_  & ~\new_[3034]_ );
  assign n976 = (~\new_[2574]_  & ~\new_[3097]_ ) | (~\new_[2371]_  & ~\new_[1919]_ );
  assign n1001 = ~\new_[2237]_  | (~\new_[2680]_  & ~\new_[3031]_ );
  assign n1096 = ~\new_[2257]_  | (~\new_[2680]_  & ~\new_[3098]_ );
  assign n1061 = ~\new_[2254]_  | (~\new_[2680]_  & ~\new_[3073]_ );
  assign n1086 = ~\new_[2252]_  | (~\new_[2680]_  & ~\new_[3056]_ );
  assign n1041 = (~\new_[2574]_  & ~\new_[3075]_ ) | (~\new_[2371]_  & ~\new_[3319]_ );
  assign n966 = (~\new_[2574]_  & ~\new_[3073]_ ) | (~\new_[2371]_  & ~\new_[3140]_ );
  assign n1066 = (~\new_[2574]_  & ~\new_[3094]_ ) | (~\new_[2371]_  & ~\new_[3124]_ );
  assign n1071 = (~\new_[2574]_  & ~\new_[3102]_ ) | (~\new_[2371]_  & ~\new_[3190]_ );
  assign n991 = (~\new_[2574]_  & ~\new_[3098]_ ) | (~\new_[2371]_  & ~\new_[3175]_ );
  assign n1076 = (~\new_[2574]_  & ~\new_[3107]_ ) | (~\new_[2371]_  & ~\new_[3095]_ );
  assign n1081 = ~\new_[2251]_  | (~\new_[2680]_  & ~\new_[3051]_ );
  assign n951 = ~\new_[2284]_  | (~\new_[2680]_  & ~\new_[3052]_ );
  assign n1046 = ~\new_[2247]_  | (~\new_[2680]_  & ~\new_[3060]_ );
  assign n971 = ~\new_[2255]_  | (~\new_[2680]_  & ~\new_[3090]_ );
  assign n986 = ~\new_[2260]_  | (~\new_[2680]_  & ~\new_[3054]_ );
  assign n1056 = ~\new_[2250]_  | (~\new_[2680]_  & ~\new_[3075]_ );
  assign n1101 = ~\new_[2258]_  | (~\new_[2680]_  & ~\new_[3107]_ );
  assign n1091 = ~\new_[2256]_  | (~\new_[2680]_  & ~\new_[3094]_ );
  assign n1106 = ~\new_[2259]_  | (~\new_[2680]_  & ~\new_[3097]_ );
  assign n1111 = ~\new_[2261]_  | (~\new_[2680]_  & ~\new_[3072]_ );
  assign \wb_dat_o[4]  = \\wb_dat_o_reg[4] ;
  assign \new_[2177]_  = ~\new_[2377]_  | ~\new_[383]_ ;
  assign \new_[2178]_  = ~\new_[2377]_  | ~\new_[386]_ ;
  assign \new_[2179]_  = ~\new_[2244]_ ;
  assign \new_[2180]_  = ~\new_[2244]_ ;
  assign \new_[2181]_  = \new_[3310]_ ;
  assign \new_[2182]_  = ~\new_[3500]_ ;
  assign \new_[2183]_  = ~\new_[3500]_ ;
  assign \new_[2184]_  = ~\new_[2377]_  | ~\new_[382]_ ;
  assign \new_[2185]_  = \new_[2371]_  | \new_[3122]_ ;
  assign \new_[2186]_  = ~\new_[2377]_  | ~\new_[390]_ ;
  assign \new_[2187]_  = ~\new_[2377]_  | ~\new_[376]_ ;
  assign \new_[2188]_  = ~\new_[2377]_  | ~\new_[375]_ ;
  assign \new_[2189]_  = ~\new_[2386]_  | (~\new_[2638]_  & ~\new_[2573]_ );
  assign \new_[2190]_  = \new_[2671]_  | \new_[2573]_  | \new_[2850]_  | \new_[2638]_ ;
  assign \new_[2191]_  = ~\new_[2581]_  & (~\new_[2489]_  | ~\new_[2582]_ );
  assign \new_[2192]_  = \new_[437]_  ? \new_[2498]_  : \new_[493]_ ;
  assign \new_[2193]_  = ~\new_[2279]_ ;
  assign \new_[2194]_  = ~\new_[2597]_  | ~\new_[3176]_ ;
  assign \new_[2195]_  = ~\new_[2389]_  | ~\new_[3113]_ ;
  assign \new_[2196]_  = ~\new_[2389]_  | ~\new_[3084]_ ;
  assign \new_[2197]_  = ~\new_[2389]_  | ~\new_[3146]_ ;
  assign \new_[2198]_  = ~\new_[2389]_  | ~\new_[3195]_ ;
  assign \new_[2199]_  = ~\new_[2597]_  | ~\new_[3139]_ ;
  assign \new_[2200]_  = \new_[2386]_  | \new_[2671]_ ;
  assign \new_[2201]_  = ~\new_[2597]_  | ~\new_[3138]_ ;
  assign \new_[2202]_  = ~\new_[2597]_  | ~\new_[3199]_ ;
  assign \wb_dat_o[5]  = \\wb_dat_o_reg[5] ;
  assign \new_[2204]_  = ~\new_[2498]_ ;
  assign \new_[2205]_  = ~\new_[2285]_ ;
  assign \wb_dat_o[0]  = \\wb_dat_o_reg[0] ;
  assign n1141 = \new_[2586]_  ? \new_[2519]_  : \new_[1923]_ ;
  assign n1116 = \new_[2679]_  ? \new_[2519]_  : \new_[1916]_ ;
  assign \new_[2209]_  = ~\new_[2380]_  & ~\new_[2590]_ ;
  assign \new_[2210]_  = ~\new_[2381]_  | ~\new_[1941]_ ;
  assign \wb_dat_o[1]  = \\wb_dat_o_reg[1] ;
  assign \wb_dat_o[6]  = \\wb_dat_o_reg[6] ;
  assign \wb_dat_o[2]  = \\wb_dat_o_reg[2] ;
  assign \new_[2214]_  = ~\new_[2385]_  | ~\new_[1789]_ ;
  assign \new_[2215]_  = ~\new_[2385]_  & ~\new_[1694]_ ;
  assign \new_[2216]_  = ~\new_[2384]_  | ~\new_[1580]_ ;
  assign \new_[2217]_  = ~\new_[2395]_  | ~\new_[3436]_ ;
  assign n1121 = (~\new_[2623]_  & ~\new_[3319]_  & ~\new_[1658]_ ) | (~\new_[3145]_  & ~\new_[2741]_  & ~\new_[2552]_ );
  assign \new_[2219]_  = ~\new_[2307]_ ;
  assign n1131 = ~\new_[2567]_  | ~\new_[2633]_  | ~\new_[2695]_  | ~\new_[2838]_ ;
  assign n1126 = ~\new_[2566]_  | ~\new_[2631]_  | ~\new_[2688]_  | ~\new_[2791]_ ;
  assign \new_[2222]_  = \new_[3365]_  | \new_[3500]_ ;
  assign \new_[2223]_  = ~\new_[3074]_  | ~\new_[2361]_  | ~\new_[3032]_ ;
  assign n1136 = ~\new_[2599]_  | ~\new_[2356]_ ;
  assign \new_[2225]_  = \new_[2374]_  & \new_[376]_ ;
  assign \new_[2226]_  = \new_[2374]_  & \new_[378]_ ;
  assign \new_[2227]_  = \new_[2374]_  & \new_[379]_ ;
  assign \new_[2228]_  = \new_[3292]_  & \new_[351]_ ;
  assign \new_[2229]_  = \new_[3292]_  & \new_[345]_ ;
  assign \new_[2230]_  = \new_[2374]_  & \new_[347]_ ;
  assign \new_[2231]_  = \new_[3292]_  & \new_[350]_ ;
  assign \new_[2232]_  = \new_[2374]_  & \new_[353]_ ;
  assign \new_[2233]_  = \new_[2929]_  | \new_[2483]_ ;
  assign \new_[2234]_  = \new_[2876]_  | \new_[2483]_ ;
  assign \new_[2235]_  = \new_[2909]_  | \new_[2483]_ ;
  assign \new_[2236]_  = \new_[2890]_  | \new_[2483]_ ;
  assign \new_[2237]_  = ~\new_[2484]_  | ~\new_[1928]_ ;
  assign \new_[2238]_  = ~\new_[3308]_  | ~\new_[327]_ ;
  assign \new_[2239]_  = ~\new_[3308]_  | ~\new_[324]_ ;
  assign \new_[2240]_  = ~\new_[2363]_ ;
  assign \new_[2241]_  = ~\new_[2363]_ ;
  assign \new_[2242]_  = ~\new_[2363]_ ;
  assign \new_[2243]_  = ~\new_[3308]_  | ~\new_[325]_ ;
  assign \new_[2244]_  = \new_[3500]_ ;
  assign \new_[2245]_  = ~\new_[2478]_  | ~\new_[1916]_ ;
  assign \new_[2246]_  = ~\new_[3308]_  | ~\new_[326]_ ;
  assign \new_[2247]_  = ~\new_[2484]_  | ~\new_[1937]_ ;
  assign \wb_dat_o[10]  = \\wb_dat_o_reg[10] ;
  assign \new_[2249]_  = ~\new_[2372]_ ;
  assign \new_[2250]_  = ~\new_[2478]_  | ~\new_[1939]_ ;
  assign \new_[2251]_  = ~\new_[2478]_  | ~\new_[1944]_ ;
  assign \new_[2252]_  = ~\new_[2484]_  | ~\new_[1945]_ ;
  assign \new_[2253]_  = ~\new_[2484]_  | ~\new_[1938]_ ;
  assign \new_[2254]_  = ~\new_[2478]_  | ~\new_[1940]_ ;
  assign \new_[2255]_  = ~\new_[2484]_  | ~\new_[1918]_ ;
  assign \new_[2256]_  = ~\new_[2478]_  | ~\new_[1946]_ ;
  assign \new_[2257]_  = ~\new_[2478]_  | ~\new_[1947]_ ;
  assign \new_[2258]_  = ~\new_[2478]_  | ~\new_[1948]_ ;
  assign \new_[2259]_  = ~\new_[2478]_  | ~\new_[1949]_ ;
  assign \new_[2260]_  = ~\new_[2484]_  | ~\new_[1923]_ ;
  assign \new_[2261]_  = ~\new_[2484]_  | ~\new_[1950]_ ;
  assign \new_[2262]_  = \new_[3074]_  ^ \new_[2572]_ ;
  assign \new_[2263]_  = \new_[2580]_  ^ \new_[2573]_ ;
  assign \new_[2264]_  = ~\new_[2515]_  & ~\new_[3147]_ ;
  assign \new_[2265]_  = ~\new_[2515]_  & ~\new_[3115]_ ;
  assign \new_[2266]_  = ~\new_[2515]_  & ~\new_[3163]_ ;
  assign \new_[2267]_  = ~\new_[2515]_  & ~\new_[3174]_ ;
  assign \new_[2268]_  = ~\new_[2637]_  & ~\new_[3123]_ ;
  assign \new_[2269]_  = ~\new_[2487]_  & ~\new_[3168]_ ;
  assign \new_[2270]_  = ~\new_[2487]_  & ~\new_[3131]_ ;
  assign \new_[2271]_  = ~\new_[2488]_  & ~\new_[3164]_ ;
  assign \new_[2272]_  = ~\new_[2637]_  & ~\new_[3156]_ ;
  assign \new_[2273]_  = ~\new_[2488]_  & ~\new_[3161]_ ;
  assign \new_[2274]_  = ~\new_[2487]_  & ~\new_[3198]_ ;
  assign \new_[2275]_  = ~\new_[2487]_  & ~\new_[3154]_ ;
  assign \new_[2276]_  = ~\new_[3298]_ ;
  assign \new_[2277]_  = ~\new_[2637]_  & ~\new_[3162]_ ;
  assign \new_[2278]_  = ~\new_[2637]_  & ~\new_[3157]_ ;
  assign \new_[2279]_  = \new_[2635]_  & \wb_sel_i[1] ;
  assign \new_[2280]_  = \new_[2575]_  | \new_[2489]_ ;
  assign \new_[2281]_  = ~\new_[3349]_ ;
  assign \new_[2282]_  = ~\new_[2372]_ ;
  assign \new_[2283]_  = ~\new_[3219]_ ;
  assign \new_[2284]_  = ~\new_[2484]_  | ~\new_[1891]_ ;
  assign \new_[2285]_  = \new_[2491]_  | \new_[1692]_ ;
  assign \new_[2286]_  = ~\new_[3331]_  & ~\new_[3074]_ ;
  assign \wb_dat_o[13]  = \\wb_dat_o_reg[13] ;
  assign \wb_dat_o[14]  = \\wb_dat_o_reg[14] ;
  assign \wb_dat_o[12]  = \\wb_dat_o_reg[12] ;
  assign \wb_dat_o[8]  = \\wb_dat_o_reg[8] ;
  assign \wb_dat_o[15]  = \\wb_dat_o_reg[15] ;
  assign \new_[2292]_  = \new_[1854]_  ^ \new_[2593]_ ;
  assign \new_[2293]_  = \new_[1859]_  ^ \new_[2595]_ ;
  assign \new_[2294]_  = ~\new_[2519]_  | ~\new_[1947]_ ;
  assign \new_[2295]_  = ~\new_[2519]_  | ~\new_[1948]_ ;
  assign \new_[2296]_  = ~\new_[2519]_  | ~\new_[1949]_ ;
  assign \new_[2297]_  = ~\new_[2519]_  | ~\new_[1950]_ ;
  assign \new_[2298]_  = ~\new_[2519]_  | ~\new_[1944]_ ;
  assign \new_[2299]_  = ~\new_[2519]_  | ~\new_[1891]_ ;
  assign \new_[2300]_  = ~\new_[2519]_  | ~\new_[1928]_ ;
  assign \new_[2301]_  = ~\new_[2519]_  | ~\new_[1945]_ ;
  assign \new_[2302]_  = ~\new_[2519]_  | ~\new_[1918]_ ;
  assign \new_[2303]_  = ~\new_[2519]_  | ~\new_[1939]_ ;
  assign \new_[2304]_  = ~\new_[2519]_  | ~\new_[1940]_ ;
  assign \new_[2305]_  = ~\new_[2519]_  | ~\new_[1946]_ ;
  assign \new_[2306]_  = ~\new_[2677]_  | ~\new_[2521]_ ;
  assign \new_[2307]_  = ~\new_[2812]_  | ~\new_[2520]_ ;
  assign \new_[2308]_  = ~\new_[3510]_ ;
  assign \new_[2309]_  = ~\new_[3320]_ ;
  assign n1176 = (~\new_[2670]_  & ~\new_[3102]_ ) | (~\new_[2598]_  & ~\new_[2138]_ );
  assign n1161 = (~\new_[2670]_  & ~\new_[3097]_ ) | (~\new_[2598]_  & ~\new_[2135]_ );
  assign n1181 = (~\new_[2670]_  & ~\new_[3107]_ ) | (~\new_[2598]_  & ~\new_[2139]_ );
  assign n1146 = (~\new_[2670]_  & ~\new_[3098]_ ) | (~\new_[2598]_  & ~\new_[2109]_ );
  assign n1171 = (~\new_[2670]_  & ~\new_[3073]_ ) | (~\new_[2598]_  & ~\new_[2137]_ );
  assign n1166 = (~\new_[2670]_  & ~\new_[3051]_ ) | (~\new_[2598]_  & ~\new_[2136]_ );
  assign n1156 = (~\new_[2670]_  & ~\new_[3075]_ ) | (~\new_[2598]_  & ~\new_[2126]_ );
  assign n1151 = (~\new_[2670]_  & ~\new_[3094]_ ) | (~\new_[2598]_  & ~\new_[2124]_ );
  assign \new_[2318]_  = \new_[3292]_  & \new_[383]_ ;
  assign \new_[2319]_  = \new_[3292]_  & \new_[373]_ ;
  assign \new_[2320]_  = \new_[3292]_  & \new_[374]_ ;
  assign \new_[2321]_  = \new_[3292]_  & \new_[377]_ ;
  assign \new_[2322]_  = \new_[3292]_  & \new_[389]_ ;
  assign \new_[2323]_  = \new_[3292]_  & \new_[381]_ ;
  assign \new_[2324]_  = \new_[3292]_  & \new_[384]_ ;
  assign \new_[2325]_  = \new_[3292]_  & \new_[388]_ ;
  assign \new_[2326]_  = \new_[3292]_  & \new_[382]_ ;
  assign \new_[2327]_  = \new_[3292]_  & \new_[387]_ ;
  assign \new_[2328]_  = \new_[3292]_  & \new_[386]_ ;
  assign \new_[2329]_  = \new_[3292]_  & \new_[390]_ ;
  assign \new_[2330]_  = \new_[3292]_  & \new_[391]_ ;
  assign \new_[2331]_  = \new_[3292]_  & \new_[375]_ ;
  assign \new_[2332]_  = \new_[2908]_  | \new_[2565]_ ;
  assign \new_[2333]_  = \new_[2842]_  | \new_[2565]_ ;
  assign \new_[2334]_  = \new_[2882]_  | \new_[2565]_ ;
  assign \new_[2335]_  = \new_[2877]_  | \new_[2562]_ ;
  assign \new_[2336]_  = \new_[2865]_  | \new_[2565]_ ;
  assign \new_[2337]_  = \new_[2803]_  | \new_[2565]_ ;
  assign \new_[2338]_  = \new_[2854]_  | \new_[2565]_ ;
  assign \new_[2339]_  = \new_[2873]_  | \new_[2565]_ ;
  assign \new_[2340]_  = \new_[2836]_  | \new_[2565]_ ;
  assign \new_[2341]_  = \new_[2861]_  | \new_[2565]_ ;
  assign \new_[2342]_  = \new_[2897]_  | \new_[2565]_ ;
  assign \new_[2343]_  = \new_[2901]_  | \new_[2565]_ ;
  assign \new_[2344]_  = \new_[2903]_  | \new_[2565]_ ;
  assign \new_[2345]_  = \new_[2805]_  | \new_[2562]_ ;
  assign \new_[2346]_  = \new_[2866]_  | \new_[2565]_ ;
  assign \new_[2347]_  = \new_[2864]_  | \new_[2562]_ ;
  assign \new_[2348]_  = \new_[2910]_  | \new_[2565]_ ;
  assign \new_[2349]_  = \new_[2863]_  | \new_[2562]_ ;
  assign \new_[2350]_  = \new_[2892]_  | \new_[2562]_ ;
  assign \new_[2351]_  = \new_[2931]_  | \new_[2562]_ ;
  assign \new_[2352]_  = \new_[2888]_  | \new_[2562]_ ;
  assign \new_[2353]_  = \new_[2875]_  | \new_[2565]_ ;
  assign \new_[2354]_  = \new_[2798]_  | \new_[2562]_ ;
  assign \new_[2355]_  = \new_[2849]_  | \new_[2565]_ ;
  assign \new_[2356]_  = ~\new_[3145]_  | ~\new_[2557]_  | ~\new_[1860]_ ;
  assign \new_[2357]_  = \new_[2758]_  & \new_[2579]_ ;
  assign \new_[2358]_  = ~\new_[3145]_  | ~\new_[2557]_  | ~\new_[1941]_ ;
  assign \new_[2359]_  = ~\new_[3145]_  | ~\new_[2557]_  | ~\new_[1942]_ ;
  assign \new_[2360]_  = ~\new_[2465]_ ;
  assign \new_[2361]_  = ~\new_[2563]_  & ~\new_[1665]_ ;
  assign \new_[2362]_  = ~\new_[2498]_ ;
  assign \new_[2363]_  = ~\new_[2465]_ ;
  assign \new_[2364]_  = \new_[2597]_  & \new_[327]_ ;
  assign \new_[2365]_  = \new_[2597]_  & \new_[324]_ ;
  assign \new_[2366]_  = \new_[2597]_  & \new_[325]_ ;
  assign \new_[2367]_  = \new_[2578]_  & \new_[328]_ ;
  assign \new_[2368]_  = \new_[2578]_  & \new_[358]_ ;
  assign \new_[2369]_  = \new_[2578]_  & \new_[362]_ ;
  assign \new_[2370]_  = \new_[2596]_  & \new_[333]_ ;
  assign \new_[2371]_  = ~\new_[2574]_  & ~\new_[3188]_ ;
  assign \new_[2372]_  = ~\new_[3424]_ ;
  assign \new_[2373]_  = ~\new_[2575]_  | ~\new_[2582]_ ;
  assign \new_[2374]_  = ~\new_[3293]_ ;
  assign \new_[2375]_  = \new_[2596]_  & \new_[371]_ ;
  assign \new_[2376]_  = \new_[2578]_  & \new_[369]_ ;
  assign \new_[2377]_  = \new_[3424]_ ;
  assign \new_[2378]_  = ~\new_[2587]_  & ~\new_[2585]_ ;
  assign \new_[2379]_  = \new_[1892]_  ^ \new_[2647]_ ;
  assign \new_[2380]_  = \new_[1665]_  ^ \new_[2656]_ ;
  assign \new_[2381]_  = (~\new_[3448]_  | ~\new_[3436]_ ) & (~\new_[3435]_  | ~\new_[3061]_ );
  assign n1211 = ~\new_[2715]_  | ~\new_[2787]_  | ~\new_[2556]_  | ~\new_[2661]_ ;
  assign \new_[2383]_  = \new_[3170]_  ^ \new_[2657]_ ;
  assign \new_[2384]_  = ~\new_[2754]_  | ~\new_[2822]_  | ~\new_[2817]_ ;
  assign \new_[2385]_  = \new_[2594]_  & \new_[2656]_ ;
  assign \new_[2386]_  = ~\new_[2685]_  & (~\new_[2650]_  | ~\new_[2747]_ );
  assign \new_[2387]_  = \new_[2601]_  & \new_[1789]_ ;
  assign \new_[2388]_  = ~\new_[2601]_  & ~\new_[1694]_ ;
  assign \new_[2389]_  = ~\new_[2488]_ ;
  assign n1191 = ~\new_[2703]_  | ~\new_[2792]_  | ~\new_[2571]_  | ~\new_[2655]_ ;
  assign n1206 = ~\new_[2706]_  | ~\new_[2826]_  | ~\new_[2570]_  | ~\new_[2658]_ ;
  assign n1186 = ~\new_[2709]_  | ~\new_[2840]_  | ~\new_[2568]_  | ~\new_[2649]_ ;
  assign n1196 = ~\new_[2724]_  | ~\new_[2790]_  | ~\new_[2589]_  | ~\new_[2663]_ ;
  assign n1201 = ~\new_[2727]_  | ~\new_[2829]_  | ~\new_[2569]_  | ~\new_[2629]_ ;
  assign \new_[2395]_  = \new_[3074]_  ? \new_[2621]_  : \new_[1690]_ ;
  assign \new_[2396]_  = ~\new_[3484]_ ;
  assign \new_[2397]_  = ~\new_[2553]_  & (~\new_[2942]_  | ~\new_[3051]_ );
  assign \new_[2398]_  = \new_[2800]_  | \new_[2553]_ ;
  assign \new_[2399]_  = \new_[2781]_  | \new_[2553]_ ;
  assign \new_[2400]_  = \new_[2831]_  | \new_[2553]_ ;
  assign \new_[2401]_  = \new_[2913]_  | \new_[2553]_ ;
  assign \new_[2402]_  = \new_[2894]_  | \new_[2553]_ ;
  assign \new_[2403]_  = \new_[2834]_  | \new_[2553]_ ;
  assign \new_[2404]_  = ~\new_[2553]_  & (~\new_[2944]_  | ~\new_[3097]_ );
  assign \new_[2405]_  = \new_[2860]_  | \new_[2553]_ ;
  assign \new_[2406]_  = \new_[2867]_  | \new_[2553]_ ;
  assign \new_[2407]_  = \new_[2869]_  | \new_[2553]_ ;
  assign \new_[2408]_  = \new_[2797]_  | \new_[2553]_ ;
  assign \new_[2409]_  = \new_[2870]_  | \new_[2553]_ ;
  assign \new_[2410]_  = \new_[2923]_  | \new_[2553]_ ;
  assign \new_[2411]_  = \new_[2852]_  | \new_[2553]_ ;
  assign \new_[2412]_  = \new_[2846]_  | \new_[2553]_ ;
  assign \new_[2413]_  = \new_[2917]_  | \new_[2553]_ ;
  assign \new_[2414]_  = \new_[2872]_  | \new_[2553]_ ;
  assign \new_[2415]_  = \new_[2874]_  | \new_[2553]_ ;
  assign \new_[2416]_  = \new_[2891]_  | \new_[2553]_ ;
  assign \new_[2417]_  = \new_[2921]_  | \new_[2553]_ ;
  assign \new_[2418]_  = \new_[2916]_  | \new_[2553]_ ;
  assign \new_[2419]_  = ~\new_[2554]_  & ~\new_[2918]_ ;
  assign \new_[2420]_  = ~\new_[2553]_  & (~\new_[2958]_  | ~\new_[3088]_ );
  assign \new_[2421]_  = \new_[2871]_  | \new_[2553]_ ;
  assign \new_[2422]_  = \new_[2883]_  | \new_[2553]_ ;
  assign \new_[2423]_  = ~\new_[2807]_  | ~\new_[2602]_ ;
  assign \new_[2424]_  = \new_[2898]_  | \new_[2553]_ ;
  assign \new_[2425]_  = \new_[2885]_  | \new_[2553]_ ;
  assign \new_[2426]_  = \new_[2830]_  | \new_[2553]_ ;
  assign \new_[2427]_  = \new_[2899]_  | \new_[2553]_ ;
  assign \new_[2428]_  = ~\new_[2553]_  & (~\new_[2811]_  | ~\new_[3078]_ );
  assign \new_[2429]_  = ~\new_[2809]_  | ~\new_[2602]_ ;
  assign \new_[2430]_  = ~\new_[2879]_  | ~\new_[2602]_ ;
  assign \new_[2431]_  = ~\new_[2804]_  | ~\new_[2602]_ ;
  assign \new_[2432]_  = ~\new_[2893]_  | ~\new_[2602]_ ;
  assign \new_[2433]_  = ~\new_[2784]_  | ~\new_[2602]_ ;
  assign \new_[2434]_  = ~\new_[2887]_  | ~\new_[2602]_ ;
  assign \new_[2435]_  = ~\new_[2926]_  | ~\new_[2602]_ ;
  assign \new_[2436]_  = ~\new_[2782]_  | ~\new_[2602]_ ;
  assign \new_[2437]_  = ~\new_[2828]_  | ~\new_[2602]_ ;
  assign \new_[2438]_  = ~\new_[2934]_  | ~\new_[2602]_ ;
  assign \new_[2439]_  = ~\new_[2802]_  | ~\new_[2602]_ ;
  assign \new_[2440]_  = ~\new_[2919]_  | ~\new_[2602]_ ;
  assign \new_[2441]_  = ~\new_[2884]_  | ~\new_[2602]_ ;
  assign \new_[2442]_  = ~\new_[2853]_  | ~\new_[2602]_ ;
  assign \new_[2443]_  = ~\new_[2799]_  | ~\new_[2602]_ ;
  assign \new_[2444]_  = ~\new_[2932]_  | ~\new_[2602]_ ;
  assign \new_[2445]_  = ~\new_[2835]_  | ~\new_[2602]_ ;
  assign \new_[2446]_  = ~\new_[2819]_  | ~\new_[2602]_ ;
  assign \new_[2447]_  = ~\new_[2868]_  | ~\new_[2602]_ ;
  assign \new_[2448]_  = ~\new_[2806]_  | ~\new_[2602]_ ;
  assign \new_[2449]_  = ~\new_[2889]_  | ~\new_[2602]_ ;
  assign \new_[2450]_  = ~\new_[2880]_  | ~\new_[2602]_ ;
  assign \new_[2451]_  = ~\new_[2896]_  | ~\new_[2602]_ ;
  assign \new_[2452]_  = ~\new_[2801]_  | ~\new_[2602]_ ;
  assign \new_[2453]_  = ~\new_[2808]_  | ~\new_[2602]_ ;
  assign \new_[2454]_  = ~\new_[2902]_  | ~\new_[2602]_ ;
  assign \new_[2455]_  = ~\new_[2848]_  | ~\new_[2602]_ ;
  assign \new_[2456]_  = ~\new_[2895]_  | ~\new_[2602]_ ;
  assign \new_[2457]_  = ~\new_[2878]_  | ~\new_[2602]_ ;
  assign \new_[2458]_  = \new_[2881]_  | \new_[2553]_ ;
  assign \new_[2459]_  = ~\new_[2810]_  | ~\new_[2602]_ ;
  assign \new_[2460]_  = ~\new_[2862]_  | ~\new_[2602]_ ;
  assign \new_[2461]_  = \new_[2900]_  | \new_[2565]_ ;
  assign \new_[2462]_  = \new_[2847]_  | \new_[2565]_ ;
  assign \new_[2463]_  = \new_[2928]_  | \new_[2565]_ ;
  assign \new_[2464]_  = \new_[2886]_  | \new_[2565]_ ;
  assign \new_[2465]_  = ~\new_[3365]_  & ~\new_[3292]_ ;
  assign \wb_dat_o[26]  = \\wb_dat_o_reg[26] ;
  assign \new_[2467]_  = \new_[2648]_  & \new_[363]_ ;
  assign \new_[2468]_  = \new_[2648]_  & \new_[360]_ ;
  assign \new_[2469]_  = \new_[2648]_  & \new_[339]_ ;
  assign \new_[2470]_  = \new_[2648]_  & \new_[367]_ ;
  assign \new_[2471]_  = \new_[2648]_  & \new_[335]_ ;
  assign \new_[2472]_  = \new_[2648]_  & \new_[336]_ ;
  assign \new_[2473]_  = \new_[2648]_  & \new_[337]_ ;
  assign \new_[2474]_  = \new_[2648]_  & \new_[368]_ ;
  assign \new_[2475]_  = \new_[2648]_  & \new_[359]_ ;
  assign \new_[2476]_  = \new_[2648]_  & \new_[370]_ ;
  assign \new_[2477]_  = \new_[2648]_  & \new_[366]_ ;
  assign \new_[2478]_  = ~\new_[2636]_  | ~\wb_sel_i[0] ;
  assign \new_[2479]_  = ~\new_[3364]_  | ~\new_[327]_ ;
  assign \new_[2480]_  = ~\new_[3364]_  | ~\new_[324]_ ;
  assign \new_[2481]_  = ~\new_[3364]_  | ~\new_[325]_ ;
  assign \wb_dat_o[16]  = \\wb_dat_o_reg[16] ;
  assign \new_[2483]_  = ~\new_[3308]_ ;
  assign \new_[2484]_  = ~\new_[2636]_  | ~\wb_sel_i[1] ;
  assign \ss_pad_o[0]  = ~\new_[2641]_  | ~\new_[3151]_ ;
  assign \ss_pad_o[1]  = ~\new_[2641]_  | ~\new_[3148]_ ;
  assign \new_[2487]_  = ~\new_[2597]_ ;
  assign \new_[2488]_  = ~\new_[2597]_ ;
  assign \new_[2489]_  = ~\new_[2639]_  | ~\new_[2676]_ ;
  assign \ss_pad_o[4]  = ~\new_[2641]_  | ~\new_[3135]_ ;
  assign \new_[2491]_  = ~\new_[3170]_  | ~\new_[2646]_  | ~\new_[3048]_ ;
  assign \ss_pad_o[2]  = ~\new_[2641]_  | ~\new_[3165]_ ;
  assign \new_[2493]_  = ~\new_[3331]_  & ~\new_[3143]_ ;
  assign \wb_dat_o[18]  = \\wb_dat_o_reg[18] ;
  assign \new_[2495]_  = ~\new_[2646]_  & (~\new_[2745]_  | ~\new_[1932]_ );
  assign \wb_dat_o[17]  = \\wb_dat_o_reg[17] ;
  assign \wb_dat_o[19]  = \\wb_dat_o_reg[19] ;
  assign \new_[2498]_  = ~\new_[2576]_ ;
  assign \wb_dat_o[22]  = \\wb_dat_o_reg[22] ;
  assign \wb_dat_o[27]  = \\wb_dat_o_reg[27] ;
  assign \wb_dat_o[21]  = \\wb_dat_o_reg[21] ;
  assign \wb_dat_o[31]  = \\wb_dat_o_reg[31] ;
  assign \wb_dat_o[28]  = \\wb_dat_o_reg[28] ;
  assign \wb_dat_o[24]  = \\wb_dat_o_reg[24] ;
  assign \wb_dat_o[23]  = \\wb_dat_o_reg[23] ;
  assign \wb_dat_o[30]  = \\wb_dat_o_reg[30] ;
  assign \wb_dat_o[20]  = \\wb_dat_o_reg[20] ;
  assign \wb_dat_o[29]  = \\wb_dat_o_reg[29] ;
  assign \wb_dat_o[25]  = \\wb_dat_o_reg[25] ;
  assign \ss_pad_o[7]  = ~\new_[2641]_  | ~\new_[3136]_ ;
  assign \ss_pad_o[6]  = ~\new_[2641]_  | ~\new_[3172]_ ;
  assign \ss_pad_o[5]  = ~\new_[2641]_  | ~\new_[3141]_ ;
  assign \ss_pad_o[3]  = ~\new_[2641]_  | ~\new_[3193]_ ;
  assign \new_[2514]_  = ~\new_[2591]_ ;
  assign \new_[2515]_  = ~\new_[2597]_ ;
  assign \new_[2516]_  = ~\new_[2818]_  | ~\new_[2651]_ ;
  assign n1236 = ~\new_[2711]_  | ~\new_[2789]_  | ~\new_[2628]_  | ~\new_[2763]_ ;
  assign n1216 = ~\new_[2696]_  | ~\new_[2825]_  | ~\new_[2634]_  | ~\new_[2762]_ ;
  assign \new_[2519]_  = ~\new_[2662]_  | ~\new_[1658]_ ;
  assign \new_[2520]_  = ~\new_[2664]_  | ~\new_[3436]_ ;
  assign \new_[2521]_  = ~\new_[2620]_  | ~\new_[3331]_ ;
  assign n1231 = ~\new_[2719]_  | ~\new_[2823]_  | ~\new_[2645]_  | ~\new_[2765]_ ;
  assign n1221 = ~\new_[2716]_  | ~\new_[2841]_  | ~\new_[2630]_  | ~\new_[2755]_ ;
  assign \new_[2524]_  = ~\new_[2591]_ ;
  assign \new_[2525]_  = \new_[2648]_  & \new_[341]_ ;
  assign n1226 = ~\new_[2666]_  | ~\new_[2753]_  | ~\new_[2767]_ ;
  assign n1241 = ~\new_[2669]_  | ~\new_[2714]_  | ~\new_[2779]_ ;
  assign \new_[2528]_  = ~\new_[2772]_  | ~\new_[2612]_ ;
  assign \new_[2529]_  = ~\new_[2667]_  & (~\new_[3025]_  | ~\new_[3075]_ );
  assign \new_[2530]_  = ~\new_[2667]_  & (~\new_[3021]_  | ~\new_[3055]_ );
  assign \new_[2531]_  = ~\new_[2667]_  & (~\new_[2961]_  | ~\new_[3058]_ );
  assign \new_[2532]_  = ~\new_[2667]_  & (~\new_[2993]_  | ~\new_[3093]_ );
  assign \new_[2533]_  = ~\new_[2667]_  & (~\new_[2979]_  | ~\new_[3094]_ );
  assign \new_[2534]_  = ~\new_[2667]_  & (~\new_[2945]_  | ~\new_[3054]_ );
  assign \new_[2535]_  = ~\new_[2667]_  & (~\new_[3017]_  | ~\new_[3072]_ );
  assign \new_[2536]_  = ~\new_[2667]_  & (~\new_[2943]_  | ~\new_[3034]_ );
  assign \new_[2537]_  = ~\new_[2667]_  & (~\new_[2998]_  | ~\new_[3052]_ );
  assign \new_[2538]_  = ~\new_[2667]_  & (~\new_[3013]_  | ~\new_[3060]_ );
  assign \new_[2539]_  = ~\new_[2667]_  & (~\new_[2972]_  | ~\new_[3090]_ );
  assign \new_[2540]_  = ~\new_[2667]_  & (~\new_[3028]_  | ~\new_[3078]_ );
  assign \new_[2541]_  = ~\new_[2667]_  & (~\new_[3020]_  | ~\new_[3105]_ );
  assign \new_[2542]_  = ~\new_[2667]_  & (~\new_[3023]_  | ~\new_[3041]_ );
  assign \new_[2543]_  = ~\new_[2667]_  & (~\new_[3026]_  | ~\new_[3092]_ );
  assign \new_[2544]_  = ~\new_[2667]_  & (~\new_[2975]_  | ~\new_[3083]_ );
  assign \new_[2545]_  = ~\new_[2667]_  & (~\new_[3027]_  | ~\new_[3051]_ );
  assign \new_[2546]_  = ~\new_[2667]_  & (~\new_[3006]_  | ~\new_[3070]_ );
  assign \new_[2547]_  = ~\new_[2667]_  & (~\new_[2980]_  | ~\new_[3091]_ );
  assign \new_[2548]_  = ~\new_[2667]_  & (~\new_[3016]_  | ~\new_[3073]_ );
  assign \new_[2549]_  = ~\new_[2667]_  & (~\new_[3015]_  | ~\new_[3108]_ );
  assign \new_[2550]_  = ~\new_[2667]_  & (~\new_[3029]_  | ~\new_[3047]_ );
  assign \new_[2551]_  = ~\new_[2667]_  & (~\new_[3005]_  | ~\new_[3088]_ );
  assign \new_[2552]_  = \new_[3382]_  & \new_[1789]_ ;
  assign \new_[2553]_  = ~\new_[2627]_  | ~\new_[3292]_ ;
  assign \new_[2554]_  = \new_[2668]_  | \new_[1935]_ ;
  assign \new_[2555]_  = ~\new_[3318]_ ;
  assign \new_[2556]_  = (~\new_[2832]_  | ~\new_[1940]_ ) & (~\new_[2731]_  | ~\new_[3165]_ );
  assign \new_[2557]_  = ~\new_[2623]_ ;
  assign \new_[2558]_  = ~\new_[2624]_ ;
  assign \new_[2559]_  = \new_[2627]_ ;
  assign \new_[2560]_  = ~\new_[3306]_ ;
  assign \new_[2561]_  = \new_[2624]_ ;
  assign \new_[2562]_  = ~\new_[3311]_ ;
  assign \new_[2563]_  = \new_[2912]_  | \new_[2678]_ ;
  assign \new_[2564]_  = \new_[2627]_ ;
  assign \new_[2565]_  = ~\new_[3308]_ ;
  assign \new_[2566]_  = (~\new_[2832]_  | ~\new_[1949]_ ) & (~\new_[2731]_  | ~\new_[3136]_ );
  assign \new_[2567]_  = (~\new_[2832]_  | ~\new_[1946]_ ) & (~\new_[2731]_  | ~\new_[3193]_ );
  assign \new_[2568]_  = (~\new_[2832]_  | ~\new_[1916]_ ) & (~\new_[2731]_  | ~\new_[3135]_ );
  assign \new_[2569]_  = (~\new_[2832]_  | ~\new_[1939]_ ) & (~\new_[2731]_  | ~\new_[3148]_ );
  assign \new_[2570]_  = (~\new_[2832]_  | ~\new_[1948]_ ) & (~\new_[2731]_  | ~\new_[3172]_ );
  assign \new_[2571]_  = (~\new_[2832]_  | ~\new_[1947]_ ) & (~\new_[2731]_  | ~\new_[3141]_ );
  assign \new_[2572]_  = ~\new_[2915]_  | ~\new_[2924]_  | ~\new_[2817]_  | ~\new_[2954]_ ;
  assign \new_[2573]_  = ~\new_[2672]_  & ~\new_[2824]_ ;
  assign \new_[2574]_  = ~\new_[2635]_ ;
  assign \new_[2575]_  = \new_[2735]_  & \new_[2672]_ ;
  assign \new_[2576]_  = ~\new_[2743]_  & (~\new_[3388]_  | ~\new_[1694]_ );
  assign \new_[2577]_  = ~\new_[2659]_ ;
  assign \new_[2578]_  = ~\new_[2637]_ ;
  assign \new_[2579]_  = ~\new_[2678]_  & ~\new_[1690]_ ;
  assign \new_[2580]_  = ~\new_[2676]_  | ~\new_[2735]_ ;
  assign \new_[2581]_  = ~\new_[2671]_  & ~\new_[2674]_ ;
  assign \new_[2582]_  = ~\new_[2671]_  & ~\new_[2775]_ ;
  assign \new_[2583]_  = ~\new_[2667]_  & (~\new_[2999]_  | ~\new_[3102]_ );
  assign \new_[2584]_  = ~\new_[2667]_  & (~\new_[2978]_  | ~\new_[3038]_ );
  assign \new_[2585]_  = ~\new_[2622]_ ;
  assign \new_[2586]_  = \new_[2076]_  ^ \new_[2746]_ ;
  assign \new_[2587]_  = ~\new_[2739]_  | ~\new_[2675]_ ;
  assign \new_[2588]_  = \new_[2617]_ ;
  assign \new_[2589]_  = (~\new_[2832]_  | ~\new_[1944]_ ) & (~\new_[2731]_  | ~\new_[3151]_ );
  assign \new_[2590]_  = ~\new_[3331]_ ;
  assign \new_[2591]_  = ~\new_[3222]_ ;
  assign \new_[2592]_  = ~\new_[2681]_  | ~\new_[1597]_ ;
  assign \new_[2593]_  = ~\new_[3081]_  | ~\new_[2682]_  | ~\new_[3053]_ ;
  assign \new_[2594]_  = ~\new_[2778]_  | ~\new_[1693]_ ;
  assign \new_[2595]_  = ~\new_[3053]_  | ~\new_[3049]_  | ~\new_[2730]_ ;
  assign \new_[2596]_  = ~\new_[2637]_ ;
  assign \new_[2597]_  = ~\new_[2637]_ ;
  assign \new_[2598]_  = ~\new_[2670]_  & ~\new_[3188]_ ;
  assign \new_[2599]_  = ~\new_[2673]_  | ~\new_[1658]_ ;
  assign \new_[2600]_  = ~\new_[2659]_ ;
  assign \new_[2601]_  = ~\new_[2620]_ ;
  assign \new_[2602]_  = ~\new_[3367]_  & ~\new_[3292]_ ;
  assign n1296 = ~\new_[2693]_  | ~\new_[2736]_ ;
  assign n1246 = ~\new_[2697]_  | ~\new_[2723]_ ;
  assign n1316 = ~\new_[2738]_  | ~\new_[2686]_ ;
  assign n1306 = ~\new_[2712]_  | ~\new_[2701]_ ;
  assign n1286 = ~\new_[2752]_  | ~\new_[2684]_ ;
  assign n1321 = ~\new_[2718]_  | ~\new_[2720]_ ;
  assign n1276 = ~\new_[2694]_  | ~\new_[2750]_ ;
  assign n1291 = ~\new_[2721]_  | ~\new_[2749]_ ;
  assign n1256 = ~\new_[2726]_  | ~\new_[2704]_ ;
  assign \new_[2612]_  = ~\new_[3383]_  | ~\new_[2820]_ ;
  assign n1311 = ~\new_[2700]_  | ~\new_[2705]_ ;
  assign n1251 = ~\new_[2717]_  | ~\new_[2708]_ ;
  assign n1261 = ~\new_[2733]_  | ~\new_[2725]_ ;
  assign n1266 = ~\new_[2702]_  | ~\new_[2734]_ ;
  assign \new_[2617]_  = ~\new_[3308]_ ;
  assign n1281 = ~\new_[2699]_  | ~\new_[2722]_ ;
  assign n1271 = ~\new_[2710]_  | ~\new_[2692]_ ;
  assign \new_[2620]_  = ~\new_[2689]_  | ~\new_[2778]_ ;
  assign \new_[2621]_  = ~\new_[1665]_  | ~\new_[2911]_  | ~\new_[2776]_ ;
  assign \new_[2622]_  = ~\new_[3459]_ ;
  assign \new_[2623]_  = \new_[2729]_  & \new_[2947]_ ;
  assign \new_[2624]_  = ~\new_[3306]_ ;
  assign \new_[2625]_  = ~\new_[3312]_ ;
  assign \new_[2626]_  = \new_[3308]_ ;
  assign \new_[2627]_  = ~\new_[3306]_ ;
  assign \new_[2628]_  = (~\new_[2832]_  | ~\new_[1923]_ ) & (~\new_[3158]_  | ~\new_[2768]_ );
  assign \new_[2629]_  = (~\new_[1936]_  | ~\new_[2768]_ ) & (~\new_[442]_  | ~\new_[2858]_ );
  assign \new_[2630]_  = (~\new_[2832]_  | ~\new_[1928]_ ) & (~\new_[2768]_  | ~\new_[3119]_ );
  assign \new_[2631]_  = (~\new_[3173]_  | ~\new_[2768]_ ) & (~\new_[505]_  | ~\new_[2858]_ );
  assign \new_[2632]_  = ~\new_[3312]_ ;
  assign \new_[2633]_  = (~\new_[1941]_  | ~\new_[2768]_ ) & (~\new_[509]_  | ~\new_[2858]_ );
  assign \new_[2634]_  = (~\new_[2832]_  | ~\new_[1938]_ ) & (~\new_[1712]_  | ~\new_[2768]_ );
  assign \new_[2635]_  = ~\new_[2857]_  & ~\new_[2742]_ ;
  assign \new_[2636]_  = ~\new_[2680]_ ;
  assign \new_[2637]_  = ~\new_[3225]_ ;
  assign \new_[2638]_  = ~\new_[2735]_  | ~\new_[2747]_ ;
  assign \new_[2639]_  = ~\new_[2735]_  | ~\new_[2824]_ ;
  assign \new_[2640]_  = ~\new_[2775]_  & ~\new_[2685]_ ;
  assign \new_[2641]_  = ~\new_[3145]_  | ~\new_[3119]_ ;
  assign \new_[2642]_  = ~\new_[1665]_  & ~\new_[1789]_ ;
  assign \new_[2643]_  = \new_[3451]_  | \new_[3150]_ ;
  assign \new_[2644]_  = ~\new_[3112]_  & ~\new_[1789]_ ;
  assign \new_[2645]_  = (~\new_[2832]_  | ~\new_[1937]_ ) & (~\new_[2768]_  | ~\new_[3159]_ );
  assign \new_[2646]_  = ~\new_[2745]_  & ~\new_[1932]_ ;
  assign \new_[2647]_  = \new_[2953]_  & \new_[2746]_ ;
  assign \new_[2648]_  = \new_[3225]_ ;
  assign \new_[2649]_  = (~\new_[1942]_  | ~\new_[2768]_ ) & (~\new_[506]_  | ~\new_[2858]_ );
  assign \new_[2650]_  = ~\new_[2676]_ ;
  assign \new_[2651]_  = ~\new_[2728]_  | ~\new_[3436]_ ;
  assign \new_[2652]_  = ~\new_[3331]_  | ~\new_[1690]_ ;
  assign \new_[2653]_  = ~\new_[2690]_  | ~\new_[2761]_ ;
  assign n1301 = ~\new_[2713]_  | ~\new_[2751]_ ;
  assign \new_[2655]_  = (~\new_[1926]_  | ~\new_[2768]_ ) & (~\new_[557]_  | ~\new_[2858]_ );
  assign \new_[2656]_  = ~\new_[2754]_  | ~\new_[3150]_ ;
  assign \new_[2657]_  = ~\new_[2682]_ ;
  assign \new_[2658]_  = (~\new_[1943]_  | ~\new_[2768]_ ) & (~\new_[558]_  | ~\new_[2858]_ );
  assign \new_[2659]_  = ~\new_[3225]_ ;
  assign \new_[2660]_  = \new_[1934]_  ^ \new_[2757]_ ;
  assign \new_[2661]_  = (~\new_[1917]_  | ~\new_[2768]_ ) & (~\new_[465]_  | ~\new_[2858]_ );
  assign \new_[2662]_  = \new_[2788]_  | \new_[1930]_  | \new_[2918]_  | \new_[1935]_ ;
  assign \new_[2663]_  = (~\new_[1860]_  | ~\new_[2768]_ ) & (~\new_[508]_  | ~\new_[2858]_ );
  assign \new_[2664]_  = \new_[3143]_  ? \new_[2760]_  : \new_[1665]_ ;
  assign \new_[2665]_  = ~\new_[3486]_ ;
  assign \new_[2666]_  = (~\new_[2832]_  | ~\new_[1945]_ ) & (~\new_[347]_  | ~\new_[2955]_ );
  assign \new_[2667]_  = \new_[3222]_  | \new_[3365]_ ;
  assign \new_[2668]_  = ~\new_[2766]_  | ~\new_[1930]_ ;
  assign \new_[2669]_  = (~\new_[2832]_  | ~\new_[1918]_ ) & (~\new_[348]_  | ~\new_[2955]_ );
  assign \new_[2670]_  = ~\wb_adr_i[3]  | ~\wb_adr_i[4]  | ~\new_[2774]_  | ~wb_we_i;
  assign \new_[2671]_  = ~\new_[2739]_ ;
  assign \new_[2672]_  = ~\new_[2771]_  & ~\new_[3386]_ ;
  assign \new_[2673]_  = \new_[3137]_  ^ \new_[2954]_ ;
  assign \new_[2674]_  = ~\new_[2685]_ ;
  assign \new_[2675]_  = ~\new_[1942]_  | ~\new_[3143]_ ;
  assign \new_[2676]_  = ~\new_[1917]_  | ~\new_[2924]_ ;
  assign \new_[2677]_  = \new_[2820]_  | \new_[2924]_ ;
  assign \new_[2678]_  = ~\new_[3150]_  | ~\new_[2924]_ ;
  assign \new_[2679]_  = \new_[2004]_  ^ \new_[2837]_ ;
  assign \new_[2680]_  = ~\new_[2920]_  | ~wb_we_i | ~\new_[2814]_  | ~\new_[2946]_ ;
  assign \new_[2681]_  = ~\new_[1665]_  | ~\new_[2827]_  | ~\new_[2786]_ ;
  assign \new_[2682]_  = \new_[3048]_  & \new_[2777]_ ;
  assign \new_[2683]_  = ~\new_[2756]_  & ~\new_[3122]_ ;
  assign \new_[2684]_  = (~\new_[447]_  | ~\new_[2858]_ ) & (~\new_[341]_  | ~\new_[2951]_ );
  assign \new_[2685]_  = ~\new_[3124]_  & ~\new_[1693]_ ;
  assign \new_[2686]_  = (~\new_[444]_  | ~\new_[2858]_ ) & (~\new_[339]_  | ~\new_[2951]_ );
  assign \new_[2687]_  = \new_[1929]_  ^ \new_[2925]_ ;
  assign \new_[2688]_  = (~\new_[331]_  | ~\new_[2951]_ ) & (~\new_[324]_  | ~\new_[2856]_ );
  assign \new_[2689]_  = ~\new_[2912]_  | ~\new_[3112]_ ;
  assign \new_[2690]_  = ~\new_[2794]_  & ~\new_[2795]_ ;
  assign \new_[2691]_  = ~\new_[2759]_ ;
  assign \new_[2692]_  = (~\new_[391]_  | ~\new_[2955]_ ) & (~\new_[393]_  | ~\new_[2856]_ );
  assign \new_[2693]_  = (~\new_[375]_  | ~\new_[2955]_ ) & (~\new_[325]_  | ~\new_[2856]_ );
  assign \new_[2694]_  = (~\new_[374]_  | ~\new_[2955]_ ) & (~\new_[434]_  | ~\new_[2856]_ );
  assign \new_[2695]_  = (~\new_[358]_  | ~\new_[2951]_ ) & (~\new_[426]_  | ~\new_[2856]_ );
  assign \new_[2696]_  = (~\new_[332]_  | ~\new_[2951]_ ) & (~\new_[499]_  | ~\new_[2856]_ );
  assign \new_[2697]_  = (~\new_[433]_  | ~\new_[2856]_ ) & (~\new_[370]_  | ~\new_[2951]_ );
  assign \new_[2698]_  = (~\new_[2951]_  | ~\new_[362]_ ) & (~\new_[2856]_  | ~\new_[486]_ );
  assign \new_[2699]_  = (~\new_[390]_  | ~\new_[2955]_ ) & (~\new_[392]_  | ~\new_[2856]_ );
  assign \new_[2700]_  = (~\new_[353]_  | ~\new_[2955]_ ) & (~\new_[503]_  | ~\new_[2856]_ );
  assign \new_[2701]_  = (~\new_[445]_  | ~\new_[2858]_ ) & (~\new_[340]_  | ~\new_[2951]_ );
  assign \new_[2702]_  = (~\new_[528]_  | ~\new_[2858]_ ) & (~\new_[365]_  | ~\new_[2951]_ );
  assign \new_[2703]_  = (~\new_[359]_  | ~\new_[2951]_ ) & (~\new_[496]_  | ~\new_[2856]_ );
  assign \new_[2704]_  = (~\new_[468]_  | ~\new_[2858]_ ) & (~\new_[369]_  | ~\new_[2951]_ );
  assign \new_[2705]_  = (~\new_[498]_  | ~\new_[2858]_ ) & (~\new_[366]_  | ~\new_[2951]_ );
  assign \new_[2706]_  = (~\new_[360]_  | ~\new_[2951]_ ) & (~\new_[497]_  | ~\new_[2856]_ );
  assign \new_[2707]_  = (~\new_[333]_  | ~\new_[2951]_ ) & (~\new_[428]_  | ~\new_[2856]_ );
  assign \new_[2708]_  = (~\new_[349]_  | ~\new_[2955]_ ) & (~\new_[482]_  | ~\new_[2856]_ );
  assign \new_[2709]_  = (~\new_[330]_  | ~\new_[2951]_ ) & (~\new_[427]_  | ~\new_[2856]_ );
  assign \new_[2710]_  = (~\new_[524]_  | ~\new_[2858]_ ) & (~\new_[336]_  | ~\new_[2951]_ );
  assign \new_[2711]_  = (~\new_[361]_  | ~\new_[2951]_ ) & (~\new_[488]_  | ~\new_[2856]_ );
  assign \new_[2712]_  = (~\new_[378]_  | ~\new_[2955]_ ) & (~\new_[436]_  | ~\new_[2856]_ );
  assign \new_[2713]_  = (~\new_[354]_  | ~\new_[2955]_ ) & (~\new_[504]_  | ~\new_[2856]_ );
  assign \new_[2714]_  = (~\new_[438]_  | ~\new_[2858]_ ) & (~\new_[371]_  | ~\new_[2951]_ );
  assign \new_[2715]_  = (~\new_[329]_  | ~\new_[2951]_ ) & (~\new_[425]_  | ~\new_[2856]_ );
  assign \new_[2716]_  = (~\new_[363]_  | ~\new_[2951]_ ) & (~\new_[429]_  | ~\new_[2856]_ );
  assign \new_[2717]_  = (~\new_[439]_  | ~\new_[2858]_ ) & (~\new_[364]_  | ~\new_[2951]_ );
  assign \new_[2718]_  = (~\new_[383]_  | ~\new_[2955]_ ) & (~\new_[432]_  | ~\new_[2856]_ );
  assign \new_[2719]_  = (~\new_[334]_  | ~\new_[2951]_ ) & (~\new_[502]_  | ~\new_[2856]_ );
  assign \new_[2720]_  = (~\new_[441]_  | ~\new_[2858]_ ) & (~\new_[356]_  | ~\new_[2951]_ );
  assign \new_[2721]_  = (~\new_[377]_  | ~\new_[2955]_ ) & (~\new_[474]_  | ~\new_[2856]_ );
  assign \new_[2722]_  = (~\new_[562]_  | ~\new_[2858]_ ) & (~\new_[335]_  | ~\new_[2951]_ );
  assign \new_[2723]_  = (~\new_[446]_  | ~\new_[2858]_ ) & (~\new_[373]_  | ~\new_[2955]_ );
  assign \new_[2724]_  = (~\new_[357]_  | ~\new_[2951]_ ) & (~\new_[327]_  | ~\new_[2856]_ );
  assign \new_[2725]_  = (~\new_[350]_  | ~\new_[2955]_ ) & (~\new_[500]_  | ~\new_[2856]_ );
  assign \new_[2726]_  = (~\new_[351]_  | ~\new_[2955]_ ) & (~\new_[501]_  | ~\new_[2856]_ );
  assign \new_[2727]_  = (~\new_[328]_  | ~\new_[2951]_ ) & (~\new_[424]_  | ~\new_[2856]_ );
  assign \new_[2728]_  = ~\new_[2833]_  | ~\new_[2851]_ ;
  assign \new_[2729]_  = ~\new_[2796]_  & ~\new_[1860]_ ;
  assign \new_[2730]_  = ~\new_[2757]_ ;
  assign \new_[2731]_  = ~\new_[2904]_  & ~\new_[3189]_ ;
  assign \new_[2732]_  = ~\new_[2850]_  & ~\new_[2813]_ ;
  assign \new_[2733]_  = (~\new_[494]_  | ~\new_[2858]_ ) & (~\new_[367]_  | ~\new_[2951]_ );
  assign \new_[2734]_  = (~\new_[389]_  | ~\new_[2955]_ ) & (~\new_[394]_  | ~\new_[2856]_ );
  assign \new_[2735]_  = ~\new_[3140]_  | ~\new_[3112]_ ;
  assign \new_[2736]_  = (~\new_[492]_  | ~\new_[2858]_ ) & (~\new_[368]_  | ~\new_[2951]_ );
  assign \new_[2737]_  = ~sclk_pad_o & ~\new_[3145]_ ;
  assign \new_[2738]_  = (~\new_[376]_  | ~\new_[2955]_ ) & (~\new_[435]_  | ~\new_[2856]_ );
  assign \new_[2739]_  = ~\new_[3190]_  | ~\new_[1665]_ ;
  assign \new_[2740]_  = ~\new_[2964]_  & (~\wb_sel_i[0]  | ~\new_[1860]_ );
  assign \new_[2741]_  = ~\new_[2952]_  & ~\new_[1789]_ ;
  assign \new_[2742]_  = ~\new_[2814]_  | ~\new_[2920]_ ;
  assign \new_[2743]_  = ~\new_[2927]_  & (~\new_[3122]_  | ~\new_[1694]_ );
  assign \new_[2744]_  = \new_[1933]_  ^ \new_[2845]_ ;
  assign \new_[2745]_  = ~\new_[3196]_  | ~\new_[2837]_  | ~\new_[3059]_ ;
  assign \new_[2746]_  = \new_[2837]_  & \new_[2938]_ ;
  assign \new_[2747]_  = ~\new_[2775]_ ;
  assign \new_[2748]_  = ~\new_[2837]_  & (~\new_[2936]_  | ~\new_[1927]_ );
  assign \new_[2749]_  = (~\new_[464]_  | ~\new_[2858]_ ) & (~\new_[355]_  | ~\new_[2951]_ );
  assign \new_[2750]_  = (~\new_[443]_  | ~\new_[2858]_ ) & (~\new_[338]_  | ~\new_[2951]_ );
  assign \new_[2751]_  = (~\new_[440]_  | ~\new_[2858]_ ) & (~\new_[337]_  | ~\new_[2951]_ );
  assign \new_[2752]_  = (~\new_[379]_  | ~\new_[2955]_ ) & (~\new_[326]_  | ~\new_[2856]_ );
  assign \new_[2753]_  = (~\new_[561]_  | ~\new_[2858]_ ) & (~\new_[372]_  | ~\new_[2951]_ );
  assign \new_[2754]_  = ~\new_[2778]_ ;
  assign \new_[2755]_  = ~\new_[560]_  | ~\new_[2858]_ ;
  assign \new_[2756]_  = ~\new_[2855]_  | ~\new_[2941]_ ;
  assign \new_[2757]_  = \new_[1929]_  | \new_[2076]_  | \new_[2925]_  | \new_[2959]_ ;
  assign \new_[2758]_  = ~\new_[1665]_  & ~\new_[2912]_ ;
  assign \new_[2759]_  = ~\new_[3451]_  & (~\new_[2935]_  | ~\new_[2957]_ );
  assign \new_[2760]_  = ~\new_[2911]_  | ~\new_[3244]_ ;
  assign \new_[2761]_  = ~\new_[1581]_  & ~\new_[1658]_ ;
  assign \new_[2762]_  = ~\new_[507]_  | ~\new_[2858]_ ;
  assign \new_[2763]_  = ~\new_[437]_  | ~\new_[2858]_ ;
  assign \new_[2764]_  = ~\new_[559]_  | ~\new_[2858]_ ;
  assign \new_[2765]_  = ~\new_[495]_  | ~\new_[2858]_ ;
  assign \new_[2766]_  = ~\new_[2788]_ ;
  assign \new_[2767]_  = ~\new_[430]_  | ~\new_[2856]_ ;
  assign \new_[2768]_  = ~\new_[2904]_  & ~\wb_adr_i[3] ;
  assign wb_ack_o = wb_ack_o_reg;
  assign \new_[2770]_  = ~\new_[2818]_ ;
  assign \new_[2771]_  = ~\new_[1936]_  & ~\new_[3014]_ ;
  assign \new_[2772]_  = \new_[3435]_  | \new_[2915]_ ;
  assign \new_[2773]_  = ~\new_[2858]_  | ~\new_[493]_ ;
  assign \new_[2774]_  = \new_[2920]_  & \new_[3009]_ ;
  assign \new_[2775]_  = ~\new_[1941]_  & ~\new_[3150]_ ;
  assign \new_[2776]_  = ~\new_[2815]_ ;
  assign \new_[2777]_  = ~\new_[2845]_  & ~\new_[2959]_ ;
  assign \new_[2778]_  = ~\new_[3014]_  | ~\new_[2924]_  | ~\new_[3012]_ ;
  assign \new_[2779]_  = ~\new_[431]_  | ~\new_[2856]_ ;
  assign \new_[2780]_  = ~\new_[2955]_  | ~\new_[388]_ ;
  assign \new_[2781]_  = ~\new_[2960]_  & (~\new_[3188]_  | ~\new_[425]_ );
  assign \new_[2782]_  = ~\new_[3097]_  | (~\wb_sel_i[0]  & ~\new_[3123]_ );
  assign \new_[2783]_  = ~\new_[2843]_ ;
  assign \new_[2784]_  = ~\new_[3102]_  | (~\wb_sel_i[0]  & ~\new_[3174]_ );
  assign \new_[2785]_  = \new_[2949]_  & \new_[2936]_ ;
  assign \new_[2786]_  = ~\new_[2933]_ ;
  assign \new_[2787]_  = ~\new_[343]_  | ~\new_[2955]_ ;
  assign \new_[2788]_  = ~\new_[2953]_  | ~\new_[2938]_ ;
  assign \new_[2789]_  = ~\new_[346]_  | ~\new_[2955]_ ;
  assign \new_[2790]_  = ~\new_[342]_  | ~\new_[2955]_ ;
  assign \new_[2791]_  = ~\new_[345]_  | ~\new_[2955]_ ;
  assign \new_[2792]_  = ~\new_[382]_  | ~\new_[2955]_ ;
  assign \new_[2793]_  = ~\new_[2933]_ ;
  assign \new_[2794]_  = ~\new_[3039]_  | ~\new_[3063]_  | ~\new_[3110]_  | ~\new_[3085]_ ;
  assign \new_[2795]_  = ~\new_[3076]_  | ~\new_[3066]_  | ~\new_[3101]_  | ~\new_[3064]_ ;
  assign \new_[2796]_  = ~\new_[3175]_  | ~\new_[3095]_  | ~\new_[3124]_  | ~\new_[3190]_ ;
  assign \new_[2797]_  = ~\new_[3002]_  & (~\new_[3106]_  | ~\new_[428]_ );
  assign \new_[2798]_  = ~\new_[2987]_  & (~\new_[3080]_  | ~\new_[390]_ );
  assign \new_[2799]_  = ~\new_[3060]_  | (~\wb_sel_i[1]  & ~\new_[3164]_ );
  assign \new_[2800]_  = ~\new_[3018]_  & (~\new_[3188]_  | ~\new_[424]_ );
  assign \new_[2801]_  = ~\new_[3108]_  | (~\wb_sel_i[3]  & ~\new_[3157]_ );
  assign \new_[2802]_  = ~\new_[3034]_  | (~\wb_sel_i[1]  & ~\new_[3131]_ );
  assign \new_[2803]_  = ~\new_[2985]_  & (~\new_[3080]_  | ~\new_[349]_ );
  assign \new_[2804]_  = ~\new_[3073]_  | (~\wb_sel_i[0]  & ~\new_[3163]_ );
  assign \new_[2805]_  = ~\new_[2996]_  & (~\new_[3188]_  | ~\new_[345]_ );
  assign \new_[2806]_  = ~\new_[3043]_  | (~\wb_sel_i[2]  & ~\new_[3198]_ );
  assign \new_[2807]_  = ~\new_[3091]_  | (~\wb_sel_i[3]  & ~\new_[3154]_ );
  assign \new_[2808]_  = ~\new_[3087]_  | (~\wb_sel_i[3]  & ~\new_[3147]_ );
  assign \new_[2809]_  = ~\new_[3051]_  | (~\wb_sel_i[0]  & ~\new_[3115]_ );
  assign \new_[2810]_  = ~\new_[3047]_  | (~\wb_sel_i[3]  & ~\new_[3162]_ );
  assign \new_[2811]_  = ~\new_[3120]_  | ~\new_[326]_ ;
  assign \new_[2812]_  = ~\new_[3435]_  | ~\new_[1665]_ ;
  assign \new_[2813]_  = ~\new_[3175]_  & ~\new_[1690]_ ;
  assign \new_[2814]_  = \new_[3189]_  & \wb_adr_i[4] ;
  assign \new_[2815]_  = ~\new_[2956]_  | ~\new_[2952]_ ;
  assign \new_[2816]_  = ~\new_[1690]_  & ~\new_[1789]_ ;
  assign \new_[2817]_  = \new_[3143]_  & \new_[3150]_ ;
  assign \new_[2818]_  = ~\new_[3332]_  | ~\new_[3112]_ ;
  assign \new_[2819]_  = ~\new_[3105]_  | (~\wb_sel_i[2]  & ~\new_[3161]_ );
  assign \new_[2820]_  = ~\new_[3436]_ ;
  assign \new_[2821]_  = ~\new_[1597]_  & ~\new_[1789]_ ;
  assign \new_[2822]_  = ~\new_[1690]_  & ~\new_[1597]_ ;
  assign \new_[2823]_  = ~\new_[385]_  | ~\new_[2955]_ ;
  assign \new_[2824]_  = ~\new_[3319]_  & ~\new_[2952]_ ;
  assign \new_[2825]_  = ~\new_[380]_  | ~\new_[2955]_ ;
  assign \new_[2826]_  = ~\new_[384]_  | ~\new_[2955]_ ;
  assign \new_[2827]_  = ~\new_[3150]_  & ~\new_[3074]_ ;
  assign \new_[2828]_  = ~\new_[3054]_  | (~\wb_sel_i[1]  & ~\new_[3168]_ );
  assign \new_[2829]_  = ~\new_[352]_  | ~\new_[2955]_ ;
  assign \new_[2830]_  = ~\new_[2992]_  & (~\new_[3120]_  | ~\new_[435]_ );
  assign \new_[2831]_  = ~\new_[2984]_  & (~\new_[3188]_  | ~\new_[426]_ );
  assign \new_[2832]_  = ~\new_[2939]_  & ~\wb_adr_i[3] ;
  assign \new_[2833]_  = ~\new_[2937]_  | ~\new_[3112]_ ;
  assign \new_[2834]_  = ~\new_[2962]_  & (~\new_[3188]_  | ~\new_[497]_ );
  assign \new_[2835]_  = ~\new_[3056]_  | (~\wb_sel_i[1]  & ~\new_[3156]_ );
  assign \new_[2836]_  = ~\new_[2997]_  & (~\new_[3120]_  | ~\new_[374]_ );
  assign \new_[2837]_  = ~\new_[2936]_  & ~\new_[1927]_ ;
  assign \new_[2838]_  = ~\new_[381]_  | ~\new_[2955]_ ;
  assign \new_[2839]_  = ~\new_[387]_  | ~\new_[2955]_ ;
  assign \new_[2840]_  = ~\new_[344]_  | ~\new_[2955]_ ;
  assign \new_[2841]_  = ~\new_[386]_  | ~\new_[2955]_ ;
  assign \new_[2842]_  = ~\new_[2967]_  & (~\new_[3120]_  | ~\new_[378]_ );
  assign \new_[2843]_  = ~wb_we_i | ~\new_[3033]_  | ~\new_[3082]_ ;
  assign \new_[2844]_  = ~\new_[3003]_  & (~\new_[3080]_  | ~\new_[504]_ );
  assign \new_[2845]_  = ~\new_[3062]_  | ~\new_[3059]_  | ~\new_[3036]_ ;
  assign \new_[2846]_  = ~\new_[2986]_  & (~\new_[3106]_  | ~\new_[431]_ );
  assign \new_[2847]_  = ~\new_[2982]_  & (~\new_[3120]_  | ~\new_[373]_ );
  assign \new_[2848]_  = ~\new_[3078]_  | (~\wb_sel_i[3]  & ~\new_[3045]_ );
  assign \new_[2849]_  = ~\new_[2991]_  & (~\new_[3120]_  | ~\new_[375]_ );
  assign \new_[2850]_  = ~\new_[1926]_  & ~\new_[3074]_ ;
  assign \new_[2851]_  = ~\new_[3244]_  | ~\new_[3127]_ ;
  assign \new_[2852]_  = ~\new_[2968]_  & (~\new_[3106]_  | ~\new_[430]_ );
  assign \new_[2853]_  = ~\new_[3088]_  | (~\wb_sel_i[3]  & ~\new_[3037]_ );
  assign \new_[2854]_  = ~\new_[2964]_  & (~\new_[3188]_  | ~\new_[342]_ );
  assign \new_[2855]_  = ~\new_[2940]_ ;
  assign \new_[2856]_  = ~\new_[3000]_  & ~\wb_adr_i[3] ;
  assign \new_[2857]_  = ~\new_[3009]_  | ~wb_we_i;
  assign \new_[2858]_  = ~\new_[3000]_  & ~\new_[3189]_ ;
  assign \new_[2859]_  = ~\new_[3022]_  | ~\new_[3019]_ ;
  assign \new_[2860]_  = ~\new_[3004]_  & (~\new_[3106]_  | ~\new_[488]_ );
  assign \new_[2861]_  = ~\new_[2986]_  & (~\new_[3106]_  | ~\new_[348]_ );
  assign \new_[2862]_  = ~\new_[3083]_  | (~\wb_sel_i[2]  & ~\new_[3096]_ );
  assign \new_[2863]_  = ~\new_[3002]_  & (~\new_[3106]_  | ~\new_[387]_ );
  assign \new_[2864]_  = ~\new_[2990]_  & (~\new_[3080]_  | ~\new_[353]_ );
  assign \new_[2865]_  = ~\new_[2984]_  & (~\new_[3188]_  | ~\new_[381]_ );
  assign \new_[2866]_  = ~\new_[2962]_  & (~\new_[3188]_  | ~\new_[384]_ );
  assign \new_[2867]_  = ~\new_[3001]_  & (~\new_[3106]_  | ~\new_[486]_ );
  assign \new_[2868]_  = ~\new_[3092]_  | (~\wb_sel_i[2]  & ~\new_[3065]_ );
  assign \new_[2869]_  = ~\new_[3007]_  & (~\new_[3106]_  | ~\new_[499]_ );
  assign \new_[2870]_  = ~\new_[2974]_  & (~\new_[3106]_  | ~\new_[502]_ );
  assign \new_[2871]_  = ~\new_[2983]_  & (~\new_[3120]_  | ~\new_[432]_ );
  assign \new_[2872]_  = ~\new_[3008]_  & (~\new_[3080]_  | ~\new_[500]_ );
  assign \new_[2873]_  = ~\new_[2971]_  & (~\new_[3188]_  | ~\new_[344]_ );
  assign \new_[2874]_  = ~\new_[2969]_  & (~\new_[3080]_  | ~\new_[501]_ );
  assign \new_[2875]_  = ~\new_[2995]_  & (~\new_[3080]_  | ~\new_[389]_ );
  assign \new_[2876]_  = ~\new_[3010]_  & (~\new_[3080]_  | ~\new_[391]_ );
  assign \new_[2877]_  = ~\new_[2969]_  & (~\new_[3080]_  | ~\new_[351]_ );
  assign \new_[2878]_  = ~\new_[3041]_  | (~\wb_sel_i[2]  & ~\new_[3035]_ );
  assign \new_[2879]_  = ~\new_[3075]_  | (~\wb_sel_i[0]  & ~\new_[3086]_ );
  assign \new_[2880]_  = ~\new_[3038]_  | (~\wb_sel_i[2]  & ~\new_[3030]_ );
  assign \new_[2881]_  = ~\new_[3010]_  & (~\new_[3080]_  | ~\new_[393]_ );
  assign \new_[2882]_  = ~\new_[2988]_  & (~\new_[3120]_  | ~\new_[379]_ );
  assign \new_[2883]_  = ~\new_[2982]_  & (~\new_[3120]_  | ~\new_[433]_ );
  assign \new_[2884]_  = ~\new_[3090]_  | (~\wb_sel_i[1]  & ~\new_[3111]_ );
  assign \new_[2885]_  = ~\new_[2989]_  & (~\new_[3120]_  | ~\new_[474]_ );
  assign \new_[2886]_  = ~\new_[2992]_  & (~\new_[3120]_  | ~\new_[376]_ );
  assign \new_[2887]_  = ~\new_[3098]_  | (~\wb_sel_i[0]  & ~\new_[3089]_ );
  assign \new_[2888]_  = ~\new_[3008]_  & (~\new_[3080]_  | ~\new_[350]_ );
  assign \new_[2889]_  = ~\new_[3070]_  | (~\wb_sel_i[2]  & ~\new_[3050]_ );
  assign \new_[2890]_  = ~\new_[3018]_  & (~\new_[3188]_  | ~\new_[352]_ );
  assign \new_[2891]_  = ~\new_[2995]_  & (~\new_[3080]_  | ~\new_[394]_ );
  assign \new_[2892]_  = ~\new_[3001]_  & (~\new_[3106]_  | ~\new_[388]_ );
  assign \new_[2893]_  = ~\new_[3094]_  | (~\wb_sel_i[0]  & ~\new_[3079]_ );
  assign \new_[2894]_  = ~\new_[2966]_  & (~\new_[3188]_  | ~\new_[496]_ );
  assign \new_[2895]_  = ~\new_[3055]_  | (~\wb_sel_i[2]  & ~\new_[3067]_ );
  assign \new_[2896]_  = ~\new_[3058]_  | (~\wb_sel_i[3]  & ~\new_[3046]_ );
  assign \new_[2897]_  = ~\new_[2963]_  & (~\new_[3106]_  | ~\new_[386]_ );
  assign \new_[2898]_  = ~\new_[2997]_  & (~\new_[3120]_  | ~\new_[434]_ );
  assign \new_[2899]_  = ~\new_[2967]_  & (~\new_[3120]_  | ~\new_[436]_ );
  assign \new_[2900]_  = ~\new_[2983]_  & (~\new_[3120]_  | ~\new_[383]_ );
  assign \new_[2901]_  = ~\new_[2966]_  & (~\new_[3188]_  | ~\new_[382]_ );
  assign \new_[2902]_  = ~\new_[3093]_  | (~\wb_sel_i[3]  & ~\new_[3071]_ );
  assign \new_[2903]_  = ~\new_[3003]_  & (~\new_[3080]_  | ~\new_[354]_ );
  assign \new_[2904]_  = ~\new_[3129]_  | ~\wb_adr_i[4] ;
  assign \new_[2905]_  = ~\new_[2820]_  | ~\new_[3099]_ ;
  assign \new_[2906]_  = \new_[3332]_  & \new_[3012]_ ;
  assign \new_[2907]_  = ~\new_[3332]_  & ~\new_[3012]_ ;
  assign \new_[2908]_  = ~\new_[2960]_  & (~\new_[3188]_  | ~\new_[343]_ );
  assign \new_[2909]_  = ~\new_[2974]_  & (~\new_[3106]_  | ~\new_[385]_ );
  assign \new_[2910]_  = ~\new_[3004]_  & (~\new_[3106]_  | ~\new_[346]_ );
  assign \new_[2911]_  = ~\new_[3150]_  & ~\new_[3127]_ ;
  assign \new_[2912]_  = ~\new_[3012]_  | ~\new_[3014]_ ;
  assign \new_[2913]_  = ~\new_[2971]_  & (~\new_[3188]_  | ~\new_[427]_ );
  assign \new_[2914]_  = ~\new_[3036]_  & (~\new_[1935]_  | ~\new_[1930]_ );
  assign \new_[2915]_  = ~\new_[2952]_ ;
  assign \new_[2916]_  = ~\new_[2987]_  & (~\new_[3080]_  | ~\new_[392]_ );
  assign \new_[2917]_  = ~\new_[2985]_  & (~\new_[3080]_  | ~\new_[482]_ );
  assign \new_[2918]_  = ~\new_[3081]_  | ~\new_[3062]_  | ~\new_[3040]_ ;
  assign \new_[2919]_  = ~\new_[3052]_  | (~\wb_sel_i[1]  & ~\new_[3044]_ );
  assign \new_[2920]_  = wb_cyc_i & \new_[3145]_ ;
  assign \new_[2921]_  = ~\new_[2990]_  & (~\new_[3080]_  | ~\new_[503]_ );
  assign n1326 = ~\new_[3011]_  & ~wb_ack_o;
  assign \new_[2923]_  = ~\new_[2963]_  & (~\new_[3106]_  | ~\new_[429]_ );
  assign \new_[2924]_  = ~\new_[3112]_ ;
  assign \new_[2925]_  = ~\new_[3116]_  | ~\new_[3069]_  | ~\new_[3062]_ ;
  assign \new_[2926]_  = ~\new_[3107]_  | (~\wb_sel_i[0]  & ~\new_[3109]_ );
  assign \new_[2927]_  = ~\new_[2954]_ ;
  assign \new_[2928]_  = ~\new_[2989]_  & (~\new_[3120]_  | ~\new_[377]_ );
  assign \new_[2929]_  = ~\new_[3007]_  & (~\new_[3106]_  | ~\new_[380]_ );
  assign \new_[2930]_  = ~\new_[3004]_  & (~\new_[3106]_  | ~\new_[3158]_ );
  assign \new_[2931]_  = ~\new_[2968]_  & (~\new_[3106]_  | ~\new_[347]_ );
  assign \new_[2932]_  = ~\new_[3031]_  | (~\wb_sel_i[1]  & ~\new_[3077]_ );
  assign \new_[2933]_  = ~\new_[3244]_  | ~\new_[3112]_ ;
  assign \new_[2934]_  = ~\new_[3072]_  | (~\wb_sel_i[1]  & ~\new_[3104]_ );
  assign \new_[2935]_  = \new_[3245]_  | \new_[3057]_ ;
  assign \new_[2936]_  = ~\new_[3036]_  | ~\new_[3130]_ ;
  assign \new_[2937]_  = ~\new_[3244]_ ;
  assign \new_[2938]_  = \new_[3059]_  & \new_[3042]_ ;
  assign \new_[2939]_  = ~\wb_adr_i[2]  | ~\wb_adr_i[4] ;
  assign \new_[2940]_  = ~\new_[3451]_  & ~\new_[3068]_ ;
  assign \new_[2941]_  = ~\new_[3451]_  | ~\new_[3068]_ ;
  assign \new_[2942]_  = ~\new_[3188]_  | ~\new_[327]_ ;
  assign \new_[2943]_  = ~\new_[3106]_  | ~\new_[507]_ ;
  assign \new_[2944]_  = ~\new_[3188]_  | ~\new_[324]_ ;
  assign \new_[2945]_  = ~\new_[3106]_  | ~\new_[437]_ ;
  assign \new_[2946]_  = wb_stb_i & \wb_adr_i[2] ;
  assign \new_[2947]_  = ~\new_[1936]_  & ~\new_[1917]_ ;
  assign \new_[2948]_  = ~\new_[3106]_  | ~\new_[560]_ ;
  assign \new_[2949]_  = \new_[3036]_  | \new_[3130]_ ;
  assign \new_[2950]_  = \new_[1943]_  ^ \new_[1597]_ ;
  assign \new_[2951]_  = ~\new_[3189]_  & ~\new_[3103]_ ;
  assign \new_[2952]_  = ~\new_[3014]_ ;
  assign \new_[2953]_  = \new_[3048]_  & \new_[3053]_ ;
  assign \new_[2954]_  = \new_[3012]_ ;
  assign \new_[2955]_  = ~\wb_adr_i[3]  & ~\new_[3103]_ ;
  assign \new_[2956]_  = ~\new_[3012]_ ;
  assign \new_[2957]_  = ~\new_[3245]_  | ~\new_[3099]_ ;
  assign \new_[2958]_  = ~\new_[3120]_  | ~\new_[325]_ ;
  assign \new_[2959]_  = ~\new_[3042]_ ;
  assign \new_[2960]_  = ~\new_[3073]_ ;
  assign \new_[2961]_  = ~\new_[3120]_  | ~\new_[446]_ ;
  assign \new_[2962]_  = ~\new_[3107]_ ;
  assign \new_[2963]_  = ~\new_[3031]_ ;
  assign \new_[2964]_  = ~\new_[3051]_ ;
  assign \new_[2965]_  = ~\new_[3129]_  | ~\new_[3145]_ ;
  assign \new_[2966]_  = ~\new_[3098]_ ;
  assign \new_[2967]_  = ~\new_[3047]_ ;
  assign \new_[2968]_  = ~\new_[3056]_ ;
  assign \new_[2969]_  = ~\new_[3092]_ ;
  assign \new_[2970]_  = ~\new_[3490]_ ;
  assign \new_[2971]_  = ~\new_[3102]_ ;
  assign \new_[2972]_  = ~\new_[3106]_  | ~\new_[438]_ ;
  assign \new_[2973]_  = ~\new_[3120]_  | ~\new_[464]_ ;
  assign \new_[2974]_  = ~\new_[3060]_ ;
  assign \new_[2975]_  = ~\new_[3080]_  | ~\new_[562]_ ;
  assign \new_[2976]_  = ~\new_[3106]_  | ~\new_[561]_ ;
  assign \new_[2977]_  = ~\new_[3080]_  | ~\new_[528]_ ;
  assign \new_[2978]_  = ~\new_[3080]_  | ~\new_[440]_ ;
  assign \new_[2979]_  = ~\new_[3188]_  | ~\new_[509]_ ;
  assign \new_[2980]_  = ~\new_[3120]_  | ~\new_[441]_ ;
  assign \new_[2981]_  = ~\new_[3188]_  | ~\new_[505]_ ;
  assign \new_[2982]_  = ~\new_[3058]_ ;
  assign \new_[2983]_  = ~\new_[3091]_ ;
  assign \new_[2984]_  = ~\new_[3094]_ ;
  assign \new_[2985]_  = ~\new_[3105]_ ;
  assign \new_[2986]_  = ~\new_[3090]_ ;
  assign \new_[2987]_  = ~\new_[3083]_ ;
  assign \new_[2988]_  = ~\new_[3078]_ ;
  assign \new_[2989]_  = ~\new_[3087]_ ;
  assign \new_[2990]_  = ~\new_[3070]_ ;
  assign \new_[2991]_  = ~\new_[3088]_ ;
  assign \new_[2992]_  = ~\new_[3093]_ ;
  assign \new_[2993]_  = ~\new_[3120]_  | ~\new_[444]_ ;
  assign \new_[2994]_  = ~\new_[3188]_  | ~\new_[557]_ ;
  assign \new_[2995]_  = ~\new_[3043]_ ;
  assign \new_[2996]_  = ~\new_[3097]_ ;
  assign \new_[2997]_  = ~\new_[3108]_ ;
  assign \new_[2998]_  = ~\new_[3106]_  | ~\new_[559]_ ;
  assign \new_[2999]_  = ~\new_[3188]_  | ~\new_[506]_ ;
  assign \new_[3000]_  = \new_[3129]_  | \wb_adr_i[4] ;
  assign \new_[3001]_  = ~\new_[3072]_ ;
  assign \new_[3002]_  = ~\new_[3052]_ ;
  assign \new_[3003]_  = ~\new_[3038]_ ;
  assign \new_[3004]_  = ~\new_[3054]_ ;
  assign \new_[3005]_  = ~\new_[3120]_  | ~\new_[492]_ ;
  assign \new_[3006]_  = ~\new_[3080]_  | ~\new_[498]_ ;
  assign \new_[3007]_  = ~\new_[3034]_ ;
  assign \new_[3008]_  = ~\new_[3041]_ ;
  assign \new_[3009]_  = wb_stb_i & \new_[3129]_ ;
  assign \new_[3010]_  = ~\new_[3055]_ ;
  assign \new_[3011]_  = ~\new_[3033]_ ;
  assign \new_[3012]_  = ~\new_[3068]_ ;
  assign \new_[3013]_  = ~\new_[3106]_  | ~\new_[495]_ ;
  assign \new_[3014]_  = ~\new_[3099]_ ;
  assign \new_[3015]_  = ~\new_[3120]_  | ~\new_[443]_ ;
  assign \new_[3016]_  = ~\new_[3188]_  | ~\new_[465]_ ;
  assign \new_[3017]_  = ~\new_[3106]_  | ~\new_[493]_ ;
  assign \new_[3018]_  = ~\new_[3075]_ ;
  assign \new_[3019]_  = ~\new_[3177]_  & ~\wb_adr_i[4] ;
  assign \new_[3020]_  = ~\new_[3080]_  | ~\new_[439]_ ;
  assign \new_[3021]_  = ~\new_[3080]_  | ~\new_[524]_ ;
  assign \new_[3022]_  = ~\new_[3189]_  & ~\new_[1658]_ ;
  assign \new_[3023]_  = ~\new_[3080]_  | ~\new_[494]_ ;
  assign \new_[3024]_  = ~\new_[3188]_  | ~\new_[558]_ ;
  assign \new_[3025]_  = ~\new_[3188]_  | ~\new_[442]_ ;
  assign \new_[3026]_  = ~\new_[3080]_  | ~\new_[468]_ ;
  assign \new_[3027]_  = ~\new_[3188]_  | ~\new_[508]_ ;
  assign \new_[3028]_  = ~\new_[3120]_  | ~\new_[447]_ ;
  assign \new_[3029]_  = ~\new_[3120]_  | ~\new_[445]_ ;
  assign \new_[3030]_  = ~\new_[337]_ ;
  assign \new_[3031]_  = ~\wb_dat_i[13]  | ~\wb_sel_i[1] ;
  assign \new_[3032]_  = ~\new_[1597]_  & ~\new_[1580]_ ;
  assign \new_[3033]_  = wb_stb_i & wb_cyc_i;
  assign \new_[3034]_  = ~\wb_dat_i[10]  | ~\wb_sel_i[1] ;
  assign \new_[3035]_  = ~\new_[367]_ ;
  assign \new_[3036]_  = ~\new_[1935]_  & ~\new_[1930]_ ;
  assign \new_[3037]_  = ~\new_[368]_ ;
  assign \new_[3038]_  = ~\wb_dat_i[23]  | ~\wb_sel_i[2] ;
  assign \new_[3039]_  = ~\new_[1938]_  & ~\new_[1891]_ ;
  assign \new_[3040]_  = ~\new_[1854]_  & ~\new_[1583]_ ;
  assign \new_[3041]_  = ~\wb_dat_i[17]  | ~\wb_sel_i[2] ;
  assign \new_[3042]_  = ~\new_[1932]_  & ~\new_[1933]_ ;
  assign \new_[3043]_  = ~\wb_dat_i[19]  | ~\wb_sel_i[2] ;
  assign \new_[3044]_  = ~\new_[333]_ ;
  assign \new_[3045]_  = ~\new_[341]_ ;
  assign \new_[3046]_  = ~\new_[370]_ ;
  assign \new_[3047]_  = ~\wb_dat_i[30]  | ~\wb_sel_i[3] ;
  assign \new_[3048]_  = ~\new_[1934]_  & ~\new_[2076]_ ;
  assign \new_[3049]_  = ~\new_[1934]_  & ~\new_[1892]_ ;
  assign \new_[3050]_  = ~\new_[366]_ ;
  assign \new_[3051]_  = ~\wb_dat_i[0]  | ~\wb_sel_i[0] ;
  assign \new_[3052]_  = ~\wb_dat_i[11]  | ~\wb_sel_i[1] ;
  assign \new_[3053]_  = ~\new_[1692]_  & ~\new_[1922]_ ;
  assign \new_[3054]_  = ~\wb_dat_i[8]  | ~\wb_sel_i[1] ;
  assign \new_[3055]_  = ~\wb_dat_i[22]  | ~\wb_sel_i[2] ;
  assign \new_[3056]_  = ~\wb_dat_i[14]  | ~\wb_sel_i[1] ;
  assign \new_[3057]_  = ~\new_[3246]_ ;
  assign \new_[3058]_  = ~\wb_dat_i[26]  | ~\wb_sel_i[3] ;
  assign \new_[3059]_  = ~\new_[1929]_  & ~\new_[2004]_ ;
  assign \new_[3060]_  = ~\wb_dat_i[12]  | ~\wb_sel_i[1] ;
  assign \new_[3061]_  = ~\new_[3150]_ ;
  assign \new_[3062]_  = ~\new_[1927]_  & ~\new_[1931]_ ;
  assign \new_[3063]_  = ~\new_[1923]_  & ~\new_[1950]_ ;
  assign \new_[3064]_  = ~\new_[1948]_  & ~\new_[1949]_ ;
  assign \new_[3065]_  = ~\new_[369]_ ;
  assign \new_[3066]_  = ~\new_[1940]_  & ~\new_[1946]_ ;
  assign \new_[3067]_  = ~\new_[336]_ ;
  assign \new_[3068]_  = ~\new_[3245]_ ;
  assign \new_[3069]_  = ~\new_[2004]_  & ~\new_[1930]_ ;
  assign \new_[3070]_  = ~\wb_dat_i[20]  | ~\wb_sel_i[2] ;
  assign \new_[3071]_  = ~\new_[339]_ ;
  assign \new_[3072]_  = ~\wb_dat_i[9]  | ~\wb_sel_i[1] ;
  assign \new_[3073]_  = ~\wb_dat_i[2]  | ~\wb_sel_i[0] ;
  assign \new_[3074]_  = ~\new_[1690]_ ;
  assign \new_[3075]_  = ~\wb_dat_i[1]  | ~\wb_sel_i[0] ;
  assign \new_[3076]_  = ~\new_[1944]_  & ~\new_[1939]_ ;
  assign \new_[3077]_  = ~\new_[363]_ ;
  assign \new_[3078]_  = ~\wb_dat_i[31]  | ~\wb_sel_i[3] ;
  assign \new_[3079]_  = ~\new_[358]_ ;
  assign \new_[3080]_  = ~\wb_sel_i[2] ;
  assign \new_[3081]_  = ~\new_[1892]_  & ~\new_[1859]_ ;
  assign \new_[3082]_  = ~\wb_adr_i[3]  & ~\wb_adr_i[4] ;
  assign \new_[3083]_  = ~\wb_dat_i[21]  | ~\wb_sel_i[2] ;
  assign \new_[3084]_  = ~\new_[349]_ ;
  assign \new_[3085]_  = ~\new_[1945]_  & ~\new_[1918]_ ;
  assign \new_[3086]_  = ~\new_[328]_ ;
  assign \new_[3087]_  = ~\wb_dat_i[28]  | ~\wb_sel_i[3] ;
  assign \new_[3088]_  = ~\wb_dat_i[24]  | ~\wb_sel_i[3] ;
  assign \new_[3089]_  = ~\new_[359]_ ;
  assign \new_[3090]_  = ~\wb_dat_i[15]  | ~\wb_sel_i[1] ;
  assign \new_[3091]_  = ~\wb_dat_i[25]  | ~\wb_sel_i[3] ;
  assign \new_[3092]_  = ~\wb_dat_i[18]  | ~\wb_sel_i[2] ;
  assign \new_[3093]_  = ~\wb_dat_i[29]  | ~\wb_sel_i[3] ;
  assign \new_[3094]_  = ~\wb_dat_i[3]  | ~\wb_sel_i[0] ;
  assign \new_[3095]_  = ~\new_[1943]_ ;
  assign \new_[3096]_  = ~\new_[335]_ ;
  assign \new_[3097]_  = ~\wb_dat_i[7]  | ~\wb_sel_i[0] ;
  assign \new_[3098]_  = ~\wb_dat_i[5]  | ~\wb_sel_i[0] ;
  assign \new_[3099]_  = ~\new_[3246]_ ;
  assign \new_[3100]_  = ~\new_[3319]_ ;
  assign \new_[3101]_  = ~\new_[1916]_  & ~\new_[1947]_ ;
  assign \new_[3102]_  = ~\wb_dat_i[4]  | ~\wb_sel_i[0] ;
  assign \new_[3103]_  = \wb_adr_i[2]  | \wb_adr_i[4] ;
  assign \new_[3104]_  = ~\new_[362]_ ;
  assign \new_[3105]_  = ~\wb_dat_i[16]  | ~\wb_sel_i[2] ;
  assign \new_[3106]_  = ~\wb_sel_i[1] ;
  assign \new_[3107]_  = ~\wb_dat_i[6]  | ~\wb_sel_i[0] ;
  assign \new_[3108]_  = ~\wb_dat_i[27]  | ~\wb_sel_i[3] ;
  assign \new_[3109]_  = ~\new_[360]_ ;
  assign \new_[3110]_  = ~\new_[1937]_  & ~\new_[1928]_ ;
  assign \new_[3111]_  = ~\new_[371]_ ;
  assign \new_[3112]_  = ~\new_[3127]_ ;
  assign \new_[3113]_  = ~\new_[346]_ ;
  assign \new_[3114]_  = ~\new_[501]_ ;
  assign \new_[3115]_  = ~\new_[357]_ ;
  assign \new_[3116]_  = ~\new_[1935]_ ;
  assign \new_[3117]_  = ~\new_[444]_ ;
  assign \new_[3118]_  = ~\new_[437]_ ;
  assign \new_[3119]_  = ~\new_[1862]_ ;
  assign \new_[3120]_  = ~\wb_sel_i[3] ;
  assign \new_[3121]_  = ~sclk_pad_o;
  assign \new_[3122]_  = ~\new_[1860]_ ;
  assign \new_[3123]_  = ~\new_[331]_ ;
  assign \new_[3124]_  = ~\new_[1941]_ ;
  assign \new_[3125]_  = ~\new_[509]_ ;
  assign \new_[3127]_  = ~\new_[1856]_ ;
  assign \new_[3128]_  = ~\new_[497]_ ;
  assign \new_[3129]_  = ~\wb_adr_i[2] ;
  assign \new_[3130]_  = ~\new_[1931]_ ;
  assign \new_[3131]_  = ~\new_[332]_ ;
  assign \new_[3132]_  = ~\new_[390]_ ;
  assign \new_[3133]_  = ~\new_[474]_ ;
  assign \new_[3134]_  = ~\new_[528]_ ;
  assign \new_[3135]_  = ~\new_[2138]_ ;
  assign \new_[3136]_  = ~\new_[2135]_ ;
  assign \new_[3137]_  = ~\new_[1789]_ ;
  assign \new_[3138]_  = ~\new_[348]_ ;
  assign \new_[3139]_  = ~\new_[352]_ ;
  assign \new_[3140]_  = ~\new_[1917]_ ;
  assign \new_[3141]_  = ~\new_[2109]_ ;
  assign \new_[3142]_  = ~\new_[424]_ ;
  assign \new_[3143]_  = ~\new_[1665]_ ;
  assign \new_[3144]_  = ~\new_[500]_ ;
  assign \new_[3145]_  = ~\new_[1658]_ ;
  assign \new_[3146]_  = ~\new_[342]_ ;
  assign \new_[3147]_  = ~\new_[355]_ ;
  assign \new_[3148]_  = ~\new_[2126]_ ;
  assign \new_[3149]_  = ~\new_[1941]_ ;
  assign \new_[3150]_  = ~\new_[1693]_ ;
  assign \new_[3151]_  = ~\new_[2136]_ ;
  assign \new_[3152]_  = ~\new_[347]_ ;
  assign \new_[3153]_  = ~\new_[488]_ ;
  assign \new_[3154]_  = ~\new_[356]_ ;
  assign \new_[3155]_  = ~\new_[560]_ ;
  assign \new_[3156]_  = ~\new_[372]_ ;
  assign \new_[3157]_  = ~\new_[338]_ ;
  assign \new_[3158]_  = ~\new_[1581]_ ;
  assign \new_[3159]_  = ~\new_[1861]_ ;
  assign \new_[3160]_  = ~\new_[499]_ ;
  assign \new_[3161]_  = ~\new_[364]_ ;
  assign \new_[3162]_  = ~\new_[340]_ ;
  assign \new_[3163]_  = ~\new_[329]_ ;
  assign \new_[3164]_  = ~\new_[334]_ ;
  assign \new_[3165]_  = ~\new_[2137]_ ;
  assign \new_[3166]_  = ~\new_[427]_ ;
  assign \new_[3167]_  = ~\new_[438]_ ;
  assign \new_[3168]_  = ~\new_[361]_ ;
  assign \new_[3169]_  = ~\new_[482]_ ;
  assign \new_[3170]_  = ~\new_[1922]_ ;
  assign \new_[3171]_  = ~wb_int_o;
  assign \new_[3172]_  = ~\new_[2139]_ ;
  assign \new_[3173]_  = ~\new_[1919]_ ;
  assign \new_[3174]_  = ~\new_[330]_ ;
  assign \new_[3175]_  = ~\new_[1926]_ ;
  assign \new_[3176]_  = ~\new_[343]_ ;
  assign \new_[3177]_  = ~wb_cyc_i;
  assign \new_[3178]_  = ~\new_[558]_ ;
  assign \new_[3179]_  = ~\new_[496]_ ;
  assign \new_[3180]_  = ~\new_[439]_ ;
  assign \new_[3181]_  = ~\new_[508]_ ;
  assign \new_[3182]_  = ~\new_[506]_ ;
  assign \new_[3183]_  = ~\new_[428]_ ;
  assign \new_[3184]_  = ~\new_[374]_ ;
  assign \new_[3185]_  = ~\new_[503]_ ;
  assign \new_[3186]_  = ~\new_[326]_ ;
  assign \new_[3187]_  = ~\new_[375]_ ;
  assign \new_[3188]_  = ~\wb_sel_i[0] ;
  assign \new_[3189]_  = ~\wb_adr_i[3] ;
  assign \new_[3190]_  = ~\new_[1942]_ ;
  assign \new_[3191]_  = ~\new_[435]_ ;
  assign \new_[3192]_  = ~\new_[507]_ ;
  assign \new_[3193]_  = ~\new_[2124]_ ;
  assign \new_[3194]_  = ~\new_[486]_ ;
  assign \new_[3195]_  = ~\new_[354]_ ;
  assign \new_[3196]_  = ~\new_[1933]_ ;
  assign \new_[3197]_  = ~\new_[426]_ ;
  assign \new_[3198]_  = ~\new_[365]_ ;
  assign \new_[3199]_  = ~\new_[344]_ ;
  assign \new_[3200]_  = ~\new_[502]_ ;
  assign \new_[3201]_  = ~\new_[3393]_  | ~\new_[3248]_ ;
  assign \new_[3202]_  = ~\new_[3203]_  & ~\new_[1438]_ ;
  assign \new_[3203]_  = ~\new_[3422]_ ;
  assign \new_[3204]_  = \new_[3203]_  & miso_pad_i;
  assign \new_[3205]_  = ~\new_[3412]_  & ~\new_[3206]_ ;
  assign \new_[3206]_  = ~\new_[3207]_  | ~\new_[3208]_ ;
  assign \new_[3207]_  = \new_[1447]_  & \new_[3543]_ ;
  assign \new_[3208]_  = ~\new_[3532]_ ;
  assign \new_[3209]_  = ~\new_[3208]_ ;
  assign \new_[3210]_  = ~\new_[3218]_  | (~\new_[3211]_  & ~\new_[3215]_ );
  assign \new_[3211]_  = ~\new_[3214]_  & (~\new_[3212]_  | ~\new_[3213]_ );
  assign \new_[3212]_  = ~\new_[1030]_ ;
  assign \new_[3213]_  = ~\new_[464]_  | ~\new_[1095]_ ;
  assign \new_[3214]_  = \new_[3424]_ ;
  assign \new_[3215]_  = \new_[3216]_  & \new_[3217]_ ;
  assign \new_[3216]_  = ~\new_[2667]_ ;
  assign \new_[3217]_  = ~\new_[2973]_  | ~\new_[3087]_ ;
  assign \new_[3218]_  = ~\new_[3500]_ ;
  assign \new_[3219]_  = ~\new_[3214]_ ;
  assign \new_[3220]_  = ~\new_[3221]_  | ~\new_[3223]_ ;
  assign \new_[3221]_  = ~\new_[3222]_  | ~\new_[1317]_  | ~\new_[1088]_  | ~\new_[1390]_ ;
  assign \new_[3222]_  = ~wb_we_i | ~\new_[3019]_  | ~\new_[3022]_  | ~\new_[2946]_ ;
  assign \new_[3223]_  = ~\new_[360]_  | ~\new_[3224]_  | ~\new_[3222]_ ;
  assign \new_[3224]_  = ~\new_[1390]_  | ~\new_[1317]_ ;
  assign \new_[3225]_  = ~\new_[3222]_ ;
  assign \new_[3226]_  = ~\new_[3310]_  | ~\new_[3227]_  | ~\new_[3231]_ ;
  assign \new_[3227]_  = ~\new_[3228]_  | ~\new_[3229]_ ;
  assign \new_[3228]_  = ~\new_[1010]_ ;
  assign \new_[3229]_  = ~\new_[3230]_  & (~\new_[505]_  | ~\new_[1250]_ );
  assign \new_[3230]_  = ~\new_[2667]_  & (~\new_[2981]_  | ~\new_[3097]_ );
  assign \new_[3231]_  = \new_[3230]_  | \new_[3349]_ ;
  assign \new_[3232]_  = ~\new_[3233]_  & ~\new_[3237]_ ;
  assign \new_[3233]_  = ~\new_[3277]_  | ~\new_[3234]_ ;
  assign \new_[3234]_  = ~\new_[3235]_ ;
  assign \new_[3235]_  = ~\new_[3548]_ ;
  assign \new_[3236]_  = ~\new_[1969]_  | ~\new_[3459]_ ;
  assign \new_[3237]_  = ~\new_[1482]_  | ~\new_[3315]_  | ~\new_[3412]_ ;
  assign \new_[3238]_  = ~\new_[3496]_  | ~\new_[3239]_  | ~\new_[3243]_ ;
  assign \new_[3239]_  = ~\new_[3240]_  | ~\new_[3241]_ ;
  assign \new_[3240]_  = ~\new_[3430]_  | ~\new_[1265]_ ;
  assign \new_[3241]_  = ~\new_[3242]_  & (~\new_[1330]_  | ~\new_[558]_ );
  assign \new_[3242]_  = ~\new_[2667]_  & (~\new_[3024]_  | ~\new_[3107]_ );
  assign \new_[3243]_  = \new_[3349]_  | \new_[3242]_ ;
  assign \new_[3244]_  = ~\new_[3245]_  & ~\new_[3246]_ ;
  assign \new_[3245]_  = ~\new_[2032]_ ;
  assign \new_[3246]_  = ~\new_[2029]_ ;
  assign \new_[3247]_  = ~\new_[1699]_  | ~\new_[1429]_  | ~\new_[1477]_ ;
  assign \new_[3248]_  = ~\new_[3538]_  | ~\new_[3249]_  | ~\new_[3250]_ ;
  assign \new_[3249]_  = ~\new_[3397]_  | ~\new_[1468]_  | ~\new_[1469]_ ;
  assign \new_[3250]_  = ~\new_[3507]_  | ~\new_[3251]_  | ~\new_[3252]_ ;
  assign \new_[3251]_  = ~\new_[3445]_  | (~\new_[1491]_  & ~\new_[1499]_ );
  assign \new_[3252]_  = ~\new_[3544]_  | (~\new_[1498]_  & ~\new_[1490]_ );
  assign \new_[3253]_  = ~\new_[3257]_  & (~\new_[3254]_  | ~\new_[562]_ );
  assign \new_[3254]_  = \new_[3255]_  | \new_[3256]_ ;
  assign \new_[3255]_  = \new_[1459]_  | \new_[1424]_ ;
  assign \new_[3256]_  = ~\new_[1593]_  | ~\new_[1429]_  | ~\new_[1476]_ ;
  assign \new_[3257]_  = ~\new_[3254]_  & ~\new_[1066]_ ;
  assign \new_[3258]_  = \new_[1459]_  | \new_[1424]_ ;
  assign \new_[3259]_  = ~\new_[3430]_  | ~\new_[1264]_ ;
  assign \new_[3260]_  = ~\new_[3261]_  & (~\new_[1329]_  | ~\new_[557]_ );
  assign \new_[3261]_  = ~\new_[2667]_  & (~\new_[2994]_  | ~\new_[3098]_ );
  assign \new_[3262]_  = ~\new_[3523]_  | ~\new_[3417]_ ;
  assign \new_[3263]_  = ~\new_[3419]_ ;
  assign \new_[3264]_  = ~\new_[3496]_  | ~\new_[3265]_  | ~\new_[3269]_ ;
  assign \new_[3265]_  = ~\new_[3266]_  | ~\new_[3267]_ ;
  assign \new_[3266]_  = ~\new_[3430]_  | ~\new_[1171]_ ;
  assign \new_[3267]_  = ~\new_[3268]_  & (~\new_[528]_  | ~\new_[1237]_ );
  assign \new_[3268]_  = ~\new_[2667]_  & (~\new_[2977]_  | ~\new_[3043]_ );
  assign \new_[3269]_  = \new_[3268]_  | \new_[3349]_ ;
  assign \new_[3270]_  = ~\new_[3401]_  | ~\new_[3271]_  | ~\new_[3273]_ ;
  assign \new_[3271]_  = \new_[3272]_ ;
  assign \new_[3272]_  = \new_[3208]_  & \new_[1452]_ ;
  assign \new_[3273]_  = ~\new_[1472]_  & ~\new_[3276]_ ;
  assign \new_[3274]_  = \new_[3275]_ ;
  assign \new_[3275]_  = ~\new_[3353]_ ;
  assign \new_[3276]_  = ~\new_[3277]_ ;
  assign \new_[3277]_  = \new_[3546]_ ;
  assign \new_[3278]_  = ~\new_[3279]_ ;
  assign \new_[3279]_  = ~\new_[3282]_  & (~\new_[3280]_  | ~\new_[3281]_ );
  assign \new_[3280]_  = ~\new_[3298]_  | ~\new_[1118]_  | ~\new_[1016]_ ;
  assign \new_[3281]_  = ~\new_[380]_  | (~\new_[2377]_  & ~\new_[3292]_ );
  assign \new_[3282]_  = ~\new_[3283]_  | ~\new_[3312]_ ;
  assign \new_[3283]_  = ~\new_[3284]_  | ~\new_[3292]_ ;
  assign \new_[3284]_  = ~\new_[3292]_  | ~\new_[380]_ ;
  assign \new_[3285]_  = ~\new_[3286]_ ;
  assign \new_[3286]_  = ~\new_[3289]_  & (~\new_[3287]_  | ~\new_[3288]_ );
  assign \new_[3287]_  = ~\new_[3298]_  | ~\new_[1120]_  | ~\new_[1031]_ ;
  assign \new_[3288]_  = ~\new_[385]_  | (~\new_[2377]_  & ~\new_[3292]_ );
  assign \new_[3289]_  = ~\new_[3290]_  | ~\new_[3312]_ ;
  assign \new_[3290]_  = ~\new_[3291]_  | ~\new_[3292]_ ;
  assign \new_[3291]_  = ~\new_[3292]_  | ~\new_[385]_ ;
  assign \new_[3292]_  = ~\new_[3293]_ ;
  assign \new_[3293]_  = ~\wb_adr_i[2]  | ~\new_[2783]_  | ~\new_[3145]_ ;
  assign \new_[3294]_  = ~\new_[3298]_  | ~\new_[3295]_  | ~\new_[3297]_ ;
  assign \new_[3295]_  = ~\new_[1066]_  | ~\new_[3296]_ ;
  assign \new_[3296]_  = \new_[1314]_  & \new_[1382]_ ;
  assign \new_[3297]_  = \new_[388]_  | \new_[3296]_ ;
  assign \new_[3298]_  = \new_[3349]_ ;
  assign \new_[3299]_  = ~\new_[3301]_  & (~\new_[3300]_  | ~\new_[524]_ );
  assign \new_[3300]_  = \new_[3247]_  | \new_[3258]_ ;
  assign \new_[3301]_  = ~\new_[1066]_  & ~\new_[3300]_ ;
  assign n756 = ~\new_[3303]_  | ~\new_[3307]_ ;
  assign \new_[3303]_  = ~\new_[3304]_  | (~\new_[952]_  & ~\new_[2249]_ );
  assign \new_[3304]_  = ~\new_[3500]_  & (~\new_[2249]_  | ~\new_[3305]_ );
  assign \new_[3305]_  = ~\new_[504]_ ;
  assign \new_[3306]_  = ~\new_[2843]_  & ~\new_[2965]_ ;
  assign \new_[3307]_  = ~\new_[3309]_  & (~\new_[3308]_  | ~\new_[504]_ );
  assign \new_[3308]_  = \new_[3306]_ ;
  assign \new_[3309]_  = ~\new_[2844]_  & ~\new_[2553]_ ;
  assign \new_[3310]_  = ~\new_[3500]_ ;
  assign \new_[3311]_  = \new_[3308]_ ;
  assign \new_[3312]_  = ~\new_[3308]_ ;
  assign \new_[3313]_  = ~\new_[3314]_  & ~\new_[3550]_ ;
  assign \new_[3314]_  = ~\new_[1467]_  | ~\new_[3532]_ ;
  assign \new_[3315]_  = ~\new_[3314]_ ;
  assign \new_[3316]_  = ~\new_[3317]_ ;
  assign \new_[3317]_  = ~\new_[3318]_  | ~\new_[3319]_ ;
  assign \new_[3318]_  = ~\new_[2691]_  | ~\new_[2905]_ ;
  assign \new_[3319]_  = ~\new_[1936]_ ;
  assign \new_[3320]_  = ~\new_[3321]_ ;
  assign \new_[3321]_  = \new_[3317]_ ;
  assign \new_[3322]_  = ~\new_[1694]_  | ~\new_[3262]_  | ~\new_[3263]_ ;
  assign \new_[3323]_  = \new_[2209]_  | \new_[3324]_ ;
  assign \new_[3324]_  = \new_[1694]_  | \new_[2493]_ ;
  assign \new_[3325]_  = ~\new_[3342]_  | ~\new_[3326]_  | ~\new_[2210]_ ;
  assign \new_[3326]_  = \new_[3528]_ ;
  assign \new_[3327]_  = ~\new_[3342]_ ;
  assign \new_[3328]_  = \new_[3095]_  ? \new_[3329]_  : \new_[1943]_ ;
  assign \new_[3329]_  = (~\new_[3436]_  & ~\new_[1597]_ ) | (~\new_[3330]_  & ~\new_[3331]_ );
  assign \new_[3330]_  = ~\new_[2592]_  | (~\new_[2681]_  & ~\new_[1597]_ );
  assign \new_[3331]_  = ~\new_[3436]_ ;
  assign \new_[3332]_  = ~\new_[3436]_ ;
  assign \new_[3333]_  = ~\new_[3477]_  & (~\new_[3334]_  | ~\new_[3335]_ );
  assign \new_[3334]_  = ~\new_[1638]_  | ~\new_[3411]_ ;
  assign \new_[3335]_  = ~\new_[1639]_  | ~\new_[1617]_ ;
  assign \new_[3336]_  = ~\new_[3508]_  | ~\new_[3342]_ ;
  assign \new_[3337]_  = ~\new_[2306]_  | ~\new_[3490]_ ;
  assign \new_[3338]_  = \new_[3339]_  | \new_[3325]_ ;
  assign \new_[3339]_  = ~\new_[2026]_  | ~\new_[1925]_ ;
  assign \new_[3340]_  = ~\new_[3342]_  | ~\new_[3341]_  | ~\new_[3339]_ ;
  assign \new_[3341]_  = ~\new_[2210]_  | ~\new_[3326]_ ;
  assign \new_[3342]_  = \new_[1694]_ ;
  assign \new_[3343]_  = ~\new_[2133]_  | ~\new_[3327]_ ;
  assign \new_[3344]_  = ~\new_[3350]_  | (~\new_[3345]_  & ~\new_[3346]_ );
  assign \new_[3345]_  = \new_[1068]_ ;
  assign \new_[3346]_  = ~\new_[3349]_  | ~\new_[3347]_  | ~\new_[3348]_ ;
  assign \new_[3347]_  = \new_[1367]_ ;
  assign \new_[3348]_  = \new_[1451]_  & \new_[3406]_ ;
  assign \new_[3349]_  = ~\new_[3424]_ ;
  assign \new_[3350]_  = ~\new_[492]_  | ~\new_[3351]_  | ~\new_[3349]_ ;
  assign \new_[3351]_  = ~\new_[3347]_  | ~\new_[3348]_ ;
  assign \new_[3352]_  = \new_[3336]_ ;
  assign \new_[3353]_  = ~\new_[3352]_  | ~\new_[3337]_ ;
  assign \new_[3354]_  = ~\new_[3357]_  & (~\new_[3355]_  | ~\new_[3356]_ );
  assign \new_[3355]_  = ~\new_[3472]_  | ~\new_[1636]_ ;
  assign \new_[3356]_  = ~\new_[1635]_  | ~\new_[3411]_ ;
  assign \new_[3357]_  = \new_[3352]_  & \new_[3337]_ ;
  assign \new_[3358]_  = ~\new_[3522]_  & (~\new_[1532]_  | ~\new_[1566]_ );
  assign \new_[3359]_  = ~\new_[3366]_  | (~\new_[3360]_  & ~\new_[3364]_ );
  assign \new_[3360]_  = ~\new_[3361]_  & ~\new_[3363]_ ;
  assign \new_[3361]_  = ~\new_[3362]_  | (~\new_[1195]_  & ~\new_[2596]_ );
  assign \new_[3362]_  = \new_[3186]_  | \new_[3222]_ ;
  assign \new_[3363]_  = ~\new_[2596]_  & ~\new_[1045]_ ;
  assign \new_[3364]_  = \new_[3365]_ ;
  assign \new_[3365]_  = ~\new_[2857]_  & ~\new_[2859]_ ;
  assign \new_[3366]_  = ~\new_[3364]_  | ~\new_[326]_ ;
  assign \new_[3367]_  = ~\new_[3365]_ ;
  assign \new_[3368]_  = ~\new_[3406]_  | ~\new_[344]_ ;
  assign \new_[3369]_  = ~\new_[2907]_  & ~\new_[2906]_ ;
  assign \new_[3370]_  = ~\new_[3489]_  | (~\new_[3371]_  & ~\new_[2683]_ );
  assign \new_[3371]_  = ~\new_[3372]_ ;
  assign \new_[3372]_  = ~\new_[2665]_ ;
  assign \new_[3373]_  = \new_[3374]_ ;
  assign \new_[3374]_  = ~\new_[3375]_  | ~\new_[3378]_ ;
  assign \new_[3375]_  = ~\new_[3372]_  | ~\new_[3376]_ ;
  assign \new_[3376]_  = ~\new_[3377]_  & ~\new_[2683]_ ;
  assign \new_[3377]_  = ~\new_[1694]_ ;
  assign \new_[3378]_  = ~\new_[3379]_  | ~\new_[3380]_ ;
  assign \new_[3379]_  = ~\new_[2906]_ ;
  assign \new_[3380]_  = ~\new_[1694]_  & ~\new_[2907]_ ;
  assign \new_[3381]_  = \new_[3382]_  ? \new_[1694]_  : \new_[3384]_ ;
  assign \new_[3382]_  = ~\new_[3383]_ ;
  assign \new_[3383]_  = ~\new_[2912]_  | ~\new_[2815]_ ;
  assign \new_[3384]_  = ~\new_[3387]_  & (~\new_[3385]_  | ~\new_[3386]_ );
  assign \new_[3385]_  = ~\new_[2824]_  & ~\new_[2771]_ ;
  assign \new_[3386]_  = ~\new_[1860]_  & ~\new_[2954]_ ;
  assign \new_[3387]_  = ~\new_[3388]_  & ~\new_[3385]_ ;
  assign \new_[3388]_  = ~\new_[1860]_  & ~\new_[2954]_ ;
  assign \new_[3389]_  = ~\new_[3440]_  & (~\new_[3390]_  | ~\new_[3391]_ );
  assign \new_[3390]_  = ~\new_[1685]_  | ~\new_[3410]_ ;
  assign \new_[3391]_  = ~\new_[1619]_  | ~\new_[1686]_ ;
  assign \new_[3392]_  = ~\new_[3353]_  & (~\new_[1590]_  | ~\new_[1536]_ );
  assign \new_[3393]_  = ~\new_[3537]_  | ~\new_[3394]_  | ~\new_[3398]_ ;
  assign \new_[3394]_  = ~\new_[3397]_  | ~\new_[3395]_  | ~\new_[3396]_ ;
  assign \new_[3395]_  = ~\new_[3445]_  | (~\new_[3358]_  & ~\new_[3354]_ );
  assign \new_[3396]_  = ~\new_[3520]_  | (~\new_[1500]_  & ~\new_[3333]_ );
  assign \new_[3397]_  = ~\new_[3507]_ ;
  assign \new_[3398]_  = ~\new_[3507]_  | ~\new_[3399]_  | ~\new_[3400]_ ;
  assign \new_[3399]_  = ~\new_[3544]_  | (~\new_[3389]_  & ~\new_[3392]_ );
  assign \new_[3400]_  = ~\new_[3445]_  | (~\new_[1501]_  & ~\new_[1492]_ );
  assign \new_[3401]_  = ~\new_[3402]_  & ~\new_[3413]_ ;
  assign \new_[3402]_  = \new_[3403]_ ;
  assign \new_[3403]_  = ~\new_[3370]_  | (~\new_[3369]_  & ~\new_[3489]_ );
  assign \new_[3404]_  = ~\new_[3482]_  | ~\new_[3405]_ ;
  assign \new_[3405]_  = ~\new_[2528]_  | ~\new_[3490]_ ;
  assign \new_[3406]_  = ~\new_[3402]_ ;
  assign \new_[3407]_  = ~\new_[3140]_  | ~\new_[2516]_ ;
  assign \new_[3408]_  = ~\new_[2651]_  | ~\new_[3409]_ ;
  assign \new_[3409]_  = ~\new_[3140]_  & ~\new_[2770]_ ;
  assign \new_[3410]_  = \new_[3404]_ ;
  assign \new_[3411]_  = ~\new_[3415]_ ;
  assign \new_[3412]_  = \new_[3413]_ ;
  assign \new_[3413]_  = \new_[3414]_ ;
  assign \new_[3414]_  = ~\new_[3415]_ ;
  assign \new_[3415]_  = ~\new_[3404]_ ;
  assign \new_[3416]_  = ~\new_[3418]_  | ~\new_[3417]_  | ~\new_[3523]_ ;
  assign \new_[3417]_  = ~\new_[2131]_  & (~\new_[2141]_  | ~\new_[3528]_ );
  assign \new_[3418]_  = \new_[3419]_  & \new_[1694]_ ;
  assign \new_[3419]_  = ~\new_[2037]_  | ~\new_[2140]_ ;
  assign \new_[3420]_  = ~\new_[3204]_  & (~\new_[3201]_  | ~\new_[3202]_ );
  assign \new_[3421]_  = ~\new_[3422]_  | ~\new_[3533]_  | ~\new_[3549]_ ;
  assign \new_[3422]_  = ~\new_[1672]_  | ~\new_[2047]_  | ~\new_[1921]_ ;
  assign \new_[3423]_  = ~\new_[3424]_  & ~\new_[3425]_ ;
  assign \new_[3424]_  = \new_[3365]_  | \new_[3225]_ ;
  assign \new_[3425]_  = ~\new_[3427]_  & (~\new_[3426]_  | ~\new_[559]_ );
  assign \new_[3426]_  = \new_[1413]_  | \new_[1355]_ ;
  assign \new_[3427]_  = ~\new_[1066]_  & ~\new_[3426]_ ;
  assign \new_[3428]_  = \new_[3429]_ ;
  assign \new_[3429]_  = ~\new_[3420]_  | ~\new_[3421]_ ;
  assign \new_[3430]_  = ~\new_[1066]_ ;
  assign \new_[3431]_  = ~\new_[3477]_  & (~\new_[1523]_  | ~\new_[1557]_ );
  assign \new_[3432]_  = ~\new_[3518]_  & (~\new_[3433]_  | ~\new_[3434]_ );
  assign \new_[3433]_  = ~\new_[1676]_  | ~\new_[1619]_ ;
  assign \new_[3434]_  = ~\new_[1675]_  | ~\new_[3410]_ ;
  assign \new_[3435]_  = ~\new_[3436]_ ;
  assign \new_[3436]_  = ~\new_[3451]_ ;
  assign \new_[3437]_  = ~\new_[3440]_  & (~\new_[3438]_  | ~\new_[3439]_ );
  assign \new_[3438]_  = ~\new_[1689]_  | ~\new_[1618]_ ;
  assign \new_[3439]_  = ~\new_[1688]_  | ~\new_[3410]_ ;
  assign \new_[3440]_  = ~\new_[3441]_ ;
  assign \new_[3441]_  = \new_[3478]_ ;
  assign \new_[3442]_  = ~\new_[1521]_  & (~\new_[1541]_  | ~\new_[1572]_ );
  assign \new_[3443]_  = ~\new_[3444]_ ;
  assign \new_[3444]_  = \new_[3521]_ ;
  assign \new_[3445]_  = ~\new_[3444]_ ;
  assign \new_[3446]_  = ~\new_[3452]_  | (~\new_[3447]_  & ~\new_[3451]_ );
  assign \new_[3447]_  = ~\new_[3448]_ ;
  assign \new_[3448]_  = ~\new_[3449]_  | ~\new_[3450]_ ;
  assign \new_[3449]_  = ~\new_[2793]_  | ~\new_[3150]_ ;
  assign \new_[3450]_  = ~\new_[2933]_  | ~\new_[3061]_ ;
  assign \new_[3451]_  = ~\new_[1662]_ ;
  assign \new_[3452]_  = ~\new_[3435]_  | ~\new_[3061]_ ;
  assign \new_[3453]_  = ~\new_[1694]_  | ~\new_[3454]_  | ~\new_[3458]_ ;
  assign \new_[3454]_  = ~\new_[3455]_  | ~\new_[3456]_ ;
  assign \new_[3455]_  = ~\new_[1668]_  | ~\new_[1669]_ ;
  assign \new_[3456]_  = ~\new_[3457]_ ;
  assign \new_[3457]_  = ~\new_[1865]_  | ~\new_[1864]_ ;
  assign \new_[3458]_  = ~\new_[3457]_  | ~\new_[1668]_  | ~\new_[1669]_ ;
  assign \new_[3459]_  = ~\new_[1694]_ ;
  assign \new_[3460]_  = ~\new_[3275]_  & (~\new_[1574]_  | ~\new_[1543]_ );
  assign \new_[3461]_  = ~\new_[3477]_  & (~\new_[1575]_  | ~\new_[1537]_ );
  assign \new_[3462]_  = ~\new_[3544]_ ;
  assign n796 = ~\new_[3464]_  | ~\new_[3468]_ ;
  assign \new_[3464]_  = ~\new_[3465]_  | ~\new_[3467]_ ;
  assign \new_[3465]_  = ~\new_[3500]_  & ~\new_[3466]_ ;
  assign \new_[3466]_  = ~\new_[3349]_  & ~\new_[3261]_ ;
  assign \new_[3467]_  = ~\new_[3259]_  | ~\new_[3260]_ ;
  assign \new_[3468]_  = ~\new_[2222]_  | ~\new_[557]_ ;
  assign \new_[3469]_  = ~\new_[3477]_  & (~\new_[3470]_  | ~\new_[3471]_ );
  assign \new_[3470]_  = ~\new_[3414]_  | ~\new_[1647]_ ;
  assign \new_[3471]_  = ~\new_[3472]_  | ~\new_[3476]_ ;
  assign \new_[3472]_  = ~\new_[3473]_ ;
  assign \new_[3473]_  = ~\new_[3474]_ ;
  assign \new_[3474]_  = ~\new_[3475]_  & (~\new_[3483]_  | ~\new_[2970]_ );
  assign \new_[3475]_  = \new_[2528]_  & \new_[3490]_ ;
  assign \new_[3476]_  = ~\new_[1743]_  | ~\new_[1815]_ ;
  assign \new_[3477]_  = \new_[3478]_ ;
  assign \new_[3478]_  = ~\new_[3336]_  | ~\new_[3337]_ ;
  assign \new_[3479]_  = ~\new_[3443]_  | (~\new_[3442]_  & ~\new_[3437]_ );
  assign \new_[3480]_  = ~\new_[3520]_  | (~\new_[3469]_  & ~\new_[1503]_ );
  assign \new_[3481]_  = ~\new_[3462]_  | (~\new_[1502]_  & ~\new_[1493]_ );
  assign \new_[3482]_  = ~\new_[3483]_  | ~\new_[3489]_ ;
  assign \new_[3483]_  = \new_[3484]_  ? \new_[3488]_  : \new_[3487]_ ;
  assign \new_[3484]_  = \new_[3485]_ ;
  assign \new_[3485]_  = ~\new_[3486]_ ;
  assign \new_[3486]_  = ~\new_[3122]_  | ~\new_[2756]_ ;
  assign \new_[3487]_  = ~\new_[3484]_ ;
  assign \new_[3488]_  = ~\new_[3321]_  | ~\new_[3510]_ ;
  assign \new_[3489]_  = \new_[1694]_ ;
  assign \new_[3490]_  = ~\new_[3489]_ ;
  assign n811 = ~\new_[3493]_  | (~\new_[3492]_  & ~\new_[953]_ );
  assign \new_[3492]_  = \new_[3500]_  | \new_[2283]_ ;
  assign \new_[3493]_  = ~\new_[3494]_  & (~\new_[2222]_  | ~\new_[560]_ );
  assign \new_[3494]_  = ~\new_[2667]_  & ~\new_[3495]_ ;
  assign \new_[3495]_  = ~\new_[3496]_  | ~\new_[3497]_ ;
  assign \new_[3496]_  = ~\new_[3500]_ ;
  assign \new_[3497]_  = ~\new_[2948]_  | ~\new_[3031]_ ;
  assign n816 = ~\new_[3501]_  | (~\new_[3499]_  & ~\new_[954]_ );
  assign \new_[3499]_  = \new_[3500]_  | \new_[2283]_ ;
  assign \new_[3500]_  = \new_[3306]_  | \new_[3292]_ ;
  assign \new_[3501]_  = ~\new_[3502]_  & (~\new_[2222]_  | ~\new_[561]_ );
  assign \new_[3502]_  = ~\new_[2667]_  & ~\new_[3503]_ ;
  assign \new_[3503]_  = ~\new_[2098]_  | ~\new_[3504]_ ;
  assign \new_[3504]_  = ~\new_[2976]_  | ~\new_[3056]_ ;
  assign \new_[3505]_  = ~\new_[3462]_  | (~\new_[3460]_  & ~\new_[3461]_ );
  assign \new_[3506]_  = ~\new_[3520]_  | (~\new_[1494]_  & ~\new_[1505]_ );
  assign \new_[3507]_  = \new_[3532]_ ;
  assign \new_[3508]_  = \new_[3509]_  ^ \new_[3527]_ ;
  assign \new_[3509]_  = ~\new_[3407]_  | ~\new_[3408]_ ;
  assign \new_[3510]_  = ~\new_[2555]_  | ~\new_[3100]_ ;
  assign \new_[3511]_  = ~\new_[3485]_  & ~\new_[3316]_ ;
  assign \new_[3512]_  = ~\new_[3520]_  | (~\new_[3513]_  & ~\new_[3514]_ );
  assign \new_[3513]_  = ~\new_[3440]_  & (~\new_[1542]_  | ~\new_[1573]_ );
  assign \new_[3514]_  = ~\new_[3517]_  & (~\new_[3515]_  | ~\new_[3516]_ );
  assign \new_[3515]_  = ~\new_[1629]_  | ~\new_[1619]_ ;
  assign \new_[3516]_  = ~\new_[1691]_  | ~\new_[3410]_ ;
  assign \new_[3517]_  = ~\new_[3518]_ ;
  assign \new_[3518]_  = ~\new_[3519]_ ;
  assign \new_[3519]_  = ~\new_[3336]_  | ~\new_[3337]_ ;
  assign \new_[3520]_  = \new_[3521]_ ;
  assign \new_[3521]_  = ~\new_[3343]_  | ~\new_[3338]_  | ~\new_[3340]_ ;
  assign \new_[3522]_  = ~\new_[3518]_ ;
  assign \new_[3523]_  = ~\new_[3524]_  | ~\new_[3528]_ ;
  assign \new_[3524]_  = ~\new_[3525]_  & ~\new_[3527]_ ;
  assign \new_[3525]_  = ~\new_[3526]_ ;
  assign \new_[3526]_  = ~\new_[2516]_  | ~\new_[3140]_ ;
  assign \new_[3527]_  = ~\new_[2308]_  & ~\new_[3511]_ ;
  assign \new_[3528]_  = ~\new_[3446]_  | ~\new_[3149]_ ;
  assign \new_[3529]_  = ~\new_[3524]_ ;
  assign \new_[3530]_  = ~\new_[3520]_  | (~\new_[1506]_  & ~\new_[1495]_ );
  assign \new_[3531]_  = ~\new_[3443]_  | (~\new_[3431]_  & ~\new_[3432]_ );
  assign \new_[3532]_  = ~\new_[3323]_  | ~\new_[3322]_  | ~\new_[3416]_ ;
  assign \new_[3533]_  = ~\new_[3534]_  | ~\new_[3539]_ ;
  assign \new_[3534]_  = ~\new_[3537]_  | (~\new_[3535]_  & ~\new_[3536]_ );
  assign \new_[3535]_  = ~\new_[3208]_  & (~\new_[3480]_  | ~\new_[3481]_ );
  assign \new_[3536]_  = ~\new_[3507]_  & (~\new_[3479]_  | ~\new_[3512]_ );
  assign \new_[3537]_  = ~\new_[3538]_ ;
  assign \new_[3538]_  = ~\new_[3453]_  | ~\new_[3236]_ ;
  assign \new_[3539]_  = ~\new_[3538]_  | (~\new_[3540]_  & ~\new_[3541]_ );
  assign \new_[3540]_  = ~\new_[3507]_  & (~\new_[3505]_  | ~\new_[3506]_ );
  assign \new_[3541]_  = ~\new_[3208]_  & (~\new_[3530]_  | ~\new_[3531]_ );
  assign \new_[3542]_  = ~\new_[3543]_  & ~\new_[3545]_ ;
  assign \new_[3543]_  = \new_[3544]_ ;
  assign \new_[3544]_  = ~\new_[3338]_  | ~\new_[3343]_  | ~\new_[3340]_ ;
  assign \new_[3545]_  = ~\new_[3546]_  | ~\new_[3235]_ ;
  assign \new_[3546]_  = ~\new_[3547]_ ;
  assign \new_[3547]_  = ~\new_[1758]_  | (~\new_[1480]_  & ~\new_[3459]_ );
  assign \new_[3548]_  = ~\new_[3453]_  | ~\new_[3236]_ ;
  assign \new_[3549]_  = ~\new_[3550]_ ;
  assign \new_[3550]_  = ~\new_[3546]_ ;
  always @ (posedge clock) begin
    \\shift_data_reg[39]  <= n186;
    \\shift_data_reg[56]  <= n191;
    \\shift_data_reg[63]  <= n196;
    \\shift_data_reg[32]  <= n201;
    \\shift_data_reg[65]  <= n206;
    \\shift_data_reg[66]  <= n211;
    \\shift_data_reg[68]  <= n216;
    \\shift_data_reg[71]  <= n221;
    \\shift_data_reg[74]  <= n226;
    \\shift_data_reg[75]  <= n231;
    \\shift_data_reg[76]  <= n236;
    \\shift_data_reg[85]  <= n241;
    \\shift_data_reg[86]  <= n246;
    \\shift_data_reg[87]  <= n251;
    \\shift_data_reg[91]  <= n256;
    \\shift_data_reg[93]  <= n261;
    \\shift_data_reg[94]  <= n266;
    \\shift_data_reg[95]  <= n271;
    \\shift_data_reg[0]  <= n276;
    \\shift_data_reg[2]  <= n281;
    \\shift_data_reg[4]  <= n286;
    \\shift_data_reg[7]  <= n291;
    \\shift_data_reg[8]  <= n296;
    \\shift_data_reg[14]  <= n301;
    \\shift_data_reg[15]  <= n306;
    \\shift_data_reg[16]  <= n311;
    \\shift_data_reg[17]  <= n316;
    \\shift_data_reg[18]  <= n321;
    \\shift_data_reg[1]  <= n326;
    \\shift_data_reg[20]  <= n331;
    \\shift_data_reg[23]  <= n336;
    \\shift_data_reg[92]  <= n341;
    \\shift_data_reg[89]  <= n346;
    \\shift_data_reg[64]  <= n351;
    \\shift_data_reg[67]  <= n356;
    \\shift_data_reg[69]  <= n361;
    \\shift_data_reg[70]  <= n366;
    \\shift_data_reg[72]  <= n371;
    \\shift_data_reg[73]  <= n376;
    \\shift_data_reg[77]  <= n381;
    \\shift_data_reg[80]  <= n386;
    \\shift_data_reg[83]  <= n391;
    \\shift_data_reg[84]  <= n396;
    \\shift_data_reg[81]  <= n401;
    \\shift_data_reg[88]  <= n406;
    \\shift_data_reg[82]  <= n411;
    \\shift_data_reg[90]  <= n416;
    \\shift_data_reg[79]  <= n421;
    \\shift_data_reg[78]  <= n426;
    \\shift_data_reg[26]  <= n431;
    \\shift_data_reg[27]  <= n436;
    \\shift_data_reg[24]  <= n441;
    \\shift_data_reg[29]  <= n446;
    \\shift_data_reg[28]  <= n451;
    \\shift_data_reg[30]  <= n456;
    \\shift_data_reg[31]  <= n461;
    \\shift_data_reg[10]  <= n466;
    \\shift_data_reg[3]  <= n471;
    \\shift_data_reg[5]  <= n476;
    \\shift_data_reg[25]  <= n481;
    \\shift_data_reg[6]  <= n486;
    \\shift_data_reg[12]  <= n491;
    \\shift_data_reg[13]  <= n496;
    \\shift_data_reg[11]  <= n501;
    \\shift_data_reg[9]  <= n506;
    \\shift_data_reg[19]  <= n511;
    \\shift_data_reg[21]  <= n516;
    \\shift_data_reg[22]  <= n521;
    \\shift_data_reg[53]  <= n526;
    \\shift_data_reg[54]  <= n531;
    \\shift_data_reg[51]  <= n536;
    \\shift_data_reg[33]  <= n541;
    \\shift_data_reg[34]  <= n546;
    \\shift_data_reg[35]  <= n551;
    \\shift_data_reg[36]  <= n556;
    \\shift_data_reg[43]  <= n561;
    \\shift_data_reg[45]  <= n566;
    \\shift_data_reg[46]  <= n571;
    \\shift_data_reg[47]  <= n576;
    \\shift_data_reg[57]  <= n581;
    \\shift_data_reg[58]  <= n586;
    \\shift_data_reg[59]  <= n591;
    \\shift_data_reg[61]  <= n596;
    \\shift_data_reg[62]  <= n601;
    \\shift_data_reg[104]  <= n606;
    \\shift_data_reg[111]  <= n611;
    \\shift_data_reg[112]  <= n616;
    \\shift_data_reg[119]  <= n621;
    \\shift_data_reg[121]  <= n626;
    \\shift_data_reg[97]  <= n631;
    \\shift_data_reg[123]  <= n636;
    \\shift_data_reg[125]  <= n641;
    \\shift_data_reg[126]  <= n646;
    \\shift_data_reg[122]  <= n651;
    \\shift_data_reg[127]  <= n656;
    \\shift_data_reg[124]  <= n661;
    \\shift_data_reg[98]  <= n666;
    \\shift_data_reg[114]  <= n671;
    \\shift_data_reg[60]  <= n676;
    \\shift_data_reg[48]  <= n681;
    \\shift_data_reg[41]  <= n686;
    \\shift_data_reg[40]  <= n691;
    \\shift_data_reg[120]  <= n696;
    \\shift_data_reg[105]  <= n701;
    \\shift_data_reg[113]  <= n706;
    \\shift_data_reg[108]  <= n711;
    \\shift_data_reg[37]  <= n716;
    \\shift_data_reg[38]  <= n721;
    \\shift_data_reg[116]  <= n726;
    \\shift_data_reg[42]  <= n731;
    \\shift_data_reg[49]  <= n736;
    \\shift_data_reg[50]  <= n741;
    \\shift_data_reg[44]  <= n746;
    \\shift_data_reg[52]  <= n751;
    \\shift_data_reg[55]  <= n756;
    \\shift_data_reg[103]  <= n761;
    \\shift_data_reg[100]  <= n766;
    \\shift_data_reg[106]  <= n771;
    \\shift_data_reg[96]  <= n776;
    \\shift_data_reg[99]  <= n781;
    \\shift_data_reg[118]  <= n786;
    \\shift_data_reg[115]  <= n791;
    \\shift_data_reg[101]  <= n796;
    \\shift_data_reg[102]  <= n801;
    \\shift_data_reg[107]  <= n806;
    \\shift_data_reg[109]  <= n811;
    \\shift_data_reg[110]  <= n816;
    \\shift_data_reg[117]  <= n821;
    shift_s_out_reg <= n826;
    clgen_clk_out_reg <= n831;
    \\shift_cnt_reg[7]  <= n836;
    \\ctrl_reg[8]  <= n841;
    \\clgen_cnt_reg[15]  <= n846;
    \\shift_cnt_reg[6]  <= n851;
    wb_int_o_reg <= n856;
    \\wb_dat_o_reg[9]  <= n861;
    shift_tip_reg <= n866;
    \\wb_dat_o_reg[11]  <= n871;
    \\ctrl_reg[9]  <= n876;
    \\shift_cnt_reg[4]  <= n881;
    \\shift_cnt_reg[5]  <= n886;
    \\clgen_cnt_reg[11]  <= n891;
    \\shift_cnt_reg[3]  <= n896;
    \\ctrl_reg[11]  <= n901;
    \\ctrl_reg[10]  <= n906;
    clgen_pos_edge_reg <= n911;
    clgen_neg_edge_reg <= n916;
    \\clgen_cnt_reg[14]  <= n921;
    \\shift_cnt_reg[2]  <= n926;
    \\clgen_cnt_reg[13]  <= n931;
    \\ctrl_reg[0]  <= n936;
    \\ctrl_reg[12]  <= n941;
    \\ctrl_reg[13]  <= n946;
    \\divider_reg[11]  <= n951;
    \\clgen_cnt_reg[12]  <= n956;
    \\divider_reg[4]  <= n961;
    \\ctrl_reg[2]  <= n966;
    \\divider_reg[15]  <= n971;
    \\ctrl_reg[7]  <= n976;
    \\clgen_cnt_reg[10]  <= n981;
    \\divider_reg[8]  <= n986;
    \\ctrl_reg[5]  <= n991;
    \\clgen_cnt_reg[3]  <= n996;
    \\divider_reg[13]  <= n1001;
    \\clgen_cnt_reg[5]  <= n1006;
    \\clgen_cnt_reg[0]  <= n1011;
    \\clgen_cnt_reg[2]  <= n1016;
    \\clgen_cnt_reg[7]  <= n1021;
    \\clgen_cnt_reg[6]  <= n1026;
    \\clgen_cnt_reg[9]  <= n1031;
    \\clgen_cnt_reg[1]  <= n1036;
    \\ctrl_reg[1]  <= n1041;
    \\divider_reg[12]  <= n1046;
    \\divider_reg[10]  <= n1051;
    \\divider_reg[1]  <= n1056;
    \\divider_reg[2]  <= n1061;
    \\ctrl_reg[3]  <= n1066;
    \\ctrl_reg[4]  <= n1071;
    \\ctrl_reg[6]  <= n1076;
    \\divider_reg[0]  <= n1081;
    \\divider_reg[14]  <= n1086;
    \\divider_reg[3]  <= n1091;
    \\divider_reg[5]  <= n1096;
    \\divider_reg[6]  <= n1101;
    \\divider_reg[7]  <= n1106;
    \\divider_reg[9]  <= n1111;
    \\clgen_cnt_reg[4]  <= n1116;
    \\shift_cnt_reg[1]  <= n1121;
    \\wb_dat_o_reg[7]  <= n1126;
    \\wb_dat_o_reg[3]  <= n1131;
    \\shift_cnt_reg[0]  <= n1136;
    \\clgen_cnt_reg[8]  <= n1141;
    \\ss_reg[5]  <= n1146;
    \\ss_reg[3]  <= n1151;
    \\ss_reg[1]  <= n1156;
    \\ss_reg[7]  <= n1161;
    \\ss_reg[0]  <= n1166;
    \\ss_reg[2]  <= n1171;
    \\ss_reg[4]  <= n1176;
    \\ss_reg[6]  <= n1181;
    \\wb_dat_o_reg[4]  <= n1186;
    \\wb_dat_o_reg[5]  <= n1191;
    \\wb_dat_o_reg[0]  <= n1196;
    \\wb_dat_o_reg[1]  <= n1201;
    \\wb_dat_o_reg[6]  <= n1206;
    \\wb_dat_o_reg[2]  <= n1211;
    \\wb_dat_o_reg[10]  <= n1216;
    \\wb_dat_o_reg[13]  <= n1221;
    \\wb_dat_o_reg[14]  <= n1226;
    \\wb_dat_o_reg[12]  <= n1231;
    \\wb_dat_o_reg[8]  <= n1236;
    \\wb_dat_o_reg[15]  <= n1241;
    \\wb_dat_o_reg[26]  <= n1246;
    \\wb_dat_o_reg[16]  <= n1251;
    \\wb_dat_o_reg[18]  <= n1256;
    \\wb_dat_o_reg[17]  <= n1261;
    \\wb_dat_o_reg[19]  <= n1266;
    \\wb_dat_o_reg[22]  <= n1271;
    \\wb_dat_o_reg[27]  <= n1276;
    \\wb_dat_o_reg[21]  <= n1281;
    \\wb_dat_o_reg[31]  <= n1286;
    \\wb_dat_o_reg[28]  <= n1291;
    \\wb_dat_o_reg[24]  <= n1296;
    \\wb_dat_o_reg[23]  <= n1301;
    \\wb_dat_o_reg[30]  <= n1306;
    \\wb_dat_o_reg[20]  <= n1311;
    \\wb_dat_o_reg[29]  <= n1316;
    \\wb_dat_o_reg[25]  <= n1321;
    wb_ack_o_reg <= n1326;
  end
  initial begin
    \\shift_data_reg[39]  <= 1'b0;
    \\shift_data_reg[56]  <= 1'b0;
    \\shift_data_reg[63]  <= 1'b0;
    \\shift_data_reg[32]  <= 1'b0;
    \\shift_data_reg[65]  <= 1'b0;
    \\shift_data_reg[66]  <= 1'b0;
    \\shift_data_reg[68]  <= 1'b0;
    \\shift_data_reg[71]  <= 1'b0;
    \\shift_data_reg[74]  <= 1'b0;
    \\shift_data_reg[75]  <= 1'b0;
    \\shift_data_reg[76]  <= 1'b0;
    \\shift_data_reg[85]  <= 1'b0;
    \\shift_data_reg[86]  <= 1'b0;
    \\shift_data_reg[87]  <= 1'b0;
    \\shift_data_reg[91]  <= 1'b0;
    \\shift_data_reg[93]  <= 1'b0;
    \\shift_data_reg[94]  <= 1'b0;
    \\shift_data_reg[95]  <= 1'b0;
    \\shift_data_reg[0]  <= 1'b0;
    \\shift_data_reg[2]  <= 1'b0;
    \\shift_data_reg[4]  <= 1'b0;
    \\shift_data_reg[7]  <= 1'b0;
    \\shift_data_reg[8]  <= 1'b0;
    \\shift_data_reg[14]  <= 1'b0;
    \\shift_data_reg[15]  <= 1'b0;
    \\shift_data_reg[16]  <= 1'b0;
    \\shift_data_reg[17]  <= 1'b0;
    \\shift_data_reg[18]  <= 1'b0;
    \\shift_data_reg[1]  <= 1'b0;
    \\shift_data_reg[20]  <= 1'b0;
    \\shift_data_reg[23]  <= 1'b0;
    \\shift_data_reg[92]  <= 1'b0;
    \\shift_data_reg[89]  <= 1'b0;
    \\shift_data_reg[64]  <= 1'b0;
    \\shift_data_reg[67]  <= 1'b0;
    \\shift_data_reg[69]  <= 1'b0;
    \\shift_data_reg[70]  <= 1'b0;
    \\shift_data_reg[72]  <= 1'b0;
    \\shift_data_reg[73]  <= 1'b0;
    \\shift_data_reg[77]  <= 1'b0;
    \\shift_data_reg[80]  <= 1'b0;
    \\shift_data_reg[83]  <= 1'b0;
    \\shift_data_reg[84]  <= 1'b0;
    \\shift_data_reg[81]  <= 1'b0;
    \\shift_data_reg[88]  <= 1'b0;
    \\shift_data_reg[82]  <= 1'b0;
    \\shift_data_reg[90]  <= 1'b0;
    \\shift_data_reg[79]  <= 1'b0;
    \\shift_data_reg[78]  <= 1'b0;
    \\shift_data_reg[26]  <= 1'b0;
    \\shift_data_reg[27]  <= 1'b0;
    \\shift_data_reg[24]  <= 1'b0;
    \\shift_data_reg[29]  <= 1'b0;
    \\shift_data_reg[28]  <= 1'b0;
    \\shift_data_reg[30]  <= 1'b0;
    \\shift_data_reg[31]  <= 1'b0;
    \\shift_data_reg[10]  <= 1'b0;
    \\shift_data_reg[3]  <= 1'b0;
    \\shift_data_reg[5]  <= 1'b0;
    \\shift_data_reg[25]  <= 1'b0;
    \\shift_data_reg[6]  <= 1'b0;
    \\shift_data_reg[12]  <= 1'b0;
    \\shift_data_reg[13]  <= 1'b0;
    \\shift_data_reg[11]  <= 1'b0;
    \\shift_data_reg[9]  <= 1'b0;
    \\shift_data_reg[19]  <= 1'b0;
    \\shift_data_reg[21]  <= 1'b0;
    \\shift_data_reg[22]  <= 1'b0;
    \\shift_data_reg[53]  <= 1'b0;
    \\shift_data_reg[54]  <= 1'b0;
    \\shift_data_reg[51]  <= 1'b0;
    \\shift_data_reg[33]  <= 1'b0;
    \\shift_data_reg[34]  <= 1'b0;
    \\shift_data_reg[35]  <= 1'b0;
    \\shift_data_reg[36]  <= 1'b0;
    \\shift_data_reg[43]  <= 1'b0;
    \\shift_data_reg[45]  <= 1'b0;
    \\shift_data_reg[46]  <= 1'b0;
    \\shift_data_reg[47]  <= 1'b0;
    \\shift_data_reg[57]  <= 1'b0;
    \\shift_data_reg[58]  <= 1'b0;
    \\shift_data_reg[59]  <= 1'b0;
    \\shift_data_reg[61]  <= 1'b0;
    \\shift_data_reg[62]  <= 1'b0;
    \\shift_data_reg[104]  <= 1'b0;
    \\shift_data_reg[111]  <= 1'b0;
    \\shift_data_reg[112]  <= 1'b0;
    \\shift_data_reg[119]  <= 1'b0;
    \\shift_data_reg[121]  <= 1'b0;
    \\shift_data_reg[97]  <= 1'b0;
    \\shift_data_reg[123]  <= 1'b0;
    \\shift_data_reg[125]  <= 1'b0;
    \\shift_data_reg[126]  <= 1'b0;
    \\shift_data_reg[122]  <= 1'b0;
    \\shift_data_reg[127]  <= 1'b0;
    \\shift_data_reg[124]  <= 1'b0;
    \\shift_data_reg[98]  <= 1'b0;
    \\shift_data_reg[114]  <= 1'b0;
    \\shift_data_reg[60]  <= 1'b0;
    \\shift_data_reg[48]  <= 1'b0;
    \\shift_data_reg[41]  <= 1'b0;
    \\shift_data_reg[40]  <= 1'b0;
    \\shift_data_reg[120]  <= 1'b0;
    \\shift_data_reg[105]  <= 1'b0;
    \\shift_data_reg[113]  <= 1'b0;
    \\shift_data_reg[108]  <= 1'b0;
    \\shift_data_reg[37]  <= 1'b0;
    \\shift_data_reg[38]  <= 1'b0;
    \\shift_data_reg[116]  <= 1'b0;
    \\shift_data_reg[42]  <= 1'b0;
    \\shift_data_reg[49]  <= 1'b0;
    \\shift_data_reg[50]  <= 1'b0;
    \\shift_data_reg[44]  <= 1'b0;
    \\shift_data_reg[52]  <= 1'b0;
    \\shift_data_reg[55]  <= 1'b0;
    \\shift_data_reg[103]  <= 1'b0;
    \\shift_data_reg[100]  <= 1'b0;
    \\shift_data_reg[106]  <= 1'b0;
    \\shift_data_reg[96]  <= 1'b0;
    \\shift_data_reg[99]  <= 1'b0;
    \\shift_data_reg[118]  <= 1'b0;
    \\shift_data_reg[115]  <= 1'b0;
    \\shift_data_reg[101]  <= 1'b0;
    \\shift_data_reg[102]  <= 1'b0;
    \\shift_data_reg[107]  <= 1'b0;
    \\shift_data_reg[109]  <= 1'b0;
    \\shift_data_reg[110]  <= 1'b0;
    \\shift_data_reg[117]  <= 1'b0;
    shift_s_out_reg <= 1'b0;
    clgen_clk_out_reg <= 1'b0;
    \\shift_cnt_reg[7]  <= 1'b0;
    \\ctrl_reg[8]  <= 1'b0;
    \\clgen_cnt_reg[15]  <= 1'b1;
    \\shift_cnt_reg[6]  <= 1'b0;
    wb_int_o_reg <= 1'b0;
    \\wb_dat_o_reg[9]  <= 1'b0;
    shift_tip_reg <= 1'b0;
    \\wb_dat_o_reg[11]  <= 1'b0;
    \\ctrl_reg[9]  <= 1'b0;
    \\shift_cnt_reg[4]  <= 1'b0;
    \\shift_cnt_reg[5]  <= 1'b0;
    \\clgen_cnt_reg[11]  <= 1'b1;
    \\shift_cnt_reg[3]  <= 1'b0;
    \\ctrl_reg[11]  <= 1'b0;
    \\ctrl_reg[10]  <= 1'b0;
    clgen_pos_edge_reg <= 1'b0;
    clgen_neg_edge_reg <= 1'b0;
    \\clgen_cnt_reg[14]  <= 1'b1;
    \\shift_cnt_reg[2]  <= 1'b0;
    \\clgen_cnt_reg[13]  <= 1'b1;
    \\ctrl_reg[0]  <= 1'b0;
    \\ctrl_reg[12]  <= 1'b0;
    \\ctrl_reg[13]  <= 1'b0;
    \\divider_reg[11]  <= 1'b0;
    \\clgen_cnt_reg[12]  <= 1'b1;
    \\divider_reg[4]  <= 1'b0;
    \\ctrl_reg[2]  <= 1'b0;
    \\divider_reg[15]  <= 1'b0;
    \\ctrl_reg[7]  <= 1'b0;
    \\clgen_cnt_reg[10]  <= 1'b1;
    \\divider_reg[8]  <= 1'b0;
    \\ctrl_reg[5]  <= 1'b0;
    \\clgen_cnt_reg[3]  <= 1'b1;
    \\divider_reg[13]  <= 1'b0;
    \\clgen_cnt_reg[5]  <= 1'b1;
    \\clgen_cnt_reg[0]  <= 1'b1;
    \\clgen_cnt_reg[2]  <= 1'b1;
    \\clgen_cnt_reg[7]  <= 1'b1;
    \\clgen_cnt_reg[6]  <= 1'b1;
    \\clgen_cnt_reg[9]  <= 1'b1;
    \\clgen_cnt_reg[1]  <= 1'b1;
    \\ctrl_reg[1]  <= 1'b0;
    \\divider_reg[12]  <= 1'b0;
    \\divider_reg[10]  <= 1'b0;
    \\divider_reg[1]  <= 1'b0;
    \\divider_reg[2]  <= 1'b0;
    \\ctrl_reg[3]  <= 1'b0;
    \\ctrl_reg[4]  <= 1'b0;
    \\ctrl_reg[6]  <= 1'b0;
    \\divider_reg[0]  <= 1'b0;
    \\divider_reg[14]  <= 1'b0;
    \\divider_reg[3]  <= 1'b0;
    \\divider_reg[5]  <= 1'b0;
    \\divider_reg[6]  <= 1'b0;
    \\divider_reg[7]  <= 1'b0;
    \\divider_reg[9]  <= 1'b0;
    \\clgen_cnt_reg[4]  <= 1'b1;
    \\shift_cnt_reg[1]  <= 1'b0;
    \\wb_dat_o_reg[7]  <= 1'b0;
    \\wb_dat_o_reg[3]  <= 1'b0;
    \\shift_cnt_reg[0]  <= 1'b0;
    \\clgen_cnt_reg[8]  <= 1'b1;
    \\ss_reg[5]  <= 1'b0;
    \\ss_reg[3]  <= 1'b0;
    \\ss_reg[1]  <= 1'b0;
    \\ss_reg[7]  <= 1'b0;
    \\ss_reg[0]  <= 1'b0;
    \\ss_reg[2]  <= 1'b0;
    \\ss_reg[4]  <= 1'b0;
    \\ss_reg[6]  <= 1'b0;
    \\wb_dat_o_reg[4]  <= 1'b0;
    \\wb_dat_o_reg[5]  <= 1'b0;
    \\wb_dat_o_reg[0]  <= 1'b0;
    \\wb_dat_o_reg[1]  <= 1'b0;
    \\wb_dat_o_reg[6]  <= 1'b0;
    \\wb_dat_o_reg[2]  <= 1'b0;
    \\wb_dat_o_reg[10]  <= 1'b0;
    \\wb_dat_o_reg[13]  <= 1'b0;
    \\wb_dat_o_reg[14]  <= 1'b0;
    \\wb_dat_o_reg[12]  <= 1'b0;
    \\wb_dat_o_reg[8]  <= 1'b0;
    \\wb_dat_o_reg[15]  <= 1'b0;
    \\wb_dat_o_reg[26]  <= 1'b0;
    \\wb_dat_o_reg[16]  <= 1'b0;
    \\wb_dat_o_reg[18]  <= 1'b0;
    \\wb_dat_o_reg[17]  <= 1'b0;
    \\wb_dat_o_reg[19]  <= 1'b0;
    \\wb_dat_o_reg[22]  <= 1'b0;
    \\wb_dat_o_reg[27]  <= 1'b0;
    \\wb_dat_o_reg[21]  <= 1'b0;
    \\wb_dat_o_reg[31]  <= 1'b0;
    \\wb_dat_o_reg[28]  <= 1'b0;
    \\wb_dat_o_reg[24]  <= 1'b0;
    \\wb_dat_o_reg[23]  <= 1'b0;
    \\wb_dat_o_reg[30]  <= 1'b0;
    \\wb_dat_o_reg[20]  <= 1'b0;
    \\wb_dat_o_reg[29]  <= 1'b0;
    \\wb_dat_o_reg[25]  <= 1'b0;
    wb_ack_o_reg <= 1'b0;
  end
endmodule


