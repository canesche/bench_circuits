module pair ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, y,
    z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0,
    r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1,
    j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2,
    b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2,
    t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3,
    l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4,
    d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4,
    v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5,
    n5, o5, p5, q5, r5,
    s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6,
    k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7,
    c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7,
    u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8,
    m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9,
    e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9,
    w9, x9, y9, z9, a10, b10, c10, d10, e10, f10, g10, h10, i10, j10, k10,
    l10, m10, n10, o10, p10, q10, r10, s10, t10, u10, v10, w10, x10, y10  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0,
    p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1,
    h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1,
    z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2,
    r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3,
    j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4,
    b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4,
    t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5,
    l5, m5, n5, o5, p5, q5, r5;
  output s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6,
    j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7,
    b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7,
    t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8,
    l8, m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9,
    d9, e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9,
    v9, w9, x9, y9, z9, a10, b10, c10, d10, e10, f10, g10, h10, i10, j10,
    k10, l10, m10, n10, o10, p10, q10, r10, s10, t10, u10, v10, w10, x10,
    y10;
  wire new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_,
    new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_,
    new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n942_, new_n943_, new_n945_, new_n946_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n965_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n996_,
    new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_,
    new_n1003_, new_n1004_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1042_, new_n1043_,
    new_n1044_, new_n1046_, new_n1047_, new_n1048_, new_n1050_, new_n1051_,
    new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_,
    new_n1058_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1098_, new_n1099_, new_n1100_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_,
    new_n1124_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1188_, new_n1189_,
    new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1213_, new_n1214_, new_n1215_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1245_, new_n1246_, new_n1247_, new_n1248_,
    new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_,
    new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1268_,
    new_n1269_, new_n1270_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1307_, new_n1308_,
    new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1368_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1383_, new_n1384_, new_n1385_, new_n1386_,
    new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_, new_n1392_,
    new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_,
    new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1482_,
    new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_, new_n1488_,
    new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_, new_n1494_,
    new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_, new_n1501_,
    new_n1502_, new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_,
    new_n1508_, new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_,
    new_n1514_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1533_, new_n1534_,
    new_n1536_, new_n1537_, new_n1539_, new_n1540_, new_n1541_, new_n1542_,
    new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_, new_n1548_,
    new_n1549_, new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_,
    new_n1556_, new_n1557_, new_n1559_, new_n1560_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1600_, new_n1601_, new_n1602_, new_n1603_,
    new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1648_, new_n1649_, new_n1650_,
    new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1683_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1697_, new_n1698_, new_n1699_, new_n1701_,
    new_n1702_, new_n1703_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1730_,
    new_n1731_, new_n1732_, new_n1734_, new_n1735_, new_n1736_, new_n1737_,
    new_n1738_, new_n1739_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1789_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1800_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_,
    new_n1809_;
  assign new_n311_ = w & y0;
  assign new_n312_ = v & d1;
  assign new_n313_ = u & g2;
  assign new_n314_ = t & j2;
  assign new_n315_ = ~new_n311_ & ~new_n312_;
  assign new_n316_ = ~new_n313_ & ~new_n314_;
  assign new_n317_ = new_n315_ & new_n316_;
  assign new_n318_ = s & o2;
  assign new_n319_ = r & u1;
  assign new_n320_ = q & x1;
  assign new_n321_ = p & a2;
  assign new_n322_ = ~new_n318_ & ~new_n319_;
  assign new_n323_ = ~new_n320_ & ~new_n321_;
  assign new_n324_ = new_n322_ & new_n323_;
  assign new_n325_ = o & t2;
  assign new_n326_ = n & a3;
  assign new_n327_ = m & e3;
  assign new_n328_ = ~new_n325_ & ~new_n326_;
  assign new_n329_ = ~new_n327_ & new_n328_;
  assign new_n330_ = new_n317_ & new_n324_;
  assign s5 = ~new_n329_ | ~new_n330_;
  assign new_n332_ = w & x0;
  assign new_n333_ = v & c1;
  assign new_n334_ = u & d2;
  assign new_n335_ = t & i2;
  assign new_n336_ = ~new_n332_ & ~new_n333_;
  assign new_n337_ = ~new_n334_ & ~new_n335_;
  assign new_n338_ = new_n336_ & new_n337_;
  assign new_n339_ = s & m2;
  assign new_n340_ = r & t1;
  assign new_n341_ = q & w1;
  assign new_n342_ = p & z1;
  assign new_n343_ = ~new_n339_ & ~new_n340_;
  assign new_n344_ = ~new_n341_ & ~new_n342_;
  assign new_n345_ = new_n343_ & new_n344_;
  assign new_n346_ = o & s2;
  assign new_n347_ = n & z2;
  assign new_n348_ = m & d3;
  assign new_n349_ = ~new_n346_ & ~new_n347_;
  assign new_n350_ = ~new_n348_ & new_n349_;
  assign new_n351_ = new_n338_ & new_n345_;
  assign t5 = ~new_n350_ | ~new_n351_;
  assign new_n353_ = w & w0;
  assign new_n354_ = v & b1;
  assign new_n355_ = u & c2;
  assign new_n356_ = t & h2;
  assign new_n357_ = ~new_n353_ & ~new_n354_;
  assign new_n358_ = ~new_n355_ & ~new_n356_;
  assign new_n359_ = new_n357_ & new_n358_;
  assign new_n360_ = s & l2;
  assign new_n361_ = r & s1;
  assign new_n362_ = q & v1;
  assign new_n363_ = p & y1;
  assign new_n364_ = ~new_n360_ & ~new_n361_;
  assign new_n365_ = ~new_n362_ & ~new_n363_;
  assign new_n366_ = new_n364_ & new_n365_;
  assign new_n367_ = o & r2;
  assign new_n368_ = n & y2;
  assign new_n369_ = m & c3;
  assign new_n370_ = ~new_n367_ & ~new_n368_;
  assign new_n371_ = ~new_n369_ & new_n370_;
  assign new_n372_ = new_n359_ & new_n366_;
  assign u5 = ~new_n371_ | ~new_n372_;
  assign new_n374_ = w & v0;
  assign new_n375_ = v & a1;
  assign new_n376_ = u & b2;
  assign new_n377_ = t & f2;
  assign new_n378_ = ~new_n374_ & ~new_n375_;
  assign new_n379_ = ~new_n376_ & ~new_n377_;
  assign new_n380_ = new_n378_ & new_n379_;
  assign new_n381_ = s & k2;
  assign new_n382_ = r & m1;
  assign new_n383_ = q & r1;
  assign new_n384_ = p & p1;
  assign new_n385_ = ~new_n381_ & ~new_n382_;
  assign new_n386_ = ~new_n383_ & ~new_n384_;
  assign new_n387_ = new_n385_ & new_n386_;
  assign new_n388_ = o & q2;
  assign new_n389_ = n & x2;
  assign new_n390_ = m & b3;
  assign new_n391_ = ~new_n388_ & ~new_n389_;
  assign new_n392_ = ~new_n390_ & new_n391_;
  assign new_n393_ = new_n380_ & new_n387_;
  assign v5 = ~new_n392_ | ~new_n393_;
  assign new_n395_ = w & l1;
  assign new_n396_ = v & z0;
  assign new_n397_ = ~h1 & ~i1;
  assign new_n398_ = e1 & ~f1;
  assign new_n399_ = ~k1 & o1;
  assign new_n400_ = ~j1 & ~o1;
  assign new_n401_ = ~new_n399_ & ~new_n400_;
  assign new_n402_ = j1 & ~new_n401_;
  assign new_n403_ = ~new_n398_ & new_n402_;
  assign new_n404_ = new_n398_ & ~new_n402_;
  assign new_n405_ = ~new_n403_ & ~new_n404_;
  assign new_n406_ = new_n397_ & ~new_n405_;
  assign new_n407_ = new_n402_ & new_n406_;
  assign new_n408_ = ~h1 & ~new_n407_;
  assign new_n409_ = new_n398_ & ~new_n405_;
  assign new_n410_ = new_n397_ & new_n409_;
  assign n6 = i1 | new_n410_;
  assign new_n412_ = ~g1 & ~n6;
  assign new_n413_ = ~x0 & ~y0;
  assign new_n414_ = ~z0 & new_n413_;
  assign new_n415_ = ~a1 & new_n414_;
  assign new_n416_ = ~b1 & new_n415_;
  assign new_n417_ = ~c1 & new_n416_;
  assign new_n418_ = ~w0 & new_n417_;
  assign new_n419_ = ~d1 & new_n418_;
  assign new_n420_ = ~v0 & new_n419_;
  assign new_n421_ = new_n408_ & new_n412_;
  assign new_n422_ = new_n420_ & ~new_n421_;
  assign new_n423_ = l1 & m1;
  assign new_n424_ = ~b & ~n1;
  assign new_n425_ = new_n423_ & new_n424_;
  assign new_n426_ = ~l1 & ~m1;
  assign new_n427_ = ~n1 & new_n426_;
  assign v6 = b | new_n427_;
  assign new_n429_ = new_n422_ & v6;
  assign new_n430_ = ~v0 & r1;
  assign new_n431_ = new_n425_ & ~new_n430_;
  assign new_n432_ = ~new_n429_ & ~new_n431_;
  assign new_n433_ = ~f & new_n432_;
  assign new_n434_ = u & new_n433_;
  assign new_n435_ = t & e2;
  assign new_n436_ = ~new_n395_ & ~new_n396_;
  assign new_n437_ = ~new_n434_ & ~new_n435_;
  assign new_n438_ = new_n436_ & new_n437_;
  assign new_n439_ = ~l & q1;
  assign new_n440_ = b2 & c2;
  assign new_n441_ = d2 & new_n440_;
  assign new_n442_ = ~new_n439_ & ~new_n441_;
  assign new_n443_ = g2 & ~new_n442_;
  assign new_n444_ = ~l & ~p1;
  assign new_n445_ = ~new_n443_ & new_n444_;
  assign new_n446_ = e2 & ~new_n445_;
  assign new_n447_ = n2 & new_n446_;
  assign new_n448_ = s & new_n447_;
  assign new_n449_ = r & n1;
  assign new_n450_ = ~l1 & m1;
  assign new_n451_ = ~n1 & new_n450_;
  assign new_n452_ = ~b & new_n451_;
  assign new_n453_ = ~b & ~new_n452_;
  assign new_n454_ = q & ~new_n453_;
  assign new_n455_ = p & q1;
  assign new_n456_ = ~new_n448_ & ~new_n449_;
  assign new_n457_ = ~new_n454_ & ~new_n455_;
  assign new_n458_ = new_n456_ & new_n457_;
  assign new_n459_ = d3 & e3;
  assign new_n460_ = c3 & new_n459_;
  assign new_n461_ = o & new_n460_;
  assign new_n462_ = n & w2;
  assign new_n463_ = y2 & ~z2;
  assign new_n464_ = ~a3 & new_n463_;
  assign new_n465_ = ~b3 & ~c3;
  assign new_n466_ = ~d3 & ~e3;
  assign new_n467_ = new_n465_ & new_n466_;
  assign new_n468_ = new_n464_ & new_n467_;
  assign new_n469_ = m & new_n468_;
  assign new_n470_ = ~new_n461_ & ~new_n462_;
  assign new_n471_ = ~new_n469_ & new_n470_;
  assign new_n472_ = new_n438_ & new_n458_;
  assign w5 = ~new_n471_ | ~new_n472_;
  assign new_n474_ = u0 & u4;
  assign new_n475_ = t0 & z4;
  assign new_n476_ = s0 & i4;
  assign new_n477_ = r0 & l4;
  assign new_n478_ = ~new_n474_ & ~new_n475_;
  assign new_n479_ = ~new_n476_ & ~new_n477_;
  assign new_n480_ = new_n478_ & new_n479_;
  assign new_n481_ = q0 & q4;
  assign new_n482_ = p0 & w3;
  assign new_n483_ = o0 & z3;
  assign new_n484_ = n0 & c4;
  assign new_n485_ = ~new_n481_ & ~new_n482_;
  assign new_n486_ = ~new_n483_ & ~new_n484_;
  assign new_n487_ = new_n485_ & new_n486_;
  assign new_n488_ = m0 & i3;
  assign new_n489_ = l0 & p3;
  assign new_n490_ = k0 & t3;
  assign new_n491_ = ~new_n488_ & ~new_n489_;
  assign new_n492_ = ~new_n490_ & new_n491_;
  assign new_n493_ = new_n480_ & new_n487_;
  assign x5 = ~new_n492_ | ~new_n493_;
  assign new_n495_ = u0 & t4;
  assign new_n496_ = t0 & y4;
  assign new_n497_ = s0 & f4;
  assign new_n498_ = r0 & k4;
  assign new_n499_ = ~new_n495_ & ~new_n496_;
  assign new_n500_ = ~new_n497_ & ~new_n498_;
  assign new_n501_ = new_n499_ & new_n500_;
  assign new_n502_ = q0 & o4;
  assign new_n503_ = p0 & v3;
  assign new_n504_ = o0 & y3;
  assign new_n505_ = n0 & b4;
  assign new_n506_ = ~new_n502_ & ~new_n503_;
  assign new_n507_ = ~new_n504_ & ~new_n505_;
  assign new_n508_ = new_n506_ & new_n507_;
  assign new_n509_ = m0 & h3;
  assign new_n510_ = l0 & o3;
  assign new_n511_ = k0 & s3;
  assign new_n512_ = ~new_n509_ & ~new_n510_;
  assign new_n513_ = ~new_n511_ & new_n512_;
  assign new_n514_ = new_n501_ & new_n508_;
  assign y5 = ~new_n513_ | ~new_n514_;
  assign new_n516_ = u0 & s4;
  assign new_n517_ = t0 & x4;
  assign new_n518_ = s0 & e4;
  assign new_n519_ = r0 & j4;
  assign new_n520_ = ~new_n516_ & ~new_n517_;
  assign new_n521_ = ~new_n518_ & ~new_n519_;
  assign new_n522_ = new_n520_ & new_n521_;
  assign new_n523_ = q0 & n4;
  assign new_n524_ = p0 & u3;
  assign new_n525_ = o0 & x3;
  assign new_n526_ = n0 & a4;
  assign new_n527_ = ~new_n523_ & ~new_n524_;
  assign new_n528_ = ~new_n525_ & ~new_n526_;
  assign new_n529_ = new_n527_ & new_n528_;
  assign new_n530_ = m0 & g3;
  assign new_n531_ = l0 & n3;
  assign new_n532_ = k0 & r3;
  assign new_n533_ = ~new_n530_ & ~new_n531_;
  assign new_n534_ = ~new_n532_ & new_n533_;
  assign new_n535_ = new_n522_ & new_n529_;
  assign z5 = ~new_n534_ | ~new_n535_;
  assign new_n537_ = u0 & r4;
  assign new_n538_ = t0 & w4;
  assign new_n539_ = s0 & d4;
  assign new_n540_ = r0 & h4;
  assign new_n541_ = ~new_n537_ & ~new_n538_;
  assign new_n542_ = ~new_n539_ & ~new_n540_;
  assign new_n543_ = new_n541_ & new_n542_;
  assign new_n544_ = q0 & m4;
  assign new_n545_ = p0 & m5;
  assign new_n546_ = o0 & r5;
  assign new_n547_ = n0 & p5;
  assign new_n548_ = ~new_n544_ & ~new_n545_;
  assign new_n549_ = ~new_n546_ & ~new_n547_;
  assign new_n550_ = new_n548_ & new_n549_;
  assign new_n551_ = m0 & f3;
  assign new_n552_ = l0 & m3;
  assign new_n553_ = k0 & q3;
  assign new_n554_ = ~new_n551_ & ~new_n552_;
  assign new_n555_ = ~new_n553_ & new_n554_;
  assign new_n556_ = new_n543_ & new_n550_;
  assign a6 = ~new_n555_ | ~new_n556_;
  assign new_n558_ = u0 & l5;
  assign new_n559_ = t0 & v4;
  assign new_n560_ = ~j5 & k5;
  assign new_n561_ = ~d5 & ~e5;
  assign new_n562_ = a5 & ~b5;
  assign new_n563_ = ~i5 & o5;
  assign new_n564_ = ~g5 & ~o5;
  assign new_n565_ = ~new_n563_ & ~new_n564_;
  assign new_n566_ = g5 & ~new_n565_;
  assign new_n567_ = ~new_n562_ & new_n566_;
  assign new_n568_ = new_n562_ & ~new_n566_;
  assign new_n569_ = ~new_n567_ & ~new_n568_;
  assign new_n570_ = new_n561_ & ~new_n569_;
  assign new_n571_ = new_n566_ & new_n570_;
  assign new_n572_ = ~d5 & ~new_n571_;
  assign new_n573_ = new_n562_ & ~new_n569_;
  assign new_n574_ = new_n561_ & new_n573_;
  assign j10 = e5 | new_n574_;
  assign new_n576_ = ~c5 & ~j10;
  assign new_n577_ = ~t4 & ~u4;
  assign new_n578_ = ~v4 & new_n577_;
  assign new_n579_ = ~w4 & new_n578_;
  assign new_n580_ = ~x4 & new_n579_;
  assign new_n581_ = ~y4 & new_n580_;
  assign new_n582_ = ~s4 & new_n581_;
  assign new_n583_ = ~z4 & new_n582_;
  assign new_n584_ = ~r4 & new_n583_;
  assign new_n585_ = new_n572_ & new_n576_;
  assign new_n586_ = new_n584_ & ~new_n585_;
  assign new_n587_ = ~l5 & ~m5;
  assign new_n588_ = ~n5 & new_n587_;
  assign v10 = z | new_n588_;
  assign new_n590_ = new_n586_ & v10;
  assign new_n591_ = ~r4 & r5;
  assign new_n592_ = new_n560_ & ~new_n591_;
  assign new_n593_ = ~new_n590_ & ~new_n592_;
  assign new_n594_ = ~d0 & new_n593_;
  assign new_n595_ = s0 & new_n594_;
  assign new_n596_ = r0 & g4;
  assign new_n597_ = ~new_n558_ & ~new_n559_;
  assign new_n598_ = ~new_n595_ & ~new_n596_;
  assign new_n599_ = new_n597_ & new_n598_;
  assign new_n600_ = ~j0 & q5;
  assign new_n601_ = d4 & e4;
  assign new_n602_ = f4 & new_n601_;
  assign new_n603_ = ~new_n600_ & ~new_n602_;
  assign new_n604_ = i4 & ~new_n603_;
  assign new_n605_ = ~j0 & ~p5;
  assign new_n606_ = ~new_n604_ & new_n605_;
  assign new_n607_ = g4 & ~new_n606_;
  assign new_n608_ = p4 & new_n607_;
  assign new_n609_ = q0 & new_n608_;
  assign new_n610_ = p0 & n5;
  assign new_n611_ = ~l5 & m5;
  assign new_n612_ = ~n5 & new_n611_;
  assign new_n613_ = ~z & new_n612_;
  assign new_n614_ = ~z & ~new_n613_;
  assign new_n615_ = o0 & ~new_n614_;
  assign new_n616_ = n0 & q5;
  assign new_n617_ = ~new_n609_ & ~new_n610_;
  assign new_n618_ = ~new_n615_ & ~new_n616_;
  assign new_n619_ = new_n617_ & new_n618_;
  assign new_n620_ = p3 & q3;
  assign new_n621_ = s3 & t3;
  assign new_n622_ = r3 & new_n621_;
  assign new_n623_ = new_n620_ & new_n622_;
  assign new_n624_ = m0 & new_n623_;
  assign new_n625_ = l0 & l3;
  assign new_n626_ = n3 & ~o3;
  assign new_n627_ = ~p3 & new_n626_;
  assign new_n628_ = ~q3 & ~r3;
  assign new_n629_ = ~s3 & ~t3;
  assign new_n630_ = new_n628_ & new_n629_;
  assign new_n631_ = new_n627_ & new_n630_;
  assign new_n632_ = k0 & new_n631_;
  assign new_n633_ = ~new_n624_ & ~new_n625_;
  assign new_n634_ = ~new_n632_ & new_n633_;
  assign new_n635_ = new_n599_ & new_n619_;
  assign b6 = ~new_n634_ | ~new_n635_;
  assign new_n637_ = r1 & new_n425_;
  assign new_n638_ = new_n412_ & ~new_n637_;
  assign new_n639_ = new_n408_ & new_n638_;
  assign new_n640_ = ~v0 & new_n639_;
  assign new_n641_ = v0 & ~new_n639_;
  assign new_n642_ = ~new_n640_ & ~new_n641_;
  assign new_n643_ = new_n421_ & v6;
  assign new_n644_ = v0 & new_n637_;
  assign new_n645_ = ~m1 & n1;
  assign new_n646_ = ~b & l1;
  assign new_n647_ = new_n645_ & new_n646_;
  assign new_n648_ = ~new_n643_ & ~new_n644_;
  assign new_n649_ = ~b & ~new_n647_;
  assign new_n650_ = new_n648_ & new_n649_;
  assign c6 = new_n642_ & new_n650_;
  assign new_n652_ = ~w0 & ~new_n641_;
  assign new_n653_ = w0 & new_n641_;
  assign new_n654_ = ~new_n652_ & ~new_n653_;
  assign d6 = new_n650_ & new_n654_;
  assign new_n656_ = v0 & w0;
  assign new_n657_ = ~new_n639_ & new_n656_;
  assign new_n658_ = ~x0 & ~new_n657_;
  assign new_n659_ = x0 & new_n657_;
  assign new_n660_ = ~new_n658_ & ~new_n659_;
  assign e6 = new_n650_ & new_n660_;
  assign new_n662_ = x0 & new_n656_;
  assign new_n663_ = ~new_n639_ & new_n662_;
  assign new_n664_ = ~y0 & ~new_n663_;
  assign new_n665_ = y0 & new_n663_;
  assign new_n666_ = ~new_n664_ & ~new_n665_;
  assign f6 = new_n650_ & new_n666_;
  assign new_n668_ = x0 & y0;
  assign new_n669_ = new_n656_ & new_n668_;
  assign new_n670_ = ~new_n639_ & new_n669_;
  assign new_n671_ = ~z0 & ~new_n670_;
  assign new_n672_ = z0 & new_n670_;
  assign new_n673_ = ~new_n671_ & ~new_n672_;
  assign g6 = new_n650_ & new_n673_;
  assign new_n675_ = z0 & new_n669_;
  assign new_n676_ = ~new_n639_ & new_n675_;
  assign new_n677_ = ~a1 & ~new_n676_;
  assign new_n678_ = a1 & new_n676_;
  assign new_n679_ = ~new_n677_ & ~new_n678_;
  assign h6 = new_n650_ & new_n679_;
  assign new_n681_ = a1 & new_n675_;
  assign new_n682_ = ~new_n639_ & new_n681_;
  assign new_n683_ = ~b1 & ~new_n682_;
  assign new_n684_ = b1 & new_n682_;
  assign new_n685_ = ~new_n683_ & ~new_n684_;
  assign i6 = new_n650_ & new_n685_;
  assign new_n687_ = z0 & a1;
  assign new_n688_ = b1 & new_n687_;
  assign new_n689_ = new_n669_ & new_n688_;
  assign new_n690_ = ~new_n639_ & new_n689_;
  assign new_n691_ = ~c1 & ~new_n690_;
  assign new_n692_ = c1 & new_n690_;
  assign new_n693_ = ~new_n691_ & ~new_n692_;
  assign j6 = new_n650_ & new_n693_;
  assign new_n695_ = c1 & ~new_n639_;
  assign new_n696_ = new_n689_ & new_n695_;
  assign new_n697_ = d1 & new_n696_;
  assign new_n698_ = ~d1 & ~new_n696_;
  assign new_n699_ = ~new_n697_ & ~new_n698_;
  assign k6 = new_n650_ & new_n699_;
  assign new_n701_ = h1 & new_n398_;
  assign new_n702_ = new_n649_ & ~new_n701_;
  assign new_n703_ = h1 & new_n702_;
  assign o6 = new_n407_ | new_n703_;
  assign new_n705_ = i1 & new_n402_;
  assign new_n706_ = new_n649_ & ~new_n705_;
  assign new_n707_ = i1 & new_n706_;
  assign p6 = new_n410_ | new_n707_;
  assign new_n709_ = j1 & new_n447_;
  assign new_n710_ = ~j1 & ~new_n447_;
  assign new_n711_ = ~new_n709_ & ~new_n710_;
  assign new_n712_ = ~b & new_n711_;
  assign new_n713_ = l1 & ~m1;
  assign new_n714_ = ~n1 & new_n713_;
  assign new_n715_ = ~b & new_n714_;
  assign new_n716_ = ~new_n647_ & ~new_n715_;
  assign q6 = new_n712_ | ~new_n716_;
  assign new_n718_ = new_n398_ & ~new_n468_;
  assign new_n719_ = new_n460_ & new_n718_;
  assign new_n720_ = new_n425_ & ~new_n719_;
  assign new_n721_ = new_n398_ & new_n452_;
  assign new_n722_ = ~new_n715_ & ~new_n720_;
  assign new_n723_ = ~new_n721_ & new_n722_;
  assign s6 = ~b & ~new_n723_;
  assign new_n725_ = r1 & ~new_n697_;
  assign new_n726_ = r1 & new_n697_;
  assign new_n727_ = ~d1 & ~new_n726_;
  assign new_n728_ = ~new_n725_ & ~new_n727_;
  assign new_n729_ = ~c & ~new_n728_;
  assign new_n730_ = v6 & ~new_n729_;
  assign new_n731_ = new_n425_ & new_n468_;
  assign new_n732_ = ~new_n730_ & ~new_n731_;
  assign new_n733_ = n1 & new_n426_;
  assign new_n734_ = ~b & new_n733_;
  assign new_n735_ = ~new_n452_ & new_n732_;
  assign new_n736_ = ~new_n734_ & new_n735_;
  assign new_n737_ = n1 & new_n423_;
  assign new_n738_ = ~b & new_n737_;
  assign new_n739_ = m1 & n1;
  assign new_n740_ = ~new_n398_ & ~new_n468_;
  assign new_n741_ = new_n425_ & new_n740_;
  assign new_n742_ = ~new_n739_ & ~new_n741_;
  assign new_n743_ = ~new_n738_ & new_n742_;
  assign new_n744_ = new_n736_ & new_n743_;
  assign t6 = ~b & ~new_n744_;
  assign new_n746_ = ~new_n731_ & ~new_n734_;
  assign new_n747_ = ~new_n715_ & new_n746_;
  assign new_n748_ = new_n398_ & new_n425_;
  assign new_n749_ = new_n460_ & ~new_n468_;
  assign new_n750_ = new_n748_ & new_n749_;
  assign new_n751_ = ~new_n738_ & ~new_n750_;
  assign new_n752_ = new_n747_ & new_n751_;
  assign u6 = ~b & ~new_n752_;
  assign new_n754_ = q1 & r1;
  assign new_n755_ = ~p1 & ~new_n754_;
  assign new_n756_ = ~q1 & ~r1;
  assign new_n757_ = ~new_n755_ & ~new_n756_;
  assign new_n758_ = ~p1 & new_n756_;
  assign new_n759_ = ~b & ~new_n758_;
  assign new_n760_ = ~new_n757_ & new_n759_;
  assign new_n761_ = ~e & ~new_n738_;
  assign new_n762_ = ~d & ~new_n734_;
  assign new_n763_ = q1 & ~new_n762_;
  assign new_n764_ = r1 & ~new_n761_;
  assign new_n765_ = ~p1 & ~new_n764_;
  assign new_n766_ = ~r1 & ~new_n761_;
  assign new_n767_ = ~new_n765_ & ~new_n766_;
  assign new_n768_ = ~new_n763_ & ~new_n767_;
  assign new_n769_ = ~new_n762_ & ~new_n764_;
  assign new_n770_ = ~q1 & new_n769_;
  assign new_n771_ = ~new_n768_ & ~new_n770_;
  assign w6 = ~new_n760_ | new_n771_;
  assign new_n773_ = r1 & ~new_n762_;
  assign new_n774_ = q1 & new_n761_;
  assign new_n775_ = ~p1 & ~new_n774_;
  assign new_n776_ = ~q1 & new_n761_;
  assign new_n777_ = ~new_n775_ & ~new_n776_;
  assign new_n778_ = ~new_n773_ & ~new_n777_;
  assign new_n779_ = p1 & ~new_n761_;
  assign new_n780_ = ~new_n762_ & ~new_n779_;
  assign new_n781_ = ~r1 & new_n780_;
  assign new_n782_ = ~new_n778_ & ~new_n781_;
  assign x6 = new_n760_ & new_n782_;
  assign new_n784_ = p1 & ~new_n762_;
  assign new_n785_ = ~r1 & new_n761_;
  assign new_n786_ = r1 & new_n761_;
  assign new_n787_ = ~q1 & ~new_n786_;
  assign new_n788_ = ~new_n785_ & ~new_n787_;
  assign new_n789_ = ~new_n784_ & ~new_n788_;
  assign new_n790_ = q1 & ~new_n761_;
  assign new_n791_ = ~new_n762_ & ~new_n790_;
  assign new_n792_ = ~p1 & new_n791_;
  assign new_n793_ = ~new_n789_ & ~new_n792_;
  assign y6 = new_n760_ & new_n793_;
  assign new_n795_ = v0 & new_n419_;
  assign new_n796_ = v6 & new_n795_;
  assign new_n797_ = ~new_n715_ & ~new_n796_;
  assign new_n798_ = ~v0 & w0;
  assign new_n799_ = q1 & new_n414_;
  assign new_n800_ = r1 & new_n417_;
  assign new_n801_ = p1 & new_n413_;
  assign new_n802_ = ~new_n800_ & ~new_n801_;
  assign new_n803_ = ~new_n799_ & new_n802_;
  assign new_n804_ = new_n798_ & ~new_n803_;
  assign new_n805_ = v6 & new_n804_;
  assign new_n806_ = ~h & ~new_n805_;
  assign new_n807_ = ~s1 & ~new_n806_;
  assign new_n808_ = s1 & new_n806_;
  assign new_n809_ = ~new_n807_ & ~new_n808_;
  assign new_n810_ = new_n797_ & new_n809_;
  assign new_n811_ = new_n797_ & ~new_n809_;
  assign new_n812_ = ~w2 & ~new_n811_;
  assign new_n813_ = ~new_n810_ & ~new_n812_;
  assign z6 = ~b & new_n813_;
  assign new_n815_ = ~i & new_n412_;
  assign new_n816_ = ~s1 & ~new_n815_;
  assign new_n817_ = s1 & new_n815_;
  assign new_n818_ = ~new_n816_ & ~new_n817_;
  assign new_n819_ = ~new_n806_ & new_n818_;
  assign new_n820_ = ~t1 & new_n819_;
  assign new_n821_ = t1 & ~new_n819_;
  assign new_n822_ = ~new_n820_ & ~new_n821_;
  assign new_n823_ = new_n797_ & new_n822_;
  assign new_n824_ = new_n797_ & ~new_n822_;
  assign new_n825_ = ~x2 & ~new_n824_;
  assign new_n826_ = ~new_n823_ & ~new_n825_;
  assign a7 = ~b & new_n826_;
  assign new_n828_ = ~s1 & ~t1;
  assign new_n829_ = s1 & t1;
  assign new_n830_ = ~new_n815_ & new_n829_;
  assign new_n831_ = ~new_n828_ & ~new_n830_;
  assign new_n832_ = ~new_n815_ & ~new_n829_;
  assign new_n833_ = ~new_n831_ & ~new_n832_;
  assign new_n834_ = ~new_n806_ & new_n833_;
  assign new_n835_ = ~u1 & new_n834_;
  assign new_n836_ = u1 & ~new_n834_;
  assign new_n837_ = ~new_n835_ & ~new_n836_;
  assign new_n838_ = new_n797_ & new_n837_;
  assign new_n839_ = new_n797_ & ~new_n837_;
  assign new_n840_ = ~y2 & ~new_n839_;
  assign new_n841_ = ~new_n838_ & ~new_n840_;
  assign b7 = ~b & new_n841_;
  assign new_n843_ = ~u1 & new_n828_;
  assign new_n844_ = ~k & ~new_n843_;
  assign new_n845_ = u1 & new_n829_;
  assign new_n846_ = ~k & ~new_n845_;
  assign new_n847_ = ~new_n815_ & ~new_n846_;
  assign new_n848_ = new_n844_ & ~new_n847_;
  assign new_n849_ = ~new_n815_ & new_n846_;
  assign new_n850_ = ~new_n848_ & ~new_n849_;
  assign new_n851_ = ~new_n806_ & new_n850_;
  assign new_n852_ = ~v1 & new_n851_;
  assign new_n853_ = v1 & ~new_n851_;
  assign new_n854_ = ~new_n852_ & ~new_n853_;
  assign new_n855_ = new_n797_ & new_n854_;
  assign new_n856_ = new_n797_ & ~new_n854_;
  assign new_n857_ = ~z2 & ~new_n856_;
  assign new_n858_ = ~new_n855_ & ~new_n857_;
  assign c7 = b | new_n858_;
  assign new_n860_ = ~v1 & ~new_n844_;
  assign new_n861_ = v1 & ~new_n846_;
  assign new_n862_ = ~new_n815_ & new_n861_;
  assign new_n863_ = ~new_n860_ & ~new_n862_;
  assign new_n864_ = ~new_n815_ & ~new_n861_;
  assign new_n865_ = ~new_n863_ & ~new_n864_;
  assign new_n866_ = ~new_n806_ & new_n865_;
  assign new_n867_ = ~w1 & new_n866_;
  assign new_n868_ = w1 & ~new_n866_;
  assign new_n869_ = ~new_n867_ & ~new_n868_;
  assign new_n870_ = new_n797_ & new_n869_;
  assign new_n871_ = new_n797_ & ~new_n869_;
  assign new_n872_ = ~a3 & ~new_n871_;
  assign new_n873_ = ~new_n870_ & ~new_n872_;
  assign d7 = b | new_n873_;
  assign new_n875_ = ~w1 & new_n860_;
  assign new_n876_ = v1 & w1;
  assign new_n877_ = ~new_n846_ & new_n876_;
  assign new_n878_ = ~new_n815_ & new_n877_;
  assign new_n879_ = ~new_n875_ & ~new_n878_;
  assign new_n880_ = ~new_n815_ & ~new_n877_;
  assign new_n881_ = ~new_n879_ & ~new_n880_;
  assign new_n882_ = ~new_n806_ & new_n881_;
  assign new_n883_ = ~x1 & new_n882_;
  assign new_n884_ = x1 & ~new_n882_;
  assign new_n885_ = ~new_n883_ & ~new_n884_;
  assign new_n886_ = new_n797_ & new_n885_;
  assign new_n887_ = new_n797_ & ~new_n885_;
  assign new_n888_ = ~b3 & ~new_n887_;
  assign new_n889_ = ~new_n886_ & ~new_n888_;
  assign e7 = b | new_n889_;
  assign new_n891_ = ~w1 & ~x1;
  assign new_n892_ = new_n860_ & new_n891_;
  assign new_n893_ = ~k & ~new_n892_;
  assign new_n894_ = w1 & x1;
  assign new_n895_ = new_n861_ & new_n894_;
  assign new_n896_ = ~k & ~new_n895_;
  assign new_n897_ = ~new_n815_ & ~new_n896_;
  assign new_n898_ = new_n893_ & ~new_n897_;
  assign new_n899_ = ~new_n815_ & new_n896_;
  assign new_n900_ = ~new_n898_ & ~new_n899_;
  assign new_n901_ = ~new_n806_ & new_n900_;
  assign new_n902_ = ~y1 & new_n901_;
  assign new_n903_ = y1 & ~new_n901_;
  assign new_n904_ = ~new_n902_ & ~new_n903_;
  assign new_n905_ = new_n797_ & new_n904_;
  assign new_n906_ = new_n797_ & ~new_n904_;
  assign new_n907_ = ~c3 & ~new_n906_;
  assign new_n908_ = ~new_n905_ & ~new_n907_;
  assign f7 = ~b & new_n908_;
  assign new_n910_ = ~y1 & ~new_n893_;
  assign new_n911_ = y1 & ~new_n896_;
  assign new_n912_ = ~new_n815_ & new_n911_;
  assign new_n913_ = ~new_n910_ & ~new_n912_;
  assign new_n914_ = ~new_n815_ & ~new_n911_;
  assign new_n915_ = ~new_n913_ & ~new_n914_;
  assign new_n916_ = ~new_n806_ & new_n915_;
  assign new_n917_ = ~z1 & new_n916_;
  assign new_n918_ = z1 & ~new_n916_;
  assign new_n919_ = ~new_n917_ & ~new_n918_;
  assign new_n920_ = new_n797_ & new_n919_;
  assign new_n921_ = new_n797_ & ~new_n919_;
  assign new_n922_ = ~d3 & ~new_n921_;
  assign new_n923_ = ~new_n920_ & ~new_n922_;
  assign g7 = b | new_n923_;
  assign new_n925_ = ~z1 & new_n910_;
  assign new_n926_ = y1 & z1;
  assign new_n927_ = ~new_n896_ & new_n926_;
  assign new_n928_ = ~new_n815_ & new_n927_;
  assign new_n929_ = ~new_n925_ & ~new_n928_;
  assign new_n930_ = ~new_n815_ & ~new_n927_;
  assign new_n931_ = ~new_n929_ & ~new_n930_;
  assign new_n932_ = ~new_n806_ & new_n931_;
  assign new_n933_ = ~a2 & new_n932_;
  assign new_n934_ = a2 & ~new_n932_;
  assign new_n935_ = ~new_n933_ & ~new_n934_;
  assign new_n936_ = new_n797_ & new_n935_;
  assign new_n937_ = new_n797_ & ~new_n935_;
  assign new_n938_ = ~e3 & ~new_n937_;
  assign new_n939_ = ~new_n936_ & ~new_n938_;
  assign h7 = b | new_n939_;
  assign i7 = b | ~b2;
  assign new_n942_ = ~b2 & ~c2;
  assign new_n943_ = ~new_n440_ & ~new_n942_;
  assign j7 = b | new_n943_;
  assign new_n945_ = ~d2 & ~new_n440_;
  assign new_n946_ = ~new_n441_ & ~new_n945_;
  assign k7 = b | new_n946_;
  assign new_n948_ = ~new_n447_ & ~new_n647_;
  assign new_n949_ = ~e2 & ~new_n445_;
  assign new_n950_ = e2 & new_n445_;
  assign new_n951_ = ~new_n949_ & ~new_n950_;
  assign new_n952_ = new_n948_ & ~new_n951_;
  assign new_n953_ = ~s1 & ~new_n952_;
  assign new_n954_ = new_n948_ & new_n951_;
  assign new_n955_ = ~new_n953_ & ~new_n954_;
  assign l7 = b | new_n955_;
  assign new_n957_ = ~f2 & new_n446_;
  assign new_n958_ = f2 & ~new_n446_;
  assign new_n959_ = ~new_n957_ & ~new_n958_;
  assign new_n960_ = new_n948_ & ~new_n959_;
  assign new_n961_ = ~t1 & ~new_n960_;
  assign new_n962_ = new_n948_ & new_n959_;
  assign new_n963_ = ~new_n961_ & ~new_n962_;
  assign m7 = b | new_n963_;
  assign new_n965_ = ~g2 & new_n442_;
  assign new_n966_ = ~new_n443_ & ~new_n965_;
  assign n7 = b | new_n966_;
  assign new_n968_ = f2 & new_n446_;
  assign new_n969_ = ~h2 & new_n968_;
  assign new_n970_ = h2 & ~new_n968_;
  assign new_n971_ = ~new_n969_ & ~new_n970_;
  assign new_n972_ = new_n948_ & ~new_n971_;
  assign new_n973_ = ~u1 & ~new_n972_;
  assign new_n974_ = new_n948_ & new_n971_;
  assign new_n975_ = ~new_n973_ & ~new_n974_;
  assign o7 = b | new_n975_;
  assign new_n977_ = f2 & h2;
  assign new_n978_ = new_n446_ & new_n977_;
  assign new_n979_ = ~i2 & new_n978_;
  assign new_n980_ = i2 & ~new_n978_;
  assign new_n981_ = ~new_n979_ & ~new_n980_;
  assign new_n982_ = new_n948_ & ~new_n981_;
  assign new_n983_ = ~v1 & ~new_n982_;
  assign new_n984_ = new_n948_ & new_n981_;
  assign new_n985_ = ~new_n983_ & ~new_n984_;
  assign p7 = b | new_n985_;
  assign new_n987_ = i2 & new_n978_;
  assign new_n988_ = ~j2 & new_n987_;
  assign new_n989_ = j2 & ~new_n987_;
  assign new_n990_ = ~new_n988_ & ~new_n989_;
  assign new_n991_ = new_n948_ & ~new_n990_;
  assign new_n992_ = ~w1 & ~new_n991_;
  assign new_n993_ = new_n948_ & new_n990_;
  assign new_n994_ = ~new_n992_ & ~new_n993_;
  assign q7 = b | new_n994_;
  assign new_n996_ = j2 & new_n987_;
  assign new_n997_ = ~l & ~new_n996_;
  assign new_n998_ = ~k2 & ~new_n997_;
  assign new_n999_ = k2 & new_n997_;
  assign new_n1000_ = ~new_n998_ & ~new_n999_;
  assign new_n1001_ = new_n948_ & ~new_n1000_;
  assign new_n1002_ = ~x1 & ~new_n1001_;
  assign new_n1003_ = new_n948_ & new_n1000_;
  assign new_n1004_ = ~new_n1002_ & ~new_n1003_;
  assign r7 = b | new_n1004_;
  assign new_n1006_ = k2 & ~new_n997_;
  assign new_n1007_ = ~l2 & new_n1006_;
  assign new_n1008_ = l2 & ~new_n1006_;
  assign new_n1009_ = ~new_n1007_ & ~new_n1008_;
  assign new_n1010_ = new_n948_ & ~new_n1009_;
  assign new_n1011_ = ~y1 & ~new_n1010_;
  assign new_n1012_ = new_n948_ & new_n1009_;
  assign new_n1013_ = ~new_n1011_ & ~new_n1012_;
  assign s7 = b | new_n1013_;
  assign new_n1015_ = k2 & l2;
  assign new_n1016_ = ~new_n997_ & new_n1015_;
  assign new_n1017_ = ~m2 & new_n1016_;
  assign new_n1018_ = m2 & ~new_n1016_;
  assign new_n1019_ = ~new_n1017_ & ~new_n1018_;
  assign new_n1020_ = new_n948_ & ~new_n1019_;
  assign new_n1021_ = ~z1 & ~new_n1020_;
  assign new_n1022_ = new_n948_ & new_n1019_;
  assign new_n1023_ = ~new_n1021_ & ~new_n1022_;
  assign t7 = b | new_n1023_;
  assign new_n1025_ = m2 & o2;
  assign new_n1026_ = l2 & new_n1025_;
  assign new_n1027_ = j2 & k2;
  assign new_n1028_ = i2 & new_n1027_;
  assign new_n1029_ = ~b & ~new_n948_;
  assign new_n1030_ = new_n1026_ & new_n1028_;
  assign new_n1031_ = new_n977_ & new_n1030_;
  assign u7 = ~new_n1029_ & new_n1031_;
  assign new_n1033_ = m2 & new_n1016_;
  assign new_n1034_ = ~o2 & new_n1033_;
  assign new_n1035_ = o2 & ~new_n1033_;
  assign new_n1036_ = ~new_n1034_ & ~new_n1035_;
  assign new_n1037_ = new_n948_ & ~new_n1036_;
  assign new_n1038_ = ~a2 & ~new_n1037_;
  assign new_n1039_ = new_n948_ & new_n1036_;
  assign new_n1040_ = ~new_n1038_ & ~new_n1039_;
  assign v7 = b | new_n1040_;
  assign new_n1042_ = ~p2 & ~new_n709_;
  assign new_n1043_ = ~a & ~new_n1042_;
  assign new_n1044_ = p2 & ~new_n709_;
  assign w7 = new_n1043_ | new_n1044_;
  assign new_n1046_ = ~q2 & new_n433_;
  assign new_n1047_ = q2 & ~new_n433_;
  assign new_n1048_ = ~new_n1046_ & ~new_n1047_;
  assign x7 = new_n453_ & new_n1048_;
  assign new_n1050_ = ~new_n412_ & v6;
  assign new_n1051_ = ~g & ~new_n1050_;
  assign new_n1052_ = ~q2 & ~new_n1051_;
  assign new_n1053_ = q2 & new_n1051_;
  assign new_n1054_ = ~new_n1052_ & ~new_n1053_;
  assign new_n1055_ = ~new_n433_ & new_n1054_;
  assign new_n1056_ = ~r2 & ~new_n1055_;
  assign new_n1057_ = r2 & new_n1055_;
  assign new_n1058_ = ~new_n1056_ & ~new_n1057_;
  assign y7 = new_n453_ & new_n1058_;
  assign new_n1060_ = q1 & new_n425_;
  assign new_n1061_ = ~j & new_n1060_;
  assign new_n1062_ = ~q2 & ~r2;
  assign new_n1063_ = ~new_n1061_ & ~new_n1062_;
  assign new_n1064_ = q2 & r2;
  assign new_n1065_ = ~new_n1061_ & ~new_n1064_;
  assign new_n1066_ = ~new_n1051_ & ~new_n1065_;
  assign new_n1067_ = new_n1063_ & ~new_n1066_;
  assign new_n1068_ = ~new_n1051_ & new_n1065_;
  assign new_n1069_ = ~new_n1067_ & ~new_n1068_;
  assign new_n1070_ = ~new_n433_ & new_n1069_;
  assign new_n1071_ = ~s2 & ~new_n1070_;
  assign new_n1072_ = s2 & new_n1070_;
  assign new_n1073_ = ~new_n1071_ & ~new_n1072_;
  assign z7 = new_n453_ & new_n1073_;
  assign new_n1075_ = p1 & new_n425_;
  assign new_n1076_ = ~j & new_n1075_;
  assign new_n1077_ = ~s2 & ~new_n1063_;
  assign new_n1078_ = ~new_n1076_ & ~new_n1077_;
  assign new_n1079_ = s2 & ~new_n1065_;
  assign new_n1080_ = ~new_n1076_ & ~new_n1079_;
  assign new_n1081_ = new_n1051_ & ~new_n1078_;
  assign new_n1082_ = ~new_n1051_ & ~new_n1080_;
  assign new_n1083_ = ~new_n1081_ & ~new_n1082_;
  assign new_n1084_ = ~new_n433_ & ~new_n1083_;
  assign new_n1085_ = ~t2 & new_n1084_;
  assign new_n1086_ = t2 & ~new_n1084_;
  assign new_n1087_ = ~new_n1085_ & ~new_n1086_;
  assign new_n1088_ = new_n453_ & ~new_n1087_;
  assign new_n1089_ = ~new_n453_ & ~new_n1051_;
  assign a8 = new_n1088_ | new_n1089_;
  assign new_n1091_ = ~w2 & ~x2;
  assign new_n1092_ = ~y2 & ~z2;
  assign new_n1093_ = new_n1091_ & new_n1092_;
  assign new_n1094_ = new_n453_ & ~new_n1093_;
  assign new_n1095_ = new_n1051_ & ~new_n1094_;
  assign new_n1096_ = new_n453_ & new_n1093_;
  assign b8 = new_n1095_ | new_n1096_;
  assign new_n1098_ = w2 & x2;
  assign new_n1099_ = y2 & z2;
  assign new_n1100_ = new_n1098_ & new_n1099_;
  assign c8 = new_n453_ & new_n1100_;
  assign new_n1102_ = ~t2 & ~new_n1078_;
  assign new_n1103_ = ~j & ~new_n1102_;
  assign new_n1104_ = t2 & ~new_n1080_;
  assign new_n1105_ = ~j & ~new_n1104_;
  assign new_n1106_ = ~new_n1051_ & ~new_n1105_;
  assign new_n1107_ = new_n1103_ & ~new_n1106_;
  assign new_n1108_ = ~new_n1051_ & new_n1105_;
  assign new_n1109_ = ~new_n1107_ & ~new_n1108_;
  assign new_n1110_ = ~new_n433_ & new_n1109_;
  assign new_n1111_ = ~w2 & ~new_n1110_;
  assign new_n1112_ = w2 & new_n1110_;
  assign new_n1113_ = ~new_n1111_ & ~new_n1112_;
  assign d8 = new_n453_ & new_n1113_;
  assign new_n1115_ = ~w2 & ~new_n1103_;
  assign new_n1116_ = w2 & ~new_n1105_;
  assign new_n1117_ = ~new_n1051_ & new_n1116_;
  assign new_n1118_ = ~new_n1115_ & ~new_n1117_;
  assign new_n1119_ = ~new_n1051_ & ~new_n1116_;
  assign new_n1120_ = ~new_n1118_ & ~new_n1119_;
  assign new_n1121_ = ~new_n433_ & new_n1120_;
  assign new_n1122_ = ~x2 & ~new_n1121_;
  assign new_n1123_ = x2 & new_n1121_;
  assign new_n1124_ = ~new_n1122_ & ~new_n1123_;
  assign e8 = new_n453_ & new_n1124_;
  assign new_n1126_ = ~x2 & new_n1115_;
  assign new_n1127_ = new_n1098_ & ~new_n1105_;
  assign new_n1128_ = ~new_n1051_ & new_n1127_;
  assign new_n1129_ = ~new_n1126_ & ~new_n1128_;
  assign new_n1130_ = ~new_n1051_ & ~new_n1127_;
  assign new_n1131_ = ~new_n1129_ & ~new_n1130_;
  assign new_n1132_ = ~new_n433_ & new_n1131_;
  assign new_n1133_ = ~y2 & ~new_n1132_;
  assign new_n1134_ = y2 & new_n1132_;
  assign new_n1135_ = ~new_n1133_ & ~new_n1134_;
  assign f8 = new_n453_ & new_n1135_;
  assign new_n1137_ = ~y2 & new_n1126_;
  assign new_n1138_ = x2 & y2;
  assign new_n1139_ = w2 & new_n1138_;
  assign new_n1140_ = ~new_n1105_ & new_n1139_;
  assign new_n1141_ = ~new_n1051_ & new_n1140_;
  assign new_n1142_ = ~new_n1137_ & ~new_n1141_;
  assign new_n1143_ = ~new_n1051_ & ~new_n1140_;
  assign new_n1144_ = ~new_n1142_ & ~new_n1143_;
  assign new_n1145_ = ~new_n433_ & new_n1144_;
  assign new_n1146_ = ~z2 & new_n1145_;
  assign new_n1147_ = z2 & ~new_n1145_;
  assign new_n1148_ = ~new_n1146_ & ~new_n1147_;
  assign new_n1149_ = new_n453_ & ~new_n1148_;
  assign g8 = new_n1089_ | new_n1149_;
  assign new_n1151_ = u2 & ~new_n1103_;
  assign new_n1152_ = v2 & ~new_n1105_;
  assign new_n1153_ = ~new_n1051_ & new_n1152_;
  assign new_n1154_ = ~new_n1151_ & ~new_n1153_;
  assign new_n1155_ = ~new_n1051_ & ~new_n1152_;
  assign new_n1156_ = ~new_n1154_ & ~new_n1155_;
  assign new_n1157_ = ~new_n433_ & new_n1156_;
  assign new_n1158_ = ~a3 & new_n1157_;
  assign new_n1159_ = a3 & ~new_n1157_;
  assign new_n1160_ = ~new_n1158_ & ~new_n1159_;
  assign new_n1161_ = new_n453_ & ~new_n1160_;
  assign h8 = new_n1089_ | new_n1161_;
  assign new_n1163_ = ~a3 & new_n1151_;
  assign new_n1164_ = ~j & ~new_n1163_;
  assign new_n1165_ = a3 & new_n1152_;
  assign new_n1166_ = ~j & ~new_n1165_;
  assign new_n1167_ = ~new_n1051_ & ~new_n1166_;
  assign new_n1168_ = new_n1164_ & ~new_n1167_;
  assign new_n1169_ = ~new_n1051_ & new_n1166_;
  assign new_n1170_ = ~new_n1168_ & ~new_n1169_;
  assign new_n1171_ = ~new_n433_ & new_n1170_;
  assign new_n1172_ = ~b3 & new_n1171_;
  assign new_n1173_ = b3 & ~new_n1171_;
  assign new_n1174_ = ~new_n1172_ & ~new_n1173_;
  assign new_n1175_ = new_n453_ & ~new_n1174_;
  assign i8 = new_n1089_ | new_n1175_;
  assign new_n1177_ = ~b3 & ~new_n1164_;
  assign new_n1178_ = b3 & ~new_n1166_;
  assign new_n1179_ = ~new_n1051_ & ~new_n1178_;
  assign new_n1180_ = ~new_n1051_ & new_n1178_;
  assign new_n1181_ = ~new_n1177_ & ~new_n1180_;
  assign new_n1182_ = ~new_n1179_ & ~new_n1181_;
  assign new_n1183_ = ~new_n433_ & new_n1182_;
  assign new_n1184_ = ~c3 & ~new_n1183_;
  assign new_n1185_ = c3 & new_n1183_;
  assign new_n1186_ = ~new_n1184_ & ~new_n1185_;
  assign j8 = new_n453_ & new_n1186_;
  assign new_n1188_ = ~c3 & new_n1177_;
  assign new_n1189_ = c3 & new_n1178_;
  assign new_n1190_ = ~new_n1051_ & new_n1189_;
  assign new_n1191_ = ~new_n1188_ & ~new_n1190_;
  assign new_n1192_ = ~new_n1051_ & ~new_n1189_;
  assign new_n1193_ = ~new_n1191_ & ~new_n1192_;
  assign new_n1194_ = ~new_n433_ & new_n1193_;
  assign new_n1195_ = ~d3 & new_n1194_;
  assign new_n1196_ = d3 & ~new_n1194_;
  assign new_n1197_ = ~new_n1195_ & ~new_n1196_;
  assign new_n1198_ = new_n453_ & ~new_n1197_;
  assign k8 = new_n1089_ | new_n1198_;
  assign new_n1200_ = ~d3 & new_n1188_;
  assign new_n1201_ = c3 & d3;
  assign new_n1202_ = new_n1178_ & new_n1201_;
  assign new_n1203_ = ~new_n1051_ & new_n1202_;
  assign new_n1204_ = ~new_n1200_ & ~new_n1203_;
  assign new_n1205_ = ~new_n1051_ & ~new_n1202_;
  assign new_n1206_ = ~new_n1204_ & ~new_n1205_;
  assign new_n1207_ = ~new_n433_ & new_n1206_;
  assign new_n1208_ = ~e3 & new_n1207_;
  assign new_n1209_ = e3 & ~new_n1207_;
  assign new_n1210_ = ~new_n1208_ & ~new_n1209_;
  assign new_n1211_ = new_n453_ & ~new_n1210_;
  assign l8 = new_n1089_ | new_n1211_;
  assign new_n1213_ = ~f3 & new_n594_;
  assign new_n1214_ = f3 & ~new_n594_;
  assign new_n1215_ = ~new_n1213_ & ~new_n1214_;
  assign m8 = new_n614_ & new_n1215_;
  assign new_n1217_ = ~new_n576_ & v10;
  assign new_n1218_ = ~e0 & ~new_n1217_;
  assign new_n1219_ = ~f3 & ~new_n1218_;
  assign new_n1220_ = f3 & new_n1218_;
  assign new_n1221_ = ~new_n1219_ & ~new_n1220_;
  assign new_n1222_ = ~new_n594_ & new_n1221_;
  assign new_n1223_ = ~g3 & ~new_n1222_;
  assign new_n1224_ = g3 & new_n1222_;
  assign new_n1225_ = ~new_n1223_ & ~new_n1224_;
  assign n8 = new_n614_ & new_n1225_;
  assign new_n1227_ = l5 & m5;
  assign new_n1228_ = ~z & ~n5;
  assign new_n1229_ = new_n1227_ & new_n1228_;
  assign new_n1230_ = q5 & new_n1229_;
  assign new_n1231_ = ~h0 & new_n1230_;
  assign new_n1232_ = ~f3 & ~g3;
  assign new_n1233_ = ~new_n1231_ & ~new_n1232_;
  assign new_n1234_ = f3 & g3;
  assign new_n1235_ = ~new_n1231_ & ~new_n1234_;
  assign new_n1236_ = ~new_n1218_ & new_n1235_;
  assign new_n1237_ = ~new_n1218_ & ~new_n1235_;
  assign new_n1238_ = new_n1233_ & ~new_n1237_;
  assign new_n1239_ = ~new_n1236_ & ~new_n1238_;
  assign new_n1240_ = ~new_n594_ & new_n1239_;
  assign new_n1241_ = ~h3 & ~new_n1240_;
  assign new_n1242_ = h3 & new_n1240_;
  assign new_n1243_ = ~new_n1241_ & ~new_n1242_;
  assign o8 = new_n614_ & new_n1243_;
  assign new_n1245_ = p5 & new_n1229_;
  assign new_n1246_ = ~h0 & new_n1245_;
  assign new_n1247_ = ~h3 & ~new_n1233_;
  assign new_n1248_ = ~new_n1246_ & ~new_n1247_;
  assign new_n1249_ = h3 & ~new_n1235_;
  assign new_n1250_ = ~new_n1246_ & ~new_n1249_;
  assign new_n1251_ = new_n1218_ & ~new_n1248_;
  assign new_n1252_ = ~new_n1218_ & ~new_n1250_;
  assign new_n1253_ = ~new_n1251_ & ~new_n1252_;
  assign new_n1254_ = ~new_n594_ & ~new_n1253_;
  assign new_n1255_ = ~i3 & new_n1254_;
  assign new_n1256_ = i3 & ~new_n1254_;
  assign new_n1257_ = ~new_n1255_ & ~new_n1256_;
  assign new_n1258_ = new_n614_ & ~new_n1257_;
  assign new_n1259_ = ~new_n614_ & ~new_n1218_;
  assign p8 = new_n1258_ | new_n1259_;
  assign new_n1261_ = ~l3 & ~m3;
  assign new_n1262_ = ~n3 & ~o3;
  assign new_n1263_ = new_n1261_ & new_n1262_;
  assign new_n1264_ = new_n614_ & new_n1263_;
  assign new_n1265_ = new_n614_ & ~new_n1263_;
  assign new_n1266_ = new_n1218_ & ~new_n1265_;
  assign q8 = new_n1264_ | new_n1266_;
  assign new_n1268_ = l3 & m3;
  assign new_n1269_ = n3 & o3;
  assign new_n1270_ = new_n1268_ & new_n1269_;
  assign r8 = new_n614_ & new_n1270_;
  assign new_n1272_ = ~i3 & ~new_n1248_;
  assign new_n1273_ = ~h0 & ~new_n1272_;
  assign new_n1274_ = i3 & ~new_n1250_;
  assign new_n1275_ = ~h0 & ~new_n1274_;
  assign new_n1276_ = ~new_n1218_ & new_n1275_;
  assign new_n1277_ = ~new_n1218_ & ~new_n1275_;
  assign new_n1278_ = new_n1273_ & ~new_n1277_;
  assign new_n1279_ = ~new_n1276_ & ~new_n1278_;
  assign new_n1280_ = ~new_n594_ & new_n1279_;
  assign new_n1281_ = ~l3 & ~new_n1280_;
  assign new_n1282_ = l3 & new_n1280_;
  assign new_n1283_ = ~new_n1281_ & ~new_n1282_;
  assign s8 = new_n614_ & new_n1283_;
  assign new_n1285_ = ~l3 & ~new_n1273_;
  assign new_n1286_ = l3 & ~new_n1275_;
  assign new_n1287_ = ~new_n1218_ & ~new_n1286_;
  assign new_n1288_ = ~new_n1218_ & new_n1286_;
  assign new_n1289_ = ~new_n1285_ & ~new_n1288_;
  assign new_n1290_ = ~new_n1287_ & ~new_n1289_;
  assign new_n1291_ = ~new_n594_ & new_n1290_;
  assign new_n1292_ = ~m3 & ~new_n1291_;
  assign new_n1293_ = m3 & new_n1291_;
  assign new_n1294_ = ~new_n1292_ & ~new_n1293_;
  assign t8 = new_n614_ & new_n1294_;
  assign new_n1296_ = ~m3 & new_n1285_;
  assign new_n1297_ = new_n1268_ & ~new_n1275_;
  assign new_n1298_ = ~new_n1218_ & ~new_n1297_;
  assign new_n1299_ = ~new_n1218_ & new_n1297_;
  assign new_n1300_ = ~new_n1296_ & ~new_n1299_;
  assign new_n1301_ = ~new_n1298_ & ~new_n1300_;
  assign new_n1302_ = ~new_n594_ & new_n1301_;
  assign new_n1303_ = ~n3 & ~new_n1302_;
  assign new_n1304_ = n3 & new_n1302_;
  assign new_n1305_ = ~new_n1303_ & ~new_n1304_;
  assign u8 = new_n614_ & new_n1305_;
  assign new_n1307_ = ~n3 & new_n1296_;
  assign new_n1308_ = m3 & n3;
  assign new_n1309_ = l3 & new_n1308_;
  assign new_n1310_ = ~new_n1275_ & new_n1309_;
  assign new_n1311_ = ~new_n1218_ & ~new_n1310_;
  assign new_n1312_ = ~new_n1218_ & new_n1310_;
  assign new_n1313_ = ~new_n1307_ & ~new_n1312_;
  assign new_n1314_ = ~new_n1311_ & ~new_n1313_;
  assign new_n1315_ = ~new_n594_ & new_n1314_;
  assign new_n1316_ = ~o3 & new_n1315_;
  assign new_n1317_ = o3 & ~new_n1315_;
  assign new_n1318_ = ~new_n1316_ & ~new_n1317_;
  assign new_n1319_ = new_n614_ & ~new_n1318_;
  assign v8 = new_n1259_ | new_n1319_;
  assign new_n1321_ = j3 & ~new_n1273_;
  assign new_n1322_ = k3 & ~new_n1275_;
  assign new_n1323_ = ~new_n1218_ & ~new_n1322_;
  assign new_n1324_ = ~new_n1218_ & new_n1322_;
  assign new_n1325_ = ~new_n1321_ & ~new_n1324_;
  assign new_n1326_ = ~new_n1323_ & ~new_n1325_;
  assign new_n1327_ = ~new_n594_ & new_n1326_;
  assign new_n1328_ = ~p3 & new_n1327_;
  assign new_n1329_ = p3 & ~new_n1327_;
  assign new_n1330_ = ~new_n1328_ & ~new_n1329_;
  assign new_n1331_ = new_n614_ & ~new_n1330_;
  assign w8 = new_n1259_ | new_n1331_;
  assign new_n1333_ = ~p3 & new_n1321_;
  assign new_n1334_ = ~h0 & ~new_n1333_;
  assign new_n1335_ = p3 & new_n1322_;
  assign new_n1336_ = ~h0 & ~new_n1335_;
  assign new_n1337_ = ~new_n1218_ & new_n1336_;
  assign new_n1338_ = ~new_n1218_ & ~new_n1336_;
  assign new_n1339_ = new_n1334_ & ~new_n1338_;
  assign new_n1340_ = ~new_n1337_ & ~new_n1339_;
  assign new_n1341_ = ~new_n594_ & new_n1340_;
  assign new_n1342_ = ~q3 & new_n1341_;
  assign new_n1343_ = q3 & ~new_n1341_;
  assign new_n1344_ = ~new_n1342_ & ~new_n1343_;
  assign new_n1345_ = new_n614_ & ~new_n1344_;
  assign x8 = new_n1259_ | new_n1345_;
  assign new_n1347_ = ~q3 & ~new_n1334_;
  assign new_n1348_ = q3 & ~new_n1336_;
  assign new_n1349_ = ~new_n1218_ & ~new_n1348_;
  assign new_n1350_ = ~new_n1218_ & new_n1348_;
  assign new_n1351_ = ~new_n1347_ & ~new_n1350_;
  assign new_n1352_ = ~new_n1349_ & ~new_n1351_;
  assign new_n1353_ = ~new_n594_ & new_n1352_;
  assign new_n1354_ = ~r3 & ~new_n1353_;
  assign new_n1355_ = r3 & new_n1353_;
  assign new_n1356_ = ~new_n1354_ & ~new_n1355_;
  assign y8 = new_n614_ & new_n1356_;
  assign new_n1358_ = ~r3 & new_n1347_;
  assign new_n1359_ = r3 & new_n1348_;
  assign new_n1360_ = ~new_n1218_ & ~new_n1359_;
  assign new_n1361_ = ~new_n1218_ & new_n1359_;
  assign new_n1362_ = ~new_n1358_ & ~new_n1361_;
  assign new_n1363_ = ~new_n1360_ & ~new_n1362_;
  assign new_n1364_ = ~new_n594_ & new_n1363_;
  assign new_n1365_ = ~s3 & new_n1364_;
  assign new_n1366_ = s3 & ~new_n1364_;
  assign new_n1367_ = ~new_n1365_ & ~new_n1366_;
  assign new_n1368_ = new_n614_ & ~new_n1367_;
  assign z8 = new_n1259_ | new_n1368_;
  assign new_n1370_ = ~s3 & new_n1358_;
  assign new_n1371_ = r3 & s3;
  assign new_n1372_ = new_n1348_ & new_n1371_;
  assign new_n1373_ = ~new_n1218_ & ~new_n1372_;
  assign new_n1374_ = ~new_n1218_ & new_n1372_;
  assign new_n1375_ = ~new_n1370_ & ~new_n1374_;
  assign new_n1376_ = ~new_n1373_ & ~new_n1375_;
  assign new_n1377_ = ~new_n594_ & new_n1376_;
  assign new_n1378_ = ~t3 & new_n1377_;
  assign new_n1379_ = t3 & ~new_n1377_;
  assign new_n1380_ = ~new_n1378_ & ~new_n1379_;
  assign new_n1381_ = new_n614_ & ~new_n1380_;
  assign a9 = new_n1259_ | new_n1381_;
  assign new_n1383_ = ~r4 & s4;
  assign new_n1384_ = r5 & new_n581_;
  assign new_n1385_ = p5 & new_n577_;
  assign new_n1386_ = q5 & new_n578_;
  assign new_n1387_ = ~new_n1385_ & ~new_n1386_;
  assign new_n1388_ = ~new_n1384_ & new_n1387_;
  assign new_n1389_ = new_n1383_ & ~new_n1388_;
  assign new_n1390_ = v10 & new_n1389_;
  assign new_n1391_ = ~f0 & ~new_n1390_;
  assign new_n1392_ = ~u3 & ~new_n1391_;
  assign new_n1393_ = u3 & new_n1391_;
  assign new_n1394_ = ~new_n1392_ & ~new_n1393_;
  assign new_n1395_ = r4 & new_n583_;
  assign new_n1396_ = l5 & ~m5;
  assign new_n1397_ = ~n5 & new_n1396_;
  assign new_n1398_ = ~z & new_n1397_;
  assign new_n1399_ = v10 & new_n1395_;
  assign new_n1400_ = ~new_n1398_ & ~new_n1399_;
  assign new_n1401_ = new_n1394_ & new_n1400_;
  assign new_n1402_ = ~new_n1394_ & new_n1400_;
  assign new_n1403_ = ~l3 & ~new_n1402_;
  assign new_n1404_ = ~new_n1401_ & ~new_n1403_;
  assign b9 = ~z & new_n1404_;
  assign new_n1406_ = ~g0 & new_n576_;
  assign new_n1407_ = ~u3 & ~new_n1406_;
  assign new_n1408_ = u3 & new_n1406_;
  assign new_n1409_ = ~new_n1407_ & ~new_n1408_;
  assign new_n1410_ = ~new_n1391_ & new_n1409_;
  assign new_n1411_ = ~v3 & new_n1410_;
  assign new_n1412_ = v3 & ~new_n1410_;
  assign new_n1413_ = ~new_n1411_ & ~new_n1412_;
  assign new_n1414_ = new_n1400_ & new_n1413_;
  assign new_n1415_ = new_n1400_ & ~new_n1413_;
  assign new_n1416_ = ~m3 & ~new_n1415_;
  assign new_n1417_ = ~new_n1414_ & ~new_n1416_;
  assign c9 = ~z & new_n1417_;
  assign new_n1419_ = ~u3 & ~v3;
  assign new_n1420_ = u3 & v3;
  assign new_n1421_ = ~new_n1406_ & ~new_n1420_;
  assign new_n1422_ = ~new_n1406_ & new_n1420_;
  assign new_n1423_ = ~new_n1419_ & ~new_n1422_;
  assign new_n1424_ = ~new_n1421_ & ~new_n1423_;
  assign new_n1425_ = ~new_n1391_ & new_n1424_;
  assign new_n1426_ = ~w3 & new_n1425_;
  assign new_n1427_ = w3 & ~new_n1425_;
  assign new_n1428_ = ~new_n1426_ & ~new_n1427_;
  assign new_n1429_ = new_n1400_ & new_n1428_;
  assign new_n1430_ = new_n1400_ & ~new_n1428_;
  assign new_n1431_ = ~n3 & ~new_n1430_;
  assign new_n1432_ = ~new_n1429_ & ~new_n1431_;
  assign d9 = ~z & new_n1432_;
  assign new_n1434_ = ~w3 & new_n1419_;
  assign new_n1435_ = ~i0 & ~new_n1434_;
  assign new_n1436_ = w3 & new_n1420_;
  assign new_n1437_ = ~i0 & ~new_n1436_;
  assign new_n1438_ = ~new_n1406_ & new_n1437_;
  assign new_n1439_ = ~new_n1406_ & ~new_n1437_;
  assign new_n1440_ = new_n1435_ & ~new_n1439_;
  assign new_n1441_ = ~new_n1438_ & ~new_n1440_;
  assign new_n1442_ = ~new_n1391_ & new_n1441_;
  assign new_n1443_ = ~x3 & new_n1442_;
  assign new_n1444_ = x3 & ~new_n1442_;
  assign new_n1445_ = ~new_n1443_ & ~new_n1444_;
  assign new_n1446_ = new_n1400_ & new_n1445_;
  assign new_n1447_ = new_n1400_ & ~new_n1445_;
  assign new_n1448_ = ~o3 & ~new_n1447_;
  assign new_n1449_ = ~new_n1446_ & ~new_n1448_;
  assign e9 = z | new_n1449_;
  assign new_n1451_ = ~x3 & ~new_n1435_;
  assign new_n1452_ = x3 & ~new_n1437_;
  assign new_n1453_ = ~new_n1406_ & ~new_n1452_;
  assign new_n1454_ = ~new_n1406_ & new_n1452_;
  assign new_n1455_ = ~new_n1451_ & ~new_n1454_;
  assign new_n1456_ = ~new_n1453_ & ~new_n1455_;
  assign new_n1457_ = ~new_n1391_ & new_n1456_;
  assign new_n1458_ = ~y3 & new_n1457_;
  assign new_n1459_ = y3 & ~new_n1457_;
  assign new_n1460_ = ~new_n1458_ & ~new_n1459_;
  assign new_n1461_ = new_n1400_ & new_n1460_;
  assign new_n1462_ = new_n1400_ & ~new_n1460_;
  assign new_n1463_ = ~p3 & ~new_n1462_;
  assign new_n1464_ = ~new_n1461_ & ~new_n1463_;
  assign f9 = z | new_n1464_;
  assign new_n1466_ = ~y3 & new_n1451_;
  assign new_n1467_ = x3 & y3;
  assign new_n1468_ = ~new_n1437_ & new_n1467_;
  assign new_n1469_ = ~new_n1406_ & ~new_n1468_;
  assign new_n1470_ = ~new_n1406_ & new_n1468_;
  assign new_n1471_ = ~new_n1466_ & ~new_n1470_;
  assign new_n1472_ = ~new_n1469_ & ~new_n1471_;
  assign new_n1473_ = ~new_n1391_ & new_n1472_;
  assign new_n1474_ = ~z3 & new_n1473_;
  assign new_n1475_ = z3 & ~new_n1473_;
  assign new_n1476_ = ~new_n1474_ & ~new_n1475_;
  assign new_n1477_ = new_n1400_ & new_n1476_;
  assign new_n1478_ = new_n1400_ & ~new_n1476_;
  assign new_n1479_ = ~q3 & ~new_n1478_;
  assign new_n1480_ = ~new_n1477_ & ~new_n1479_;
  assign g9 = z | new_n1480_;
  assign new_n1482_ = ~y3 & ~z3;
  assign new_n1483_ = new_n1451_ & new_n1482_;
  assign new_n1484_ = ~i0 & ~new_n1483_;
  assign new_n1485_ = y3 & z3;
  assign new_n1486_ = new_n1452_ & new_n1485_;
  assign new_n1487_ = ~i0 & ~new_n1486_;
  assign new_n1488_ = ~new_n1406_ & new_n1487_;
  assign new_n1489_ = ~new_n1406_ & ~new_n1487_;
  assign new_n1490_ = new_n1484_ & ~new_n1489_;
  assign new_n1491_ = ~new_n1488_ & ~new_n1490_;
  assign new_n1492_ = ~new_n1391_ & new_n1491_;
  assign new_n1493_ = ~a4 & new_n1492_;
  assign new_n1494_ = a4 & ~new_n1492_;
  assign new_n1495_ = ~new_n1493_ & ~new_n1494_;
  assign new_n1496_ = new_n1400_ & new_n1495_;
  assign new_n1497_ = new_n1400_ & ~new_n1495_;
  assign new_n1498_ = ~r3 & ~new_n1497_;
  assign new_n1499_ = ~new_n1496_ & ~new_n1498_;
  assign h9 = ~z & new_n1499_;
  assign new_n1501_ = ~a4 & ~new_n1484_;
  assign new_n1502_ = a4 & ~new_n1487_;
  assign new_n1503_ = ~new_n1406_ & ~new_n1502_;
  assign new_n1504_ = ~new_n1406_ & new_n1502_;
  assign new_n1505_ = ~new_n1501_ & ~new_n1504_;
  assign new_n1506_ = ~new_n1503_ & ~new_n1505_;
  assign new_n1507_ = ~new_n1391_ & new_n1506_;
  assign new_n1508_ = ~b4 & new_n1507_;
  assign new_n1509_ = b4 & ~new_n1507_;
  assign new_n1510_ = ~new_n1508_ & ~new_n1509_;
  assign new_n1511_ = new_n1400_ & new_n1510_;
  assign new_n1512_ = new_n1400_ & ~new_n1510_;
  assign new_n1513_ = ~s3 & ~new_n1512_;
  assign new_n1514_ = ~new_n1511_ & ~new_n1513_;
  assign i9 = z | new_n1514_;
  assign new_n1516_ = ~b4 & new_n1501_;
  assign new_n1517_ = a4 & b4;
  assign new_n1518_ = ~new_n1487_ & new_n1517_;
  assign new_n1519_ = ~new_n1406_ & ~new_n1518_;
  assign new_n1520_ = ~new_n1406_ & new_n1518_;
  assign new_n1521_ = ~new_n1516_ & ~new_n1520_;
  assign new_n1522_ = ~new_n1519_ & ~new_n1521_;
  assign new_n1523_ = ~new_n1391_ & new_n1522_;
  assign new_n1524_ = ~c4 & new_n1523_;
  assign new_n1525_ = c4 & ~new_n1523_;
  assign new_n1526_ = ~new_n1524_ & ~new_n1525_;
  assign new_n1527_ = new_n1400_ & new_n1526_;
  assign new_n1528_ = new_n1400_ & ~new_n1526_;
  assign new_n1529_ = ~t3 & ~new_n1528_;
  assign new_n1530_ = ~new_n1527_ & ~new_n1529_;
  assign j9 = z | new_n1530_;
  assign k9 = z | ~d4;
  assign new_n1533_ = ~d4 & ~e4;
  assign new_n1534_ = ~new_n601_ & ~new_n1533_;
  assign l9 = z | new_n1534_;
  assign new_n1536_ = ~f4 & ~new_n601_;
  assign new_n1537_ = ~new_n602_ & ~new_n1536_;
  assign m9 = z | new_n1537_;
  assign new_n1539_ = ~g4 & ~new_n606_;
  assign new_n1540_ = g4 & new_n606_;
  assign new_n1541_ = ~new_n1539_ & ~new_n1540_;
  assign new_n1542_ = ~m5 & n5;
  assign new_n1543_ = ~z & l5;
  assign new_n1544_ = new_n1542_ & new_n1543_;
  assign new_n1545_ = ~new_n608_ & ~new_n1544_;
  assign new_n1546_ = new_n1541_ & new_n1545_;
  assign new_n1547_ = ~new_n1541_ & new_n1545_;
  assign new_n1548_ = ~u3 & ~new_n1547_;
  assign new_n1549_ = ~new_n1546_ & ~new_n1548_;
  assign n9 = z | new_n1549_;
  assign new_n1551_ = ~h4 & new_n607_;
  assign new_n1552_ = h4 & ~new_n607_;
  assign new_n1553_ = ~new_n1551_ & ~new_n1552_;
  assign new_n1554_ = new_n1545_ & new_n1553_;
  assign new_n1555_ = new_n1545_ & ~new_n1553_;
  assign new_n1556_ = ~v3 & ~new_n1555_;
  assign new_n1557_ = ~new_n1554_ & ~new_n1556_;
  assign o9 = z | new_n1557_;
  assign new_n1559_ = ~i4 & new_n603_;
  assign new_n1560_ = ~new_n604_ & ~new_n1559_;
  assign p9 = z | new_n1560_;
  assign new_n1562_ = h4 & new_n607_;
  assign new_n1563_ = ~j4 & new_n1562_;
  assign new_n1564_ = j4 & ~new_n1562_;
  assign new_n1565_ = ~new_n1563_ & ~new_n1564_;
  assign new_n1566_ = new_n1545_ & new_n1565_;
  assign new_n1567_ = new_n1545_ & ~new_n1565_;
  assign new_n1568_ = ~w3 & ~new_n1567_;
  assign new_n1569_ = ~new_n1566_ & ~new_n1568_;
  assign q9 = z | new_n1569_;
  assign new_n1571_ = h4 & j4;
  assign new_n1572_ = new_n607_ & new_n1571_;
  assign new_n1573_ = ~k4 & new_n1572_;
  assign new_n1574_ = k4 & ~new_n1572_;
  assign new_n1575_ = ~new_n1573_ & ~new_n1574_;
  assign new_n1576_ = new_n1545_ & new_n1575_;
  assign new_n1577_ = new_n1545_ & ~new_n1575_;
  assign new_n1578_ = ~x3 & ~new_n1577_;
  assign new_n1579_ = ~new_n1576_ & ~new_n1578_;
  assign r9 = z | new_n1579_;
  assign new_n1581_ = k4 & new_n1572_;
  assign new_n1582_ = ~l4 & new_n1581_;
  assign new_n1583_ = l4 & ~new_n1581_;
  assign new_n1584_ = ~new_n1582_ & ~new_n1583_;
  assign new_n1585_ = new_n1545_ & new_n1584_;
  assign new_n1586_ = new_n1545_ & ~new_n1584_;
  assign new_n1587_ = ~y3 & ~new_n1586_;
  assign new_n1588_ = ~new_n1585_ & ~new_n1587_;
  assign s9 = z | new_n1588_;
  assign new_n1590_ = l4 & new_n1581_;
  assign new_n1591_ = ~j0 & ~new_n1590_;
  assign new_n1592_ = ~m4 & ~new_n1591_;
  assign new_n1593_ = m4 & new_n1591_;
  assign new_n1594_ = ~new_n1592_ & ~new_n1593_;
  assign new_n1595_ = new_n1545_ & new_n1594_;
  assign new_n1596_ = new_n1545_ & ~new_n1594_;
  assign new_n1597_ = ~z3 & ~new_n1596_;
  assign new_n1598_ = ~new_n1595_ & ~new_n1597_;
  assign t9 = z | new_n1598_;
  assign new_n1600_ = m4 & ~new_n1591_;
  assign new_n1601_ = ~n4 & new_n1600_;
  assign new_n1602_ = n4 & ~new_n1600_;
  assign new_n1603_ = ~new_n1601_ & ~new_n1602_;
  assign new_n1604_ = new_n1545_ & new_n1603_;
  assign new_n1605_ = new_n1545_ & ~new_n1603_;
  assign new_n1606_ = ~a4 & ~new_n1605_;
  assign new_n1607_ = ~new_n1604_ & ~new_n1606_;
  assign u9 = z | new_n1607_;
  assign new_n1609_ = m4 & n4;
  assign new_n1610_ = ~new_n1591_ & new_n1609_;
  assign new_n1611_ = ~o4 & new_n1610_;
  assign new_n1612_ = o4 & ~new_n1610_;
  assign new_n1613_ = ~new_n1611_ & ~new_n1612_;
  assign new_n1614_ = new_n1545_ & new_n1613_;
  assign new_n1615_ = new_n1545_ & ~new_n1613_;
  assign new_n1616_ = ~b4 & ~new_n1615_;
  assign new_n1617_ = ~new_n1614_ & ~new_n1616_;
  assign v9 = z | new_n1617_;
  assign new_n1619_ = o4 & q4;
  assign new_n1620_ = n4 & new_n1619_;
  assign new_n1621_ = l4 & m4;
  assign new_n1622_ = k4 & new_n1621_;
  assign new_n1623_ = ~z & ~new_n1545_;
  assign new_n1624_ = new_n1620_ & new_n1622_;
  assign new_n1625_ = new_n1571_ & new_n1624_;
  assign w9 = ~new_n1623_ & new_n1625_;
  assign new_n1627_ = o4 & new_n1610_;
  assign new_n1628_ = ~q4 & new_n1627_;
  assign new_n1629_ = q4 & ~new_n1627_;
  assign new_n1630_ = ~new_n1628_ & ~new_n1629_;
  assign new_n1631_ = new_n1545_ & new_n1630_;
  assign new_n1632_ = new_n1545_ & ~new_n1630_;
  assign new_n1633_ = ~c4 & ~new_n1632_;
  assign new_n1634_ = ~new_n1631_ & ~new_n1633_;
  assign x9 = z | new_n1634_;
  assign new_n1636_ = r5 & new_n1229_;
  assign new_n1637_ = new_n576_ & ~new_n1636_;
  assign new_n1638_ = new_n572_ & new_n1637_;
  assign new_n1639_ = ~r4 & new_n1638_;
  assign new_n1640_ = r4 & ~new_n1638_;
  assign new_n1641_ = ~new_n1639_ & ~new_n1640_;
  assign new_n1642_ = new_n585_ & v10;
  assign new_n1643_ = r4 & new_n1636_;
  assign new_n1644_ = ~new_n1642_ & ~new_n1643_;
  assign new_n1645_ = ~z & ~new_n1544_;
  assign new_n1646_ = new_n1644_ & new_n1645_;
  assign y9 = new_n1641_ & new_n1646_;
  assign new_n1648_ = ~s4 & ~new_n1640_;
  assign new_n1649_ = s4 & new_n1640_;
  assign new_n1650_ = ~new_n1648_ & ~new_n1649_;
  assign z9 = new_n1646_ & new_n1650_;
  assign new_n1652_ = r4 & s4;
  assign new_n1653_ = ~new_n1638_ & new_n1652_;
  assign new_n1654_ = ~t4 & ~new_n1653_;
  assign new_n1655_ = t4 & new_n1653_;
  assign new_n1656_ = ~new_n1654_ & ~new_n1655_;
  assign a10 = new_n1646_ & new_n1656_;
  assign new_n1658_ = t4 & new_n1652_;
  assign new_n1659_ = ~new_n1638_ & new_n1658_;
  assign new_n1660_ = ~u4 & ~new_n1659_;
  assign new_n1661_ = u4 & new_n1659_;
  assign new_n1662_ = ~new_n1660_ & ~new_n1661_;
  assign b10 = new_n1646_ & new_n1662_;
  assign new_n1664_ = t4 & u4;
  assign new_n1665_ = new_n1652_ & new_n1664_;
  assign new_n1666_ = ~new_n1638_ & new_n1665_;
  assign new_n1667_ = ~v4 & ~new_n1666_;
  assign new_n1668_ = v4 & new_n1666_;
  assign new_n1669_ = ~new_n1667_ & ~new_n1668_;
  assign c10 = new_n1646_ & new_n1669_;
  assign new_n1671_ = v4 & new_n1665_;
  assign new_n1672_ = ~new_n1638_ & new_n1671_;
  assign new_n1673_ = ~w4 & ~new_n1672_;
  assign new_n1674_ = w4 & new_n1672_;
  assign new_n1675_ = ~new_n1673_ & ~new_n1674_;
  assign d10 = new_n1646_ & new_n1675_;
  assign new_n1677_ = w4 & new_n1671_;
  assign new_n1678_ = ~new_n1638_ & new_n1677_;
  assign new_n1679_ = ~x4 & ~new_n1678_;
  assign new_n1680_ = x4 & new_n1678_;
  assign new_n1681_ = ~new_n1679_ & ~new_n1680_;
  assign e10 = new_n1646_ & new_n1681_;
  assign new_n1683_ = v4 & w4;
  assign new_n1684_ = x4 & new_n1683_;
  assign new_n1685_ = new_n1665_ & new_n1684_;
  assign new_n1686_ = ~new_n1638_ & new_n1685_;
  assign new_n1687_ = ~y4 & ~new_n1686_;
  assign new_n1688_ = y4 & new_n1686_;
  assign new_n1689_ = ~new_n1687_ & ~new_n1688_;
  assign f10 = new_n1646_ & new_n1689_;
  assign new_n1691_ = y4 & ~new_n1638_;
  assign new_n1692_ = new_n1685_ & new_n1691_;
  assign new_n1693_ = z4 & new_n1692_;
  assign new_n1694_ = ~z4 & ~new_n1692_;
  assign new_n1695_ = ~new_n1693_ & ~new_n1694_;
  assign g10 = new_n1646_ & new_n1695_;
  assign new_n1697_ = d5 & new_n562_;
  assign new_n1698_ = new_n1645_ & ~new_n1697_;
  assign new_n1699_ = d5 & new_n1698_;
  assign k10 = new_n571_ | new_n1699_;
  assign new_n1701_ = e5 & new_n566_;
  assign new_n1702_ = new_n1645_ & ~new_n1701_;
  assign new_n1703_ = e5 & new_n1702_;
  assign l10 = new_n574_ | new_n1703_;
  assign new_n1705_ = h5 & new_n608_;
  assign new_n1706_ = ~h5 & ~new_n608_;
  assign new_n1707_ = ~new_n1705_ & ~new_n1706_;
  assign new_n1708_ = ~z & new_n1707_;
  assign new_n1709_ = ~new_n1398_ & ~new_n1544_;
  assign o10 = new_n1708_ | ~new_n1709_;
  assign new_n1711_ = ~h5 & o10;
  assign new_n1712_ = ~f5 & ~g5;
  assign new_n1713_ = new_n1711_ & ~new_n1712_;
  assign new_n1714_ = new_n1711_ & new_n1712_;
  assign new_n1715_ = ~f5 & ~new_n1714_;
  assign new_n1716_ = ~new_n1713_ & ~new_n1715_;
  assign new_n1717_ = ~z & ~new_n1716_;
  assign m10 = new_n1709_ & ~new_n1717_;
  assign new_n1719_ = ~g5 & ~new_n1711_;
  assign new_n1720_ = g5 & ~new_n1711_;
  assign new_n1721_ = ~f5 & ~new_n1720_;
  assign new_n1722_ = ~new_n1719_ & ~new_n1721_;
  assign new_n1723_ = new_n1709_ & ~new_n1722_;
  assign n10 = ~z & ~new_n1723_;
  assign new_n1725_ = j5 & new_n1229_;
  assign new_n1726_ = ~j5 & ~new_n1229_;
  assign new_n1727_ = ~new_n1725_ & ~new_n1726_;
  assign new_n1728_ = ~z & ~new_n560_;
  assign q10 = new_n1727_ & new_n1728_;
  assign new_n1730_ = ~k5 & ~new_n1725_;
  assign new_n1731_ = k5 & new_n1725_;
  assign new_n1732_ = ~new_n1730_ & ~new_n1731_;
  assign r10 = new_n1728_ & new_n1732_;
  assign new_n1734_ = new_n562_ & ~new_n631_;
  assign new_n1735_ = new_n623_ & new_n1734_;
  assign new_n1736_ = new_n1229_ & ~new_n1735_;
  assign new_n1737_ = new_n562_ & new_n613_;
  assign new_n1738_ = ~new_n1398_ & ~new_n1736_;
  assign new_n1739_ = ~new_n1737_ & new_n1738_;
  assign s10 = ~z & ~new_n1739_;
  assign new_n1741_ = r5 & ~new_n1693_;
  assign new_n1742_ = r5 & new_n1693_;
  assign new_n1743_ = ~z4 & ~new_n1742_;
  assign new_n1744_ = ~new_n1741_ & ~new_n1743_;
  assign new_n1745_ = ~a0 & ~new_n1744_;
  assign new_n1746_ = v10 & ~new_n1745_;
  assign new_n1747_ = new_n631_ & new_n1229_;
  assign new_n1748_ = ~new_n1746_ & ~new_n1747_;
  assign new_n1749_ = n5 & new_n587_;
  assign new_n1750_ = ~z & new_n1749_;
  assign new_n1751_ = ~new_n613_ & new_n1748_;
  assign new_n1752_ = ~new_n1750_ & new_n1751_;
  assign new_n1753_ = n5 & new_n1227_;
  assign new_n1754_ = ~z & new_n1753_;
  assign new_n1755_ = m5 & n5;
  assign new_n1756_ = ~new_n562_ & ~new_n631_;
  assign new_n1757_ = new_n1229_ & new_n1756_;
  assign new_n1758_ = ~new_n1755_ & ~new_n1757_;
  assign new_n1759_ = ~new_n1754_ & new_n1758_;
  assign new_n1760_ = new_n1752_ & new_n1759_;
  assign t10 = ~z & ~new_n1760_;
  assign new_n1762_ = ~new_n1747_ & ~new_n1750_;
  assign new_n1763_ = ~new_n1398_ & new_n1762_;
  assign new_n1764_ = new_n562_ & new_n1229_;
  assign new_n1765_ = new_n623_ & ~new_n631_;
  assign new_n1766_ = new_n1764_ & new_n1765_;
  assign new_n1767_ = ~new_n1754_ & ~new_n1766_;
  assign new_n1768_ = new_n1763_ & new_n1767_;
  assign u10 = ~z & ~new_n1768_;
  assign new_n1770_ = q5 & r5;
  assign new_n1771_ = ~p5 & ~new_n1770_;
  assign new_n1772_ = ~q5 & ~r5;
  assign new_n1773_ = ~new_n1771_ & ~new_n1772_;
  assign new_n1774_ = ~p5 & new_n1772_;
  assign new_n1775_ = ~z & ~new_n1774_;
  assign new_n1776_ = ~new_n1773_ & new_n1775_;
  assign new_n1777_ = ~c0 & ~new_n1754_;
  assign new_n1778_ = ~b0 & ~new_n1750_;
  assign new_n1779_ = q5 & ~new_n1778_;
  assign new_n1780_ = r5 & ~new_n1777_;
  assign new_n1781_ = ~p5 & ~new_n1780_;
  assign new_n1782_ = ~r5 & ~new_n1777_;
  assign new_n1783_ = ~new_n1781_ & ~new_n1782_;
  assign new_n1784_ = ~new_n1779_ & ~new_n1783_;
  assign new_n1785_ = ~new_n1778_ & ~new_n1780_;
  assign new_n1786_ = ~q5 & new_n1785_;
  assign new_n1787_ = ~new_n1784_ & ~new_n1786_;
  assign w10 = ~new_n1776_ | new_n1787_;
  assign new_n1789_ = r5 & ~new_n1778_;
  assign new_n1790_ = q5 & new_n1777_;
  assign new_n1791_ = ~p5 & ~new_n1790_;
  assign new_n1792_ = ~q5 & new_n1777_;
  assign new_n1793_ = ~new_n1791_ & ~new_n1792_;
  assign new_n1794_ = ~new_n1789_ & ~new_n1793_;
  assign new_n1795_ = p5 & ~new_n1777_;
  assign new_n1796_ = ~new_n1778_ & ~new_n1795_;
  assign new_n1797_ = ~r5 & new_n1796_;
  assign new_n1798_ = ~new_n1794_ & ~new_n1797_;
  assign x10 = new_n1776_ & new_n1798_;
  assign new_n1800_ = p5 & ~new_n1778_;
  assign new_n1801_ = ~r5 & new_n1777_;
  assign new_n1802_ = r5 & new_n1777_;
  assign new_n1803_ = ~q5 & ~new_n1802_;
  assign new_n1804_ = ~new_n1801_ & ~new_n1803_;
  assign new_n1805_ = ~new_n1800_ & ~new_n1804_;
  assign new_n1806_ = q5 & ~new_n1777_;
  assign new_n1807_ = ~new_n1778_ & ~new_n1806_;
  assign new_n1808_ = ~p5 & new_n1807_;
  assign new_n1809_ = ~new_n1805_ & ~new_n1808_;
  assign y10 = new_n1776_ & new_n1809_;
  assign l6 = a;
  assign m6 = e1;
  assign r6 = j1;
  assign h10 = y;
  assign i10 = a5;
  assign p10 = g5;
endmodule

