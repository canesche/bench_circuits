// Benchmark "testing" written by ABC on Thu Oct  8 22:16:31 2020

module testing ( 
    A302, A301, A300, A299, A298, A269, A268, A267, A266, A265, A236, A235,
    A234, A233, A232, A203, A202, A201, A200, A199, A166, A167, A168, A169,
    A170,
    A72  );
  input  A302, A301, A300, A299, A298, A269, A268, A267, A266, A265,
    A236, A235, A234, A233, A232, A203, A202, A201, A200, A199, A166, A167,
    A168, A169, A170;
  output A72;
  wire \new_[1]_ , \new_[2]_ , \new_[3]_ , \new_[4]_ , \new_[5]_ ,
    \new_[6]_ , \new_[7]_ , \new_[8]_ , \new_[9]_ , \new_[10]_ ,
    \new_[11]_ , \new_[12]_ , \new_[13]_ , \new_[14]_ , \new_[15]_ ,
    \new_[16]_ , \new_[17]_ , \new_[18]_ , \new_[19]_ , \new_[20]_ ,
    \new_[21]_ , \new_[22]_ , \new_[23]_ , \new_[24]_ , \new_[25]_ ,
    \new_[26]_ , \new_[27]_ , \new_[28]_ , \new_[29]_ , \new_[30]_ ,
    \new_[31]_ , \new_[32]_ , \new_[33]_ , \new_[34]_ , \new_[35]_ ,
    \new_[36]_ , \new_[37]_ , \new_[38]_ , \new_[39]_ , \new_[40]_ ,
    \new_[41]_ , \new_[42]_ , \new_[43]_ , \new_[44]_ , \new_[45]_ ,
    \new_[46]_ , \new_[47]_ , \new_[48]_ , \new_[49]_ , \new_[50]_ ,
    \new_[51]_ , \new_[52]_ , \new_[53]_ , \new_[54]_ , \new_[55]_ ,
    \new_[56]_ , \new_[57]_ , \new_[58]_ , \new_[59]_ , \new_[60]_ ,
    \new_[61]_ , \new_[62]_ , \new_[63]_ , \new_[64]_ , \new_[65]_ ,
    \new_[66]_ , \new_[67]_ , \new_[68]_ , \new_[69]_ , \new_[70]_ ,
    \new_[71]_ , \new_[72]_ , \new_[73]_ , \new_[74]_ , \new_[75]_ ,
    \new_[76]_ , \new_[77]_ , \new_[78]_ , \new_[79]_ , \new_[80]_ ,
    \new_[81]_ , \new_[82]_ , \new_[83]_ , \new_[84]_ , \new_[85]_ ,
    \new_[86]_ , \new_[87]_ , \new_[88]_ , \new_[89]_ , \new_[90]_ ,
    \new_[91]_ , \new_[92]_ , \new_[93]_ , \new_[94]_ , \new_[95]_ ,
    \new_[96]_ , \new_[97]_ , \new_[98]_ , \new_[99]_ , \new_[100]_ ,
    \new_[101]_ , \new_[102]_ , \new_[103]_ , \new_[104]_ , \new_[105]_ ,
    \new_[106]_ , \new_[107]_ , \new_[108]_ , \new_[109]_ , \new_[110]_ ,
    \new_[111]_ , \new_[112]_ , \new_[113]_ , \new_[114]_ , \new_[115]_ ,
    \new_[116]_ , \new_[117]_ , \new_[118]_ , \new_[119]_ , \new_[120]_ ,
    \new_[121]_ , \new_[122]_ , \new_[123]_ , \new_[124]_ , \new_[125]_ ,
    \new_[126]_ , \new_[127]_ , \new_[128]_ , \new_[129]_ , \new_[130]_ ,
    \new_[131]_ , \new_[132]_ , \new_[133]_ , \new_[134]_ , \new_[135]_ ,
    \new_[136]_ , \new_[137]_ , \new_[138]_ , \new_[139]_ , \new_[140]_ ,
    \new_[141]_ , \new_[142]_ , \new_[143]_ , \new_[144]_ , \new_[145]_ ,
    \new_[146]_ , \new_[147]_ , \new_[148]_ , \new_[149]_ , \new_[150]_ ,
    \new_[151]_ , \new_[152]_ , \new_[153]_ , \new_[154]_ , \new_[155]_ ,
    \new_[156]_ , \new_[157]_ , \new_[158]_ , \new_[159]_ , \new_[160]_ ,
    \new_[161]_ , \new_[162]_ , \new_[163]_ , \new_[164]_ , \new_[165]_ ,
    \new_[166]_ , \new_[167]_ , \new_[168]_ , \new_[169]_ , \new_[170]_ ,
    \new_[171]_ , \new_[172]_ , \new_[173]_ , \new_[174]_ , \new_[175]_ ,
    \new_[176]_ , \new_[177]_ , \new_[178]_ , \new_[179]_ , \new_[180]_ ,
    \new_[181]_ , \new_[182]_ , \new_[183]_ , \new_[184]_ , \new_[185]_ ,
    \new_[186]_ , \new_[187]_ , \new_[188]_ , \new_[189]_ , \new_[190]_ ,
    \new_[191]_ , \new_[192]_ , \new_[193]_ , \new_[194]_ , \new_[195]_ ,
    \new_[196]_ , \new_[197]_ , \new_[198]_ , \new_[199]_ , \new_[200]_ ,
    \new_[201]_ , \new_[202]_ , \new_[203]_ , \new_[204]_ , \new_[205]_ ,
    \new_[206]_ , \new_[207]_ , \new_[208]_ , \new_[209]_ , \new_[210]_ ,
    \new_[211]_ , \new_[212]_ , \new_[213]_ , \new_[214]_ , \new_[215]_ ,
    \new_[216]_ , \new_[217]_ , \new_[218]_ , \new_[219]_ , \new_[220]_ ,
    \new_[221]_ , \new_[222]_ , \new_[223]_ , \new_[224]_ , \new_[225]_ ,
    \new_[226]_ , \new_[227]_ , \new_[228]_ , \new_[229]_ , \new_[230]_ ,
    \new_[231]_ , \new_[232]_ , \new_[233]_ , \new_[234]_ , \new_[235]_ ,
    \new_[236]_ , \new_[237]_ , \new_[238]_ , \new_[239]_ , \new_[240]_ ,
    \new_[241]_ , \new_[242]_ , \new_[243]_ , \new_[244]_ , \new_[245]_ ,
    \new_[246]_ , \new_[247]_ , \new_[248]_ , \new_[249]_ , \new_[250]_ ,
    \new_[251]_ , \new_[252]_ , \new_[253]_ , \new_[254]_ , \new_[255]_ ,
    \new_[256]_ , \new_[257]_ , \new_[258]_ , \new_[259]_ , \new_[260]_ ,
    \new_[261]_ , \new_[262]_ , \new_[263]_ , \new_[264]_ , \new_[265]_ ,
    \new_[266]_ , \new_[267]_ , \new_[268]_ , \new_[269]_ , \new_[270]_ ,
    \new_[271]_ , \new_[272]_ , \new_[273]_ , \new_[274]_ , \new_[275]_ ,
    \new_[276]_ , \new_[277]_ , \new_[278]_ , \new_[279]_ , \new_[280]_ ,
    \new_[281]_ , \new_[282]_ , \new_[283]_ , \new_[284]_ , \new_[285]_ ,
    \new_[286]_ , \new_[287]_ , \new_[288]_ , \new_[289]_ , \new_[290]_ ,
    \new_[291]_ , \new_[292]_ , \new_[293]_ , \new_[294]_ , \new_[295]_ ,
    \new_[296]_ , \new_[297]_ , \new_[298]_ , \new_[299]_ , \new_[300]_ ,
    \new_[301]_ , \new_[302]_ , \new_[303]_ , \new_[304]_ , \new_[305]_ ,
    \new_[306]_ , \new_[307]_ , \new_[308]_ , \new_[309]_ , \new_[310]_ ,
    \new_[311]_ , \new_[312]_ , \new_[313]_ , \new_[314]_ , \new_[315]_ ,
    \new_[316]_ , \new_[317]_ , \new_[318]_ , \new_[319]_ , \new_[320]_ ,
    \new_[321]_ , \new_[322]_ , \new_[323]_ , \new_[324]_ , \new_[325]_ ,
    \new_[326]_ , \new_[327]_ , \new_[328]_ , \new_[329]_ , \new_[330]_ ,
    \new_[331]_ , \new_[332]_ , \new_[333]_ , \new_[334]_ , \new_[335]_ ,
    \new_[336]_ , \new_[337]_ , \new_[338]_ , \new_[339]_ , \new_[340]_ ,
    \new_[341]_ , \new_[342]_ , \new_[343]_ , \new_[344]_ , \new_[345]_ ,
    \new_[346]_ , \new_[347]_ , \new_[348]_ , \new_[349]_ , \new_[350]_ ,
    \new_[351]_ , \new_[352]_ , \new_[353]_ , \new_[354]_ , \new_[355]_ ,
    \new_[356]_ , \new_[357]_ , \new_[358]_ , \new_[359]_ , \new_[360]_ ,
    \new_[361]_ , \new_[362]_ , \new_[363]_ , \new_[364]_ , \new_[365]_ ,
    \new_[366]_ , \new_[367]_ , \new_[368]_ , \new_[369]_ , \new_[370]_ ,
    \new_[371]_ , \new_[372]_ , \new_[373]_ , \new_[374]_ , \new_[375]_ ,
    \new_[376]_ , \new_[377]_ , \new_[378]_ , \new_[379]_ , \new_[380]_ ,
    \new_[381]_ , \new_[382]_ , \new_[383]_ , \new_[384]_ , \new_[385]_ ,
    \new_[386]_ , \new_[387]_ , \new_[388]_ , \new_[389]_ , \new_[390]_ ,
    \new_[391]_ , \new_[392]_ , \new_[393]_ , \new_[394]_ , \new_[395]_ ,
    \new_[396]_ , \new_[397]_ , \new_[398]_ , \new_[399]_ , \new_[400]_ ,
    \new_[401]_ , \new_[402]_ , \new_[403]_ , \new_[404]_ , \new_[405]_ ,
    \new_[406]_ , \new_[407]_ , \new_[408]_ , \new_[409]_ , \new_[410]_ ,
    \new_[411]_ , \new_[412]_ , \new_[413]_ , \new_[414]_ , \new_[415]_ ,
    \new_[416]_ , \new_[417]_ , \new_[418]_ , \new_[419]_ , \new_[420]_ ,
    \new_[421]_ , \new_[422]_ , \new_[423]_ , \new_[424]_ , \new_[425]_ ,
    \new_[426]_ , \new_[427]_ , \new_[428]_ , \new_[429]_ , \new_[430]_ ,
    \new_[431]_ , \new_[432]_ , \new_[433]_ , \new_[434]_ , \new_[435]_ ,
    \new_[436]_ , \new_[437]_ , \new_[438]_ , \new_[439]_ , \new_[440]_ ,
    \new_[441]_ , \new_[442]_ , \new_[443]_ , \new_[444]_ , \new_[445]_ ,
    \new_[446]_ , \new_[447]_ , \new_[448]_ , \new_[449]_ , \new_[450]_ ,
    \new_[451]_ , \new_[452]_ , \new_[453]_ , \new_[454]_ , \new_[455]_ ,
    \new_[456]_ , \new_[457]_ , \new_[458]_ , \new_[459]_ , \new_[460]_ ,
    \new_[461]_ , \new_[462]_ , \new_[463]_ , \new_[464]_ , \new_[465]_ ,
    \new_[466]_ , \new_[467]_ , \new_[468]_ , \new_[469]_ , \new_[470]_ ,
    \new_[471]_ , \new_[472]_ , \new_[473]_ , \new_[474]_ , \new_[475]_ ,
    \new_[476]_ , \new_[477]_ , \new_[478]_ , \new_[479]_ , \new_[480]_ ,
    \new_[481]_ , \new_[482]_ , \new_[483]_ , \new_[484]_ , \new_[485]_ ,
    \new_[486]_ , \new_[487]_ , \new_[488]_ , \new_[489]_ , \new_[490]_ ,
    \new_[491]_ , \new_[492]_ , \new_[493]_ , \new_[494]_ , \new_[495]_ ,
    \new_[496]_ , \new_[497]_ , \new_[498]_ , \new_[499]_ , \new_[500]_ ,
    \new_[501]_ , \new_[502]_ , \new_[503]_ , \new_[504]_ , \new_[505]_ ,
    \new_[506]_ , \new_[507]_ , \new_[508]_ , \new_[509]_ , \new_[510]_ ,
    \new_[511]_ , \new_[512]_ , \new_[513]_ , \new_[514]_ , \new_[515]_ ,
    \new_[516]_ , \new_[517]_ , \new_[518]_ , \new_[519]_ , \new_[520]_ ,
    \new_[521]_ , \new_[522]_ , \new_[523]_ , \new_[524]_ , \new_[525]_ ,
    \new_[526]_ , \new_[527]_ , \new_[528]_ , \new_[529]_ , \new_[530]_ ,
    \new_[531]_ , \new_[532]_ , \new_[533]_ , \new_[534]_ , \new_[535]_ ,
    \new_[536]_ , \new_[537]_ , \new_[538]_ , \new_[539]_ , \new_[540]_ ,
    \new_[541]_ , \new_[542]_ , \new_[543]_ , \new_[544]_ , \new_[545]_ ,
    \new_[546]_ , \new_[547]_ , \new_[548]_ , \new_[549]_ , \new_[550]_ ,
    \new_[551]_ , \new_[552]_ , \new_[553]_ , \new_[554]_ , \new_[555]_ ,
    \new_[556]_ , \new_[557]_ , \new_[558]_ , \new_[559]_ , \new_[560]_ ,
    \new_[561]_ , \new_[562]_ , \new_[563]_ , \new_[564]_ , \new_[565]_ ,
    \new_[566]_ , \new_[567]_ , \new_[568]_ , \new_[569]_ , \new_[570]_ ,
    \new_[571]_ , \new_[572]_ , \new_[573]_ , \new_[574]_ , \new_[575]_ ,
    \new_[576]_ , \new_[577]_ , \new_[578]_ , \new_[579]_ , \new_[580]_ ,
    \new_[581]_ , \new_[582]_ , \new_[583]_ , \new_[584]_ , \new_[585]_ ,
    \new_[586]_ , \new_[587]_ , \new_[588]_ , \new_[589]_ , \new_[590]_ ,
    \new_[591]_ , \new_[592]_ , \new_[593]_ , \new_[594]_ , \new_[595]_ ,
    \new_[596]_ , \new_[597]_ , \new_[598]_ , \new_[599]_ , \new_[600]_ ,
    \new_[601]_ , \new_[602]_ , \new_[603]_ , \new_[604]_ , \new_[605]_ ,
    \new_[606]_ , \new_[607]_ , \new_[608]_ , \new_[609]_ , \new_[610]_ ,
    \new_[611]_ , \new_[612]_ , \new_[613]_ , \new_[614]_ , \new_[615]_ ,
    \new_[616]_ , \new_[617]_ , \new_[618]_ , \new_[619]_ , \new_[620]_ ,
    \new_[621]_ , \new_[622]_ , \new_[623]_ , \new_[624]_ , \new_[625]_ ,
    \new_[626]_ , \new_[627]_ , \new_[628]_ , \new_[629]_ , \new_[630]_ ,
    \new_[631]_ , \new_[632]_ , \new_[633]_ , \new_[634]_ , \new_[635]_ ,
    \new_[636]_ , \new_[637]_ , \new_[638]_ , \new_[639]_ , \new_[640]_ ,
    \new_[641]_ , \new_[642]_ , \new_[643]_ , \new_[644]_ , \new_[645]_ ,
    \new_[646]_ , \new_[647]_ , \new_[648]_ , \new_[649]_ , \new_[650]_ ,
    \new_[651]_ , \new_[652]_ , \new_[653]_ , \new_[654]_ , \new_[655]_ ,
    \new_[656]_ , \new_[657]_ , \new_[658]_ , \new_[659]_ , \new_[660]_ ,
    \new_[661]_ , \new_[662]_ , \new_[663]_ , \new_[664]_ , \new_[665]_ ,
    \new_[666]_ , \new_[667]_ , \new_[668]_ , \new_[669]_ , \new_[670]_ ,
    \new_[671]_ , \new_[672]_ , \new_[673]_ , \new_[674]_ , \new_[675]_ ,
    \new_[676]_ , \new_[677]_ , \new_[678]_ , \new_[679]_ , \new_[680]_ ,
    \new_[681]_ , \new_[682]_ , \new_[683]_ , \new_[684]_ , \new_[685]_ ,
    \new_[686]_ , \new_[687]_ , \new_[688]_ , \new_[689]_ , \new_[690]_ ,
    \new_[691]_ , \new_[692]_ , \new_[693]_ , \new_[694]_ , \new_[695]_ ,
    \new_[696]_ , \new_[697]_ , \new_[698]_ , \new_[699]_ , \new_[700]_ ,
    \new_[701]_ , \new_[702]_ , \new_[703]_ , \new_[704]_ , \new_[705]_ ,
    \new_[706]_ , \new_[707]_ , \new_[708]_ , \new_[709]_ , \new_[710]_ ,
    \new_[711]_ , \new_[712]_ , \new_[713]_ , \new_[714]_ , \new_[715]_ ,
    \new_[716]_ , \new_[717]_ , \new_[718]_ , \new_[719]_ , \new_[720]_ ,
    \new_[721]_ , \new_[722]_ , \new_[723]_ , \new_[724]_ , \new_[725]_ ,
    \new_[726]_ , \new_[727]_ , \new_[728]_ , \new_[729]_ , \new_[730]_ ,
    \new_[731]_ , \new_[732]_ , \new_[733]_ , \new_[734]_ , \new_[735]_ ,
    \new_[736]_ , \new_[737]_ , \new_[738]_ , \new_[739]_ , \new_[740]_ ,
    \new_[741]_ , \new_[742]_ , \new_[743]_ , \new_[744]_ , \new_[745]_ ,
    \new_[746]_ , \new_[747]_ , \new_[748]_ , \new_[749]_ , \new_[750]_ ,
    \new_[751]_ , \new_[752]_ , \new_[753]_ , \new_[754]_ , \new_[755]_ ,
    \new_[756]_ , \new_[757]_ , \new_[758]_ , \new_[759]_ , \new_[760]_ ,
    \new_[761]_ , \new_[762]_ , \new_[763]_ , \new_[764]_ , \new_[765]_ ,
    \new_[766]_ , \new_[767]_ , \new_[768]_ , \new_[769]_ , \new_[770]_ ,
    \new_[771]_ , \new_[772]_ , \new_[773]_ , \new_[774]_ , \new_[775]_ ,
    \new_[776]_ , \new_[777]_ , \new_[778]_ , \new_[779]_ , \new_[780]_ ,
    \new_[781]_ , \new_[782]_ , \new_[783]_ , \new_[784]_ , \new_[785]_ ,
    \new_[786]_ , \new_[787]_ , \new_[788]_ , \new_[789]_ , \new_[790]_ ,
    \new_[791]_ , \new_[792]_ , \new_[793]_ , \new_[794]_ , \new_[795]_ ,
    \new_[796]_ , \new_[797]_ , \new_[798]_ , \new_[799]_ , \new_[800]_ ,
    \new_[801]_ , \new_[802]_ , \new_[803]_ , \new_[804]_ , \new_[805]_ ,
    \new_[806]_ , \new_[807]_ , \new_[808]_ , \new_[809]_ , \new_[810]_ ,
    \new_[811]_ , \new_[812]_ , \new_[813]_ , \new_[814]_ , \new_[815]_ ,
    \new_[816]_ , \new_[817]_ , \new_[818]_ , \new_[819]_ , \new_[820]_ ,
    \new_[821]_ , \new_[822]_ , \new_[823]_ , \new_[824]_ , \new_[825]_ ,
    \new_[826]_ , \new_[827]_ , \new_[828]_ , \new_[829]_ , \new_[830]_ ,
    \new_[831]_ , \new_[832]_ , \new_[833]_ , \new_[834]_ , \new_[835]_ ,
    \new_[836]_ , \new_[837]_ , \new_[838]_ , \new_[839]_ , \new_[840]_ ,
    \new_[841]_ , \new_[842]_ , \new_[843]_ , \new_[844]_ , \new_[845]_ ,
    \new_[846]_ , \new_[847]_ , \new_[848]_ , \new_[849]_ , \new_[850]_ ,
    \new_[851]_ , \new_[852]_ , \new_[853]_ , \new_[854]_ , \new_[855]_ ,
    \new_[856]_ , \new_[857]_ , \new_[858]_ , \new_[859]_ , \new_[860]_ ,
    \new_[861]_ , \new_[862]_ , \new_[863]_ , \new_[864]_ , \new_[865]_ ,
    \new_[866]_ , \new_[867]_ , \new_[868]_ , \new_[869]_ , \new_[870]_ ,
    \new_[871]_ , \new_[872]_ , \new_[873]_ , \new_[874]_ , \new_[875]_ ,
    \new_[876]_ , \new_[877]_ , \new_[878]_ , \new_[879]_ , \new_[880]_ ,
    \new_[881]_ , \new_[882]_ , \new_[883]_ , \new_[884]_ , \new_[885]_ ,
    \new_[886]_ , \new_[887]_ , \new_[888]_ , \new_[889]_ , \new_[890]_ ,
    \new_[891]_ , \new_[892]_ , \new_[893]_ , \new_[894]_ , \new_[895]_ ,
    \new_[896]_ , \new_[897]_ , \new_[898]_ , \new_[899]_ , \new_[900]_ ,
    \new_[901]_ , \new_[902]_ , \new_[903]_ , \new_[904]_ , \new_[905]_ ,
    \new_[906]_ , \new_[907]_ , \new_[908]_ , \new_[909]_ , \new_[910]_ ,
    \new_[911]_ , \new_[912]_ , \new_[913]_ , \new_[914]_ , \new_[915]_ ,
    \new_[916]_ , \new_[917]_ , \new_[918]_ , \new_[919]_ , \new_[920]_ ,
    \new_[921]_ , \new_[922]_ , \new_[923]_ , \new_[924]_ , \new_[925]_ ,
    \new_[926]_ , \new_[927]_ , \new_[928]_ , \new_[929]_ , \new_[930]_ ,
    \new_[931]_ , \new_[932]_ , \new_[933]_ , \new_[934]_ , \new_[935]_ ,
    \new_[936]_ , \new_[937]_ , \new_[938]_ , \new_[939]_ , \new_[940]_ ,
    \new_[941]_ , \new_[942]_ , \new_[943]_ , \new_[944]_ , \new_[945]_ ,
    \new_[946]_ , \new_[947]_ , \new_[948]_ , \new_[949]_ , \new_[950]_ ,
    \new_[951]_ , \new_[952]_ , \new_[953]_ , \new_[954]_ , \new_[955]_ ,
    \new_[956]_ , \new_[957]_ , \new_[958]_ , \new_[959]_ , \new_[960]_ ,
    \new_[961]_ , \new_[962]_ , \new_[963]_ , \new_[964]_ , \new_[965]_ ,
    \new_[966]_ , \new_[967]_ , \new_[968]_ , \new_[969]_ , \new_[970]_ ,
    \new_[971]_ , \new_[972]_ , \new_[973]_ , \new_[974]_ , \new_[975]_ ,
    \new_[976]_ , \new_[977]_ , \new_[978]_ , \new_[979]_ , \new_[980]_ ,
    \new_[981]_ , \new_[982]_ , \new_[983]_ , \new_[984]_ , \new_[985]_ ,
    \new_[986]_ , \new_[987]_ , \new_[988]_ , \new_[989]_ , \new_[990]_ ,
    \new_[991]_ , \new_[992]_ , \new_[993]_ , \new_[994]_ , \new_[995]_ ,
    \new_[996]_ , \new_[997]_ , \new_[998]_ , \new_[999]_ , \new_[1000]_ ,
    \new_[1001]_ , \new_[1002]_ , \new_[1003]_ , \new_[1004]_ ,
    \new_[1005]_ , \new_[1006]_ , \new_[1007]_ , \new_[1008]_ ,
    \new_[1009]_ , \new_[1010]_ , \new_[1011]_ , \new_[1012]_ ,
    \new_[1013]_ , \new_[1014]_ , \new_[1015]_ , \new_[1016]_ ,
    \new_[1017]_ , \new_[1018]_ , \new_[1019]_ , \new_[1020]_ ,
    \new_[1021]_ , \new_[1022]_ , \new_[1023]_ , \new_[1024]_ ,
    \new_[1025]_ , \new_[1026]_ , \new_[1027]_ , \new_[1028]_ ,
    \new_[1029]_ , \new_[1030]_ , \new_[1031]_ , \new_[1032]_ ,
    \new_[1033]_ , \new_[1034]_ , \new_[1035]_ , \new_[1036]_ ,
    \new_[1037]_ , \new_[1038]_ , \new_[1039]_ , \new_[1040]_ ,
    \new_[1041]_ , \new_[1042]_ , \new_[1043]_ , \new_[1044]_ ,
    \new_[1045]_ , \new_[1046]_ , \new_[1047]_ , \new_[1048]_ ,
    \new_[1049]_ , \new_[1050]_ , \new_[1051]_ , \new_[1052]_ ,
    \new_[1053]_ , \new_[1054]_ , \new_[1055]_ , \new_[1056]_ ,
    \new_[1057]_ , \new_[1058]_ , \new_[1059]_ , \new_[1060]_ ,
    \new_[1061]_ , \new_[1062]_ , \new_[1063]_ , \new_[1064]_ ,
    \new_[1065]_ , \new_[1066]_ , \new_[1067]_ , \new_[1068]_ ,
    \new_[1069]_ , \new_[1070]_ , \new_[1071]_ , \new_[1072]_ ,
    \new_[1073]_ , \new_[1074]_ , \new_[1075]_ , \new_[1076]_ ,
    \new_[1077]_ , \new_[1078]_ , \new_[1079]_ , \new_[1080]_ ,
    \new_[1081]_ , \new_[1082]_ , \new_[1083]_ , \new_[1084]_ ,
    \new_[1085]_ , \new_[1086]_ , \new_[1087]_ , \new_[1088]_ ,
    \new_[1089]_ , \new_[1090]_ , \new_[1091]_ , \new_[1092]_ ,
    \new_[1093]_ , \new_[1094]_ , \new_[1095]_ , \new_[1096]_ ,
    \new_[1097]_ , \new_[1098]_ , \new_[1099]_ , \new_[1100]_ ,
    \new_[1101]_ , \new_[1102]_ , \new_[1103]_ , \new_[1104]_ ,
    \new_[1105]_ , \new_[1106]_ , \new_[1107]_ , \new_[1108]_ ,
    \new_[1109]_ , \new_[1110]_ , \new_[1111]_ , \new_[1112]_ ,
    \new_[1113]_ , \new_[1114]_ , \new_[1115]_ , \new_[1116]_ ,
    \new_[1117]_ , \new_[1118]_ , \new_[1119]_ , \new_[1120]_ ,
    \new_[1121]_ , \new_[1122]_ , \new_[1123]_ , \new_[1124]_ ,
    \new_[1125]_ , \new_[1126]_ , \new_[1127]_ , \new_[1128]_ ,
    \new_[1129]_ , \new_[1130]_ , \new_[1131]_ , \new_[1132]_ ,
    \new_[1133]_ , \new_[1134]_ , \new_[1135]_ , \new_[1136]_ ,
    \new_[1137]_ , \new_[1138]_ , \new_[1139]_ , \new_[1140]_ ,
    \new_[1141]_ , \new_[1142]_ , \new_[1143]_ , \new_[1144]_ ,
    \new_[1145]_ , \new_[1146]_ , \new_[1147]_ , \new_[1148]_ ,
    \new_[1149]_ , \new_[1150]_ , \new_[1151]_ , \new_[1152]_ ,
    \new_[1153]_ , \new_[1154]_ , \new_[1155]_ , \new_[1156]_ ,
    \new_[1157]_ , \new_[1158]_ , \new_[1159]_ , \new_[1160]_ ,
    \new_[1161]_ , \new_[1162]_ , \new_[1163]_ , \new_[1164]_ ,
    \new_[1165]_ , \new_[1166]_ , \new_[1167]_ , \new_[1168]_ ,
    \new_[1169]_ , \new_[1170]_ , \new_[1171]_ , \new_[1172]_ ,
    \new_[1173]_ , \new_[1174]_ , \new_[1175]_ , \new_[1176]_ ,
    \new_[1177]_ , \new_[1178]_ , \new_[1179]_ , \new_[1180]_ ,
    \new_[1181]_ , \new_[1182]_ , \new_[1183]_ , \new_[1184]_ ,
    \new_[1185]_ , \new_[1186]_ , \new_[1187]_ , \new_[1188]_ ,
    \new_[1189]_ , \new_[1190]_ , \new_[1191]_ , \new_[1192]_ ,
    \new_[1193]_ , \new_[1194]_ , \new_[1195]_ , \new_[1196]_ ,
    \new_[1197]_ , \new_[1198]_ , \new_[1199]_ , \new_[1200]_ ,
    \new_[1201]_ , \new_[1202]_ , \new_[1203]_ , \new_[1204]_ ,
    \new_[1205]_ , \new_[1206]_ , \new_[1207]_ , \new_[1208]_ ,
    \new_[1209]_ , \new_[1210]_ , \new_[1211]_ , \new_[1212]_ ,
    \new_[1213]_ , \new_[1214]_ , \new_[1215]_ , \new_[1216]_ ,
    \new_[1217]_ , \new_[1218]_ , \new_[1219]_ , \new_[1220]_ ,
    \new_[1221]_ , \new_[1222]_ , \new_[1223]_ , \new_[1224]_ ,
    \new_[1225]_ , \new_[1226]_ , \new_[1227]_ , \new_[1228]_ ,
    \new_[1229]_ , \new_[1230]_ , \new_[1231]_ , \new_[1232]_ ,
    \new_[1233]_ , \new_[1234]_ , \new_[1235]_ , \new_[1236]_ ,
    \new_[1237]_ , \new_[1238]_ , \new_[1239]_ , \new_[1240]_ ,
    \new_[1241]_ , \new_[1242]_ , \new_[1243]_ , \new_[1244]_ ,
    \new_[1245]_ , \new_[1246]_ , \new_[1247]_ , \new_[1248]_ ,
    \new_[1249]_ , \new_[1250]_ , \new_[1251]_ , \new_[1252]_ ,
    \new_[1253]_ , \new_[1254]_ , \new_[1255]_ , \new_[1256]_ ,
    \new_[1257]_ , \new_[1258]_ , \new_[1259]_ , \new_[1260]_ ,
    \new_[1261]_ , \new_[1262]_ , \new_[1263]_ , \new_[1264]_ ,
    \new_[1265]_ , \new_[1266]_ , \new_[1267]_ , \new_[1268]_ ,
    \new_[1269]_ , \new_[1270]_ , \new_[1271]_ , \new_[1272]_ ,
    \new_[1273]_ , \new_[1274]_ , \new_[1275]_ , \new_[1276]_ ,
    \new_[1277]_ , \new_[1278]_ , \new_[1279]_ , \new_[1280]_ ,
    \new_[1281]_ , \new_[1282]_ , \new_[1283]_ , \new_[1284]_ ,
    \new_[1285]_ , \new_[1286]_ , \new_[1287]_ , \new_[1288]_ ,
    \new_[1289]_ , \new_[1290]_ , \new_[1291]_ , \new_[1292]_ ,
    \new_[1293]_ , \new_[1294]_ , \new_[1295]_ , \new_[1296]_ ,
    \new_[1297]_ , \new_[1298]_ , \new_[1299]_ , \new_[1300]_ ,
    \new_[1301]_ , \new_[1302]_ , \new_[1303]_ , \new_[1304]_ ,
    \new_[1305]_ , \new_[1306]_ , \new_[1307]_ , \new_[1308]_ ,
    \new_[1309]_ , \new_[1310]_ , \new_[1311]_ , \new_[1312]_ ,
    \new_[1313]_ , \new_[1314]_ , \new_[1315]_ , \new_[1316]_ ,
    \new_[1317]_ , \new_[1318]_ , \new_[1319]_ , \new_[1320]_ ,
    \new_[1321]_ , \new_[1322]_ , \new_[1323]_ , \new_[1324]_ ,
    \new_[1325]_ , \new_[1326]_ , \new_[1327]_ , \new_[1328]_ ,
    \new_[1329]_ , \new_[1330]_ , \new_[1331]_ , \new_[1332]_ ,
    \new_[1333]_ , \new_[1334]_ , \new_[1335]_ , \new_[1336]_ ,
    \new_[1337]_ , \new_[1338]_ , \new_[1339]_ , \new_[1340]_ ,
    \new_[1341]_ , \new_[1342]_ , \new_[1343]_ , \new_[1344]_ ,
    \new_[1345]_ , \new_[1346]_ , \new_[1347]_ , \new_[1348]_ ,
    \new_[1349]_ , \new_[1350]_ , \new_[1351]_ , \new_[1352]_ ,
    \new_[1353]_ , \new_[1354]_ , \new_[1355]_ , \new_[1356]_ ,
    \new_[1357]_ , \new_[1358]_ , \new_[1359]_ , \new_[1360]_ ,
    \new_[1361]_ , \new_[1362]_ , \new_[1363]_ , \new_[1364]_ ,
    \new_[1365]_ , \new_[1366]_ , \new_[1367]_ , \new_[1368]_ ,
    \new_[1369]_ , \new_[1370]_ , \new_[1371]_ , \new_[1372]_ ,
    \new_[1373]_ , \new_[1374]_ , \new_[1375]_ , \new_[1376]_ ,
    \new_[1377]_ , \new_[1378]_ , \new_[1379]_ , \new_[1380]_ ,
    \new_[1381]_ , \new_[1382]_ , \new_[1383]_ , \new_[1384]_ ,
    \new_[1385]_ , \new_[1386]_ , \new_[1387]_ , \new_[1388]_ ,
    \new_[1389]_ , \new_[1390]_ , \new_[1391]_ , \new_[1392]_ ,
    \new_[1393]_ , \new_[1394]_ , \new_[1395]_ , \new_[1396]_ ,
    \new_[1397]_ , \new_[1398]_ , \new_[1399]_ , \new_[1400]_ ,
    \new_[1401]_ , \new_[1402]_ , \new_[1403]_ , \new_[1404]_ ,
    \new_[1405]_ , \new_[1406]_ , \new_[1407]_ , \new_[1408]_ ,
    \new_[1409]_ , \new_[1410]_ , \new_[1411]_ , \new_[1412]_ ,
    \new_[1413]_ , \new_[1414]_ , \new_[1415]_ , \new_[1416]_ ,
    \new_[1417]_ , \new_[1418]_ , \new_[1419]_ , \new_[1420]_ ,
    \new_[1421]_ , \new_[1422]_ , \new_[1423]_ , \new_[1424]_ ,
    \new_[1425]_ , \new_[1426]_ , \new_[1427]_ , \new_[1428]_ ,
    \new_[1429]_ , \new_[1430]_ , \new_[1431]_ , \new_[1432]_ ,
    \new_[1433]_ , \new_[1434]_ , \new_[1435]_ , \new_[1436]_ ,
    \new_[1437]_ , \new_[1438]_ , \new_[1439]_ , \new_[1440]_ ,
    \new_[1441]_ , \new_[1442]_ , \new_[1443]_ , \new_[1444]_ ,
    \new_[1445]_ , \new_[1446]_ , \new_[1447]_ , \new_[1448]_ ,
    \new_[1449]_ , \new_[1450]_ , \new_[1451]_ , \new_[1452]_ ,
    \new_[1453]_ , \new_[1454]_ , \new_[1455]_ , \new_[1456]_ ,
    \new_[1457]_ , \new_[1458]_ , \new_[1459]_ , \new_[1460]_ ,
    \new_[1461]_ , \new_[1462]_ , \new_[1463]_ , \new_[1464]_ ,
    \new_[1465]_ , \new_[1466]_ , \new_[1467]_ , \new_[1468]_ ,
    \new_[1469]_ , \new_[1470]_ , \new_[1471]_ , \new_[1472]_ ,
    \new_[1473]_ , \new_[1474]_ , \new_[1475]_ , \new_[1476]_ ,
    \new_[1477]_ , \new_[1478]_ , \new_[1479]_ , \new_[1480]_ ,
    \new_[1481]_ , \new_[1482]_ , \new_[1483]_ , \new_[1484]_ ,
    \new_[1485]_ , \new_[1486]_ , \new_[1487]_ , \new_[1488]_ ,
    \new_[1489]_ , \new_[1490]_ , \new_[1491]_ , \new_[1492]_ ,
    \new_[1493]_ , \new_[1494]_ , \new_[1495]_ , \new_[1496]_ ,
    \new_[1497]_ , \new_[1498]_ , \new_[1499]_ , \new_[1500]_ ,
    \new_[1501]_ , \new_[1502]_ , \new_[1503]_ , \new_[1504]_ ,
    \new_[1505]_ , \new_[1506]_ , \new_[1507]_ , \new_[1508]_ ,
    \new_[1509]_ , \new_[1510]_ , \new_[1511]_ , \new_[1512]_ ,
    \new_[1513]_ , \new_[1514]_ , \new_[1515]_ , \new_[1516]_ ,
    \new_[1517]_ , \new_[1518]_ , \new_[1519]_ , \new_[1520]_ ,
    \new_[1521]_ , \new_[1522]_ , \new_[1523]_ , \new_[1524]_ ,
    \new_[1525]_ , \new_[1526]_ , \new_[1527]_ , \new_[1528]_ ,
    \new_[1529]_ , \new_[1530]_ , \new_[1531]_ , \new_[1532]_ ,
    \new_[1533]_ , \new_[1534]_ , \new_[1535]_ , \new_[1536]_ ,
    \new_[1537]_ , \new_[1538]_ , \new_[1539]_ , \new_[1540]_ ,
    \new_[1541]_ , \new_[1542]_ , \new_[1543]_ , \new_[1544]_ ,
    \new_[1545]_ , \new_[1546]_ , \new_[1547]_ , \new_[1548]_ ,
    \new_[1549]_ , \new_[1550]_ , \new_[1551]_ , \new_[1552]_ ,
    \new_[1553]_ , \new_[1554]_ , \new_[1555]_ , \new_[1556]_ ,
    \new_[1557]_ , \new_[1558]_ , \new_[1559]_ , \new_[1560]_ ,
    \new_[1561]_ , \new_[1562]_ , \new_[1563]_ , \new_[1564]_ ,
    \new_[1565]_ , \new_[1566]_ , \new_[1567]_ , \new_[1568]_ ,
    \new_[1569]_ , \new_[1570]_ , \new_[1571]_ , \new_[1572]_ ,
    \new_[1573]_ , \new_[1574]_ , \new_[1575]_ , \new_[1576]_ ,
    \new_[1577]_ , \new_[1578]_ , \new_[1579]_ , \new_[1580]_ ,
    \new_[1581]_ , \new_[1582]_ , \new_[1583]_ , \new_[1584]_ ,
    \new_[1585]_ , \new_[1586]_ , \new_[1587]_ , \new_[1588]_ ,
    \new_[1589]_ , \new_[1590]_ , \new_[1591]_ , \new_[1592]_ ,
    \new_[1593]_ , \new_[1594]_ , \new_[1595]_ , \new_[1596]_ ,
    \new_[1597]_ , \new_[1598]_ , \new_[1599]_ , \new_[1600]_ ,
    \new_[1601]_ , \new_[1602]_ , \new_[1603]_ , \new_[1604]_ ,
    \new_[1605]_ , \new_[1606]_ , \new_[1607]_ , \new_[1608]_ ,
    \new_[1609]_ , \new_[1610]_ , \new_[1611]_ , \new_[1612]_ ,
    \new_[1613]_ , \new_[1614]_ , \new_[1615]_ , \new_[1616]_ ,
    \new_[1617]_ , \new_[1618]_ , \new_[1619]_ , \new_[1620]_ ,
    \new_[1621]_ , \new_[1622]_ , \new_[1623]_ , \new_[1624]_ ,
    \new_[1625]_ , \new_[1626]_ , \new_[1627]_ , \new_[1628]_ ,
    \new_[1629]_ , \new_[1630]_ , \new_[1631]_ , \new_[1632]_ ,
    \new_[1633]_ , \new_[1634]_ , \new_[1635]_ , \new_[1636]_ ,
    \new_[1637]_ , \new_[1638]_ , \new_[1639]_ , \new_[1640]_ ,
    \new_[1641]_ , \new_[1642]_ , \new_[1643]_ , \new_[1644]_ ,
    \new_[1645]_ , \new_[1646]_ , \new_[1647]_ , \new_[1648]_ ,
    \new_[1649]_ , \new_[1650]_ , \new_[1651]_ , \new_[1652]_ ,
    \new_[1653]_ , \new_[1654]_ , \new_[1655]_ , \new_[1656]_ ,
    \new_[1657]_ , \new_[1658]_ , \new_[1659]_ , \new_[1660]_ ,
    \new_[1661]_ , \new_[1662]_ , \new_[1663]_ , \new_[1664]_ ,
    \new_[1665]_ , \new_[1666]_ , \new_[1667]_ , \new_[1668]_ ,
    \new_[1669]_ , \new_[1670]_ , \new_[1671]_ , \new_[1672]_ ,
    \new_[1673]_ , \new_[1674]_ , \new_[1675]_ , \new_[1676]_ ,
    \new_[1677]_ , \new_[1678]_ , \new_[1679]_ , \new_[1680]_ ,
    \new_[1681]_ , \new_[1682]_ , \new_[1683]_ , \new_[1684]_ ,
    \new_[1685]_ , \new_[1686]_ , \new_[1687]_ , \new_[1688]_ ,
    \new_[1689]_ , \new_[1690]_ , \new_[1691]_ , \new_[1692]_ ,
    \new_[1693]_ , \new_[1694]_ , \new_[1695]_ , \new_[1696]_ ,
    \new_[1697]_ , \new_[1698]_ , \new_[1699]_ , \new_[1700]_ ,
    \new_[1701]_ , \new_[1702]_ , \new_[1703]_ , \new_[1704]_ ,
    \new_[1705]_ , \new_[1706]_ , \new_[1707]_ , \new_[1708]_ ,
    \new_[1709]_ , \new_[1710]_ , \new_[1711]_ , \new_[1712]_ ,
    \new_[1713]_ , \new_[1714]_ , \new_[1715]_ , \new_[1716]_ ,
    \new_[1717]_ , \new_[1718]_ , \new_[1719]_ , \new_[1720]_ ,
    \new_[1721]_ , \new_[1722]_ , \new_[1723]_ , \new_[1724]_ ,
    \new_[1725]_ , \new_[1726]_ , \new_[1727]_ , \new_[1728]_ ,
    \new_[1729]_ , \new_[1730]_ , \new_[1731]_ , \new_[1732]_ ,
    \new_[1733]_ , \new_[1734]_ , \new_[1735]_ , \new_[1736]_ ,
    \new_[1737]_ , \new_[1738]_ , \new_[1739]_ , \new_[1740]_ ,
    \new_[1741]_ , \new_[1742]_ , \new_[1743]_ , \new_[1744]_ ,
    \new_[1745]_ , \new_[1746]_ , \new_[1747]_ , \new_[1748]_ ,
    \new_[1749]_ , \new_[1750]_ , \new_[1751]_ , \new_[1752]_ ,
    \new_[1753]_ , \new_[1754]_ , \new_[1755]_ , \new_[1756]_ ,
    \new_[1757]_ , \new_[1758]_ , \new_[1759]_ , \new_[1760]_ ,
    \new_[1761]_ , \new_[1762]_ , \new_[1763]_ , \new_[1764]_ ,
    \new_[1765]_ , \new_[1766]_ , \new_[1767]_ , \new_[1768]_ ,
    \new_[1769]_ , \new_[1770]_ , \new_[1771]_ , \new_[1772]_ ,
    \new_[1773]_ , \new_[1774]_ , \new_[1775]_ , \new_[1776]_ ,
    \new_[1777]_ , \new_[1778]_ , \new_[1779]_ , \new_[1780]_ ,
    \new_[1781]_ , \new_[1782]_ , \new_[1783]_ , \new_[1784]_ ,
    \new_[1785]_ , \new_[1786]_ , \new_[1787]_ , \new_[1788]_ ,
    \new_[1789]_ , \new_[1790]_ , \new_[1791]_ , \new_[1792]_ ,
    \new_[1793]_ , \new_[1794]_ , \new_[1795]_ , \new_[1796]_ ,
    \new_[1797]_ , \new_[1798]_ , \new_[1799]_ , \new_[1800]_ ,
    \new_[1801]_ , \new_[1802]_ , \new_[1803]_ , \new_[1804]_ ,
    \new_[1805]_ , \new_[1806]_ , \new_[1807]_ , \new_[1808]_ ,
    \new_[1809]_ , \new_[1810]_ , \new_[1811]_ , \new_[1812]_ ,
    \new_[1813]_ , \new_[1814]_ , \new_[1815]_ , \new_[1816]_ ,
    \new_[1817]_ , \new_[1818]_ , \new_[1819]_ , \new_[1820]_ ,
    \new_[1821]_ , \new_[1822]_ , \new_[1823]_ , \new_[1824]_ ,
    \new_[1825]_ , \new_[1826]_ , \new_[1827]_ , \new_[1828]_ ,
    \new_[1829]_ , \new_[1830]_ , \new_[1831]_ , \new_[1832]_ ,
    \new_[1833]_ , \new_[1834]_ , \new_[1835]_ , \new_[1836]_ ,
    \new_[1837]_ , \new_[1838]_ , \new_[1839]_ , \new_[1840]_ ,
    \new_[1841]_ , \new_[1842]_ , \new_[1843]_ , \new_[1844]_ ,
    \new_[1845]_ , \new_[1846]_ , \new_[1847]_ , \new_[1848]_ ,
    \new_[1849]_ , \new_[1850]_ , \new_[1851]_ , \new_[1852]_ ,
    \new_[1853]_ , \new_[1854]_ , \new_[1855]_ , \new_[1856]_ ,
    \new_[1857]_ , \new_[1858]_ , \new_[1859]_ , \new_[1860]_ ,
    \new_[1861]_ , \new_[1862]_ , \new_[1863]_ , \new_[1864]_ ,
    \new_[1865]_ , \new_[1866]_ , \new_[1867]_ , \new_[1868]_ ,
    \new_[1869]_ , \new_[1870]_ , \new_[1871]_ , \new_[1872]_ ,
    \new_[1873]_ , \new_[1874]_ , \new_[1875]_ , \new_[1876]_ ,
    \new_[1877]_ , \new_[1878]_ , \new_[1879]_ , \new_[1880]_ ,
    \new_[1881]_ , \new_[1882]_ , \new_[1883]_ , \new_[1884]_ ,
    \new_[1885]_ , \new_[1886]_ , \new_[1887]_ , \new_[1888]_ ,
    \new_[1889]_ , \new_[1890]_ , \new_[1891]_ , \new_[1892]_ ,
    \new_[1893]_ , \new_[1894]_ , \new_[1895]_ , \new_[1896]_ ,
    \new_[1897]_ , \new_[1898]_ , \new_[1899]_ , \new_[1900]_ ,
    \new_[1901]_ , \new_[1902]_ , \new_[1903]_ , \new_[1904]_ ,
    \new_[1905]_ , \new_[1906]_ , \new_[1907]_ , \new_[1908]_ ,
    \new_[1909]_ , \new_[1910]_ , \new_[1911]_ , \new_[1912]_ ,
    \new_[1913]_ , \new_[1914]_ , \new_[1915]_ , \new_[1916]_ ,
    \new_[1917]_ , \new_[1918]_ , \new_[1919]_ , \new_[1920]_ ,
    \new_[1921]_ , \new_[1922]_ , \new_[1923]_ , \new_[1924]_ ,
    \new_[1925]_ , \new_[1926]_ , \new_[1927]_ , \new_[1928]_ ,
    \new_[1929]_ , \new_[1930]_ , \new_[1931]_ , \new_[1932]_ ,
    \new_[1933]_ , \new_[1934]_ , \new_[1935]_ , \new_[1936]_ ,
    \new_[1937]_ , \new_[1938]_ , \new_[1939]_ , \new_[1940]_ ,
    \new_[1941]_ , \new_[1942]_ , \new_[1943]_ , \new_[1944]_ ,
    \new_[1945]_ , \new_[1946]_ , \new_[1947]_ , \new_[1948]_ ,
    \new_[1949]_ , \new_[1950]_ , \new_[1951]_ , \new_[1952]_ ,
    \new_[1953]_ , \new_[1954]_ , \new_[1955]_ , \new_[1956]_ ,
    \new_[1957]_ , \new_[1958]_ , \new_[1959]_ , \new_[1960]_ ,
    \new_[1961]_ , \new_[1962]_ , \new_[1963]_ , \new_[1964]_ ,
    \new_[1965]_ , \new_[1966]_ , \new_[1967]_ , \new_[1968]_ ,
    \new_[1969]_ , \new_[1970]_ , \new_[1971]_ , \new_[1972]_ ,
    \new_[1973]_ , \new_[1974]_ , \new_[1975]_ , \new_[1976]_ ,
    \new_[1977]_ , \new_[1978]_ , \new_[1979]_ , \new_[1980]_ ,
    \new_[1981]_ , \new_[1982]_ , \new_[1983]_ , \new_[1984]_ ,
    \new_[1985]_ , \new_[1986]_ , \new_[1987]_ , \new_[1988]_ ,
    \new_[1989]_ , \new_[1990]_ , \new_[1991]_ , \new_[1992]_ ,
    \new_[1993]_ , \new_[1994]_ , \new_[1995]_ , \new_[1996]_ ,
    \new_[1997]_ , \new_[1998]_ , \new_[1999]_ , \new_[2000]_ ,
    \new_[2001]_ , \new_[2002]_ , \new_[2003]_ , \new_[2004]_ ,
    \new_[2005]_ , \new_[2006]_ , \new_[2007]_ , \new_[2008]_ ,
    \new_[2009]_ , \new_[2010]_ , \new_[2011]_ , \new_[2012]_ ,
    \new_[2013]_ , \new_[2014]_ , \new_[2015]_ , \new_[2016]_ ,
    \new_[2017]_ , \new_[2018]_ , \new_[2019]_ , \new_[2020]_ ,
    \new_[2021]_ , \new_[2022]_ , \new_[2023]_ , \new_[2024]_ ,
    \new_[2025]_ , \new_[2026]_ , \new_[2027]_ , \new_[2028]_ ,
    \new_[2029]_ , \new_[2030]_ , \new_[2031]_ , \new_[2032]_ ,
    \new_[2033]_ , \new_[2034]_ , \new_[2035]_ , \new_[2036]_ ,
    \new_[2037]_ , \new_[2038]_ , \new_[2039]_ , \new_[2040]_ ,
    \new_[2041]_ , \new_[2042]_ , \new_[2043]_ , \new_[2044]_ ,
    \new_[2045]_ , \new_[2046]_ , \new_[2047]_ , \new_[2048]_ ,
    \new_[2049]_ , \new_[2050]_ , \new_[2051]_ , \new_[2052]_ ,
    \new_[2053]_ , \new_[2054]_ , \new_[2055]_ , \new_[2056]_ ,
    \new_[2057]_ , \new_[2058]_ , \new_[2059]_ , \new_[2060]_ ,
    \new_[2061]_ , \new_[2062]_ , \new_[2063]_ , \new_[2064]_ ,
    \new_[2065]_ , \new_[2066]_ , \new_[2067]_ , \new_[2068]_ ,
    \new_[2069]_ , \new_[2070]_ , \new_[2071]_ , \new_[2072]_ ,
    \new_[2073]_ , \new_[2074]_ , \new_[2075]_ , \new_[2076]_ ,
    \new_[2077]_ , \new_[2078]_ , \new_[2079]_ , \new_[2080]_ ,
    \new_[2081]_ , \new_[2082]_ , \new_[2083]_ , \new_[2084]_ ,
    \new_[2085]_ , \new_[2086]_ , \new_[2087]_ , \new_[2088]_ ,
    \new_[2089]_ , \new_[2090]_ , \new_[2091]_ , \new_[2092]_ ,
    \new_[2093]_ , \new_[2094]_ , \new_[2095]_ , \new_[2096]_ ,
    \new_[2097]_ , \new_[2098]_ , \new_[2099]_ , \new_[2100]_ ,
    \new_[2101]_ , \new_[2102]_ , \new_[2103]_ , \new_[2104]_ ,
    \new_[2105]_ , \new_[2106]_ , \new_[2107]_ , \new_[2108]_ ,
    \new_[2109]_ , \new_[2110]_ , \new_[2111]_ , \new_[2112]_ ,
    \new_[2113]_ , \new_[2114]_ , \new_[2115]_ , \new_[2116]_ ,
    \new_[2117]_ , \new_[2118]_ , \new_[2119]_ , \new_[2120]_ ,
    \new_[2121]_ , \new_[2122]_ , \new_[2123]_ , \new_[2124]_ ,
    \new_[2125]_ , \new_[2126]_ , \new_[2127]_ , \new_[2128]_ ,
    \new_[2129]_ , \new_[2130]_ , \new_[2131]_ , \new_[2132]_ ,
    \new_[2133]_ , \new_[2134]_ , \new_[2135]_ , \new_[2136]_ ,
    \new_[2137]_ , \new_[2138]_ , \new_[2139]_ , \new_[2140]_ ,
    \new_[2141]_ , \new_[2142]_ , \new_[2143]_ , \new_[2144]_ ,
    \new_[2145]_ , \new_[2146]_ , \new_[2147]_ , \new_[2148]_ ,
    \new_[2149]_ , \new_[2150]_ , \new_[2151]_ , \new_[2152]_ ,
    \new_[2153]_ , \new_[2154]_ , \new_[2155]_ , \new_[2156]_ ,
    \new_[2157]_ , \new_[2158]_ , \new_[2159]_ , \new_[2160]_ ,
    \new_[2161]_ , \new_[2162]_ , \new_[2163]_ , \new_[2164]_ ,
    \new_[2165]_ , \new_[2166]_ , \new_[2167]_ , \new_[2168]_ ,
    \new_[2169]_ , \new_[2170]_ , \new_[2171]_ , \new_[2172]_ ,
    \new_[2173]_ , \new_[2174]_ , \new_[2175]_ , \new_[2176]_ ,
    \new_[2177]_ , \new_[2178]_ , \new_[2179]_ , \new_[2180]_ ,
    \new_[2181]_ , \new_[2182]_ , \new_[2183]_ , \new_[2184]_ ,
    \new_[2185]_ , \new_[2186]_ , \new_[2187]_ , \new_[2188]_ ,
    \new_[2189]_ , \new_[2190]_ , \new_[2191]_ , \new_[2192]_ ,
    \new_[2193]_ , \new_[2194]_ , \new_[2195]_ , \new_[2196]_ ,
    \new_[2197]_ , \new_[2198]_ , \new_[2199]_ , \new_[2200]_ ,
    \new_[2201]_ , \new_[2202]_ , \new_[2203]_ , \new_[2204]_ ,
    \new_[2205]_ , \new_[2206]_ , \new_[2207]_ , \new_[2208]_ ,
    \new_[2209]_ , \new_[2210]_ , \new_[2211]_ , \new_[2212]_ ,
    \new_[2213]_ , \new_[2214]_ , \new_[2215]_ , \new_[2216]_ ,
    \new_[2217]_ , \new_[2218]_ , \new_[2219]_ , \new_[2220]_ ,
    \new_[2221]_ , \new_[2222]_ , \new_[2223]_ , \new_[2224]_ ,
    \new_[2225]_ , \new_[2226]_ , \new_[2227]_ , \new_[2228]_ ,
    \new_[2229]_ , \new_[2230]_ , \new_[2231]_ , \new_[2232]_ ,
    \new_[2233]_ , \new_[2234]_ , \new_[2235]_ , \new_[2236]_ ,
    \new_[2237]_ , \new_[2238]_ , \new_[2239]_ , \new_[2240]_ ,
    \new_[2241]_ , \new_[2242]_ , \new_[2243]_ , \new_[2244]_ ,
    \new_[2245]_ , \new_[2246]_ , \new_[2247]_ , \new_[2248]_ ,
    \new_[2249]_ , \new_[2250]_ , \new_[2251]_ , \new_[2252]_ ,
    \new_[2253]_ , \new_[2254]_ , \new_[2255]_ , \new_[2256]_ ,
    \new_[2257]_ , \new_[2258]_ , \new_[2259]_ , \new_[2260]_ ,
    \new_[2261]_ , \new_[2262]_ , \new_[2263]_ , \new_[2264]_ ,
    \new_[2265]_ , \new_[2266]_ , \new_[2267]_ , \new_[2268]_ ,
    \new_[2269]_ , \new_[2270]_ , \new_[2271]_ , \new_[2272]_ ,
    \new_[2273]_ , \new_[2274]_ , \new_[2275]_ , \new_[2276]_ ,
    \new_[2277]_ , \new_[2278]_ , \new_[2279]_ , \new_[2280]_ ,
    \new_[2281]_ , \new_[2282]_ , \new_[2283]_ , \new_[2284]_ ,
    \new_[2285]_ , \new_[2286]_ , \new_[2287]_ , \new_[2288]_ ,
    \new_[2289]_ , \new_[2290]_ , \new_[2291]_ , \new_[2292]_ ,
    \new_[2293]_ , \new_[2294]_ , \new_[2295]_ , \new_[2296]_ ,
    \new_[2297]_ , \new_[2298]_ , \new_[2299]_ , \new_[2300]_ ,
    \new_[2301]_ , \new_[2302]_ , \new_[2303]_ , \new_[2304]_ ,
    \new_[2305]_ , \new_[2306]_ , \new_[2307]_ , \new_[2308]_ ,
    \new_[2309]_ , \new_[2310]_ , \new_[2311]_ , \new_[2312]_ ,
    \new_[2313]_ , \new_[2314]_ , \new_[2315]_ , \new_[2316]_ ,
    \new_[2317]_ , \new_[2318]_ , \new_[2319]_ , \new_[2320]_ ,
    \new_[2321]_ , \new_[2322]_ , \new_[2323]_ , \new_[2324]_ ,
    \new_[2325]_ , \new_[2326]_ , \new_[2327]_ , \new_[2328]_ ,
    \new_[2329]_ , \new_[2330]_ , \new_[2331]_ , \new_[2332]_ ,
    \new_[2333]_ , \new_[2334]_ , \new_[2335]_ , \new_[2336]_ ,
    \new_[2337]_ , \new_[2338]_ , \new_[2339]_ , \new_[2340]_ ,
    \new_[2341]_ , \new_[2342]_ , \new_[2343]_ , \new_[2344]_ ,
    \new_[2345]_ , \new_[2346]_ , \new_[2347]_ , \new_[2348]_ ,
    \new_[2349]_ , \new_[2350]_ , \new_[2351]_ , \new_[2352]_ ,
    \new_[2353]_ , \new_[2354]_ , \new_[2355]_ , \new_[2356]_ ,
    \new_[2357]_ , \new_[2358]_ , \new_[2359]_ , \new_[2360]_ ,
    \new_[2361]_ , \new_[2362]_ , \new_[2363]_ , \new_[2364]_ ,
    \new_[2365]_ , \new_[2366]_ , \new_[2367]_ , \new_[2368]_ ,
    \new_[2369]_ , \new_[2370]_ , \new_[2371]_ , \new_[2372]_ ,
    \new_[2373]_ , \new_[2374]_ , \new_[2375]_ , \new_[2376]_ ,
    \new_[2377]_ , \new_[2378]_ , \new_[2379]_ , \new_[2380]_ ,
    \new_[2381]_ , \new_[2382]_ , \new_[2383]_ , \new_[2384]_ ,
    \new_[2385]_ , \new_[2386]_ , \new_[2387]_ , \new_[2388]_ ,
    \new_[2389]_ , \new_[2390]_ , \new_[2391]_ , \new_[2392]_ ,
    \new_[2393]_ , \new_[2394]_ , \new_[2395]_ , \new_[2396]_ ,
    \new_[2397]_ , \new_[2398]_ , \new_[2399]_ , \new_[2400]_ ,
    \new_[2401]_ , \new_[2402]_ , \new_[2403]_ , \new_[2404]_ ,
    \new_[2405]_ , \new_[2406]_ , \new_[2407]_ , \new_[2408]_ ,
    \new_[2409]_ , \new_[2410]_ , \new_[2411]_ , \new_[2412]_ ,
    \new_[2413]_ , \new_[2414]_ , \new_[2415]_ , \new_[2416]_ ,
    \new_[2417]_ , \new_[2418]_ , \new_[2419]_ , \new_[2420]_ ,
    \new_[2421]_ , \new_[2422]_ , \new_[2423]_ , \new_[2424]_ ,
    \new_[2425]_ , \new_[2426]_ , \new_[2427]_ , \new_[2428]_ ,
    \new_[2429]_ , \new_[2430]_ , \new_[2431]_ , \new_[2432]_ ,
    \new_[2433]_ , \new_[2434]_ , \new_[2435]_ , \new_[2436]_ ,
    \new_[2437]_ , \new_[2438]_ , \new_[2439]_ , \new_[2440]_ ,
    \new_[2441]_ , \new_[2442]_ , \new_[2443]_ , \new_[2444]_ ,
    \new_[2445]_ , \new_[2446]_ , \new_[2447]_ , \new_[2448]_ ,
    \new_[2449]_ , \new_[2450]_ , \new_[2451]_ , \new_[2452]_ ,
    \new_[2453]_ , \new_[2454]_ , \new_[2455]_ , \new_[2456]_ ,
    \new_[2457]_ , \new_[2458]_ , \new_[2459]_ , \new_[2460]_ ,
    \new_[2461]_ , \new_[2462]_ , \new_[2463]_ , \new_[2464]_ ,
    \new_[2465]_ , \new_[2466]_ , \new_[2467]_ , \new_[2468]_ ,
    \new_[2469]_ , \new_[2470]_ , \new_[2471]_ , \new_[2472]_ ,
    \new_[2473]_ , \new_[2474]_ , \new_[2475]_ , \new_[2476]_ ,
    \new_[2477]_ , \new_[2478]_ , \new_[2479]_ , \new_[2480]_ ,
    \new_[2481]_ , \new_[2482]_ , \new_[2483]_ , \new_[2484]_ ,
    \new_[2485]_ , \new_[2486]_ , \new_[2487]_ , \new_[2488]_ ,
    \new_[2489]_ , \new_[2490]_ , \new_[2491]_ , \new_[2492]_ ,
    \new_[2493]_ , \new_[2494]_ , \new_[2495]_ , \new_[2496]_ ,
    \new_[2497]_ , \new_[2498]_ , \new_[2499]_ , \new_[2500]_ ,
    \new_[2501]_ , \new_[2502]_ , \new_[2503]_ , \new_[2504]_ ,
    \new_[2505]_ , \new_[2506]_ , \new_[2507]_ , \new_[2508]_ ,
    \new_[2509]_ , \new_[2510]_ , \new_[2511]_ , \new_[2512]_ ,
    \new_[2513]_ , \new_[2514]_ , \new_[2515]_ , \new_[2516]_ ,
    \new_[2517]_ , \new_[2518]_ , \new_[2519]_ , \new_[2520]_ ,
    \new_[2521]_ , \new_[2522]_ , \new_[2523]_ , \new_[2524]_ ,
    \new_[2525]_ , \new_[2526]_ , \new_[2527]_ , \new_[2528]_ ,
    \new_[2529]_ , \new_[2530]_ , \new_[2531]_ , \new_[2532]_ ,
    \new_[2533]_ , \new_[2534]_ , \new_[2535]_ , \new_[2536]_ ,
    \new_[2537]_ , \new_[2538]_ , \new_[2539]_ , \new_[2540]_ ,
    \new_[2541]_ , \new_[2542]_ , \new_[2543]_ , \new_[2544]_ ,
    \new_[2545]_ , \new_[2546]_ , \new_[2547]_ , \new_[2548]_ ,
    \new_[2549]_ , \new_[2550]_ , \new_[2553]_ , \new_[2556]_ ,
    \new_[2557]_ , \new_[2560]_ , \new_[2564]_ , \new_[2565]_ ,
    \new_[2566]_ , \new_[2567]_ , \new_[2570]_ , \new_[2574]_ ,
    \new_[2575]_ , \new_[2576]_ , \new_[2579]_ , \new_[2583]_ ,
    \new_[2584]_ , \new_[2585]_ , \new_[2586]_ , \new_[2587]_ ,
    \new_[2590]_ , \new_[2594]_ , \new_[2595]_ , \new_[2596]_ ,
    \new_[2599]_ , \new_[2603]_ , \new_[2604]_ , \new_[2605]_ ,
    \new_[2606]_ , \new_[2609]_ , \new_[2613]_ , \new_[2614]_ ,
    \new_[2615]_ , \new_[2618]_ , \new_[2622]_ , \new_[2623]_ ,
    \new_[2624]_ , \new_[2625]_ , \new_[2626]_ , \new_[2627]_ ,
    \new_[2630]_ , \new_[2634]_ , \new_[2635]_ , \new_[2636]_ ,
    \new_[2639]_ , \new_[2643]_ , \new_[2644]_ , \new_[2645]_ ,
    \new_[2646]_ , \new_[2649]_ , \new_[2653]_ , \new_[2654]_ ,
    \new_[2655]_ , \new_[2658]_ , \new_[2662]_ , \new_[2663]_ ,
    \new_[2664]_ , \new_[2665]_ , \new_[2666]_ , \new_[2669]_ ,
    \new_[2673]_ , \new_[2674]_ , \new_[2675]_ , \new_[2678]_ ,
    \new_[2682]_ , \new_[2683]_ , \new_[2684]_ , \new_[2685]_ ,
    \new_[2688]_ , \new_[2692]_ , \new_[2693]_ , \new_[2694]_ ,
    \new_[2697]_ , \new_[2701]_ , \new_[2702]_ , \new_[2703]_ ,
    \new_[2704]_ , \new_[2705]_ , \new_[2706]_ , \new_[2707]_ ,
    \new_[2710]_ , \new_[2714]_ , \new_[2715]_ , \new_[2716]_ ,
    \new_[2719]_ , \new_[2723]_ , \new_[2724]_ , \new_[2725]_ ,
    \new_[2726]_ , \new_[2729]_ , \new_[2733]_ , \new_[2734]_ ,
    \new_[2735]_ , \new_[2738]_ , \new_[2742]_ , \new_[2743]_ ,
    \new_[2744]_ , \new_[2745]_ , \new_[2746]_ , \new_[2749]_ ,
    \new_[2753]_ , \new_[2754]_ , \new_[2755]_ , \new_[2758]_ ,
    \new_[2762]_ , \new_[2763]_ , \new_[2764]_ , \new_[2765]_ ,
    \new_[2768]_ , \new_[2772]_ , \new_[2773]_ , \new_[2774]_ ,
    \new_[2777]_ , \new_[2781]_ , \new_[2782]_ , \new_[2783]_ ,
    \new_[2784]_ , \new_[2785]_ , \new_[2786]_ , \new_[2789]_ ,
    \new_[2793]_ , \new_[2794]_ , \new_[2795]_ , \new_[2798]_ ,
    \new_[2802]_ , \new_[2803]_ , \new_[2804]_ , \new_[2805]_ ,
    \new_[2808]_ , \new_[2812]_ , \new_[2813]_ , \new_[2814]_ ,
    \new_[2817]_ , \new_[2821]_ , \new_[2822]_ , \new_[2823]_ ,
    \new_[2824]_ , \new_[2825]_ , \new_[2828]_ , \new_[2832]_ ,
    \new_[2833]_ , \new_[2834]_ , \new_[2837]_ , \new_[2841]_ ,
    \new_[2842]_ , \new_[2843]_ , \new_[2844]_ , \new_[2847]_ ,
    \new_[2851]_ , \new_[2852]_ , \new_[2853]_ , \new_[2856]_ ,
    \new_[2860]_ , \new_[2861]_ , \new_[2862]_ , \new_[2863]_ ,
    \new_[2864]_ , \new_[2865]_ , \new_[2866]_ , \new_[2867]_ ,
    \new_[2870]_ , \new_[2873]_ , \new_[2874]_ , \new_[2877]_ ,
    \new_[2881]_ , \new_[2882]_ , \new_[2883]_ , \new_[2884]_ ,
    \new_[2887]_ , \new_[2891]_ , \new_[2892]_ , \new_[2893]_ ,
    \new_[2896]_ , \new_[2900]_ , \new_[2901]_ , \new_[2902]_ ,
    \new_[2903]_ , \new_[2904]_ , \new_[2907]_ , \new_[2911]_ ,
    \new_[2912]_ , \new_[2913]_ , \new_[2916]_ , \new_[2920]_ ,
    \new_[2921]_ , \new_[2922]_ , \new_[2923]_ , \new_[2926]_ ,
    \new_[2930]_ , \new_[2931]_ , \new_[2932]_ , \new_[2935]_ ,
    \new_[2939]_ , \new_[2940]_ , \new_[2941]_ , \new_[2942]_ ,
    \new_[2943]_ , \new_[2944]_ , \new_[2947]_ , \new_[2951]_ ,
    \new_[2952]_ , \new_[2953]_ , \new_[2956]_ , \new_[2960]_ ,
    \new_[2961]_ , \new_[2962]_ , \new_[2963]_ , \new_[2966]_ ,
    \new_[2970]_ , \new_[2971]_ , \new_[2972]_ , \new_[2975]_ ,
    \new_[2979]_ , \new_[2980]_ , \new_[2981]_ , \new_[2982]_ ,
    \new_[2983]_ , \new_[2986]_ , \new_[2990]_ , \new_[2991]_ ,
    \new_[2992]_ , \new_[2995]_ , \new_[2999]_ , \new_[3000]_ ,
    \new_[3001]_ , \new_[3002]_ , \new_[3005]_ , \new_[3009]_ ,
    \new_[3010]_ , \new_[3011]_ , \new_[3014]_ , \new_[3018]_ ,
    \new_[3019]_ , \new_[3020]_ , \new_[3021]_ , \new_[3022]_ ,
    \new_[3023]_ , \new_[3024]_ , \new_[3027]_ , \new_[3031]_ ,
    \new_[3032]_ , \new_[3033]_ , \new_[3036]_ , \new_[3040]_ ,
    \new_[3041]_ , \new_[3042]_ , \new_[3043]_ , \new_[3046]_ ,
    \new_[3050]_ , \new_[3051]_ , \new_[3052]_ , \new_[3055]_ ,
    \new_[3059]_ , \new_[3060]_ , \new_[3061]_ , \new_[3062]_ ,
    \new_[3063]_ , \new_[3066]_ , \new_[3070]_ , \new_[3071]_ ,
    \new_[3072]_ , \new_[3075]_ , \new_[3079]_ , \new_[3080]_ ,
    \new_[3081]_ , \new_[3082]_ , \new_[3085]_ , \new_[3089]_ ,
    \new_[3090]_ , \new_[3091]_ , \new_[3094]_ , \new_[3098]_ ,
    \new_[3099]_ , \new_[3100]_ , \new_[3101]_ , \new_[3102]_ ,
    \new_[3103]_ , \new_[3106]_ , \new_[3110]_ , \new_[3111]_ ,
    \new_[3112]_ , \new_[3115]_ , \new_[3119]_ , \new_[3120]_ ,
    \new_[3121]_ , \new_[3122]_ , \new_[3125]_ , \new_[3129]_ ,
    \new_[3130]_ , \new_[3131]_ , \new_[3134]_ , \new_[3138]_ ,
    \new_[3139]_ , \new_[3140]_ , \new_[3141]_ , \new_[3142]_ ,
    \new_[3145]_ , \new_[3149]_ , \new_[3150]_ , \new_[3151]_ ,
    \new_[3154]_ , \new_[3158]_ , \new_[3159]_ , \new_[3160]_ ,
    \new_[3161]_ , \new_[3164]_ , \new_[3168]_ , \new_[3169]_ ,
    \new_[3170]_ , \new_[3173]_ , \new_[3177]_ , \new_[3178]_ ,
    \new_[3179]_ , \new_[3180]_ , \new_[3181]_ , \new_[3182]_ ,
    \new_[3183]_ , \new_[3184]_ , \new_[3185]_ , \new_[3188]_ ,
    \new_[3191]_ , \new_[3192]_ , \new_[3195]_ , \new_[3199]_ ,
    \new_[3200]_ , \new_[3201]_ , \new_[3202]_ , \new_[3205]_ ,
    \new_[3209]_ , \new_[3210]_ , \new_[3211]_ , \new_[3214]_ ,
    \new_[3218]_ , \new_[3219]_ , \new_[3220]_ , \new_[3221]_ ,
    \new_[3222]_ , \new_[3225]_ , \new_[3229]_ , \new_[3230]_ ,
    \new_[3231]_ , \new_[3234]_ , \new_[3238]_ , \new_[3239]_ ,
    \new_[3240]_ , \new_[3241]_ , \new_[3244]_ , \new_[3248]_ ,
    \new_[3249]_ , \new_[3250]_ , \new_[3253]_ , \new_[3257]_ ,
    \new_[3258]_ , \new_[3259]_ , \new_[3260]_ , \new_[3261]_ ,
    \new_[3262]_ , \new_[3265]_ , \new_[3269]_ , \new_[3270]_ ,
    \new_[3271]_ , \new_[3274]_ , \new_[3278]_ , \new_[3279]_ ,
    \new_[3280]_ , \new_[3281]_ , \new_[3284]_ , \new_[3288]_ ,
    \new_[3289]_ , \new_[3290]_ , \new_[3293]_ , \new_[3297]_ ,
    \new_[3298]_ , \new_[3299]_ , \new_[3300]_ , \new_[3301]_ ,
    \new_[3304]_ , \new_[3308]_ , \new_[3309]_ , \new_[3310]_ ,
    \new_[3313]_ , \new_[3317]_ , \new_[3318]_ , \new_[3319]_ ,
    \new_[3320]_ , \new_[3323]_ , \new_[3327]_ , \new_[3328]_ ,
    \new_[3329]_ , \new_[3332]_ , \new_[3336]_ , \new_[3337]_ ,
    \new_[3338]_ , \new_[3339]_ , \new_[3340]_ , \new_[3341]_ ,
    \new_[3342]_ , \new_[3345]_ , \new_[3349]_ , \new_[3350]_ ,
    \new_[3351]_ , \new_[3354]_ , \new_[3358]_ , \new_[3359]_ ,
    \new_[3360]_ , \new_[3361]_ , \new_[3364]_ , \new_[3368]_ ,
    \new_[3369]_ , \new_[3370]_ , \new_[3373]_ , \new_[3377]_ ,
    \new_[3378]_ , \new_[3379]_ , \new_[3380]_ , \new_[3381]_ ,
    \new_[3384]_ , \new_[3388]_ , \new_[3389]_ , \new_[3390]_ ,
    \new_[3393]_ , \new_[3397]_ , \new_[3398]_ , \new_[3399]_ ,
    \new_[3400]_ , \new_[3403]_ , \new_[3407]_ , \new_[3408]_ ,
    \new_[3409]_ , \new_[3412]_ , \new_[3416]_ , \new_[3417]_ ,
    \new_[3418]_ , \new_[3419]_ , \new_[3420]_ , \new_[3421]_ ,
    \new_[3424]_ , \new_[3428]_ , \new_[3429]_ , \new_[3430]_ ,
    \new_[3433]_ , \new_[3437]_ , \new_[3438]_ , \new_[3439]_ ,
    \new_[3440]_ , \new_[3443]_ , \new_[3447]_ , \new_[3448]_ ,
    \new_[3449]_ , \new_[3452]_ , \new_[3456]_ , \new_[3457]_ ,
    \new_[3458]_ , \new_[3459]_ , \new_[3460]_ , \new_[3463]_ ,
    \new_[3467]_ , \new_[3468]_ , \new_[3469]_ , \new_[3472]_ ,
    \new_[3476]_ , \new_[3477]_ , \new_[3478]_ , \new_[3479]_ ,
    \new_[3482]_ , \new_[3486]_ , \new_[3487]_ , \new_[3488]_ ,
    \new_[3491]_ , \new_[3495]_ , \new_[3496]_ , \new_[3497]_ ,
    \new_[3498]_ , \new_[3499]_ , \new_[3500]_ , \new_[3501]_ ,
    \new_[3502]_ , \new_[3505]_ , \new_[3509]_ , \new_[3510]_ ,
    \new_[3511]_ , \new_[3514]_ , \new_[3518]_ , \new_[3519]_ ,
    \new_[3520]_ , \new_[3521]_ , \new_[3524]_ , \new_[3528]_ ,
    \new_[3529]_ , \new_[3530]_ , \new_[3533]_ , \new_[3537]_ ,
    \new_[3538]_ , \new_[3539]_ , \new_[3540]_ , \new_[3541]_ ,
    \new_[3544]_ , \new_[3548]_ , \new_[3549]_ , \new_[3550]_ ,
    \new_[3553]_ , \new_[3557]_ , \new_[3558]_ , \new_[3559]_ ,
    \new_[3560]_ , \new_[3563]_ , \new_[3567]_ , \new_[3568]_ ,
    \new_[3569]_ , \new_[3572]_ , \new_[3576]_ , \new_[3577]_ ,
    \new_[3578]_ , \new_[3579]_ , \new_[3580]_ , \new_[3581]_ ,
    \new_[3584]_ , \new_[3588]_ , \new_[3589]_ , \new_[3590]_ ,
    \new_[3593]_ , \new_[3597]_ , \new_[3598]_ , \new_[3599]_ ,
    \new_[3600]_ , \new_[3603]_ , \new_[3607]_ , \new_[3608]_ ,
    \new_[3609]_ , \new_[3612]_ , \new_[3616]_ , \new_[3617]_ ,
    \new_[3618]_ , \new_[3619]_ , \new_[3620]_ , \new_[3623]_ ,
    \new_[3627]_ , \new_[3628]_ , \new_[3629]_ , \new_[3632]_ ,
    \new_[3636]_ , \new_[3637]_ , \new_[3638]_ , \new_[3639]_ ,
    \new_[3642]_ , \new_[3646]_ , \new_[3647]_ , \new_[3648]_ ,
    \new_[3651]_ , \new_[3655]_ , \new_[3656]_ , \new_[3657]_ ,
    \new_[3658]_ , \new_[3659]_ , \new_[3660]_ , \new_[3661]_ ,
    \new_[3664]_ , \new_[3668]_ , \new_[3669]_ , \new_[3670]_ ,
    \new_[3673]_ , \new_[3677]_ , \new_[3678]_ , \new_[3679]_ ,
    \new_[3680]_ , \new_[3683]_ , \new_[3687]_ , \new_[3688]_ ,
    \new_[3689]_ , \new_[3692]_ , \new_[3696]_ , \new_[3697]_ ,
    \new_[3698]_ , \new_[3699]_ , \new_[3700]_ , \new_[3703]_ ,
    \new_[3707]_ , \new_[3708]_ , \new_[3709]_ , \new_[3712]_ ,
    \new_[3716]_ , \new_[3717]_ , \new_[3718]_ , \new_[3719]_ ,
    \new_[3722]_ , \new_[3726]_ , \new_[3727]_ , \new_[3728]_ ,
    \new_[3731]_ , \new_[3735]_ , \new_[3736]_ , \new_[3737]_ ,
    \new_[3738]_ , \new_[3739]_ , \new_[3740]_ , \new_[3743]_ ,
    \new_[3747]_ , \new_[3748]_ , \new_[3749]_ , \new_[3752]_ ,
    \new_[3756]_ , \new_[3757]_ , \new_[3758]_ , \new_[3759]_ ,
    \new_[3762]_ , \new_[3766]_ , \new_[3767]_ , \new_[3768]_ ,
    \new_[3771]_ , \new_[3775]_ , \new_[3776]_ , \new_[3777]_ ,
    \new_[3778]_ , \new_[3779]_ , \new_[3782]_ , \new_[3786]_ ,
    \new_[3787]_ , \new_[3788]_ , \new_[3791]_ , \new_[3795]_ ,
    \new_[3796]_ , \new_[3797]_ , \new_[3798]_ , \new_[3801]_ ,
    \new_[3805]_ , \new_[3806]_ , \new_[3807]_ , \new_[3810]_ ,
    \new_[3814]_ , \new_[3815]_ , \new_[3816]_ , \new_[3817]_ ,
    \new_[3818]_ , \new_[3819]_ , \new_[3820]_ , \new_[3821]_ ,
    \new_[3822]_ , \new_[3823]_ , \new_[3826]_ , \new_[3829]_ ,
    \new_[3830]_ , \new_[3833]_ , \new_[3837]_ , \new_[3838]_ ,
    \new_[3839]_ , \new_[3840]_ , \new_[3843]_ , \new_[3847]_ ,
    \new_[3848]_ , \new_[3849]_ , \new_[3852]_ , \new_[3856]_ ,
    \new_[3857]_ , \new_[3858]_ , \new_[3859]_ , \new_[3860]_ ,
    \new_[3863]_ , \new_[3867]_ , \new_[3868]_ , \new_[3869]_ ,
    \new_[3872]_ , \new_[3876]_ , \new_[3877]_ , \new_[3878]_ ,
    \new_[3879]_ , \new_[3882]_ , \new_[3886]_ , \new_[3887]_ ,
    \new_[3888]_ , \new_[3891]_ , \new_[3895]_ , \new_[3896]_ ,
    \new_[3897]_ , \new_[3898]_ , \new_[3899]_ , \new_[3900]_ ,
    \new_[3903]_ , \new_[3907]_ , \new_[3908]_ , \new_[3909]_ ,
    \new_[3912]_ , \new_[3916]_ , \new_[3917]_ , \new_[3918]_ ,
    \new_[3919]_ , \new_[3922]_ , \new_[3926]_ , \new_[3927]_ ,
    \new_[3928]_ , \new_[3931]_ , \new_[3935]_ , \new_[3936]_ ,
    \new_[3937]_ , \new_[3938]_ , \new_[3939]_ , \new_[3942]_ ,
    \new_[3946]_ , \new_[3947]_ , \new_[3948]_ , \new_[3951]_ ,
    \new_[3955]_ , \new_[3956]_ , \new_[3957]_ , \new_[3958]_ ,
    \new_[3961]_ , \new_[3965]_ , \new_[3966]_ , \new_[3967]_ ,
    \new_[3970]_ , \new_[3974]_ , \new_[3975]_ , \new_[3976]_ ,
    \new_[3977]_ , \new_[3978]_ , \new_[3979]_ , \new_[3980]_ ,
    \new_[3983]_ , \new_[3987]_ , \new_[3988]_ , \new_[3989]_ ,
    \new_[3992]_ , \new_[3996]_ , \new_[3997]_ , \new_[3998]_ ,
    \new_[3999]_ , \new_[4002]_ , \new_[4006]_ , \new_[4007]_ ,
    \new_[4008]_ , \new_[4011]_ , \new_[4015]_ , \new_[4016]_ ,
    \new_[4017]_ , \new_[4018]_ , \new_[4019]_ , \new_[4022]_ ,
    \new_[4026]_ , \new_[4027]_ , \new_[4028]_ , \new_[4031]_ ,
    \new_[4035]_ , \new_[4036]_ , \new_[4037]_ , \new_[4038]_ ,
    \new_[4041]_ , \new_[4045]_ , \new_[4046]_ , \new_[4047]_ ,
    \new_[4050]_ , \new_[4054]_ , \new_[4055]_ , \new_[4056]_ ,
    \new_[4057]_ , \new_[4058]_ , \new_[4059]_ , \new_[4062]_ ,
    \new_[4066]_ , \new_[4067]_ , \new_[4068]_ , \new_[4071]_ ,
    \new_[4075]_ , \new_[4076]_ , \new_[4077]_ , \new_[4078]_ ,
    \new_[4081]_ , \new_[4085]_ , \new_[4086]_ , \new_[4087]_ ,
    \new_[4090]_ , \new_[4094]_ , \new_[4095]_ , \new_[4096]_ ,
    \new_[4097]_ , \new_[4098]_ , \new_[4101]_ , \new_[4105]_ ,
    \new_[4106]_ , \new_[4107]_ , \new_[4110]_ , \new_[4114]_ ,
    \new_[4115]_ , \new_[4116]_ , \new_[4117]_ , \new_[4120]_ ,
    \new_[4124]_ , \new_[4125]_ , \new_[4126]_ , \new_[4129]_ ,
    \new_[4133]_ , \new_[4134]_ , \new_[4135]_ , \new_[4136]_ ,
    \new_[4137]_ , \new_[4138]_ , \new_[4139]_ , \new_[4140]_ ,
    \new_[4143]_ , \new_[4147]_ , \new_[4148]_ , \new_[4149]_ ,
    \new_[4152]_ , \new_[4156]_ , \new_[4157]_ , \new_[4158]_ ,
    \new_[4159]_ , \new_[4162]_ , \new_[4166]_ , \new_[4167]_ ,
    \new_[4168]_ , \new_[4171]_ , \new_[4175]_ , \new_[4176]_ ,
    \new_[4177]_ , \new_[4178]_ , \new_[4179]_ , \new_[4182]_ ,
    \new_[4186]_ , \new_[4187]_ , \new_[4188]_ , \new_[4191]_ ,
    \new_[4195]_ , \new_[4196]_ , \new_[4197]_ , \new_[4198]_ ,
    \new_[4201]_ , \new_[4205]_ , \new_[4206]_ , \new_[4207]_ ,
    \new_[4210]_ , \new_[4214]_ , \new_[4215]_ , \new_[4216]_ ,
    \new_[4217]_ , \new_[4218]_ , \new_[4219]_ , \new_[4222]_ ,
    \new_[4226]_ , \new_[4227]_ , \new_[4228]_ , \new_[4231]_ ,
    \new_[4235]_ , \new_[4236]_ , \new_[4237]_ , \new_[4238]_ ,
    \new_[4241]_ , \new_[4245]_ , \new_[4246]_ , \new_[4247]_ ,
    \new_[4250]_ , \new_[4254]_ , \new_[4255]_ , \new_[4256]_ ,
    \new_[4257]_ , \new_[4258]_ , \new_[4261]_ , \new_[4265]_ ,
    \new_[4266]_ , \new_[4267]_ , \new_[4270]_ , \new_[4274]_ ,
    \new_[4275]_ , \new_[4276]_ , \new_[4277]_ , \new_[4280]_ ,
    \new_[4284]_ , \new_[4285]_ , \new_[4286]_ , \new_[4289]_ ,
    \new_[4293]_ , \new_[4294]_ , \new_[4295]_ , \new_[4296]_ ,
    \new_[4297]_ , \new_[4298]_ , \new_[4299]_ , \new_[4302]_ ,
    \new_[4306]_ , \new_[4307]_ , \new_[4308]_ , \new_[4311]_ ,
    \new_[4315]_ , \new_[4316]_ , \new_[4317]_ , \new_[4318]_ ,
    \new_[4321]_ , \new_[4325]_ , \new_[4326]_ , \new_[4327]_ ,
    \new_[4330]_ , \new_[4334]_ , \new_[4335]_ , \new_[4336]_ ,
    \new_[4337]_ , \new_[4338]_ , \new_[4341]_ , \new_[4345]_ ,
    \new_[4346]_ , \new_[4347]_ , \new_[4350]_ , \new_[4354]_ ,
    \new_[4355]_ , \new_[4356]_ , \new_[4357]_ , \new_[4360]_ ,
    \new_[4364]_ , \new_[4365]_ , \new_[4366]_ , \new_[4369]_ ,
    \new_[4373]_ , \new_[4374]_ , \new_[4375]_ , \new_[4376]_ ,
    \new_[4377]_ , \new_[4378]_ , \new_[4381]_ , \new_[4385]_ ,
    \new_[4386]_ , \new_[4387]_ , \new_[4390]_ , \new_[4394]_ ,
    \new_[4395]_ , \new_[4396]_ , \new_[4397]_ , \new_[4400]_ ,
    \new_[4404]_ , \new_[4405]_ , \new_[4406]_ , \new_[4409]_ ,
    \new_[4413]_ , \new_[4414]_ , \new_[4415]_ , \new_[4416]_ ,
    \new_[4417]_ , \new_[4420]_ , \new_[4424]_ , \new_[4425]_ ,
    \new_[4426]_ , \new_[4429]_ , \new_[4433]_ , \new_[4434]_ ,
    \new_[4435]_ , \new_[4436]_ , \new_[4439]_ , \new_[4443]_ ,
    \new_[4444]_ , \new_[4445]_ , \new_[4448]_ , \new_[4452]_ ,
    \new_[4453]_ , \new_[4454]_ , \new_[4455]_ , \new_[4456]_ ,
    \new_[4457]_ , \new_[4458]_ , \new_[4459]_ , \new_[4460]_ ,
    \new_[4463]_ , \new_[4466]_ , \new_[4467]_ , \new_[4470]_ ,
    \new_[4474]_ , \new_[4475]_ , \new_[4476]_ , \new_[4477]_ ,
    \new_[4480]_ , \new_[4484]_ , \new_[4485]_ , \new_[4486]_ ,
    \new_[4489]_ , \new_[4493]_ , \new_[4494]_ , \new_[4495]_ ,
    \new_[4496]_ , \new_[4497]_ , \new_[4500]_ , \new_[4504]_ ,
    \new_[4505]_ , \new_[4506]_ , \new_[4509]_ , \new_[4513]_ ,
    \new_[4514]_ , \new_[4515]_ , \new_[4516]_ , \new_[4519]_ ,
    \new_[4523]_ , \new_[4524]_ , \new_[4525]_ , \new_[4528]_ ,
    \new_[4532]_ , \new_[4533]_ , \new_[4534]_ , \new_[4535]_ ,
    \new_[4536]_ , \new_[4537]_ , \new_[4540]_ , \new_[4544]_ ,
    \new_[4545]_ , \new_[4546]_ , \new_[4549]_ , \new_[4553]_ ,
    \new_[4554]_ , \new_[4555]_ , \new_[4556]_ , \new_[4559]_ ,
    \new_[4563]_ , \new_[4564]_ , \new_[4565]_ , \new_[4568]_ ,
    \new_[4572]_ , \new_[4573]_ , \new_[4574]_ , \new_[4575]_ ,
    \new_[4576]_ , \new_[4579]_ , \new_[4583]_ , \new_[4584]_ ,
    \new_[4585]_ , \new_[4588]_ , \new_[4592]_ , \new_[4593]_ ,
    \new_[4594]_ , \new_[4595]_ , \new_[4598]_ , \new_[4602]_ ,
    \new_[4603]_ , \new_[4604]_ , \new_[4607]_ , \new_[4611]_ ,
    \new_[4612]_ , \new_[4613]_ , \new_[4614]_ , \new_[4615]_ ,
    \new_[4616]_ , \new_[4617]_ , \new_[4620]_ , \new_[4624]_ ,
    \new_[4625]_ , \new_[4626]_ , \new_[4629]_ , \new_[4633]_ ,
    \new_[4634]_ , \new_[4635]_ , \new_[4636]_ , \new_[4639]_ ,
    \new_[4643]_ , \new_[4644]_ , \new_[4645]_ , \new_[4648]_ ,
    \new_[4652]_ , \new_[4653]_ , \new_[4654]_ , \new_[4655]_ ,
    \new_[4656]_ , \new_[4659]_ , \new_[4663]_ , \new_[4664]_ ,
    \new_[4665]_ , \new_[4668]_ , \new_[4672]_ , \new_[4673]_ ,
    \new_[4674]_ , \new_[4675]_ , \new_[4678]_ , \new_[4682]_ ,
    \new_[4683]_ , \new_[4684]_ , \new_[4687]_ , \new_[4691]_ ,
    \new_[4692]_ , \new_[4693]_ , \new_[4694]_ , \new_[4695]_ ,
    \new_[4696]_ , \new_[4699]_ , \new_[4703]_ , \new_[4704]_ ,
    \new_[4705]_ , \new_[4708]_ , \new_[4712]_ , \new_[4713]_ ,
    \new_[4714]_ , \new_[4715]_ , \new_[4718]_ , \new_[4722]_ ,
    \new_[4723]_ , \new_[4724]_ , \new_[4727]_ , \new_[4731]_ ,
    \new_[4732]_ , \new_[4733]_ , \new_[4734]_ , \new_[4735]_ ,
    \new_[4738]_ , \new_[4742]_ , \new_[4743]_ , \new_[4744]_ ,
    \new_[4747]_ , \new_[4751]_ , \new_[4752]_ , \new_[4753]_ ,
    \new_[4754]_ , \new_[4757]_ , \new_[4761]_ , \new_[4762]_ ,
    \new_[4763]_ , \new_[4766]_ , \new_[4770]_ , \new_[4771]_ ,
    \new_[4772]_ , \new_[4773]_ , \new_[4774]_ , \new_[4775]_ ,
    \new_[4776]_ , \new_[4777]_ , \new_[4780]_ , \new_[4784]_ ,
    \new_[4785]_ , \new_[4786]_ , \new_[4789]_ , \new_[4793]_ ,
    \new_[4794]_ , \new_[4795]_ , \new_[4796]_ , \new_[4799]_ ,
    \new_[4803]_ , \new_[4804]_ , \new_[4805]_ , \new_[4808]_ ,
    \new_[4812]_ , \new_[4813]_ , \new_[4814]_ , \new_[4815]_ ,
    \new_[4816]_ , \new_[4819]_ , \new_[4823]_ , \new_[4824]_ ,
    \new_[4825]_ , \new_[4828]_ , \new_[4832]_ , \new_[4833]_ ,
    \new_[4834]_ , \new_[4835]_ , \new_[4838]_ , \new_[4842]_ ,
    \new_[4843]_ , \new_[4844]_ , \new_[4847]_ , \new_[4851]_ ,
    \new_[4852]_ , \new_[4853]_ , \new_[4854]_ , \new_[4855]_ ,
    \new_[4856]_ , \new_[4859]_ , \new_[4863]_ , \new_[4864]_ ,
    \new_[4865]_ , \new_[4868]_ , \new_[4872]_ , \new_[4873]_ ,
    \new_[4874]_ , \new_[4875]_ , \new_[4878]_ , \new_[4882]_ ,
    \new_[4883]_ , \new_[4884]_ , \new_[4887]_ , \new_[4891]_ ,
    \new_[4892]_ , \new_[4893]_ , \new_[4894]_ , \new_[4895]_ ,
    \new_[4898]_ , \new_[4902]_ , \new_[4903]_ , \new_[4904]_ ,
    \new_[4907]_ , \new_[4911]_ , \new_[4912]_ , \new_[4913]_ ,
    \new_[4914]_ , \new_[4917]_ , \new_[4921]_ , \new_[4922]_ ,
    \new_[4923]_ , \new_[4926]_ , \new_[4930]_ , \new_[4931]_ ,
    \new_[4932]_ , \new_[4933]_ , \new_[4934]_ , \new_[4935]_ ,
    \new_[4936]_ , \new_[4939]_ , \new_[4943]_ , \new_[4944]_ ,
    \new_[4945]_ , \new_[4948]_ , \new_[4952]_ , \new_[4953]_ ,
    \new_[4954]_ , \new_[4955]_ , \new_[4958]_ , \new_[4962]_ ,
    \new_[4963]_ , \new_[4964]_ , \new_[4967]_ , \new_[4971]_ ,
    \new_[4972]_ , \new_[4973]_ , \new_[4974]_ , \new_[4975]_ ,
    \new_[4978]_ , \new_[4982]_ , \new_[4983]_ , \new_[4984]_ ,
    \new_[4987]_ , \new_[4991]_ , \new_[4992]_ , \new_[4993]_ ,
    \new_[4994]_ , \new_[4997]_ , \new_[5001]_ , \new_[5002]_ ,
    \new_[5003]_ , \new_[5006]_ , \new_[5010]_ , \new_[5011]_ ,
    \new_[5012]_ , \new_[5013]_ , \new_[5014]_ , \new_[5015]_ ,
    \new_[5018]_ , \new_[5022]_ , \new_[5023]_ , \new_[5024]_ ,
    \new_[5027]_ , \new_[5031]_ , \new_[5032]_ , \new_[5033]_ ,
    \new_[5034]_ , \new_[5037]_ , \new_[5041]_ , \new_[5042]_ ,
    \new_[5043]_ , \new_[5046]_ , \new_[5050]_ , \new_[5051]_ ,
    \new_[5052]_ , \new_[5053]_ , \new_[5054]_ , \new_[5057]_ ,
    \new_[5061]_ , \new_[5062]_ , \new_[5063]_ , \new_[5066]_ ,
    \new_[5070]_ , \new_[5071]_ , \new_[5072]_ , \new_[5073]_ ,
    \new_[5076]_ , \new_[5080]_ , \new_[5081]_ , \new_[5082]_ ,
    \new_[5085]_ , \new_[5089]_ , \new_[5090]_ , \new_[5091]_ ,
    \new_[5092]_ , \new_[5093]_ , \new_[5094]_ , \new_[5095]_ ,
    \new_[5096]_ , \new_[5097]_ , \new_[5098]_ , \new_[5099]_ ,
    \new_[5102]_ , \new_[5105]_ , \new_[5106]_ , \new_[5109]_ ,
    \new_[5113]_ , \new_[5114]_ , \new_[5115]_ , \new_[5116]_ ,
    \new_[5119]_ , \new_[5123]_ , \new_[5124]_ , \new_[5125]_ ,
    \new_[5128]_ , \new_[5132]_ , \new_[5133]_ , \new_[5134]_ ,
    \new_[5135]_ , \new_[5136]_ , \new_[5139]_ , \new_[5143]_ ,
    \new_[5144]_ , \new_[5145]_ , \new_[5148]_ , \new_[5152]_ ,
    \new_[5153]_ , \new_[5154]_ , \new_[5155]_ , \new_[5158]_ ,
    \new_[5162]_ , \new_[5163]_ , \new_[5164]_ , \new_[5167]_ ,
    \new_[5171]_ , \new_[5172]_ , \new_[5173]_ , \new_[5174]_ ,
    \new_[5175]_ , \new_[5176]_ , \new_[5179]_ , \new_[5183]_ ,
    \new_[5184]_ , \new_[5185]_ , \new_[5188]_ , \new_[5192]_ ,
    \new_[5193]_ , \new_[5194]_ , \new_[5195]_ , \new_[5198]_ ,
    \new_[5202]_ , \new_[5203]_ , \new_[5204]_ , \new_[5207]_ ,
    \new_[5211]_ , \new_[5212]_ , \new_[5213]_ , \new_[5214]_ ,
    \new_[5215]_ , \new_[5218]_ , \new_[5222]_ , \new_[5223]_ ,
    \new_[5224]_ , \new_[5227]_ , \new_[5231]_ , \new_[5232]_ ,
    \new_[5233]_ , \new_[5234]_ , \new_[5237]_ , \new_[5241]_ ,
    \new_[5242]_ , \new_[5243]_ , \new_[5246]_ , \new_[5250]_ ,
    \new_[5251]_ , \new_[5252]_ , \new_[5253]_ , \new_[5254]_ ,
    \new_[5255]_ , \new_[5256]_ , \new_[5259]_ , \new_[5263]_ ,
    \new_[5264]_ , \new_[5265]_ , \new_[5268]_ , \new_[5272]_ ,
    \new_[5273]_ , \new_[5274]_ , \new_[5275]_ , \new_[5278]_ ,
    \new_[5282]_ , \new_[5283]_ , \new_[5284]_ , \new_[5287]_ ,
    \new_[5291]_ , \new_[5292]_ , \new_[5293]_ , \new_[5294]_ ,
    \new_[5295]_ , \new_[5298]_ , \new_[5302]_ , \new_[5303]_ ,
    \new_[5304]_ , \new_[5307]_ , \new_[5311]_ , \new_[5312]_ ,
    \new_[5313]_ , \new_[5314]_ , \new_[5317]_ , \new_[5321]_ ,
    \new_[5322]_ , \new_[5323]_ , \new_[5326]_ , \new_[5330]_ ,
    \new_[5331]_ , \new_[5332]_ , \new_[5333]_ , \new_[5334]_ ,
    \new_[5335]_ , \new_[5338]_ , \new_[5342]_ , \new_[5343]_ ,
    \new_[5344]_ , \new_[5347]_ , \new_[5351]_ , \new_[5352]_ ,
    \new_[5353]_ , \new_[5354]_ , \new_[5357]_ , \new_[5361]_ ,
    \new_[5362]_ , \new_[5363]_ , \new_[5366]_ , \new_[5370]_ ,
    \new_[5371]_ , \new_[5372]_ , \new_[5373]_ , \new_[5374]_ ,
    \new_[5377]_ , \new_[5381]_ , \new_[5382]_ , \new_[5383]_ ,
    \new_[5386]_ , \new_[5390]_ , \new_[5391]_ , \new_[5392]_ ,
    \new_[5393]_ , \new_[5396]_ , \new_[5400]_ , \new_[5401]_ ,
    \new_[5402]_ , \new_[5405]_ , \new_[5409]_ , \new_[5410]_ ,
    \new_[5411]_ , \new_[5412]_ , \new_[5413]_ , \new_[5414]_ ,
    \new_[5415]_ , \new_[5416]_ , \new_[5419]_ , \new_[5422]_ ,
    \new_[5423]_ , \new_[5426]_ , \new_[5430]_ , \new_[5431]_ ,
    \new_[5432]_ , \new_[5433]_ , \new_[5436]_ , \new_[5440]_ ,
    \new_[5441]_ , \new_[5442]_ , \new_[5445]_ , \new_[5449]_ ,
    \new_[5450]_ , \new_[5451]_ , \new_[5452]_ , \new_[5453]_ ,
    \new_[5456]_ , \new_[5460]_ , \new_[5461]_ , \new_[5462]_ ,
    \new_[5465]_ , \new_[5469]_ , \new_[5470]_ , \new_[5471]_ ,
    \new_[5472]_ , \new_[5475]_ , \new_[5479]_ , \new_[5480]_ ,
    \new_[5481]_ , \new_[5484]_ , \new_[5488]_ , \new_[5489]_ ,
    \new_[5490]_ , \new_[5491]_ , \new_[5492]_ , \new_[5493]_ ,
    \new_[5496]_ , \new_[5500]_ , \new_[5501]_ , \new_[5502]_ ,
    \new_[5505]_ , \new_[5509]_ , \new_[5510]_ , \new_[5511]_ ,
    \new_[5512]_ , \new_[5515]_ , \new_[5519]_ , \new_[5520]_ ,
    \new_[5521]_ , \new_[5524]_ , \new_[5528]_ , \new_[5529]_ ,
    \new_[5530]_ , \new_[5531]_ , \new_[5532]_ , \new_[5535]_ ,
    \new_[5539]_ , \new_[5540]_ , \new_[5541]_ , \new_[5544]_ ,
    \new_[5548]_ , \new_[5549]_ , \new_[5550]_ , \new_[5551]_ ,
    \new_[5554]_ , \new_[5558]_ , \new_[5559]_ , \new_[5560]_ ,
    \new_[5563]_ , \new_[5567]_ , \new_[5568]_ , \new_[5569]_ ,
    \new_[5570]_ , \new_[5571]_ , \new_[5572]_ , \new_[5573]_ ,
    \new_[5576]_ , \new_[5580]_ , \new_[5581]_ , \new_[5582]_ ,
    \new_[5585]_ , \new_[5589]_ , \new_[5590]_ , \new_[5591]_ ,
    \new_[5592]_ , \new_[5595]_ , \new_[5599]_ , \new_[5600]_ ,
    \new_[5601]_ , \new_[5604]_ , \new_[5608]_ , \new_[5609]_ ,
    \new_[5610]_ , \new_[5611]_ , \new_[5612]_ , \new_[5615]_ ,
    \new_[5619]_ , \new_[5620]_ , \new_[5621]_ , \new_[5624]_ ,
    \new_[5628]_ , \new_[5629]_ , \new_[5630]_ , \new_[5631]_ ,
    \new_[5634]_ , \new_[5638]_ , \new_[5639]_ , \new_[5640]_ ,
    \new_[5643]_ , \new_[5647]_ , \new_[5648]_ , \new_[5649]_ ,
    \new_[5650]_ , \new_[5651]_ , \new_[5652]_ , \new_[5655]_ ,
    \new_[5659]_ , \new_[5660]_ , \new_[5661]_ , \new_[5664]_ ,
    \new_[5668]_ , \new_[5669]_ , \new_[5670]_ , \new_[5671]_ ,
    \new_[5674]_ , \new_[5678]_ , \new_[5679]_ , \new_[5680]_ ,
    \new_[5683]_ , \new_[5687]_ , \new_[5688]_ , \new_[5689]_ ,
    \new_[5690]_ , \new_[5691]_ , \new_[5694]_ , \new_[5698]_ ,
    \new_[5699]_ , \new_[5700]_ , \new_[5703]_ , \new_[5707]_ ,
    \new_[5708]_ , \new_[5709]_ , \new_[5710]_ , \new_[5713]_ ,
    \new_[5717]_ , \new_[5718]_ , \new_[5719]_ , \new_[5722]_ ,
    \new_[5726]_ , \new_[5727]_ , \new_[5728]_ , \new_[5729]_ ,
    \new_[5730]_ , \new_[5731]_ , \new_[5732]_ , \new_[5733]_ ,
    \new_[5734]_ , \new_[5737]_ , \new_[5740]_ , \new_[5741]_ ,
    \new_[5744]_ , \new_[5748]_ , \new_[5749]_ , \new_[5750]_ ,
    \new_[5751]_ , \new_[5754]_ , \new_[5758]_ , \new_[5759]_ ,
    \new_[5760]_ , \new_[5763]_ , \new_[5767]_ , \new_[5768]_ ,
    \new_[5769]_ , \new_[5770]_ , \new_[5771]_ , \new_[5774]_ ,
    \new_[5778]_ , \new_[5779]_ , \new_[5780]_ , \new_[5783]_ ,
    \new_[5787]_ , \new_[5788]_ , \new_[5789]_ , \new_[5790]_ ,
    \new_[5793]_ , \new_[5797]_ , \new_[5798]_ , \new_[5799]_ ,
    \new_[5802]_ , \new_[5806]_ , \new_[5807]_ , \new_[5808]_ ,
    \new_[5809]_ , \new_[5810]_ , \new_[5811]_ , \new_[5814]_ ,
    \new_[5818]_ , \new_[5819]_ , \new_[5820]_ , \new_[5823]_ ,
    \new_[5827]_ , \new_[5828]_ , \new_[5829]_ , \new_[5830]_ ,
    \new_[5833]_ , \new_[5837]_ , \new_[5838]_ , \new_[5839]_ ,
    \new_[5842]_ , \new_[5846]_ , \new_[5847]_ , \new_[5848]_ ,
    \new_[5849]_ , \new_[5850]_ , \new_[5853]_ , \new_[5857]_ ,
    \new_[5858]_ , \new_[5859]_ , \new_[5862]_ , \new_[5866]_ ,
    \new_[5867]_ , \new_[5868]_ , \new_[5869]_ , \new_[5872]_ ,
    \new_[5876]_ , \new_[5877]_ , \new_[5878]_ , \new_[5881]_ ,
    \new_[5885]_ , \new_[5886]_ , \new_[5887]_ , \new_[5888]_ ,
    \new_[5889]_ , \new_[5890]_ , \new_[5891]_ , \new_[5894]_ ,
    \new_[5898]_ , \new_[5899]_ , \new_[5900]_ , \new_[5903]_ ,
    \new_[5907]_ , \new_[5908]_ , \new_[5909]_ , \new_[5910]_ ,
    \new_[5913]_ , \new_[5917]_ , \new_[5918]_ , \new_[5919]_ ,
    \new_[5922]_ , \new_[5926]_ , \new_[5927]_ , \new_[5928]_ ,
    \new_[5929]_ , \new_[5930]_ , \new_[5933]_ , \new_[5937]_ ,
    \new_[5938]_ , \new_[5939]_ , \new_[5942]_ , \new_[5946]_ ,
    \new_[5947]_ , \new_[5948]_ , \new_[5949]_ , \new_[5952]_ ,
    \new_[5956]_ , \new_[5957]_ , \new_[5958]_ , \new_[5961]_ ,
    \new_[5965]_ , \new_[5966]_ , \new_[5967]_ , \new_[5968]_ ,
    \new_[5969]_ , \new_[5970]_ , \new_[5973]_ , \new_[5977]_ ,
    \new_[5978]_ , \new_[5979]_ , \new_[5982]_ , \new_[5986]_ ,
    \new_[5987]_ , \new_[5988]_ , \new_[5989]_ , \new_[5992]_ ,
    \new_[5996]_ , \new_[5997]_ , \new_[5998]_ , \new_[6001]_ ,
    \new_[6005]_ , \new_[6006]_ , \new_[6007]_ , \new_[6008]_ ,
    \new_[6009]_ , \new_[6012]_ , \new_[6016]_ , \new_[6017]_ ,
    \new_[6018]_ , \new_[6021]_ , \new_[6025]_ , \new_[6026]_ ,
    \new_[6027]_ , \new_[6028]_ , \new_[6031]_ , \new_[6035]_ ,
    \new_[6036]_ , \new_[6037]_ , \new_[6040]_ , \new_[6044]_ ,
    \new_[6045]_ , \new_[6046]_ , \new_[6047]_ , \new_[6048]_ ,
    \new_[6049]_ , \new_[6050]_ , \new_[6051]_ , \new_[6054]_ ,
    \new_[6058]_ , \new_[6059]_ , \new_[6060]_ , \new_[6063]_ ,
    \new_[6067]_ , \new_[6068]_ , \new_[6069]_ , \new_[6070]_ ,
    \new_[6073]_ , \new_[6077]_ , \new_[6078]_ , \new_[6079]_ ,
    \new_[6082]_ , \new_[6086]_ , \new_[6087]_ , \new_[6088]_ ,
    \new_[6089]_ , \new_[6090]_ , \new_[6093]_ , \new_[6097]_ ,
    \new_[6098]_ , \new_[6099]_ , \new_[6102]_ , \new_[6106]_ ,
    \new_[6107]_ , \new_[6108]_ , \new_[6109]_ , \new_[6112]_ ,
    \new_[6116]_ , \new_[6117]_ , \new_[6118]_ , \new_[6121]_ ,
    \new_[6125]_ , \new_[6126]_ , \new_[6127]_ , \new_[6128]_ ,
    \new_[6129]_ , \new_[6130]_ , \new_[6133]_ , \new_[6137]_ ,
    \new_[6138]_ , \new_[6139]_ , \new_[6142]_ , \new_[6146]_ ,
    \new_[6147]_ , \new_[6148]_ , \new_[6149]_ , \new_[6152]_ ,
    \new_[6156]_ , \new_[6157]_ , \new_[6158]_ , \new_[6161]_ ,
    \new_[6165]_ , \new_[6166]_ , \new_[6167]_ , \new_[6168]_ ,
    \new_[6169]_ , \new_[6172]_ , \new_[6176]_ , \new_[6177]_ ,
    \new_[6178]_ , \new_[6181]_ , \new_[6185]_ , \new_[6186]_ ,
    \new_[6187]_ , \new_[6188]_ , \new_[6191]_ , \new_[6195]_ ,
    \new_[6196]_ , \new_[6197]_ , \new_[6200]_ , \new_[6204]_ ,
    \new_[6205]_ , \new_[6206]_ , \new_[6207]_ , \new_[6208]_ ,
    \new_[6209]_ , \new_[6210]_ , \new_[6213]_ , \new_[6217]_ ,
    \new_[6218]_ , \new_[6219]_ , \new_[6222]_ , \new_[6226]_ ,
    \new_[6227]_ , \new_[6228]_ , \new_[6229]_ , \new_[6232]_ ,
    \new_[6236]_ , \new_[6237]_ , \new_[6238]_ , \new_[6241]_ ,
    \new_[6245]_ , \new_[6246]_ , \new_[6247]_ , \new_[6248]_ ,
    \new_[6249]_ , \new_[6252]_ , \new_[6256]_ , \new_[6257]_ ,
    \new_[6258]_ , \new_[6261]_ , \new_[6265]_ , \new_[6266]_ ,
    \new_[6267]_ , \new_[6268]_ , \new_[6271]_ , \new_[6275]_ ,
    \new_[6276]_ , \new_[6277]_ , \new_[6280]_ , \new_[6284]_ ,
    \new_[6285]_ , \new_[6286]_ , \new_[6287]_ , \new_[6288]_ ,
    \new_[6289]_ , \new_[6292]_ , \new_[6296]_ , \new_[6297]_ ,
    \new_[6298]_ , \new_[6301]_ , \new_[6305]_ , \new_[6306]_ ,
    \new_[6307]_ , \new_[6308]_ , \new_[6311]_ , \new_[6315]_ ,
    \new_[6316]_ , \new_[6317]_ , \new_[6320]_ , \new_[6324]_ ,
    \new_[6325]_ , \new_[6326]_ , \new_[6327]_ , \new_[6328]_ ,
    \new_[6331]_ , \new_[6335]_ , \new_[6336]_ , \new_[6337]_ ,
    \new_[6340]_ , \new_[6344]_ , \new_[6345]_ , \new_[6346]_ ,
    \new_[6347]_ , \new_[6350]_ , \new_[6354]_ , \new_[6355]_ ,
    \new_[6356]_ , \new_[6359]_ , \new_[6363]_ , \new_[6364]_ ,
    \new_[6365]_ , \new_[6366]_ , \new_[6367]_ , \new_[6368]_ ,
    \new_[6369]_ , \new_[6370]_ , \new_[6371]_ , \new_[6372]_ ,
    \new_[6375]_ , \new_[6378]_ , \new_[6379]_ , \new_[6382]_ ,
    \new_[6386]_ , \new_[6387]_ , \new_[6388]_ , \new_[6389]_ ,
    \new_[6392]_ , \new_[6396]_ , \new_[6397]_ , \new_[6398]_ ,
    \new_[6401]_ , \new_[6405]_ , \new_[6406]_ , \new_[6407]_ ,
    \new_[6408]_ , \new_[6409]_ , \new_[6412]_ , \new_[6416]_ ,
    \new_[6417]_ , \new_[6418]_ , \new_[6421]_ , \new_[6425]_ ,
    \new_[6426]_ , \new_[6427]_ , \new_[6428]_ , \new_[6431]_ ,
    \new_[6435]_ , \new_[6436]_ , \new_[6437]_ , \new_[6440]_ ,
    \new_[6444]_ , \new_[6445]_ , \new_[6446]_ , \new_[6447]_ ,
    \new_[6448]_ , \new_[6449]_ , \new_[6452]_ , \new_[6456]_ ,
    \new_[6457]_ , \new_[6458]_ , \new_[6461]_ , \new_[6465]_ ,
    \new_[6466]_ , \new_[6467]_ , \new_[6468]_ , \new_[6471]_ ,
    \new_[6475]_ , \new_[6476]_ , \new_[6477]_ , \new_[6480]_ ,
    \new_[6484]_ , \new_[6485]_ , \new_[6486]_ , \new_[6487]_ ,
    \new_[6488]_ , \new_[6491]_ , \new_[6495]_ , \new_[6496]_ ,
    \new_[6497]_ , \new_[6500]_ , \new_[6504]_ , \new_[6505]_ ,
    \new_[6506]_ , \new_[6507]_ , \new_[6510]_ , \new_[6514]_ ,
    \new_[6515]_ , \new_[6516]_ , \new_[6519]_ , \new_[6523]_ ,
    \new_[6524]_ , \new_[6525]_ , \new_[6526]_ , \new_[6527]_ ,
    \new_[6528]_ , \new_[6529]_ , \new_[6532]_ , \new_[6536]_ ,
    \new_[6537]_ , \new_[6538]_ , \new_[6541]_ , \new_[6545]_ ,
    \new_[6546]_ , \new_[6547]_ , \new_[6548]_ , \new_[6551]_ ,
    \new_[6555]_ , \new_[6556]_ , \new_[6557]_ , \new_[6560]_ ,
    \new_[6564]_ , \new_[6565]_ , \new_[6566]_ , \new_[6567]_ ,
    \new_[6568]_ , \new_[6571]_ , \new_[6575]_ , \new_[6576]_ ,
    \new_[6577]_ , \new_[6580]_ , \new_[6584]_ , \new_[6585]_ ,
    \new_[6586]_ , \new_[6587]_ , \new_[6590]_ , \new_[6594]_ ,
    \new_[6595]_ , \new_[6596]_ , \new_[6599]_ , \new_[6603]_ ,
    \new_[6604]_ , \new_[6605]_ , \new_[6606]_ , \new_[6607]_ ,
    \new_[6608]_ , \new_[6611]_ , \new_[6615]_ , \new_[6616]_ ,
    \new_[6617]_ , \new_[6620]_ , \new_[6624]_ , \new_[6625]_ ,
    \new_[6626]_ , \new_[6627]_ , \new_[6630]_ , \new_[6634]_ ,
    \new_[6635]_ , \new_[6636]_ , \new_[6639]_ , \new_[6643]_ ,
    \new_[6644]_ , \new_[6645]_ , \new_[6646]_ , \new_[6647]_ ,
    \new_[6650]_ , \new_[6654]_ , \new_[6655]_ , \new_[6656]_ ,
    \new_[6659]_ , \new_[6663]_ , \new_[6664]_ , \new_[6665]_ ,
    \new_[6666]_ , \new_[6669]_ , \new_[6673]_ , \new_[6674]_ ,
    \new_[6675]_ , \new_[6678]_ , \new_[6682]_ , \new_[6683]_ ,
    \new_[6684]_ , \new_[6685]_ , \new_[6686]_ , \new_[6687]_ ,
    \new_[6688]_ , \new_[6689]_ , \new_[6692]_ , \new_[6696]_ ,
    \new_[6697]_ , \new_[6698]_ , \new_[6701]_ , \new_[6705]_ ,
    \new_[6706]_ , \new_[6707]_ , \new_[6708]_ , \new_[6711]_ ,
    \new_[6715]_ , \new_[6716]_ , \new_[6717]_ , \new_[6720]_ ,
    \new_[6724]_ , \new_[6725]_ , \new_[6726]_ , \new_[6727]_ ,
    \new_[6728]_ , \new_[6731]_ , \new_[6735]_ , \new_[6736]_ ,
    \new_[6737]_ , \new_[6740]_ , \new_[6744]_ , \new_[6745]_ ,
    \new_[6746]_ , \new_[6747]_ , \new_[6750]_ , \new_[6754]_ ,
    \new_[6755]_ , \new_[6756]_ , \new_[6759]_ , \new_[6763]_ ,
    \new_[6764]_ , \new_[6765]_ , \new_[6766]_ , \new_[6767]_ ,
    \new_[6768]_ , \new_[6771]_ , \new_[6775]_ , \new_[6776]_ ,
    \new_[6777]_ , \new_[6780]_ , \new_[6784]_ , \new_[6785]_ ,
    \new_[6786]_ , \new_[6787]_ , \new_[6790]_ , \new_[6794]_ ,
    \new_[6795]_ , \new_[6796]_ , \new_[6799]_ , \new_[6803]_ ,
    \new_[6804]_ , \new_[6805]_ , \new_[6806]_ , \new_[6807]_ ,
    \new_[6810]_ , \new_[6814]_ , \new_[6815]_ , \new_[6816]_ ,
    \new_[6819]_ , \new_[6823]_ , \new_[6824]_ , \new_[6825]_ ,
    \new_[6826]_ , \new_[6829]_ , \new_[6833]_ , \new_[6834]_ ,
    \new_[6835]_ , \new_[6838]_ , \new_[6842]_ , \new_[6843]_ ,
    \new_[6844]_ , \new_[6845]_ , \new_[6846]_ , \new_[6847]_ ,
    \new_[6848]_ , \new_[6851]_ , \new_[6855]_ , \new_[6856]_ ,
    \new_[6857]_ , \new_[6860]_ , \new_[6864]_ , \new_[6865]_ ,
    \new_[6866]_ , \new_[6867]_ , \new_[6870]_ , \new_[6874]_ ,
    \new_[6875]_ , \new_[6876]_ , \new_[6879]_ , \new_[6883]_ ,
    \new_[6884]_ , \new_[6885]_ , \new_[6886]_ , \new_[6887]_ ,
    \new_[6890]_ , \new_[6894]_ , \new_[6895]_ , \new_[6896]_ ,
    \new_[6899]_ , \new_[6903]_ , \new_[6904]_ , \new_[6905]_ ,
    \new_[6906]_ , \new_[6909]_ , \new_[6913]_ , \new_[6914]_ ,
    \new_[6915]_ , \new_[6918]_ , \new_[6922]_ , \new_[6923]_ ,
    \new_[6924]_ , \new_[6925]_ , \new_[6926]_ , \new_[6927]_ ,
    \new_[6930]_ , \new_[6934]_ , \new_[6935]_ , \new_[6936]_ ,
    \new_[6939]_ , \new_[6943]_ , \new_[6944]_ , \new_[6945]_ ,
    \new_[6946]_ , \new_[6949]_ , \new_[6953]_ , \new_[6954]_ ,
    \new_[6955]_ , \new_[6958]_ , \new_[6962]_ , \new_[6963]_ ,
    \new_[6964]_ , \new_[6965]_ , \new_[6966]_ , \new_[6969]_ ,
    \new_[6973]_ , \new_[6974]_ , \new_[6975]_ , \new_[6978]_ ,
    \new_[6982]_ , \new_[6983]_ , \new_[6984]_ , \new_[6985]_ ,
    \new_[6988]_ , \new_[6992]_ , \new_[6993]_ , \new_[6994]_ ,
    \new_[6997]_ , \new_[7001]_ , \new_[7002]_ , \new_[7003]_ ,
    \new_[7004]_ , \new_[7005]_ , \new_[7006]_ , \new_[7007]_ ,
    \new_[7008]_ , \new_[7009]_ , \new_[7012]_ , \new_[7015]_ ,
    \new_[7016]_ , \new_[7019]_ , \new_[7023]_ , \new_[7024]_ ,
    \new_[7025]_ , \new_[7026]_ , \new_[7029]_ , \new_[7033]_ ,
    \new_[7034]_ , \new_[7035]_ , \new_[7038]_ , \new_[7042]_ ,
    \new_[7043]_ , \new_[7044]_ , \new_[7045]_ , \new_[7046]_ ,
    \new_[7049]_ , \new_[7053]_ , \new_[7054]_ , \new_[7055]_ ,
    \new_[7058]_ , \new_[7062]_ , \new_[7063]_ , \new_[7064]_ ,
    \new_[7065]_ , \new_[7068]_ , \new_[7072]_ , \new_[7073]_ ,
    \new_[7074]_ , \new_[7077]_ , \new_[7081]_ , \new_[7082]_ ,
    \new_[7083]_ , \new_[7084]_ , \new_[7085]_ , \new_[7086]_ ,
    \new_[7089]_ , \new_[7093]_ , \new_[7094]_ , \new_[7095]_ ,
    \new_[7098]_ , \new_[7102]_ , \new_[7103]_ , \new_[7104]_ ,
    \new_[7105]_ , \new_[7108]_ , \new_[7112]_ , \new_[7113]_ ,
    \new_[7114]_ , \new_[7117]_ , \new_[7121]_ , \new_[7122]_ ,
    \new_[7123]_ , \new_[7124]_ , \new_[7125]_ , \new_[7128]_ ,
    \new_[7132]_ , \new_[7133]_ , \new_[7134]_ , \new_[7137]_ ,
    \new_[7141]_ , \new_[7142]_ , \new_[7143]_ , \new_[7144]_ ,
    \new_[7147]_ , \new_[7151]_ , \new_[7152]_ , \new_[7153]_ ,
    \new_[7156]_ , \new_[7160]_ , \new_[7161]_ , \new_[7162]_ ,
    \new_[7163]_ , \new_[7164]_ , \new_[7165]_ , \new_[7166]_ ,
    \new_[7169]_ , \new_[7173]_ , \new_[7174]_ , \new_[7175]_ ,
    \new_[7178]_ , \new_[7182]_ , \new_[7183]_ , \new_[7184]_ ,
    \new_[7185]_ , \new_[7188]_ , \new_[7192]_ , \new_[7193]_ ,
    \new_[7194]_ , \new_[7197]_ , \new_[7201]_ , \new_[7202]_ ,
    \new_[7203]_ , \new_[7204]_ , \new_[7205]_ , \new_[7208]_ ,
    \new_[7212]_ , \new_[7213]_ , \new_[7214]_ , \new_[7217]_ ,
    \new_[7221]_ , \new_[7222]_ , \new_[7223]_ , \new_[7224]_ ,
    \new_[7227]_ , \new_[7231]_ , \new_[7232]_ , \new_[7233]_ ,
    \new_[7236]_ , \new_[7240]_ , \new_[7241]_ , \new_[7242]_ ,
    \new_[7243]_ , \new_[7244]_ , \new_[7245]_ , \new_[7248]_ ,
    \new_[7252]_ , \new_[7253]_ , \new_[7254]_ , \new_[7257]_ ,
    \new_[7261]_ , \new_[7262]_ , \new_[7263]_ , \new_[7264]_ ,
    \new_[7267]_ , \new_[7271]_ , \new_[7272]_ , \new_[7273]_ ,
    \new_[7276]_ , \new_[7280]_ , \new_[7281]_ , \new_[7282]_ ,
    \new_[7283]_ , \new_[7284]_ , \new_[7287]_ , \new_[7291]_ ,
    \new_[7292]_ , \new_[7293]_ , \new_[7296]_ , \new_[7300]_ ,
    \new_[7301]_ , \new_[7302]_ , \new_[7303]_ , \new_[7306]_ ,
    \new_[7310]_ , \new_[7311]_ , \new_[7312]_ , \new_[7315]_ ,
    \new_[7319]_ , \new_[7320]_ , \new_[7321]_ , \new_[7322]_ ,
    \new_[7323]_ , \new_[7324]_ , \new_[7325]_ , \new_[7326]_ ,
    \new_[7329]_ , \new_[7333]_ , \new_[7334]_ , \new_[7335]_ ,
    \new_[7338]_ , \new_[7342]_ , \new_[7343]_ , \new_[7344]_ ,
    \new_[7345]_ , \new_[7348]_ , \new_[7352]_ , \new_[7353]_ ,
    \new_[7354]_ , \new_[7357]_ , \new_[7361]_ , \new_[7362]_ ,
    \new_[7363]_ , \new_[7364]_ , \new_[7365]_ , \new_[7368]_ ,
    \new_[7372]_ , \new_[7373]_ , \new_[7374]_ , \new_[7377]_ ,
    \new_[7381]_ , \new_[7382]_ , \new_[7383]_ , \new_[7384]_ ,
    \new_[7387]_ , \new_[7391]_ , \new_[7392]_ , \new_[7393]_ ,
    \new_[7396]_ , \new_[7400]_ , \new_[7401]_ , \new_[7402]_ ,
    \new_[7403]_ , \new_[7404]_ , \new_[7405]_ , \new_[7408]_ ,
    \new_[7412]_ , \new_[7413]_ , \new_[7414]_ , \new_[7417]_ ,
    \new_[7421]_ , \new_[7422]_ , \new_[7423]_ , \new_[7424]_ ,
    \new_[7427]_ , \new_[7431]_ , \new_[7432]_ , \new_[7433]_ ,
    \new_[7436]_ , \new_[7440]_ , \new_[7441]_ , \new_[7442]_ ,
    \new_[7443]_ , \new_[7444]_ , \new_[7447]_ , \new_[7451]_ ,
    \new_[7452]_ , \new_[7453]_ , \new_[7456]_ , \new_[7460]_ ,
    \new_[7461]_ , \new_[7462]_ , \new_[7463]_ , \new_[7466]_ ,
    \new_[7470]_ , \new_[7471]_ , \new_[7472]_ , \new_[7475]_ ,
    \new_[7479]_ , \new_[7480]_ , \new_[7481]_ , \new_[7482]_ ,
    \new_[7483]_ , \new_[7484]_ , \new_[7485]_ , \new_[7488]_ ,
    \new_[7492]_ , \new_[7493]_ , \new_[7494]_ , \new_[7497]_ ,
    \new_[7501]_ , \new_[7502]_ , \new_[7503]_ , \new_[7504]_ ,
    \new_[7507]_ , \new_[7511]_ , \new_[7512]_ , \new_[7513]_ ,
    \new_[7516]_ , \new_[7520]_ , \new_[7521]_ , \new_[7522]_ ,
    \new_[7523]_ , \new_[7524]_ , \new_[7527]_ , \new_[7531]_ ,
    \new_[7532]_ , \new_[7533]_ , \new_[7536]_ , \new_[7540]_ ,
    \new_[7541]_ , \new_[7542]_ , \new_[7543]_ , \new_[7546]_ ,
    \new_[7550]_ , \new_[7551]_ , \new_[7552]_ , \new_[7555]_ ,
    \new_[7559]_ , \new_[7560]_ , \new_[7561]_ , \new_[7562]_ ,
    \new_[7563]_ , \new_[7564]_ , \new_[7567]_ , \new_[7571]_ ,
    \new_[7572]_ , \new_[7573]_ , \new_[7576]_ , \new_[7580]_ ,
    \new_[7581]_ , \new_[7582]_ , \new_[7583]_ , \new_[7586]_ ,
    \new_[7590]_ , \new_[7591]_ , \new_[7592]_ , \new_[7595]_ ,
    \new_[7599]_ , \new_[7600]_ , \new_[7601]_ , \new_[7602]_ ,
    \new_[7603]_ , \new_[7606]_ , \new_[7610]_ , \new_[7611]_ ,
    \new_[7612]_ , \new_[7615]_ , \new_[7619]_ , \new_[7620]_ ,
    \new_[7621]_ , \new_[7622]_ , \new_[7625]_ , \new_[7629]_ ,
    \new_[7630]_ , \new_[7631]_ , \new_[7634]_ , \new_[7638]_ ,
    \new_[7639]_ , \new_[7640]_ , \new_[7641]_ , \new_[7642]_ ,
    \new_[7643]_ , \new_[7644]_ , \new_[7645]_ , \new_[7646]_ ,
    \new_[7647]_ , \new_[7648]_ , \new_[7652]_ , \new_[7653]_ ,
    \new_[7657]_ , \new_[7658]_ , \new_[7662]_ , \new_[7663]_ ,
    \new_[7667]_ , \new_[7668]_ , \new_[7672]_ , \new_[7673]_ ,
    \new_[7677]_ , \new_[7678]_ , \new_[7682]_ , \new_[7683]_ ,
    \new_[7687]_ , \new_[7688]_ , \new_[7692]_ , \new_[7693]_ ,
    \new_[7696]_ , \new_[7699]_ , \new_[7700]_ , \new_[7704]_ ,
    \new_[7705]_ , \new_[7708]_ , \new_[7711]_ , \new_[7712]_ ,
    \new_[7716]_ , \new_[7717]_ , \new_[7720]_ , \new_[7723]_ ,
    \new_[7724]_ , \new_[7728]_ , \new_[7729]_ , \new_[7732]_ ,
    \new_[7735]_ , \new_[7736]_ , \new_[7740]_ , \new_[7741]_ ,
    \new_[7744]_ , \new_[7747]_ , \new_[7748]_ , \new_[7752]_ ,
    \new_[7753]_ , \new_[7756]_ , \new_[7759]_ , \new_[7760]_ ,
    \new_[7764]_ , \new_[7765]_ , \new_[7768]_ , \new_[7771]_ ,
    \new_[7772]_ , \new_[7776]_ , \new_[7777]_ , \new_[7780]_ ,
    \new_[7783]_ , \new_[7784]_ , \new_[7788]_ , \new_[7789]_ ,
    \new_[7792]_ , \new_[7795]_ , \new_[7796]_ , \new_[7800]_ ,
    \new_[7801]_ , \new_[7804]_ , \new_[7807]_ , \new_[7808]_ ,
    \new_[7812]_ , \new_[7813]_ , \new_[7816]_ , \new_[7819]_ ,
    \new_[7820]_ , \new_[7824]_ , \new_[7825]_ , \new_[7828]_ ,
    \new_[7831]_ , \new_[7832]_ , \new_[7836]_ , \new_[7837]_ ,
    \new_[7840]_ , \new_[7843]_ , \new_[7844]_ , \new_[7848]_ ,
    \new_[7849]_ , \new_[7852]_ , \new_[7855]_ , \new_[7856]_ ,
    \new_[7860]_ , \new_[7861]_ , \new_[7864]_ , \new_[7867]_ ,
    \new_[7868]_ , \new_[7872]_ , \new_[7873]_ , \new_[7876]_ ,
    \new_[7879]_ , \new_[7880]_ , \new_[7884]_ , \new_[7885]_ ,
    \new_[7888]_ , \new_[7891]_ , \new_[7892]_ , \new_[7896]_ ,
    \new_[7897]_ , \new_[7900]_ , \new_[7903]_ , \new_[7904]_ ,
    \new_[7908]_ , \new_[7909]_ , \new_[7912]_ , \new_[7915]_ ,
    \new_[7916]_ , \new_[7920]_ , \new_[7921]_ , \new_[7924]_ ,
    \new_[7927]_ , \new_[7928]_ , \new_[7932]_ , \new_[7933]_ ,
    \new_[7936]_ , \new_[7939]_ , \new_[7940]_ , \new_[7944]_ ,
    \new_[7945]_ , \new_[7948]_ , \new_[7951]_ , \new_[7952]_ ,
    \new_[7956]_ , \new_[7957]_ , \new_[7960]_ , \new_[7963]_ ,
    \new_[7964]_ , \new_[7968]_ , \new_[7969]_ , \new_[7972]_ ,
    \new_[7975]_ , \new_[7976]_ , \new_[7980]_ , \new_[7981]_ ,
    \new_[7984]_ , \new_[7987]_ , \new_[7988]_ , \new_[7992]_ ,
    \new_[7993]_ , \new_[7996]_ , \new_[7999]_ , \new_[8000]_ ,
    \new_[8003]_ , \new_[8006]_ , \new_[8007]_ , \new_[8010]_ ,
    \new_[8013]_ , \new_[8014]_ , \new_[8017]_ , \new_[8020]_ ,
    \new_[8021]_ , \new_[8024]_ , \new_[8027]_ , \new_[8028]_ ,
    \new_[8031]_ , \new_[8034]_ , \new_[8035]_ , \new_[8038]_ ,
    \new_[8041]_ , \new_[8042]_ , \new_[8045]_ , \new_[8048]_ ,
    \new_[8049]_ , \new_[8052]_ , \new_[8055]_ , \new_[8056]_ ,
    \new_[8059]_ , \new_[8062]_ , \new_[8063]_ , \new_[8066]_ ,
    \new_[8069]_ , \new_[8070]_ , \new_[8073]_ , \new_[8076]_ ,
    \new_[8077]_ , \new_[8080]_ , \new_[8083]_ , \new_[8084]_ ,
    \new_[8087]_ , \new_[8090]_ , \new_[8091]_ , \new_[8094]_ ,
    \new_[8097]_ , \new_[8098]_ , \new_[8101]_ , \new_[8104]_ ,
    \new_[8105]_ , \new_[8108]_ , \new_[8111]_ , \new_[8112]_ ,
    \new_[8115]_ , \new_[8118]_ , \new_[8119]_ , \new_[8122]_ ,
    \new_[8125]_ , \new_[8126]_ , \new_[8129]_ , \new_[8132]_ ,
    \new_[8133]_ , \new_[8136]_ , \new_[8139]_ , \new_[8140]_ ,
    \new_[8143]_ , \new_[8146]_ , \new_[8147]_ , \new_[8150]_ ,
    \new_[8153]_ , \new_[8154]_ , \new_[8157]_ , \new_[8160]_ ,
    \new_[8161]_ , \new_[8164]_ , \new_[8167]_ , \new_[8168]_ ,
    \new_[8171]_ , \new_[8174]_ , \new_[8175]_ , \new_[8178]_ ,
    \new_[8181]_ , \new_[8182]_ , \new_[8185]_ , \new_[8188]_ ,
    \new_[8189]_ , \new_[8192]_ , \new_[8195]_ , \new_[8196]_ ,
    \new_[8199]_ , \new_[8202]_ , \new_[8203]_ , \new_[8206]_ ,
    \new_[8209]_ , \new_[8210]_ , \new_[8213]_ , \new_[8216]_ ,
    \new_[8217]_ , \new_[8220]_ , \new_[8223]_ , \new_[8224]_ ,
    \new_[8227]_ , \new_[8230]_ , \new_[8231]_ , \new_[8234]_ ,
    \new_[8237]_ , \new_[8238]_ , \new_[8241]_ , \new_[8244]_ ,
    \new_[8245]_ , \new_[8248]_ , \new_[8251]_ , \new_[8252]_ ,
    \new_[8255]_ , \new_[8258]_ , \new_[8259]_ , \new_[8262]_ ,
    \new_[8265]_ , \new_[8266]_ , \new_[8269]_ , \new_[8272]_ ,
    \new_[8273]_ , \new_[8276]_ , \new_[8279]_ , \new_[8280]_ ,
    \new_[8283]_ , \new_[8286]_ , \new_[8287]_ , \new_[8290]_ ,
    \new_[8293]_ , \new_[8294]_ , \new_[8297]_ , \new_[8300]_ ,
    \new_[8301]_ , \new_[8304]_ , \new_[8307]_ , \new_[8308]_ ,
    \new_[8311]_ , \new_[8314]_ , \new_[8315]_ , \new_[8318]_ ,
    \new_[8321]_ , \new_[8322]_ , \new_[8325]_ , \new_[8328]_ ,
    \new_[8329]_ , \new_[8332]_ , \new_[8335]_ , \new_[8336]_ ,
    \new_[8339]_ , \new_[8342]_ , \new_[8343]_ , \new_[8346]_ ,
    \new_[8349]_ , \new_[8350]_ , \new_[8353]_ , \new_[8356]_ ,
    \new_[8357]_ , \new_[8360]_ , \new_[8363]_ , \new_[8364]_ ,
    \new_[8367]_ , \new_[8370]_ , \new_[8371]_ , \new_[8374]_ ,
    \new_[8377]_ , \new_[8378]_ , \new_[8381]_ , \new_[8384]_ ,
    \new_[8385]_ , \new_[8388]_ , \new_[8391]_ , \new_[8392]_ ,
    \new_[8395]_ , \new_[8398]_ , \new_[8399]_ , \new_[8402]_ ,
    \new_[8405]_ , \new_[8406]_ , \new_[8409]_ , \new_[8412]_ ,
    \new_[8413]_ , \new_[8416]_ , \new_[8419]_ , \new_[8420]_ ,
    \new_[8423]_ , \new_[8426]_ , \new_[8427]_ , \new_[8430]_ ,
    \new_[8433]_ , \new_[8434]_ , \new_[8437]_ , \new_[8440]_ ,
    \new_[8441]_ , \new_[8444]_ , \new_[8447]_ , \new_[8448]_ ,
    \new_[8451]_ , \new_[8454]_ , \new_[8455]_ , \new_[8458]_ ,
    \new_[8461]_ , \new_[8462]_ , \new_[8465]_ , \new_[8468]_ ,
    \new_[8469]_ , \new_[8472]_ , \new_[8475]_ , \new_[8476]_ ,
    \new_[8479]_ , \new_[8482]_ , \new_[8483]_ , \new_[8486]_ ,
    \new_[8489]_ , \new_[8490]_ , \new_[8493]_ , \new_[8496]_ ,
    \new_[8497]_ , \new_[8500]_ , \new_[8503]_ , \new_[8504]_ ,
    \new_[8507]_ , \new_[8510]_ , \new_[8511]_ , \new_[8514]_ ,
    \new_[8517]_ , \new_[8518]_ , \new_[8521]_ , \new_[8524]_ ,
    \new_[8525]_ , \new_[8528]_ , \new_[8531]_ , \new_[8532]_ ,
    \new_[8535]_ , \new_[8538]_ , \new_[8539]_ , \new_[8542]_ ,
    \new_[8545]_ , \new_[8546]_ , \new_[8549]_ , \new_[8552]_ ,
    \new_[8553]_ , \new_[8556]_ , \new_[8559]_ , \new_[8560]_ ,
    \new_[8563]_ , \new_[8566]_ , \new_[8567]_ , \new_[8570]_ ,
    \new_[8573]_ , \new_[8574]_ , \new_[8577]_ , \new_[8580]_ ,
    \new_[8581]_ , \new_[8584]_ , \new_[8587]_ , \new_[8588]_ ,
    \new_[8591]_ , \new_[8594]_ , \new_[8595]_ , \new_[8598]_ ,
    \new_[8601]_ , \new_[8602]_ , \new_[8605]_ , \new_[8608]_ ,
    \new_[8609]_ , \new_[8612]_ , \new_[8615]_ , \new_[8616]_ ,
    \new_[8619]_ , \new_[8622]_ , \new_[8623]_ , \new_[8626]_ ,
    \new_[8629]_ , \new_[8630]_ , \new_[8633]_ , \new_[8636]_ ,
    \new_[8637]_ , \new_[8640]_ , \new_[8643]_ , \new_[8644]_ ,
    \new_[8647]_ , \new_[8650]_ , \new_[8651]_ , \new_[8654]_ ,
    \new_[8657]_ , \new_[8658]_ , \new_[8661]_ , \new_[8664]_ ,
    \new_[8665]_ , \new_[8668]_ , \new_[8671]_ , \new_[8672]_ ,
    \new_[8675]_ , \new_[8678]_ , \new_[8679]_ , \new_[8682]_ ,
    \new_[8685]_ , \new_[8686]_ , \new_[8689]_ , \new_[8692]_ ,
    \new_[8693]_ , \new_[8696]_ , \new_[8699]_ , \new_[8700]_ ,
    \new_[8703]_ , \new_[8706]_ , \new_[8707]_ , \new_[8710]_ ,
    \new_[8713]_ , \new_[8714]_ , \new_[8717]_ , \new_[8720]_ ,
    \new_[8721]_ , \new_[8724]_ , \new_[8727]_ , \new_[8728]_ ,
    \new_[8731]_ , \new_[8734]_ , \new_[8735]_ , \new_[8738]_ ,
    \new_[8741]_ , \new_[8742]_ , \new_[8745]_ , \new_[8748]_ ,
    \new_[8749]_ , \new_[8752]_ , \new_[8755]_ , \new_[8756]_ ,
    \new_[8759]_ , \new_[8762]_ , \new_[8763]_ , \new_[8766]_ ,
    \new_[8769]_ , \new_[8770]_ , \new_[8773]_ , \new_[8776]_ ,
    \new_[8777]_ , \new_[8780]_ , \new_[8783]_ , \new_[8784]_ ,
    \new_[8787]_ , \new_[8790]_ , \new_[8791]_ , \new_[8794]_ ,
    \new_[8797]_ , \new_[8798]_ , \new_[8801]_ , \new_[8804]_ ,
    \new_[8805]_ , \new_[8808]_ , \new_[8811]_ , \new_[8812]_ ,
    \new_[8815]_ , \new_[8818]_ , \new_[8819]_ , \new_[8822]_ ,
    \new_[8825]_ , \new_[8826]_ , \new_[8829]_ , \new_[8832]_ ,
    \new_[8833]_ , \new_[8836]_ , \new_[8839]_ , \new_[8840]_ ,
    \new_[8843]_ , \new_[8846]_ , \new_[8847]_ , \new_[8850]_ ,
    \new_[8853]_ , \new_[8854]_ , \new_[8857]_ , \new_[8860]_ ,
    \new_[8861]_ , \new_[8864]_ , \new_[8867]_ , \new_[8868]_ ,
    \new_[8871]_ , \new_[8874]_ , \new_[8875]_ , \new_[8878]_ ,
    \new_[8881]_ , \new_[8882]_ , \new_[8885]_ , \new_[8888]_ ,
    \new_[8889]_ , \new_[8892]_ , \new_[8895]_ , \new_[8896]_ ,
    \new_[8899]_ , \new_[8902]_ , \new_[8903]_ , \new_[8906]_ ,
    \new_[8909]_ , \new_[8910]_ , \new_[8913]_ , \new_[8916]_ ,
    \new_[8917]_ , \new_[8920]_ , \new_[8923]_ , \new_[8924]_ ,
    \new_[8927]_ , \new_[8930]_ , \new_[8931]_ , \new_[8934]_ ,
    \new_[8937]_ , \new_[8938]_ , \new_[8941]_ , \new_[8944]_ ,
    \new_[8945]_ , \new_[8948]_ , \new_[8951]_ , \new_[8952]_ ,
    \new_[8955]_ , \new_[8958]_ , \new_[8959]_ , \new_[8962]_ ,
    \new_[8965]_ , \new_[8966]_ , \new_[8969]_ , \new_[8972]_ ,
    \new_[8973]_ , \new_[8976]_ , \new_[8979]_ , \new_[8980]_ ,
    \new_[8983]_ , \new_[8986]_ , \new_[8987]_ , \new_[8990]_ ,
    \new_[8993]_ , \new_[8994]_ , \new_[8997]_ , \new_[9000]_ ,
    \new_[9001]_ , \new_[9004]_ , \new_[9007]_ , \new_[9008]_ ,
    \new_[9011]_ , \new_[9014]_ , \new_[9015]_ , \new_[9018]_ ,
    \new_[9021]_ , \new_[9022]_ , \new_[9025]_ , \new_[9028]_ ,
    \new_[9029]_ , \new_[9032]_ , \new_[9035]_ , \new_[9036]_ ,
    \new_[9039]_ , \new_[9042]_ , \new_[9043]_ , \new_[9046]_ ,
    \new_[9049]_ , \new_[9050]_ , \new_[9053]_ , \new_[9056]_ ,
    \new_[9057]_ , \new_[9060]_ , \new_[9063]_ , \new_[9064]_ ,
    \new_[9067]_ , \new_[9070]_ , \new_[9071]_ , \new_[9074]_ ,
    \new_[9077]_ , \new_[9078]_ , \new_[9081]_ , \new_[9084]_ ,
    \new_[9085]_ , \new_[9088]_ , \new_[9091]_ , \new_[9092]_ ,
    \new_[9095]_ , \new_[9098]_ , \new_[9099]_ , \new_[9102]_ ,
    \new_[9105]_ , \new_[9106]_ , \new_[9109]_ , \new_[9112]_ ,
    \new_[9113]_ , \new_[9116]_ , \new_[9119]_ , \new_[9120]_ ,
    \new_[9123]_ , \new_[9126]_ , \new_[9127]_ , \new_[9130]_ ,
    \new_[9133]_ , \new_[9134]_ , \new_[9137]_ , \new_[9140]_ ,
    \new_[9141]_ , \new_[9144]_ , \new_[9147]_ , \new_[9148]_ ,
    \new_[9151]_ , \new_[9154]_ , \new_[9155]_ , \new_[9158]_ ,
    \new_[9161]_ , \new_[9162]_ , \new_[9165]_ , \new_[9168]_ ,
    \new_[9169]_ , \new_[9172]_ , \new_[9175]_ , \new_[9176]_ ,
    \new_[9179]_ , \new_[9182]_ , \new_[9183]_ , \new_[9186]_ ,
    \new_[9189]_ , \new_[9190]_ , \new_[9193]_ , \new_[9196]_ ,
    \new_[9197]_ , \new_[9200]_ , \new_[9203]_ , \new_[9204]_ ,
    \new_[9207]_ , \new_[9210]_ , \new_[9211]_ , \new_[9214]_ ,
    \new_[9217]_ , \new_[9218]_ , \new_[9221]_ , \new_[9224]_ ,
    \new_[9225]_ , \new_[9228]_ , \new_[9231]_ , \new_[9232]_ ,
    \new_[9235]_ , \new_[9238]_ , \new_[9239]_ , \new_[9242]_ ,
    \new_[9245]_ , \new_[9246]_ , \new_[9249]_ , \new_[9252]_ ,
    \new_[9253]_ , \new_[9256]_ , \new_[9259]_ , \new_[9260]_ ,
    \new_[9263]_ , \new_[9266]_ , \new_[9267]_ , \new_[9270]_ ,
    \new_[9273]_ , \new_[9274]_ , \new_[9277]_ , \new_[9280]_ ,
    \new_[9281]_ , \new_[9284]_ , \new_[9287]_ , \new_[9288]_ ,
    \new_[9291]_ , \new_[9294]_ , \new_[9295]_ , \new_[9298]_ ,
    \new_[9302]_ , \new_[9303]_ , \new_[9304]_ , \new_[9307]_ ,
    \new_[9310]_ , \new_[9311]_ , \new_[9314]_ , \new_[9318]_ ,
    \new_[9319]_ , \new_[9320]_ , \new_[9323]_ , \new_[9326]_ ,
    \new_[9327]_ , \new_[9330]_ , \new_[9334]_ , \new_[9335]_ ,
    \new_[9336]_ , \new_[9339]_ , \new_[9342]_ , \new_[9343]_ ,
    \new_[9346]_ , \new_[9350]_ , \new_[9351]_ , \new_[9352]_ ,
    \new_[9355]_ , \new_[9358]_ , \new_[9359]_ , \new_[9362]_ ,
    \new_[9366]_ , \new_[9367]_ , \new_[9368]_ , \new_[9371]_ ,
    \new_[9374]_ , \new_[9375]_ , \new_[9378]_ , \new_[9382]_ ,
    \new_[9383]_ , \new_[9384]_ , \new_[9387]_ , \new_[9390]_ ,
    \new_[9391]_ , \new_[9394]_ , \new_[9398]_ , \new_[9399]_ ,
    \new_[9400]_ , \new_[9403]_ , \new_[9406]_ , \new_[9407]_ ,
    \new_[9410]_ , \new_[9414]_ , \new_[9415]_ , \new_[9416]_ ,
    \new_[9419]_ , \new_[9422]_ , \new_[9423]_ , \new_[9426]_ ,
    \new_[9430]_ , \new_[9431]_ , \new_[9432]_ , \new_[9435]_ ,
    \new_[9438]_ , \new_[9439]_ , \new_[9442]_ , \new_[9446]_ ,
    \new_[9447]_ , \new_[9448]_ , \new_[9451]_ , \new_[9454]_ ,
    \new_[9455]_ , \new_[9458]_ , \new_[9462]_ , \new_[9463]_ ,
    \new_[9464]_ , \new_[9467]_ , \new_[9470]_ , \new_[9471]_ ,
    \new_[9474]_ , \new_[9478]_ , \new_[9479]_ , \new_[9480]_ ,
    \new_[9483]_ , \new_[9486]_ , \new_[9487]_ , \new_[9490]_ ,
    \new_[9494]_ , \new_[9495]_ , \new_[9496]_ , \new_[9499]_ ,
    \new_[9502]_ , \new_[9503]_ , \new_[9506]_ , \new_[9510]_ ,
    \new_[9511]_ , \new_[9512]_ , \new_[9515]_ , \new_[9518]_ ,
    \new_[9519]_ , \new_[9522]_ , \new_[9526]_ , \new_[9527]_ ,
    \new_[9528]_ , \new_[9531]_ , \new_[9534]_ , \new_[9535]_ ,
    \new_[9538]_ , \new_[9542]_ , \new_[9543]_ , \new_[9544]_ ,
    \new_[9547]_ , \new_[9550]_ , \new_[9551]_ , \new_[9554]_ ,
    \new_[9558]_ , \new_[9559]_ , \new_[9560]_ , \new_[9563]_ ,
    \new_[9566]_ , \new_[9567]_ , \new_[9570]_ , \new_[9574]_ ,
    \new_[9575]_ , \new_[9576]_ , \new_[9579]_ , \new_[9582]_ ,
    \new_[9583]_ , \new_[9586]_ , \new_[9590]_ , \new_[9591]_ ,
    \new_[9592]_ , \new_[9595]_ , \new_[9598]_ , \new_[9599]_ ,
    \new_[9602]_ , \new_[9606]_ , \new_[9607]_ , \new_[9608]_ ,
    \new_[9611]_ , \new_[9614]_ , \new_[9615]_ , \new_[9618]_ ,
    \new_[9622]_ , \new_[9623]_ , \new_[9624]_ , \new_[9627]_ ,
    \new_[9630]_ , \new_[9631]_ , \new_[9634]_ , \new_[9638]_ ,
    \new_[9639]_ , \new_[9640]_ , \new_[9643]_ , \new_[9646]_ ,
    \new_[9647]_ , \new_[9650]_ , \new_[9654]_ , \new_[9655]_ ,
    \new_[9656]_ , \new_[9659]_ , \new_[9662]_ , \new_[9663]_ ,
    \new_[9666]_ , \new_[9670]_ , \new_[9671]_ , \new_[9672]_ ,
    \new_[9675]_ , \new_[9678]_ , \new_[9679]_ , \new_[9682]_ ,
    \new_[9686]_ , \new_[9687]_ , \new_[9688]_ , \new_[9691]_ ,
    \new_[9694]_ , \new_[9695]_ , \new_[9698]_ , \new_[9702]_ ,
    \new_[9703]_ , \new_[9704]_ , \new_[9707]_ , \new_[9710]_ ,
    \new_[9711]_ , \new_[9714]_ , \new_[9718]_ , \new_[9719]_ ,
    \new_[9720]_ , \new_[9723]_ , \new_[9726]_ , \new_[9727]_ ,
    \new_[9730]_ , \new_[9734]_ , \new_[9735]_ , \new_[9736]_ ,
    \new_[9739]_ , \new_[9742]_ , \new_[9743]_ , \new_[9746]_ ,
    \new_[9750]_ , \new_[9751]_ , \new_[9752]_ , \new_[9755]_ ,
    \new_[9758]_ , \new_[9759]_ , \new_[9762]_ , \new_[9766]_ ,
    \new_[9767]_ , \new_[9768]_ , \new_[9771]_ , \new_[9774]_ ,
    \new_[9775]_ , \new_[9778]_ , \new_[9782]_ , \new_[9783]_ ,
    \new_[9784]_ , \new_[9787]_ , \new_[9790]_ , \new_[9791]_ ,
    \new_[9794]_ , \new_[9798]_ , \new_[9799]_ , \new_[9800]_ ,
    \new_[9803]_ , \new_[9806]_ , \new_[9807]_ , \new_[9810]_ ,
    \new_[9814]_ , \new_[9815]_ , \new_[9816]_ , \new_[9819]_ ,
    \new_[9822]_ , \new_[9823]_ , \new_[9826]_ , \new_[9830]_ ,
    \new_[9831]_ , \new_[9832]_ , \new_[9835]_ , \new_[9838]_ ,
    \new_[9839]_ , \new_[9842]_ , \new_[9846]_ , \new_[9847]_ ,
    \new_[9848]_ , \new_[9851]_ , \new_[9854]_ , \new_[9855]_ ,
    \new_[9858]_ , \new_[9862]_ , \new_[9863]_ , \new_[9864]_ ,
    \new_[9867]_ , \new_[9870]_ , \new_[9871]_ , \new_[9874]_ ,
    \new_[9878]_ , \new_[9879]_ , \new_[9880]_ , \new_[9883]_ ,
    \new_[9886]_ , \new_[9887]_ , \new_[9890]_ , \new_[9894]_ ,
    \new_[9895]_ , \new_[9896]_ , \new_[9899]_ , \new_[9902]_ ,
    \new_[9903]_ , \new_[9906]_ , \new_[9910]_ , \new_[9911]_ ,
    \new_[9912]_ , \new_[9915]_ , \new_[9918]_ , \new_[9919]_ ,
    \new_[9922]_ , \new_[9926]_ , \new_[9927]_ , \new_[9928]_ ,
    \new_[9931]_ , \new_[9934]_ , \new_[9935]_ , \new_[9938]_ ,
    \new_[9942]_ , \new_[9943]_ , \new_[9944]_ , \new_[9947]_ ,
    \new_[9950]_ , \new_[9951]_ , \new_[9954]_ , \new_[9958]_ ,
    \new_[9959]_ , \new_[9960]_ , \new_[9963]_ , \new_[9966]_ ,
    \new_[9967]_ , \new_[9970]_ , \new_[9974]_ , \new_[9975]_ ,
    \new_[9976]_ , \new_[9979]_ , \new_[9982]_ , \new_[9983]_ ,
    \new_[9986]_ , \new_[9990]_ , \new_[9991]_ , \new_[9992]_ ,
    \new_[9995]_ , \new_[9998]_ , \new_[9999]_ , \new_[10002]_ ,
    \new_[10006]_ , \new_[10007]_ , \new_[10008]_ , \new_[10011]_ ,
    \new_[10014]_ , \new_[10015]_ , \new_[10018]_ , \new_[10022]_ ,
    \new_[10023]_ , \new_[10024]_ , \new_[10027]_ , \new_[10030]_ ,
    \new_[10031]_ , \new_[10034]_ , \new_[10038]_ , \new_[10039]_ ,
    \new_[10040]_ , \new_[10043]_ , \new_[10046]_ , \new_[10047]_ ,
    \new_[10050]_ , \new_[10054]_ , \new_[10055]_ , \new_[10056]_ ,
    \new_[10059]_ , \new_[10062]_ , \new_[10063]_ , \new_[10066]_ ,
    \new_[10070]_ , \new_[10071]_ , \new_[10072]_ , \new_[10075]_ ,
    \new_[10078]_ , \new_[10079]_ , \new_[10082]_ , \new_[10086]_ ,
    \new_[10087]_ , \new_[10088]_ , \new_[10091]_ , \new_[10094]_ ,
    \new_[10095]_ , \new_[10098]_ , \new_[10102]_ , \new_[10103]_ ,
    \new_[10104]_ , \new_[10107]_ , \new_[10110]_ , \new_[10111]_ ,
    \new_[10114]_ , \new_[10118]_ , \new_[10119]_ , \new_[10120]_ ,
    \new_[10123]_ , \new_[10126]_ , \new_[10127]_ , \new_[10130]_ ,
    \new_[10134]_ , \new_[10135]_ , \new_[10136]_ , \new_[10139]_ ,
    \new_[10142]_ , \new_[10143]_ , \new_[10146]_ , \new_[10150]_ ,
    \new_[10151]_ , \new_[10152]_ , \new_[10155]_ , \new_[10158]_ ,
    \new_[10159]_ , \new_[10162]_ , \new_[10166]_ , \new_[10167]_ ,
    \new_[10168]_ , \new_[10171]_ , \new_[10174]_ , \new_[10175]_ ,
    \new_[10178]_ , \new_[10182]_ , \new_[10183]_ , \new_[10184]_ ,
    \new_[10187]_ , \new_[10190]_ , \new_[10191]_ , \new_[10194]_ ,
    \new_[10198]_ , \new_[10199]_ , \new_[10200]_ , \new_[10203]_ ,
    \new_[10206]_ , \new_[10207]_ , \new_[10210]_ , \new_[10214]_ ,
    \new_[10215]_ , \new_[10216]_ , \new_[10219]_ , \new_[10222]_ ,
    \new_[10223]_ , \new_[10226]_ , \new_[10230]_ , \new_[10231]_ ,
    \new_[10232]_ , \new_[10235]_ , \new_[10238]_ , \new_[10239]_ ,
    \new_[10242]_ , \new_[10246]_ , \new_[10247]_ , \new_[10248]_ ,
    \new_[10251]_ , \new_[10254]_ , \new_[10255]_ , \new_[10258]_ ,
    \new_[10262]_ , \new_[10263]_ , \new_[10264]_ , \new_[10267]_ ,
    \new_[10270]_ , \new_[10271]_ , \new_[10274]_ , \new_[10278]_ ,
    \new_[10279]_ , \new_[10280]_ , \new_[10283]_ , \new_[10286]_ ,
    \new_[10287]_ , \new_[10290]_ , \new_[10294]_ , \new_[10295]_ ,
    \new_[10296]_ , \new_[10299]_ , \new_[10302]_ , \new_[10303]_ ,
    \new_[10306]_ , \new_[10310]_ , \new_[10311]_ , \new_[10312]_ ,
    \new_[10315]_ , \new_[10318]_ , \new_[10319]_ , \new_[10322]_ ,
    \new_[10326]_ , \new_[10327]_ , \new_[10328]_ , \new_[10331]_ ,
    \new_[10334]_ , \new_[10335]_ , \new_[10338]_ , \new_[10342]_ ,
    \new_[10343]_ , \new_[10344]_ , \new_[10347]_ , \new_[10350]_ ,
    \new_[10351]_ , \new_[10354]_ , \new_[10358]_ , \new_[10359]_ ,
    \new_[10360]_ , \new_[10363]_ , \new_[10366]_ , \new_[10367]_ ,
    \new_[10370]_ , \new_[10374]_ , \new_[10375]_ , \new_[10376]_ ,
    \new_[10379]_ , \new_[10382]_ , \new_[10383]_ , \new_[10386]_ ,
    \new_[10390]_ , \new_[10391]_ , \new_[10392]_ , \new_[10395]_ ,
    \new_[10398]_ , \new_[10399]_ , \new_[10402]_ , \new_[10406]_ ,
    \new_[10407]_ , \new_[10408]_ , \new_[10411]_ , \new_[10414]_ ,
    \new_[10415]_ , \new_[10418]_ , \new_[10422]_ , \new_[10423]_ ,
    \new_[10424]_ , \new_[10427]_ , \new_[10430]_ , \new_[10431]_ ,
    \new_[10434]_ , \new_[10438]_ , \new_[10439]_ , \new_[10440]_ ,
    \new_[10443]_ , \new_[10446]_ , \new_[10447]_ , \new_[10450]_ ,
    \new_[10454]_ , \new_[10455]_ , \new_[10456]_ , \new_[10459]_ ,
    \new_[10462]_ , \new_[10463]_ , \new_[10466]_ , \new_[10470]_ ,
    \new_[10471]_ , \new_[10472]_ , \new_[10475]_ , \new_[10478]_ ,
    \new_[10479]_ , \new_[10482]_ , \new_[10486]_ , \new_[10487]_ ,
    \new_[10488]_ , \new_[10491]_ , \new_[10494]_ , \new_[10495]_ ,
    \new_[10498]_ , \new_[10502]_ , \new_[10503]_ , \new_[10504]_ ,
    \new_[10507]_ , \new_[10510]_ , \new_[10511]_ , \new_[10514]_ ,
    \new_[10518]_ , \new_[10519]_ , \new_[10520]_ , \new_[10523]_ ,
    \new_[10526]_ , \new_[10527]_ , \new_[10530]_ , \new_[10534]_ ,
    \new_[10535]_ , \new_[10536]_ , \new_[10539]_ , \new_[10542]_ ,
    \new_[10543]_ , \new_[10546]_ , \new_[10550]_ , \new_[10551]_ ,
    \new_[10552]_ , \new_[10555]_ , \new_[10558]_ , \new_[10559]_ ,
    \new_[10562]_ , \new_[10566]_ , \new_[10567]_ , \new_[10568]_ ,
    \new_[10571]_ , \new_[10574]_ , \new_[10575]_ , \new_[10578]_ ,
    \new_[10582]_ , \new_[10583]_ , \new_[10584]_ , \new_[10587]_ ,
    \new_[10590]_ , \new_[10591]_ , \new_[10594]_ , \new_[10598]_ ,
    \new_[10599]_ , \new_[10600]_ , \new_[10603]_ , \new_[10606]_ ,
    \new_[10607]_ , \new_[10610]_ , \new_[10614]_ , \new_[10615]_ ,
    \new_[10616]_ , \new_[10619]_ , \new_[10622]_ , \new_[10623]_ ,
    \new_[10626]_ , \new_[10630]_ , \new_[10631]_ , \new_[10632]_ ,
    \new_[10635]_ , \new_[10638]_ , \new_[10639]_ , \new_[10642]_ ,
    \new_[10646]_ , \new_[10647]_ , \new_[10648]_ , \new_[10651]_ ,
    \new_[10654]_ , \new_[10655]_ , \new_[10658]_ , \new_[10662]_ ,
    \new_[10663]_ , \new_[10664]_ , \new_[10667]_ , \new_[10670]_ ,
    \new_[10671]_ , \new_[10674]_ , \new_[10678]_ , \new_[10679]_ ,
    \new_[10680]_ , \new_[10683]_ , \new_[10686]_ , \new_[10687]_ ,
    \new_[10690]_ , \new_[10694]_ , \new_[10695]_ , \new_[10696]_ ,
    \new_[10699]_ , \new_[10702]_ , \new_[10703]_ , \new_[10706]_ ,
    \new_[10710]_ , \new_[10711]_ , \new_[10712]_ , \new_[10715]_ ,
    \new_[10718]_ , \new_[10719]_ , \new_[10722]_ , \new_[10726]_ ,
    \new_[10727]_ , \new_[10728]_ , \new_[10731]_ , \new_[10734]_ ,
    \new_[10735]_ , \new_[10738]_ , \new_[10742]_ , \new_[10743]_ ,
    \new_[10744]_ , \new_[10747]_ , \new_[10750]_ , \new_[10751]_ ,
    \new_[10754]_ , \new_[10758]_ , \new_[10759]_ , \new_[10760]_ ,
    \new_[10763]_ , \new_[10766]_ , \new_[10767]_ , \new_[10770]_ ,
    \new_[10774]_ , \new_[10775]_ , \new_[10776]_ , \new_[10779]_ ,
    \new_[10782]_ , \new_[10783]_ , \new_[10786]_ , \new_[10790]_ ,
    \new_[10791]_ , \new_[10792]_ , \new_[10795]_ , \new_[10798]_ ,
    \new_[10799]_ , \new_[10802]_ , \new_[10806]_ , \new_[10807]_ ,
    \new_[10808]_ , \new_[10811]_ , \new_[10814]_ , \new_[10815]_ ,
    \new_[10818]_ , \new_[10822]_ , \new_[10823]_ , \new_[10824]_ ,
    \new_[10827]_ , \new_[10830]_ , \new_[10831]_ , \new_[10834]_ ,
    \new_[10838]_ , \new_[10839]_ , \new_[10840]_ , \new_[10843]_ ,
    \new_[10846]_ , \new_[10847]_ , \new_[10850]_ , \new_[10854]_ ,
    \new_[10855]_ , \new_[10856]_ , \new_[10859]_ , \new_[10862]_ ,
    \new_[10863]_ , \new_[10866]_ , \new_[10870]_ , \new_[10871]_ ,
    \new_[10872]_ , \new_[10875]_ , \new_[10878]_ , \new_[10879]_ ,
    \new_[10882]_ , \new_[10886]_ , \new_[10887]_ , \new_[10888]_ ,
    \new_[10891]_ , \new_[10894]_ , \new_[10895]_ , \new_[10898]_ ,
    \new_[10902]_ , \new_[10903]_ , \new_[10904]_ , \new_[10907]_ ,
    \new_[10910]_ , \new_[10911]_ , \new_[10914]_ , \new_[10918]_ ,
    \new_[10919]_ , \new_[10920]_ , \new_[10923]_ , \new_[10926]_ ,
    \new_[10927]_ , \new_[10930]_ , \new_[10934]_ , \new_[10935]_ ,
    \new_[10936]_ , \new_[10939]_ , \new_[10942]_ , \new_[10943]_ ,
    \new_[10946]_ , \new_[10950]_ , \new_[10951]_ , \new_[10952]_ ,
    \new_[10955]_ , \new_[10958]_ , \new_[10959]_ , \new_[10962]_ ,
    \new_[10966]_ , \new_[10967]_ , \new_[10968]_ , \new_[10971]_ ,
    \new_[10974]_ , \new_[10975]_ , \new_[10978]_ , \new_[10982]_ ,
    \new_[10983]_ , \new_[10984]_ , \new_[10987]_ , \new_[10990]_ ,
    \new_[10991]_ , \new_[10994]_ , \new_[10998]_ , \new_[10999]_ ,
    \new_[11000]_ , \new_[11003]_ , \new_[11006]_ , \new_[11007]_ ,
    \new_[11010]_ , \new_[11014]_ , \new_[11015]_ , \new_[11016]_ ,
    \new_[11019]_ , \new_[11022]_ , \new_[11023]_ , \new_[11026]_ ,
    \new_[11030]_ , \new_[11031]_ , \new_[11032]_ , \new_[11035]_ ,
    \new_[11038]_ , \new_[11039]_ , \new_[11042]_ , \new_[11046]_ ,
    \new_[11047]_ , \new_[11048]_ , \new_[11051]_ , \new_[11054]_ ,
    \new_[11055]_ , \new_[11058]_ , \new_[11062]_ , \new_[11063]_ ,
    \new_[11064]_ , \new_[11067]_ , \new_[11070]_ , \new_[11071]_ ,
    \new_[11074]_ , \new_[11078]_ , \new_[11079]_ , \new_[11080]_ ,
    \new_[11083]_ , \new_[11086]_ , \new_[11087]_ , \new_[11090]_ ,
    \new_[11094]_ , \new_[11095]_ , \new_[11096]_ , \new_[11099]_ ,
    \new_[11102]_ , \new_[11103]_ , \new_[11106]_ , \new_[11110]_ ,
    \new_[11111]_ , \new_[11112]_ , \new_[11115]_ , \new_[11118]_ ,
    \new_[11119]_ , \new_[11122]_ , \new_[11126]_ , \new_[11127]_ ,
    \new_[11128]_ , \new_[11131]_ , \new_[11134]_ , \new_[11135]_ ,
    \new_[11138]_ , \new_[11142]_ , \new_[11143]_ , \new_[11144]_ ,
    \new_[11147]_ , \new_[11150]_ , \new_[11151]_ , \new_[11154]_ ,
    \new_[11158]_ , \new_[11159]_ , \new_[11160]_ , \new_[11163]_ ,
    \new_[11166]_ , \new_[11167]_ , \new_[11170]_ , \new_[11174]_ ,
    \new_[11175]_ , \new_[11176]_ , \new_[11179]_ , \new_[11182]_ ,
    \new_[11183]_ , \new_[11186]_ , \new_[11190]_ , \new_[11191]_ ,
    \new_[11192]_ , \new_[11195]_ , \new_[11198]_ , \new_[11199]_ ,
    \new_[11202]_ , \new_[11206]_ , \new_[11207]_ , \new_[11208]_ ,
    \new_[11211]_ , \new_[11214]_ , \new_[11215]_ , \new_[11218]_ ,
    \new_[11222]_ , \new_[11223]_ , \new_[11224]_ , \new_[11227]_ ,
    \new_[11230]_ , \new_[11231]_ , \new_[11234]_ , \new_[11238]_ ,
    \new_[11239]_ , \new_[11240]_ , \new_[11243]_ , \new_[11246]_ ,
    \new_[11247]_ , \new_[11250]_ , \new_[11254]_ , \new_[11255]_ ,
    \new_[11256]_ , \new_[11259]_ , \new_[11262]_ , \new_[11263]_ ,
    \new_[11266]_ , \new_[11270]_ , \new_[11271]_ , \new_[11272]_ ,
    \new_[11275]_ , \new_[11278]_ , \new_[11279]_ , \new_[11282]_ ,
    \new_[11286]_ , \new_[11287]_ , \new_[11288]_ , \new_[11291]_ ,
    \new_[11294]_ , \new_[11295]_ , \new_[11298]_ , \new_[11302]_ ,
    \new_[11303]_ , \new_[11304]_ , \new_[11307]_ , \new_[11310]_ ,
    \new_[11311]_ , \new_[11314]_ , \new_[11318]_ , \new_[11319]_ ,
    \new_[11320]_ , \new_[11323]_ , \new_[11326]_ , \new_[11327]_ ,
    \new_[11330]_ , \new_[11334]_ , \new_[11335]_ , \new_[11336]_ ,
    \new_[11339]_ , \new_[11342]_ , \new_[11343]_ , \new_[11346]_ ,
    \new_[11350]_ , \new_[11351]_ , \new_[11352]_ , \new_[11355]_ ,
    \new_[11358]_ , \new_[11359]_ , \new_[11362]_ , \new_[11366]_ ,
    \new_[11367]_ , \new_[11368]_ , \new_[11371]_ , \new_[11374]_ ,
    \new_[11375]_ , \new_[11378]_ , \new_[11382]_ , \new_[11383]_ ,
    \new_[11384]_ , \new_[11387]_ , \new_[11390]_ , \new_[11391]_ ,
    \new_[11394]_ , \new_[11398]_ , \new_[11399]_ , \new_[11400]_ ,
    \new_[11403]_ , \new_[11406]_ , \new_[11407]_ , \new_[11410]_ ,
    \new_[11414]_ , \new_[11415]_ , \new_[11416]_ , \new_[11419]_ ,
    \new_[11422]_ , \new_[11423]_ , \new_[11426]_ , \new_[11430]_ ,
    \new_[11431]_ , \new_[11432]_ , \new_[11435]_ , \new_[11438]_ ,
    \new_[11439]_ , \new_[11442]_ , \new_[11446]_ , \new_[11447]_ ,
    \new_[11448]_ , \new_[11451]_ , \new_[11454]_ , \new_[11455]_ ,
    \new_[11458]_ , \new_[11462]_ , \new_[11463]_ , \new_[11464]_ ,
    \new_[11467]_ , \new_[11470]_ , \new_[11471]_ , \new_[11474]_ ,
    \new_[11478]_ , \new_[11479]_ , \new_[11480]_ , \new_[11483]_ ,
    \new_[11486]_ , \new_[11487]_ , \new_[11490]_ , \new_[11494]_ ,
    \new_[11495]_ , \new_[11496]_ , \new_[11499]_ , \new_[11502]_ ,
    \new_[11503]_ , \new_[11506]_ , \new_[11510]_ , \new_[11511]_ ,
    \new_[11512]_ , \new_[11515]_ , \new_[11518]_ , \new_[11519]_ ,
    \new_[11522]_ , \new_[11526]_ , \new_[11527]_ , \new_[11528]_ ,
    \new_[11531]_ , \new_[11534]_ , \new_[11535]_ , \new_[11538]_ ,
    \new_[11542]_ , \new_[11543]_ , \new_[11544]_ , \new_[11547]_ ,
    \new_[11550]_ , \new_[11551]_ , \new_[11554]_ , \new_[11558]_ ,
    \new_[11559]_ , \new_[11560]_ , \new_[11563]_ , \new_[11566]_ ,
    \new_[11567]_ , \new_[11570]_ , \new_[11574]_ , \new_[11575]_ ,
    \new_[11576]_ , \new_[11579]_ , \new_[11582]_ , \new_[11583]_ ,
    \new_[11586]_ , \new_[11590]_ , \new_[11591]_ , \new_[11592]_ ,
    \new_[11595]_ , \new_[11598]_ , \new_[11599]_ , \new_[11602]_ ,
    \new_[11606]_ , \new_[11607]_ , \new_[11608]_ , \new_[11611]_ ,
    \new_[11614]_ , \new_[11615]_ , \new_[11618]_ , \new_[11622]_ ,
    \new_[11623]_ , \new_[11624]_ , \new_[11627]_ , \new_[11630]_ ,
    \new_[11631]_ , \new_[11634]_ , \new_[11638]_ , \new_[11639]_ ,
    \new_[11640]_ , \new_[11643]_ , \new_[11646]_ , \new_[11647]_ ,
    \new_[11650]_ , \new_[11654]_ , \new_[11655]_ , \new_[11656]_ ,
    \new_[11659]_ , \new_[11662]_ , \new_[11663]_ , \new_[11666]_ ,
    \new_[11670]_ , \new_[11671]_ , \new_[11672]_ , \new_[11675]_ ,
    \new_[11678]_ , \new_[11679]_ , \new_[11682]_ , \new_[11686]_ ,
    \new_[11687]_ , \new_[11688]_ , \new_[11691]_ , \new_[11694]_ ,
    \new_[11695]_ , \new_[11698]_ , \new_[11702]_ , \new_[11703]_ ,
    \new_[11704]_ , \new_[11707]_ , \new_[11710]_ , \new_[11711]_ ,
    \new_[11714]_ , \new_[11718]_ , \new_[11719]_ , \new_[11720]_ ,
    \new_[11723]_ , \new_[11726]_ , \new_[11727]_ , \new_[11730]_ ,
    \new_[11734]_ , \new_[11735]_ , \new_[11736]_ , \new_[11739]_ ,
    \new_[11742]_ , \new_[11743]_ , \new_[11746]_ , \new_[11750]_ ,
    \new_[11751]_ , \new_[11752]_ , \new_[11755]_ , \new_[11758]_ ,
    \new_[11759]_ , \new_[11762]_ , \new_[11766]_ , \new_[11767]_ ,
    \new_[11768]_ , \new_[11771]_ , \new_[11774]_ , \new_[11775]_ ,
    \new_[11778]_ , \new_[11782]_ , \new_[11783]_ , \new_[11784]_ ,
    \new_[11787]_ , \new_[11790]_ , \new_[11791]_ , \new_[11794]_ ,
    \new_[11798]_ , \new_[11799]_ , \new_[11800]_ , \new_[11803]_ ,
    \new_[11806]_ , \new_[11807]_ , \new_[11810]_ , \new_[11814]_ ,
    \new_[11815]_ , \new_[11816]_ , \new_[11819]_ , \new_[11822]_ ,
    \new_[11823]_ , \new_[11826]_ , \new_[11830]_ , \new_[11831]_ ,
    \new_[11832]_ , \new_[11835]_ , \new_[11838]_ , \new_[11839]_ ,
    \new_[11842]_ , \new_[11846]_ , \new_[11847]_ , \new_[11848]_ ,
    \new_[11851]_ , \new_[11854]_ , \new_[11855]_ , \new_[11858]_ ,
    \new_[11862]_ , \new_[11863]_ , \new_[11864]_ , \new_[11867]_ ,
    \new_[11870]_ , \new_[11871]_ , \new_[11874]_ , \new_[11878]_ ,
    \new_[11879]_ , \new_[11880]_ , \new_[11883]_ , \new_[11886]_ ,
    \new_[11887]_ , \new_[11890]_ , \new_[11894]_ , \new_[11895]_ ,
    \new_[11896]_ , \new_[11899]_ , \new_[11902]_ , \new_[11903]_ ,
    \new_[11906]_ , \new_[11910]_ , \new_[11911]_ , \new_[11912]_ ,
    \new_[11915]_ , \new_[11918]_ , \new_[11919]_ , \new_[11922]_ ,
    \new_[11926]_ , \new_[11927]_ , \new_[11928]_ , \new_[11931]_ ,
    \new_[11934]_ , \new_[11935]_ , \new_[11938]_ , \new_[11942]_ ,
    \new_[11943]_ , \new_[11944]_ , \new_[11947]_ , \new_[11950]_ ,
    \new_[11951]_ , \new_[11954]_ , \new_[11958]_ , \new_[11959]_ ,
    \new_[11960]_ , \new_[11963]_ , \new_[11966]_ , \new_[11967]_ ,
    \new_[11970]_ , \new_[11974]_ , \new_[11975]_ , \new_[11976]_ ,
    \new_[11979]_ , \new_[11982]_ , \new_[11983]_ , \new_[11986]_ ,
    \new_[11990]_ , \new_[11991]_ , \new_[11992]_ , \new_[11995]_ ,
    \new_[11998]_ , \new_[11999]_ , \new_[12002]_ , \new_[12006]_ ,
    \new_[12007]_ , \new_[12008]_ , \new_[12011]_ , \new_[12014]_ ,
    \new_[12015]_ , \new_[12018]_ , \new_[12022]_ , \new_[12023]_ ,
    \new_[12024]_ , \new_[12027]_ , \new_[12030]_ , \new_[12031]_ ,
    \new_[12034]_ , \new_[12038]_ , \new_[12039]_ , \new_[12040]_ ,
    \new_[12043]_ , \new_[12046]_ , \new_[12047]_ , \new_[12050]_ ,
    \new_[12054]_ , \new_[12055]_ , \new_[12056]_ , \new_[12059]_ ,
    \new_[12062]_ , \new_[12063]_ , \new_[12066]_ , \new_[12070]_ ,
    \new_[12071]_ , \new_[12072]_ , \new_[12075]_ , \new_[12078]_ ,
    \new_[12079]_ , \new_[12082]_ , \new_[12086]_ , \new_[12087]_ ,
    \new_[12088]_ , \new_[12091]_ , \new_[12094]_ , \new_[12095]_ ,
    \new_[12098]_ , \new_[12102]_ , \new_[12103]_ , \new_[12104]_ ,
    \new_[12107]_ , \new_[12110]_ , \new_[12111]_ , \new_[12114]_ ,
    \new_[12118]_ , \new_[12119]_ , \new_[12120]_ , \new_[12123]_ ,
    \new_[12126]_ , \new_[12127]_ , \new_[12130]_ , \new_[12134]_ ,
    \new_[12135]_ , \new_[12136]_ , \new_[12139]_ , \new_[12142]_ ,
    \new_[12143]_ , \new_[12146]_ , \new_[12150]_ , \new_[12151]_ ,
    \new_[12152]_ , \new_[12155]_ , \new_[12158]_ , \new_[12159]_ ,
    \new_[12162]_ , \new_[12166]_ , \new_[12167]_ , \new_[12168]_ ,
    \new_[12171]_ , \new_[12174]_ , \new_[12175]_ , \new_[12178]_ ,
    \new_[12182]_ , \new_[12183]_ , \new_[12184]_ , \new_[12187]_ ,
    \new_[12190]_ , \new_[12191]_ , \new_[12194]_ , \new_[12198]_ ,
    \new_[12199]_ , \new_[12200]_ , \new_[12203]_ , \new_[12206]_ ,
    \new_[12207]_ , \new_[12210]_ , \new_[12214]_ , \new_[12215]_ ,
    \new_[12216]_ , \new_[12219]_ , \new_[12222]_ , \new_[12223]_ ,
    \new_[12226]_ , \new_[12230]_ , \new_[12231]_ , \new_[12232]_ ,
    \new_[12235]_ , \new_[12238]_ , \new_[12239]_ , \new_[12242]_ ,
    \new_[12246]_ , \new_[12247]_ , \new_[12248]_ , \new_[12251]_ ,
    \new_[12254]_ , \new_[12255]_ , \new_[12258]_ , \new_[12262]_ ,
    \new_[12263]_ , \new_[12264]_ , \new_[12267]_ , \new_[12270]_ ,
    \new_[12271]_ , \new_[12274]_ , \new_[12278]_ , \new_[12279]_ ,
    \new_[12280]_ , \new_[12283]_ , \new_[12286]_ , \new_[12287]_ ,
    \new_[12290]_ , \new_[12294]_ , \new_[12295]_ , \new_[12296]_ ,
    \new_[12299]_ , \new_[12302]_ , \new_[12303]_ , \new_[12306]_ ,
    \new_[12310]_ , \new_[12311]_ , \new_[12312]_ , \new_[12315]_ ,
    \new_[12318]_ , \new_[12319]_ , \new_[12322]_ , \new_[12326]_ ,
    \new_[12327]_ , \new_[12328]_ , \new_[12331]_ , \new_[12334]_ ,
    \new_[12335]_ , \new_[12338]_ , \new_[12342]_ , \new_[12343]_ ,
    \new_[12344]_ , \new_[12347]_ , \new_[12350]_ , \new_[12351]_ ,
    \new_[12354]_ , \new_[12358]_ , \new_[12359]_ , \new_[12360]_ ,
    \new_[12363]_ , \new_[12366]_ , \new_[12367]_ , \new_[12370]_ ,
    \new_[12374]_ , \new_[12375]_ , \new_[12376]_ , \new_[12379]_ ,
    \new_[12382]_ , \new_[12383]_ , \new_[12386]_ , \new_[12390]_ ,
    \new_[12391]_ , \new_[12392]_ , \new_[12395]_ , \new_[12398]_ ,
    \new_[12399]_ , \new_[12402]_ , \new_[12406]_ , \new_[12407]_ ,
    \new_[12408]_ , \new_[12411]_ , \new_[12414]_ , \new_[12415]_ ,
    \new_[12418]_ , \new_[12422]_ , \new_[12423]_ , \new_[12424]_ ,
    \new_[12427]_ , \new_[12430]_ , \new_[12431]_ , \new_[12434]_ ,
    \new_[12438]_ , \new_[12439]_ , \new_[12440]_ , \new_[12443]_ ,
    \new_[12446]_ , \new_[12447]_ , \new_[12450]_ , \new_[12454]_ ,
    \new_[12455]_ , \new_[12456]_ , \new_[12459]_ , \new_[12462]_ ,
    \new_[12463]_ , \new_[12466]_ , \new_[12470]_ , \new_[12471]_ ,
    \new_[12472]_ , \new_[12475]_ , \new_[12478]_ , \new_[12479]_ ,
    \new_[12482]_ , \new_[12486]_ , \new_[12487]_ , \new_[12488]_ ,
    \new_[12491]_ , \new_[12494]_ , \new_[12495]_ , \new_[12498]_ ,
    \new_[12502]_ , \new_[12503]_ , \new_[12504]_ , \new_[12507]_ ,
    \new_[12510]_ , \new_[12511]_ , \new_[12514]_ , \new_[12518]_ ,
    \new_[12519]_ , \new_[12520]_ , \new_[12523]_ , \new_[12526]_ ,
    \new_[12527]_ , \new_[12530]_ , \new_[12534]_ , \new_[12535]_ ,
    \new_[12536]_ , \new_[12539]_ , \new_[12542]_ , \new_[12543]_ ,
    \new_[12546]_ , \new_[12550]_ , \new_[12551]_ , \new_[12552]_ ,
    \new_[12555]_ , \new_[12559]_ , \new_[12560]_ , \new_[12561]_ ,
    \new_[12564]_ , \new_[12568]_ , \new_[12569]_ , \new_[12570]_ ,
    \new_[12573]_ , \new_[12577]_ , \new_[12578]_ , \new_[12579]_ ,
    \new_[12582]_ , \new_[12586]_ , \new_[12587]_ , \new_[12588]_ ,
    \new_[12591]_ , \new_[12595]_ , \new_[12596]_ , \new_[12597]_ ,
    \new_[12600]_ , \new_[12604]_ , \new_[12605]_ , \new_[12606]_ ,
    \new_[12609]_ , \new_[12613]_ , \new_[12614]_ , \new_[12615]_ ,
    \new_[12618]_ , \new_[12622]_ , \new_[12623]_ , \new_[12624]_ ,
    \new_[12627]_ , \new_[12631]_ , \new_[12632]_ , \new_[12633]_ ,
    \new_[12636]_ , \new_[12640]_ , \new_[12641]_ , \new_[12642]_ ,
    \new_[12645]_ , \new_[12649]_ , \new_[12650]_ , \new_[12651]_ ,
    \new_[12654]_ , \new_[12658]_ , \new_[12659]_ , \new_[12660]_ ,
    \new_[12663]_ , \new_[12667]_ , \new_[12668]_ , \new_[12669]_ ,
    \new_[12672]_ , \new_[12676]_ , \new_[12677]_ , \new_[12678]_ ,
    \new_[12681]_ , \new_[12685]_ , \new_[12686]_ , \new_[12687]_ ,
    \new_[12690]_ , \new_[12694]_ , \new_[12695]_ , \new_[12696]_ ,
    \new_[12699]_ , \new_[12703]_ , \new_[12704]_ , \new_[12705]_ ,
    \new_[12708]_ , \new_[12712]_ , \new_[12713]_ , \new_[12714]_ ,
    \new_[12717]_ , \new_[12721]_ , \new_[12722]_ , \new_[12723]_ ,
    \new_[12726]_ , \new_[12730]_ , \new_[12731]_ , \new_[12732]_ ,
    \new_[12735]_ , \new_[12739]_ , \new_[12740]_ , \new_[12741]_ ,
    \new_[12744]_ , \new_[12748]_ , \new_[12749]_ , \new_[12750]_ ,
    \new_[12753]_ , \new_[12757]_ , \new_[12758]_ , \new_[12759]_ ,
    \new_[12762]_ , \new_[12766]_ , \new_[12767]_ , \new_[12768]_ ,
    \new_[12771]_ , \new_[12775]_ , \new_[12776]_ , \new_[12777]_ ,
    \new_[12780]_ , \new_[12784]_ , \new_[12785]_ , \new_[12786]_ ,
    \new_[12789]_ , \new_[12793]_ , \new_[12794]_ , \new_[12795]_ ,
    \new_[12798]_ , \new_[12802]_ , \new_[12803]_ , \new_[12804]_ ,
    \new_[12807]_ , \new_[12811]_ , \new_[12812]_ , \new_[12813]_ ,
    \new_[12816]_ , \new_[12820]_ , \new_[12821]_ , \new_[12822]_ ,
    \new_[12825]_ , \new_[12829]_ , \new_[12830]_ , \new_[12831]_ ,
    \new_[12834]_ , \new_[12838]_ , \new_[12839]_ , \new_[12840]_ ,
    \new_[12843]_ , \new_[12847]_ , \new_[12848]_ , \new_[12849]_ ,
    \new_[12852]_ , \new_[12856]_ , \new_[12857]_ , \new_[12858]_ ,
    \new_[12861]_ , \new_[12865]_ , \new_[12866]_ , \new_[12867]_ ,
    \new_[12870]_ , \new_[12874]_ , \new_[12875]_ , \new_[12876]_ ,
    \new_[12879]_ , \new_[12883]_ , \new_[12884]_ , \new_[12885]_ ,
    \new_[12888]_ , \new_[12892]_ , \new_[12893]_ , \new_[12894]_ ,
    \new_[12897]_ , \new_[12901]_ , \new_[12902]_ , \new_[12903]_ ,
    \new_[12906]_ , \new_[12910]_ , \new_[12911]_ , \new_[12912]_ ,
    \new_[12915]_ , \new_[12919]_ , \new_[12920]_ , \new_[12921]_ ,
    \new_[12924]_ , \new_[12928]_ , \new_[12929]_ , \new_[12930]_ ,
    \new_[12933]_ , \new_[12937]_ , \new_[12938]_ , \new_[12939]_ ,
    \new_[12942]_ , \new_[12946]_ , \new_[12947]_ , \new_[12948]_ ,
    \new_[12951]_ , \new_[12955]_ , \new_[12956]_ , \new_[12957]_ ,
    \new_[12960]_ , \new_[12964]_ , \new_[12965]_ , \new_[12966]_ ,
    \new_[12969]_ , \new_[12973]_ , \new_[12974]_ , \new_[12975]_ ,
    \new_[12978]_ , \new_[12982]_ , \new_[12983]_ , \new_[12984]_ ,
    \new_[12987]_ , \new_[12991]_ , \new_[12992]_ , \new_[12993]_ ,
    \new_[12996]_ , \new_[13000]_ , \new_[13001]_ , \new_[13002]_ ,
    \new_[13005]_ , \new_[13009]_ , \new_[13010]_ , \new_[13011]_ ,
    \new_[13014]_ , \new_[13018]_ , \new_[13019]_ , \new_[13020]_ ,
    \new_[13023]_ , \new_[13027]_ , \new_[13028]_ , \new_[13029]_ ,
    \new_[13032]_ , \new_[13036]_ , \new_[13037]_ , \new_[13038]_ ,
    \new_[13041]_ , \new_[13045]_ , \new_[13046]_ , \new_[13047]_ ,
    \new_[13050]_ , \new_[13054]_ , \new_[13055]_ , \new_[13056]_ ,
    \new_[13059]_ , \new_[13063]_ , \new_[13064]_ , \new_[13065]_ ,
    \new_[13068]_ , \new_[13072]_ , \new_[13073]_ , \new_[13074]_ ,
    \new_[13077]_ , \new_[13081]_ , \new_[13082]_ , \new_[13083]_ ,
    \new_[13086]_ , \new_[13090]_ , \new_[13091]_ , \new_[13092]_ ,
    \new_[13095]_ , \new_[13099]_ , \new_[13100]_ , \new_[13101]_ ,
    \new_[13104]_ , \new_[13108]_ , \new_[13109]_ , \new_[13110]_ ,
    \new_[13113]_ , \new_[13117]_ , \new_[13118]_ , \new_[13119]_ ,
    \new_[13122]_ , \new_[13126]_ , \new_[13127]_ , \new_[13128]_ ,
    \new_[13131]_ , \new_[13135]_ , \new_[13136]_ , \new_[13137]_ ,
    \new_[13140]_ , \new_[13144]_ , \new_[13145]_ , \new_[13146]_ ,
    \new_[13149]_ , \new_[13153]_ , \new_[13154]_ , \new_[13155]_ ,
    \new_[13158]_ , \new_[13162]_ , \new_[13163]_ , \new_[13164]_ ,
    \new_[13167]_ , \new_[13171]_ , \new_[13172]_ , \new_[13173]_ ,
    \new_[13176]_ , \new_[13180]_ , \new_[13181]_ , \new_[13182]_ ,
    \new_[13185]_ , \new_[13189]_ , \new_[13190]_ , \new_[13191]_ ,
    \new_[13194]_ , \new_[13198]_ , \new_[13199]_ , \new_[13200]_ ,
    \new_[13203]_ , \new_[13207]_ , \new_[13208]_ , \new_[13209]_ ,
    \new_[13212]_ , \new_[13216]_ , \new_[13217]_ , \new_[13218]_ ,
    \new_[13221]_ , \new_[13225]_ , \new_[13226]_ , \new_[13227]_ ,
    \new_[13230]_ , \new_[13234]_ , \new_[13235]_ , \new_[13236]_ ,
    \new_[13239]_ , \new_[13243]_ , \new_[13244]_ , \new_[13245]_ ,
    \new_[13248]_ , \new_[13252]_ , \new_[13253]_ , \new_[13254]_ ,
    \new_[13257]_ , \new_[13261]_ , \new_[13262]_ , \new_[13263]_ ,
    \new_[13266]_ , \new_[13270]_ , \new_[13271]_ , \new_[13272]_ ,
    \new_[13275]_ , \new_[13279]_ , \new_[13280]_ , \new_[13281]_ ,
    \new_[13284]_ , \new_[13288]_ , \new_[13289]_ , \new_[13290]_ ,
    \new_[13293]_ , \new_[13297]_ , \new_[13298]_ , \new_[13299]_ ,
    \new_[13302]_ , \new_[13306]_ , \new_[13307]_ , \new_[13308]_ ,
    \new_[13311]_ , \new_[13315]_ , \new_[13316]_ , \new_[13317]_ ,
    \new_[13320]_ , \new_[13324]_ , \new_[13325]_ , \new_[13326]_ ,
    \new_[13329]_ , \new_[13333]_ , \new_[13334]_ , \new_[13335]_ ,
    \new_[13338]_ , \new_[13342]_ , \new_[13343]_ , \new_[13344]_ ,
    \new_[13347]_ , \new_[13351]_ , \new_[13352]_ , \new_[13353]_ ,
    \new_[13356]_ , \new_[13360]_ , \new_[13361]_ , \new_[13362]_ ,
    \new_[13365]_ , \new_[13369]_ , \new_[13370]_ , \new_[13371]_ ,
    \new_[13374]_ , \new_[13378]_ , \new_[13379]_ , \new_[13380]_ ,
    \new_[13383]_ , \new_[13387]_ , \new_[13388]_ , \new_[13389]_ ,
    \new_[13392]_ , \new_[13396]_ , \new_[13397]_ , \new_[13398]_ ,
    \new_[13401]_ , \new_[13405]_ , \new_[13406]_ , \new_[13407]_ ,
    \new_[13410]_ , \new_[13414]_ , \new_[13415]_ , \new_[13416]_ ,
    \new_[13419]_ , \new_[13423]_ , \new_[13424]_ , \new_[13425]_ ,
    \new_[13428]_ , \new_[13432]_ , \new_[13433]_ , \new_[13434]_ ,
    \new_[13437]_ , \new_[13441]_ , \new_[13442]_ , \new_[13443]_ ,
    \new_[13446]_ , \new_[13450]_ , \new_[13451]_ , \new_[13452]_ ,
    \new_[13455]_ , \new_[13459]_ , \new_[13460]_ , \new_[13461]_ ,
    \new_[13464]_ , \new_[13468]_ , \new_[13469]_ , \new_[13470]_ ,
    \new_[13473]_ , \new_[13477]_ , \new_[13478]_ , \new_[13479]_ ,
    \new_[13482]_ , \new_[13486]_ , \new_[13487]_ , \new_[13488]_ ,
    \new_[13491]_ , \new_[13495]_ , \new_[13496]_ , \new_[13497]_ ,
    \new_[13500]_ , \new_[13504]_ , \new_[13505]_ , \new_[13506]_ ,
    \new_[13509]_ , \new_[13513]_ , \new_[13514]_ , \new_[13515]_ ,
    \new_[13518]_ , \new_[13522]_ , \new_[13523]_ , \new_[13524]_ ,
    \new_[13527]_ , \new_[13531]_ , \new_[13532]_ , \new_[13533]_ ,
    \new_[13536]_ , \new_[13540]_ , \new_[13541]_ , \new_[13542]_ ,
    \new_[13545]_ , \new_[13549]_ , \new_[13550]_ , \new_[13551]_ ,
    \new_[13554]_ , \new_[13558]_ , \new_[13559]_ , \new_[13560]_ ,
    \new_[13563]_ , \new_[13567]_ , \new_[13568]_ , \new_[13569]_ ,
    \new_[13572]_ , \new_[13576]_ , \new_[13577]_ , \new_[13578]_ ,
    \new_[13581]_ , \new_[13585]_ , \new_[13586]_ , \new_[13587]_ ,
    \new_[13590]_ , \new_[13594]_ , \new_[13595]_ , \new_[13596]_ ,
    \new_[13599]_ , \new_[13603]_ , \new_[13604]_ , \new_[13605]_ ,
    \new_[13608]_ , \new_[13612]_ , \new_[13613]_ , \new_[13614]_ ,
    \new_[13617]_ , \new_[13621]_ , \new_[13622]_ , \new_[13623]_ ,
    \new_[13626]_ , \new_[13630]_ , \new_[13631]_ , \new_[13632]_ ,
    \new_[13635]_ , \new_[13639]_ , \new_[13640]_ , \new_[13641]_ ,
    \new_[13644]_ , \new_[13648]_ , \new_[13649]_ , \new_[13650]_ ,
    \new_[13653]_ , \new_[13657]_ , \new_[13658]_ , \new_[13659]_ ,
    \new_[13662]_ , \new_[13666]_ , \new_[13667]_ , \new_[13668]_ ,
    \new_[13671]_ , \new_[13675]_ , \new_[13676]_ , \new_[13677]_ ,
    \new_[13680]_ , \new_[13684]_ , \new_[13685]_ , \new_[13686]_ ,
    \new_[13689]_ , \new_[13693]_ , \new_[13694]_ , \new_[13695]_ ,
    \new_[13698]_ , \new_[13702]_ , \new_[13703]_ , \new_[13704]_ ,
    \new_[13707]_ , \new_[13711]_ , \new_[13712]_ , \new_[13713]_ ,
    \new_[13716]_ , \new_[13720]_ , \new_[13721]_ , \new_[13722]_ ,
    \new_[13725]_ , \new_[13729]_ , \new_[13730]_ , \new_[13731]_ ,
    \new_[13734]_ , \new_[13738]_ , \new_[13739]_ , \new_[13740]_ ,
    \new_[13743]_ , \new_[13747]_ , \new_[13748]_ , \new_[13749]_ ,
    \new_[13752]_ , \new_[13756]_ , \new_[13757]_ , \new_[13758]_ ,
    \new_[13761]_ , \new_[13765]_ , \new_[13766]_ , \new_[13767]_ ,
    \new_[13770]_ , \new_[13774]_ , \new_[13775]_ , \new_[13776]_ ,
    \new_[13779]_ , \new_[13783]_ , \new_[13784]_ , \new_[13785]_ ,
    \new_[13788]_ , \new_[13792]_ , \new_[13793]_ , \new_[13794]_ ,
    \new_[13797]_ , \new_[13801]_ , \new_[13802]_ , \new_[13803]_ ,
    \new_[13806]_ , \new_[13810]_ , \new_[13811]_ , \new_[13812]_ ,
    \new_[13815]_ , \new_[13819]_ , \new_[13820]_ , \new_[13821]_ ,
    \new_[13824]_ , \new_[13828]_ , \new_[13829]_ , \new_[13830]_ ,
    \new_[13833]_ , \new_[13837]_ , \new_[13838]_ , \new_[13839]_ ,
    \new_[13842]_ , \new_[13846]_ , \new_[13847]_ , \new_[13848]_ ,
    \new_[13851]_ , \new_[13855]_ , \new_[13856]_ , \new_[13857]_ ,
    \new_[13860]_ , \new_[13864]_ , \new_[13865]_ , \new_[13866]_ ,
    \new_[13869]_ , \new_[13873]_ , \new_[13874]_ , \new_[13875]_ ,
    \new_[13878]_ , \new_[13882]_ , \new_[13883]_ , \new_[13884]_ ,
    \new_[13887]_ , \new_[13891]_ , \new_[13892]_ , \new_[13893]_ ,
    \new_[13896]_ , \new_[13900]_ , \new_[13901]_ , \new_[13902]_ ,
    \new_[13905]_ , \new_[13909]_ , \new_[13910]_ , \new_[13911]_ ,
    \new_[13914]_ , \new_[13918]_ , \new_[13919]_ , \new_[13920]_ ,
    \new_[13923]_ , \new_[13927]_ , \new_[13928]_ , \new_[13929]_ ,
    \new_[13932]_ , \new_[13936]_ , \new_[13937]_ , \new_[13938]_ ,
    \new_[13941]_ , \new_[13945]_ , \new_[13946]_ , \new_[13947]_ ,
    \new_[13950]_ , \new_[13954]_ , \new_[13955]_ , \new_[13956]_ ,
    \new_[13959]_ , \new_[13963]_ , \new_[13964]_ , \new_[13965]_ ,
    \new_[13968]_ , \new_[13972]_ , \new_[13973]_ , \new_[13974]_ ,
    \new_[13977]_ , \new_[13981]_ , \new_[13982]_ , \new_[13983]_ ,
    \new_[13986]_ , \new_[13990]_ , \new_[13991]_ , \new_[13992]_ ,
    \new_[13995]_ , \new_[13999]_ , \new_[14000]_ , \new_[14001]_ ,
    \new_[14004]_ , \new_[14008]_ , \new_[14009]_ , \new_[14010]_ ,
    \new_[14013]_ , \new_[14017]_ , \new_[14018]_ , \new_[14019]_ ,
    \new_[14022]_ , \new_[14026]_ , \new_[14027]_ , \new_[14028]_ ,
    \new_[14031]_ , \new_[14035]_ , \new_[14036]_ , \new_[14037]_ ,
    \new_[14040]_ , \new_[14044]_ , \new_[14045]_ , \new_[14046]_ ,
    \new_[14049]_ , \new_[14053]_ , \new_[14054]_ , \new_[14055]_ ,
    \new_[14058]_ , \new_[14062]_ , \new_[14063]_ , \new_[14064]_ ,
    \new_[14067]_ , \new_[14071]_ , \new_[14072]_ , \new_[14073]_ ,
    \new_[14076]_ , \new_[14080]_ , \new_[14081]_ , \new_[14082]_ ,
    \new_[14085]_ , \new_[14089]_ , \new_[14090]_ , \new_[14091]_ ,
    \new_[14094]_ , \new_[14098]_ , \new_[14099]_ , \new_[14100]_ ,
    \new_[14103]_ , \new_[14107]_ , \new_[14108]_ , \new_[14109]_ ,
    \new_[14112]_ , \new_[14116]_ , \new_[14117]_ , \new_[14118]_ ,
    \new_[14121]_ , \new_[14125]_ , \new_[14126]_ , \new_[14127]_ ,
    \new_[14130]_ , \new_[14134]_ , \new_[14135]_ , \new_[14136]_ ,
    \new_[14139]_ , \new_[14143]_ , \new_[14144]_ , \new_[14145]_ ,
    \new_[14148]_ , \new_[14152]_ , \new_[14153]_ , \new_[14154]_ ,
    \new_[14157]_ , \new_[14161]_ , \new_[14162]_ , \new_[14163]_ ,
    \new_[14166]_ , \new_[14170]_ , \new_[14171]_ , \new_[14172]_ ,
    \new_[14175]_ , \new_[14179]_ , \new_[14180]_ , \new_[14181]_ ,
    \new_[14184]_ , \new_[14188]_ , \new_[14189]_ , \new_[14190]_ ,
    \new_[14193]_ , \new_[14197]_ , \new_[14198]_ , \new_[14199]_ ,
    \new_[14202]_ , \new_[14206]_ , \new_[14207]_ , \new_[14208]_ ,
    \new_[14211]_ , \new_[14215]_ , \new_[14216]_ , \new_[14217]_ ,
    \new_[14220]_ , \new_[14224]_ , \new_[14225]_ , \new_[14226]_ ,
    \new_[14229]_ , \new_[14233]_ , \new_[14234]_ , \new_[14235]_ ,
    \new_[14238]_ , \new_[14242]_ , \new_[14243]_ , \new_[14244]_ ,
    \new_[14247]_ , \new_[14251]_ , \new_[14252]_ , \new_[14253]_ ,
    \new_[14256]_ , \new_[14260]_ , \new_[14261]_ , \new_[14262]_ ,
    \new_[14265]_ , \new_[14269]_ , \new_[14270]_ , \new_[14271]_ ,
    \new_[14274]_ , \new_[14278]_ , \new_[14279]_ , \new_[14280]_ ,
    \new_[14283]_ , \new_[14287]_ , \new_[14288]_ , \new_[14289]_ ,
    \new_[14292]_ , \new_[14296]_ , \new_[14297]_ , \new_[14298]_ ,
    \new_[14301]_ , \new_[14305]_ , \new_[14306]_ , \new_[14307]_ ,
    \new_[14310]_ , \new_[14314]_ , \new_[14315]_ , \new_[14316]_ ,
    \new_[14319]_ , \new_[14323]_ , \new_[14324]_ , \new_[14325]_ ,
    \new_[14328]_ , \new_[14332]_ , \new_[14333]_ , \new_[14334]_ ,
    \new_[14337]_ , \new_[14341]_ , \new_[14342]_ , \new_[14343]_ ,
    \new_[14346]_ , \new_[14350]_ , \new_[14351]_ , \new_[14352]_ ,
    \new_[14355]_ , \new_[14359]_ , \new_[14360]_ , \new_[14361]_ ,
    \new_[14364]_ , \new_[14368]_ , \new_[14369]_ , \new_[14370]_ ,
    \new_[14373]_ , \new_[14377]_ , \new_[14378]_ , \new_[14379]_ ,
    \new_[14382]_ , \new_[14386]_ , \new_[14387]_ , \new_[14388]_ ,
    \new_[14391]_ , \new_[14395]_ , \new_[14396]_ , \new_[14397]_ ,
    \new_[14400]_ , \new_[14404]_ , \new_[14405]_ , \new_[14406]_ ,
    \new_[14409]_ , \new_[14413]_ , \new_[14414]_ , \new_[14415]_ ,
    \new_[14418]_ , \new_[14422]_ , \new_[14423]_ , \new_[14424]_ ,
    \new_[14427]_ , \new_[14431]_ , \new_[14432]_ , \new_[14433]_ ,
    \new_[14436]_ , \new_[14440]_ , \new_[14441]_ , \new_[14442]_ ,
    \new_[14445]_ , \new_[14449]_ , \new_[14450]_ , \new_[14451]_ ,
    \new_[14454]_ , \new_[14458]_ , \new_[14459]_ , \new_[14460]_ ,
    \new_[14463]_ , \new_[14467]_ , \new_[14468]_ , \new_[14469]_ ,
    \new_[14472]_ , \new_[14476]_ , \new_[14477]_ , \new_[14478]_ ,
    \new_[14481]_ , \new_[14485]_ , \new_[14486]_ , \new_[14487]_ ,
    \new_[14490]_ , \new_[14494]_ , \new_[14495]_ , \new_[14496]_ ,
    \new_[14499]_ , \new_[14503]_ , \new_[14504]_ , \new_[14505]_ ,
    \new_[14508]_ , \new_[14512]_ , \new_[14513]_ , \new_[14514]_ ,
    \new_[14517]_ , \new_[14521]_ , \new_[14522]_ , \new_[14523]_ ,
    \new_[14526]_ , \new_[14530]_ , \new_[14531]_ , \new_[14532]_ ,
    \new_[14535]_ , \new_[14539]_ , \new_[14540]_ , \new_[14541]_ ,
    \new_[14544]_ , \new_[14548]_ , \new_[14549]_ , \new_[14550]_ ,
    \new_[14553]_ , \new_[14557]_ , \new_[14558]_ , \new_[14559]_ ,
    \new_[14562]_ , \new_[14566]_ , \new_[14567]_ , \new_[14568]_ ,
    \new_[14571]_ , \new_[14575]_ , \new_[14576]_ , \new_[14577]_ ,
    \new_[14580]_ , \new_[14584]_ , \new_[14585]_ , \new_[14586]_ ,
    \new_[14589]_ , \new_[14593]_ , \new_[14594]_ , \new_[14595]_ ,
    \new_[14598]_ , \new_[14602]_ , \new_[14603]_ , \new_[14604]_ ,
    \new_[14607]_ , \new_[14611]_ , \new_[14612]_ , \new_[14613]_ ,
    \new_[14616]_ , \new_[14620]_ , \new_[14621]_ , \new_[14622]_ ,
    \new_[14625]_ , \new_[14629]_ , \new_[14630]_ , \new_[14631]_ ,
    \new_[14634]_ , \new_[14638]_ , \new_[14639]_ , \new_[14640]_ ,
    \new_[14643]_ , \new_[14647]_ , \new_[14648]_ , \new_[14649]_ ,
    \new_[14652]_ , \new_[14656]_ , \new_[14657]_ , \new_[14658]_ ,
    \new_[14661]_ , \new_[14665]_ , \new_[14666]_ , \new_[14667]_ ,
    \new_[14670]_ , \new_[14674]_ , \new_[14675]_ , \new_[14676]_ ,
    \new_[14679]_ , \new_[14683]_ , \new_[14684]_ , \new_[14685]_ ,
    \new_[14688]_ , \new_[14692]_ , \new_[14693]_ , \new_[14694]_ ,
    \new_[14697]_ , \new_[14701]_ , \new_[14702]_ , \new_[14703]_ ,
    \new_[14706]_ , \new_[14710]_ , \new_[14711]_ , \new_[14712]_ ,
    \new_[14715]_ , \new_[14719]_ , \new_[14720]_ , \new_[14721]_ ,
    \new_[14724]_ , \new_[14728]_ , \new_[14729]_ , \new_[14730]_ ,
    \new_[14733]_ , \new_[14737]_ , \new_[14738]_ , \new_[14739]_ ,
    \new_[14742]_ , \new_[14746]_ , \new_[14747]_ , \new_[14748]_ ,
    \new_[14751]_ , \new_[14755]_ , \new_[14756]_ , \new_[14757]_ ,
    \new_[14760]_ , \new_[14764]_ , \new_[14765]_ , \new_[14766]_ ,
    \new_[14769]_ , \new_[14773]_ , \new_[14774]_ , \new_[14775]_ ,
    \new_[14778]_ , \new_[14782]_ , \new_[14783]_ , \new_[14784]_ ,
    \new_[14787]_ , \new_[14791]_ , \new_[14792]_ , \new_[14793]_ ,
    \new_[14796]_ , \new_[14800]_ , \new_[14801]_ , \new_[14802]_ ,
    \new_[14805]_ , \new_[14809]_ , \new_[14810]_ , \new_[14811]_ ,
    \new_[14814]_ , \new_[14818]_ , \new_[14819]_ , \new_[14820]_ ,
    \new_[14823]_ , \new_[14827]_ , \new_[14828]_ , \new_[14829]_ ,
    \new_[14832]_ , \new_[14836]_ , \new_[14837]_ , \new_[14838]_ ,
    \new_[14841]_ , \new_[14845]_ , \new_[14846]_ , \new_[14847]_ ,
    \new_[14850]_ , \new_[14854]_ , \new_[14855]_ , \new_[14856]_ ,
    \new_[14859]_ , \new_[14863]_ , \new_[14864]_ , \new_[14865]_ ,
    \new_[14868]_ , \new_[14872]_ , \new_[14873]_ , \new_[14874]_ ,
    \new_[14877]_ , \new_[14881]_ , \new_[14882]_ , \new_[14883]_ ,
    \new_[14886]_ , \new_[14890]_ , \new_[14891]_ , \new_[14892]_ ,
    \new_[14895]_ , \new_[14899]_ , \new_[14900]_ , \new_[14901]_ ,
    \new_[14904]_ , \new_[14908]_ , \new_[14909]_ , \new_[14910]_ ,
    \new_[14913]_ , \new_[14917]_ , \new_[14918]_ , \new_[14919]_ ,
    \new_[14922]_ , \new_[14926]_ , \new_[14927]_ , \new_[14928]_ ,
    \new_[14931]_ , \new_[14935]_ , \new_[14936]_ , \new_[14937]_ ,
    \new_[14940]_ , \new_[14944]_ , \new_[14945]_ , \new_[14946]_ ,
    \new_[14949]_ , \new_[14953]_ , \new_[14954]_ , \new_[14955]_ ,
    \new_[14958]_ , \new_[14962]_ , \new_[14963]_ , \new_[14964]_ ,
    \new_[14967]_ , \new_[14971]_ , \new_[14972]_ , \new_[14973]_ ,
    \new_[14976]_ , \new_[14980]_ , \new_[14981]_ , \new_[14982]_ ,
    \new_[14985]_ , \new_[14989]_ , \new_[14990]_ , \new_[14991]_ ,
    \new_[14994]_ , \new_[14998]_ , \new_[14999]_ , \new_[15000]_ ,
    \new_[15003]_ , \new_[15007]_ , \new_[15008]_ , \new_[15009]_ ,
    \new_[15012]_ , \new_[15016]_ , \new_[15017]_ , \new_[15018]_ ,
    \new_[15021]_ , \new_[15025]_ , \new_[15026]_ , \new_[15027]_ ,
    \new_[15030]_ , \new_[15034]_ , \new_[15035]_ , \new_[15036]_ ,
    \new_[15039]_ , \new_[15043]_ , \new_[15044]_ , \new_[15045]_ ,
    \new_[15048]_ , \new_[15052]_ , \new_[15053]_ , \new_[15054]_ ,
    \new_[15057]_ , \new_[15061]_ , \new_[15062]_ , \new_[15063]_ ,
    \new_[15066]_ , \new_[15070]_ , \new_[15071]_ , \new_[15072]_ ,
    \new_[15075]_ , \new_[15079]_ , \new_[15080]_ , \new_[15081]_ ,
    \new_[15084]_ , \new_[15088]_ , \new_[15089]_ , \new_[15090]_ ,
    \new_[15093]_ , \new_[15097]_ , \new_[15098]_ , \new_[15099]_ ,
    \new_[15102]_ , \new_[15106]_ , \new_[15107]_ , \new_[15108]_ ,
    \new_[15111]_ , \new_[15115]_ , \new_[15116]_ , \new_[15117]_ ,
    \new_[15120]_ , \new_[15124]_ , \new_[15125]_ , \new_[15126]_ ,
    \new_[15129]_ , \new_[15133]_ , \new_[15134]_ , \new_[15135]_ ,
    \new_[15138]_ , \new_[15142]_ , \new_[15143]_ , \new_[15144]_ ,
    \new_[15147]_ , \new_[15151]_ , \new_[15152]_ , \new_[15153]_ ,
    \new_[15156]_ , \new_[15160]_ , \new_[15161]_ , \new_[15162]_ ,
    \new_[15165]_ , \new_[15169]_ , \new_[15170]_ , \new_[15171]_ ,
    \new_[15174]_ , \new_[15178]_ , \new_[15179]_ , \new_[15180]_ ,
    \new_[15183]_ , \new_[15187]_ , \new_[15188]_ , \new_[15189]_ ,
    \new_[15192]_ , \new_[15196]_ , \new_[15197]_ , \new_[15198]_ ,
    \new_[15201]_ , \new_[15205]_ , \new_[15206]_ , \new_[15207]_ ,
    \new_[15210]_ , \new_[15214]_ , \new_[15215]_ , \new_[15216]_ ,
    \new_[15219]_ , \new_[15223]_ , \new_[15224]_ , \new_[15225]_ ,
    \new_[15228]_ , \new_[15232]_ , \new_[15233]_ , \new_[15234]_ ,
    \new_[15237]_ , \new_[15241]_ , \new_[15242]_ , \new_[15243]_ ,
    \new_[15246]_ , \new_[15250]_ , \new_[15251]_ , \new_[15252]_ ,
    \new_[15255]_ , \new_[15259]_ , \new_[15260]_ , \new_[15261]_ ,
    \new_[15264]_ , \new_[15268]_ , \new_[15269]_ , \new_[15270]_ ,
    \new_[15273]_ , \new_[15277]_ , \new_[15278]_ , \new_[15279]_ ,
    \new_[15282]_ , \new_[15286]_ , \new_[15287]_ , \new_[15288]_ ,
    \new_[15291]_ , \new_[15295]_ , \new_[15296]_ , \new_[15297]_ ,
    \new_[15300]_ , \new_[15304]_ , \new_[15305]_ , \new_[15306]_ ,
    \new_[15309]_ , \new_[15313]_ , \new_[15314]_ , \new_[15315]_ ,
    \new_[15318]_ , \new_[15322]_ , \new_[15323]_ , \new_[15324]_ ,
    \new_[15327]_ , \new_[15331]_ , \new_[15332]_ , \new_[15333]_ ,
    \new_[15336]_ , \new_[15340]_ , \new_[15341]_ , \new_[15342]_ ,
    \new_[15345]_ , \new_[15349]_ , \new_[15350]_ , \new_[15351]_ ,
    \new_[15354]_ , \new_[15358]_ , \new_[15359]_ , \new_[15360]_ ,
    \new_[15363]_ , \new_[15367]_ , \new_[15368]_ , \new_[15369]_ ,
    \new_[15372]_ , \new_[15376]_ , \new_[15377]_ , \new_[15378]_ ,
    \new_[15381]_ , \new_[15385]_ , \new_[15386]_ , \new_[15387]_ ,
    \new_[15390]_ , \new_[15394]_ , \new_[15395]_ , \new_[15396]_ ,
    \new_[15399]_ , \new_[15403]_ , \new_[15404]_ , \new_[15405]_ ,
    \new_[15408]_ , \new_[15412]_ , \new_[15413]_ , \new_[15414]_ ,
    \new_[15417]_ , \new_[15421]_ , \new_[15422]_ , \new_[15423]_ ,
    \new_[15426]_ , \new_[15430]_ , \new_[15431]_ , \new_[15432]_ ,
    \new_[15435]_ , \new_[15439]_ , \new_[15440]_ , \new_[15441]_ ,
    \new_[15444]_ , \new_[15448]_ , \new_[15449]_ , \new_[15450]_ ,
    \new_[15453]_ , \new_[15457]_ , \new_[15458]_ , \new_[15459]_ ,
    \new_[15462]_ , \new_[15466]_ , \new_[15467]_ , \new_[15468]_ ,
    \new_[15471]_ , \new_[15475]_ , \new_[15476]_ , \new_[15477]_ ,
    \new_[15480]_ , \new_[15484]_ , \new_[15485]_ , \new_[15486]_ ,
    \new_[15489]_ , \new_[15493]_ , \new_[15494]_ , \new_[15495]_ ,
    \new_[15498]_ , \new_[15502]_ , \new_[15503]_ , \new_[15504]_ ,
    \new_[15507]_ , \new_[15511]_ , \new_[15512]_ , \new_[15513]_ ,
    \new_[15516]_ , \new_[15520]_ , \new_[15521]_ , \new_[15522]_ ,
    \new_[15525]_ , \new_[15529]_ , \new_[15530]_ , \new_[15531]_ ,
    \new_[15534]_ , \new_[15538]_ , \new_[15539]_ , \new_[15540]_ ,
    \new_[15543]_ , \new_[15547]_ , \new_[15548]_ , \new_[15549]_ ,
    \new_[15552]_ , \new_[15556]_ , \new_[15557]_ , \new_[15558]_ ,
    \new_[15561]_ , \new_[15565]_ , \new_[15566]_ , \new_[15567]_ ,
    \new_[15570]_ , \new_[15574]_ , \new_[15575]_ , \new_[15576]_ ,
    \new_[15579]_ , \new_[15583]_ , \new_[15584]_ , \new_[15585]_ ,
    \new_[15588]_ , \new_[15592]_ , \new_[15593]_ , \new_[15594]_ ,
    \new_[15597]_ , \new_[15601]_ , \new_[15602]_ , \new_[15603]_ ,
    \new_[15606]_ , \new_[15610]_ , \new_[15611]_ , \new_[15612]_ ,
    \new_[15615]_ , \new_[15619]_ , \new_[15620]_ , \new_[15621]_ ,
    \new_[15624]_ , \new_[15628]_ , \new_[15629]_ , \new_[15630]_ ,
    \new_[15633]_ , \new_[15637]_ , \new_[15638]_ , \new_[15639]_ ,
    \new_[15642]_ , \new_[15646]_ , \new_[15647]_ , \new_[15648]_ ,
    \new_[15651]_ , \new_[15655]_ , \new_[15656]_ , \new_[15657]_ ,
    \new_[15660]_ , \new_[15664]_ , \new_[15665]_ , \new_[15666]_ ,
    \new_[15669]_ , \new_[15673]_ , \new_[15674]_ , \new_[15675]_ ,
    \new_[15678]_ , \new_[15682]_ , \new_[15683]_ , \new_[15684]_ ,
    \new_[15687]_ , \new_[15691]_ , \new_[15692]_ , \new_[15693]_ ,
    \new_[15696]_ , \new_[15700]_ , \new_[15701]_ , \new_[15702]_ ,
    \new_[15705]_ , \new_[15709]_ , \new_[15710]_ , \new_[15711]_ ,
    \new_[15714]_ , \new_[15718]_ , \new_[15719]_ , \new_[15720]_ ,
    \new_[15723]_ , \new_[15727]_ , \new_[15728]_ , \new_[15729]_ ,
    \new_[15732]_ , \new_[15736]_ , \new_[15737]_ , \new_[15738]_ ,
    \new_[15741]_ , \new_[15745]_ , \new_[15746]_ , \new_[15747]_ ,
    \new_[15750]_ , \new_[15754]_ , \new_[15755]_ , \new_[15756]_ ,
    \new_[15759]_ , \new_[15763]_ , \new_[15764]_ , \new_[15765]_ ,
    \new_[15768]_ , \new_[15772]_ , \new_[15773]_ , \new_[15774]_ ,
    \new_[15777]_ , \new_[15781]_ , \new_[15782]_ , \new_[15783]_ ,
    \new_[15786]_ , \new_[15790]_ , \new_[15791]_ , \new_[15792]_ ,
    \new_[15795]_ , \new_[15799]_ , \new_[15800]_ , \new_[15801]_ ,
    \new_[15804]_ , \new_[15808]_ , \new_[15809]_ , \new_[15810]_ ,
    \new_[15813]_ , \new_[15817]_ , \new_[15818]_ , \new_[15819]_ ,
    \new_[15822]_ , \new_[15826]_ , \new_[15827]_ , \new_[15828]_ ,
    \new_[15831]_ , \new_[15835]_ , \new_[15836]_ , \new_[15837]_ ,
    \new_[15840]_ , \new_[15844]_ , \new_[15845]_ , \new_[15846]_ ,
    \new_[15849]_ , \new_[15853]_ , \new_[15854]_ , \new_[15855]_ ,
    \new_[15858]_ , \new_[15862]_ , \new_[15863]_ , \new_[15864]_ ,
    \new_[15867]_ , \new_[15871]_ , \new_[15872]_ , \new_[15873]_ ,
    \new_[15876]_ , \new_[15880]_ , \new_[15881]_ , \new_[15882]_ ,
    \new_[15885]_ , \new_[15889]_ , \new_[15890]_ , \new_[15891]_ ,
    \new_[15894]_ , \new_[15898]_ , \new_[15899]_ , \new_[15900]_ ,
    \new_[15903]_ , \new_[15907]_ , \new_[15908]_ , \new_[15909]_ ,
    \new_[15912]_ , \new_[15916]_ , \new_[15917]_ , \new_[15918]_ ,
    \new_[15921]_ , \new_[15925]_ , \new_[15926]_ , \new_[15927]_ ,
    \new_[15930]_ , \new_[15934]_ , \new_[15935]_ , \new_[15936]_ ,
    \new_[15939]_ , \new_[15943]_ , \new_[15944]_ , \new_[15945]_ ,
    \new_[15948]_ , \new_[15952]_ , \new_[15953]_ , \new_[15954]_ ,
    \new_[15957]_ , \new_[15961]_ , \new_[15962]_ , \new_[15963]_ ,
    \new_[15966]_ , \new_[15970]_ , \new_[15971]_ , \new_[15972]_ ,
    \new_[15975]_ , \new_[15979]_ , \new_[15980]_ , \new_[15981]_ ,
    \new_[15984]_ , \new_[15988]_ , \new_[15989]_ , \new_[15990]_ ,
    \new_[15993]_ , \new_[15997]_ , \new_[15998]_ , \new_[15999]_ ,
    \new_[16002]_ , \new_[16006]_ , \new_[16007]_ , \new_[16008]_ ,
    \new_[16011]_ , \new_[16015]_ , \new_[16016]_ , \new_[16017]_ ,
    \new_[16020]_ , \new_[16024]_ , \new_[16025]_ , \new_[16026]_ ,
    \new_[16029]_ , \new_[16033]_ , \new_[16034]_ , \new_[16035]_ ,
    \new_[16038]_ , \new_[16042]_ , \new_[16043]_ , \new_[16044]_ ,
    \new_[16047]_ , \new_[16051]_ , \new_[16052]_ , \new_[16053]_ ,
    \new_[16056]_ , \new_[16060]_ , \new_[16061]_ , \new_[16062]_ ,
    \new_[16065]_ , \new_[16069]_ , \new_[16070]_ , \new_[16071]_ ,
    \new_[16074]_ , \new_[16078]_ , \new_[16079]_ , \new_[16080]_ ,
    \new_[16083]_ , \new_[16087]_ , \new_[16088]_ , \new_[16089]_ ,
    \new_[16092]_ , \new_[16096]_ , \new_[16097]_ , \new_[16098]_ ,
    \new_[16101]_ , \new_[16105]_ , \new_[16106]_ , \new_[16107]_ ,
    \new_[16110]_ , \new_[16114]_ , \new_[16115]_ , \new_[16116]_ ,
    \new_[16119]_ , \new_[16123]_ , \new_[16124]_ , \new_[16125]_ ,
    \new_[16128]_ , \new_[16132]_ , \new_[16133]_ , \new_[16134]_ ,
    \new_[16137]_ , \new_[16141]_ , \new_[16142]_ , \new_[16143]_ ,
    \new_[16146]_ , \new_[16150]_ , \new_[16151]_ , \new_[16152]_ ,
    \new_[16155]_ , \new_[16159]_ , \new_[16160]_ , \new_[16161]_ ,
    \new_[16164]_ , \new_[16168]_ , \new_[16169]_ , \new_[16170]_ ,
    \new_[16173]_ , \new_[16177]_ , \new_[16178]_ , \new_[16179]_ ,
    \new_[16182]_ , \new_[16186]_ , \new_[16187]_ , \new_[16188]_ ,
    \new_[16191]_ , \new_[16195]_ , \new_[16196]_ , \new_[16197]_ ,
    \new_[16200]_ , \new_[16204]_ , \new_[16205]_ , \new_[16206]_ ,
    \new_[16209]_ , \new_[16213]_ , \new_[16214]_ , \new_[16215]_ ,
    \new_[16218]_ , \new_[16222]_ , \new_[16223]_ , \new_[16224]_ ,
    \new_[16227]_ , \new_[16231]_ , \new_[16232]_ , \new_[16233]_ ,
    \new_[16236]_ , \new_[16240]_ , \new_[16241]_ , \new_[16242]_ ,
    \new_[16245]_ , \new_[16249]_ , \new_[16250]_ , \new_[16251]_ ,
    \new_[16254]_ , \new_[16258]_ , \new_[16259]_ , \new_[16260]_ ,
    \new_[16263]_ , \new_[16267]_ , \new_[16268]_ , \new_[16269]_ ,
    \new_[16272]_ , \new_[16276]_ , \new_[16277]_ , \new_[16278]_ ,
    \new_[16281]_ , \new_[16285]_ , \new_[16286]_ , \new_[16287]_ ,
    \new_[16290]_ , \new_[16294]_ , \new_[16295]_ , \new_[16296]_ ,
    \new_[16299]_ , \new_[16303]_ , \new_[16304]_ , \new_[16305]_ ,
    \new_[16308]_ , \new_[16312]_ , \new_[16313]_ , \new_[16314]_ ,
    \new_[16317]_ , \new_[16321]_ , \new_[16322]_ , \new_[16323]_ ,
    \new_[16326]_ , \new_[16330]_ , \new_[16331]_ , \new_[16332]_ ,
    \new_[16335]_ , \new_[16339]_ , \new_[16340]_ , \new_[16341]_ ,
    \new_[16344]_ , \new_[16348]_ , \new_[16349]_ , \new_[16350]_ ,
    \new_[16353]_ , \new_[16357]_ , \new_[16358]_ , \new_[16359]_ ,
    \new_[16362]_ , \new_[16366]_ , \new_[16367]_ , \new_[16368]_ ,
    \new_[16371]_ , \new_[16375]_ , \new_[16376]_ , \new_[16377]_ ,
    \new_[16380]_ , \new_[16384]_ , \new_[16385]_ , \new_[16386]_ ,
    \new_[16389]_ , \new_[16393]_ , \new_[16394]_ , \new_[16395]_ ,
    \new_[16398]_ , \new_[16402]_ , \new_[16403]_ , \new_[16404]_ ,
    \new_[16407]_ , \new_[16411]_ , \new_[16412]_ , \new_[16413]_ ,
    \new_[16416]_ , \new_[16420]_ , \new_[16421]_ , \new_[16422]_ ,
    \new_[16425]_ , \new_[16429]_ , \new_[16430]_ , \new_[16431]_ ,
    \new_[16434]_ , \new_[16438]_ , \new_[16439]_ , \new_[16440]_ ,
    \new_[16443]_ , \new_[16447]_ , \new_[16448]_ , \new_[16449]_ ,
    \new_[16452]_ , \new_[16456]_ , \new_[16457]_ , \new_[16458]_ ,
    \new_[16461]_ , \new_[16465]_ , \new_[16466]_ , \new_[16467]_ ,
    \new_[16470]_ , \new_[16474]_ , \new_[16475]_ , \new_[16476]_ ,
    \new_[16479]_ , \new_[16483]_ , \new_[16484]_ , \new_[16485]_ ,
    \new_[16488]_ , \new_[16492]_ , \new_[16493]_ , \new_[16494]_ ,
    \new_[16497]_ , \new_[16501]_ , \new_[16502]_ , \new_[16503]_ ,
    \new_[16506]_ , \new_[16510]_ , \new_[16511]_ , \new_[16512]_ ,
    \new_[16515]_ , \new_[16519]_ , \new_[16520]_ , \new_[16521]_ ,
    \new_[16524]_ , \new_[16528]_ , \new_[16529]_ , \new_[16530]_ ,
    \new_[16533]_ , \new_[16537]_ , \new_[16538]_ , \new_[16539]_ ,
    \new_[16542]_ , \new_[16546]_ , \new_[16547]_ , \new_[16548]_ ,
    \new_[16551]_ , \new_[16555]_ , \new_[16556]_ , \new_[16557]_ ,
    \new_[16560]_ , \new_[16564]_ , \new_[16565]_ , \new_[16566]_ ,
    \new_[16569]_ , \new_[16573]_ , \new_[16574]_ , \new_[16575]_ ,
    \new_[16578]_ , \new_[16582]_ , \new_[16583]_ , \new_[16584]_ ,
    \new_[16587]_ , \new_[16591]_ , \new_[16592]_ , \new_[16593]_ ,
    \new_[16596]_ , \new_[16600]_ , \new_[16601]_ , \new_[16602]_ ,
    \new_[16605]_ , \new_[16609]_ , \new_[16610]_ , \new_[16611]_ ,
    \new_[16614]_ , \new_[16618]_ , \new_[16619]_ , \new_[16620]_ ,
    \new_[16623]_ , \new_[16627]_ , \new_[16628]_ , \new_[16629]_ ,
    \new_[16632]_ , \new_[16636]_ , \new_[16637]_ , \new_[16638]_ ,
    \new_[16641]_ , \new_[16645]_ , \new_[16646]_ , \new_[16647]_ ,
    \new_[16650]_ , \new_[16654]_ , \new_[16655]_ , \new_[16656]_ ,
    \new_[16659]_ , \new_[16663]_ , \new_[16664]_ , \new_[16665]_ ,
    \new_[16668]_ , \new_[16672]_ , \new_[16673]_ , \new_[16674]_ ,
    \new_[16677]_ , \new_[16681]_ , \new_[16682]_ , \new_[16683]_ ,
    \new_[16686]_ , \new_[16690]_ , \new_[16691]_ , \new_[16692]_ ,
    \new_[16695]_ , \new_[16699]_ , \new_[16700]_ , \new_[16701]_ ,
    \new_[16704]_ , \new_[16708]_ , \new_[16709]_ , \new_[16710]_ ,
    \new_[16713]_ , \new_[16717]_ , \new_[16718]_ , \new_[16719]_ ,
    \new_[16722]_ , \new_[16726]_ , \new_[16727]_ , \new_[16728]_ ,
    \new_[16731]_ , \new_[16735]_ , \new_[16736]_ , \new_[16737]_ ,
    \new_[16740]_ , \new_[16744]_ , \new_[16745]_ , \new_[16746]_ ,
    \new_[16749]_ , \new_[16753]_ , \new_[16754]_ , \new_[16755]_ ,
    \new_[16758]_ , \new_[16762]_ , \new_[16763]_ , \new_[16764]_ ,
    \new_[16767]_ , \new_[16771]_ , \new_[16772]_ , \new_[16773]_ ,
    \new_[16776]_ , \new_[16780]_ , \new_[16781]_ , \new_[16782]_ ,
    \new_[16785]_ , \new_[16789]_ , \new_[16790]_ , \new_[16791]_ ,
    \new_[16794]_ , \new_[16798]_ , \new_[16799]_ , \new_[16800]_ ,
    \new_[16803]_ , \new_[16807]_ , \new_[16808]_ , \new_[16809]_ ,
    \new_[16812]_ , \new_[16816]_ , \new_[16817]_ , \new_[16818]_ ,
    \new_[16821]_ , \new_[16825]_ , \new_[16826]_ , \new_[16827]_ ,
    \new_[16830]_ , \new_[16834]_ , \new_[16835]_ , \new_[16836]_ ,
    \new_[16839]_ , \new_[16843]_ , \new_[16844]_ , \new_[16845]_ ,
    \new_[16848]_ , \new_[16852]_ , \new_[16853]_ , \new_[16854]_ ,
    \new_[16857]_ , \new_[16861]_ , \new_[16862]_ , \new_[16863]_ ,
    \new_[16866]_ , \new_[16870]_ , \new_[16871]_ , \new_[16872]_ ,
    \new_[16875]_ , \new_[16879]_ , \new_[16880]_ , \new_[16881]_ ,
    \new_[16884]_ , \new_[16888]_ , \new_[16889]_ , \new_[16890]_ ,
    \new_[16893]_ , \new_[16897]_ , \new_[16898]_ , \new_[16899]_ ,
    \new_[16902]_ , \new_[16906]_ , \new_[16907]_ , \new_[16908]_ ,
    \new_[16911]_ , \new_[16915]_ , \new_[16916]_ , \new_[16917]_ ,
    \new_[16920]_ , \new_[16924]_ , \new_[16925]_ , \new_[16926]_ ,
    \new_[16929]_ , \new_[16933]_ , \new_[16934]_ , \new_[16935]_ ,
    \new_[16938]_ , \new_[16942]_ , \new_[16943]_ , \new_[16944]_ ,
    \new_[16947]_ , \new_[16951]_ , \new_[16952]_ , \new_[16953]_ ,
    \new_[16956]_ , \new_[16960]_ , \new_[16961]_ , \new_[16962]_ ,
    \new_[16965]_ , \new_[16969]_ , \new_[16970]_ , \new_[16971]_ ,
    \new_[16974]_ , \new_[16978]_ , \new_[16979]_ , \new_[16980]_ ,
    \new_[16983]_ , \new_[16987]_ , \new_[16988]_ , \new_[16989]_ ,
    \new_[16992]_ , \new_[16996]_ , \new_[16997]_ , \new_[16998]_ ,
    \new_[17001]_ , \new_[17005]_ , \new_[17006]_ , \new_[17007]_ ,
    \new_[17010]_ , \new_[17014]_ , \new_[17015]_ , \new_[17016]_ ,
    \new_[17019]_ , \new_[17023]_ , \new_[17024]_ , \new_[17025]_ ,
    \new_[17028]_ , \new_[17032]_ , \new_[17033]_ , \new_[17034]_ ,
    \new_[17037]_ , \new_[17041]_ , \new_[17042]_ , \new_[17043]_ ,
    \new_[17046]_ , \new_[17050]_ , \new_[17051]_ , \new_[17052]_ ,
    \new_[17055]_ , \new_[17059]_ , \new_[17060]_ , \new_[17061]_ ,
    \new_[17064]_ , \new_[17068]_ , \new_[17069]_ , \new_[17070]_ ,
    \new_[17073]_ , \new_[17077]_ , \new_[17078]_ , \new_[17079]_ ,
    \new_[17082]_ , \new_[17086]_ , \new_[17087]_ , \new_[17088]_ ,
    \new_[17091]_ , \new_[17095]_ , \new_[17096]_ , \new_[17097]_ ,
    \new_[17100]_ , \new_[17104]_ , \new_[17105]_ , \new_[17106]_ ,
    \new_[17109]_ , \new_[17113]_ , \new_[17114]_ , \new_[17115]_ ,
    \new_[17118]_ , \new_[17122]_ , \new_[17123]_ , \new_[17124]_ ,
    \new_[17127]_ , \new_[17131]_ , \new_[17132]_ , \new_[17133]_ ,
    \new_[17136]_ , \new_[17140]_ , \new_[17141]_ , \new_[17142]_ ,
    \new_[17145]_ , \new_[17149]_ , \new_[17150]_ , \new_[17151]_ ,
    \new_[17154]_ , \new_[17158]_ , \new_[17159]_ , \new_[17160]_ ,
    \new_[17163]_ , \new_[17167]_ , \new_[17168]_ , \new_[17169]_ ,
    \new_[17172]_ , \new_[17176]_ , \new_[17177]_ , \new_[17178]_ ,
    \new_[17181]_ , \new_[17185]_ , \new_[17186]_ , \new_[17187]_ ,
    \new_[17190]_ , \new_[17194]_ , \new_[17195]_ , \new_[17196]_ ,
    \new_[17199]_ , \new_[17203]_ , \new_[17204]_ , \new_[17205]_ ,
    \new_[17208]_ , \new_[17212]_ , \new_[17213]_ , \new_[17214]_ ,
    \new_[17217]_ , \new_[17221]_ , \new_[17222]_ , \new_[17223]_ ,
    \new_[17226]_ , \new_[17230]_ , \new_[17231]_ , \new_[17232]_ ,
    \new_[17235]_ , \new_[17239]_ , \new_[17240]_ , \new_[17241]_ ,
    \new_[17244]_ , \new_[17248]_ , \new_[17249]_ , \new_[17250]_ ,
    \new_[17253]_ , \new_[17257]_ , \new_[17258]_ , \new_[17259]_ ,
    \new_[17262]_ , \new_[17266]_ , \new_[17267]_ , \new_[17268]_ ,
    \new_[17271]_ , \new_[17275]_ , \new_[17276]_ , \new_[17277]_ ,
    \new_[17280]_ , \new_[17284]_ , \new_[17285]_ , \new_[17286]_ ,
    \new_[17289]_ , \new_[17293]_ , \new_[17294]_ , \new_[17295]_ ,
    \new_[17298]_ , \new_[17302]_ , \new_[17303]_ , \new_[17304]_ ,
    \new_[17307]_ , \new_[17311]_ , \new_[17312]_ , \new_[17313]_ ,
    \new_[17316]_ , \new_[17320]_ , \new_[17321]_ , \new_[17322]_ ,
    \new_[17325]_ , \new_[17329]_ , \new_[17330]_ , \new_[17331]_ ,
    \new_[17334]_ , \new_[17338]_ , \new_[17339]_ , \new_[17340]_ ,
    \new_[17343]_ , \new_[17347]_ , \new_[17348]_ , \new_[17349]_ ,
    \new_[17352]_ , \new_[17356]_ , \new_[17357]_ , \new_[17358]_ ,
    \new_[17361]_ , \new_[17365]_ , \new_[17366]_ , \new_[17367]_ ,
    \new_[17370]_ , \new_[17374]_ , \new_[17375]_ , \new_[17376]_ ,
    \new_[17379]_ , \new_[17383]_ , \new_[17384]_ , \new_[17385]_ ,
    \new_[17388]_ , \new_[17392]_ , \new_[17393]_ , \new_[17394]_ ,
    \new_[17397]_ , \new_[17401]_ , \new_[17402]_ , \new_[17403]_ ,
    \new_[17406]_ , \new_[17410]_ , \new_[17411]_ , \new_[17412]_ ,
    \new_[17415]_ , \new_[17419]_ , \new_[17420]_ , \new_[17421]_ ,
    \new_[17424]_ , \new_[17428]_ , \new_[17429]_ , \new_[17430]_ ,
    \new_[17433]_ , \new_[17437]_ , \new_[17438]_ , \new_[17439]_ ,
    \new_[17442]_ , \new_[17446]_ , \new_[17447]_ , \new_[17448]_ ,
    \new_[17451]_ , \new_[17455]_ , \new_[17456]_ , \new_[17457]_ ,
    \new_[17460]_ , \new_[17464]_ , \new_[17465]_ , \new_[17466]_ ,
    \new_[17469]_ , \new_[17473]_ , \new_[17474]_ , \new_[17475]_ ,
    \new_[17478]_ , \new_[17482]_ , \new_[17483]_ , \new_[17484]_ ,
    \new_[17487]_ , \new_[17491]_ , \new_[17492]_ , \new_[17493]_ ,
    \new_[17496]_ , \new_[17500]_ , \new_[17501]_ , \new_[17502]_ ,
    \new_[17505]_ , \new_[17509]_ , \new_[17510]_ , \new_[17511]_ ,
    \new_[17514]_ , \new_[17518]_ , \new_[17519]_ , \new_[17520]_ ,
    \new_[17523]_ , \new_[17527]_ , \new_[17528]_ , \new_[17529]_ ,
    \new_[17532]_ , \new_[17536]_ , \new_[17537]_ , \new_[17538]_ ,
    \new_[17541]_ , \new_[17545]_ , \new_[17546]_ , \new_[17547]_ ,
    \new_[17550]_ , \new_[17554]_ , \new_[17555]_ , \new_[17556]_ ,
    \new_[17559]_ , \new_[17563]_ , \new_[17564]_ , \new_[17565]_ ,
    \new_[17568]_ , \new_[17572]_ , \new_[17573]_ , \new_[17574]_ ,
    \new_[17577]_ , \new_[17581]_ , \new_[17582]_ , \new_[17583]_ ,
    \new_[17586]_ , \new_[17590]_ , \new_[17591]_ , \new_[17592]_ ,
    \new_[17595]_ , \new_[17599]_ , \new_[17600]_ , \new_[17601]_ ,
    \new_[17604]_ , \new_[17608]_ , \new_[17609]_ , \new_[17610]_ ,
    \new_[17613]_ , \new_[17617]_ , \new_[17618]_ , \new_[17619]_ ,
    \new_[17622]_ , \new_[17626]_ , \new_[17627]_ , \new_[17628]_ ,
    \new_[17631]_ , \new_[17635]_ , \new_[17636]_ , \new_[17637]_ ,
    \new_[17640]_ , \new_[17644]_ , \new_[17645]_ , \new_[17646]_ ,
    \new_[17649]_ , \new_[17653]_ , \new_[17654]_ , \new_[17655]_ ,
    \new_[17658]_ , \new_[17662]_ , \new_[17663]_ , \new_[17664]_ ,
    \new_[17667]_ , \new_[17671]_ , \new_[17672]_ , \new_[17673]_ ,
    \new_[17676]_ , \new_[17680]_ , \new_[17681]_ , \new_[17682]_ ,
    \new_[17685]_ , \new_[17689]_ , \new_[17690]_ , \new_[17691]_ ,
    \new_[17694]_ , \new_[17698]_ , \new_[17699]_ , \new_[17700]_ ,
    \new_[17703]_ , \new_[17707]_ , \new_[17708]_ , \new_[17709]_ ,
    \new_[17712]_ , \new_[17716]_ , \new_[17717]_ , \new_[17718]_ ,
    \new_[17721]_ , \new_[17725]_ , \new_[17726]_ , \new_[17727]_ ,
    \new_[17730]_ , \new_[17734]_ , \new_[17735]_ , \new_[17736]_ ,
    \new_[17739]_ , \new_[17743]_ , \new_[17744]_ , \new_[17745]_ ,
    \new_[17748]_ , \new_[17752]_ , \new_[17753]_ , \new_[17754]_ ,
    \new_[17757]_ , \new_[17761]_ , \new_[17762]_ , \new_[17763]_ ,
    \new_[17766]_ , \new_[17770]_ , \new_[17771]_ , \new_[17772]_ ,
    \new_[17775]_ , \new_[17779]_ , \new_[17780]_ , \new_[17781]_ ,
    \new_[17784]_ , \new_[17788]_ , \new_[17789]_ , \new_[17790]_ ,
    \new_[17793]_ , \new_[17797]_ , \new_[17798]_ , \new_[17799]_ ,
    \new_[17802]_ , \new_[17806]_ , \new_[17807]_ , \new_[17808]_ ,
    \new_[17811]_ , \new_[17815]_ , \new_[17816]_ , \new_[17817]_ ,
    \new_[17820]_ , \new_[17824]_ , \new_[17825]_ , \new_[17826]_ ,
    \new_[17829]_ , \new_[17833]_ , \new_[17834]_ , \new_[17835]_ ,
    \new_[17838]_ , \new_[17842]_ , \new_[17843]_ , \new_[17844]_ ,
    \new_[17847]_ , \new_[17851]_ , \new_[17852]_ , \new_[17853]_ ,
    \new_[17856]_ , \new_[17860]_ , \new_[17861]_ , \new_[17862]_ ,
    \new_[17865]_ , \new_[17869]_ , \new_[17870]_ , \new_[17871]_ ,
    \new_[17874]_ , \new_[17878]_ , \new_[17879]_ , \new_[17880]_ ,
    \new_[17883]_ , \new_[17887]_ , \new_[17888]_ , \new_[17889]_ ,
    \new_[17892]_ , \new_[17896]_ , \new_[17897]_ , \new_[17898]_ ,
    \new_[17901]_ , \new_[17905]_ , \new_[17906]_ , \new_[17907]_ ,
    \new_[17910]_ , \new_[17914]_ , \new_[17915]_ , \new_[17916]_ ,
    \new_[17919]_ , \new_[17923]_ , \new_[17924]_ , \new_[17925]_ ,
    \new_[17928]_ , \new_[17932]_ , \new_[17933]_ , \new_[17934]_ ,
    \new_[17937]_ , \new_[17941]_ , \new_[17942]_ , \new_[17943]_ ,
    \new_[17946]_ , \new_[17950]_ , \new_[17951]_ , \new_[17952]_ ,
    \new_[17955]_ , \new_[17959]_ , \new_[17960]_ , \new_[17961]_ ,
    \new_[17964]_ , \new_[17968]_ , \new_[17969]_ , \new_[17970]_ ,
    \new_[17973]_ , \new_[17977]_ , \new_[17978]_ , \new_[17979]_ ,
    \new_[17982]_ , \new_[17986]_ , \new_[17987]_ , \new_[17988]_ ,
    \new_[17991]_ , \new_[17995]_ , \new_[17996]_ , \new_[17997]_ ,
    \new_[18000]_ , \new_[18004]_ , \new_[18005]_ , \new_[18006]_ ,
    \new_[18009]_ , \new_[18013]_ , \new_[18014]_ , \new_[18015]_ ,
    \new_[18018]_ , \new_[18022]_ , \new_[18023]_ , \new_[18024]_ ,
    \new_[18027]_ , \new_[18031]_ , \new_[18032]_ , \new_[18033]_ ,
    \new_[18036]_ , \new_[18040]_ , \new_[18041]_ , \new_[18042]_ ,
    \new_[18045]_ , \new_[18049]_ , \new_[18050]_ , \new_[18051]_ ,
    \new_[18054]_ , \new_[18058]_ , \new_[18059]_ , \new_[18060]_ ,
    \new_[18063]_ , \new_[18067]_ , \new_[18068]_ , \new_[18069]_ ,
    \new_[18073]_ , \new_[18074]_ , \new_[18078]_ , \new_[18079]_ ,
    \new_[18080]_ , \new_[18083]_ , \new_[18087]_ , \new_[18088]_ ,
    \new_[18089]_ , \new_[18093]_ , \new_[18094]_ , \new_[18098]_ ,
    \new_[18099]_ , \new_[18100]_ , \new_[18103]_ , \new_[18107]_ ,
    \new_[18108]_ , \new_[18109]_ , \new_[18113]_ , \new_[18114]_ ,
    \new_[18118]_ , \new_[18119]_ , \new_[18120]_ , \new_[18123]_ ,
    \new_[18127]_ , \new_[18128]_ , \new_[18129]_ , \new_[18133]_ ,
    \new_[18134]_ , \new_[18138]_ , \new_[18139]_ , \new_[18140]_ ,
    \new_[18143]_ , \new_[18147]_ , \new_[18148]_ , \new_[18149]_ ,
    \new_[18153]_ , \new_[18154]_ , \new_[18158]_ , \new_[18159]_ ,
    \new_[18160]_ , \new_[18163]_ , \new_[18167]_ , \new_[18168]_ ,
    \new_[18169]_ , \new_[18173]_ , \new_[18174]_ , \new_[18178]_ ,
    \new_[18179]_ , \new_[18180]_ , \new_[18183]_ , \new_[18187]_ ,
    \new_[18188]_ , \new_[18189]_ , \new_[18193]_ , \new_[18194]_ ,
    \new_[18198]_ , \new_[18199]_ , \new_[18200]_ , \new_[18203]_ ,
    \new_[18207]_ , \new_[18208]_ , \new_[18209]_ , \new_[18213]_ ,
    \new_[18214]_ , \new_[18218]_ , \new_[18219]_ , \new_[18220]_ ,
    \new_[18223]_ , \new_[18227]_ , \new_[18228]_ , \new_[18229]_ ,
    \new_[18233]_ , \new_[18234]_ , \new_[18238]_ , \new_[18239]_ ,
    \new_[18240]_ , \new_[18243]_ , \new_[18247]_ , \new_[18248]_ ,
    \new_[18249]_ , \new_[18253]_ , \new_[18254]_ , \new_[18258]_ ,
    \new_[18259]_ , \new_[18260]_ , \new_[18263]_ , \new_[18267]_ ,
    \new_[18268]_ , \new_[18269]_ , \new_[18273]_ , \new_[18274]_ ,
    \new_[18278]_ , \new_[18279]_ , \new_[18280]_ , \new_[18283]_ ,
    \new_[18287]_ , \new_[18288]_ , \new_[18289]_ , \new_[18293]_ ,
    \new_[18294]_ , \new_[18298]_ , \new_[18299]_ , \new_[18300]_ ,
    \new_[18303]_ , \new_[18307]_ , \new_[18308]_ , \new_[18309]_ ,
    \new_[18313]_ , \new_[18314]_ , \new_[18318]_ , \new_[18319]_ ,
    \new_[18320]_ , \new_[18323]_ , \new_[18327]_ , \new_[18328]_ ,
    \new_[18329]_ , \new_[18333]_ , \new_[18334]_ , \new_[18338]_ ,
    \new_[18339]_ , \new_[18340]_ , \new_[18343]_ , \new_[18347]_ ,
    \new_[18348]_ , \new_[18349]_ , \new_[18353]_ , \new_[18354]_ ,
    \new_[18358]_ , \new_[18359]_ , \new_[18360]_ , \new_[18363]_ ,
    \new_[18367]_ , \new_[18368]_ , \new_[18369]_ , \new_[18373]_ ,
    \new_[18374]_ , \new_[18378]_ , \new_[18379]_ , \new_[18380]_ ,
    \new_[18383]_ , \new_[18387]_ , \new_[18388]_ , \new_[18389]_ ,
    \new_[18393]_ , \new_[18394]_ , \new_[18398]_ , \new_[18399]_ ,
    \new_[18400]_ , \new_[18403]_ , \new_[18407]_ , \new_[18408]_ ,
    \new_[18409]_ , \new_[18413]_ , \new_[18414]_ , \new_[18418]_ ,
    \new_[18419]_ , \new_[18420]_ , \new_[18423]_ , \new_[18427]_ ,
    \new_[18428]_ , \new_[18429]_ , \new_[18433]_ , \new_[18434]_ ,
    \new_[18438]_ , \new_[18439]_ , \new_[18440]_ , \new_[18443]_ ,
    \new_[18447]_ , \new_[18448]_ , \new_[18449]_ , \new_[18453]_ ,
    \new_[18454]_ , \new_[18458]_ , \new_[18459]_ , \new_[18460]_ ,
    \new_[18463]_ , \new_[18467]_ , \new_[18468]_ , \new_[18469]_ ,
    \new_[18473]_ , \new_[18474]_ , \new_[18478]_ , \new_[18479]_ ,
    \new_[18480]_ , \new_[18483]_ , \new_[18487]_ , \new_[18488]_ ,
    \new_[18489]_ , \new_[18493]_ , \new_[18494]_ , \new_[18498]_ ,
    \new_[18499]_ , \new_[18500]_ , \new_[18503]_ , \new_[18507]_ ,
    \new_[18508]_ , \new_[18509]_ , \new_[18513]_ , \new_[18514]_ ,
    \new_[18518]_ , \new_[18519]_ , \new_[18520]_ , \new_[18523]_ ,
    \new_[18527]_ , \new_[18528]_ , \new_[18529]_ , \new_[18533]_ ,
    \new_[18534]_ , \new_[18538]_ , \new_[18539]_ , \new_[18540]_ ,
    \new_[18543]_ , \new_[18547]_ , \new_[18548]_ , \new_[18549]_ ,
    \new_[18553]_ , \new_[18554]_ , \new_[18558]_ , \new_[18559]_ ,
    \new_[18560]_ , \new_[18563]_ , \new_[18567]_ , \new_[18568]_ ,
    \new_[18569]_ , \new_[18573]_ , \new_[18574]_ , \new_[18578]_ ,
    \new_[18579]_ , \new_[18580]_ , \new_[18583]_ , \new_[18587]_ ,
    \new_[18588]_ , \new_[18589]_ , \new_[18593]_ , \new_[18594]_ ,
    \new_[18598]_ , \new_[18599]_ , \new_[18600]_ , \new_[18603]_ ,
    \new_[18607]_ , \new_[18608]_ , \new_[18609]_ , \new_[18613]_ ,
    \new_[18614]_ , \new_[18618]_ , \new_[18619]_ , \new_[18620]_ ,
    \new_[18623]_ , \new_[18627]_ , \new_[18628]_ , \new_[18629]_ ,
    \new_[18633]_ , \new_[18634]_ , \new_[18638]_ , \new_[18639]_ ,
    \new_[18640]_ , \new_[18643]_ , \new_[18647]_ , \new_[18648]_ ,
    \new_[18649]_ , \new_[18653]_ , \new_[18654]_ , \new_[18658]_ ,
    \new_[18659]_ , \new_[18660]_ , \new_[18663]_ , \new_[18667]_ ,
    \new_[18668]_ , \new_[18669]_ , \new_[18673]_ , \new_[18674]_ ,
    \new_[18678]_ , \new_[18679]_ , \new_[18680]_ , \new_[18683]_ ,
    \new_[18687]_ , \new_[18688]_ , \new_[18689]_ , \new_[18693]_ ,
    \new_[18694]_ , \new_[18698]_ , \new_[18699]_ , \new_[18700]_ ,
    \new_[18703]_ , \new_[18707]_ , \new_[18708]_ , \new_[18709]_ ,
    \new_[18713]_ , \new_[18714]_ , \new_[18718]_ , \new_[18719]_ ,
    \new_[18720]_ , \new_[18723]_ , \new_[18727]_ , \new_[18728]_ ,
    \new_[18729]_ , \new_[18733]_ , \new_[18734]_ , \new_[18738]_ ,
    \new_[18739]_ , \new_[18740]_ , \new_[18743]_ , \new_[18747]_ ,
    \new_[18748]_ , \new_[18749]_ , \new_[18753]_ , \new_[18754]_ ,
    \new_[18758]_ , \new_[18759]_ , \new_[18760]_ , \new_[18763]_ ,
    \new_[18767]_ , \new_[18768]_ , \new_[18769]_ , \new_[18773]_ ,
    \new_[18774]_ , \new_[18778]_ , \new_[18779]_ , \new_[18780]_ ,
    \new_[18783]_ , \new_[18787]_ , \new_[18788]_ , \new_[18789]_ ,
    \new_[18793]_ , \new_[18794]_ , \new_[18798]_ , \new_[18799]_ ,
    \new_[18800]_ , \new_[18803]_ , \new_[18807]_ , \new_[18808]_ ,
    \new_[18809]_ , \new_[18813]_ , \new_[18814]_ , \new_[18818]_ ,
    \new_[18819]_ , \new_[18820]_ , \new_[18823]_ , \new_[18827]_ ,
    \new_[18828]_ , \new_[18829]_ , \new_[18833]_ , \new_[18834]_ ,
    \new_[18838]_ , \new_[18839]_ , \new_[18840]_ , \new_[18843]_ ,
    \new_[18847]_ , \new_[18848]_ , \new_[18849]_ , \new_[18853]_ ,
    \new_[18854]_ , \new_[18858]_ , \new_[18859]_ , \new_[18860]_ ,
    \new_[18863]_ , \new_[18867]_ , \new_[18868]_ , \new_[18869]_ ,
    \new_[18873]_ , \new_[18874]_ , \new_[18878]_ , \new_[18879]_ ,
    \new_[18880]_ , \new_[18883]_ , \new_[18887]_ , \new_[18888]_ ,
    \new_[18889]_ , \new_[18893]_ , \new_[18894]_ , \new_[18898]_ ,
    \new_[18899]_ , \new_[18900]_ , \new_[18903]_ , \new_[18907]_ ,
    \new_[18908]_ , \new_[18909]_ , \new_[18913]_ , \new_[18914]_ ,
    \new_[18918]_ , \new_[18919]_ , \new_[18920]_ , \new_[18923]_ ,
    \new_[18927]_ , \new_[18928]_ , \new_[18929]_ , \new_[18933]_ ,
    \new_[18934]_ , \new_[18938]_ , \new_[18939]_ , \new_[18940]_ ,
    \new_[18943]_ , \new_[18947]_ , \new_[18948]_ , \new_[18949]_ ,
    \new_[18953]_ , \new_[18954]_ , \new_[18958]_ , \new_[18959]_ ,
    \new_[18960]_ , \new_[18963]_ , \new_[18967]_ , \new_[18968]_ ,
    \new_[18969]_ , \new_[18973]_ , \new_[18974]_ , \new_[18978]_ ,
    \new_[18979]_ , \new_[18980]_ , \new_[18983]_ , \new_[18987]_ ,
    \new_[18988]_ , \new_[18989]_ , \new_[18993]_ , \new_[18994]_ ,
    \new_[18998]_ , \new_[18999]_ , \new_[19000]_ , \new_[19003]_ ,
    \new_[19007]_ , \new_[19008]_ , \new_[19009]_ , \new_[19013]_ ,
    \new_[19014]_ , \new_[19018]_ , \new_[19019]_ , \new_[19020]_ ,
    \new_[19023]_ , \new_[19027]_ , \new_[19028]_ , \new_[19029]_ ,
    \new_[19033]_ , \new_[19034]_ , \new_[19038]_ , \new_[19039]_ ,
    \new_[19040]_ , \new_[19043]_ , \new_[19047]_ , \new_[19048]_ ,
    \new_[19049]_ , \new_[19053]_ , \new_[19054]_ , \new_[19058]_ ,
    \new_[19059]_ , \new_[19060]_ , \new_[19063]_ , \new_[19067]_ ,
    \new_[19068]_ , \new_[19069]_ , \new_[19073]_ , \new_[19074]_ ,
    \new_[19078]_ , \new_[19079]_ , \new_[19080]_ , \new_[19083]_ ,
    \new_[19087]_ , \new_[19088]_ , \new_[19089]_ , \new_[19093]_ ,
    \new_[19094]_ , \new_[19098]_ , \new_[19099]_ , \new_[19100]_ ,
    \new_[19103]_ , \new_[19107]_ , \new_[19108]_ , \new_[19109]_ ,
    \new_[19113]_ , \new_[19114]_ , \new_[19118]_ , \new_[19119]_ ,
    \new_[19120]_ , \new_[19123]_ , \new_[19127]_ , \new_[19128]_ ,
    \new_[19129]_ , \new_[19133]_ , \new_[19134]_ , \new_[19138]_ ,
    \new_[19139]_ , \new_[19140]_ , \new_[19143]_ , \new_[19147]_ ,
    \new_[19148]_ , \new_[19149]_ , \new_[19153]_ , \new_[19154]_ ,
    \new_[19158]_ , \new_[19159]_ , \new_[19160]_ , \new_[19163]_ ,
    \new_[19167]_ , \new_[19168]_ , \new_[19169]_ , \new_[19173]_ ,
    \new_[19174]_ , \new_[19178]_ , \new_[19179]_ , \new_[19180]_ ,
    \new_[19183]_ , \new_[19187]_ , \new_[19188]_ , \new_[19189]_ ,
    \new_[19193]_ , \new_[19194]_ , \new_[19198]_ , \new_[19199]_ ,
    \new_[19200]_ , \new_[19203]_ , \new_[19207]_ , \new_[19208]_ ,
    \new_[19209]_ , \new_[19213]_ , \new_[19214]_ , \new_[19218]_ ,
    \new_[19219]_ , \new_[19220]_ , \new_[19223]_ , \new_[19227]_ ,
    \new_[19228]_ , \new_[19229]_ , \new_[19233]_ , \new_[19234]_ ,
    \new_[19238]_ , \new_[19239]_ , \new_[19240]_ , \new_[19243]_ ,
    \new_[19247]_ , \new_[19248]_ , \new_[19249]_ , \new_[19253]_ ,
    \new_[19254]_ , \new_[19258]_ , \new_[19259]_ , \new_[19260]_ ,
    \new_[19263]_ , \new_[19267]_ , \new_[19268]_ , \new_[19269]_ ,
    \new_[19273]_ , \new_[19274]_ , \new_[19278]_ , \new_[19279]_ ,
    \new_[19280]_ , \new_[19283]_ , \new_[19287]_ , \new_[19288]_ ,
    \new_[19289]_ , \new_[19293]_ , \new_[19294]_ , \new_[19298]_ ,
    \new_[19299]_ , \new_[19300]_ , \new_[19303]_ , \new_[19307]_ ,
    \new_[19308]_ , \new_[19309]_ , \new_[19313]_ , \new_[19314]_ ,
    \new_[19318]_ , \new_[19319]_ , \new_[19320]_ , \new_[19323]_ ,
    \new_[19327]_ , \new_[19328]_ , \new_[19329]_ , \new_[19333]_ ,
    \new_[19334]_ , \new_[19338]_ , \new_[19339]_ , \new_[19340]_ ,
    \new_[19343]_ , \new_[19347]_ , \new_[19348]_ , \new_[19349]_ ,
    \new_[19353]_ , \new_[19354]_ , \new_[19358]_ , \new_[19359]_ ,
    \new_[19360]_ , \new_[19363]_ , \new_[19367]_ , \new_[19368]_ ,
    \new_[19369]_ , \new_[19373]_ , \new_[19374]_ , \new_[19378]_ ,
    \new_[19379]_ , \new_[19380]_ , \new_[19383]_ , \new_[19387]_ ,
    \new_[19388]_ , \new_[19389]_ , \new_[19393]_ , \new_[19394]_ ,
    \new_[19398]_ , \new_[19399]_ , \new_[19400]_ , \new_[19403]_ ,
    \new_[19407]_ , \new_[19408]_ , \new_[19409]_ , \new_[19413]_ ,
    \new_[19414]_ , \new_[19418]_ , \new_[19419]_ , \new_[19420]_ ,
    \new_[19423]_ , \new_[19427]_ , \new_[19428]_ , \new_[19429]_ ,
    \new_[19433]_ , \new_[19434]_ , \new_[19438]_ , \new_[19439]_ ,
    \new_[19440]_ , \new_[19443]_ , \new_[19447]_ , \new_[19448]_ ,
    \new_[19449]_ , \new_[19453]_ , \new_[19454]_ , \new_[19458]_ ,
    \new_[19459]_ , \new_[19460]_ , \new_[19463]_ , \new_[19467]_ ,
    \new_[19468]_ , \new_[19469]_ , \new_[19473]_ , \new_[19474]_ ,
    \new_[19478]_ , \new_[19479]_ , \new_[19480]_ , \new_[19483]_ ,
    \new_[19487]_ , \new_[19488]_ , \new_[19489]_ , \new_[19493]_ ,
    \new_[19494]_ , \new_[19498]_ , \new_[19499]_ , \new_[19500]_ ,
    \new_[19503]_ , \new_[19507]_ , \new_[19508]_ , \new_[19509]_ ,
    \new_[19513]_ , \new_[19514]_ , \new_[19518]_ , \new_[19519]_ ,
    \new_[19520]_ , \new_[19523]_ , \new_[19527]_ , \new_[19528]_ ,
    \new_[19529]_ , \new_[19533]_ , \new_[19534]_ , \new_[19538]_ ,
    \new_[19539]_ , \new_[19540]_ , \new_[19543]_ , \new_[19547]_ ,
    \new_[19548]_ , \new_[19549]_ , \new_[19553]_ , \new_[19554]_ ,
    \new_[19558]_ , \new_[19559]_ , \new_[19560]_ , \new_[19563]_ ,
    \new_[19567]_ , \new_[19568]_ , \new_[19569]_ , \new_[19573]_ ,
    \new_[19574]_ , \new_[19578]_ , \new_[19579]_ , \new_[19580]_ ,
    \new_[19583]_ , \new_[19587]_ , \new_[19588]_ , \new_[19589]_ ,
    \new_[19593]_ , \new_[19594]_ , \new_[19598]_ , \new_[19599]_ ,
    \new_[19600]_ , \new_[19603]_ , \new_[19607]_ , \new_[19608]_ ,
    \new_[19609]_ , \new_[19613]_ , \new_[19614]_ , \new_[19618]_ ,
    \new_[19619]_ , \new_[19620]_ , \new_[19623]_ , \new_[19627]_ ,
    \new_[19628]_ , \new_[19629]_ , \new_[19633]_ , \new_[19634]_ ,
    \new_[19638]_ , \new_[19639]_ , \new_[19640]_ , \new_[19643]_ ,
    \new_[19647]_ , \new_[19648]_ , \new_[19649]_ , \new_[19653]_ ,
    \new_[19654]_ , \new_[19658]_ , \new_[19659]_ , \new_[19660]_ ,
    \new_[19663]_ , \new_[19667]_ , \new_[19668]_ , \new_[19669]_ ,
    \new_[19673]_ , \new_[19674]_ , \new_[19678]_ , \new_[19679]_ ,
    \new_[19680]_ , \new_[19683]_ , \new_[19687]_ , \new_[19688]_ ,
    \new_[19689]_ , \new_[19693]_ , \new_[19694]_ , \new_[19698]_ ,
    \new_[19699]_ , \new_[19700]_ , \new_[19703]_ , \new_[19707]_ ,
    \new_[19708]_ , \new_[19709]_ , \new_[19713]_ , \new_[19714]_ ,
    \new_[19718]_ , \new_[19719]_ , \new_[19720]_ , \new_[19723]_ ,
    \new_[19727]_ , \new_[19728]_ , \new_[19729]_ , \new_[19733]_ ,
    \new_[19734]_ , \new_[19738]_ , \new_[19739]_ , \new_[19740]_ ,
    \new_[19743]_ , \new_[19747]_ , \new_[19748]_ , \new_[19749]_ ,
    \new_[19753]_ , \new_[19754]_ , \new_[19758]_ , \new_[19759]_ ,
    \new_[19760]_ , \new_[19763]_ , \new_[19767]_ , \new_[19768]_ ,
    \new_[19769]_ , \new_[19773]_ , \new_[19774]_ , \new_[19778]_ ,
    \new_[19779]_ , \new_[19780]_ , \new_[19783]_ , \new_[19787]_ ,
    \new_[19788]_ , \new_[19789]_ , \new_[19793]_ , \new_[19794]_ ,
    \new_[19798]_ , \new_[19799]_ , \new_[19800]_ , \new_[19803]_ ,
    \new_[19807]_ , \new_[19808]_ , \new_[19809]_ , \new_[19813]_ ,
    \new_[19814]_ , \new_[19818]_ , \new_[19819]_ , \new_[19820]_ ,
    \new_[19823]_ , \new_[19827]_ , \new_[19828]_ , \new_[19829]_ ,
    \new_[19833]_ , \new_[19834]_ , \new_[19838]_ , \new_[19839]_ ,
    \new_[19840]_ , \new_[19843]_ , \new_[19847]_ , \new_[19848]_ ,
    \new_[19849]_ , \new_[19853]_ , \new_[19854]_ , \new_[19858]_ ,
    \new_[19859]_ , \new_[19860]_ , \new_[19863]_ , \new_[19867]_ ,
    \new_[19868]_ , \new_[19869]_ , \new_[19873]_ , \new_[19874]_ ,
    \new_[19878]_ , \new_[19879]_ , \new_[19880]_ , \new_[19883]_ ,
    \new_[19887]_ , \new_[19888]_ , \new_[19889]_ , \new_[19893]_ ,
    \new_[19894]_ , \new_[19898]_ , \new_[19899]_ , \new_[19900]_ ,
    \new_[19903]_ , \new_[19907]_ , \new_[19908]_ , \new_[19909]_ ,
    \new_[19913]_ , \new_[19914]_ , \new_[19918]_ , \new_[19919]_ ,
    \new_[19920]_ , \new_[19923]_ , \new_[19927]_ , \new_[19928]_ ,
    \new_[19929]_ , \new_[19933]_ , \new_[19934]_ , \new_[19938]_ ,
    \new_[19939]_ , \new_[19940]_ , \new_[19943]_ , \new_[19947]_ ,
    \new_[19948]_ , \new_[19949]_ , \new_[19953]_ , \new_[19954]_ ,
    \new_[19958]_ , \new_[19959]_ , \new_[19960]_ , \new_[19963]_ ,
    \new_[19967]_ , \new_[19968]_ , \new_[19969]_ , \new_[19973]_ ,
    \new_[19974]_ , \new_[19978]_ , \new_[19979]_ , \new_[19980]_ ,
    \new_[19983]_ , \new_[19987]_ , \new_[19988]_ , \new_[19989]_ ,
    \new_[19993]_ , \new_[19994]_ , \new_[19998]_ , \new_[19999]_ ,
    \new_[20000]_ , \new_[20003]_ , \new_[20007]_ , \new_[20008]_ ,
    \new_[20009]_ , \new_[20013]_ , \new_[20014]_ , \new_[20018]_ ,
    \new_[20019]_ , \new_[20020]_ , \new_[20023]_ , \new_[20027]_ ,
    \new_[20028]_ , \new_[20029]_ , \new_[20033]_ , \new_[20034]_ ,
    \new_[20038]_ , \new_[20039]_ , \new_[20040]_ , \new_[20043]_ ,
    \new_[20047]_ , \new_[20048]_ , \new_[20049]_ , \new_[20053]_ ,
    \new_[20054]_ , \new_[20058]_ , \new_[20059]_ , \new_[20060]_ ,
    \new_[20063]_ , \new_[20067]_ , \new_[20068]_ , \new_[20069]_ ,
    \new_[20073]_ , \new_[20074]_ , \new_[20078]_ , \new_[20079]_ ,
    \new_[20080]_ , \new_[20083]_ , \new_[20087]_ , \new_[20088]_ ,
    \new_[20089]_ , \new_[20093]_ , \new_[20094]_ , \new_[20098]_ ,
    \new_[20099]_ , \new_[20100]_ , \new_[20103]_ , \new_[20107]_ ,
    \new_[20108]_ , \new_[20109]_ , \new_[20113]_ , \new_[20114]_ ,
    \new_[20118]_ , \new_[20119]_ , \new_[20120]_ , \new_[20123]_ ,
    \new_[20127]_ , \new_[20128]_ , \new_[20129]_ , \new_[20133]_ ,
    \new_[20134]_ , \new_[20138]_ , \new_[20139]_ , \new_[20140]_ ,
    \new_[20143]_ , \new_[20147]_ , \new_[20148]_ , \new_[20149]_ ,
    \new_[20153]_ , \new_[20154]_ , \new_[20158]_ , \new_[20159]_ ,
    \new_[20160]_ , \new_[20163]_ , \new_[20167]_ , \new_[20168]_ ,
    \new_[20169]_ , \new_[20173]_ , \new_[20174]_ , \new_[20178]_ ,
    \new_[20179]_ , \new_[20180]_ , \new_[20183]_ , \new_[20187]_ ,
    \new_[20188]_ , \new_[20189]_ , \new_[20193]_ , \new_[20194]_ ,
    \new_[20198]_ , \new_[20199]_ , \new_[20200]_ , \new_[20203]_ ,
    \new_[20207]_ , \new_[20208]_ , \new_[20209]_ , \new_[20213]_ ,
    \new_[20214]_ , \new_[20218]_ , \new_[20219]_ , \new_[20220]_ ,
    \new_[20223]_ , \new_[20227]_ , \new_[20228]_ , \new_[20229]_ ,
    \new_[20233]_ , \new_[20234]_ , \new_[20238]_ , \new_[20239]_ ,
    \new_[20240]_ , \new_[20243]_ , \new_[20247]_ , \new_[20248]_ ,
    \new_[20249]_ , \new_[20253]_ , \new_[20254]_ , \new_[20258]_ ,
    \new_[20259]_ , \new_[20260]_ , \new_[20263]_ , \new_[20267]_ ,
    \new_[20268]_ , \new_[20269]_ , \new_[20273]_ , \new_[20274]_ ,
    \new_[20278]_ , \new_[20279]_ , \new_[20280]_ , \new_[20283]_ ,
    \new_[20287]_ , \new_[20288]_ , \new_[20289]_ , \new_[20293]_ ,
    \new_[20294]_ , \new_[20298]_ , \new_[20299]_ , \new_[20300]_ ,
    \new_[20303]_ , \new_[20307]_ , \new_[20308]_ , \new_[20309]_ ,
    \new_[20313]_ , \new_[20314]_ , \new_[20318]_ , \new_[20319]_ ,
    \new_[20320]_ , \new_[20323]_ , \new_[20327]_ , \new_[20328]_ ,
    \new_[20329]_ , \new_[20333]_ , \new_[20334]_ , \new_[20338]_ ,
    \new_[20339]_ , \new_[20340]_ , \new_[20343]_ , \new_[20347]_ ,
    \new_[20348]_ , \new_[20349]_ , \new_[20353]_ , \new_[20354]_ ,
    \new_[20358]_ , \new_[20359]_ , \new_[20360]_ , \new_[20363]_ ,
    \new_[20367]_ , \new_[20368]_ , \new_[20369]_ , \new_[20373]_ ,
    \new_[20374]_ , \new_[20378]_ , \new_[20379]_ , \new_[20380]_ ,
    \new_[20383]_ , \new_[20387]_ , \new_[20388]_ , \new_[20389]_ ,
    \new_[20393]_ , \new_[20394]_ , \new_[20398]_ , \new_[20399]_ ,
    \new_[20400]_ , \new_[20403]_ , \new_[20407]_ , \new_[20408]_ ,
    \new_[20409]_ , \new_[20413]_ , \new_[20414]_ , \new_[20418]_ ,
    \new_[20419]_ , \new_[20420]_ , \new_[20423]_ , \new_[20427]_ ,
    \new_[20428]_ , \new_[20429]_ , \new_[20433]_ , \new_[20434]_ ,
    \new_[20438]_ , \new_[20439]_ , \new_[20440]_ , \new_[20443]_ ,
    \new_[20447]_ , \new_[20448]_ , \new_[20449]_ , \new_[20453]_ ,
    \new_[20454]_ , \new_[20458]_ , \new_[20459]_ , \new_[20460]_ ,
    \new_[20463]_ , \new_[20467]_ , \new_[20468]_ , \new_[20469]_ ,
    \new_[20473]_ , \new_[20474]_ , \new_[20478]_ , \new_[20479]_ ,
    \new_[20480]_ , \new_[20483]_ , \new_[20487]_ , \new_[20488]_ ,
    \new_[20489]_ , \new_[20493]_ , \new_[20494]_ , \new_[20498]_ ,
    \new_[20499]_ , \new_[20500]_ , \new_[20503]_ , \new_[20507]_ ,
    \new_[20508]_ , \new_[20509]_ , \new_[20513]_ , \new_[20514]_ ,
    \new_[20518]_ , \new_[20519]_ , \new_[20520]_ , \new_[20523]_ ,
    \new_[20527]_ , \new_[20528]_ , \new_[20529]_ , \new_[20533]_ ,
    \new_[20534]_ , \new_[20538]_ , \new_[20539]_ , \new_[20540]_ ,
    \new_[20543]_ , \new_[20547]_ , \new_[20548]_ , \new_[20549]_ ,
    \new_[20553]_ , \new_[20554]_ , \new_[20558]_ , \new_[20559]_ ,
    \new_[20560]_ , \new_[20563]_ , \new_[20567]_ , \new_[20568]_ ,
    \new_[20569]_ , \new_[20573]_ , \new_[20574]_ , \new_[20578]_ ,
    \new_[20579]_ , \new_[20580]_ , \new_[20583]_ , \new_[20587]_ ,
    \new_[20588]_ , \new_[20589]_ , \new_[20593]_ , \new_[20594]_ ,
    \new_[20598]_ , \new_[20599]_ , \new_[20600]_ , \new_[20603]_ ,
    \new_[20607]_ , \new_[20608]_ , \new_[20609]_ , \new_[20613]_ ,
    \new_[20614]_ , \new_[20618]_ , \new_[20619]_ , \new_[20620]_ ,
    \new_[20623]_ , \new_[20627]_ , \new_[20628]_ , \new_[20629]_ ,
    \new_[20633]_ , \new_[20634]_ , \new_[20638]_ , \new_[20639]_ ,
    \new_[20640]_ , \new_[20643]_ , \new_[20647]_ , \new_[20648]_ ,
    \new_[20649]_ , \new_[20653]_ , \new_[20654]_ , \new_[20658]_ ,
    \new_[20659]_ , \new_[20660]_ , \new_[20663]_ , \new_[20667]_ ,
    \new_[20668]_ , \new_[20669]_ , \new_[20673]_ , \new_[20674]_ ,
    \new_[20678]_ , \new_[20679]_ , \new_[20680]_ , \new_[20683]_ ,
    \new_[20687]_ , \new_[20688]_ , \new_[20689]_ , \new_[20693]_ ,
    \new_[20694]_ , \new_[20698]_ , \new_[20699]_ , \new_[20700]_ ,
    \new_[20703]_ , \new_[20707]_ , \new_[20708]_ , \new_[20709]_ ,
    \new_[20713]_ , \new_[20714]_ , \new_[20718]_ , \new_[20719]_ ,
    \new_[20720]_ , \new_[20723]_ , \new_[20727]_ , \new_[20728]_ ,
    \new_[20729]_ , \new_[20733]_ , \new_[20734]_ , \new_[20738]_ ,
    \new_[20739]_ , \new_[20740]_ , \new_[20743]_ , \new_[20747]_ ,
    \new_[20748]_ , \new_[20749]_ , \new_[20753]_ , \new_[20754]_ ,
    \new_[20758]_ , \new_[20759]_ , \new_[20760]_ , \new_[20763]_ ,
    \new_[20767]_ , \new_[20768]_ , \new_[20769]_ , \new_[20773]_ ,
    \new_[20774]_ , \new_[20778]_ , \new_[20779]_ , \new_[20780]_ ,
    \new_[20783]_ , \new_[20787]_ , \new_[20788]_ , \new_[20789]_ ,
    \new_[20793]_ , \new_[20794]_ , \new_[20798]_ , \new_[20799]_ ,
    \new_[20800]_ , \new_[20803]_ , \new_[20807]_ , \new_[20808]_ ,
    \new_[20809]_ , \new_[20813]_ , \new_[20814]_ , \new_[20818]_ ,
    \new_[20819]_ , \new_[20820]_ , \new_[20823]_ , \new_[20827]_ ,
    \new_[20828]_ , \new_[20829]_ , \new_[20833]_ , \new_[20834]_ ,
    \new_[20838]_ , \new_[20839]_ , \new_[20840]_ , \new_[20843]_ ,
    \new_[20847]_ , \new_[20848]_ , \new_[20849]_ , \new_[20853]_ ,
    \new_[20854]_ , \new_[20858]_ , \new_[20859]_ , \new_[20860]_ ,
    \new_[20863]_ , \new_[20867]_ , \new_[20868]_ , \new_[20869]_ ,
    \new_[20873]_ , \new_[20874]_ , \new_[20878]_ , \new_[20879]_ ,
    \new_[20880]_ , \new_[20883]_ , \new_[20887]_ , \new_[20888]_ ,
    \new_[20889]_ , \new_[20893]_ , \new_[20894]_ , \new_[20898]_ ,
    \new_[20899]_ , \new_[20900]_ , \new_[20903]_ , \new_[20907]_ ,
    \new_[20908]_ , \new_[20909]_ , \new_[20913]_ , \new_[20914]_ ,
    \new_[20918]_ , \new_[20919]_ , \new_[20920]_ , \new_[20923]_ ,
    \new_[20927]_ , \new_[20928]_ , \new_[20929]_ , \new_[20933]_ ,
    \new_[20934]_ , \new_[20938]_ , \new_[20939]_ , \new_[20940]_ ,
    \new_[20943]_ , \new_[20947]_ , \new_[20948]_ , \new_[20949]_ ,
    \new_[20953]_ , \new_[20954]_ , \new_[20958]_ , \new_[20959]_ ,
    \new_[20960]_ , \new_[20963]_ , \new_[20967]_ , \new_[20968]_ ,
    \new_[20969]_ , \new_[20973]_ , \new_[20974]_ , \new_[20978]_ ,
    \new_[20979]_ , \new_[20980]_ , \new_[20983]_ , \new_[20987]_ ,
    \new_[20988]_ , \new_[20989]_ , \new_[20993]_ , \new_[20994]_ ,
    \new_[20998]_ , \new_[20999]_ , \new_[21000]_ , \new_[21003]_ ,
    \new_[21007]_ , \new_[21008]_ , \new_[21009]_ , \new_[21013]_ ,
    \new_[21014]_ , \new_[21018]_ , \new_[21019]_ , \new_[21020]_ ,
    \new_[21023]_ , \new_[21027]_ , \new_[21028]_ , \new_[21029]_ ,
    \new_[21033]_ , \new_[21034]_ , \new_[21038]_ , \new_[21039]_ ,
    \new_[21040]_ , \new_[21043]_ , \new_[21047]_ , \new_[21048]_ ,
    \new_[21049]_ , \new_[21053]_ , \new_[21054]_ , \new_[21058]_ ,
    \new_[21059]_ , \new_[21060]_ , \new_[21063]_ , \new_[21067]_ ,
    \new_[21068]_ , \new_[21069]_ , \new_[21073]_ , \new_[21074]_ ,
    \new_[21078]_ , \new_[21079]_ , \new_[21080]_ , \new_[21083]_ ,
    \new_[21087]_ , \new_[21088]_ , \new_[21089]_ , \new_[21093]_ ,
    \new_[21094]_ , \new_[21098]_ , \new_[21099]_ , \new_[21100]_ ,
    \new_[21103]_ , \new_[21107]_ , \new_[21108]_ , \new_[21109]_ ,
    \new_[21113]_ , \new_[21114]_ , \new_[21118]_ , \new_[21119]_ ,
    \new_[21120]_ , \new_[21123]_ , \new_[21127]_ , \new_[21128]_ ,
    \new_[21129]_ , \new_[21133]_ , \new_[21134]_ , \new_[21138]_ ,
    \new_[21139]_ , \new_[21140]_ , \new_[21143]_ , \new_[21147]_ ,
    \new_[21148]_ , \new_[21149]_ , \new_[21153]_ , \new_[21154]_ ,
    \new_[21158]_ , \new_[21159]_ , \new_[21160]_ , \new_[21163]_ ,
    \new_[21167]_ , \new_[21168]_ , \new_[21169]_ , \new_[21173]_ ,
    \new_[21174]_ , \new_[21178]_ , \new_[21179]_ , \new_[21180]_ ,
    \new_[21183]_ , \new_[21187]_ , \new_[21188]_ , \new_[21189]_ ,
    \new_[21193]_ , \new_[21194]_ , \new_[21198]_ , \new_[21199]_ ,
    \new_[21200]_ , \new_[21203]_ , \new_[21207]_ , \new_[21208]_ ,
    \new_[21209]_ , \new_[21213]_ , \new_[21214]_ , \new_[21218]_ ,
    \new_[21219]_ , \new_[21220]_ , \new_[21223]_ , \new_[21227]_ ,
    \new_[21228]_ , \new_[21229]_ , \new_[21233]_ , \new_[21234]_ ,
    \new_[21238]_ , \new_[21239]_ , \new_[21240]_ , \new_[21243]_ ,
    \new_[21247]_ , \new_[21248]_ , \new_[21249]_ , \new_[21253]_ ,
    \new_[21254]_ , \new_[21258]_ , \new_[21259]_ , \new_[21260]_ ,
    \new_[21263]_ , \new_[21267]_ , \new_[21268]_ , \new_[21269]_ ,
    \new_[21273]_ , \new_[21274]_ , \new_[21278]_ , \new_[21279]_ ,
    \new_[21280]_ , \new_[21283]_ , \new_[21287]_ , \new_[21288]_ ,
    \new_[21289]_ , \new_[21293]_ , \new_[21294]_ , \new_[21298]_ ,
    \new_[21299]_ , \new_[21300]_ , \new_[21303]_ , \new_[21307]_ ,
    \new_[21308]_ , \new_[21309]_ , \new_[21313]_ , \new_[21314]_ ,
    \new_[21318]_ , \new_[21319]_ , \new_[21320]_ , \new_[21323]_ ,
    \new_[21327]_ , \new_[21328]_ , \new_[21329]_ , \new_[21333]_ ,
    \new_[21334]_ , \new_[21338]_ , \new_[21339]_ , \new_[21340]_ ,
    \new_[21343]_ , \new_[21347]_ , \new_[21348]_ , \new_[21349]_ ,
    \new_[21353]_ , \new_[21354]_ , \new_[21358]_ , \new_[21359]_ ,
    \new_[21360]_ , \new_[21363]_ , \new_[21367]_ , \new_[21368]_ ,
    \new_[21369]_ , \new_[21373]_ , \new_[21374]_ , \new_[21378]_ ,
    \new_[21379]_ , \new_[21380]_ , \new_[21383]_ , \new_[21387]_ ,
    \new_[21388]_ , \new_[21389]_ , \new_[21393]_ , \new_[21394]_ ,
    \new_[21398]_ , \new_[21399]_ , \new_[21400]_ , \new_[21403]_ ,
    \new_[21407]_ , \new_[21408]_ , \new_[21409]_ , \new_[21413]_ ,
    \new_[21414]_ , \new_[21418]_ , \new_[21419]_ , \new_[21420]_ ,
    \new_[21423]_ , \new_[21427]_ , \new_[21428]_ , \new_[21429]_ ,
    \new_[21433]_ , \new_[21434]_ , \new_[21438]_ , \new_[21439]_ ,
    \new_[21440]_ , \new_[21443]_ , \new_[21447]_ , \new_[21448]_ ,
    \new_[21449]_ , \new_[21453]_ , \new_[21454]_ , \new_[21458]_ ,
    \new_[21459]_ , \new_[21460]_ , \new_[21463]_ , \new_[21467]_ ,
    \new_[21468]_ , \new_[21469]_ , \new_[21473]_ , \new_[21474]_ ,
    \new_[21478]_ , \new_[21479]_ , \new_[21480]_ , \new_[21483]_ ,
    \new_[21487]_ , \new_[21488]_ , \new_[21489]_ , \new_[21493]_ ,
    \new_[21494]_ , \new_[21498]_ , \new_[21499]_ , \new_[21500]_ ,
    \new_[21503]_ , \new_[21507]_ , \new_[21508]_ , \new_[21509]_ ,
    \new_[21513]_ , \new_[21514]_ , \new_[21518]_ , \new_[21519]_ ,
    \new_[21520]_ , \new_[21523]_ , \new_[21527]_ , \new_[21528]_ ,
    \new_[21529]_ , \new_[21533]_ , \new_[21534]_ , \new_[21538]_ ,
    \new_[21539]_ , \new_[21540]_ , \new_[21543]_ , \new_[21547]_ ,
    \new_[21548]_ , \new_[21549]_ , \new_[21553]_ , \new_[21554]_ ,
    \new_[21558]_ , \new_[21559]_ , \new_[21560]_ , \new_[21563]_ ,
    \new_[21567]_ , \new_[21568]_ , \new_[21569]_ , \new_[21573]_ ,
    \new_[21574]_ , \new_[21578]_ , \new_[21579]_ , \new_[21580]_ ,
    \new_[21583]_ , \new_[21587]_ , \new_[21588]_ , \new_[21589]_ ,
    \new_[21593]_ , \new_[21594]_ , \new_[21598]_ , \new_[21599]_ ,
    \new_[21600]_ , \new_[21603]_ , \new_[21607]_ , \new_[21608]_ ,
    \new_[21609]_ , \new_[21613]_ , \new_[21614]_ , \new_[21618]_ ,
    \new_[21619]_ , \new_[21620]_ , \new_[21623]_ , \new_[21627]_ ,
    \new_[21628]_ , \new_[21629]_ , \new_[21633]_ , \new_[21634]_ ,
    \new_[21638]_ , \new_[21639]_ , \new_[21640]_ , \new_[21643]_ ,
    \new_[21647]_ , \new_[21648]_ , \new_[21649]_ , \new_[21653]_ ,
    \new_[21654]_ , \new_[21658]_ , \new_[21659]_ , \new_[21660]_ ,
    \new_[21663]_ , \new_[21667]_ , \new_[21668]_ , \new_[21669]_ ,
    \new_[21673]_ , \new_[21674]_ , \new_[21678]_ , \new_[21679]_ ,
    \new_[21680]_ , \new_[21683]_ , \new_[21687]_ , \new_[21688]_ ,
    \new_[21689]_ , \new_[21693]_ , \new_[21694]_ , \new_[21698]_ ,
    \new_[21699]_ , \new_[21700]_ , \new_[21703]_ , \new_[21707]_ ,
    \new_[21708]_ , \new_[21709]_ , \new_[21713]_ , \new_[21714]_ ,
    \new_[21718]_ , \new_[21719]_ , \new_[21720]_ , \new_[21723]_ ,
    \new_[21727]_ , \new_[21728]_ , \new_[21729]_ , \new_[21733]_ ,
    \new_[21734]_ , \new_[21738]_ , \new_[21739]_ , \new_[21740]_ ,
    \new_[21743]_ , \new_[21747]_ , \new_[21748]_ , \new_[21749]_ ,
    \new_[21753]_ , \new_[21754]_ , \new_[21758]_ , \new_[21759]_ ,
    \new_[21760]_ , \new_[21763]_ , \new_[21767]_ , \new_[21768]_ ,
    \new_[21769]_ , \new_[21773]_ , \new_[21774]_ , \new_[21778]_ ,
    \new_[21779]_ , \new_[21780]_ , \new_[21783]_ , \new_[21787]_ ,
    \new_[21788]_ , \new_[21789]_ , \new_[21793]_ , \new_[21794]_ ,
    \new_[21798]_ , \new_[21799]_ , \new_[21800]_ , \new_[21803]_ ,
    \new_[21807]_ , \new_[21808]_ , \new_[21809]_ , \new_[21813]_ ,
    \new_[21814]_ , \new_[21818]_ , \new_[21819]_ , \new_[21820]_ ,
    \new_[21823]_ , \new_[21827]_ , \new_[21828]_ , \new_[21829]_ ,
    \new_[21833]_ , \new_[21834]_ , \new_[21838]_ , \new_[21839]_ ,
    \new_[21840]_ , \new_[21843]_ , \new_[21847]_ , \new_[21848]_ ,
    \new_[21849]_ , \new_[21853]_ , \new_[21854]_ , \new_[21858]_ ,
    \new_[21859]_ , \new_[21860]_ , \new_[21863]_ , \new_[21867]_ ,
    \new_[21868]_ , \new_[21869]_ , \new_[21873]_ , \new_[21874]_ ,
    \new_[21878]_ , \new_[21879]_ , \new_[21880]_ , \new_[21883]_ ,
    \new_[21887]_ , \new_[21888]_ , \new_[21889]_ , \new_[21893]_ ,
    \new_[21894]_ , \new_[21898]_ , \new_[21899]_ , \new_[21900]_ ,
    \new_[21903]_ , \new_[21907]_ , \new_[21908]_ , \new_[21909]_ ,
    \new_[21913]_ , \new_[21914]_ , \new_[21918]_ , \new_[21919]_ ,
    \new_[21920]_ , \new_[21923]_ , \new_[21927]_ , \new_[21928]_ ,
    \new_[21929]_ , \new_[21933]_ , \new_[21934]_ , \new_[21938]_ ,
    \new_[21939]_ , \new_[21940]_ , \new_[21943]_ , \new_[21947]_ ,
    \new_[21948]_ , \new_[21949]_ , \new_[21953]_ , \new_[21954]_ ,
    \new_[21958]_ , \new_[21959]_ , \new_[21960]_ , \new_[21963]_ ,
    \new_[21967]_ , \new_[21968]_ , \new_[21969]_ , \new_[21973]_ ,
    \new_[21974]_ , \new_[21978]_ , \new_[21979]_ , \new_[21980]_ ,
    \new_[21983]_ , \new_[21987]_ , \new_[21988]_ , \new_[21989]_ ,
    \new_[21993]_ , \new_[21994]_ , \new_[21998]_ , \new_[21999]_ ,
    \new_[22000]_ , \new_[22003]_ , \new_[22007]_ , \new_[22008]_ ,
    \new_[22009]_ , \new_[22013]_ , \new_[22014]_ , \new_[22018]_ ,
    \new_[22019]_ , \new_[22020]_ , \new_[22023]_ , \new_[22027]_ ,
    \new_[22028]_ , \new_[22029]_ , \new_[22033]_ , \new_[22034]_ ,
    \new_[22038]_ , \new_[22039]_ , \new_[22040]_ , \new_[22043]_ ,
    \new_[22047]_ , \new_[22048]_ , \new_[22049]_ , \new_[22053]_ ,
    \new_[22054]_ , \new_[22058]_ , \new_[22059]_ , \new_[22060]_ ,
    \new_[22063]_ , \new_[22067]_ , \new_[22068]_ , \new_[22069]_ ,
    \new_[22073]_ , \new_[22074]_ , \new_[22078]_ , \new_[22079]_ ,
    \new_[22080]_ , \new_[22083]_ , \new_[22087]_ , \new_[22088]_ ,
    \new_[22089]_ , \new_[22093]_ , \new_[22094]_ , \new_[22098]_ ,
    \new_[22099]_ , \new_[22100]_ , \new_[22103]_ , \new_[22107]_ ,
    \new_[22108]_ , \new_[22109]_ , \new_[22113]_ , \new_[22114]_ ,
    \new_[22118]_ , \new_[22119]_ , \new_[22120]_ , \new_[22123]_ ,
    \new_[22127]_ , \new_[22128]_ , \new_[22129]_ , \new_[22133]_ ,
    \new_[22134]_ , \new_[22138]_ , \new_[22139]_ , \new_[22140]_ ,
    \new_[22143]_ , \new_[22147]_ , \new_[22148]_ , \new_[22149]_ ,
    \new_[22153]_ , \new_[22154]_ , \new_[22158]_ , \new_[22159]_ ,
    \new_[22160]_ , \new_[22163]_ , \new_[22167]_ , \new_[22168]_ ,
    \new_[22169]_ , \new_[22173]_ , \new_[22174]_ , \new_[22178]_ ,
    \new_[22179]_ , \new_[22180]_ , \new_[22183]_ , \new_[22187]_ ,
    \new_[22188]_ , \new_[22189]_ , \new_[22193]_ , \new_[22194]_ ,
    \new_[22198]_ , \new_[22199]_ , \new_[22200]_ , \new_[22203]_ ,
    \new_[22207]_ , \new_[22208]_ , \new_[22209]_ , \new_[22213]_ ,
    \new_[22214]_ , \new_[22218]_ , \new_[22219]_ , \new_[22220]_ ,
    \new_[22223]_ , \new_[22227]_ , \new_[22228]_ , \new_[22229]_ ,
    \new_[22233]_ , \new_[22234]_ , \new_[22238]_ , \new_[22239]_ ,
    \new_[22240]_ , \new_[22243]_ , \new_[22247]_ , \new_[22248]_ ,
    \new_[22249]_ , \new_[22253]_ , \new_[22254]_ , \new_[22258]_ ,
    \new_[22259]_ , \new_[22260]_ , \new_[22263]_ , \new_[22267]_ ,
    \new_[22268]_ , \new_[22269]_ , \new_[22273]_ , \new_[22274]_ ,
    \new_[22278]_ , \new_[22279]_ , \new_[22280]_ , \new_[22283]_ ,
    \new_[22287]_ , \new_[22288]_ , \new_[22289]_ , \new_[22293]_ ,
    \new_[22294]_ , \new_[22298]_ , \new_[22299]_ , \new_[22300]_ ,
    \new_[22303]_ , \new_[22307]_ , \new_[22308]_ , \new_[22309]_ ,
    \new_[22313]_ , \new_[22314]_ , \new_[22318]_ , \new_[22319]_ ,
    \new_[22320]_ , \new_[22323]_ , \new_[22327]_ , \new_[22328]_ ,
    \new_[22329]_ , \new_[22333]_ , \new_[22334]_ , \new_[22338]_ ,
    \new_[22339]_ , \new_[22340]_ , \new_[22343]_ , \new_[22347]_ ,
    \new_[22348]_ , \new_[22349]_ , \new_[22353]_ , \new_[22354]_ ,
    \new_[22358]_ , \new_[22359]_ , \new_[22360]_ , \new_[22363]_ ,
    \new_[22367]_ , \new_[22368]_ , \new_[22369]_ , \new_[22373]_ ,
    \new_[22374]_ , \new_[22378]_ , \new_[22379]_ , \new_[22380]_ ,
    \new_[22383]_ , \new_[22387]_ , \new_[22388]_ , \new_[22389]_ ,
    \new_[22393]_ , \new_[22394]_ , \new_[22398]_ , \new_[22399]_ ,
    \new_[22400]_ , \new_[22403]_ , \new_[22407]_ , \new_[22408]_ ,
    \new_[22409]_ , \new_[22413]_ , \new_[22414]_ , \new_[22418]_ ,
    \new_[22419]_ , \new_[22420]_ , \new_[22423]_ , \new_[22427]_ ,
    \new_[22428]_ , \new_[22429]_ , \new_[22433]_ , \new_[22434]_ ,
    \new_[22438]_ , \new_[22439]_ , \new_[22440]_ , \new_[22443]_ ,
    \new_[22447]_ , \new_[22448]_ , \new_[22449]_ , \new_[22453]_ ,
    \new_[22454]_ , \new_[22458]_ , \new_[22459]_ , \new_[22460]_ ,
    \new_[22463]_ , \new_[22467]_ , \new_[22468]_ , \new_[22469]_ ,
    \new_[22473]_ , \new_[22474]_ , \new_[22478]_ , \new_[22479]_ ,
    \new_[22480]_ , \new_[22483]_ , \new_[22487]_ , \new_[22488]_ ,
    \new_[22489]_ , \new_[22493]_ , \new_[22494]_ , \new_[22498]_ ,
    \new_[22499]_ , \new_[22500]_ , \new_[22503]_ , \new_[22507]_ ,
    \new_[22508]_ , \new_[22509]_ , \new_[22513]_ , \new_[22514]_ ,
    \new_[22518]_ , \new_[22519]_ , \new_[22520]_ , \new_[22523]_ ,
    \new_[22527]_ , \new_[22528]_ , \new_[22529]_ , \new_[22533]_ ,
    \new_[22534]_ , \new_[22538]_ , \new_[22539]_ , \new_[22540]_ ,
    \new_[22543]_ , \new_[22547]_ , \new_[22548]_ , \new_[22549]_ ,
    \new_[22553]_ , \new_[22554]_ , \new_[22558]_ , \new_[22559]_ ,
    \new_[22560]_ , \new_[22563]_ , \new_[22567]_ , \new_[22568]_ ,
    \new_[22569]_ , \new_[22573]_ , \new_[22574]_ , \new_[22578]_ ,
    \new_[22579]_ , \new_[22580]_ , \new_[22583]_ , \new_[22587]_ ,
    \new_[22588]_ , \new_[22589]_ , \new_[22593]_ , \new_[22594]_ ,
    \new_[22598]_ , \new_[22599]_ , \new_[22600]_ , \new_[22603]_ ,
    \new_[22607]_ , \new_[22608]_ , \new_[22609]_ , \new_[22613]_ ,
    \new_[22614]_ , \new_[22618]_ , \new_[22619]_ , \new_[22620]_ ,
    \new_[22623]_ , \new_[22627]_ , \new_[22628]_ , \new_[22629]_ ,
    \new_[22633]_ , \new_[22634]_ , \new_[22638]_ , \new_[22639]_ ,
    \new_[22640]_ , \new_[22643]_ , \new_[22647]_ , \new_[22648]_ ,
    \new_[22649]_ , \new_[22653]_ , \new_[22654]_ , \new_[22658]_ ,
    \new_[22659]_ , \new_[22660]_ , \new_[22663]_ , \new_[22667]_ ,
    \new_[22668]_ , \new_[22669]_ , \new_[22673]_ , \new_[22674]_ ,
    \new_[22678]_ , \new_[22679]_ , \new_[22680]_ , \new_[22683]_ ,
    \new_[22687]_ , \new_[22688]_ , \new_[22689]_ , \new_[22693]_ ,
    \new_[22694]_ , \new_[22698]_ , \new_[22699]_ , \new_[22700]_ ,
    \new_[22703]_ , \new_[22707]_ , \new_[22708]_ , \new_[22709]_ ,
    \new_[22713]_ , \new_[22714]_ , \new_[22718]_ , \new_[22719]_ ,
    \new_[22720]_ , \new_[22723]_ , \new_[22727]_ , \new_[22728]_ ,
    \new_[22729]_ , \new_[22733]_ , \new_[22734]_ , \new_[22738]_ ,
    \new_[22739]_ , \new_[22740]_ , \new_[22743]_ , \new_[22747]_ ,
    \new_[22748]_ , \new_[22749]_ , \new_[22753]_ , \new_[22754]_ ,
    \new_[22758]_ , \new_[22759]_ , \new_[22760]_ , \new_[22763]_ ,
    \new_[22767]_ , \new_[22768]_ , \new_[22769]_ , \new_[22773]_ ,
    \new_[22774]_ , \new_[22778]_ , \new_[22779]_ , \new_[22780]_ ,
    \new_[22783]_ , \new_[22787]_ , \new_[22788]_ , \new_[22789]_ ,
    \new_[22793]_ , \new_[22794]_ , \new_[22798]_ , \new_[22799]_ ,
    \new_[22800]_ , \new_[22803]_ , \new_[22807]_ , \new_[22808]_ ,
    \new_[22809]_ , \new_[22813]_ , \new_[22814]_ , \new_[22818]_ ,
    \new_[22819]_ , \new_[22820]_ , \new_[22823]_ , \new_[22827]_ ,
    \new_[22828]_ , \new_[22829]_ , \new_[22833]_ , \new_[22834]_ ,
    \new_[22838]_ , \new_[22839]_ , \new_[22840]_ , \new_[22843]_ ,
    \new_[22847]_ , \new_[22848]_ , \new_[22849]_ , \new_[22853]_ ,
    \new_[22854]_ , \new_[22858]_ , \new_[22859]_ , \new_[22860]_ ,
    \new_[22863]_ , \new_[22867]_ , \new_[22868]_ , \new_[22869]_ ,
    \new_[22873]_ , \new_[22874]_ , \new_[22878]_ , \new_[22879]_ ,
    \new_[22880]_ , \new_[22883]_ , \new_[22887]_ , \new_[22888]_ ,
    \new_[22889]_ , \new_[22893]_ , \new_[22894]_ , \new_[22898]_ ,
    \new_[22899]_ , \new_[22900]_ , \new_[22903]_ , \new_[22907]_ ,
    \new_[22908]_ , \new_[22909]_ , \new_[22913]_ , \new_[22914]_ ,
    \new_[22918]_ , \new_[22919]_ , \new_[22920]_ , \new_[22923]_ ,
    \new_[22927]_ , \new_[22928]_ , \new_[22929]_ , \new_[22933]_ ,
    \new_[22934]_ , \new_[22938]_ , \new_[22939]_ , \new_[22940]_ ,
    \new_[22943]_ , \new_[22947]_ , \new_[22948]_ , \new_[22949]_ ,
    \new_[22953]_ , \new_[22954]_ , \new_[22958]_ , \new_[22959]_ ,
    \new_[22960]_ , \new_[22963]_ , \new_[22967]_ , \new_[22968]_ ,
    \new_[22969]_ , \new_[22973]_ , \new_[22974]_ , \new_[22978]_ ,
    \new_[22979]_ , \new_[22980]_ , \new_[22983]_ , \new_[22987]_ ,
    \new_[22988]_ , \new_[22989]_ , \new_[22993]_ , \new_[22994]_ ,
    \new_[22998]_ , \new_[22999]_ , \new_[23000]_ , \new_[23003]_ ,
    \new_[23007]_ , \new_[23008]_ , \new_[23009]_ , \new_[23013]_ ,
    \new_[23014]_ , \new_[23018]_ , \new_[23019]_ , \new_[23020]_ ,
    \new_[23023]_ , \new_[23027]_ , \new_[23028]_ , \new_[23029]_ ,
    \new_[23033]_ , \new_[23034]_ , \new_[23038]_ , \new_[23039]_ ,
    \new_[23040]_ , \new_[23043]_ , \new_[23047]_ , \new_[23048]_ ,
    \new_[23049]_ , \new_[23053]_ , \new_[23054]_ , \new_[23058]_ ,
    \new_[23059]_ , \new_[23060]_ , \new_[23063]_ , \new_[23067]_ ,
    \new_[23068]_ , \new_[23069]_ , \new_[23073]_ , \new_[23074]_ ,
    \new_[23078]_ , \new_[23079]_ , \new_[23080]_ , \new_[23083]_ ,
    \new_[23087]_ , \new_[23088]_ , \new_[23089]_ , \new_[23093]_ ,
    \new_[23094]_ , \new_[23098]_ , \new_[23099]_ , \new_[23100]_ ,
    \new_[23103]_ , \new_[23107]_ , \new_[23108]_ , \new_[23109]_ ,
    \new_[23113]_ , \new_[23114]_ , \new_[23118]_ , \new_[23119]_ ,
    \new_[23120]_ , \new_[23123]_ , \new_[23127]_ , \new_[23128]_ ,
    \new_[23129]_ , \new_[23133]_ , \new_[23134]_ , \new_[23138]_ ,
    \new_[23139]_ , \new_[23140]_ , \new_[23143]_ , \new_[23147]_ ,
    \new_[23148]_ , \new_[23149]_ , \new_[23153]_ , \new_[23154]_ ,
    \new_[23158]_ , \new_[23159]_ , \new_[23160]_ , \new_[23163]_ ,
    \new_[23167]_ , \new_[23168]_ , \new_[23169]_ , \new_[23173]_ ,
    \new_[23174]_ , \new_[23178]_ , \new_[23179]_ , \new_[23180]_ ,
    \new_[23183]_ , \new_[23187]_ , \new_[23188]_ , \new_[23189]_ ,
    \new_[23193]_ , \new_[23194]_ , \new_[23198]_ , \new_[23199]_ ,
    \new_[23200]_ , \new_[23203]_ , \new_[23207]_ , \new_[23208]_ ,
    \new_[23209]_ , \new_[23213]_ , \new_[23214]_ , \new_[23218]_ ,
    \new_[23219]_ , \new_[23220]_ , \new_[23223]_ , \new_[23227]_ ,
    \new_[23228]_ , \new_[23229]_ , \new_[23233]_ , \new_[23234]_ ,
    \new_[23238]_ , \new_[23239]_ , \new_[23240]_ , \new_[23243]_ ,
    \new_[23247]_ , \new_[23248]_ , \new_[23249]_ , \new_[23253]_ ,
    \new_[23254]_ , \new_[23258]_ , \new_[23259]_ , \new_[23260]_ ,
    \new_[23263]_ , \new_[23267]_ , \new_[23268]_ , \new_[23269]_ ,
    \new_[23273]_ , \new_[23274]_ , \new_[23278]_ , \new_[23279]_ ,
    \new_[23280]_ , \new_[23283]_ , \new_[23287]_ , \new_[23288]_ ,
    \new_[23289]_ , \new_[23293]_ , \new_[23294]_ , \new_[23298]_ ,
    \new_[23299]_ , \new_[23300]_ , \new_[23303]_ , \new_[23307]_ ,
    \new_[23308]_ , \new_[23309]_ , \new_[23313]_ , \new_[23314]_ ,
    \new_[23318]_ , \new_[23319]_ , \new_[23320]_ , \new_[23323]_ ,
    \new_[23327]_ , \new_[23328]_ , \new_[23329]_ , \new_[23333]_ ,
    \new_[23334]_ , \new_[23338]_ , \new_[23339]_ , \new_[23340]_ ,
    \new_[23343]_ , \new_[23347]_ , \new_[23348]_ , \new_[23349]_ ,
    \new_[23353]_ , \new_[23354]_ , \new_[23358]_ , \new_[23359]_ ,
    \new_[23360]_ , \new_[23363]_ , \new_[23367]_ , \new_[23368]_ ,
    \new_[23369]_ , \new_[23373]_ , \new_[23374]_ , \new_[23378]_ ,
    \new_[23379]_ , \new_[23380]_ , \new_[23383]_ , \new_[23387]_ ,
    \new_[23388]_ , \new_[23389]_ , \new_[23393]_ , \new_[23394]_ ,
    \new_[23398]_ , \new_[23399]_ , \new_[23400]_ , \new_[23403]_ ,
    \new_[23407]_ , \new_[23408]_ , \new_[23409]_ , \new_[23413]_ ,
    \new_[23414]_ , \new_[23418]_ , \new_[23419]_ , \new_[23420]_ ,
    \new_[23423]_ , \new_[23427]_ , \new_[23428]_ , \new_[23429]_ ,
    \new_[23433]_ , \new_[23434]_ , \new_[23438]_ , \new_[23439]_ ,
    \new_[23440]_ , \new_[23443]_ , \new_[23447]_ , \new_[23448]_ ,
    \new_[23449]_ , \new_[23453]_ , \new_[23454]_ , \new_[23458]_ ,
    \new_[23459]_ , \new_[23460]_ , \new_[23463]_ , \new_[23467]_ ,
    \new_[23468]_ , \new_[23469]_ , \new_[23473]_ , \new_[23474]_ ,
    \new_[23478]_ , \new_[23479]_ , \new_[23480]_ , \new_[23483]_ ,
    \new_[23487]_ , \new_[23488]_ , \new_[23489]_ , \new_[23493]_ ,
    \new_[23494]_ , \new_[23498]_ , \new_[23499]_ , \new_[23500]_ ,
    \new_[23503]_ , \new_[23507]_ , \new_[23508]_ , \new_[23509]_ ,
    \new_[23513]_ , \new_[23514]_ , \new_[23518]_ , \new_[23519]_ ,
    \new_[23520]_ , \new_[23523]_ , \new_[23527]_ , \new_[23528]_ ,
    \new_[23529]_ , \new_[23533]_ , \new_[23534]_ , \new_[23538]_ ,
    \new_[23539]_ , \new_[23540]_ , \new_[23543]_ , \new_[23547]_ ,
    \new_[23548]_ , \new_[23549]_ , \new_[23553]_ , \new_[23554]_ ,
    \new_[23558]_ , \new_[23559]_ , \new_[23560]_ , \new_[23563]_ ,
    \new_[23567]_ , \new_[23568]_ , \new_[23569]_ , \new_[23573]_ ,
    \new_[23574]_ , \new_[23578]_ , \new_[23579]_ , \new_[23580]_ ,
    \new_[23583]_ , \new_[23587]_ , \new_[23588]_ , \new_[23589]_ ,
    \new_[23593]_ , \new_[23594]_ , \new_[23598]_ , \new_[23599]_ ,
    \new_[23600]_ , \new_[23603]_ , \new_[23607]_ , \new_[23608]_ ,
    \new_[23609]_ , \new_[23613]_ , \new_[23614]_ , \new_[23618]_ ,
    \new_[23619]_ , \new_[23620]_ , \new_[23623]_ , \new_[23627]_ ,
    \new_[23628]_ , \new_[23629]_ , \new_[23633]_ , \new_[23634]_ ,
    \new_[23638]_ , \new_[23639]_ , \new_[23640]_ , \new_[23643]_ ,
    \new_[23647]_ , \new_[23648]_ , \new_[23649]_ , \new_[23653]_ ,
    \new_[23654]_ , \new_[23658]_ , \new_[23659]_ , \new_[23660]_ ,
    \new_[23663]_ , \new_[23667]_ , \new_[23668]_ , \new_[23669]_ ,
    \new_[23673]_ , \new_[23674]_ , \new_[23678]_ , \new_[23679]_ ,
    \new_[23680]_ , \new_[23683]_ , \new_[23687]_ , \new_[23688]_ ,
    \new_[23689]_ , \new_[23693]_ , \new_[23694]_ , \new_[23698]_ ,
    \new_[23699]_ , \new_[23700]_ , \new_[23703]_ , \new_[23707]_ ,
    \new_[23708]_ , \new_[23709]_ , \new_[23713]_ , \new_[23714]_ ,
    \new_[23718]_ , \new_[23719]_ , \new_[23720]_ , \new_[23723]_ ,
    \new_[23727]_ , \new_[23728]_ , \new_[23729]_ , \new_[23733]_ ,
    \new_[23734]_ , \new_[23738]_ , \new_[23739]_ , \new_[23740]_ ,
    \new_[23743]_ , \new_[23747]_ , \new_[23748]_ , \new_[23749]_ ,
    \new_[23753]_ , \new_[23754]_ , \new_[23758]_ , \new_[23759]_ ,
    \new_[23760]_ , \new_[23763]_ , \new_[23767]_ , \new_[23768]_ ,
    \new_[23769]_ , \new_[23773]_ , \new_[23774]_ , \new_[23778]_ ,
    \new_[23779]_ , \new_[23780]_ , \new_[23783]_ , \new_[23787]_ ,
    \new_[23788]_ , \new_[23789]_ , \new_[23793]_ , \new_[23794]_ ,
    \new_[23798]_ , \new_[23799]_ , \new_[23800]_ , \new_[23803]_ ,
    \new_[23807]_ , \new_[23808]_ , \new_[23809]_ , \new_[23813]_ ,
    \new_[23814]_ , \new_[23818]_ , \new_[23819]_ , \new_[23820]_ ,
    \new_[23823]_ , \new_[23827]_ , \new_[23828]_ , \new_[23829]_ ,
    \new_[23833]_ , \new_[23834]_ , \new_[23838]_ , \new_[23839]_ ,
    \new_[23840]_ , \new_[23843]_ , \new_[23847]_ , \new_[23848]_ ,
    \new_[23849]_ , \new_[23853]_ , \new_[23854]_ , \new_[23858]_ ,
    \new_[23859]_ , \new_[23860]_ , \new_[23863]_ , \new_[23867]_ ,
    \new_[23868]_ , \new_[23869]_ , \new_[23873]_ , \new_[23874]_ ,
    \new_[23878]_ , \new_[23879]_ , \new_[23880]_ , \new_[23883]_ ,
    \new_[23887]_ , \new_[23888]_ , \new_[23889]_ , \new_[23893]_ ,
    \new_[23894]_ , \new_[23898]_ , \new_[23899]_ , \new_[23900]_ ,
    \new_[23903]_ , \new_[23907]_ , \new_[23908]_ , \new_[23909]_ ,
    \new_[23913]_ , \new_[23914]_ , \new_[23918]_ , \new_[23919]_ ,
    \new_[23920]_ , \new_[23923]_ , \new_[23927]_ , \new_[23928]_ ,
    \new_[23929]_ , \new_[23933]_ , \new_[23934]_ , \new_[23938]_ ,
    \new_[23939]_ , \new_[23940]_ , \new_[23943]_ , \new_[23947]_ ,
    \new_[23948]_ , \new_[23949]_ , \new_[23953]_ , \new_[23954]_ ,
    \new_[23958]_ , \new_[23959]_ , \new_[23960]_ , \new_[23963]_ ,
    \new_[23967]_ , \new_[23968]_ , \new_[23969]_ , \new_[23973]_ ,
    \new_[23974]_ , \new_[23978]_ , \new_[23979]_ , \new_[23980]_ ,
    \new_[23983]_ , \new_[23987]_ , \new_[23988]_ , \new_[23989]_ ,
    \new_[23993]_ , \new_[23994]_ , \new_[23998]_ , \new_[23999]_ ,
    \new_[24000]_ , \new_[24003]_ , \new_[24007]_ , \new_[24008]_ ,
    \new_[24009]_ , \new_[24013]_ , \new_[24014]_ , \new_[24018]_ ,
    \new_[24019]_ , \new_[24020]_ , \new_[24023]_ , \new_[24027]_ ,
    \new_[24028]_ , \new_[24029]_ , \new_[24033]_ , \new_[24034]_ ,
    \new_[24038]_ , \new_[24039]_ , \new_[24040]_ , \new_[24043]_ ,
    \new_[24047]_ , \new_[24048]_ , \new_[24049]_ , \new_[24053]_ ,
    \new_[24054]_ , \new_[24058]_ , \new_[24059]_ , \new_[24060]_ ,
    \new_[24063]_ , \new_[24067]_ , \new_[24068]_ , \new_[24069]_ ,
    \new_[24073]_ , \new_[24074]_ , \new_[24078]_ , \new_[24079]_ ,
    \new_[24080]_ , \new_[24083]_ , \new_[24087]_ , \new_[24088]_ ,
    \new_[24089]_ , \new_[24093]_ , \new_[24094]_ , \new_[24098]_ ,
    \new_[24099]_ , \new_[24100]_ , \new_[24103]_ , \new_[24107]_ ,
    \new_[24108]_ , \new_[24109]_ , \new_[24113]_ , \new_[24114]_ ,
    \new_[24118]_ , \new_[24119]_ , \new_[24120]_ , \new_[24123]_ ,
    \new_[24127]_ , \new_[24128]_ , \new_[24129]_ , \new_[24133]_ ,
    \new_[24134]_ , \new_[24138]_ , \new_[24139]_ , \new_[24140]_ ,
    \new_[24143]_ , \new_[24147]_ , \new_[24148]_ , \new_[24149]_ ,
    \new_[24153]_ , \new_[24154]_ , \new_[24158]_ , \new_[24159]_ ,
    \new_[24160]_ , \new_[24163]_ , \new_[24167]_ , \new_[24168]_ ,
    \new_[24169]_ , \new_[24173]_ , \new_[24174]_ , \new_[24178]_ ,
    \new_[24179]_ , \new_[24180]_ , \new_[24183]_ , \new_[24187]_ ,
    \new_[24188]_ , \new_[24189]_ , \new_[24193]_ , \new_[24194]_ ,
    \new_[24198]_ , \new_[24199]_ , \new_[24200]_ , \new_[24203]_ ,
    \new_[24207]_ , \new_[24208]_ , \new_[24209]_ , \new_[24213]_ ,
    \new_[24214]_ , \new_[24218]_ , \new_[24219]_ , \new_[24220]_ ,
    \new_[24223]_ , \new_[24227]_ , \new_[24228]_ , \new_[24229]_ ,
    \new_[24233]_ , \new_[24234]_ , \new_[24238]_ , \new_[24239]_ ,
    \new_[24240]_ , \new_[24243]_ , \new_[24247]_ , \new_[24248]_ ,
    \new_[24249]_ , \new_[24253]_ , \new_[24254]_ , \new_[24258]_ ,
    \new_[24259]_ , \new_[24260]_ , \new_[24263]_ , \new_[24267]_ ,
    \new_[24268]_ , \new_[24269]_ , \new_[24273]_ , \new_[24274]_ ,
    \new_[24278]_ , \new_[24279]_ , \new_[24280]_ , \new_[24283]_ ,
    \new_[24287]_ , \new_[24288]_ , \new_[24289]_ , \new_[24293]_ ,
    \new_[24294]_ , \new_[24298]_ , \new_[24299]_ , \new_[24300]_ ,
    \new_[24303]_ , \new_[24307]_ , \new_[24308]_ , \new_[24309]_ ,
    \new_[24313]_ , \new_[24314]_ , \new_[24318]_ , \new_[24319]_ ,
    \new_[24320]_ , \new_[24323]_ , \new_[24327]_ , \new_[24328]_ ,
    \new_[24329]_ , \new_[24333]_ , \new_[24334]_ , \new_[24338]_ ,
    \new_[24339]_ , \new_[24340]_ , \new_[24343]_ , \new_[24347]_ ,
    \new_[24348]_ , \new_[24349]_ , \new_[24353]_ , \new_[24354]_ ,
    \new_[24358]_ , \new_[24359]_ , \new_[24360]_ , \new_[24363]_ ,
    \new_[24367]_ , \new_[24368]_ , \new_[24369]_ , \new_[24373]_ ,
    \new_[24374]_ , \new_[24378]_ , \new_[24379]_ , \new_[24380]_ ,
    \new_[24383]_ , \new_[24387]_ , \new_[24388]_ , \new_[24389]_ ,
    \new_[24393]_ , \new_[24394]_ , \new_[24398]_ , \new_[24399]_ ,
    \new_[24400]_ , \new_[24403]_ , \new_[24407]_ , \new_[24408]_ ,
    \new_[24409]_ , \new_[24413]_ , \new_[24414]_ , \new_[24418]_ ,
    \new_[24419]_ , \new_[24420]_ , \new_[24423]_ , \new_[24427]_ ,
    \new_[24428]_ , \new_[24429]_ , \new_[24433]_ , \new_[24434]_ ,
    \new_[24438]_ , \new_[24439]_ , \new_[24440]_ , \new_[24443]_ ,
    \new_[24447]_ , \new_[24448]_ , \new_[24449]_ , \new_[24453]_ ,
    \new_[24454]_ , \new_[24458]_ , \new_[24459]_ , \new_[24460]_ ,
    \new_[24464]_ , \new_[24465]_ , \new_[24469]_ , \new_[24470]_ ,
    \new_[24471]_ , \new_[24475]_ , \new_[24476]_ , \new_[24480]_ ,
    \new_[24481]_ , \new_[24482]_ , \new_[24486]_ , \new_[24487]_ ,
    \new_[24491]_ , \new_[24492]_ , \new_[24493]_ , \new_[24497]_ ,
    \new_[24498]_ , \new_[24502]_ , \new_[24503]_ , \new_[24504]_ ,
    \new_[24508]_ , \new_[24509]_ , \new_[24513]_ , \new_[24514]_ ,
    \new_[24515]_ , \new_[24519]_ , \new_[24520]_ , \new_[24524]_ ,
    \new_[24525]_ , \new_[24526]_ , \new_[24530]_ , \new_[24531]_ ,
    \new_[24535]_ , \new_[24536]_ , \new_[24537]_ , \new_[24541]_ ,
    \new_[24542]_ , \new_[24546]_ , \new_[24547]_ , \new_[24548]_ ,
    \new_[24552]_ , \new_[24553]_ , \new_[24557]_ , \new_[24558]_ ,
    \new_[24559]_ , \new_[24563]_ , \new_[24564]_ , \new_[24568]_ ,
    \new_[24569]_ , \new_[24570]_ , \new_[24574]_ , \new_[24575]_ ,
    \new_[24579]_ , \new_[24580]_ , \new_[24581]_ , \new_[24585]_ ,
    \new_[24586]_ , \new_[24590]_ , \new_[24591]_ , \new_[24592]_ ,
    \new_[24596]_ , \new_[24597]_ , \new_[24601]_ , \new_[24602]_ ,
    \new_[24603]_ , \new_[24607]_ , \new_[24608]_ , \new_[24612]_ ,
    \new_[24613]_ , \new_[24614]_ , \new_[24618]_ , \new_[24619]_ ,
    \new_[24623]_ , \new_[24624]_ , \new_[24625]_ , \new_[24629]_ ,
    \new_[24630]_ , \new_[24634]_ , \new_[24635]_ , \new_[24636]_ ,
    \new_[24640]_ , \new_[24641]_ , \new_[24645]_ , \new_[24646]_ ,
    \new_[24647]_ , \new_[24651]_ , \new_[24652]_ , \new_[24656]_ ,
    \new_[24657]_ , \new_[24658]_ , \new_[24662]_ , \new_[24663]_ ,
    \new_[24667]_ , \new_[24668]_ , \new_[24669]_ , \new_[24673]_ ,
    \new_[24674]_ , \new_[24678]_ , \new_[24679]_ , \new_[24680]_ ,
    \new_[24684]_ , \new_[24685]_ , \new_[24689]_ , \new_[24690]_ ,
    \new_[24691]_ , \new_[24695]_ , \new_[24696]_ , \new_[24700]_ ,
    \new_[24701]_ , \new_[24702]_ , \new_[24706]_ , \new_[24707]_ ,
    \new_[24711]_ , \new_[24712]_ , \new_[24713]_ , \new_[24717]_ ,
    \new_[24718]_ , \new_[24722]_ , \new_[24723]_ , \new_[24724]_ ,
    \new_[24728]_ , \new_[24729]_ , \new_[24733]_ , \new_[24734]_ ,
    \new_[24735]_ , \new_[24739]_ , \new_[24740]_ , \new_[24744]_ ,
    \new_[24745]_ , \new_[24746]_ , \new_[24750]_ , \new_[24751]_ ,
    \new_[24755]_ , \new_[24756]_ , \new_[24757]_ , \new_[24761]_ ,
    \new_[24762]_ , \new_[24766]_ , \new_[24767]_ , \new_[24768]_ ,
    \new_[24772]_ , \new_[24773]_ , \new_[24777]_ , \new_[24778]_ ,
    \new_[24779]_ , \new_[24783]_ , \new_[24784]_ , \new_[24788]_ ,
    \new_[24789]_ , \new_[24790]_ , \new_[24794]_ , \new_[24795]_ ,
    \new_[24799]_ , \new_[24800]_ , \new_[24801]_ , \new_[24805]_ ,
    \new_[24806]_ , \new_[24810]_ , \new_[24811]_ , \new_[24812]_ ,
    \new_[24816]_ , \new_[24817]_ , \new_[24821]_ , \new_[24822]_ ,
    \new_[24823]_ , \new_[24827]_ , \new_[24828]_ , \new_[24832]_ ,
    \new_[24833]_ , \new_[24834]_ , \new_[24838]_ , \new_[24839]_ ,
    \new_[24843]_ , \new_[24844]_ , \new_[24845]_ , \new_[24849]_ ,
    \new_[24850]_ , \new_[24854]_ , \new_[24855]_ , \new_[24856]_ ,
    \new_[24860]_ , \new_[24861]_ , \new_[24865]_ , \new_[24866]_ ,
    \new_[24867]_ , \new_[24871]_ , \new_[24872]_ , \new_[24876]_ ,
    \new_[24877]_ , \new_[24878]_ , \new_[24882]_ , \new_[24883]_ ,
    \new_[24887]_ , \new_[24888]_ , \new_[24889]_ , \new_[24893]_ ,
    \new_[24894]_ , \new_[24898]_ , \new_[24899]_ , \new_[24900]_ ,
    \new_[24904]_ , \new_[24905]_ , \new_[24909]_ , \new_[24910]_ ,
    \new_[24911]_ , \new_[24915]_ , \new_[24916]_ , \new_[24920]_ ,
    \new_[24921]_ , \new_[24922]_ , \new_[24926]_ , \new_[24927]_ ,
    \new_[24931]_ , \new_[24932]_ , \new_[24933]_ , \new_[24937]_ ,
    \new_[24938]_ , \new_[24942]_ , \new_[24943]_ , \new_[24944]_ ,
    \new_[24948]_ , \new_[24949]_ , \new_[24953]_ , \new_[24954]_ ,
    \new_[24955]_ , \new_[24959]_ , \new_[24960]_ , \new_[24964]_ ,
    \new_[24965]_ , \new_[24966]_ , \new_[24970]_ , \new_[24971]_ ,
    \new_[24975]_ , \new_[24976]_ , \new_[24977]_ , \new_[24981]_ ,
    \new_[24982]_ , \new_[24986]_ , \new_[24987]_ , \new_[24988]_ ,
    \new_[24992]_ , \new_[24993]_ , \new_[24997]_ , \new_[24998]_ ,
    \new_[24999]_ , \new_[25003]_ , \new_[25004]_ , \new_[25008]_ ,
    \new_[25009]_ , \new_[25010]_ , \new_[25014]_ , \new_[25015]_ ,
    \new_[25019]_ , \new_[25020]_ , \new_[25021]_ , \new_[25025]_ ,
    \new_[25026]_ , \new_[25030]_ , \new_[25031]_ , \new_[25032]_ ,
    \new_[25036]_ , \new_[25037]_ , \new_[25041]_ , \new_[25042]_ ,
    \new_[25043]_ , \new_[25047]_ , \new_[25048]_ , \new_[25052]_ ,
    \new_[25053]_ , \new_[25054]_ , \new_[25058]_ , \new_[25059]_ ,
    \new_[25063]_ , \new_[25064]_ , \new_[25065]_ , \new_[25069]_ ,
    \new_[25070]_ , \new_[25074]_ , \new_[25075]_ , \new_[25076]_ ,
    \new_[25080]_ , \new_[25081]_ , \new_[25085]_ , \new_[25086]_ ,
    \new_[25087]_ , \new_[25091]_ , \new_[25092]_ , \new_[25096]_ ,
    \new_[25097]_ , \new_[25098]_ , \new_[25102]_ , \new_[25103]_ ,
    \new_[25107]_ , \new_[25108]_ , \new_[25109]_ , \new_[25113]_ ,
    \new_[25114]_ , \new_[25118]_ , \new_[25119]_ , \new_[25120]_ ,
    \new_[25124]_ , \new_[25125]_ , \new_[25129]_ , \new_[25130]_ ,
    \new_[25131]_ , \new_[25135]_ , \new_[25136]_ , \new_[25140]_ ,
    \new_[25141]_ , \new_[25142]_ , \new_[25146]_ , \new_[25147]_ ,
    \new_[25151]_ , \new_[25152]_ , \new_[25153]_ , \new_[25157]_ ,
    \new_[25158]_ , \new_[25162]_ , \new_[25163]_ , \new_[25164]_ ,
    \new_[25168]_ , \new_[25169]_ , \new_[25173]_ , \new_[25174]_ ,
    \new_[25175]_ , \new_[25179]_ , \new_[25180]_ , \new_[25184]_ ,
    \new_[25185]_ , \new_[25186]_ , \new_[25190]_ , \new_[25191]_ ,
    \new_[25195]_ , \new_[25196]_ , \new_[25197]_ , \new_[25201]_ ,
    \new_[25202]_ , \new_[25206]_ , \new_[25207]_ , \new_[25208]_ ,
    \new_[25212]_ , \new_[25213]_ , \new_[25217]_ , \new_[25218]_ ,
    \new_[25219]_ , \new_[25223]_ , \new_[25224]_ , \new_[25228]_ ,
    \new_[25229]_ , \new_[25230]_ , \new_[25234]_ , \new_[25235]_ ,
    \new_[25239]_ , \new_[25240]_ , \new_[25241]_ , \new_[25245]_ ,
    \new_[25246]_ , \new_[25250]_ , \new_[25251]_ , \new_[25252]_ ,
    \new_[25256]_ , \new_[25257]_ , \new_[25261]_ , \new_[25262]_ ,
    \new_[25263]_ , \new_[25267]_ , \new_[25268]_ , \new_[25272]_ ,
    \new_[25273]_ , \new_[25274]_ , \new_[25278]_ , \new_[25279]_ ,
    \new_[25283]_ , \new_[25284]_ , \new_[25285]_ , \new_[25289]_ ,
    \new_[25290]_ , \new_[25294]_ , \new_[25295]_ , \new_[25296]_ ,
    \new_[25300]_ , \new_[25301]_ , \new_[25305]_ , \new_[25306]_ ,
    \new_[25307]_ , \new_[25311]_ , \new_[25312]_ , \new_[25316]_ ,
    \new_[25317]_ , \new_[25318]_ , \new_[25322]_ , \new_[25323]_ ,
    \new_[25327]_ , \new_[25328]_ , \new_[25329]_ , \new_[25333]_ ,
    \new_[25334]_ , \new_[25338]_ , \new_[25339]_ , \new_[25340]_ ,
    \new_[25344]_ , \new_[25345]_ , \new_[25349]_ , \new_[25350]_ ,
    \new_[25351]_ , \new_[25355]_ , \new_[25356]_ , \new_[25360]_ ,
    \new_[25361]_ , \new_[25362]_ , \new_[25366]_ , \new_[25367]_ ,
    \new_[25371]_ , \new_[25372]_ , \new_[25373]_ , \new_[25377]_ ,
    \new_[25378]_ , \new_[25382]_ , \new_[25383]_ , \new_[25384]_ ,
    \new_[25388]_ , \new_[25389]_ , \new_[25393]_ , \new_[25394]_ ,
    \new_[25395]_ , \new_[25399]_ , \new_[25400]_ , \new_[25404]_ ,
    \new_[25405]_ , \new_[25406]_ , \new_[25410]_ , \new_[25411]_ ,
    \new_[25415]_ , \new_[25416]_ , \new_[25417]_ , \new_[25421]_ ,
    \new_[25422]_ , \new_[25426]_ , \new_[25427]_ , \new_[25428]_ ,
    \new_[25432]_ , \new_[25433]_ , \new_[25437]_ , \new_[25438]_ ,
    \new_[25439]_ , \new_[25443]_ , \new_[25444]_ , \new_[25448]_ ,
    \new_[25449]_ , \new_[25450]_ , \new_[25454]_ , \new_[25455]_ ,
    \new_[25459]_ , \new_[25460]_ , \new_[25461]_ , \new_[25465]_ ,
    \new_[25466]_ , \new_[25470]_ , \new_[25471]_ , \new_[25472]_ ,
    \new_[25476]_ , \new_[25477]_ , \new_[25481]_ , \new_[25482]_ ,
    \new_[25483]_ , \new_[25487]_ , \new_[25488]_ , \new_[25492]_ ,
    \new_[25493]_ , \new_[25494]_ , \new_[25498]_ , \new_[25499]_ ,
    \new_[25503]_ , \new_[25504]_ , \new_[25505]_ , \new_[25509]_ ,
    \new_[25510]_ , \new_[25514]_ , \new_[25515]_ , \new_[25516]_ ,
    \new_[25520]_ , \new_[25521]_ , \new_[25525]_ , \new_[25526]_ ,
    \new_[25527]_ , \new_[25531]_ , \new_[25532]_ , \new_[25536]_ ,
    \new_[25537]_ , \new_[25538]_ , \new_[25542]_ , \new_[25543]_ ,
    \new_[25547]_ , \new_[25548]_ , \new_[25549]_ , \new_[25553]_ ,
    \new_[25554]_ , \new_[25558]_ , \new_[25559]_ , \new_[25560]_ ,
    \new_[25564]_ , \new_[25565]_ , \new_[25569]_ , \new_[25570]_ ,
    \new_[25571]_ , \new_[25575]_ , \new_[25576]_ , \new_[25580]_ ,
    \new_[25581]_ , \new_[25582]_ , \new_[25586]_ , \new_[25587]_ ,
    \new_[25591]_ , \new_[25592]_ , \new_[25593]_ , \new_[25597]_ ,
    \new_[25598]_ , \new_[25602]_ , \new_[25603]_ , \new_[25604]_ ,
    \new_[25608]_ , \new_[25609]_ , \new_[25613]_ , \new_[25614]_ ,
    \new_[25615]_ , \new_[25619]_ , \new_[25620]_ , \new_[25624]_ ,
    \new_[25625]_ , \new_[25626]_ , \new_[25630]_ , \new_[25631]_ ,
    \new_[25635]_ , \new_[25636]_ , \new_[25637]_ , \new_[25641]_ ,
    \new_[25642]_ , \new_[25646]_ , \new_[25647]_ , \new_[25648]_ ,
    \new_[25652]_ , \new_[25653]_ , \new_[25657]_ , \new_[25658]_ ,
    \new_[25659]_ , \new_[25663]_ , \new_[25664]_ , \new_[25668]_ ,
    \new_[25669]_ , \new_[25670]_ , \new_[25674]_ , \new_[25675]_ ,
    \new_[25679]_ , \new_[25680]_ , \new_[25681]_ , \new_[25685]_ ,
    \new_[25686]_ , \new_[25690]_ , \new_[25691]_ , \new_[25692]_ ,
    \new_[25696]_ , \new_[25697]_ , \new_[25701]_ , \new_[25702]_ ,
    \new_[25703]_ , \new_[25707]_ , \new_[25708]_ , \new_[25712]_ ,
    \new_[25713]_ , \new_[25714]_ , \new_[25718]_ , \new_[25719]_ ,
    \new_[25723]_ , \new_[25724]_ , \new_[25725]_ , \new_[25729]_ ,
    \new_[25730]_ , \new_[25734]_ , \new_[25735]_ , \new_[25736]_ ,
    \new_[25740]_ , \new_[25741]_ , \new_[25745]_ , \new_[25746]_ ,
    \new_[25747]_ , \new_[25751]_ , \new_[25752]_ , \new_[25756]_ ,
    \new_[25757]_ , \new_[25758]_ , \new_[25762]_ , \new_[25763]_ ,
    \new_[25767]_ , \new_[25768]_ , \new_[25769]_ , \new_[25773]_ ,
    \new_[25774]_ , \new_[25778]_ , \new_[25779]_ , \new_[25780]_ ,
    \new_[25784]_ , \new_[25785]_ , \new_[25789]_ , \new_[25790]_ ,
    \new_[25791]_ , \new_[25795]_ , \new_[25796]_ , \new_[25800]_ ,
    \new_[25801]_ , \new_[25802]_ , \new_[25806]_ , \new_[25807]_ ,
    \new_[25811]_ , \new_[25812]_ , \new_[25813]_ , \new_[25817]_ ,
    \new_[25818]_ , \new_[25822]_ , \new_[25823]_ , \new_[25824]_ ,
    \new_[25828]_ , \new_[25829]_ , \new_[25833]_ , \new_[25834]_ ,
    \new_[25835]_ , \new_[25839]_ , \new_[25840]_ , \new_[25844]_ ,
    \new_[25845]_ , \new_[25846]_ , \new_[25850]_ , \new_[25851]_ ,
    \new_[25855]_ , \new_[25856]_ , \new_[25857]_ , \new_[25861]_ ,
    \new_[25862]_ , \new_[25866]_ , \new_[25867]_ , \new_[25868]_ ,
    \new_[25872]_ , \new_[25873]_ , \new_[25877]_ , \new_[25878]_ ,
    \new_[25879]_ , \new_[25883]_ , \new_[25884]_ , \new_[25888]_ ,
    \new_[25889]_ , \new_[25890]_ , \new_[25894]_ , \new_[25895]_ ,
    \new_[25899]_ , \new_[25900]_ , \new_[25901]_ , \new_[25905]_ ,
    \new_[25906]_ , \new_[25910]_ , \new_[25911]_ , \new_[25912]_ ,
    \new_[25916]_ , \new_[25917]_ , \new_[25921]_ , \new_[25922]_ ,
    \new_[25923]_ , \new_[25927]_ , \new_[25928]_ , \new_[25932]_ ,
    \new_[25933]_ , \new_[25934]_ , \new_[25938]_ , \new_[25939]_ ,
    \new_[25943]_ , \new_[25944]_ , \new_[25945]_ , \new_[25949]_ ,
    \new_[25950]_ , \new_[25954]_ , \new_[25955]_ , \new_[25956]_ ,
    \new_[25960]_ , \new_[25961]_ , \new_[25965]_ , \new_[25966]_ ,
    \new_[25967]_ , \new_[25971]_ , \new_[25972]_ , \new_[25976]_ ,
    \new_[25977]_ , \new_[25978]_ , \new_[25982]_ , \new_[25983]_ ,
    \new_[25987]_ , \new_[25988]_ , \new_[25989]_ , \new_[25993]_ ,
    \new_[25994]_ , \new_[25998]_ , \new_[25999]_ , \new_[26000]_ ,
    \new_[26004]_ , \new_[26005]_ , \new_[26009]_ , \new_[26010]_ ,
    \new_[26011]_ , \new_[26015]_ , \new_[26016]_ , \new_[26020]_ ,
    \new_[26021]_ , \new_[26022]_ , \new_[26026]_ , \new_[26027]_ ,
    \new_[26031]_ , \new_[26032]_ , \new_[26033]_ , \new_[26037]_ ,
    \new_[26038]_ , \new_[26042]_ , \new_[26043]_ , \new_[26044]_ ,
    \new_[26048]_ , \new_[26049]_ , \new_[26053]_ , \new_[26054]_ ,
    \new_[26055]_ , \new_[26059]_ , \new_[26060]_ , \new_[26064]_ ,
    \new_[26065]_ , \new_[26066]_ , \new_[26070]_ , \new_[26071]_ ,
    \new_[26075]_ , \new_[26076]_ , \new_[26077]_ , \new_[26081]_ ,
    \new_[26082]_ , \new_[26086]_ , \new_[26087]_ , \new_[26088]_ ,
    \new_[26092]_ , \new_[26093]_ , \new_[26097]_ , \new_[26098]_ ,
    \new_[26099]_ , \new_[26103]_ , \new_[26104]_ , \new_[26108]_ ,
    \new_[26109]_ , \new_[26110]_ , \new_[26114]_ , \new_[26115]_ ,
    \new_[26119]_ , \new_[26120]_ , \new_[26121]_ , \new_[26125]_ ,
    \new_[26126]_ , \new_[26130]_ , \new_[26131]_ , \new_[26132]_ ,
    \new_[26136]_ , \new_[26137]_ , \new_[26141]_ , \new_[26142]_ ,
    \new_[26143]_ , \new_[26147]_ , \new_[26148]_ , \new_[26152]_ ,
    \new_[26153]_ , \new_[26154]_ , \new_[26158]_ , \new_[26159]_ ,
    \new_[26163]_ , \new_[26164]_ , \new_[26165]_ , \new_[26169]_ ,
    \new_[26170]_ , \new_[26174]_ , \new_[26175]_ , \new_[26176]_ ,
    \new_[26180]_ , \new_[26181]_ , \new_[26185]_ , \new_[26186]_ ,
    \new_[26187]_ , \new_[26191]_ , \new_[26192]_ , \new_[26196]_ ,
    \new_[26197]_ , \new_[26198]_ , \new_[26202]_ , \new_[26203]_ ,
    \new_[26207]_ , \new_[26208]_ , \new_[26209]_ , \new_[26213]_ ,
    \new_[26214]_ , \new_[26218]_ , \new_[26219]_ , \new_[26220]_ ,
    \new_[26224]_ , \new_[26225]_ , \new_[26229]_ , \new_[26230]_ ,
    \new_[26231]_ , \new_[26235]_ , \new_[26236]_ , \new_[26240]_ ,
    \new_[26241]_ , \new_[26242]_ , \new_[26246]_ , \new_[26247]_ ,
    \new_[26251]_ , \new_[26252]_ , \new_[26253]_ , \new_[26257]_ ,
    \new_[26258]_ , \new_[26262]_ , \new_[26263]_ , \new_[26264]_ ,
    \new_[26268]_ , \new_[26269]_ , \new_[26273]_ , \new_[26274]_ ,
    \new_[26275]_ , \new_[26279]_ , \new_[26280]_ , \new_[26284]_ ,
    \new_[26285]_ , \new_[26286]_ , \new_[26290]_ , \new_[26291]_ ,
    \new_[26295]_ , \new_[26296]_ , \new_[26297]_ , \new_[26301]_ ,
    \new_[26302]_ , \new_[26306]_ , \new_[26307]_ , \new_[26308]_ ,
    \new_[26312]_ , \new_[26313]_ , \new_[26317]_ , \new_[26318]_ ,
    \new_[26319]_ , \new_[26323]_ , \new_[26324]_ , \new_[26328]_ ,
    \new_[26329]_ , \new_[26330]_ , \new_[26334]_ , \new_[26335]_ ,
    \new_[26339]_ , \new_[26340]_ , \new_[26341]_ , \new_[26345]_ ,
    \new_[26346]_ , \new_[26350]_ , \new_[26351]_ , \new_[26352]_ ,
    \new_[26356]_ , \new_[26357]_ , \new_[26361]_ , \new_[26362]_ ,
    \new_[26363]_ , \new_[26367]_ , \new_[26368]_ , \new_[26372]_ ,
    \new_[26373]_ , \new_[26374]_ , \new_[26378]_ , \new_[26379]_ ,
    \new_[26383]_ , \new_[26384]_ , \new_[26385]_ , \new_[26389]_ ,
    \new_[26390]_ , \new_[26394]_ , \new_[26395]_ , \new_[26396]_ ,
    \new_[26400]_ , \new_[26401]_ , \new_[26405]_ , \new_[26406]_ ,
    \new_[26407]_ , \new_[26411]_ , \new_[26412]_ , \new_[26416]_ ,
    \new_[26417]_ , \new_[26418]_ , \new_[26422]_ , \new_[26423]_ ,
    \new_[26427]_ , \new_[26428]_ , \new_[26429]_ , \new_[26433]_ ,
    \new_[26434]_ , \new_[26438]_ , \new_[26439]_ , \new_[26440]_ ,
    \new_[26444]_ , \new_[26445]_ , \new_[26449]_ , \new_[26450]_ ,
    \new_[26451]_ , \new_[26455]_ , \new_[26456]_ , \new_[26460]_ ,
    \new_[26461]_ , \new_[26462]_ , \new_[26466]_ , \new_[26467]_ ,
    \new_[26471]_ , \new_[26472]_ , \new_[26473]_ , \new_[26477]_ ,
    \new_[26478]_ , \new_[26482]_ , \new_[26483]_ , \new_[26484]_ ,
    \new_[26488]_ , \new_[26489]_ , \new_[26493]_ , \new_[26494]_ ,
    \new_[26495]_ , \new_[26499]_ , \new_[26500]_ , \new_[26504]_ ,
    \new_[26505]_ , \new_[26506]_ , \new_[26510]_ , \new_[26511]_ ,
    \new_[26515]_ , \new_[26516]_ , \new_[26517]_ , \new_[26521]_ ,
    \new_[26522]_ , \new_[26526]_ , \new_[26527]_ , \new_[26528]_ ,
    \new_[26532]_ , \new_[26533]_ , \new_[26537]_ , \new_[26538]_ ,
    \new_[26539]_ , \new_[26543]_ , \new_[26544]_ , \new_[26548]_ ,
    \new_[26549]_ , \new_[26550]_ , \new_[26554]_ , \new_[26555]_ ,
    \new_[26559]_ , \new_[26560]_ , \new_[26561]_ , \new_[26565]_ ,
    \new_[26566]_ , \new_[26570]_ , \new_[26571]_ , \new_[26572]_ ,
    \new_[26576]_ , \new_[26577]_ , \new_[26581]_ , \new_[26582]_ ,
    \new_[26583]_ , \new_[26587]_ , \new_[26588]_ , \new_[26592]_ ,
    \new_[26593]_ , \new_[26594]_ , \new_[26598]_ , \new_[26599]_ ,
    \new_[26603]_ , \new_[26604]_ , \new_[26605]_ , \new_[26609]_ ,
    \new_[26610]_ , \new_[26614]_ , \new_[26615]_ , \new_[26616]_ ,
    \new_[26620]_ , \new_[26621]_ , \new_[26625]_ , \new_[26626]_ ,
    \new_[26627]_ , \new_[26631]_ , \new_[26632]_ , \new_[26636]_ ,
    \new_[26637]_ , \new_[26638]_ , \new_[26642]_ , \new_[26643]_ ,
    \new_[26647]_ , \new_[26648]_ , \new_[26649]_ , \new_[26653]_ ,
    \new_[26654]_ , \new_[26658]_ , \new_[26659]_ , \new_[26660]_ ,
    \new_[26664]_ , \new_[26665]_ , \new_[26669]_ , \new_[26670]_ ,
    \new_[26671]_ , \new_[26675]_ , \new_[26676]_ , \new_[26680]_ ,
    \new_[26681]_ , \new_[26682]_ , \new_[26686]_ , \new_[26687]_ ,
    \new_[26691]_ , \new_[26692]_ , \new_[26693]_ , \new_[26697]_ ,
    \new_[26698]_ , \new_[26702]_ , \new_[26703]_ , \new_[26704]_ ,
    \new_[26708]_ , \new_[26709]_ , \new_[26713]_ , \new_[26714]_ ,
    \new_[26715]_ , \new_[26719]_ , \new_[26720]_ , \new_[26724]_ ,
    \new_[26725]_ , \new_[26726]_ , \new_[26730]_ , \new_[26731]_ ,
    \new_[26735]_ , \new_[26736]_ , \new_[26737]_ , \new_[26741]_ ,
    \new_[26742]_ , \new_[26746]_ , \new_[26747]_ , \new_[26748]_ ,
    \new_[26752]_ , \new_[26753]_ , \new_[26757]_ , \new_[26758]_ ,
    \new_[26759]_ , \new_[26763]_ , \new_[26764]_ , \new_[26768]_ ,
    \new_[26769]_ , \new_[26770]_ , \new_[26774]_ , \new_[26775]_ ,
    \new_[26779]_ , \new_[26780]_ , \new_[26781]_ , \new_[26785]_ ,
    \new_[26786]_ , \new_[26790]_ , \new_[26791]_ , \new_[26792]_ ,
    \new_[26796]_ , \new_[26797]_ , \new_[26801]_ , \new_[26802]_ ,
    \new_[26803]_ , \new_[26807]_ , \new_[26808]_ , \new_[26812]_ ,
    \new_[26813]_ , \new_[26814]_ , \new_[26818]_ , \new_[26819]_ ,
    \new_[26823]_ , \new_[26824]_ , \new_[26825]_ , \new_[26829]_ ,
    \new_[26830]_ , \new_[26834]_ , \new_[26835]_ , \new_[26836]_ ,
    \new_[26840]_ , \new_[26841]_ , \new_[26845]_ , \new_[26846]_ ,
    \new_[26847]_ , \new_[26851]_ , \new_[26852]_ , \new_[26856]_ ,
    \new_[26857]_ , \new_[26858]_ , \new_[26862]_ , \new_[26863]_ ,
    \new_[26867]_ , \new_[26868]_ , \new_[26869]_ , \new_[26873]_ ,
    \new_[26874]_ , \new_[26878]_ , \new_[26879]_ , \new_[26880]_ ,
    \new_[26884]_ , \new_[26885]_ , \new_[26889]_ , \new_[26890]_ ,
    \new_[26891]_ , \new_[26895]_ , \new_[26896]_ , \new_[26900]_ ,
    \new_[26901]_ , \new_[26902]_ , \new_[26906]_ , \new_[26907]_ ,
    \new_[26911]_ , \new_[26912]_ , \new_[26913]_ , \new_[26917]_ ,
    \new_[26918]_ , \new_[26922]_ , \new_[26923]_ , \new_[26924]_ ,
    \new_[26928]_ , \new_[26929]_ , \new_[26933]_ , \new_[26934]_ ,
    \new_[26935]_ , \new_[26939]_ , \new_[26940]_ , \new_[26944]_ ,
    \new_[26945]_ , \new_[26946]_ , \new_[26950]_ , \new_[26951]_ ,
    \new_[26955]_ , \new_[26956]_ , \new_[26957]_ , \new_[26961]_ ,
    \new_[26962]_ , \new_[26966]_ , \new_[26967]_ , \new_[26968]_ ,
    \new_[26972]_ , \new_[26973]_ , \new_[26977]_ , \new_[26978]_ ,
    \new_[26979]_ , \new_[26983]_ , \new_[26984]_ , \new_[26988]_ ,
    \new_[26989]_ , \new_[26990]_ , \new_[26994]_ , \new_[26995]_ ,
    \new_[26999]_ , \new_[27000]_ , \new_[27001]_ , \new_[27005]_ ,
    \new_[27006]_ , \new_[27010]_ , \new_[27011]_ , \new_[27012]_ ,
    \new_[27016]_ , \new_[27017]_ , \new_[27021]_ , \new_[27022]_ ,
    \new_[27023]_ , \new_[27027]_ , \new_[27028]_ , \new_[27032]_ ,
    \new_[27033]_ , \new_[27034]_ , \new_[27038]_ , \new_[27039]_ ,
    \new_[27043]_ , \new_[27044]_ , \new_[27045]_ , \new_[27049]_ ,
    \new_[27050]_ , \new_[27054]_ , \new_[27055]_ , \new_[27056]_ ,
    \new_[27060]_ , \new_[27061]_ , \new_[27065]_ , \new_[27066]_ ,
    \new_[27067]_ , \new_[27071]_ , \new_[27072]_ , \new_[27076]_ ,
    \new_[27077]_ , \new_[27078]_ , \new_[27082]_ , \new_[27083]_ ,
    \new_[27087]_ , \new_[27088]_ , \new_[27089]_ , \new_[27093]_ ,
    \new_[27094]_ , \new_[27098]_ , \new_[27099]_ , \new_[27100]_ ,
    \new_[27104]_ , \new_[27105]_ , \new_[27109]_ , \new_[27110]_ ,
    \new_[27111]_ , \new_[27115]_ , \new_[27116]_ , \new_[27120]_ ,
    \new_[27121]_ , \new_[27122]_ , \new_[27126]_ , \new_[27127]_ ,
    \new_[27131]_ , \new_[27132]_ , \new_[27133]_ , \new_[27137]_ ,
    \new_[27138]_ , \new_[27142]_ , \new_[27143]_ , \new_[27144]_ ,
    \new_[27148]_ , \new_[27149]_ , \new_[27153]_ , \new_[27154]_ ,
    \new_[27155]_ , \new_[27159]_ , \new_[27160]_ , \new_[27164]_ ,
    \new_[27165]_ , \new_[27166]_ , \new_[27170]_ , \new_[27171]_ ,
    \new_[27175]_ , \new_[27176]_ , \new_[27177]_ , \new_[27181]_ ,
    \new_[27182]_ , \new_[27186]_ , \new_[27187]_ , \new_[27188]_ ,
    \new_[27192]_ , \new_[27193]_ , \new_[27197]_ , \new_[27198]_ ,
    \new_[27199]_ , \new_[27203]_ , \new_[27204]_ , \new_[27208]_ ,
    \new_[27209]_ , \new_[27210]_ , \new_[27214]_ , \new_[27215]_ ,
    \new_[27219]_ , \new_[27220]_ , \new_[27221]_ , \new_[27225]_ ,
    \new_[27226]_ , \new_[27230]_ , \new_[27231]_ , \new_[27232]_ ,
    \new_[27236]_ , \new_[27237]_ , \new_[27241]_ , \new_[27242]_ ,
    \new_[27243]_ , \new_[27247]_ , \new_[27248]_ , \new_[27252]_ ,
    \new_[27253]_ , \new_[27254]_ , \new_[27258]_ , \new_[27259]_ ,
    \new_[27263]_ , \new_[27264]_ , \new_[27265]_ , \new_[27269]_ ,
    \new_[27270]_ , \new_[27274]_ , \new_[27275]_ , \new_[27276]_ ,
    \new_[27280]_ , \new_[27281]_ , \new_[27285]_ , \new_[27286]_ ,
    \new_[27287]_ , \new_[27291]_ , \new_[27292]_ , \new_[27296]_ ,
    \new_[27297]_ , \new_[27298]_ , \new_[27302]_ , \new_[27303]_ ,
    \new_[27307]_ , \new_[27308]_ , \new_[27309]_ , \new_[27313]_ ,
    \new_[27314]_ , \new_[27318]_ , \new_[27319]_ , \new_[27320]_ ,
    \new_[27324]_ , \new_[27325]_ , \new_[27329]_ , \new_[27330]_ ,
    \new_[27331]_ , \new_[27335]_ , \new_[27336]_ , \new_[27340]_ ,
    \new_[27341]_ , \new_[27342]_ , \new_[27346]_ , \new_[27347]_ ,
    \new_[27351]_ , \new_[27352]_ , \new_[27353]_ , \new_[27357]_ ,
    \new_[27358]_ , \new_[27362]_ , \new_[27363]_ , \new_[27364]_ ,
    \new_[27368]_ , \new_[27369]_ , \new_[27373]_ , \new_[27374]_ ,
    \new_[27375]_ , \new_[27379]_ , \new_[27380]_ , \new_[27384]_ ,
    \new_[27385]_ , \new_[27386]_ , \new_[27390]_ , \new_[27391]_ ,
    \new_[27395]_ , \new_[27396]_ , \new_[27397]_ , \new_[27401]_ ,
    \new_[27402]_ , \new_[27406]_ , \new_[27407]_ , \new_[27408]_ ,
    \new_[27412]_ , \new_[27413]_ , \new_[27417]_ , \new_[27418]_ ,
    \new_[27419]_ , \new_[27423]_ , \new_[27424]_ , \new_[27428]_ ,
    \new_[27429]_ , \new_[27430]_ , \new_[27434]_ , \new_[27435]_ ,
    \new_[27439]_ , \new_[27440]_ , \new_[27441]_ , \new_[27445]_ ,
    \new_[27446]_ , \new_[27450]_ , \new_[27451]_ , \new_[27452]_ ,
    \new_[27456]_ , \new_[27457]_ , \new_[27461]_ , \new_[27462]_ ,
    \new_[27463]_ , \new_[27467]_ , \new_[27468]_ , \new_[27472]_ ,
    \new_[27473]_ , \new_[27474]_ , \new_[27478]_ , \new_[27479]_ ,
    \new_[27483]_ , \new_[27484]_ , \new_[27485]_ , \new_[27489]_ ,
    \new_[27490]_ , \new_[27494]_ , \new_[27495]_ , \new_[27496]_ ,
    \new_[27500]_ , \new_[27501]_ , \new_[27505]_ , \new_[27506]_ ,
    \new_[27507]_ , \new_[27511]_ , \new_[27512]_ , \new_[27516]_ ,
    \new_[27517]_ , \new_[27518]_ , \new_[27522]_ , \new_[27523]_ ,
    \new_[27527]_ , \new_[27528]_ , \new_[27529]_ , \new_[27533]_ ,
    \new_[27534]_ , \new_[27538]_ , \new_[27539]_ , \new_[27540]_ ,
    \new_[27544]_ , \new_[27545]_ , \new_[27549]_ , \new_[27550]_ ,
    \new_[27551]_ , \new_[27555]_ , \new_[27556]_ , \new_[27560]_ ,
    \new_[27561]_ , \new_[27562]_ , \new_[27566]_ , \new_[27567]_ ,
    \new_[27571]_ , \new_[27572]_ , \new_[27573]_ , \new_[27577]_ ,
    \new_[27578]_ , \new_[27582]_ , \new_[27583]_ , \new_[27584]_ ,
    \new_[27588]_ , \new_[27589]_ , \new_[27593]_ , \new_[27594]_ ,
    \new_[27595]_ , \new_[27599]_ , \new_[27600]_ , \new_[27604]_ ,
    \new_[27605]_ , \new_[27606]_ , \new_[27610]_ , \new_[27611]_ ,
    \new_[27615]_ , \new_[27616]_ , \new_[27617]_ , \new_[27621]_ ,
    \new_[27622]_ , \new_[27626]_ , \new_[27627]_ , \new_[27628]_ ,
    \new_[27632]_ , \new_[27633]_ , \new_[27637]_ , \new_[27638]_ ,
    \new_[27639]_ , \new_[27643]_ , \new_[27644]_ , \new_[27648]_ ,
    \new_[27649]_ , \new_[27650]_ , \new_[27654]_ , \new_[27655]_ ,
    \new_[27659]_ , \new_[27660]_ , \new_[27661]_ , \new_[27665]_ ,
    \new_[27666]_ , \new_[27670]_ , \new_[27671]_ , \new_[27672]_ ,
    \new_[27676]_ , \new_[27677]_ , \new_[27681]_ , \new_[27682]_ ,
    \new_[27683]_ , \new_[27687]_ , \new_[27688]_ , \new_[27692]_ ,
    \new_[27693]_ , \new_[27694]_ , \new_[27698]_ , \new_[27699]_ ,
    \new_[27703]_ , \new_[27704]_ , \new_[27705]_ , \new_[27709]_ ,
    \new_[27710]_ , \new_[27714]_ , \new_[27715]_ , \new_[27716]_ ,
    \new_[27720]_ , \new_[27721]_ , \new_[27725]_ , \new_[27726]_ ,
    \new_[27727]_ , \new_[27731]_ , \new_[27732]_ , \new_[27736]_ ,
    \new_[27737]_ , \new_[27738]_ , \new_[27742]_ , \new_[27743]_ ,
    \new_[27747]_ , \new_[27748]_ , \new_[27749]_ , \new_[27753]_ ,
    \new_[27754]_ , \new_[27758]_ , \new_[27759]_ , \new_[27760]_ ,
    \new_[27764]_ , \new_[27765]_ , \new_[27769]_ , \new_[27770]_ ,
    \new_[27771]_ , \new_[27775]_ , \new_[27776]_ , \new_[27780]_ ,
    \new_[27781]_ , \new_[27782]_ , \new_[27786]_ , \new_[27787]_ ,
    \new_[27791]_ , \new_[27792]_ , \new_[27793]_ , \new_[27797]_ ,
    \new_[27798]_ , \new_[27802]_ , \new_[27803]_ , \new_[27804]_ ,
    \new_[27808]_ , \new_[27809]_ , \new_[27813]_ , \new_[27814]_ ,
    \new_[27815]_ , \new_[27819]_ , \new_[27820]_ , \new_[27824]_ ,
    \new_[27825]_ , \new_[27826]_ , \new_[27830]_ , \new_[27831]_ ,
    \new_[27835]_ , \new_[27836]_ , \new_[27837]_ , \new_[27841]_ ,
    \new_[27842]_ , \new_[27846]_ , \new_[27847]_ , \new_[27848]_ ,
    \new_[27852]_ , \new_[27853]_ , \new_[27857]_ , \new_[27858]_ ,
    \new_[27859]_ , \new_[27863]_ , \new_[27864]_ , \new_[27868]_ ,
    \new_[27869]_ , \new_[27870]_ , \new_[27874]_ , \new_[27875]_ ,
    \new_[27879]_ , \new_[27880]_ , \new_[27881]_ , \new_[27885]_ ,
    \new_[27886]_ , \new_[27890]_ , \new_[27891]_ , \new_[27892]_ ,
    \new_[27896]_ , \new_[27897]_ , \new_[27901]_ , \new_[27902]_ ,
    \new_[27903]_ , \new_[27907]_ , \new_[27908]_ , \new_[27912]_ ,
    \new_[27913]_ , \new_[27914]_ , \new_[27918]_ , \new_[27919]_ ,
    \new_[27923]_ , \new_[27924]_ , \new_[27925]_ , \new_[27929]_ ,
    \new_[27930]_ , \new_[27934]_ , \new_[27935]_ , \new_[27936]_ ,
    \new_[27940]_ , \new_[27941]_ , \new_[27945]_ , \new_[27946]_ ,
    \new_[27947]_ , \new_[27951]_ , \new_[27952]_ , \new_[27956]_ ,
    \new_[27957]_ , \new_[27958]_ , \new_[27962]_ , \new_[27963]_ ,
    \new_[27967]_ , \new_[27968]_ , \new_[27969]_ , \new_[27973]_ ,
    \new_[27974]_ , \new_[27978]_ , \new_[27979]_ , \new_[27980]_ ,
    \new_[27984]_ , \new_[27985]_ , \new_[27989]_ , \new_[27990]_ ,
    \new_[27991]_ , \new_[27995]_ , \new_[27996]_ , \new_[28000]_ ,
    \new_[28001]_ , \new_[28002]_ , \new_[28006]_ , \new_[28007]_ ,
    \new_[28011]_ , \new_[28012]_ , \new_[28013]_ , \new_[28017]_ ,
    \new_[28018]_ , \new_[28022]_ , \new_[28023]_ , \new_[28024]_ ,
    \new_[28028]_ , \new_[28029]_ , \new_[28033]_ , \new_[28034]_ ,
    \new_[28035]_ , \new_[28039]_ , \new_[28040]_ , \new_[28044]_ ,
    \new_[28045]_ , \new_[28046]_ , \new_[28050]_ , \new_[28051]_ ,
    \new_[28055]_ , \new_[28056]_ , \new_[28057]_ , \new_[28061]_ ,
    \new_[28062]_ , \new_[28066]_ , \new_[28067]_ , \new_[28068]_ ,
    \new_[28072]_ , \new_[28073]_ , \new_[28077]_ , \new_[28078]_ ,
    \new_[28079]_ , \new_[28083]_ , \new_[28084]_ , \new_[28088]_ ,
    \new_[28089]_ , \new_[28090]_ , \new_[28094]_ , \new_[28095]_ ,
    \new_[28099]_ , \new_[28100]_ , \new_[28101]_ , \new_[28105]_ ,
    \new_[28106]_ , \new_[28110]_ , \new_[28111]_ , \new_[28112]_ ,
    \new_[28116]_ , \new_[28117]_ , \new_[28121]_ , \new_[28122]_ ,
    \new_[28123]_ , \new_[28127]_ , \new_[28128]_ , \new_[28132]_ ,
    \new_[28133]_ , \new_[28134]_ , \new_[28138]_ , \new_[28139]_ ,
    \new_[28143]_ , \new_[28144]_ , \new_[28145]_ , \new_[28149]_ ,
    \new_[28150]_ , \new_[28154]_ , \new_[28155]_ , \new_[28156]_ ,
    \new_[28160]_ , \new_[28161]_ , \new_[28165]_ , \new_[28166]_ ,
    \new_[28167]_ , \new_[28171]_ , \new_[28172]_ , \new_[28176]_ ,
    \new_[28177]_ , \new_[28178]_ , \new_[28182]_ , \new_[28183]_ ,
    \new_[28187]_ , \new_[28188]_ , \new_[28189]_ , \new_[28193]_ ,
    \new_[28194]_ , \new_[28198]_ , \new_[28199]_ , \new_[28200]_ ,
    \new_[28204]_ , \new_[28205]_ , \new_[28209]_ , \new_[28210]_ ,
    \new_[28211]_ , \new_[28215]_ , \new_[28216]_ , \new_[28220]_ ,
    \new_[28221]_ , \new_[28222]_ , \new_[28226]_ , \new_[28227]_ ,
    \new_[28231]_ , \new_[28232]_ , \new_[28233]_ , \new_[28237]_ ,
    \new_[28238]_ , \new_[28242]_ , \new_[28243]_ , \new_[28244]_ ,
    \new_[28248]_ , \new_[28249]_ , \new_[28253]_ , \new_[28254]_ ,
    \new_[28255]_ , \new_[28259]_ , \new_[28260]_ , \new_[28264]_ ,
    \new_[28265]_ , \new_[28266]_ , \new_[28270]_ , \new_[28271]_ ,
    \new_[28275]_ , \new_[28276]_ , \new_[28277]_ , \new_[28281]_ ,
    \new_[28282]_ , \new_[28286]_ , \new_[28287]_ , \new_[28288]_ ,
    \new_[28292]_ , \new_[28293]_ , \new_[28297]_ , \new_[28298]_ ,
    \new_[28299]_ , \new_[28303]_ , \new_[28304]_ , \new_[28308]_ ,
    \new_[28309]_ , \new_[28310]_ , \new_[28314]_ , \new_[28315]_ ,
    \new_[28319]_ , \new_[28320]_ , \new_[28321]_ , \new_[28325]_ ,
    \new_[28326]_ , \new_[28330]_ , \new_[28331]_ , \new_[28332]_ ,
    \new_[28336]_ , \new_[28337]_ , \new_[28341]_ , \new_[28342]_ ,
    \new_[28343]_ , \new_[28347]_ , \new_[28348]_ , \new_[28352]_ ,
    \new_[28353]_ , \new_[28354]_ , \new_[28358]_ , \new_[28359]_ ,
    \new_[28363]_ , \new_[28364]_ , \new_[28365]_ , \new_[28369]_ ,
    \new_[28370]_ , \new_[28374]_ , \new_[28375]_ , \new_[28376]_ ,
    \new_[28380]_ , \new_[28381]_ , \new_[28385]_ , \new_[28386]_ ,
    \new_[28387]_ , \new_[28391]_ , \new_[28392]_ , \new_[28396]_ ,
    \new_[28397]_ , \new_[28398]_ , \new_[28402]_ , \new_[28403]_ ,
    \new_[28407]_ , \new_[28408]_ , \new_[28409]_ , \new_[28413]_ ,
    \new_[28414]_ , \new_[28418]_ , \new_[28419]_ , \new_[28420]_ ,
    \new_[28424]_ , \new_[28425]_ , \new_[28429]_ , \new_[28430]_ ,
    \new_[28431]_ , \new_[28435]_ , \new_[28436]_ , \new_[28440]_ ,
    \new_[28441]_ , \new_[28442]_ , \new_[28446]_ , \new_[28447]_ ,
    \new_[28451]_ , \new_[28452]_ , \new_[28453]_ , \new_[28457]_ ,
    \new_[28458]_ , \new_[28462]_ , \new_[28463]_ , \new_[28464]_ ,
    \new_[28468]_ , \new_[28469]_ , \new_[28473]_ , \new_[28474]_ ,
    \new_[28475]_ , \new_[28479]_ , \new_[28480]_ , \new_[28484]_ ,
    \new_[28485]_ , \new_[28486]_ , \new_[28490]_ , \new_[28491]_ ,
    \new_[28495]_ , \new_[28496]_ , \new_[28497]_ , \new_[28501]_ ,
    \new_[28502]_ , \new_[28506]_ , \new_[28507]_ , \new_[28508]_ ,
    \new_[28512]_ , \new_[28513]_ , \new_[28517]_ , \new_[28518]_ ,
    \new_[28519]_ , \new_[28523]_ , \new_[28524]_ , \new_[28528]_ ,
    \new_[28529]_ , \new_[28530]_ , \new_[28534]_ , \new_[28535]_ ,
    \new_[28539]_ , \new_[28540]_ , \new_[28541]_ , \new_[28545]_ ,
    \new_[28546]_ , \new_[28550]_ , \new_[28551]_ , \new_[28552]_ ,
    \new_[28556]_ , \new_[28557]_ , \new_[28561]_ , \new_[28562]_ ,
    \new_[28563]_ , \new_[28567]_ , \new_[28568]_ , \new_[28572]_ ,
    \new_[28573]_ , \new_[28574]_ , \new_[28578]_ , \new_[28579]_ ,
    \new_[28583]_ , \new_[28584]_ , \new_[28585]_ , \new_[28589]_ ,
    \new_[28590]_ , \new_[28594]_ , \new_[28595]_ , \new_[28596]_ ,
    \new_[28600]_ , \new_[28601]_ , \new_[28605]_ , \new_[28606]_ ,
    \new_[28607]_ , \new_[28611]_ , \new_[28612]_ , \new_[28616]_ ,
    \new_[28617]_ , \new_[28618]_ , \new_[28622]_ , \new_[28623]_ ,
    \new_[28627]_ , \new_[28628]_ , \new_[28629]_ , \new_[28633]_ ,
    \new_[28634]_ , \new_[28638]_ , \new_[28639]_ , \new_[28640]_ ,
    \new_[28644]_ , \new_[28645]_ , \new_[28649]_ , \new_[28650]_ ,
    \new_[28651]_ , \new_[28655]_ , \new_[28656]_ , \new_[28660]_ ,
    \new_[28661]_ , \new_[28662]_ , \new_[28666]_ , \new_[28667]_ ,
    \new_[28671]_ , \new_[28672]_ , \new_[28673]_ , \new_[28677]_ ,
    \new_[28678]_ , \new_[28682]_ , \new_[28683]_ , \new_[28684]_ ,
    \new_[28688]_ , \new_[28689]_ , \new_[28693]_ , \new_[28694]_ ,
    \new_[28695]_ , \new_[28699]_ , \new_[28700]_ , \new_[28704]_ ,
    \new_[28705]_ , \new_[28706]_ , \new_[28710]_ , \new_[28711]_ ,
    \new_[28715]_ , \new_[28716]_ , \new_[28717]_ , \new_[28721]_ ,
    \new_[28722]_ , \new_[28726]_ , \new_[28727]_ , \new_[28728]_ ,
    \new_[28732]_ , \new_[28733]_ , \new_[28737]_ , \new_[28738]_ ,
    \new_[28739]_ , \new_[28743]_ , \new_[28744]_ , \new_[28748]_ ,
    \new_[28749]_ , \new_[28750]_ , \new_[28754]_ , \new_[28755]_ ,
    \new_[28759]_ , \new_[28760]_ , \new_[28761]_ , \new_[28765]_ ,
    \new_[28766]_ , \new_[28770]_ , \new_[28771]_ , \new_[28772]_ ,
    \new_[28776]_ , \new_[28777]_ , \new_[28781]_ , \new_[28782]_ ,
    \new_[28783]_ , \new_[28787]_ , \new_[28788]_ , \new_[28792]_ ,
    \new_[28793]_ , \new_[28794]_ , \new_[28798]_ , \new_[28799]_ ,
    \new_[28803]_ , \new_[28804]_ , \new_[28805]_ , \new_[28809]_ ,
    \new_[28810]_ , \new_[28814]_ , \new_[28815]_ , \new_[28816]_ ,
    \new_[28820]_ , \new_[28821]_ , \new_[28825]_ , \new_[28826]_ ,
    \new_[28827]_ , \new_[28831]_ , \new_[28832]_ , \new_[28836]_ ,
    \new_[28837]_ , \new_[28838]_ , \new_[28842]_ , \new_[28843]_ ,
    \new_[28847]_ , \new_[28848]_ , \new_[28849]_ , \new_[28853]_ ,
    \new_[28854]_ , \new_[28858]_ , \new_[28859]_ , \new_[28860]_ ,
    \new_[28864]_ , \new_[28865]_ , \new_[28869]_ , \new_[28870]_ ,
    \new_[28871]_ , \new_[28875]_ , \new_[28876]_ , \new_[28880]_ ,
    \new_[28881]_ , \new_[28882]_ , \new_[28886]_ , \new_[28887]_ ,
    \new_[28891]_ , \new_[28892]_ , \new_[28893]_ , \new_[28897]_ ,
    \new_[28898]_ , \new_[28902]_ , \new_[28903]_ , \new_[28904]_ ,
    \new_[28908]_ , \new_[28909]_ , \new_[28913]_ , \new_[28914]_ ,
    \new_[28915]_ , \new_[28919]_ , \new_[28920]_ , \new_[28924]_ ,
    \new_[28925]_ , \new_[28926]_ , \new_[28930]_ , \new_[28931]_ ,
    \new_[28935]_ , \new_[28936]_ , \new_[28937]_ , \new_[28941]_ ,
    \new_[28942]_ , \new_[28946]_ , \new_[28947]_ , \new_[28948]_ ,
    \new_[28952]_ , \new_[28953]_ , \new_[28957]_ , \new_[28958]_ ,
    \new_[28959]_ , \new_[28963]_ , \new_[28964]_ , \new_[28968]_ ,
    \new_[28969]_ , \new_[28970]_ , \new_[28974]_ , \new_[28975]_ ,
    \new_[28979]_ , \new_[28980]_ , \new_[28981]_ , \new_[28985]_ ,
    \new_[28986]_ , \new_[28990]_ , \new_[28991]_ , \new_[28992]_ ,
    \new_[28996]_ , \new_[28997]_ , \new_[29001]_ , \new_[29002]_ ,
    \new_[29003]_ , \new_[29007]_ , \new_[29008]_ , \new_[29012]_ ,
    \new_[29013]_ , \new_[29014]_ , \new_[29018]_ , \new_[29019]_ ,
    \new_[29023]_ , \new_[29024]_ , \new_[29025]_ , \new_[29029]_ ,
    \new_[29030]_ , \new_[29034]_ , \new_[29035]_ , \new_[29036]_ ,
    \new_[29040]_ , \new_[29041]_ , \new_[29045]_ , \new_[29046]_ ,
    \new_[29047]_ , \new_[29051]_ , \new_[29052]_ , \new_[29056]_ ,
    \new_[29057]_ , \new_[29058]_ , \new_[29062]_ , \new_[29063]_ ,
    \new_[29067]_ , \new_[29068]_ , \new_[29069]_ , \new_[29073]_ ,
    \new_[29074]_ , \new_[29078]_ , \new_[29079]_ , \new_[29080]_ ,
    \new_[29084]_ , \new_[29085]_ , \new_[29089]_ , \new_[29090]_ ,
    \new_[29091]_ , \new_[29095]_ , \new_[29096]_ , \new_[29100]_ ,
    \new_[29101]_ , \new_[29102]_ , \new_[29106]_ , \new_[29107]_ ,
    \new_[29111]_ , \new_[29112]_ , \new_[29113]_ , \new_[29117]_ ,
    \new_[29118]_ , \new_[29122]_ , \new_[29123]_ , \new_[29124]_ ,
    \new_[29128]_ , \new_[29129]_ , \new_[29133]_ , \new_[29134]_ ,
    \new_[29135]_ , \new_[29139]_ , \new_[29140]_ , \new_[29144]_ ,
    \new_[29145]_ , \new_[29146]_ , \new_[29150]_ , \new_[29151]_ ,
    \new_[29155]_ , \new_[29156]_ , \new_[29157]_ , \new_[29161]_ ,
    \new_[29162]_ , \new_[29166]_ , \new_[29167]_ , \new_[29168]_ ,
    \new_[29172]_ , \new_[29173]_ , \new_[29177]_ , \new_[29178]_ ,
    \new_[29179]_ , \new_[29183]_ , \new_[29184]_ , \new_[29188]_ ,
    \new_[29189]_ , \new_[29190]_ , \new_[29194]_ , \new_[29195]_ ,
    \new_[29199]_ , \new_[29200]_ , \new_[29201]_ , \new_[29205]_ ,
    \new_[29206]_ , \new_[29210]_ , \new_[29211]_ , \new_[29212]_ ,
    \new_[29216]_ , \new_[29217]_ , \new_[29221]_ , \new_[29222]_ ,
    \new_[29223]_ , \new_[29227]_ , \new_[29228]_ , \new_[29232]_ ,
    \new_[29233]_ , \new_[29234]_ , \new_[29238]_ , \new_[29239]_ ,
    \new_[29243]_ , \new_[29244]_ , \new_[29245]_ , \new_[29249]_ ,
    \new_[29250]_ , \new_[29254]_ , \new_[29255]_ , \new_[29256]_ ,
    \new_[29260]_ , \new_[29261]_ , \new_[29265]_ , \new_[29266]_ ,
    \new_[29267]_ , \new_[29271]_ , \new_[29272]_ , \new_[29276]_ ,
    \new_[29277]_ , \new_[29278]_ , \new_[29282]_ , \new_[29283]_ ,
    \new_[29287]_ , \new_[29288]_ , \new_[29289]_ , \new_[29293]_ ,
    \new_[29294]_ , \new_[29298]_ , \new_[29299]_ , \new_[29300]_ ,
    \new_[29304]_ , \new_[29305]_ , \new_[29309]_ , \new_[29310]_ ,
    \new_[29311]_ , \new_[29315]_ , \new_[29316]_ , \new_[29320]_ ,
    \new_[29321]_ , \new_[29322]_ , \new_[29326]_ , \new_[29327]_ ,
    \new_[29331]_ , \new_[29332]_ , \new_[29333]_ , \new_[29337]_ ,
    \new_[29338]_ , \new_[29342]_ , \new_[29343]_ , \new_[29344]_ ,
    \new_[29348]_ , \new_[29349]_ , \new_[29353]_ , \new_[29354]_ ,
    \new_[29355]_ , \new_[29359]_ , \new_[29360]_ , \new_[29364]_ ,
    \new_[29365]_ , \new_[29366]_ , \new_[29370]_ , \new_[29371]_ ,
    \new_[29375]_ , \new_[29376]_ , \new_[29377]_ , \new_[29381]_ ,
    \new_[29382]_ , \new_[29386]_ , \new_[29387]_ , \new_[29388]_ ,
    \new_[29392]_ , \new_[29393]_ , \new_[29397]_ , \new_[29398]_ ,
    \new_[29399]_ , \new_[29403]_ , \new_[29404]_ , \new_[29408]_ ,
    \new_[29409]_ , \new_[29410]_ , \new_[29414]_ , \new_[29415]_ ,
    \new_[29419]_ , \new_[29420]_ , \new_[29421]_ , \new_[29425]_ ,
    \new_[29426]_ , \new_[29430]_ , \new_[29431]_ , \new_[29432]_ ,
    \new_[29436]_ , \new_[29437]_ , \new_[29441]_ , \new_[29442]_ ,
    \new_[29443]_ , \new_[29447]_ , \new_[29448]_ , \new_[29452]_ ,
    \new_[29453]_ , \new_[29454]_ , \new_[29458]_ , \new_[29459]_ ,
    \new_[29463]_ , \new_[29464]_ , \new_[29465]_ , \new_[29469]_ ,
    \new_[29470]_ , \new_[29474]_ , \new_[29475]_ , \new_[29476]_ ,
    \new_[29480]_ , \new_[29481]_ , \new_[29485]_ , \new_[29486]_ ,
    \new_[29487]_ , \new_[29491]_ , \new_[29492]_ , \new_[29496]_ ,
    \new_[29497]_ , \new_[29498]_ , \new_[29502]_ , \new_[29503]_ ,
    \new_[29507]_ , \new_[29508]_ , \new_[29509]_ , \new_[29513]_ ,
    \new_[29514]_ , \new_[29518]_ , \new_[29519]_ , \new_[29520]_ ,
    \new_[29524]_ , \new_[29525]_ , \new_[29529]_ , \new_[29530]_ ,
    \new_[29531]_ , \new_[29535]_ , \new_[29536]_ , \new_[29540]_ ,
    \new_[29541]_ , \new_[29542]_ , \new_[29546]_ , \new_[29547]_ ,
    \new_[29551]_ , \new_[29552]_ , \new_[29553]_ , \new_[29557]_ ,
    \new_[29558]_ , \new_[29562]_ , \new_[29563]_ , \new_[29564]_ ,
    \new_[29568]_ , \new_[29569]_ , \new_[29573]_ , \new_[29574]_ ,
    \new_[29575]_ , \new_[29579]_ , \new_[29580]_ , \new_[29584]_ ,
    \new_[29585]_ , \new_[29586]_ , \new_[29590]_ , \new_[29591]_ ,
    \new_[29595]_ , \new_[29596]_ , \new_[29597]_ , \new_[29601]_ ,
    \new_[29602]_ , \new_[29606]_ , \new_[29607]_ , \new_[29608]_ ,
    \new_[29612]_ , \new_[29613]_ , \new_[29617]_ , \new_[29618]_ ,
    \new_[29619]_ , \new_[29623]_ , \new_[29624]_ , \new_[29628]_ ,
    \new_[29629]_ , \new_[29630]_ , \new_[29634]_ , \new_[29635]_ ,
    \new_[29639]_ , \new_[29640]_ , \new_[29641]_ , \new_[29645]_ ,
    \new_[29646]_ , \new_[29650]_ , \new_[29651]_ , \new_[29652]_ ,
    \new_[29656]_ , \new_[29657]_ , \new_[29661]_ , \new_[29662]_ ,
    \new_[29663]_ , \new_[29667]_ , \new_[29668]_ , \new_[29672]_ ,
    \new_[29673]_ , \new_[29674]_ , \new_[29678]_ , \new_[29679]_ ,
    \new_[29683]_ , \new_[29684]_ , \new_[29685]_ , \new_[29689]_ ,
    \new_[29690]_ , \new_[29694]_ , \new_[29695]_ , \new_[29696]_ ,
    \new_[29700]_ , \new_[29701]_ , \new_[29705]_ , \new_[29706]_ ,
    \new_[29707]_ , \new_[29711]_ , \new_[29712]_ , \new_[29716]_ ,
    \new_[29717]_ , \new_[29718]_ , \new_[29722]_ , \new_[29723]_ ,
    \new_[29727]_ , \new_[29728]_ , \new_[29729]_ , \new_[29733]_ ,
    \new_[29734]_ , \new_[29738]_ , \new_[29739]_ , \new_[29740]_ ,
    \new_[29744]_ , \new_[29745]_ , \new_[29749]_ , \new_[29750]_ ,
    \new_[29751]_ , \new_[29755]_ , \new_[29756]_ , \new_[29760]_ ,
    \new_[29761]_ , \new_[29762]_ , \new_[29766]_ , \new_[29767]_ ,
    \new_[29771]_ , \new_[29772]_ , \new_[29773]_ , \new_[29777]_ ,
    \new_[29778]_ , \new_[29782]_ , \new_[29783]_ , \new_[29784]_ ,
    \new_[29788]_ , \new_[29789]_ , \new_[29793]_ , \new_[29794]_ ,
    \new_[29795]_ , \new_[29799]_ , \new_[29800]_ , \new_[29804]_ ,
    \new_[29805]_ , \new_[29806]_ , \new_[29810]_ , \new_[29811]_ ,
    \new_[29815]_ , \new_[29816]_ , \new_[29817]_ , \new_[29821]_ ,
    \new_[29822]_ , \new_[29826]_ , \new_[29827]_ , \new_[29828]_ ,
    \new_[29832]_ , \new_[29833]_ , \new_[29837]_ , \new_[29838]_ ,
    \new_[29839]_ , \new_[29843]_ , \new_[29844]_ , \new_[29848]_ ,
    \new_[29849]_ , \new_[29850]_ , \new_[29854]_ , \new_[29855]_ ,
    \new_[29859]_ , \new_[29860]_ , \new_[29861]_ , \new_[29865]_ ,
    \new_[29866]_ , \new_[29870]_ , \new_[29871]_ , \new_[29872]_ ,
    \new_[29876]_ , \new_[29877]_ , \new_[29881]_ , \new_[29882]_ ,
    \new_[29883]_ , \new_[29887]_ , \new_[29888]_ , \new_[29892]_ ,
    \new_[29893]_ , \new_[29894]_ , \new_[29898]_ , \new_[29899]_ ,
    \new_[29903]_ , \new_[29904]_ , \new_[29905]_ , \new_[29909]_ ,
    \new_[29910]_ , \new_[29914]_ , \new_[29915]_ , \new_[29916]_ ,
    \new_[29920]_ , \new_[29921]_ , \new_[29925]_ , \new_[29926]_ ,
    \new_[29927]_ , \new_[29931]_ , \new_[29932]_ , \new_[29936]_ ,
    \new_[29937]_ , \new_[29938]_ , \new_[29942]_ , \new_[29943]_ ,
    \new_[29947]_ , \new_[29948]_ , \new_[29949]_ , \new_[29953]_ ,
    \new_[29954]_ , \new_[29958]_ , \new_[29959]_ , \new_[29960]_ ,
    \new_[29964]_ , \new_[29965]_ , \new_[29969]_ , \new_[29970]_ ,
    \new_[29971]_ , \new_[29975]_ , \new_[29976]_ , \new_[29980]_ ,
    \new_[29981]_ , \new_[29982]_ , \new_[29986]_ , \new_[29987]_ ,
    \new_[29991]_ , \new_[29992]_ , \new_[29993]_ , \new_[29997]_ ,
    \new_[29998]_ , \new_[30002]_ , \new_[30003]_ , \new_[30004]_ ,
    \new_[30008]_ , \new_[30009]_ , \new_[30013]_ , \new_[30014]_ ,
    \new_[30015]_ , \new_[30019]_ , \new_[30020]_ , \new_[30024]_ ,
    \new_[30025]_ , \new_[30026]_ , \new_[30030]_ , \new_[30031]_ ,
    \new_[30035]_ , \new_[30036]_ , \new_[30037]_ , \new_[30041]_ ,
    \new_[30042]_ , \new_[30046]_ , \new_[30047]_ , \new_[30048]_ ,
    \new_[30052]_ , \new_[30053]_ , \new_[30057]_ , \new_[30058]_ ,
    \new_[30059]_ , \new_[30063]_ , \new_[30064]_ , \new_[30068]_ ,
    \new_[30069]_ , \new_[30070]_ , \new_[30074]_ , \new_[30075]_ ,
    \new_[30079]_ , \new_[30080]_ , \new_[30081]_ , \new_[30085]_ ,
    \new_[30086]_ , \new_[30090]_ , \new_[30091]_ , \new_[30092]_ ,
    \new_[30096]_ , \new_[30097]_ , \new_[30101]_ , \new_[30102]_ ,
    \new_[30103]_ , \new_[30107]_ , \new_[30108]_ , \new_[30112]_ ,
    \new_[30113]_ , \new_[30114]_ , \new_[30118]_ , \new_[30119]_ ,
    \new_[30123]_ , \new_[30124]_ , \new_[30125]_ , \new_[30129]_ ,
    \new_[30130]_ , \new_[30134]_ , \new_[30135]_ , \new_[30136]_ ,
    \new_[30140]_ , \new_[30141]_ , \new_[30145]_ , \new_[30146]_ ,
    \new_[30147]_ , \new_[30151]_ , \new_[30152]_ , \new_[30156]_ ,
    \new_[30157]_ , \new_[30158]_ , \new_[30162]_ , \new_[30163]_ ,
    \new_[30167]_ , \new_[30168]_ , \new_[30169]_ , \new_[30173]_ ,
    \new_[30174]_ , \new_[30178]_ , \new_[30179]_ , \new_[30180]_ ,
    \new_[30184]_ , \new_[30185]_ , \new_[30189]_ , \new_[30190]_ ,
    \new_[30191]_ , \new_[30195]_ , \new_[30196]_ , \new_[30200]_ ,
    \new_[30201]_ , \new_[30202]_ , \new_[30206]_ , \new_[30207]_ ,
    \new_[30211]_ , \new_[30212]_ , \new_[30213]_ , \new_[30217]_ ,
    \new_[30218]_ , \new_[30222]_ , \new_[30223]_ , \new_[30224]_ ,
    \new_[30228]_ , \new_[30229]_ , \new_[30233]_ , \new_[30234]_ ,
    \new_[30235]_ , \new_[30239]_ , \new_[30240]_ , \new_[30244]_ ,
    \new_[30245]_ , \new_[30246]_ , \new_[30250]_ , \new_[30251]_ ,
    \new_[30255]_ , \new_[30256]_ , \new_[30257]_ , \new_[30261]_ ,
    \new_[30262]_ , \new_[30266]_ , \new_[30267]_ , \new_[30268]_ ,
    \new_[30272]_ , \new_[30273]_ , \new_[30277]_ , \new_[30278]_ ,
    \new_[30279]_ , \new_[30283]_ , \new_[30284]_ , \new_[30288]_ ,
    \new_[30289]_ , \new_[30290]_ , \new_[30294]_ , \new_[30295]_ ,
    \new_[30299]_ , \new_[30300]_ , \new_[30301]_ , \new_[30305]_ ,
    \new_[30306]_ , \new_[30310]_ , \new_[30311]_ , \new_[30312]_ ,
    \new_[30316]_ , \new_[30317]_ , \new_[30321]_ , \new_[30322]_ ,
    \new_[30323]_ , \new_[30327]_ , \new_[30328]_ , \new_[30332]_ ,
    \new_[30333]_ , \new_[30334]_ , \new_[30338]_ , \new_[30339]_ ,
    \new_[30343]_ , \new_[30344]_ , \new_[30345]_ , \new_[30349]_ ,
    \new_[30350]_ , \new_[30354]_ , \new_[30355]_ , \new_[30356]_ ,
    \new_[30360]_ , \new_[30361]_ , \new_[30365]_ , \new_[30366]_ ,
    \new_[30367]_ , \new_[30371]_ , \new_[30372]_ , \new_[30376]_ ,
    \new_[30377]_ , \new_[30378]_ , \new_[30382]_ , \new_[30383]_ ,
    \new_[30387]_ , \new_[30388]_ , \new_[30389]_ , \new_[30393]_ ,
    \new_[30394]_ , \new_[30398]_ , \new_[30399]_ , \new_[30400]_ ,
    \new_[30404]_ , \new_[30405]_ , \new_[30409]_ , \new_[30410]_ ,
    \new_[30411]_ , \new_[30415]_ , \new_[30416]_ , \new_[30420]_ ,
    \new_[30421]_ , \new_[30422]_ , \new_[30426]_ , \new_[30427]_ ,
    \new_[30431]_ , \new_[30432]_ , \new_[30433]_ , \new_[30437]_ ,
    \new_[30438]_ , \new_[30442]_ , \new_[30443]_ , \new_[30444]_ ,
    \new_[30448]_ , \new_[30449]_ , \new_[30453]_ , \new_[30454]_ ,
    \new_[30455]_ , \new_[30459]_ , \new_[30460]_ , \new_[30464]_ ,
    \new_[30465]_ , \new_[30466]_ , \new_[30470]_ , \new_[30471]_ ,
    \new_[30475]_ , \new_[30476]_ , \new_[30477]_ , \new_[30481]_ ,
    \new_[30482]_ , \new_[30486]_ , \new_[30487]_ , \new_[30488]_ ,
    \new_[30492]_ , \new_[30493]_ , \new_[30497]_ , \new_[30498]_ ,
    \new_[30499]_ , \new_[30503]_ , \new_[30504]_ , \new_[30508]_ ,
    \new_[30509]_ , \new_[30510]_ , \new_[30514]_ , \new_[30515]_ ,
    \new_[30519]_ , \new_[30520]_ , \new_[30521]_ , \new_[30525]_ ,
    \new_[30526]_ , \new_[30530]_ , \new_[30531]_ , \new_[30532]_ ,
    \new_[30536]_ , \new_[30537]_ , \new_[30541]_ , \new_[30542]_ ,
    \new_[30543]_ , \new_[30547]_ , \new_[30548]_ , \new_[30552]_ ,
    \new_[30553]_ , \new_[30554]_ , \new_[30558]_ , \new_[30559]_ ,
    \new_[30563]_ , \new_[30564]_ , \new_[30565]_ , \new_[30569]_ ,
    \new_[30570]_ , \new_[30574]_ , \new_[30575]_ , \new_[30576]_ ,
    \new_[30580]_ , \new_[30581]_ , \new_[30585]_ , \new_[30586]_ ,
    \new_[30587]_ , \new_[30591]_ , \new_[30592]_ , \new_[30596]_ ,
    \new_[30597]_ , \new_[30598]_ , \new_[30602]_ , \new_[30603]_ ,
    \new_[30607]_ , \new_[30608]_ , \new_[30609]_ , \new_[30613]_ ,
    \new_[30614]_ , \new_[30618]_ , \new_[30619]_ , \new_[30620]_ ,
    \new_[30624]_ , \new_[30625]_ , \new_[30629]_ , \new_[30630]_ ,
    \new_[30631]_ , \new_[30635]_ , \new_[30636]_ , \new_[30639]_ ,
    \new_[30642]_ , \new_[30643]_ , \new_[30644]_ , \new_[30648]_ ,
    \new_[30649]_ , \new_[30653]_ , \new_[30654]_ , \new_[30655]_ ,
    \new_[30659]_ , \new_[30660]_ , \new_[30663]_ , \new_[30666]_ ,
    \new_[30667]_ , \new_[30668]_ , \new_[30672]_ , \new_[30673]_ ,
    \new_[30677]_ , \new_[30678]_ , \new_[30679]_ , \new_[30683]_ ,
    \new_[30684]_ , \new_[30687]_ , \new_[30690]_ , \new_[30691]_ ,
    \new_[30692]_ , \new_[30696]_ , \new_[30697]_ , \new_[30701]_ ,
    \new_[30702]_ , \new_[30703]_ , \new_[30707]_ , \new_[30708]_ ,
    \new_[30711]_ , \new_[30714]_ , \new_[30715]_ , \new_[30716]_ ,
    \new_[30720]_ , \new_[30721]_ , \new_[30725]_ , \new_[30726]_ ,
    \new_[30727]_ , \new_[30731]_ , \new_[30732]_ , \new_[30735]_ ,
    \new_[30738]_ , \new_[30739]_ , \new_[30740]_ , \new_[30744]_ ,
    \new_[30745]_ , \new_[30749]_ , \new_[30750]_ , \new_[30751]_ ,
    \new_[30755]_ , \new_[30756]_ , \new_[30759]_ , \new_[30762]_ ,
    \new_[30763]_ , \new_[30764]_ , \new_[30768]_ , \new_[30769]_ ,
    \new_[30773]_ , \new_[30774]_ , \new_[30775]_ , \new_[30779]_ ,
    \new_[30780]_ , \new_[30783]_ , \new_[30786]_ , \new_[30787]_ ,
    \new_[30788]_ , \new_[30792]_ , \new_[30793]_ , \new_[30797]_ ,
    \new_[30798]_ , \new_[30799]_ , \new_[30803]_ , \new_[30804]_ ,
    \new_[30807]_ , \new_[30810]_ , \new_[30811]_ , \new_[30812]_ ,
    \new_[30816]_ , \new_[30817]_ , \new_[30821]_ , \new_[30822]_ ,
    \new_[30823]_ , \new_[30827]_ , \new_[30828]_ , \new_[30831]_ ,
    \new_[30834]_ , \new_[30835]_ , \new_[30836]_ , \new_[30840]_ ,
    \new_[30841]_ , \new_[30845]_ , \new_[30846]_ , \new_[30847]_ ,
    \new_[30851]_ , \new_[30852]_ , \new_[30855]_ , \new_[30858]_ ,
    \new_[30859]_ , \new_[30860]_ , \new_[30864]_ , \new_[30865]_ ,
    \new_[30869]_ , \new_[30870]_ , \new_[30871]_ , \new_[30875]_ ,
    \new_[30876]_ , \new_[30879]_ , \new_[30882]_ , \new_[30883]_ ,
    \new_[30884]_ , \new_[30888]_ , \new_[30889]_ , \new_[30893]_ ,
    \new_[30894]_ , \new_[30895]_ , \new_[30899]_ , \new_[30900]_ ,
    \new_[30903]_ , \new_[30906]_ , \new_[30907]_ , \new_[30908]_ ,
    \new_[30912]_ , \new_[30913]_ , \new_[30917]_ , \new_[30918]_ ,
    \new_[30919]_ , \new_[30923]_ , \new_[30924]_ , \new_[30927]_ ,
    \new_[30930]_ , \new_[30931]_ , \new_[30932]_ , \new_[30936]_ ,
    \new_[30937]_ , \new_[30941]_ , \new_[30942]_ , \new_[30943]_ ,
    \new_[30947]_ , \new_[30948]_ , \new_[30951]_ , \new_[30954]_ ,
    \new_[30955]_ , \new_[30956]_ , \new_[30960]_ , \new_[30961]_ ,
    \new_[30965]_ , \new_[30966]_ , \new_[30967]_ , \new_[30971]_ ,
    \new_[30972]_ , \new_[30975]_ , \new_[30978]_ , \new_[30979]_ ,
    \new_[30980]_ , \new_[30984]_ , \new_[30985]_ , \new_[30989]_ ,
    \new_[30990]_ , \new_[30991]_ , \new_[30995]_ , \new_[30996]_ ,
    \new_[30999]_ , \new_[31002]_ , \new_[31003]_ , \new_[31004]_ ,
    \new_[31008]_ , \new_[31009]_ , \new_[31013]_ , \new_[31014]_ ,
    \new_[31015]_ , \new_[31019]_ , \new_[31020]_ , \new_[31023]_ ,
    \new_[31026]_ , \new_[31027]_ , \new_[31028]_ , \new_[31032]_ ,
    \new_[31033]_ , \new_[31037]_ , \new_[31038]_ , \new_[31039]_ ,
    \new_[31043]_ , \new_[31044]_ , \new_[31047]_ , \new_[31050]_ ,
    \new_[31051]_ , \new_[31052]_ , \new_[31056]_ , \new_[31057]_ ,
    \new_[31061]_ , \new_[31062]_ , \new_[31063]_ , \new_[31067]_ ,
    \new_[31068]_ , \new_[31071]_ , \new_[31074]_ , \new_[31075]_ ,
    \new_[31076]_ , \new_[31080]_ , \new_[31081]_ , \new_[31085]_ ,
    \new_[31086]_ , \new_[31087]_ , \new_[31091]_ , \new_[31092]_ ,
    \new_[31095]_ , \new_[31098]_ , \new_[31099]_ , \new_[31100]_ ,
    \new_[31104]_ , \new_[31105]_ , \new_[31109]_ , \new_[31110]_ ,
    \new_[31111]_ , \new_[31115]_ , \new_[31116]_ , \new_[31119]_ ,
    \new_[31122]_ , \new_[31123]_ , \new_[31124]_ , \new_[31128]_ ,
    \new_[31129]_ , \new_[31133]_ , \new_[31134]_ , \new_[31135]_ ,
    \new_[31139]_ , \new_[31140]_ , \new_[31143]_ , \new_[31146]_ ,
    \new_[31147]_ , \new_[31148]_ , \new_[31152]_ , \new_[31153]_ ,
    \new_[31157]_ , \new_[31158]_ , \new_[31159]_ , \new_[31163]_ ,
    \new_[31164]_ , \new_[31167]_ , \new_[31170]_ , \new_[31171]_ ,
    \new_[31172]_ , \new_[31176]_ , \new_[31177]_ , \new_[31181]_ ,
    \new_[31182]_ , \new_[31183]_ , \new_[31187]_ , \new_[31188]_ ,
    \new_[31191]_ , \new_[31194]_ , \new_[31195]_ , \new_[31196]_ ,
    \new_[31200]_ , \new_[31201]_ , \new_[31205]_ , \new_[31206]_ ,
    \new_[31207]_ , \new_[31211]_ , \new_[31212]_ , \new_[31215]_ ,
    \new_[31218]_ , \new_[31219]_ , \new_[31220]_ , \new_[31224]_ ,
    \new_[31225]_ , \new_[31229]_ , \new_[31230]_ , \new_[31231]_ ,
    \new_[31235]_ , \new_[31236]_ , \new_[31239]_ , \new_[31242]_ ,
    \new_[31243]_ , \new_[31244]_ , \new_[31248]_ , \new_[31249]_ ,
    \new_[31253]_ , \new_[31254]_ , \new_[31255]_ , \new_[31259]_ ,
    \new_[31260]_ , \new_[31263]_ , \new_[31266]_ , \new_[31267]_ ,
    \new_[31268]_ , \new_[31272]_ , \new_[31273]_ , \new_[31277]_ ,
    \new_[31278]_ , \new_[31279]_ , \new_[31283]_ , \new_[31284]_ ,
    \new_[31287]_ , \new_[31290]_ , \new_[31291]_ , \new_[31292]_ ,
    \new_[31296]_ , \new_[31297]_ , \new_[31301]_ , \new_[31302]_ ,
    \new_[31303]_ , \new_[31307]_ , \new_[31308]_ , \new_[31311]_ ,
    \new_[31314]_ , \new_[31315]_ , \new_[31316]_ , \new_[31320]_ ,
    \new_[31321]_ , \new_[31325]_ , \new_[31326]_ , \new_[31327]_ ,
    \new_[31331]_ , \new_[31332]_ , \new_[31335]_ , \new_[31338]_ ,
    \new_[31339]_ , \new_[31340]_ , \new_[31344]_ , \new_[31345]_ ,
    \new_[31349]_ , \new_[31350]_ , \new_[31351]_ , \new_[31355]_ ,
    \new_[31356]_ , \new_[31359]_ , \new_[31362]_ , \new_[31363]_ ,
    \new_[31364]_ , \new_[31368]_ , \new_[31369]_ , \new_[31373]_ ,
    \new_[31374]_ , \new_[31375]_ , \new_[31379]_ , \new_[31380]_ ,
    \new_[31383]_ , \new_[31386]_ , \new_[31387]_ , \new_[31388]_ ,
    \new_[31392]_ , \new_[31393]_ , \new_[31397]_ , \new_[31398]_ ,
    \new_[31399]_ , \new_[31403]_ , \new_[31404]_ , \new_[31407]_ ,
    \new_[31410]_ , \new_[31411]_ , \new_[31412]_ , \new_[31416]_ ,
    \new_[31417]_ , \new_[31421]_ , \new_[31422]_ , \new_[31423]_ ,
    \new_[31427]_ , \new_[31428]_ , \new_[31431]_ , \new_[31434]_ ,
    \new_[31435]_ , \new_[31436]_ , \new_[31440]_ , \new_[31441]_ ,
    \new_[31445]_ , \new_[31446]_ , \new_[31447]_ , \new_[31451]_ ,
    \new_[31452]_ , \new_[31455]_ , \new_[31458]_ , \new_[31459]_ ,
    \new_[31460]_ , \new_[31464]_ , \new_[31465]_ , \new_[31469]_ ,
    \new_[31470]_ , \new_[31471]_ , \new_[31475]_ , \new_[31476]_ ,
    \new_[31479]_ , \new_[31482]_ , \new_[31483]_ , \new_[31484]_ ,
    \new_[31488]_ , \new_[31489]_ , \new_[31493]_ , \new_[31494]_ ,
    \new_[31495]_ , \new_[31499]_ , \new_[31500]_ , \new_[31503]_ ,
    \new_[31506]_ , \new_[31507]_ , \new_[31508]_ , \new_[31512]_ ,
    \new_[31513]_ , \new_[31517]_ , \new_[31518]_ , \new_[31519]_ ,
    \new_[31523]_ , \new_[31524]_ , \new_[31527]_ , \new_[31530]_ ,
    \new_[31531]_ , \new_[31532]_ , \new_[31536]_ , \new_[31537]_ ,
    \new_[31541]_ , \new_[31542]_ , \new_[31543]_ , \new_[31547]_ ,
    \new_[31548]_ , \new_[31551]_ , \new_[31554]_ , \new_[31555]_ ,
    \new_[31556]_ , \new_[31560]_ , \new_[31561]_ , \new_[31565]_ ,
    \new_[31566]_ , \new_[31567]_ , \new_[31571]_ , \new_[31572]_ ,
    \new_[31575]_ , \new_[31578]_ , \new_[31579]_ , \new_[31580]_ ,
    \new_[31584]_ , \new_[31585]_ , \new_[31589]_ , \new_[31590]_ ,
    \new_[31591]_ , \new_[31595]_ , \new_[31596]_ , \new_[31599]_ ,
    \new_[31602]_ , \new_[31603]_ , \new_[31604]_ , \new_[31608]_ ,
    \new_[31609]_ , \new_[31613]_ , \new_[31614]_ , \new_[31615]_ ,
    \new_[31619]_ , \new_[31620]_ , \new_[31623]_ , \new_[31626]_ ,
    \new_[31627]_ , \new_[31628]_ , \new_[31632]_ , \new_[31633]_ ,
    \new_[31637]_ , \new_[31638]_ , \new_[31639]_ , \new_[31643]_ ,
    \new_[31644]_ , \new_[31647]_ , \new_[31650]_ , \new_[31651]_ ,
    \new_[31652]_ , \new_[31656]_ , \new_[31657]_ , \new_[31661]_ ,
    \new_[31662]_ , \new_[31663]_ , \new_[31667]_ , \new_[31668]_ ,
    \new_[31671]_ , \new_[31674]_ , \new_[31675]_ , \new_[31676]_ ,
    \new_[31680]_ , \new_[31681]_ , \new_[31685]_ , \new_[31686]_ ,
    \new_[31687]_ , \new_[31691]_ , \new_[31692]_ , \new_[31695]_ ,
    \new_[31698]_ , \new_[31699]_ , \new_[31700]_ , \new_[31704]_ ,
    \new_[31705]_ , \new_[31709]_ , \new_[31710]_ , \new_[31711]_ ,
    \new_[31715]_ , \new_[31716]_ , \new_[31719]_ , \new_[31722]_ ,
    \new_[31723]_ , \new_[31724]_ , \new_[31728]_ , \new_[31729]_ ,
    \new_[31733]_ , \new_[31734]_ , \new_[31735]_ , \new_[31739]_ ,
    \new_[31740]_ , \new_[31743]_ , \new_[31746]_ , \new_[31747]_ ,
    \new_[31748]_ , \new_[31752]_ , \new_[31753]_ , \new_[31757]_ ,
    \new_[31758]_ , \new_[31759]_ , \new_[31763]_ , \new_[31764]_ ,
    \new_[31767]_ , \new_[31770]_ , \new_[31771]_ , \new_[31772]_ ,
    \new_[31776]_ , \new_[31777]_ , \new_[31781]_ , \new_[31782]_ ,
    \new_[31783]_ , \new_[31787]_ , \new_[31788]_ , \new_[31791]_ ,
    \new_[31794]_ , \new_[31795]_ , \new_[31796]_ , \new_[31800]_ ,
    \new_[31801]_ , \new_[31805]_ , \new_[31806]_ , \new_[31807]_ ,
    \new_[31811]_ , \new_[31812]_ , \new_[31815]_ , \new_[31818]_ ,
    \new_[31819]_ , \new_[31820]_ , \new_[31824]_ , \new_[31825]_ ,
    \new_[31829]_ , \new_[31830]_ , \new_[31831]_ , \new_[31835]_ ,
    \new_[31836]_ , \new_[31839]_ , \new_[31842]_ , \new_[31843]_ ,
    \new_[31844]_ , \new_[31848]_ , \new_[31849]_ , \new_[31853]_ ,
    \new_[31854]_ , \new_[31855]_ , \new_[31859]_ , \new_[31860]_ ,
    \new_[31863]_ , \new_[31866]_ , \new_[31867]_ , \new_[31868]_ ,
    \new_[31872]_ , \new_[31873]_ , \new_[31877]_ , \new_[31878]_ ,
    \new_[31879]_ , \new_[31883]_ , \new_[31884]_ , \new_[31887]_ ,
    \new_[31890]_ , \new_[31891]_ , \new_[31892]_ , \new_[31896]_ ,
    \new_[31897]_ , \new_[31901]_ , \new_[31902]_ , \new_[31903]_ ,
    \new_[31907]_ , \new_[31908]_ , \new_[31911]_ , \new_[31914]_ ,
    \new_[31915]_ , \new_[31916]_ , \new_[31920]_ , \new_[31921]_ ,
    \new_[31925]_ , \new_[31926]_ , \new_[31927]_ , \new_[31931]_ ,
    \new_[31932]_ , \new_[31935]_ , \new_[31938]_ , \new_[31939]_ ,
    \new_[31940]_ , \new_[31944]_ , \new_[31945]_ , \new_[31949]_ ,
    \new_[31950]_ , \new_[31951]_ , \new_[31955]_ , \new_[31956]_ ,
    \new_[31959]_ , \new_[31962]_ , \new_[31963]_ , \new_[31964]_ ,
    \new_[31968]_ , \new_[31969]_ , \new_[31973]_ , \new_[31974]_ ,
    \new_[31975]_ , \new_[31979]_ , \new_[31980]_ , \new_[31983]_ ,
    \new_[31986]_ , \new_[31987]_ , \new_[31988]_ , \new_[31992]_ ,
    \new_[31993]_ , \new_[31997]_ , \new_[31998]_ , \new_[31999]_ ,
    \new_[32003]_ , \new_[32004]_ , \new_[32007]_ , \new_[32010]_ ,
    \new_[32011]_ , \new_[32012]_ , \new_[32016]_ , \new_[32017]_ ,
    \new_[32021]_ , \new_[32022]_ , \new_[32023]_ , \new_[32027]_ ,
    \new_[32028]_ , \new_[32031]_ , \new_[32034]_ , \new_[32035]_ ,
    \new_[32036]_ , \new_[32040]_ , \new_[32041]_ , \new_[32045]_ ,
    \new_[32046]_ , \new_[32047]_ , \new_[32051]_ , \new_[32052]_ ,
    \new_[32055]_ , \new_[32058]_ , \new_[32059]_ , \new_[32060]_ ,
    \new_[32064]_ , \new_[32065]_ , \new_[32069]_ , \new_[32070]_ ,
    \new_[32071]_ , \new_[32075]_ , \new_[32076]_ , \new_[32079]_ ,
    \new_[32082]_ , \new_[32083]_ , \new_[32084]_ , \new_[32088]_ ,
    \new_[32089]_ , \new_[32093]_ , \new_[32094]_ , \new_[32095]_ ,
    \new_[32099]_ , \new_[32100]_ , \new_[32103]_ , \new_[32106]_ ,
    \new_[32107]_ , \new_[32108]_ , \new_[32112]_ , \new_[32113]_ ,
    \new_[32117]_ , \new_[32118]_ , \new_[32119]_ , \new_[32123]_ ,
    \new_[32124]_ , \new_[32127]_ , \new_[32130]_ , \new_[32131]_ ,
    \new_[32132]_ , \new_[32136]_ , \new_[32137]_ , \new_[32141]_ ,
    \new_[32142]_ , \new_[32143]_ , \new_[32147]_ , \new_[32148]_ ,
    \new_[32151]_ , \new_[32154]_ , \new_[32155]_ , \new_[32156]_ ,
    \new_[32160]_ , \new_[32161]_ , \new_[32165]_ , \new_[32166]_ ,
    \new_[32167]_ , \new_[32171]_ , \new_[32172]_ , \new_[32175]_ ,
    \new_[32178]_ , \new_[32179]_ , \new_[32180]_ , \new_[32184]_ ,
    \new_[32185]_ , \new_[32189]_ , \new_[32190]_ , \new_[32191]_ ,
    \new_[32195]_ , \new_[32196]_ , \new_[32199]_ , \new_[32202]_ ,
    \new_[32203]_ , \new_[32204]_ , \new_[32208]_ , \new_[32209]_ ,
    \new_[32213]_ , \new_[32214]_ , \new_[32215]_ , \new_[32219]_ ,
    \new_[32220]_ , \new_[32223]_ , \new_[32226]_ , \new_[32227]_ ,
    \new_[32228]_ , \new_[32232]_ , \new_[32233]_ , \new_[32237]_ ,
    \new_[32238]_ , \new_[32239]_ , \new_[32243]_ , \new_[32244]_ ,
    \new_[32247]_ , \new_[32250]_ , \new_[32251]_ , \new_[32252]_ ,
    \new_[32256]_ , \new_[32257]_ , \new_[32261]_ , \new_[32262]_ ,
    \new_[32263]_ , \new_[32267]_ , \new_[32268]_ , \new_[32271]_ ,
    \new_[32274]_ , \new_[32275]_ , \new_[32276]_ , \new_[32280]_ ,
    \new_[32281]_ , \new_[32285]_ , \new_[32286]_ , \new_[32287]_ ,
    \new_[32291]_ , \new_[32292]_ , \new_[32295]_ , \new_[32298]_ ,
    \new_[32299]_ , \new_[32300]_ , \new_[32304]_ , \new_[32305]_ ,
    \new_[32309]_ , \new_[32310]_ , \new_[32311]_ , \new_[32315]_ ,
    \new_[32316]_ , \new_[32319]_ , \new_[32322]_ , \new_[32323]_ ,
    \new_[32324]_ , \new_[32328]_ , \new_[32329]_ , \new_[32333]_ ,
    \new_[32334]_ , \new_[32335]_ , \new_[32339]_ , \new_[32340]_ ,
    \new_[32343]_ , \new_[32346]_ , \new_[32347]_ , \new_[32348]_ ,
    \new_[32352]_ , \new_[32353]_ , \new_[32357]_ , \new_[32358]_ ,
    \new_[32359]_ , \new_[32363]_ , \new_[32364]_ , \new_[32367]_ ,
    \new_[32370]_ , \new_[32371]_ , \new_[32372]_ , \new_[32376]_ ,
    \new_[32377]_ , \new_[32381]_ , \new_[32382]_ , \new_[32383]_ ,
    \new_[32387]_ , \new_[32388]_ , \new_[32391]_ , \new_[32394]_ ,
    \new_[32395]_ , \new_[32396]_ , \new_[32400]_ , \new_[32401]_ ,
    \new_[32405]_ , \new_[32406]_ , \new_[32407]_ , \new_[32411]_ ,
    \new_[32412]_ , \new_[32415]_ , \new_[32418]_ , \new_[32419]_ ,
    \new_[32420]_ , \new_[32424]_ , \new_[32425]_ , \new_[32429]_ ,
    \new_[32430]_ , \new_[32431]_ , \new_[32435]_ , \new_[32436]_ ,
    \new_[32439]_ , \new_[32442]_ , \new_[32443]_ , \new_[32444]_ ,
    \new_[32448]_ , \new_[32449]_ , \new_[32453]_ , \new_[32454]_ ,
    \new_[32455]_ , \new_[32459]_ , \new_[32460]_ , \new_[32463]_ ,
    \new_[32466]_ , \new_[32467]_ , \new_[32468]_ , \new_[32472]_ ,
    \new_[32473]_ , \new_[32477]_ , \new_[32478]_ , \new_[32479]_ ,
    \new_[32483]_ , \new_[32484]_ , \new_[32487]_ , \new_[32490]_ ,
    \new_[32491]_ , \new_[32492]_ , \new_[32496]_ , \new_[32497]_ ,
    \new_[32501]_ , \new_[32502]_ , \new_[32503]_ , \new_[32507]_ ,
    \new_[32508]_ , \new_[32511]_ , \new_[32514]_ , \new_[32515]_ ,
    \new_[32516]_ , \new_[32520]_ , \new_[32521]_ , \new_[32525]_ ,
    \new_[32526]_ , \new_[32527]_ , \new_[32531]_ , \new_[32532]_ ,
    \new_[32535]_ , \new_[32538]_ , \new_[32539]_ , \new_[32540]_ ,
    \new_[32544]_ , \new_[32545]_ , \new_[32549]_ , \new_[32550]_ ,
    \new_[32551]_ , \new_[32555]_ , \new_[32556]_ , \new_[32559]_ ,
    \new_[32562]_ , \new_[32563]_ , \new_[32564]_ , \new_[32568]_ ,
    \new_[32569]_ , \new_[32573]_ , \new_[32574]_ , \new_[32575]_ ,
    \new_[32579]_ , \new_[32580]_ , \new_[32583]_ , \new_[32586]_ ,
    \new_[32587]_ , \new_[32588]_ , \new_[32592]_ , \new_[32593]_ ,
    \new_[32597]_ , \new_[32598]_ , \new_[32599]_ , \new_[32603]_ ,
    \new_[32604]_ , \new_[32607]_ , \new_[32610]_ , \new_[32611]_ ,
    \new_[32612]_ , \new_[32616]_ , \new_[32617]_ , \new_[32621]_ ,
    \new_[32622]_ , \new_[32623]_ , \new_[32627]_ , \new_[32628]_ ,
    \new_[32631]_ , \new_[32634]_ , \new_[32635]_ , \new_[32636]_ ,
    \new_[32640]_ , \new_[32641]_ , \new_[32645]_ , \new_[32646]_ ,
    \new_[32647]_ , \new_[32651]_ , \new_[32652]_ , \new_[32655]_ ,
    \new_[32658]_ , \new_[32659]_ , \new_[32660]_ , \new_[32664]_ ,
    \new_[32665]_ , \new_[32669]_ , \new_[32670]_ , \new_[32671]_ ,
    \new_[32675]_ , \new_[32676]_ , \new_[32679]_ , \new_[32682]_ ,
    \new_[32683]_ , \new_[32684]_ , \new_[32688]_ , \new_[32689]_ ,
    \new_[32693]_ , \new_[32694]_ , \new_[32695]_ , \new_[32699]_ ,
    \new_[32700]_ , \new_[32703]_ , \new_[32706]_ , \new_[32707]_ ,
    \new_[32708]_ , \new_[32712]_ , \new_[32713]_ , \new_[32717]_ ,
    \new_[32718]_ , \new_[32719]_ , \new_[32723]_ , \new_[32724]_ ,
    \new_[32727]_ , \new_[32730]_ , \new_[32731]_ , \new_[32732]_ ,
    \new_[32736]_ , \new_[32737]_ , \new_[32741]_ , \new_[32742]_ ,
    \new_[32743]_ , \new_[32747]_ , \new_[32748]_ , \new_[32751]_ ,
    \new_[32754]_ , \new_[32755]_ , \new_[32756]_ , \new_[32760]_ ,
    \new_[32761]_ , \new_[32765]_ , \new_[32766]_ , \new_[32767]_ ,
    \new_[32771]_ , \new_[32772]_ , \new_[32775]_ , \new_[32778]_ ,
    \new_[32779]_ , \new_[32780]_ , \new_[32784]_ , \new_[32785]_ ,
    \new_[32789]_ , \new_[32790]_ , \new_[32791]_ , \new_[32795]_ ,
    \new_[32796]_ , \new_[32799]_ , \new_[32802]_ , \new_[32803]_ ,
    \new_[32804]_ , \new_[32808]_ , \new_[32809]_ , \new_[32813]_ ,
    \new_[32814]_ , \new_[32815]_ , \new_[32819]_ , \new_[32820]_ ,
    \new_[32823]_ , \new_[32826]_ , \new_[32827]_ , \new_[32828]_ ,
    \new_[32832]_ , \new_[32833]_ , \new_[32837]_ , \new_[32838]_ ,
    \new_[32839]_ , \new_[32843]_ , \new_[32844]_ , \new_[32847]_ ,
    \new_[32850]_ , \new_[32851]_ , \new_[32852]_ , \new_[32856]_ ,
    \new_[32857]_ , \new_[32861]_ , \new_[32862]_ , \new_[32863]_ ,
    \new_[32867]_ , \new_[32868]_ , \new_[32871]_ , \new_[32874]_ ,
    \new_[32875]_ , \new_[32876]_ , \new_[32880]_ , \new_[32881]_ ,
    \new_[32885]_ , \new_[32886]_ , \new_[32887]_ , \new_[32891]_ ,
    \new_[32892]_ , \new_[32895]_ , \new_[32898]_ , \new_[32899]_ ,
    \new_[32900]_ , \new_[32904]_ , \new_[32905]_ , \new_[32909]_ ,
    \new_[32910]_ , \new_[32911]_ , \new_[32915]_ , \new_[32916]_ ,
    \new_[32919]_ , \new_[32922]_ , \new_[32923]_ , \new_[32924]_ ,
    \new_[32928]_ , \new_[32929]_ , \new_[32933]_ , \new_[32934]_ ,
    \new_[32935]_ , \new_[32939]_ , \new_[32940]_ , \new_[32943]_ ,
    \new_[32946]_ , \new_[32947]_ , \new_[32948]_ , \new_[32952]_ ,
    \new_[32953]_ , \new_[32957]_ , \new_[32958]_ , \new_[32959]_ ,
    \new_[32963]_ , \new_[32964]_ , \new_[32967]_ , \new_[32970]_ ,
    \new_[32971]_ , \new_[32972]_ , \new_[32976]_ , \new_[32977]_ ,
    \new_[32981]_ , \new_[32982]_ , \new_[32983]_ , \new_[32987]_ ,
    \new_[32988]_ , \new_[32991]_ , \new_[32994]_ , \new_[32995]_ ,
    \new_[32996]_ , \new_[33000]_ , \new_[33001]_ , \new_[33005]_ ,
    \new_[33006]_ , \new_[33007]_ , \new_[33011]_ , \new_[33012]_ ,
    \new_[33015]_ , \new_[33018]_ , \new_[33019]_ , \new_[33020]_ ,
    \new_[33024]_ , \new_[33025]_ , \new_[33029]_ , \new_[33030]_ ,
    \new_[33031]_ , \new_[33035]_ , \new_[33036]_ , \new_[33039]_ ,
    \new_[33042]_ , \new_[33043]_ , \new_[33044]_ , \new_[33048]_ ,
    \new_[33049]_ , \new_[33053]_ , \new_[33054]_ , \new_[33055]_ ,
    \new_[33059]_ , \new_[33060]_ , \new_[33063]_ , \new_[33066]_ ,
    \new_[33067]_ , \new_[33068]_ , \new_[33072]_ , \new_[33073]_ ,
    \new_[33077]_ , \new_[33078]_ , \new_[33079]_ , \new_[33083]_ ,
    \new_[33084]_ , \new_[33087]_ , \new_[33090]_ , \new_[33091]_ ,
    \new_[33092]_ , \new_[33096]_ , \new_[33097]_ , \new_[33101]_ ,
    \new_[33102]_ , \new_[33103]_ , \new_[33107]_ , \new_[33108]_ ,
    \new_[33111]_ , \new_[33114]_ , \new_[33115]_ , \new_[33116]_ ,
    \new_[33120]_ , \new_[33121]_ , \new_[33125]_ , \new_[33126]_ ,
    \new_[33127]_ , \new_[33131]_ , \new_[33132]_ , \new_[33135]_ ,
    \new_[33138]_ , \new_[33139]_ , \new_[33140]_ , \new_[33144]_ ,
    \new_[33145]_ , \new_[33149]_ , \new_[33150]_ , \new_[33151]_ ,
    \new_[33155]_ , \new_[33156]_ , \new_[33159]_ , \new_[33162]_ ,
    \new_[33163]_ , \new_[33164]_ , \new_[33168]_ , \new_[33169]_ ,
    \new_[33173]_ , \new_[33174]_ , \new_[33175]_ , \new_[33179]_ ,
    \new_[33180]_ , \new_[33183]_ , \new_[33186]_ , \new_[33187]_ ,
    \new_[33188]_ , \new_[33192]_ , \new_[33193]_ , \new_[33197]_ ,
    \new_[33198]_ , \new_[33199]_ , \new_[33203]_ , \new_[33204]_ ,
    \new_[33207]_ , \new_[33210]_ , \new_[33211]_ , \new_[33212]_ ,
    \new_[33216]_ , \new_[33217]_ , \new_[33221]_ , \new_[33222]_ ,
    \new_[33223]_ , \new_[33227]_ , \new_[33228]_ , \new_[33231]_ ,
    \new_[33234]_ , \new_[33235]_ , \new_[33236]_ , \new_[33240]_ ,
    \new_[33241]_ , \new_[33245]_ , \new_[33246]_ , \new_[33247]_ ,
    \new_[33251]_ , \new_[33252]_ , \new_[33255]_ , \new_[33258]_ ,
    \new_[33259]_ , \new_[33260]_ , \new_[33264]_ , \new_[33265]_ ,
    \new_[33269]_ , \new_[33270]_ , \new_[33271]_ , \new_[33275]_ ,
    \new_[33276]_ , \new_[33279]_ , \new_[33282]_ , \new_[33283]_ ,
    \new_[33284]_ , \new_[33288]_ , \new_[33289]_ , \new_[33293]_ ,
    \new_[33294]_ , \new_[33295]_ , \new_[33299]_ , \new_[33300]_ ,
    \new_[33303]_ , \new_[33306]_ , \new_[33307]_ , \new_[33308]_ ,
    \new_[33312]_ , \new_[33313]_ , \new_[33317]_ , \new_[33318]_ ,
    \new_[33319]_ , \new_[33323]_ , \new_[33324]_ , \new_[33327]_ ,
    \new_[33330]_ , \new_[33331]_ , \new_[33332]_ , \new_[33336]_ ,
    \new_[33337]_ , \new_[33341]_ , \new_[33342]_ , \new_[33343]_ ,
    \new_[33347]_ , \new_[33348]_ , \new_[33351]_ , \new_[33354]_ ,
    \new_[33355]_ , \new_[33356]_ , \new_[33360]_ , \new_[33361]_ ,
    \new_[33365]_ , \new_[33366]_ , \new_[33367]_ , \new_[33371]_ ,
    \new_[33372]_ , \new_[33375]_ , \new_[33378]_ , \new_[33379]_ ,
    \new_[33380]_ , \new_[33384]_ , \new_[33385]_ , \new_[33389]_ ,
    \new_[33390]_ , \new_[33391]_ , \new_[33395]_ , \new_[33396]_ ,
    \new_[33399]_ , \new_[33402]_ , \new_[33403]_ , \new_[33404]_ ,
    \new_[33408]_ , \new_[33409]_ , \new_[33413]_ , \new_[33414]_ ,
    \new_[33415]_ , \new_[33419]_ , \new_[33420]_ , \new_[33423]_ ,
    \new_[33426]_ , \new_[33427]_ , \new_[33428]_ , \new_[33432]_ ,
    \new_[33433]_ , \new_[33437]_ , \new_[33438]_ , \new_[33439]_ ,
    \new_[33443]_ , \new_[33444]_ , \new_[33447]_ , \new_[33450]_ ,
    \new_[33451]_ , \new_[33452]_ , \new_[33456]_ , \new_[33457]_ ,
    \new_[33461]_ , \new_[33462]_ , \new_[33463]_ , \new_[33467]_ ,
    \new_[33468]_ , \new_[33471]_ , \new_[33474]_ , \new_[33475]_ ,
    \new_[33476]_ , \new_[33480]_ , \new_[33481]_ , \new_[33485]_ ,
    \new_[33486]_ , \new_[33487]_ , \new_[33491]_ , \new_[33492]_ ,
    \new_[33495]_ , \new_[33498]_ , \new_[33499]_ , \new_[33500]_ ,
    \new_[33504]_ , \new_[33505]_ , \new_[33509]_ , \new_[33510]_ ,
    \new_[33511]_ , \new_[33515]_ , \new_[33516]_ , \new_[33519]_ ,
    \new_[33522]_ , \new_[33523]_ , \new_[33524]_ , \new_[33528]_ ,
    \new_[33529]_ , \new_[33533]_ , \new_[33534]_ , \new_[33535]_ ,
    \new_[33539]_ , \new_[33540]_ , \new_[33543]_ , \new_[33546]_ ,
    \new_[33547]_ , \new_[33548]_ , \new_[33552]_ , \new_[33553]_ ,
    \new_[33557]_ , \new_[33558]_ , \new_[33559]_ , \new_[33563]_ ,
    \new_[33564]_ , \new_[33567]_ , \new_[33570]_ , \new_[33571]_ ,
    \new_[33572]_ , \new_[33576]_ , \new_[33577]_ , \new_[33581]_ ,
    \new_[33582]_ , \new_[33583]_ , \new_[33587]_ , \new_[33588]_ ,
    \new_[33591]_ , \new_[33594]_ , \new_[33595]_ , \new_[33596]_ ,
    \new_[33600]_ , \new_[33601]_ , \new_[33605]_ , \new_[33606]_ ,
    \new_[33607]_ , \new_[33611]_ , \new_[33612]_ , \new_[33615]_ ,
    \new_[33618]_ , \new_[33619]_ , \new_[33620]_ , \new_[33624]_ ,
    \new_[33625]_ , \new_[33629]_ , \new_[33630]_ , \new_[33631]_ ,
    \new_[33635]_ , \new_[33636]_ , \new_[33639]_ , \new_[33642]_ ,
    \new_[33643]_ , \new_[33644]_ , \new_[33648]_ , \new_[33649]_ ,
    \new_[33653]_ , \new_[33654]_ , \new_[33655]_ , \new_[33659]_ ,
    \new_[33660]_ , \new_[33663]_ , \new_[33666]_ , \new_[33667]_ ,
    \new_[33668]_ , \new_[33672]_ , \new_[33673]_ , \new_[33677]_ ,
    \new_[33678]_ , \new_[33679]_ , \new_[33683]_ , \new_[33684]_ ,
    \new_[33687]_ , \new_[33690]_ , \new_[33691]_ , \new_[33692]_ ,
    \new_[33696]_ , \new_[33697]_ , \new_[33701]_ , \new_[33702]_ ,
    \new_[33703]_ , \new_[33707]_ , \new_[33708]_ , \new_[33711]_ ,
    \new_[33714]_ , \new_[33715]_ , \new_[33716]_ , \new_[33720]_ ,
    \new_[33721]_ , \new_[33725]_ , \new_[33726]_ , \new_[33727]_ ,
    \new_[33731]_ , \new_[33732]_ , \new_[33735]_ , \new_[33738]_ ,
    \new_[33739]_ , \new_[33740]_ , \new_[33744]_ , \new_[33745]_ ,
    \new_[33749]_ , \new_[33750]_ , \new_[33751]_ , \new_[33755]_ ,
    \new_[33756]_ , \new_[33759]_ , \new_[33762]_ , \new_[33763]_ ,
    \new_[33764]_ , \new_[33768]_ , \new_[33769]_ , \new_[33773]_ ,
    \new_[33774]_ , \new_[33775]_ , \new_[33779]_ , \new_[33780]_ ,
    \new_[33783]_ , \new_[33786]_ , \new_[33787]_ , \new_[33788]_ ,
    \new_[33792]_ , \new_[33793]_ , \new_[33797]_ , \new_[33798]_ ,
    \new_[33799]_ , \new_[33803]_ , \new_[33804]_ , \new_[33807]_ ,
    \new_[33810]_ , \new_[33811]_ , \new_[33812]_ , \new_[33816]_ ,
    \new_[33817]_ , \new_[33821]_ , \new_[33822]_ , \new_[33823]_ ,
    \new_[33827]_ , \new_[33828]_ , \new_[33831]_ , \new_[33834]_ ,
    \new_[33835]_ , \new_[33836]_ , \new_[33840]_ , \new_[33841]_ ,
    \new_[33845]_ , \new_[33846]_ , \new_[33847]_ , \new_[33851]_ ,
    \new_[33852]_ , \new_[33855]_ , \new_[33858]_ , \new_[33859]_ ,
    \new_[33860]_ , \new_[33864]_ , \new_[33865]_ , \new_[33869]_ ,
    \new_[33870]_ , \new_[33871]_ , \new_[33875]_ , \new_[33876]_ ,
    \new_[33879]_ , \new_[33882]_ , \new_[33883]_ , \new_[33884]_ ,
    \new_[33888]_ , \new_[33889]_ , \new_[33893]_ , \new_[33894]_ ,
    \new_[33895]_ , \new_[33899]_ , \new_[33900]_ , \new_[33903]_ ,
    \new_[33906]_ , \new_[33907]_ , \new_[33908]_ , \new_[33912]_ ,
    \new_[33913]_ , \new_[33917]_ , \new_[33918]_ , \new_[33919]_ ,
    \new_[33923]_ , \new_[33924]_ , \new_[33927]_ , \new_[33930]_ ,
    \new_[33931]_ , \new_[33932]_ , \new_[33936]_ , \new_[33937]_ ,
    \new_[33941]_ , \new_[33942]_ , \new_[33943]_ , \new_[33947]_ ,
    \new_[33948]_ , \new_[33951]_ , \new_[33954]_ , \new_[33955]_ ,
    \new_[33956]_ , \new_[33960]_ , \new_[33961]_ , \new_[33965]_ ,
    \new_[33966]_ , \new_[33967]_ , \new_[33971]_ , \new_[33972]_ ,
    \new_[33975]_ , \new_[33978]_ , \new_[33979]_ , \new_[33980]_ ,
    \new_[33984]_ , \new_[33985]_ , \new_[33989]_ , \new_[33990]_ ,
    \new_[33991]_ , \new_[33995]_ , \new_[33996]_ , \new_[33999]_ ,
    \new_[34002]_ , \new_[34003]_ , \new_[34004]_ , \new_[34008]_ ,
    \new_[34009]_ , \new_[34013]_ , \new_[34014]_ , \new_[34015]_ ,
    \new_[34019]_ , \new_[34020]_ , \new_[34023]_ , \new_[34026]_ ,
    \new_[34027]_ , \new_[34028]_ , \new_[34032]_ , \new_[34033]_ ,
    \new_[34037]_ , \new_[34038]_ , \new_[34039]_ , \new_[34043]_ ,
    \new_[34044]_ , \new_[34047]_ , \new_[34050]_ , \new_[34051]_ ,
    \new_[34052]_ , \new_[34056]_ , \new_[34057]_ , \new_[34061]_ ,
    \new_[34062]_ , \new_[34063]_ , \new_[34067]_ , \new_[34068]_ ,
    \new_[34071]_ , \new_[34074]_ , \new_[34075]_ , \new_[34076]_ ,
    \new_[34080]_ , \new_[34081]_ , \new_[34085]_ , \new_[34086]_ ,
    \new_[34087]_ , \new_[34091]_ , \new_[34092]_ , \new_[34095]_ ,
    \new_[34098]_ , \new_[34099]_ , \new_[34100]_ , \new_[34104]_ ,
    \new_[34105]_ , \new_[34109]_ , \new_[34110]_ , \new_[34111]_ ,
    \new_[34115]_ , \new_[34116]_ , \new_[34119]_ , \new_[34122]_ ,
    \new_[34123]_ , \new_[34124]_ , \new_[34128]_ , \new_[34129]_ ,
    \new_[34133]_ , \new_[34134]_ , \new_[34135]_ , \new_[34139]_ ,
    \new_[34140]_ , \new_[34143]_ , \new_[34146]_ , \new_[34147]_ ,
    \new_[34148]_ , \new_[34152]_ , \new_[34153]_ , \new_[34157]_ ,
    \new_[34158]_ , \new_[34159]_ , \new_[34163]_ , \new_[34164]_ ,
    \new_[34167]_ , \new_[34170]_ , \new_[34171]_ , \new_[34172]_ ,
    \new_[34176]_ , \new_[34177]_ , \new_[34181]_ , \new_[34182]_ ,
    \new_[34183]_ , \new_[34187]_ , \new_[34188]_ , \new_[34191]_ ,
    \new_[34194]_ , \new_[34195]_ , \new_[34196]_ , \new_[34200]_ ,
    \new_[34201]_ , \new_[34205]_ , \new_[34206]_ , \new_[34207]_ ,
    \new_[34211]_ , \new_[34212]_ , \new_[34215]_ , \new_[34218]_ ,
    \new_[34219]_ , \new_[34220]_ , \new_[34224]_ , \new_[34225]_ ,
    \new_[34229]_ , \new_[34230]_ , \new_[34231]_ , \new_[34235]_ ,
    \new_[34236]_ , \new_[34239]_ , \new_[34242]_ , \new_[34243]_ ,
    \new_[34244]_ , \new_[34248]_ , \new_[34249]_ , \new_[34253]_ ,
    \new_[34254]_ , \new_[34255]_ , \new_[34259]_ , \new_[34260]_ ,
    \new_[34263]_ , \new_[34266]_ , \new_[34267]_ , \new_[34268]_ ,
    \new_[34272]_ , \new_[34273]_ , \new_[34277]_ , \new_[34278]_ ,
    \new_[34279]_ , \new_[34283]_ , \new_[34284]_ , \new_[34287]_ ,
    \new_[34290]_ , \new_[34291]_ , \new_[34292]_ , \new_[34296]_ ,
    \new_[34297]_ , \new_[34301]_ , \new_[34302]_ , \new_[34303]_ ,
    \new_[34307]_ , \new_[34308]_ , \new_[34311]_ , \new_[34314]_ ,
    \new_[34315]_ , \new_[34316]_ , \new_[34320]_ , \new_[34321]_ ,
    \new_[34325]_ , \new_[34326]_ , \new_[34327]_ , \new_[34331]_ ,
    \new_[34332]_ , \new_[34335]_ , \new_[34338]_ , \new_[34339]_ ,
    \new_[34340]_ , \new_[34344]_ , \new_[34345]_ , \new_[34349]_ ,
    \new_[34350]_ , \new_[34351]_ , \new_[34355]_ , \new_[34356]_ ,
    \new_[34359]_ , \new_[34362]_ , \new_[34363]_ , \new_[34364]_ ,
    \new_[34368]_ , \new_[34369]_ , \new_[34373]_ , \new_[34374]_ ,
    \new_[34375]_ , \new_[34379]_ , \new_[34380]_ , \new_[34383]_ ,
    \new_[34386]_ , \new_[34387]_ , \new_[34388]_ , \new_[34392]_ ,
    \new_[34393]_ , \new_[34397]_ , \new_[34398]_ , \new_[34399]_ ,
    \new_[34403]_ , \new_[34404]_ , \new_[34407]_ , \new_[34410]_ ,
    \new_[34411]_ , \new_[34412]_ , \new_[34416]_ , \new_[34417]_ ,
    \new_[34421]_ , \new_[34422]_ , \new_[34423]_ , \new_[34427]_ ,
    \new_[34428]_ , \new_[34431]_ , \new_[34434]_ , \new_[34435]_ ,
    \new_[34436]_ , \new_[34440]_ , \new_[34441]_ , \new_[34445]_ ,
    \new_[34446]_ , \new_[34447]_ , \new_[34451]_ , \new_[34452]_ ,
    \new_[34455]_ , \new_[34458]_ , \new_[34459]_ , \new_[34460]_ ,
    \new_[34464]_ , \new_[34465]_ , \new_[34469]_ , \new_[34470]_ ,
    \new_[34471]_ , \new_[34475]_ , \new_[34476]_ , \new_[34479]_ ,
    \new_[34482]_ , \new_[34483]_ , \new_[34484]_ , \new_[34488]_ ,
    \new_[34489]_ , \new_[34493]_ , \new_[34494]_ , \new_[34495]_ ,
    \new_[34499]_ , \new_[34500]_ , \new_[34503]_ , \new_[34506]_ ,
    \new_[34507]_ , \new_[34508]_ , \new_[34512]_ , \new_[34513]_ ,
    \new_[34517]_ , \new_[34518]_ , \new_[34519]_ , \new_[34523]_ ,
    \new_[34524]_ , \new_[34527]_ , \new_[34530]_ , \new_[34531]_ ,
    \new_[34532]_ , \new_[34536]_ , \new_[34537]_ , \new_[34541]_ ,
    \new_[34542]_ , \new_[34543]_ , \new_[34547]_ , \new_[34548]_ ,
    \new_[34551]_ , \new_[34554]_ , \new_[34555]_ , \new_[34556]_ ,
    \new_[34560]_ , \new_[34561]_ , \new_[34565]_ , \new_[34566]_ ,
    \new_[34567]_ , \new_[34571]_ , \new_[34572]_ , \new_[34575]_ ,
    \new_[34578]_ , \new_[34579]_ , \new_[34580]_ , \new_[34584]_ ,
    \new_[34585]_ , \new_[34589]_ , \new_[34590]_ , \new_[34591]_ ,
    \new_[34595]_ , \new_[34596]_ , \new_[34599]_ , \new_[34602]_ ,
    \new_[34603]_ , \new_[34604]_ , \new_[34608]_ , \new_[34609]_ ,
    \new_[34613]_ , \new_[34614]_ , \new_[34615]_ , \new_[34619]_ ,
    \new_[34620]_ , \new_[34623]_ , \new_[34626]_ , \new_[34627]_ ,
    \new_[34628]_ , \new_[34632]_ , \new_[34633]_ , \new_[34637]_ ,
    \new_[34638]_ , \new_[34639]_ , \new_[34643]_ , \new_[34644]_ ,
    \new_[34647]_ , \new_[34650]_ , \new_[34651]_ , \new_[34652]_ ,
    \new_[34656]_ , \new_[34657]_ , \new_[34661]_ , \new_[34662]_ ,
    \new_[34663]_ , \new_[34667]_ , \new_[34668]_ , \new_[34671]_ ,
    \new_[34674]_ , \new_[34675]_ , \new_[34676]_ , \new_[34680]_ ,
    \new_[34681]_ , \new_[34685]_ , \new_[34686]_ , \new_[34687]_ ,
    \new_[34691]_ , \new_[34692]_ , \new_[34695]_ , \new_[34698]_ ,
    \new_[34699]_ , \new_[34700]_ , \new_[34704]_ , \new_[34705]_ ,
    \new_[34709]_ , \new_[34710]_ , \new_[34711]_ , \new_[34715]_ ,
    \new_[34716]_ , \new_[34719]_ , \new_[34722]_ , \new_[34723]_ ,
    \new_[34724]_ , \new_[34728]_ , \new_[34729]_ , \new_[34733]_ ,
    \new_[34734]_ , \new_[34735]_ , \new_[34739]_ , \new_[34740]_ ,
    \new_[34743]_ , \new_[34746]_ , \new_[34747]_ , \new_[34748]_ ,
    \new_[34752]_ , \new_[34753]_ , \new_[34757]_ , \new_[34758]_ ,
    \new_[34759]_ , \new_[34763]_ , \new_[34764]_ , \new_[34767]_ ,
    \new_[34770]_ , \new_[34771]_ , \new_[34772]_ , \new_[34776]_ ,
    \new_[34777]_ , \new_[34781]_ , \new_[34782]_ , \new_[34783]_ ,
    \new_[34787]_ , \new_[34788]_ , \new_[34791]_ , \new_[34794]_ ,
    \new_[34795]_ , \new_[34796]_ , \new_[34800]_ , \new_[34801]_ ,
    \new_[34805]_ , \new_[34806]_ , \new_[34807]_ , \new_[34811]_ ,
    \new_[34812]_ , \new_[34815]_ , \new_[34818]_ , \new_[34819]_ ,
    \new_[34820]_ , \new_[34824]_ , \new_[34825]_ , \new_[34829]_ ,
    \new_[34830]_ , \new_[34831]_ , \new_[34835]_ , \new_[34836]_ ,
    \new_[34839]_ , \new_[34842]_ , \new_[34843]_ , \new_[34844]_ ,
    \new_[34848]_ , \new_[34849]_ , \new_[34853]_ , \new_[34854]_ ,
    \new_[34855]_ , \new_[34859]_ , \new_[34860]_ , \new_[34863]_ ,
    \new_[34866]_ , \new_[34867]_ , \new_[34868]_ , \new_[34872]_ ,
    \new_[34873]_ , \new_[34877]_ , \new_[34878]_ , \new_[34879]_ ,
    \new_[34883]_ , \new_[34884]_ , \new_[34887]_ , \new_[34890]_ ,
    \new_[34891]_ , \new_[34892]_ , \new_[34896]_ , \new_[34897]_ ,
    \new_[34901]_ , \new_[34902]_ , \new_[34903]_ , \new_[34907]_ ,
    \new_[34908]_ , \new_[34911]_ , \new_[34914]_ , \new_[34915]_ ,
    \new_[34916]_ , \new_[34920]_ , \new_[34921]_ , \new_[34925]_ ,
    \new_[34926]_ , \new_[34927]_ , \new_[34931]_ , \new_[34932]_ ,
    \new_[34935]_ , \new_[34938]_ , \new_[34939]_ , \new_[34940]_ ,
    \new_[34944]_ , \new_[34945]_ , \new_[34949]_ , \new_[34950]_ ,
    \new_[34951]_ , \new_[34955]_ , \new_[34956]_ , \new_[34959]_ ,
    \new_[34962]_ , \new_[34963]_ , \new_[34964]_ , \new_[34968]_ ,
    \new_[34969]_ , \new_[34973]_ , \new_[34974]_ , \new_[34975]_ ,
    \new_[34979]_ , \new_[34980]_ , \new_[34983]_ , \new_[34986]_ ,
    \new_[34987]_ , \new_[34988]_ , \new_[34992]_ , \new_[34993]_ ,
    \new_[34997]_ , \new_[34998]_ , \new_[34999]_ , \new_[35003]_ ,
    \new_[35004]_ , \new_[35007]_ , \new_[35010]_ , \new_[35011]_ ,
    \new_[35012]_ , \new_[35016]_ , \new_[35017]_ , \new_[35021]_ ,
    \new_[35022]_ , \new_[35023]_ , \new_[35027]_ , \new_[35028]_ ,
    \new_[35031]_ , \new_[35034]_ , \new_[35035]_ , \new_[35036]_ ,
    \new_[35040]_ , \new_[35041]_ , \new_[35045]_ , \new_[35046]_ ,
    \new_[35047]_ , \new_[35051]_ , \new_[35052]_ , \new_[35055]_ ,
    \new_[35058]_ , \new_[35059]_ , \new_[35060]_ , \new_[35064]_ ,
    \new_[35065]_ , \new_[35069]_ , \new_[35070]_ , \new_[35071]_ ,
    \new_[35075]_ , \new_[35076]_ , \new_[35079]_ , \new_[35082]_ ,
    \new_[35083]_ , \new_[35084]_ , \new_[35088]_ , \new_[35089]_ ,
    \new_[35093]_ , \new_[35094]_ , \new_[35095]_ , \new_[35099]_ ,
    \new_[35100]_ , \new_[35103]_ , \new_[35106]_ , \new_[35107]_ ,
    \new_[35108]_ , \new_[35112]_ , \new_[35113]_ , \new_[35117]_ ,
    \new_[35118]_ , \new_[35119]_ , \new_[35123]_ , \new_[35124]_ ,
    \new_[35127]_ , \new_[35130]_ , \new_[35131]_ , \new_[35132]_ ,
    \new_[35136]_ , \new_[35137]_ , \new_[35141]_ , \new_[35142]_ ,
    \new_[35143]_ , \new_[35147]_ , \new_[35148]_ , \new_[35151]_ ,
    \new_[35154]_ , \new_[35155]_ , \new_[35156]_ , \new_[35160]_ ,
    \new_[35161]_ , \new_[35165]_ , \new_[35166]_ , \new_[35167]_ ,
    \new_[35171]_ , \new_[35172]_ , \new_[35175]_ , \new_[35178]_ ,
    \new_[35179]_ , \new_[35180]_ , \new_[35184]_ , \new_[35185]_ ,
    \new_[35189]_ , \new_[35190]_ , \new_[35191]_ , \new_[35195]_ ,
    \new_[35196]_ , \new_[35199]_ , \new_[35202]_ , \new_[35203]_ ,
    \new_[35204]_ , \new_[35208]_ , \new_[35209]_ , \new_[35213]_ ,
    \new_[35214]_ , \new_[35215]_ , \new_[35219]_ , \new_[35220]_ ,
    \new_[35223]_ , \new_[35226]_ , \new_[35227]_ , \new_[35228]_ ,
    \new_[35232]_ , \new_[35233]_ , \new_[35237]_ , \new_[35238]_ ,
    \new_[35239]_ , \new_[35243]_ , \new_[35244]_ , \new_[35247]_ ,
    \new_[35250]_ , \new_[35251]_ , \new_[35252]_ , \new_[35256]_ ,
    \new_[35257]_ , \new_[35261]_ , \new_[35262]_ , \new_[35263]_ ,
    \new_[35267]_ , \new_[35268]_ , \new_[35271]_ , \new_[35274]_ ,
    \new_[35275]_ , \new_[35276]_ , \new_[35280]_ , \new_[35281]_ ,
    \new_[35285]_ , \new_[35286]_ , \new_[35287]_ , \new_[35291]_ ,
    \new_[35292]_ , \new_[35295]_ , \new_[35298]_ , \new_[35299]_ ,
    \new_[35300]_ , \new_[35304]_ , \new_[35305]_ , \new_[35309]_ ,
    \new_[35310]_ , \new_[35311]_ , \new_[35315]_ , \new_[35316]_ ,
    \new_[35319]_ , \new_[35322]_ , \new_[35323]_ , \new_[35324]_ ,
    \new_[35328]_ , \new_[35329]_ , \new_[35333]_ , \new_[35334]_ ,
    \new_[35335]_ , \new_[35339]_ , \new_[35340]_ , \new_[35343]_ ,
    \new_[35346]_ , \new_[35347]_ , \new_[35348]_ , \new_[35352]_ ,
    \new_[35353]_ , \new_[35357]_ , \new_[35358]_ , \new_[35359]_ ,
    \new_[35363]_ , \new_[35364]_ , \new_[35367]_ , \new_[35370]_ ,
    \new_[35371]_ , \new_[35372]_ , \new_[35376]_ , \new_[35377]_ ,
    \new_[35381]_ , \new_[35382]_ , \new_[35383]_ , \new_[35387]_ ,
    \new_[35388]_ , \new_[35391]_ , \new_[35394]_ , \new_[35395]_ ,
    \new_[35396]_ , \new_[35400]_ , \new_[35401]_ , \new_[35405]_ ,
    \new_[35406]_ , \new_[35407]_ , \new_[35411]_ , \new_[35412]_ ,
    \new_[35415]_ , \new_[35418]_ , \new_[35419]_ , \new_[35420]_ ,
    \new_[35424]_ , \new_[35425]_ , \new_[35429]_ , \new_[35430]_ ,
    \new_[35431]_ , \new_[35435]_ , \new_[35436]_ , \new_[35439]_ ,
    \new_[35442]_ , \new_[35443]_ , \new_[35444]_ , \new_[35448]_ ,
    \new_[35449]_ , \new_[35453]_ , \new_[35454]_ , \new_[35455]_ ,
    \new_[35459]_ , \new_[35460]_ , \new_[35463]_ , \new_[35466]_ ,
    \new_[35467]_ , \new_[35468]_ , \new_[35472]_ , \new_[35473]_ ,
    \new_[35477]_ , \new_[35478]_ , \new_[35479]_ , \new_[35483]_ ,
    \new_[35484]_ , \new_[35487]_ , \new_[35490]_ , \new_[35491]_ ,
    \new_[35492]_ , \new_[35496]_ , \new_[35497]_ , \new_[35501]_ ,
    \new_[35502]_ , \new_[35503]_ , \new_[35507]_ , \new_[35508]_ ,
    \new_[35511]_ , \new_[35514]_ , \new_[35515]_ , \new_[35516]_ ,
    \new_[35520]_ , \new_[35521]_ , \new_[35525]_ , \new_[35526]_ ,
    \new_[35527]_ , \new_[35531]_ , \new_[35532]_ , \new_[35535]_ ,
    \new_[35538]_ , \new_[35539]_ , \new_[35540]_ , \new_[35544]_ ,
    \new_[35545]_ , \new_[35549]_ , \new_[35550]_ , \new_[35551]_ ,
    \new_[35555]_ , \new_[35556]_ , \new_[35559]_ , \new_[35562]_ ,
    \new_[35563]_ , \new_[35564]_ , \new_[35568]_ , \new_[35569]_ ,
    \new_[35573]_ , \new_[35574]_ , \new_[35575]_ , \new_[35579]_ ,
    \new_[35580]_ , \new_[35583]_ , \new_[35586]_ , \new_[35587]_ ,
    \new_[35588]_ , \new_[35592]_ , \new_[35593]_ , \new_[35597]_ ,
    \new_[35598]_ , \new_[35599]_ , \new_[35603]_ , \new_[35604]_ ,
    \new_[35607]_ , \new_[35610]_ , \new_[35611]_ , \new_[35612]_ ,
    \new_[35616]_ , \new_[35617]_ , \new_[35621]_ , \new_[35622]_ ,
    \new_[35623]_ , \new_[35627]_ , \new_[35628]_ , \new_[35631]_ ,
    \new_[35634]_ , \new_[35635]_ , \new_[35636]_ , \new_[35640]_ ,
    \new_[35641]_ , \new_[35645]_ , \new_[35646]_ , \new_[35647]_ ,
    \new_[35651]_ , \new_[35652]_ , \new_[35655]_ , \new_[35658]_ ,
    \new_[35659]_ , \new_[35660]_ , \new_[35664]_ , \new_[35665]_ ,
    \new_[35669]_ , \new_[35670]_ , \new_[35671]_ , \new_[35675]_ ,
    \new_[35676]_ , \new_[35679]_ , \new_[35682]_ , \new_[35683]_ ,
    \new_[35684]_ , \new_[35688]_ , \new_[35689]_ , \new_[35693]_ ,
    \new_[35694]_ , \new_[35695]_ , \new_[35699]_ , \new_[35700]_ ,
    \new_[35703]_ , \new_[35706]_ , \new_[35707]_ , \new_[35708]_ ,
    \new_[35712]_ , \new_[35713]_ , \new_[35717]_ , \new_[35718]_ ,
    \new_[35719]_ , \new_[35723]_ , \new_[35724]_ , \new_[35727]_ ,
    \new_[35730]_ , \new_[35731]_ , \new_[35732]_ , \new_[35736]_ ,
    \new_[35737]_ , \new_[35741]_ , \new_[35742]_ , \new_[35743]_ ,
    \new_[35747]_ , \new_[35748]_ , \new_[35751]_ , \new_[35754]_ ,
    \new_[35755]_ , \new_[35756]_ , \new_[35760]_ , \new_[35761]_ ,
    \new_[35765]_ , \new_[35766]_ , \new_[35767]_ , \new_[35771]_ ,
    \new_[35772]_ , \new_[35775]_ , \new_[35778]_ , \new_[35779]_ ,
    \new_[35780]_ , \new_[35784]_ , \new_[35785]_ , \new_[35789]_ ,
    \new_[35790]_ , \new_[35791]_ , \new_[35795]_ , \new_[35796]_ ,
    \new_[35799]_ , \new_[35802]_ , \new_[35803]_ , \new_[35804]_ ,
    \new_[35808]_ , \new_[35809]_ , \new_[35813]_ , \new_[35814]_ ,
    \new_[35815]_ , \new_[35819]_ , \new_[35820]_ , \new_[35823]_ ,
    \new_[35826]_ , \new_[35827]_ , \new_[35828]_ , \new_[35832]_ ,
    \new_[35833]_ , \new_[35837]_ , \new_[35838]_ , \new_[35839]_ ,
    \new_[35843]_ , \new_[35844]_ , \new_[35847]_ , \new_[35850]_ ,
    \new_[35851]_ , \new_[35852]_ , \new_[35856]_ , \new_[35857]_ ,
    \new_[35861]_ , \new_[35862]_ , \new_[35863]_ , \new_[35867]_ ,
    \new_[35868]_ , \new_[35871]_ , \new_[35874]_ , \new_[35875]_ ,
    \new_[35876]_ , \new_[35880]_ , \new_[35881]_ , \new_[35885]_ ,
    \new_[35886]_ , \new_[35887]_ , \new_[35891]_ , \new_[35892]_ ,
    \new_[35895]_ , \new_[35898]_ , \new_[35899]_ , \new_[35900]_ ,
    \new_[35904]_ , \new_[35905]_ , \new_[35909]_ , \new_[35910]_ ,
    \new_[35911]_ , \new_[35915]_ , \new_[35916]_ , \new_[35919]_ ,
    \new_[35922]_ , \new_[35923]_ , \new_[35924]_ , \new_[35928]_ ,
    \new_[35929]_ , \new_[35933]_ , \new_[35934]_ , \new_[35935]_ ,
    \new_[35939]_ , \new_[35940]_ , \new_[35943]_ , \new_[35946]_ ,
    \new_[35947]_ , \new_[35948]_ , \new_[35952]_ , \new_[35953]_ ,
    \new_[35957]_ , \new_[35958]_ , \new_[35959]_ , \new_[35963]_ ,
    \new_[35964]_ , \new_[35967]_ , \new_[35970]_ , \new_[35971]_ ,
    \new_[35972]_ , \new_[35976]_ , \new_[35977]_ , \new_[35981]_ ,
    \new_[35982]_ , \new_[35983]_ , \new_[35987]_ , \new_[35988]_ ,
    \new_[35991]_ , \new_[35994]_ , \new_[35995]_ , \new_[35996]_ ,
    \new_[36000]_ , \new_[36001]_ , \new_[36005]_ , \new_[36006]_ ,
    \new_[36007]_ , \new_[36011]_ , \new_[36012]_ , \new_[36015]_ ,
    \new_[36018]_ , \new_[36019]_ , \new_[36020]_ , \new_[36024]_ ,
    \new_[36025]_ , \new_[36029]_ , \new_[36030]_ , \new_[36031]_ ,
    \new_[36035]_ , \new_[36036]_ , \new_[36039]_ , \new_[36042]_ ,
    \new_[36043]_ , \new_[36044]_ , \new_[36048]_ , \new_[36049]_ ,
    \new_[36053]_ , \new_[36054]_ , \new_[36055]_ , \new_[36059]_ ,
    \new_[36060]_ , \new_[36063]_ , \new_[36066]_ , \new_[36067]_ ,
    \new_[36068]_ , \new_[36072]_ , \new_[36073]_ , \new_[36077]_ ,
    \new_[36078]_ , \new_[36079]_ , \new_[36083]_ , \new_[36084]_ ,
    \new_[36087]_ , \new_[36090]_ , \new_[36091]_ , \new_[36092]_ ,
    \new_[36096]_ , \new_[36097]_ , \new_[36101]_ , \new_[36102]_ ,
    \new_[36103]_ , \new_[36107]_ , \new_[36108]_ , \new_[36111]_ ,
    \new_[36114]_ , \new_[36115]_ , \new_[36116]_ , \new_[36120]_ ,
    \new_[36121]_ , \new_[36125]_ , \new_[36126]_ , \new_[36127]_ ,
    \new_[36131]_ , \new_[36132]_ , \new_[36135]_ , \new_[36138]_ ,
    \new_[36139]_ , \new_[36140]_ , \new_[36144]_ , \new_[36145]_ ,
    \new_[36149]_ , \new_[36150]_ , \new_[36151]_ , \new_[36155]_ ,
    \new_[36156]_ , \new_[36159]_ , \new_[36162]_ , \new_[36163]_ ,
    \new_[36164]_ , \new_[36168]_ , \new_[36169]_ , \new_[36173]_ ,
    \new_[36174]_ , \new_[36175]_ , \new_[36179]_ , \new_[36180]_ ,
    \new_[36183]_ , \new_[36186]_ , \new_[36187]_ , \new_[36188]_ ,
    \new_[36192]_ , \new_[36193]_ , \new_[36197]_ , \new_[36198]_ ,
    \new_[36199]_ , \new_[36203]_ , \new_[36204]_ , \new_[36207]_ ,
    \new_[36210]_ , \new_[36211]_ , \new_[36212]_ , \new_[36216]_ ,
    \new_[36217]_ , \new_[36221]_ , \new_[36222]_ , \new_[36223]_ ,
    \new_[36227]_ , \new_[36228]_ , \new_[36231]_ , \new_[36234]_ ,
    \new_[36235]_ , \new_[36236]_ , \new_[36240]_ , \new_[36241]_ ,
    \new_[36245]_ , \new_[36246]_ , \new_[36247]_ , \new_[36251]_ ,
    \new_[36252]_ , \new_[36255]_ , \new_[36258]_ , \new_[36259]_ ,
    \new_[36260]_ , \new_[36264]_ , \new_[36265]_ , \new_[36269]_ ,
    \new_[36270]_ , \new_[36271]_ , \new_[36275]_ , \new_[36276]_ ,
    \new_[36279]_ , \new_[36282]_ , \new_[36283]_ , \new_[36284]_ ,
    \new_[36288]_ , \new_[36289]_ , \new_[36293]_ , \new_[36294]_ ,
    \new_[36295]_ , \new_[36299]_ , \new_[36300]_ , \new_[36303]_ ,
    \new_[36306]_ , \new_[36307]_ , \new_[36308]_ , \new_[36312]_ ,
    \new_[36313]_ , \new_[36317]_ , \new_[36318]_ , \new_[36319]_ ,
    \new_[36323]_ , \new_[36324]_ , \new_[36327]_ , \new_[36330]_ ,
    \new_[36331]_ , \new_[36332]_ , \new_[36336]_ , \new_[36337]_ ,
    \new_[36341]_ , \new_[36342]_ , \new_[36343]_ , \new_[36347]_ ,
    \new_[36348]_ , \new_[36351]_ , \new_[36354]_ , \new_[36355]_ ,
    \new_[36356]_ , \new_[36360]_ , \new_[36361]_ , \new_[36365]_ ,
    \new_[36366]_ , \new_[36367]_ , \new_[36371]_ , \new_[36372]_ ,
    \new_[36375]_ , \new_[36378]_ , \new_[36379]_ , \new_[36380]_ ,
    \new_[36384]_ , \new_[36385]_ , \new_[36389]_ , \new_[36390]_ ,
    \new_[36391]_ , \new_[36395]_ , \new_[36396]_ , \new_[36399]_ ,
    \new_[36402]_ , \new_[36403]_ , \new_[36404]_ , \new_[36408]_ ,
    \new_[36409]_ , \new_[36413]_ , \new_[36414]_ , \new_[36415]_ ,
    \new_[36419]_ , \new_[36420]_ , \new_[36423]_ , \new_[36426]_ ,
    \new_[36427]_ , \new_[36428]_ , \new_[36432]_ , \new_[36433]_ ,
    \new_[36437]_ , \new_[36438]_ , \new_[36439]_ , \new_[36443]_ ,
    \new_[36444]_ , \new_[36447]_ , \new_[36450]_ , \new_[36451]_ ,
    \new_[36452]_ , \new_[36456]_ , \new_[36457]_ , \new_[36461]_ ,
    \new_[36462]_ , \new_[36463]_ , \new_[36467]_ , \new_[36468]_ ,
    \new_[36471]_ , \new_[36474]_ , \new_[36475]_ , \new_[36476]_ ,
    \new_[36480]_ , \new_[36481]_ , \new_[36485]_ , \new_[36486]_ ,
    \new_[36487]_ , \new_[36491]_ , \new_[36492]_ , \new_[36495]_ ,
    \new_[36498]_ , \new_[36499]_ , \new_[36500]_ , \new_[36504]_ ,
    \new_[36505]_ , \new_[36509]_ , \new_[36510]_ , \new_[36511]_ ,
    \new_[36515]_ , \new_[36516]_ , \new_[36519]_ , \new_[36522]_ ,
    \new_[36523]_ , \new_[36524]_ , \new_[36528]_ , \new_[36529]_ ,
    \new_[36533]_ , \new_[36534]_ , \new_[36535]_ , \new_[36539]_ ,
    \new_[36540]_ , \new_[36543]_ , \new_[36546]_ , \new_[36547]_ ,
    \new_[36548]_ , \new_[36552]_ , \new_[36553]_ , \new_[36557]_ ,
    \new_[36558]_ , \new_[36559]_ , \new_[36563]_ , \new_[36564]_ ,
    \new_[36567]_ , \new_[36570]_ , \new_[36571]_ , \new_[36572]_ ,
    \new_[36576]_ , \new_[36577]_ , \new_[36581]_ , \new_[36582]_ ,
    \new_[36583]_ , \new_[36587]_ , \new_[36588]_ , \new_[36591]_ ,
    \new_[36594]_ , \new_[36595]_ , \new_[36596]_ , \new_[36600]_ ,
    \new_[36601]_ , \new_[36605]_ , \new_[36606]_ , \new_[36607]_ ,
    \new_[36611]_ , \new_[36612]_ , \new_[36615]_ , \new_[36618]_ ,
    \new_[36619]_ , \new_[36620]_ , \new_[36624]_ , \new_[36625]_ ,
    \new_[36629]_ , \new_[36630]_ , \new_[36631]_ , \new_[36635]_ ,
    \new_[36636]_ , \new_[36639]_ , \new_[36642]_ , \new_[36643]_ ,
    \new_[36644]_ , \new_[36648]_ , \new_[36649]_ , \new_[36653]_ ,
    \new_[36654]_ , \new_[36655]_ , \new_[36659]_ , \new_[36660]_ ,
    \new_[36663]_ , \new_[36666]_ , \new_[36667]_ , \new_[36668]_ ,
    \new_[36672]_ , \new_[36673]_ , \new_[36677]_ , \new_[36678]_ ,
    \new_[36679]_ , \new_[36683]_ , \new_[36684]_ , \new_[36687]_ ,
    \new_[36690]_ , \new_[36691]_ , \new_[36692]_ , \new_[36696]_ ,
    \new_[36697]_ , \new_[36701]_ , \new_[36702]_ , \new_[36703]_ ,
    \new_[36707]_ , \new_[36708]_ , \new_[36711]_ , \new_[36714]_ ,
    \new_[36715]_ , \new_[36716]_ , \new_[36720]_ , \new_[36721]_ ,
    \new_[36725]_ , \new_[36726]_ , \new_[36727]_ , \new_[36731]_ ,
    \new_[36732]_ , \new_[36735]_ , \new_[36738]_ , \new_[36739]_ ,
    \new_[36740]_ , \new_[36744]_ , \new_[36745]_ , \new_[36749]_ ,
    \new_[36750]_ , \new_[36751]_ , \new_[36755]_ , \new_[36756]_ ,
    \new_[36759]_ , \new_[36762]_ , \new_[36763]_ , \new_[36764]_ ,
    \new_[36768]_ , \new_[36769]_ , \new_[36773]_ , \new_[36774]_ ,
    \new_[36775]_ , \new_[36779]_ , \new_[36780]_ , \new_[36783]_ ,
    \new_[36786]_ , \new_[36787]_ , \new_[36788]_ , \new_[36792]_ ,
    \new_[36793]_ , \new_[36797]_ , \new_[36798]_ , \new_[36799]_ ,
    \new_[36803]_ , \new_[36804]_ , \new_[36807]_ , \new_[36810]_ ,
    \new_[36811]_ , \new_[36812]_ , \new_[36816]_ , \new_[36817]_ ,
    \new_[36821]_ , \new_[36822]_ , \new_[36823]_ , \new_[36827]_ ,
    \new_[36828]_ , \new_[36831]_ , \new_[36834]_ , \new_[36835]_ ,
    \new_[36836]_ , \new_[36840]_ , \new_[36841]_ , \new_[36845]_ ,
    \new_[36846]_ , \new_[36847]_ , \new_[36851]_ , \new_[36852]_ ,
    \new_[36855]_ , \new_[36858]_ , \new_[36859]_ , \new_[36860]_ ,
    \new_[36864]_ , \new_[36865]_ , \new_[36869]_ , \new_[36870]_ ,
    \new_[36871]_ , \new_[36875]_ , \new_[36876]_ , \new_[36879]_ ,
    \new_[36882]_ , \new_[36883]_ , \new_[36884]_ , \new_[36888]_ ,
    \new_[36889]_ , \new_[36893]_ , \new_[36894]_ , \new_[36895]_ ,
    \new_[36899]_ , \new_[36900]_ , \new_[36903]_ , \new_[36906]_ ,
    \new_[36907]_ , \new_[36908]_ , \new_[36912]_ , \new_[36913]_ ,
    \new_[36917]_ , \new_[36918]_ , \new_[36919]_ , \new_[36923]_ ,
    \new_[36924]_ , \new_[36927]_ , \new_[36930]_ , \new_[36931]_ ,
    \new_[36932]_ , \new_[36936]_ , \new_[36937]_ , \new_[36941]_ ,
    \new_[36942]_ , \new_[36943]_ , \new_[36947]_ , \new_[36948]_ ,
    \new_[36951]_ , \new_[36954]_ , \new_[36955]_ , \new_[36956]_ ,
    \new_[36960]_ , \new_[36961]_ , \new_[36965]_ , \new_[36966]_ ,
    \new_[36967]_ , \new_[36971]_ , \new_[36972]_ , \new_[36975]_ ,
    \new_[36978]_ , \new_[36979]_ , \new_[36980]_ , \new_[36984]_ ,
    \new_[36985]_ , \new_[36989]_ , \new_[36990]_ , \new_[36991]_ ,
    \new_[36995]_ , \new_[36996]_ , \new_[36999]_ , \new_[37002]_ ,
    \new_[37003]_ , \new_[37004]_ , \new_[37008]_ , \new_[37009]_ ,
    \new_[37013]_ , \new_[37014]_ , \new_[37015]_ , \new_[37019]_ ,
    \new_[37020]_ , \new_[37023]_ , \new_[37026]_ , \new_[37027]_ ,
    \new_[37028]_ , \new_[37032]_ , \new_[37033]_ , \new_[37037]_ ,
    \new_[37038]_ , \new_[37039]_ , \new_[37043]_ , \new_[37044]_ ,
    \new_[37047]_ , \new_[37050]_ , \new_[37051]_ , \new_[37052]_ ,
    \new_[37056]_ , \new_[37057]_ , \new_[37061]_ , \new_[37062]_ ,
    \new_[37063]_ , \new_[37067]_ , \new_[37068]_ , \new_[37071]_ ,
    \new_[37074]_ , \new_[37075]_ , \new_[37076]_ , \new_[37080]_ ,
    \new_[37081]_ , \new_[37085]_ , \new_[37086]_ , \new_[37087]_ ,
    \new_[37091]_ , \new_[37092]_ , \new_[37095]_ , \new_[37098]_ ,
    \new_[37099]_ , \new_[37100]_ , \new_[37104]_ , \new_[37105]_ ,
    \new_[37109]_ , \new_[37110]_ , \new_[37111]_ , \new_[37115]_ ,
    \new_[37116]_ , \new_[37119]_ , \new_[37122]_ , \new_[37123]_ ,
    \new_[37124]_ , \new_[37128]_ , \new_[37129]_ , \new_[37133]_ ,
    \new_[37134]_ , \new_[37135]_ , \new_[37139]_ , \new_[37140]_ ,
    \new_[37143]_ , \new_[37146]_ , \new_[37147]_ , \new_[37148]_ ,
    \new_[37152]_ , \new_[37153]_ , \new_[37157]_ , \new_[37158]_ ,
    \new_[37159]_ , \new_[37163]_ , \new_[37164]_ , \new_[37167]_ ,
    \new_[37170]_ , \new_[37171]_ , \new_[37172]_ , \new_[37176]_ ,
    \new_[37177]_ , \new_[37181]_ , \new_[37182]_ , \new_[37183]_ ,
    \new_[37187]_ , \new_[37188]_ , \new_[37191]_ , \new_[37194]_ ,
    \new_[37195]_ , \new_[37196]_ , \new_[37200]_ , \new_[37201]_ ,
    \new_[37205]_ , \new_[37206]_ , \new_[37207]_ , \new_[37211]_ ,
    \new_[37212]_ , \new_[37215]_ , \new_[37218]_ , \new_[37219]_ ,
    \new_[37220]_ , \new_[37224]_ , \new_[37225]_ , \new_[37229]_ ,
    \new_[37230]_ , \new_[37231]_ , \new_[37235]_ , \new_[37236]_ ,
    \new_[37239]_ , \new_[37242]_ , \new_[37243]_ , \new_[37244]_ ,
    \new_[37248]_ , \new_[37249]_ , \new_[37253]_ , \new_[37254]_ ,
    \new_[37255]_ , \new_[37259]_ , \new_[37260]_ , \new_[37263]_ ,
    \new_[37266]_ , \new_[37267]_ , \new_[37268]_ , \new_[37272]_ ,
    \new_[37273]_ , \new_[37277]_ , \new_[37278]_ , \new_[37279]_ ,
    \new_[37283]_ , \new_[37284]_ , \new_[37287]_ , \new_[37290]_ ,
    \new_[37291]_ , \new_[37292]_ , \new_[37296]_ , \new_[37297]_ ,
    \new_[37301]_ , \new_[37302]_ , \new_[37303]_ , \new_[37307]_ ,
    \new_[37308]_ , \new_[37311]_ , \new_[37314]_ , \new_[37315]_ ,
    \new_[37316]_ , \new_[37320]_ , \new_[37321]_ , \new_[37325]_ ,
    \new_[37326]_ , \new_[37327]_ , \new_[37331]_ , \new_[37332]_ ,
    \new_[37335]_ , \new_[37338]_ , \new_[37339]_ , \new_[37340]_ ,
    \new_[37344]_ , \new_[37345]_ , \new_[37349]_ , \new_[37350]_ ,
    \new_[37351]_ , \new_[37355]_ , \new_[37356]_ , \new_[37359]_ ,
    \new_[37362]_ , \new_[37363]_ , \new_[37364]_ , \new_[37368]_ ,
    \new_[37369]_ , \new_[37373]_ , \new_[37374]_ , \new_[37375]_ ,
    \new_[37379]_ , \new_[37380]_ , \new_[37383]_ , \new_[37386]_ ,
    \new_[37387]_ , \new_[37388]_ , \new_[37392]_ , \new_[37393]_ ,
    \new_[37397]_ , \new_[37398]_ , \new_[37399]_ , \new_[37403]_ ,
    \new_[37404]_ , \new_[37407]_ , \new_[37410]_ , \new_[37411]_ ,
    \new_[37412]_ , \new_[37416]_ , \new_[37417]_ , \new_[37421]_ ,
    \new_[37422]_ , \new_[37423]_ , \new_[37427]_ , \new_[37428]_ ,
    \new_[37431]_ , \new_[37434]_ , \new_[37435]_ , \new_[37436]_ ,
    \new_[37440]_ , \new_[37441]_ , \new_[37445]_ , \new_[37446]_ ,
    \new_[37447]_ , \new_[37451]_ , \new_[37452]_ , \new_[37455]_ ,
    \new_[37458]_ , \new_[37459]_ , \new_[37460]_ , \new_[37464]_ ,
    \new_[37465]_ , \new_[37469]_ , \new_[37470]_ , \new_[37471]_ ,
    \new_[37475]_ , \new_[37476]_ , \new_[37479]_ , \new_[37482]_ ,
    \new_[37483]_ , \new_[37484]_ , \new_[37488]_ , \new_[37489]_ ,
    \new_[37493]_ , \new_[37494]_ , \new_[37495]_ , \new_[37499]_ ,
    \new_[37500]_ , \new_[37503]_ , \new_[37506]_ , \new_[37507]_ ,
    \new_[37508]_ , \new_[37512]_ , \new_[37513]_ , \new_[37517]_ ,
    \new_[37518]_ , \new_[37519]_ , \new_[37523]_ , \new_[37524]_ ,
    \new_[37527]_ , \new_[37530]_ , \new_[37531]_ , \new_[37532]_ ,
    \new_[37536]_ , \new_[37537]_ , \new_[37541]_ , \new_[37542]_ ,
    \new_[37543]_ , \new_[37547]_ , \new_[37548]_ , \new_[37551]_ ,
    \new_[37554]_ , \new_[37555]_ , \new_[37556]_ , \new_[37560]_ ,
    \new_[37561]_ , \new_[37565]_ , \new_[37566]_ , \new_[37567]_ ,
    \new_[37571]_ , \new_[37572]_ , \new_[37575]_ , \new_[37578]_ ,
    \new_[37579]_ , \new_[37580]_ , \new_[37584]_ , \new_[37585]_ ,
    \new_[37589]_ , \new_[37590]_ , \new_[37591]_ , \new_[37595]_ ,
    \new_[37596]_ , \new_[37599]_ , \new_[37602]_ , \new_[37603]_ ,
    \new_[37604]_ , \new_[37608]_ , \new_[37609]_ , \new_[37613]_ ,
    \new_[37614]_ , \new_[37615]_ , \new_[37619]_ , \new_[37620]_ ,
    \new_[37623]_ , \new_[37626]_ , \new_[37627]_ , \new_[37628]_ ,
    \new_[37632]_ , \new_[37633]_ , \new_[37637]_ , \new_[37638]_ ,
    \new_[37639]_ , \new_[37643]_ , \new_[37644]_ , \new_[37647]_ ,
    \new_[37650]_ , \new_[37651]_ , \new_[37652]_ , \new_[37656]_ ,
    \new_[37657]_ , \new_[37661]_ , \new_[37662]_ , \new_[37663]_ ,
    \new_[37667]_ , \new_[37668]_ , \new_[37671]_ , \new_[37674]_ ,
    \new_[37675]_ , \new_[37676]_ , \new_[37680]_ , \new_[37681]_ ,
    \new_[37685]_ , \new_[37686]_ , \new_[37687]_ , \new_[37691]_ ,
    \new_[37692]_ , \new_[37695]_ , \new_[37698]_ , \new_[37699]_ ,
    \new_[37700]_ , \new_[37704]_ , \new_[37705]_ , \new_[37709]_ ,
    \new_[37710]_ , \new_[37711]_ , \new_[37715]_ , \new_[37716]_ ,
    \new_[37719]_ , \new_[37722]_ , \new_[37723]_ , \new_[37724]_ ,
    \new_[37728]_ , \new_[37729]_ , \new_[37733]_ , \new_[37734]_ ,
    \new_[37735]_ , \new_[37739]_ , \new_[37740]_ , \new_[37743]_ ,
    \new_[37746]_ , \new_[37747]_ , \new_[37748]_ , \new_[37752]_ ,
    \new_[37753]_ , \new_[37757]_ , \new_[37758]_ , \new_[37759]_ ,
    \new_[37763]_ , \new_[37764]_ , \new_[37767]_ , \new_[37770]_ ,
    \new_[37771]_ , \new_[37772]_ , \new_[37776]_ , \new_[37777]_ ,
    \new_[37781]_ , \new_[37782]_ , \new_[37783]_ , \new_[37787]_ ,
    \new_[37788]_ , \new_[37791]_ , \new_[37794]_ , \new_[37795]_ ,
    \new_[37796]_ , \new_[37800]_ , \new_[37801]_ , \new_[37805]_ ,
    \new_[37806]_ , \new_[37807]_ , \new_[37811]_ , \new_[37812]_ ,
    \new_[37815]_ , \new_[37818]_ , \new_[37819]_ , \new_[37820]_ ,
    \new_[37824]_ , \new_[37825]_ , \new_[37828]_ , \new_[37831]_ ,
    \new_[37832]_ , \new_[37833]_ , \new_[37837]_ , \new_[37838]_ ,
    \new_[37841]_ , \new_[37844]_ , \new_[37845]_ , \new_[37846]_ ,
    \new_[37850]_ , \new_[37851]_ , \new_[37854]_ , \new_[37857]_ ,
    \new_[37858]_ , \new_[37859]_ , \new_[37863]_ , \new_[37864]_ ,
    \new_[37867]_ , \new_[37870]_ , \new_[37871]_ , \new_[37872]_ ,
    \new_[37876]_ , \new_[37877]_ , \new_[37880]_ , \new_[37883]_ ,
    \new_[37884]_ , \new_[37885]_ , \new_[37889]_ , \new_[37890]_ ,
    \new_[37893]_ , \new_[37896]_ , \new_[37897]_ , \new_[37898]_ ,
    \new_[37902]_ , \new_[37903]_ , \new_[37906]_ , \new_[37909]_ ,
    \new_[37910]_ , \new_[37911]_ , \new_[37915]_ , \new_[37916]_ ,
    \new_[37919]_ , \new_[37922]_ , \new_[37923]_ , \new_[37924]_ ,
    \new_[37928]_ , \new_[37929]_ , \new_[37932]_ , \new_[37935]_ ,
    \new_[37936]_ , \new_[37937]_ , \new_[37941]_ , \new_[37942]_ ,
    \new_[37945]_ , \new_[37948]_ , \new_[37949]_ , \new_[37950]_ ,
    \new_[37954]_ , \new_[37955]_ , \new_[37958]_ , \new_[37961]_ ,
    \new_[37962]_ , \new_[37963]_ , \new_[37967]_ , \new_[37968]_ ,
    \new_[37971]_ , \new_[37974]_ , \new_[37975]_ , \new_[37976]_ ,
    \new_[37980]_ , \new_[37981]_ , \new_[37984]_ , \new_[37987]_ ,
    \new_[37988]_ , \new_[37989]_ , \new_[37993]_ , \new_[37994]_ ,
    \new_[37997]_ , \new_[38000]_ , \new_[38001]_ , \new_[38002]_ ,
    \new_[38006]_ , \new_[38007]_ , \new_[38010]_ , \new_[38013]_ ,
    \new_[38014]_ , \new_[38015]_ , \new_[38019]_ , \new_[38020]_ ,
    \new_[38023]_ , \new_[38026]_ , \new_[38027]_ , \new_[38028]_ ,
    \new_[38032]_ , \new_[38033]_ , \new_[38036]_ , \new_[38039]_ ,
    \new_[38040]_ , \new_[38041]_ , \new_[38045]_ , \new_[38046]_ ,
    \new_[38049]_ , \new_[38052]_ , \new_[38053]_ , \new_[38054]_ ,
    \new_[38058]_ , \new_[38059]_ , \new_[38062]_ , \new_[38065]_ ,
    \new_[38066]_ , \new_[38067]_ , \new_[38071]_ , \new_[38072]_ ,
    \new_[38075]_ , \new_[38078]_ , \new_[38079]_ , \new_[38080]_ ,
    \new_[38084]_ , \new_[38085]_ , \new_[38088]_ , \new_[38091]_ ,
    \new_[38092]_ , \new_[38093]_ , \new_[38097]_ , \new_[38098]_ ,
    \new_[38101]_ , \new_[38104]_ , \new_[38105]_ , \new_[38106]_ ,
    \new_[38110]_ , \new_[38111]_ , \new_[38114]_ , \new_[38117]_ ,
    \new_[38118]_ , \new_[38119]_ , \new_[38123]_ , \new_[38124]_ ,
    \new_[38127]_ , \new_[38130]_ , \new_[38131]_ , \new_[38132]_ ,
    \new_[38136]_ , \new_[38137]_ , \new_[38140]_ , \new_[38143]_ ,
    \new_[38144]_ , \new_[38145]_ , \new_[38149]_ , \new_[38150]_ ,
    \new_[38153]_ , \new_[38156]_ , \new_[38157]_ , \new_[38158]_ ,
    \new_[38162]_ , \new_[38163]_ , \new_[38166]_ , \new_[38169]_ ,
    \new_[38170]_ , \new_[38171]_ , \new_[38175]_ , \new_[38176]_ ,
    \new_[38179]_ , \new_[38182]_ , \new_[38183]_ , \new_[38184]_ ,
    \new_[38188]_ , \new_[38189]_ , \new_[38192]_ , \new_[38195]_ ,
    \new_[38196]_ , \new_[38197]_ , \new_[38201]_ , \new_[38202]_ ,
    \new_[38205]_ , \new_[38208]_ , \new_[38209]_ , \new_[38210]_ ,
    \new_[38214]_ , \new_[38215]_ , \new_[38218]_ , \new_[38221]_ ,
    \new_[38222]_ , \new_[38223]_ , \new_[38227]_ , \new_[38228]_ ,
    \new_[38231]_ , \new_[38234]_ , \new_[38235]_ , \new_[38236]_ ,
    \new_[38240]_ , \new_[38241]_ , \new_[38244]_ , \new_[38247]_ ,
    \new_[38248]_ , \new_[38249]_ , \new_[38253]_ , \new_[38254]_ ,
    \new_[38257]_ , \new_[38260]_ , \new_[38261]_ , \new_[38262]_ ,
    \new_[38266]_ , \new_[38267]_ , \new_[38270]_ , \new_[38273]_ ,
    \new_[38274]_ , \new_[38275]_ , \new_[38279]_ , \new_[38280]_ ,
    \new_[38283]_ , \new_[38286]_ , \new_[38287]_ , \new_[38288]_ ,
    \new_[38292]_ , \new_[38293]_ , \new_[38296]_ , \new_[38299]_ ,
    \new_[38300]_ , \new_[38301]_ , \new_[38305]_ , \new_[38306]_ ,
    \new_[38309]_ , \new_[38312]_ , \new_[38313]_ , \new_[38314]_ ,
    \new_[38318]_ , \new_[38319]_ , \new_[38322]_ , \new_[38325]_ ,
    \new_[38326]_ , \new_[38327]_ , \new_[38331]_ , \new_[38332]_ ,
    \new_[38335]_ , \new_[38338]_ , \new_[38339]_ , \new_[38340]_ ,
    \new_[38344]_ , \new_[38345]_ , \new_[38348]_ , \new_[38351]_ ,
    \new_[38352]_ , \new_[38353]_ , \new_[38357]_ , \new_[38358]_ ,
    \new_[38361]_ , \new_[38364]_ , \new_[38365]_ , \new_[38366]_ ,
    \new_[38370]_ , \new_[38371]_ , \new_[38374]_ , \new_[38377]_ ,
    \new_[38378]_ , \new_[38379]_ , \new_[38383]_ , \new_[38384]_ ,
    \new_[38387]_ , \new_[38390]_ , \new_[38391]_ , \new_[38392]_ ,
    \new_[38396]_ , \new_[38397]_ , \new_[38400]_ , \new_[38403]_ ,
    \new_[38404]_ , \new_[38405]_ , \new_[38409]_ , \new_[38410]_ ,
    \new_[38413]_ , \new_[38416]_ , \new_[38417]_ , \new_[38418]_ ,
    \new_[38422]_ , \new_[38423]_ , \new_[38426]_ , \new_[38429]_ ,
    \new_[38430]_ , \new_[38431]_ , \new_[38435]_ , \new_[38436]_ ,
    \new_[38439]_ , \new_[38442]_ , \new_[38443]_ , \new_[38444]_ ,
    \new_[38448]_ , \new_[38449]_ , \new_[38452]_ , \new_[38455]_ ,
    \new_[38456]_ , \new_[38457]_ , \new_[38461]_ , \new_[38462]_ ,
    \new_[38465]_ , \new_[38468]_ , \new_[38469]_ , \new_[38470]_ ,
    \new_[38474]_ , \new_[38475]_ , \new_[38478]_ , \new_[38481]_ ,
    \new_[38482]_ , \new_[38483]_ , \new_[38487]_ , \new_[38488]_ ,
    \new_[38491]_ , \new_[38494]_ , \new_[38495]_ , \new_[38496]_ ,
    \new_[38500]_ , \new_[38501]_ , \new_[38504]_ , \new_[38507]_ ,
    \new_[38508]_ , \new_[38509]_ , \new_[38513]_ , \new_[38514]_ ,
    \new_[38517]_ , \new_[38520]_ , \new_[38521]_ , \new_[38522]_ ,
    \new_[38526]_ , \new_[38527]_ , \new_[38530]_ , \new_[38533]_ ,
    \new_[38534]_ , \new_[38535]_ , \new_[38539]_ , \new_[38540]_ ,
    \new_[38543]_ , \new_[38546]_ , \new_[38547]_ , \new_[38548]_ ,
    \new_[38552]_ , \new_[38553]_ , \new_[38556]_ , \new_[38559]_ ,
    \new_[38560]_ , \new_[38561]_ , \new_[38565]_ , \new_[38566]_ ,
    \new_[38569]_ , \new_[38572]_ , \new_[38573]_ , \new_[38574]_ ,
    \new_[38578]_ , \new_[38579]_ , \new_[38582]_ , \new_[38585]_ ,
    \new_[38586]_ , \new_[38587]_ , \new_[38591]_ , \new_[38592]_ ,
    \new_[38595]_ , \new_[38598]_ , \new_[38599]_ , \new_[38600]_ ,
    \new_[38604]_ , \new_[38605]_ , \new_[38608]_ , \new_[38611]_ ,
    \new_[38612]_ , \new_[38613]_ , \new_[38617]_ , \new_[38618]_ ,
    \new_[38621]_ , \new_[38624]_ , \new_[38625]_ , \new_[38626]_ ,
    \new_[38630]_ , \new_[38631]_ , \new_[38634]_ , \new_[38637]_ ,
    \new_[38638]_ , \new_[38639]_ , \new_[38643]_ , \new_[38644]_ ,
    \new_[38647]_ , \new_[38650]_ , \new_[38651]_ , \new_[38652]_ ,
    \new_[38656]_ , \new_[38657]_ , \new_[38660]_ , \new_[38663]_ ,
    \new_[38664]_ , \new_[38665]_ , \new_[38669]_ , \new_[38670]_ ,
    \new_[38673]_ , \new_[38676]_ , \new_[38677]_ , \new_[38678]_ ,
    \new_[38682]_ , \new_[38683]_ , \new_[38686]_ , \new_[38689]_ ,
    \new_[38690]_ , \new_[38691]_ , \new_[38695]_ , \new_[38696]_ ,
    \new_[38699]_ , \new_[38702]_ , \new_[38703]_ , \new_[38704]_ ,
    \new_[38708]_ , \new_[38709]_ , \new_[38712]_ , \new_[38715]_ ,
    \new_[38716]_ , \new_[38717]_ , \new_[38721]_ , \new_[38722]_ ,
    \new_[38725]_ , \new_[38728]_ , \new_[38729]_ , \new_[38730]_ ,
    \new_[38734]_ , \new_[38735]_ , \new_[38738]_ , \new_[38741]_ ,
    \new_[38742]_ , \new_[38743]_ , \new_[38747]_ , \new_[38748]_ ,
    \new_[38751]_ , \new_[38754]_ , \new_[38755]_ , \new_[38756]_ ,
    \new_[38760]_ , \new_[38761]_ , \new_[38764]_ , \new_[38767]_ ,
    \new_[38768]_ , \new_[38769]_ , \new_[38773]_ , \new_[38774]_ ,
    \new_[38777]_ , \new_[38780]_ , \new_[38781]_ , \new_[38782]_ ,
    \new_[38786]_ , \new_[38787]_ , \new_[38790]_ , \new_[38793]_ ,
    \new_[38794]_ , \new_[38795]_ , \new_[38799]_ , \new_[38800]_ ,
    \new_[38803]_ , \new_[38806]_ , \new_[38807]_ , \new_[38808]_ ,
    \new_[38812]_ , \new_[38813]_ , \new_[38816]_ , \new_[38819]_ ,
    \new_[38820]_ , \new_[38821]_ , \new_[38825]_ , \new_[38826]_ ,
    \new_[38829]_ , \new_[38832]_ , \new_[38833]_ , \new_[38834]_ ,
    \new_[38838]_ , \new_[38839]_ , \new_[38842]_ , \new_[38845]_ ,
    \new_[38846]_ , \new_[38847]_ , \new_[38851]_ , \new_[38852]_ ,
    \new_[38855]_ , \new_[38858]_ , \new_[38859]_ , \new_[38860]_ ,
    \new_[38864]_ , \new_[38865]_ , \new_[38868]_ , \new_[38871]_ ,
    \new_[38872]_ , \new_[38873]_ , \new_[38877]_ , \new_[38878]_ ,
    \new_[38881]_ , \new_[38884]_ , \new_[38885]_ , \new_[38886]_ ,
    \new_[38890]_ , \new_[38891]_ , \new_[38894]_ , \new_[38897]_ ,
    \new_[38898]_ , \new_[38899]_ , \new_[38903]_ , \new_[38904]_ ,
    \new_[38907]_ , \new_[38910]_ , \new_[38911]_ , \new_[38912]_ ,
    \new_[38916]_ , \new_[38917]_ , \new_[38920]_ , \new_[38923]_ ,
    \new_[38924]_ , \new_[38925]_ , \new_[38929]_ , \new_[38930]_ ,
    \new_[38933]_ , \new_[38936]_ , \new_[38937]_ , \new_[38938]_ ,
    \new_[38942]_ , \new_[38943]_ , \new_[38946]_ , \new_[38949]_ ,
    \new_[38950]_ , \new_[38951]_ , \new_[38955]_ , \new_[38956]_ ,
    \new_[38959]_ , \new_[38962]_ , \new_[38963]_ , \new_[38964]_ ,
    \new_[38968]_ , \new_[38969]_ , \new_[38972]_ , \new_[38975]_ ,
    \new_[38976]_ , \new_[38977]_ , \new_[38981]_ , \new_[38982]_ ,
    \new_[38985]_ , \new_[38988]_ , \new_[38989]_ , \new_[38990]_ ,
    \new_[38994]_ , \new_[38995]_ , \new_[38998]_ , \new_[39001]_ ,
    \new_[39002]_ , \new_[39003]_ , \new_[39007]_ , \new_[39008]_ ,
    \new_[39011]_ , \new_[39014]_ , \new_[39015]_ , \new_[39016]_ ,
    \new_[39020]_ , \new_[39021]_ , \new_[39024]_ , \new_[39027]_ ,
    \new_[39028]_ , \new_[39029]_ , \new_[39033]_ , \new_[39034]_ ,
    \new_[39037]_ , \new_[39040]_ , \new_[39041]_ , \new_[39042]_ ,
    \new_[39046]_ , \new_[39047]_ , \new_[39050]_ , \new_[39053]_ ,
    \new_[39054]_ , \new_[39055]_ , \new_[39059]_ , \new_[39060]_ ,
    \new_[39063]_ , \new_[39066]_ , \new_[39067]_ , \new_[39068]_ ,
    \new_[39072]_ , \new_[39073]_ , \new_[39076]_ , \new_[39079]_ ,
    \new_[39080]_ , \new_[39081]_ , \new_[39085]_ , \new_[39086]_ ,
    \new_[39089]_ , \new_[39092]_ , \new_[39093]_ , \new_[39094]_ ,
    \new_[39098]_ , \new_[39099]_ , \new_[39102]_ , \new_[39105]_ ,
    \new_[39106]_ , \new_[39107]_ , \new_[39111]_ , \new_[39112]_ ,
    \new_[39115]_ , \new_[39118]_ , \new_[39119]_ , \new_[39120]_ ,
    \new_[39124]_ , \new_[39125]_ , \new_[39128]_ , \new_[39131]_ ,
    \new_[39132]_ , \new_[39133]_ , \new_[39137]_ , \new_[39138]_ ,
    \new_[39141]_ , \new_[39144]_ , \new_[39145]_ , \new_[39146]_ ,
    \new_[39150]_ , \new_[39151]_ , \new_[39154]_ , \new_[39157]_ ,
    \new_[39158]_ , \new_[39159]_ , \new_[39163]_ , \new_[39164]_ ,
    \new_[39167]_ , \new_[39170]_ , \new_[39171]_ , \new_[39172]_ ,
    \new_[39176]_ , \new_[39177]_ , \new_[39180]_ , \new_[39183]_ ,
    \new_[39184]_ , \new_[39185]_ , \new_[39189]_ , \new_[39190]_ ,
    \new_[39193]_ , \new_[39196]_ , \new_[39197]_ , \new_[39198]_ ,
    \new_[39202]_ , \new_[39203]_ , \new_[39206]_ , \new_[39209]_ ,
    \new_[39210]_ , \new_[39211]_ , \new_[39215]_ , \new_[39216]_ ,
    \new_[39219]_ , \new_[39222]_ , \new_[39223]_ , \new_[39224]_ ,
    \new_[39228]_ , \new_[39229]_ , \new_[39232]_ , \new_[39235]_ ,
    \new_[39236]_ , \new_[39237]_ , \new_[39241]_ , \new_[39242]_ ,
    \new_[39245]_ , \new_[39248]_ , \new_[39249]_ , \new_[39250]_ ,
    \new_[39254]_ , \new_[39255]_ , \new_[39258]_ , \new_[39261]_ ,
    \new_[39262]_ , \new_[39263]_ , \new_[39267]_ , \new_[39268]_ ,
    \new_[39271]_ , \new_[39274]_ , \new_[39275]_ , \new_[39276]_ ,
    \new_[39280]_ , \new_[39281]_ , \new_[39284]_ , \new_[39287]_ ,
    \new_[39288]_ , \new_[39289]_ , \new_[39293]_ , \new_[39294]_ ,
    \new_[39297]_ , \new_[39300]_ , \new_[39301]_ , \new_[39302]_ ,
    \new_[39306]_ , \new_[39307]_ , \new_[39310]_ , \new_[39313]_ ,
    \new_[39314]_ , \new_[39315]_ , \new_[39319]_ , \new_[39320]_ ,
    \new_[39323]_ , \new_[39326]_ , \new_[39327]_ , \new_[39328]_ ,
    \new_[39332]_ , \new_[39333]_ , \new_[39336]_ , \new_[39339]_ ,
    \new_[39340]_ , \new_[39341]_ , \new_[39345]_ , \new_[39346]_ ,
    \new_[39349]_ , \new_[39352]_ , \new_[39353]_ , \new_[39354]_ ,
    \new_[39358]_ , \new_[39359]_ , \new_[39362]_ , \new_[39365]_ ,
    \new_[39366]_ , \new_[39367]_ , \new_[39371]_ , \new_[39372]_ ,
    \new_[39375]_ , \new_[39378]_ , \new_[39379]_ , \new_[39380]_ ,
    \new_[39384]_ , \new_[39385]_ , \new_[39388]_ , \new_[39391]_ ,
    \new_[39392]_ , \new_[39393]_ , \new_[39397]_ , \new_[39398]_ ,
    \new_[39401]_ , \new_[39404]_ , \new_[39405]_ , \new_[39406]_ ,
    \new_[39410]_ , \new_[39411]_ , \new_[39414]_ , \new_[39417]_ ,
    \new_[39418]_ , \new_[39419]_ , \new_[39423]_ , \new_[39424]_ ,
    \new_[39427]_ , \new_[39430]_ , \new_[39431]_ , \new_[39432]_ ,
    \new_[39436]_ , \new_[39437]_ , \new_[39440]_ , \new_[39443]_ ,
    \new_[39444]_ , \new_[39445]_ , \new_[39449]_ , \new_[39450]_ ,
    \new_[39453]_ , \new_[39456]_ , \new_[39457]_ , \new_[39458]_ ,
    \new_[39462]_ , \new_[39463]_ , \new_[39466]_ , \new_[39469]_ ,
    \new_[39470]_ , \new_[39471]_ , \new_[39475]_ , \new_[39476]_ ,
    \new_[39479]_ , \new_[39482]_ , \new_[39483]_ , \new_[39484]_ ,
    \new_[39488]_ , \new_[39489]_ , \new_[39492]_ , \new_[39495]_ ,
    \new_[39496]_ , \new_[39497]_ , \new_[39501]_ , \new_[39502]_ ,
    \new_[39505]_ , \new_[39508]_ , \new_[39509]_ , \new_[39510]_ ,
    \new_[39514]_ , \new_[39515]_ , \new_[39518]_ , \new_[39521]_ ,
    \new_[39522]_ , \new_[39523]_ , \new_[39527]_ , \new_[39528]_ ,
    \new_[39531]_ , \new_[39534]_ , \new_[39535]_ , \new_[39536]_ ,
    \new_[39540]_ , \new_[39541]_ , \new_[39544]_ , \new_[39547]_ ,
    \new_[39548]_ , \new_[39549]_ , \new_[39553]_ , \new_[39554]_ ,
    \new_[39557]_ , \new_[39560]_ , \new_[39561]_ , \new_[39562]_ ,
    \new_[39566]_ , \new_[39567]_ , \new_[39570]_ , \new_[39573]_ ,
    \new_[39574]_ , \new_[39575]_ , \new_[39579]_ , \new_[39580]_ ,
    \new_[39583]_ , \new_[39586]_ , \new_[39587]_ , \new_[39588]_ ,
    \new_[39592]_ , \new_[39593]_ , \new_[39596]_ , \new_[39599]_ ,
    \new_[39600]_ , \new_[39601]_ , \new_[39605]_ , \new_[39606]_ ,
    \new_[39609]_ , \new_[39612]_ , \new_[39613]_ , \new_[39614]_ ,
    \new_[39618]_ , \new_[39619]_ , \new_[39622]_ , \new_[39625]_ ,
    \new_[39626]_ , \new_[39627]_ , \new_[39631]_ , \new_[39632]_ ,
    \new_[39635]_ , \new_[39638]_ , \new_[39639]_ , \new_[39640]_ ,
    \new_[39644]_ , \new_[39645]_ , \new_[39648]_ , \new_[39651]_ ,
    \new_[39652]_ , \new_[39653]_ , \new_[39657]_ , \new_[39658]_ ,
    \new_[39661]_ , \new_[39664]_ , \new_[39665]_ , \new_[39666]_ ,
    \new_[39670]_ , \new_[39671]_ , \new_[39674]_ , \new_[39677]_ ,
    \new_[39678]_ , \new_[39679]_ , \new_[39683]_ , \new_[39684]_ ,
    \new_[39687]_ , \new_[39690]_ , \new_[39691]_ , \new_[39692]_ ,
    \new_[39696]_ , \new_[39697]_ , \new_[39700]_ , \new_[39703]_ ,
    \new_[39704]_ , \new_[39705]_ , \new_[39709]_ , \new_[39710]_ ,
    \new_[39713]_ , \new_[39716]_ , \new_[39717]_ , \new_[39718]_ ,
    \new_[39722]_ , \new_[39723]_ , \new_[39726]_ , \new_[39729]_ ,
    \new_[39730]_ , \new_[39731]_ , \new_[39735]_ , \new_[39736]_ ,
    \new_[39739]_ , \new_[39742]_ , \new_[39743]_ , \new_[39744]_ ,
    \new_[39748]_ , \new_[39749]_ , \new_[39752]_ , \new_[39755]_ ,
    \new_[39756]_ , \new_[39757]_ , \new_[39761]_ , \new_[39762]_ ,
    \new_[39765]_ , \new_[39768]_ , \new_[39769]_ , \new_[39770]_ ,
    \new_[39774]_ , \new_[39775]_ , \new_[39778]_ , \new_[39781]_ ,
    \new_[39782]_ , \new_[39783]_ , \new_[39787]_ , \new_[39788]_ ,
    \new_[39791]_ , \new_[39794]_ , \new_[39795]_ , \new_[39796]_ ,
    \new_[39800]_ , \new_[39801]_ , \new_[39804]_ , \new_[39807]_ ,
    \new_[39808]_ , \new_[39809]_ , \new_[39813]_ , \new_[39814]_ ,
    \new_[39817]_ , \new_[39820]_ , \new_[39821]_ , \new_[39822]_ ,
    \new_[39826]_ , \new_[39827]_ , \new_[39830]_ , \new_[39833]_ ,
    \new_[39834]_ , \new_[39835]_ , \new_[39839]_ , \new_[39840]_ ,
    \new_[39843]_ , \new_[39846]_ , \new_[39847]_ , \new_[39848]_ ,
    \new_[39852]_ , \new_[39853]_ , \new_[39856]_ , \new_[39859]_ ,
    \new_[39860]_ , \new_[39861]_ , \new_[39865]_ , \new_[39866]_ ,
    \new_[39869]_ , \new_[39872]_ , \new_[39873]_ , \new_[39874]_ ,
    \new_[39878]_ , \new_[39879]_ , \new_[39882]_ , \new_[39885]_ ,
    \new_[39886]_ , \new_[39887]_ , \new_[39891]_ , \new_[39892]_ ,
    \new_[39895]_ , \new_[39898]_ , \new_[39899]_ , \new_[39900]_ ,
    \new_[39904]_ , \new_[39905]_ , \new_[39908]_ , \new_[39911]_ ,
    \new_[39912]_ , \new_[39913]_ , \new_[39917]_ , \new_[39918]_ ,
    \new_[39921]_ , \new_[39924]_ , \new_[39925]_ , \new_[39926]_ ,
    \new_[39930]_ , \new_[39931]_ , \new_[39934]_ , \new_[39937]_ ,
    \new_[39938]_ , \new_[39939]_ , \new_[39943]_ , \new_[39944]_ ,
    \new_[39947]_ , \new_[39950]_ , \new_[39951]_ , \new_[39952]_ ,
    \new_[39956]_ , \new_[39957]_ , \new_[39960]_ , \new_[39963]_ ,
    \new_[39964]_ , \new_[39965]_ , \new_[39969]_ , \new_[39970]_ ,
    \new_[39973]_ , \new_[39976]_ , \new_[39977]_ , \new_[39978]_ ,
    \new_[39982]_ , \new_[39983]_ , \new_[39986]_ , \new_[39989]_ ,
    \new_[39990]_ , \new_[39991]_ , \new_[39995]_ , \new_[39996]_ ,
    \new_[39999]_ , \new_[40002]_ , \new_[40003]_ , \new_[40004]_ ,
    \new_[40008]_ , \new_[40009]_ , \new_[40012]_ , \new_[40015]_ ,
    \new_[40016]_ , \new_[40017]_ , \new_[40021]_ , \new_[40022]_ ,
    \new_[40025]_ , \new_[40028]_ , \new_[40029]_ , \new_[40030]_ ,
    \new_[40034]_ , \new_[40035]_ , \new_[40038]_ , \new_[40041]_ ,
    \new_[40042]_ , \new_[40043]_ , \new_[40047]_ , \new_[40048]_ ,
    \new_[40051]_ , \new_[40054]_ , \new_[40055]_ , \new_[40056]_ ,
    \new_[40060]_ , \new_[40061]_ , \new_[40064]_ , \new_[40067]_ ,
    \new_[40068]_ , \new_[40069]_ , \new_[40073]_ , \new_[40074]_ ,
    \new_[40077]_ , \new_[40080]_ , \new_[40081]_ , \new_[40082]_ ,
    \new_[40086]_ , \new_[40087]_ , \new_[40090]_ , \new_[40093]_ ,
    \new_[40094]_ , \new_[40095]_ , \new_[40099]_ , \new_[40100]_ ,
    \new_[40103]_ , \new_[40106]_ , \new_[40107]_ , \new_[40108]_ ,
    \new_[40112]_ , \new_[40113]_ , \new_[40116]_ , \new_[40119]_ ,
    \new_[40120]_ , \new_[40121]_ , \new_[40125]_ , \new_[40126]_ ,
    \new_[40129]_ , \new_[40132]_ , \new_[40133]_ , \new_[40134]_ ,
    \new_[40138]_ , \new_[40139]_ , \new_[40142]_ , \new_[40145]_ ,
    \new_[40146]_ , \new_[40147]_ , \new_[40151]_ , \new_[40152]_ ,
    \new_[40155]_ , \new_[40158]_ , \new_[40159]_ , \new_[40160]_ ,
    \new_[40164]_ , \new_[40165]_ , \new_[40168]_ , \new_[40171]_ ,
    \new_[40172]_ , \new_[40173]_ , \new_[40177]_ , \new_[40178]_ ,
    \new_[40181]_ , \new_[40184]_ , \new_[40185]_ , \new_[40186]_ ,
    \new_[40190]_ , \new_[40191]_ , \new_[40194]_ , \new_[40197]_ ,
    \new_[40198]_ , \new_[40199]_ , \new_[40203]_ , \new_[40204]_ ,
    \new_[40207]_ , \new_[40210]_ , \new_[40211]_ , \new_[40212]_ ,
    \new_[40216]_ , \new_[40217]_ , \new_[40220]_ , \new_[40223]_ ,
    \new_[40224]_ , \new_[40225]_ , \new_[40229]_ , \new_[40230]_ ,
    \new_[40233]_ , \new_[40236]_ , \new_[40237]_ , \new_[40238]_ ,
    \new_[40242]_ , \new_[40243]_ , \new_[40246]_ , \new_[40249]_ ,
    \new_[40250]_ , \new_[40251]_ , \new_[40255]_ , \new_[40256]_ ,
    \new_[40259]_ , \new_[40262]_ , \new_[40263]_ , \new_[40264]_ ,
    \new_[40268]_ , \new_[40269]_ , \new_[40272]_ , \new_[40275]_ ,
    \new_[40276]_ , \new_[40277]_ , \new_[40281]_ , \new_[40282]_ ,
    \new_[40285]_ , \new_[40288]_ , \new_[40289]_ , \new_[40290]_ ,
    \new_[40294]_ , \new_[40295]_ , \new_[40298]_ , \new_[40301]_ ,
    \new_[40302]_ , \new_[40303]_ , \new_[40307]_ , \new_[40308]_ ,
    \new_[40311]_ , \new_[40314]_ , \new_[40315]_ , \new_[40316]_ ,
    \new_[40320]_ , \new_[40321]_ , \new_[40324]_ , \new_[40327]_ ,
    \new_[40328]_ , \new_[40329]_ , \new_[40333]_ , \new_[40334]_ ,
    \new_[40337]_ , \new_[40340]_ , \new_[40341]_ , \new_[40342]_ ,
    \new_[40346]_ , \new_[40347]_ , \new_[40350]_ , \new_[40353]_ ,
    \new_[40354]_ , \new_[40355]_ , \new_[40359]_ , \new_[40360]_ ,
    \new_[40363]_ , \new_[40366]_ , \new_[40367]_ , \new_[40368]_ ,
    \new_[40372]_ , \new_[40373]_ , \new_[40376]_ , \new_[40379]_ ,
    \new_[40380]_ , \new_[40381]_ , \new_[40385]_ , \new_[40386]_ ,
    \new_[40389]_ , \new_[40392]_ , \new_[40393]_ , \new_[40394]_ ,
    \new_[40398]_ , \new_[40399]_ , \new_[40402]_ , \new_[40405]_ ,
    \new_[40406]_ , \new_[40407]_ , \new_[40411]_ , \new_[40412]_ ,
    \new_[40415]_ , \new_[40418]_ , \new_[40419]_ , \new_[40420]_ ,
    \new_[40424]_ , \new_[40425]_ , \new_[40428]_ , \new_[40431]_ ,
    \new_[40432]_ , \new_[40433]_ , \new_[40437]_ , \new_[40438]_ ,
    \new_[40441]_ , \new_[40444]_ , \new_[40445]_ , \new_[40446]_ ,
    \new_[40450]_ , \new_[40451]_ , \new_[40454]_ , \new_[40457]_ ,
    \new_[40458]_ , \new_[40459]_ , \new_[40463]_ , \new_[40464]_ ,
    \new_[40467]_ , \new_[40470]_ , \new_[40471]_ , \new_[40472]_ ,
    \new_[40476]_ , \new_[40477]_ , \new_[40480]_ , \new_[40483]_ ,
    \new_[40484]_ , \new_[40485]_ , \new_[40489]_ , \new_[40490]_ ,
    \new_[40493]_ , \new_[40496]_ , \new_[40497]_ , \new_[40498]_ ,
    \new_[40502]_ , \new_[40503]_ , \new_[40506]_ , \new_[40509]_ ,
    \new_[40510]_ , \new_[40511]_ , \new_[40515]_ , \new_[40516]_ ,
    \new_[40519]_ , \new_[40522]_ , \new_[40523]_ , \new_[40524]_ ,
    \new_[40528]_ , \new_[40529]_ , \new_[40532]_ , \new_[40535]_ ,
    \new_[40536]_ , \new_[40537]_ , \new_[40541]_ , \new_[40542]_ ,
    \new_[40545]_ , \new_[40548]_ , \new_[40549]_ , \new_[40550]_ ,
    \new_[40554]_ , \new_[40555]_ , \new_[40558]_ , \new_[40561]_ ,
    \new_[40562]_ , \new_[40563]_ , \new_[40567]_ , \new_[40568]_ ,
    \new_[40571]_ , \new_[40574]_ , \new_[40575]_ , \new_[40576]_ ,
    \new_[40580]_ , \new_[40581]_ , \new_[40584]_ , \new_[40587]_ ,
    \new_[40588]_ , \new_[40589]_ , \new_[40593]_ , \new_[40594]_ ,
    \new_[40597]_ , \new_[40600]_ , \new_[40601]_ , \new_[40602]_ ,
    \new_[40606]_ , \new_[40607]_ , \new_[40610]_ , \new_[40613]_ ,
    \new_[40614]_ , \new_[40615]_ , \new_[40619]_ , \new_[40620]_ ,
    \new_[40623]_ , \new_[40626]_ , \new_[40627]_ , \new_[40628]_ ,
    \new_[40632]_ , \new_[40633]_ , \new_[40636]_ , \new_[40639]_ ,
    \new_[40640]_ , \new_[40641]_ , \new_[40645]_ , \new_[40646]_ ,
    \new_[40649]_ , \new_[40652]_ , \new_[40653]_ , \new_[40654]_ ,
    \new_[40658]_ , \new_[40659]_ , \new_[40662]_ , \new_[40665]_ ,
    \new_[40666]_ , \new_[40667]_ , \new_[40671]_ , \new_[40672]_ ,
    \new_[40675]_ , \new_[40678]_ , \new_[40679]_ , \new_[40680]_ ,
    \new_[40684]_ , \new_[40685]_ , \new_[40688]_ , \new_[40691]_ ,
    \new_[40692]_ , \new_[40693]_ , \new_[40697]_ , \new_[40698]_ ,
    \new_[40701]_ , \new_[40704]_ , \new_[40705]_ , \new_[40706]_ ,
    \new_[40710]_ , \new_[40711]_ , \new_[40714]_ , \new_[40717]_ ,
    \new_[40718]_ , \new_[40719]_ , \new_[40723]_ , \new_[40724]_ ,
    \new_[40727]_ , \new_[40730]_ , \new_[40731]_ , \new_[40732]_ ,
    \new_[40736]_ , \new_[40737]_ , \new_[40740]_ , \new_[40743]_ ,
    \new_[40744]_ , \new_[40745]_ , \new_[40749]_ , \new_[40750]_ ,
    \new_[40753]_ , \new_[40756]_ , \new_[40757]_ , \new_[40758]_ ,
    \new_[40762]_ , \new_[40763]_ , \new_[40766]_ , \new_[40769]_ ,
    \new_[40770]_ , \new_[40771]_ , \new_[40775]_ , \new_[40776]_ ,
    \new_[40779]_ , \new_[40782]_ , \new_[40783]_ , \new_[40784]_ ,
    \new_[40788]_ , \new_[40789]_ , \new_[40792]_ , \new_[40795]_ ,
    \new_[40796]_ , \new_[40797]_ , \new_[40801]_ , \new_[40802]_ ,
    \new_[40805]_ , \new_[40808]_ , \new_[40809]_ , \new_[40810]_ ,
    \new_[40814]_ , \new_[40815]_ , \new_[40818]_ , \new_[40821]_ ,
    \new_[40822]_ , \new_[40823]_ , \new_[40827]_ , \new_[40828]_ ,
    \new_[40831]_ , \new_[40834]_ , \new_[40835]_ , \new_[40836]_ ,
    \new_[40840]_ , \new_[40841]_ , \new_[40844]_ , \new_[40847]_ ,
    \new_[40848]_ , \new_[40849]_ , \new_[40853]_ , \new_[40854]_ ,
    \new_[40857]_ , \new_[40860]_ , \new_[40861]_ , \new_[40862]_ ,
    \new_[40866]_ , \new_[40867]_ , \new_[40870]_ , \new_[40873]_ ,
    \new_[40874]_ , \new_[40875]_ , \new_[40879]_ , \new_[40880]_ ,
    \new_[40883]_ , \new_[40886]_ , \new_[40887]_ , \new_[40888]_ ,
    \new_[40892]_ , \new_[40893]_ , \new_[40896]_ , \new_[40899]_ ,
    \new_[40900]_ , \new_[40901]_ , \new_[40905]_ , \new_[40906]_ ,
    \new_[40909]_ , \new_[40912]_ , \new_[40913]_ , \new_[40914]_ ,
    \new_[40918]_ , \new_[40919]_ , \new_[40922]_ , \new_[40925]_ ,
    \new_[40926]_ , \new_[40927]_ , \new_[40931]_ , \new_[40932]_ ,
    \new_[40935]_ , \new_[40938]_ , \new_[40939]_ , \new_[40940]_ ,
    \new_[40944]_ , \new_[40945]_ , \new_[40948]_ , \new_[40951]_ ,
    \new_[40952]_ , \new_[40953]_ , \new_[40957]_ , \new_[40958]_ ,
    \new_[40961]_ , \new_[40964]_ , \new_[40965]_ , \new_[40966]_ ,
    \new_[40970]_ , \new_[40971]_ , \new_[40974]_ , \new_[40977]_ ,
    \new_[40978]_ , \new_[40979]_ , \new_[40983]_ , \new_[40984]_ ,
    \new_[40987]_ , \new_[40990]_ , \new_[40991]_ , \new_[40992]_ ,
    \new_[40996]_ , \new_[40997]_ , \new_[41000]_ , \new_[41003]_ ,
    \new_[41004]_ , \new_[41005]_ , \new_[41009]_ , \new_[41010]_ ,
    \new_[41013]_ , \new_[41016]_ , \new_[41017]_ , \new_[41018]_ ,
    \new_[41022]_ , \new_[41023]_ , \new_[41026]_ , \new_[41029]_ ,
    \new_[41030]_ , \new_[41031]_ , \new_[41035]_ , \new_[41036]_ ,
    \new_[41039]_ , \new_[41042]_ , \new_[41043]_ , \new_[41044]_ ,
    \new_[41048]_ , \new_[41049]_ , \new_[41052]_ , \new_[41055]_ ,
    \new_[41056]_ , \new_[41057]_ , \new_[41061]_ , \new_[41062]_ ,
    \new_[41065]_ , \new_[41068]_ , \new_[41069]_ , \new_[41070]_ ,
    \new_[41074]_ , \new_[41075]_ , \new_[41078]_ , \new_[41081]_ ,
    \new_[41082]_ , \new_[41083]_ , \new_[41087]_ , \new_[41088]_ ,
    \new_[41091]_ , \new_[41094]_ , \new_[41095]_ , \new_[41096]_ ,
    \new_[41100]_ , \new_[41101]_ , \new_[41104]_ , \new_[41107]_ ,
    \new_[41108]_ , \new_[41109]_ , \new_[41113]_ , \new_[41114]_ ,
    \new_[41117]_ , \new_[41120]_ , \new_[41121]_ , \new_[41122]_ ,
    \new_[41126]_ , \new_[41127]_ , \new_[41130]_ , \new_[41133]_ ,
    \new_[41134]_ , \new_[41135]_ , \new_[41139]_ , \new_[41140]_ ,
    \new_[41143]_ , \new_[41146]_ , \new_[41147]_ , \new_[41148]_ ,
    \new_[41152]_ , \new_[41153]_ , \new_[41156]_ , \new_[41159]_ ,
    \new_[41160]_ , \new_[41161]_ , \new_[41165]_ , \new_[41166]_ ,
    \new_[41169]_ , \new_[41172]_ , \new_[41173]_ , \new_[41174]_ ,
    \new_[41178]_ , \new_[41179]_ , \new_[41182]_ , \new_[41185]_ ,
    \new_[41186]_ , \new_[41187]_ , \new_[41191]_ , \new_[41192]_ ,
    \new_[41195]_ , \new_[41198]_ , \new_[41199]_ , \new_[41200]_ ,
    \new_[41204]_ , \new_[41205]_ , \new_[41208]_ , \new_[41211]_ ,
    \new_[41212]_ , \new_[41213]_ , \new_[41217]_ , \new_[41218]_ ,
    \new_[41221]_ , \new_[41224]_ , \new_[41225]_ , \new_[41226]_ ,
    \new_[41230]_ , \new_[41231]_ , \new_[41234]_ , \new_[41237]_ ,
    \new_[41238]_ , \new_[41239]_ , \new_[41243]_ , \new_[41244]_ ,
    \new_[41247]_ , \new_[41250]_ , \new_[41251]_ , \new_[41252]_ ,
    \new_[41256]_ , \new_[41257]_ , \new_[41260]_ , \new_[41263]_ ,
    \new_[41264]_ , \new_[41265]_ , \new_[41269]_ , \new_[41270]_ ,
    \new_[41273]_ , \new_[41276]_ , \new_[41277]_ , \new_[41278]_ ,
    \new_[41282]_ , \new_[41283]_ , \new_[41286]_ , \new_[41289]_ ,
    \new_[41290]_ , \new_[41291]_ , \new_[41295]_ , \new_[41296]_ ,
    \new_[41299]_ , \new_[41302]_ , \new_[41303]_ , \new_[41304]_ ,
    \new_[41308]_ , \new_[41309]_ , \new_[41312]_ , \new_[41315]_ ,
    \new_[41316]_ , \new_[41317]_ , \new_[41321]_ , \new_[41322]_ ,
    \new_[41325]_ , \new_[41328]_ , \new_[41329]_ , \new_[41330]_ ,
    \new_[41334]_ , \new_[41335]_ , \new_[41338]_ , \new_[41341]_ ,
    \new_[41342]_ , \new_[41343]_ , \new_[41347]_ , \new_[41348]_ ,
    \new_[41351]_ , \new_[41354]_ , \new_[41355]_ , \new_[41356]_ ,
    \new_[41360]_ , \new_[41361]_ , \new_[41364]_ , \new_[41367]_ ,
    \new_[41368]_ , \new_[41369]_ , \new_[41373]_ , \new_[41374]_ ,
    \new_[41377]_ , \new_[41380]_ , \new_[41381]_ , \new_[41382]_ ,
    \new_[41386]_ , \new_[41387]_ , \new_[41390]_ , \new_[41393]_ ,
    \new_[41394]_ , \new_[41395]_ , \new_[41399]_ , \new_[41400]_ ,
    \new_[41403]_ , \new_[41406]_ , \new_[41407]_ , \new_[41408]_ ,
    \new_[41412]_ , \new_[41413]_ , \new_[41416]_ , \new_[41419]_ ,
    \new_[41420]_ , \new_[41421]_ , \new_[41425]_ , \new_[41426]_ ,
    \new_[41429]_ , \new_[41432]_ , \new_[41433]_ , \new_[41434]_ ,
    \new_[41438]_ , \new_[41439]_ , \new_[41442]_ , \new_[41445]_ ,
    \new_[41446]_ , \new_[41447]_ , \new_[41451]_ , \new_[41452]_ ,
    \new_[41455]_ , \new_[41458]_ , \new_[41459]_ , \new_[41460]_ ,
    \new_[41464]_ , \new_[41465]_ , \new_[41468]_ , \new_[41471]_ ,
    \new_[41472]_ , \new_[41473]_ , \new_[41477]_ , \new_[41478]_ ,
    \new_[41481]_ , \new_[41484]_ , \new_[41485]_ , \new_[41486]_ ,
    \new_[41490]_ , \new_[41491]_ , \new_[41494]_ , \new_[41497]_ ,
    \new_[41498]_ , \new_[41499]_ , \new_[41503]_ , \new_[41504]_ ,
    \new_[41507]_ , \new_[41510]_ , \new_[41511]_ , \new_[41512]_ ,
    \new_[41516]_ , \new_[41517]_ , \new_[41520]_ , \new_[41523]_ ,
    \new_[41524]_ , \new_[41525]_ , \new_[41529]_ , \new_[41530]_ ,
    \new_[41533]_ , \new_[41536]_ , \new_[41537]_ , \new_[41538]_ ,
    \new_[41542]_ , \new_[41543]_ , \new_[41546]_ , \new_[41549]_ ,
    \new_[41550]_ , \new_[41551]_ , \new_[41555]_ , \new_[41556]_ ,
    \new_[41559]_ , \new_[41562]_ , \new_[41563]_ , \new_[41564]_ ,
    \new_[41568]_ , \new_[41569]_ , \new_[41572]_ , \new_[41575]_ ,
    \new_[41576]_ , \new_[41577]_ , \new_[41581]_ , \new_[41582]_ ,
    \new_[41585]_ , \new_[41588]_ , \new_[41589]_ , \new_[41590]_ ,
    \new_[41594]_ , \new_[41595]_ , \new_[41598]_ , \new_[41601]_ ,
    \new_[41602]_ , \new_[41603]_ , \new_[41607]_ , \new_[41608]_ ,
    \new_[41611]_ , \new_[41614]_ , \new_[41615]_ , \new_[41616]_ ,
    \new_[41620]_ , \new_[41621]_ , \new_[41624]_ , \new_[41627]_ ,
    \new_[41628]_ , \new_[41629]_ , \new_[41633]_ , \new_[41634]_ ,
    \new_[41637]_ , \new_[41640]_ , \new_[41641]_ , \new_[41642]_ ,
    \new_[41646]_ , \new_[41647]_ , \new_[41650]_ , \new_[41653]_ ,
    \new_[41654]_ , \new_[41655]_ , \new_[41659]_ , \new_[41660]_ ,
    \new_[41663]_ , \new_[41666]_ , \new_[41667]_ , \new_[41668]_ ,
    \new_[41672]_ , \new_[41673]_ , \new_[41676]_ , \new_[41679]_ ,
    \new_[41680]_ , \new_[41681]_ , \new_[41685]_ , \new_[41686]_ ,
    \new_[41689]_ , \new_[41692]_ , \new_[41693]_ , \new_[41694]_ ,
    \new_[41698]_ , \new_[41699]_ , \new_[41702]_ , \new_[41705]_ ,
    \new_[41706]_ , \new_[41707]_ , \new_[41711]_ , \new_[41712]_ ,
    \new_[41715]_ , \new_[41718]_ , \new_[41719]_ , \new_[41720]_ ,
    \new_[41724]_ , \new_[41725]_ , \new_[41728]_ , \new_[41731]_ ,
    \new_[41732]_ , \new_[41733]_ , \new_[41737]_ , \new_[41738]_ ,
    \new_[41741]_ , \new_[41744]_ , \new_[41745]_ , \new_[41746]_ ,
    \new_[41750]_ , \new_[41751]_ , \new_[41754]_ , \new_[41757]_ ,
    \new_[41758]_ , \new_[41759]_ , \new_[41763]_ , \new_[41764]_ ,
    \new_[41767]_ , \new_[41770]_ , \new_[41771]_ , \new_[41772]_ ,
    \new_[41776]_ , \new_[41777]_ , \new_[41780]_ , \new_[41783]_ ,
    \new_[41784]_ , \new_[41785]_ , \new_[41789]_ , \new_[41790]_ ,
    \new_[41793]_ , \new_[41796]_ , \new_[41797]_ , \new_[41798]_ ,
    \new_[41802]_ , \new_[41803]_ , \new_[41806]_ , \new_[41809]_ ,
    \new_[41810]_ , \new_[41811]_ , \new_[41815]_ , \new_[41816]_ ,
    \new_[41819]_ , \new_[41822]_ , \new_[41823]_ , \new_[41824]_ ,
    \new_[41828]_ , \new_[41829]_ , \new_[41832]_ , \new_[41835]_ ,
    \new_[41836]_ , \new_[41837]_ , \new_[41841]_ , \new_[41842]_ ,
    \new_[41845]_ , \new_[41848]_ , \new_[41849]_ , \new_[41850]_ ,
    \new_[41854]_ , \new_[41855]_ , \new_[41858]_ , \new_[41861]_ ,
    \new_[41862]_ , \new_[41863]_ , \new_[41867]_ , \new_[41868]_ ,
    \new_[41871]_ , \new_[41874]_ , \new_[41875]_ , \new_[41876]_ ,
    \new_[41880]_ , \new_[41881]_ , \new_[41884]_ , \new_[41887]_ ,
    \new_[41888]_ , \new_[41889]_ , \new_[41893]_ , \new_[41894]_ ,
    \new_[41897]_ , \new_[41900]_ , \new_[41901]_ , \new_[41902]_ ,
    \new_[41906]_ , \new_[41907]_ , \new_[41910]_ , \new_[41913]_ ,
    \new_[41914]_ , \new_[41915]_ , \new_[41919]_ , \new_[41920]_ ,
    \new_[41923]_ , \new_[41926]_ , \new_[41927]_ , \new_[41928]_ ,
    \new_[41932]_ , \new_[41933]_ , \new_[41936]_ , \new_[41939]_ ,
    \new_[41940]_ , \new_[41941]_ , \new_[41945]_ , \new_[41946]_ ,
    \new_[41949]_ , \new_[41952]_ , \new_[41953]_ , \new_[41954]_ ,
    \new_[41958]_ , \new_[41959]_ , \new_[41962]_ , \new_[41965]_ ,
    \new_[41966]_ , \new_[41967]_ , \new_[41971]_ , \new_[41972]_ ,
    \new_[41975]_ , \new_[41978]_ , \new_[41979]_ , \new_[41980]_ ,
    \new_[41984]_ , \new_[41985]_ , \new_[41988]_ , \new_[41991]_ ,
    \new_[41992]_ , \new_[41993]_ , \new_[41997]_ , \new_[41998]_ ,
    \new_[42001]_ , \new_[42004]_ , \new_[42005]_ , \new_[42006]_ ,
    \new_[42010]_ , \new_[42011]_ , \new_[42014]_ , \new_[42017]_ ,
    \new_[42018]_ , \new_[42019]_ , \new_[42023]_ , \new_[42024]_ ,
    \new_[42027]_ , \new_[42030]_ , \new_[42031]_ , \new_[42032]_ ,
    \new_[42036]_ , \new_[42037]_ , \new_[42040]_ , \new_[42043]_ ,
    \new_[42044]_ , \new_[42045]_ , \new_[42049]_ , \new_[42050]_ ,
    \new_[42053]_ , \new_[42056]_ , \new_[42057]_ , \new_[42058]_ ,
    \new_[42062]_ , \new_[42063]_ , \new_[42066]_ , \new_[42069]_ ,
    \new_[42070]_ , \new_[42071]_ , \new_[42075]_ , \new_[42076]_ ,
    \new_[42079]_ , \new_[42082]_ , \new_[42083]_ , \new_[42084]_ ,
    \new_[42088]_ , \new_[42089]_ , \new_[42092]_ , \new_[42095]_ ,
    \new_[42096]_ , \new_[42097]_ , \new_[42101]_ , \new_[42102]_ ,
    \new_[42105]_ , \new_[42108]_ , \new_[42109]_ , \new_[42110]_ ,
    \new_[42114]_ , \new_[42115]_ , \new_[42118]_ , \new_[42121]_ ,
    \new_[42122]_ , \new_[42123]_ , \new_[42127]_ , \new_[42128]_ ,
    \new_[42131]_ , \new_[42134]_ , \new_[42135]_ , \new_[42136]_ ,
    \new_[42140]_ , \new_[42141]_ , \new_[42144]_ , \new_[42147]_ ,
    \new_[42148]_ , \new_[42149]_ , \new_[42153]_ , \new_[42154]_ ,
    \new_[42157]_ , \new_[42160]_ , \new_[42161]_ , \new_[42162]_ ,
    \new_[42166]_ , \new_[42167]_ , \new_[42170]_ , \new_[42173]_ ,
    \new_[42174]_ , \new_[42175]_ , \new_[42179]_ , \new_[42180]_ ,
    \new_[42183]_ , \new_[42186]_ , \new_[42187]_ , \new_[42188]_ ,
    \new_[42192]_ , \new_[42193]_ , \new_[42196]_ , \new_[42199]_ ,
    \new_[42200]_ , \new_[42201]_ , \new_[42205]_ , \new_[42206]_ ,
    \new_[42209]_ , \new_[42212]_ , \new_[42213]_ , \new_[42214]_ ,
    \new_[42218]_ , \new_[42219]_ , \new_[42222]_ , \new_[42225]_ ,
    \new_[42226]_ , \new_[42227]_ , \new_[42231]_ , \new_[42232]_ ,
    \new_[42235]_ , \new_[42238]_ , \new_[42239]_ , \new_[42240]_ ,
    \new_[42244]_ , \new_[42245]_ , \new_[42248]_ , \new_[42251]_ ,
    \new_[42252]_ , \new_[42253]_ , \new_[42257]_ , \new_[42258]_ ,
    \new_[42261]_ , \new_[42264]_ , \new_[42265]_ , \new_[42266]_ ,
    \new_[42270]_ , \new_[42271]_ , \new_[42274]_ , \new_[42277]_ ,
    \new_[42278]_ , \new_[42279]_ , \new_[42283]_ , \new_[42284]_ ,
    \new_[42287]_ , \new_[42290]_ , \new_[42291]_ , \new_[42292]_ ,
    \new_[42296]_ , \new_[42297]_ , \new_[42300]_ , \new_[42303]_ ,
    \new_[42304]_ , \new_[42305]_ , \new_[42309]_ , \new_[42310]_ ,
    \new_[42313]_ , \new_[42316]_ , \new_[42317]_ , \new_[42318]_ ,
    \new_[42322]_ , \new_[42323]_ , \new_[42326]_ , \new_[42329]_ ,
    \new_[42330]_ , \new_[42331]_ , \new_[42335]_ , \new_[42336]_ ,
    \new_[42339]_ , \new_[42342]_ , \new_[42343]_ , \new_[42344]_ ,
    \new_[42348]_ , \new_[42349]_ , \new_[42352]_ , \new_[42355]_ ,
    \new_[42356]_ , \new_[42357]_ , \new_[42361]_ , \new_[42362]_ ,
    \new_[42365]_ , \new_[42368]_ , \new_[42369]_ , \new_[42370]_ ,
    \new_[42374]_ , \new_[42375]_ , \new_[42378]_ , \new_[42381]_ ,
    \new_[42382]_ , \new_[42383]_ , \new_[42387]_ , \new_[42388]_ ,
    \new_[42391]_ , \new_[42394]_ , \new_[42395]_ , \new_[42396]_ ,
    \new_[42400]_ , \new_[42401]_ , \new_[42404]_ , \new_[42407]_ ,
    \new_[42408]_ , \new_[42409]_ , \new_[42413]_ , \new_[42414]_ ,
    \new_[42417]_ , \new_[42420]_ , \new_[42421]_ , \new_[42422]_ ,
    \new_[42426]_ , \new_[42427]_ , \new_[42430]_ , \new_[42433]_ ,
    \new_[42434]_ , \new_[42435]_ , \new_[42439]_ , \new_[42440]_ ,
    \new_[42443]_ , \new_[42446]_ , \new_[42447]_ , \new_[42448]_ ,
    \new_[42452]_ , \new_[42453]_ , \new_[42456]_ , \new_[42459]_ ,
    \new_[42460]_ , \new_[42461]_ , \new_[42465]_ , \new_[42466]_ ,
    \new_[42469]_ , \new_[42472]_ , \new_[42473]_ , \new_[42474]_ ,
    \new_[42478]_ , \new_[42479]_ , \new_[42482]_ , \new_[42485]_ ,
    \new_[42486]_ , \new_[42487]_ , \new_[42491]_ , \new_[42492]_ ,
    \new_[42495]_ , \new_[42498]_ , \new_[42499]_ , \new_[42500]_ ,
    \new_[42504]_ , \new_[42505]_ , \new_[42508]_ , \new_[42511]_ ,
    \new_[42512]_ , \new_[42513]_ , \new_[42517]_ , \new_[42518]_ ,
    \new_[42521]_ , \new_[42524]_ , \new_[42525]_ , \new_[42526]_ ,
    \new_[42530]_ , \new_[42531]_ , \new_[42534]_ , \new_[42537]_ ,
    \new_[42538]_ , \new_[42539]_ , \new_[42543]_ , \new_[42544]_ ,
    \new_[42547]_ , \new_[42550]_ , \new_[42551]_ , \new_[42552]_ ,
    \new_[42556]_ , \new_[42557]_ , \new_[42560]_ , \new_[42563]_ ,
    \new_[42564]_ , \new_[42565]_ , \new_[42569]_ , \new_[42570]_ ,
    \new_[42573]_ , \new_[42576]_ , \new_[42577]_ , \new_[42578]_ ,
    \new_[42582]_ , \new_[42583]_ , \new_[42586]_ , \new_[42589]_ ,
    \new_[42590]_ , \new_[42591]_ , \new_[42595]_ , \new_[42596]_ ,
    \new_[42599]_ , \new_[42602]_ , \new_[42603]_ , \new_[42604]_ ,
    \new_[42608]_ , \new_[42609]_ , \new_[42612]_ , \new_[42615]_ ,
    \new_[42616]_ , \new_[42617]_ , \new_[42621]_ , \new_[42622]_ ,
    \new_[42625]_ , \new_[42628]_ , \new_[42629]_ , \new_[42630]_ ,
    \new_[42634]_ , \new_[42635]_ , \new_[42638]_ , \new_[42641]_ ,
    \new_[42642]_ , \new_[42643]_ , \new_[42647]_ , \new_[42648]_ ,
    \new_[42651]_ , \new_[42654]_ , \new_[42655]_ , \new_[42656]_ ,
    \new_[42660]_ , \new_[42661]_ , \new_[42664]_ , \new_[42667]_ ,
    \new_[42668]_ , \new_[42669]_ , \new_[42673]_ , \new_[42674]_ ,
    \new_[42677]_ , \new_[42680]_ , \new_[42681]_ , \new_[42682]_ ,
    \new_[42686]_ , \new_[42687]_ , \new_[42690]_ , \new_[42693]_ ,
    \new_[42694]_ , \new_[42695]_ , \new_[42699]_ , \new_[42700]_ ,
    \new_[42703]_ , \new_[42706]_ , \new_[42707]_ , \new_[42708]_ ,
    \new_[42712]_ , \new_[42713]_ , \new_[42716]_ , \new_[42719]_ ,
    \new_[42720]_ , \new_[42721]_ , \new_[42725]_ , \new_[42726]_ ,
    \new_[42729]_ , \new_[42732]_ , \new_[42733]_ , \new_[42734]_ ,
    \new_[42738]_ , \new_[42739]_ , \new_[42742]_ , \new_[42745]_ ,
    \new_[42746]_ , \new_[42747]_ , \new_[42751]_ , \new_[42752]_ ,
    \new_[42755]_ , \new_[42758]_ , \new_[42759]_ , \new_[42760]_ ,
    \new_[42764]_ , \new_[42765]_ , \new_[42768]_ , \new_[42771]_ ,
    \new_[42772]_ , \new_[42773]_ , \new_[42777]_ , \new_[42778]_ ,
    \new_[42781]_ , \new_[42784]_ , \new_[42785]_ , \new_[42786]_ ,
    \new_[42790]_ , \new_[42791]_ , \new_[42794]_ , \new_[42797]_ ,
    \new_[42798]_ , \new_[42799]_ , \new_[42803]_ , \new_[42804]_ ,
    \new_[42807]_ , \new_[42810]_ , \new_[42811]_ , \new_[42812]_ ,
    \new_[42816]_ , \new_[42817]_ , \new_[42820]_ , \new_[42823]_ ,
    \new_[42824]_ , \new_[42825]_ , \new_[42829]_ , \new_[42830]_ ,
    \new_[42833]_ , \new_[42836]_ , \new_[42837]_ , \new_[42838]_ ,
    \new_[42842]_ , \new_[42843]_ , \new_[42846]_ , \new_[42849]_ ,
    \new_[42850]_ , \new_[42851]_ , \new_[42855]_ , \new_[42856]_ ,
    \new_[42859]_ , \new_[42862]_ , \new_[42863]_ , \new_[42864]_ ,
    \new_[42868]_ , \new_[42869]_ , \new_[42872]_ , \new_[42875]_ ,
    \new_[42876]_ , \new_[42877]_ , \new_[42881]_ , \new_[42882]_ ,
    \new_[42885]_ , \new_[42888]_ , \new_[42889]_ , \new_[42890]_ ,
    \new_[42894]_ , \new_[42895]_ , \new_[42898]_ , \new_[42901]_ ,
    \new_[42902]_ , \new_[42903]_ , \new_[42907]_ , \new_[42908]_ ,
    \new_[42911]_ , \new_[42914]_ , \new_[42915]_ , \new_[42916]_ ,
    \new_[42920]_ , \new_[42921]_ , \new_[42924]_ , \new_[42927]_ ,
    \new_[42928]_ , \new_[42929]_ , \new_[42933]_ , \new_[42934]_ ,
    \new_[42937]_ , \new_[42940]_ , \new_[42941]_ , \new_[42942]_ ,
    \new_[42946]_ , \new_[42947]_ , \new_[42950]_ , \new_[42953]_ ,
    \new_[42954]_ , \new_[42955]_ , \new_[42959]_ , \new_[42960]_ ,
    \new_[42963]_ , \new_[42966]_ , \new_[42967]_ , \new_[42968]_ ,
    \new_[42972]_ , \new_[42973]_ , \new_[42976]_ , \new_[42979]_ ,
    \new_[42980]_ , \new_[42981]_ , \new_[42985]_ , \new_[42986]_ ,
    \new_[42989]_ , \new_[42992]_ , \new_[42993]_ , \new_[42994]_ ,
    \new_[42998]_ , \new_[42999]_ , \new_[43002]_ , \new_[43005]_ ,
    \new_[43006]_ , \new_[43007]_ , \new_[43011]_ , \new_[43012]_ ,
    \new_[43015]_ , \new_[43018]_ , \new_[43019]_ , \new_[43020]_ ,
    \new_[43024]_ , \new_[43025]_ , \new_[43028]_ , \new_[43031]_ ,
    \new_[43032]_ , \new_[43033]_ , \new_[43037]_ , \new_[43038]_ ,
    \new_[43041]_ , \new_[43044]_ , \new_[43045]_ , \new_[43046]_ ,
    \new_[43050]_ , \new_[43051]_ , \new_[43054]_ , \new_[43057]_ ,
    \new_[43058]_ , \new_[43059]_ , \new_[43063]_ , \new_[43064]_ ,
    \new_[43067]_ , \new_[43070]_ , \new_[43071]_ , \new_[43072]_ ,
    \new_[43076]_ , \new_[43077]_ , \new_[43080]_ , \new_[43083]_ ,
    \new_[43084]_ , \new_[43085]_ , \new_[43089]_ , \new_[43090]_ ,
    \new_[43093]_ , \new_[43096]_ , \new_[43097]_ , \new_[43098]_ ,
    \new_[43102]_ , \new_[43103]_ , \new_[43106]_ , \new_[43109]_ ,
    \new_[43110]_ , \new_[43111]_ , \new_[43115]_ , \new_[43116]_ ,
    \new_[43119]_ , \new_[43122]_ , \new_[43123]_ , \new_[43124]_ ,
    \new_[43128]_ , \new_[43129]_ , \new_[43132]_ , \new_[43135]_ ,
    \new_[43136]_ , \new_[43137]_ , \new_[43141]_ , \new_[43142]_ ,
    \new_[43145]_ , \new_[43148]_ , \new_[43149]_ , \new_[43150]_ ,
    \new_[43154]_ , \new_[43155]_ , \new_[43158]_ , \new_[43161]_ ,
    \new_[43162]_ , \new_[43163]_ , \new_[43167]_ , \new_[43168]_ ,
    \new_[43171]_ , \new_[43174]_ , \new_[43175]_ , \new_[43176]_ ,
    \new_[43180]_ , \new_[43181]_ , \new_[43184]_ , \new_[43187]_ ,
    \new_[43188]_ , \new_[43189]_ , \new_[43193]_ , \new_[43194]_ ,
    \new_[43197]_ , \new_[43200]_ , \new_[43201]_ , \new_[43202]_ ,
    \new_[43206]_ , \new_[43207]_ , \new_[43210]_ , \new_[43213]_ ,
    \new_[43214]_ , \new_[43215]_ , \new_[43219]_ , \new_[43220]_ ,
    \new_[43223]_ , \new_[43226]_ , \new_[43227]_ , \new_[43228]_ ,
    \new_[43232]_ , \new_[43233]_ , \new_[43236]_ , \new_[43239]_ ,
    \new_[43240]_ , \new_[43241]_ , \new_[43245]_ , \new_[43246]_ ,
    \new_[43249]_ , \new_[43252]_ , \new_[43253]_ , \new_[43254]_ ,
    \new_[43258]_ , \new_[43259]_ , \new_[43262]_ , \new_[43265]_ ,
    \new_[43266]_ , \new_[43267]_ , \new_[43271]_ , \new_[43272]_ ,
    \new_[43275]_ , \new_[43278]_ , \new_[43279]_ , \new_[43280]_ ,
    \new_[43284]_ , \new_[43285]_ , \new_[43288]_ , \new_[43291]_ ,
    \new_[43292]_ , \new_[43293]_ , \new_[43297]_ , \new_[43298]_ ,
    \new_[43301]_ , \new_[43304]_ , \new_[43305]_ , \new_[43306]_ ,
    \new_[43310]_ , \new_[43311]_ , \new_[43314]_ , \new_[43317]_ ,
    \new_[43318]_ , \new_[43319]_ , \new_[43323]_ , \new_[43324]_ ,
    \new_[43327]_ , \new_[43330]_ , \new_[43331]_ , \new_[43332]_ ,
    \new_[43336]_ , \new_[43337]_ , \new_[43340]_ , \new_[43343]_ ,
    \new_[43344]_ , \new_[43345]_ , \new_[43349]_ , \new_[43350]_ ,
    \new_[43353]_ , \new_[43356]_ , \new_[43357]_ , \new_[43358]_ ,
    \new_[43362]_ , \new_[43363]_ , \new_[43366]_ , \new_[43369]_ ,
    \new_[43370]_ , \new_[43371]_ , \new_[43375]_ , \new_[43376]_ ,
    \new_[43379]_ , \new_[43382]_ , \new_[43383]_ , \new_[43384]_ ,
    \new_[43388]_ , \new_[43389]_ , \new_[43392]_ , \new_[43395]_ ,
    \new_[43396]_ , \new_[43397]_ , \new_[43401]_ , \new_[43402]_ ,
    \new_[43405]_ , \new_[43408]_ , \new_[43409]_ , \new_[43410]_ ,
    \new_[43414]_ , \new_[43415]_ , \new_[43418]_ , \new_[43421]_ ,
    \new_[43422]_ , \new_[43423]_ , \new_[43427]_ , \new_[43428]_ ,
    \new_[43431]_ , \new_[43434]_ , \new_[43435]_ , \new_[43436]_ ,
    \new_[43440]_ , \new_[43441]_ , \new_[43444]_ , \new_[43447]_ ,
    \new_[43448]_ , \new_[43449]_ , \new_[43453]_ , \new_[43454]_ ,
    \new_[43457]_ , \new_[43460]_ , \new_[43461]_ , \new_[43462]_ ,
    \new_[43466]_ , \new_[43467]_ , \new_[43470]_ , \new_[43473]_ ,
    \new_[43474]_ , \new_[43475]_ , \new_[43479]_ , \new_[43480]_ ,
    \new_[43483]_ , \new_[43486]_ , \new_[43487]_ , \new_[43488]_ ,
    \new_[43492]_ , \new_[43493]_ , \new_[43496]_ , \new_[43499]_ ,
    \new_[43500]_ , \new_[43501]_ , \new_[43505]_ , \new_[43506]_ ,
    \new_[43509]_ , \new_[43512]_ , \new_[43513]_ , \new_[43514]_ ,
    \new_[43518]_ , \new_[43519]_ , \new_[43522]_ , \new_[43525]_ ,
    \new_[43526]_ , \new_[43527]_ , \new_[43531]_ , \new_[43532]_ ,
    \new_[43535]_ , \new_[43538]_ , \new_[43539]_ , \new_[43540]_ ,
    \new_[43544]_ , \new_[43545]_ , \new_[43548]_ , \new_[43551]_ ,
    \new_[43552]_ , \new_[43553]_ , \new_[43557]_ , \new_[43558]_ ,
    \new_[43561]_ , \new_[43564]_ , \new_[43565]_ , \new_[43566]_ ,
    \new_[43570]_ , \new_[43571]_ , \new_[43574]_ , \new_[43577]_ ,
    \new_[43578]_ , \new_[43579]_ , \new_[43583]_ , \new_[43584]_ ,
    \new_[43587]_ , \new_[43590]_ , \new_[43591]_ , \new_[43592]_ ,
    \new_[43596]_ , \new_[43597]_ , \new_[43600]_ , \new_[43603]_ ,
    \new_[43604]_ , \new_[43605]_ , \new_[43609]_ , \new_[43610]_ ,
    \new_[43613]_ , \new_[43616]_ , \new_[43617]_ , \new_[43618]_ ,
    \new_[43622]_ , \new_[43623]_ , \new_[43626]_ , \new_[43629]_ ,
    \new_[43630]_ , \new_[43631]_ , \new_[43635]_ , \new_[43636]_ ,
    \new_[43639]_ , \new_[43642]_ , \new_[43643]_ , \new_[43644]_ ,
    \new_[43648]_ , \new_[43649]_ , \new_[43652]_ , \new_[43655]_ ,
    \new_[43656]_ , \new_[43657]_ , \new_[43661]_ , \new_[43662]_ ,
    \new_[43665]_ , \new_[43668]_ , \new_[43669]_ , \new_[43670]_ ,
    \new_[43674]_ , \new_[43675]_ , \new_[43678]_ , \new_[43681]_ ,
    \new_[43682]_ , \new_[43683]_ , \new_[43687]_ , \new_[43688]_ ,
    \new_[43691]_ , \new_[43694]_ , \new_[43695]_ , \new_[43696]_ ,
    \new_[43700]_ , \new_[43701]_ , \new_[43704]_ , \new_[43707]_ ,
    \new_[43708]_ , \new_[43709]_ , \new_[43713]_ , \new_[43714]_ ,
    \new_[43717]_ , \new_[43720]_ , \new_[43721]_ , \new_[43722]_ ,
    \new_[43726]_ , \new_[43727]_ , \new_[43730]_ , \new_[43733]_ ,
    \new_[43734]_ , \new_[43735]_ , \new_[43739]_ , \new_[43740]_ ,
    \new_[43743]_ , \new_[43746]_ , \new_[43747]_ , \new_[43748]_ ,
    \new_[43752]_ , \new_[43753]_ , \new_[43756]_ , \new_[43759]_ ,
    \new_[43760]_ , \new_[43761]_ , \new_[43765]_ , \new_[43766]_ ,
    \new_[43769]_ , \new_[43772]_ , \new_[43773]_ , \new_[43774]_ ,
    \new_[43778]_ , \new_[43779]_ , \new_[43782]_ , \new_[43785]_ ,
    \new_[43786]_ , \new_[43787]_ , \new_[43791]_ , \new_[43792]_ ,
    \new_[43795]_ , \new_[43798]_ , \new_[43799]_ , \new_[43800]_ ,
    \new_[43804]_ , \new_[43805]_ , \new_[43808]_ , \new_[43811]_ ,
    \new_[43812]_ , \new_[43813]_ , \new_[43817]_ , \new_[43818]_ ,
    \new_[43821]_ , \new_[43824]_ , \new_[43825]_ , \new_[43826]_ ,
    \new_[43830]_ , \new_[43831]_ , \new_[43834]_ , \new_[43837]_ ,
    \new_[43838]_ , \new_[43839]_ , \new_[43843]_ , \new_[43844]_ ,
    \new_[43847]_ , \new_[43850]_ , \new_[43851]_ , \new_[43852]_ ,
    \new_[43856]_ , \new_[43857]_ , \new_[43860]_ , \new_[43863]_ ,
    \new_[43864]_ , \new_[43865]_ , \new_[43869]_ , \new_[43870]_ ,
    \new_[43873]_ , \new_[43876]_ , \new_[43877]_ , \new_[43878]_ ,
    \new_[43882]_ , \new_[43883]_ , \new_[43886]_ , \new_[43889]_ ,
    \new_[43890]_ , \new_[43891]_ , \new_[43895]_ , \new_[43896]_ ,
    \new_[43899]_ , \new_[43902]_ , \new_[43903]_ , \new_[43904]_ ,
    \new_[43908]_ , \new_[43909]_ , \new_[43912]_ , \new_[43915]_ ,
    \new_[43916]_ , \new_[43917]_ , \new_[43921]_ , \new_[43922]_ ,
    \new_[43925]_ , \new_[43928]_ , \new_[43929]_ , \new_[43930]_ ,
    \new_[43934]_ , \new_[43935]_ , \new_[43938]_ , \new_[43941]_ ,
    \new_[43942]_ , \new_[43943]_ , \new_[43947]_ , \new_[43948]_ ,
    \new_[43951]_ , \new_[43954]_ , \new_[43955]_ , \new_[43956]_ ,
    \new_[43960]_ , \new_[43961]_ , \new_[43964]_ , \new_[43967]_ ,
    \new_[43968]_ , \new_[43969]_ , \new_[43973]_ , \new_[43974]_ ,
    \new_[43977]_ , \new_[43980]_ , \new_[43981]_ , \new_[43982]_ ,
    \new_[43986]_ , \new_[43987]_ , \new_[43990]_ , \new_[43993]_ ,
    \new_[43994]_ , \new_[43995]_ , \new_[43999]_ , \new_[44000]_ ,
    \new_[44003]_ , \new_[44006]_ , \new_[44007]_ , \new_[44008]_ ,
    \new_[44012]_ , \new_[44013]_ , \new_[44016]_ , \new_[44019]_ ,
    \new_[44020]_ , \new_[44021]_ , \new_[44025]_ , \new_[44026]_ ,
    \new_[44029]_ , \new_[44032]_ , \new_[44033]_ , \new_[44034]_ ,
    \new_[44038]_ , \new_[44039]_ , \new_[44042]_ , \new_[44045]_ ,
    \new_[44046]_ , \new_[44047]_ , \new_[44051]_ , \new_[44052]_ ,
    \new_[44055]_ , \new_[44058]_ , \new_[44059]_ , \new_[44060]_ ,
    \new_[44064]_ , \new_[44065]_ , \new_[44068]_ , \new_[44071]_ ,
    \new_[44072]_ , \new_[44073]_ , \new_[44077]_ , \new_[44078]_ ,
    \new_[44081]_ , \new_[44084]_ , \new_[44085]_ , \new_[44086]_ ,
    \new_[44090]_ , \new_[44091]_ , \new_[44094]_ , \new_[44097]_ ,
    \new_[44098]_ , \new_[44099]_ , \new_[44103]_ , \new_[44104]_ ,
    \new_[44107]_ , \new_[44110]_ , \new_[44111]_ , \new_[44112]_ ,
    \new_[44116]_ , \new_[44117]_ , \new_[44120]_ , \new_[44123]_ ,
    \new_[44124]_ , \new_[44125]_ , \new_[44129]_ , \new_[44130]_ ,
    \new_[44133]_ , \new_[44136]_ , \new_[44137]_ , \new_[44138]_ ,
    \new_[44142]_ , \new_[44143]_ , \new_[44146]_ , \new_[44149]_ ,
    \new_[44150]_ , \new_[44151]_ , \new_[44155]_ , \new_[44156]_ ,
    \new_[44159]_ , \new_[44162]_ , \new_[44163]_ , \new_[44164]_ ,
    \new_[44168]_ , \new_[44169]_ , \new_[44172]_ , \new_[44175]_ ,
    \new_[44176]_ , \new_[44177]_ , \new_[44181]_ , \new_[44182]_ ,
    \new_[44185]_ , \new_[44188]_ , \new_[44189]_ , \new_[44190]_ ,
    \new_[44194]_ , \new_[44195]_ , \new_[44198]_ , \new_[44201]_ ,
    \new_[44202]_ , \new_[44203]_ , \new_[44207]_ , \new_[44208]_ ,
    \new_[44211]_ , \new_[44214]_ , \new_[44215]_ , \new_[44216]_ ,
    \new_[44220]_ , \new_[44221]_ , \new_[44224]_ , \new_[44227]_ ,
    \new_[44228]_ , \new_[44229]_ , \new_[44233]_ , \new_[44234]_ ,
    \new_[44237]_ , \new_[44240]_ , \new_[44241]_ , \new_[44242]_ ,
    \new_[44246]_ , \new_[44247]_ , \new_[44250]_ , \new_[44253]_ ,
    \new_[44254]_ , \new_[44255]_ , \new_[44259]_ , \new_[44260]_ ,
    \new_[44263]_ , \new_[44266]_ , \new_[44267]_ , \new_[44268]_ ,
    \new_[44272]_ , \new_[44273]_ , \new_[44276]_ , \new_[44279]_ ,
    \new_[44280]_ , \new_[44281]_ , \new_[44285]_ , \new_[44286]_ ,
    \new_[44289]_ , \new_[44292]_ , \new_[44293]_ , \new_[44294]_ ,
    \new_[44298]_ , \new_[44299]_ , \new_[44302]_ , \new_[44305]_ ,
    \new_[44306]_ , \new_[44307]_ , \new_[44311]_ , \new_[44312]_ ,
    \new_[44315]_ , \new_[44318]_ , \new_[44319]_ , \new_[44320]_ ,
    \new_[44324]_ , \new_[44325]_ , \new_[44328]_ , \new_[44331]_ ,
    \new_[44332]_ , \new_[44333]_ , \new_[44337]_ , \new_[44338]_ ,
    \new_[44341]_ , \new_[44344]_ , \new_[44345]_ , \new_[44346]_ ,
    \new_[44350]_ , \new_[44351]_ , \new_[44354]_ , \new_[44357]_ ,
    \new_[44358]_ , \new_[44359]_ , \new_[44363]_ , \new_[44364]_ ,
    \new_[44367]_ , \new_[44370]_ , \new_[44371]_ , \new_[44372]_ ,
    \new_[44376]_ , \new_[44377]_ , \new_[44380]_ , \new_[44383]_ ,
    \new_[44384]_ , \new_[44385]_ , \new_[44389]_ , \new_[44390]_ ,
    \new_[44393]_ , \new_[44396]_ , \new_[44397]_ , \new_[44398]_ ,
    \new_[44402]_ , \new_[44403]_ , \new_[44406]_ , \new_[44409]_ ,
    \new_[44410]_ , \new_[44411]_ , \new_[44415]_ , \new_[44416]_ ,
    \new_[44419]_ , \new_[44422]_ , \new_[44423]_ , \new_[44424]_ ,
    \new_[44428]_ , \new_[44429]_ , \new_[44432]_ , \new_[44435]_ ,
    \new_[44436]_ , \new_[44437]_ , \new_[44441]_ , \new_[44442]_ ,
    \new_[44445]_ , \new_[44448]_ , \new_[44449]_ , \new_[44450]_ ,
    \new_[44454]_ , \new_[44455]_ , \new_[44458]_ , \new_[44461]_ ,
    \new_[44462]_ , \new_[44463]_ , \new_[44467]_ , \new_[44468]_ ,
    \new_[44471]_ , \new_[44474]_ , \new_[44475]_ , \new_[44476]_ ,
    \new_[44480]_ , \new_[44481]_ , \new_[44484]_ , \new_[44487]_ ,
    \new_[44488]_ , \new_[44489]_ , \new_[44493]_ , \new_[44494]_ ,
    \new_[44497]_ , \new_[44500]_ , \new_[44501]_ , \new_[44502]_ ,
    \new_[44506]_ , \new_[44507]_ , \new_[44510]_ , \new_[44513]_ ,
    \new_[44514]_ , \new_[44515]_ , \new_[44519]_ , \new_[44520]_ ,
    \new_[44523]_ , \new_[44526]_ , \new_[44527]_ , \new_[44528]_ ,
    \new_[44532]_ , \new_[44533]_ , \new_[44536]_ , \new_[44539]_ ,
    \new_[44540]_ , \new_[44541]_ , \new_[44545]_ , \new_[44546]_ ,
    \new_[44549]_ , \new_[44552]_ , \new_[44553]_ , \new_[44554]_ ,
    \new_[44558]_ , \new_[44559]_ , \new_[44562]_ , \new_[44565]_ ,
    \new_[44566]_ , \new_[44567]_ , \new_[44571]_ , \new_[44572]_ ,
    \new_[44575]_ , \new_[44578]_ , \new_[44579]_ , \new_[44580]_ ,
    \new_[44584]_ , \new_[44585]_ , \new_[44588]_ , \new_[44591]_ ,
    \new_[44592]_ , \new_[44593]_ , \new_[44597]_ , \new_[44598]_ ,
    \new_[44601]_ , \new_[44604]_ , \new_[44605]_ , \new_[44606]_ ,
    \new_[44610]_ , \new_[44611]_ , \new_[44614]_ , \new_[44617]_ ,
    \new_[44618]_ , \new_[44619]_ , \new_[44623]_ , \new_[44624]_ ,
    \new_[44627]_ , \new_[44630]_ , \new_[44631]_ , \new_[44632]_ ,
    \new_[44636]_ , \new_[44637]_ , \new_[44640]_ , \new_[44643]_ ,
    \new_[44644]_ , \new_[44645]_ , \new_[44649]_ , \new_[44650]_ ,
    \new_[44653]_ , \new_[44656]_ , \new_[44657]_ , \new_[44658]_ ,
    \new_[44662]_ , \new_[44663]_ , \new_[44666]_ , \new_[44669]_ ,
    \new_[44670]_ , \new_[44671]_ , \new_[44675]_ , \new_[44676]_ ,
    \new_[44679]_ , \new_[44682]_ , \new_[44683]_ , \new_[44684]_ ,
    \new_[44688]_ , \new_[44689]_ , \new_[44692]_ , \new_[44695]_ ,
    \new_[44696]_ , \new_[44697]_ , \new_[44701]_ , \new_[44702]_ ,
    \new_[44705]_ , \new_[44708]_ , \new_[44709]_ , \new_[44710]_ ,
    \new_[44714]_ , \new_[44715]_ , \new_[44718]_ , \new_[44721]_ ,
    \new_[44722]_ , \new_[44723]_ , \new_[44727]_ , \new_[44728]_ ,
    \new_[44731]_ , \new_[44734]_ , \new_[44735]_ , \new_[44736]_ ,
    \new_[44740]_ , \new_[44741]_ , \new_[44744]_ , \new_[44747]_ ,
    \new_[44748]_ , \new_[44749]_ , \new_[44753]_ , \new_[44754]_ ,
    \new_[44757]_ , \new_[44760]_ , \new_[44761]_ , \new_[44762]_ ,
    \new_[44766]_ , \new_[44767]_ , \new_[44770]_ , \new_[44773]_ ,
    \new_[44774]_ , \new_[44775]_ , \new_[44779]_ , \new_[44780]_ ,
    \new_[44783]_ , \new_[44786]_ , \new_[44787]_ , \new_[44788]_ ,
    \new_[44792]_ , \new_[44793]_ , \new_[44796]_ , \new_[44799]_ ,
    \new_[44800]_ , \new_[44801]_ , \new_[44805]_ , \new_[44806]_ ,
    \new_[44809]_ , \new_[44812]_ , \new_[44813]_ , \new_[44814]_ ,
    \new_[44818]_ , \new_[44819]_ , \new_[44822]_ , \new_[44825]_ ,
    \new_[44826]_ , \new_[44827]_ , \new_[44831]_ , \new_[44832]_ ,
    \new_[44835]_ , \new_[44838]_ , \new_[44839]_ , \new_[44840]_ ,
    \new_[44844]_ , \new_[44845]_ , \new_[44848]_ , \new_[44851]_ ,
    \new_[44852]_ , \new_[44853]_ , \new_[44857]_ , \new_[44858]_ ,
    \new_[44861]_ , \new_[44864]_ , \new_[44865]_ , \new_[44866]_ ,
    \new_[44870]_ , \new_[44871]_ , \new_[44874]_ , \new_[44877]_ ,
    \new_[44878]_ , \new_[44879]_ , \new_[44883]_ , \new_[44884]_ ,
    \new_[44887]_ , \new_[44890]_ , \new_[44891]_ , \new_[44892]_ ,
    \new_[44896]_ , \new_[44897]_ , \new_[44900]_ , \new_[44903]_ ,
    \new_[44904]_ , \new_[44905]_ , \new_[44909]_ , \new_[44910]_ ,
    \new_[44913]_ , \new_[44916]_ , \new_[44917]_ , \new_[44918]_ ,
    \new_[44922]_ , \new_[44923]_ , \new_[44926]_ , \new_[44929]_ ,
    \new_[44930]_ , \new_[44931]_ , \new_[44935]_ , \new_[44936]_ ,
    \new_[44939]_ , \new_[44942]_ , \new_[44943]_ , \new_[44944]_ ,
    \new_[44948]_ , \new_[44949]_ , \new_[44952]_ , \new_[44955]_ ,
    \new_[44956]_ , \new_[44957]_ , \new_[44961]_ , \new_[44962]_ ,
    \new_[44965]_ , \new_[44968]_ , \new_[44969]_ , \new_[44970]_ ,
    \new_[44974]_ , \new_[44975]_ , \new_[44978]_ , \new_[44981]_ ,
    \new_[44982]_ , \new_[44983]_ , \new_[44987]_ , \new_[44988]_ ,
    \new_[44991]_ , \new_[44994]_ , \new_[44995]_ , \new_[44996]_ ,
    \new_[45000]_ , \new_[45001]_ , \new_[45004]_ , \new_[45007]_ ,
    \new_[45008]_ , \new_[45009]_ , \new_[45013]_ , \new_[45014]_ ,
    \new_[45017]_ , \new_[45020]_ , \new_[45021]_ , \new_[45022]_ ,
    \new_[45026]_ , \new_[45027]_ , \new_[45030]_ , \new_[45033]_ ,
    \new_[45034]_ , \new_[45035]_ , \new_[45039]_ , \new_[45040]_ ,
    \new_[45043]_ , \new_[45046]_ , \new_[45047]_ , \new_[45048]_ ,
    \new_[45052]_ , \new_[45053]_ , \new_[45056]_ , \new_[45059]_ ,
    \new_[45060]_ , \new_[45061]_ , \new_[45065]_ , \new_[45066]_ ,
    \new_[45069]_ , \new_[45072]_ , \new_[45073]_ , \new_[45074]_ ,
    \new_[45078]_ , \new_[45079]_ , \new_[45082]_ , \new_[45085]_ ,
    \new_[45086]_ , \new_[45087]_ , \new_[45091]_ , \new_[45092]_ ,
    \new_[45095]_ , \new_[45098]_ , \new_[45099]_ , \new_[45100]_ ,
    \new_[45104]_ , \new_[45105]_ , \new_[45108]_ , \new_[45111]_ ,
    \new_[45112]_ , \new_[45113]_ , \new_[45117]_ , \new_[45118]_ ,
    \new_[45121]_ , \new_[45124]_ , \new_[45125]_ , \new_[45126]_ ,
    \new_[45130]_ , \new_[45131]_ , \new_[45134]_ , \new_[45137]_ ,
    \new_[45138]_ , \new_[45139]_ , \new_[45143]_ , \new_[45144]_ ,
    \new_[45147]_ , \new_[45150]_ , \new_[45151]_ , \new_[45152]_ ,
    \new_[45156]_ , \new_[45157]_ , \new_[45160]_ , \new_[45163]_ ,
    \new_[45164]_ , \new_[45165]_ , \new_[45169]_ , \new_[45170]_ ,
    \new_[45173]_ , \new_[45176]_ , \new_[45177]_ , \new_[45178]_ ,
    \new_[45182]_ , \new_[45183]_ , \new_[45186]_ , \new_[45189]_ ,
    \new_[45190]_ , \new_[45191]_ , \new_[45195]_ , \new_[45196]_ ,
    \new_[45199]_ , \new_[45202]_ , \new_[45203]_ , \new_[45204]_ ,
    \new_[45208]_ , \new_[45209]_ , \new_[45212]_ , \new_[45215]_ ,
    \new_[45216]_ , \new_[45217]_ , \new_[45221]_ , \new_[45222]_ ,
    \new_[45225]_ , \new_[45228]_ , \new_[45229]_ , \new_[45230]_ ,
    \new_[45234]_ , \new_[45235]_ , \new_[45238]_ , \new_[45241]_ ,
    \new_[45242]_ , \new_[45243]_ , \new_[45247]_ , \new_[45248]_ ,
    \new_[45251]_ , \new_[45254]_ , \new_[45255]_ , \new_[45256]_ ,
    \new_[45260]_ , \new_[45261]_ , \new_[45264]_ , \new_[45267]_ ,
    \new_[45268]_ , \new_[45269]_ , \new_[45273]_ , \new_[45274]_ ,
    \new_[45277]_ , \new_[45280]_ , \new_[45281]_ , \new_[45282]_ ,
    \new_[45286]_ , \new_[45287]_ , \new_[45290]_ , \new_[45293]_ ,
    \new_[45294]_ , \new_[45295]_ , \new_[45299]_ , \new_[45300]_ ,
    \new_[45303]_ , \new_[45306]_ , \new_[45307]_ , \new_[45308]_ ,
    \new_[45312]_ , \new_[45313]_ , \new_[45316]_ , \new_[45319]_ ,
    \new_[45320]_ , \new_[45321]_ , \new_[45325]_ , \new_[45326]_ ,
    \new_[45329]_ , \new_[45332]_ , \new_[45333]_ , \new_[45334]_ ,
    \new_[45338]_ , \new_[45339]_ , \new_[45342]_ , \new_[45345]_ ,
    \new_[45346]_ , \new_[45347]_ , \new_[45351]_ , \new_[45352]_ ,
    \new_[45355]_ , \new_[45358]_ , \new_[45359]_ , \new_[45360]_ ,
    \new_[45364]_ , \new_[45365]_ , \new_[45368]_ , \new_[45371]_ ,
    \new_[45372]_ , \new_[45373]_ , \new_[45377]_ , \new_[45378]_ ,
    \new_[45381]_ , \new_[45384]_ , \new_[45385]_ , \new_[45386]_ ,
    \new_[45390]_ , \new_[45391]_ , \new_[45394]_ , \new_[45397]_ ,
    \new_[45398]_ , \new_[45399]_ , \new_[45403]_ , \new_[45404]_ ,
    \new_[45407]_ , \new_[45410]_ , \new_[45411]_ , \new_[45412]_ ,
    \new_[45416]_ , \new_[45417]_ , \new_[45420]_ , \new_[45423]_ ,
    \new_[45424]_ , \new_[45425]_ , \new_[45429]_ , \new_[45430]_ ,
    \new_[45433]_ , \new_[45436]_ , \new_[45437]_ , \new_[45438]_ ,
    \new_[45442]_ , \new_[45443]_ , \new_[45446]_ , \new_[45449]_ ,
    \new_[45450]_ , \new_[45451]_ , \new_[45455]_ , \new_[45456]_ ,
    \new_[45459]_ , \new_[45462]_ , \new_[45463]_ , \new_[45464]_ ,
    \new_[45468]_ , \new_[45469]_ , \new_[45472]_ , \new_[45475]_ ,
    \new_[45476]_ , \new_[45477]_ , \new_[45481]_ , \new_[45482]_ ,
    \new_[45485]_ , \new_[45488]_ , \new_[45489]_ , \new_[45490]_ ,
    \new_[45494]_ , \new_[45495]_ , \new_[45498]_ , \new_[45501]_ ,
    \new_[45502]_ , \new_[45503]_ , \new_[45507]_ , \new_[45508]_ ,
    \new_[45511]_ , \new_[45514]_ , \new_[45515]_ , \new_[45516]_ ,
    \new_[45520]_ , \new_[45521]_ , \new_[45524]_ , \new_[45527]_ ,
    \new_[45528]_ , \new_[45529]_ , \new_[45533]_ , \new_[45534]_ ,
    \new_[45537]_ , \new_[45540]_ , \new_[45541]_ , \new_[45542]_ ,
    \new_[45546]_ , \new_[45547]_ , \new_[45550]_ , \new_[45553]_ ,
    \new_[45554]_ , \new_[45555]_ , \new_[45559]_ , \new_[45560]_ ,
    \new_[45563]_ , \new_[45566]_ , \new_[45567]_ , \new_[45568]_ ,
    \new_[45572]_ , \new_[45573]_ , \new_[45576]_ , \new_[45579]_ ,
    \new_[45580]_ , \new_[45581]_ , \new_[45585]_ , \new_[45586]_ ,
    \new_[45589]_ , \new_[45592]_ , \new_[45593]_ , \new_[45594]_ ,
    \new_[45598]_ , \new_[45599]_ , \new_[45602]_ , \new_[45605]_ ,
    \new_[45606]_ , \new_[45607]_ , \new_[45611]_ , \new_[45612]_ ,
    \new_[45615]_ , \new_[45618]_ , \new_[45619]_ , \new_[45620]_ ,
    \new_[45624]_ , \new_[45625]_ , \new_[45628]_ , \new_[45631]_ ,
    \new_[45632]_ , \new_[45633]_ , \new_[45637]_ , \new_[45638]_ ,
    \new_[45641]_ , \new_[45644]_ , \new_[45645]_ , \new_[45646]_ ,
    \new_[45650]_ , \new_[45651]_ , \new_[45654]_ , \new_[45657]_ ,
    \new_[45658]_ , \new_[45659]_ , \new_[45663]_ , \new_[45664]_ ,
    \new_[45667]_ , \new_[45670]_ , \new_[45671]_ , \new_[45672]_ ,
    \new_[45676]_ , \new_[45677]_ , \new_[45680]_ , \new_[45683]_ ,
    \new_[45684]_ , \new_[45685]_ , \new_[45689]_ , \new_[45690]_ ,
    \new_[45693]_ , \new_[45696]_ , \new_[45697]_ , \new_[45698]_ ,
    \new_[45702]_ , \new_[45703]_ , \new_[45706]_ , \new_[45709]_ ,
    \new_[45710]_ , \new_[45711]_ , \new_[45715]_ , \new_[45716]_ ,
    \new_[45719]_ , \new_[45722]_ , \new_[45723]_ , \new_[45724]_ ,
    \new_[45728]_ , \new_[45729]_ , \new_[45732]_ , \new_[45735]_ ,
    \new_[45736]_ , \new_[45737]_ , \new_[45741]_ , \new_[45742]_ ,
    \new_[45745]_ , \new_[45748]_ , \new_[45749]_ , \new_[45750]_ ,
    \new_[45754]_ , \new_[45755]_ , \new_[45758]_ , \new_[45761]_ ,
    \new_[45762]_ , \new_[45763]_ , \new_[45767]_ , \new_[45768]_ ,
    \new_[45771]_ , \new_[45774]_ , \new_[45775]_ , \new_[45776]_ ,
    \new_[45780]_ , \new_[45781]_ , \new_[45784]_ , \new_[45787]_ ,
    \new_[45788]_ , \new_[45789]_ , \new_[45793]_ , \new_[45794]_ ,
    \new_[45797]_ , \new_[45800]_ , \new_[45801]_ , \new_[45802]_ ,
    \new_[45806]_ , \new_[45807]_ , \new_[45810]_ , \new_[45813]_ ,
    \new_[45814]_ , \new_[45815]_ , \new_[45819]_ , \new_[45820]_ ,
    \new_[45823]_ , \new_[45826]_ , \new_[45827]_ , \new_[45828]_ ,
    \new_[45832]_ , \new_[45833]_ , \new_[45836]_ , \new_[45839]_ ,
    \new_[45840]_ , \new_[45841]_ , \new_[45845]_ , \new_[45846]_ ,
    \new_[45849]_ , \new_[45852]_ , \new_[45853]_ , \new_[45854]_ ,
    \new_[45858]_ , \new_[45859]_ , \new_[45862]_ , \new_[45865]_ ,
    \new_[45866]_ , \new_[45867]_ , \new_[45871]_ , \new_[45872]_ ,
    \new_[45875]_ , \new_[45878]_ , \new_[45879]_ , \new_[45880]_ ,
    \new_[45884]_ , \new_[45885]_ , \new_[45888]_ , \new_[45891]_ ,
    \new_[45892]_ , \new_[45893]_ , \new_[45897]_ , \new_[45898]_ ,
    \new_[45901]_ , \new_[45904]_ , \new_[45905]_ , \new_[45906]_ ,
    \new_[45910]_ , \new_[45911]_ , \new_[45914]_ , \new_[45917]_ ,
    \new_[45918]_ , \new_[45919]_ , \new_[45923]_ , \new_[45924]_ ,
    \new_[45927]_ , \new_[45930]_ , \new_[45931]_ , \new_[45932]_ ,
    \new_[45936]_ , \new_[45937]_ , \new_[45940]_ , \new_[45943]_ ,
    \new_[45944]_ , \new_[45945]_ , \new_[45949]_ , \new_[45950]_ ,
    \new_[45953]_ , \new_[45956]_ , \new_[45957]_ , \new_[45958]_ ,
    \new_[45962]_ , \new_[45963]_ , \new_[45966]_ , \new_[45969]_ ,
    \new_[45970]_ , \new_[45971]_ , \new_[45975]_ , \new_[45976]_ ,
    \new_[45979]_ , \new_[45982]_ , \new_[45983]_ , \new_[45984]_ ,
    \new_[45988]_ , \new_[45989]_ , \new_[45992]_ , \new_[45995]_ ,
    \new_[45996]_ , \new_[45997]_ , \new_[46001]_ , \new_[46002]_ ,
    \new_[46005]_ , \new_[46008]_ , \new_[46009]_ , \new_[46010]_ ,
    \new_[46014]_ , \new_[46015]_ , \new_[46018]_ , \new_[46021]_ ,
    \new_[46022]_ , \new_[46023]_ , \new_[46027]_ , \new_[46028]_ ,
    \new_[46031]_ , \new_[46034]_ , \new_[46035]_ , \new_[46036]_ ,
    \new_[46040]_ , \new_[46041]_ , \new_[46044]_ , \new_[46047]_ ,
    \new_[46048]_ , \new_[46049]_ , \new_[46053]_ , \new_[46054]_ ,
    \new_[46057]_ , \new_[46060]_ , \new_[46061]_ , \new_[46062]_ ,
    \new_[46066]_ , \new_[46067]_ , \new_[46070]_ , \new_[46073]_ ,
    \new_[46074]_ , \new_[46075]_ , \new_[46079]_ , \new_[46080]_ ,
    \new_[46083]_ , \new_[46086]_ , \new_[46087]_ , \new_[46088]_ ,
    \new_[46092]_ , \new_[46093]_ , \new_[46096]_ , \new_[46099]_ ,
    \new_[46100]_ , \new_[46101]_ , \new_[46105]_ , \new_[46106]_ ,
    \new_[46109]_ , \new_[46112]_ , \new_[46113]_ , \new_[46114]_ ,
    \new_[46118]_ , \new_[46119]_ , \new_[46122]_ , \new_[46125]_ ,
    \new_[46126]_ , \new_[46127]_ , \new_[46131]_ , \new_[46132]_ ,
    \new_[46135]_ , \new_[46138]_ , \new_[46139]_ , \new_[46140]_ ,
    \new_[46144]_ , \new_[46145]_ , \new_[46148]_ , \new_[46151]_ ,
    \new_[46152]_ , \new_[46153]_ , \new_[46157]_ , \new_[46158]_ ,
    \new_[46161]_ , \new_[46164]_ , \new_[46165]_ , \new_[46166]_ ,
    \new_[46170]_ , \new_[46171]_ , \new_[46174]_ , \new_[46177]_ ,
    \new_[46178]_ , \new_[46179]_ , \new_[46183]_ , \new_[46184]_ ,
    \new_[46187]_ , \new_[46190]_ , \new_[46191]_ , \new_[46192]_ ,
    \new_[46196]_ , \new_[46197]_ , \new_[46200]_ , \new_[46203]_ ,
    \new_[46204]_ , \new_[46205]_ , \new_[46209]_ , \new_[46210]_ ,
    \new_[46213]_ , \new_[46216]_ , \new_[46217]_ , \new_[46218]_ ,
    \new_[46222]_ , \new_[46223]_ , \new_[46226]_ , \new_[46229]_ ,
    \new_[46230]_ , \new_[46231]_ , \new_[46235]_ , \new_[46236]_ ,
    \new_[46239]_ , \new_[46242]_ , \new_[46243]_ , \new_[46244]_ ,
    \new_[46248]_ , \new_[46249]_ , \new_[46252]_ , \new_[46255]_ ,
    \new_[46256]_ , \new_[46257]_ , \new_[46261]_ , \new_[46262]_ ,
    \new_[46265]_ , \new_[46268]_ , \new_[46269]_ , \new_[46270]_ ,
    \new_[46274]_ , \new_[46275]_ , \new_[46278]_ , \new_[46281]_ ,
    \new_[46282]_ , \new_[46283]_ , \new_[46287]_ , \new_[46288]_ ,
    \new_[46291]_ , \new_[46294]_ , \new_[46295]_ , \new_[46296]_ ,
    \new_[46300]_ , \new_[46301]_ , \new_[46304]_ , \new_[46307]_ ,
    \new_[46308]_ , \new_[46309]_ , \new_[46313]_ , \new_[46314]_ ,
    \new_[46317]_ , \new_[46320]_ , \new_[46321]_ , \new_[46322]_ ,
    \new_[46326]_ , \new_[46327]_ , \new_[46330]_ , \new_[46333]_ ,
    \new_[46334]_ , \new_[46335]_ , \new_[46339]_ , \new_[46340]_ ,
    \new_[46343]_ , \new_[46346]_ , \new_[46347]_ , \new_[46348]_ ,
    \new_[46352]_ , \new_[46353]_ , \new_[46356]_ , \new_[46359]_ ,
    \new_[46360]_ , \new_[46361]_ , \new_[46365]_ , \new_[46366]_ ,
    \new_[46369]_ , \new_[46372]_ , \new_[46373]_ , \new_[46374]_ ,
    \new_[46378]_ , \new_[46379]_ , \new_[46382]_ , \new_[46385]_ ,
    \new_[46386]_ , \new_[46387]_ , \new_[46391]_ , \new_[46392]_ ,
    \new_[46395]_ , \new_[46398]_ , \new_[46399]_ , \new_[46400]_ ,
    \new_[46404]_ , \new_[46405]_ , \new_[46408]_ , \new_[46411]_ ,
    \new_[46412]_ , \new_[46413]_ , \new_[46417]_ , \new_[46418]_ ,
    \new_[46421]_ , \new_[46424]_ , \new_[46425]_ , \new_[46426]_ ,
    \new_[46430]_ , \new_[46431]_ , \new_[46434]_ , \new_[46437]_ ,
    \new_[46438]_ , \new_[46439]_ , \new_[46443]_ , \new_[46444]_ ,
    \new_[46447]_ , \new_[46450]_ , \new_[46451]_ , \new_[46452]_ ,
    \new_[46456]_ , \new_[46457]_ , \new_[46460]_ , \new_[46463]_ ,
    \new_[46464]_ , \new_[46465]_ , \new_[46469]_ , \new_[46470]_ ,
    \new_[46473]_ , \new_[46476]_ , \new_[46477]_ , \new_[46478]_ ,
    \new_[46482]_ , \new_[46483]_ , \new_[46486]_ , \new_[46489]_ ,
    \new_[46490]_ , \new_[46491]_ , \new_[46495]_ , \new_[46496]_ ,
    \new_[46499]_ , \new_[46502]_ , \new_[46503]_ , \new_[46504]_ ,
    \new_[46508]_ , \new_[46509]_ , \new_[46512]_ , \new_[46515]_ ,
    \new_[46516]_ , \new_[46517]_ , \new_[46521]_ , \new_[46522]_ ,
    \new_[46525]_ , \new_[46528]_ , \new_[46529]_ , \new_[46530]_ ,
    \new_[46534]_ , \new_[46535]_ , \new_[46538]_ , \new_[46541]_ ,
    \new_[46542]_ , \new_[46543]_ , \new_[46547]_ , \new_[46548]_ ,
    \new_[46551]_ , \new_[46554]_ , \new_[46555]_ , \new_[46556]_ ,
    \new_[46560]_ , \new_[46561]_ , \new_[46564]_ , \new_[46567]_ ,
    \new_[46568]_ , \new_[46569]_ , \new_[46573]_ , \new_[46574]_ ,
    \new_[46577]_ , \new_[46580]_ , \new_[46581]_ , \new_[46582]_ ,
    \new_[46586]_ , \new_[46587]_ , \new_[46590]_ , \new_[46593]_ ,
    \new_[46594]_ , \new_[46595]_ , \new_[46599]_ , \new_[46600]_ ,
    \new_[46603]_ , \new_[46606]_ , \new_[46607]_ , \new_[46608]_ ,
    \new_[46612]_ , \new_[46613]_ , \new_[46616]_ , \new_[46619]_ ,
    \new_[46620]_ , \new_[46621]_ , \new_[46625]_ , \new_[46626]_ ,
    \new_[46629]_ , \new_[46632]_ , \new_[46633]_ , \new_[46634]_ ,
    \new_[46638]_ , \new_[46639]_ , \new_[46642]_ , \new_[46645]_ ,
    \new_[46646]_ , \new_[46647]_ , \new_[46651]_ , \new_[46652]_ ,
    \new_[46655]_ , \new_[46658]_ , \new_[46659]_ , \new_[46660]_ ,
    \new_[46664]_ , \new_[46665]_ , \new_[46668]_ , \new_[46671]_ ,
    \new_[46672]_ , \new_[46673]_ , \new_[46677]_ , \new_[46678]_ ,
    \new_[46681]_ , \new_[46684]_ , \new_[46685]_ , \new_[46686]_ ,
    \new_[46690]_ , \new_[46691]_ , \new_[46694]_ , \new_[46697]_ ,
    \new_[46698]_ , \new_[46699]_ , \new_[46703]_ , \new_[46704]_ ,
    \new_[46707]_ , \new_[46710]_ , \new_[46711]_ , \new_[46712]_ ,
    \new_[46716]_ , \new_[46717]_ , \new_[46720]_ , \new_[46723]_ ,
    \new_[46724]_ , \new_[46725]_ , \new_[46729]_ , \new_[46730]_ ,
    \new_[46733]_ , \new_[46736]_ , \new_[46737]_ , \new_[46738]_ ,
    \new_[46742]_ , \new_[46743]_ , \new_[46746]_ , \new_[46749]_ ,
    \new_[46750]_ , \new_[46751]_ , \new_[46755]_ , \new_[46756]_ ,
    \new_[46759]_ , \new_[46762]_ , \new_[46763]_ , \new_[46764]_ ,
    \new_[46768]_ , \new_[46769]_ , \new_[46772]_ , \new_[46775]_ ,
    \new_[46776]_ , \new_[46777]_ , \new_[46781]_ , \new_[46782]_ ,
    \new_[46785]_ , \new_[46788]_ , \new_[46789]_ , \new_[46790]_ ,
    \new_[46794]_ , \new_[46795]_ , \new_[46798]_ , \new_[46801]_ ,
    \new_[46802]_ , \new_[46803]_ , \new_[46807]_ , \new_[46808]_ ,
    \new_[46811]_ , \new_[46814]_ , \new_[46815]_ , \new_[46816]_ ,
    \new_[46820]_ , \new_[46821]_ , \new_[46824]_ , \new_[46827]_ ,
    \new_[46828]_ , \new_[46829]_ , \new_[46833]_ , \new_[46834]_ ,
    \new_[46837]_ , \new_[46840]_ , \new_[46841]_ , \new_[46842]_ ,
    \new_[46846]_ , \new_[46847]_ , \new_[46850]_ , \new_[46853]_ ,
    \new_[46854]_ , \new_[46855]_ , \new_[46859]_ , \new_[46860]_ ,
    \new_[46863]_ , \new_[46866]_ , \new_[46867]_ , \new_[46868]_ ,
    \new_[46872]_ , \new_[46873]_ , \new_[46876]_ , \new_[46879]_ ,
    \new_[46880]_ , \new_[46881]_ , \new_[46885]_ , \new_[46886]_ ,
    \new_[46889]_ , \new_[46892]_ , \new_[46893]_ , \new_[46894]_ ,
    \new_[46898]_ , \new_[46899]_ , \new_[46902]_ , \new_[46905]_ ,
    \new_[46906]_ , \new_[46907]_ , \new_[46911]_ , \new_[46912]_ ,
    \new_[46915]_ , \new_[46918]_ , \new_[46919]_ , \new_[46920]_ ,
    \new_[46924]_ , \new_[46925]_ , \new_[46928]_ , \new_[46931]_ ,
    \new_[46932]_ , \new_[46933]_ , \new_[46937]_ , \new_[46938]_ ,
    \new_[46941]_ , \new_[46944]_ , \new_[46945]_ , \new_[46946]_ ,
    \new_[46950]_ , \new_[46951]_ , \new_[46954]_ , \new_[46957]_ ,
    \new_[46958]_ , \new_[46959]_ , \new_[46963]_ , \new_[46964]_ ,
    \new_[46967]_ , \new_[46970]_ , \new_[46971]_ , \new_[46972]_ ,
    \new_[46976]_ , \new_[46977]_ , \new_[46980]_ , \new_[46983]_ ,
    \new_[46984]_ , \new_[46985]_ , \new_[46989]_ , \new_[46990]_ ,
    \new_[46993]_ , \new_[46996]_ , \new_[46997]_ , \new_[46998]_ ,
    \new_[47002]_ , \new_[47003]_ , \new_[47006]_ , \new_[47009]_ ,
    \new_[47010]_ , \new_[47011]_ , \new_[47015]_ , \new_[47016]_ ,
    \new_[47019]_ , \new_[47022]_ , \new_[47023]_ , \new_[47024]_ ,
    \new_[47028]_ , \new_[47029]_ , \new_[47032]_ , \new_[47035]_ ,
    \new_[47036]_ , \new_[47037]_ , \new_[47041]_ , \new_[47042]_ ,
    \new_[47045]_ , \new_[47048]_ , \new_[47049]_ , \new_[47050]_ ,
    \new_[47054]_ , \new_[47055]_ , \new_[47058]_ , \new_[47061]_ ,
    \new_[47062]_ , \new_[47063]_ , \new_[47067]_ , \new_[47068]_ ,
    \new_[47071]_ , \new_[47074]_ , \new_[47075]_ , \new_[47076]_ ,
    \new_[47080]_ , \new_[47081]_ , \new_[47084]_ , \new_[47087]_ ,
    \new_[47088]_ , \new_[47089]_ , \new_[47093]_ , \new_[47094]_ ,
    \new_[47097]_ , \new_[47100]_ , \new_[47101]_ , \new_[47102]_ ,
    \new_[47106]_ , \new_[47107]_ , \new_[47110]_ , \new_[47113]_ ,
    \new_[47114]_ , \new_[47115]_ , \new_[47119]_ , \new_[47120]_ ,
    \new_[47123]_ , \new_[47126]_ , \new_[47127]_ , \new_[47128]_ ,
    \new_[47132]_ , \new_[47133]_ , \new_[47136]_ , \new_[47139]_ ,
    \new_[47140]_ , \new_[47141]_ , \new_[47145]_ , \new_[47146]_ ,
    \new_[47149]_ , \new_[47152]_ , \new_[47153]_ , \new_[47154]_ ,
    \new_[47158]_ , \new_[47159]_ , \new_[47162]_ , \new_[47165]_ ,
    \new_[47166]_ , \new_[47167]_ , \new_[47171]_ , \new_[47172]_ ,
    \new_[47175]_ , \new_[47178]_ , \new_[47179]_ , \new_[47180]_ ,
    \new_[47184]_ , \new_[47185]_ , \new_[47188]_ , \new_[47191]_ ,
    \new_[47192]_ , \new_[47193]_ , \new_[47197]_ , \new_[47198]_ ,
    \new_[47201]_ , \new_[47204]_ , \new_[47205]_ , \new_[47206]_ ,
    \new_[47210]_ , \new_[47211]_ , \new_[47214]_ , \new_[47217]_ ,
    \new_[47218]_ , \new_[47219]_ , \new_[47223]_ , \new_[47224]_ ,
    \new_[47227]_ , \new_[47230]_ , \new_[47231]_ , \new_[47232]_ ,
    \new_[47236]_ , \new_[47237]_ , \new_[47240]_ , \new_[47243]_ ,
    \new_[47244]_ , \new_[47245]_ , \new_[47249]_ , \new_[47250]_ ,
    \new_[47253]_ , \new_[47256]_ , \new_[47257]_ , \new_[47258]_ ,
    \new_[47262]_ , \new_[47263]_ , \new_[47266]_ , \new_[47269]_ ,
    \new_[47270]_ , \new_[47271]_ , \new_[47275]_ , \new_[47276]_ ,
    \new_[47279]_ , \new_[47282]_ , \new_[47283]_ , \new_[47284]_ ,
    \new_[47288]_ , \new_[47289]_ , \new_[47292]_ , \new_[47295]_ ,
    \new_[47296]_ , \new_[47297]_ , \new_[47301]_ , \new_[47302]_ ,
    \new_[47305]_ , \new_[47308]_ , \new_[47309]_ , \new_[47310]_ ,
    \new_[47314]_ , \new_[47315]_ , \new_[47318]_ , \new_[47321]_ ,
    \new_[47322]_ , \new_[47323]_ , \new_[47327]_ , \new_[47328]_ ,
    \new_[47331]_ , \new_[47334]_ , \new_[47335]_ , \new_[47336]_ ,
    \new_[47340]_ , \new_[47341]_ , \new_[47344]_ , \new_[47347]_ ,
    \new_[47348]_ , \new_[47349]_ , \new_[47353]_ , \new_[47354]_ ,
    \new_[47357]_ , \new_[47360]_ , \new_[47361]_ , \new_[47362]_ ,
    \new_[47366]_ , \new_[47367]_ , \new_[47370]_ , \new_[47373]_ ,
    \new_[47374]_ , \new_[47375]_ , \new_[47379]_ , \new_[47380]_ ,
    \new_[47383]_ , \new_[47386]_ , \new_[47387]_ , \new_[47388]_ ,
    \new_[47392]_ , \new_[47393]_ , \new_[47396]_ , \new_[47399]_ ,
    \new_[47400]_ , \new_[47401]_ , \new_[47405]_ , \new_[47406]_ ,
    \new_[47409]_ , \new_[47412]_ , \new_[47413]_ , \new_[47414]_ ,
    \new_[47418]_ , \new_[47419]_ , \new_[47422]_ , \new_[47425]_ ,
    \new_[47426]_ , \new_[47427]_ , \new_[47431]_ , \new_[47432]_ ,
    \new_[47435]_ , \new_[47438]_ , \new_[47439]_ , \new_[47440]_ ,
    \new_[47444]_ , \new_[47445]_ , \new_[47448]_ , \new_[47451]_ ,
    \new_[47452]_ , \new_[47453]_ , \new_[47457]_ , \new_[47458]_ ,
    \new_[47461]_ , \new_[47464]_ , \new_[47465]_ , \new_[47466]_ ,
    \new_[47470]_ , \new_[47471]_ , \new_[47474]_ , \new_[47477]_ ,
    \new_[47478]_ , \new_[47479]_ , \new_[47483]_ , \new_[47484]_ ,
    \new_[47487]_ , \new_[47490]_ , \new_[47491]_ , \new_[47492]_ ,
    \new_[47496]_ , \new_[47497]_ , \new_[47500]_ , \new_[47503]_ ,
    \new_[47504]_ , \new_[47505]_ , \new_[47509]_ , \new_[47510]_ ,
    \new_[47513]_ , \new_[47516]_ , \new_[47517]_ , \new_[47518]_ ,
    \new_[47522]_ , \new_[47523]_ , \new_[47526]_ , \new_[47529]_ ,
    \new_[47530]_ , \new_[47531]_ , \new_[47535]_ , \new_[47536]_ ,
    \new_[47539]_ , \new_[47542]_ , \new_[47543]_ , \new_[47544]_ ,
    \new_[47548]_ , \new_[47549]_ , \new_[47552]_ , \new_[47555]_ ,
    \new_[47556]_ , \new_[47557]_ , \new_[47561]_ , \new_[47562]_ ,
    \new_[47565]_ , \new_[47568]_ , \new_[47569]_ , \new_[47570]_ ,
    \new_[47574]_ , \new_[47575]_ , \new_[47578]_ , \new_[47581]_ ,
    \new_[47582]_ , \new_[47583]_ , \new_[47587]_ , \new_[47588]_ ,
    \new_[47591]_ , \new_[47594]_ , \new_[47595]_ , \new_[47596]_ ,
    \new_[47600]_ , \new_[47601]_ , \new_[47604]_ , \new_[47607]_ ,
    \new_[47608]_ , \new_[47609]_ , \new_[47613]_ , \new_[47614]_ ,
    \new_[47617]_ , \new_[47620]_ , \new_[47621]_ , \new_[47622]_ ,
    \new_[47626]_ , \new_[47627]_ , \new_[47630]_ , \new_[47633]_ ,
    \new_[47634]_ , \new_[47635]_ , \new_[47639]_ , \new_[47640]_ ,
    \new_[47643]_ , \new_[47646]_ , \new_[47647]_ , \new_[47648]_ ,
    \new_[47652]_ , \new_[47653]_ , \new_[47656]_ , \new_[47659]_ ,
    \new_[47660]_ , \new_[47661]_ , \new_[47664]_ , \new_[47667]_ ,
    \new_[47668]_ , \new_[47671]_ , \new_[47674]_ , \new_[47675]_ ,
    \new_[47676]_ , \new_[47680]_ , \new_[47681]_ , \new_[47684]_ ,
    \new_[47687]_ , \new_[47688]_ , \new_[47689]_ , \new_[47692]_ ,
    \new_[47695]_ , \new_[47696]_ , \new_[47699]_ , \new_[47702]_ ,
    \new_[47703]_ , \new_[47704]_ , \new_[47708]_ , \new_[47709]_ ,
    \new_[47712]_ , \new_[47715]_ , \new_[47716]_ , \new_[47717]_ ,
    \new_[47720]_ , \new_[47723]_ , \new_[47724]_ , \new_[47727]_ ,
    \new_[47730]_ , \new_[47731]_ , \new_[47732]_ , \new_[47736]_ ,
    \new_[47737]_ , \new_[47740]_ , \new_[47743]_ , \new_[47744]_ ,
    \new_[47745]_ , \new_[47748]_ , \new_[47751]_ , \new_[47752]_ ,
    \new_[47755]_ , \new_[47758]_ , \new_[47759]_ , \new_[47760]_ ,
    \new_[47764]_ , \new_[47765]_ , \new_[47768]_ , \new_[47771]_ ,
    \new_[47772]_ , \new_[47773]_ , \new_[47776]_ , \new_[47779]_ ,
    \new_[47780]_ , \new_[47783]_ , \new_[47786]_ , \new_[47787]_ ,
    \new_[47788]_ , \new_[47792]_ , \new_[47793]_ , \new_[47796]_ ,
    \new_[47799]_ , \new_[47800]_ , \new_[47801]_ , \new_[47804]_ ,
    \new_[47807]_ , \new_[47808]_ , \new_[47811]_ , \new_[47814]_ ,
    \new_[47815]_ , \new_[47816]_ , \new_[47820]_ , \new_[47821]_ ,
    \new_[47824]_ , \new_[47827]_ , \new_[47828]_ , \new_[47829]_ ,
    \new_[47832]_ , \new_[47835]_ , \new_[47836]_ , \new_[47839]_ ,
    \new_[47842]_ , \new_[47843]_ , \new_[47844]_ , \new_[47848]_ ,
    \new_[47849]_ , \new_[47852]_ , \new_[47855]_ , \new_[47856]_ ,
    \new_[47857]_ , \new_[47860]_ , \new_[47863]_ , \new_[47864]_ ,
    \new_[47867]_ , \new_[47870]_ , \new_[47871]_ , \new_[47872]_ ,
    \new_[47876]_ , \new_[47877]_ , \new_[47880]_ , \new_[47883]_ ,
    \new_[47884]_ , \new_[47885]_ , \new_[47888]_ , \new_[47891]_ ,
    \new_[47892]_ , \new_[47895]_ , \new_[47898]_ , \new_[47899]_ ,
    \new_[47900]_ , \new_[47904]_ , \new_[47905]_ , \new_[47908]_ ,
    \new_[47911]_ , \new_[47912]_ , \new_[47913]_ , \new_[47916]_ ,
    \new_[47919]_ , \new_[47920]_ , \new_[47923]_ , \new_[47926]_ ,
    \new_[47927]_ , \new_[47928]_ , \new_[47932]_ , \new_[47933]_ ,
    \new_[47936]_ , \new_[47939]_ , \new_[47940]_ , \new_[47941]_ ,
    \new_[47944]_ , \new_[47947]_ , \new_[47948]_ , \new_[47951]_ ,
    \new_[47954]_ , \new_[47955]_ , \new_[47956]_ , \new_[47960]_ ,
    \new_[47961]_ , \new_[47964]_ , \new_[47967]_ , \new_[47968]_ ,
    \new_[47969]_ , \new_[47972]_ , \new_[47975]_ , \new_[47976]_ ,
    \new_[47979]_ , \new_[47982]_ , \new_[47983]_ , \new_[47984]_ ,
    \new_[47988]_ , \new_[47989]_ , \new_[47992]_ , \new_[47995]_ ,
    \new_[47996]_ , \new_[47997]_ , \new_[48000]_ , \new_[48003]_ ,
    \new_[48004]_ , \new_[48007]_ , \new_[48010]_ , \new_[48011]_ ,
    \new_[48012]_ , \new_[48016]_ , \new_[48017]_ , \new_[48020]_ ,
    \new_[48023]_ , \new_[48024]_ , \new_[48025]_ , \new_[48028]_ ,
    \new_[48031]_ , \new_[48032]_ , \new_[48035]_ , \new_[48038]_ ,
    \new_[48039]_ , \new_[48040]_ , \new_[48044]_ , \new_[48045]_ ,
    \new_[48048]_ , \new_[48051]_ , \new_[48052]_ , \new_[48053]_ ,
    \new_[48056]_ , \new_[48059]_ , \new_[48060]_ , \new_[48063]_ ,
    \new_[48066]_ , \new_[48067]_ , \new_[48068]_ , \new_[48072]_ ,
    \new_[48073]_ , \new_[48076]_ , \new_[48079]_ , \new_[48080]_ ,
    \new_[48081]_ , \new_[48084]_ , \new_[48087]_ , \new_[48088]_ ,
    \new_[48091]_ , \new_[48094]_ , \new_[48095]_ , \new_[48096]_ ,
    \new_[48100]_ , \new_[48101]_ , \new_[48104]_ , \new_[48107]_ ,
    \new_[48108]_ , \new_[48109]_ , \new_[48112]_ , \new_[48115]_ ,
    \new_[48116]_ , \new_[48119]_ , \new_[48122]_ , \new_[48123]_ ,
    \new_[48124]_ , \new_[48128]_ , \new_[48129]_ , \new_[48132]_ ,
    \new_[48135]_ , \new_[48136]_ , \new_[48137]_ , \new_[48140]_ ,
    \new_[48143]_ , \new_[48144]_ , \new_[48147]_ , \new_[48150]_ ,
    \new_[48151]_ , \new_[48152]_ , \new_[48156]_ , \new_[48157]_ ,
    \new_[48160]_ , \new_[48163]_ , \new_[48164]_ , \new_[48165]_ ,
    \new_[48168]_ , \new_[48171]_ , \new_[48172]_ , \new_[48175]_ ,
    \new_[48178]_ , \new_[48179]_ , \new_[48180]_ , \new_[48184]_ ,
    \new_[48185]_ , \new_[48188]_ , \new_[48191]_ , \new_[48192]_ ,
    \new_[48193]_ , \new_[48196]_ , \new_[48199]_ , \new_[48200]_ ,
    \new_[48203]_ , \new_[48206]_ , \new_[48207]_ , \new_[48208]_ ,
    \new_[48212]_ , \new_[48213]_ , \new_[48216]_ , \new_[48219]_ ,
    \new_[48220]_ , \new_[48221]_ , \new_[48224]_ , \new_[48227]_ ,
    \new_[48228]_ , \new_[48231]_ , \new_[48234]_ , \new_[48235]_ ,
    \new_[48236]_ , \new_[48240]_ , \new_[48241]_ , \new_[48244]_ ,
    \new_[48247]_ , \new_[48248]_ , \new_[48249]_ , \new_[48252]_ ,
    \new_[48255]_ , \new_[48256]_ , \new_[48259]_ , \new_[48262]_ ,
    \new_[48263]_ , \new_[48264]_ , \new_[48268]_ , \new_[48269]_ ,
    \new_[48272]_ , \new_[48275]_ , \new_[48276]_ , \new_[48277]_ ,
    \new_[48280]_ , \new_[48283]_ , \new_[48284]_ , \new_[48287]_ ,
    \new_[48290]_ , \new_[48291]_ , \new_[48292]_ , \new_[48296]_ ,
    \new_[48297]_ , \new_[48300]_ , \new_[48303]_ , \new_[48304]_ ,
    \new_[48305]_ , \new_[48308]_ , \new_[48311]_ , \new_[48312]_ ,
    \new_[48315]_ , \new_[48318]_ , \new_[48319]_ , \new_[48320]_ ,
    \new_[48324]_ , \new_[48325]_ , \new_[48328]_ , \new_[48331]_ ,
    \new_[48332]_ , \new_[48333]_ , \new_[48336]_ , \new_[48339]_ ,
    \new_[48340]_ , \new_[48343]_ , \new_[48346]_ , \new_[48347]_ ,
    \new_[48348]_ , \new_[48352]_ , \new_[48353]_ , \new_[48356]_ ,
    \new_[48359]_ , \new_[48360]_ , \new_[48361]_ , \new_[48364]_ ,
    \new_[48367]_ , \new_[48368]_ , \new_[48371]_ , \new_[48374]_ ,
    \new_[48375]_ , \new_[48376]_ , \new_[48380]_ , \new_[48381]_ ,
    \new_[48384]_ , \new_[48387]_ , \new_[48388]_ , \new_[48389]_ ,
    \new_[48392]_ , \new_[48395]_ , \new_[48396]_ , \new_[48399]_ ,
    \new_[48402]_ , \new_[48403]_ , \new_[48404]_ , \new_[48408]_ ,
    \new_[48409]_ , \new_[48412]_ , \new_[48415]_ , \new_[48416]_ ,
    \new_[48417]_ , \new_[48420]_ , \new_[48423]_ , \new_[48424]_ ,
    \new_[48427]_ , \new_[48430]_ , \new_[48431]_ , \new_[48432]_ ,
    \new_[48436]_ , \new_[48437]_ , \new_[48440]_ , \new_[48443]_ ,
    \new_[48444]_ , \new_[48445]_ , \new_[48448]_ , \new_[48451]_ ,
    \new_[48452]_ , \new_[48455]_ , \new_[48458]_ , \new_[48459]_ ,
    \new_[48460]_ , \new_[48464]_ , \new_[48465]_ , \new_[48468]_ ,
    \new_[48471]_ , \new_[48472]_ , \new_[48473]_ , \new_[48476]_ ,
    \new_[48479]_ , \new_[48480]_ , \new_[48483]_ , \new_[48486]_ ,
    \new_[48487]_ , \new_[48488]_ , \new_[48492]_ , \new_[48493]_ ,
    \new_[48496]_ , \new_[48499]_ , \new_[48500]_ , \new_[48501]_ ,
    \new_[48504]_ , \new_[48507]_ , \new_[48508]_ , \new_[48511]_ ,
    \new_[48514]_ , \new_[48515]_ , \new_[48516]_ , \new_[48520]_ ,
    \new_[48521]_ , \new_[48524]_ , \new_[48527]_ , \new_[48528]_ ,
    \new_[48529]_ , \new_[48532]_ , \new_[48535]_ , \new_[48536]_ ,
    \new_[48539]_ , \new_[48542]_ , \new_[48543]_ , \new_[48544]_ ,
    \new_[48548]_ , \new_[48549]_ , \new_[48552]_ , \new_[48555]_ ,
    \new_[48556]_ , \new_[48557]_ , \new_[48560]_ , \new_[48563]_ ,
    \new_[48564]_ , \new_[48567]_ , \new_[48570]_ , \new_[48571]_ ,
    \new_[48572]_ , \new_[48576]_ , \new_[48577]_ , \new_[48580]_ ,
    \new_[48583]_ , \new_[48584]_ , \new_[48585]_ , \new_[48588]_ ,
    \new_[48591]_ , \new_[48592]_ , \new_[48595]_ , \new_[48598]_ ,
    \new_[48599]_ , \new_[48600]_ , \new_[48604]_ , \new_[48605]_ ,
    \new_[48608]_ , \new_[48611]_ , \new_[48612]_ , \new_[48613]_ ,
    \new_[48616]_ , \new_[48619]_ , \new_[48620]_ , \new_[48623]_ ,
    \new_[48626]_ , \new_[48627]_ , \new_[48628]_ , \new_[48632]_ ,
    \new_[48633]_ , \new_[48636]_ , \new_[48639]_ , \new_[48640]_ ,
    \new_[48641]_ , \new_[48644]_ , \new_[48647]_ , \new_[48648]_ ,
    \new_[48651]_ , \new_[48654]_ , \new_[48655]_ , \new_[48656]_ ,
    \new_[48660]_ , \new_[48661]_ , \new_[48664]_ , \new_[48667]_ ,
    \new_[48668]_ , \new_[48669]_ , \new_[48672]_ , \new_[48675]_ ,
    \new_[48676]_ , \new_[48679]_ , \new_[48682]_ , \new_[48683]_ ,
    \new_[48684]_ , \new_[48688]_ , \new_[48689]_ , \new_[48692]_ ,
    \new_[48695]_ , \new_[48696]_ , \new_[48697]_ , \new_[48700]_ ,
    \new_[48703]_ , \new_[48704]_ , \new_[48707]_ , \new_[48710]_ ,
    \new_[48711]_ , \new_[48712]_ , \new_[48716]_ , \new_[48717]_ ,
    \new_[48720]_ , \new_[48723]_ , \new_[48724]_ , \new_[48725]_ ,
    \new_[48728]_ , \new_[48731]_ , \new_[48732]_ , \new_[48735]_ ,
    \new_[48738]_ , \new_[48739]_ , \new_[48740]_ , \new_[48744]_ ,
    \new_[48745]_ , \new_[48748]_ , \new_[48751]_ , \new_[48752]_ ,
    \new_[48753]_ , \new_[48756]_ , \new_[48759]_ , \new_[48760]_ ,
    \new_[48763]_ , \new_[48766]_ , \new_[48767]_ , \new_[48768]_ ,
    \new_[48772]_ , \new_[48773]_ , \new_[48776]_ , \new_[48779]_ ,
    \new_[48780]_ , \new_[48781]_ , \new_[48784]_ , \new_[48787]_ ,
    \new_[48788]_ , \new_[48791]_ , \new_[48794]_ , \new_[48795]_ ,
    \new_[48796]_ , \new_[48800]_ , \new_[48801]_ , \new_[48804]_ ,
    \new_[48807]_ , \new_[48808]_ , \new_[48809]_ , \new_[48812]_ ,
    \new_[48815]_ , \new_[48816]_ , \new_[48819]_ , \new_[48822]_ ,
    \new_[48823]_ , \new_[48824]_ , \new_[48828]_ , \new_[48829]_ ,
    \new_[48832]_ , \new_[48835]_ , \new_[48836]_ , \new_[48837]_ ,
    \new_[48840]_ , \new_[48843]_ , \new_[48844]_ , \new_[48847]_ ,
    \new_[48850]_ , \new_[48851]_ , \new_[48852]_ , \new_[48856]_ ,
    \new_[48857]_ , \new_[48860]_ , \new_[48863]_ , \new_[48864]_ ,
    \new_[48865]_ , \new_[48868]_ , \new_[48871]_ , \new_[48872]_ ,
    \new_[48875]_ , \new_[48878]_ , \new_[48879]_ , \new_[48880]_ ,
    \new_[48884]_ , \new_[48885]_ , \new_[48888]_ , \new_[48891]_ ,
    \new_[48892]_ , \new_[48893]_ , \new_[48896]_ , \new_[48899]_ ,
    \new_[48900]_ , \new_[48903]_ , \new_[48906]_ , \new_[48907]_ ,
    \new_[48908]_ , \new_[48912]_ , \new_[48913]_ , \new_[48916]_ ,
    \new_[48919]_ , \new_[48920]_ , \new_[48921]_ , \new_[48924]_ ,
    \new_[48927]_ , \new_[48928]_ , \new_[48931]_ , \new_[48934]_ ,
    \new_[48935]_ , \new_[48936]_ , \new_[48940]_ , \new_[48941]_ ,
    \new_[48944]_ , \new_[48947]_ , \new_[48948]_ , \new_[48949]_ ,
    \new_[48952]_ , \new_[48955]_ , \new_[48956]_ , \new_[48959]_ ,
    \new_[48962]_ , \new_[48963]_ , \new_[48964]_ , \new_[48968]_ ,
    \new_[48969]_ , \new_[48972]_ , \new_[48975]_ , \new_[48976]_ ,
    \new_[48977]_ , \new_[48980]_ , \new_[48983]_ , \new_[48984]_ ,
    \new_[48987]_ , \new_[48990]_ , \new_[48991]_ , \new_[48992]_ ,
    \new_[48996]_ , \new_[48997]_ , \new_[49000]_ , \new_[49003]_ ,
    \new_[49004]_ , \new_[49005]_ , \new_[49008]_ , \new_[49011]_ ,
    \new_[49012]_ , \new_[49015]_ , \new_[49018]_ , \new_[49019]_ ,
    \new_[49020]_ , \new_[49024]_ , \new_[49025]_ , \new_[49028]_ ,
    \new_[49031]_ , \new_[49032]_ , \new_[49033]_ , \new_[49036]_ ,
    \new_[49039]_ , \new_[49040]_ , \new_[49043]_ , \new_[49046]_ ,
    \new_[49047]_ , \new_[49048]_ , \new_[49052]_ , \new_[49053]_ ,
    \new_[49056]_ , \new_[49059]_ , \new_[49060]_ , \new_[49061]_ ,
    \new_[49064]_ , \new_[49067]_ , \new_[49068]_ , \new_[49071]_ ,
    \new_[49074]_ , \new_[49075]_ , \new_[49076]_ , \new_[49080]_ ,
    \new_[49081]_ , \new_[49084]_ , \new_[49087]_ , \new_[49088]_ ,
    \new_[49089]_ , \new_[49092]_ , \new_[49095]_ , \new_[49096]_ ,
    \new_[49099]_ , \new_[49102]_ , \new_[49103]_ , \new_[49104]_ ,
    \new_[49108]_ , \new_[49109]_ , \new_[49112]_ , \new_[49115]_ ,
    \new_[49116]_ , \new_[49117]_ , \new_[49120]_ , \new_[49123]_ ,
    \new_[49124]_ , \new_[49127]_ , \new_[49130]_ , \new_[49131]_ ,
    \new_[49132]_ , \new_[49136]_ , \new_[49137]_ , \new_[49140]_ ,
    \new_[49143]_ , \new_[49144]_ , \new_[49145]_ , \new_[49148]_ ,
    \new_[49151]_ , \new_[49152]_ , \new_[49155]_ , \new_[49158]_ ,
    \new_[49159]_ , \new_[49160]_ , \new_[49164]_ , \new_[49165]_ ,
    \new_[49168]_ , \new_[49171]_ , \new_[49172]_ , \new_[49173]_ ,
    \new_[49176]_ , \new_[49179]_ , \new_[49180]_ , \new_[49183]_ ,
    \new_[49186]_ , \new_[49187]_ , \new_[49188]_ , \new_[49192]_ ,
    \new_[49193]_ , \new_[49196]_ , \new_[49199]_ , \new_[49200]_ ,
    \new_[49201]_ , \new_[49204]_ , \new_[49207]_ , \new_[49208]_ ,
    \new_[49211]_ , \new_[49214]_ , \new_[49215]_ , \new_[49216]_ ,
    \new_[49220]_ , \new_[49221]_ , \new_[49224]_ , \new_[49227]_ ,
    \new_[49228]_ , \new_[49229]_ , \new_[49232]_ , \new_[49235]_ ,
    \new_[49236]_ , \new_[49239]_ , \new_[49242]_ , \new_[49243]_ ,
    \new_[49244]_ , \new_[49248]_ , \new_[49249]_ , \new_[49252]_ ,
    \new_[49255]_ , \new_[49256]_ , \new_[49257]_ , \new_[49260]_ ,
    \new_[49263]_ , \new_[49264]_ , \new_[49267]_ , \new_[49270]_ ,
    \new_[49271]_ , \new_[49272]_ , \new_[49276]_ , \new_[49277]_ ,
    \new_[49280]_ , \new_[49283]_ , \new_[49284]_ , \new_[49285]_ ,
    \new_[49288]_ , \new_[49291]_ , \new_[49292]_ , \new_[49295]_ ,
    \new_[49298]_ , \new_[49299]_ , \new_[49300]_ , \new_[49304]_ ,
    \new_[49305]_ , \new_[49308]_ , \new_[49311]_ , \new_[49312]_ ,
    \new_[49313]_ , \new_[49316]_ , \new_[49319]_ , \new_[49320]_ ,
    \new_[49323]_ , \new_[49326]_ , \new_[49327]_ , \new_[49328]_ ,
    \new_[49332]_ , \new_[49333]_ , \new_[49336]_ , \new_[49339]_ ,
    \new_[49340]_ , \new_[49341]_ , \new_[49344]_ , \new_[49347]_ ,
    \new_[49348]_ , \new_[49351]_ , \new_[49354]_ , \new_[49355]_ ,
    \new_[49356]_ , \new_[49360]_ , \new_[49361]_ , \new_[49364]_ ,
    \new_[49367]_ , \new_[49368]_ , \new_[49369]_ , \new_[49372]_ ,
    \new_[49375]_ , \new_[49376]_ , \new_[49379]_ , \new_[49382]_ ,
    \new_[49383]_ , \new_[49384]_ , \new_[49388]_ , \new_[49389]_ ,
    \new_[49392]_ , \new_[49395]_ , \new_[49396]_ , \new_[49397]_ ,
    \new_[49400]_ , \new_[49403]_ , \new_[49404]_ , \new_[49407]_ ,
    \new_[49410]_ , \new_[49411]_ , \new_[49412]_ , \new_[49416]_ ,
    \new_[49417]_ , \new_[49420]_ , \new_[49423]_ , \new_[49424]_ ,
    \new_[49425]_ , \new_[49428]_ , \new_[49431]_ , \new_[49432]_ ,
    \new_[49435]_ , \new_[49438]_ , \new_[49439]_ , \new_[49440]_ ,
    \new_[49444]_ , \new_[49445]_ , \new_[49448]_ , \new_[49451]_ ,
    \new_[49452]_ , \new_[49453]_ , \new_[49456]_ , \new_[49459]_ ,
    \new_[49460]_ , \new_[49463]_ , \new_[49466]_ , \new_[49467]_ ,
    \new_[49468]_ , \new_[49472]_ , \new_[49473]_ , \new_[49476]_ ,
    \new_[49479]_ , \new_[49480]_ , \new_[49481]_ , \new_[49484]_ ,
    \new_[49487]_ , \new_[49488]_ , \new_[49491]_ , \new_[49494]_ ,
    \new_[49495]_ , \new_[49496]_ , \new_[49500]_ , \new_[49501]_ ,
    \new_[49504]_ , \new_[49507]_ , \new_[49508]_ , \new_[49509]_ ,
    \new_[49512]_ , \new_[49515]_ , \new_[49516]_ , \new_[49519]_ ,
    \new_[49522]_ , \new_[49523]_ , \new_[49524]_ , \new_[49528]_ ,
    \new_[49529]_ , \new_[49532]_ , \new_[49535]_ , \new_[49536]_ ,
    \new_[49537]_ , \new_[49540]_ , \new_[49543]_ , \new_[49544]_ ,
    \new_[49547]_ , \new_[49550]_ , \new_[49551]_ , \new_[49552]_ ,
    \new_[49556]_ , \new_[49557]_ , \new_[49560]_ , \new_[49563]_ ,
    \new_[49564]_ , \new_[49565]_ , \new_[49568]_ , \new_[49571]_ ,
    \new_[49572]_ , \new_[49575]_ , \new_[49578]_ , \new_[49579]_ ,
    \new_[49580]_ , \new_[49584]_ , \new_[49585]_ , \new_[49588]_ ,
    \new_[49591]_ , \new_[49592]_ , \new_[49593]_ , \new_[49596]_ ,
    \new_[49599]_ , \new_[49600]_ , \new_[49603]_ , \new_[49606]_ ,
    \new_[49607]_ , \new_[49608]_ , \new_[49612]_ , \new_[49613]_ ,
    \new_[49616]_ , \new_[49619]_ , \new_[49620]_ , \new_[49621]_ ,
    \new_[49624]_ , \new_[49627]_ , \new_[49628]_ , \new_[49631]_ ,
    \new_[49634]_ , \new_[49635]_ , \new_[49636]_ , \new_[49640]_ ,
    \new_[49641]_ , \new_[49644]_ , \new_[49647]_ , \new_[49648]_ ,
    \new_[49649]_ , \new_[49652]_ , \new_[49655]_ , \new_[49656]_ ,
    \new_[49659]_ , \new_[49662]_ , \new_[49663]_ , \new_[49664]_ ,
    \new_[49668]_ , \new_[49669]_ , \new_[49672]_ , \new_[49675]_ ,
    \new_[49676]_ , \new_[49677]_ , \new_[49680]_ , \new_[49683]_ ,
    \new_[49684]_ , \new_[49687]_ , \new_[49690]_ , \new_[49691]_ ,
    \new_[49692]_ , \new_[49696]_ , \new_[49697]_ , \new_[49700]_ ,
    \new_[49703]_ , \new_[49704]_ , \new_[49705]_ , \new_[49708]_ ,
    \new_[49711]_ , \new_[49712]_ , \new_[49715]_ , \new_[49718]_ ,
    \new_[49719]_ , \new_[49720]_ , \new_[49724]_ , \new_[49725]_ ,
    \new_[49728]_ , \new_[49731]_ , \new_[49732]_ , \new_[49733]_ ,
    \new_[49736]_ , \new_[49739]_ , \new_[49740]_ , \new_[49743]_ ,
    \new_[49746]_ , \new_[49747]_ , \new_[49748]_ , \new_[49752]_ ,
    \new_[49753]_ , \new_[49756]_ , \new_[49759]_ , \new_[49760]_ ,
    \new_[49761]_ , \new_[49764]_ , \new_[49767]_ , \new_[49768]_ ,
    \new_[49771]_ , \new_[49774]_ , \new_[49775]_ , \new_[49776]_ ,
    \new_[49780]_ , \new_[49781]_ , \new_[49784]_ , \new_[49787]_ ,
    \new_[49788]_ , \new_[49789]_ , \new_[49792]_ , \new_[49795]_ ,
    \new_[49796]_ , \new_[49799]_ , \new_[49802]_ , \new_[49803]_ ,
    \new_[49804]_ , \new_[49808]_ , \new_[49809]_ , \new_[49812]_ ,
    \new_[49815]_ , \new_[49816]_ , \new_[49817]_ , \new_[49820]_ ,
    \new_[49823]_ , \new_[49824]_ , \new_[49827]_ , \new_[49830]_ ,
    \new_[49831]_ , \new_[49832]_ , \new_[49836]_ , \new_[49837]_ ,
    \new_[49840]_ , \new_[49843]_ , \new_[49844]_ , \new_[49845]_ ,
    \new_[49848]_ , \new_[49851]_ , \new_[49852]_ , \new_[49855]_ ,
    \new_[49858]_ , \new_[49859]_ , \new_[49860]_ , \new_[49864]_ ,
    \new_[49865]_ , \new_[49868]_ , \new_[49871]_ , \new_[49872]_ ,
    \new_[49873]_ , \new_[49876]_ , \new_[49879]_ , \new_[49880]_ ,
    \new_[49883]_ , \new_[49886]_ , \new_[49887]_ , \new_[49888]_ ,
    \new_[49892]_ , \new_[49893]_ , \new_[49896]_ , \new_[49899]_ ,
    \new_[49900]_ , \new_[49901]_ , \new_[49904]_ , \new_[49907]_ ,
    \new_[49908]_ , \new_[49911]_ , \new_[49914]_ , \new_[49915]_ ,
    \new_[49916]_ , \new_[49920]_ , \new_[49921]_ , \new_[49924]_ ,
    \new_[49927]_ , \new_[49928]_ , \new_[49929]_ , \new_[49932]_ ,
    \new_[49935]_ , \new_[49936]_ , \new_[49939]_ , \new_[49942]_ ,
    \new_[49943]_ , \new_[49944]_ , \new_[49948]_ , \new_[49949]_ ,
    \new_[49952]_ , \new_[49955]_ , \new_[49956]_ , \new_[49957]_ ,
    \new_[49960]_ , \new_[49963]_ , \new_[49964]_ , \new_[49967]_ ,
    \new_[49970]_ , \new_[49971]_ , \new_[49972]_ , \new_[49976]_ ,
    \new_[49977]_ , \new_[49980]_ , \new_[49983]_ , \new_[49984]_ ,
    \new_[49985]_ , \new_[49988]_ , \new_[49991]_ , \new_[49992]_ ,
    \new_[49995]_ , \new_[49998]_ , \new_[49999]_ , \new_[50000]_ ,
    \new_[50004]_ , \new_[50005]_ , \new_[50008]_ , \new_[50011]_ ,
    \new_[50012]_ , \new_[50013]_ , \new_[50016]_ , \new_[50019]_ ,
    \new_[50020]_ , \new_[50023]_ , \new_[50026]_ , \new_[50027]_ ,
    \new_[50028]_ , \new_[50032]_ , \new_[50033]_ , \new_[50036]_ ,
    \new_[50039]_ , \new_[50040]_ , \new_[50041]_ , \new_[50044]_ ,
    \new_[50047]_ , \new_[50048]_ , \new_[50051]_ , \new_[50054]_ ,
    \new_[50055]_ , \new_[50056]_ , \new_[50060]_ , \new_[50061]_ ,
    \new_[50064]_ , \new_[50067]_ , \new_[50068]_ , \new_[50069]_ ,
    \new_[50072]_ , \new_[50075]_ , \new_[50076]_ , \new_[50079]_ ,
    \new_[50082]_ , \new_[50083]_ , \new_[50084]_ , \new_[50088]_ ,
    \new_[50089]_ , \new_[50092]_ , \new_[50095]_ , \new_[50096]_ ,
    \new_[50097]_ , \new_[50100]_ , \new_[50103]_ , \new_[50104]_ ,
    \new_[50107]_ , \new_[50110]_ , \new_[50111]_ , \new_[50112]_ ,
    \new_[50116]_ , \new_[50117]_ , \new_[50120]_ , \new_[50123]_ ,
    \new_[50124]_ , \new_[50125]_ , \new_[50128]_ , \new_[50131]_ ,
    \new_[50132]_ , \new_[50135]_ , \new_[50138]_ , \new_[50139]_ ,
    \new_[50140]_ , \new_[50144]_ , \new_[50145]_ , \new_[50148]_ ,
    \new_[50151]_ , \new_[50152]_ , \new_[50153]_ , \new_[50156]_ ,
    \new_[50159]_ , \new_[50160]_ , \new_[50163]_ , \new_[50166]_ ,
    \new_[50167]_ , \new_[50168]_ , \new_[50172]_ , \new_[50173]_ ,
    \new_[50176]_ , \new_[50179]_ , \new_[50180]_ , \new_[50181]_ ,
    \new_[50184]_ , \new_[50187]_ , \new_[50188]_ , \new_[50191]_ ,
    \new_[50194]_ , \new_[50195]_ , \new_[50196]_ , \new_[50200]_ ,
    \new_[50201]_ , \new_[50204]_ , \new_[50207]_ , \new_[50208]_ ,
    \new_[50209]_ , \new_[50212]_ , \new_[50215]_ , \new_[50216]_ ,
    \new_[50219]_ , \new_[50222]_ , \new_[50223]_ , \new_[50224]_ ,
    \new_[50228]_ , \new_[50229]_ , \new_[50232]_ , \new_[50235]_ ,
    \new_[50236]_ , \new_[50237]_ , \new_[50240]_ , \new_[50243]_ ,
    \new_[50244]_ , \new_[50247]_ , \new_[50250]_ , \new_[50251]_ ,
    \new_[50252]_ , \new_[50256]_ , \new_[50257]_ , \new_[50260]_ ,
    \new_[50263]_ , \new_[50264]_ , \new_[50265]_ , \new_[50268]_ ,
    \new_[50271]_ , \new_[50272]_ , \new_[50275]_ , \new_[50278]_ ,
    \new_[50279]_ , \new_[50280]_ , \new_[50284]_ , \new_[50285]_ ,
    \new_[50288]_ , \new_[50291]_ , \new_[50292]_ , \new_[50293]_ ,
    \new_[50296]_ , \new_[50299]_ , \new_[50300]_ , \new_[50303]_ ,
    \new_[50306]_ , \new_[50307]_ , \new_[50308]_ , \new_[50312]_ ,
    \new_[50313]_ , \new_[50316]_ , \new_[50319]_ , \new_[50320]_ ,
    \new_[50321]_ , \new_[50324]_ , \new_[50327]_ , \new_[50328]_ ,
    \new_[50331]_ , \new_[50334]_ , \new_[50335]_ , \new_[50336]_ ,
    \new_[50340]_ , \new_[50341]_ , \new_[50344]_ , \new_[50347]_ ,
    \new_[50348]_ , \new_[50349]_ , \new_[50352]_ , \new_[50355]_ ,
    \new_[50356]_ , \new_[50359]_ , \new_[50362]_ , \new_[50363]_ ,
    \new_[50364]_ , \new_[50368]_ , \new_[50369]_ , \new_[50372]_ ,
    \new_[50375]_ , \new_[50376]_ , \new_[50377]_ , \new_[50380]_ ,
    \new_[50383]_ , \new_[50384]_ , \new_[50387]_ , \new_[50390]_ ,
    \new_[50391]_ , \new_[50392]_ , \new_[50396]_ , \new_[50397]_ ,
    \new_[50400]_ , \new_[50403]_ , \new_[50404]_ , \new_[50405]_ ,
    \new_[50408]_ , \new_[50411]_ , \new_[50412]_ , \new_[50415]_ ,
    \new_[50418]_ , \new_[50419]_ , \new_[50420]_ , \new_[50424]_ ,
    \new_[50425]_ , \new_[50428]_ , \new_[50431]_ , \new_[50432]_ ,
    \new_[50433]_ , \new_[50436]_ , \new_[50439]_ , \new_[50440]_ ,
    \new_[50443]_ , \new_[50446]_ , \new_[50447]_ , \new_[50448]_ ,
    \new_[50452]_ , \new_[50453]_ , \new_[50456]_ , \new_[50459]_ ,
    \new_[50460]_ , \new_[50461]_ , \new_[50464]_ , \new_[50467]_ ,
    \new_[50468]_ , \new_[50471]_ , \new_[50474]_ , \new_[50475]_ ,
    \new_[50476]_ , \new_[50480]_ , \new_[50481]_ , \new_[50484]_ ,
    \new_[50487]_ , \new_[50488]_ , \new_[50489]_ , \new_[50492]_ ,
    \new_[50495]_ , \new_[50496]_ , \new_[50499]_ , \new_[50502]_ ,
    \new_[50503]_ , \new_[50504]_ , \new_[50508]_ , \new_[50509]_ ,
    \new_[50512]_ , \new_[50515]_ , \new_[50516]_ , \new_[50517]_ ,
    \new_[50520]_ , \new_[50523]_ , \new_[50524]_ , \new_[50527]_ ,
    \new_[50530]_ , \new_[50531]_ , \new_[50532]_ , \new_[50536]_ ,
    \new_[50537]_ , \new_[50540]_ , \new_[50543]_ , \new_[50544]_ ,
    \new_[50545]_ , \new_[50548]_ , \new_[50551]_ , \new_[50552]_ ,
    \new_[50555]_ , \new_[50558]_ , \new_[50559]_ , \new_[50560]_ ,
    \new_[50564]_ , \new_[50565]_ , \new_[50568]_ , \new_[50571]_ ,
    \new_[50572]_ , \new_[50573]_ , \new_[50576]_ , \new_[50579]_ ,
    \new_[50580]_ , \new_[50583]_ , \new_[50586]_ , \new_[50587]_ ,
    \new_[50588]_ , \new_[50592]_ , \new_[50593]_ , \new_[50596]_ ,
    \new_[50599]_ , \new_[50600]_ , \new_[50601]_ , \new_[50604]_ ,
    \new_[50607]_ , \new_[50608]_ , \new_[50611]_ , \new_[50614]_ ,
    \new_[50615]_ , \new_[50616]_ , \new_[50620]_ , \new_[50621]_ ,
    \new_[50624]_ , \new_[50627]_ , \new_[50628]_ , \new_[50629]_ ,
    \new_[50632]_ , \new_[50635]_ , \new_[50636]_ , \new_[50639]_ ,
    \new_[50642]_ , \new_[50643]_ , \new_[50644]_ , \new_[50648]_ ,
    \new_[50649]_ , \new_[50652]_ , \new_[50655]_ , \new_[50656]_ ,
    \new_[50657]_ , \new_[50660]_ , \new_[50663]_ , \new_[50664]_ ,
    \new_[50667]_ , \new_[50670]_ , \new_[50671]_ , \new_[50672]_ ,
    \new_[50676]_ , \new_[50677]_ , \new_[50680]_ , \new_[50683]_ ,
    \new_[50684]_ , \new_[50685]_ , \new_[50688]_ , \new_[50691]_ ,
    \new_[50692]_ , \new_[50695]_ , \new_[50698]_ , \new_[50699]_ ,
    \new_[50700]_ , \new_[50704]_ , \new_[50705]_ , \new_[50708]_ ,
    \new_[50711]_ , \new_[50712]_ , \new_[50713]_ , \new_[50716]_ ,
    \new_[50719]_ , \new_[50720]_ , \new_[50723]_ , \new_[50726]_ ,
    \new_[50727]_ , \new_[50728]_ , \new_[50732]_ , \new_[50733]_ ,
    \new_[50736]_ , \new_[50739]_ , \new_[50740]_ , \new_[50741]_ ,
    \new_[50744]_ , \new_[50747]_ , \new_[50748]_ , \new_[50751]_ ,
    \new_[50754]_ , \new_[50755]_ , \new_[50756]_ , \new_[50760]_ ,
    \new_[50761]_ , \new_[50764]_ , \new_[50767]_ , \new_[50768]_ ,
    \new_[50769]_ , \new_[50772]_ , \new_[50775]_ , \new_[50776]_ ,
    \new_[50779]_ , \new_[50782]_ , \new_[50783]_ , \new_[50784]_ ,
    \new_[50788]_ , \new_[50789]_ , \new_[50792]_ , \new_[50795]_ ,
    \new_[50796]_ , \new_[50797]_ , \new_[50800]_ , \new_[50803]_ ,
    \new_[50804]_ , \new_[50807]_ , \new_[50810]_ , \new_[50811]_ ,
    \new_[50812]_ , \new_[50816]_ , \new_[50817]_ , \new_[50820]_ ,
    \new_[50823]_ , \new_[50824]_ , \new_[50825]_ , \new_[50828]_ ,
    \new_[50831]_ , \new_[50832]_ , \new_[50835]_ , \new_[50838]_ ,
    \new_[50839]_ , \new_[50840]_ , \new_[50844]_ , \new_[50845]_ ,
    \new_[50848]_ , \new_[50851]_ , \new_[50852]_ , \new_[50853]_ ,
    \new_[50856]_ , \new_[50859]_ , \new_[50860]_ , \new_[50863]_ ,
    \new_[50866]_ , \new_[50867]_ , \new_[50868]_ , \new_[50872]_ ,
    \new_[50873]_ , \new_[50876]_ , \new_[50879]_ , \new_[50880]_ ,
    \new_[50881]_ , \new_[50884]_ , \new_[50887]_ , \new_[50888]_ ,
    \new_[50891]_ , \new_[50894]_ , \new_[50895]_ , \new_[50896]_ ,
    \new_[50900]_ , \new_[50901]_ , \new_[50904]_ , \new_[50907]_ ,
    \new_[50908]_ , \new_[50909]_ , \new_[50912]_ , \new_[50915]_ ,
    \new_[50916]_ , \new_[50919]_ , \new_[50922]_ , \new_[50923]_ ,
    \new_[50924]_ , \new_[50928]_ , \new_[50929]_ , \new_[50932]_ ,
    \new_[50935]_ , \new_[50936]_ , \new_[50937]_ , \new_[50940]_ ,
    \new_[50943]_ , \new_[50944]_ , \new_[50947]_ , \new_[50950]_ ,
    \new_[50951]_ , \new_[50952]_ , \new_[50956]_ , \new_[50957]_ ,
    \new_[50960]_ , \new_[50963]_ , \new_[50964]_ , \new_[50965]_ ,
    \new_[50968]_ , \new_[50971]_ , \new_[50972]_ , \new_[50975]_ ,
    \new_[50978]_ , \new_[50979]_ , \new_[50980]_ , \new_[50984]_ ,
    \new_[50985]_ , \new_[50988]_ , \new_[50991]_ , \new_[50992]_ ,
    \new_[50993]_ , \new_[50996]_ , \new_[50999]_ , \new_[51000]_ ,
    \new_[51003]_ , \new_[51006]_ , \new_[51007]_ , \new_[51008]_ ,
    \new_[51012]_ , \new_[51013]_ , \new_[51016]_ , \new_[51019]_ ,
    \new_[51020]_ , \new_[51021]_ , \new_[51024]_ , \new_[51027]_ ,
    \new_[51028]_ , \new_[51031]_ , \new_[51034]_ , \new_[51035]_ ,
    \new_[51036]_ , \new_[51040]_ , \new_[51041]_ , \new_[51044]_ ,
    \new_[51047]_ , \new_[51048]_ , \new_[51049]_ , \new_[51052]_ ,
    \new_[51055]_ , \new_[51056]_ , \new_[51059]_ , \new_[51062]_ ,
    \new_[51063]_ , \new_[51064]_ , \new_[51068]_ , \new_[51069]_ ,
    \new_[51072]_ , \new_[51075]_ , \new_[51076]_ , \new_[51077]_ ,
    \new_[51080]_ , \new_[51083]_ , \new_[51084]_ , \new_[51087]_ ,
    \new_[51090]_ , \new_[51091]_ , \new_[51092]_ , \new_[51096]_ ,
    \new_[51097]_ , \new_[51100]_ , \new_[51103]_ , \new_[51104]_ ,
    \new_[51105]_ , \new_[51108]_ , \new_[51111]_ , \new_[51112]_ ,
    \new_[51115]_ , \new_[51118]_ , \new_[51119]_ , \new_[51120]_ ,
    \new_[51124]_ , \new_[51125]_ , \new_[51128]_ , \new_[51131]_ ,
    \new_[51132]_ , \new_[51133]_ , \new_[51136]_ , \new_[51139]_ ,
    \new_[51140]_ , \new_[51143]_ , \new_[51146]_ , \new_[51147]_ ,
    \new_[51148]_ , \new_[51152]_ , \new_[51153]_ , \new_[51156]_ ,
    \new_[51159]_ , \new_[51160]_ , \new_[51161]_ , \new_[51164]_ ,
    \new_[51167]_ , \new_[51168]_ , \new_[51171]_ , \new_[51174]_ ,
    \new_[51175]_ , \new_[51176]_ , \new_[51180]_ , \new_[51181]_ ,
    \new_[51184]_ , \new_[51187]_ , \new_[51188]_ , \new_[51189]_ ,
    \new_[51192]_ , \new_[51195]_ , \new_[51196]_ , \new_[51199]_ ,
    \new_[51202]_ , \new_[51203]_ , \new_[51204]_ , \new_[51208]_ ,
    \new_[51209]_ , \new_[51212]_ , \new_[51215]_ , \new_[51216]_ ,
    \new_[51217]_ , \new_[51220]_ , \new_[51223]_ , \new_[51224]_ ,
    \new_[51227]_ , \new_[51230]_ , \new_[51231]_ , \new_[51232]_ ,
    \new_[51236]_ , \new_[51237]_ , \new_[51240]_ , \new_[51243]_ ,
    \new_[51244]_ , \new_[51245]_ , \new_[51248]_ , \new_[51251]_ ,
    \new_[51252]_ , \new_[51255]_ , \new_[51258]_ , \new_[51259]_ ,
    \new_[51260]_ , \new_[51264]_ , \new_[51265]_ , \new_[51268]_ ,
    \new_[51271]_ , \new_[51272]_ , \new_[51273]_ , \new_[51276]_ ,
    \new_[51279]_ , \new_[51280]_ , \new_[51283]_ , \new_[51286]_ ,
    \new_[51287]_ , \new_[51288]_ , \new_[51292]_ , \new_[51293]_ ,
    \new_[51296]_ , \new_[51299]_ , \new_[51300]_ , \new_[51301]_ ,
    \new_[51304]_ , \new_[51307]_ , \new_[51308]_ , \new_[51311]_ ,
    \new_[51314]_ , \new_[51315]_ , \new_[51316]_ , \new_[51320]_ ,
    \new_[51321]_ , \new_[51324]_ , \new_[51327]_ , \new_[51328]_ ,
    \new_[51329]_ , \new_[51332]_ , \new_[51335]_ , \new_[51336]_ ,
    \new_[51339]_ , \new_[51342]_ , \new_[51343]_ , \new_[51344]_ ,
    \new_[51348]_ , \new_[51349]_ , \new_[51352]_ , \new_[51355]_ ,
    \new_[51356]_ , \new_[51357]_ , \new_[51360]_ , \new_[51363]_ ,
    \new_[51364]_ , \new_[51367]_ , \new_[51370]_ , \new_[51371]_ ,
    \new_[51372]_ , \new_[51376]_ , \new_[51377]_ , \new_[51380]_ ,
    \new_[51383]_ , \new_[51384]_ , \new_[51385]_ , \new_[51388]_ ,
    \new_[51391]_ , \new_[51392]_ , \new_[51395]_ , \new_[51398]_ ,
    \new_[51399]_ , \new_[51400]_ , \new_[51404]_ , \new_[51405]_ ,
    \new_[51408]_ , \new_[51411]_ , \new_[51412]_ , \new_[51413]_ ,
    \new_[51416]_ , \new_[51419]_ , \new_[51420]_ , \new_[51423]_ ,
    \new_[51426]_ , \new_[51427]_ , \new_[51428]_ , \new_[51432]_ ,
    \new_[51433]_ , \new_[51436]_ , \new_[51439]_ , \new_[51440]_ ,
    \new_[51441]_ , \new_[51444]_ , \new_[51447]_ , \new_[51448]_ ,
    \new_[51451]_ , \new_[51454]_ , \new_[51455]_ , \new_[51456]_ ,
    \new_[51460]_ , \new_[51461]_ , \new_[51464]_ , \new_[51467]_ ,
    \new_[51468]_ , \new_[51469]_ , \new_[51472]_ , \new_[51475]_ ,
    \new_[51476]_ , \new_[51479]_ , \new_[51482]_ , \new_[51483]_ ,
    \new_[51484]_ , \new_[51488]_ , \new_[51489]_ , \new_[51492]_ ,
    \new_[51495]_ , \new_[51496]_ , \new_[51497]_ , \new_[51500]_ ,
    \new_[51503]_ , \new_[51504]_ , \new_[51507]_ , \new_[51510]_ ,
    \new_[51511]_ , \new_[51512]_ , \new_[51516]_ , \new_[51517]_ ,
    \new_[51520]_ , \new_[51523]_ , \new_[51524]_ , \new_[51525]_ ,
    \new_[51528]_ , \new_[51531]_ , \new_[51532]_ , \new_[51535]_ ,
    \new_[51538]_ , \new_[51539]_ , \new_[51540]_ , \new_[51544]_ ,
    \new_[51545]_ , \new_[51548]_ , \new_[51551]_ , \new_[51552]_ ,
    \new_[51553]_ , \new_[51556]_ , \new_[51559]_ , \new_[51560]_ ,
    \new_[51563]_ , \new_[51566]_ , \new_[51567]_ , \new_[51568]_ ,
    \new_[51572]_ , \new_[51573]_ , \new_[51576]_ , \new_[51579]_ ,
    \new_[51580]_ , \new_[51581]_ , \new_[51584]_ , \new_[51587]_ ,
    \new_[51588]_ , \new_[51591]_ , \new_[51594]_ , \new_[51595]_ ,
    \new_[51596]_ , \new_[51600]_ , \new_[51601]_ , \new_[51604]_ ,
    \new_[51607]_ , \new_[51608]_ , \new_[51609]_ , \new_[51612]_ ,
    \new_[51615]_ , \new_[51616]_ , \new_[51619]_ , \new_[51622]_ ,
    \new_[51623]_ , \new_[51624]_ , \new_[51628]_ , \new_[51629]_ ,
    \new_[51632]_ , \new_[51635]_ , \new_[51636]_ , \new_[51637]_ ,
    \new_[51640]_ , \new_[51643]_ , \new_[51644]_ , \new_[51647]_ ,
    \new_[51650]_ , \new_[51651]_ , \new_[51652]_ , \new_[51656]_ ,
    \new_[51657]_ , \new_[51660]_ , \new_[51663]_ , \new_[51664]_ ,
    \new_[51665]_ , \new_[51668]_ , \new_[51671]_ , \new_[51672]_ ,
    \new_[51675]_ , \new_[51678]_ , \new_[51679]_ , \new_[51680]_ ,
    \new_[51684]_ , \new_[51685]_ , \new_[51688]_ , \new_[51691]_ ,
    \new_[51692]_ , \new_[51693]_ , \new_[51696]_ , \new_[51699]_ ,
    \new_[51700]_ , \new_[51703]_ , \new_[51706]_ , \new_[51707]_ ,
    \new_[51708]_ , \new_[51712]_ , \new_[51713]_ , \new_[51716]_ ,
    \new_[51719]_ , \new_[51720]_ , \new_[51721]_ , \new_[51724]_ ,
    \new_[51727]_ , \new_[51728]_ , \new_[51731]_ , \new_[51734]_ ,
    \new_[51735]_ , \new_[51736]_ , \new_[51740]_ , \new_[51741]_ ,
    \new_[51744]_ , \new_[51747]_ , \new_[51748]_ , \new_[51749]_ ,
    \new_[51752]_ , \new_[51755]_ , \new_[51756]_ , \new_[51759]_ ,
    \new_[51762]_ , \new_[51763]_ , \new_[51764]_ , \new_[51768]_ ,
    \new_[51769]_ , \new_[51772]_ , \new_[51775]_ , \new_[51776]_ ,
    \new_[51777]_ , \new_[51780]_ , \new_[51783]_ , \new_[51784]_ ,
    \new_[51787]_ , \new_[51790]_ , \new_[51791]_ , \new_[51792]_ ,
    \new_[51796]_ , \new_[51797]_ , \new_[51800]_ , \new_[51803]_ ,
    \new_[51804]_ , \new_[51805]_ , \new_[51808]_ , \new_[51811]_ ,
    \new_[51812]_ , \new_[51815]_ , \new_[51818]_ , \new_[51819]_ ,
    \new_[51820]_ , \new_[51824]_ , \new_[51825]_ , \new_[51828]_ ,
    \new_[51831]_ , \new_[51832]_ , \new_[51833]_ , \new_[51836]_ ,
    \new_[51839]_ , \new_[51840]_ , \new_[51843]_ , \new_[51846]_ ,
    \new_[51847]_ , \new_[51848]_ , \new_[51852]_ , \new_[51853]_ ,
    \new_[51856]_ , \new_[51859]_ , \new_[51860]_ , \new_[51861]_ ,
    \new_[51864]_ , \new_[51867]_ , \new_[51868]_ , \new_[51871]_ ,
    \new_[51874]_ , \new_[51875]_ , \new_[51876]_ , \new_[51880]_ ,
    \new_[51881]_ , \new_[51884]_ , \new_[51887]_ , \new_[51888]_ ,
    \new_[51889]_ , \new_[51892]_ , \new_[51895]_ , \new_[51896]_ ,
    \new_[51899]_ , \new_[51902]_ , \new_[51903]_ , \new_[51904]_ ,
    \new_[51908]_ , \new_[51909]_ , \new_[51912]_ , \new_[51915]_ ,
    \new_[51916]_ , \new_[51917]_ , \new_[51920]_ , \new_[51923]_ ,
    \new_[51924]_ , \new_[51927]_ , \new_[51930]_ , \new_[51931]_ ,
    \new_[51932]_ , \new_[51936]_ , \new_[51937]_ , \new_[51940]_ ,
    \new_[51943]_ , \new_[51944]_ , \new_[51945]_ , \new_[51948]_ ,
    \new_[51951]_ , \new_[51952]_ , \new_[51955]_ , \new_[51958]_ ,
    \new_[51959]_ , \new_[51960]_ , \new_[51964]_ , \new_[51965]_ ,
    \new_[51968]_ , \new_[51971]_ , \new_[51972]_ , \new_[51973]_ ,
    \new_[51976]_ , \new_[51979]_ , \new_[51980]_ , \new_[51983]_ ,
    \new_[51986]_ , \new_[51987]_ , \new_[51988]_ , \new_[51992]_ ,
    \new_[51993]_ , \new_[51996]_ , \new_[51999]_ , \new_[52000]_ ,
    \new_[52001]_ , \new_[52004]_ , \new_[52007]_ , \new_[52008]_ ,
    \new_[52011]_ , \new_[52014]_ , \new_[52015]_ , \new_[52016]_ ,
    \new_[52020]_ , \new_[52021]_ , \new_[52024]_ , \new_[52027]_ ,
    \new_[52028]_ , \new_[52029]_ , \new_[52032]_ , \new_[52035]_ ,
    \new_[52036]_ , \new_[52039]_ , \new_[52042]_ , \new_[52043]_ ,
    \new_[52044]_ , \new_[52048]_ , \new_[52049]_ , \new_[52052]_ ,
    \new_[52055]_ , \new_[52056]_ , \new_[52057]_ , \new_[52060]_ ,
    \new_[52063]_ , \new_[52064]_ , \new_[52067]_ , \new_[52070]_ ,
    \new_[52071]_ , \new_[52072]_ , \new_[52076]_ , \new_[52077]_ ,
    \new_[52080]_ , \new_[52083]_ , \new_[52084]_ , \new_[52085]_ ,
    \new_[52088]_ , \new_[52091]_ , \new_[52092]_ , \new_[52095]_ ,
    \new_[52098]_ , \new_[52099]_ , \new_[52100]_ , \new_[52104]_ ,
    \new_[52105]_ , \new_[52108]_ , \new_[52111]_ , \new_[52112]_ ,
    \new_[52113]_ , \new_[52116]_ , \new_[52119]_ , \new_[52120]_ ,
    \new_[52123]_ , \new_[52126]_ , \new_[52127]_ , \new_[52128]_ ,
    \new_[52132]_ , \new_[52133]_ , \new_[52136]_ , \new_[52139]_ ,
    \new_[52140]_ , \new_[52141]_ , \new_[52144]_ , \new_[52147]_ ,
    \new_[52148]_ , \new_[52151]_ , \new_[52154]_ , \new_[52155]_ ,
    \new_[52156]_ , \new_[52160]_ , \new_[52161]_ , \new_[52164]_ ,
    \new_[52167]_ , \new_[52168]_ , \new_[52169]_ , \new_[52172]_ ,
    \new_[52175]_ , \new_[52176]_ , \new_[52179]_ , \new_[52182]_ ,
    \new_[52183]_ , \new_[52184]_ , \new_[52188]_ , \new_[52189]_ ,
    \new_[52192]_ , \new_[52195]_ , \new_[52196]_ , \new_[52197]_ ,
    \new_[52200]_ , \new_[52203]_ , \new_[52204]_ , \new_[52207]_ ,
    \new_[52210]_ , \new_[52211]_ , \new_[52212]_ , \new_[52216]_ ,
    \new_[52217]_ , \new_[52220]_ , \new_[52223]_ , \new_[52224]_ ,
    \new_[52225]_ , \new_[52228]_ , \new_[52231]_ , \new_[52232]_ ,
    \new_[52235]_ , \new_[52238]_ , \new_[52239]_ , \new_[52240]_ ,
    \new_[52244]_ , \new_[52245]_ , \new_[52248]_ , \new_[52251]_ ,
    \new_[52252]_ , \new_[52253]_ , \new_[52256]_ , \new_[52259]_ ,
    \new_[52260]_ , \new_[52263]_ , \new_[52266]_ , \new_[52267]_ ,
    \new_[52268]_ , \new_[52272]_ , \new_[52273]_ , \new_[52276]_ ,
    \new_[52279]_ , \new_[52280]_ , \new_[52281]_ , \new_[52284]_ ,
    \new_[52287]_ , \new_[52288]_ , \new_[52291]_ , \new_[52294]_ ,
    \new_[52295]_ , \new_[52296]_ , \new_[52300]_ , \new_[52301]_ ,
    \new_[52304]_ , \new_[52307]_ , \new_[52308]_ , \new_[52309]_ ,
    \new_[52312]_ , \new_[52315]_ , \new_[52316]_ , \new_[52319]_ ,
    \new_[52322]_ , \new_[52323]_ , \new_[52324]_ , \new_[52328]_ ,
    \new_[52329]_ , \new_[52332]_ , \new_[52335]_ , \new_[52336]_ ,
    \new_[52337]_ , \new_[52340]_ , \new_[52343]_ , \new_[52344]_ ,
    \new_[52347]_ , \new_[52350]_ , \new_[52351]_ , \new_[52352]_ ,
    \new_[52356]_ , \new_[52357]_ , \new_[52360]_ , \new_[52363]_ ,
    \new_[52364]_ , \new_[52365]_ , \new_[52368]_ , \new_[52371]_ ,
    \new_[52372]_ , \new_[52375]_ , \new_[52378]_ , \new_[52379]_ ,
    \new_[52380]_ , \new_[52384]_ , \new_[52385]_ , \new_[52388]_ ,
    \new_[52391]_ , \new_[52392]_ , \new_[52393]_ , \new_[52396]_ ,
    \new_[52399]_ , \new_[52400]_ , \new_[52403]_ , \new_[52406]_ ,
    \new_[52407]_ , \new_[52408]_ , \new_[52412]_ , \new_[52413]_ ,
    \new_[52416]_ , \new_[52419]_ , \new_[52420]_ , \new_[52421]_ ,
    \new_[52424]_ , \new_[52427]_ , \new_[52428]_ , \new_[52431]_ ,
    \new_[52434]_ , \new_[52435]_ , \new_[52436]_ , \new_[52440]_ ,
    \new_[52441]_ , \new_[52444]_ , \new_[52447]_ , \new_[52448]_ ,
    \new_[52449]_ , \new_[52452]_ , \new_[52455]_ , \new_[52456]_ ,
    \new_[52459]_ , \new_[52462]_ , \new_[52463]_ , \new_[52464]_ ,
    \new_[52468]_ , \new_[52469]_ , \new_[52472]_ , \new_[52475]_ ,
    \new_[52476]_ , \new_[52477]_ , \new_[52480]_ , \new_[52483]_ ,
    \new_[52484]_ , \new_[52487]_ , \new_[52490]_ , \new_[52491]_ ,
    \new_[52492]_ , \new_[52496]_ , \new_[52497]_ , \new_[52500]_ ,
    \new_[52503]_ , \new_[52504]_ , \new_[52505]_ , \new_[52508]_ ,
    \new_[52511]_ , \new_[52512]_ , \new_[52515]_ , \new_[52518]_ ,
    \new_[52519]_ , \new_[52520]_ , \new_[52524]_ , \new_[52525]_ ,
    \new_[52528]_ , \new_[52531]_ , \new_[52532]_ , \new_[52533]_ ,
    \new_[52536]_ , \new_[52539]_ , \new_[52540]_ , \new_[52543]_ ,
    \new_[52546]_ , \new_[52547]_ , \new_[52548]_ , \new_[52552]_ ,
    \new_[52553]_ , \new_[52556]_ , \new_[52559]_ , \new_[52560]_ ,
    \new_[52561]_ , \new_[52564]_ , \new_[52567]_ , \new_[52568]_ ,
    \new_[52571]_ , \new_[52574]_ , \new_[52575]_ , \new_[52576]_ ,
    \new_[52580]_ , \new_[52581]_ , \new_[52584]_ , \new_[52587]_ ,
    \new_[52588]_ , \new_[52589]_ , \new_[52592]_ , \new_[52595]_ ,
    \new_[52596]_ , \new_[52599]_ , \new_[52602]_ , \new_[52603]_ ,
    \new_[52604]_ , \new_[52608]_ , \new_[52609]_ , \new_[52612]_ ,
    \new_[52615]_ , \new_[52616]_ , \new_[52617]_ , \new_[52620]_ ,
    \new_[52623]_ , \new_[52624]_ , \new_[52627]_ , \new_[52630]_ ,
    \new_[52631]_ , \new_[52632]_ , \new_[52636]_ , \new_[52637]_ ,
    \new_[52640]_ , \new_[52643]_ , \new_[52644]_ , \new_[52645]_ ,
    \new_[52648]_ , \new_[52651]_ , \new_[52652]_ , \new_[52655]_ ,
    \new_[52658]_ , \new_[52659]_ , \new_[52660]_ , \new_[52664]_ ,
    \new_[52665]_ , \new_[52668]_ , \new_[52671]_ , \new_[52672]_ ,
    \new_[52673]_ , \new_[52676]_ , \new_[52679]_ , \new_[52680]_ ,
    \new_[52683]_ , \new_[52686]_ , \new_[52687]_ , \new_[52688]_ ,
    \new_[52692]_ , \new_[52693]_ , \new_[52696]_ , \new_[52699]_ ,
    \new_[52700]_ , \new_[52701]_ , \new_[52704]_ , \new_[52707]_ ,
    \new_[52708]_ , \new_[52711]_ , \new_[52714]_ , \new_[52715]_ ,
    \new_[52716]_ , \new_[52720]_ , \new_[52721]_ , \new_[52724]_ ,
    \new_[52727]_ , \new_[52728]_ , \new_[52729]_ , \new_[52732]_ ,
    \new_[52735]_ , \new_[52736]_ , \new_[52739]_ , \new_[52742]_ ,
    \new_[52743]_ , \new_[52744]_ , \new_[52748]_ , \new_[52749]_ ,
    \new_[52752]_ , \new_[52755]_ , \new_[52756]_ , \new_[52757]_ ,
    \new_[52760]_ , \new_[52763]_ , \new_[52764]_ , \new_[52767]_ ,
    \new_[52770]_ , \new_[52771]_ , \new_[52772]_ , \new_[52776]_ ,
    \new_[52777]_ , \new_[52780]_ , \new_[52783]_ , \new_[52784]_ ,
    \new_[52785]_ , \new_[52788]_ , \new_[52791]_ , \new_[52792]_ ,
    \new_[52795]_ , \new_[52798]_ , \new_[52799]_ , \new_[52800]_ ,
    \new_[52804]_ , \new_[52805]_ , \new_[52808]_ , \new_[52811]_ ,
    \new_[52812]_ , \new_[52813]_ , \new_[52816]_ , \new_[52819]_ ,
    \new_[52820]_ , \new_[52823]_ , \new_[52826]_ , \new_[52827]_ ,
    \new_[52828]_ , \new_[52832]_ , \new_[52833]_ , \new_[52836]_ ,
    \new_[52839]_ , \new_[52840]_ , \new_[52841]_ , \new_[52844]_ ,
    \new_[52847]_ , \new_[52848]_ , \new_[52851]_ , \new_[52854]_ ,
    \new_[52855]_ , \new_[52856]_ , \new_[52860]_ , \new_[52861]_ ,
    \new_[52864]_ , \new_[52867]_ , \new_[52868]_ , \new_[52869]_ ,
    \new_[52872]_ , \new_[52875]_ , \new_[52876]_ , \new_[52879]_ ,
    \new_[52882]_ , \new_[52883]_ , \new_[52884]_ , \new_[52888]_ ,
    \new_[52889]_ , \new_[52892]_ , \new_[52895]_ , \new_[52896]_ ,
    \new_[52897]_ , \new_[52900]_ , \new_[52903]_ , \new_[52904]_ ,
    \new_[52907]_ , \new_[52910]_ , \new_[52911]_ , \new_[52912]_ ,
    \new_[52916]_ , \new_[52917]_ , \new_[52920]_ , \new_[52923]_ ,
    \new_[52924]_ , \new_[52925]_ , \new_[52928]_ , \new_[52931]_ ,
    \new_[52932]_ , \new_[52935]_ , \new_[52938]_ , \new_[52939]_ ,
    \new_[52940]_ , \new_[52944]_ , \new_[52945]_ , \new_[52948]_ ,
    \new_[52951]_ , \new_[52952]_ , \new_[52953]_ , \new_[52956]_ ,
    \new_[52959]_ , \new_[52960]_ , \new_[52963]_ , \new_[52966]_ ,
    \new_[52967]_ , \new_[52968]_ , \new_[52972]_ , \new_[52973]_ ,
    \new_[52976]_ , \new_[52979]_ , \new_[52980]_ , \new_[52981]_ ,
    \new_[52984]_ , \new_[52987]_ , \new_[52988]_ , \new_[52991]_ ,
    \new_[52994]_ , \new_[52995]_ , \new_[52996]_ , \new_[53000]_ ,
    \new_[53001]_ , \new_[53004]_ , \new_[53007]_ , \new_[53008]_ ,
    \new_[53009]_ , \new_[53012]_ , \new_[53015]_ , \new_[53016]_ ,
    \new_[53019]_ , \new_[53022]_ , \new_[53023]_ , \new_[53024]_ ,
    \new_[53028]_ , \new_[53029]_ , \new_[53032]_ , \new_[53035]_ ,
    \new_[53036]_ , \new_[53037]_ , \new_[53040]_ , \new_[53043]_ ,
    \new_[53044]_ , \new_[53047]_ , \new_[53050]_ , \new_[53051]_ ,
    \new_[53052]_ , \new_[53056]_ , \new_[53057]_ , \new_[53060]_ ,
    \new_[53063]_ , \new_[53064]_ , \new_[53065]_ , \new_[53068]_ ,
    \new_[53071]_ , \new_[53072]_ , \new_[53075]_ , \new_[53078]_ ,
    \new_[53079]_ , \new_[53080]_ , \new_[53084]_ , \new_[53085]_ ,
    \new_[53088]_ , \new_[53091]_ , \new_[53092]_ , \new_[53093]_ ,
    \new_[53096]_ , \new_[53099]_ , \new_[53100]_ , \new_[53103]_ ,
    \new_[53106]_ , \new_[53107]_ , \new_[53108]_ , \new_[53112]_ ,
    \new_[53113]_ , \new_[53116]_ , \new_[53119]_ , \new_[53120]_ ,
    \new_[53121]_ , \new_[53124]_ , \new_[53127]_ , \new_[53128]_ ,
    \new_[53131]_ , \new_[53134]_ , \new_[53135]_ , \new_[53136]_ ,
    \new_[53140]_ , \new_[53141]_ , \new_[53144]_ , \new_[53147]_ ,
    \new_[53148]_ , \new_[53149]_ , \new_[53152]_ , \new_[53155]_ ,
    \new_[53156]_ , \new_[53159]_ , \new_[53162]_ , \new_[53163]_ ,
    \new_[53164]_ , \new_[53168]_ , \new_[53169]_ , \new_[53172]_ ,
    \new_[53175]_ , \new_[53176]_ , \new_[53177]_ , \new_[53180]_ ,
    \new_[53183]_ , \new_[53184]_ , \new_[53187]_ , \new_[53190]_ ,
    \new_[53191]_ , \new_[53192]_ , \new_[53196]_ , \new_[53197]_ ,
    \new_[53200]_ , \new_[53203]_ , \new_[53204]_ , \new_[53205]_ ,
    \new_[53208]_ , \new_[53211]_ , \new_[53212]_ , \new_[53215]_ ,
    \new_[53218]_ , \new_[53219]_ , \new_[53220]_ , \new_[53224]_ ,
    \new_[53225]_ , \new_[53228]_ , \new_[53231]_ , \new_[53232]_ ,
    \new_[53233]_ , \new_[53236]_ , \new_[53239]_ , \new_[53240]_ ,
    \new_[53243]_ , \new_[53246]_ , \new_[53247]_ , \new_[53248]_ ,
    \new_[53252]_ , \new_[53253]_ , \new_[53256]_ , \new_[53259]_ ,
    \new_[53260]_ , \new_[53261]_ , \new_[53264]_ , \new_[53267]_ ,
    \new_[53268]_ , \new_[53271]_ , \new_[53274]_ , \new_[53275]_ ,
    \new_[53276]_ , \new_[53280]_ , \new_[53281]_ , \new_[53284]_ ,
    \new_[53287]_ , \new_[53288]_ , \new_[53289]_ , \new_[53292]_ ,
    \new_[53295]_ , \new_[53296]_ , \new_[53299]_ , \new_[53302]_ ,
    \new_[53303]_ , \new_[53304]_ , \new_[53308]_ , \new_[53309]_ ,
    \new_[53312]_ , \new_[53315]_ , \new_[53316]_ , \new_[53317]_ ,
    \new_[53320]_ , \new_[53323]_ , \new_[53324]_ , \new_[53327]_ ,
    \new_[53330]_ , \new_[53331]_ , \new_[53332]_ , \new_[53336]_ ,
    \new_[53337]_ , \new_[53340]_ , \new_[53343]_ , \new_[53344]_ ,
    \new_[53345]_ , \new_[53348]_ , \new_[53351]_ , \new_[53352]_ ,
    \new_[53355]_ , \new_[53358]_ , \new_[53359]_ , \new_[53360]_ ,
    \new_[53364]_ , \new_[53365]_ , \new_[53368]_ , \new_[53371]_ ,
    \new_[53372]_ , \new_[53373]_ , \new_[53376]_ , \new_[53379]_ ,
    \new_[53380]_ , \new_[53383]_ , \new_[53386]_ , \new_[53387]_ ,
    \new_[53388]_ , \new_[53392]_ , \new_[53393]_ , \new_[53396]_ ,
    \new_[53399]_ , \new_[53400]_ , \new_[53401]_ , \new_[53404]_ ,
    \new_[53407]_ , \new_[53408]_ , \new_[53411]_ , \new_[53414]_ ,
    \new_[53415]_ , \new_[53416]_ , \new_[53420]_ , \new_[53421]_ ,
    \new_[53424]_ , \new_[53427]_ , \new_[53428]_ , \new_[53429]_ ,
    \new_[53432]_ , \new_[53435]_ , \new_[53436]_ , \new_[53439]_ ,
    \new_[53442]_ , \new_[53443]_ , \new_[53444]_ , \new_[53448]_ ,
    \new_[53449]_ , \new_[53452]_ , \new_[53455]_ , \new_[53456]_ ,
    \new_[53457]_ , \new_[53460]_ , \new_[53463]_ , \new_[53464]_ ,
    \new_[53467]_ , \new_[53470]_ , \new_[53471]_ , \new_[53472]_ ,
    \new_[53476]_ , \new_[53477]_ , \new_[53480]_ , \new_[53483]_ ,
    \new_[53484]_ , \new_[53485]_ , \new_[53488]_ , \new_[53491]_ ,
    \new_[53492]_ , \new_[53495]_ , \new_[53498]_ , \new_[53499]_ ,
    \new_[53500]_ , \new_[53504]_ , \new_[53505]_ , \new_[53508]_ ,
    \new_[53511]_ , \new_[53512]_ , \new_[53513]_ , \new_[53516]_ ,
    \new_[53519]_ , \new_[53520]_ , \new_[53523]_ , \new_[53526]_ ,
    \new_[53527]_ , \new_[53528]_ , \new_[53532]_ , \new_[53533]_ ,
    \new_[53536]_ , \new_[53539]_ , \new_[53540]_ , \new_[53541]_ ,
    \new_[53544]_ , \new_[53547]_ , \new_[53548]_ , \new_[53551]_ ,
    \new_[53554]_ , \new_[53555]_ , \new_[53556]_ , \new_[53560]_ ,
    \new_[53561]_ , \new_[53564]_ , \new_[53567]_ , \new_[53568]_ ,
    \new_[53569]_ , \new_[53572]_ , \new_[53575]_ , \new_[53576]_ ,
    \new_[53579]_ , \new_[53582]_ , \new_[53583]_ , \new_[53584]_ ,
    \new_[53588]_ , \new_[53589]_ , \new_[53592]_ , \new_[53595]_ ,
    \new_[53596]_ , \new_[53597]_ , \new_[53600]_ , \new_[53603]_ ,
    \new_[53604]_ , \new_[53607]_ , \new_[53610]_ , \new_[53611]_ ,
    \new_[53612]_ , \new_[53616]_ , \new_[53617]_ , \new_[53620]_ ,
    \new_[53623]_ , \new_[53624]_ , \new_[53625]_ , \new_[53628]_ ,
    \new_[53631]_ , \new_[53632]_ , \new_[53635]_ , \new_[53638]_ ,
    \new_[53639]_ , \new_[53640]_ , \new_[53644]_ , \new_[53645]_ ,
    \new_[53648]_ , \new_[53651]_ , \new_[53652]_ , \new_[53653]_ ,
    \new_[53656]_ , \new_[53659]_ , \new_[53660]_ , \new_[53663]_ ,
    \new_[53666]_ , \new_[53667]_ , \new_[53668]_ , \new_[53672]_ ,
    \new_[53673]_ , \new_[53676]_ , \new_[53679]_ , \new_[53680]_ ,
    \new_[53681]_ , \new_[53684]_ , \new_[53687]_ , \new_[53688]_ ,
    \new_[53691]_ , \new_[53694]_ , \new_[53695]_ , \new_[53696]_ ,
    \new_[53700]_ , \new_[53701]_ , \new_[53704]_ , \new_[53707]_ ,
    \new_[53708]_ , \new_[53709]_ , \new_[53712]_ , \new_[53715]_ ,
    \new_[53716]_ , \new_[53719]_ , \new_[53722]_ , \new_[53723]_ ,
    \new_[53724]_ , \new_[53728]_ , \new_[53729]_ , \new_[53732]_ ,
    \new_[53735]_ , \new_[53736]_ , \new_[53737]_ , \new_[53740]_ ,
    \new_[53743]_ , \new_[53744]_ , \new_[53747]_ , \new_[53750]_ ,
    \new_[53751]_ , \new_[53752]_ , \new_[53756]_ , \new_[53757]_ ,
    \new_[53760]_ , \new_[53763]_ , \new_[53764]_ , \new_[53765]_ ,
    \new_[53768]_ , \new_[53771]_ , \new_[53772]_ , \new_[53775]_ ,
    \new_[53778]_ , \new_[53779]_ , \new_[53780]_ , \new_[53784]_ ,
    \new_[53785]_ , \new_[53788]_ , \new_[53791]_ , \new_[53792]_ ,
    \new_[53793]_ , \new_[53796]_ , \new_[53799]_ , \new_[53800]_ ,
    \new_[53803]_ , \new_[53806]_ , \new_[53807]_ , \new_[53808]_ ,
    \new_[53812]_ , \new_[53813]_ , \new_[53816]_ , \new_[53819]_ ,
    \new_[53820]_ , \new_[53821]_ , \new_[53824]_ , \new_[53827]_ ,
    \new_[53828]_ , \new_[53831]_ , \new_[53834]_ , \new_[53835]_ ,
    \new_[53836]_ , \new_[53840]_ , \new_[53841]_ , \new_[53844]_ ,
    \new_[53847]_ , \new_[53848]_ , \new_[53849]_ , \new_[53852]_ ,
    \new_[53855]_ , \new_[53856]_ , \new_[53859]_ , \new_[53862]_ ,
    \new_[53863]_ , \new_[53864]_ , \new_[53868]_ , \new_[53869]_ ,
    \new_[53872]_ , \new_[53875]_ , \new_[53876]_ , \new_[53877]_ ,
    \new_[53880]_ , \new_[53883]_ , \new_[53884]_ , \new_[53887]_ ,
    \new_[53890]_ , \new_[53891]_ , \new_[53892]_ , \new_[53896]_ ,
    \new_[53897]_ , \new_[53900]_ , \new_[53903]_ , \new_[53904]_ ,
    \new_[53905]_ , \new_[53908]_ , \new_[53911]_ , \new_[53912]_ ,
    \new_[53915]_ , \new_[53918]_ , \new_[53919]_ , \new_[53920]_ ,
    \new_[53924]_ , \new_[53925]_ , \new_[53928]_ , \new_[53931]_ ,
    \new_[53932]_ , \new_[53933]_ , \new_[53936]_ , \new_[53939]_ ,
    \new_[53940]_ , \new_[53943]_ , \new_[53946]_ , \new_[53947]_ ,
    \new_[53948]_ , \new_[53952]_ , \new_[53953]_ , \new_[53956]_ ,
    \new_[53959]_ , \new_[53960]_ , \new_[53961]_ , \new_[53964]_ ,
    \new_[53967]_ , \new_[53968]_ , \new_[53971]_ , \new_[53974]_ ,
    \new_[53975]_ , \new_[53976]_ , \new_[53980]_ , \new_[53981]_ ,
    \new_[53984]_ , \new_[53987]_ , \new_[53988]_ , \new_[53989]_ ,
    \new_[53992]_ , \new_[53995]_ , \new_[53996]_ , \new_[53999]_ ,
    \new_[54002]_ , \new_[54003]_ , \new_[54004]_ , \new_[54008]_ ,
    \new_[54009]_ , \new_[54012]_ , \new_[54015]_ , \new_[54016]_ ,
    \new_[54017]_ , \new_[54020]_ , \new_[54023]_ , \new_[54024]_ ,
    \new_[54027]_ , \new_[54030]_ , \new_[54031]_ , \new_[54032]_ ,
    \new_[54036]_ , \new_[54037]_ , \new_[54040]_ , \new_[54043]_ ,
    \new_[54044]_ , \new_[54045]_ , \new_[54048]_ , \new_[54051]_ ,
    \new_[54052]_ , \new_[54055]_ , \new_[54058]_ , \new_[54059]_ ,
    \new_[54060]_ , \new_[54064]_ , \new_[54065]_ , \new_[54068]_ ,
    \new_[54071]_ , \new_[54072]_ , \new_[54073]_ , \new_[54076]_ ,
    \new_[54079]_ , \new_[54080]_ , \new_[54083]_ , \new_[54086]_ ,
    \new_[54087]_ , \new_[54088]_ , \new_[54092]_ , \new_[54093]_ ,
    \new_[54096]_ , \new_[54099]_ , \new_[54100]_ , \new_[54101]_ ,
    \new_[54104]_ , \new_[54107]_ , \new_[54108]_ , \new_[54111]_ ,
    \new_[54114]_ , \new_[54115]_ , \new_[54116]_ , \new_[54120]_ ,
    \new_[54121]_ , \new_[54124]_ , \new_[54127]_ , \new_[54128]_ ,
    \new_[54129]_ , \new_[54132]_ , \new_[54135]_ , \new_[54136]_ ,
    \new_[54139]_ , \new_[54142]_ , \new_[54143]_ , \new_[54144]_ ,
    \new_[54148]_ , \new_[54149]_ , \new_[54152]_ , \new_[54155]_ ,
    \new_[54156]_ , \new_[54157]_ , \new_[54160]_ , \new_[54163]_ ,
    \new_[54164]_ , \new_[54167]_ , \new_[54170]_ , \new_[54171]_ ,
    \new_[54172]_ , \new_[54176]_ , \new_[54177]_ , \new_[54180]_ ,
    \new_[54183]_ , \new_[54184]_ , \new_[54185]_ , \new_[54188]_ ,
    \new_[54191]_ , \new_[54192]_ , \new_[54195]_ , \new_[54198]_ ,
    \new_[54199]_ , \new_[54200]_ , \new_[54204]_ , \new_[54205]_ ,
    \new_[54208]_ , \new_[54211]_ , \new_[54212]_ , \new_[54213]_ ,
    \new_[54216]_ , \new_[54219]_ , \new_[54220]_ , \new_[54223]_ ,
    \new_[54226]_ , \new_[54227]_ , \new_[54228]_ , \new_[54232]_ ,
    \new_[54233]_ , \new_[54236]_ , \new_[54239]_ , \new_[54240]_ ,
    \new_[54241]_ , \new_[54244]_ , \new_[54247]_ , \new_[54248]_ ,
    \new_[54251]_ , \new_[54254]_ , \new_[54255]_ , \new_[54256]_ ,
    \new_[54260]_ , \new_[54261]_ , \new_[54264]_ , \new_[54267]_ ,
    \new_[54268]_ , \new_[54269]_ , \new_[54272]_ , \new_[54275]_ ,
    \new_[54276]_ , \new_[54279]_ , \new_[54282]_ , \new_[54283]_ ,
    \new_[54284]_ , \new_[54288]_ , \new_[54289]_ , \new_[54292]_ ,
    \new_[54295]_ , \new_[54296]_ , \new_[54297]_ , \new_[54300]_ ,
    \new_[54303]_ , \new_[54304]_ , \new_[54307]_ , \new_[54310]_ ,
    \new_[54311]_ , \new_[54312]_ , \new_[54316]_ , \new_[54317]_ ,
    \new_[54320]_ , \new_[54323]_ , \new_[54324]_ , \new_[54325]_ ,
    \new_[54328]_ , \new_[54331]_ , \new_[54332]_ , \new_[54335]_ ,
    \new_[54338]_ , \new_[54339]_ , \new_[54340]_ , \new_[54344]_ ,
    \new_[54345]_ , \new_[54348]_ , \new_[54351]_ , \new_[54352]_ ,
    \new_[54353]_ , \new_[54356]_ , \new_[54359]_ , \new_[54360]_ ,
    \new_[54363]_ , \new_[54366]_ , \new_[54367]_ , \new_[54368]_ ,
    \new_[54372]_ , \new_[54373]_ , \new_[54376]_ , \new_[54379]_ ,
    \new_[54380]_ , \new_[54381]_ , \new_[54384]_ , \new_[54387]_ ,
    \new_[54388]_ , \new_[54391]_ , \new_[54394]_ , \new_[54395]_ ,
    \new_[54396]_ , \new_[54400]_ , \new_[54401]_ , \new_[54404]_ ,
    \new_[54407]_ , \new_[54408]_ , \new_[54409]_ , \new_[54412]_ ,
    \new_[54415]_ , \new_[54416]_ , \new_[54419]_ , \new_[54422]_ ,
    \new_[54423]_ , \new_[54424]_ , \new_[54428]_ , \new_[54429]_ ,
    \new_[54432]_ , \new_[54435]_ , \new_[54436]_ , \new_[54437]_ ,
    \new_[54440]_ , \new_[54443]_ , \new_[54444]_ , \new_[54447]_ ,
    \new_[54450]_ , \new_[54451]_ , \new_[54452]_ , \new_[54456]_ ,
    \new_[54457]_ , \new_[54460]_ , \new_[54463]_ , \new_[54464]_ ,
    \new_[54465]_ , \new_[54468]_ , \new_[54471]_ , \new_[54472]_ ,
    \new_[54475]_ , \new_[54478]_ , \new_[54479]_ , \new_[54480]_ ,
    \new_[54484]_ , \new_[54485]_ , \new_[54488]_ , \new_[54491]_ ,
    \new_[54492]_ , \new_[54493]_ , \new_[54496]_ , \new_[54499]_ ,
    \new_[54500]_ , \new_[54503]_ , \new_[54506]_ , \new_[54507]_ ,
    \new_[54508]_ , \new_[54512]_ , \new_[54513]_ , \new_[54516]_ ,
    \new_[54519]_ , \new_[54520]_ , \new_[54521]_ , \new_[54524]_ ,
    \new_[54527]_ , \new_[54528]_ , \new_[54531]_ , \new_[54534]_ ,
    \new_[54535]_ , \new_[54536]_ , \new_[54540]_ , \new_[54541]_ ,
    \new_[54544]_ , \new_[54547]_ , \new_[54548]_ , \new_[54549]_ ,
    \new_[54552]_ , \new_[54555]_ , \new_[54556]_ , \new_[54559]_ ,
    \new_[54562]_ , \new_[54563]_ , \new_[54564]_ , \new_[54568]_ ,
    \new_[54569]_ , \new_[54572]_ , \new_[54575]_ , \new_[54576]_ ,
    \new_[54577]_ , \new_[54580]_ , \new_[54583]_ , \new_[54584]_ ,
    \new_[54587]_ , \new_[54590]_ , \new_[54591]_ , \new_[54592]_ ,
    \new_[54596]_ , \new_[54597]_ , \new_[54600]_ , \new_[54603]_ ,
    \new_[54604]_ , \new_[54605]_ , \new_[54608]_ , \new_[54611]_ ,
    \new_[54612]_ , \new_[54615]_ , \new_[54618]_ , \new_[54619]_ ,
    \new_[54620]_ , \new_[54624]_ , \new_[54625]_ , \new_[54628]_ ,
    \new_[54631]_ , \new_[54632]_ , \new_[54633]_ , \new_[54636]_ ,
    \new_[54639]_ , \new_[54640]_ , \new_[54643]_ , \new_[54646]_ ,
    \new_[54647]_ , \new_[54648]_ , \new_[54652]_ , \new_[54653]_ ,
    \new_[54656]_ , \new_[54659]_ , \new_[54660]_ , \new_[54661]_ ,
    \new_[54664]_ , \new_[54667]_ , \new_[54668]_ , \new_[54671]_ ,
    \new_[54674]_ , \new_[54675]_ , \new_[54676]_ , \new_[54680]_ ,
    \new_[54681]_ , \new_[54684]_ , \new_[54687]_ , \new_[54688]_ ,
    \new_[54689]_ , \new_[54692]_ , \new_[54695]_ , \new_[54696]_ ,
    \new_[54699]_ , \new_[54702]_ , \new_[54703]_ , \new_[54704]_ ,
    \new_[54708]_ , \new_[54709]_ , \new_[54712]_ , \new_[54715]_ ,
    \new_[54716]_ , \new_[54717]_ , \new_[54720]_ , \new_[54723]_ ,
    \new_[54724]_ , \new_[54727]_ , \new_[54730]_ , \new_[54731]_ ,
    \new_[54732]_ , \new_[54736]_ , \new_[54737]_ , \new_[54740]_ ,
    \new_[54743]_ , \new_[54744]_ , \new_[54745]_ , \new_[54748]_ ,
    \new_[54751]_ , \new_[54752]_ , \new_[54755]_ , \new_[54758]_ ,
    \new_[54759]_ , \new_[54760]_ , \new_[54764]_ , \new_[54765]_ ,
    \new_[54768]_ , \new_[54771]_ , \new_[54772]_ , \new_[54773]_ ,
    \new_[54776]_ , \new_[54779]_ , \new_[54780]_ , \new_[54783]_ ,
    \new_[54786]_ , \new_[54787]_ , \new_[54788]_ , \new_[54792]_ ,
    \new_[54793]_ , \new_[54796]_ , \new_[54799]_ , \new_[54800]_ ,
    \new_[54801]_ , \new_[54804]_ , \new_[54807]_ , \new_[54808]_ ,
    \new_[54811]_ , \new_[54814]_ , \new_[54815]_ , \new_[54816]_ ,
    \new_[54820]_ , \new_[54821]_ , \new_[54824]_ , \new_[54827]_ ,
    \new_[54828]_ , \new_[54829]_ , \new_[54832]_ , \new_[54835]_ ,
    \new_[54836]_ , \new_[54839]_ , \new_[54842]_ , \new_[54843]_ ,
    \new_[54844]_ , \new_[54848]_ , \new_[54849]_ , \new_[54852]_ ,
    \new_[54855]_ , \new_[54856]_ , \new_[54857]_ , \new_[54860]_ ,
    \new_[54863]_ , \new_[54864]_ , \new_[54867]_ , \new_[54870]_ ,
    \new_[54871]_ , \new_[54872]_ , \new_[54876]_ , \new_[54877]_ ,
    \new_[54880]_ , \new_[54883]_ , \new_[54884]_ , \new_[54885]_ ,
    \new_[54888]_ , \new_[54891]_ , \new_[54892]_ , \new_[54895]_ ,
    \new_[54898]_ , \new_[54899]_ , \new_[54900]_ , \new_[54904]_ ,
    \new_[54905]_ , \new_[54908]_ , \new_[54911]_ , \new_[54912]_ ,
    \new_[54913]_ , \new_[54916]_ , \new_[54919]_ , \new_[54920]_ ,
    \new_[54923]_ , \new_[54926]_ , \new_[54927]_ , \new_[54928]_ ,
    \new_[54932]_ , \new_[54933]_ , \new_[54936]_ , \new_[54939]_ ,
    \new_[54940]_ , \new_[54941]_ , \new_[54944]_ , \new_[54947]_ ,
    \new_[54948]_ , \new_[54951]_ , \new_[54954]_ , \new_[54955]_ ,
    \new_[54956]_ , \new_[54960]_ , \new_[54961]_ , \new_[54964]_ ,
    \new_[54967]_ , \new_[54968]_ , \new_[54969]_ , \new_[54972]_ ,
    \new_[54975]_ , \new_[54976]_ , \new_[54979]_ , \new_[54982]_ ,
    \new_[54983]_ , \new_[54984]_ , \new_[54988]_ , \new_[54989]_ ,
    \new_[54992]_ , \new_[54995]_ , \new_[54996]_ , \new_[54997]_ ,
    \new_[55000]_ , \new_[55003]_ , \new_[55004]_ , \new_[55007]_ ,
    \new_[55010]_ , \new_[55011]_ , \new_[55012]_ , \new_[55016]_ ,
    \new_[55017]_ , \new_[55020]_ , \new_[55023]_ , \new_[55024]_ ,
    \new_[55025]_ , \new_[55028]_ , \new_[55031]_ , \new_[55032]_ ,
    \new_[55035]_ , \new_[55038]_ , \new_[55039]_ , \new_[55040]_ ,
    \new_[55044]_ , \new_[55045]_ , \new_[55048]_ , \new_[55051]_ ,
    \new_[55052]_ , \new_[55053]_ , \new_[55056]_ , \new_[55059]_ ,
    \new_[55060]_ , \new_[55063]_ , \new_[55066]_ , \new_[55067]_ ,
    \new_[55068]_ , \new_[55072]_ , \new_[55073]_ , \new_[55076]_ ,
    \new_[55079]_ , \new_[55080]_ , \new_[55081]_ , \new_[55084]_ ,
    \new_[55087]_ , \new_[55088]_ , \new_[55091]_ , \new_[55094]_ ,
    \new_[55095]_ , \new_[55096]_ , \new_[55100]_ , \new_[55101]_ ,
    \new_[55104]_ , \new_[55107]_ , \new_[55108]_ , \new_[55109]_ ,
    \new_[55112]_ , \new_[55115]_ , \new_[55116]_ , \new_[55119]_ ,
    \new_[55122]_ , \new_[55123]_ , \new_[55124]_ , \new_[55128]_ ,
    \new_[55129]_ , \new_[55132]_ , \new_[55135]_ , \new_[55136]_ ,
    \new_[55137]_ , \new_[55140]_ , \new_[55143]_ , \new_[55144]_ ,
    \new_[55147]_ , \new_[55150]_ , \new_[55151]_ , \new_[55152]_ ,
    \new_[55156]_ , \new_[55157]_ , \new_[55160]_ , \new_[55163]_ ,
    \new_[55164]_ , \new_[55165]_ , \new_[55168]_ , \new_[55171]_ ,
    \new_[55172]_ , \new_[55175]_ , \new_[55178]_ , \new_[55179]_ ,
    \new_[55180]_ , \new_[55184]_ , \new_[55185]_ , \new_[55188]_ ,
    \new_[55191]_ , \new_[55192]_ , \new_[55193]_ , \new_[55196]_ ,
    \new_[55199]_ , \new_[55200]_ , \new_[55203]_ , \new_[55206]_ ,
    \new_[55207]_ , \new_[55208]_ , \new_[55212]_ , \new_[55213]_ ,
    \new_[55216]_ , \new_[55219]_ , \new_[55220]_ , \new_[55221]_ ,
    \new_[55224]_ , \new_[55227]_ , \new_[55228]_ , \new_[55231]_ ,
    \new_[55234]_ , \new_[55235]_ , \new_[55236]_ , \new_[55240]_ ,
    \new_[55241]_ , \new_[55244]_ , \new_[55247]_ , \new_[55248]_ ,
    \new_[55249]_ , \new_[55252]_ , \new_[55255]_ , \new_[55256]_ ,
    \new_[55259]_ , \new_[55262]_ , \new_[55263]_ , \new_[55264]_ ,
    \new_[55268]_ , \new_[55269]_ , \new_[55272]_ , \new_[55275]_ ,
    \new_[55276]_ , \new_[55277]_ , \new_[55280]_ , \new_[55283]_ ,
    \new_[55284]_ , \new_[55287]_ , \new_[55290]_ , \new_[55291]_ ,
    \new_[55292]_ , \new_[55296]_ , \new_[55297]_ , \new_[55300]_ ,
    \new_[55303]_ , \new_[55304]_ , \new_[55305]_ , \new_[55308]_ ,
    \new_[55311]_ , \new_[55312]_ , \new_[55315]_ , \new_[55318]_ ,
    \new_[55319]_ , \new_[55320]_ , \new_[55324]_ , \new_[55325]_ ,
    \new_[55328]_ , \new_[55331]_ , \new_[55332]_ , \new_[55333]_ ,
    \new_[55336]_ , \new_[55339]_ , \new_[55340]_ , \new_[55343]_ ,
    \new_[55346]_ , \new_[55347]_ , \new_[55348]_ , \new_[55352]_ ,
    \new_[55353]_ , \new_[55356]_ , \new_[55359]_ , \new_[55360]_ ,
    \new_[55361]_ , \new_[55364]_ , \new_[55367]_ , \new_[55368]_ ,
    \new_[55371]_ , \new_[55374]_ , \new_[55375]_ , \new_[55376]_ ,
    \new_[55380]_ , \new_[55381]_ , \new_[55384]_ , \new_[55387]_ ,
    \new_[55388]_ , \new_[55389]_ , \new_[55392]_ , \new_[55395]_ ,
    \new_[55396]_ , \new_[55399]_ , \new_[55402]_ , \new_[55403]_ ,
    \new_[55404]_ , \new_[55408]_ , \new_[55409]_ , \new_[55412]_ ,
    \new_[55415]_ , \new_[55416]_ , \new_[55417]_ , \new_[55420]_ ,
    \new_[55423]_ , \new_[55424]_ , \new_[55427]_ , \new_[55430]_ ,
    \new_[55431]_ , \new_[55432]_ , \new_[55436]_ , \new_[55437]_ ,
    \new_[55440]_ , \new_[55443]_ , \new_[55444]_ , \new_[55445]_ ,
    \new_[55448]_ , \new_[55451]_ , \new_[55452]_ , \new_[55455]_ ,
    \new_[55458]_ , \new_[55459]_ , \new_[55460]_ , \new_[55464]_ ,
    \new_[55465]_ , \new_[55468]_ , \new_[55471]_ , \new_[55472]_ ,
    \new_[55473]_ , \new_[55476]_ , \new_[55479]_ , \new_[55480]_ ,
    \new_[55483]_ , \new_[55486]_ , \new_[55487]_ , \new_[55488]_ ,
    \new_[55492]_ , \new_[55493]_ , \new_[55496]_ , \new_[55499]_ ,
    \new_[55500]_ , \new_[55501]_ , \new_[55504]_ , \new_[55507]_ ,
    \new_[55508]_ , \new_[55511]_ , \new_[55514]_ , \new_[55515]_ ,
    \new_[55516]_ , \new_[55520]_ , \new_[55521]_ , \new_[55524]_ ,
    \new_[55527]_ , \new_[55528]_ , \new_[55529]_ , \new_[55532]_ ,
    \new_[55535]_ , \new_[55536]_ , \new_[55539]_ , \new_[55542]_ ,
    \new_[55543]_ , \new_[55544]_ , \new_[55548]_ , \new_[55549]_ ,
    \new_[55552]_ , \new_[55555]_ , \new_[55556]_ , \new_[55557]_ ,
    \new_[55560]_ , \new_[55563]_ , \new_[55564]_ , \new_[55567]_ ,
    \new_[55570]_ , \new_[55571]_ , \new_[55572]_ , \new_[55576]_ ,
    \new_[55577]_ , \new_[55580]_ , \new_[55583]_ , \new_[55584]_ ,
    \new_[55585]_ , \new_[55588]_ , \new_[55591]_ , \new_[55592]_ ,
    \new_[55595]_ , \new_[55598]_ , \new_[55599]_ , \new_[55600]_ ,
    \new_[55604]_ , \new_[55605]_ , \new_[55608]_ , \new_[55611]_ ,
    \new_[55612]_ , \new_[55613]_ , \new_[55616]_ , \new_[55619]_ ,
    \new_[55620]_ , \new_[55623]_ , \new_[55626]_ , \new_[55627]_ ,
    \new_[55628]_ , \new_[55632]_ , \new_[55633]_ , \new_[55636]_ ,
    \new_[55639]_ , \new_[55640]_ , \new_[55641]_ , \new_[55644]_ ,
    \new_[55647]_ , \new_[55648]_ , \new_[55651]_ , \new_[55654]_ ,
    \new_[55655]_ , \new_[55656]_ , \new_[55660]_ , \new_[55661]_ ,
    \new_[55664]_ , \new_[55667]_ , \new_[55668]_ , \new_[55669]_ ,
    \new_[55672]_ , \new_[55675]_ , \new_[55676]_ , \new_[55679]_ ,
    \new_[55682]_ , \new_[55683]_ , \new_[55684]_ , \new_[55688]_ ,
    \new_[55689]_ , \new_[55692]_ , \new_[55695]_ , \new_[55696]_ ,
    \new_[55697]_ , \new_[55700]_ , \new_[55703]_ , \new_[55704]_ ,
    \new_[55707]_ , \new_[55710]_ , \new_[55711]_ , \new_[55712]_ ,
    \new_[55716]_ , \new_[55717]_ , \new_[55720]_ , \new_[55723]_ ,
    \new_[55724]_ , \new_[55725]_ , \new_[55728]_ , \new_[55731]_ ,
    \new_[55732]_ , \new_[55735]_ , \new_[55738]_ , \new_[55739]_ ,
    \new_[55740]_ , \new_[55744]_ , \new_[55745]_ , \new_[55748]_ ,
    \new_[55751]_ , \new_[55752]_ , \new_[55753]_ , \new_[55756]_ ,
    \new_[55759]_ , \new_[55760]_ , \new_[55763]_ , \new_[55766]_ ,
    \new_[55767]_ , \new_[55768]_ , \new_[55772]_ , \new_[55773]_ ,
    \new_[55776]_ , \new_[55779]_ , \new_[55780]_ , \new_[55781]_ ,
    \new_[55784]_ , \new_[55787]_ , \new_[55788]_ , \new_[55791]_ ,
    \new_[55794]_ , \new_[55795]_ , \new_[55796]_ , \new_[55800]_ ,
    \new_[55801]_ , \new_[55804]_ , \new_[55807]_ , \new_[55808]_ ,
    \new_[55809]_ , \new_[55812]_ , \new_[55815]_ , \new_[55816]_ ,
    \new_[55819]_ , \new_[55822]_ , \new_[55823]_ , \new_[55824]_ ,
    \new_[55828]_ , \new_[55829]_ , \new_[55832]_ , \new_[55835]_ ,
    \new_[55836]_ , \new_[55837]_ , \new_[55840]_ , \new_[55843]_ ,
    \new_[55844]_ , \new_[55847]_ , \new_[55850]_ , \new_[55851]_ ,
    \new_[55852]_ , \new_[55856]_ , \new_[55857]_ , \new_[55860]_ ,
    \new_[55863]_ , \new_[55864]_ , \new_[55865]_ , \new_[55868]_ ,
    \new_[55871]_ , \new_[55872]_ , \new_[55875]_ , \new_[55878]_ ,
    \new_[55879]_ , \new_[55880]_ , \new_[55884]_ , \new_[55885]_ ,
    \new_[55888]_ , \new_[55891]_ , \new_[55892]_ , \new_[55893]_ ,
    \new_[55896]_ , \new_[55899]_ , \new_[55900]_ , \new_[55903]_ ,
    \new_[55906]_ , \new_[55907]_ , \new_[55908]_ , \new_[55912]_ ,
    \new_[55913]_ , \new_[55916]_ , \new_[55919]_ , \new_[55920]_ ,
    \new_[55921]_ , \new_[55924]_ , \new_[55927]_ , \new_[55928]_ ,
    \new_[55931]_ , \new_[55934]_ , \new_[55935]_ , \new_[55936]_ ,
    \new_[55940]_ , \new_[55941]_ , \new_[55944]_ , \new_[55947]_ ,
    \new_[55948]_ , \new_[55949]_ , \new_[55952]_ , \new_[55955]_ ,
    \new_[55956]_ , \new_[55959]_ , \new_[55962]_ , \new_[55963]_ ,
    \new_[55964]_ , \new_[55968]_ , \new_[55969]_ , \new_[55972]_ ,
    \new_[55975]_ , \new_[55976]_ , \new_[55977]_ , \new_[55980]_ ,
    \new_[55983]_ , \new_[55984]_ , \new_[55987]_ , \new_[55990]_ ,
    \new_[55991]_ , \new_[55992]_ , \new_[55996]_ , \new_[55997]_ ,
    \new_[56000]_ , \new_[56003]_ , \new_[56004]_ , \new_[56005]_ ,
    \new_[56008]_ , \new_[56011]_ , \new_[56012]_ , \new_[56015]_ ,
    \new_[56018]_ , \new_[56019]_ , \new_[56020]_ , \new_[56024]_ ,
    \new_[56025]_ , \new_[56028]_ , \new_[56031]_ , \new_[56032]_ ,
    \new_[56033]_ , \new_[56036]_ , \new_[56039]_ , \new_[56040]_ ,
    \new_[56043]_ , \new_[56046]_ , \new_[56047]_ , \new_[56048]_ ,
    \new_[56052]_ , \new_[56053]_ , \new_[56056]_ , \new_[56059]_ ,
    \new_[56060]_ , \new_[56061]_ , \new_[56064]_ , \new_[56067]_ ,
    \new_[56068]_ , \new_[56071]_ , \new_[56074]_ , \new_[56075]_ ,
    \new_[56076]_ , \new_[56080]_ , \new_[56081]_ , \new_[56084]_ ,
    \new_[56087]_ , \new_[56088]_ , \new_[56089]_ , \new_[56092]_ ,
    \new_[56095]_ , \new_[56096]_ , \new_[56099]_ , \new_[56102]_ ,
    \new_[56103]_ , \new_[56104]_ , \new_[56108]_ , \new_[56109]_ ,
    \new_[56112]_ , \new_[56115]_ , \new_[56116]_ , \new_[56117]_ ,
    \new_[56120]_ , \new_[56123]_ , \new_[56124]_ , \new_[56127]_ ,
    \new_[56130]_ , \new_[56131]_ , \new_[56132]_ , \new_[56136]_ ,
    \new_[56137]_ , \new_[56140]_ , \new_[56143]_ , \new_[56144]_ ,
    \new_[56145]_ , \new_[56148]_ , \new_[56151]_ , \new_[56152]_ ,
    \new_[56155]_ , \new_[56158]_ , \new_[56159]_ , \new_[56160]_ ,
    \new_[56164]_ , \new_[56165]_ , \new_[56168]_ , \new_[56171]_ ,
    \new_[56172]_ , \new_[56173]_ , \new_[56176]_ , \new_[56179]_ ,
    \new_[56180]_ , \new_[56183]_ , \new_[56186]_ , \new_[56187]_ ,
    \new_[56188]_ , \new_[56192]_ , \new_[56193]_ , \new_[56196]_ ,
    \new_[56199]_ , \new_[56200]_ , \new_[56201]_ , \new_[56204]_ ,
    \new_[56207]_ , \new_[56208]_ , \new_[56211]_ , \new_[56214]_ ,
    \new_[56215]_ , \new_[56216]_ , \new_[56220]_ , \new_[56221]_ ,
    \new_[56224]_ , \new_[56227]_ , \new_[56228]_ , \new_[56229]_ ,
    \new_[56232]_ , \new_[56235]_ , \new_[56236]_ , \new_[56239]_ ,
    \new_[56242]_ , \new_[56243]_ , \new_[56244]_ , \new_[56248]_ ,
    \new_[56249]_ , \new_[56252]_ , \new_[56255]_ , \new_[56256]_ ,
    \new_[56257]_ , \new_[56260]_ , \new_[56263]_ , \new_[56264]_ ,
    \new_[56267]_ , \new_[56270]_ , \new_[56271]_ , \new_[56272]_ ,
    \new_[56276]_ , \new_[56277]_ , \new_[56280]_ , \new_[56283]_ ,
    \new_[56284]_ , \new_[56285]_ , \new_[56288]_ , \new_[56291]_ ,
    \new_[56292]_ , \new_[56295]_ , \new_[56298]_ , \new_[56299]_ ,
    \new_[56300]_ , \new_[56304]_ , \new_[56305]_ , \new_[56308]_ ,
    \new_[56311]_ , \new_[56312]_ , \new_[56313]_ , \new_[56316]_ ,
    \new_[56319]_ , \new_[56320]_ , \new_[56323]_ , \new_[56326]_ ,
    \new_[56327]_ , \new_[56328]_ , \new_[56332]_ , \new_[56333]_ ,
    \new_[56336]_ , \new_[56339]_ , \new_[56340]_ , \new_[56341]_ ,
    \new_[56344]_ , \new_[56347]_ , \new_[56348]_ , \new_[56351]_ ,
    \new_[56354]_ , \new_[56355]_ , \new_[56356]_ , \new_[56360]_ ,
    \new_[56361]_ , \new_[56364]_ , \new_[56367]_ , \new_[56368]_ ,
    \new_[56369]_ , \new_[56372]_ , \new_[56375]_ , \new_[56376]_ ,
    \new_[56379]_ , \new_[56382]_ , \new_[56383]_ , \new_[56384]_ ,
    \new_[56388]_ , \new_[56389]_ , \new_[56392]_ , \new_[56395]_ ,
    \new_[56396]_ , \new_[56397]_ , \new_[56400]_ , \new_[56403]_ ,
    \new_[56404]_ , \new_[56407]_ , \new_[56410]_ , \new_[56411]_ ,
    \new_[56412]_ , \new_[56416]_ , \new_[56417]_ , \new_[56420]_ ,
    \new_[56423]_ , \new_[56424]_ , \new_[56425]_ , \new_[56428]_ ,
    \new_[56431]_ , \new_[56432]_ , \new_[56435]_ , \new_[56438]_ ,
    \new_[56439]_ , \new_[56440]_ , \new_[56444]_ , \new_[56445]_ ,
    \new_[56448]_ , \new_[56451]_ , \new_[56452]_ , \new_[56453]_ ,
    \new_[56456]_ , \new_[56459]_ , \new_[56460]_ , \new_[56463]_ ,
    \new_[56466]_ , \new_[56467]_ , \new_[56468]_ , \new_[56472]_ ,
    \new_[56473]_ , \new_[56476]_ , \new_[56479]_ , \new_[56480]_ ,
    \new_[56481]_ , \new_[56484]_ , \new_[56487]_ , \new_[56488]_ ,
    \new_[56491]_ , \new_[56494]_ , \new_[56495]_ , \new_[56496]_ ,
    \new_[56500]_ , \new_[56501]_ , \new_[56504]_ , \new_[56507]_ ,
    \new_[56508]_ , \new_[56509]_ , \new_[56512]_ , \new_[56515]_ ,
    \new_[56516]_ , \new_[56519]_ , \new_[56522]_ , \new_[56523]_ ,
    \new_[56524]_ , \new_[56528]_ , \new_[56529]_ , \new_[56532]_ ,
    \new_[56535]_ , \new_[56536]_ , \new_[56537]_ , \new_[56540]_ ,
    \new_[56543]_ , \new_[56544]_ , \new_[56547]_ , \new_[56550]_ ,
    \new_[56551]_ , \new_[56552]_ , \new_[56556]_ , \new_[56557]_ ,
    \new_[56560]_ , \new_[56563]_ , \new_[56564]_ , \new_[56565]_ ,
    \new_[56568]_ , \new_[56571]_ , \new_[56572]_ , \new_[56575]_ ,
    \new_[56578]_ , \new_[56579]_ , \new_[56580]_ , \new_[56584]_ ,
    \new_[56585]_ , \new_[56588]_ , \new_[56591]_ , \new_[56592]_ ,
    \new_[56593]_ , \new_[56596]_ , \new_[56599]_ , \new_[56600]_ ,
    \new_[56603]_ , \new_[56606]_ , \new_[56607]_ , \new_[56608]_ ,
    \new_[56612]_ , \new_[56613]_ , \new_[56616]_ , \new_[56619]_ ,
    \new_[56620]_ , \new_[56621]_ , \new_[56624]_ , \new_[56627]_ ,
    \new_[56628]_ , \new_[56631]_ , \new_[56634]_ , \new_[56635]_ ,
    \new_[56636]_ , \new_[56640]_ , \new_[56641]_ , \new_[56644]_ ,
    \new_[56647]_ , \new_[56648]_ , \new_[56649]_ , \new_[56652]_ ,
    \new_[56655]_ , \new_[56656]_ , \new_[56659]_ , \new_[56662]_ ,
    \new_[56663]_ , \new_[56664]_ , \new_[56668]_ , \new_[56669]_ ,
    \new_[56672]_ , \new_[56675]_ , \new_[56676]_ , \new_[56677]_ ,
    \new_[56680]_ , \new_[56683]_ , \new_[56684]_ , \new_[56687]_ ,
    \new_[56690]_ , \new_[56691]_ , \new_[56692]_ , \new_[56696]_ ,
    \new_[56697]_ , \new_[56700]_ , \new_[56703]_ , \new_[56704]_ ,
    \new_[56705]_ , \new_[56708]_ , \new_[56711]_ , \new_[56712]_ ,
    \new_[56715]_ , \new_[56718]_ , \new_[56719]_ , \new_[56720]_ ,
    \new_[56724]_ , \new_[56725]_ , \new_[56728]_ , \new_[56731]_ ,
    \new_[56732]_ , \new_[56733]_ , \new_[56736]_ , \new_[56739]_ ,
    \new_[56740]_ , \new_[56743]_ , \new_[56746]_ , \new_[56747]_ ,
    \new_[56748]_ , \new_[56752]_ , \new_[56753]_ , \new_[56756]_ ,
    \new_[56759]_ , \new_[56760]_ , \new_[56761]_ , \new_[56764]_ ,
    \new_[56767]_ , \new_[56768]_ , \new_[56771]_ , \new_[56774]_ ,
    \new_[56775]_ , \new_[56776]_ , \new_[56780]_ , \new_[56781]_ ,
    \new_[56784]_ , \new_[56787]_ , \new_[56788]_ , \new_[56789]_ ,
    \new_[56792]_ , \new_[56795]_ , \new_[56796]_ , \new_[56799]_ ,
    \new_[56802]_ , \new_[56803]_ , \new_[56804]_ , \new_[56808]_ ,
    \new_[56809]_ , \new_[56812]_ , \new_[56815]_ , \new_[56816]_ ,
    \new_[56817]_ , \new_[56820]_ , \new_[56823]_ , \new_[56824]_ ,
    \new_[56827]_ , \new_[56830]_ , \new_[56831]_ , \new_[56832]_ ,
    \new_[56836]_ , \new_[56837]_ , \new_[56840]_ , \new_[56843]_ ,
    \new_[56844]_ , \new_[56845]_ , \new_[56848]_ , \new_[56851]_ ,
    \new_[56852]_ , \new_[56855]_ , \new_[56858]_ , \new_[56859]_ ,
    \new_[56860]_ , \new_[56864]_ , \new_[56865]_ , \new_[56868]_ ,
    \new_[56871]_ , \new_[56872]_ , \new_[56873]_ , \new_[56876]_ ,
    \new_[56879]_ , \new_[56880]_ , \new_[56883]_ , \new_[56886]_ ,
    \new_[56887]_ , \new_[56888]_ , \new_[56892]_ , \new_[56893]_ ,
    \new_[56896]_ , \new_[56899]_ , \new_[56900]_ , \new_[56901]_ ,
    \new_[56904]_ , \new_[56907]_ , \new_[56908]_ , \new_[56911]_ ,
    \new_[56914]_ , \new_[56915]_ , \new_[56916]_ , \new_[56920]_ ,
    \new_[56921]_ , \new_[56924]_ , \new_[56927]_ , \new_[56928]_ ,
    \new_[56929]_ , \new_[56932]_ , \new_[56935]_ , \new_[56936]_ ,
    \new_[56939]_ , \new_[56942]_ , \new_[56943]_ , \new_[56944]_ ,
    \new_[56948]_ , \new_[56949]_ , \new_[56952]_ , \new_[56955]_ ,
    \new_[56956]_ , \new_[56957]_ , \new_[56960]_ , \new_[56963]_ ,
    \new_[56964]_ , \new_[56967]_ , \new_[56970]_ , \new_[56971]_ ,
    \new_[56972]_ , \new_[56976]_ , \new_[56977]_ , \new_[56980]_ ,
    \new_[56983]_ , \new_[56984]_ , \new_[56985]_ , \new_[56988]_ ,
    \new_[56991]_ , \new_[56992]_ , \new_[56995]_ , \new_[56998]_ ,
    \new_[56999]_ , \new_[57000]_ , \new_[57004]_ , \new_[57005]_ ,
    \new_[57008]_ , \new_[57011]_ , \new_[57012]_ , \new_[57013]_ ,
    \new_[57016]_ , \new_[57019]_ , \new_[57020]_ , \new_[57023]_ ,
    \new_[57026]_ , \new_[57027]_ , \new_[57028]_ , \new_[57032]_ ,
    \new_[57033]_ , \new_[57036]_ , \new_[57039]_ , \new_[57040]_ ,
    \new_[57041]_ , \new_[57044]_ , \new_[57047]_ , \new_[57048]_ ,
    \new_[57051]_ , \new_[57054]_ , \new_[57055]_ , \new_[57056]_ ,
    \new_[57060]_ , \new_[57061]_ , \new_[57064]_ , \new_[57067]_ ,
    \new_[57068]_ , \new_[57069]_ , \new_[57072]_ , \new_[57075]_ ,
    \new_[57076]_ , \new_[57079]_ , \new_[57082]_ , \new_[57083]_ ,
    \new_[57084]_ , \new_[57088]_ , \new_[57089]_ , \new_[57092]_ ,
    \new_[57095]_ , \new_[57096]_ , \new_[57097]_ , \new_[57100]_ ,
    \new_[57103]_ , \new_[57104]_ , \new_[57107]_ , \new_[57110]_ ,
    \new_[57111]_ , \new_[57112]_ , \new_[57116]_ , \new_[57117]_ ,
    \new_[57120]_ , \new_[57123]_ , \new_[57124]_ , \new_[57125]_ ,
    \new_[57128]_ , \new_[57131]_ , \new_[57132]_ , \new_[57135]_ ,
    \new_[57138]_ , \new_[57139]_ , \new_[57140]_ , \new_[57144]_ ,
    \new_[57145]_ , \new_[57148]_ , \new_[57151]_ , \new_[57152]_ ,
    \new_[57153]_ , \new_[57156]_ , \new_[57159]_ , \new_[57160]_ ,
    \new_[57163]_ , \new_[57166]_ , \new_[57167]_ , \new_[57168]_ ,
    \new_[57172]_ , \new_[57173]_ , \new_[57176]_ , \new_[57179]_ ,
    \new_[57180]_ , \new_[57181]_ , \new_[57184]_ , \new_[57187]_ ,
    \new_[57188]_ , \new_[57191]_ , \new_[57194]_ , \new_[57195]_ ,
    \new_[57196]_ , \new_[57200]_ , \new_[57201]_ , \new_[57204]_ ,
    \new_[57207]_ , \new_[57208]_ , \new_[57209]_ , \new_[57212]_ ,
    \new_[57215]_ , \new_[57216]_ , \new_[57219]_ , \new_[57222]_ ,
    \new_[57223]_ , \new_[57224]_ , \new_[57228]_ , \new_[57229]_ ,
    \new_[57232]_ , \new_[57235]_ , \new_[57236]_ , \new_[57237]_ ,
    \new_[57240]_ , \new_[57243]_ , \new_[57244]_ , \new_[57247]_ ,
    \new_[57250]_ , \new_[57251]_ , \new_[57252]_ , \new_[57256]_ ,
    \new_[57257]_ , \new_[57260]_ , \new_[57263]_ , \new_[57264]_ ,
    \new_[57265]_ , \new_[57268]_ , \new_[57271]_ , \new_[57272]_ ,
    \new_[57275]_ , \new_[57278]_ , \new_[57279]_ , \new_[57280]_ ,
    \new_[57284]_ , \new_[57285]_ , \new_[57288]_ , \new_[57291]_ ,
    \new_[57292]_ , \new_[57293]_ , \new_[57296]_ , \new_[57299]_ ,
    \new_[57300]_ , \new_[57303]_ , \new_[57306]_ , \new_[57307]_ ,
    \new_[57308]_ , \new_[57312]_ , \new_[57313]_ , \new_[57316]_ ,
    \new_[57319]_ , \new_[57320]_ , \new_[57321]_ , \new_[57324]_ ,
    \new_[57327]_ , \new_[57328]_ , \new_[57331]_ , \new_[57334]_ ,
    \new_[57335]_ , \new_[57336]_ , \new_[57340]_ , \new_[57341]_ ,
    \new_[57344]_ , \new_[57347]_ , \new_[57348]_ , \new_[57349]_ ,
    \new_[57352]_ , \new_[57355]_ , \new_[57356]_ , \new_[57359]_ ,
    \new_[57362]_ , \new_[57363]_ , \new_[57364]_ , \new_[57368]_ ,
    \new_[57369]_ , \new_[57372]_ , \new_[57375]_ , \new_[57376]_ ,
    \new_[57377]_ , \new_[57380]_ , \new_[57383]_ , \new_[57384]_ ,
    \new_[57387]_ , \new_[57390]_ , \new_[57391]_ , \new_[57392]_ ,
    \new_[57396]_ , \new_[57397]_ , \new_[57400]_ , \new_[57403]_ ,
    \new_[57404]_ , \new_[57405]_ , \new_[57408]_ , \new_[57411]_ ,
    \new_[57412]_ , \new_[57415]_ , \new_[57418]_ , \new_[57419]_ ,
    \new_[57420]_ , \new_[57424]_ , \new_[57425]_ , \new_[57428]_ ,
    \new_[57431]_ , \new_[57432]_ , \new_[57433]_ , \new_[57436]_ ,
    \new_[57439]_ , \new_[57440]_ , \new_[57443]_ , \new_[57446]_ ,
    \new_[57447]_ , \new_[57448]_ , \new_[57452]_ , \new_[57453]_ ,
    \new_[57456]_ , \new_[57459]_ , \new_[57460]_ , \new_[57461]_ ,
    \new_[57464]_ , \new_[57467]_ , \new_[57468]_ , \new_[57471]_ ,
    \new_[57474]_ , \new_[57475]_ , \new_[57476]_ , \new_[57480]_ ,
    \new_[57481]_ , \new_[57484]_ , \new_[57487]_ , \new_[57488]_ ,
    \new_[57489]_ , \new_[57492]_ , \new_[57495]_ , \new_[57496]_ ,
    \new_[57499]_ , \new_[57502]_ , \new_[57503]_ , \new_[57504]_ ,
    \new_[57508]_ , \new_[57509]_ , \new_[57512]_ , \new_[57515]_ ,
    \new_[57516]_ , \new_[57517]_ , \new_[57520]_ , \new_[57523]_ ,
    \new_[57524]_ , \new_[57527]_ , \new_[57530]_ , \new_[57531]_ ,
    \new_[57532]_ , \new_[57536]_ , \new_[57537]_ , \new_[57540]_ ,
    \new_[57543]_ , \new_[57544]_ , \new_[57545]_ , \new_[57548]_ ,
    \new_[57551]_ , \new_[57552]_ , \new_[57555]_ , \new_[57558]_ ,
    \new_[57559]_ , \new_[57560]_ , \new_[57564]_ , \new_[57565]_ ,
    \new_[57568]_ , \new_[57571]_ , \new_[57572]_ , \new_[57573]_ ,
    \new_[57576]_ , \new_[57579]_ , \new_[57580]_ , \new_[57583]_ ,
    \new_[57586]_ , \new_[57587]_ , \new_[57588]_ , \new_[57592]_ ,
    \new_[57593]_ , \new_[57596]_ , \new_[57599]_ , \new_[57600]_ ,
    \new_[57601]_ , \new_[57604]_ , \new_[57607]_ , \new_[57608]_ ,
    \new_[57611]_ , \new_[57614]_ , \new_[57615]_ , \new_[57616]_ ,
    \new_[57620]_ , \new_[57621]_ , \new_[57624]_ , \new_[57627]_ ,
    \new_[57628]_ , \new_[57629]_ , \new_[57632]_ , \new_[57635]_ ,
    \new_[57636]_ , \new_[57639]_ , \new_[57642]_ , \new_[57643]_ ,
    \new_[57644]_ , \new_[57648]_ , \new_[57649]_ , \new_[57652]_ ,
    \new_[57655]_ , \new_[57656]_ , \new_[57657]_ , \new_[57660]_ ,
    \new_[57663]_ , \new_[57664]_ , \new_[57667]_ , \new_[57670]_ ,
    \new_[57671]_ , \new_[57672]_ , \new_[57676]_ , \new_[57677]_ ,
    \new_[57680]_ , \new_[57683]_ , \new_[57684]_ , \new_[57685]_ ,
    \new_[57688]_ , \new_[57691]_ , \new_[57692]_ , \new_[57695]_ ,
    \new_[57698]_ , \new_[57699]_ , \new_[57700]_ , \new_[57704]_ ,
    \new_[57705]_ , \new_[57708]_ , \new_[57711]_ , \new_[57712]_ ,
    \new_[57713]_ , \new_[57716]_ , \new_[57719]_ , \new_[57720]_ ,
    \new_[57723]_ , \new_[57726]_ , \new_[57727]_ , \new_[57728]_ ,
    \new_[57731]_ , \new_[57734]_ , \new_[57735]_ , \new_[57738]_ ,
    \new_[57741]_ , \new_[57742]_ , \new_[57743]_ , \new_[57746]_ ,
    \new_[57749]_ , \new_[57750]_ , \new_[57753]_ , \new_[57756]_ ,
    \new_[57757]_ , \new_[57758]_ , \new_[57761]_ , \new_[57764]_ ,
    \new_[57765]_ , \new_[57768]_ , \new_[57771]_ , \new_[57772]_ ,
    \new_[57773]_ , \new_[57776]_ , \new_[57779]_ , \new_[57780]_ ,
    \new_[57783]_ , \new_[57786]_ , \new_[57787]_ , \new_[57788]_ ,
    \new_[57791]_ , \new_[57794]_ , \new_[57795]_ , \new_[57798]_ ,
    \new_[57801]_ , \new_[57802]_ , \new_[57803]_ , \new_[57806]_ ,
    \new_[57809]_ , \new_[57810]_ , \new_[57813]_ , \new_[57816]_ ,
    \new_[57817]_ , \new_[57818]_ , \new_[57821]_ , \new_[57824]_ ,
    \new_[57825]_ , \new_[57828]_ , \new_[57831]_ , \new_[57832]_ ,
    \new_[57833]_ , \new_[57836]_ , \new_[57839]_ , \new_[57840]_ ,
    \new_[57843]_ , \new_[57846]_ , \new_[57847]_ , \new_[57848]_ ,
    \new_[57851]_ , \new_[57854]_ , \new_[57855]_ , \new_[57858]_ ,
    \new_[57861]_ , \new_[57862]_ , \new_[57863]_ , \new_[57866]_ ,
    \new_[57869]_ , \new_[57870]_ , \new_[57873]_ , \new_[57876]_ ,
    \new_[57877]_ , \new_[57878]_ , \new_[57881]_ , \new_[57884]_ ,
    \new_[57885]_ , \new_[57888]_ , \new_[57891]_ , \new_[57892]_ ,
    \new_[57893]_ , \new_[57896]_ , \new_[57899]_ , \new_[57900]_ ,
    \new_[57903]_ , \new_[57906]_ , \new_[57907]_ , \new_[57908]_ ,
    \new_[57911]_ , \new_[57914]_ , \new_[57915]_ , \new_[57918]_ ,
    \new_[57921]_ , \new_[57922]_ , \new_[57923]_ , \new_[57926]_ ,
    \new_[57929]_ , \new_[57930]_ , \new_[57933]_ , \new_[57936]_ ,
    \new_[57937]_ , \new_[57938]_ , \new_[57941]_ , \new_[57944]_ ,
    \new_[57945]_ , \new_[57948]_ , \new_[57951]_ , \new_[57952]_ ,
    \new_[57953]_ , \new_[57956]_ , \new_[57959]_ , \new_[57960]_ ,
    \new_[57963]_ , \new_[57966]_ , \new_[57967]_ , \new_[57968]_ ,
    \new_[57971]_ , \new_[57974]_ , \new_[57975]_ , \new_[57978]_ ,
    \new_[57981]_ , \new_[57982]_ , \new_[57983]_ , \new_[57986]_ ,
    \new_[57989]_ , \new_[57990]_ , \new_[57993]_ , \new_[57996]_ ,
    \new_[57997]_ , \new_[57998]_ , \new_[58001]_ , \new_[58004]_ ,
    \new_[58005]_ , \new_[58008]_ , \new_[58011]_ , \new_[58012]_ ,
    \new_[58013]_ , \new_[58016]_ , \new_[58019]_ , \new_[58020]_ ,
    \new_[58023]_ , \new_[58026]_ , \new_[58027]_ , \new_[58028]_ ,
    \new_[58031]_ , \new_[58034]_ , \new_[58035]_ , \new_[58038]_ ,
    \new_[58041]_ , \new_[58042]_ , \new_[58043]_ , \new_[58046]_ ,
    \new_[58049]_ , \new_[58050]_ , \new_[58053]_ , \new_[58056]_ ,
    \new_[58057]_ , \new_[58058]_ , \new_[58061]_ , \new_[58064]_ ,
    \new_[58065]_ , \new_[58068]_ , \new_[58071]_ , \new_[58072]_ ,
    \new_[58073]_ , \new_[58076]_ , \new_[58079]_ , \new_[58080]_ ,
    \new_[58083]_ , \new_[58086]_ , \new_[58087]_ , \new_[58088]_ ,
    \new_[58091]_ , \new_[58094]_ , \new_[58095]_ , \new_[58098]_ ,
    \new_[58101]_ , \new_[58102]_ , \new_[58103]_ , \new_[58106]_ ,
    \new_[58109]_ , \new_[58110]_ , \new_[58113]_ , \new_[58116]_ ,
    \new_[58117]_ , \new_[58118]_ , \new_[58121]_ , \new_[58124]_ ,
    \new_[58125]_ , \new_[58128]_ , \new_[58131]_ , \new_[58132]_ ,
    \new_[58133]_ , \new_[58136]_ , \new_[58139]_ , \new_[58140]_ ,
    \new_[58143]_ , \new_[58146]_ , \new_[58147]_ , \new_[58148]_ ,
    \new_[58151]_ , \new_[58154]_ , \new_[58155]_ , \new_[58158]_ ,
    \new_[58161]_ , \new_[58162]_ , \new_[58163]_ , \new_[58166]_ ,
    \new_[58169]_ , \new_[58170]_ , \new_[58173]_ , \new_[58176]_ ,
    \new_[58177]_ , \new_[58178]_ , \new_[58181]_ , \new_[58184]_ ,
    \new_[58185]_ , \new_[58188]_ , \new_[58191]_ , \new_[58192]_ ,
    \new_[58193]_ , \new_[58196]_ , \new_[58199]_ , \new_[58200]_ ,
    \new_[58203]_ , \new_[58206]_ , \new_[58207]_ , \new_[58208]_ ,
    \new_[58211]_ , \new_[58214]_ , \new_[58215]_ , \new_[58218]_ ,
    \new_[58221]_ , \new_[58222]_ , \new_[58223]_ , \new_[58226]_ ,
    \new_[58229]_ , \new_[58230]_ , \new_[58233]_ , \new_[58236]_ ,
    \new_[58237]_ , \new_[58238]_ , \new_[58241]_ , \new_[58244]_ ,
    \new_[58245]_ , \new_[58248]_ , \new_[58251]_ , \new_[58252]_ ,
    \new_[58253]_ , \new_[58256]_ , \new_[58259]_ , \new_[58260]_ ,
    \new_[58263]_ , \new_[58266]_ , \new_[58267]_ , \new_[58268]_ ,
    \new_[58271]_ , \new_[58274]_ , \new_[58275]_ , \new_[58278]_ ,
    \new_[58281]_ , \new_[58282]_ , \new_[58283]_ , \new_[58286]_ ,
    \new_[58289]_ , \new_[58290]_ , \new_[58293]_ , \new_[58296]_ ,
    \new_[58297]_ , \new_[58298]_ , \new_[58301]_ , \new_[58304]_ ,
    \new_[58305]_ , \new_[58308]_ , \new_[58311]_ , \new_[58312]_ ,
    \new_[58313]_ , \new_[58316]_ , \new_[58319]_ , \new_[58320]_ ,
    \new_[58323]_ , \new_[58326]_ , \new_[58327]_ , \new_[58328]_ ,
    \new_[58331]_ , \new_[58334]_ , \new_[58335]_ , \new_[58338]_ ,
    \new_[58341]_ , \new_[58342]_ , \new_[58343]_ , \new_[58346]_ ,
    \new_[58349]_ , \new_[58350]_ , \new_[58353]_ , \new_[58356]_ ,
    \new_[58357]_ , \new_[58358]_ , \new_[58361]_ , \new_[58364]_ ,
    \new_[58365]_ , \new_[58368]_ , \new_[58371]_ , \new_[58372]_ ,
    \new_[58373]_ , \new_[58376]_ , \new_[58379]_ , \new_[58380]_ ,
    \new_[58383]_ , \new_[58386]_ , \new_[58387]_ , \new_[58388]_ ,
    \new_[58391]_ , \new_[58394]_ , \new_[58395]_ , \new_[58398]_ ,
    \new_[58401]_ , \new_[58402]_ , \new_[58403]_ , \new_[58406]_ ,
    \new_[58409]_ , \new_[58410]_ , \new_[58413]_ , \new_[58416]_ ,
    \new_[58417]_ , \new_[58418]_ , \new_[58421]_ , \new_[58424]_ ,
    \new_[58425]_ , \new_[58428]_ , \new_[58431]_ , \new_[58432]_ ,
    \new_[58433]_ , \new_[58436]_ , \new_[58439]_ , \new_[58440]_ ,
    \new_[58443]_ , \new_[58446]_ , \new_[58447]_ , \new_[58448]_ ,
    \new_[58451]_ , \new_[58454]_ , \new_[58455]_ , \new_[58458]_ ,
    \new_[58461]_ , \new_[58462]_ , \new_[58463]_ , \new_[58466]_ ,
    \new_[58469]_ , \new_[58470]_ , \new_[58473]_ , \new_[58476]_ ,
    \new_[58477]_ , \new_[58478]_ , \new_[58481]_ , \new_[58484]_ ,
    \new_[58485]_ , \new_[58488]_ , \new_[58491]_ , \new_[58492]_ ,
    \new_[58493]_ , \new_[58496]_ , \new_[58499]_ , \new_[58500]_ ,
    \new_[58503]_ , \new_[58506]_ , \new_[58507]_ , \new_[58508]_ ,
    \new_[58511]_ , \new_[58514]_ , \new_[58515]_ , \new_[58518]_ ,
    \new_[58521]_ , \new_[58522]_ , \new_[58523]_ , \new_[58526]_ ,
    \new_[58529]_ , \new_[58530]_ , \new_[58533]_ , \new_[58536]_ ,
    \new_[58537]_ , \new_[58538]_ , \new_[58541]_ , \new_[58544]_ ,
    \new_[58545]_ , \new_[58548]_ , \new_[58551]_ , \new_[58552]_ ,
    \new_[58553]_ , \new_[58556]_ , \new_[58559]_ , \new_[58560]_ ,
    \new_[58563]_ , \new_[58566]_ , \new_[58567]_ , \new_[58568]_ ,
    \new_[58571]_ , \new_[58574]_ , \new_[58575]_ , \new_[58578]_ ,
    \new_[58581]_ , \new_[58582]_ , \new_[58583]_ , \new_[58586]_ ,
    \new_[58589]_ , \new_[58590]_ , \new_[58593]_ , \new_[58596]_ ,
    \new_[58597]_ , \new_[58598]_ , \new_[58601]_ , \new_[58604]_ ,
    \new_[58605]_ , \new_[58608]_ , \new_[58611]_ , \new_[58612]_ ,
    \new_[58613]_ , \new_[58616]_ , \new_[58619]_ , \new_[58620]_ ,
    \new_[58623]_ , \new_[58626]_ , \new_[58627]_ , \new_[58628]_ ,
    \new_[58631]_ , \new_[58634]_ , \new_[58635]_ , \new_[58638]_ ,
    \new_[58641]_ , \new_[58642]_ , \new_[58643]_ , \new_[58646]_ ,
    \new_[58649]_ , \new_[58650]_ , \new_[58653]_ , \new_[58656]_ ,
    \new_[58657]_ , \new_[58658]_ , \new_[58661]_ , \new_[58664]_ ,
    \new_[58665]_ , \new_[58668]_ , \new_[58671]_ , \new_[58672]_ ,
    \new_[58673]_ , \new_[58676]_ , \new_[58679]_ , \new_[58680]_ ,
    \new_[58683]_ , \new_[58686]_ , \new_[58687]_ , \new_[58688]_ ,
    \new_[58691]_ , \new_[58694]_ , \new_[58695]_ , \new_[58698]_ ,
    \new_[58701]_ , \new_[58702]_ , \new_[58703]_ , \new_[58706]_ ,
    \new_[58709]_ , \new_[58710]_ , \new_[58713]_ , \new_[58716]_ ,
    \new_[58717]_ , \new_[58718]_ , \new_[58721]_ , \new_[58724]_ ,
    \new_[58725]_ , \new_[58728]_ , \new_[58731]_ , \new_[58732]_ ,
    \new_[58733]_ , \new_[58736]_ , \new_[58739]_ , \new_[58740]_ ,
    \new_[58743]_ , \new_[58746]_ , \new_[58747]_ , \new_[58748]_ ,
    \new_[58751]_ , \new_[58754]_ , \new_[58755]_ , \new_[58758]_ ,
    \new_[58761]_ , \new_[58762]_ , \new_[58763]_ , \new_[58766]_ ,
    \new_[58769]_ , \new_[58770]_ , \new_[58773]_ , \new_[58776]_ ,
    \new_[58777]_ , \new_[58778]_ , \new_[58781]_ , \new_[58784]_ ,
    \new_[58785]_ , \new_[58788]_ , \new_[58791]_ , \new_[58792]_ ,
    \new_[58793]_ , \new_[58796]_ , \new_[58799]_ , \new_[58800]_ ,
    \new_[58803]_ , \new_[58806]_ , \new_[58807]_ , \new_[58808]_ ,
    \new_[58811]_ , \new_[58814]_ , \new_[58815]_ , \new_[58818]_ ,
    \new_[58821]_ , \new_[58822]_ , \new_[58823]_ , \new_[58826]_ ,
    \new_[58829]_ , \new_[58830]_ , \new_[58833]_ , \new_[58836]_ ,
    \new_[58837]_ , \new_[58838]_ , \new_[58841]_ , \new_[58844]_ ,
    \new_[58845]_ , \new_[58848]_ , \new_[58851]_ , \new_[58852]_ ,
    \new_[58853]_ , \new_[58856]_ , \new_[58859]_ , \new_[58860]_ ,
    \new_[58863]_ , \new_[58866]_ , \new_[58867]_ , \new_[58868]_ ,
    \new_[58871]_ , \new_[58874]_ , \new_[58875]_ , \new_[58878]_ ,
    \new_[58881]_ , \new_[58882]_ , \new_[58883]_ , \new_[58886]_ ,
    \new_[58889]_ , \new_[58890]_ , \new_[58893]_ , \new_[58896]_ ,
    \new_[58897]_ , \new_[58898]_ , \new_[58901]_ , \new_[58904]_ ,
    \new_[58905]_ , \new_[58908]_ , \new_[58911]_ , \new_[58912]_ ,
    \new_[58913]_ , \new_[58916]_ , \new_[58919]_ , \new_[58920]_ ,
    \new_[58923]_ , \new_[58926]_ , \new_[58927]_ , \new_[58928]_ ,
    \new_[58931]_ , \new_[58934]_ , \new_[58935]_ , \new_[58938]_ ,
    \new_[58941]_ , \new_[58942]_ , \new_[58943]_ , \new_[58946]_ ,
    \new_[58949]_ , \new_[58950]_ , \new_[58953]_ , \new_[58956]_ ,
    \new_[58957]_ , \new_[58958]_ , \new_[58961]_ , \new_[58964]_ ,
    \new_[58965]_ , \new_[58968]_ , \new_[58971]_ , \new_[58972]_ ,
    \new_[58973]_ , \new_[58976]_ , \new_[58979]_ , \new_[58980]_ ,
    \new_[58983]_ , \new_[58986]_ , \new_[58987]_ , \new_[58988]_ ,
    \new_[58991]_ , \new_[58994]_ , \new_[58995]_ , \new_[58998]_ ,
    \new_[59001]_ , \new_[59002]_ , \new_[59003]_ , \new_[59006]_ ,
    \new_[59009]_ , \new_[59010]_ , \new_[59013]_ , \new_[59016]_ ,
    \new_[59017]_ , \new_[59018]_ , \new_[59021]_ , \new_[59024]_ ,
    \new_[59025]_ , \new_[59028]_ , \new_[59031]_ , \new_[59032]_ ,
    \new_[59033]_ , \new_[59036]_ , \new_[59039]_ , \new_[59040]_ ,
    \new_[59043]_ , \new_[59046]_ , \new_[59047]_ , \new_[59048]_ ,
    \new_[59051]_ , \new_[59054]_ , \new_[59055]_ , \new_[59058]_ ,
    \new_[59061]_ , \new_[59062]_ , \new_[59063]_ , \new_[59066]_ ,
    \new_[59069]_ , \new_[59070]_ , \new_[59073]_ , \new_[59076]_ ,
    \new_[59077]_ , \new_[59078]_ , \new_[59081]_ , \new_[59084]_ ,
    \new_[59085]_ , \new_[59088]_ , \new_[59091]_ , \new_[59092]_ ,
    \new_[59093]_ , \new_[59096]_ , \new_[59099]_ , \new_[59100]_ ,
    \new_[59103]_ , \new_[59106]_ , \new_[59107]_ , \new_[59108]_ ,
    \new_[59111]_ , \new_[59114]_ , \new_[59115]_ , \new_[59118]_ ,
    \new_[59121]_ , \new_[59122]_ , \new_[59123]_ , \new_[59126]_ ,
    \new_[59129]_ , \new_[59130]_ , \new_[59133]_ , \new_[59136]_ ,
    \new_[59137]_ , \new_[59138]_ , \new_[59141]_ , \new_[59144]_ ,
    \new_[59145]_ , \new_[59148]_ , \new_[59151]_ , \new_[59152]_ ,
    \new_[59153]_ , \new_[59156]_ , \new_[59159]_ , \new_[59160]_ ,
    \new_[59163]_ , \new_[59166]_ , \new_[59167]_ , \new_[59168]_ ,
    \new_[59171]_ , \new_[59174]_ , \new_[59175]_ , \new_[59178]_ ,
    \new_[59181]_ , \new_[59182]_ , \new_[59183]_ , \new_[59186]_ ,
    \new_[59189]_ , \new_[59190]_ , \new_[59193]_ , \new_[59196]_ ,
    \new_[59197]_ , \new_[59198]_ , \new_[59201]_ , \new_[59204]_ ,
    \new_[59205]_ , \new_[59208]_ , \new_[59211]_ , \new_[59212]_ ,
    \new_[59213]_ , \new_[59216]_ , \new_[59219]_ , \new_[59220]_ ,
    \new_[59223]_ , \new_[59226]_ , \new_[59227]_ , \new_[59228]_ ,
    \new_[59231]_ , \new_[59234]_ , \new_[59235]_ , \new_[59238]_ ,
    \new_[59241]_ , \new_[59242]_ , \new_[59243]_ , \new_[59246]_ ,
    \new_[59249]_ , \new_[59250]_ , \new_[59253]_ , \new_[59256]_ ,
    \new_[59257]_ , \new_[59258]_ , \new_[59261]_ , \new_[59264]_ ,
    \new_[59265]_ , \new_[59268]_ , \new_[59271]_ , \new_[59272]_ ,
    \new_[59273]_ , \new_[59276]_ , \new_[59279]_ , \new_[59280]_ ,
    \new_[59283]_ , \new_[59286]_ , \new_[59287]_ , \new_[59288]_ ,
    \new_[59291]_ , \new_[59294]_ , \new_[59295]_ , \new_[59298]_ ,
    \new_[59301]_ , \new_[59302]_ , \new_[59303]_ , \new_[59306]_ ,
    \new_[59309]_ , \new_[59310]_ , \new_[59313]_ , \new_[59316]_ ,
    \new_[59317]_ , \new_[59318]_ , \new_[59321]_ , \new_[59324]_ ,
    \new_[59325]_ , \new_[59328]_ , \new_[59331]_ , \new_[59332]_ ,
    \new_[59333]_ , \new_[59336]_ , \new_[59339]_ , \new_[59340]_ ,
    \new_[59343]_ , \new_[59346]_ , \new_[59347]_ , \new_[59348]_ ,
    \new_[59351]_ , \new_[59354]_ , \new_[59355]_ , \new_[59358]_ ,
    \new_[59361]_ , \new_[59362]_ , \new_[59363]_ , \new_[59366]_ ,
    \new_[59369]_ , \new_[59370]_ , \new_[59373]_ , \new_[59376]_ ,
    \new_[59377]_ , \new_[59378]_ , \new_[59381]_ , \new_[59384]_ ,
    \new_[59385]_ , \new_[59388]_ , \new_[59391]_ , \new_[59392]_ ,
    \new_[59393]_ , \new_[59396]_ , \new_[59399]_ , \new_[59400]_ ,
    \new_[59403]_ , \new_[59406]_ , \new_[59407]_ , \new_[59408]_ ,
    \new_[59411]_ , \new_[59414]_ , \new_[59415]_ , \new_[59418]_ ,
    \new_[59421]_ , \new_[59422]_ , \new_[59423]_ , \new_[59426]_ ,
    \new_[59429]_ , \new_[59430]_ , \new_[59433]_ , \new_[59436]_ ,
    \new_[59437]_ , \new_[59438]_ , \new_[59441]_ , \new_[59444]_ ,
    \new_[59445]_ , \new_[59448]_ , \new_[59451]_ , \new_[59452]_ ,
    \new_[59453]_ , \new_[59456]_ , \new_[59459]_ , \new_[59460]_ ,
    \new_[59463]_ , \new_[59466]_ , \new_[59467]_ , \new_[59468]_ ,
    \new_[59471]_ , \new_[59474]_ , \new_[59475]_ , \new_[59478]_ ,
    \new_[59481]_ , \new_[59482]_ , \new_[59483]_ , \new_[59486]_ ,
    \new_[59489]_ , \new_[59490]_ , \new_[59493]_ , \new_[59496]_ ,
    \new_[59497]_ , \new_[59498]_ , \new_[59501]_ , \new_[59504]_ ,
    \new_[59505]_ , \new_[59508]_ , \new_[59511]_ , \new_[59512]_ ,
    \new_[59513]_ , \new_[59516]_ , \new_[59519]_ , \new_[59520]_ ,
    \new_[59523]_ , \new_[59526]_ , \new_[59527]_ , \new_[59528]_ ,
    \new_[59531]_ , \new_[59534]_ , \new_[59535]_ , \new_[59538]_ ,
    \new_[59541]_ , \new_[59542]_ , \new_[59543]_ , \new_[59546]_ ,
    \new_[59549]_ , \new_[59550]_ , \new_[59553]_ , \new_[59556]_ ,
    \new_[59557]_ , \new_[59558]_ , \new_[59561]_ , \new_[59564]_ ,
    \new_[59565]_ , \new_[59568]_ , \new_[59571]_ , \new_[59572]_ ,
    \new_[59573]_ , \new_[59576]_ , \new_[59579]_ , \new_[59580]_ ,
    \new_[59583]_ , \new_[59586]_ , \new_[59587]_ , \new_[59588]_ ,
    \new_[59591]_ , \new_[59594]_ , \new_[59595]_ , \new_[59598]_ ,
    \new_[59601]_ , \new_[59602]_ , \new_[59603]_ , \new_[59606]_ ,
    \new_[59609]_ , \new_[59610]_ , \new_[59613]_ , \new_[59616]_ ,
    \new_[59617]_ , \new_[59618]_ , \new_[59621]_ , \new_[59624]_ ,
    \new_[59625]_ , \new_[59628]_ , \new_[59631]_ , \new_[59632]_ ,
    \new_[59633]_ , \new_[59636]_ , \new_[59639]_ , \new_[59640]_ ,
    \new_[59643]_ , \new_[59646]_ , \new_[59647]_ , \new_[59648]_ ,
    \new_[59651]_ , \new_[59654]_ , \new_[59655]_ , \new_[59658]_ ,
    \new_[59661]_ , \new_[59662]_ , \new_[59663]_ , \new_[59666]_ ,
    \new_[59669]_ , \new_[59670]_ , \new_[59673]_ , \new_[59676]_ ,
    \new_[59677]_ , \new_[59678]_ , \new_[59681]_ , \new_[59684]_ ,
    \new_[59685]_ , \new_[59688]_ , \new_[59691]_ , \new_[59692]_ ,
    \new_[59693]_ , \new_[59696]_ , \new_[59699]_ , \new_[59700]_ ,
    \new_[59703]_ , \new_[59706]_ , \new_[59707]_ , \new_[59708]_ ,
    \new_[59711]_ , \new_[59714]_ , \new_[59715]_ , \new_[59718]_ ,
    \new_[59721]_ , \new_[59722]_ , \new_[59723]_ , \new_[59726]_ ,
    \new_[59729]_ , \new_[59730]_ , \new_[59733]_ , \new_[59736]_ ,
    \new_[59737]_ , \new_[59738]_ , \new_[59741]_ , \new_[59744]_ ,
    \new_[59745]_ , \new_[59748]_ , \new_[59751]_ , \new_[59752]_ ,
    \new_[59753]_ , \new_[59756]_ , \new_[59759]_ , \new_[59760]_ ,
    \new_[59763]_ , \new_[59766]_ , \new_[59767]_ , \new_[59768]_ ,
    \new_[59771]_ , \new_[59774]_ , \new_[59775]_ , \new_[59778]_ ,
    \new_[59781]_ , \new_[59782]_ , \new_[59783]_ , \new_[59786]_ ,
    \new_[59789]_ , \new_[59790]_ , \new_[59793]_ , \new_[59796]_ ,
    \new_[59797]_ , \new_[59798]_ , \new_[59801]_ , \new_[59804]_ ,
    \new_[59805]_ , \new_[59808]_ , \new_[59811]_ , \new_[59812]_ ,
    \new_[59813]_ , \new_[59816]_ , \new_[59819]_ , \new_[59820]_ ,
    \new_[59823]_ , \new_[59826]_ , \new_[59827]_ , \new_[59828]_ ,
    \new_[59831]_ , \new_[59834]_ , \new_[59835]_ , \new_[59838]_ ,
    \new_[59841]_ , \new_[59842]_ , \new_[59843]_ , \new_[59846]_ ,
    \new_[59849]_ , \new_[59850]_ , \new_[59853]_ , \new_[59856]_ ,
    \new_[59857]_ , \new_[59858]_ , \new_[59861]_ , \new_[59864]_ ,
    \new_[59865]_ , \new_[59868]_ , \new_[59871]_ , \new_[59872]_ ,
    \new_[59873]_ , \new_[59876]_ , \new_[59879]_ , \new_[59880]_ ,
    \new_[59883]_ , \new_[59886]_ , \new_[59887]_ , \new_[59888]_ ,
    \new_[59891]_ , \new_[59894]_ , \new_[59895]_ , \new_[59898]_ ,
    \new_[59901]_ , \new_[59902]_ , \new_[59903]_ , \new_[59906]_ ,
    \new_[59909]_ , \new_[59910]_ , \new_[59913]_ , \new_[59916]_ ,
    \new_[59917]_ , \new_[59918]_ , \new_[59921]_ , \new_[59924]_ ,
    \new_[59925]_ , \new_[59928]_ , \new_[59931]_ , \new_[59932]_ ,
    \new_[59933]_ , \new_[59936]_ , \new_[59939]_ , \new_[59940]_ ,
    \new_[59943]_ , \new_[59946]_ , \new_[59947]_ , \new_[59948]_ ,
    \new_[59951]_ , \new_[59954]_ , \new_[59955]_ , \new_[59958]_ ,
    \new_[59961]_ , \new_[59962]_ , \new_[59963]_ , \new_[59966]_ ,
    \new_[59969]_ , \new_[59970]_ , \new_[59973]_ , \new_[59976]_ ,
    \new_[59977]_ , \new_[59978]_ , \new_[59981]_ , \new_[59984]_ ,
    \new_[59985]_ , \new_[59988]_ , \new_[59991]_ , \new_[59992]_ ,
    \new_[59993]_ , \new_[59996]_ , \new_[59999]_ , \new_[60000]_ ,
    \new_[60003]_ , \new_[60006]_ , \new_[60007]_ , \new_[60008]_ ,
    \new_[60011]_ , \new_[60014]_ , \new_[60015]_ , \new_[60018]_ ,
    \new_[60021]_ , \new_[60022]_ , \new_[60023]_ , \new_[60026]_ ,
    \new_[60029]_ , \new_[60030]_ , \new_[60033]_ , \new_[60036]_ ,
    \new_[60037]_ , \new_[60038]_ , \new_[60041]_ , \new_[60044]_ ,
    \new_[60045]_ , \new_[60048]_ , \new_[60051]_ , \new_[60052]_ ,
    \new_[60053]_ , \new_[60056]_ , \new_[60059]_ , \new_[60060]_ ,
    \new_[60063]_ , \new_[60066]_ , \new_[60067]_ , \new_[60068]_ ,
    \new_[60071]_ , \new_[60074]_ , \new_[60075]_ , \new_[60078]_ ,
    \new_[60081]_ , \new_[60082]_ , \new_[60083]_ , \new_[60086]_ ,
    \new_[60089]_ , \new_[60090]_ , \new_[60093]_ , \new_[60096]_ ,
    \new_[60097]_ , \new_[60098]_ , \new_[60101]_ , \new_[60104]_ ,
    \new_[60105]_ , \new_[60108]_ , \new_[60111]_ , \new_[60112]_ ,
    \new_[60113]_ , \new_[60116]_ , \new_[60119]_ , \new_[60120]_ ,
    \new_[60123]_ , \new_[60126]_ , \new_[60127]_ , \new_[60128]_ ,
    \new_[60131]_ , \new_[60134]_ , \new_[60135]_ , \new_[60138]_ ,
    \new_[60141]_ , \new_[60142]_ , \new_[60143]_ , \new_[60146]_ ,
    \new_[60149]_ , \new_[60150]_ , \new_[60153]_ , \new_[60156]_ ,
    \new_[60157]_ , \new_[60158]_ , \new_[60161]_ , \new_[60164]_ ,
    \new_[60165]_ , \new_[60168]_ , \new_[60171]_ , \new_[60172]_ ,
    \new_[60173]_ , \new_[60176]_ , \new_[60179]_ , \new_[60180]_ ,
    \new_[60183]_ , \new_[60186]_ , \new_[60187]_ , \new_[60188]_ ,
    \new_[60191]_ , \new_[60194]_ , \new_[60195]_ , \new_[60198]_ ,
    \new_[60201]_ , \new_[60202]_ , \new_[60203]_ , \new_[60206]_ ,
    \new_[60209]_ , \new_[60210]_ , \new_[60213]_ , \new_[60216]_ ,
    \new_[60217]_ , \new_[60218]_ , \new_[60221]_ , \new_[60224]_ ,
    \new_[60225]_ , \new_[60228]_ , \new_[60231]_ , \new_[60232]_ ,
    \new_[60233]_ , \new_[60236]_ , \new_[60239]_ , \new_[60240]_ ,
    \new_[60243]_ , \new_[60246]_ , \new_[60247]_ , \new_[60248]_ ,
    \new_[60251]_ , \new_[60254]_ , \new_[60255]_ , \new_[60258]_ ,
    \new_[60261]_ , \new_[60262]_ , \new_[60263]_ , \new_[60266]_ ,
    \new_[60269]_ , \new_[60270]_ , \new_[60273]_ , \new_[60276]_ ,
    \new_[60277]_ , \new_[60278]_ , \new_[60281]_ , \new_[60284]_ ,
    \new_[60285]_ , \new_[60288]_ , \new_[60291]_ , \new_[60292]_ ,
    \new_[60293]_ , \new_[60296]_ , \new_[60299]_ , \new_[60300]_ ,
    \new_[60303]_ , \new_[60306]_ , \new_[60307]_ , \new_[60308]_ ,
    \new_[60311]_ , \new_[60314]_ , \new_[60315]_ , \new_[60318]_ ,
    \new_[60321]_ , \new_[60322]_ , \new_[60323]_ , \new_[60326]_ ,
    \new_[60329]_ , \new_[60330]_ , \new_[60333]_ , \new_[60336]_ ,
    \new_[60337]_ , \new_[60338]_ , \new_[60341]_ , \new_[60344]_ ,
    \new_[60345]_ , \new_[60348]_ , \new_[60351]_ , \new_[60352]_ ,
    \new_[60353]_ , \new_[60356]_ , \new_[60359]_ , \new_[60360]_ ,
    \new_[60363]_ , \new_[60366]_ , \new_[60367]_ , \new_[60368]_ ,
    \new_[60371]_ , \new_[60374]_ , \new_[60375]_ , \new_[60378]_ ,
    \new_[60381]_ , \new_[60382]_ , \new_[60383]_ , \new_[60386]_ ,
    \new_[60389]_ , \new_[60390]_ , \new_[60393]_ , \new_[60396]_ ,
    \new_[60397]_ , \new_[60398]_ , \new_[60401]_ , \new_[60404]_ ,
    \new_[60405]_ , \new_[60408]_ , \new_[60411]_ , \new_[60412]_ ,
    \new_[60413]_ , \new_[60416]_ , \new_[60419]_ , \new_[60420]_ ,
    \new_[60423]_ , \new_[60426]_ , \new_[60427]_ , \new_[60428]_ ,
    \new_[60431]_ , \new_[60434]_ , \new_[60435]_ , \new_[60438]_ ,
    \new_[60441]_ , \new_[60442]_ , \new_[60443]_ , \new_[60446]_ ,
    \new_[60449]_ , \new_[60450]_ , \new_[60453]_ , \new_[60456]_ ,
    \new_[60457]_ , \new_[60458]_ , \new_[60461]_ , \new_[60464]_ ,
    \new_[60465]_ , \new_[60468]_ , \new_[60471]_ , \new_[60472]_ ,
    \new_[60473]_ , \new_[60476]_ , \new_[60479]_ , \new_[60480]_ ,
    \new_[60483]_ , \new_[60486]_ , \new_[60487]_ , \new_[60488]_ ,
    \new_[60491]_ , \new_[60494]_ , \new_[60495]_ , \new_[60498]_ ,
    \new_[60501]_ , \new_[60502]_ , \new_[60503]_ , \new_[60506]_ ,
    \new_[60509]_ , \new_[60510]_ , \new_[60513]_ , \new_[60516]_ ,
    \new_[60517]_ , \new_[60518]_ , \new_[60521]_ , \new_[60524]_ ,
    \new_[60525]_ , \new_[60528]_ , \new_[60531]_ , \new_[60532]_ ,
    \new_[60533]_ , \new_[60536]_ , \new_[60539]_ , \new_[60540]_ ,
    \new_[60543]_ , \new_[60546]_ , \new_[60547]_ , \new_[60548]_ ,
    \new_[60551]_ , \new_[60554]_ , \new_[60555]_ , \new_[60558]_ ,
    \new_[60561]_ , \new_[60562]_ , \new_[60563]_ , \new_[60566]_ ,
    \new_[60569]_ , \new_[60570]_ , \new_[60573]_ , \new_[60576]_ ,
    \new_[60577]_ , \new_[60578]_ , \new_[60581]_ , \new_[60584]_ ,
    \new_[60585]_ , \new_[60588]_ , \new_[60591]_ , \new_[60592]_ ,
    \new_[60593]_ , \new_[60596]_ , \new_[60599]_ , \new_[60600]_ ,
    \new_[60603]_ , \new_[60606]_ , \new_[60607]_ , \new_[60608]_ ,
    \new_[60611]_ , \new_[60614]_ , \new_[60615]_ , \new_[60618]_ ,
    \new_[60621]_ , \new_[60622]_ , \new_[60623]_ , \new_[60626]_ ,
    \new_[60629]_ , \new_[60630]_ , \new_[60633]_ , \new_[60636]_ ,
    \new_[60637]_ , \new_[60638]_ , \new_[60641]_ , \new_[60644]_ ,
    \new_[60645]_ , \new_[60648]_ , \new_[60651]_ , \new_[60652]_ ,
    \new_[60653]_ , \new_[60656]_ , \new_[60659]_ , \new_[60660]_ ,
    \new_[60663]_ , \new_[60666]_ , \new_[60667]_ , \new_[60668]_ ,
    \new_[60671]_ , \new_[60674]_ , \new_[60675]_ , \new_[60678]_ ,
    \new_[60681]_ , \new_[60682]_ , \new_[60683]_ , \new_[60686]_ ,
    \new_[60689]_ , \new_[60690]_ , \new_[60693]_ , \new_[60696]_ ,
    \new_[60697]_ , \new_[60698]_ , \new_[60701]_ , \new_[60704]_ ,
    \new_[60705]_ , \new_[60708]_ , \new_[60711]_ , \new_[60712]_ ,
    \new_[60713]_ , \new_[60716]_ , \new_[60719]_ , \new_[60720]_ ,
    \new_[60723]_ , \new_[60726]_ , \new_[60727]_ , \new_[60728]_ ,
    \new_[60731]_ , \new_[60734]_ , \new_[60735]_ , \new_[60738]_ ,
    \new_[60741]_ , \new_[60742]_ , \new_[60743]_ , \new_[60746]_ ,
    \new_[60749]_ , \new_[60750]_ , \new_[60753]_ , \new_[60756]_ ,
    \new_[60757]_ , \new_[60758]_ , \new_[60761]_ , \new_[60764]_ ,
    \new_[60765]_ , \new_[60768]_ , \new_[60771]_ , \new_[60772]_ ,
    \new_[60773]_ , \new_[60776]_ , \new_[60779]_ , \new_[60780]_ ,
    \new_[60783]_ , \new_[60786]_ , \new_[60787]_ , \new_[60788]_ ,
    \new_[60791]_ , \new_[60794]_ , \new_[60795]_ , \new_[60798]_ ,
    \new_[60801]_ , \new_[60802]_ , \new_[60803]_ , \new_[60806]_ ,
    \new_[60809]_ , \new_[60810]_ , \new_[60813]_ , \new_[60816]_ ,
    \new_[60817]_ , \new_[60818]_ , \new_[60821]_ , \new_[60824]_ ,
    \new_[60825]_ , \new_[60828]_ , \new_[60831]_ , \new_[60832]_ ,
    \new_[60833]_ , \new_[60836]_ , \new_[60839]_ , \new_[60840]_ ,
    \new_[60843]_ , \new_[60846]_ , \new_[60847]_ , \new_[60848]_ ,
    \new_[60851]_ , \new_[60854]_ , \new_[60855]_ , \new_[60858]_ ,
    \new_[60861]_ , \new_[60862]_ , \new_[60863]_ , \new_[60866]_ ,
    \new_[60869]_ , \new_[60870]_ , \new_[60873]_ , \new_[60876]_ ,
    \new_[60877]_ , \new_[60878]_ , \new_[60881]_ , \new_[60884]_ ,
    \new_[60885]_ , \new_[60888]_ , \new_[60891]_ , \new_[60892]_ ,
    \new_[60893]_ , \new_[60896]_ , \new_[60899]_ , \new_[60900]_ ,
    \new_[60903]_ , \new_[60906]_ , \new_[60907]_ , \new_[60908]_ ,
    \new_[60911]_ , \new_[60914]_ , \new_[60915]_ , \new_[60918]_ ,
    \new_[60921]_ , \new_[60922]_ , \new_[60923]_ , \new_[60926]_ ,
    \new_[60929]_ , \new_[60930]_ , \new_[60933]_ , \new_[60936]_ ,
    \new_[60937]_ , \new_[60938]_ , \new_[60941]_ , \new_[60944]_ ,
    \new_[60945]_ , \new_[60948]_ , \new_[60951]_ , \new_[60952]_ ,
    \new_[60953]_ , \new_[60956]_ , \new_[60959]_ , \new_[60960]_ ,
    \new_[60963]_ , \new_[60966]_ , \new_[60967]_ , \new_[60968]_ ,
    \new_[60971]_ , \new_[60974]_ , \new_[60975]_ , \new_[60978]_ ,
    \new_[60981]_ , \new_[60982]_ , \new_[60983]_ , \new_[60986]_ ,
    \new_[60989]_ , \new_[60990]_ , \new_[60993]_ , \new_[60996]_ ,
    \new_[60997]_ , \new_[60998]_ , \new_[61001]_ , \new_[61004]_ ,
    \new_[61005]_ , \new_[61008]_ , \new_[61011]_ , \new_[61012]_ ,
    \new_[61013]_ , \new_[61016]_ , \new_[61019]_ , \new_[61020]_ ,
    \new_[61023]_ , \new_[61026]_ , \new_[61027]_ , \new_[61028]_ ,
    \new_[61031]_ , \new_[61034]_ , \new_[61035]_ , \new_[61038]_ ,
    \new_[61041]_ , \new_[61042]_ , \new_[61043]_ , \new_[61046]_ ,
    \new_[61049]_ , \new_[61050]_ , \new_[61053]_ , \new_[61056]_ ,
    \new_[61057]_ , \new_[61058]_ , \new_[61061]_ , \new_[61064]_ ,
    \new_[61065]_ , \new_[61068]_ , \new_[61071]_ , \new_[61072]_ ,
    \new_[61073]_ , \new_[61076]_ , \new_[61079]_ , \new_[61080]_ ,
    \new_[61083]_ , \new_[61086]_ , \new_[61087]_ , \new_[61088]_ ,
    \new_[61091]_ , \new_[61094]_ , \new_[61095]_ , \new_[61098]_ ,
    \new_[61101]_ , \new_[61102]_ , \new_[61103]_ , \new_[61106]_ ,
    \new_[61109]_ , \new_[61110]_ , \new_[61113]_ , \new_[61116]_ ,
    \new_[61117]_ , \new_[61118]_ , \new_[61121]_ , \new_[61124]_ ,
    \new_[61125]_ , \new_[61128]_ , \new_[61131]_ , \new_[61132]_ ,
    \new_[61133]_ , \new_[61136]_ , \new_[61139]_ , \new_[61140]_ ,
    \new_[61143]_ , \new_[61146]_ , \new_[61147]_ , \new_[61148]_ ,
    \new_[61151]_ , \new_[61154]_ , \new_[61155]_ , \new_[61158]_ ,
    \new_[61161]_ , \new_[61162]_ , \new_[61163]_ , \new_[61166]_ ,
    \new_[61169]_ , \new_[61170]_ , \new_[61173]_ , \new_[61176]_ ,
    \new_[61177]_ , \new_[61178]_ , \new_[61181]_ , \new_[61184]_ ,
    \new_[61185]_ , \new_[61188]_ , \new_[61191]_ , \new_[61192]_ ,
    \new_[61193]_ , \new_[61196]_ , \new_[61199]_ , \new_[61200]_ ,
    \new_[61203]_ , \new_[61206]_ , \new_[61207]_ , \new_[61208]_ ,
    \new_[61211]_ , \new_[61214]_ , \new_[61215]_ , \new_[61218]_ ,
    \new_[61221]_ , \new_[61222]_ , \new_[61223]_ , \new_[61226]_ ,
    \new_[61229]_ , \new_[61230]_ , \new_[61233]_ , \new_[61236]_ ,
    \new_[61237]_ , \new_[61238]_ , \new_[61241]_ , \new_[61244]_ ,
    \new_[61245]_ , \new_[61248]_ , \new_[61251]_ , \new_[61252]_ ,
    \new_[61253]_ , \new_[61256]_ , \new_[61259]_ , \new_[61260]_ ,
    \new_[61263]_ , \new_[61266]_ , \new_[61267]_ , \new_[61268]_ ,
    \new_[61271]_ , \new_[61274]_ , \new_[61275]_ , \new_[61278]_ ,
    \new_[61281]_ , \new_[61282]_ , \new_[61283]_ , \new_[61286]_ ,
    \new_[61289]_ , \new_[61290]_ , \new_[61293]_ , \new_[61296]_ ,
    \new_[61297]_ , \new_[61298]_ , \new_[61301]_ , \new_[61304]_ ,
    \new_[61305]_ , \new_[61308]_ , \new_[61311]_ , \new_[61312]_ ,
    \new_[61313]_ , \new_[61316]_ , \new_[61319]_ , \new_[61320]_ ,
    \new_[61323]_ , \new_[61326]_ , \new_[61327]_ , \new_[61328]_ ,
    \new_[61331]_ , \new_[61334]_ , \new_[61335]_ , \new_[61338]_ ,
    \new_[61341]_ , \new_[61342]_ , \new_[61343]_ , \new_[61346]_ ,
    \new_[61349]_ , \new_[61350]_ , \new_[61353]_ , \new_[61356]_ ,
    \new_[61357]_ , \new_[61358]_ , \new_[61361]_ , \new_[61364]_ ,
    \new_[61365]_ , \new_[61368]_ , \new_[61371]_ , \new_[61372]_ ,
    \new_[61373]_ , \new_[61376]_ , \new_[61379]_ , \new_[61380]_ ,
    \new_[61383]_ , \new_[61386]_ , \new_[61387]_ , \new_[61388]_ ,
    \new_[61391]_ , \new_[61394]_ , \new_[61395]_ , \new_[61398]_ ,
    \new_[61401]_ , \new_[61402]_ , \new_[61403]_ , \new_[61406]_ ,
    \new_[61409]_ , \new_[61410]_ , \new_[61413]_ , \new_[61416]_ ,
    \new_[61417]_ , \new_[61418]_ , \new_[61421]_ , \new_[61424]_ ,
    \new_[61425]_ , \new_[61428]_ , \new_[61431]_ , \new_[61432]_ ,
    \new_[61433]_ , \new_[61436]_ , \new_[61439]_ , \new_[61440]_ ,
    \new_[61443]_ , \new_[61446]_ , \new_[61447]_ , \new_[61448]_ ,
    \new_[61451]_ , \new_[61454]_ , \new_[61455]_ , \new_[61458]_ ,
    \new_[61461]_ , \new_[61462]_ , \new_[61463]_ , \new_[61466]_ ,
    \new_[61469]_ , \new_[61470]_ , \new_[61473]_ , \new_[61476]_ ,
    \new_[61477]_ , \new_[61478]_ , \new_[61481]_ , \new_[61484]_ ,
    \new_[61485]_ , \new_[61488]_ , \new_[61491]_ , \new_[61492]_ ,
    \new_[61493]_ , \new_[61496]_ , \new_[61499]_ , \new_[61500]_ ,
    \new_[61503]_ , \new_[61506]_ , \new_[61507]_ , \new_[61508]_ ,
    \new_[61511]_ , \new_[61514]_ , \new_[61515]_ , \new_[61518]_ ,
    \new_[61521]_ , \new_[61522]_ , \new_[61523]_ , \new_[61526]_ ,
    \new_[61529]_ , \new_[61530]_ , \new_[61533]_ , \new_[61536]_ ,
    \new_[61537]_ , \new_[61538]_ , \new_[61541]_ , \new_[61544]_ ,
    \new_[61545]_ , \new_[61548]_ , \new_[61551]_ , \new_[61552]_ ,
    \new_[61553]_ , \new_[61556]_ , \new_[61559]_ , \new_[61560]_ ,
    \new_[61563]_ , \new_[61566]_ , \new_[61567]_ , \new_[61568]_ ,
    \new_[61571]_ , \new_[61574]_ , \new_[61575]_ , \new_[61578]_ ,
    \new_[61581]_ , \new_[61582]_ , \new_[61583]_ , \new_[61586]_ ,
    \new_[61589]_ , \new_[61590]_ , \new_[61593]_ , \new_[61596]_ ,
    \new_[61597]_ , \new_[61598]_ , \new_[61601]_ , \new_[61604]_ ,
    \new_[61605]_ , \new_[61608]_ , \new_[61611]_ , \new_[61612]_ ,
    \new_[61613]_ , \new_[61616]_ , \new_[61619]_ , \new_[61620]_ ,
    \new_[61623]_ , \new_[61626]_ , \new_[61627]_ , \new_[61628]_ ,
    \new_[61631]_ , \new_[61634]_ , \new_[61635]_ , \new_[61638]_ ,
    \new_[61641]_ , \new_[61642]_ , \new_[61643]_ , \new_[61646]_ ,
    \new_[61649]_ , \new_[61650]_ , \new_[61653]_ , \new_[61656]_ ,
    \new_[61657]_ , \new_[61658]_ , \new_[61661]_ , \new_[61664]_ ,
    \new_[61665]_ , \new_[61668]_ , \new_[61671]_ , \new_[61672]_ ,
    \new_[61673]_ , \new_[61676]_ , \new_[61679]_ , \new_[61680]_ ,
    \new_[61683]_ , \new_[61686]_ , \new_[61687]_ , \new_[61688]_ ,
    \new_[61691]_ , \new_[61694]_ , \new_[61695]_ , \new_[61698]_ ,
    \new_[61701]_ , \new_[61702]_ , \new_[61703]_ , \new_[61706]_ ,
    \new_[61709]_ , \new_[61710]_ , \new_[61713]_ , \new_[61716]_ ,
    \new_[61717]_ , \new_[61718]_ , \new_[61721]_ , \new_[61724]_ ,
    \new_[61725]_ , \new_[61728]_ , \new_[61731]_ , \new_[61732]_ ,
    \new_[61733]_ , \new_[61736]_ , \new_[61739]_ , \new_[61740]_ ,
    \new_[61743]_ , \new_[61746]_ , \new_[61747]_ , \new_[61748]_ ,
    \new_[61751]_ , \new_[61754]_ , \new_[61755]_ , \new_[61758]_ ,
    \new_[61761]_ , \new_[61762]_ , \new_[61763]_ , \new_[61766]_ ,
    \new_[61769]_ , \new_[61770]_ , \new_[61773]_ , \new_[61776]_ ,
    \new_[61777]_ , \new_[61778]_ , \new_[61781]_ , \new_[61784]_ ,
    \new_[61785]_ , \new_[61788]_ , \new_[61791]_ , \new_[61792]_ ,
    \new_[61793]_ , \new_[61796]_ , \new_[61799]_ , \new_[61800]_ ,
    \new_[61803]_ , \new_[61806]_ , \new_[61807]_ , \new_[61808]_ ,
    \new_[61811]_ , \new_[61814]_ , \new_[61815]_ , \new_[61818]_ ,
    \new_[61821]_ , \new_[61822]_ , \new_[61823]_ , \new_[61826]_ ,
    \new_[61829]_ , \new_[61830]_ , \new_[61833]_ , \new_[61836]_ ,
    \new_[61837]_ , \new_[61838]_ , \new_[61841]_ , \new_[61844]_ ,
    \new_[61845]_ , \new_[61848]_ , \new_[61851]_ , \new_[61852]_ ,
    \new_[61853]_ , \new_[61856]_ , \new_[61859]_ , \new_[61860]_ ,
    \new_[61863]_ , \new_[61866]_ , \new_[61867]_ , \new_[61868]_ ,
    \new_[61871]_ , \new_[61874]_ , \new_[61875]_ , \new_[61878]_ ,
    \new_[61881]_ , \new_[61882]_ , \new_[61883]_ , \new_[61886]_ ,
    \new_[61889]_ , \new_[61890]_ , \new_[61893]_ , \new_[61896]_ ,
    \new_[61897]_ , \new_[61898]_ , \new_[61901]_ , \new_[61904]_ ,
    \new_[61905]_ , \new_[61908]_ , \new_[61911]_ , \new_[61912]_ ,
    \new_[61913]_ , \new_[61916]_ , \new_[61919]_ , \new_[61920]_ ,
    \new_[61923]_ , \new_[61926]_ , \new_[61927]_ , \new_[61928]_ ,
    \new_[61931]_ , \new_[61934]_ , \new_[61935]_ , \new_[61938]_ ,
    \new_[61941]_ , \new_[61942]_ , \new_[61943]_ , \new_[61946]_ ,
    \new_[61949]_ , \new_[61950]_ , \new_[61953]_ , \new_[61956]_ ,
    \new_[61957]_ , \new_[61958]_ , \new_[61961]_ , \new_[61964]_ ,
    \new_[61965]_ , \new_[61968]_ , \new_[61971]_ , \new_[61972]_ ,
    \new_[61973]_ , \new_[61976]_ , \new_[61979]_ , \new_[61980]_ ,
    \new_[61983]_ , \new_[61986]_ , \new_[61987]_ , \new_[61988]_ ,
    \new_[61991]_ , \new_[61994]_ , \new_[61995]_ , \new_[61998]_ ,
    \new_[62001]_ , \new_[62002]_ , \new_[62003]_ , \new_[62006]_ ,
    \new_[62009]_ , \new_[62010]_ , \new_[62013]_ , \new_[62016]_ ,
    \new_[62017]_ , \new_[62018]_ , \new_[62021]_ , \new_[62024]_ ,
    \new_[62025]_ , \new_[62028]_ , \new_[62031]_ , \new_[62032]_ ,
    \new_[62033]_ , \new_[62036]_ , \new_[62039]_ , \new_[62040]_ ,
    \new_[62043]_ , \new_[62046]_ , \new_[62047]_ , \new_[62048]_ ,
    \new_[62051]_ , \new_[62054]_ , \new_[62055]_ , \new_[62058]_ ,
    \new_[62061]_ , \new_[62062]_ , \new_[62063]_ , \new_[62066]_ ,
    \new_[62069]_ , \new_[62070]_ , \new_[62073]_ , \new_[62076]_ ,
    \new_[62077]_ , \new_[62078]_ , \new_[62081]_ , \new_[62084]_ ,
    \new_[62085]_ , \new_[62088]_ , \new_[62091]_ , \new_[62092]_ ,
    \new_[62093]_ , \new_[62096]_ , \new_[62099]_ , \new_[62100]_ ,
    \new_[62103]_ , \new_[62106]_ , \new_[62107]_ , \new_[62108]_ ,
    \new_[62111]_ , \new_[62114]_ , \new_[62115]_ , \new_[62118]_ ,
    \new_[62121]_ , \new_[62122]_ , \new_[62123]_ , \new_[62126]_ ,
    \new_[62129]_ , \new_[62130]_ , \new_[62133]_ , \new_[62136]_ ,
    \new_[62137]_ , \new_[62138]_ , \new_[62141]_ , \new_[62144]_ ,
    \new_[62145]_ , \new_[62148]_ , \new_[62151]_ , \new_[62152]_ ,
    \new_[62153]_ , \new_[62156]_ , \new_[62159]_ , \new_[62160]_ ,
    \new_[62163]_ , \new_[62166]_ , \new_[62167]_ , \new_[62168]_ ,
    \new_[62171]_ , \new_[62174]_ , \new_[62175]_ , \new_[62178]_ ,
    \new_[62181]_ , \new_[62182]_ , \new_[62183]_ , \new_[62186]_ ,
    \new_[62189]_ , \new_[62190]_ , \new_[62193]_ , \new_[62196]_ ,
    \new_[62197]_ , \new_[62198]_ , \new_[62201]_ , \new_[62204]_ ,
    \new_[62205]_ , \new_[62208]_ , \new_[62211]_ , \new_[62212]_ ,
    \new_[62213]_ , \new_[62216]_ , \new_[62219]_ , \new_[62220]_ ,
    \new_[62223]_ , \new_[62226]_ , \new_[62227]_ , \new_[62228]_ ,
    \new_[62231]_ , \new_[62234]_ , \new_[62235]_ , \new_[62238]_ ,
    \new_[62241]_ , \new_[62242]_ , \new_[62243]_ , \new_[62246]_ ,
    \new_[62249]_ , \new_[62250]_ , \new_[62253]_ , \new_[62256]_ ,
    \new_[62257]_ , \new_[62258]_ , \new_[62261]_ , \new_[62264]_ ,
    \new_[62265]_ , \new_[62268]_ , \new_[62271]_ , \new_[62272]_ ,
    \new_[62273]_ , \new_[62276]_ , \new_[62279]_ , \new_[62280]_ ,
    \new_[62283]_ , \new_[62286]_ , \new_[62287]_ , \new_[62288]_ ,
    \new_[62291]_ , \new_[62294]_ , \new_[62295]_ , \new_[62298]_ ,
    \new_[62301]_ , \new_[62302]_ , \new_[62303]_ , \new_[62306]_ ,
    \new_[62309]_ , \new_[62310]_ , \new_[62313]_ , \new_[62316]_ ,
    \new_[62317]_ , \new_[62318]_ , \new_[62321]_ , \new_[62324]_ ,
    \new_[62325]_ , \new_[62328]_ , \new_[62331]_ , \new_[62332]_ ,
    \new_[62333]_ , \new_[62336]_ , \new_[62339]_ , \new_[62340]_ ,
    \new_[62343]_ , \new_[62346]_ , \new_[62347]_ , \new_[62348]_ ,
    \new_[62351]_ , \new_[62354]_ , \new_[62355]_ , \new_[62358]_ ,
    \new_[62361]_ , \new_[62362]_ , \new_[62363]_ , \new_[62366]_ ,
    \new_[62369]_ , \new_[62370]_ , \new_[62373]_ , \new_[62376]_ ,
    \new_[62377]_ , \new_[62378]_ , \new_[62381]_ , \new_[62384]_ ,
    \new_[62385]_ , \new_[62388]_ , \new_[62391]_ , \new_[62392]_ ,
    \new_[62393]_ , \new_[62396]_ , \new_[62399]_ , \new_[62400]_ ,
    \new_[62403]_ , \new_[62406]_ , \new_[62407]_ , \new_[62408]_ ,
    \new_[62411]_ , \new_[62414]_ , \new_[62415]_ , \new_[62418]_ ,
    \new_[62421]_ , \new_[62422]_ , \new_[62423]_ , \new_[62426]_ ,
    \new_[62429]_ , \new_[62430]_ , \new_[62433]_ , \new_[62436]_ ,
    \new_[62437]_ , \new_[62438]_ , \new_[62441]_ , \new_[62444]_ ,
    \new_[62445]_ , \new_[62448]_ , \new_[62451]_ , \new_[62452]_ ,
    \new_[62453]_ , \new_[62456]_ , \new_[62459]_ , \new_[62460]_ ,
    \new_[62463]_ , \new_[62466]_ , \new_[62467]_ , \new_[62468]_ ,
    \new_[62471]_ , \new_[62474]_ , \new_[62475]_ , \new_[62478]_ ,
    \new_[62481]_ , \new_[62482]_ , \new_[62483]_ , \new_[62486]_ ,
    \new_[62489]_ , \new_[62490]_ , \new_[62493]_ , \new_[62496]_ ,
    \new_[62497]_ , \new_[62498]_ , \new_[62501]_ , \new_[62504]_ ,
    \new_[62505]_ , \new_[62508]_ , \new_[62511]_ , \new_[62512]_ ,
    \new_[62513]_ , \new_[62516]_ , \new_[62519]_ , \new_[62520]_ ,
    \new_[62523]_ , \new_[62526]_ , \new_[62527]_ , \new_[62528]_ ,
    \new_[62531]_ , \new_[62534]_ , \new_[62535]_ , \new_[62538]_ ,
    \new_[62541]_ , \new_[62542]_ , \new_[62543]_ , \new_[62546]_ ,
    \new_[62549]_ , \new_[62550]_ , \new_[62553]_ , \new_[62556]_ ,
    \new_[62557]_ , \new_[62558]_ , \new_[62561]_ , \new_[62564]_ ,
    \new_[62565]_ , \new_[62568]_ , \new_[62571]_ , \new_[62572]_ ,
    \new_[62573]_ , \new_[62576]_ , \new_[62579]_ , \new_[62580]_ ,
    \new_[62583]_ , \new_[62586]_ , \new_[62587]_ , \new_[62588]_ ,
    \new_[62591]_ , \new_[62594]_ , \new_[62595]_ , \new_[62598]_ ,
    \new_[62601]_ , \new_[62602]_ , \new_[62603]_ , \new_[62606]_ ,
    \new_[62609]_ , \new_[62610]_ , \new_[62613]_ , \new_[62616]_ ,
    \new_[62617]_ , \new_[62618]_ , \new_[62621]_ , \new_[62624]_ ,
    \new_[62625]_ , \new_[62628]_ , \new_[62631]_ , \new_[62632]_ ,
    \new_[62633]_ , \new_[62636]_ , \new_[62639]_ , \new_[62640]_ ,
    \new_[62643]_ , \new_[62646]_ , \new_[62647]_ , \new_[62648]_ ,
    \new_[62651]_ , \new_[62654]_ , \new_[62655]_ , \new_[62658]_ ,
    \new_[62661]_ , \new_[62662]_ , \new_[62663]_ , \new_[62666]_ ,
    \new_[62669]_ , \new_[62670]_ , \new_[62673]_ , \new_[62676]_ ,
    \new_[62677]_ , \new_[62678]_ , \new_[62681]_ , \new_[62684]_ ,
    \new_[62685]_ , \new_[62688]_ , \new_[62691]_ , \new_[62692]_ ,
    \new_[62693]_ , \new_[62696]_ , \new_[62699]_ , \new_[62700]_ ,
    \new_[62703]_ , \new_[62706]_ , \new_[62707]_ , \new_[62708]_ ,
    \new_[62711]_ , \new_[62714]_ , \new_[62715]_ , \new_[62718]_ ,
    \new_[62721]_ , \new_[62722]_ , \new_[62723]_ , \new_[62726]_ ,
    \new_[62729]_ , \new_[62730]_ , \new_[62733]_ , \new_[62736]_ ,
    \new_[62737]_ , \new_[62738]_ , \new_[62741]_ , \new_[62744]_ ,
    \new_[62745]_ , \new_[62748]_ , \new_[62751]_ , \new_[62752]_ ,
    \new_[62753]_ , \new_[62756]_ , \new_[62759]_ , \new_[62760]_ ,
    \new_[62763]_ , \new_[62766]_ , \new_[62767]_ , \new_[62768]_ ,
    \new_[62771]_ , \new_[62774]_ , \new_[62775]_ , \new_[62778]_ ,
    \new_[62781]_ , \new_[62782]_ , \new_[62783]_ , \new_[62786]_ ,
    \new_[62789]_ , \new_[62790]_ , \new_[62793]_ , \new_[62796]_ ,
    \new_[62797]_ , \new_[62798]_ , \new_[62801]_ , \new_[62804]_ ,
    \new_[62805]_ , \new_[62808]_ , \new_[62811]_ , \new_[62812]_ ,
    \new_[62813]_ , \new_[62816]_ , \new_[62819]_ , \new_[62820]_ ,
    \new_[62823]_ , \new_[62826]_ , \new_[62827]_ , \new_[62828]_ ,
    \new_[62831]_ , \new_[62834]_ , \new_[62835]_ , \new_[62838]_ ,
    \new_[62841]_ , \new_[62842]_ , \new_[62843]_ , \new_[62846]_ ,
    \new_[62849]_ , \new_[62850]_ , \new_[62853]_ , \new_[62856]_ ,
    \new_[62857]_ , \new_[62858]_ , \new_[62861]_ , \new_[62864]_ ,
    \new_[62865]_ , \new_[62868]_ , \new_[62871]_ , \new_[62872]_ ,
    \new_[62873]_ , \new_[62876]_ , \new_[62879]_ , \new_[62880]_ ,
    \new_[62883]_ , \new_[62886]_ , \new_[62887]_ , \new_[62888]_ ,
    \new_[62891]_ , \new_[62894]_ , \new_[62895]_ , \new_[62898]_ ,
    \new_[62901]_ , \new_[62902]_ , \new_[62903]_ , \new_[62906]_ ,
    \new_[62909]_ , \new_[62910]_ , \new_[62913]_ , \new_[62916]_ ,
    \new_[62917]_ , \new_[62918]_ , \new_[62921]_ , \new_[62924]_ ,
    \new_[62925]_ , \new_[62928]_ , \new_[62931]_ , \new_[62932]_ ,
    \new_[62933]_ , \new_[62936]_ , \new_[62939]_ , \new_[62940]_ ,
    \new_[62943]_ , \new_[62946]_ , \new_[62947]_ , \new_[62948]_ ,
    \new_[62951]_ , \new_[62954]_ , \new_[62955]_ , \new_[62958]_ ,
    \new_[62961]_ , \new_[62962]_ , \new_[62963]_ , \new_[62966]_ ,
    \new_[62969]_ , \new_[62970]_ , \new_[62973]_ , \new_[62976]_ ,
    \new_[62977]_ , \new_[62978]_ , \new_[62981]_ , \new_[62984]_ ,
    \new_[62985]_ , \new_[62988]_ , \new_[62991]_ , \new_[62992]_ ,
    \new_[62993]_ , \new_[62996]_ , \new_[62999]_ , \new_[63000]_ ,
    \new_[63003]_ , \new_[63006]_ , \new_[63007]_ , \new_[63008]_ ,
    \new_[63011]_ , \new_[63014]_ , \new_[63015]_ , \new_[63018]_ ,
    \new_[63021]_ , \new_[63022]_ , \new_[63023]_ , \new_[63026]_ ,
    \new_[63029]_ , \new_[63030]_ , \new_[63033]_ , \new_[63036]_ ,
    \new_[63037]_ , \new_[63038]_ , \new_[63041]_ , \new_[63044]_ ,
    \new_[63045]_ , \new_[63048]_ , \new_[63051]_ , \new_[63052]_ ,
    \new_[63053]_ , \new_[63056]_ , \new_[63059]_ , \new_[63060]_ ,
    \new_[63063]_ , \new_[63066]_ , \new_[63067]_ , \new_[63068]_ ,
    \new_[63071]_ , \new_[63074]_ , \new_[63075]_ , \new_[63078]_ ,
    \new_[63081]_ , \new_[63082]_ , \new_[63083]_ , \new_[63086]_ ,
    \new_[63089]_ , \new_[63090]_ , \new_[63093]_ , \new_[63096]_ ,
    \new_[63097]_ , \new_[63098]_ , \new_[63101]_ , \new_[63104]_ ,
    \new_[63105]_ , \new_[63108]_ , \new_[63111]_ , \new_[63112]_ ,
    \new_[63113]_ , \new_[63116]_ , \new_[63119]_ , \new_[63120]_ ,
    \new_[63123]_ , \new_[63126]_ , \new_[63127]_ , \new_[63128]_ ,
    \new_[63131]_ , \new_[63134]_ , \new_[63135]_ , \new_[63138]_ ,
    \new_[63141]_ , \new_[63142]_ , \new_[63143]_ , \new_[63146]_ ,
    \new_[63149]_ , \new_[63150]_ , \new_[63153]_ , \new_[63156]_ ,
    \new_[63157]_ , \new_[63158]_ , \new_[63161]_ , \new_[63164]_ ,
    \new_[63165]_ , \new_[63168]_ , \new_[63171]_ , \new_[63172]_ ,
    \new_[63173]_ , \new_[63176]_ , \new_[63179]_ , \new_[63180]_ ,
    \new_[63183]_ , \new_[63186]_ , \new_[63187]_ , \new_[63188]_ ,
    \new_[63191]_ , \new_[63194]_ , \new_[63195]_ , \new_[63198]_ ,
    \new_[63201]_ , \new_[63202]_ , \new_[63203]_ , \new_[63206]_ ,
    \new_[63209]_ , \new_[63210]_ , \new_[63213]_ , \new_[63216]_ ,
    \new_[63217]_ , \new_[63218]_ , \new_[63221]_ , \new_[63224]_ ,
    \new_[63225]_ , \new_[63228]_ , \new_[63231]_ , \new_[63232]_ ,
    \new_[63233]_ , \new_[63236]_ , \new_[63239]_ , \new_[63240]_ ,
    \new_[63243]_ , \new_[63246]_ , \new_[63247]_ , \new_[63248]_ ,
    \new_[63251]_ , \new_[63254]_ , \new_[63255]_ , \new_[63258]_ ,
    \new_[63261]_ , \new_[63262]_ , \new_[63263]_ , \new_[63266]_ ,
    \new_[63269]_ , \new_[63270]_ , \new_[63273]_ , \new_[63276]_ ,
    \new_[63277]_ , \new_[63278]_ , \new_[63281]_ , \new_[63284]_ ,
    \new_[63285]_ , \new_[63288]_ , \new_[63291]_ , \new_[63292]_ ,
    \new_[63293]_ , \new_[63296]_ , \new_[63299]_ , \new_[63300]_ ,
    \new_[63303]_ , \new_[63306]_ , \new_[63307]_ , \new_[63308]_ ,
    \new_[63311]_ , \new_[63314]_ , \new_[63315]_ , \new_[63318]_ ,
    \new_[63321]_ , \new_[63322]_ , \new_[63323]_ , \new_[63326]_ ,
    \new_[63329]_ , \new_[63330]_ , \new_[63333]_ , \new_[63336]_ ,
    \new_[63337]_ , \new_[63338]_ , \new_[63341]_ , \new_[63344]_ ,
    \new_[63345]_ , \new_[63348]_ , \new_[63351]_ , \new_[63352]_ ,
    \new_[63353]_ , \new_[63356]_ , \new_[63359]_ , \new_[63360]_ ,
    \new_[63363]_ , \new_[63366]_ , \new_[63367]_ , \new_[63368]_ ,
    \new_[63371]_ , \new_[63374]_ , \new_[63375]_ , \new_[63378]_ ,
    \new_[63381]_ , \new_[63382]_ , \new_[63383]_ , \new_[63386]_ ,
    \new_[63389]_ , \new_[63390]_ , \new_[63393]_ , \new_[63396]_ ,
    \new_[63397]_ , \new_[63398]_ , \new_[63401]_ , \new_[63404]_ ,
    \new_[63405]_ , \new_[63408]_ , \new_[63411]_ , \new_[63412]_ ,
    \new_[63413]_ , \new_[63416]_ , \new_[63419]_ , \new_[63420]_ ,
    \new_[63423]_ , \new_[63426]_ , \new_[63427]_ , \new_[63428]_ ,
    \new_[63431]_ , \new_[63434]_ , \new_[63435]_ , \new_[63438]_ ,
    \new_[63441]_ , \new_[63442]_ , \new_[63443]_ , \new_[63446]_ ,
    \new_[63449]_ , \new_[63450]_ , \new_[63453]_ , \new_[63456]_ ,
    \new_[63457]_ , \new_[63458]_ , \new_[63461]_ , \new_[63464]_ ,
    \new_[63465]_ , \new_[63468]_ , \new_[63471]_ , \new_[63472]_ ,
    \new_[63473]_ , \new_[63476]_ , \new_[63479]_ , \new_[63480]_ ,
    \new_[63483]_ , \new_[63486]_ , \new_[63487]_ , \new_[63488]_ ,
    \new_[63491]_ , \new_[63494]_ , \new_[63495]_ , \new_[63498]_ ,
    \new_[63501]_ , \new_[63502]_ , \new_[63503]_ , \new_[63506]_ ,
    \new_[63509]_ , \new_[63510]_ , \new_[63513]_ , \new_[63516]_ ,
    \new_[63517]_ , \new_[63518]_ , \new_[63521]_ , \new_[63524]_ ,
    \new_[63525]_ , \new_[63528]_ , \new_[63531]_ , \new_[63532]_ ,
    \new_[63533]_ , \new_[63536]_ , \new_[63539]_ , \new_[63540]_ ,
    \new_[63543]_ , \new_[63546]_ , \new_[63547]_ , \new_[63548]_ ,
    \new_[63551]_ , \new_[63554]_ , \new_[63555]_ , \new_[63558]_ ,
    \new_[63561]_ , \new_[63562]_ , \new_[63563]_ , \new_[63566]_ ,
    \new_[63569]_ , \new_[63570]_ , \new_[63573]_ , \new_[63576]_ ,
    \new_[63577]_ , \new_[63578]_ , \new_[63581]_ , \new_[63584]_ ,
    \new_[63585]_ , \new_[63588]_ , \new_[63591]_ , \new_[63592]_ ,
    \new_[63593]_ , \new_[63596]_ , \new_[63599]_ , \new_[63600]_ ,
    \new_[63603]_ , \new_[63606]_ , \new_[63607]_ , \new_[63608]_ ,
    \new_[63611]_ , \new_[63614]_ , \new_[63615]_ , \new_[63618]_ ,
    \new_[63621]_ , \new_[63622]_ , \new_[63623]_ , \new_[63626]_ ,
    \new_[63629]_ , \new_[63630]_ , \new_[63633]_ , \new_[63636]_ ,
    \new_[63637]_ , \new_[63638]_ , \new_[63641]_ , \new_[63644]_ ,
    \new_[63645]_ , \new_[63648]_ , \new_[63651]_ , \new_[63652]_ ,
    \new_[63653]_ , \new_[63656]_ , \new_[63659]_ , \new_[63660]_ ,
    \new_[63663]_ , \new_[63666]_ , \new_[63667]_ , \new_[63668]_ ,
    \new_[63671]_ , \new_[63674]_ , \new_[63675]_ , \new_[63678]_ ,
    \new_[63681]_ , \new_[63682]_ , \new_[63683]_ , \new_[63686]_ ,
    \new_[63689]_ , \new_[63690]_ , \new_[63693]_ , \new_[63696]_ ,
    \new_[63697]_ , \new_[63698]_ , \new_[63701]_ , \new_[63704]_ ,
    \new_[63705]_ , \new_[63708]_ , \new_[63711]_ , \new_[63712]_ ,
    \new_[63713]_ , \new_[63716]_ , \new_[63719]_ , \new_[63720]_ ,
    \new_[63723]_ , \new_[63726]_ , \new_[63727]_ , \new_[63728]_ ,
    \new_[63731]_ , \new_[63734]_ , \new_[63735]_ , \new_[63738]_ ,
    \new_[63741]_ , \new_[63742]_ , \new_[63743]_ , \new_[63746]_ ,
    \new_[63749]_ , \new_[63750]_ , \new_[63753]_ , \new_[63756]_ ,
    \new_[63757]_ , \new_[63758]_ , \new_[63761]_ , \new_[63764]_ ,
    \new_[63765]_ , \new_[63768]_ , \new_[63771]_ , \new_[63772]_ ,
    \new_[63773]_ , \new_[63776]_ , \new_[63779]_ , \new_[63780]_ ,
    \new_[63783]_ , \new_[63786]_ , \new_[63787]_ , \new_[63788]_ ,
    \new_[63791]_ , \new_[63794]_ , \new_[63795]_ , \new_[63798]_ ,
    \new_[63801]_ , \new_[63802]_ , \new_[63803]_ , \new_[63806]_ ,
    \new_[63809]_ , \new_[63810]_ , \new_[63813]_ , \new_[63816]_ ,
    \new_[63817]_ , \new_[63818]_ , \new_[63821]_ , \new_[63824]_ ,
    \new_[63825]_ , \new_[63828]_ , \new_[63831]_ , \new_[63832]_ ,
    \new_[63833]_ , \new_[63836]_ , \new_[63839]_ , \new_[63840]_ ,
    \new_[63843]_ , \new_[63846]_ , \new_[63847]_ , \new_[63848]_ ,
    \new_[63851]_ , \new_[63854]_ , \new_[63855]_ , \new_[63858]_ ,
    \new_[63861]_ , \new_[63862]_ , \new_[63863]_ , \new_[63866]_ ,
    \new_[63869]_ , \new_[63870]_ , \new_[63873]_ , \new_[63876]_ ,
    \new_[63877]_ , \new_[63878]_ , \new_[63881]_ , \new_[63884]_ ,
    \new_[63885]_ , \new_[63888]_ , \new_[63891]_ , \new_[63892]_ ,
    \new_[63893]_ , \new_[63896]_ , \new_[63899]_ , \new_[63900]_ ,
    \new_[63903]_ , \new_[63906]_ , \new_[63907]_ , \new_[63908]_ ,
    \new_[63911]_ , \new_[63914]_ , \new_[63915]_ , \new_[63918]_ ,
    \new_[63921]_ , \new_[63922]_ , \new_[63923]_ , \new_[63926]_ ,
    \new_[63929]_ , \new_[63930]_ , \new_[63933]_ , \new_[63936]_ ,
    \new_[63937]_ , \new_[63938]_ , \new_[63941]_ , \new_[63944]_ ,
    \new_[63945]_ , \new_[63948]_ , \new_[63951]_ , \new_[63952]_ ,
    \new_[63953]_ , \new_[63956]_ , \new_[63959]_ , \new_[63960]_ ,
    \new_[63963]_ , \new_[63966]_ , \new_[63967]_ , \new_[63968]_ ,
    \new_[63971]_ , \new_[63974]_ , \new_[63975]_ , \new_[63978]_ ,
    \new_[63981]_ , \new_[63982]_ , \new_[63983]_ , \new_[63986]_ ,
    \new_[63989]_ , \new_[63990]_ , \new_[63993]_ , \new_[63997]_ ,
    \new_[63998]_ , \new_[63999]_ , \new_[64000]_ , \new_[64003]_ ,
    \new_[64006]_ , \new_[64007]_ , \new_[64010]_ , \new_[64013]_ ,
    \new_[64014]_ , \new_[64015]_ , \new_[64018]_ , \new_[64021]_ ,
    \new_[64022]_ , \new_[64025]_ , \new_[64029]_ , \new_[64030]_ ,
    \new_[64031]_ , \new_[64032]_ , \new_[64035]_ , \new_[64038]_ ,
    \new_[64039]_ , \new_[64042]_ , \new_[64045]_ , \new_[64046]_ ,
    \new_[64047]_ , \new_[64050]_ , \new_[64053]_ , \new_[64054]_ ,
    \new_[64057]_ , \new_[64061]_ , \new_[64062]_ , \new_[64063]_ ,
    \new_[64064]_ , \new_[64067]_ , \new_[64070]_ , \new_[64071]_ ,
    \new_[64074]_ , \new_[64077]_ , \new_[64078]_ , \new_[64079]_ ,
    \new_[64082]_ , \new_[64085]_ , \new_[64086]_ , \new_[64089]_ ,
    \new_[64093]_ , \new_[64094]_ , \new_[64095]_ , \new_[64096]_ ,
    \new_[64099]_ , \new_[64102]_ , \new_[64103]_ , \new_[64106]_ ,
    \new_[64109]_ , \new_[64110]_ , \new_[64111]_ , \new_[64114]_ ,
    \new_[64117]_ , \new_[64118]_ , \new_[64121]_ , \new_[64125]_ ,
    \new_[64126]_ , \new_[64127]_ , \new_[64128]_ , \new_[64131]_ ,
    \new_[64134]_ , \new_[64135]_ , \new_[64138]_ , \new_[64141]_ ,
    \new_[64142]_ , \new_[64143]_ , \new_[64146]_ , \new_[64149]_ ,
    \new_[64150]_ , \new_[64153]_ , \new_[64157]_ , \new_[64158]_ ,
    \new_[64159]_ , \new_[64160]_ , \new_[64163]_ , \new_[64166]_ ,
    \new_[64167]_ , \new_[64170]_ , \new_[64173]_ , \new_[64174]_ ,
    \new_[64175]_ , \new_[64178]_ , \new_[64181]_ , \new_[64182]_ ,
    \new_[64185]_ , \new_[64189]_ , \new_[64190]_ , \new_[64191]_ ,
    \new_[64192]_ , \new_[64195]_ , \new_[64198]_ , \new_[64199]_ ,
    \new_[64202]_ , \new_[64205]_ , \new_[64206]_ , \new_[64207]_ ,
    \new_[64210]_ , \new_[64213]_ , \new_[64214]_ , \new_[64217]_ ,
    \new_[64221]_ , \new_[64222]_ , \new_[64223]_ , \new_[64224]_ ,
    \new_[64227]_ , \new_[64230]_ , \new_[64231]_ , \new_[64234]_ ,
    \new_[64237]_ , \new_[64238]_ , \new_[64239]_ , \new_[64242]_ ,
    \new_[64245]_ , \new_[64246]_ , \new_[64249]_ , \new_[64253]_ ,
    \new_[64254]_ , \new_[64255]_ , \new_[64256]_ , \new_[64259]_ ,
    \new_[64262]_ , \new_[64263]_ , \new_[64266]_ , \new_[64269]_ ,
    \new_[64270]_ , \new_[64271]_ , \new_[64274]_ , \new_[64277]_ ,
    \new_[64278]_ , \new_[64281]_ , \new_[64285]_ , \new_[64286]_ ,
    \new_[64287]_ , \new_[64288]_ , \new_[64291]_ , \new_[64294]_ ,
    \new_[64295]_ , \new_[64298]_ , \new_[64301]_ , \new_[64302]_ ,
    \new_[64303]_ , \new_[64306]_ , \new_[64309]_ , \new_[64310]_ ,
    \new_[64313]_ , \new_[64317]_ , \new_[64318]_ , \new_[64319]_ ,
    \new_[64320]_ , \new_[64323]_ , \new_[64326]_ , \new_[64327]_ ,
    \new_[64330]_ , \new_[64333]_ , \new_[64334]_ , \new_[64335]_ ,
    \new_[64338]_ , \new_[64341]_ , \new_[64342]_ , \new_[64345]_ ,
    \new_[64349]_ , \new_[64350]_ , \new_[64351]_ , \new_[64352]_ ,
    \new_[64355]_ , \new_[64358]_ , \new_[64359]_ , \new_[64362]_ ,
    \new_[64365]_ , \new_[64366]_ , \new_[64367]_ , \new_[64370]_ ,
    \new_[64373]_ , \new_[64374]_ , \new_[64377]_ , \new_[64381]_ ,
    \new_[64382]_ , \new_[64383]_ , \new_[64384]_ , \new_[64387]_ ,
    \new_[64390]_ , \new_[64391]_ , \new_[64394]_ , \new_[64397]_ ,
    \new_[64398]_ , \new_[64399]_ , \new_[64402]_ , \new_[64405]_ ,
    \new_[64406]_ , \new_[64409]_ , \new_[64413]_ , \new_[64414]_ ,
    \new_[64415]_ , \new_[64416]_ , \new_[64419]_ , \new_[64422]_ ,
    \new_[64423]_ , \new_[64426]_ , \new_[64429]_ , \new_[64430]_ ,
    \new_[64431]_ , \new_[64434]_ , \new_[64437]_ , \new_[64438]_ ,
    \new_[64441]_ , \new_[64445]_ , \new_[64446]_ , \new_[64447]_ ,
    \new_[64448]_ , \new_[64451]_ , \new_[64454]_ , \new_[64455]_ ,
    \new_[64458]_ , \new_[64461]_ , \new_[64462]_ , \new_[64463]_ ,
    \new_[64466]_ , \new_[64469]_ , \new_[64470]_ , \new_[64473]_ ,
    \new_[64477]_ , \new_[64478]_ , \new_[64479]_ , \new_[64480]_ ,
    \new_[64483]_ , \new_[64486]_ , \new_[64487]_ , \new_[64490]_ ,
    \new_[64493]_ , \new_[64494]_ , \new_[64495]_ , \new_[64498]_ ,
    \new_[64501]_ , \new_[64502]_ , \new_[64505]_ , \new_[64509]_ ,
    \new_[64510]_ , \new_[64511]_ , \new_[64512]_ , \new_[64515]_ ,
    \new_[64518]_ , \new_[64519]_ , \new_[64522]_ , \new_[64525]_ ,
    \new_[64526]_ , \new_[64527]_ , \new_[64530]_ , \new_[64533]_ ,
    \new_[64534]_ , \new_[64537]_ , \new_[64541]_ , \new_[64542]_ ,
    \new_[64543]_ , \new_[64544]_ , \new_[64547]_ , \new_[64550]_ ,
    \new_[64551]_ , \new_[64554]_ , \new_[64557]_ , \new_[64558]_ ,
    \new_[64559]_ , \new_[64562]_ , \new_[64565]_ , \new_[64566]_ ,
    \new_[64569]_ , \new_[64573]_ , \new_[64574]_ , \new_[64575]_ ,
    \new_[64576]_ , \new_[64579]_ , \new_[64582]_ , \new_[64583]_ ,
    \new_[64586]_ , \new_[64589]_ , \new_[64590]_ , \new_[64591]_ ,
    \new_[64594]_ , \new_[64597]_ , \new_[64598]_ , \new_[64601]_ ,
    \new_[64605]_ , \new_[64606]_ , \new_[64607]_ , \new_[64608]_ ,
    \new_[64611]_ , \new_[64614]_ , \new_[64615]_ , \new_[64618]_ ,
    \new_[64621]_ , \new_[64622]_ , \new_[64623]_ , \new_[64626]_ ,
    \new_[64629]_ , \new_[64630]_ , \new_[64633]_ , \new_[64637]_ ,
    \new_[64638]_ , \new_[64639]_ , \new_[64640]_ , \new_[64643]_ ,
    \new_[64646]_ , \new_[64647]_ , \new_[64650]_ , \new_[64653]_ ,
    \new_[64654]_ , \new_[64655]_ , \new_[64658]_ , \new_[64661]_ ,
    \new_[64662]_ , \new_[64665]_ , \new_[64669]_ , \new_[64670]_ ,
    \new_[64671]_ , \new_[64672]_ , \new_[64675]_ , \new_[64678]_ ,
    \new_[64679]_ , \new_[64682]_ , \new_[64685]_ , \new_[64686]_ ,
    \new_[64687]_ , \new_[64690]_ , \new_[64693]_ , \new_[64694]_ ,
    \new_[64697]_ , \new_[64701]_ , \new_[64702]_ , \new_[64703]_ ,
    \new_[64704]_ , \new_[64707]_ , \new_[64710]_ , \new_[64711]_ ,
    \new_[64714]_ , \new_[64717]_ , \new_[64718]_ , \new_[64719]_ ,
    \new_[64722]_ , \new_[64725]_ , \new_[64726]_ , \new_[64729]_ ,
    \new_[64733]_ , \new_[64734]_ , \new_[64735]_ , \new_[64736]_ ,
    \new_[64739]_ , \new_[64742]_ , \new_[64743]_ , \new_[64746]_ ,
    \new_[64749]_ , \new_[64750]_ , \new_[64751]_ , \new_[64754]_ ,
    \new_[64757]_ , \new_[64758]_ , \new_[64761]_ , \new_[64765]_ ,
    \new_[64766]_ , \new_[64767]_ , \new_[64768]_ , \new_[64771]_ ,
    \new_[64774]_ , \new_[64775]_ , \new_[64778]_ , \new_[64781]_ ,
    \new_[64782]_ , \new_[64783]_ , \new_[64786]_ , \new_[64789]_ ,
    \new_[64790]_ , \new_[64793]_ , \new_[64797]_ , \new_[64798]_ ,
    \new_[64799]_ , \new_[64800]_ , \new_[64803]_ , \new_[64806]_ ,
    \new_[64807]_ , \new_[64810]_ , \new_[64813]_ , \new_[64814]_ ,
    \new_[64815]_ , \new_[64818]_ , \new_[64821]_ , \new_[64822]_ ,
    \new_[64825]_ , \new_[64829]_ , \new_[64830]_ , \new_[64831]_ ,
    \new_[64832]_ , \new_[64835]_ , \new_[64838]_ , \new_[64839]_ ,
    \new_[64842]_ , \new_[64845]_ , \new_[64846]_ , \new_[64847]_ ,
    \new_[64850]_ , \new_[64853]_ , \new_[64854]_ , \new_[64857]_ ,
    \new_[64861]_ , \new_[64862]_ , \new_[64863]_ , \new_[64864]_ ,
    \new_[64867]_ , \new_[64870]_ , \new_[64871]_ , \new_[64874]_ ,
    \new_[64877]_ , \new_[64878]_ , \new_[64879]_ , \new_[64882]_ ,
    \new_[64885]_ , \new_[64886]_ , \new_[64889]_ , \new_[64893]_ ,
    \new_[64894]_ , \new_[64895]_ , \new_[64896]_ , \new_[64899]_ ,
    \new_[64902]_ , \new_[64903]_ , \new_[64906]_ , \new_[64909]_ ,
    \new_[64910]_ , \new_[64911]_ , \new_[64914]_ , \new_[64917]_ ,
    \new_[64918]_ , \new_[64921]_ , \new_[64925]_ , \new_[64926]_ ,
    \new_[64927]_ , \new_[64928]_ , \new_[64931]_ , \new_[64934]_ ,
    \new_[64935]_ , \new_[64938]_ , \new_[64941]_ , \new_[64942]_ ,
    \new_[64943]_ , \new_[64946]_ , \new_[64949]_ , \new_[64950]_ ,
    \new_[64953]_ , \new_[64957]_ , \new_[64958]_ , \new_[64959]_ ,
    \new_[64960]_ , \new_[64963]_ , \new_[64966]_ , \new_[64967]_ ,
    \new_[64970]_ , \new_[64973]_ , \new_[64974]_ , \new_[64975]_ ,
    \new_[64978]_ , \new_[64981]_ , \new_[64982]_ , \new_[64985]_ ,
    \new_[64989]_ , \new_[64990]_ , \new_[64991]_ , \new_[64992]_ ,
    \new_[64995]_ , \new_[64998]_ , \new_[64999]_ , \new_[65002]_ ,
    \new_[65005]_ , \new_[65006]_ , \new_[65007]_ , \new_[65010]_ ,
    \new_[65013]_ , \new_[65014]_ , \new_[65017]_ , \new_[65021]_ ,
    \new_[65022]_ , \new_[65023]_ , \new_[65024]_ , \new_[65027]_ ,
    \new_[65030]_ , \new_[65031]_ , \new_[65034]_ , \new_[65037]_ ,
    \new_[65038]_ , \new_[65039]_ , \new_[65042]_ , \new_[65045]_ ,
    \new_[65046]_ , \new_[65049]_ , \new_[65053]_ , \new_[65054]_ ,
    \new_[65055]_ , \new_[65056]_ , \new_[65059]_ , \new_[65062]_ ,
    \new_[65063]_ , \new_[65066]_ , \new_[65069]_ , \new_[65070]_ ,
    \new_[65071]_ , \new_[65074]_ , \new_[65077]_ , \new_[65078]_ ,
    \new_[65081]_ , \new_[65085]_ , \new_[65086]_ , \new_[65087]_ ,
    \new_[65088]_ , \new_[65091]_ , \new_[65094]_ , \new_[65095]_ ,
    \new_[65098]_ , \new_[65101]_ , \new_[65102]_ , \new_[65103]_ ,
    \new_[65106]_ , \new_[65109]_ , \new_[65110]_ , \new_[65113]_ ,
    \new_[65117]_ , \new_[65118]_ , \new_[65119]_ , \new_[65120]_ ,
    \new_[65123]_ , \new_[65126]_ , \new_[65127]_ , \new_[65130]_ ,
    \new_[65133]_ , \new_[65134]_ , \new_[65135]_ , \new_[65138]_ ,
    \new_[65141]_ , \new_[65142]_ , \new_[65145]_ , \new_[65149]_ ,
    \new_[65150]_ , \new_[65151]_ , \new_[65152]_ , \new_[65155]_ ,
    \new_[65158]_ , \new_[65159]_ , \new_[65162]_ , \new_[65165]_ ,
    \new_[65166]_ , \new_[65167]_ , \new_[65170]_ , \new_[65173]_ ,
    \new_[65174]_ , \new_[65177]_ , \new_[65181]_ , \new_[65182]_ ,
    \new_[65183]_ , \new_[65184]_ , \new_[65187]_ , \new_[65190]_ ,
    \new_[65191]_ , \new_[65194]_ , \new_[65197]_ , \new_[65198]_ ,
    \new_[65199]_ , \new_[65202]_ , \new_[65205]_ , \new_[65206]_ ,
    \new_[65209]_ , \new_[65213]_ , \new_[65214]_ , \new_[65215]_ ,
    \new_[65216]_ , \new_[65219]_ , \new_[65222]_ , \new_[65223]_ ,
    \new_[65226]_ , \new_[65229]_ , \new_[65230]_ , \new_[65231]_ ,
    \new_[65234]_ , \new_[65237]_ , \new_[65238]_ , \new_[65241]_ ,
    \new_[65245]_ , \new_[65246]_ , \new_[65247]_ , \new_[65248]_ ,
    \new_[65251]_ , \new_[65254]_ , \new_[65255]_ , \new_[65258]_ ,
    \new_[65261]_ , \new_[65262]_ , \new_[65263]_ , \new_[65266]_ ,
    \new_[65269]_ , \new_[65270]_ , \new_[65273]_ , \new_[65277]_ ,
    \new_[65278]_ , \new_[65279]_ , \new_[65280]_ , \new_[65283]_ ,
    \new_[65286]_ , \new_[65287]_ , \new_[65290]_ , \new_[65293]_ ,
    \new_[65294]_ , \new_[65295]_ , \new_[65298]_ , \new_[65301]_ ,
    \new_[65302]_ , \new_[65305]_ , \new_[65309]_ , \new_[65310]_ ,
    \new_[65311]_ , \new_[65312]_ , \new_[65315]_ , \new_[65318]_ ,
    \new_[65319]_ , \new_[65322]_ , \new_[65325]_ , \new_[65326]_ ,
    \new_[65327]_ , \new_[65330]_ , \new_[65333]_ , \new_[65334]_ ,
    \new_[65337]_ , \new_[65341]_ , \new_[65342]_ , \new_[65343]_ ,
    \new_[65344]_ , \new_[65347]_ , \new_[65350]_ , \new_[65351]_ ,
    \new_[65354]_ , \new_[65357]_ , \new_[65358]_ , \new_[65359]_ ,
    \new_[65362]_ , \new_[65365]_ , \new_[65366]_ , \new_[65369]_ ,
    \new_[65373]_ , \new_[65374]_ , \new_[65375]_ , \new_[65376]_ ,
    \new_[65379]_ , \new_[65382]_ , \new_[65383]_ , \new_[65386]_ ,
    \new_[65389]_ , \new_[65390]_ , \new_[65391]_ , \new_[65394]_ ,
    \new_[65397]_ , \new_[65398]_ , \new_[65401]_ , \new_[65405]_ ,
    \new_[65406]_ , \new_[65407]_ , \new_[65408]_ , \new_[65411]_ ,
    \new_[65414]_ , \new_[65415]_ , \new_[65418]_ , \new_[65421]_ ,
    \new_[65422]_ , \new_[65423]_ , \new_[65426]_ , \new_[65429]_ ,
    \new_[65430]_ , \new_[65433]_ , \new_[65437]_ , \new_[65438]_ ,
    \new_[65439]_ , \new_[65440]_ , \new_[65443]_ , \new_[65446]_ ,
    \new_[65447]_ , \new_[65450]_ , \new_[65453]_ , \new_[65454]_ ,
    \new_[65455]_ , \new_[65458]_ , \new_[65461]_ , \new_[65462]_ ,
    \new_[65465]_ , \new_[65469]_ , \new_[65470]_ , \new_[65471]_ ,
    \new_[65472]_ , \new_[65475]_ , \new_[65478]_ , \new_[65479]_ ,
    \new_[65482]_ , \new_[65485]_ , \new_[65486]_ , \new_[65487]_ ,
    \new_[65490]_ , \new_[65493]_ , \new_[65494]_ , \new_[65497]_ ,
    \new_[65501]_ , \new_[65502]_ , \new_[65503]_ , \new_[65504]_ ,
    \new_[65507]_ , \new_[65510]_ , \new_[65511]_ , \new_[65514]_ ,
    \new_[65517]_ , \new_[65518]_ , \new_[65519]_ , \new_[65522]_ ,
    \new_[65525]_ , \new_[65526]_ , \new_[65529]_ , \new_[65533]_ ,
    \new_[65534]_ , \new_[65535]_ , \new_[65536]_ , \new_[65539]_ ,
    \new_[65542]_ , \new_[65543]_ , \new_[65546]_ , \new_[65549]_ ,
    \new_[65550]_ , \new_[65551]_ , \new_[65554]_ , \new_[65557]_ ,
    \new_[65558]_ , \new_[65561]_ , \new_[65565]_ , \new_[65566]_ ,
    \new_[65567]_ , \new_[65568]_ , \new_[65571]_ , \new_[65574]_ ,
    \new_[65575]_ , \new_[65578]_ , \new_[65581]_ , \new_[65582]_ ,
    \new_[65583]_ , \new_[65586]_ , \new_[65589]_ , \new_[65590]_ ,
    \new_[65593]_ , \new_[65597]_ , \new_[65598]_ , \new_[65599]_ ,
    \new_[65600]_ , \new_[65603]_ , \new_[65606]_ , \new_[65607]_ ,
    \new_[65610]_ , \new_[65613]_ , \new_[65614]_ , \new_[65615]_ ,
    \new_[65618]_ , \new_[65621]_ , \new_[65622]_ , \new_[65625]_ ,
    \new_[65629]_ , \new_[65630]_ , \new_[65631]_ , \new_[65632]_ ,
    \new_[65635]_ , \new_[65638]_ , \new_[65639]_ , \new_[65642]_ ,
    \new_[65645]_ , \new_[65646]_ , \new_[65647]_ , \new_[65650]_ ,
    \new_[65653]_ , \new_[65654]_ , \new_[65657]_ , \new_[65661]_ ,
    \new_[65662]_ , \new_[65663]_ , \new_[65664]_ , \new_[65667]_ ,
    \new_[65670]_ , \new_[65671]_ , \new_[65674]_ , \new_[65677]_ ,
    \new_[65678]_ , \new_[65679]_ , \new_[65682]_ , \new_[65685]_ ,
    \new_[65686]_ , \new_[65689]_ , \new_[65693]_ , \new_[65694]_ ,
    \new_[65695]_ , \new_[65696]_ , \new_[65699]_ , \new_[65702]_ ,
    \new_[65703]_ , \new_[65706]_ , \new_[65709]_ , \new_[65710]_ ,
    \new_[65711]_ , \new_[65714]_ , \new_[65717]_ , \new_[65718]_ ,
    \new_[65721]_ , \new_[65725]_ , \new_[65726]_ , \new_[65727]_ ,
    \new_[65728]_ , \new_[65731]_ , \new_[65734]_ , \new_[65735]_ ,
    \new_[65738]_ , \new_[65741]_ , \new_[65742]_ , \new_[65743]_ ,
    \new_[65746]_ , \new_[65749]_ , \new_[65750]_ , \new_[65753]_ ,
    \new_[65757]_ , \new_[65758]_ , \new_[65759]_ , \new_[65760]_ ,
    \new_[65763]_ , \new_[65766]_ , \new_[65767]_ , \new_[65770]_ ,
    \new_[65773]_ , \new_[65774]_ , \new_[65775]_ , \new_[65778]_ ,
    \new_[65781]_ , \new_[65782]_ , \new_[65785]_ , \new_[65789]_ ,
    \new_[65790]_ , \new_[65791]_ , \new_[65792]_ , \new_[65795]_ ,
    \new_[65798]_ , \new_[65799]_ , \new_[65802]_ , \new_[65805]_ ,
    \new_[65806]_ , \new_[65807]_ , \new_[65810]_ , \new_[65813]_ ,
    \new_[65814]_ , \new_[65817]_ , \new_[65821]_ , \new_[65822]_ ,
    \new_[65823]_ , \new_[65824]_ , \new_[65827]_ , \new_[65830]_ ,
    \new_[65831]_ , \new_[65834]_ , \new_[65837]_ , \new_[65838]_ ,
    \new_[65839]_ , \new_[65842]_ , \new_[65845]_ , \new_[65846]_ ,
    \new_[65849]_ , \new_[65853]_ , \new_[65854]_ , \new_[65855]_ ,
    \new_[65856]_ , \new_[65859]_ , \new_[65862]_ , \new_[65863]_ ,
    \new_[65866]_ , \new_[65869]_ , \new_[65870]_ , \new_[65871]_ ,
    \new_[65874]_ , \new_[65877]_ , \new_[65878]_ , \new_[65881]_ ,
    \new_[65885]_ , \new_[65886]_ , \new_[65887]_ , \new_[65888]_ ,
    \new_[65891]_ , \new_[65894]_ , \new_[65895]_ , \new_[65898]_ ,
    \new_[65901]_ , \new_[65902]_ , \new_[65903]_ , \new_[65906]_ ,
    \new_[65909]_ , \new_[65910]_ , \new_[65913]_ , \new_[65917]_ ,
    \new_[65918]_ , \new_[65919]_ , \new_[65920]_ , \new_[65923]_ ,
    \new_[65926]_ , \new_[65927]_ , \new_[65930]_ , \new_[65933]_ ,
    \new_[65934]_ , \new_[65935]_ , \new_[65938]_ , \new_[65941]_ ,
    \new_[65942]_ , \new_[65945]_ , \new_[65949]_ , \new_[65950]_ ,
    \new_[65951]_ , \new_[65952]_ , \new_[65955]_ , \new_[65958]_ ,
    \new_[65959]_ , \new_[65962]_ , \new_[65965]_ , \new_[65966]_ ,
    \new_[65967]_ , \new_[65970]_ , \new_[65973]_ , \new_[65974]_ ,
    \new_[65977]_ , \new_[65981]_ , \new_[65982]_ , \new_[65983]_ ,
    \new_[65984]_ , \new_[65987]_ , \new_[65990]_ , \new_[65991]_ ,
    \new_[65994]_ , \new_[65997]_ , \new_[65998]_ , \new_[65999]_ ,
    \new_[66002]_ , \new_[66005]_ , \new_[66006]_ , \new_[66009]_ ,
    \new_[66013]_ , \new_[66014]_ , \new_[66015]_ , \new_[66016]_ ,
    \new_[66019]_ , \new_[66022]_ , \new_[66023]_ , \new_[66026]_ ,
    \new_[66030]_ , \new_[66031]_ , \new_[66032]_ , \new_[66033]_ ,
    \new_[66036]_ , \new_[66039]_ , \new_[66040]_ , \new_[66043]_ ,
    \new_[66047]_ , \new_[66048]_ , \new_[66049]_ , \new_[66050]_ ,
    \new_[66053]_ , \new_[66056]_ , \new_[66057]_ , \new_[66060]_ ,
    \new_[66064]_ , \new_[66065]_ , \new_[66066]_ , \new_[66067]_ ,
    \new_[66070]_ , \new_[66073]_ , \new_[66074]_ , \new_[66077]_ ,
    \new_[66081]_ , \new_[66082]_ , \new_[66083]_ , \new_[66084]_ ,
    \new_[66087]_ , \new_[66090]_ , \new_[66091]_ , \new_[66094]_ ,
    \new_[66098]_ , \new_[66099]_ , \new_[66100]_ , \new_[66101]_ ,
    \new_[66104]_ , \new_[66107]_ , \new_[66108]_ , \new_[66111]_ ,
    \new_[66115]_ , \new_[66116]_ , \new_[66117]_ , \new_[66118]_ ,
    \new_[66121]_ , \new_[66124]_ , \new_[66125]_ , \new_[66128]_ ,
    \new_[66132]_ , \new_[66133]_ , \new_[66134]_ , \new_[66135]_ ,
    \new_[66138]_ , \new_[66141]_ , \new_[66142]_ , \new_[66145]_ ,
    \new_[66149]_ , \new_[66150]_ , \new_[66151]_ , \new_[66152]_ ,
    \new_[66155]_ , \new_[66158]_ , \new_[66159]_ , \new_[66162]_ ,
    \new_[66166]_ , \new_[66167]_ , \new_[66168]_ , \new_[66169]_ ,
    \new_[66172]_ , \new_[66175]_ , \new_[66176]_ , \new_[66179]_ ,
    \new_[66183]_ , \new_[66184]_ , \new_[66185]_ , \new_[66186]_ ,
    \new_[66189]_ , \new_[66192]_ , \new_[66193]_ , \new_[66196]_ ,
    \new_[66200]_ , \new_[66201]_ , \new_[66202]_ , \new_[66203]_ ,
    \new_[66206]_ , \new_[66209]_ , \new_[66210]_ , \new_[66213]_ ,
    \new_[66217]_ , \new_[66218]_ , \new_[66219]_ , \new_[66220]_ ,
    \new_[66223]_ , \new_[66226]_ , \new_[66227]_ , \new_[66230]_ ,
    \new_[66234]_ , \new_[66235]_ , \new_[66236]_ , \new_[66237]_ ,
    \new_[66240]_ , \new_[66243]_ , \new_[66244]_ , \new_[66247]_ ,
    \new_[66251]_ , \new_[66252]_ , \new_[66253]_ , \new_[66254]_ ,
    \new_[66257]_ , \new_[66260]_ , \new_[66261]_ , \new_[66264]_ ,
    \new_[66268]_ , \new_[66269]_ , \new_[66270]_ , \new_[66271]_ ,
    \new_[66274]_ , \new_[66277]_ , \new_[66278]_ , \new_[66281]_ ,
    \new_[66285]_ , \new_[66286]_ , \new_[66287]_ , \new_[66288]_ ;
  assign A72 = \new_[7648]_  | \new_[5099]_ ;
  assign \new_[1]_  = \new_[66288]_  & \new_[66271]_ ;
  assign \new_[2]_  = \new_[66254]_  & \new_[66237]_ ;
  assign \new_[3]_  = \new_[66220]_  & \new_[66203]_ ;
  assign \new_[4]_  = \new_[66186]_  & \new_[66169]_ ;
  assign \new_[5]_  = \new_[66152]_  & \new_[66135]_ ;
  assign \new_[6]_  = \new_[66118]_  & \new_[66101]_ ;
  assign \new_[7]_  = \new_[66084]_  & \new_[66067]_ ;
  assign \new_[8]_  = \new_[66050]_  & \new_[66033]_ ;
  assign \new_[9]_  = \new_[66016]_  & \new_[65999]_ ;
  assign \new_[10]_  = \new_[65984]_  & \new_[65967]_ ;
  assign \new_[11]_  = \new_[65952]_  & \new_[65935]_ ;
  assign \new_[12]_  = \new_[65920]_  & \new_[65903]_ ;
  assign \new_[13]_  = \new_[65888]_  & \new_[65871]_ ;
  assign \new_[14]_  = \new_[65856]_  & \new_[65839]_ ;
  assign \new_[15]_  = \new_[65824]_  & \new_[65807]_ ;
  assign \new_[16]_  = \new_[65792]_  & \new_[65775]_ ;
  assign \new_[17]_  = \new_[65760]_  & \new_[65743]_ ;
  assign \new_[18]_  = \new_[65728]_  & \new_[65711]_ ;
  assign \new_[19]_  = \new_[65696]_  & \new_[65679]_ ;
  assign \new_[20]_  = \new_[65664]_  & \new_[65647]_ ;
  assign \new_[21]_  = \new_[65632]_  & \new_[65615]_ ;
  assign \new_[22]_  = \new_[65600]_  & \new_[65583]_ ;
  assign \new_[23]_  = \new_[65568]_  & \new_[65551]_ ;
  assign \new_[24]_  = \new_[65536]_  & \new_[65519]_ ;
  assign \new_[25]_  = \new_[65504]_  & \new_[65487]_ ;
  assign \new_[26]_  = \new_[65472]_  & \new_[65455]_ ;
  assign \new_[27]_  = \new_[65440]_  & \new_[65423]_ ;
  assign \new_[28]_  = \new_[65408]_  & \new_[65391]_ ;
  assign \new_[29]_  = \new_[65376]_  & \new_[65359]_ ;
  assign \new_[30]_  = \new_[65344]_  & \new_[65327]_ ;
  assign \new_[31]_  = \new_[65312]_  & \new_[65295]_ ;
  assign \new_[32]_  = \new_[65280]_  & \new_[65263]_ ;
  assign \new_[33]_  = \new_[65248]_  & \new_[65231]_ ;
  assign \new_[34]_  = \new_[65216]_  & \new_[65199]_ ;
  assign \new_[35]_  = \new_[65184]_  & \new_[65167]_ ;
  assign \new_[36]_  = \new_[65152]_  & \new_[65135]_ ;
  assign \new_[37]_  = \new_[65120]_  & \new_[65103]_ ;
  assign \new_[38]_  = \new_[65088]_  & \new_[65071]_ ;
  assign \new_[39]_  = \new_[65056]_  & \new_[65039]_ ;
  assign \new_[40]_  = \new_[65024]_  & \new_[65007]_ ;
  assign \new_[41]_  = \new_[64992]_  & \new_[64975]_ ;
  assign \new_[42]_  = \new_[64960]_  & \new_[64943]_ ;
  assign \new_[43]_  = \new_[64928]_  & \new_[64911]_ ;
  assign \new_[44]_  = \new_[64896]_  & \new_[64879]_ ;
  assign \new_[45]_  = \new_[64864]_  & \new_[64847]_ ;
  assign \new_[46]_  = \new_[64832]_  & \new_[64815]_ ;
  assign \new_[47]_  = \new_[64800]_  & \new_[64783]_ ;
  assign \new_[48]_  = \new_[64768]_  & \new_[64751]_ ;
  assign \new_[49]_  = \new_[64736]_  & \new_[64719]_ ;
  assign \new_[50]_  = \new_[64704]_  & \new_[64687]_ ;
  assign \new_[51]_  = \new_[64672]_  & \new_[64655]_ ;
  assign \new_[52]_  = \new_[64640]_  & \new_[64623]_ ;
  assign \new_[53]_  = \new_[64608]_  & \new_[64591]_ ;
  assign \new_[54]_  = \new_[64576]_  & \new_[64559]_ ;
  assign \new_[55]_  = \new_[64544]_  & \new_[64527]_ ;
  assign \new_[56]_  = \new_[64512]_  & \new_[64495]_ ;
  assign \new_[57]_  = \new_[64480]_  & \new_[64463]_ ;
  assign \new_[58]_  = \new_[64448]_  & \new_[64431]_ ;
  assign \new_[59]_  = \new_[64416]_  & \new_[64399]_ ;
  assign \new_[60]_  = \new_[64384]_  & \new_[64367]_ ;
  assign \new_[61]_  = \new_[64352]_  & \new_[64335]_ ;
  assign \new_[62]_  = \new_[64320]_  & \new_[64303]_ ;
  assign \new_[63]_  = \new_[64288]_  & \new_[64271]_ ;
  assign \new_[64]_  = \new_[64256]_  & \new_[64239]_ ;
  assign \new_[65]_  = \new_[64224]_  & \new_[64207]_ ;
  assign \new_[66]_  = \new_[64192]_  & \new_[64175]_ ;
  assign \new_[67]_  = \new_[64160]_  & \new_[64143]_ ;
  assign \new_[68]_  = \new_[64128]_  & \new_[64111]_ ;
  assign \new_[69]_  = \new_[64096]_  & \new_[64079]_ ;
  assign \new_[70]_  = \new_[64064]_  & \new_[64047]_ ;
  assign \new_[71]_  = \new_[64032]_  & \new_[64015]_ ;
  assign \new_[72]_  = \new_[64000]_  & \new_[63983]_ ;
  assign \new_[73]_  = \new_[63968]_  & \new_[63953]_ ;
  assign \new_[74]_  = \new_[63938]_  & \new_[63923]_ ;
  assign \new_[75]_  = \new_[63908]_  & \new_[63893]_ ;
  assign \new_[76]_  = \new_[63878]_  & \new_[63863]_ ;
  assign \new_[77]_  = \new_[63848]_  & \new_[63833]_ ;
  assign \new_[78]_  = \new_[63818]_  & \new_[63803]_ ;
  assign \new_[79]_  = \new_[63788]_  & \new_[63773]_ ;
  assign \new_[80]_  = \new_[63758]_  & \new_[63743]_ ;
  assign \new_[81]_  = \new_[63728]_  & \new_[63713]_ ;
  assign \new_[82]_  = \new_[63698]_  & \new_[63683]_ ;
  assign \new_[83]_  = \new_[63668]_  & \new_[63653]_ ;
  assign \new_[84]_  = \new_[63638]_  & \new_[63623]_ ;
  assign \new_[85]_  = \new_[63608]_  & \new_[63593]_ ;
  assign \new_[86]_  = \new_[63578]_  & \new_[63563]_ ;
  assign \new_[87]_  = \new_[63548]_  & \new_[63533]_ ;
  assign \new_[88]_  = \new_[63518]_  & \new_[63503]_ ;
  assign \new_[89]_  = \new_[63488]_  & \new_[63473]_ ;
  assign \new_[90]_  = \new_[63458]_  & \new_[63443]_ ;
  assign \new_[91]_  = \new_[63428]_  & \new_[63413]_ ;
  assign \new_[92]_  = \new_[63398]_  & \new_[63383]_ ;
  assign \new_[93]_  = \new_[63368]_  & \new_[63353]_ ;
  assign \new_[94]_  = \new_[63338]_  & \new_[63323]_ ;
  assign \new_[95]_  = \new_[63308]_  & \new_[63293]_ ;
  assign \new_[96]_  = \new_[63278]_  & \new_[63263]_ ;
  assign \new_[97]_  = \new_[63248]_  & \new_[63233]_ ;
  assign \new_[98]_  = \new_[63218]_  & \new_[63203]_ ;
  assign \new_[99]_  = \new_[63188]_  & \new_[63173]_ ;
  assign \new_[100]_  = \new_[63158]_  & \new_[63143]_ ;
  assign \new_[101]_  = \new_[63128]_  & \new_[63113]_ ;
  assign \new_[102]_  = \new_[63098]_  & \new_[63083]_ ;
  assign \new_[103]_  = \new_[63068]_  & \new_[63053]_ ;
  assign \new_[104]_  = \new_[63038]_  & \new_[63023]_ ;
  assign \new_[105]_  = \new_[63008]_  & \new_[62993]_ ;
  assign \new_[106]_  = \new_[62978]_  & \new_[62963]_ ;
  assign \new_[107]_  = \new_[62948]_  & \new_[62933]_ ;
  assign \new_[108]_  = \new_[62918]_  & \new_[62903]_ ;
  assign \new_[109]_  = \new_[62888]_  & \new_[62873]_ ;
  assign \new_[110]_  = \new_[62858]_  & \new_[62843]_ ;
  assign \new_[111]_  = \new_[62828]_  & \new_[62813]_ ;
  assign \new_[112]_  = \new_[62798]_  & \new_[62783]_ ;
  assign \new_[113]_  = \new_[62768]_  & \new_[62753]_ ;
  assign \new_[114]_  = \new_[62738]_  & \new_[62723]_ ;
  assign \new_[115]_  = \new_[62708]_  & \new_[62693]_ ;
  assign \new_[116]_  = \new_[62678]_  & \new_[62663]_ ;
  assign \new_[117]_  = \new_[62648]_  & \new_[62633]_ ;
  assign \new_[118]_  = \new_[62618]_  & \new_[62603]_ ;
  assign \new_[119]_  = \new_[62588]_  & \new_[62573]_ ;
  assign \new_[120]_  = \new_[62558]_  & \new_[62543]_ ;
  assign \new_[121]_  = \new_[62528]_  & \new_[62513]_ ;
  assign \new_[122]_  = \new_[62498]_  & \new_[62483]_ ;
  assign \new_[123]_  = \new_[62468]_  & \new_[62453]_ ;
  assign \new_[124]_  = \new_[62438]_  & \new_[62423]_ ;
  assign \new_[125]_  = \new_[62408]_  & \new_[62393]_ ;
  assign \new_[126]_  = \new_[62378]_  & \new_[62363]_ ;
  assign \new_[127]_  = \new_[62348]_  & \new_[62333]_ ;
  assign \new_[128]_  = \new_[62318]_  & \new_[62303]_ ;
  assign \new_[129]_  = \new_[62288]_  & \new_[62273]_ ;
  assign \new_[130]_  = \new_[62258]_  & \new_[62243]_ ;
  assign \new_[131]_  = \new_[62228]_  & \new_[62213]_ ;
  assign \new_[132]_  = \new_[62198]_  & \new_[62183]_ ;
  assign \new_[133]_  = \new_[62168]_  & \new_[62153]_ ;
  assign \new_[134]_  = \new_[62138]_  & \new_[62123]_ ;
  assign \new_[135]_  = \new_[62108]_  & \new_[62093]_ ;
  assign \new_[136]_  = \new_[62078]_  & \new_[62063]_ ;
  assign \new_[137]_  = \new_[62048]_  & \new_[62033]_ ;
  assign \new_[138]_  = \new_[62018]_  & \new_[62003]_ ;
  assign \new_[139]_  = \new_[61988]_  & \new_[61973]_ ;
  assign \new_[140]_  = \new_[61958]_  & \new_[61943]_ ;
  assign \new_[141]_  = \new_[61928]_  & \new_[61913]_ ;
  assign \new_[142]_  = \new_[61898]_  & \new_[61883]_ ;
  assign \new_[143]_  = \new_[61868]_  & \new_[61853]_ ;
  assign \new_[144]_  = \new_[61838]_  & \new_[61823]_ ;
  assign \new_[145]_  = \new_[61808]_  & \new_[61793]_ ;
  assign \new_[146]_  = \new_[61778]_  & \new_[61763]_ ;
  assign \new_[147]_  = \new_[61748]_  & \new_[61733]_ ;
  assign \new_[148]_  = \new_[61718]_  & \new_[61703]_ ;
  assign \new_[149]_  = \new_[61688]_  & \new_[61673]_ ;
  assign \new_[150]_  = \new_[61658]_  & \new_[61643]_ ;
  assign \new_[151]_  = \new_[61628]_  & \new_[61613]_ ;
  assign \new_[152]_  = \new_[61598]_  & \new_[61583]_ ;
  assign \new_[153]_  = \new_[61568]_  & \new_[61553]_ ;
  assign \new_[154]_  = \new_[61538]_  & \new_[61523]_ ;
  assign \new_[155]_  = \new_[61508]_  & \new_[61493]_ ;
  assign \new_[156]_  = \new_[61478]_  & \new_[61463]_ ;
  assign \new_[157]_  = \new_[61448]_  & \new_[61433]_ ;
  assign \new_[158]_  = \new_[61418]_  & \new_[61403]_ ;
  assign \new_[159]_  = \new_[61388]_  & \new_[61373]_ ;
  assign \new_[160]_  = \new_[61358]_  & \new_[61343]_ ;
  assign \new_[161]_  = \new_[61328]_  & \new_[61313]_ ;
  assign \new_[162]_  = \new_[61298]_  & \new_[61283]_ ;
  assign \new_[163]_  = \new_[61268]_  & \new_[61253]_ ;
  assign \new_[164]_  = \new_[61238]_  & \new_[61223]_ ;
  assign \new_[165]_  = \new_[61208]_  & \new_[61193]_ ;
  assign \new_[166]_  = \new_[61178]_  & \new_[61163]_ ;
  assign \new_[167]_  = \new_[61148]_  & \new_[61133]_ ;
  assign \new_[168]_  = \new_[61118]_  & \new_[61103]_ ;
  assign \new_[169]_  = \new_[61088]_  & \new_[61073]_ ;
  assign \new_[170]_  = \new_[61058]_  & \new_[61043]_ ;
  assign \new_[171]_  = \new_[61028]_  & \new_[61013]_ ;
  assign \new_[172]_  = \new_[60998]_  & \new_[60983]_ ;
  assign \new_[173]_  = \new_[60968]_  & \new_[60953]_ ;
  assign \new_[174]_  = \new_[60938]_  & \new_[60923]_ ;
  assign \new_[175]_  = \new_[60908]_  & \new_[60893]_ ;
  assign \new_[176]_  = \new_[60878]_  & \new_[60863]_ ;
  assign \new_[177]_  = \new_[60848]_  & \new_[60833]_ ;
  assign \new_[178]_  = \new_[60818]_  & \new_[60803]_ ;
  assign \new_[179]_  = \new_[60788]_  & \new_[60773]_ ;
  assign \new_[180]_  = \new_[60758]_  & \new_[60743]_ ;
  assign \new_[181]_  = \new_[60728]_  & \new_[60713]_ ;
  assign \new_[182]_  = \new_[60698]_  & \new_[60683]_ ;
  assign \new_[183]_  = \new_[60668]_  & \new_[60653]_ ;
  assign \new_[184]_  = \new_[60638]_  & \new_[60623]_ ;
  assign \new_[185]_  = \new_[60608]_  & \new_[60593]_ ;
  assign \new_[186]_  = \new_[60578]_  & \new_[60563]_ ;
  assign \new_[187]_  = \new_[60548]_  & \new_[60533]_ ;
  assign \new_[188]_  = \new_[60518]_  & \new_[60503]_ ;
  assign \new_[189]_  = \new_[60488]_  & \new_[60473]_ ;
  assign \new_[190]_  = \new_[60458]_  & \new_[60443]_ ;
  assign \new_[191]_  = \new_[60428]_  & \new_[60413]_ ;
  assign \new_[192]_  = \new_[60398]_  & \new_[60383]_ ;
  assign \new_[193]_  = \new_[60368]_  & \new_[60353]_ ;
  assign \new_[194]_  = \new_[60338]_  & \new_[60323]_ ;
  assign \new_[195]_  = \new_[60308]_  & \new_[60293]_ ;
  assign \new_[196]_  = \new_[60278]_  & \new_[60263]_ ;
  assign \new_[197]_  = \new_[60248]_  & \new_[60233]_ ;
  assign \new_[198]_  = \new_[60218]_  & \new_[60203]_ ;
  assign \new_[199]_  = \new_[60188]_  & \new_[60173]_ ;
  assign \new_[200]_  = \new_[60158]_  & \new_[60143]_ ;
  assign \new_[201]_  = \new_[60128]_  & \new_[60113]_ ;
  assign \new_[202]_  = \new_[60098]_  & \new_[60083]_ ;
  assign \new_[203]_  = \new_[60068]_  & \new_[60053]_ ;
  assign \new_[204]_  = \new_[60038]_  & \new_[60023]_ ;
  assign \new_[205]_  = \new_[60008]_  & \new_[59993]_ ;
  assign \new_[206]_  = \new_[59978]_  & \new_[59963]_ ;
  assign \new_[207]_  = \new_[59948]_  & \new_[59933]_ ;
  assign \new_[208]_  = \new_[59918]_  & \new_[59903]_ ;
  assign \new_[209]_  = \new_[59888]_  & \new_[59873]_ ;
  assign \new_[210]_  = \new_[59858]_  & \new_[59843]_ ;
  assign \new_[211]_  = \new_[59828]_  & \new_[59813]_ ;
  assign \new_[212]_  = \new_[59798]_  & \new_[59783]_ ;
  assign \new_[213]_  = \new_[59768]_  & \new_[59753]_ ;
  assign \new_[214]_  = \new_[59738]_  & \new_[59723]_ ;
  assign \new_[215]_  = \new_[59708]_  & \new_[59693]_ ;
  assign \new_[216]_  = \new_[59678]_  & \new_[59663]_ ;
  assign \new_[217]_  = \new_[59648]_  & \new_[59633]_ ;
  assign \new_[218]_  = \new_[59618]_  & \new_[59603]_ ;
  assign \new_[219]_  = \new_[59588]_  & \new_[59573]_ ;
  assign \new_[220]_  = \new_[59558]_  & \new_[59543]_ ;
  assign \new_[221]_  = \new_[59528]_  & \new_[59513]_ ;
  assign \new_[222]_  = \new_[59498]_  & \new_[59483]_ ;
  assign \new_[223]_  = \new_[59468]_  & \new_[59453]_ ;
  assign \new_[224]_  = \new_[59438]_  & \new_[59423]_ ;
  assign \new_[225]_  = \new_[59408]_  & \new_[59393]_ ;
  assign \new_[226]_  = \new_[59378]_  & \new_[59363]_ ;
  assign \new_[227]_  = \new_[59348]_  & \new_[59333]_ ;
  assign \new_[228]_  = \new_[59318]_  & \new_[59303]_ ;
  assign \new_[229]_  = \new_[59288]_  & \new_[59273]_ ;
  assign \new_[230]_  = \new_[59258]_  & \new_[59243]_ ;
  assign \new_[231]_  = \new_[59228]_  & \new_[59213]_ ;
  assign \new_[232]_  = \new_[59198]_  & \new_[59183]_ ;
  assign \new_[233]_  = \new_[59168]_  & \new_[59153]_ ;
  assign \new_[234]_  = \new_[59138]_  & \new_[59123]_ ;
  assign \new_[235]_  = \new_[59108]_  & \new_[59093]_ ;
  assign \new_[236]_  = \new_[59078]_  & \new_[59063]_ ;
  assign \new_[237]_  = \new_[59048]_  & \new_[59033]_ ;
  assign \new_[238]_  = \new_[59018]_  & \new_[59003]_ ;
  assign \new_[239]_  = \new_[58988]_  & \new_[58973]_ ;
  assign \new_[240]_  = \new_[58958]_  & \new_[58943]_ ;
  assign \new_[241]_  = \new_[58928]_  & \new_[58913]_ ;
  assign \new_[242]_  = \new_[58898]_  & \new_[58883]_ ;
  assign \new_[243]_  = \new_[58868]_  & \new_[58853]_ ;
  assign \new_[244]_  = \new_[58838]_  & \new_[58823]_ ;
  assign \new_[245]_  = \new_[58808]_  & \new_[58793]_ ;
  assign \new_[246]_  = \new_[58778]_  & \new_[58763]_ ;
  assign \new_[247]_  = \new_[58748]_  & \new_[58733]_ ;
  assign \new_[248]_  = \new_[58718]_  & \new_[58703]_ ;
  assign \new_[249]_  = \new_[58688]_  & \new_[58673]_ ;
  assign \new_[250]_  = \new_[58658]_  & \new_[58643]_ ;
  assign \new_[251]_  = \new_[58628]_  & \new_[58613]_ ;
  assign \new_[252]_  = \new_[58598]_  & \new_[58583]_ ;
  assign \new_[253]_  = \new_[58568]_  & \new_[58553]_ ;
  assign \new_[254]_  = \new_[58538]_  & \new_[58523]_ ;
  assign \new_[255]_  = \new_[58508]_  & \new_[58493]_ ;
  assign \new_[256]_  = \new_[58478]_  & \new_[58463]_ ;
  assign \new_[257]_  = \new_[58448]_  & \new_[58433]_ ;
  assign \new_[258]_  = \new_[58418]_  & \new_[58403]_ ;
  assign \new_[259]_  = \new_[58388]_  & \new_[58373]_ ;
  assign \new_[260]_  = \new_[58358]_  & \new_[58343]_ ;
  assign \new_[261]_  = \new_[58328]_  & \new_[58313]_ ;
  assign \new_[262]_  = \new_[58298]_  & \new_[58283]_ ;
  assign \new_[263]_  = \new_[58268]_  & \new_[58253]_ ;
  assign \new_[264]_  = \new_[58238]_  & \new_[58223]_ ;
  assign \new_[265]_  = \new_[58208]_  & \new_[58193]_ ;
  assign \new_[266]_  = \new_[58178]_  & \new_[58163]_ ;
  assign \new_[267]_  = \new_[58148]_  & \new_[58133]_ ;
  assign \new_[268]_  = \new_[58118]_  & \new_[58103]_ ;
  assign \new_[269]_  = \new_[58088]_  & \new_[58073]_ ;
  assign \new_[270]_  = \new_[58058]_  & \new_[58043]_ ;
  assign \new_[271]_  = \new_[58028]_  & \new_[58013]_ ;
  assign \new_[272]_  = \new_[57998]_  & \new_[57983]_ ;
  assign \new_[273]_  = \new_[57968]_  & \new_[57953]_ ;
  assign \new_[274]_  = \new_[57938]_  & \new_[57923]_ ;
  assign \new_[275]_  = \new_[57908]_  & \new_[57893]_ ;
  assign \new_[276]_  = \new_[57878]_  & \new_[57863]_ ;
  assign \new_[277]_  = \new_[57848]_  & \new_[57833]_ ;
  assign \new_[278]_  = \new_[57818]_  & \new_[57803]_ ;
  assign \new_[279]_  = \new_[57788]_  & \new_[57773]_ ;
  assign \new_[280]_  = \new_[57758]_  & \new_[57743]_ ;
  assign \new_[281]_  = \new_[57728]_  & \new_[57713]_ ;
  assign \new_[282]_  = \new_[57700]_  & \new_[57685]_ ;
  assign \new_[283]_  = \new_[57672]_  & \new_[57657]_ ;
  assign \new_[284]_  = \new_[57644]_  & \new_[57629]_ ;
  assign \new_[285]_  = \new_[57616]_  & \new_[57601]_ ;
  assign \new_[286]_  = \new_[57588]_  & \new_[57573]_ ;
  assign \new_[287]_  = \new_[57560]_  & \new_[57545]_ ;
  assign \new_[288]_  = \new_[57532]_  & \new_[57517]_ ;
  assign \new_[289]_  = \new_[57504]_  & \new_[57489]_ ;
  assign \new_[290]_  = \new_[57476]_  & \new_[57461]_ ;
  assign \new_[291]_  = \new_[57448]_  & \new_[57433]_ ;
  assign \new_[292]_  = \new_[57420]_  & \new_[57405]_ ;
  assign \new_[293]_  = \new_[57392]_  & \new_[57377]_ ;
  assign \new_[294]_  = \new_[57364]_  & \new_[57349]_ ;
  assign \new_[295]_  = \new_[57336]_  & \new_[57321]_ ;
  assign \new_[296]_  = \new_[57308]_  & \new_[57293]_ ;
  assign \new_[297]_  = \new_[57280]_  & \new_[57265]_ ;
  assign \new_[298]_  = \new_[57252]_  & \new_[57237]_ ;
  assign \new_[299]_  = \new_[57224]_  & \new_[57209]_ ;
  assign \new_[300]_  = \new_[57196]_  & \new_[57181]_ ;
  assign \new_[301]_  = \new_[57168]_  & \new_[57153]_ ;
  assign \new_[302]_  = \new_[57140]_  & \new_[57125]_ ;
  assign \new_[303]_  = \new_[57112]_  & \new_[57097]_ ;
  assign \new_[304]_  = \new_[57084]_  & \new_[57069]_ ;
  assign \new_[305]_  = \new_[57056]_  & \new_[57041]_ ;
  assign \new_[306]_  = \new_[57028]_  & \new_[57013]_ ;
  assign \new_[307]_  = \new_[57000]_  & \new_[56985]_ ;
  assign \new_[308]_  = \new_[56972]_  & \new_[56957]_ ;
  assign \new_[309]_  = \new_[56944]_  & \new_[56929]_ ;
  assign \new_[310]_  = \new_[56916]_  & \new_[56901]_ ;
  assign \new_[311]_  = \new_[56888]_  & \new_[56873]_ ;
  assign \new_[312]_  = \new_[56860]_  & \new_[56845]_ ;
  assign \new_[313]_  = \new_[56832]_  & \new_[56817]_ ;
  assign \new_[314]_  = \new_[56804]_  & \new_[56789]_ ;
  assign \new_[315]_  = \new_[56776]_  & \new_[56761]_ ;
  assign \new_[316]_  = \new_[56748]_  & \new_[56733]_ ;
  assign \new_[317]_  = \new_[56720]_  & \new_[56705]_ ;
  assign \new_[318]_  = \new_[56692]_  & \new_[56677]_ ;
  assign \new_[319]_  = \new_[56664]_  & \new_[56649]_ ;
  assign \new_[320]_  = \new_[56636]_  & \new_[56621]_ ;
  assign \new_[321]_  = \new_[56608]_  & \new_[56593]_ ;
  assign \new_[322]_  = \new_[56580]_  & \new_[56565]_ ;
  assign \new_[323]_  = \new_[56552]_  & \new_[56537]_ ;
  assign \new_[324]_  = \new_[56524]_  & \new_[56509]_ ;
  assign \new_[325]_  = \new_[56496]_  & \new_[56481]_ ;
  assign \new_[326]_  = \new_[56468]_  & \new_[56453]_ ;
  assign \new_[327]_  = \new_[56440]_  & \new_[56425]_ ;
  assign \new_[328]_  = \new_[56412]_  & \new_[56397]_ ;
  assign \new_[329]_  = \new_[56384]_  & \new_[56369]_ ;
  assign \new_[330]_  = \new_[56356]_  & \new_[56341]_ ;
  assign \new_[331]_  = \new_[56328]_  & \new_[56313]_ ;
  assign \new_[332]_  = \new_[56300]_  & \new_[56285]_ ;
  assign \new_[333]_  = \new_[56272]_  & \new_[56257]_ ;
  assign \new_[334]_  = \new_[56244]_  & \new_[56229]_ ;
  assign \new_[335]_  = \new_[56216]_  & \new_[56201]_ ;
  assign \new_[336]_  = \new_[56188]_  & \new_[56173]_ ;
  assign \new_[337]_  = \new_[56160]_  & \new_[56145]_ ;
  assign \new_[338]_  = \new_[56132]_  & \new_[56117]_ ;
  assign \new_[339]_  = \new_[56104]_  & \new_[56089]_ ;
  assign \new_[340]_  = \new_[56076]_  & \new_[56061]_ ;
  assign \new_[341]_  = \new_[56048]_  & \new_[56033]_ ;
  assign \new_[342]_  = \new_[56020]_  & \new_[56005]_ ;
  assign \new_[343]_  = \new_[55992]_  & \new_[55977]_ ;
  assign \new_[344]_  = \new_[55964]_  & \new_[55949]_ ;
  assign \new_[345]_  = \new_[55936]_  & \new_[55921]_ ;
  assign \new_[346]_  = \new_[55908]_  & \new_[55893]_ ;
  assign \new_[347]_  = \new_[55880]_  & \new_[55865]_ ;
  assign \new_[348]_  = \new_[55852]_  & \new_[55837]_ ;
  assign \new_[349]_  = \new_[55824]_  & \new_[55809]_ ;
  assign \new_[350]_  = \new_[55796]_  & \new_[55781]_ ;
  assign \new_[351]_  = \new_[55768]_  & \new_[55753]_ ;
  assign \new_[352]_  = \new_[55740]_  & \new_[55725]_ ;
  assign \new_[353]_  = \new_[55712]_  & \new_[55697]_ ;
  assign \new_[354]_  = \new_[55684]_  & \new_[55669]_ ;
  assign \new_[355]_  = \new_[55656]_  & \new_[55641]_ ;
  assign \new_[356]_  = \new_[55628]_  & \new_[55613]_ ;
  assign \new_[357]_  = \new_[55600]_  & \new_[55585]_ ;
  assign \new_[358]_  = \new_[55572]_  & \new_[55557]_ ;
  assign \new_[359]_  = \new_[55544]_  & \new_[55529]_ ;
  assign \new_[360]_  = \new_[55516]_  & \new_[55501]_ ;
  assign \new_[361]_  = \new_[55488]_  & \new_[55473]_ ;
  assign \new_[362]_  = \new_[55460]_  & \new_[55445]_ ;
  assign \new_[363]_  = \new_[55432]_  & \new_[55417]_ ;
  assign \new_[364]_  = \new_[55404]_  & \new_[55389]_ ;
  assign \new_[365]_  = \new_[55376]_  & \new_[55361]_ ;
  assign \new_[366]_  = \new_[55348]_  & \new_[55333]_ ;
  assign \new_[367]_  = \new_[55320]_  & \new_[55305]_ ;
  assign \new_[368]_  = \new_[55292]_  & \new_[55277]_ ;
  assign \new_[369]_  = \new_[55264]_  & \new_[55249]_ ;
  assign \new_[370]_  = \new_[55236]_  & \new_[55221]_ ;
  assign \new_[371]_  = \new_[55208]_  & \new_[55193]_ ;
  assign \new_[372]_  = \new_[55180]_  & \new_[55165]_ ;
  assign \new_[373]_  = \new_[55152]_  & \new_[55137]_ ;
  assign \new_[374]_  = \new_[55124]_  & \new_[55109]_ ;
  assign \new_[375]_  = \new_[55096]_  & \new_[55081]_ ;
  assign \new_[376]_  = \new_[55068]_  & \new_[55053]_ ;
  assign \new_[377]_  = \new_[55040]_  & \new_[55025]_ ;
  assign \new_[378]_  = \new_[55012]_  & \new_[54997]_ ;
  assign \new_[379]_  = \new_[54984]_  & \new_[54969]_ ;
  assign \new_[380]_  = \new_[54956]_  & \new_[54941]_ ;
  assign \new_[381]_  = \new_[54928]_  & \new_[54913]_ ;
  assign \new_[382]_  = \new_[54900]_  & \new_[54885]_ ;
  assign \new_[383]_  = \new_[54872]_  & \new_[54857]_ ;
  assign \new_[384]_  = \new_[54844]_  & \new_[54829]_ ;
  assign \new_[385]_  = \new_[54816]_  & \new_[54801]_ ;
  assign \new_[386]_  = \new_[54788]_  & \new_[54773]_ ;
  assign \new_[387]_  = \new_[54760]_  & \new_[54745]_ ;
  assign \new_[388]_  = \new_[54732]_  & \new_[54717]_ ;
  assign \new_[389]_  = \new_[54704]_  & \new_[54689]_ ;
  assign \new_[390]_  = \new_[54676]_  & \new_[54661]_ ;
  assign \new_[391]_  = \new_[54648]_  & \new_[54633]_ ;
  assign \new_[392]_  = \new_[54620]_  & \new_[54605]_ ;
  assign \new_[393]_  = \new_[54592]_  & \new_[54577]_ ;
  assign \new_[394]_  = \new_[54564]_  & \new_[54549]_ ;
  assign \new_[395]_  = \new_[54536]_  & \new_[54521]_ ;
  assign \new_[396]_  = \new_[54508]_  & \new_[54493]_ ;
  assign \new_[397]_  = \new_[54480]_  & \new_[54465]_ ;
  assign \new_[398]_  = \new_[54452]_  & \new_[54437]_ ;
  assign \new_[399]_  = \new_[54424]_  & \new_[54409]_ ;
  assign \new_[400]_  = \new_[54396]_  & \new_[54381]_ ;
  assign \new_[401]_  = \new_[54368]_  & \new_[54353]_ ;
  assign \new_[402]_  = \new_[54340]_  & \new_[54325]_ ;
  assign \new_[403]_  = \new_[54312]_  & \new_[54297]_ ;
  assign \new_[404]_  = \new_[54284]_  & \new_[54269]_ ;
  assign \new_[405]_  = \new_[54256]_  & \new_[54241]_ ;
  assign \new_[406]_  = \new_[54228]_  & \new_[54213]_ ;
  assign \new_[407]_  = \new_[54200]_  & \new_[54185]_ ;
  assign \new_[408]_  = \new_[54172]_  & \new_[54157]_ ;
  assign \new_[409]_  = \new_[54144]_  & \new_[54129]_ ;
  assign \new_[410]_  = \new_[54116]_  & \new_[54101]_ ;
  assign \new_[411]_  = \new_[54088]_  & \new_[54073]_ ;
  assign \new_[412]_  = \new_[54060]_  & \new_[54045]_ ;
  assign \new_[413]_  = \new_[54032]_  & \new_[54017]_ ;
  assign \new_[414]_  = \new_[54004]_  & \new_[53989]_ ;
  assign \new_[415]_  = \new_[53976]_  & \new_[53961]_ ;
  assign \new_[416]_  = \new_[53948]_  & \new_[53933]_ ;
  assign \new_[417]_  = \new_[53920]_  & \new_[53905]_ ;
  assign \new_[418]_  = \new_[53892]_  & \new_[53877]_ ;
  assign \new_[419]_  = \new_[53864]_  & \new_[53849]_ ;
  assign \new_[420]_  = \new_[53836]_  & \new_[53821]_ ;
  assign \new_[421]_  = \new_[53808]_  & \new_[53793]_ ;
  assign \new_[422]_  = \new_[53780]_  & \new_[53765]_ ;
  assign \new_[423]_  = \new_[53752]_  & \new_[53737]_ ;
  assign \new_[424]_  = \new_[53724]_  & \new_[53709]_ ;
  assign \new_[425]_  = \new_[53696]_  & \new_[53681]_ ;
  assign \new_[426]_  = \new_[53668]_  & \new_[53653]_ ;
  assign \new_[427]_  = \new_[53640]_  & \new_[53625]_ ;
  assign \new_[428]_  = \new_[53612]_  & \new_[53597]_ ;
  assign \new_[429]_  = \new_[53584]_  & \new_[53569]_ ;
  assign \new_[430]_  = \new_[53556]_  & \new_[53541]_ ;
  assign \new_[431]_  = \new_[53528]_  & \new_[53513]_ ;
  assign \new_[432]_  = \new_[53500]_  & \new_[53485]_ ;
  assign \new_[433]_  = \new_[53472]_  & \new_[53457]_ ;
  assign \new_[434]_  = \new_[53444]_  & \new_[53429]_ ;
  assign \new_[435]_  = \new_[53416]_  & \new_[53401]_ ;
  assign \new_[436]_  = \new_[53388]_  & \new_[53373]_ ;
  assign \new_[437]_  = \new_[53360]_  & \new_[53345]_ ;
  assign \new_[438]_  = \new_[53332]_  & \new_[53317]_ ;
  assign \new_[439]_  = \new_[53304]_  & \new_[53289]_ ;
  assign \new_[440]_  = \new_[53276]_  & \new_[53261]_ ;
  assign \new_[441]_  = \new_[53248]_  & \new_[53233]_ ;
  assign \new_[442]_  = \new_[53220]_  & \new_[53205]_ ;
  assign \new_[443]_  = \new_[53192]_  & \new_[53177]_ ;
  assign \new_[444]_  = \new_[53164]_  & \new_[53149]_ ;
  assign \new_[445]_  = \new_[53136]_  & \new_[53121]_ ;
  assign \new_[446]_  = \new_[53108]_  & \new_[53093]_ ;
  assign \new_[447]_  = \new_[53080]_  & \new_[53065]_ ;
  assign \new_[448]_  = \new_[53052]_  & \new_[53037]_ ;
  assign \new_[449]_  = \new_[53024]_  & \new_[53009]_ ;
  assign \new_[450]_  = \new_[52996]_  & \new_[52981]_ ;
  assign \new_[451]_  = \new_[52968]_  & \new_[52953]_ ;
  assign \new_[452]_  = \new_[52940]_  & \new_[52925]_ ;
  assign \new_[453]_  = \new_[52912]_  & \new_[52897]_ ;
  assign \new_[454]_  = \new_[52884]_  & \new_[52869]_ ;
  assign \new_[455]_  = \new_[52856]_  & \new_[52841]_ ;
  assign \new_[456]_  = \new_[52828]_  & \new_[52813]_ ;
  assign \new_[457]_  = \new_[52800]_  & \new_[52785]_ ;
  assign \new_[458]_  = \new_[52772]_  & \new_[52757]_ ;
  assign \new_[459]_  = \new_[52744]_  & \new_[52729]_ ;
  assign \new_[460]_  = \new_[52716]_  & \new_[52701]_ ;
  assign \new_[461]_  = \new_[52688]_  & \new_[52673]_ ;
  assign \new_[462]_  = \new_[52660]_  & \new_[52645]_ ;
  assign \new_[463]_  = \new_[52632]_  & \new_[52617]_ ;
  assign \new_[464]_  = \new_[52604]_  & \new_[52589]_ ;
  assign \new_[465]_  = \new_[52576]_  & \new_[52561]_ ;
  assign \new_[466]_  = \new_[52548]_  & \new_[52533]_ ;
  assign \new_[467]_  = \new_[52520]_  & \new_[52505]_ ;
  assign \new_[468]_  = \new_[52492]_  & \new_[52477]_ ;
  assign \new_[469]_  = \new_[52464]_  & \new_[52449]_ ;
  assign \new_[470]_  = \new_[52436]_  & \new_[52421]_ ;
  assign \new_[471]_  = \new_[52408]_  & \new_[52393]_ ;
  assign \new_[472]_  = \new_[52380]_  & \new_[52365]_ ;
  assign \new_[473]_  = \new_[52352]_  & \new_[52337]_ ;
  assign \new_[474]_  = \new_[52324]_  & \new_[52309]_ ;
  assign \new_[475]_  = \new_[52296]_  & \new_[52281]_ ;
  assign \new_[476]_  = \new_[52268]_  & \new_[52253]_ ;
  assign \new_[477]_  = \new_[52240]_  & \new_[52225]_ ;
  assign \new_[478]_  = \new_[52212]_  & \new_[52197]_ ;
  assign \new_[479]_  = \new_[52184]_  & \new_[52169]_ ;
  assign \new_[480]_  = \new_[52156]_  & \new_[52141]_ ;
  assign \new_[481]_  = \new_[52128]_  & \new_[52113]_ ;
  assign \new_[482]_  = \new_[52100]_  & \new_[52085]_ ;
  assign \new_[483]_  = \new_[52072]_  & \new_[52057]_ ;
  assign \new_[484]_  = \new_[52044]_  & \new_[52029]_ ;
  assign \new_[485]_  = \new_[52016]_  & \new_[52001]_ ;
  assign \new_[486]_  = \new_[51988]_  & \new_[51973]_ ;
  assign \new_[487]_  = \new_[51960]_  & \new_[51945]_ ;
  assign \new_[488]_  = \new_[51932]_  & \new_[51917]_ ;
  assign \new_[489]_  = \new_[51904]_  & \new_[51889]_ ;
  assign \new_[490]_  = \new_[51876]_  & \new_[51861]_ ;
  assign \new_[491]_  = \new_[51848]_  & \new_[51833]_ ;
  assign \new_[492]_  = \new_[51820]_  & \new_[51805]_ ;
  assign \new_[493]_  = \new_[51792]_  & \new_[51777]_ ;
  assign \new_[494]_  = \new_[51764]_  & \new_[51749]_ ;
  assign \new_[495]_  = \new_[51736]_  & \new_[51721]_ ;
  assign \new_[496]_  = \new_[51708]_  & \new_[51693]_ ;
  assign \new_[497]_  = \new_[51680]_  & \new_[51665]_ ;
  assign \new_[498]_  = \new_[51652]_  & \new_[51637]_ ;
  assign \new_[499]_  = \new_[51624]_  & \new_[51609]_ ;
  assign \new_[500]_  = \new_[51596]_  & \new_[51581]_ ;
  assign \new_[501]_  = \new_[51568]_  & \new_[51553]_ ;
  assign \new_[502]_  = \new_[51540]_  & \new_[51525]_ ;
  assign \new_[503]_  = \new_[51512]_  & \new_[51497]_ ;
  assign \new_[504]_  = \new_[51484]_  & \new_[51469]_ ;
  assign \new_[505]_  = \new_[51456]_  & \new_[51441]_ ;
  assign \new_[506]_  = \new_[51428]_  & \new_[51413]_ ;
  assign \new_[507]_  = \new_[51400]_  & \new_[51385]_ ;
  assign \new_[508]_  = \new_[51372]_  & \new_[51357]_ ;
  assign \new_[509]_  = \new_[51344]_  & \new_[51329]_ ;
  assign \new_[510]_  = \new_[51316]_  & \new_[51301]_ ;
  assign \new_[511]_  = \new_[51288]_  & \new_[51273]_ ;
  assign \new_[512]_  = \new_[51260]_  & \new_[51245]_ ;
  assign \new_[513]_  = \new_[51232]_  & \new_[51217]_ ;
  assign \new_[514]_  = \new_[51204]_  & \new_[51189]_ ;
  assign \new_[515]_  = \new_[51176]_  & \new_[51161]_ ;
  assign \new_[516]_  = \new_[51148]_  & \new_[51133]_ ;
  assign \new_[517]_  = \new_[51120]_  & \new_[51105]_ ;
  assign \new_[518]_  = \new_[51092]_  & \new_[51077]_ ;
  assign \new_[519]_  = \new_[51064]_  & \new_[51049]_ ;
  assign \new_[520]_  = \new_[51036]_  & \new_[51021]_ ;
  assign \new_[521]_  = \new_[51008]_  & \new_[50993]_ ;
  assign \new_[522]_  = \new_[50980]_  & \new_[50965]_ ;
  assign \new_[523]_  = \new_[50952]_  & \new_[50937]_ ;
  assign \new_[524]_  = \new_[50924]_  & \new_[50909]_ ;
  assign \new_[525]_  = \new_[50896]_  & \new_[50881]_ ;
  assign \new_[526]_  = \new_[50868]_  & \new_[50853]_ ;
  assign \new_[527]_  = \new_[50840]_  & \new_[50825]_ ;
  assign \new_[528]_  = \new_[50812]_  & \new_[50797]_ ;
  assign \new_[529]_  = \new_[50784]_  & \new_[50769]_ ;
  assign \new_[530]_  = \new_[50756]_  & \new_[50741]_ ;
  assign \new_[531]_  = \new_[50728]_  & \new_[50713]_ ;
  assign \new_[532]_  = \new_[50700]_  & \new_[50685]_ ;
  assign \new_[533]_  = \new_[50672]_  & \new_[50657]_ ;
  assign \new_[534]_  = \new_[50644]_  & \new_[50629]_ ;
  assign \new_[535]_  = \new_[50616]_  & \new_[50601]_ ;
  assign \new_[536]_  = \new_[50588]_  & \new_[50573]_ ;
  assign \new_[537]_  = \new_[50560]_  & \new_[50545]_ ;
  assign \new_[538]_  = \new_[50532]_  & \new_[50517]_ ;
  assign \new_[539]_  = \new_[50504]_  & \new_[50489]_ ;
  assign \new_[540]_  = \new_[50476]_  & \new_[50461]_ ;
  assign \new_[541]_  = \new_[50448]_  & \new_[50433]_ ;
  assign \new_[542]_  = \new_[50420]_  & \new_[50405]_ ;
  assign \new_[543]_  = \new_[50392]_  & \new_[50377]_ ;
  assign \new_[544]_  = \new_[50364]_  & \new_[50349]_ ;
  assign \new_[545]_  = \new_[50336]_  & \new_[50321]_ ;
  assign \new_[546]_  = \new_[50308]_  & \new_[50293]_ ;
  assign \new_[547]_  = \new_[50280]_  & \new_[50265]_ ;
  assign \new_[548]_  = \new_[50252]_  & \new_[50237]_ ;
  assign \new_[549]_  = \new_[50224]_  & \new_[50209]_ ;
  assign \new_[550]_  = \new_[50196]_  & \new_[50181]_ ;
  assign \new_[551]_  = \new_[50168]_  & \new_[50153]_ ;
  assign \new_[552]_  = \new_[50140]_  & \new_[50125]_ ;
  assign \new_[553]_  = \new_[50112]_  & \new_[50097]_ ;
  assign \new_[554]_  = \new_[50084]_  & \new_[50069]_ ;
  assign \new_[555]_  = \new_[50056]_  & \new_[50041]_ ;
  assign \new_[556]_  = \new_[50028]_  & \new_[50013]_ ;
  assign \new_[557]_  = \new_[50000]_  & \new_[49985]_ ;
  assign \new_[558]_  = \new_[49972]_  & \new_[49957]_ ;
  assign \new_[559]_  = \new_[49944]_  & \new_[49929]_ ;
  assign \new_[560]_  = \new_[49916]_  & \new_[49901]_ ;
  assign \new_[561]_  = \new_[49888]_  & \new_[49873]_ ;
  assign \new_[562]_  = \new_[49860]_  & \new_[49845]_ ;
  assign \new_[563]_  = \new_[49832]_  & \new_[49817]_ ;
  assign \new_[564]_  = \new_[49804]_  & \new_[49789]_ ;
  assign \new_[565]_  = \new_[49776]_  & \new_[49761]_ ;
  assign \new_[566]_  = \new_[49748]_  & \new_[49733]_ ;
  assign \new_[567]_  = \new_[49720]_  & \new_[49705]_ ;
  assign \new_[568]_  = \new_[49692]_  & \new_[49677]_ ;
  assign \new_[569]_  = \new_[49664]_  & \new_[49649]_ ;
  assign \new_[570]_  = \new_[49636]_  & \new_[49621]_ ;
  assign \new_[571]_  = \new_[49608]_  & \new_[49593]_ ;
  assign \new_[572]_  = \new_[49580]_  & \new_[49565]_ ;
  assign \new_[573]_  = \new_[49552]_  & \new_[49537]_ ;
  assign \new_[574]_  = \new_[49524]_  & \new_[49509]_ ;
  assign \new_[575]_  = \new_[49496]_  & \new_[49481]_ ;
  assign \new_[576]_  = \new_[49468]_  & \new_[49453]_ ;
  assign \new_[577]_  = \new_[49440]_  & \new_[49425]_ ;
  assign \new_[578]_  = \new_[49412]_  & \new_[49397]_ ;
  assign \new_[579]_  = \new_[49384]_  & \new_[49369]_ ;
  assign \new_[580]_  = \new_[49356]_  & \new_[49341]_ ;
  assign \new_[581]_  = \new_[49328]_  & \new_[49313]_ ;
  assign \new_[582]_  = \new_[49300]_  & \new_[49285]_ ;
  assign \new_[583]_  = \new_[49272]_  & \new_[49257]_ ;
  assign \new_[584]_  = \new_[49244]_  & \new_[49229]_ ;
  assign \new_[585]_  = \new_[49216]_  & \new_[49201]_ ;
  assign \new_[586]_  = \new_[49188]_  & \new_[49173]_ ;
  assign \new_[587]_  = \new_[49160]_  & \new_[49145]_ ;
  assign \new_[588]_  = \new_[49132]_  & \new_[49117]_ ;
  assign \new_[589]_  = \new_[49104]_  & \new_[49089]_ ;
  assign \new_[590]_  = \new_[49076]_  & \new_[49061]_ ;
  assign \new_[591]_  = \new_[49048]_  & \new_[49033]_ ;
  assign \new_[592]_  = \new_[49020]_  & \new_[49005]_ ;
  assign \new_[593]_  = \new_[48992]_  & \new_[48977]_ ;
  assign \new_[594]_  = \new_[48964]_  & \new_[48949]_ ;
  assign \new_[595]_  = \new_[48936]_  & \new_[48921]_ ;
  assign \new_[596]_  = \new_[48908]_  & \new_[48893]_ ;
  assign \new_[597]_  = \new_[48880]_  & \new_[48865]_ ;
  assign \new_[598]_  = \new_[48852]_  & \new_[48837]_ ;
  assign \new_[599]_  = \new_[48824]_  & \new_[48809]_ ;
  assign \new_[600]_  = \new_[48796]_  & \new_[48781]_ ;
  assign \new_[601]_  = \new_[48768]_  & \new_[48753]_ ;
  assign \new_[602]_  = \new_[48740]_  & \new_[48725]_ ;
  assign \new_[603]_  = \new_[48712]_  & \new_[48697]_ ;
  assign \new_[604]_  = \new_[48684]_  & \new_[48669]_ ;
  assign \new_[605]_  = \new_[48656]_  & \new_[48641]_ ;
  assign \new_[606]_  = \new_[48628]_  & \new_[48613]_ ;
  assign \new_[607]_  = \new_[48600]_  & \new_[48585]_ ;
  assign \new_[608]_  = \new_[48572]_  & \new_[48557]_ ;
  assign \new_[609]_  = \new_[48544]_  & \new_[48529]_ ;
  assign \new_[610]_  = \new_[48516]_  & \new_[48501]_ ;
  assign \new_[611]_  = \new_[48488]_  & \new_[48473]_ ;
  assign \new_[612]_  = \new_[48460]_  & \new_[48445]_ ;
  assign \new_[613]_  = \new_[48432]_  & \new_[48417]_ ;
  assign \new_[614]_  = \new_[48404]_  & \new_[48389]_ ;
  assign \new_[615]_  = \new_[48376]_  & \new_[48361]_ ;
  assign \new_[616]_  = \new_[48348]_  & \new_[48333]_ ;
  assign \new_[617]_  = \new_[48320]_  & \new_[48305]_ ;
  assign \new_[618]_  = \new_[48292]_  & \new_[48277]_ ;
  assign \new_[619]_  = \new_[48264]_  & \new_[48249]_ ;
  assign \new_[620]_  = \new_[48236]_  & \new_[48221]_ ;
  assign \new_[621]_  = \new_[48208]_  & \new_[48193]_ ;
  assign \new_[622]_  = \new_[48180]_  & \new_[48165]_ ;
  assign \new_[623]_  = \new_[48152]_  & \new_[48137]_ ;
  assign \new_[624]_  = \new_[48124]_  & \new_[48109]_ ;
  assign \new_[625]_  = \new_[48096]_  & \new_[48081]_ ;
  assign \new_[626]_  = \new_[48068]_  & \new_[48053]_ ;
  assign \new_[627]_  = \new_[48040]_  & \new_[48025]_ ;
  assign \new_[628]_  = \new_[48012]_  & \new_[47997]_ ;
  assign \new_[629]_  = \new_[47984]_  & \new_[47969]_ ;
  assign \new_[630]_  = \new_[47956]_  & \new_[47941]_ ;
  assign \new_[631]_  = \new_[47928]_  & \new_[47913]_ ;
  assign \new_[632]_  = \new_[47900]_  & \new_[47885]_ ;
  assign \new_[633]_  = \new_[47872]_  & \new_[47857]_ ;
  assign \new_[634]_  = \new_[47844]_  & \new_[47829]_ ;
  assign \new_[635]_  = \new_[47816]_  & \new_[47801]_ ;
  assign \new_[636]_  = \new_[47788]_  & \new_[47773]_ ;
  assign \new_[637]_  = \new_[47760]_  & \new_[47745]_ ;
  assign \new_[638]_  = \new_[47732]_  & \new_[47717]_ ;
  assign \new_[639]_  = \new_[47704]_  & \new_[47689]_ ;
  assign \new_[640]_  = \new_[47676]_  & \new_[47661]_ ;
  assign \new_[641]_  = \new_[47648]_  & \new_[47635]_ ;
  assign \new_[642]_  = \new_[47622]_  & \new_[47609]_ ;
  assign \new_[643]_  = \new_[47596]_  & \new_[47583]_ ;
  assign \new_[644]_  = \new_[47570]_  & \new_[47557]_ ;
  assign \new_[645]_  = \new_[47544]_  & \new_[47531]_ ;
  assign \new_[646]_  = \new_[47518]_  & \new_[47505]_ ;
  assign \new_[647]_  = \new_[47492]_  & \new_[47479]_ ;
  assign \new_[648]_  = \new_[47466]_  & \new_[47453]_ ;
  assign \new_[649]_  = \new_[47440]_  & \new_[47427]_ ;
  assign \new_[650]_  = \new_[47414]_  & \new_[47401]_ ;
  assign \new_[651]_  = \new_[47388]_  & \new_[47375]_ ;
  assign \new_[652]_  = \new_[47362]_  & \new_[47349]_ ;
  assign \new_[653]_  = \new_[47336]_  & \new_[47323]_ ;
  assign \new_[654]_  = \new_[47310]_  & \new_[47297]_ ;
  assign \new_[655]_  = \new_[47284]_  & \new_[47271]_ ;
  assign \new_[656]_  = \new_[47258]_  & \new_[47245]_ ;
  assign \new_[657]_  = \new_[47232]_  & \new_[47219]_ ;
  assign \new_[658]_  = \new_[47206]_  & \new_[47193]_ ;
  assign \new_[659]_  = \new_[47180]_  & \new_[47167]_ ;
  assign \new_[660]_  = \new_[47154]_  & \new_[47141]_ ;
  assign \new_[661]_  = \new_[47128]_  & \new_[47115]_ ;
  assign \new_[662]_  = \new_[47102]_  & \new_[47089]_ ;
  assign \new_[663]_  = \new_[47076]_  & \new_[47063]_ ;
  assign \new_[664]_  = \new_[47050]_  & \new_[47037]_ ;
  assign \new_[665]_  = \new_[47024]_  & \new_[47011]_ ;
  assign \new_[666]_  = \new_[46998]_  & \new_[46985]_ ;
  assign \new_[667]_  = \new_[46972]_  & \new_[46959]_ ;
  assign \new_[668]_  = \new_[46946]_  & \new_[46933]_ ;
  assign \new_[669]_  = \new_[46920]_  & \new_[46907]_ ;
  assign \new_[670]_  = \new_[46894]_  & \new_[46881]_ ;
  assign \new_[671]_  = \new_[46868]_  & \new_[46855]_ ;
  assign \new_[672]_  = \new_[46842]_  & \new_[46829]_ ;
  assign \new_[673]_  = \new_[46816]_  & \new_[46803]_ ;
  assign \new_[674]_  = \new_[46790]_  & \new_[46777]_ ;
  assign \new_[675]_  = \new_[46764]_  & \new_[46751]_ ;
  assign \new_[676]_  = \new_[46738]_  & \new_[46725]_ ;
  assign \new_[677]_  = \new_[46712]_  & \new_[46699]_ ;
  assign \new_[678]_  = \new_[46686]_  & \new_[46673]_ ;
  assign \new_[679]_  = \new_[46660]_  & \new_[46647]_ ;
  assign \new_[680]_  = \new_[46634]_  & \new_[46621]_ ;
  assign \new_[681]_  = \new_[46608]_  & \new_[46595]_ ;
  assign \new_[682]_  = \new_[46582]_  & \new_[46569]_ ;
  assign \new_[683]_  = \new_[46556]_  & \new_[46543]_ ;
  assign \new_[684]_  = \new_[46530]_  & \new_[46517]_ ;
  assign \new_[685]_  = \new_[46504]_  & \new_[46491]_ ;
  assign \new_[686]_  = \new_[46478]_  & \new_[46465]_ ;
  assign \new_[687]_  = \new_[46452]_  & \new_[46439]_ ;
  assign \new_[688]_  = \new_[46426]_  & \new_[46413]_ ;
  assign \new_[689]_  = \new_[46400]_  & \new_[46387]_ ;
  assign \new_[690]_  = \new_[46374]_  & \new_[46361]_ ;
  assign \new_[691]_  = \new_[46348]_  & \new_[46335]_ ;
  assign \new_[692]_  = \new_[46322]_  & \new_[46309]_ ;
  assign \new_[693]_  = \new_[46296]_  & \new_[46283]_ ;
  assign \new_[694]_  = \new_[46270]_  & \new_[46257]_ ;
  assign \new_[695]_  = \new_[46244]_  & \new_[46231]_ ;
  assign \new_[696]_  = \new_[46218]_  & \new_[46205]_ ;
  assign \new_[697]_  = \new_[46192]_  & \new_[46179]_ ;
  assign \new_[698]_  = \new_[46166]_  & \new_[46153]_ ;
  assign \new_[699]_  = \new_[46140]_  & \new_[46127]_ ;
  assign \new_[700]_  = \new_[46114]_  & \new_[46101]_ ;
  assign \new_[701]_  = \new_[46088]_  & \new_[46075]_ ;
  assign \new_[702]_  = \new_[46062]_  & \new_[46049]_ ;
  assign \new_[703]_  = \new_[46036]_  & \new_[46023]_ ;
  assign \new_[704]_  = \new_[46010]_  & \new_[45997]_ ;
  assign \new_[705]_  = \new_[45984]_  & \new_[45971]_ ;
  assign \new_[706]_  = \new_[45958]_  & \new_[45945]_ ;
  assign \new_[707]_  = \new_[45932]_  & \new_[45919]_ ;
  assign \new_[708]_  = \new_[45906]_  & \new_[45893]_ ;
  assign \new_[709]_  = \new_[45880]_  & \new_[45867]_ ;
  assign \new_[710]_  = \new_[45854]_  & \new_[45841]_ ;
  assign \new_[711]_  = \new_[45828]_  & \new_[45815]_ ;
  assign \new_[712]_  = \new_[45802]_  & \new_[45789]_ ;
  assign \new_[713]_  = \new_[45776]_  & \new_[45763]_ ;
  assign \new_[714]_  = \new_[45750]_  & \new_[45737]_ ;
  assign \new_[715]_  = \new_[45724]_  & \new_[45711]_ ;
  assign \new_[716]_  = \new_[45698]_  & \new_[45685]_ ;
  assign \new_[717]_  = \new_[45672]_  & \new_[45659]_ ;
  assign \new_[718]_  = \new_[45646]_  & \new_[45633]_ ;
  assign \new_[719]_  = \new_[45620]_  & \new_[45607]_ ;
  assign \new_[720]_  = \new_[45594]_  & \new_[45581]_ ;
  assign \new_[721]_  = \new_[45568]_  & \new_[45555]_ ;
  assign \new_[722]_  = \new_[45542]_  & \new_[45529]_ ;
  assign \new_[723]_  = \new_[45516]_  & \new_[45503]_ ;
  assign \new_[724]_  = \new_[45490]_  & \new_[45477]_ ;
  assign \new_[725]_  = \new_[45464]_  & \new_[45451]_ ;
  assign \new_[726]_  = \new_[45438]_  & \new_[45425]_ ;
  assign \new_[727]_  = \new_[45412]_  & \new_[45399]_ ;
  assign \new_[728]_  = \new_[45386]_  & \new_[45373]_ ;
  assign \new_[729]_  = \new_[45360]_  & \new_[45347]_ ;
  assign \new_[730]_  = \new_[45334]_  & \new_[45321]_ ;
  assign \new_[731]_  = \new_[45308]_  & \new_[45295]_ ;
  assign \new_[732]_  = \new_[45282]_  & \new_[45269]_ ;
  assign \new_[733]_  = \new_[45256]_  & \new_[45243]_ ;
  assign \new_[734]_  = \new_[45230]_  & \new_[45217]_ ;
  assign \new_[735]_  = \new_[45204]_  & \new_[45191]_ ;
  assign \new_[736]_  = \new_[45178]_  & \new_[45165]_ ;
  assign \new_[737]_  = \new_[45152]_  & \new_[45139]_ ;
  assign \new_[738]_  = \new_[45126]_  & \new_[45113]_ ;
  assign \new_[739]_  = \new_[45100]_  & \new_[45087]_ ;
  assign \new_[740]_  = \new_[45074]_  & \new_[45061]_ ;
  assign \new_[741]_  = \new_[45048]_  & \new_[45035]_ ;
  assign \new_[742]_  = \new_[45022]_  & \new_[45009]_ ;
  assign \new_[743]_  = \new_[44996]_  & \new_[44983]_ ;
  assign \new_[744]_  = \new_[44970]_  & \new_[44957]_ ;
  assign \new_[745]_  = \new_[44944]_  & \new_[44931]_ ;
  assign \new_[746]_  = \new_[44918]_  & \new_[44905]_ ;
  assign \new_[747]_  = \new_[44892]_  & \new_[44879]_ ;
  assign \new_[748]_  = \new_[44866]_  & \new_[44853]_ ;
  assign \new_[749]_  = \new_[44840]_  & \new_[44827]_ ;
  assign \new_[750]_  = \new_[44814]_  & \new_[44801]_ ;
  assign \new_[751]_  = \new_[44788]_  & \new_[44775]_ ;
  assign \new_[752]_  = \new_[44762]_  & \new_[44749]_ ;
  assign \new_[753]_  = \new_[44736]_  & \new_[44723]_ ;
  assign \new_[754]_  = \new_[44710]_  & \new_[44697]_ ;
  assign \new_[755]_  = \new_[44684]_  & \new_[44671]_ ;
  assign \new_[756]_  = \new_[44658]_  & \new_[44645]_ ;
  assign \new_[757]_  = \new_[44632]_  & \new_[44619]_ ;
  assign \new_[758]_  = \new_[44606]_  & \new_[44593]_ ;
  assign \new_[759]_  = \new_[44580]_  & \new_[44567]_ ;
  assign \new_[760]_  = \new_[44554]_  & \new_[44541]_ ;
  assign \new_[761]_  = \new_[44528]_  & \new_[44515]_ ;
  assign \new_[762]_  = \new_[44502]_  & \new_[44489]_ ;
  assign \new_[763]_  = \new_[44476]_  & \new_[44463]_ ;
  assign \new_[764]_  = \new_[44450]_  & \new_[44437]_ ;
  assign \new_[765]_  = \new_[44424]_  & \new_[44411]_ ;
  assign \new_[766]_  = \new_[44398]_  & \new_[44385]_ ;
  assign \new_[767]_  = \new_[44372]_  & \new_[44359]_ ;
  assign \new_[768]_  = \new_[44346]_  & \new_[44333]_ ;
  assign \new_[769]_  = \new_[44320]_  & \new_[44307]_ ;
  assign \new_[770]_  = \new_[44294]_  & \new_[44281]_ ;
  assign \new_[771]_  = \new_[44268]_  & \new_[44255]_ ;
  assign \new_[772]_  = \new_[44242]_  & \new_[44229]_ ;
  assign \new_[773]_  = \new_[44216]_  & \new_[44203]_ ;
  assign \new_[774]_  = \new_[44190]_  & \new_[44177]_ ;
  assign \new_[775]_  = \new_[44164]_  & \new_[44151]_ ;
  assign \new_[776]_  = \new_[44138]_  & \new_[44125]_ ;
  assign \new_[777]_  = \new_[44112]_  & \new_[44099]_ ;
  assign \new_[778]_  = \new_[44086]_  & \new_[44073]_ ;
  assign \new_[779]_  = \new_[44060]_  & \new_[44047]_ ;
  assign \new_[780]_  = \new_[44034]_  & \new_[44021]_ ;
  assign \new_[781]_  = \new_[44008]_  & \new_[43995]_ ;
  assign \new_[782]_  = \new_[43982]_  & \new_[43969]_ ;
  assign \new_[783]_  = \new_[43956]_  & \new_[43943]_ ;
  assign \new_[784]_  = \new_[43930]_  & \new_[43917]_ ;
  assign \new_[785]_  = \new_[43904]_  & \new_[43891]_ ;
  assign \new_[786]_  = \new_[43878]_  & \new_[43865]_ ;
  assign \new_[787]_  = \new_[43852]_  & \new_[43839]_ ;
  assign \new_[788]_  = \new_[43826]_  & \new_[43813]_ ;
  assign \new_[789]_  = \new_[43800]_  & \new_[43787]_ ;
  assign \new_[790]_  = \new_[43774]_  & \new_[43761]_ ;
  assign \new_[791]_  = \new_[43748]_  & \new_[43735]_ ;
  assign \new_[792]_  = \new_[43722]_  & \new_[43709]_ ;
  assign \new_[793]_  = \new_[43696]_  & \new_[43683]_ ;
  assign \new_[794]_  = \new_[43670]_  & \new_[43657]_ ;
  assign \new_[795]_  = \new_[43644]_  & \new_[43631]_ ;
  assign \new_[796]_  = \new_[43618]_  & \new_[43605]_ ;
  assign \new_[797]_  = \new_[43592]_  & \new_[43579]_ ;
  assign \new_[798]_  = \new_[43566]_  & \new_[43553]_ ;
  assign \new_[799]_  = \new_[43540]_  & \new_[43527]_ ;
  assign \new_[800]_  = \new_[43514]_  & \new_[43501]_ ;
  assign \new_[801]_  = \new_[43488]_  & \new_[43475]_ ;
  assign \new_[802]_  = \new_[43462]_  & \new_[43449]_ ;
  assign \new_[803]_  = \new_[43436]_  & \new_[43423]_ ;
  assign \new_[804]_  = \new_[43410]_  & \new_[43397]_ ;
  assign \new_[805]_  = \new_[43384]_  & \new_[43371]_ ;
  assign \new_[806]_  = \new_[43358]_  & \new_[43345]_ ;
  assign \new_[807]_  = \new_[43332]_  & \new_[43319]_ ;
  assign \new_[808]_  = \new_[43306]_  & \new_[43293]_ ;
  assign \new_[809]_  = \new_[43280]_  & \new_[43267]_ ;
  assign \new_[810]_  = \new_[43254]_  & \new_[43241]_ ;
  assign \new_[811]_  = \new_[43228]_  & \new_[43215]_ ;
  assign \new_[812]_  = \new_[43202]_  & \new_[43189]_ ;
  assign \new_[813]_  = \new_[43176]_  & \new_[43163]_ ;
  assign \new_[814]_  = \new_[43150]_  & \new_[43137]_ ;
  assign \new_[815]_  = \new_[43124]_  & \new_[43111]_ ;
  assign \new_[816]_  = \new_[43098]_  & \new_[43085]_ ;
  assign \new_[817]_  = \new_[43072]_  & \new_[43059]_ ;
  assign \new_[818]_  = \new_[43046]_  & \new_[43033]_ ;
  assign \new_[819]_  = \new_[43020]_  & \new_[43007]_ ;
  assign \new_[820]_  = \new_[42994]_  & \new_[42981]_ ;
  assign \new_[821]_  = \new_[42968]_  & \new_[42955]_ ;
  assign \new_[822]_  = \new_[42942]_  & \new_[42929]_ ;
  assign \new_[823]_  = \new_[42916]_  & \new_[42903]_ ;
  assign \new_[824]_  = \new_[42890]_  & \new_[42877]_ ;
  assign \new_[825]_  = \new_[42864]_  & \new_[42851]_ ;
  assign \new_[826]_  = \new_[42838]_  & \new_[42825]_ ;
  assign \new_[827]_  = \new_[42812]_  & \new_[42799]_ ;
  assign \new_[828]_  = \new_[42786]_  & \new_[42773]_ ;
  assign \new_[829]_  = \new_[42760]_  & \new_[42747]_ ;
  assign \new_[830]_  = \new_[42734]_  & \new_[42721]_ ;
  assign \new_[831]_  = \new_[42708]_  & \new_[42695]_ ;
  assign \new_[832]_  = \new_[42682]_  & \new_[42669]_ ;
  assign \new_[833]_  = \new_[42656]_  & \new_[42643]_ ;
  assign \new_[834]_  = \new_[42630]_  & \new_[42617]_ ;
  assign \new_[835]_  = \new_[42604]_  & \new_[42591]_ ;
  assign \new_[836]_  = \new_[42578]_  & \new_[42565]_ ;
  assign \new_[837]_  = \new_[42552]_  & \new_[42539]_ ;
  assign \new_[838]_  = \new_[42526]_  & \new_[42513]_ ;
  assign \new_[839]_  = \new_[42500]_  & \new_[42487]_ ;
  assign \new_[840]_  = \new_[42474]_  & \new_[42461]_ ;
  assign \new_[841]_  = \new_[42448]_  & \new_[42435]_ ;
  assign \new_[842]_  = \new_[42422]_  & \new_[42409]_ ;
  assign \new_[843]_  = \new_[42396]_  & \new_[42383]_ ;
  assign \new_[844]_  = \new_[42370]_  & \new_[42357]_ ;
  assign \new_[845]_  = \new_[42344]_  & \new_[42331]_ ;
  assign \new_[846]_  = \new_[42318]_  & \new_[42305]_ ;
  assign \new_[847]_  = \new_[42292]_  & \new_[42279]_ ;
  assign \new_[848]_  = \new_[42266]_  & \new_[42253]_ ;
  assign \new_[849]_  = \new_[42240]_  & \new_[42227]_ ;
  assign \new_[850]_  = \new_[42214]_  & \new_[42201]_ ;
  assign \new_[851]_  = \new_[42188]_  & \new_[42175]_ ;
  assign \new_[852]_  = \new_[42162]_  & \new_[42149]_ ;
  assign \new_[853]_  = \new_[42136]_  & \new_[42123]_ ;
  assign \new_[854]_  = \new_[42110]_  & \new_[42097]_ ;
  assign \new_[855]_  = \new_[42084]_  & \new_[42071]_ ;
  assign \new_[856]_  = \new_[42058]_  & \new_[42045]_ ;
  assign \new_[857]_  = \new_[42032]_  & \new_[42019]_ ;
  assign \new_[858]_  = \new_[42006]_  & \new_[41993]_ ;
  assign \new_[859]_  = \new_[41980]_  & \new_[41967]_ ;
  assign \new_[860]_  = \new_[41954]_  & \new_[41941]_ ;
  assign \new_[861]_  = \new_[41928]_  & \new_[41915]_ ;
  assign \new_[862]_  = \new_[41902]_  & \new_[41889]_ ;
  assign \new_[863]_  = \new_[41876]_  & \new_[41863]_ ;
  assign \new_[864]_  = \new_[41850]_  & \new_[41837]_ ;
  assign \new_[865]_  = \new_[41824]_  & \new_[41811]_ ;
  assign \new_[866]_  = \new_[41798]_  & \new_[41785]_ ;
  assign \new_[867]_  = \new_[41772]_  & \new_[41759]_ ;
  assign \new_[868]_  = \new_[41746]_  & \new_[41733]_ ;
  assign \new_[869]_  = \new_[41720]_  & \new_[41707]_ ;
  assign \new_[870]_  = \new_[41694]_  & \new_[41681]_ ;
  assign \new_[871]_  = \new_[41668]_  & \new_[41655]_ ;
  assign \new_[872]_  = \new_[41642]_  & \new_[41629]_ ;
  assign \new_[873]_  = \new_[41616]_  & \new_[41603]_ ;
  assign \new_[874]_  = \new_[41590]_  & \new_[41577]_ ;
  assign \new_[875]_  = \new_[41564]_  & \new_[41551]_ ;
  assign \new_[876]_  = \new_[41538]_  & \new_[41525]_ ;
  assign \new_[877]_  = \new_[41512]_  & \new_[41499]_ ;
  assign \new_[878]_  = \new_[41486]_  & \new_[41473]_ ;
  assign \new_[879]_  = \new_[41460]_  & \new_[41447]_ ;
  assign \new_[880]_  = \new_[41434]_  & \new_[41421]_ ;
  assign \new_[881]_  = \new_[41408]_  & \new_[41395]_ ;
  assign \new_[882]_  = \new_[41382]_  & \new_[41369]_ ;
  assign \new_[883]_  = \new_[41356]_  & \new_[41343]_ ;
  assign \new_[884]_  = \new_[41330]_  & \new_[41317]_ ;
  assign \new_[885]_  = \new_[41304]_  & \new_[41291]_ ;
  assign \new_[886]_  = \new_[41278]_  & \new_[41265]_ ;
  assign \new_[887]_  = \new_[41252]_  & \new_[41239]_ ;
  assign \new_[888]_  = \new_[41226]_  & \new_[41213]_ ;
  assign \new_[889]_  = \new_[41200]_  & \new_[41187]_ ;
  assign \new_[890]_  = \new_[41174]_  & \new_[41161]_ ;
  assign \new_[891]_  = \new_[41148]_  & \new_[41135]_ ;
  assign \new_[892]_  = \new_[41122]_  & \new_[41109]_ ;
  assign \new_[893]_  = \new_[41096]_  & \new_[41083]_ ;
  assign \new_[894]_  = \new_[41070]_  & \new_[41057]_ ;
  assign \new_[895]_  = \new_[41044]_  & \new_[41031]_ ;
  assign \new_[896]_  = \new_[41018]_  & \new_[41005]_ ;
  assign \new_[897]_  = \new_[40992]_  & \new_[40979]_ ;
  assign \new_[898]_  = \new_[40966]_  & \new_[40953]_ ;
  assign \new_[899]_  = \new_[40940]_  & \new_[40927]_ ;
  assign \new_[900]_  = \new_[40914]_  & \new_[40901]_ ;
  assign \new_[901]_  = \new_[40888]_  & \new_[40875]_ ;
  assign \new_[902]_  = \new_[40862]_  & \new_[40849]_ ;
  assign \new_[903]_  = \new_[40836]_  & \new_[40823]_ ;
  assign \new_[904]_  = \new_[40810]_  & \new_[40797]_ ;
  assign \new_[905]_  = \new_[40784]_  & \new_[40771]_ ;
  assign \new_[906]_  = \new_[40758]_  & \new_[40745]_ ;
  assign \new_[907]_  = \new_[40732]_  & \new_[40719]_ ;
  assign \new_[908]_  = \new_[40706]_  & \new_[40693]_ ;
  assign \new_[909]_  = \new_[40680]_  & \new_[40667]_ ;
  assign \new_[910]_  = \new_[40654]_  & \new_[40641]_ ;
  assign \new_[911]_  = \new_[40628]_  & \new_[40615]_ ;
  assign \new_[912]_  = \new_[40602]_  & \new_[40589]_ ;
  assign \new_[913]_  = \new_[40576]_  & \new_[40563]_ ;
  assign \new_[914]_  = \new_[40550]_  & \new_[40537]_ ;
  assign \new_[915]_  = \new_[40524]_  & \new_[40511]_ ;
  assign \new_[916]_  = \new_[40498]_  & \new_[40485]_ ;
  assign \new_[917]_  = \new_[40472]_  & \new_[40459]_ ;
  assign \new_[918]_  = \new_[40446]_  & \new_[40433]_ ;
  assign \new_[919]_  = \new_[40420]_  & \new_[40407]_ ;
  assign \new_[920]_  = \new_[40394]_  & \new_[40381]_ ;
  assign \new_[921]_  = \new_[40368]_  & \new_[40355]_ ;
  assign \new_[922]_  = \new_[40342]_  & \new_[40329]_ ;
  assign \new_[923]_  = \new_[40316]_  & \new_[40303]_ ;
  assign \new_[924]_  = \new_[40290]_  & \new_[40277]_ ;
  assign \new_[925]_  = \new_[40264]_  & \new_[40251]_ ;
  assign \new_[926]_  = \new_[40238]_  & \new_[40225]_ ;
  assign \new_[927]_  = \new_[40212]_  & \new_[40199]_ ;
  assign \new_[928]_  = \new_[40186]_  & \new_[40173]_ ;
  assign \new_[929]_  = \new_[40160]_  & \new_[40147]_ ;
  assign \new_[930]_  = \new_[40134]_  & \new_[40121]_ ;
  assign \new_[931]_  = \new_[40108]_  & \new_[40095]_ ;
  assign \new_[932]_  = \new_[40082]_  & \new_[40069]_ ;
  assign \new_[933]_  = \new_[40056]_  & \new_[40043]_ ;
  assign \new_[934]_  = \new_[40030]_  & \new_[40017]_ ;
  assign \new_[935]_  = \new_[40004]_  & \new_[39991]_ ;
  assign \new_[936]_  = \new_[39978]_  & \new_[39965]_ ;
  assign \new_[937]_  = \new_[39952]_  & \new_[39939]_ ;
  assign \new_[938]_  = \new_[39926]_  & \new_[39913]_ ;
  assign \new_[939]_  = \new_[39900]_  & \new_[39887]_ ;
  assign \new_[940]_  = \new_[39874]_  & \new_[39861]_ ;
  assign \new_[941]_  = \new_[39848]_  & \new_[39835]_ ;
  assign \new_[942]_  = \new_[39822]_  & \new_[39809]_ ;
  assign \new_[943]_  = \new_[39796]_  & \new_[39783]_ ;
  assign \new_[944]_  = \new_[39770]_  & \new_[39757]_ ;
  assign \new_[945]_  = \new_[39744]_  & \new_[39731]_ ;
  assign \new_[946]_  = \new_[39718]_  & \new_[39705]_ ;
  assign \new_[947]_  = \new_[39692]_  & \new_[39679]_ ;
  assign \new_[948]_  = \new_[39666]_  & \new_[39653]_ ;
  assign \new_[949]_  = \new_[39640]_  & \new_[39627]_ ;
  assign \new_[950]_  = \new_[39614]_  & \new_[39601]_ ;
  assign \new_[951]_  = \new_[39588]_  & \new_[39575]_ ;
  assign \new_[952]_  = \new_[39562]_  & \new_[39549]_ ;
  assign \new_[953]_  = \new_[39536]_  & \new_[39523]_ ;
  assign \new_[954]_  = \new_[39510]_  & \new_[39497]_ ;
  assign \new_[955]_  = \new_[39484]_  & \new_[39471]_ ;
  assign \new_[956]_  = \new_[39458]_  & \new_[39445]_ ;
  assign \new_[957]_  = \new_[39432]_  & \new_[39419]_ ;
  assign \new_[958]_  = \new_[39406]_  & \new_[39393]_ ;
  assign \new_[959]_  = \new_[39380]_  & \new_[39367]_ ;
  assign \new_[960]_  = \new_[39354]_  & \new_[39341]_ ;
  assign \new_[961]_  = \new_[39328]_  & \new_[39315]_ ;
  assign \new_[962]_  = \new_[39302]_  & \new_[39289]_ ;
  assign \new_[963]_  = \new_[39276]_  & \new_[39263]_ ;
  assign \new_[964]_  = \new_[39250]_  & \new_[39237]_ ;
  assign \new_[965]_  = \new_[39224]_  & \new_[39211]_ ;
  assign \new_[966]_  = \new_[39198]_  & \new_[39185]_ ;
  assign \new_[967]_  = \new_[39172]_  & \new_[39159]_ ;
  assign \new_[968]_  = \new_[39146]_  & \new_[39133]_ ;
  assign \new_[969]_  = \new_[39120]_  & \new_[39107]_ ;
  assign \new_[970]_  = \new_[39094]_  & \new_[39081]_ ;
  assign \new_[971]_  = \new_[39068]_  & \new_[39055]_ ;
  assign \new_[972]_  = \new_[39042]_  & \new_[39029]_ ;
  assign \new_[973]_  = \new_[39016]_  & \new_[39003]_ ;
  assign \new_[974]_  = \new_[38990]_  & \new_[38977]_ ;
  assign \new_[975]_  = \new_[38964]_  & \new_[38951]_ ;
  assign \new_[976]_  = \new_[38938]_  & \new_[38925]_ ;
  assign \new_[977]_  = \new_[38912]_  & \new_[38899]_ ;
  assign \new_[978]_  = \new_[38886]_  & \new_[38873]_ ;
  assign \new_[979]_  = \new_[38860]_  & \new_[38847]_ ;
  assign \new_[980]_  = \new_[38834]_  & \new_[38821]_ ;
  assign \new_[981]_  = \new_[38808]_  & \new_[38795]_ ;
  assign \new_[982]_  = \new_[38782]_  & \new_[38769]_ ;
  assign \new_[983]_  = \new_[38756]_  & \new_[38743]_ ;
  assign \new_[984]_  = \new_[38730]_  & \new_[38717]_ ;
  assign \new_[985]_  = \new_[38704]_  & \new_[38691]_ ;
  assign \new_[986]_  = \new_[38678]_  & \new_[38665]_ ;
  assign \new_[987]_  = \new_[38652]_  & \new_[38639]_ ;
  assign \new_[988]_  = \new_[38626]_  & \new_[38613]_ ;
  assign \new_[989]_  = \new_[38600]_  & \new_[38587]_ ;
  assign \new_[990]_  = \new_[38574]_  & \new_[38561]_ ;
  assign \new_[991]_  = \new_[38548]_  & \new_[38535]_ ;
  assign \new_[992]_  = \new_[38522]_  & \new_[38509]_ ;
  assign \new_[993]_  = \new_[38496]_  & \new_[38483]_ ;
  assign \new_[994]_  = \new_[38470]_  & \new_[38457]_ ;
  assign \new_[995]_  = \new_[38444]_  & \new_[38431]_ ;
  assign \new_[996]_  = \new_[38418]_  & \new_[38405]_ ;
  assign \new_[997]_  = \new_[38392]_  & \new_[38379]_ ;
  assign \new_[998]_  = \new_[38366]_  & \new_[38353]_ ;
  assign \new_[999]_  = \new_[38340]_  & \new_[38327]_ ;
  assign \new_[1000]_  = \new_[38314]_  & \new_[38301]_ ;
  assign \new_[1001]_  = \new_[38288]_  & \new_[38275]_ ;
  assign \new_[1002]_  = \new_[38262]_  & \new_[38249]_ ;
  assign \new_[1003]_  = \new_[38236]_  & \new_[38223]_ ;
  assign \new_[1004]_  = \new_[38210]_  & \new_[38197]_ ;
  assign \new_[1005]_  = \new_[38184]_  & \new_[38171]_ ;
  assign \new_[1006]_  = \new_[38158]_  & \new_[38145]_ ;
  assign \new_[1007]_  = \new_[38132]_  & \new_[38119]_ ;
  assign \new_[1008]_  = \new_[38106]_  & \new_[38093]_ ;
  assign \new_[1009]_  = \new_[38080]_  & \new_[38067]_ ;
  assign \new_[1010]_  = \new_[38054]_  & \new_[38041]_ ;
  assign \new_[1011]_  = \new_[38028]_  & \new_[38015]_ ;
  assign \new_[1012]_  = \new_[38002]_  & \new_[37989]_ ;
  assign \new_[1013]_  = \new_[37976]_  & \new_[37963]_ ;
  assign \new_[1014]_  = \new_[37950]_  & \new_[37937]_ ;
  assign \new_[1015]_  = \new_[37924]_  & \new_[37911]_ ;
  assign \new_[1016]_  = \new_[37898]_  & \new_[37885]_ ;
  assign \new_[1017]_  = \new_[37872]_  & \new_[37859]_ ;
  assign \new_[1018]_  = \new_[37846]_  & \new_[37833]_ ;
  assign \new_[1019]_  = \new_[37820]_  & \new_[37807]_ ;
  assign \new_[1020]_  = \new_[37796]_  & \new_[37783]_ ;
  assign \new_[1021]_  = \new_[37772]_  & \new_[37759]_ ;
  assign \new_[1022]_  = \new_[37748]_  & \new_[37735]_ ;
  assign \new_[1023]_  = \new_[37724]_  & \new_[37711]_ ;
  assign \new_[1024]_  = \new_[37700]_  & \new_[37687]_ ;
  assign \new_[1025]_  = \new_[37676]_  & \new_[37663]_ ;
  assign \new_[1026]_  = \new_[37652]_  & \new_[37639]_ ;
  assign \new_[1027]_  = \new_[37628]_  & \new_[37615]_ ;
  assign \new_[1028]_  = \new_[37604]_  & \new_[37591]_ ;
  assign \new_[1029]_  = \new_[37580]_  & \new_[37567]_ ;
  assign \new_[1030]_  = \new_[37556]_  & \new_[37543]_ ;
  assign \new_[1031]_  = \new_[37532]_  & \new_[37519]_ ;
  assign \new_[1032]_  = \new_[37508]_  & \new_[37495]_ ;
  assign \new_[1033]_  = \new_[37484]_  & \new_[37471]_ ;
  assign \new_[1034]_  = \new_[37460]_  & \new_[37447]_ ;
  assign \new_[1035]_  = \new_[37436]_  & \new_[37423]_ ;
  assign \new_[1036]_  = \new_[37412]_  & \new_[37399]_ ;
  assign \new_[1037]_  = \new_[37388]_  & \new_[37375]_ ;
  assign \new_[1038]_  = \new_[37364]_  & \new_[37351]_ ;
  assign \new_[1039]_  = \new_[37340]_  & \new_[37327]_ ;
  assign \new_[1040]_  = \new_[37316]_  & \new_[37303]_ ;
  assign \new_[1041]_  = \new_[37292]_  & \new_[37279]_ ;
  assign \new_[1042]_  = \new_[37268]_  & \new_[37255]_ ;
  assign \new_[1043]_  = \new_[37244]_  & \new_[37231]_ ;
  assign \new_[1044]_  = \new_[37220]_  & \new_[37207]_ ;
  assign \new_[1045]_  = \new_[37196]_  & \new_[37183]_ ;
  assign \new_[1046]_  = \new_[37172]_  & \new_[37159]_ ;
  assign \new_[1047]_  = \new_[37148]_  & \new_[37135]_ ;
  assign \new_[1048]_  = \new_[37124]_  & \new_[37111]_ ;
  assign \new_[1049]_  = \new_[37100]_  & \new_[37087]_ ;
  assign \new_[1050]_  = \new_[37076]_  & \new_[37063]_ ;
  assign \new_[1051]_  = \new_[37052]_  & \new_[37039]_ ;
  assign \new_[1052]_  = \new_[37028]_  & \new_[37015]_ ;
  assign \new_[1053]_  = \new_[37004]_  & \new_[36991]_ ;
  assign \new_[1054]_  = \new_[36980]_  & \new_[36967]_ ;
  assign \new_[1055]_  = \new_[36956]_  & \new_[36943]_ ;
  assign \new_[1056]_  = \new_[36932]_  & \new_[36919]_ ;
  assign \new_[1057]_  = \new_[36908]_  & \new_[36895]_ ;
  assign \new_[1058]_  = \new_[36884]_  & \new_[36871]_ ;
  assign \new_[1059]_  = \new_[36860]_  & \new_[36847]_ ;
  assign \new_[1060]_  = \new_[36836]_  & \new_[36823]_ ;
  assign \new_[1061]_  = \new_[36812]_  & \new_[36799]_ ;
  assign \new_[1062]_  = \new_[36788]_  & \new_[36775]_ ;
  assign \new_[1063]_  = \new_[36764]_  & \new_[36751]_ ;
  assign \new_[1064]_  = \new_[36740]_  & \new_[36727]_ ;
  assign \new_[1065]_  = \new_[36716]_  & \new_[36703]_ ;
  assign \new_[1066]_  = \new_[36692]_  & \new_[36679]_ ;
  assign \new_[1067]_  = \new_[36668]_  & \new_[36655]_ ;
  assign \new_[1068]_  = \new_[36644]_  & \new_[36631]_ ;
  assign \new_[1069]_  = \new_[36620]_  & \new_[36607]_ ;
  assign \new_[1070]_  = \new_[36596]_  & \new_[36583]_ ;
  assign \new_[1071]_  = \new_[36572]_  & \new_[36559]_ ;
  assign \new_[1072]_  = \new_[36548]_  & \new_[36535]_ ;
  assign \new_[1073]_  = \new_[36524]_  & \new_[36511]_ ;
  assign \new_[1074]_  = \new_[36500]_  & \new_[36487]_ ;
  assign \new_[1075]_  = \new_[36476]_  & \new_[36463]_ ;
  assign \new_[1076]_  = \new_[36452]_  & \new_[36439]_ ;
  assign \new_[1077]_  = \new_[36428]_  & \new_[36415]_ ;
  assign \new_[1078]_  = \new_[36404]_  & \new_[36391]_ ;
  assign \new_[1079]_  = \new_[36380]_  & \new_[36367]_ ;
  assign \new_[1080]_  = \new_[36356]_  & \new_[36343]_ ;
  assign \new_[1081]_  = \new_[36332]_  & \new_[36319]_ ;
  assign \new_[1082]_  = \new_[36308]_  & \new_[36295]_ ;
  assign \new_[1083]_  = \new_[36284]_  & \new_[36271]_ ;
  assign \new_[1084]_  = \new_[36260]_  & \new_[36247]_ ;
  assign \new_[1085]_  = \new_[36236]_  & \new_[36223]_ ;
  assign \new_[1086]_  = \new_[36212]_  & \new_[36199]_ ;
  assign \new_[1087]_  = \new_[36188]_  & \new_[36175]_ ;
  assign \new_[1088]_  = \new_[36164]_  & \new_[36151]_ ;
  assign \new_[1089]_  = \new_[36140]_  & \new_[36127]_ ;
  assign \new_[1090]_  = \new_[36116]_  & \new_[36103]_ ;
  assign \new_[1091]_  = \new_[36092]_  & \new_[36079]_ ;
  assign \new_[1092]_  = \new_[36068]_  & \new_[36055]_ ;
  assign \new_[1093]_  = \new_[36044]_  & \new_[36031]_ ;
  assign \new_[1094]_  = \new_[36020]_  & \new_[36007]_ ;
  assign \new_[1095]_  = \new_[35996]_  & \new_[35983]_ ;
  assign \new_[1096]_  = \new_[35972]_  & \new_[35959]_ ;
  assign \new_[1097]_  = \new_[35948]_  & \new_[35935]_ ;
  assign \new_[1098]_  = \new_[35924]_  & \new_[35911]_ ;
  assign \new_[1099]_  = \new_[35900]_  & \new_[35887]_ ;
  assign \new_[1100]_  = \new_[35876]_  & \new_[35863]_ ;
  assign \new_[1101]_  = \new_[35852]_  & \new_[35839]_ ;
  assign \new_[1102]_  = \new_[35828]_  & \new_[35815]_ ;
  assign \new_[1103]_  = \new_[35804]_  & \new_[35791]_ ;
  assign \new_[1104]_  = \new_[35780]_  & \new_[35767]_ ;
  assign \new_[1105]_  = \new_[35756]_  & \new_[35743]_ ;
  assign \new_[1106]_  = \new_[35732]_  & \new_[35719]_ ;
  assign \new_[1107]_  = \new_[35708]_  & \new_[35695]_ ;
  assign \new_[1108]_  = \new_[35684]_  & \new_[35671]_ ;
  assign \new_[1109]_  = \new_[35660]_  & \new_[35647]_ ;
  assign \new_[1110]_  = \new_[35636]_  & \new_[35623]_ ;
  assign \new_[1111]_  = \new_[35612]_  & \new_[35599]_ ;
  assign \new_[1112]_  = \new_[35588]_  & \new_[35575]_ ;
  assign \new_[1113]_  = \new_[35564]_  & \new_[35551]_ ;
  assign \new_[1114]_  = \new_[35540]_  & \new_[35527]_ ;
  assign \new_[1115]_  = \new_[35516]_  & \new_[35503]_ ;
  assign \new_[1116]_  = \new_[35492]_  & \new_[35479]_ ;
  assign \new_[1117]_  = \new_[35468]_  & \new_[35455]_ ;
  assign \new_[1118]_  = \new_[35444]_  & \new_[35431]_ ;
  assign \new_[1119]_  = \new_[35420]_  & \new_[35407]_ ;
  assign \new_[1120]_  = \new_[35396]_  & \new_[35383]_ ;
  assign \new_[1121]_  = \new_[35372]_  & \new_[35359]_ ;
  assign \new_[1122]_  = \new_[35348]_  & \new_[35335]_ ;
  assign \new_[1123]_  = \new_[35324]_  & \new_[35311]_ ;
  assign \new_[1124]_  = \new_[35300]_  & \new_[35287]_ ;
  assign \new_[1125]_  = \new_[35276]_  & \new_[35263]_ ;
  assign \new_[1126]_  = \new_[35252]_  & \new_[35239]_ ;
  assign \new_[1127]_  = \new_[35228]_  & \new_[35215]_ ;
  assign \new_[1128]_  = \new_[35204]_  & \new_[35191]_ ;
  assign \new_[1129]_  = \new_[35180]_  & \new_[35167]_ ;
  assign \new_[1130]_  = \new_[35156]_  & \new_[35143]_ ;
  assign \new_[1131]_  = \new_[35132]_  & \new_[35119]_ ;
  assign \new_[1132]_  = \new_[35108]_  & \new_[35095]_ ;
  assign \new_[1133]_  = \new_[35084]_  & \new_[35071]_ ;
  assign \new_[1134]_  = \new_[35060]_  & \new_[35047]_ ;
  assign \new_[1135]_  = \new_[35036]_  & \new_[35023]_ ;
  assign \new_[1136]_  = \new_[35012]_  & \new_[34999]_ ;
  assign \new_[1137]_  = \new_[34988]_  & \new_[34975]_ ;
  assign \new_[1138]_  = \new_[34964]_  & \new_[34951]_ ;
  assign \new_[1139]_  = \new_[34940]_  & \new_[34927]_ ;
  assign \new_[1140]_  = \new_[34916]_  & \new_[34903]_ ;
  assign \new_[1141]_  = \new_[34892]_  & \new_[34879]_ ;
  assign \new_[1142]_  = \new_[34868]_  & \new_[34855]_ ;
  assign \new_[1143]_  = \new_[34844]_  & \new_[34831]_ ;
  assign \new_[1144]_  = \new_[34820]_  & \new_[34807]_ ;
  assign \new_[1145]_  = \new_[34796]_  & \new_[34783]_ ;
  assign \new_[1146]_  = \new_[34772]_  & \new_[34759]_ ;
  assign \new_[1147]_  = \new_[34748]_  & \new_[34735]_ ;
  assign \new_[1148]_  = \new_[34724]_  & \new_[34711]_ ;
  assign \new_[1149]_  = \new_[34700]_  & \new_[34687]_ ;
  assign \new_[1150]_  = \new_[34676]_  & \new_[34663]_ ;
  assign \new_[1151]_  = \new_[34652]_  & \new_[34639]_ ;
  assign \new_[1152]_  = \new_[34628]_  & \new_[34615]_ ;
  assign \new_[1153]_  = \new_[34604]_  & \new_[34591]_ ;
  assign \new_[1154]_  = \new_[34580]_  & \new_[34567]_ ;
  assign \new_[1155]_  = \new_[34556]_  & \new_[34543]_ ;
  assign \new_[1156]_  = \new_[34532]_  & \new_[34519]_ ;
  assign \new_[1157]_  = \new_[34508]_  & \new_[34495]_ ;
  assign \new_[1158]_  = \new_[34484]_  & \new_[34471]_ ;
  assign \new_[1159]_  = \new_[34460]_  & \new_[34447]_ ;
  assign \new_[1160]_  = \new_[34436]_  & \new_[34423]_ ;
  assign \new_[1161]_  = \new_[34412]_  & \new_[34399]_ ;
  assign \new_[1162]_  = \new_[34388]_  & \new_[34375]_ ;
  assign \new_[1163]_  = \new_[34364]_  & \new_[34351]_ ;
  assign \new_[1164]_  = \new_[34340]_  & \new_[34327]_ ;
  assign \new_[1165]_  = \new_[34316]_  & \new_[34303]_ ;
  assign \new_[1166]_  = \new_[34292]_  & \new_[34279]_ ;
  assign \new_[1167]_  = \new_[34268]_  & \new_[34255]_ ;
  assign \new_[1168]_  = \new_[34244]_  & \new_[34231]_ ;
  assign \new_[1169]_  = \new_[34220]_  & \new_[34207]_ ;
  assign \new_[1170]_  = \new_[34196]_  & \new_[34183]_ ;
  assign \new_[1171]_  = \new_[34172]_  & \new_[34159]_ ;
  assign \new_[1172]_  = \new_[34148]_  & \new_[34135]_ ;
  assign \new_[1173]_  = \new_[34124]_  & \new_[34111]_ ;
  assign \new_[1174]_  = \new_[34100]_  & \new_[34087]_ ;
  assign \new_[1175]_  = \new_[34076]_  & \new_[34063]_ ;
  assign \new_[1176]_  = \new_[34052]_  & \new_[34039]_ ;
  assign \new_[1177]_  = \new_[34028]_  & \new_[34015]_ ;
  assign \new_[1178]_  = \new_[34004]_  & \new_[33991]_ ;
  assign \new_[1179]_  = \new_[33980]_  & \new_[33967]_ ;
  assign \new_[1180]_  = \new_[33956]_  & \new_[33943]_ ;
  assign \new_[1181]_  = \new_[33932]_  & \new_[33919]_ ;
  assign \new_[1182]_  = \new_[33908]_  & \new_[33895]_ ;
  assign \new_[1183]_  = \new_[33884]_  & \new_[33871]_ ;
  assign \new_[1184]_  = \new_[33860]_  & \new_[33847]_ ;
  assign \new_[1185]_  = \new_[33836]_  & \new_[33823]_ ;
  assign \new_[1186]_  = \new_[33812]_  & \new_[33799]_ ;
  assign \new_[1187]_  = \new_[33788]_  & \new_[33775]_ ;
  assign \new_[1188]_  = \new_[33764]_  & \new_[33751]_ ;
  assign \new_[1189]_  = \new_[33740]_  & \new_[33727]_ ;
  assign \new_[1190]_  = \new_[33716]_  & \new_[33703]_ ;
  assign \new_[1191]_  = \new_[33692]_  & \new_[33679]_ ;
  assign \new_[1192]_  = \new_[33668]_  & \new_[33655]_ ;
  assign \new_[1193]_  = \new_[33644]_  & \new_[33631]_ ;
  assign \new_[1194]_  = \new_[33620]_  & \new_[33607]_ ;
  assign \new_[1195]_  = \new_[33596]_  & \new_[33583]_ ;
  assign \new_[1196]_  = \new_[33572]_  & \new_[33559]_ ;
  assign \new_[1197]_  = \new_[33548]_  & \new_[33535]_ ;
  assign \new_[1198]_  = \new_[33524]_  & \new_[33511]_ ;
  assign \new_[1199]_  = \new_[33500]_  & \new_[33487]_ ;
  assign \new_[1200]_  = \new_[33476]_  & \new_[33463]_ ;
  assign \new_[1201]_  = \new_[33452]_  & \new_[33439]_ ;
  assign \new_[1202]_  = \new_[33428]_  & \new_[33415]_ ;
  assign \new_[1203]_  = \new_[33404]_  & \new_[33391]_ ;
  assign \new_[1204]_  = \new_[33380]_  & \new_[33367]_ ;
  assign \new_[1205]_  = \new_[33356]_  & \new_[33343]_ ;
  assign \new_[1206]_  = \new_[33332]_  & \new_[33319]_ ;
  assign \new_[1207]_  = \new_[33308]_  & \new_[33295]_ ;
  assign \new_[1208]_  = \new_[33284]_  & \new_[33271]_ ;
  assign \new_[1209]_  = \new_[33260]_  & \new_[33247]_ ;
  assign \new_[1210]_  = \new_[33236]_  & \new_[33223]_ ;
  assign \new_[1211]_  = \new_[33212]_  & \new_[33199]_ ;
  assign \new_[1212]_  = \new_[33188]_  & \new_[33175]_ ;
  assign \new_[1213]_  = \new_[33164]_  & \new_[33151]_ ;
  assign \new_[1214]_  = \new_[33140]_  & \new_[33127]_ ;
  assign \new_[1215]_  = \new_[33116]_  & \new_[33103]_ ;
  assign \new_[1216]_  = \new_[33092]_  & \new_[33079]_ ;
  assign \new_[1217]_  = \new_[33068]_  & \new_[33055]_ ;
  assign \new_[1218]_  = \new_[33044]_  & \new_[33031]_ ;
  assign \new_[1219]_  = \new_[33020]_  & \new_[33007]_ ;
  assign \new_[1220]_  = \new_[32996]_  & \new_[32983]_ ;
  assign \new_[1221]_  = \new_[32972]_  & \new_[32959]_ ;
  assign \new_[1222]_  = \new_[32948]_  & \new_[32935]_ ;
  assign \new_[1223]_  = \new_[32924]_  & \new_[32911]_ ;
  assign \new_[1224]_  = \new_[32900]_  & \new_[32887]_ ;
  assign \new_[1225]_  = \new_[32876]_  & \new_[32863]_ ;
  assign \new_[1226]_  = \new_[32852]_  & \new_[32839]_ ;
  assign \new_[1227]_  = \new_[32828]_  & \new_[32815]_ ;
  assign \new_[1228]_  = \new_[32804]_  & \new_[32791]_ ;
  assign \new_[1229]_  = \new_[32780]_  & \new_[32767]_ ;
  assign \new_[1230]_  = \new_[32756]_  & \new_[32743]_ ;
  assign \new_[1231]_  = \new_[32732]_  & \new_[32719]_ ;
  assign \new_[1232]_  = \new_[32708]_  & \new_[32695]_ ;
  assign \new_[1233]_  = \new_[32684]_  & \new_[32671]_ ;
  assign \new_[1234]_  = \new_[32660]_  & \new_[32647]_ ;
  assign \new_[1235]_  = \new_[32636]_  & \new_[32623]_ ;
  assign \new_[1236]_  = \new_[32612]_  & \new_[32599]_ ;
  assign \new_[1237]_  = \new_[32588]_  & \new_[32575]_ ;
  assign \new_[1238]_  = \new_[32564]_  & \new_[32551]_ ;
  assign \new_[1239]_  = \new_[32540]_  & \new_[32527]_ ;
  assign \new_[1240]_  = \new_[32516]_  & \new_[32503]_ ;
  assign \new_[1241]_  = \new_[32492]_  & \new_[32479]_ ;
  assign \new_[1242]_  = \new_[32468]_  & \new_[32455]_ ;
  assign \new_[1243]_  = \new_[32444]_  & \new_[32431]_ ;
  assign \new_[1244]_  = \new_[32420]_  & \new_[32407]_ ;
  assign \new_[1245]_  = \new_[32396]_  & \new_[32383]_ ;
  assign \new_[1246]_  = \new_[32372]_  & \new_[32359]_ ;
  assign \new_[1247]_  = \new_[32348]_  & \new_[32335]_ ;
  assign \new_[1248]_  = \new_[32324]_  & \new_[32311]_ ;
  assign \new_[1249]_  = \new_[32300]_  & \new_[32287]_ ;
  assign \new_[1250]_  = \new_[32276]_  & \new_[32263]_ ;
  assign \new_[1251]_  = \new_[32252]_  & \new_[32239]_ ;
  assign \new_[1252]_  = \new_[32228]_  & \new_[32215]_ ;
  assign \new_[1253]_  = \new_[32204]_  & \new_[32191]_ ;
  assign \new_[1254]_  = \new_[32180]_  & \new_[32167]_ ;
  assign \new_[1255]_  = \new_[32156]_  & \new_[32143]_ ;
  assign \new_[1256]_  = \new_[32132]_  & \new_[32119]_ ;
  assign \new_[1257]_  = \new_[32108]_  & \new_[32095]_ ;
  assign \new_[1258]_  = \new_[32084]_  & \new_[32071]_ ;
  assign \new_[1259]_  = \new_[32060]_  & \new_[32047]_ ;
  assign \new_[1260]_  = \new_[32036]_  & \new_[32023]_ ;
  assign \new_[1261]_  = \new_[32012]_  & \new_[31999]_ ;
  assign \new_[1262]_  = \new_[31988]_  & \new_[31975]_ ;
  assign \new_[1263]_  = \new_[31964]_  & \new_[31951]_ ;
  assign \new_[1264]_  = \new_[31940]_  & \new_[31927]_ ;
  assign \new_[1265]_  = \new_[31916]_  & \new_[31903]_ ;
  assign \new_[1266]_  = \new_[31892]_  & \new_[31879]_ ;
  assign \new_[1267]_  = \new_[31868]_  & \new_[31855]_ ;
  assign \new_[1268]_  = \new_[31844]_  & \new_[31831]_ ;
  assign \new_[1269]_  = \new_[31820]_  & \new_[31807]_ ;
  assign \new_[1270]_  = \new_[31796]_  & \new_[31783]_ ;
  assign \new_[1271]_  = \new_[31772]_  & \new_[31759]_ ;
  assign \new_[1272]_  = \new_[31748]_  & \new_[31735]_ ;
  assign \new_[1273]_  = \new_[31724]_  & \new_[31711]_ ;
  assign \new_[1274]_  = \new_[31700]_  & \new_[31687]_ ;
  assign \new_[1275]_  = \new_[31676]_  & \new_[31663]_ ;
  assign \new_[1276]_  = \new_[31652]_  & \new_[31639]_ ;
  assign \new_[1277]_  = \new_[31628]_  & \new_[31615]_ ;
  assign \new_[1278]_  = \new_[31604]_  & \new_[31591]_ ;
  assign \new_[1279]_  = \new_[31580]_  & \new_[31567]_ ;
  assign \new_[1280]_  = \new_[31556]_  & \new_[31543]_ ;
  assign \new_[1281]_  = \new_[31532]_  & \new_[31519]_ ;
  assign \new_[1282]_  = \new_[31508]_  & \new_[31495]_ ;
  assign \new_[1283]_  = \new_[31484]_  & \new_[31471]_ ;
  assign \new_[1284]_  = \new_[31460]_  & \new_[31447]_ ;
  assign \new_[1285]_  = \new_[31436]_  & \new_[31423]_ ;
  assign \new_[1286]_  = \new_[31412]_  & \new_[31399]_ ;
  assign \new_[1287]_  = \new_[31388]_  & \new_[31375]_ ;
  assign \new_[1288]_  = \new_[31364]_  & \new_[31351]_ ;
  assign \new_[1289]_  = \new_[31340]_  & \new_[31327]_ ;
  assign \new_[1290]_  = \new_[31316]_  & \new_[31303]_ ;
  assign \new_[1291]_  = \new_[31292]_  & \new_[31279]_ ;
  assign \new_[1292]_  = \new_[31268]_  & \new_[31255]_ ;
  assign \new_[1293]_  = \new_[31244]_  & \new_[31231]_ ;
  assign \new_[1294]_  = \new_[31220]_  & \new_[31207]_ ;
  assign \new_[1295]_  = \new_[31196]_  & \new_[31183]_ ;
  assign \new_[1296]_  = \new_[31172]_  & \new_[31159]_ ;
  assign \new_[1297]_  = \new_[31148]_  & \new_[31135]_ ;
  assign \new_[1298]_  = \new_[31124]_  & \new_[31111]_ ;
  assign \new_[1299]_  = \new_[31100]_  & \new_[31087]_ ;
  assign \new_[1300]_  = \new_[31076]_  & \new_[31063]_ ;
  assign \new_[1301]_  = \new_[31052]_  & \new_[31039]_ ;
  assign \new_[1302]_  = \new_[31028]_  & \new_[31015]_ ;
  assign \new_[1303]_  = \new_[31004]_  & \new_[30991]_ ;
  assign \new_[1304]_  = \new_[30980]_  & \new_[30967]_ ;
  assign \new_[1305]_  = \new_[30956]_  & \new_[30943]_ ;
  assign \new_[1306]_  = \new_[30932]_  & \new_[30919]_ ;
  assign \new_[1307]_  = \new_[30908]_  & \new_[30895]_ ;
  assign \new_[1308]_  = \new_[30884]_  & \new_[30871]_ ;
  assign \new_[1309]_  = \new_[30860]_  & \new_[30847]_ ;
  assign \new_[1310]_  = \new_[30836]_  & \new_[30823]_ ;
  assign \new_[1311]_  = \new_[30812]_  & \new_[30799]_ ;
  assign \new_[1312]_  = \new_[30788]_  & \new_[30775]_ ;
  assign \new_[1313]_  = \new_[30764]_  & \new_[30751]_ ;
  assign \new_[1314]_  = \new_[30740]_  & \new_[30727]_ ;
  assign \new_[1315]_  = \new_[30716]_  & \new_[30703]_ ;
  assign \new_[1316]_  = \new_[30692]_  & \new_[30679]_ ;
  assign \new_[1317]_  = \new_[30668]_  & \new_[30655]_ ;
  assign \new_[1318]_  = \new_[30644]_  & \new_[30631]_ ;
  assign \new_[1319]_  = \new_[30620]_  & \new_[30609]_ ;
  assign \new_[1320]_  = \new_[30598]_  & \new_[30587]_ ;
  assign \new_[1321]_  = \new_[30576]_  & \new_[30565]_ ;
  assign \new_[1322]_  = \new_[30554]_  & \new_[30543]_ ;
  assign \new_[1323]_  = \new_[30532]_  & \new_[30521]_ ;
  assign \new_[1324]_  = \new_[30510]_  & \new_[30499]_ ;
  assign \new_[1325]_  = \new_[30488]_  & \new_[30477]_ ;
  assign \new_[1326]_  = \new_[30466]_  & \new_[30455]_ ;
  assign \new_[1327]_  = \new_[30444]_  & \new_[30433]_ ;
  assign \new_[1328]_  = \new_[30422]_  & \new_[30411]_ ;
  assign \new_[1329]_  = \new_[30400]_  & \new_[30389]_ ;
  assign \new_[1330]_  = \new_[30378]_  & \new_[30367]_ ;
  assign \new_[1331]_  = \new_[30356]_  & \new_[30345]_ ;
  assign \new_[1332]_  = \new_[30334]_  & \new_[30323]_ ;
  assign \new_[1333]_  = \new_[30312]_  & \new_[30301]_ ;
  assign \new_[1334]_  = \new_[30290]_  & \new_[30279]_ ;
  assign \new_[1335]_  = \new_[30268]_  & \new_[30257]_ ;
  assign \new_[1336]_  = \new_[30246]_  & \new_[30235]_ ;
  assign \new_[1337]_  = \new_[30224]_  & \new_[30213]_ ;
  assign \new_[1338]_  = \new_[30202]_  & \new_[30191]_ ;
  assign \new_[1339]_  = \new_[30180]_  & \new_[30169]_ ;
  assign \new_[1340]_  = \new_[30158]_  & \new_[30147]_ ;
  assign \new_[1341]_  = \new_[30136]_  & \new_[30125]_ ;
  assign \new_[1342]_  = \new_[30114]_  & \new_[30103]_ ;
  assign \new_[1343]_  = \new_[30092]_  & \new_[30081]_ ;
  assign \new_[1344]_  = \new_[30070]_  & \new_[30059]_ ;
  assign \new_[1345]_  = \new_[30048]_  & \new_[30037]_ ;
  assign \new_[1346]_  = \new_[30026]_  & \new_[30015]_ ;
  assign \new_[1347]_  = \new_[30004]_  & \new_[29993]_ ;
  assign \new_[1348]_  = \new_[29982]_  & \new_[29971]_ ;
  assign \new_[1349]_  = \new_[29960]_  & \new_[29949]_ ;
  assign \new_[1350]_  = \new_[29938]_  & \new_[29927]_ ;
  assign \new_[1351]_  = \new_[29916]_  & \new_[29905]_ ;
  assign \new_[1352]_  = \new_[29894]_  & \new_[29883]_ ;
  assign \new_[1353]_  = \new_[29872]_  & \new_[29861]_ ;
  assign \new_[1354]_  = \new_[29850]_  & \new_[29839]_ ;
  assign \new_[1355]_  = \new_[29828]_  & \new_[29817]_ ;
  assign \new_[1356]_  = \new_[29806]_  & \new_[29795]_ ;
  assign \new_[1357]_  = \new_[29784]_  & \new_[29773]_ ;
  assign \new_[1358]_  = \new_[29762]_  & \new_[29751]_ ;
  assign \new_[1359]_  = \new_[29740]_  & \new_[29729]_ ;
  assign \new_[1360]_  = \new_[29718]_  & \new_[29707]_ ;
  assign \new_[1361]_  = \new_[29696]_  & \new_[29685]_ ;
  assign \new_[1362]_  = \new_[29674]_  & \new_[29663]_ ;
  assign \new_[1363]_  = \new_[29652]_  & \new_[29641]_ ;
  assign \new_[1364]_  = \new_[29630]_  & \new_[29619]_ ;
  assign \new_[1365]_  = \new_[29608]_  & \new_[29597]_ ;
  assign \new_[1366]_  = \new_[29586]_  & \new_[29575]_ ;
  assign \new_[1367]_  = \new_[29564]_  & \new_[29553]_ ;
  assign \new_[1368]_  = \new_[29542]_  & \new_[29531]_ ;
  assign \new_[1369]_  = \new_[29520]_  & \new_[29509]_ ;
  assign \new_[1370]_  = \new_[29498]_  & \new_[29487]_ ;
  assign \new_[1371]_  = \new_[29476]_  & \new_[29465]_ ;
  assign \new_[1372]_  = \new_[29454]_  & \new_[29443]_ ;
  assign \new_[1373]_  = \new_[29432]_  & \new_[29421]_ ;
  assign \new_[1374]_  = \new_[29410]_  & \new_[29399]_ ;
  assign \new_[1375]_  = \new_[29388]_  & \new_[29377]_ ;
  assign \new_[1376]_  = \new_[29366]_  & \new_[29355]_ ;
  assign \new_[1377]_  = \new_[29344]_  & \new_[29333]_ ;
  assign \new_[1378]_  = \new_[29322]_  & \new_[29311]_ ;
  assign \new_[1379]_  = \new_[29300]_  & \new_[29289]_ ;
  assign \new_[1380]_  = \new_[29278]_  & \new_[29267]_ ;
  assign \new_[1381]_  = \new_[29256]_  & \new_[29245]_ ;
  assign \new_[1382]_  = \new_[29234]_  & \new_[29223]_ ;
  assign \new_[1383]_  = \new_[29212]_  & \new_[29201]_ ;
  assign \new_[1384]_  = \new_[29190]_  & \new_[29179]_ ;
  assign \new_[1385]_  = \new_[29168]_  & \new_[29157]_ ;
  assign \new_[1386]_  = \new_[29146]_  & \new_[29135]_ ;
  assign \new_[1387]_  = \new_[29124]_  & \new_[29113]_ ;
  assign \new_[1388]_  = \new_[29102]_  & \new_[29091]_ ;
  assign \new_[1389]_  = \new_[29080]_  & \new_[29069]_ ;
  assign \new_[1390]_  = \new_[29058]_  & \new_[29047]_ ;
  assign \new_[1391]_  = \new_[29036]_  & \new_[29025]_ ;
  assign \new_[1392]_  = \new_[29014]_  & \new_[29003]_ ;
  assign \new_[1393]_  = \new_[28992]_  & \new_[28981]_ ;
  assign \new_[1394]_  = \new_[28970]_  & \new_[28959]_ ;
  assign \new_[1395]_  = \new_[28948]_  & \new_[28937]_ ;
  assign \new_[1396]_  = \new_[28926]_  & \new_[28915]_ ;
  assign \new_[1397]_  = \new_[28904]_  & \new_[28893]_ ;
  assign \new_[1398]_  = \new_[28882]_  & \new_[28871]_ ;
  assign \new_[1399]_  = \new_[28860]_  & \new_[28849]_ ;
  assign \new_[1400]_  = \new_[28838]_  & \new_[28827]_ ;
  assign \new_[1401]_  = \new_[28816]_  & \new_[28805]_ ;
  assign \new_[1402]_  = \new_[28794]_  & \new_[28783]_ ;
  assign \new_[1403]_  = \new_[28772]_  & \new_[28761]_ ;
  assign \new_[1404]_  = \new_[28750]_  & \new_[28739]_ ;
  assign \new_[1405]_  = \new_[28728]_  & \new_[28717]_ ;
  assign \new_[1406]_  = \new_[28706]_  & \new_[28695]_ ;
  assign \new_[1407]_  = \new_[28684]_  & \new_[28673]_ ;
  assign \new_[1408]_  = \new_[28662]_  & \new_[28651]_ ;
  assign \new_[1409]_  = \new_[28640]_  & \new_[28629]_ ;
  assign \new_[1410]_  = \new_[28618]_  & \new_[28607]_ ;
  assign \new_[1411]_  = \new_[28596]_  & \new_[28585]_ ;
  assign \new_[1412]_  = \new_[28574]_  & \new_[28563]_ ;
  assign \new_[1413]_  = \new_[28552]_  & \new_[28541]_ ;
  assign \new_[1414]_  = \new_[28530]_  & \new_[28519]_ ;
  assign \new_[1415]_  = \new_[28508]_  & \new_[28497]_ ;
  assign \new_[1416]_  = \new_[28486]_  & \new_[28475]_ ;
  assign \new_[1417]_  = \new_[28464]_  & \new_[28453]_ ;
  assign \new_[1418]_  = \new_[28442]_  & \new_[28431]_ ;
  assign \new_[1419]_  = \new_[28420]_  & \new_[28409]_ ;
  assign \new_[1420]_  = \new_[28398]_  & \new_[28387]_ ;
  assign \new_[1421]_  = \new_[28376]_  & \new_[28365]_ ;
  assign \new_[1422]_  = \new_[28354]_  & \new_[28343]_ ;
  assign \new_[1423]_  = \new_[28332]_  & \new_[28321]_ ;
  assign \new_[1424]_  = \new_[28310]_  & \new_[28299]_ ;
  assign \new_[1425]_  = \new_[28288]_  & \new_[28277]_ ;
  assign \new_[1426]_  = \new_[28266]_  & \new_[28255]_ ;
  assign \new_[1427]_  = \new_[28244]_  & \new_[28233]_ ;
  assign \new_[1428]_  = \new_[28222]_  & \new_[28211]_ ;
  assign \new_[1429]_  = \new_[28200]_  & \new_[28189]_ ;
  assign \new_[1430]_  = \new_[28178]_  & \new_[28167]_ ;
  assign \new_[1431]_  = \new_[28156]_  & \new_[28145]_ ;
  assign \new_[1432]_  = \new_[28134]_  & \new_[28123]_ ;
  assign \new_[1433]_  = \new_[28112]_  & \new_[28101]_ ;
  assign \new_[1434]_  = \new_[28090]_  & \new_[28079]_ ;
  assign \new_[1435]_  = \new_[28068]_  & \new_[28057]_ ;
  assign \new_[1436]_  = \new_[28046]_  & \new_[28035]_ ;
  assign \new_[1437]_  = \new_[28024]_  & \new_[28013]_ ;
  assign \new_[1438]_  = \new_[28002]_  & \new_[27991]_ ;
  assign \new_[1439]_  = \new_[27980]_  & \new_[27969]_ ;
  assign \new_[1440]_  = \new_[27958]_  & \new_[27947]_ ;
  assign \new_[1441]_  = \new_[27936]_  & \new_[27925]_ ;
  assign \new_[1442]_  = \new_[27914]_  & \new_[27903]_ ;
  assign \new_[1443]_  = \new_[27892]_  & \new_[27881]_ ;
  assign \new_[1444]_  = \new_[27870]_  & \new_[27859]_ ;
  assign \new_[1445]_  = \new_[27848]_  & \new_[27837]_ ;
  assign \new_[1446]_  = \new_[27826]_  & \new_[27815]_ ;
  assign \new_[1447]_  = \new_[27804]_  & \new_[27793]_ ;
  assign \new_[1448]_  = \new_[27782]_  & \new_[27771]_ ;
  assign \new_[1449]_  = \new_[27760]_  & \new_[27749]_ ;
  assign \new_[1450]_  = \new_[27738]_  & \new_[27727]_ ;
  assign \new_[1451]_  = \new_[27716]_  & \new_[27705]_ ;
  assign \new_[1452]_  = \new_[27694]_  & \new_[27683]_ ;
  assign \new_[1453]_  = \new_[27672]_  & \new_[27661]_ ;
  assign \new_[1454]_  = \new_[27650]_  & \new_[27639]_ ;
  assign \new_[1455]_  = \new_[27628]_  & \new_[27617]_ ;
  assign \new_[1456]_  = \new_[27606]_  & \new_[27595]_ ;
  assign \new_[1457]_  = \new_[27584]_  & \new_[27573]_ ;
  assign \new_[1458]_  = \new_[27562]_  & \new_[27551]_ ;
  assign \new_[1459]_  = \new_[27540]_  & \new_[27529]_ ;
  assign \new_[1460]_  = \new_[27518]_  & \new_[27507]_ ;
  assign \new_[1461]_  = \new_[27496]_  & \new_[27485]_ ;
  assign \new_[1462]_  = \new_[27474]_  & \new_[27463]_ ;
  assign \new_[1463]_  = \new_[27452]_  & \new_[27441]_ ;
  assign \new_[1464]_  = \new_[27430]_  & \new_[27419]_ ;
  assign \new_[1465]_  = \new_[27408]_  & \new_[27397]_ ;
  assign \new_[1466]_  = \new_[27386]_  & \new_[27375]_ ;
  assign \new_[1467]_  = \new_[27364]_  & \new_[27353]_ ;
  assign \new_[1468]_  = \new_[27342]_  & \new_[27331]_ ;
  assign \new_[1469]_  = \new_[27320]_  & \new_[27309]_ ;
  assign \new_[1470]_  = \new_[27298]_  & \new_[27287]_ ;
  assign \new_[1471]_  = \new_[27276]_  & \new_[27265]_ ;
  assign \new_[1472]_  = \new_[27254]_  & \new_[27243]_ ;
  assign \new_[1473]_  = \new_[27232]_  & \new_[27221]_ ;
  assign \new_[1474]_  = \new_[27210]_  & \new_[27199]_ ;
  assign \new_[1475]_  = \new_[27188]_  & \new_[27177]_ ;
  assign \new_[1476]_  = \new_[27166]_  & \new_[27155]_ ;
  assign \new_[1477]_  = \new_[27144]_  & \new_[27133]_ ;
  assign \new_[1478]_  = \new_[27122]_  & \new_[27111]_ ;
  assign \new_[1479]_  = \new_[27100]_  & \new_[27089]_ ;
  assign \new_[1480]_  = \new_[27078]_  & \new_[27067]_ ;
  assign \new_[1481]_  = \new_[27056]_  & \new_[27045]_ ;
  assign \new_[1482]_  = \new_[27034]_  & \new_[27023]_ ;
  assign \new_[1483]_  = \new_[27012]_  & \new_[27001]_ ;
  assign \new_[1484]_  = \new_[26990]_  & \new_[26979]_ ;
  assign \new_[1485]_  = \new_[26968]_  & \new_[26957]_ ;
  assign \new_[1486]_  = \new_[26946]_  & \new_[26935]_ ;
  assign \new_[1487]_  = \new_[26924]_  & \new_[26913]_ ;
  assign \new_[1488]_  = \new_[26902]_  & \new_[26891]_ ;
  assign \new_[1489]_  = \new_[26880]_  & \new_[26869]_ ;
  assign \new_[1490]_  = \new_[26858]_  & \new_[26847]_ ;
  assign \new_[1491]_  = \new_[26836]_  & \new_[26825]_ ;
  assign \new_[1492]_  = \new_[26814]_  & \new_[26803]_ ;
  assign \new_[1493]_  = \new_[26792]_  & \new_[26781]_ ;
  assign \new_[1494]_  = \new_[26770]_  & \new_[26759]_ ;
  assign \new_[1495]_  = \new_[26748]_  & \new_[26737]_ ;
  assign \new_[1496]_  = \new_[26726]_  & \new_[26715]_ ;
  assign \new_[1497]_  = \new_[26704]_  & \new_[26693]_ ;
  assign \new_[1498]_  = \new_[26682]_  & \new_[26671]_ ;
  assign \new_[1499]_  = \new_[26660]_  & \new_[26649]_ ;
  assign \new_[1500]_  = \new_[26638]_  & \new_[26627]_ ;
  assign \new_[1501]_  = \new_[26616]_  & \new_[26605]_ ;
  assign \new_[1502]_  = \new_[26594]_  & \new_[26583]_ ;
  assign \new_[1503]_  = \new_[26572]_  & \new_[26561]_ ;
  assign \new_[1504]_  = \new_[26550]_  & \new_[26539]_ ;
  assign \new_[1505]_  = \new_[26528]_  & \new_[26517]_ ;
  assign \new_[1506]_  = \new_[26506]_  & \new_[26495]_ ;
  assign \new_[1507]_  = \new_[26484]_  & \new_[26473]_ ;
  assign \new_[1508]_  = \new_[26462]_  & \new_[26451]_ ;
  assign \new_[1509]_  = \new_[26440]_  & \new_[26429]_ ;
  assign \new_[1510]_  = \new_[26418]_  & \new_[26407]_ ;
  assign \new_[1511]_  = \new_[26396]_  & \new_[26385]_ ;
  assign \new_[1512]_  = \new_[26374]_  & \new_[26363]_ ;
  assign \new_[1513]_  = \new_[26352]_  & \new_[26341]_ ;
  assign \new_[1514]_  = \new_[26330]_  & \new_[26319]_ ;
  assign \new_[1515]_  = \new_[26308]_  & \new_[26297]_ ;
  assign \new_[1516]_  = \new_[26286]_  & \new_[26275]_ ;
  assign \new_[1517]_  = \new_[26264]_  & \new_[26253]_ ;
  assign \new_[1518]_  = \new_[26242]_  & \new_[26231]_ ;
  assign \new_[1519]_  = \new_[26220]_  & \new_[26209]_ ;
  assign \new_[1520]_  = \new_[26198]_  & \new_[26187]_ ;
  assign \new_[1521]_  = \new_[26176]_  & \new_[26165]_ ;
  assign \new_[1522]_  = \new_[26154]_  & \new_[26143]_ ;
  assign \new_[1523]_  = \new_[26132]_  & \new_[26121]_ ;
  assign \new_[1524]_  = \new_[26110]_  & \new_[26099]_ ;
  assign \new_[1525]_  = \new_[26088]_  & \new_[26077]_ ;
  assign \new_[1526]_  = \new_[26066]_  & \new_[26055]_ ;
  assign \new_[1527]_  = \new_[26044]_  & \new_[26033]_ ;
  assign \new_[1528]_  = \new_[26022]_  & \new_[26011]_ ;
  assign \new_[1529]_  = \new_[26000]_  & \new_[25989]_ ;
  assign \new_[1530]_  = \new_[25978]_  & \new_[25967]_ ;
  assign \new_[1531]_  = \new_[25956]_  & \new_[25945]_ ;
  assign \new_[1532]_  = \new_[25934]_  & \new_[25923]_ ;
  assign \new_[1533]_  = \new_[25912]_  & \new_[25901]_ ;
  assign \new_[1534]_  = \new_[25890]_  & \new_[25879]_ ;
  assign \new_[1535]_  = \new_[25868]_  & \new_[25857]_ ;
  assign \new_[1536]_  = \new_[25846]_  & \new_[25835]_ ;
  assign \new_[1537]_  = \new_[25824]_  & \new_[25813]_ ;
  assign \new_[1538]_  = \new_[25802]_  & \new_[25791]_ ;
  assign \new_[1539]_  = \new_[25780]_  & \new_[25769]_ ;
  assign \new_[1540]_  = \new_[25758]_  & \new_[25747]_ ;
  assign \new_[1541]_  = \new_[25736]_  & \new_[25725]_ ;
  assign \new_[1542]_  = \new_[25714]_  & \new_[25703]_ ;
  assign \new_[1543]_  = \new_[25692]_  & \new_[25681]_ ;
  assign \new_[1544]_  = \new_[25670]_  & \new_[25659]_ ;
  assign \new_[1545]_  = \new_[25648]_  & \new_[25637]_ ;
  assign \new_[1546]_  = \new_[25626]_  & \new_[25615]_ ;
  assign \new_[1547]_  = \new_[25604]_  & \new_[25593]_ ;
  assign \new_[1548]_  = \new_[25582]_  & \new_[25571]_ ;
  assign \new_[1549]_  = \new_[25560]_  & \new_[25549]_ ;
  assign \new_[1550]_  = \new_[25538]_  & \new_[25527]_ ;
  assign \new_[1551]_  = \new_[25516]_  & \new_[25505]_ ;
  assign \new_[1552]_  = \new_[25494]_  & \new_[25483]_ ;
  assign \new_[1553]_  = \new_[25472]_  & \new_[25461]_ ;
  assign \new_[1554]_  = \new_[25450]_  & \new_[25439]_ ;
  assign \new_[1555]_  = \new_[25428]_  & \new_[25417]_ ;
  assign \new_[1556]_  = \new_[25406]_  & \new_[25395]_ ;
  assign \new_[1557]_  = \new_[25384]_  & \new_[25373]_ ;
  assign \new_[1558]_  = \new_[25362]_  & \new_[25351]_ ;
  assign \new_[1559]_  = \new_[25340]_  & \new_[25329]_ ;
  assign \new_[1560]_  = \new_[25318]_  & \new_[25307]_ ;
  assign \new_[1561]_  = \new_[25296]_  & \new_[25285]_ ;
  assign \new_[1562]_  = \new_[25274]_  & \new_[25263]_ ;
  assign \new_[1563]_  = \new_[25252]_  & \new_[25241]_ ;
  assign \new_[1564]_  = \new_[25230]_  & \new_[25219]_ ;
  assign \new_[1565]_  = \new_[25208]_  & \new_[25197]_ ;
  assign \new_[1566]_  = \new_[25186]_  & \new_[25175]_ ;
  assign \new_[1567]_  = \new_[25164]_  & \new_[25153]_ ;
  assign \new_[1568]_  = \new_[25142]_  & \new_[25131]_ ;
  assign \new_[1569]_  = \new_[25120]_  & \new_[25109]_ ;
  assign \new_[1570]_  = \new_[25098]_  & \new_[25087]_ ;
  assign \new_[1571]_  = \new_[25076]_  & \new_[25065]_ ;
  assign \new_[1572]_  = \new_[25054]_  & \new_[25043]_ ;
  assign \new_[1573]_  = \new_[25032]_  & \new_[25021]_ ;
  assign \new_[1574]_  = \new_[25010]_  & \new_[24999]_ ;
  assign \new_[1575]_  = \new_[24988]_  & \new_[24977]_ ;
  assign \new_[1576]_  = \new_[24966]_  & \new_[24955]_ ;
  assign \new_[1577]_  = \new_[24944]_  & \new_[24933]_ ;
  assign \new_[1578]_  = \new_[24922]_  & \new_[24911]_ ;
  assign \new_[1579]_  = \new_[24900]_  & \new_[24889]_ ;
  assign \new_[1580]_  = \new_[24878]_  & \new_[24867]_ ;
  assign \new_[1581]_  = \new_[24856]_  & \new_[24845]_ ;
  assign \new_[1582]_  = \new_[24834]_  & \new_[24823]_ ;
  assign \new_[1583]_  = \new_[24812]_  & \new_[24801]_ ;
  assign \new_[1584]_  = \new_[24790]_  & \new_[24779]_ ;
  assign \new_[1585]_  = \new_[24768]_  & \new_[24757]_ ;
  assign \new_[1586]_  = \new_[24746]_  & \new_[24735]_ ;
  assign \new_[1587]_  = \new_[24724]_  & \new_[24713]_ ;
  assign \new_[1588]_  = \new_[24702]_  & \new_[24691]_ ;
  assign \new_[1589]_  = \new_[24680]_  & \new_[24669]_ ;
  assign \new_[1590]_  = \new_[24658]_  & \new_[24647]_ ;
  assign \new_[1591]_  = \new_[24636]_  & \new_[24625]_ ;
  assign \new_[1592]_  = \new_[24614]_  & \new_[24603]_ ;
  assign \new_[1593]_  = \new_[24592]_  & \new_[24581]_ ;
  assign \new_[1594]_  = \new_[24570]_  & \new_[24559]_ ;
  assign \new_[1595]_  = \new_[24548]_  & \new_[24537]_ ;
  assign \new_[1596]_  = \new_[24526]_  & \new_[24515]_ ;
  assign \new_[1597]_  = \new_[24504]_  & \new_[24493]_ ;
  assign \new_[1598]_  = \new_[24482]_  & \new_[24471]_ ;
  assign \new_[1599]_  = \new_[24460]_  & \new_[24449]_ ;
  assign \new_[1600]_  = \new_[24440]_  & \new_[24429]_ ;
  assign \new_[1601]_  = \new_[24420]_  & \new_[24409]_ ;
  assign \new_[1602]_  = \new_[24400]_  & \new_[24389]_ ;
  assign \new_[1603]_  = \new_[24380]_  & \new_[24369]_ ;
  assign \new_[1604]_  = \new_[24360]_  & \new_[24349]_ ;
  assign \new_[1605]_  = \new_[24340]_  & \new_[24329]_ ;
  assign \new_[1606]_  = \new_[24320]_  & \new_[24309]_ ;
  assign \new_[1607]_  = \new_[24300]_  & \new_[24289]_ ;
  assign \new_[1608]_  = \new_[24280]_  & \new_[24269]_ ;
  assign \new_[1609]_  = \new_[24260]_  & \new_[24249]_ ;
  assign \new_[1610]_  = \new_[24240]_  & \new_[24229]_ ;
  assign \new_[1611]_  = \new_[24220]_  & \new_[24209]_ ;
  assign \new_[1612]_  = \new_[24200]_  & \new_[24189]_ ;
  assign \new_[1613]_  = \new_[24180]_  & \new_[24169]_ ;
  assign \new_[1614]_  = \new_[24160]_  & \new_[24149]_ ;
  assign \new_[1615]_  = \new_[24140]_  & \new_[24129]_ ;
  assign \new_[1616]_  = \new_[24120]_  & \new_[24109]_ ;
  assign \new_[1617]_  = \new_[24100]_  & \new_[24089]_ ;
  assign \new_[1618]_  = \new_[24080]_  & \new_[24069]_ ;
  assign \new_[1619]_  = \new_[24060]_  & \new_[24049]_ ;
  assign \new_[1620]_  = \new_[24040]_  & \new_[24029]_ ;
  assign \new_[1621]_  = \new_[24020]_  & \new_[24009]_ ;
  assign \new_[1622]_  = \new_[24000]_  & \new_[23989]_ ;
  assign \new_[1623]_  = \new_[23980]_  & \new_[23969]_ ;
  assign \new_[1624]_  = \new_[23960]_  & \new_[23949]_ ;
  assign \new_[1625]_  = \new_[23940]_  & \new_[23929]_ ;
  assign \new_[1626]_  = \new_[23920]_  & \new_[23909]_ ;
  assign \new_[1627]_  = \new_[23900]_  & \new_[23889]_ ;
  assign \new_[1628]_  = \new_[23880]_  & \new_[23869]_ ;
  assign \new_[1629]_  = \new_[23860]_  & \new_[23849]_ ;
  assign \new_[1630]_  = \new_[23840]_  & \new_[23829]_ ;
  assign \new_[1631]_  = \new_[23820]_  & \new_[23809]_ ;
  assign \new_[1632]_  = \new_[23800]_  & \new_[23789]_ ;
  assign \new_[1633]_  = \new_[23780]_  & \new_[23769]_ ;
  assign \new_[1634]_  = \new_[23760]_  & \new_[23749]_ ;
  assign \new_[1635]_  = \new_[23740]_  & \new_[23729]_ ;
  assign \new_[1636]_  = \new_[23720]_  & \new_[23709]_ ;
  assign \new_[1637]_  = \new_[23700]_  & \new_[23689]_ ;
  assign \new_[1638]_  = \new_[23680]_  & \new_[23669]_ ;
  assign \new_[1639]_  = \new_[23660]_  & \new_[23649]_ ;
  assign \new_[1640]_  = \new_[23640]_  & \new_[23629]_ ;
  assign \new_[1641]_  = \new_[23620]_  & \new_[23609]_ ;
  assign \new_[1642]_  = \new_[23600]_  & \new_[23589]_ ;
  assign \new_[1643]_  = \new_[23580]_  & \new_[23569]_ ;
  assign \new_[1644]_  = \new_[23560]_  & \new_[23549]_ ;
  assign \new_[1645]_  = \new_[23540]_  & \new_[23529]_ ;
  assign \new_[1646]_  = \new_[23520]_  & \new_[23509]_ ;
  assign \new_[1647]_  = \new_[23500]_  & \new_[23489]_ ;
  assign \new_[1648]_  = \new_[23480]_  & \new_[23469]_ ;
  assign \new_[1649]_  = \new_[23460]_  & \new_[23449]_ ;
  assign \new_[1650]_  = \new_[23440]_  & \new_[23429]_ ;
  assign \new_[1651]_  = \new_[23420]_  & \new_[23409]_ ;
  assign \new_[1652]_  = \new_[23400]_  & \new_[23389]_ ;
  assign \new_[1653]_  = \new_[23380]_  & \new_[23369]_ ;
  assign \new_[1654]_  = \new_[23360]_  & \new_[23349]_ ;
  assign \new_[1655]_  = \new_[23340]_  & \new_[23329]_ ;
  assign \new_[1656]_  = \new_[23320]_  & \new_[23309]_ ;
  assign \new_[1657]_  = \new_[23300]_  & \new_[23289]_ ;
  assign \new_[1658]_  = \new_[23280]_  & \new_[23269]_ ;
  assign \new_[1659]_  = \new_[23260]_  & \new_[23249]_ ;
  assign \new_[1660]_  = \new_[23240]_  & \new_[23229]_ ;
  assign \new_[1661]_  = \new_[23220]_  & \new_[23209]_ ;
  assign \new_[1662]_  = \new_[23200]_  & \new_[23189]_ ;
  assign \new_[1663]_  = \new_[23180]_  & \new_[23169]_ ;
  assign \new_[1664]_  = \new_[23160]_  & \new_[23149]_ ;
  assign \new_[1665]_  = \new_[23140]_  & \new_[23129]_ ;
  assign \new_[1666]_  = \new_[23120]_  & \new_[23109]_ ;
  assign \new_[1667]_  = \new_[23100]_  & \new_[23089]_ ;
  assign \new_[1668]_  = \new_[23080]_  & \new_[23069]_ ;
  assign \new_[1669]_  = \new_[23060]_  & \new_[23049]_ ;
  assign \new_[1670]_  = \new_[23040]_  & \new_[23029]_ ;
  assign \new_[1671]_  = \new_[23020]_  & \new_[23009]_ ;
  assign \new_[1672]_  = \new_[23000]_  & \new_[22989]_ ;
  assign \new_[1673]_  = \new_[22980]_  & \new_[22969]_ ;
  assign \new_[1674]_  = \new_[22960]_  & \new_[22949]_ ;
  assign \new_[1675]_  = \new_[22940]_  & \new_[22929]_ ;
  assign \new_[1676]_  = \new_[22920]_  & \new_[22909]_ ;
  assign \new_[1677]_  = \new_[22900]_  & \new_[22889]_ ;
  assign \new_[1678]_  = \new_[22880]_  & \new_[22869]_ ;
  assign \new_[1679]_  = \new_[22860]_  & \new_[22849]_ ;
  assign \new_[1680]_  = \new_[22840]_  & \new_[22829]_ ;
  assign \new_[1681]_  = \new_[22820]_  & \new_[22809]_ ;
  assign \new_[1682]_  = \new_[22800]_  & \new_[22789]_ ;
  assign \new_[1683]_  = \new_[22780]_  & \new_[22769]_ ;
  assign \new_[1684]_  = \new_[22760]_  & \new_[22749]_ ;
  assign \new_[1685]_  = \new_[22740]_  & \new_[22729]_ ;
  assign \new_[1686]_  = \new_[22720]_  & \new_[22709]_ ;
  assign \new_[1687]_  = \new_[22700]_  & \new_[22689]_ ;
  assign \new_[1688]_  = \new_[22680]_  & \new_[22669]_ ;
  assign \new_[1689]_  = \new_[22660]_  & \new_[22649]_ ;
  assign \new_[1690]_  = \new_[22640]_  & \new_[22629]_ ;
  assign \new_[1691]_  = \new_[22620]_  & \new_[22609]_ ;
  assign \new_[1692]_  = \new_[22600]_  & \new_[22589]_ ;
  assign \new_[1693]_  = \new_[22580]_  & \new_[22569]_ ;
  assign \new_[1694]_  = \new_[22560]_  & \new_[22549]_ ;
  assign \new_[1695]_  = \new_[22540]_  & \new_[22529]_ ;
  assign \new_[1696]_  = \new_[22520]_  & \new_[22509]_ ;
  assign \new_[1697]_  = \new_[22500]_  & \new_[22489]_ ;
  assign \new_[1698]_  = \new_[22480]_  & \new_[22469]_ ;
  assign \new_[1699]_  = \new_[22460]_  & \new_[22449]_ ;
  assign \new_[1700]_  = \new_[22440]_  & \new_[22429]_ ;
  assign \new_[1701]_  = \new_[22420]_  & \new_[22409]_ ;
  assign \new_[1702]_  = \new_[22400]_  & \new_[22389]_ ;
  assign \new_[1703]_  = \new_[22380]_  & \new_[22369]_ ;
  assign \new_[1704]_  = \new_[22360]_  & \new_[22349]_ ;
  assign \new_[1705]_  = \new_[22340]_  & \new_[22329]_ ;
  assign \new_[1706]_  = \new_[22320]_  & \new_[22309]_ ;
  assign \new_[1707]_  = \new_[22300]_  & \new_[22289]_ ;
  assign \new_[1708]_  = \new_[22280]_  & \new_[22269]_ ;
  assign \new_[1709]_  = \new_[22260]_  & \new_[22249]_ ;
  assign \new_[1710]_  = \new_[22240]_  & \new_[22229]_ ;
  assign \new_[1711]_  = \new_[22220]_  & \new_[22209]_ ;
  assign \new_[1712]_  = \new_[22200]_  & \new_[22189]_ ;
  assign \new_[1713]_  = \new_[22180]_  & \new_[22169]_ ;
  assign \new_[1714]_  = \new_[22160]_  & \new_[22149]_ ;
  assign \new_[1715]_  = \new_[22140]_  & \new_[22129]_ ;
  assign \new_[1716]_  = \new_[22120]_  & \new_[22109]_ ;
  assign \new_[1717]_  = \new_[22100]_  & \new_[22089]_ ;
  assign \new_[1718]_  = \new_[22080]_  & \new_[22069]_ ;
  assign \new_[1719]_  = \new_[22060]_  & \new_[22049]_ ;
  assign \new_[1720]_  = \new_[22040]_  & \new_[22029]_ ;
  assign \new_[1721]_  = \new_[22020]_  & \new_[22009]_ ;
  assign \new_[1722]_  = \new_[22000]_  & \new_[21989]_ ;
  assign \new_[1723]_  = \new_[21980]_  & \new_[21969]_ ;
  assign \new_[1724]_  = \new_[21960]_  & \new_[21949]_ ;
  assign \new_[1725]_  = \new_[21940]_  & \new_[21929]_ ;
  assign \new_[1726]_  = \new_[21920]_  & \new_[21909]_ ;
  assign \new_[1727]_  = \new_[21900]_  & \new_[21889]_ ;
  assign \new_[1728]_  = \new_[21880]_  & \new_[21869]_ ;
  assign \new_[1729]_  = \new_[21860]_  & \new_[21849]_ ;
  assign \new_[1730]_  = \new_[21840]_  & \new_[21829]_ ;
  assign \new_[1731]_  = \new_[21820]_  & \new_[21809]_ ;
  assign \new_[1732]_  = \new_[21800]_  & \new_[21789]_ ;
  assign \new_[1733]_  = \new_[21780]_  & \new_[21769]_ ;
  assign \new_[1734]_  = \new_[21760]_  & \new_[21749]_ ;
  assign \new_[1735]_  = \new_[21740]_  & \new_[21729]_ ;
  assign \new_[1736]_  = \new_[21720]_  & \new_[21709]_ ;
  assign \new_[1737]_  = \new_[21700]_  & \new_[21689]_ ;
  assign \new_[1738]_  = \new_[21680]_  & \new_[21669]_ ;
  assign \new_[1739]_  = \new_[21660]_  & \new_[21649]_ ;
  assign \new_[1740]_  = \new_[21640]_  & \new_[21629]_ ;
  assign \new_[1741]_  = \new_[21620]_  & \new_[21609]_ ;
  assign \new_[1742]_  = \new_[21600]_  & \new_[21589]_ ;
  assign \new_[1743]_  = \new_[21580]_  & \new_[21569]_ ;
  assign \new_[1744]_  = \new_[21560]_  & \new_[21549]_ ;
  assign \new_[1745]_  = \new_[21540]_  & \new_[21529]_ ;
  assign \new_[1746]_  = \new_[21520]_  & \new_[21509]_ ;
  assign \new_[1747]_  = \new_[21500]_  & \new_[21489]_ ;
  assign \new_[1748]_  = \new_[21480]_  & \new_[21469]_ ;
  assign \new_[1749]_  = \new_[21460]_  & \new_[21449]_ ;
  assign \new_[1750]_  = \new_[21440]_  & \new_[21429]_ ;
  assign \new_[1751]_  = \new_[21420]_  & \new_[21409]_ ;
  assign \new_[1752]_  = \new_[21400]_  & \new_[21389]_ ;
  assign \new_[1753]_  = \new_[21380]_  & \new_[21369]_ ;
  assign \new_[1754]_  = \new_[21360]_  & \new_[21349]_ ;
  assign \new_[1755]_  = \new_[21340]_  & \new_[21329]_ ;
  assign \new_[1756]_  = \new_[21320]_  & \new_[21309]_ ;
  assign \new_[1757]_  = \new_[21300]_  & \new_[21289]_ ;
  assign \new_[1758]_  = \new_[21280]_  & \new_[21269]_ ;
  assign \new_[1759]_  = \new_[21260]_  & \new_[21249]_ ;
  assign \new_[1760]_  = \new_[21240]_  & \new_[21229]_ ;
  assign \new_[1761]_  = \new_[21220]_  & \new_[21209]_ ;
  assign \new_[1762]_  = \new_[21200]_  & \new_[21189]_ ;
  assign \new_[1763]_  = \new_[21180]_  & \new_[21169]_ ;
  assign \new_[1764]_  = \new_[21160]_  & \new_[21149]_ ;
  assign \new_[1765]_  = \new_[21140]_  & \new_[21129]_ ;
  assign \new_[1766]_  = \new_[21120]_  & \new_[21109]_ ;
  assign \new_[1767]_  = \new_[21100]_  & \new_[21089]_ ;
  assign \new_[1768]_  = \new_[21080]_  & \new_[21069]_ ;
  assign \new_[1769]_  = \new_[21060]_  & \new_[21049]_ ;
  assign \new_[1770]_  = \new_[21040]_  & \new_[21029]_ ;
  assign \new_[1771]_  = \new_[21020]_  & \new_[21009]_ ;
  assign \new_[1772]_  = \new_[21000]_  & \new_[20989]_ ;
  assign \new_[1773]_  = \new_[20980]_  & \new_[20969]_ ;
  assign \new_[1774]_  = \new_[20960]_  & \new_[20949]_ ;
  assign \new_[1775]_  = \new_[20940]_  & \new_[20929]_ ;
  assign \new_[1776]_  = \new_[20920]_  & \new_[20909]_ ;
  assign \new_[1777]_  = \new_[20900]_  & \new_[20889]_ ;
  assign \new_[1778]_  = \new_[20880]_  & \new_[20869]_ ;
  assign \new_[1779]_  = \new_[20860]_  & \new_[20849]_ ;
  assign \new_[1780]_  = \new_[20840]_  & \new_[20829]_ ;
  assign \new_[1781]_  = \new_[20820]_  & \new_[20809]_ ;
  assign \new_[1782]_  = \new_[20800]_  & \new_[20789]_ ;
  assign \new_[1783]_  = \new_[20780]_  & \new_[20769]_ ;
  assign \new_[1784]_  = \new_[20760]_  & \new_[20749]_ ;
  assign \new_[1785]_  = \new_[20740]_  & \new_[20729]_ ;
  assign \new_[1786]_  = \new_[20720]_  & \new_[20709]_ ;
  assign \new_[1787]_  = \new_[20700]_  & \new_[20689]_ ;
  assign \new_[1788]_  = \new_[20680]_  & \new_[20669]_ ;
  assign \new_[1789]_  = \new_[20660]_  & \new_[20649]_ ;
  assign \new_[1790]_  = \new_[20640]_  & \new_[20629]_ ;
  assign \new_[1791]_  = \new_[20620]_  & \new_[20609]_ ;
  assign \new_[1792]_  = \new_[20600]_  & \new_[20589]_ ;
  assign \new_[1793]_  = \new_[20580]_  & \new_[20569]_ ;
  assign \new_[1794]_  = \new_[20560]_  & \new_[20549]_ ;
  assign \new_[1795]_  = \new_[20540]_  & \new_[20529]_ ;
  assign \new_[1796]_  = \new_[20520]_  & \new_[20509]_ ;
  assign \new_[1797]_  = \new_[20500]_  & \new_[20489]_ ;
  assign \new_[1798]_  = \new_[20480]_  & \new_[20469]_ ;
  assign \new_[1799]_  = \new_[20460]_  & \new_[20449]_ ;
  assign \new_[1800]_  = \new_[20440]_  & \new_[20429]_ ;
  assign \new_[1801]_  = \new_[20420]_  & \new_[20409]_ ;
  assign \new_[1802]_  = \new_[20400]_  & \new_[20389]_ ;
  assign \new_[1803]_  = \new_[20380]_  & \new_[20369]_ ;
  assign \new_[1804]_  = \new_[20360]_  & \new_[20349]_ ;
  assign \new_[1805]_  = \new_[20340]_  & \new_[20329]_ ;
  assign \new_[1806]_  = \new_[20320]_  & \new_[20309]_ ;
  assign \new_[1807]_  = \new_[20300]_  & \new_[20289]_ ;
  assign \new_[1808]_  = \new_[20280]_  & \new_[20269]_ ;
  assign \new_[1809]_  = \new_[20260]_  & \new_[20249]_ ;
  assign \new_[1810]_  = \new_[20240]_  & \new_[20229]_ ;
  assign \new_[1811]_  = \new_[20220]_  & \new_[20209]_ ;
  assign \new_[1812]_  = \new_[20200]_  & \new_[20189]_ ;
  assign \new_[1813]_  = \new_[20180]_  & \new_[20169]_ ;
  assign \new_[1814]_  = \new_[20160]_  & \new_[20149]_ ;
  assign \new_[1815]_  = \new_[20140]_  & \new_[20129]_ ;
  assign \new_[1816]_  = \new_[20120]_  & \new_[20109]_ ;
  assign \new_[1817]_  = \new_[20100]_  & \new_[20089]_ ;
  assign \new_[1818]_  = \new_[20080]_  & \new_[20069]_ ;
  assign \new_[1819]_  = \new_[20060]_  & \new_[20049]_ ;
  assign \new_[1820]_  = \new_[20040]_  & \new_[20029]_ ;
  assign \new_[1821]_  = \new_[20020]_  & \new_[20009]_ ;
  assign \new_[1822]_  = \new_[20000]_  & \new_[19989]_ ;
  assign \new_[1823]_  = \new_[19980]_  & \new_[19969]_ ;
  assign \new_[1824]_  = \new_[19960]_  & \new_[19949]_ ;
  assign \new_[1825]_  = \new_[19940]_  & \new_[19929]_ ;
  assign \new_[1826]_  = \new_[19920]_  & \new_[19909]_ ;
  assign \new_[1827]_  = \new_[19900]_  & \new_[19889]_ ;
  assign \new_[1828]_  = \new_[19880]_  & \new_[19869]_ ;
  assign \new_[1829]_  = \new_[19860]_  & \new_[19849]_ ;
  assign \new_[1830]_  = \new_[19840]_  & \new_[19829]_ ;
  assign \new_[1831]_  = \new_[19820]_  & \new_[19809]_ ;
  assign \new_[1832]_  = \new_[19800]_  & \new_[19789]_ ;
  assign \new_[1833]_  = \new_[19780]_  & \new_[19769]_ ;
  assign \new_[1834]_  = \new_[19760]_  & \new_[19749]_ ;
  assign \new_[1835]_  = \new_[19740]_  & \new_[19729]_ ;
  assign \new_[1836]_  = \new_[19720]_  & \new_[19709]_ ;
  assign \new_[1837]_  = \new_[19700]_  & \new_[19689]_ ;
  assign \new_[1838]_  = \new_[19680]_  & \new_[19669]_ ;
  assign \new_[1839]_  = \new_[19660]_  & \new_[19649]_ ;
  assign \new_[1840]_  = \new_[19640]_  & \new_[19629]_ ;
  assign \new_[1841]_  = \new_[19620]_  & \new_[19609]_ ;
  assign \new_[1842]_  = \new_[19600]_  & \new_[19589]_ ;
  assign \new_[1843]_  = \new_[19580]_  & \new_[19569]_ ;
  assign \new_[1844]_  = \new_[19560]_  & \new_[19549]_ ;
  assign \new_[1845]_  = \new_[19540]_  & \new_[19529]_ ;
  assign \new_[1846]_  = \new_[19520]_  & \new_[19509]_ ;
  assign \new_[1847]_  = \new_[19500]_  & \new_[19489]_ ;
  assign \new_[1848]_  = \new_[19480]_  & \new_[19469]_ ;
  assign \new_[1849]_  = \new_[19460]_  & \new_[19449]_ ;
  assign \new_[1850]_  = \new_[19440]_  & \new_[19429]_ ;
  assign \new_[1851]_  = \new_[19420]_  & \new_[19409]_ ;
  assign \new_[1852]_  = \new_[19400]_  & \new_[19389]_ ;
  assign \new_[1853]_  = \new_[19380]_  & \new_[19369]_ ;
  assign \new_[1854]_  = \new_[19360]_  & \new_[19349]_ ;
  assign \new_[1855]_  = \new_[19340]_  & \new_[19329]_ ;
  assign \new_[1856]_  = \new_[19320]_  & \new_[19309]_ ;
  assign \new_[1857]_  = \new_[19300]_  & \new_[19289]_ ;
  assign \new_[1858]_  = \new_[19280]_  & \new_[19269]_ ;
  assign \new_[1859]_  = \new_[19260]_  & \new_[19249]_ ;
  assign \new_[1860]_  = \new_[19240]_  & \new_[19229]_ ;
  assign \new_[1861]_  = \new_[19220]_  & \new_[19209]_ ;
  assign \new_[1862]_  = \new_[19200]_  & \new_[19189]_ ;
  assign \new_[1863]_  = \new_[19180]_  & \new_[19169]_ ;
  assign \new_[1864]_  = \new_[19160]_  & \new_[19149]_ ;
  assign \new_[1865]_  = \new_[19140]_  & \new_[19129]_ ;
  assign \new_[1866]_  = \new_[19120]_  & \new_[19109]_ ;
  assign \new_[1867]_  = \new_[19100]_  & \new_[19089]_ ;
  assign \new_[1868]_  = \new_[19080]_  & \new_[19069]_ ;
  assign \new_[1869]_  = \new_[19060]_  & \new_[19049]_ ;
  assign \new_[1870]_  = \new_[19040]_  & \new_[19029]_ ;
  assign \new_[1871]_  = \new_[19020]_  & \new_[19009]_ ;
  assign \new_[1872]_  = \new_[19000]_  & \new_[18989]_ ;
  assign \new_[1873]_  = \new_[18980]_  & \new_[18969]_ ;
  assign \new_[1874]_  = \new_[18960]_  & \new_[18949]_ ;
  assign \new_[1875]_  = \new_[18940]_  & \new_[18929]_ ;
  assign \new_[1876]_  = \new_[18920]_  & \new_[18909]_ ;
  assign \new_[1877]_  = \new_[18900]_  & \new_[18889]_ ;
  assign \new_[1878]_  = \new_[18880]_  & \new_[18869]_ ;
  assign \new_[1879]_  = \new_[18860]_  & \new_[18849]_ ;
  assign \new_[1880]_  = \new_[18840]_  & \new_[18829]_ ;
  assign \new_[1881]_  = \new_[18820]_  & \new_[18809]_ ;
  assign \new_[1882]_  = \new_[18800]_  & \new_[18789]_ ;
  assign \new_[1883]_  = \new_[18780]_  & \new_[18769]_ ;
  assign \new_[1884]_  = \new_[18760]_  & \new_[18749]_ ;
  assign \new_[1885]_  = \new_[18740]_  & \new_[18729]_ ;
  assign \new_[1886]_  = \new_[18720]_  & \new_[18709]_ ;
  assign \new_[1887]_  = \new_[18700]_  & \new_[18689]_ ;
  assign \new_[1888]_  = \new_[18680]_  & \new_[18669]_ ;
  assign \new_[1889]_  = \new_[18660]_  & \new_[18649]_ ;
  assign \new_[1890]_  = \new_[18640]_  & \new_[18629]_ ;
  assign \new_[1891]_  = \new_[18620]_  & \new_[18609]_ ;
  assign \new_[1892]_  = \new_[18600]_  & \new_[18589]_ ;
  assign \new_[1893]_  = \new_[18580]_  & \new_[18569]_ ;
  assign \new_[1894]_  = \new_[18560]_  & \new_[18549]_ ;
  assign \new_[1895]_  = \new_[18540]_  & \new_[18529]_ ;
  assign \new_[1896]_  = \new_[18520]_  & \new_[18509]_ ;
  assign \new_[1897]_  = \new_[18500]_  & \new_[18489]_ ;
  assign \new_[1898]_  = \new_[18480]_  & \new_[18469]_ ;
  assign \new_[1899]_  = \new_[18460]_  & \new_[18449]_ ;
  assign \new_[1900]_  = \new_[18440]_  & \new_[18429]_ ;
  assign \new_[1901]_  = \new_[18420]_  & \new_[18409]_ ;
  assign \new_[1902]_  = \new_[18400]_  & \new_[18389]_ ;
  assign \new_[1903]_  = \new_[18380]_  & \new_[18369]_ ;
  assign \new_[1904]_  = \new_[18360]_  & \new_[18349]_ ;
  assign \new_[1905]_  = \new_[18340]_  & \new_[18329]_ ;
  assign \new_[1906]_  = \new_[18320]_  & \new_[18309]_ ;
  assign \new_[1907]_  = \new_[18300]_  & \new_[18289]_ ;
  assign \new_[1908]_  = \new_[18280]_  & \new_[18269]_ ;
  assign \new_[1909]_  = \new_[18260]_  & \new_[18249]_ ;
  assign \new_[1910]_  = \new_[18240]_  & \new_[18229]_ ;
  assign \new_[1911]_  = \new_[18220]_  & \new_[18209]_ ;
  assign \new_[1912]_  = \new_[18200]_  & \new_[18189]_ ;
  assign \new_[1913]_  = \new_[18180]_  & \new_[18169]_ ;
  assign \new_[1914]_  = \new_[18160]_  & \new_[18149]_ ;
  assign \new_[1915]_  = \new_[18140]_  & \new_[18129]_ ;
  assign \new_[1916]_  = \new_[18120]_  & \new_[18109]_ ;
  assign \new_[1917]_  = \new_[18100]_  & \new_[18089]_ ;
  assign \new_[1918]_  = \new_[18080]_  & \new_[18069]_ ;
  assign \new_[1919]_  = \new_[18060]_  & \new_[18051]_ ;
  assign \new_[1920]_  = \new_[18042]_  & \new_[18033]_ ;
  assign \new_[1921]_  = \new_[18024]_  & \new_[18015]_ ;
  assign \new_[1922]_  = \new_[18006]_  & \new_[17997]_ ;
  assign \new_[1923]_  = \new_[17988]_  & \new_[17979]_ ;
  assign \new_[1924]_  = \new_[17970]_  & \new_[17961]_ ;
  assign \new_[1925]_  = \new_[17952]_  & \new_[17943]_ ;
  assign \new_[1926]_  = \new_[17934]_  & \new_[17925]_ ;
  assign \new_[1927]_  = \new_[17916]_  & \new_[17907]_ ;
  assign \new_[1928]_  = \new_[17898]_  & \new_[17889]_ ;
  assign \new_[1929]_  = \new_[17880]_  & \new_[17871]_ ;
  assign \new_[1930]_  = \new_[17862]_  & \new_[17853]_ ;
  assign \new_[1931]_  = \new_[17844]_  & \new_[17835]_ ;
  assign \new_[1932]_  = \new_[17826]_  & \new_[17817]_ ;
  assign \new_[1933]_  = \new_[17808]_  & \new_[17799]_ ;
  assign \new_[1934]_  = \new_[17790]_  & \new_[17781]_ ;
  assign \new_[1935]_  = \new_[17772]_  & \new_[17763]_ ;
  assign \new_[1936]_  = \new_[17754]_  & \new_[17745]_ ;
  assign \new_[1937]_  = \new_[17736]_  & \new_[17727]_ ;
  assign \new_[1938]_  = \new_[17718]_  & \new_[17709]_ ;
  assign \new_[1939]_  = \new_[17700]_  & \new_[17691]_ ;
  assign \new_[1940]_  = \new_[17682]_  & \new_[17673]_ ;
  assign \new_[1941]_  = \new_[17664]_  & \new_[17655]_ ;
  assign \new_[1942]_  = \new_[17646]_  & \new_[17637]_ ;
  assign \new_[1943]_  = \new_[17628]_  & \new_[17619]_ ;
  assign \new_[1944]_  = \new_[17610]_  & \new_[17601]_ ;
  assign \new_[1945]_  = \new_[17592]_  & \new_[17583]_ ;
  assign \new_[1946]_  = \new_[17574]_  & \new_[17565]_ ;
  assign \new_[1947]_  = \new_[17556]_  & \new_[17547]_ ;
  assign \new_[1948]_  = \new_[17538]_  & \new_[17529]_ ;
  assign \new_[1949]_  = \new_[17520]_  & \new_[17511]_ ;
  assign \new_[1950]_  = \new_[17502]_  & \new_[17493]_ ;
  assign \new_[1951]_  = \new_[17484]_  & \new_[17475]_ ;
  assign \new_[1952]_  = \new_[17466]_  & \new_[17457]_ ;
  assign \new_[1953]_  = \new_[17448]_  & \new_[17439]_ ;
  assign \new_[1954]_  = \new_[17430]_  & \new_[17421]_ ;
  assign \new_[1955]_  = \new_[17412]_  & \new_[17403]_ ;
  assign \new_[1956]_  = \new_[17394]_  & \new_[17385]_ ;
  assign \new_[1957]_  = \new_[17376]_  & \new_[17367]_ ;
  assign \new_[1958]_  = \new_[17358]_  & \new_[17349]_ ;
  assign \new_[1959]_  = \new_[17340]_  & \new_[17331]_ ;
  assign \new_[1960]_  = \new_[17322]_  & \new_[17313]_ ;
  assign \new_[1961]_  = \new_[17304]_  & \new_[17295]_ ;
  assign \new_[1962]_  = \new_[17286]_  & \new_[17277]_ ;
  assign \new_[1963]_  = \new_[17268]_  & \new_[17259]_ ;
  assign \new_[1964]_  = \new_[17250]_  & \new_[17241]_ ;
  assign \new_[1965]_  = \new_[17232]_  & \new_[17223]_ ;
  assign \new_[1966]_  = \new_[17214]_  & \new_[17205]_ ;
  assign \new_[1967]_  = \new_[17196]_  & \new_[17187]_ ;
  assign \new_[1968]_  = \new_[17178]_  & \new_[17169]_ ;
  assign \new_[1969]_  = \new_[17160]_  & \new_[17151]_ ;
  assign \new_[1970]_  = \new_[17142]_  & \new_[17133]_ ;
  assign \new_[1971]_  = \new_[17124]_  & \new_[17115]_ ;
  assign \new_[1972]_  = \new_[17106]_  & \new_[17097]_ ;
  assign \new_[1973]_  = \new_[17088]_  & \new_[17079]_ ;
  assign \new_[1974]_  = \new_[17070]_  & \new_[17061]_ ;
  assign \new_[1975]_  = \new_[17052]_  & \new_[17043]_ ;
  assign \new_[1976]_  = \new_[17034]_  & \new_[17025]_ ;
  assign \new_[1977]_  = \new_[17016]_  & \new_[17007]_ ;
  assign \new_[1978]_  = \new_[16998]_  & \new_[16989]_ ;
  assign \new_[1979]_  = \new_[16980]_  & \new_[16971]_ ;
  assign \new_[1980]_  = \new_[16962]_  & \new_[16953]_ ;
  assign \new_[1981]_  = \new_[16944]_  & \new_[16935]_ ;
  assign \new_[1982]_  = \new_[16926]_  & \new_[16917]_ ;
  assign \new_[1983]_  = \new_[16908]_  & \new_[16899]_ ;
  assign \new_[1984]_  = \new_[16890]_  & \new_[16881]_ ;
  assign \new_[1985]_  = \new_[16872]_  & \new_[16863]_ ;
  assign \new_[1986]_  = \new_[16854]_  & \new_[16845]_ ;
  assign \new_[1987]_  = \new_[16836]_  & \new_[16827]_ ;
  assign \new_[1988]_  = \new_[16818]_  & \new_[16809]_ ;
  assign \new_[1989]_  = \new_[16800]_  & \new_[16791]_ ;
  assign \new_[1990]_  = \new_[16782]_  & \new_[16773]_ ;
  assign \new_[1991]_  = \new_[16764]_  & \new_[16755]_ ;
  assign \new_[1992]_  = \new_[16746]_  & \new_[16737]_ ;
  assign \new_[1993]_  = \new_[16728]_  & \new_[16719]_ ;
  assign \new_[1994]_  = \new_[16710]_  & \new_[16701]_ ;
  assign \new_[1995]_  = \new_[16692]_  & \new_[16683]_ ;
  assign \new_[1996]_  = \new_[16674]_  & \new_[16665]_ ;
  assign \new_[1997]_  = \new_[16656]_  & \new_[16647]_ ;
  assign \new_[1998]_  = \new_[16638]_  & \new_[16629]_ ;
  assign \new_[1999]_  = \new_[16620]_  & \new_[16611]_ ;
  assign \new_[2000]_  = \new_[16602]_  & \new_[16593]_ ;
  assign \new_[2001]_  = \new_[16584]_  & \new_[16575]_ ;
  assign \new_[2002]_  = \new_[16566]_  & \new_[16557]_ ;
  assign \new_[2003]_  = \new_[16548]_  & \new_[16539]_ ;
  assign \new_[2004]_  = \new_[16530]_  & \new_[16521]_ ;
  assign \new_[2005]_  = \new_[16512]_  & \new_[16503]_ ;
  assign \new_[2006]_  = \new_[16494]_  & \new_[16485]_ ;
  assign \new_[2007]_  = \new_[16476]_  & \new_[16467]_ ;
  assign \new_[2008]_  = \new_[16458]_  & \new_[16449]_ ;
  assign \new_[2009]_  = \new_[16440]_  & \new_[16431]_ ;
  assign \new_[2010]_  = \new_[16422]_  & \new_[16413]_ ;
  assign \new_[2011]_  = \new_[16404]_  & \new_[16395]_ ;
  assign \new_[2012]_  = \new_[16386]_  & \new_[16377]_ ;
  assign \new_[2013]_  = \new_[16368]_  & \new_[16359]_ ;
  assign \new_[2014]_  = \new_[16350]_  & \new_[16341]_ ;
  assign \new_[2015]_  = \new_[16332]_  & \new_[16323]_ ;
  assign \new_[2016]_  = \new_[16314]_  & \new_[16305]_ ;
  assign \new_[2017]_  = \new_[16296]_  & \new_[16287]_ ;
  assign \new_[2018]_  = \new_[16278]_  & \new_[16269]_ ;
  assign \new_[2019]_  = \new_[16260]_  & \new_[16251]_ ;
  assign \new_[2020]_  = \new_[16242]_  & \new_[16233]_ ;
  assign \new_[2021]_  = \new_[16224]_  & \new_[16215]_ ;
  assign \new_[2022]_  = \new_[16206]_  & \new_[16197]_ ;
  assign \new_[2023]_  = \new_[16188]_  & \new_[16179]_ ;
  assign \new_[2024]_  = \new_[16170]_  & \new_[16161]_ ;
  assign \new_[2025]_  = \new_[16152]_  & \new_[16143]_ ;
  assign \new_[2026]_  = \new_[16134]_  & \new_[16125]_ ;
  assign \new_[2027]_  = \new_[16116]_  & \new_[16107]_ ;
  assign \new_[2028]_  = \new_[16098]_  & \new_[16089]_ ;
  assign \new_[2029]_  = \new_[16080]_  & \new_[16071]_ ;
  assign \new_[2030]_  = \new_[16062]_  & \new_[16053]_ ;
  assign \new_[2031]_  = \new_[16044]_  & \new_[16035]_ ;
  assign \new_[2032]_  = \new_[16026]_  & \new_[16017]_ ;
  assign \new_[2033]_  = \new_[16008]_  & \new_[15999]_ ;
  assign \new_[2034]_  = \new_[15990]_  & \new_[15981]_ ;
  assign \new_[2035]_  = \new_[15972]_  & \new_[15963]_ ;
  assign \new_[2036]_  = \new_[15954]_  & \new_[15945]_ ;
  assign \new_[2037]_  = \new_[15936]_  & \new_[15927]_ ;
  assign \new_[2038]_  = \new_[15918]_  & \new_[15909]_ ;
  assign \new_[2039]_  = \new_[15900]_  & \new_[15891]_ ;
  assign \new_[2040]_  = \new_[15882]_  & \new_[15873]_ ;
  assign \new_[2041]_  = \new_[15864]_  & \new_[15855]_ ;
  assign \new_[2042]_  = \new_[15846]_  & \new_[15837]_ ;
  assign \new_[2043]_  = \new_[15828]_  & \new_[15819]_ ;
  assign \new_[2044]_  = \new_[15810]_  & \new_[15801]_ ;
  assign \new_[2045]_  = \new_[15792]_  & \new_[15783]_ ;
  assign \new_[2046]_  = \new_[15774]_  & \new_[15765]_ ;
  assign \new_[2047]_  = \new_[15756]_  & \new_[15747]_ ;
  assign \new_[2048]_  = \new_[15738]_  & \new_[15729]_ ;
  assign \new_[2049]_  = \new_[15720]_  & \new_[15711]_ ;
  assign \new_[2050]_  = \new_[15702]_  & \new_[15693]_ ;
  assign \new_[2051]_  = \new_[15684]_  & \new_[15675]_ ;
  assign \new_[2052]_  = \new_[15666]_  & \new_[15657]_ ;
  assign \new_[2053]_  = \new_[15648]_  & \new_[15639]_ ;
  assign \new_[2054]_  = \new_[15630]_  & \new_[15621]_ ;
  assign \new_[2055]_  = \new_[15612]_  & \new_[15603]_ ;
  assign \new_[2056]_  = \new_[15594]_  & \new_[15585]_ ;
  assign \new_[2057]_  = \new_[15576]_  & \new_[15567]_ ;
  assign \new_[2058]_  = \new_[15558]_  & \new_[15549]_ ;
  assign \new_[2059]_  = \new_[15540]_  & \new_[15531]_ ;
  assign \new_[2060]_  = \new_[15522]_  & \new_[15513]_ ;
  assign \new_[2061]_  = \new_[15504]_  & \new_[15495]_ ;
  assign \new_[2062]_  = \new_[15486]_  & \new_[15477]_ ;
  assign \new_[2063]_  = \new_[15468]_  & \new_[15459]_ ;
  assign \new_[2064]_  = \new_[15450]_  & \new_[15441]_ ;
  assign \new_[2065]_  = \new_[15432]_  & \new_[15423]_ ;
  assign \new_[2066]_  = \new_[15414]_  & \new_[15405]_ ;
  assign \new_[2067]_  = \new_[15396]_  & \new_[15387]_ ;
  assign \new_[2068]_  = \new_[15378]_  & \new_[15369]_ ;
  assign \new_[2069]_  = \new_[15360]_  & \new_[15351]_ ;
  assign \new_[2070]_  = \new_[15342]_  & \new_[15333]_ ;
  assign \new_[2071]_  = \new_[15324]_  & \new_[15315]_ ;
  assign \new_[2072]_  = \new_[15306]_  & \new_[15297]_ ;
  assign \new_[2073]_  = \new_[15288]_  & \new_[15279]_ ;
  assign \new_[2074]_  = \new_[15270]_  & \new_[15261]_ ;
  assign \new_[2075]_  = \new_[15252]_  & \new_[15243]_ ;
  assign \new_[2076]_  = \new_[15234]_  & \new_[15225]_ ;
  assign \new_[2077]_  = \new_[15216]_  & \new_[15207]_ ;
  assign \new_[2078]_  = \new_[15198]_  & \new_[15189]_ ;
  assign \new_[2079]_  = \new_[15180]_  & \new_[15171]_ ;
  assign \new_[2080]_  = \new_[15162]_  & \new_[15153]_ ;
  assign \new_[2081]_  = \new_[15144]_  & \new_[15135]_ ;
  assign \new_[2082]_  = \new_[15126]_  & \new_[15117]_ ;
  assign \new_[2083]_  = \new_[15108]_  & \new_[15099]_ ;
  assign \new_[2084]_  = \new_[15090]_  & \new_[15081]_ ;
  assign \new_[2085]_  = \new_[15072]_  & \new_[15063]_ ;
  assign \new_[2086]_  = \new_[15054]_  & \new_[15045]_ ;
  assign \new_[2087]_  = \new_[15036]_  & \new_[15027]_ ;
  assign \new_[2088]_  = \new_[15018]_  & \new_[15009]_ ;
  assign \new_[2089]_  = \new_[15000]_  & \new_[14991]_ ;
  assign \new_[2090]_  = \new_[14982]_  & \new_[14973]_ ;
  assign \new_[2091]_  = \new_[14964]_  & \new_[14955]_ ;
  assign \new_[2092]_  = \new_[14946]_  & \new_[14937]_ ;
  assign \new_[2093]_  = \new_[14928]_  & \new_[14919]_ ;
  assign \new_[2094]_  = \new_[14910]_  & \new_[14901]_ ;
  assign \new_[2095]_  = \new_[14892]_  & \new_[14883]_ ;
  assign \new_[2096]_  = \new_[14874]_  & \new_[14865]_ ;
  assign \new_[2097]_  = \new_[14856]_  & \new_[14847]_ ;
  assign \new_[2098]_  = \new_[14838]_  & \new_[14829]_ ;
  assign \new_[2099]_  = \new_[14820]_  & \new_[14811]_ ;
  assign \new_[2100]_  = \new_[14802]_  & \new_[14793]_ ;
  assign \new_[2101]_  = \new_[14784]_  & \new_[14775]_ ;
  assign \new_[2102]_  = \new_[14766]_  & \new_[14757]_ ;
  assign \new_[2103]_  = \new_[14748]_  & \new_[14739]_ ;
  assign \new_[2104]_  = \new_[14730]_  & \new_[14721]_ ;
  assign \new_[2105]_  = \new_[14712]_  & \new_[14703]_ ;
  assign \new_[2106]_  = \new_[14694]_  & \new_[14685]_ ;
  assign \new_[2107]_  = \new_[14676]_  & \new_[14667]_ ;
  assign \new_[2108]_  = \new_[14658]_  & \new_[14649]_ ;
  assign \new_[2109]_  = \new_[14640]_  & \new_[14631]_ ;
  assign \new_[2110]_  = \new_[14622]_  & \new_[14613]_ ;
  assign \new_[2111]_  = \new_[14604]_  & \new_[14595]_ ;
  assign \new_[2112]_  = \new_[14586]_  & \new_[14577]_ ;
  assign \new_[2113]_  = \new_[14568]_  & \new_[14559]_ ;
  assign \new_[2114]_  = \new_[14550]_  & \new_[14541]_ ;
  assign \new_[2115]_  = \new_[14532]_  & \new_[14523]_ ;
  assign \new_[2116]_  = \new_[14514]_  & \new_[14505]_ ;
  assign \new_[2117]_  = \new_[14496]_  & \new_[14487]_ ;
  assign \new_[2118]_  = \new_[14478]_  & \new_[14469]_ ;
  assign \new_[2119]_  = \new_[14460]_  & \new_[14451]_ ;
  assign \new_[2120]_  = \new_[14442]_  & \new_[14433]_ ;
  assign \new_[2121]_  = \new_[14424]_  & \new_[14415]_ ;
  assign \new_[2122]_  = \new_[14406]_  & \new_[14397]_ ;
  assign \new_[2123]_  = \new_[14388]_  & \new_[14379]_ ;
  assign \new_[2124]_  = \new_[14370]_  & \new_[14361]_ ;
  assign \new_[2125]_  = \new_[14352]_  & \new_[14343]_ ;
  assign \new_[2126]_  = \new_[14334]_  & \new_[14325]_ ;
  assign \new_[2127]_  = \new_[14316]_  & \new_[14307]_ ;
  assign \new_[2128]_  = \new_[14298]_  & \new_[14289]_ ;
  assign \new_[2129]_  = \new_[14280]_  & \new_[14271]_ ;
  assign \new_[2130]_  = \new_[14262]_  & \new_[14253]_ ;
  assign \new_[2131]_  = \new_[14244]_  & \new_[14235]_ ;
  assign \new_[2132]_  = \new_[14226]_  & \new_[14217]_ ;
  assign \new_[2133]_  = \new_[14208]_  & \new_[14199]_ ;
  assign \new_[2134]_  = \new_[14190]_  & \new_[14181]_ ;
  assign \new_[2135]_  = \new_[14172]_  & \new_[14163]_ ;
  assign \new_[2136]_  = \new_[14154]_  & \new_[14145]_ ;
  assign \new_[2137]_  = \new_[14136]_  & \new_[14127]_ ;
  assign \new_[2138]_  = \new_[14118]_  & \new_[14109]_ ;
  assign \new_[2139]_  = \new_[14100]_  & \new_[14091]_ ;
  assign \new_[2140]_  = \new_[14082]_  & \new_[14073]_ ;
  assign \new_[2141]_  = \new_[14064]_  & \new_[14055]_ ;
  assign \new_[2142]_  = \new_[14046]_  & \new_[14037]_ ;
  assign \new_[2143]_  = \new_[14028]_  & \new_[14019]_ ;
  assign \new_[2144]_  = \new_[14010]_  & \new_[14001]_ ;
  assign \new_[2145]_  = \new_[13992]_  & \new_[13983]_ ;
  assign \new_[2146]_  = \new_[13974]_  & \new_[13965]_ ;
  assign \new_[2147]_  = \new_[13956]_  & \new_[13947]_ ;
  assign \new_[2148]_  = \new_[13938]_  & \new_[13929]_ ;
  assign \new_[2149]_  = \new_[13920]_  & \new_[13911]_ ;
  assign \new_[2150]_  = \new_[13902]_  & \new_[13893]_ ;
  assign \new_[2151]_  = \new_[13884]_  & \new_[13875]_ ;
  assign \new_[2152]_  = \new_[13866]_  & \new_[13857]_ ;
  assign \new_[2153]_  = \new_[13848]_  & \new_[13839]_ ;
  assign \new_[2154]_  = \new_[13830]_  & \new_[13821]_ ;
  assign \new_[2155]_  = \new_[13812]_  & \new_[13803]_ ;
  assign \new_[2156]_  = \new_[13794]_  & \new_[13785]_ ;
  assign \new_[2157]_  = \new_[13776]_  & \new_[13767]_ ;
  assign \new_[2158]_  = \new_[13758]_  & \new_[13749]_ ;
  assign \new_[2159]_  = \new_[13740]_  & \new_[13731]_ ;
  assign \new_[2160]_  = \new_[13722]_  & \new_[13713]_ ;
  assign \new_[2161]_  = \new_[13704]_  & \new_[13695]_ ;
  assign \new_[2162]_  = \new_[13686]_  & \new_[13677]_ ;
  assign \new_[2163]_  = \new_[13668]_  & \new_[13659]_ ;
  assign \new_[2164]_  = \new_[13650]_  & \new_[13641]_ ;
  assign \new_[2165]_  = \new_[13632]_  & \new_[13623]_ ;
  assign \new_[2166]_  = \new_[13614]_  & \new_[13605]_ ;
  assign \new_[2167]_  = \new_[13596]_  & \new_[13587]_ ;
  assign \new_[2168]_  = \new_[13578]_  & \new_[13569]_ ;
  assign \new_[2169]_  = \new_[13560]_  & \new_[13551]_ ;
  assign \new_[2170]_  = \new_[13542]_  & \new_[13533]_ ;
  assign \new_[2171]_  = \new_[13524]_  & \new_[13515]_ ;
  assign \new_[2172]_  = \new_[13506]_  & \new_[13497]_ ;
  assign \new_[2173]_  = \new_[13488]_  & \new_[13479]_ ;
  assign \new_[2174]_  = \new_[13470]_  & \new_[13461]_ ;
  assign \new_[2175]_  = \new_[13452]_  & \new_[13443]_ ;
  assign \new_[2176]_  = \new_[13434]_  & \new_[13425]_ ;
  assign \new_[2177]_  = \new_[13416]_  & \new_[13407]_ ;
  assign \new_[2178]_  = \new_[13398]_  & \new_[13389]_ ;
  assign \new_[2179]_  = \new_[13380]_  & \new_[13371]_ ;
  assign \new_[2180]_  = \new_[13362]_  & \new_[13353]_ ;
  assign \new_[2181]_  = \new_[13344]_  & \new_[13335]_ ;
  assign \new_[2182]_  = \new_[13326]_  & \new_[13317]_ ;
  assign \new_[2183]_  = \new_[13308]_  & \new_[13299]_ ;
  assign \new_[2184]_  = \new_[13290]_  & \new_[13281]_ ;
  assign \new_[2185]_  = \new_[13272]_  & \new_[13263]_ ;
  assign \new_[2186]_  = \new_[13254]_  & \new_[13245]_ ;
  assign \new_[2187]_  = \new_[13236]_  & \new_[13227]_ ;
  assign \new_[2188]_  = \new_[13218]_  & \new_[13209]_ ;
  assign \new_[2189]_  = \new_[13200]_  & \new_[13191]_ ;
  assign \new_[2190]_  = \new_[13182]_  & \new_[13173]_ ;
  assign \new_[2191]_  = \new_[13164]_  & \new_[13155]_ ;
  assign \new_[2192]_  = \new_[13146]_  & \new_[13137]_ ;
  assign \new_[2193]_  = \new_[13128]_  & \new_[13119]_ ;
  assign \new_[2194]_  = \new_[13110]_  & \new_[13101]_ ;
  assign \new_[2195]_  = \new_[13092]_  & \new_[13083]_ ;
  assign \new_[2196]_  = \new_[13074]_  & \new_[13065]_ ;
  assign \new_[2197]_  = \new_[13056]_  & \new_[13047]_ ;
  assign \new_[2198]_  = \new_[13038]_  & \new_[13029]_ ;
  assign \new_[2199]_  = \new_[13020]_  & \new_[13011]_ ;
  assign \new_[2200]_  = \new_[13002]_  & \new_[12993]_ ;
  assign \new_[2201]_  = \new_[12984]_  & \new_[12975]_ ;
  assign \new_[2202]_  = \new_[12966]_  & \new_[12957]_ ;
  assign \new_[2203]_  = \new_[12948]_  & \new_[12939]_ ;
  assign \new_[2204]_  = \new_[12930]_  & \new_[12921]_ ;
  assign \new_[2205]_  = \new_[12912]_  & \new_[12903]_ ;
  assign \new_[2206]_  = \new_[12894]_  & \new_[12885]_ ;
  assign \new_[2207]_  = \new_[12876]_  & \new_[12867]_ ;
  assign \new_[2208]_  = \new_[12858]_  & \new_[12849]_ ;
  assign \new_[2209]_  = \new_[12840]_  & \new_[12831]_ ;
  assign \new_[2210]_  = \new_[12822]_  & \new_[12813]_ ;
  assign \new_[2211]_  = \new_[12804]_  & \new_[12795]_ ;
  assign \new_[2212]_  = \new_[12786]_  & \new_[12777]_ ;
  assign \new_[2213]_  = \new_[12768]_  & \new_[12759]_ ;
  assign \new_[2214]_  = \new_[12750]_  & \new_[12741]_ ;
  assign \new_[2215]_  = \new_[12732]_  & \new_[12723]_ ;
  assign \new_[2216]_  = \new_[12714]_  & \new_[12705]_ ;
  assign \new_[2217]_  = \new_[12696]_  & \new_[12687]_ ;
  assign \new_[2218]_  = \new_[12678]_  & \new_[12669]_ ;
  assign \new_[2219]_  = \new_[12660]_  & \new_[12651]_ ;
  assign \new_[2220]_  = \new_[12642]_  & \new_[12633]_ ;
  assign \new_[2221]_  = \new_[12624]_  & \new_[12615]_ ;
  assign \new_[2222]_  = \new_[12606]_  & \new_[12597]_ ;
  assign \new_[2223]_  = \new_[12588]_  & \new_[12579]_ ;
  assign \new_[2224]_  = \new_[12570]_  & \new_[12561]_ ;
  assign \new_[2225]_  = \new_[12552]_  & \new_[12543]_ ;
  assign \new_[2226]_  = \new_[12536]_  & \new_[12527]_ ;
  assign \new_[2227]_  = \new_[12520]_  & \new_[12511]_ ;
  assign \new_[2228]_  = \new_[12504]_  & \new_[12495]_ ;
  assign \new_[2229]_  = \new_[12488]_  & \new_[12479]_ ;
  assign \new_[2230]_  = \new_[12472]_  & \new_[12463]_ ;
  assign \new_[2231]_  = \new_[12456]_  & \new_[12447]_ ;
  assign \new_[2232]_  = \new_[12440]_  & \new_[12431]_ ;
  assign \new_[2233]_  = \new_[12424]_  & \new_[12415]_ ;
  assign \new_[2234]_  = \new_[12408]_  & \new_[12399]_ ;
  assign \new_[2235]_  = \new_[12392]_  & \new_[12383]_ ;
  assign \new_[2236]_  = \new_[12376]_  & \new_[12367]_ ;
  assign \new_[2237]_  = \new_[12360]_  & \new_[12351]_ ;
  assign \new_[2238]_  = \new_[12344]_  & \new_[12335]_ ;
  assign \new_[2239]_  = \new_[12328]_  & \new_[12319]_ ;
  assign \new_[2240]_  = \new_[12312]_  & \new_[12303]_ ;
  assign \new_[2241]_  = \new_[12296]_  & \new_[12287]_ ;
  assign \new_[2242]_  = \new_[12280]_  & \new_[12271]_ ;
  assign \new_[2243]_  = \new_[12264]_  & \new_[12255]_ ;
  assign \new_[2244]_  = \new_[12248]_  & \new_[12239]_ ;
  assign \new_[2245]_  = \new_[12232]_  & \new_[12223]_ ;
  assign \new_[2246]_  = \new_[12216]_  & \new_[12207]_ ;
  assign \new_[2247]_  = \new_[12200]_  & \new_[12191]_ ;
  assign \new_[2248]_  = \new_[12184]_  & \new_[12175]_ ;
  assign \new_[2249]_  = \new_[12168]_  & \new_[12159]_ ;
  assign \new_[2250]_  = \new_[12152]_  & \new_[12143]_ ;
  assign \new_[2251]_  = \new_[12136]_  & \new_[12127]_ ;
  assign \new_[2252]_  = \new_[12120]_  & \new_[12111]_ ;
  assign \new_[2253]_  = \new_[12104]_  & \new_[12095]_ ;
  assign \new_[2254]_  = \new_[12088]_  & \new_[12079]_ ;
  assign \new_[2255]_  = \new_[12072]_  & \new_[12063]_ ;
  assign \new_[2256]_  = \new_[12056]_  & \new_[12047]_ ;
  assign \new_[2257]_  = \new_[12040]_  & \new_[12031]_ ;
  assign \new_[2258]_  = \new_[12024]_  & \new_[12015]_ ;
  assign \new_[2259]_  = \new_[12008]_  & \new_[11999]_ ;
  assign \new_[2260]_  = \new_[11992]_  & \new_[11983]_ ;
  assign \new_[2261]_  = \new_[11976]_  & \new_[11967]_ ;
  assign \new_[2262]_  = \new_[11960]_  & \new_[11951]_ ;
  assign \new_[2263]_  = \new_[11944]_  & \new_[11935]_ ;
  assign \new_[2264]_  = \new_[11928]_  & \new_[11919]_ ;
  assign \new_[2265]_  = \new_[11912]_  & \new_[11903]_ ;
  assign \new_[2266]_  = \new_[11896]_  & \new_[11887]_ ;
  assign \new_[2267]_  = \new_[11880]_  & \new_[11871]_ ;
  assign \new_[2268]_  = \new_[11864]_  & \new_[11855]_ ;
  assign \new_[2269]_  = \new_[11848]_  & \new_[11839]_ ;
  assign \new_[2270]_  = \new_[11832]_  & \new_[11823]_ ;
  assign \new_[2271]_  = \new_[11816]_  & \new_[11807]_ ;
  assign \new_[2272]_  = \new_[11800]_  & \new_[11791]_ ;
  assign \new_[2273]_  = \new_[11784]_  & \new_[11775]_ ;
  assign \new_[2274]_  = \new_[11768]_  & \new_[11759]_ ;
  assign \new_[2275]_  = \new_[11752]_  & \new_[11743]_ ;
  assign \new_[2276]_  = \new_[11736]_  & \new_[11727]_ ;
  assign \new_[2277]_  = \new_[11720]_  & \new_[11711]_ ;
  assign \new_[2278]_  = \new_[11704]_  & \new_[11695]_ ;
  assign \new_[2279]_  = \new_[11688]_  & \new_[11679]_ ;
  assign \new_[2280]_  = \new_[11672]_  & \new_[11663]_ ;
  assign \new_[2281]_  = \new_[11656]_  & \new_[11647]_ ;
  assign \new_[2282]_  = \new_[11640]_  & \new_[11631]_ ;
  assign \new_[2283]_  = \new_[11624]_  & \new_[11615]_ ;
  assign \new_[2284]_  = \new_[11608]_  & \new_[11599]_ ;
  assign \new_[2285]_  = \new_[11592]_  & \new_[11583]_ ;
  assign \new_[2286]_  = \new_[11576]_  & \new_[11567]_ ;
  assign \new_[2287]_  = \new_[11560]_  & \new_[11551]_ ;
  assign \new_[2288]_  = \new_[11544]_  & \new_[11535]_ ;
  assign \new_[2289]_  = \new_[11528]_  & \new_[11519]_ ;
  assign \new_[2290]_  = \new_[11512]_  & \new_[11503]_ ;
  assign \new_[2291]_  = \new_[11496]_  & \new_[11487]_ ;
  assign \new_[2292]_  = \new_[11480]_  & \new_[11471]_ ;
  assign \new_[2293]_  = \new_[11464]_  & \new_[11455]_ ;
  assign \new_[2294]_  = \new_[11448]_  & \new_[11439]_ ;
  assign \new_[2295]_  = \new_[11432]_  & \new_[11423]_ ;
  assign \new_[2296]_  = \new_[11416]_  & \new_[11407]_ ;
  assign \new_[2297]_  = \new_[11400]_  & \new_[11391]_ ;
  assign \new_[2298]_  = \new_[11384]_  & \new_[11375]_ ;
  assign \new_[2299]_  = \new_[11368]_  & \new_[11359]_ ;
  assign \new_[2300]_  = \new_[11352]_  & \new_[11343]_ ;
  assign \new_[2301]_  = \new_[11336]_  & \new_[11327]_ ;
  assign \new_[2302]_  = \new_[11320]_  & \new_[11311]_ ;
  assign \new_[2303]_  = \new_[11304]_  & \new_[11295]_ ;
  assign \new_[2304]_  = \new_[11288]_  & \new_[11279]_ ;
  assign \new_[2305]_  = \new_[11272]_  & \new_[11263]_ ;
  assign \new_[2306]_  = \new_[11256]_  & \new_[11247]_ ;
  assign \new_[2307]_  = \new_[11240]_  & \new_[11231]_ ;
  assign \new_[2308]_  = \new_[11224]_  & \new_[11215]_ ;
  assign \new_[2309]_  = \new_[11208]_  & \new_[11199]_ ;
  assign \new_[2310]_  = \new_[11192]_  & \new_[11183]_ ;
  assign \new_[2311]_  = \new_[11176]_  & \new_[11167]_ ;
  assign \new_[2312]_  = \new_[11160]_  & \new_[11151]_ ;
  assign \new_[2313]_  = \new_[11144]_  & \new_[11135]_ ;
  assign \new_[2314]_  = \new_[11128]_  & \new_[11119]_ ;
  assign \new_[2315]_  = \new_[11112]_  & \new_[11103]_ ;
  assign \new_[2316]_  = \new_[11096]_  & \new_[11087]_ ;
  assign \new_[2317]_  = \new_[11080]_  & \new_[11071]_ ;
  assign \new_[2318]_  = \new_[11064]_  & \new_[11055]_ ;
  assign \new_[2319]_  = \new_[11048]_  & \new_[11039]_ ;
  assign \new_[2320]_  = \new_[11032]_  & \new_[11023]_ ;
  assign \new_[2321]_  = \new_[11016]_  & \new_[11007]_ ;
  assign \new_[2322]_  = \new_[11000]_  & \new_[10991]_ ;
  assign \new_[2323]_  = \new_[10984]_  & \new_[10975]_ ;
  assign \new_[2324]_  = \new_[10968]_  & \new_[10959]_ ;
  assign \new_[2325]_  = \new_[10952]_  & \new_[10943]_ ;
  assign \new_[2326]_  = \new_[10936]_  & \new_[10927]_ ;
  assign \new_[2327]_  = \new_[10920]_  & \new_[10911]_ ;
  assign \new_[2328]_  = \new_[10904]_  & \new_[10895]_ ;
  assign \new_[2329]_  = \new_[10888]_  & \new_[10879]_ ;
  assign \new_[2330]_  = \new_[10872]_  & \new_[10863]_ ;
  assign \new_[2331]_  = \new_[10856]_  & \new_[10847]_ ;
  assign \new_[2332]_  = \new_[10840]_  & \new_[10831]_ ;
  assign \new_[2333]_  = \new_[10824]_  & \new_[10815]_ ;
  assign \new_[2334]_  = \new_[10808]_  & \new_[10799]_ ;
  assign \new_[2335]_  = \new_[10792]_  & \new_[10783]_ ;
  assign \new_[2336]_  = \new_[10776]_  & \new_[10767]_ ;
  assign \new_[2337]_  = \new_[10760]_  & \new_[10751]_ ;
  assign \new_[2338]_  = \new_[10744]_  & \new_[10735]_ ;
  assign \new_[2339]_  = \new_[10728]_  & \new_[10719]_ ;
  assign \new_[2340]_  = \new_[10712]_  & \new_[10703]_ ;
  assign \new_[2341]_  = \new_[10696]_  & \new_[10687]_ ;
  assign \new_[2342]_  = \new_[10680]_  & \new_[10671]_ ;
  assign \new_[2343]_  = \new_[10664]_  & \new_[10655]_ ;
  assign \new_[2344]_  = \new_[10648]_  & \new_[10639]_ ;
  assign \new_[2345]_  = \new_[10632]_  & \new_[10623]_ ;
  assign \new_[2346]_  = \new_[10616]_  & \new_[10607]_ ;
  assign \new_[2347]_  = \new_[10600]_  & \new_[10591]_ ;
  assign \new_[2348]_  = \new_[10584]_  & \new_[10575]_ ;
  assign \new_[2349]_  = \new_[10568]_  & \new_[10559]_ ;
  assign \new_[2350]_  = \new_[10552]_  & \new_[10543]_ ;
  assign \new_[2351]_  = \new_[10536]_  & \new_[10527]_ ;
  assign \new_[2352]_  = \new_[10520]_  & \new_[10511]_ ;
  assign \new_[2353]_  = \new_[10504]_  & \new_[10495]_ ;
  assign \new_[2354]_  = \new_[10488]_  & \new_[10479]_ ;
  assign \new_[2355]_  = \new_[10472]_  & \new_[10463]_ ;
  assign \new_[2356]_  = \new_[10456]_  & \new_[10447]_ ;
  assign \new_[2357]_  = \new_[10440]_  & \new_[10431]_ ;
  assign \new_[2358]_  = \new_[10424]_  & \new_[10415]_ ;
  assign \new_[2359]_  = \new_[10408]_  & \new_[10399]_ ;
  assign \new_[2360]_  = \new_[10392]_  & \new_[10383]_ ;
  assign \new_[2361]_  = \new_[10376]_  & \new_[10367]_ ;
  assign \new_[2362]_  = \new_[10360]_  & \new_[10351]_ ;
  assign \new_[2363]_  = \new_[10344]_  & \new_[10335]_ ;
  assign \new_[2364]_  = \new_[10328]_  & \new_[10319]_ ;
  assign \new_[2365]_  = \new_[10312]_  & \new_[10303]_ ;
  assign \new_[2366]_  = \new_[10296]_  & \new_[10287]_ ;
  assign \new_[2367]_  = \new_[10280]_  & \new_[10271]_ ;
  assign \new_[2368]_  = \new_[10264]_  & \new_[10255]_ ;
  assign \new_[2369]_  = \new_[10248]_  & \new_[10239]_ ;
  assign \new_[2370]_  = \new_[10232]_  & \new_[10223]_ ;
  assign \new_[2371]_  = \new_[10216]_  & \new_[10207]_ ;
  assign \new_[2372]_  = \new_[10200]_  & \new_[10191]_ ;
  assign \new_[2373]_  = \new_[10184]_  & \new_[10175]_ ;
  assign \new_[2374]_  = \new_[10168]_  & \new_[10159]_ ;
  assign \new_[2375]_  = \new_[10152]_  & \new_[10143]_ ;
  assign \new_[2376]_  = \new_[10136]_  & \new_[10127]_ ;
  assign \new_[2377]_  = \new_[10120]_  & \new_[10111]_ ;
  assign \new_[2378]_  = \new_[10104]_  & \new_[10095]_ ;
  assign \new_[2379]_  = \new_[10088]_  & \new_[10079]_ ;
  assign \new_[2380]_  = \new_[10072]_  & \new_[10063]_ ;
  assign \new_[2381]_  = \new_[10056]_  & \new_[10047]_ ;
  assign \new_[2382]_  = \new_[10040]_  & \new_[10031]_ ;
  assign \new_[2383]_  = \new_[10024]_  & \new_[10015]_ ;
  assign \new_[2384]_  = \new_[10008]_  & \new_[9999]_ ;
  assign \new_[2385]_  = \new_[9992]_  & \new_[9983]_ ;
  assign \new_[2386]_  = \new_[9976]_  & \new_[9967]_ ;
  assign \new_[2387]_  = \new_[9960]_  & \new_[9951]_ ;
  assign \new_[2388]_  = \new_[9944]_  & \new_[9935]_ ;
  assign \new_[2389]_  = \new_[9928]_  & \new_[9919]_ ;
  assign \new_[2390]_  = \new_[9912]_  & \new_[9903]_ ;
  assign \new_[2391]_  = \new_[9896]_  & \new_[9887]_ ;
  assign \new_[2392]_  = \new_[9880]_  & \new_[9871]_ ;
  assign \new_[2393]_  = \new_[9864]_  & \new_[9855]_ ;
  assign \new_[2394]_  = \new_[9848]_  & \new_[9839]_ ;
  assign \new_[2395]_  = \new_[9832]_  & \new_[9823]_ ;
  assign \new_[2396]_  = \new_[9816]_  & \new_[9807]_ ;
  assign \new_[2397]_  = \new_[9800]_  & \new_[9791]_ ;
  assign \new_[2398]_  = \new_[9784]_  & \new_[9775]_ ;
  assign \new_[2399]_  = \new_[9768]_  & \new_[9759]_ ;
  assign \new_[2400]_  = \new_[9752]_  & \new_[9743]_ ;
  assign \new_[2401]_  = \new_[9736]_  & \new_[9727]_ ;
  assign \new_[2402]_  = \new_[9720]_  & \new_[9711]_ ;
  assign \new_[2403]_  = \new_[9704]_  & \new_[9695]_ ;
  assign \new_[2404]_  = \new_[9688]_  & \new_[9679]_ ;
  assign \new_[2405]_  = \new_[9672]_  & \new_[9663]_ ;
  assign \new_[2406]_  = \new_[9656]_  & \new_[9647]_ ;
  assign \new_[2407]_  = \new_[9640]_  & \new_[9631]_ ;
  assign \new_[2408]_  = \new_[9624]_  & \new_[9615]_ ;
  assign \new_[2409]_  = \new_[9608]_  & \new_[9599]_ ;
  assign \new_[2410]_  = \new_[9592]_  & \new_[9583]_ ;
  assign \new_[2411]_  = \new_[9576]_  & \new_[9567]_ ;
  assign \new_[2412]_  = \new_[9560]_  & \new_[9551]_ ;
  assign \new_[2413]_  = \new_[9544]_  & \new_[9535]_ ;
  assign \new_[2414]_  = \new_[9528]_  & \new_[9519]_ ;
  assign \new_[2415]_  = \new_[9512]_  & \new_[9503]_ ;
  assign \new_[2416]_  = \new_[9496]_  & \new_[9487]_ ;
  assign \new_[2417]_  = \new_[9480]_  & \new_[9471]_ ;
  assign \new_[2418]_  = \new_[9464]_  & \new_[9455]_ ;
  assign \new_[2419]_  = \new_[9448]_  & \new_[9439]_ ;
  assign \new_[2420]_  = \new_[9432]_  & \new_[9423]_ ;
  assign \new_[2421]_  = \new_[9416]_  & \new_[9407]_ ;
  assign \new_[2422]_  = \new_[9400]_  & \new_[9391]_ ;
  assign \new_[2423]_  = \new_[9384]_  & \new_[9375]_ ;
  assign \new_[2424]_  = \new_[9368]_  & \new_[9359]_ ;
  assign \new_[2425]_  = \new_[9352]_  & \new_[9343]_ ;
  assign \new_[2426]_  = \new_[9336]_  & \new_[9327]_ ;
  assign \new_[2427]_  = \new_[9320]_  & \new_[9311]_ ;
  assign \new_[2428]_  = \new_[9304]_  & \new_[9295]_ ;
  assign \new_[2429]_  = \new_[9288]_  & \new_[9281]_ ;
  assign \new_[2430]_  = \new_[9274]_  & \new_[9267]_ ;
  assign \new_[2431]_  = \new_[9260]_  & \new_[9253]_ ;
  assign \new_[2432]_  = \new_[9246]_  & \new_[9239]_ ;
  assign \new_[2433]_  = \new_[9232]_  & \new_[9225]_ ;
  assign \new_[2434]_  = \new_[9218]_  & \new_[9211]_ ;
  assign \new_[2435]_  = \new_[9204]_  & \new_[9197]_ ;
  assign \new_[2436]_  = \new_[9190]_  & \new_[9183]_ ;
  assign \new_[2437]_  = \new_[9176]_  & \new_[9169]_ ;
  assign \new_[2438]_  = \new_[9162]_  & \new_[9155]_ ;
  assign \new_[2439]_  = \new_[9148]_  & \new_[9141]_ ;
  assign \new_[2440]_  = \new_[9134]_  & \new_[9127]_ ;
  assign \new_[2441]_  = \new_[9120]_  & \new_[9113]_ ;
  assign \new_[2442]_  = \new_[9106]_  & \new_[9099]_ ;
  assign \new_[2443]_  = \new_[9092]_  & \new_[9085]_ ;
  assign \new_[2444]_  = \new_[9078]_  & \new_[9071]_ ;
  assign \new_[2445]_  = \new_[9064]_  & \new_[9057]_ ;
  assign \new_[2446]_  = \new_[9050]_  & \new_[9043]_ ;
  assign \new_[2447]_  = \new_[9036]_  & \new_[9029]_ ;
  assign \new_[2448]_  = \new_[9022]_  & \new_[9015]_ ;
  assign \new_[2449]_  = \new_[9008]_  & \new_[9001]_ ;
  assign \new_[2450]_  = \new_[8994]_  & \new_[8987]_ ;
  assign \new_[2451]_  = \new_[8980]_  & \new_[8973]_ ;
  assign \new_[2452]_  = \new_[8966]_  & \new_[8959]_ ;
  assign \new_[2453]_  = \new_[8952]_  & \new_[8945]_ ;
  assign \new_[2454]_  = \new_[8938]_  & \new_[8931]_ ;
  assign \new_[2455]_  = \new_[8924]_  & \new_[8917]_ ;
  assign \new_[2456]_  = \new_[8910]_  & \new_[8903]_ ;
  assign \new_[2457]_  = \new_[8896]_  & \new_[8889]_ ;
  assign \new_[2458]_  = \new_[8882]_  & \new_[8875]_ ;
  assign \new_[2459]_  = \new_[8868]_  & \new_[8861]_ ;
  assign \new_[2460]_  = \new_[8854]_  & \new_[8847]_ ;
  assign \new_[2461]_  = \new_[8840]_  & \new_[8833]_ ;
  assign \new_[2462]_  = \new_[8826]_  & \new_[8819]_ ;
  assign \new_[2463]_  = \new_[8812]_  & \new_[8805]_ ;
  assign \new_[2464]_  = \new_[8798]_  & \new_[8791]_ ;
  assign \new_[2465]_  = \new_[8784]_  & \new_[8777]_ ;
  assign \new_[2466]_  = \new_[8770]_  & \new_[8763]_ ;
  assign \new_[2467]_  = \new_[8756]_  & \new_[8749]_ ;
  assign \new_[2468]_  = \new_[8742]_  & \new_[8735]_ ;
  assign \new_[2469]_  = \new_[8728]_  & \new_[8721]_ ;
  assign \new_[2470]_  = \new_[8714]_  & \new_[8707]_ ;
  assign \new_[2471]_  = \new_[8700]_  & \new_[8693]_ ;
  assign \new_[2472]_  = \new_[8686]_  & \new_[8679]_ ;
  assign \new_[2473]_  = \new_[8672]_  & \new_[8665]_ ;
  assign \new_[2474]_  = \new_[8658]_  & \new_[8651]_ ;
  assign \new_[2475]_  = \new_[8644]_  & \new_[8637]_ ;
  assign \new_[2476]_  = \new_[8630]_  & \new_[8623]_ ;
  assign \new_[2477]_  = \new_[8616]_  & \new_[8609]_ ;
  assign \new_[2478]_  = \new_[8602]_  & \new_[8595]_ ;
  assign \new_[2479]_  = \new_[8588]_  & \new_[8581]_ ;
  assign \new_[2480]_  = \new_[8574]_  & \new_[8567]_ ;
  assign \new_[2481]_  = \new_[8560]_  & \new_[8553]_ ;
  assign \new_[2482]_  = \new_[8546]_  & \new_[8539]_ ;
  assign \new_[2483]_  = \new_[8532]_  & \new_[8525]_ ;
  assign \new_[2484]_  = \new_[8518]_  & \new_[8511]_ ;
  assign \new_[2485]_  = \new_[8504]_  & \new_[8497]_ ;
  assign \new_[2486]_  = \new_[8490]_  & \new_[8483]_ ;
  assign \new_[2487]_  = \new_[8476]_  & \new_[8469]_ ;
  assign \new_[2488]_  = \new_[8462]_  & \new_[8455]_ ;
  assign \new_[2489]_  = \new_[8448]_  & \new_[8441]_ ;
  assign \new_[2490]_  = \new_[8434]_  & \new_[8427]_ ;
  assign \new_[2491]_  = \new_[8420]_  & \new_[8413]_ ;
  assign \new_[2492]_  = \new_[8406]_  & \new_[8399]_ ;
  assign \new_[2493]_  = \new_[8392]_  & \new_[8385]_ ;
  assign \new_[2494]_  = \new_[8378]_  & \new_[8371]_ ;
  assign \new_[2495]_  = \new_[8364]_  & \new_[8357]_ ;
  assign \new_[2496]_  = \new_[8350]_  & \new_[8343]_ ;
  assign \new_[2497]_  = \new_[8336]_  & \new_[8329]_ ;
  assign \new_[2498]_  = \new_[8322]_  & \new_[8315]_ ;
  assign \new_[2499]_  = \new_[8308]_  & \new_[8301]_ ;
  assign \new_[2500]_  = \new_[8294]_  & \new_[8287]_ ;
  assign \new_[2501]_  = \new_[8280]_  & \new_[8273]_ ;
  assign \new_[2502]_  = \new_[8266]_  & \new_[8259]_ ;
  assign \new_[2503]_  = \new_[8252]_  & \new_[8245]_ ;
  assign \new_[2504]_  = \new_[8238]_  & \new_[8231]_ ;
  assign \new_[2505]_  = \new_[8224]_  & \new_[8217]_ ;
  assign \new_[2506]_  = \new_[8210]_  & \new_[8203]_ ;
  assign \new_[2507]_  = \new_[8196]_  & \new_[8189]_ ;
  assign \new_[2508]_  = \new_[8182]_  & \new_[8175]_ ;
  assign \new_[2509]_  = \new_[8168]_  & \new_[8161]_ ;
  assign \new_[2510]_  = \new_[8154]_  & \new_[8147]_ ;
  assign \new_[2511]_  = \new_[8140]_  & \new_[8133]_ ;
  assign \new_[2512]_  = \new_[8126]_  & \new_[8119]_ ;
  assign \new_[2513]_  = \new_[8112]_  & \new_[8105]_ ;
  assign \new_[2514]_  = \new_[8098]_  & \new_[8091]_ ;
  assign \new_[2515]_  = \new_[8084]_  & \new_[8077]_ ;
  assign \new_[2516]_  = \new_[8070]_  & \new_[8063]_ ;
  assign \new_[2517]_  = \new_[8056]_  & \new_[8049]_ ;
  assign \new_[2518]_  = \new_[8042]_  & \new_[8035]_ ;
  assign \new_[2519]_  = \new_[8028]_  & \new_[8021]_ ;
  assign \new_[2520]_  = \new_[8014]_  & \new_[8007]_ ;
  assign \new_[2521]_  = \new_[8000]_  & \new_[7993]_ ;
  assign \new_[2522]_  = \new_[7988]_  & \new_[7981]_ ;
  assign \new_[2523]_  = \new_[7976]_  & \new_[7969]_ ;
  assign \new_[2524]_  = \new_[7964]_  & \new_[7957]_ ;
  assign \new_[2525]_  = \new_[7952]_  & \new_[7945]_ ;
  assign \new_[2526]_  = \new_[7940]_  & \new_[7933]_ ;
  assign \new_[2527]_  = \new_[7928]_  & \new_[7921]_ ;
  assign \new_[2528]_  = \new_[7916]_  & \new_[7909]_ ;
  assign \new_[2529]_  = \new_[7904]_  & \new_[7897]_ ;
  assign \new_[2530]_  = \new_[7892]_  & \new_[7885]_ ;
  assign \new_[2531]_  = \new_[7880]_  & \new_[7873]_ ;
  assign \new_[2532]_  = \new_[7868]_  & \new_[7861]_ ;
  assign \new_[2533]_  = \new_[7856]_  & \new_[7849]_ ;
  assign \new_[2534]_  = \new_[7844]_  & \new_[7837]_ ;
  assign \new_[2535]_  = \new_[7832]_  & \new_[7825]_ ;
  assign \new_[2536]_  = \new_[7820]_  & \new_[7813]_ ;
  assign \new_[2537]_  = \new_[7808]_  & \new_[7801]_ ;
  assign \new_[2538]_  = \new_[7796]_  & \new_[7789]_ ;
  assign \new_[2539]_  = \new_[7784]_  & \new_[7777]_ ;
  assign \new_[2540]_  = \new_[7772]_  & \new_[7765]_ ;
  assign \new_[2541]_  = \new_[7760]_  & \new_[7753]_ ;
  assign \new_[2542]_  = \new_[7748]_  & \new_[7741]_ ;
  assign \new_[2543]_  = \new_[7736]_  & \new_[7729]_ ;
  assign \new_[2544]_  = \new_[7724]_  & \new_[7717]_ ;
  assign \new_[2545]_  = \new_[7712]_  & \new_[7705]_ ;
  assign \new_[2546]_  = \new_[7700]_  & \new_[7693]_ ;
  assign \new_[2547]_  = \new_[7688]_  & \new_[7683]_ ;
  assign \new_[2548]_  = \new_[7678]_  & \new_[7673]_ ;
  assign \new_[2549]_  = \new_[7668]_  & \new_[7663]_ ;
  assign \new_[2550]_  = \new_[7658]_  & \new_[7653]_ ;
  assign \new_[2553]_  = \new_[2549]_  | \new_[2550]_ ;
  assign \new_[2556]_  = \new_[2547]_  | \new_[2548]_ ;
  assign \new_[2557]_  = \new_[2556]_  | \new_[2553]_ ;
  assign \new_[2560]_  = \new_[2545]_  | \new_[2546]_ ;
  assign \new_[2564]_  = \new_[2542]_  | \new_[2543]_ ;
  assign \new_[2565]_  = \new_[2544]_  | \new_[2564]_ ;
  assign \new_[2566]_  = \new_[2565]_  | \new_[2560]_ ;
  assign \new_[2567]_  = \new_[2566]_  | \new_[2557]_ ;
  assign \new_[2570]_  = \new_[2540]_  | \new_[2541]_ ;
  assign \new_[2574]_  = \new_[2537]_  | \new_[2538]_ ;
  assign \new_[2575]_  = \new_[2539]_  | \new_[2574]_ ;
  assign \new_[2576]_  = \new_[2575]_  | \new_[2570]_ ;
  assign \new_[2579]_  = \new_[2535]_  | \new_[2536]_ ;
  assign \new_[2583]_  = \new_[2532]_  | \new_[2533]_ ;
  assign \new_[2584]_  = \new_[2534]_  | \new_[2583]_ ;
  assign \new_[2585]_  = \new_[2584]_  | \new_[2579]_ ;
  assign \new_[2586]_  = \new_[2585]_  | \new_[2576]_ ;
  assign \new_[2587]_  = \new_[2586]_  | \new_[2567]_ ;
  assign \new_[2590]_  = \new_[2530]_  | \new_[2531]_ ;
  assign \new_[2594]_  = \new_[2527]_  | \new_[2528]_ ;
  assign \new_[2595]_  = \new_[2529]_  | \new_[2594]_ ;
  assign \new_[2596]_  = \new_[2595]_  | \new_[2590]_ ;
  assign \new_[2599]_  = \new_[2525]_  | \new_[2526]_ ;
  assign \new_[2603]_  = \new_[2522]_  | \new_[2523]_ ;
  assign \new_[2604]_  = \new_[2524]_  | \new_[2603]_ ;
  assign \new_[2605]_  = \new_[2604]_  | \new_[2599]_ ;
  assign \new_[2606]_  = \new_[2605]_  | \new_[2596]_ ;
  assign \new_[2609]_  = \new_[2520]_  | \new_[2521]_ ;
  assign \new_[2613]_  = \new_[2517]_  | \new_[2518]_ ;
  assign \new_[2614]_  = \new_[2519]_  | \new_[2613]_ ;
  assign \new_[2615]_  = \new_[2614]_  | \new_[2609]_ ;
  assign \new_[2618]_  = \new_[2515]_  | \new_[2516]_ ;
  assign \new_[2622]_  = \new_[2512]_  | \new_[2513]_ ;
  assign \new_[2623]_  = \new_[2514]_  | \new_[2622]_ ;
  assign \new_[2624]_  = \new_[2623]_  | \new_[2618]_ ;
  assign \new_[2625]_  = \new_[2624]_  | \new_[2615]_ ;
  assign \new_[2626]_  = \new_[2625]_  | \new_[2606]_ ;
  assign \new_[2627]_  = \new_[2626]_  | \new_[2587]_ ;
  assign \new_[2630]_  = \new_[2510]_  | \new_[2511]_ ;
  assign \new_[2634]_  = \new_[2507]_  | \new_[2508]_ ;
  assign \new_[2635]_  = \new_[2509]_  | \new_[2634]_ ;
  assign \new_[2636]_  = \new_[2635]_  | \new_[2630]_ ;
  assign \new_[2639]_  = \new_[2505]_  | \new_[2506]_ ;
  assign \new_[2643]_  = \new_[2502]_  | \new_[2503]_ ;
  assign \new_[2644]_  = \new_[2504]_  | \new_[2643]_ ;
  assign \new_[2645]_  = \new_[2644]_  | \new_[2639]_ ;
  assign \new_[2646]_  = \new_[2645]_  | \new_[2636]_ ;
  assign \new_[2649]_  = \new_[2500]_  | \new_[2501]_ ;
  assign \new_[2653]_  = \new_[2497]_  | \new_[2498]_ ;
  assign \new_[2654]_  = \new_[2499]_  | \new_[2653]_ ;
  assign \new_[2655]_  = \new_[2654]_  | \new_[2649]_ ;
  assign \new_[2658]_  = \new_[2495]_  | \new_[2496]_ ;
  assign \new_[2662]_  = \new_[2492]_  | \new_[2493]_ ;
  assign \new_[2663]_  = \new_[2494]_  | \new_[2662]_ ;
  assign \new_[2664]_  = \new_[2663]_  | \new_[2658]_ ;
  assign \new_[2665]_  = \new_[2664]_  | \new_[2655]_ ;
  assign \new_[2666]_  = \new_[2665]_  | \new_[2646]_ ;
  assign \new_[2669]_  = \new_[2490]_  | \new_[2491]_ ;
  assign \new_[2673]_  = \new_[2487]_  | \new_[2488]_ ;
  assign \new_[2674]_  = \new_[2489]_  | \new_[2673]_ ;
  assign \new_[2675]_  = \new_[2674]_  | \new_[2669]_ ;
  assign \new_[2678]_  = \new_[2485]_  | \new_[2486]_ ;
  assign \new_[2682]_  = \new_[2482]_  | \new_[2483]_ ;
  assign \new_[2683]_  = \new_[2484]_  | \new_[2682]_ ;
  assign \new_[2684]_  = \new_[2683]_  | \new_[2678]_ ;
  assign \new_[2685]_  = \new_[2684]_  | \new_[2675]_ ;
  assign \new_[2688]_  = \new_[2480]_  | \new_[2481]_ ;
  assign \new_[2692]_  = \new_[2477]_  | \new_[2478]_ ;
  assign \new_[2693]_  = \new_[2479]_  | \new_[2692]_ ;
  assign \new_[2694]_  = \new_[2693]_  | \new_[2688]_ ;
  assign \new_[2697]_  = \new_[2475]_  | \new_[2476]_ ;
  assign \new_[2701]_  = \new_[2472]_  | \new_[2473]_ ;
  assign \new_[2702]_  = \new_[2474]_  | \new_[2701]_ ;
  assign \new_[2703]_  = \new_[2702]_  | \new_[2697]_ ;
  assign \new_[2704]_  = \new_[2703]_  | \new_[2694]_ ;
  assign \new_[2705]_  = \new_[2704]_  | \new_[2685]_ ;
  assign \new_[2706]_  = \new_[2705]_  | \new_[2666]_ ;
  assign \new_[2707]_  = \new_[2706]_  | \new_[2627]_ ;
  assign \new_[2710]_  = \new_[2470]_  | \new_[2471]_ ;
  assign \new_[2714]_  = \new_[2467]_  | \new_[2468]_ ;
  assign \new_[2715]_  = \new_[2469]_  | \new_[2714]_ ;
  assign \new_[2716]_  = \new_[2715]_  | \new_[2710]_ ;
  assign \new_[2719]_  = \new_[2465]_  | \new_[2466]_ ;
  assign \new_[2723]_  = \new_[2462]_  | \new_[2463]_ ;
  assign \new_[2724]_  = \new_[2464]_  | \new_[2723]_ ;
  assign \new_[2725]_  = \new_[2724]_  | \new_[2719]_ ;
  assign \new_[2726]_  = \new_[2725]_  | \new_[2716]_ ;
  assign \new_[2729]_  = \new_[2460]_  | \new_[2461]_ ;
  assign \new_[2733]_  = \new_[2457]_  | \new_[2458]_ ;
  assign \new_[2734]_  = \new_[2459]_  | \new_[2733]_ ;
  assign \new_[2735]_  = \new_[2734]_  | \new_[2729]_ ;
  assign \new_[2738]_  = \new_[2455]_  | \new_[2456]_ ;
  assign \new_[2742]_  = \new_[2452]_  | \new_[2453]_ ;
  assign \new_[2743]_  = \new_[2454]_  | \new_[2742]_ ;
  assign \new_[2744]_  = \new_[2743]_  | \new_[2738]_ ;
  assign \new_[2745]_  = \new_[2744]_  | \new_[2735]_ ;
  assign \new_[2746]_  = \new_[2745]_  | \new_[2726]_ ;
  assign \new_[2749]_  = \new_[2450]_  | \new_[2451]_ ;
  assign \new_[2753]_  = \new_[2447]_  | \new_[2448]_ ;
  assign \new_[2754]_  = \new_[2449]_  | \new_[2753]_ ;
  assign \new_[2755]_  = \new_[2754]_  | \new_[2749]_ ;
  assign \new_[2758]_  = \new_[2445]_  | \new_[2446]_ ;
  assign \new_[2762]_  = \new_[2442]_  | \new_[2443]_ ;
  assign \new_[2763]_  = \new_[2444]_  | \new_[2762]_ ;
  assign \new_[2764]_  = \new_[2763]_  | \new_[2758]_ ;
  assign \new_[2765]_  = \new_[2764]_  | \new_[2755]_ ;
  assign \new_[2768]_  = \new_[2440]_  | \new_[2441]_ ;
  assign \new_[2772]_  = \new_[2437]_  | \new_[2438]_ ;
  assign \new_[2773]_  = \new_[2439]_  | \new_[2772]_ ;
  assign \new_[2774]_  = \new_[2773]_  | \new_[2768]_ ;
  assign \new_[2777]_  = \new_[2435]_  | \new_[2436]_ ;
  assign \new_[2781]_  = \new_[2432]_  | \new_[2433]_ ;
  assign \new_[2782]_  = \new_[2434]_  | \new_[2781]_ ;
  assign \new_[2783]_  = \new_[2782]_  | \new_[2777]_ ;
  assign \new_[2784]_  = \new_[2783]_  | \new_[2774]_ ;
  assign \new_[2785]_  = \new_[2784]_  | \new_[2765]_ ;
  assign \new_[2786]_  = \new_[2785]_  | \new_[2746]_ ;
  assign \new_[2789]_  = \new_[2430]_  | \new_[2431]_ ;
  assign \new_[2793]_  = \new_[2427]_  | \new_[2428]_ ;
  assign \new_[2794]_  = \new_[2429]_  | \new_[2793]_ ;
  assign \new_[2795]_  = \new_[2794]_  | \new_[2789]_ ;
  assign \new_[2798]_  = \new_[2425]_  | \new_[2426]_ ;
  assign \new_[2802]_  = \new_[2422]_  | \new_[2423]_ ;
  assign \new_[2803]_  = \new_[2424]_  | \new_[2802]_ ;
  assign \new_[2804]_  = \new_[2803]_  | \new_[2798]_ ;
  assign \new_[2805]_  = \new_[2804]_  | \new_[2795]_ ;
  assign \new_[2808]_  = \new_[2420]_  | \new_[2421]_ ;
  assign \new_[2812]_  = \new_[2417]_  | \new_[2418]_ ;
  assign \new_[2813]_  = \new_[2419]_  | \new_[2812]_ ;
  assign \new_[2814]_  = \new_[2813]_  | \new_[2808]_ ;
  assign \new_[2817]_  = \new_[2415]_  | \new_[2416]_ ;
  assign \new_[2821]_  = \new_[2412]_  | \new_[2413]_ ;
  assign \new_[2822]_  = \new_[2414]_  | \new_[2821]_ ;
  assign \new_[2823]_  = \new_[2822]_  | \new_[2817]_ ;
  assign \new_[2824]_  = \new_[2823]_  | \new_[2814]_ ;
  assign \new_[2825]_  = \new_[2824]_  | \new_[2805]_ ;
  assign \new_[2828]_  = \new_[2410]_  | \new_[2411]_ ;
  assign \new_[2832]_  = \new_[2407]_  | \new_[2408]_ ;
  assign \new_[2833]_  = \new_[2409]_  | \new_[2832]_ ;
  assign \new_[2834]_  = \new_[2833]_  | \new_[2828]_ ;
  assign \new_[2837]_  = \new_[2405]_  | \new_[2406]_ ;
  assign \new_[2841]_  = \new_[2402]_  | \new_[2403]_ ;
  assign \new_[2842]_  = \new_[2404]_  | \new_[2841]_ ;
  assign \new_[2843]_  = \new_[2842]_  | \new_[2837]_ ;
  assign \new_[2844]_  = \new_[2843]_  | \new_[2834]_ ;
  assign \new_[2847]_  = \new_[2400]_  | \new_[2401]_ ;
  assign \new_[2851]_  = \new_[2397]_  | \new_[2398]_ ;
  assign \new_[2852]_  = \new_[2399]_  | \new_[2851]_ ;
  assign \new_[2853]_  = \new_[2852]_  | \new_[2847]_ ;
  assign \new_[2856]_  = \new_[2395]_  | \new_[2396]_ ;
  assign \new_[2860]_  = \new_[2392]_  | \new_[2393]_ ;
  assign \new_[2861]_  = \new_[2394]_  | \new_[2860]_ ;
  assign \new_[2862]_  = \new_[2861]_  | \new_[2856]_ ;
  assign \new_[2863]_  = \new_[2862]_  | \new_[2853]_ ;
  assign \new_[2864]_  = \new_[2863]_  | \new_[2844]_ ;
  assign \new_[2865]_  = \new_[2864]_  | \new_[2825]_ ;
  assign \new_[2866]_  = \new_[2865]_  | \new_[2786]_ ;
  assign \new_[2867]_  = \new_[2866]_  | \new_[2707]_ ;
  assign \new_[2870]_  = \new_[2390]_  | \new_[2391]_ ;
  assign \new_[2873]_  = \new_[2388]_  | \new_[2389]_ ;
  assign \new_[2874]_  = \new_[2873]_  | \new_[2870]_ ;
  assign \new_[2877]_  = \new_[2386]_  | \new_[2387]_ ;
  assign \new_[2881]_  = \new_[2383]_  | \new_[2384]_ ;
  assign \new_[2882]_  = \new_[2385]_  | \new_[2881]_ ;
  assign \new_[2883]_  = \new_[2882]_  | \new_[2877]_ ;
  assign \new_[2884]_  = \new_[2883]_  | \new_[2874]_ ;
  assign \new_[2887]_  = \new_[2381]_  | \new_[2382]_ ;
  assign \new_[2891]_  = \new_[2378]_  | \new_[2379]_ ;
  assign \new_[2892]_  = \new_[2380]_  | \new_[2891]_ ;
  assign \new_[2893]_  = \new_[2892]_  | \new_[2887]_ ;
  assign \new_[2896]_  = \new_[2376]_  | \new_[2377]_ ;
  assign \new_[2900]_  = \new_[2373]_  | \new_[2374]_ ;
  assign \new_[2901]_  = \new_[2375]_  | \new_[2900]_ ;
  assign \new_[2902]_  = \new_[2901]_  | \new_[2896]_ ;
  assign \new_[2903]_  = \new_[2902]_  | \new_[2893]_ ;
  assign \new_[2904]_  = \new_[2903]_  | \new_[2884]_ ;
  assign \new_[2907]_  = \new_[2371]_  | \new_[2372]_ ;
  assign \new_[2911]_  = \new_[2368]_  | \new_[2369]_ ;
  assign \new_[2912]_  = \new_[2370]_  | \new_[2911]_ ;
  assign \new_[2913]_  = \new_[2912]_  | \new_[2907]_ ;
  assign \new_[2916]_  = \new_[2366]_  | \new_[2367]_ ;
  assign \new_[2920]_  = \new_[2363]_  | \new_[2364]_ ;
  assign \new_[2921]_  = \new_[2365]_  | \new_[2920]_ ;
  assign \new_[2922]_  = \new_[2921]_  | \new_[2916]_ ;
  assign \new_[2923]_  = \new_[2922]_  | \new_[2913]_ ;
  assign \new_[2926]_  = \new_[2361]_  | \new_[2362]_ ;
  assign \new_[2930]_  = \new_[2358]_  | \new_[2359]_ ;
  assign \new_[2931]_  = \new_[2360]_  | \new_[2930]_ ;
  assign \new_[2932]_  = \new_[2931]_  | \new_[2926]_ ;
  assign \new_[2935]_  = \new_[2356]_  | \new_[2357]_ ;
  assign \new_[2939]_  = \new_[2353]_  | \new_[2354]_ ;
  assign \new_[2940]_  = \new_[2355]_  | \new_[2939]_ ;
  assign \new_[2941]_  = \new_[2940]_  | \new_[2935]_ ;
  assign \new_[2942]_  = \new_[2941]_  | \new_[2932]_ ;
  assign \new_[2943]_  = \new_[2942]_  | \new_[2923]_ ;
  assign \new_[2944]_  = \new_[2943]_  | \new_[2904]_ ;
  assign \new_[2947]_  = \new_[2351]_  | \new_[2352]_ ;
  assign \new_[2951]_  = \new_[2348]_  | \new_[2349]_ ;
  assign \new_[2952]_  = \new_[2350]_  | \new_[2951]_ ;
  assign \new_[2953]_  = \new_[2952]_  | \new_[2947]_ ;
  assign \new_[2956]_  = \new_[2346]_  | \new_[2347]_ ;
  assign \new_[2960]_  = \new_[2343]_  | \new_[2344]_ ;
  assign \new_[2961]_  = \new_[2345]_  | \new_[2960]_ ;
  assign \new_[2962]_  = \new_[2961]_  | \new_[2956]_ ;
  assign \new_[2963]_  = \new_[2962]_  | \new_[2953]_ ;
  assign \new_[2966]_  = \new_[2341]_  | \new_[2342]_ ;
  assign \new_[2970]_  = \new_[2338]_  | \new_[2339]_ ;
  assign \new_[2971]_  = \new_[2340]_  | \new_[2970]_ ;
  assign \new_[2972]_  = \new_[2971]_  | \new_[2966]_ ;
  assign \new_[2975]_  = \new_[2336]_  | \new_[2337]_ ;
  assign \new_[2979]_  = \new_[2333]_  | \new_[2334]_ ;
  assign \new_[2980]_  = \new_[2335]_  | \new_[2979]_ ;
  assign \new_[2981]_  = \new_[2980]_  | \new_[2975]_ ;
  assign \new_[2982]_  = \new_[2981]_  | \new_[2972]_ ;
  assign \new_[2983]_  = \new_[2982]_  | \new_[2963]_ ;
  assign \new_[2986]_  = \new_[2331]_  | \new_[2332]_ ;
  assign \new_[2990]_  = \new_[2328]_  | \new_[2329]_ ;
  assign \new_[2991]_  = \new_[2330]_  | \new_[2990]_ ;
  assign \new_[2992]_  = \new_[2991]_  | \new_[2986]_ ;
  assign \new_[2995]_  = \new_[2326]_  | \new_[2327]_ ;
  assign \new_[2999]_  = \new_[2323]_  | \new_[2324]_ ;
  assign \new_[3000]_  = \new_[2325]_  | \new_[2999]_ ;
  assign \new_[3001]_  = \new_[3000]_  | \new_[2995]_ ;
  assign \new_[3002]_  = \new_[3001]_  | \new_[2992]_ ;
  assign \new_[3005]_  = \new_[2321]_  | \new_[2322]_ ;
  assign \new_[3009]_  = \new_[2318]_  | \new_[2319]_ ;
  assign \new_[3010]_  = \new_[2320]_  | \new_[3009]_ ;
  assign \new_[3011]_  = \new_[3010]_  | \new_[3005]_ ;
  assign \new_[3014]_  = \new_[2316]_  | \new_[2317]_ ;
  assign \new_[3018]_  = \new_[2313]_  | \new_[2314]_ ;
  assign \new_[3019]_  = \new_[2315]_  | \new_[3018]_ ;
  assign \new_[3020]_  = \new_[3019]_  | \new_[3014]_ ;
  assign \new_[3021]_  = \new_[3020]_  | \new_[3011]_ ;
  assign \new_[3022]_  = \new_[3021]_  | \new_[3002]_ ;
  assign \new_[3023]_  = \new_[3022]_  | \new_[2983]_ ;
  assign \new_[3024]_  = \new_[3023]_  | \new_[2944]_ ;
  assign \new_[3027]_  = \new_[2311]_  | \new_[2312]_ ;
  assign \new_[3031]_  = \new_[2308]_  | \new_[2309]_ ;
  assign \new_[3032]_  = \new_[2310]_  | \new_[3031]_ ;
  assign \new_[3033]_  = \new_[3032]_  | \new_[3027]_ ;
  assign \new_[3036]_  = \new_[2306]_  | \new_[2307]_ ;
  assign \new_[3040]_  = \new_[2303]_  | \new_[2304]_ ;
  assign \new_[3041]_  = \new_[2305]_  | \new_[3040]_ ;
  assign \new_[3042]_  = \new_[3041]_  | \new_[3036]_ ;
  assign \new_[3043]_  = \new_[3042]_  | \new_[3033]_ ;
  assign \new_[3046]_  = \new_[2301]_  | \new_[2302]_ ;
  assign \new_[3050]_  = \new_[2298]_  | \new_[2299]_ ;
  assign \new_[3051]_  = \new_[2300]_  | \new_[3050]_ ;
  assign \new_[3052]_  = \new_[3051]_  | \new_[3046]_ ;
  assign \new_[3055]_  = \new_[2296]_  | \new_[2297]_ ;
  assign \new_[3059]_  = \new_[2293]_  | \new_[2294]_ ;
  assign \new_[3060]_  = \new_[2295]_  | \new_[3059]_ ;
  assign \new_[3061]_  = \new_[3060]_  | \new_[3055]_ ;
  assign \new_[3062]_  = \new_[3061]_  | \new_[3052]_ ;
  assign \new_[3063]_  = \new_[3062]_  | \new_[3043]_ ;
  assign \new_[3066]_  = \new_[2291]_  | \new_[2292]_ ;
  assign \new_[3070]_  = \new_[2288]_  | \new_[2289]_ ;
  assign \new_[3071]_  = \new_[2290]_  | \new_[3070]_ ;
  assign \new_[3072]_  = \new_[3071]_  | \new_[3066]_ ;
  assign \new_[3075]_  = \new_[2286]_  | \new_[2287]_ ;
  assign \new_[3079]_  = \new_[2283]_  | \new_[2284]_ ;
  assign \new_[3080]_  = \new_[2285]_  | \new_[3079]_ ;
  assign \new_[3081]_  = \new_[3080]_  | \new_[3075]_ ;
  assign \new_[3082]_  = \new_[3081]_  | \new_[3072]_ ;
  assign \new_[3085]_  = \new_[2281]_  | \new_[2282]_ ;
  assign \new_[3089]_  = \new_[2278]_  | \new_[2279]_ ;
  assign \new_[3090]_  = \new_[2280]_  | \new_[3089]_ ;
  assign \new_[3091]_  = \new_[3090]_  | \new_[3085]_ ;
  assign \new_[3094]_  = \new_[2276]_  | \new_[2277]_ ;
  assign \new_[3098]_  = \new_[2273]_  | \new_[2274]_ ;
  assign \new_[3099]_  = \new_[2275]_  | \new_[3098]_ ;
  assign \new_[3100]_  = \new_[3099]_  | \new_[3094]_ ;
  assign \new_[3101]_  = \new_[3100]_  | \new_[3091]_ ;
  assign \new_[3102]_  = \new_[3101]_  | \new_[3082]_ ;
  assign \new_[3103]_  = \new_[3102]_  | \new_[3063]_ ;
  assign \new_[3106]_  = \new_[2271]_  | \new_[2272]_ ;
  assign \new_[3110]_  = \new_[2268]_  | \new_[2269]_ ;
  assign \new_[3111]_  = \new_[2270]_  | \new_[3110]_ ;
  assign \new_[3112]_  = \new_[3111]_  | \new_[3106]_ ;
  assign \new_[3115]_  = \new_[2266]_  | \new_[2267]_ ;
  assign \new_[3119]_  = \new_[2263]_  | \new_[2264]_ ;
  assign \new_[3120]_  = \new_[2265]_  | \new_[3119]_ ;
  assign \new_[3121]_  = \new_[3120]_  | \new_[3115]_ ;
  assign \new_[3122]_  = \new_[3121]_  | \new_[3112]_ ;
  assign \new_[3125]_  = \new_[2261]_  | \new_[2262]_ ;
  assign \new_[3129]_  = \new_[2258]_  | \new_[2259]_ ;
  assign \new_[3130]_  = \new_[2260]_  | \new_[3129]_ ;
  assign \new_[3131]_  = \new_[3130]_  | \new_[3125]_ ;
  assign \new_[3134]_  = \new_[2256]_  | \new_[2257]_ ;
  assign \new_[3138]_  = \new_[2253]_  | \new_[2254]_ ;
  assign \new_[3139]_  = \new_[2255]_  | \new_[3138]_ ;
  assign \new_[3140]_  = \new_[3139]_  | \new_[3134]_ ;
  assign \new_[3141]_  = \new_[3140]_  | \new_[3131]_ ;
  assign \new_[3142]_  = \new_[3141]_  | \new_[3122]_ ;
  assign \new_[3145]_  = \new_[2251]_  | \new_[2252]_ ;
  assign \new_[3149]_  = \new_[2248]_  | \new_[2249]_ ;
  assign \new_[3150]_  = \new_[2250]_  | \new_[3149]_ ;
  assign \new_[3151]_  = \new_[3150]_  | \new_[3145]_ ;
  assign \new_[3154]_  = \new_[2246]_  | \new_[2247]_ ;
  assign \new_[3158]_  = \new_[2243]_  | \new_[2244]_ ;
  assign \new_[3159]_  = \new_[2245]_  | \new_[3158]_ ;
  assign \new_[3160]_  = \new_[3159]_  | \new_[3154]_ ;
  assign \new_[3161]_  = \new_[3160]_  | \new_[3151]_ ;
  assign \new_[3164]_  = \new_[2241]_  | \new_[2242]_ ;
  assign \new_[3168]_  = \new_[2238]_  | \new_[2239]_ ;
  assign \new_[3169]_  = \new_[2240]_  | \new_[3168]_ ;
  assign \new_[3170]_  = \new_[3169]_  | \new_[3164]_ ;
  assign \new_[3173]_  = \new_[2236]_  | \new_[2237]_ ;
  assign \new_[3177]_  = \new_[2233]_  | \new_[2234]_ ;
  assign \new_[3178]_  = \new_[2235]_  | \new_[3177]_ ;
  assign \new_[3179]_  = \new_[3178]_  | \new_[3173]_ ;
  assign \new_[3180]_  = \new_[3179]_  | \new_[3170]_ ;
  assign \new_[3181]_  = \new_[3180]_  | \new_[3161]_ ;
  assign \new_[3182]_  = \new_[3181]_  | \new_[3142]_ ;
  assign \new_[3183]_  = \new_[3182]_  | \new_[3103]_ ;
  assign \new_[3184]_  = \new_[3183]_  | \new_[3024]_ ;
  assign \new_[3185]_  = \new_[3184]_  | \new_[2867]_ ;
  assign \new_[3188]_  = \new_[2231]_  | \new_[2232]_ ;
  assign \new_[3191]_  = \new_[2229]_  | \new_[2230]_ ;
  assign \new_[3192]_  = \new_[3191]_  | \new_[3188]_ ;
  assign \new_[3195]_  = \new_[2227]_  | \new_[2228]_ ;
  assign \new_[3199]_  = \new_[2224]_  | \new_[2225]_ ;
  assign \new_[3200]_  = \new_[2226]_  | \new_[3199]_ ;
  assign \new_[3201]_  = \new_[3200]_  | \new_[3195]_ ;
  assign \new_[3202]_  = \new_[3201]_  | \new_[3192]_ ;
  assign \new_[3205]_  = \new_[2222]_  | \new_[2223]_ ;
  assign \new_[3209]_  = \new_[2219]_  | \new_[2220]_ ;
  assign \new_[3210]_  = \new_[2221]_  | \new_[3209]_ ;
  assign \new_[3211]_  = \new_[3210]_  | \new_[3205]_ ;
  assign \new_[3214]_  = \new_[2217]_  | \new_[2218]_ ;
  assign \new_[3218]_  = \new_[2214]_  | \new_[2215]_ ;
  assign \new_[3219]_  = \new_[2216]_  | \new_[3218]_ ;
  assign \new_[3220]_  = \new_[3219]_  | \new_[3214]_ ;
  assign \new_[3221]_  = \new_[3220]_  | \new_[3211]_ ;
  assign \new_[3222]_  = \new_[3221]_  | \new_[3202]_ ;
  assign \new_[3225]_  = \new_[2212]_  | \new_[2213]_ ;
  assign \new_[3229]_  = \new_[2209]_  | \new_[2210]_ ;
  assign \new_[3230]_  = \new_[2211]_  | \new_[3229]_ ;
  assign \new_[3231]_  = \new_[3230]_  | \new_[3225]_ ;
  assign \new_[3234]_  = \new_[2207]_  | \new_[2208]_ ;
  assign \new_[3238]_  = \new_[2204]_  | \new_[2205]_ ;
  assign \new_[3239]_  = \new_[2206]_  | \new_[3238]_ ;
  assign \new_[3240]_  = \new_[3239]_  | \new_[3234]_ ;
  assign \new_[3241]_  = \new_[3240]_  | \new_[3231]_ ;
  assign \new_[3244]_  = \new_[2202]_  | \new_[2203]_ ;
  assign \new_[3248]_  = \new_[2199]_  | \new_[2200]_ ;
  assign \new_[3249]_  = \new_[2201]_  | \new_[3248]_ ;
  assign \new_[3250]_  = \new_[3249]_  | \new_[3244]_ ;
  assign \new_[3253]_  = \new_[2197]_  | \new_[2198]_ ;
  assign \new_[3257]_  = \new_[2194]_  | \new_[2195]_ ;
  assign \new_[3258]_  = \new_[2196]_  | \new_[3257]_ ;
  assign \new_[3259]_  = \new_[3258]_  | \new_[3253]_ ;
  assign \new_[3260]_  = \new_[3259]_  | \new_[3250]_ ;
  assign \new_[3261]_  = \new_[3260]_  | \new_[3241]_ ;
  assign \new_[3262]_  = \new_[3261]_  | \new_[3222]_ ;
  assign \new_[3265]_  = \new_[2192]_  | \new_[2193]_ ;
  assign \new_[3269]_  = \new_[2189]_  | \new_[2190]_ ;
  assign \new_[3270]_  = \new_[2191]_  | \new_[3269]_ ;
  assign \new_[3271]_  = \new_[3270]_  | \new_[3265]_ ;
  assign \new_[3274]_  = \new_[2187]_  | \new_[2188]_ ;
  assign \new_[3278]_  = \new_[2184]_  | \new_[2185]_ ;
  assign \new_[3279]_  = \new_[2186]_  | \new_[3278]_ ;
  assign \new_[3280]_  = \new_[3279]_  | \new_[3274]_ ;
  assign \new_[3281]_  = \new_[3280]_  | \new_[3271]_ ;
  assign \new_[3284]_  = \new_[2182]_  | \new_[2183]_ ;
  assign \new_[3288]_  = \new_[2179]_  | \new_[2180]_ ;
  assign \new_[3289]_  = \new_[2181]_  | \new_[3288]_ ;
  assign \new_[3290]_  = \new_[3289]_  | \new_[3284]_ ;
  assign \new_[3293]_  = \new_[2177]_  | \new_[2178]_ ;
  assign \new_[3297]_  = \new_[2174]_  | \new_[2175]_ ;
  assign \new_[3298]_  = \new_[2176]_  | \new_[3297]_ ;
  assign \new_[3299]_  = \new_[3298]_  | \new_[3293]_ ;
  assign \new_[3300]_  = \new_[3299]_  | \new_[3290]_ ;
  assign \new_[3301]_  = \new_[3300]_  | \new_[3281]_ ;
  assign \new_[3304]_  = \new_[2172]_  | \new_[2173]_ ;
  assign \new_[3308]_  = \new_[2169]_  | \new_[2170]_ ;
  assign \new_[3309]_  = \new_[2171]_  | \new_[3308]_ ;
  assign \new_[3310]_  = \new_[3309]_  | \new_[3304]_ ;
  assign \new_[3313]_  = \new_[2167]_  | \new_[2168]_ ;
  assign \new_[3317]_  = \new_[2164]_  | \new_[2165]_ ;
  assign \new_[3318]_  = \new_[2166]_  | \new_[3317]_ ;
  assign \new_[3319]_  = \new_[3318]_  | \new_[3313]_ ;
  assign \new_[3320]_  = \new_[3319]_  | \new_[3310]_ ;
  assign \new_[3323]_  = \new_[2162]_  | \new_[2163]_ ;
  assign \new_[3327]_  = \new_[2159]_  | \new_[2160]_ ;
  assign \new_[3328]_  = \new_[2161]_  | \new_[3327]_ ;
  assign \new_[3329]_  = \new_[3328]_  | \new_[3323]_ ;
  assign \new_[3332]_  = \new_[2157]_  | \new_[2158]_ ;
  assign \new_[3336]_  = \new_[2154]_  | \new_[2155]_ ;
  assign \new_[3337]_  = \new_[2156]_  | \new_[3336]_ ;
  assign \new_[3338]_  = \new_[3337]_  | \new_[3332]_ ;
  assign \new_[3339]_  = \new_[3338]_  | \new_[3329]_ ;
  assign \new_[3340]_  = \new_[3339]_  | \new_[3320]_ ;
  assign \new_[3341]_  = \new_[3340]_  | \new_[3301]_ ;
  assign \new_[3342]_  = \new_[3341]_  | \new_[3262]_ ;
  assign \new_[3345]_  = \new_[2152]_  | \new_[2153]_ ;
  assign \new_[3349]_  = \new_[2149]_  | \new_[2150]_ ;
  assign \new_[3350]_  = \new_[2151]_  | \new_[3349]_ ;
  assign \new_[3351]_  = \new_[3350]_  | \new_[3345]_ ;
  assign \new_[3354]_  = \new_[2147]_  | \new_[2148]_ ;
  assign \new_[3358]_  = \new_[2144]_  | \new_[2145]_ ;
  assign \new_[3359]_  = \new_[2146]_  | \new_[3358]_ ;
  assign \new_[3360]_  = \new_[3359]_  | \new_[3354]_ ;
  assign \new_[3361]_  = \new_[3360]_  | \new_[3351]_ ;
  assign \new_[3364]_  = \new_[2142]_  | \new_[2143]_ ;
  assign \new_[3368]_  = \new_[2139]_  | \new_[2140]_ ;
  assign \new_[3369]_  = \new_[2141]_  | \new_[3368]_ ;
  assign \new_[3370]_  = \new_[3369]_  | \new_[3364]_ ;
  assign \new_[3373]_  = \new_[2137]_  | \new_[2138]_ ;
  assign \new_[3377]_  = \new_[2134]_  | \new_[2135]_ ;
  assign \new_[3378]_  = \new_[2136]_  | \new_[3377]_ ;
  assign \new_[3379]_  = \new_[3378]_  | \new_[3373]_ ;
  assign \new_[3380]_  = \new_[3379]_  | \new_[3370]_ ;
  assign \new_[3381]_  = \new_[3380]_  | \new_[3361]_ ;
  assign \new_[3384]_  = \new_[2132]_  | \new_[2133]_ ;
  assign \new_[3388]_  = \new_[2129]_  | \new_[2130]_ ;
  assign \new_[3389]_  = \new_[2131]_  | \new_[3388]_ ;
  assign \new_[3390]_  = \new_[3389]_  | \new_[3384]_ ;
  assign \new_[3393]_  = \new_[2127]_  | \new_[2128]_ ;
  assign \new_[3397]_  = \new_[2124]_  | \new_[2125]_ ;
  assign \new_[3398]_  = \new_[2126]_  | \new_[3397]_ ;
  assign \new_[3399]_  = \new_[3398]_  | \new_[3393]_ ;
  assign \new_[3400]_  = \new_[3399]_  | \new_[3390]_ ;
  assign \new_[3403]_  = \new_[2122]_  | \new_[2123]_ ;
  assign \new_[3407]_  = \new_[2119]_  | \new_[2120]_ ;
  assign \new_[3408]_  = \new_[2121]_  | \new_[3407]_ ;
  assign \new_[3409]_  = \new_[3408]_  | \new_[3403]_ ;
  assign \new_[3412]_  = \new_[2117]_  | \new_[2118]_ ;
  assign \new_[3416]_  = \new_[2114]_  | \new_[2115]_ ;
  assign \new_[3417]_  = \new_[2116]_  | \new_[3416]_ ;
  assign \new_[3418]_  = \new_[3417]_  | \new_[3412]_ ;
  assign \new_[3419]_  = \new_[3418]_  | \new_[3409]_ ;
  assign \new_[3420]_  = \new_[3419]_  | \new_[3400]_ ;
  assign \new_[3421]_  = \new_[3420]_  | \new_[3381]_ ;
  assign \new_[3424]_  = \new_[2112]_  | \new_[2113]_ ;
  assign \new_[3428]_  = \new_[2109]_  | \new_[2110]_ ;
  assign \new_[3429]_  = \new_[2111]_  | \new_[3428]_ ;
  assign \new_[3430]_  = \new_[3429]_  | \new_[3424]_ ;
  assign \new_[3433]_  = \new_[2107]_  | \new_[2108]_ ;
  assign \new_[3437]_  = \new_[2104]_  | \new_[2105]_ ;
  assign \new_[3438]_  = \new_[2106]_  | \new_[3437]_ ;
  assign \new_[3439]_  = \new_[3438]_  | \new_[3433]_ ;
  assign \new_[3440]_  = \new_[3439]_  | \new_[3430]_ ;
  assign \new_[3443]_  = \new_[2102]_  | \new_[2103]_ ;
  assign \new_[3447]_  = \new_[2099]_  | \new_[2100]_ ;
  assign \new_[3448]_  = \new_[2101]_  | \new_[3447]_ ;
  assign \new_[3449]_  = \new_[3448]_  | \new_[3443]_ ;
  assign \new_[3452]_  = \new_[2097]_  | \new_[2098]_ ;
  assign \new_[3456]_  = \new_[2094]_  | \new_[2095]_ ;
  assign \new_[3457]_  = \new_[2096]_  | \new_[3456]_ ;
  assign \new_[3458]_  = \new_[3457]_  | \new_[3452]_ ;
  assign \new_[3459]_  = \new_[3458]_  | \new_[3449]_ ;
  assign \new_[3460]_  = \new_[3459]_  | \new_[3440]_ ;
  assign \new_[3463]_  = \new_[2092]_  | \new_[2093]_ ;
  assign \new_[3467]_  = \new_[2089]_  | \new_[2090]_ ;
  assign \new_[3468]_  = \new_[2091]_  | \new_[3467]_ ;
  assign \new_[3469]_  = \new_[3468]_  | \new_[3463]_ ;
  assign \new_[3472]_  = \new_[2087]_  | \new_[2088]_ ;
  assign \new_[3476]_  = \new_[2084]_  | \new_[2085]_ ;
  assign \new_[3477]_  = \new_[2086]_  | \new_[3476]_ ;
  assign \new_[3478]_  = \new_[3477]_  | \new_[3472]_ ;
  assign \new_[3479]_  = \new_[3478]_  | \new_[3469]_ ;
  assign \new_[3482]_  = \new_[2082]_  | \new_[2083]_ ;
  assign \new_[3486]_  = \new_[2079]_  | \new_[2080]_ ;
  assign \new_[3487]_  = \new_[2081]_  | \new_[3486]_ ;
  assign \new_[3488]_  = \new_[3487]_  | \new_[3482]_ ;
  assign \new_[3491]_  = \new_[2077]_  | \new_[2078]_ ;
  assign \new_[3495]_  = \new_[2074]_  | \new_[2075]_ ;
  assign \new_[3496]_  = \new_[2076]_  | \new_[3495]_ ;
  assign \new_[3497]_  = \new_[3496]_  | \new_[3491]_ ;
  assign \new_[3498]_  = \new_[3497]_  | \new_[3488]_ ;
  assign \new_[3499]_  = \new_[3498]_  | \new_[3479]_ ;
  assign \new_[3500]_  = \new_[3499]_  | \new_[3460]_ ;
  assign \new_[3501]_  = \new_[3500]_  | \new_[3421]_ ;
  assign \new_[3502]_  = \new_[3501]_  | \new_[3342]_ ;
  assign \new_[3505]_  = \new_[2072]_  | \new_[2073]_ ;
  assign \new_[3509]_  = \new_[2069]_  | \new_[2070]_ ;
  assign \new_[3510]_  = \new_[2071]_  | \new_[3509]_ ;
  assign \new_[3511]_  = \new_[3510]_  | \new_[3505]_ ;
  assign \new_[3514]_  = \new_[2067]_  | \new_[2068]_ ;
  assign \new_[3518]_  = \new_[2064]_  | \new_[2065]_ ;
  assign \new_[3519]_  = \new_[2066]_  | \new_[3518]_ ;
  assign \new_[3520]_  = \new_[3519]_  | \new_[3514]_ ;
  assign \new_[3521]_  = \new_[3520]_  | \new_[3511]_ ;
  assign \new_[3524]_  = \new_[2062]_  | \new_[2063]_ ;
  assign \new_[3528]_  = \new_[2059]_  | \new_[2060]_ ;
  assign \new_[3529]_  = \new_[2061]_  | \new_[3528]_ ;
  assign \new_[3530]_  = \new_[3529]_  | \new_[3524]_ ;
  assign \new_[3533]_  = \new_[2057]_  | \new_[2058]_ ;
  assign \new_[3537]_  = \new_[2054]_  | \new_[2055]_ ;
  assign \new_[3538]_  = \new_[2056]_  | \new_[3537]_ ;
  assign \new_[3539]_  = \new_[3538]_  | \new_[3533]_ ;
  assign \new_[3540]_  = \new_[3539]_  | \new_[3530]_ ;
  assign \new_[3541]_  = \new_[3540]_  | \new_[3521]_ ;
  assign \new_[3544]_  = \new_[2052]_  | \new_[2053]_ ;
  assign \new_[3548]_  = \new_[2049]_  | \new_[2050]_ ;
  assign \new_[3549]_  = \new_[2051]_  | \new_[3548]_ ;
  assign \new_[3550]_  = \new_[3549]_  | \new_[3544]_ ;
  assign \new_[3553]_  = \new_[2047]_  | \new_[2048]_ ;
  assign \new_[3557]_  = \new_[2044]_  | \new_[2045]_ ;
  assign \new_[3558]_  = \new_[2046]_  | \new_[3557]_ ;
  assign \new_[3559]_  = \new_[3558]_  | \new_[3553]_ ;
  assign \new_[3560]_  = \new_[3559]_  | \new_[3550]_ ;
  assign \new_[3563]_  = \new_[2042]_  | \new_[2043]_ ;
  assign \new_[3567]_  = \new_[2039]_  | \new_[2040]_ ;
  assign \new_[3568]_  = \new_[2041]_  | \new_[3567]_ ;
  assign \new_[3569]_  = \new_[3568]_  | \new_[3563]_ ;
  assign \new_[3572]_  = \new_[2037]_  | \new_[2038]_ ;
  assign \new_[3576]_  = \new_[2034]_  | \new_[2035]_ ;
  assign \new_[3577]_  = \new_[2036]_  | \new_[3576]_ ;
  assign \new_[3578]_  = \new_[3577]_  | \new_[3572]_ ;
  assign \new_[3579]_  = \new_[3578]_  | \new_[3569]_ ;
  assign \new_[3580]_  = \new_[3579]_  | \new_[3560]_ ;
  assign \new_[3581]_  = \new_[3580]_  | \new_[3541]_ ;
  assign \new_[3584]_  = \new_[2032]_  | \new_[2033]_ ;
  assign \new_[3588]_  = \new_[2029]_  | \new_[2030]_ ;
  assign \new_[3589]_  = \new_[2031]_  | \new_[3588]_ ;
  assign \new_[3590]_  = \new_[3589]_  | \new_[3584]_ ;
  assign \new_[3593]_  = \new_[2027]_  | \new_[2028]_ ;
  assign \new_[3597]_  = \new_[2024]_  | \new_[2025]_ ;
  assign \new_[3598]_  = \new_[2026]_  | \new_[3597]_ ;
  assign \new_[3599]_  = \new_[3598]_  | \new_[3593]_ ;
  assign \new_[3600]_  = \new_[3599]_  | \new_[3590]_ ;
  assign \new_[3603]_  = \new_[2022]_  | \new_[2023]_ ;
  assign \new_[3607]_  = \new_[2019]_  | \new_[2020]_ ;
  assign \new_[3608]_  = \new_[2021]_  | \new_[3607]_ ;
  assign \new_[3609]_  = \new_[3608]_  | \new_[3603]_ ;
  assign \new_[3612]_  = \new_[2017]_  | \new_[2018]_ ;
  assign \new_[3616]_  = \new_[2014]_  | \new_[2015]_ ;
  assign \new_[3617]_  = \new_[2016]_  | \new_[3616]_ ;
  assign \new_[3618]_  = \new_[3617]_  | \new_[3612]_ ;
  assign \new_[3619]_  = \new_[3618]_  | \new_[3609]_ ;
  assign \new_[3620]_  = \new_[3619]_  | \new_[3600]_ ;
  assign \new_[3623]_  = \new_[2012]_  | \new_[2013]_ ;
  assign \new_[3627]_  = \new_[2009]_  | \new_[2010]_ ;
  assign \new_[3628]_  = \new_[2011]_  | \new_[3627]_ ;
  assign \new_[3629]_  = \new_[3628]_  | \new_[3623]_ ;
  assign \new_[3632]_  = \new_[2007]_  | \new_[2008]_ ;
  assign \new_[3636]_  = \new_[2004]_  | \new_[2005]_ ;
  assign \new_[3637]_  = \new_[2006]_  | \new_[3636]_ ;
  assign \new_[3638]_  = \new_[3637]_  | \new_[3632]_ ;
  assign \new_[3639]_  = \new_[3638]_  | \new_[3629]_ ;
  assign \new_[3642]_  = \new_[2002]_  | \new_[2003]_ ;
  assign \new_[3646]_  = \new_[1999]_  | \new_[2000]_ ;
  assign \new_[3647]_  = \new_[2001]_  | \new_[3646]_ ;
  assign \new_[3648]_  = \new_[3647]_  | \new_[3642]_ ;
  assign \new_[3651]_  = \new_[1997]_  | \new_[1998]_ ;
  assign \new_[3655]_  = \new_[1994]_  | \new_[1995]_ ;
  assign \new_[3656]_  = \new_[1996]_  | \new_[3655]_ ;
  assign \new_[3657]_  = \new_[3656]_  | \new_[3651]_ ;
  assign \new_[3658]_  = \new_[3657]_  | \new_[3648]_ ;
  assign \new_[3659]_  = \new_[3658]_  | \new_[3639]_ ;
  assign \new_[3660]_  = \new_[3659]_  | \new_[3620]_ ;
  assign \new_[3661]_  = \new_[3660]_  | \new_[3581]_ ;
  assign \new_[3664]_  = \new_[1992]_  | \new_[1993]_ ;
  assign \new_[3668]_  = \new_[1989]_  | \new_[1990]_ ;
  assign \new_[3669]_  = \new_[1991]_  | \new_[3668]_ ;
  assign \new_[3670]_  = \new_[3669]_  | \new_[3664]_ ;
  assign \new_[3673]_  = \new_[1987]_  | \new_[1988]_ ;
  assign \new_[3677]_  = \new_[1984]_  | \new_[1985]_ ;
  assign \new_[3678]_  = \new_[1986]_  | \new_[3677]_ ;
  assign \new_[3679]_  = \new_[3678]_  | \new_[3673]_ ;
  assign \new_[3680]_  = \new_[3679]_  | \new_[3670]_ ;
  assign \new_[3683]_  = \new_[1982]_  | \new_[1983]_ ;
  assign \new_[3687]_  = \new_[1979]_  | \new_[1980]_ ;
  assign \new_[3688]_  = \new_[1981]_  | \new_[3687]_ ;
  assign \new_[3689]_  = \new_[3688]_  | \new_[3683]_ ;
  assign \new_[3692]_  = \new_[1977]_  | \new_[1978]_ ;
  assign \new_[3696]_  = \new_[1974]_  | \new_[1975]_ ;
  assign \new_[3697]_  = \new_[1976]_  | \new_[3696]_ ;
  assign \new_[3698]_  = \new_[3697]_  | \new_[3692]_ ;
  assign \new_[3699]_  = \new_[3698]_  | \new_[3689]_ ;
  assign \new_[3700]_  = \new_[3699]_  | \new_[3680]_ ;
  assign \new_[3703]_  = \new_[1972]_  | \new_[1973]_ ;
  assign \new_[3707]_  = \new_[1969]_  | \new_[1970]_ ;
  assign \new_[3708]_  = \new_[1971]_  | \new_[3707]_ ;
  assign \new_[3709]_  = \new_[3708]_  | \new_[3703]_ ;
  assign \new_[3712]_  = \new_[1967]_  | \new_[1968]_ ;
  assign \new_[3716]_  = \new_[1964]_  | \new_[1965]_ ;
  assign \new_[3717]_  = \new_[1966]_  | \new_[3716]_ ;
  assign \new_[3718]_  = \new_[3717]_  | \new_[3712]_ ;
  assign \new_[3719]_  = \new_[3718]_  | \new_[3709]_ ;
  assign \new_[3722]_  = \new_[1962]_  | \new_[1963]_ ;
  assign \new_[3726]_  = \new_[1959]_  | \new_[1960]_ ;
  assign \new_[3727]_  = \new_[1961]_  | \new_[3726]_ ;
  assign \new_[3728]_  = \new_[3727]_  | \new_[3722]_ ;
  assign \new_[3731]_  = \new_[1957]_  | \new_[1958]_ ;
  assign \new_[3735]_  = \new_[1954]_  | \new_[1955]_ ;
  assign \new_[3736]_  = \new_[1956]_  | \new_[3735]_ ;
  assign \new_[3737]_  = \new_[3736]_  | \new_[3731]_ ;
  assign \new_[3738]_  = \new_[3737]_  | \new_[3728]_ ;
  assign \new_[3739]_  = \new_[3738]_  | \new_[3719]_ ;
  assign \new_[3740]_  = \new_[3739]_  | \new_[3700]_ ;
  assign \new_[3743]_  = \new_[1952]_  | \new_[1953]_ ;
  assign \new_[3747]_  = \new_[1949]_  | \new_[1950]_ ;
  assign \new_[3748]_  = \new_[1951]_  | \new_[3747]_ ;
  assign \new_[3749]_  = \new_[3748]_  | \new_[3743]_ ;
  assign \new_[3752]_  = \new_[1947]_  | \new_[1948]_ ;
  assign \new_[3756]_  = \new_[1944]_  | \new_[1945]_ ;
  assign \new_[3757]_  = \new_[1946]_  | \new_[3756]_ ;
  assign \new_[3758]_  = \new_[3757]_  | \new_[3752]_ ;
  assign \new_[3759]_  = \new_[3758]_  | \new_[3749]_ ;
  assign \new_[3762]_  = \new_[1942]_  | \new_[1943]_ ;
  assign \new_[3766]_  = \new_[1939]_  | \new_[1940]_ ;
  assign \new_[3767]_  = \new_[1941]_  | \new_[3766]_ ;
  assign \new_[3768]_  = \new_[3767]_  | \new_[3762]_ ;
  assign \new_[3771]_  = \new_[1937]_  | \new_[1938]_ ;
  assign \new_[3775]_  = \new_[1934]_  | \new_[1935]_ ;
  assign \new_[3776]_  = \new_[1936]_  | \new_[3775]_ ;
  assign \new_[3777]_  = \new_[3776]_  | \new_[3771]_ ;
  assign \new_[3778]_  = \new_[3777]_  | \new_[3768]_ ;
  assign \new_[3779]_  = \new_[3778]_  | \new_[3759]_ ;
  assign \new_[3782]_  = \new_[1932]_  | \new_[1933]_ ;
  assign \new_[3786]_  = \new_[1929]_  | \new_[1930]_ ;
  assign \new_[3787]_  = \new_[1931]_  | \new_[3786]_ ;
  assign \new_[3788]_  = \new_[3787]_  | \new_[3782]_ ;
  assign \new_[3791]_  = \new_[1927]_  | \new_[1928]_ ;
  assign \new_[3795]_  = \new_[1924]_  | \new_[1925]_ ;
  assign \new_[3796]_  = \new_[1926]_  | \new_[3795]_ ;
  assign \new_[3797]_  = \new_[3796]_  | \new_[3791]_ ;
  assign \new_[3798]_  = \new_[3797]_  | \new_[3788]_ ;
  assign \new_[3801]_  = \new_[1922]_  | \new_[1923]_ ;
  assign \new_[3805]_  = \new_[1919]_  | \new_[1920]_ ;
  assign \new_[3806]_  = \new_[1921]_  | \new_[3805]_ ;
  assign \new_[3807]_  = \new_[3806]_  | \new_[3801]_ ;
  assign \new_[3810]_  = \new_[1917]_  | \new_[1918]_ ;
  assign \new_[3814]_  = \new_[1914]_  | \new_[1915]_ ;
  assign \new_[3815]_  = \new_[1916]_  | \new_[3814]_ ;
  assign \new_[3816]_  = \new_[3815]_  | \new_[3810]_ ;
  assign \new_[3817]_  = \new_[3816]_  | \new_[3807]_ ;
  assign \new_[3818]_  = \new_[3817]_  | \new_[3798]_ ;
  assign \new_[3819]_  = \new_[3818]_  | \new_[3779]_ ;
  assign \new_[3820]_  = \new_[3819]_  | \new_[3740]_ ;
  assign \new_[3821]_  = \new_[3820]_  | \new_[3661]_ ;
  assign \new_[3822]_  = \new_[3821]_  | \new_[3502]_ ;
  assign \new_[3823]_  = \new_[3822]_  | \new_[3185]_ ;
  assign \new_[3826]_  = \new_[1912]_  | \new_[1913]_ ;
  assign \new_[3829]_  = \new_[1910]_  | \new_[1911]_ ;
  assign \new_[3830]_  = \new_[3829]_  | \new_[3826]_ ;
  assign \new_[3833]_  = \new_[1908]_  | \new_[1909]_ ;
  assign \new_[3837]_  = \new_[1905]_  | \new_[1906]_ ;
  assign \new_[3838]_  = \new_[1907]_  | \new_[3837]_ ;
  assign \new_[3839]_  = \new_[3838]_  | \new_[3833]_ ;
  assign \new_[3840]_  = \new_[3839]_  | \new_[3830]_ ;
  assign \new_[3843]_  = \new_[1903]_  | \new_[1904]_ ;
  assign \new_[3847]_  = \new_[1900]_  | \new_[1901]_ ;
  assign \new_[3848]_  = \new_[1902]_  | \new_[3847]_ ;
  assign \new_[3849]_  = \new_[3848]_  | \new_[3843]_ ;
  assign \new_[3852]_  = \new_[1898]_  | \new_[1899]_ ;
  assign \new_[3856]_  = \new_[1895]_  | \new_[1896]_ ;
  assign \new_[3857]_  = \new_[1897]_  | \new_[3856]_ ;
  assign \new_[3858]_  = \new_[3857]_  | \new_[3852]_ ;
  assign \new_[3859]_  = \new_[3858]_  | \new_[3849]_ ;
  assign \new_[3860]_  = \new_[3859]_  | \new_[3840]_ ;
  assign \new_[3863]_  = \new_[1893]_  | \new_[1894]_ ;
  assign \new_[3867]_  = \new_[1890]_  | \new_[1891]_ ;
  assign \new_[3868]_  = \new_[1892]_  | \new_[3867]_ ;
  assign \new_[3869]_  = \new_[3868]_  | \new_[3863]_ ;
  assign \new_[3872]_  = \new_[1888]_  | \new_[1889]_ ;
  assign \new_[3876]_  = \new_[1885]_  | \new_[1886]_ ;
  assign \new_[3877]_  = \new_[1887]_  | \new_[3876]_ ;
  assign \new_[3878]_  = \new_[3877]_  | \new_[3872]_ ;
  assign \new_[3879]_  = \new_[3878]_  | \new_[3869]_ ;
  assign \new_[3882]_  = \new_[1883]_  | \new_[1884]_ ;
  assign \new_[3886]_  = \new_[1880]_  | \new_[1881]_ ;
  assign \new_[3887]_  = \new_[1882]_  | \new_[3886]_ ;
  assign \new_[3888]_  = \new_[3887]_  | \new_[3882]_ ;
  assign \new_[3891]_  = \new_[1878]_  | \new_[1879]_ ;
  assign \new_[3895]_  = \new_[1875]_  | \new_[1876]_ ;
  assign \new_[3896]_  = \new_[1877]_  | \new_[3895]_ ;
  assign \new_[3897]_  = \new_[3896]_  | \new_[3891]_ ;
  assign \new_[3898]_  = \new_[3897]_  | \new_[3888]_ ;
  assign \new_[3899]_  = \new_[3898]_  | \new_[3879]_ ;
  assign \new_[3900]_  = \new_[3899]_  | \new_[3860]_ ;
  assign \new_[3903]_  = \new_[1873]_  | \new_[1874]_ ;
  assign \new_[3907]_  = \new_[1870]_  | \new_[1871]_ ;
  assign \new_[3908]_  = \new_[1872]_  | \new_[3907]_ ;
  assign \new_[3909]_  = \new_[3908]_  | \new_[3903]_ ;
  assign \new_[3912]_  = \new_[1868]_  | \new_[1869]_ ;
  assign \new_[3916]_  = \new_[1865]_  | \new_[1866]_ ;
  assign \new_[3917]_  = \new_[1867]_  | \new_[3916]_ ;
  assign \new_[3918]_  = \new_[3917]_  | \new_[3912]_ ;
  assign \new_[3919]_  = \new_[3918]_  | \new_[3909]_ ;
  assign \new_[3922]_  = \new_[1863]_  | \new_[1864]_ ;
  assign \new_[3926]_  = \new_[1860]_  | \new_[1861]_ ;
  assign \new_[3927]_  = \new_[1862]_  | \new_[3926]_ ;
  assign \new_[3928]_  = \new_[3927]_  | \new_[3922]_ ;
  assign \new_[3931]_  = \new_[1858]_  | \new_[1859]_ ;
  assign \new_[3935]_  = \new_[1855]_  | \new_[1856]_ ;
  assign \new_[3936]_  = \new_[1857]_  | \new_[3935]_ ;
  assign \new_[3937]_  = \new_[3936]_  | \new_[3931]_ ;
  assign \new_[3938]_  = \new_[3937]_  | \new_[3928]_ ;
  assign \new_[3939]_  = \new_[3938]_  | \new_[3919]_ ;
  assign \new_[3942]_  = \new_[1853]_  | \new_[1854]_ ;
  assign \new_[3946]_  = \new_[1850]_  | \new_[1851]_ ;
  assign \new_[3947]_  = \new_[1852]_  | \new_[3946]_ ;
  assign \new_[3948]_  = \new_[3947]_  | \new_[3942]_ ;
  assign \new_[3951]_  = \new_[1848]_  | \new_[1849]_ ;
  assign \new_[3955]_  = \new_[1845]_  | \new_[1846]_ ;
  assign \new_[3956]_  = \new_[1847]_  | \new_[3955]_ ;
  assign \new_[3957]_  = \new_[3956]_  | \new_[3951]_ ;
  assign \new_[3958]_  = \new_[3957]_  | \new_[3948]_ ;
  assign \new_[3961]_  = \new_[1843]_  | \new_[1844]_ ;
  assign \new_[3965]_  = \new_[1840]_  | \new_[1841]_ ;
  assign \new_[3966]_  = \new_[1842]_  | \new_[3965]_ ;
  assign \new_[3967]_  = \new_[3966]_  | \new_[3961]_ ;
  assign \new_[3970]_  = \new_[1838]_  | \new_[1839]_ ;
  assign \new_[3974]_  = \new_[1835]_  | \new_[1836]_ ;
  assign \new_[3975]_  = \new_[1837]_  | \new_[3974]_ ;
  assign \new_[3976]_  = \new_[3975]_  | \new_[3970]_ ;
  assign \new_[3977]_  = \new_[3976]_  | \new_[3967]_ ;
  assign \new_[3978]_  = \new_[3977]_  | \new_[3958]_ ;
  assign \new_[3979]_  = \new_[3978]_  | \new_[3939]_ ;
  assign \new_[3980]_  = \new_[3979]_  | \new_[3900]_ ;
  assign \new_[3983]_  = \new_[1833]_  | \new_[1834]_ ;
  assign \new_[3987]_  = \new_[1830]_  | \new_[1831]_ ;
  assign \new_[3988]_  = \new_[1832]_  | \new_[3987]_ ;
  assign \new_[3989]_  = \new_[3988]_  | \new_[3983]_ ;
  assign \new_[3992]_  = \new_[1828]_  | \new_[1829]_ ;
  assign \new_[3996]_  = \new_[1825]_  | \new_[1826]_ ;
  assign \new_[3997]_  = \new_[1827]_  | \new_[3996]_ ;
  assign \new_[3998]_  = \new_[3997]_  | \new_[3992]_ ;
  assign \new_[3999]_  = \new_[3998]_  | \new_[3989]_ ;
  assign \new_[4002]_  = \new_[1823]_  | \new_[1824]_ ;
  assign \new_[4006]_  = \new_[1820]_  | \new_[1821]_ ;
  assign \new_[4007]_  = \new_[1822]_  | \new_[4006]_ ;
  assign \new_[4008]_  = \new_[4007]_  | \new_[4002]_ ;
  assign \new_[4011]_  = \new_[1818]_  | \new_[1819]_ ;
  assign \new_[4015]_  = \new_[1815]_  | \new_[1816]_ ;
  assign \new_[4016]_  = \new_[1817]_  | \new_[4015]_ ;
  assign \new_[4017]_  = \new_[4016]_  | \new_[4011]_ ;
  assign \new_[4018]_  = \new_[4017]_  | \new_[4008]_ ;
  assign \new_[4019]_  = \new_[4018]_  | \new_[3999]_ ;
  assign \new_[4022]_  = \new_[1813]_  | \new_[1814]_ ;
  assign \new_[4026]_  = \new_[1810]_  | \new_[1811]_ ;
  assign \new_[4027]_  = \new_[1812]_  | \new_[4026]_ ;
  assign \new_[4028]_  = \new_[4027]_  | \new_[4022]_ ;
  assign \new_[4031]_  = \new_[1808]_  | \new_[1809]_ ;
  assign \new_[4035]_  = \new_[1805]_  | \new_[1806]_ ;
  assign \new_[4036]_  = \new_[1807]_  | \new_[4035]_ ;
  assign \new_[4037]_  = \new_[4036]_  | \new_[4031]_ ;
  assign \new_[4038]_  = \new_[4037]_  | \new_[4028]_ ;
  assign \new_[4041]_  = \new_[1803]_  | \new_[1804]_ ;
  assign \new_[4045]_  = \new_[1800]_  | \new_[1801]_ ;
  assign \new_[4046]_  = \new_[1802]_  | \new_[4045]_ ;
  assign \new_[4047]_  = \new_[4046]_  | \new_[4041]_ ;
  assign \new_[4050]_  = \new_[1798]_  | \new_[1799]_ ;
  assign \new_[4054]_  = \new_[1795]_  | \new_[1796]_ ;
  assign \new_[4055]_  = \new_[1797]_  | \new_[4054]_ ;
  assign \new_[4056]_  = \new_[4055]_  | \new_[4050]_ ;
  assign \new_[4057]_  = \new_[4056]_  | \new_[4047]_ ;
  assign \new_[4058]_  = \new_[4057]_  | \new_[4038]_ ;
  assign \new_[4059]_  = \new_[4058]_  | \new_[4019]_ ;
  assign \new_[4062]_  = \new_[1793]_  | \new_[1794]_ ;
  assign \new_[4066]_  = \new_[1790]_  | \new_[1791]_ ;
  assign \new_[4067]_  = \new_[1792]_  | \new_[4066]_ ;
  assign \new_[4068]_  = \new_[4067]_  | \new_[4062]_ ;
  assign \new_[4071]_  = \new_[1788]_  | \new_[1789]_ ;
  assign \new_[4075]_  = \new_[1785]_  | \new_[1786]_ ;
  assign \new_[4076]_  = \new_[1787]_  | \new_[4075]_ ;
  assign \new_[4077]_  = \new_[4076]_  | \new_[4071]_ ;
  assign \new_[4078]_  = \new_[4077]_  | \new_[4068]_ ;
  assign \new_[4081]_  = \new_[1783]_  | \new_[1784]_ ;
  assign \new_[4085]_  = \new_[1780]_  | \new_[1781]_ ;
  assign \new_[4086]_  = \new_[1782]_  | \new_[4085]_ ;
  assign \new_[4087]_  = \new_[4086]_  | \new_[4081]_ ;
  assign \new_[4090]_  = \new_[1778]_  | \new_[1779]_ ;
  assign \new_[4094]_  = \new_[1775]_  | \new_[1776]_ ;
  assign \new_[4095]_  = \new_[1777]_  | \new_[4094]_ ;
  assign \new_[4096]_  = \new_[4095]_  | \new_[4090]_ ;
  assign \new_[4097]_  = \new_[4096]_  | \new_[4087]_ ;
  assign \new_[4098]_  = \new_[4097]_  | \new_[4078]_ ;
  assign \new_[4101]_  = \new_[1773]_  | \new_[1774]_ ;
  assign \new_[4105]_  = \new_[1770]_  | \new_[1771]_ ;
  assign \new_[4106]_  = \new_[1772]_  | \new_[4105]_ ;
  assign \new_[4107]_  = \new_[4106]_  | \new_[4101]_ ;
  assign \new_[4110]_  = \new_[1768]_  | \new_[1769]_ ;
  assign \new_[4114]_  = \new_[1765]_  | \new_[1766]_ ;
  assign \new_[4115]_  = \new_[1767]_  | \new_[4114]_ ;
  assign \new_[4116]_  = \new_[4115]_  | \new_[4110]_ ;
  assign \new_[4117]_  = \new_[4116]_  | \new_[4107]_ ;
  assign \new_[4120]_  = \new_[1763]_  | \new_[1764]_ ;
  assign \new_[4124]_  = \new_[1760]_  | \new_[1761]_ ;
  assign \new_[4125]_  = \new_[1762]_  | \new_[4124]_ ;
  assign \new_[4126]_  = \new_[4125]_  | \new_[4120]_ ;
  assign \new_[4129]_  = \new_[1758]_  | \new_[1759]_ ;
  assign \new_[4133]_  = \new_[1755]_  | \new_[1756]_ ;
  assign \new_[4134]_  = \new_[1757]_  | \new_[4133]_ ;
  assign \new_[4135]_  = \new_[4134]_  | \new_[4129]_ ;
  assign \new_[4136]_  = \new_[4135]_  | \new_[4126]_ ;
  assign \new_[4137]_  = \new_[4136]_  | \new_[4117]_ ;
  assign \new_[4138]_  = \new_[4137]_  | \new_[4098]_ ;
  assign \new_[4139]_  = \new_[4138]_  | \new_[4059]_ ;
  assign \new_[4140]_  = \new_[4139]_  | \new_[3980]_ ;
  assign \new_[4143]_  = \new_[1753]_  | \new_[1754]_ ;
  assign \new_[4147]_  = \new_[1750]_  | \new_[1751]_ ;
  assign \new_[4148]_  = \new_[1752]_  | \new_[4147]_ ;
  assign \new_[4149]_  = \new_[4148]_  | \new_[4143]_ ;
  assign \new_[4152]_  = \new_[1748]_  | \new_[1749]_ ;
  assign \new_[4156]_  = \new_[1745]_  | \new_[1746]_ ;
  assign \new_[4157]_  = \new_[1747]_  | \new_[4156]_ ;
  assign \new_[4158]_  = \new_[4157]_  | \new_[4152]_ ;
  assign \new_[4159]_  = \new_[4158]_  | \new_[4149]_ ;
  assign \new_[4162]_  = \new_[1743]_  | \new_[1744]_ ;
  assign \new_[4166]_  = \new_[1740]_  | \new_[1741]_ ;
  assign \new_[4167]_  = \new_[1742]_  | \new_[4166]_ ;
  assign \new_[4168]_  = \new_[4167]_  | \new_[4162]_ ;
  assign \new_[4171]_  = \new_[1738]_  | \new_[1739]_ ;
  assign \new_[4175]_  = \new_[1735]_  | \new_[1736]_ ;
  assign \new_[4176]_  = \new_[1737]_  | \new_[4175]_ ;
  assign \new_[4177]_  = \new_[4176]_  | \new_[4171]_ ;
  assign \new_[4178]_  = \new_[4177]_  | \new_[4168]_ ;
  assign \new_[4179]_  = \new_[4178]_  | \new_[4159]_ ;
  assign \new_[4182]_  = \new_[1733]_  | \new_[1734]_ ;
  assign \new_[4186]_  = \new_[1730]_  | \new_[1731]_ ;
  assign \new_[4187]_  = \new_[1732]_  | \new_[4186]_ ;
  assign \new_[4188]_  = \new_[4187]_  | \new_[4182]_ ;
  assign \new_[4191]_  = \new_[1728]_  | \new_[1729]_ ;
  assign \new_[4195]_  = \new_[1725]_  | \new_[1726]_ ;
  assign \new_[4196]_  = \new_[1727]_  | \new_[4195]_ ;
  assign \new_[4197]_  = \new_[4196]_  | \new_[4191]_ ;
  assign \new_[4198]_  = \new_[4197]_  | \new_[4188]_ ;
  assign \new_[4201]_  = \new_[1723]_  | \new_[1724]_ ;
  assign \new_[4205]_  = \new_[1720]_  | \new_[1721]_ ;
  assign \new_[4206]_  = \new_[1722]_  | \new_[4205]_ ;
  assign \new_[4207]_  = \new_[4206]_  | \new_[4201]_ ;
  assign \new_[4210]_  = \new_[1718]_  | \new_[1719]_ ;
  assign \new_[4214]_  = \new_[1715]_  | \new_[1716]_ ;
  assign \new_[4215]_  = \new_[1717]_  | \new_[4214]_ ;
  assign \new_[4216]_  = \new_[4215]_  | \new_[4210]_ ;
  assign \new_[4217]_  = \new_[4216]_  | \new_[4207]_ ;
  assign \new_[4218]_  = \new_[4217]_  | \new_[4198]_ ;
  assign \new_[4219]_  = \new_[4218]_  | \new_[4179]_ ;
  assign \new_[4222]_  = \new_[1713]_  | \new_[1714]_ ;
  assign \new_[4226]_  = \new_[1710]_  | \new_[1711]_ ;
  assign \new_[4227]_  = \new_[1712]_  | \new_[4226]_ ;
  assign \new_[4228]_  = \new_[4227]_  | \new_[4222]_ ;
  assign \new_[4231]_  = \new_[1708]_  | \new_[1709]_ ;
  assign \new_[4235]_  = \new_[1705]_  | \new_[1706]_ ;
  assign \new_[4236]_  = \new_[1707]_  | \new_[4235]_ ;
  assign \new_[4237]_  = \new_[4236]_  | \new_[4231]_ ;
  assign \new_[4238]_  = \new_[4237]_  | \new_[4228]_ ;
  assign \new_[4241]_  = \new_[1703]_  | \new_[1704]_ ;
  assign \new_[4245]_  = \new_[1700]_  | \new_[1701]_ ;
  assign \new_[4246]_  = \new_[1702]_  | \new_[4245]_ ;
  assign \new_[4247]_  = \new_[4246]_  | \new_[4241]_ ;
  assign \new_[4250]_  = \new_[1698]_  | \new_[1699]_ ;
  assign \new_[4254]_  = \new_[1695]_  | \new_[1696]_ ;
  assign \new_[4255]_  = \new_[1697]_  | \new_[4254]_ ;
  assign \new_[4256]_  = \new_[4255]_  | \new_[4250]_ ;
  assign \new_[4257]_  = \new_[4256]_  | \new_[4247]_ ;
  assign \new_[4258]_  = \new_[4257]_  | \new_[4238]_ ;
  assign \new_[4261]_  = \new_[1693]_  | \new_[1694]_ ;
  assign \new_[4265]_  = \new_[1690]_  | \new_[1691]_ ;
  assign \new_[4266]_  = \new_[1692]_  | \new_[4265]_ ;
  assign \new_[4267]_  = \new_[4266]_  | \new_[4261]_ ;
  assign \new_[4270]_  = \new_[1688]_  | \new_[1689]_ ;
  assign \new_[4274]_  = \new_[1685]_  | \new_[1686]_ ;
  assign \new_[4275]_  = \new_[1687]_  | \new_[4274]_ ;
  assign \new_[4276]_  = \new_[4275]_  | \new_[4270]_ ;
  assign \new_[4277]_  = \new_[4276]_  | \new_[4267]_ ;
  assign \new_[4280]_  = \new_[1683]_  | \new_[1684]_ ;
  assign \new_[4284]_  = \new_[1680]_  | \new_[1681]_ ;
  assign \new_[4285]_  = \new_[1682]_  | \new_[4284]_ ;
  assign \new_[4286]_  = \new_[4285]_  | \new_[4280]_ ;
  assign \new_[4289]_  = \new_[1678]_  | \new_[1679]_ ;
  assign \new_[4293]_  = \new_[1675]_  | \new_[1676]_ ;
  assign \new_[4294]_  = \new_[1677]_  | \new_[4293]_ ;
  assign \new_[4295]_  = \new_[4294]_  | \new_[4289]_ ;
  assign \new_[4296]_  = \new_[4295]_  | \new_[4286]_ ;
  assign \new_[4297]_  = \new_[4296]_  | \new_[4277]_ ;
  assign \new_[4298]_  = \new_[4297]_  | \new_[4258]_ ;
  assign \new_[4299]_  = \new_[4298]_  | \new_[4219]_ ;
  assign \new_[4302]_  = \new_[1673]_  | \new_[1674]_ ;
  assign \new_[4306]_  = \new_[1670]_  | \new_[1671]_ ;
  assign \new_[4307]_  = \new_[1672]_  | \new_[4306]_ ;
  assign \new_[4308]_  = \new_[4307]_  | \new_[4302]_ ;
  assign \new_[4311]_  = \new_[1668]_  | \new_[1669]_ ;
  assign \new_[4315]_  = \new_[1665]_  | \new_[1666]_ ;
  assign \new_[4316]_  = \new_[1667]_  | \new_[4315]_ ;
  assign \new_[4317]_  = \new_[4316]_  | \new_[4311]_ ;
  assign \new_[4318]_  = \new_[4317]_  | \new_[4308]_ ;
  assign \new_[4321]_  = \new_[1663]_  | \new_[1664]_ ;
  assign \new_[4325]_  = \new_[1660]_  | \new_[1661]_ ;
  assign \new_[4326]_  = \new_[1662]_  | \new_[4325]_ ;
  assign \new_[4327]_  = \new_[4326]_  | \new_[4321]_ ;
  assign \new_[4330]_  = \new_[1658]_  | \new_[1659]_ ;
  assign \new_[4334]_  = \new_[1655]_  | \new_[1656]_ ;
  assign \new_[4335]_  = \new_[1657]_  | \new_[4334]_ ;
  assign \new_[4336]_  = \new_[4335]_  | \new_[4330]_ ;
  assign \new_[4337]_  = \new_[4336]_  | \new_[4327]_ ;
  assign \new_[4338]_  = \new_[4337]_  | \new_[4318]_ ;
  assign \new_[4341]_  = \new_[1653]_  | \new_[1654]_ ;
  assign \new_[4345]_  = \new_[1650]_  | \new_[1651]_ ;
  assign \new_[4346]_  = \new_[1652]_  | \new_[4345]_ ;
  assign \new_[4347]_  = \new_[4346]_  | \new_[4341]_ ;
  assign \new_[4350]_  = \new_[1648]_  | \new_[1649]_ ;
  assign \new_[4354]_  = \new_[1645]_  | \new_[1646]_ ;
  assign \new_[4355]_  = \new_[1647]_  | \new_[4354]_ ;
  assign \new_[4356]_  = \new_[4355]_  | \new_[4350]_ ;
  assign \new_[4357]_  = \new_[4356]_  | \new_[4347]_ ;
  assign \new_[4360]_  = \new_[1643]_  | \new_[1644]_ ;
  assign \new_[4364]_  = \new_[1640]_  | \new_[1641]_ ;
  assign \new_[4365]_  = \new_[1642]_  | \new_[4364]_ ;
  assign \new_[4366]_  = \new_[4365]_  | \new_[4360]_ ;
  assign \new_[4369]_  = \new_[1638]_  | \new_[1639]_ ;
  assign \new_[4373]_  = \new_[1635]_  | \new_[1636]_ ;
  assign \new_[4374]_  = \new_[1637]_  | \new_[4373]_ ;
  assign \new_[4375]_  = \new_[4374]_  | \new_[4369]_ ;
  assign \new_[4376]_  = \new_[4375]_  | \new_[4366]_ ;
  assign \new_[4377]_  = \new_[4376]_  | \new_[4357]_ ;
  assign \new_[4378]_  = \new_[4377]_  | \new_[4338]_ ;
  assign \new_[4381]_  = \new_[1633]_  | \new_[1634]_ ;
  assign \new_[4385]_  = \new_[1630]_  | \new_[1631]_ ;
  assign \new_[4386]_  = \new_[1632]_  | \new_[4385]_ ;
  assign \new_[4387]_  = \new_[4386]_  | \new_[4381]_ ;
  assign \new_[4390]_  = \new_[1628]_  | \new_[1629]_ ;
  assign \new_[4394]_  = \new_[1625]_  | \new_[1626]_ ;
  assign \new_[4395]_  = \new_[1627]_  | \new_[4394]_ ;
  assign \new_[4396]_  = \new_[4395]_  | \new_[4390]_ ;
  assign \new_[4397]_  = \new_[4396]_  | \new_[4387]_ ;
  assign \new_[4400]_  = \new_[1623]_  | \new_[1624]_ ;
  assign \new_[4404]_  = \new_[1620]_  | \new_[1621]_ ;
  assign \new_[4405]_  = \new_[1622]_  | \new_[4404]_ ;
  assign \new_[4406]_  = \new_[4405]_  | \new_[4400]_ ;
  assign \new_[4409]_  = \new_[1618]_  | \new_[1619]_ ;
  assign \new_[4413]_  = \new_[1615]_  | \new_[1616]_ ;
  assign \new_[4414]_  = \new_[1617]_  | \new_[4413]_ ;
  assign \new_[4415]_  = \new_[4414]_  | \new_[4409]_ ;
  assign \new_[4416]_  = \new_[4415]_  | \new_[4406]_ ;
  assign \new_[4417]_  = \new_[4416]_  | \new_[4397]_ ;
  assign \new_[4420]_  = \new_[1613]_  | \new_[1614]_ ;
  assign \new_[4424]_  = \new_[1610]_  | \new_[1611]_ ;
  assign \new_[4425]_  = \new_[1612]_  | \new_[4424]_ ;
  assign \new_[4426]_  = \new_[4425]_  | \new_[4420]_ ;
  assign \new_[4429]_  = \new_[1608]_  | \new_[1609]_ ;
  assign \new_[4433]_  = \new_[1605]_  | \new_[1606]_ ;
  assign \new_[4434]_  = \new_[1607]_  | \new_[4433]_ ;
  assign \new_[4435]_  = \new_[4434]_  | \new_[4429]_ ;
  assign \new_[4436]_  = \new_[4435]_  | \new_[4426]_ ;
  assign \new_[4439]_  = \new_[1603]_  | \new_[1604]_ ;
  assign \new_[4443]_  = \new_[1600]_  | \new_[1601]_ ;
  assign \new_[4444]_  = \new_[1602]_  | \new_[4443]_ ;
  assign \new_[4445]_  = \new_[4444]_  | \new_[4439]_ ;
  assign \new_[4448]_  = \new_[1598]_  | \new_[1599]_ ;
  assign \new_[4452]_  = \new_[1595]_  | \new_[1596]_ ;
  assign \new_[4453]_  = \new_[1597]_  | \new_[4452]_ ;
  assign \new_[4454]_  = \new_[4453]_  | \new_[4448]_ ;
  assign \new_[4455]_  = \new_[4454]_  | \new_[4445]_ ;
  assign \new_[4456]_  = \new_[4455]_  | \new_[4436]_ ;
  assign \new_[4457]_  = \new_[4456]_  | \new_[4417]_ ;
  assign \new_[4458]_  = \new_[4457]_  | \new_[4378]_ ;
  assign \new_[4459]_  = \new_[4458]_  | \new_[4299]_ ;
  assign \new_[4460]_  = \new_[4459]_  | \new_[4140]_ ;
  assign \new_[4463]_  = \new_[1593]_  | \new_[1594]_ ;
  assign \new_[4466]_  = \new_[1591]_  | \new_[1592]_ ;
  assign \new_[4467]_  = \new_[4466]_  | \new_[4463]_ ;
  assign \new_[4470]_  = \new_[1589]_  | \new_[1590]_ ;
  assign \new_[4474]_  = \new_[1586]_  | \new_[1587]_ ;
  assign \new_[4475]_  = \new_[1588]_  | \new_[4474]_ ;
  assign \new_[4476]_  = \new_[4475]_  | \new_[4470]_ ;
  assign \new_[4477]_  = \new_[4476]_  | \new_[4467]_ ;
  assign \new_[4480]_  = \new_[1584]_  | \new_[1585]_ ;
  assign \new_[4484]_  = \new_[1581]_  | \new_[1582]_ ;
  assign \new_[4485]_  = \new_[1583]_  | \new_[4484]_ ;
  assign \new_[4486]_  = \new_[4485]_  | \new_[4480]_ ;
  assign \new_[4489]_  = \new_[1579]_  | \new_[1580]_ ;
  assign \new_[4493]_  = \new_[1576]_  | \new_[1577]_ ;
  assign \new_[4494]_  = \new_[1578]_  | \new_[4493]_ ;
  assign \new_[4495]_  = \new_[4494]_  | \new_[4489]_ ;
  assign \new_[4496]_  = \new_[4495]_  | \new_[4486]_ ;
  assign \new_[4497]_  = \new_[4496]_  | \new_[4477]_ ;
  assign \new_[4500]_  = \new_[1574]_  | \new_[1575]_ ;
  assign \new_[4504]_  = \new_[1571]_  | \new_[1572]_ ;
  assign \new_[4505]_  = \new_[1573]_  | \new_[4504]_ ;
  assign \new_[4506]_  = \new_[4505]_  | \new_[4500]_ ;
  assign \new_[4509]_  = \new_[1569]_  | \new_[1570]_ ;
  assign \new_[4513]_  = \new_[1566]_  | \new_[1567]_ ;
  assign \new_[4514]_  = \new_[1568]_  | \new_[4513]_ ;
  assign \new_[4515]_  = \new_[4514]_  | \new_[4509]_ ;
  assign \new_[4516]_  = \new_[4515]_  | \new_[4506]_ ;
  assign \new_[4519]_  = \new_[1564]_  | \new_[1565]_ ;
  assign \new_[4523]_  = \new_[1561]_  | \new_[1562]_ ;
  assign \new_[4524]_  = \new_[1563]_  | \new_[4523]_ ;
  assign \new_[4525]_  = \new_[4524]_  | \new_[4519]_ ;
  assign \new_[4528]_  = \new_[1559]_  | \new_[1560]_ ;
  assign \new_[4532]_  = \new_[1556]_  | \new_[1557]_ ;
  assign \new_[4533]_  = \new_[1558]_  | \new_[4532]_ ;
  assign \new_[4534]_  = \new_[4533]_  | \new_[4528]_ ;
  assign \new_[4535]_  = \new_[4534]_  | \new_[4525]_ ;
  assign \new_[4536]_  = \new_[4535]_  | \new_[4516]_ ;
  assign \new_[4537]_  = \new_[4536]_  | \new_[4497]_ ;
  assign \new_[4540]_  = \new_[1554]_  | \new_[1555]_ ;
  assign \new_[4544]_  = \new_[1551]_  | \new_[1552]_ ;
  assign \new_[4545]_  = \new_[1553]_  | \new_[4544]_ ;
  assign \new_[4546]_  = \new_[4545]_  | \new_[4540]_ ;
  assign \new_[4549]_  = \new_[1549]_  | \new_[1550]_ ;
  assign \new_[4553]_  = \new_[1546]_  | \new_[1547]_ ;
  assign \new_[4554]_  = \new_[1548]_  | \new_[4553]_ ;
  assign \new_[4555]_  = \new_[4554]_  | \new_[4549]_ ;
  assign \new_[4556]_  = \new_[4555]_  | \new_[4546]_ ;
  assign \new_[4559]_  = \new_[1544]_  | \new_[1545]_ ;
  assign \new_[4563]_  = \new_[1541]_  | \new_[1542]_ ;
  assign \new_[4564]_  = \new_[1543]_  | \new_[4563]_ ;
  assign \new_[4565]_  = \new_[4564]_  | \new_[4559]_ ;
  assign \new_[4568]_  = \new_[1539]_  | \new_[1540]_ ;
  assign \new_[4572]_  = \new_[1536]_  | \new_[1537]_ ;
  assign \new_[4573]_  = \new_[1538]_  | \new_[4572]_ ;
  assign \new_[4574]_  = \new_[4573]_  | \new_[4568]_ ;
  assign \new_[4575]_  = \new_[4574]_  | \new_[4565]_ ;
  assign \new_[4576]_  = \new_[4575]_  | \new_[4556]_ ;
  assign \new_[4579]_  = \new_[1534]_  | \new_[1535]_ ;
  assign \new_[4583]_  = \new_[1531]_  | \new_[1532]_ ;
  assign \new_[4584]_  = \new_[1533]_  | \new_[4583]_ ;
  assign \new_[4585]_  = \new_[4584]_  | \new_[4579]_ ;
  assign \new_[4588]_  = \new_[1529]_  | \new_[1530]_ ;
  assign \new_[4592]_  = \new_[1526]_  | \new_[1527]_ ;
  assign \new_[4593]_  = \new_[1528]_  | \new_[4592]_ ;
  assign \new_[4594]_  = \new_[4593]_  | \new_[4588]_ ;
  assign \new_[4595]_  = \new_[4594]_  | \new_[4585]_ ;
  assign \new_[4598]_  = \new_[1524]_  | \new_[1525]_ ;
  assign \new_[4602]_  = \new_[1521]_  | \new_[1522]_ ;
  assign \new_[4603]_  = \new_[1523]_  | \new_[4602]_ ;
  assign \new_[4604]_  = \new_[4603]_  | \new_[4598]_ ;
  assign \new_[4607]_  = \new_[1519]_  | \new_[1520]_ ;
  assign \new_[4611]_  = \new_[1516]_  | \new_[1517]_ ;
  assign \new_[4612]_  = \new_[1518]_  | \new_[4611]_ ;
  assign \new_[4613]_  = \new_[4612]_  | \new_[4607]_ ;
  assign \new_[4614]_  = \new_[4613]_  | \new_[4604]_ ;
  assign \new_[4615]_  = \new_[4614]_  | \new_[4595]_ ;
  assign \new_[4616]_  = \new_[4615]_  | \new_[4576]_ ;
  assign \new_[4617]_  = \new_[4616]_  | \new_[4537]_ ;
  assign \new_[4620]_  = \new_[1514]_  | \new_[1515]_ ;
  assign \new_[4624]_  = \new_[1511]_  | \new_[1512]_ ;
  assign \new_[4625]_  = \new_[1513]_  | \new_[4624]_ ;
  assign \new_[4626]_  = \new_[4625]_  | \new_[4620]_ ;
  assign \new_[4629]_  = \new_[1509]_  | \new_[1510]_ ;
  assign \new_[4633]_  = \new_[1506]_  | \new_[1507]_ ;
  assign \new_[4634]_  = \new_[1508]_  | \new_[4633]_ ;
  assign \new_[4635]_  = \new_[4634]_  | \new_[4629]_ ;
  assign \new_[4636]_  = \new_[4635]_  | \new_[4626]_ ;
  assign \new_[4639]_  = \new_[1504]_  | \new_[1505]_ ;
  assign \new_[4643]_  = \new_[1501]_  | \new_[1502]_ ;
  assign \new_[4644]_  = \new_[1503]_  | \new_[4643]_ ;
  assign \new_[4645]_  = \new_[4644]_  | \new_[4639]_ ;
  assign \new_[4648]_  = \new_[1499]_  | \new_[1500]_ ;
  assign \new_[4652]_  = \new_[1496]_  | \new_[1497]_ ;
  assign \new_[4653]_  = \new_[1498]_  | \new_[4652]_ ;
  assign \new_[4654]_  = \new_[4653]_  | \new_[4648]_ ;
  assign \new_[4655]_  = \new_[4654]_  | \new_[4645]_ ;
  assign \new_[4656]_  = \new_[4655]_  | \new_[4636]_ ;
  assign \new_[4659]_  = \new_[1494]_  | \new_[1495]_ ;
  assign \new_[4663]_  = \new_[1491]_  | \new_[1492]_ ;
  assign \new_[4664]_  = \new_[1493]_  | \new_[4663]_ ;
  assign \new_[4665]_  = \new_[4664]_  | \new_[4659]_ ;
  assign \new_[4668]_  = \new_[1489]_  | \new_[1490]_ ;
  assign \new_[4672]_  = \new_[1486]_  | \new_[1487]_ ;
  assign \new_[4673]_  = \new_[1488]_  | \new_[4672]_ ;
  assign \new_[4674]_  = \new_[4673]_  | \new_[4668]_ ;
  assign \new_[4675]_  = \new_[4674]_  | \new_[4665]_ ;
  assign \new_[4678]_  = \new_[1484]_  | \new_[1485]_ ;
  assign \new_[4682]_  = \new_[1481]_  | \new_[1482]_ ;
  assign \new_[4683]_  = \new_[1483]_  | \new_[4682]_ ;
  assign \new_[4684]_  = \new_[4683]_  | \new_[4678]_ ;
  assign \new_[4687]_  = \new_[1479]_  | \new_[1480]_ ;
  assign \new_[4691]_  = \new_[1476]_  | \new_[1477]_ ;
  assign \new_[4692]_  = \new_[1478]_  | \new_[4691]_ ;
  assign \new_[4693]_  = \new_[4692]_  | \new_[4687]_ ;
  assign \new_[4694]_  = \new_[4693]_  | \new_[4684]_ ;
  assign \new_[4695]_  = \new_[4694]_  | \new_[4675]_ ;
  assign \new_[4696]_  = \new_[4695]_  | \new_[4656]_ ;
  assign \new_[4699]_  = \new_[1474]_  | \new_[1475]_ ;
  assign \new_[4703]_  = \new_[1471]_  | \new_[1472]_ ;
  assign \new_[4704]_  = \new_[1473]_  | \new_[4703]_ ;
  assign \new_[4705]_  = \new_[4704]_  | \new_[4699]_ ;
  assign \new_[4708]_  = \new_[1469]_  | \new_[1470]_ ;
  assign \new_[4712]_  = \new_[1466]_  | \new_[1467]_ ;
  assign \new_[4713]_  = \new_[1468]_  | \new_[4712]_ ;
  assign \new_[4714]_  = \new_[4713]_  | \new_[4708]_ ;
  assign \new_[4715]_  = \new_[4714]_  | \new_[4705]_ ;
  assign \new_[4718]_  = \new_[1464]_  | \new_[1465]_ ;
  assign \new_[4722]_  = \new_[1461]_  | \new_[1462]_ ;
  assign \new_[4723]_  = \new_[1463]_  | \new_[4722]_ ;
  assign \new_[4724]_  = \new_[4723]_  | \new_[4718]_ ;
  assign \new_[4727]_  = \new_[1459]_  | \new_[1460]_ ;
  assign \new_[4731]_  = \new_[1456]_  | \new_[1457]_ ;
  assign \new_[4732]_  = \new_[1458]_  | \new_[4731]_ ;
  assign \new_[4733]_  = \new_[4732]_  | \new_[4727]_ ;
  assign \new_[4734]_  = \new_[4733]_  | \new_[4724]_ ;
  assign \new_[4735]_  = \new_[4734]_  | \new_[4715]_ ;
  assign \new_[4738]_  = \new_[1454]_  | \new_[1455]_ ;
  assign \new_[4742]_  = \new_[1451]_  | \new_[1452]_ ;
  assign \new_[4743]_  = \new_[1453]_  | \new_[4742]_ ;
  assign \new_[4744]_  = \new_[4743]_  | \new_[4738]_ ;
  assign \new_[4747]_  = \new_[1449]_  | \new_[1450]_ ;
  assign \new_[4751]_  = \new_[1446]_  | \new_[1447]_ ;
  assign \new_[4752]_  = \new_[1448]_  | \new_[4751]_ ;
  assign \new_[4753]_  = \new_[4752]_  | \new_[4747]_ ;
  assign \new_[4754]_  = \new_[4753]_  | \new_[4744]_ ;
  assign \new_[4757]_  = \new_[1444]_  | \new_[1445]_ ;
  assign \new_[4761]_  = \new_[1441]_  | \new_[1442]_ ;
  assign \new_[4762]_  = \new_[1443]_  | \new_[4761]_ ;
  assign \new_[4763]_  = \new_[4762]_  | \new_[4757]_ ;
  assign \new_[4766]_  = \new_[1439]_  | \new_[1440]_ ;
  assign \new_[4770]_  = \new_[1436]_  | \new_[1437]_ ;
  assign \new_[4771]_  = \new_[1438]_  | \new_[4770]_ ;
  assign \new_[4772]_  = \new_[4771]_  | \new_[4766]_ ;
  assign \new_[4773]_  = \new_[4772]_  | \new_[4763]_ ;
  assign \new_[4774]_  = \new_[4773]_  | \new_[4754]_ ;
  assign \new_[4775]_  = \new_[4774]_  | \new_[4735]_ ;
  assign \new_[4776]_  = \new_[4775]_  | \new_[4696]_ ;
  assign \new_[4777]_  = \new_[4776]_  | \new_[4617]_ ;
  assign \new_[4780]_  = \new_[1434]_  | \new_[1435]_ ;
  assign \new_[4784]_  = \new_[1431]_  | \new_[1432]_ ;
  assign \new_[4785]_  = \new_[1433]_  | \new_[4784]_ ;
  assign \new_[4786]_  = \new_[4785]_  | \new_[4780]_ ;
  assign \new_[4789]_  = \new_[1429]_  | \new_[1430]_ ;
  assign \new_[4793]_  = \new_[1426]_  | \new_[1427]_ ;
  assign \new_[4794]_  = \new_[1428]_  | \new_[4793]_ ;
  assign \new_[4795]_  = \new_[4794]_  | \new_[4789]_ ;
  assign \new_[4796]_  = \new_[4795]_  | \new_[4786]_ ;
  assign \new_[4799]_  = \new_[1424]_  | \new_[1425]_ ;
  assign \new_[4803]_  = \new_[1421]_  | \new_[1422]_ ;
  assign \new_[4804]_  = \new_[1423]_  | \new_[4803]_ ;
  assign \new_[4805]_  = \new_[4804]_  | \new_[4799]_ ;
  assign \new_[4808]_  = \new_[1419]_  | \new_[1420]_ ;
  assign \new_[4812]_  = \new_[1416]_  | \new_[1417]_ ;
  assign \new_[4813]_  = \new_[1418]_  | \new_[4812]_ ;
  assign \new_[4814]_  = \new_[4813]_  | \new_[4808]_ ;
  assign \new_[4815]_  = \new_[4814]_  | \new_[4805]_ ;
  assign \new_[4816]_  = \new_[4815]_  | \new_[4796]_ ;
  assign \new_[4819]_  = \new_[1414]_  | \new_[1415]_ ;
  assign \new_[4823]_  = \new_[1411]_  | \new_[1412]_ ;
  assign \new_[4824]_  = \new_[1413]_  | \new_[4823]_ ;
  assign \new_[4825]_  = \new_[4824]_  | \new_[4819]_ ;
  assign \new_[4828]_  = \new_[1409]_  | \new_[1410]_ ;
  assign \new_[4832]_  = \new_[1406]_  | \new_[1407]_ ;
  assign \new_[4833]_  = \new_[1408]_  | \new_[4832]_ ;
  assign \new_[4834]_  = \new_[4833]_  | \new_[4828]_ ;
  assign \new_[4835]_  = \new_[4834]_  | \new_[4825]_ ;
  assign \new_[4838]_  = \new_[1404]_  | \new_[1405]_ ;
  assign \new_[4842]_  = \new_[1401]_  | \new_[1402]_ ;
  assign \new_[4843]_  = \new_[1403]_  | \new_[4842]_ ;
  assign \new_[4844]_  = \new_[4843]_  | \new_[4838]_ ;
  assign \new_[4847]_  = \new_[1399]_  | \new_[1400]_ ;
  assign \new_[4851]_  = \new_[1396]_  | \new_[1397]_ ;
  assign \new_[4852]_  = \new_[1398]_  | \new_[4851]_ ;
  assign \new_[4853]_  = \new_[4852]_  | \new_[4847]_ ;
  assign \new_[4854]_  = \new_[4853]_  | \new_[4844]_ ;
  assign \new_[4855]_  = \new_[4854]_  | \new_[4835]_ ;
  assign \new_[4856]_  = \new_[4855]_  | \new_[4816]_ ;
  assign \new_[4859]_  = \new_[1394]_  | \new_[1395]_ ;
  assign \new_[4863]_  = \new_[1391]_  | \new_[1392]_ ;
  assign \new_[4864]_  = \new_[1393]_  | \new_[4863]_ ;
  assign \new_[4865]_  = \new_[4864]_  | \new_[4859]_ ;
  assign \new_[4868]_  = \new_[1389]_  | \new_[1390]_ ;
  assign \new_[4872]_  = \new_[1386]_  | \new_[1387]_ ;
  assign \new_[4873]_  = \new_[1388]_  | \new_[4872]_ ;
  assign \new_[4874]_  = \new_[4873]_  | \new_[4868]_ ;
  assign \new_[4875]_  = \new_[4874]_  | \new_[4865]_ ;
  assign \new_[4878]_  = \new_[1384]_  | \new_[1385]_ ;
  assign \new_[4882]_  = \new_[1381]_  | \new_[1382]_ ;
  assign \new_[4883]_  = \new_[1383]_  | \new_[4882]_ ;
  assign \new_[4884]_  = \new_[4883]_  | \new_[4878]_ ;
  assign \new_[4887]_  = \new_[1379]_  | \new_[1380]_ ;
  assign \new_[4891]_  = \new_[1376]_  | \new_[1377]_ ;
  assign \new_[4892]_  = \new_[1378]_  | \new_[4891]_ ;
  assign \new_[4893]_  = \new_[4892]_  | \new_[4887]_ ;
  assign \new_[4894]_  = \new_[4893]_  | \new_[4884]_ ;
  assign \new_[4895]_  = \new_[4894]_  | \new_[4875]_ ;
  assign \new_[4898]_  = \new_[1374]_  | \new_[1375]_ ;
  assign \new_[4902]_  = \new_[1371]_  | \new_[1372]_ ;
  assign \new_[4903]_  = \new_[1373]_  | \new_[4902]_ ;
  assign \new_[4904]_  = \new_[4903]_  | \new_[4898]_ ;
  assign \new_[4907]_  = \new_[1369]_  | \new_[1370]_ ;
  assign \new_[4911]_  = \new_[1366]_  | \new_[1367]_ ;
  assign \new_[4912]_  = \new_[1368]_  | \new_[4911]_ ;
  assign \new_[4913]_  = \new_[4912]_  | \new_[4907]_ ;
  assign \new_[4914]_  = \new_[4913]_  | \new_[4904]_ ;
  assign \new_[4917]_  = \new_[1364]_  | \new_[1365]_ ;
  assign \new_[4921]_  = \new_[1361]_  | \new_[1362]_ ;
  assign \new_[4922]_  = \new_[1363]_  | \new_[4921]_ ;
  assign \new_[4923]_  = \new_[4922]_  | \new_[4917]_ ;
  assign \new_[4926]_  = \new_[1359]_  | \new_[1360]_ ;
  assign \new_[4930]_  = \new_[1356]_  | \new_[1357]_ ;
  assign \new_[4931]_  = \new_[1358]_  | \new_[4930]_ ;
  assign \new_[4932]_  = \new_[4931]_  | \new_[4926]_ ;
  assign \new_[4933]_  = \new_[4932]_  | \new_[4923]_ ;
  assign \new_[4934]_  = \new_[4933]_  | \new_[4914]_ ;
  assign \new_[4935]_  = \new_[4934]_  | \new_[4895]_ ;
  assign \new_[4936]_  = \new_[4935]_  | \new_[4856]_ ;
  assign \new_[4939]_  = \new_[1354]_  | \new_[1355]_ ;
  assign \new_[4943]_  = \new_[1351]_  | \new_[1352]_ ;
  assign \new_[4944]_  = \new_[1353]_  | \new_[4943]_ ;
  assign \new_[4945]_  = \new_[4944]_  | \new_[4939]_ ;
  assign \new_[4948]_  = \new_[1349]_  | \new_[1350]_ ;
  assign \new_[4952]_  = \new_[1346]_  | \new_[1347]_ ;
  assign \new_[4953]_  = \new_[1348]_  | \new_[4952]_ ;
  assign \new_[4954]_  = \new_[4953]_  | \new_[4948]_ ;
  assign \new_[4955]_  = \new_[4954]_  | \new_[4945]_ ;
  assign \new_[4958]_  = \new_[1344]_  | \new_[1345]_ ;
  assign \new_[4962]_  = \new_[1341]_  | \new_[1342]_ ;
  assign \new_[4963]_  = \new_[1343]_  | \new_[4962]_ ;
  assign \new_[4964]_  = \new_[4963]_  | \new_[4958]_ ;
  assign \new_[4967]_  = \new_[1339]_  | \new_[1340]_ ;
  assign \new_[4971]_  = \new_[1336]_  | \new_[1337]_ ;
  assign \new_[4972]_  = \new_[1338]_  | \new_[4971]_ ;
  assign \new_[4973]_  = \new_[4972]_  | \new_[4967]_ ;
  assign \new_[4974]_  = \new_[4973]_  | \new_[4964]_ ;
  assign \new_[4975]_  = \new_[4974]_  | \new_[4955]_ ;
  assign \new_[4978]_  = \new_[1334]_  | \new_[1335]_ ;
  assign \new_[4982]_  = \new_[1331]_  | \new_[1332]_ ;
  assign \new_[4983]_  = \new_[1333]_  | \new_[4982]_ ;
  assign \new_[4984]_  = \new_[4983]_  | \new_[4978]_ ;
  assign \new_[4987]_  = \new_[1329]_  | \new_[1330]_ ;
  assign \new_[4991]_  = \new_[1326]_  | \new_[1327]_ ;
  assign \new_[4992]_  = \new_[1328]_  | \new_[4991]_ ;
  assign \new_[4993]_  = \new_[4992]_  | \new_[4987]_ ;
  assign \new_[4994]_  = \new_[4993]_  | \new_[4984]_ ;
  assign \new_[4997]_  = \new_[1324]_  | \new_[1325]_ ;
  assign \new_[5001]_  = \new_[1321]_  | \new_[1322]_ ;
  assign \new_[5002]_  = \new_[1323]_  | \new_[5001]_ ;
  assign \new_[5003]_  = \new_[5002]_  | \new_[4997]_ ;
  assign \new_[5006]_  = \new_[1319]_  | \new_[1320]_ ;
  assign \new_[5010]_  = \new_[1316]_  | \new_[1317]_ ;
  assign \new_[5011]_  = \new_[1318]_  | \new_[5010]_ ;
  assign \new_[5012]_  = \new_[5011]_  | \new_[5006]_ ;
  assign \new_[5013]_  = \new_[5012]_  | \new_[5003]_ ;
  assign \new_[5014]_  = \new_[5013]_  | \new_[4994]_ ;
  assign \new_[5015]_  = \new_[5014]_  | \new_[4975]_ ;
  assign \new_[5018]_  = \new_[1314]_  | \new_[1315]_ ;
  assign \new_[5022]_  = \new_[1311]_  | \new_[1312]_ ;
  assign \new_[5023]_  = \new_[1313]_  | \new_[5022]_ ;
  assign \new_[5024]_  = \new_[5023]_  | \new_[5018]_ ;
  assign \new_[5027]_  = \new_[1309]_  | \new_[1310]_ ;
  assign \new_[5031]_  = \new_[1306]_  | \new_[1307]_ ;
  assign \new_[5032]_  = \new_[1308]_  | \new_[5031]_ ;
  assign \new_[5033]_  = \new_[5032]_  | \new_[5027]_ ;
  assign \new_[5034]_  = \new_[5033]_  | \new_[5024]_ ;
  assign \new_[5037]_  = \new_[1304]_  | \new_[1305]_ ;
  assign \new_[5041]_  = \new_[1301]_  | \new_[1302]_ ;
  assign \new_[5042]_  = \new_[1303]_  | \new_[5041]_ ;
  assign \new_[5043]_  = \new_[5042]_  | \new_[5037]_ ;
  assign \new_[5046]_  = \new_[1299]_  | \new_[1300]_ ;
  assign \new_[5050]_  = \new_[1296]_  | \new_[1297]_ ;
  assign \new_[5051]_  = \new_[1298]_  | \new_[5050]_ ;
  assign \new_[5052]_  = \new_[5051]_  | \new_[5046]_ ;
  assign \new_[5053]_  = \new_[5052]_  | \new_[5043]_ ;
  assign \new_[5054]_  = \new_[5053]_  | \new_[5034]_ ;
  assign \new_[5057]_  = \new_[1294]_  | \new_[1295]_ ;
  assign \new_[5061]_  = \new_[1291]_  | \new_[1292]_ ;
  assign \new_[5062]_  = \new_[1293]_  | \new_[5061]_ ;
  assign \new_[5063]_  = \new_[5062]_  | \new_[5057]_ ;
  assign \new_[5066]_  = \new_[1289]_  | \new_[1290]_ ;
  assign \new_[5070]_  = \new_[1286]_  | \new_[1287]_ ;
  assign \new_[5071]_  = \new_[1288]_  | \new_[5070]_ ;
  assign \new_[5072]_  = \new_[5071]_  | \new_[5066]_ ;
  assign \new_[5073]_  = \new_[5072]_  | \new_[5063]_ ;
  assign \new_[5076]_  = \new_[1284]_  | \new_[1285]_ ;
  assign \new_[5080]_  = \new_[1281]_  | \new_[1282]_ ;
  assign \new_[5081]_  = \new_[1283]_  | \new_[5080]_ ;
  assign \new_[5082]_  = \new_[5081]_  | \new_[5076]_ ;
  assign \new_[5085]_  = \new_[1279]_  | \new_[1280]_ ;
  assign \new_[5089]_  = \new_[1276]_  | \new_[1277]_ ;
  assign \new_[5090]_  = \new_[1278]_  | \new_[5089]_ ;
  assign \new_[5091]_  = \new_[5090]_  | \new_[5085]_ ;
  assign \new_[5092]_  = \new_[5091]_  | \new_[5082]_ ;
  assign \new_[5093]_  = \new_[5092]_  | \new_[5073]_ ;
  assign \new_[5094]_  = \new_[5093]_  | \new_[5054]_ ;
  assign \new_[5095]_  = \new_[5094]_  | \new_[5015]_ ;
  assign \new_[5096]_  = \new_[5095]_  | \new_[4936]_ ;
  assign \new_[5097]_  = \new_[5096]_  | \new_[4777]_ ;
  assign \new_[5098]_  = \new_[5097]_  | \new_[4460]_ ;
  assign \new_[5099]_  = \new_[5098]_  | \new_[3823]_ ;
  assign \new_[5102]_  = \new_[1274]_  | \new_[1275]_ ;
  assign \new_[5105]_  = \new_[1272]_  | \new_[1273]_ ;
  assign \new_[5106]_  = \new_[5105]_  | \new_[5102]_ ;
  assign \new_[5109]_  = \new_[1270]_  | \new_[1271]_ ;
  assign \new_[5113]_  = \new_[1267]_  | \new_[1268]_ ;
  assign \new_[5114]_  = \new_[1269]_  | \new_[5113]_ ;
  assign \new_[5115]_  = \new_[5114]_  | \new_[5109]_ ;
  assign \new_[5116]_  = \new_[5115]_  | \new_[5106]_ ;
  assign \new_[5119]_  = \new_[1265]_  | \new_[1266]_ ;
  assign \new_[5123]_  = \new_[1262]_  | \new_[1263]_ ;
  assign \new_[5124]_  = \new_[1264]_  | \new_[5123]_ ;
  assign \new_[5125]_  = \new_[5124]_  | \new_[5119]_ ;
  assign \new_[5128]_  = \new_[1260]_  | \new_[1261]_ ;
  assign \new_[5132]_  = \new_[1257]_  | \new_[1258]_ ;
  assign \new_[5133]_  = \new_[1259]_  | \new_[5132]_ ;
  assign \new_[5134]_  = \new_[5133]_  | \new_[5128]_ ;
  assign \new_[5135]_  = \new_[5134]_  | \new_[5125]_ ;
  assign \new_[5136]_  = \new_[5135]_  | \new_[5116]_ ;
  assign \new_[5139]_  = \new_[1255]_  | \new_[1256]_ ;
  assign \new_[5143]_  = \new_[1252]_  | \new_[1253]_ ;
  assign \new_[5144]_  = \new_[1254]_  | \new_[5143]_ ;
  assign \new_[5145]_  = \new_[5144]_  | \new_[5139]_ ;
  assign \new_[5148]_  = \new_[1250]_  | \new_[1251]_ ;
  assign \new_[5152]_  = \new_[1247]_  | \new_[1248]_ ;
  assign \new_[5153]_  = \new_[1249]_  | \new_[5152]_ ;
  assign \new_[5154]_  = \new_[5153]_  | \new_[5148]_ ;
  assign \new_[5155]_  = \new_[5154]_  | \new_[5145]_ ;
  assign \new_[5158]_  = \new_[1245]_  | \new_[1246]_ ;
  assign \new_[5162]_  = \new_[1242]_  | \new_[1243]_ ;
  assign \new_[5163]_  = \new_[1244]_  | \new_[5162]_ ;
  assign \new_[5164]_  = \new_[5163]_  | \new_[5158]_ ;
  assign \new_[5167]_  = \new_[1240]_  | \new_[1241]_ ;
  assign \new_[5171]_  = \new_[1237]_  | \new_[1238]_ ;
  assign \new_[5172]_  = \new_[1239]_  | \new_[5171]_ ;
  assign \new_[5173]_  = \new_[5172]_  | \new_[5167]_ ;
  assign \new_[5174]_  = \new_[5173]_  | \new_[5164]_ ;
  assign \new_[5175]_  = \new_[5174]_  | \new_[5155]_ ;
  assign \new_[5176]_  = \new_[5175]_  | \new_[5136]_ ;
  assign \new_[5179]_  = \new_[1235]_  | \new_[1236]_ ;
  assign \new_[5183]_  = \new_[1232]_  | \new_[1233]_ ;
  assign \new_[5184]_  = \new_[1234]_  | \new_[5183]_ ;
  assign \new_[5185]_  = \new_[5184]_  | \new_[5179]_ ;
  assign \new_[5188]_  = \new_[1230]_  | \new_[1231]_ ;
  assign \new_[5192]_  = \new_[1227]_  | \new_[1228]_ ;
  assign \new_[5193]_  = \new_[1229]_  | \new_[5192]_ ;
  assign \new_[5194]_  = \new_[5193]_  | \new_[5188]_ ;
  assign \new_[5195]_  = \new_[5194]_  | \new_[5185]_ ;
  assign \new_[5198]_  = \new_[1225]_  | \new_[1226]_ ;
  assign \new_[5202]_  = \new_[1222]_  | \new_[1223]_ ;
  assign \new_[5203]_  = \new_[1224]_  | \new_[5202]_ ;
  assign \new_[5204]_  = \new_[5203]_  | \new_[5198]_ ;
  assign \new_[5207]_  = \new_[1220]_  | \new_[1221]_ ;
  assign \new_[5211]_  = \new_[1217]_  | \new_[1218]_ ;
  assign \new_[5212]_  = \new_[1219]_  | \new_[5211]_ ;
  assign \new_[5213]_  = \new_[5212]_  | \new_[5207]_ ;
  assign \new_[5214]_  = \new_[5213]_  | \new_[5204]_ ;
  assign \new_[5215]_  = \new_[5214]_  | \new_[5195]_ ;
  assign \new_[5218]_  = \new_[1215]_  | \new_[1216]_ ;
  assign \new_[5222]_  = \new_[1212]_  | \new_[1213]_ ;
  assign \new_[5223]_  = \new_[1214]_  | \new_[5222]_ ;
  assign \new_[5224]_  = \new_[5223]_  | \new_[5218]_ ;
  assign \new_[5227]_  = \new_[1210]_  | \new_[1211]_ ;
  assign \new_[5231]_  = \new_[1207]_  | \new_[1208]_ ;
  assign \new_[5232]_  = \new_[1209]_  | \new_[5231]_ ;
  assign \new_[5233]_  = \new_[5232]_  | \new_[5227]_ ;
  assign \new_[5234]_  = \new_[5233]_  | \new_[5224]_ ;
  assign \new_[5237]_  = \new_[1205]_  | \new_[1206]_ ;
  assign \new_[5241]_  = \new_[1202]_  | \new_[1203]_ ;
  assign \new_[5242]_  = \new_[1204]_  | \new_[5241]_ ;
  assign \new_[5243]_  = \new_[5242]_  | \new_[5237]_ ;
  assign \new_[5246]_  = \new_[1200]_  | \new_[1201]_ ;
  assign \new_[5250]_  = \new_[1197]_  | \new_[1198]_ ;
  assign \new_[5251]_  = \new_[1199]_  | \new_[5250]_ ;
  assign \new_[5252]_  = \new_[5251]_  | \new_[5246]_ ;
  assign \new_[5253]_  = \new_[5252]_  | \new_[5243]_ ;
  assign \new_[5254]_  = \new_[5253]_  | \new_[5234]_ ;
  assign \new_[5255]_  = \new_[5254]_  | \new_[5215]_ ;
  assign \new_[5256]_  = \new_[5255]_  | \new_[5176]_ ;
  assign \new_[5259]_  = \new_[1195]_  | \new_[1196]_ ;
  assign \new_[5263]_  = \new_[1192]_  | \new_[1193]_ ;
  assign \new_[5264]_  = \new_[1194]_  | \new_[5263]_ ;
  assign \new_[5265]_  = \new_[5264]_  | \new_[5259]_ ;
  assign \new_[5268]_  = \new_[1190]_  | \new_[1191]_ ;
  assign \new_[5272]_  = \new_[1187]_  | \new_[1188]_ ;
  assign \new_[5273]_  = \new_[1189]_  | \new_[5272]_ ;
  assign \new_[5274]_  = \new_[5273]_  | \new_[5268]_ ;
  assign \new_[5275]_  = \new_[5274]_  | \new_[5265]_ ;
  assign \new_[5278]_  = \new_[1185]_  | \new_[1186]_ ;
  assign \new_[5282]_  = \new_[1182]_  | \new_[1183]_ ;
  assign \new_[5283]_  = \new_[1184]_  | \new_[5282]_ ;
  assign \new_[5284]_  = \new_[5283]_  | \new_[5278]_ ;
  assign \new_[5287]_  = \new_[1180]_  | \new_[1181]_ ;
  assign \new_[5291]_  = \new_[1177]_  | \new_[1178]_ ;
  assign \new_[5292]_  = \new_[1179]_  | \new_[5291]_ ;
  assign \new_[5293]_  = \new_[5292]_  | \new_[5287]_ ;
  assign \new_[5294]_  = \new_[5293]_  | \new_[5284]_ ;
  assign \new_[5295]_  = \new_[5294]_  | \new_[5275]_ ;
  assign \new_[5298]_  = \new_[1175]_  | \new_[1176]_ ;
  assign \new_[5302]_  = \new_[1172]_  | \new_[1173]_ ;
  assign \new_[5303]_  = \new_[1174]_  | \new_[5302]_ ;
  assign \new_[5304]_  = \new_[5303]_  | \new_[5298]_ ;
  assign \new_[5307]_  = \new_[1170]_  | \new_[1171]_ ;
  assign \new_[5311]_  = \new_[1167]_  | \new_[1168]_ ;
  assign \new_[5312]_  = \new_[1169]_  | \new_[5311]_ ;
  assign \new_[5313]_  = \new_[5312]_  | \new_[5307]_ ;
  assign \new_[5314]_  = \new_[5313]_  | \new_[5304]_ ;
  assign \new_[5317]_  = \new_[1165]_  | \new_[1166]_ ;
  assign \new_[5321]_  = \new_[1162]_  | \new_[1163]_ ;
  assign \new_[5322]_  = \new_[1164]_  | \new_[5321]_ ;
  assign \new_[5323]_  = \new_[5322]_  | \new_[5317]_ ;
  assign \new_[5326]_  = \new_[1160]_  | \new_[1161]_ ;
  assign \new_[5330]_  = \new_[1157]_  | \new_[1158]_ ;
  assign \new_[5331]_  = \new_[1159]_  | \new_[5330]_ ;
  assign \new_[5332]_  = \new_[5331]_  | \new_[5326]_ ;
  assign \new_[5333]_  = \new_[5332]_  | \new_[5323]_ ;
  assign \new_[5334]_  = \new_[5333]_  | \new_[5314]_ ;
  assign \new_[5335]_  = \new_[5334]_  | \new_[5295]_ ;
  assign \new_[5338]_  = \new_[1155]_  | \new_[1156]_ ;
  assign \new_[5342]_  = \new_[1152]_  | \new_[1153]_ ;
  assign \new_[5343]_  = \new_[1154]_  | \new_[5342]_ ;
  assign \new_[5344]_  = \new_[5343]_  | \new_[5338]_ ;
  assign \new_[5347]_  = \new_[1150]_  | \new_[1151]_ ;
  assign \new_[5351]_  = \new_[1147]_  | \new_[1148]_ ;
  assign \new_[5352]_  = \new_[1149]_  | \new_[5351]_ ;
  assign \new_[5353]_  = \new_[5352]_  | \new_[5347]_ ;
  assign \new_[5354]_  = \new_[5353]_  | \new_[5344]_ ;
  assign \new_[5357]_  = \new_[1145]_  | \new_[1146]_ ;
  assign \new_[5361]_  = \new_[1142]_  | \new_[1143]_ ;
  assign \new_[5362]_  = \new_[1144]_  | \new_[5361]_ ;
  assign \new_[5363]_  = \new_[5362]_  | \new_[5357]_ ;
  assign \new_[5366]_  = \new_[1140]_  | \new_[1141]_ ;
  assign \new_[5370]_  = \new_[1137]_  | \new_[1138]_ ;
  assign \new_[5371]_  = \new_[1139]_  | \new_[5370]_ ;
  assign \new_[5372]_  = \new_[5371]_  | \new_[5366]_ ;
  assign \new_[5373]_  = \new_[5372]_  | \new_[5363]_ ;
  assign \new_[5374]_  = \new_[5373]_  | \new_[5354]_ ;
  assign \new_[5377]_  = \new_[1135]_  | \new_[1136]_ ;
  assign \new_[5381]_  = \new_[1132]_  | \new_[1133]_ ;
  assign \new_[5382]_  = \new_[1134]_  | \new_[5381]_ ;
  assign \new_[5383]_  = \new_[5382]_  | \new_[5377]_ ;
  assign \new_[5386]_  = \new_[1130]_  | \new_[1131]_ ;
  assign \new_[5390]_  = \new_[1127]_  | \new_[1128]_ ;
  assign \new_[5391]_  = \new_[1129]_  | \new_[5390]_ ;
  assign \new_[5392]_  = \new_[5391]_  | \new_[5386]_ ;
  assign \new_[5393]_  = \new_[5392]_  | \new_[5383]_ ;
  assign \new_[5396]_  = \new_[1125]_  | \new_[1126]_ ;
  assign \new_[5400]_  = \new_[1122]_  | \new_[1123]_ ;
  assign \new_[5401]_  = \new_[1124]_  | \new_[5400]_ ;
  assign \new_[5402]_  = \new_[5401]_  | \new_[5396]_ ;
  assign \new_[5405]_  = \new_[1120]_  | \new_[1121]_ ;
  assign \new_[5409]_  = \new_[1117]_  | \new_[1118]_ ;
  assign \new_[5410]_  = \new_[1119]_  | \new_[5409]_ ;
  assign \new_[5411]_  = \new_[5410]_  | \new_[5405]_ ;
  assign \new_[5412]_  = \new_[5411]_  | \new_[5402]_ ;
  assign \new_[5413]_  = \new_[5412]_  | \new_[5393]_ ;
  assign \new_[5414]_  = \new_[5413]_  | \new_[5374]_ ;
  assign \new_[5415]_  = \new_[5414]_  | \new_[5335]_ ;
  assign \new_[5416]_  = \new_[5415]_  | \new_[5256]_ ;
  assign \new_[5419]_  = \new_[1115]_  | \new_[1116]_ ;
  assign \new_[5422]_  = \new_[1113]_  | \new_[1114]_ ;
  assign \new_[5423]_  = \new_[5422]_  | \new_[5419]_ ;
  assign \new_[5426]_  = \new_[1111]_  | \new_[1112]_ ;
  assign \new_[5430]_  = \new_[1108]_  | \new_[1109]_ ;
  assign \new_[5431]_  = \new_[1110]_  | \new_[5430]_ ;
  assign \new_[5432]_  = \new_[5431]_  | \new_[5426]_ ;
  assign \new_[5433]_  = \new_[5432]_  | \new_[5423]_ ;
  assign \new_[5436]_  = \new_[1106]_  | \new_[1107]_ ;
  assign \new_[5440]_  = \new_[1103]_  | \new_[1104]_ ;
  assign \new_[5441]_  = \new_[1105]_  | \new_[5440]_ ;
  assign \new_[5442]_  = \new_[5441]_  | \new_[5436]_ ;
  assign \new_[5445]_  = \new_[1101]_  | \new_[1102]_ ;
  assign \new_[5449]_  = \new_[1098]_  | \new_[1099]_ ;
  assign \new_[5450]_  = \new_[1100]_  | \new_[5449]_ ;
  assign \new_[5451]_  = \new_[5450]_  | \new_[5445]_ ;
  assign \new_[5452]_  = \new_[5451]_  | \new_[5442]_ ;
  assign \new_[5453]_  = \new_[5452]_  | \new_[5433]_ ;
  assign \new_[5456]_  = \new_[1096]_  | \new_[1097]_ ;
  assign \new_[5460]_  = \new_[1093]_  | \new_[1094]_ ;
  assign \new_[5461]_  = \new_[1095]_  | \new_[5460]_ ;
  assign \new_[5462]_  = \new_[5461]_  | \new_[5456]_ ;
  assign \new_[5465]_  = \new_[1091]_  | \new_[1092]_ ;
  assign \new_[5469]_  = \new_[1088]_  | \new_[1089]_ ;
  assign \new_[5470]_  = \new_[1090]_  | \new_[5469]_ ;
  assign \new_[5471]_  = \new_[5470]_  | \new_[5465]_ ;
  assign \new_[5472]_  = \new_[5471]_  | \new_[5462]_ ;
  assign \new_[5475]_  = \new_[1086]_  | \new_[1087]_ ;
  assign \new_[5479]_  = \new_[1083]_  | \new_[1084]_ ;
  assign \new_[5480]_  = \new_[1085]_  | \new_[5479]_ ;
  assign \new_[5481]_  = \new_[5480]_  | \new_[5475]_ ;
  assign \new_[5484]_  = \new_[1081]_  | \new_[1082]_ ;
  assign \new_[5488]_  = \new_[1078]_  | \new_[1079]_ ;
  assign \new_[5489]_  = \new_[1080]_  | \new_[5488]_ ;
  assign \new_[5490]_  = \new_[5489]_  | \new_[5484]_ ;
  assign \new_[5491]_  = \new_[5490]_  | \new_[5481]_ ;
  assign \new_[5492]_  = \new_[5491]_  | \new_[5472]_ ;
  assign \new_[5493]_  = \new_[5492]_  | \new_[5453]_ ;
  assign \new_[5496]_  = \new_[1076]_  | \new_[1077]_ ;
  assign \new_[5500]_  = \new_[1073]_  | \new_[1074]_ ;
  assign \new_[5501]_  = \new_[1075]_  | \new_[5500]_ ;
  assign \new_[5502]_  = \new_[5501]_  | \new_[5496]_ ;
  assign \new_[5505]_  = \new_[1071]_  | \new_[1072]_ ;
  assign \new_[5509]_  = \new_[1068]_  | \new_[1069]_ ;
  assign \new_[5510]_  = \new_[1070]_  | \new_[5509]_ ;
  assign \new_[5511]_  = \new_[5510]_  | \new_[5505]_ ;
  assign \new_[5512]_  = \new_[5511]_  | \new_[5502]_ ;
  assign \new_[5515]_  = \new_[1066]_  | \new_[1067]_ ;
  assign \new_[5519]_  = \new_[1063]_  | \new_[1064]_ ;
  assign \new_[5520]_  = \new_[1065]_  | \new_[5519]_ ;
  assign \new_[5521]_  = \new_[5520]_  | \new_[5515]_ ;
  assign \new_[5524]_  = \new_[1061]_  | \new_[1062]_ ;
  assign \new_[5528]_  = \new_[1058]_  | \new_[1059]_ ;
  assign \new_[5529]_  = \new_[1060]_  | \new_[5528]_ ;
  assign \new_[5530]_  = \new_[5529]_  | \new_[5524]_ ;
  assign \new_[5531]_  = \new_[5530]_  | \new_[5521]_ ;
  assign \new_[5532]_  = \new_[5531]_  | \new_[5512]_ ;
  assign \new_[5535]_  = \new_[1056]_  | \new_[1057]_ ;
  assign \new_[5539]_  = \new_[1053]_  | \new_[1054]_ ;
  assign \new_[5540]_  = \new_[1055]_  | \new_[5539]_ ;
  assign \new_[5541]_  = \new_[5540]_  | \new_[5535]_ ;
  assign \new_[5544]_  = \new_[1051]_  | \new_[1052]_ ;
  assign \new_[5548]_  = \new_[1048]_  | \new_[1049]_ ;
  assign \new_[5549]_  = \new_[1050]_  | \new_[5548]_ ;
  assign \new_[5550]_  = \new_[5549]_  | \new_[5544]_ ;
  assign \new_[5551]_  = \new_[5550]_  | \new_[5541]_ ;
  assign \new_[5554]_  = \new_[1046]_  | \new_[1047]_ ;
  assign \new_[5558]_  = \new_[1043]_  | \new_[1044]_ ;
  assign \new_[5559]_  = \new_[1045]_  | \new_[5558]_ ;
  assign \new_[5560]_  = \new_[5559]_  | \new_[5554]_ ;
  assign \new_[5563]_  = \new_[1041]_  | \new_[1042]_ ;
  assign \new_[5567]_  = \new_[1038]_  | \new_[1039]_ ;
  assign \new_[5568]_  = \new_[1040]_  | \new_[5567]_ ;
  assign \new_[5569]_  = \new_[5568]_  | \new_[5563]_ ;
  assign \new_[5570]_  = \new_[5569]_  | \new_[5560]_ ;
  assign \new_[5571]_  = \new_[5570]_  | \new_[5551]_ ;
  assign \new_[5572]_  = \new_[5571]_  | \new_[5532]_ ;
  assign \new_[5573]_  = \new_[5572]_  | \new_[5493]_ ;
  assign \new_[5576]_  = \new_[1036]_  | \new_[1037]_ ;
  assign \new_[5580]_  = \new_[1033]_  | \new_[1034]_ ;
  assign \new_[5581]_  = \new_[1035]_  | \new_[5580]_ ;
  assign \new_[5582]_  = \new_[5581]_  | \new_[5576]_ ;
  assign \new_[5585]_  = \new_[1031]_  | \new_[1032]_ ;
  assign \new_[5589]_  = \new_[1028]_  | \new_[1029]_ ;
  assign \new_[5590]_  = \new_[1030]_  | \new_[5589]_ ;
  assign \new_[5591]_  = \new_[5590]_  | \new_[5585]_ ;
  assign \new_[5592]_  = \new_[5591]_  | \new_[5582]_ ;
  assign \new_[5595]_  = \new_[1026]_  | \new_[1027]_ ;
  assign \new_[5599]_  = \new_[1023]_  | \new_[1024]_ ;
  assign \new_[5600]_  = \new_[1025]_  | \new_[5599]_ ;
  assign \new_[5601]_  = \new_[5600]_  | \new_[5595]_ ;
  assign \new_[5604]_  = \new_[1021]_  | \new_[1022]_ ;
  assign \new_[5608]_  = \new_[1018]_  | \new_[1019]_ ;
  assign \new_[5609]_  = \new_[1020]_  | \new_[5608]_ ;
  assign \new_[5610]_  = \new_[5609]_  | \new_[5604]_ ;
  assign \new_[5611]_  = \new_[5610]_  | \new_[5601]_ ;
  assign \new_[5612]_  = \new_[5611]_  | \new_[5592]_ ;
  assign \new_[5615]_  = \new_[1016]_  | \new_[1017]_ ;
  assign \new_[5619]_  = \new_[1013]_  | \new_[1014]_ ;
  assign \new_[5620]_  = \new_[1015]_  | \new_[5619]_ ;
  assign \new_[5621]_  = \new_[5620]_  | \new_[5615]_ ;
  assign \new_[5624]_  = \new_[1011]_  | \new_[1012]_ ;
  assign \new_[5628]_  = \new_[1008]_  | \new_[1009]_ ;
  assign \new_[5629]_  = \new_[1010]_  | \new_[5628]_ ;
  assign \new_[5630]_  = \new_[5629]_  | \new_[5624]_ ;
  assign \new_[5631]_  = \new_[5630]_  | \new_[5621]_ ;
  assign \new_[5634]_  = \new_[1006]_  | \new_[1007]_ ;
  assign \new_[5638]_  = \new_[1003]_  | \new_[1004]_ ;
  assign \new_[5639]_  = \new_[1005]_  | \new_[5638]_ ;
  assign \new_[5640]_  = \new_[5639]_  | \new_[5634]_ ;
  assign \new_[5643]_  = \new_[1001]_  | \new_[1002]_ ;
  assign \new_[5647]_  = \new_[998]_  | \new_[999]_ ;
  assign \new_[5648]_  = \new_[1000]_  | \new_[5647]_ ;
  assign \new_[5649]_  = \new_[5648]_  | \new_[5643]_ ;
  assign \new_[5650]_  = \new_[5649]_  | \new_[5640]_ ;
  assign \new_[5651]_  = \new_[5650]_  | \new_[5631]_ ;
  assign \new_[5652]_  = \new_[5651]_  | \new_[5612]_ ;
  assign \new_[5655]_  = \new_[996]_  | \new_[997]_ ;
  assign \new_[5659]_  = \new_[993]_  | \new_[994]_ ;
  assign \new_[5660]_  = \new_[995]_  | \new_[5659]_ ;
  assign \new_[5661]_  = \new_[5660]_  | \new_[5655]_ ;
  assign \new_[5664]_  = \new_[991]_  | \new_[992]_ ;
  assign \new_[5668]_  = \new_[988]_  | \new_[989]_ ;
  assign \new_[5669]_  = \new_[990]_  | \new_[5668]_ ;
  assign \new_[5670]_  = \new_[5669]_  | \new_[5664]_ ;
  assign \new_[5671]_  = \new_[5670]_  | \new_[5661]_ ;
  assign \new_[5674]_  = \new_[986]_  | \new_[987]_ ;
  assign \new_[5678]_  = \new_[983]_  | \new_[984]_ ;
  assign \new_[5679]_  = \new_[985]_  | \new_[5678]_ ;
  assign \new_[5680]_  = \new_[5679]_  | \new_[5674]_ ;
  assign \new_[5683]_  = \new_[981]_  | \new_[982]_ ;
  assign \new_[5687]_  = \new_[978]_  | \new_[979]_ ;
  assign \new_[5688]_  = \new_[980]_  | \new_[5687]_ ;
  assign \new_[5689]_  = \new_[5688]_  | \new_[5683]_ ;
  assign \new_[5690]_  = \new_[5689]_  | \new_[5680]_ ;
  assign \new_[5691]_  = \new_[5690]_  | \new_[5671]_ ;
  assign \new_[5694]_  = \new_[976]_  | \new_[977]_ ;
  assign \new_[5698]_  = \new_[973]_  | \new_[974]_ ;
  assign \new_[5699]_  = \new_[975]_  | \new_[5698]_ ;
  assign \new_[5700]_  = \new_[5699]_  | \new_[5694]_ ;
  assign \new_[5703]_  = \new_[971]_  | \new_[972]_ ;
  assign \new_[5707]_  = \new_[968]_  | \new_[969]_ ;
  assign \new_[5708]_  = \new_[970]_  | \new_[5707]_ ;
  assign \new_[5709]_  = \new_[5708]_  | \new_[5703]_ ;
  assign \new_[5710]_  = \new_[5709]_  | \new_[5700]_ ;
  assign \new_[5713]_  = \new_[966]_  | \new_[967]_ ;
  assign \new_[5717]_  = \new_[963]_  | \new_[964]_ ;
  assign \new_[5718]_  = \new_[965]_  | \new_[5717]_ ;
  assign \new_[5719]_  = \new_[5718]_  | \new_[5713]_ ;
  assign \new_[5722]_  = \new_[961]_  | \new_[962]_ ;
  assign \new_[5726]_  = \new_[958]_  | \new_[959]_ ;
  assign \new_[5727]_  = \new_[960]_  | \new_[5726]_ ;
  assign \new_[5728]_  = \new_[5727]_  | \new_[5722]_ ;
  assign \new_[5729]_  = \new_[5728]_  | \new_[5719]_ ;
  assign \new_[5730]_  = \new_[5729]_  | \new_[5710]_ ;
  assign \new_[5731]_  = \new_[5730]_  | \new_[5691]_ ;
  assign \new_[5732]_  = \new_[5731]_  | \new_[5652]_ ;
  assign \new_[5733]_  = \new_[5732]_  | \new_[5573]_ ;
  assign \new_[5734]_  = \new_[5733]_  | \new_[5416]_ ;
  assign \new_[5737]_  = \new_[956]_  | \new_[957]_ ;
  assign \new_[5740]_  = \new_[954]_  | \new_[955]_ ;
  assign \new_[5741]_  = \new_[5740]_  | \new_[5737]_ ;
  assign \new_[5744]_  = \new_[952]_  | \new_[953]_ ;
  assign \new_[5748]_  = \new_[949]_  | \new_[950]_ ;
  assign \new_[5749]_  = \new_[951]_  | \new_[5748]_ ;
  assign \new_[5750]_  = \new_[5749]_  | \new_[5744]_ ;
  assign \new_[5751]_  = \new_[5750]_  | \new_[5741]_ ;
  assign \new_[5754]_  = \new_[947]_  | \new_[948]_ ;
  assign \new_[5758]_  = \new_[944]_  | \new_[945]_ ;
  assign \new_[5759]_  = \new_[946]_  | \new_[5758]_ ;
  assign \new_[5760]_  = \new_[5759]_  | \new_[5754]_ ;
  assign \new_[5763]_  = \new_[942]_  | \new_[943]_ ;
  assign \new_[5767]_  = \new_[939]_  | \new_[940]_ ;
  assign \new_[5768]_  = \new_[941]_  | \new_[5767]_ ;
  assign \new_[5769]_  = \new_[5768]_  | \new_[5763]_ ;
  assign \new_[5770]_  = \new_[5769]_  | \new_[5760]_ ;
  assign \new_[5771]_  = \new_[5770]_  | \new_[5751]_ ;
  assign \new_[5774]_  = \new_[937]_  | \new_[938]_ ;
  assign \new_[5778]_  = \new_[934]_  | \new_[935]_ ;
  assign \new_[5779]_  = \new_[936]_  | \new_[5778]_ ;
  assign \new_[5780]_  = \new_[5779]_  | \new_[5774]_ ;
  assign \new_[5783]_  = \new_[932]_  | \new_[933]_ ;
  assign \new_[5787]_  = \new_[929]_  | \new_[930]_ ;
  assign \new_[5788]_  = \new_[931]_  | \new_[5787]_ ;
  assign \new_[5789]_  = \new_[5788]_  | \new_[5783]_ ;
  assign \new_[5790]_  = \new_[5789]_  | \new_[5780]_ ;
  assign \new_[5793]_  = \new_[927]_  | \new_[928]_ ;
  assign \new_[5797]_  = \new_[924]_  | \new_[925]_ ;
  assign \new_[5798]_  = \new_[926]_  | \new_[5797]_ ;
  assign \new_[5799]_  = \new_[5798]_  | \new_[5793]_ ;
  assign \new_[5802]_  = \new_[922]_  | \new_[923]_ ;
  assign \new_[5806]_  = \new_[919]_  | \new_[920]_ ;
  assign \new_[5807]_  = \new_[921]_  | \new_[5806]_ ;
  assign \new_[5808]_  = \new_[5807]_  | \new_[5802]_ ;
  assign \new_[5809]_  = \new_[5808]_  | \new_[5799]_ ;
  assign \new_[5810]_  = \new_[5809]_  | \new_[5790]_ ;
  assign \new_[5811]_  = \new_[5810]_  | \new_[5771]_ ;
  assign \new_[5814]_  = \new_[917]_  | \new_[918]_ ;
  assign \new_[5818]_  = \new_[914]_  | \new_[915]_ ;
  assign \new_[5819]_  = \new_[916]_  | \new_[5818]_ ;
  assign \new_[5820]_  = \new_[5819]_  | \new_[5814]_ ;
  assign \new_[5823]_  = \new_[912]_  | \new_[913]_ ;
  assign \new_[5827]_  = \new_[909]_  | \new_[910]_ ;
  assign \new_[5828]_  = \new_[911]_  | \new_[5827]_ ;
  assign \new_[5829]_  = \new_[5828]_  | \new_[5823]_ ;
  assign \new_[5830]_  = \new_[5829]_  | \new_[5820]_ ;
  assign \new_[5833]_  = \new_[907]_  | \new_[908]_ ;
  assign \new_[5837]_  = \new_[904]_  | \new_[905]_ ;
  assign \new_[5838]_  = \new_[906]_  | \new_[5837]_ ;
  assign \new_[5839]_  = \new_[5838]_  | \new_[5833]_ ;
  assign \new_[5842]_  = \new_[902]_  | \new_[903]_ ;
  assign \new_[5846]_  = \new_[899]_  | \new_[900]_ ;
  assign \new_[5847]_  = \new_[901]_  | \new_[5846]_ ;
  assign \new_[5848]_  = \new_[5847]_  | \new_[5842]_ ;
  assign \new_[5849]_  = \new_[5848]_  | \new_[5839]_ ;
  assign \new_[5850]_  = \new_[5849]_  | \new_[5830]_ ;
  assign \new_[5853]_  = \new_[897]_  | \new_[898]_ ;
  assign \new_[5857]_  = \new_[894]_  | \new_[895]_ ;
  assign \new_[5858]_  = \new_[896]_  | \new_[5857]_ ;
  assign \new_[5859]_  = \new_[5858]_  | \new_[5853]_ ;
  assign \new_[5862]_  = \new_[892]_  | \new_[893]_ ;
  assign \new_[5866]_  = \new_[889]_  | \new_[890]_ ;
  assign \new_[5867]_  = \new_[891]_  | \new_[5866]_ ;
  assign \new_[5868]_  = \new_[5867]_  | \new_[5862]_ ;
  assign \new_[5869]_  = \new_[5868]_  | \new_[5859]_ ;
  assign \new_[5872]_  = \new_[887]_  | \new_[888]_ ;
  assign \new_[5876]_  = \new_[884]_  | \new_[885]_ ;
  assign \new_[5877]_  = \new_[886]_  | \new_[5876]_ ;
  assign \new_[5878]_  = \new_[5877]_  | \new_[5872]_ ;
  assign \new_[5881]_  = \new_[882]_  | \new_[883]_ ;
  assign \new_[5885]_  = \new_[879]_  | \new_[880]_ ;
  assign \new_[5886]_  = \new_[881]_  | \new_[5885]_ ;
  assign \new_[5887]_  = \new_[5886]_  | \new_[5881]_ ;
  assign \new_[5888]_  = \new_[5887]_  | \new_[5878]_ ;
  assign \new_[5889]_  = \new_[5888]_  | \new_[5869]_ ;
  assign \new_[5890]_  = \new_[5889]_  | \new_[5850]_ ;
  assign \new_[5891]_  = \new_[5890]_  | \new_[5811]_ ;
  assign \new_[5894]_  = \new_[877]_  | \new_[878]_ ;
  assign \new_[5898]_  = \new_[874]_  | \new_[875]_ ;
  assign \new_[5899]_  = \new_[876]_  | \new_[5898]_ ;
  assign \new_[5900]_  = \new_[5899]_  | \new_[5894]_ ;
  assign \new_[5903]_  = \new_[872]_  | \new_[873]_ ;
  assign \new_[5907]_  = \new_[869]_  | \new_[870]_ ;
  assign \new_[5908]_  = \new_[871]_  | \new_[5907]_ ;
  assign \new_[5909]_  = \new_[5908]_  | \new_[5903]_ ;
  assign \new_[5910]_  = \new_[5909]_  | \new_[5900]_ ;
  assign \new_[5913]_  = \new_[867]_  | \new_[868]_ ;
  assign \new_[5917]_  = \new_[864]_  | \new_[865]_ ;
  assign \new_[5918]_  = \new_[866]_  | \new_[5917]_ ;
  assign \new_[5919]_  = \new_[5918]_  | \new_[5913]_ ;
  assign \new_[5922]_  = \new_[862]_  | \new_[863]_ ;
  assign \new_[5926]_  = \new_[859]_  | \new_[860]_ ;
  assign \new_[5927]_  = \new_[861]_  | \new_[5926]_ ;
  assign \new_[5928]_  = \new_[5927]_  | \new_[5922]_ ;
  assign \new_[5929]_  = \new_[5928]_  | \new_[5919]_ ;
  assign \new_[5930]_  = \new_[5929]_  | \new_[5910]_ ;
  assign \new_[5933]_  = \new_[857]_  | \new_[858]_ ;
  assign \new_[5937]_  = \new_[854]_  | \new_[855]_ ;
  assign \new_[5938]_  = \new_[856]_  | \new_[5937]_ ;
  assign \new_[5939]_  = \new_[5938]_  | \new_[5933]_ ;
  assign \new_[5942]_  = \new_[852]_  | \new_[853]_ ;
  assign \new_[5946]_  = \new_[849]_  | \new_[850]_ ;
  assign \new_[5947]_  = \new_[851]_  | \new_[5946]_ ;
  assign \new_[5948]_  = \new_[5947]_  | \new_[5942]_ ;
  assign \new_[5949]_  = \new_[5948]_  | \new_[5939]_ ;
  assign \new_[5952]_  = \new_[847]_  | \new_[848]_ ;
  assign \new_[5956]_  = \new_[844]_  | \new_[845]_ ;
  assign \new_[5957]_  = \new_[846]_  | \new_[5956]_ ;
  assign \new_[5958]_  = \new_[5957]_  | \new_[5952]_ ;
  assign \new_[5961]_  = \new_[842]_  | \new_[843]_ ;
  assign \new_[5965]_  = \new_[839]_  | \new_[840]_ ;
  assign \new_[5966]_  = \new_[841]_  | \new_[5965]_ ;
  assign \new_[5967]_  = \new_[5966]_  | \new_[5961]_ ;
  assign \new_[5968]_  = \new_[5967]_  | \new_[5958]_ ;
  assign \new_[5969]_  = \new_[5968]_  | \new_[5949]_ ;
  assign \new_[5970]_  = \new_[5969]_  | \new_[5930]_ ;
  assign \new_[5973]_  = \new_[837]_  | \new_[838]_ ;
  assign \new_[5977]_  = \new_[834]_  | \new_[835]_ ;
  assign \new_[5978]_  = \new_[836]_  | \new_[5977]_ ;
  assign \new_[5979]_  = \new_[5978]_  | \new_[5973]_ ;
  assign \new_[5982]_  = \new_[832]_  | \new_[833]_ ;
  assign \new_[5986]_  = \new_[829]_  | \new_[830]_ ;
  assign \new_[5987]_  = \new_[831]_  | \new_[5986]_ ;
  assign \new_[5988]_  = \new_[5987]_  | \new_[5982]_ ;
  assign \new_[5989]_  = \new_[5988]_  | \new_[5979]_ ;
  assign \new_[5992]_  = \new_[827]_  | \new_[828]_ ;
  assign \new_[5996]_  = \new_[824]_  | \new_[825]_ ;
  assign \new_[5997]_  = \new_[826]_  | \new_[5996]_ ;
  assign \new_[5998]_  = \new_[5997]_  | \new_[5992]_ ;
  assign \new_[6001]_  = \new_[822]_  | \new_[823]_ ;
  assign \new_[6005]_  = \new_[819]_  | \new_[820]_ ;
  assign \new_[6006]_  = \new_[821]_  | \new_[6005]_ ;
  assign \new_[6007]_  = \new_[6006]_  | \new_[6001]_ ;
  assign \new_[6008]_  = \new_[6007]_  | \new_[5998]_ ;
  assign \new_[6009]_  = \new_[6008]_  | \new_[5989]_ ;
  assign \new_[6012]_  = \new_[817]_  | \new_[818]_ ;
  assign \new_[6016]_  = \new_[814]_  | \new_[815]_ ;
  assign \new_[6017]_  = \new_[816]_  | \new_[6016]_ ;
  assign \new_[6018]_  = \new_[6017]_  | \new_[6012]_ ;
  assign \new_[6021]_  = \new_[812]_  | \new_[813]_ ;
  assign \new_[6025]_  = \new_[809]_  | \new_[810]_ ;
  assign \new_[6026]_  = \new_[811]_  | \new_[6025]_ ;
  assign \new_[6027]_  = \new_[6026]_  | \new_[6021]_ ;
  assign \new_[6028]_  = \new_[6027]_  | \new_[6018]_ ;
  assign \new_[6031]_  = \new_[807]_  | \new_[808]_ ;
  assign \new_[6035]_  = \new_[804]_  | \new_[805]_ ;
  assign \new_[6036]_  = \new_[806]_  | \new_[6035]_ ;
  assign \new_[6037]_  = \new_[6036]_  | \new_[6031]_ ;
  assign \new_[6040]_  = \new_[802]_  | \new_[803]_ ;
  assign \new_[6044]_  = \new_[799]_  | \new_[800]_ ;
  assign \new_[6045]_  = \new_[801]_  | \new_[6044]_ ;
  assign \new_[6046]_  = \new_[6045]_  | \new_[6040]_ ;
  assign \new_[6047]_  = \new_[6046]_  | \new_[6037]_ ;
  assign \new_[6048]_  = \new_[6047]_  | \new_[6028]_ ;
  assign \new_[6049]_  = \new_[6048]_  | \new_[6009]_ ;
  assign \new_[6050]_  = \new_[6049]_  | \new_[5970]_ ;
  assign \new_[6051]_  = \new_[6050]_  | \new_[5891]_ ;
  assign \new_[6054]_  = \new_[797]_  | \new_[798]_ ;
  assign \new_[6058]_  = \new_[794]_  | \new_[795]_ ;
  assign \new_[6059]_  = \new_[796]_  | \new_[6058]_ ;
  assign \new_[6060]_  = \new_[6059]_  | \new_[6054]_ ;
  assign \new_[6063]_  = \new_[792]_  | \new_[793]_ ;
  assign \new_[6067]_  = \new_[789]_  | \new_[790]_ ;
  assign \new_[6068]_  = \new_[791]_  | \new_[6067]_ ;
  assign \new_[6069]_  = \new_[6068]_  | \new_[6063]_ ;
  assign \new_[6070]_  = \new_[6069]_  | \new_[6060]_ ;
  assign \new_[6073]_  = \new_[787]_  | \new_[788]_ ;
  assign \new_[6077]_  = \new_[784]_  | \new_[785]_ ;
  assign \new_[6078]_  = \new_[786]_  | \new_[6077]_ ;
  assign \new_[6079]_  = \new_[6078]_  | \new_[6073]_ ;
  assign \new_[6082]_  = \new_[782]_  | \new_[783]_ ;
  assign \new_[6086]_  = \new_[779]_  | \new_[780]_ ;
  assign \new_[6087]_  = \new_[781]_  | \new_[6086]_ ;
  assign \new_[6088]_  = \new_[6087]_  | \new_[6082]_ ;
  assign \new_[6089]_  = \new_[6088]_  | \new_[6079]_ ;
  assign \new_[6090]_  = \new_[6089]_  | \new_[6070]_ ;
  assign \new_[6093]_  = \new_[777]_  | \new_[778]_ ;
  assign \new_[6097]_  = \new_[774]_  | \new_[775]_ ;
  assign \new_[6098]_  = \new_[776]_  | \new_[6097]_ ;
  assign \new_[6099]_  = \new_[6098]_  | \new_[6093]_ ;
  assign \new_[6102]_  = \new_[772]_  | \new_[773]_ ;
  assign \new_[6106]_  = \new_[769]_  | \new_[770]_ ;
  assign \new_[6107]_  = \new_[771]_  | \new_[6106]_ ;
  assign \new_[6108]_  = \new_[6107]_  | \new_[6102]_ ;
  assign \new_[6109]_  = \new_[6108]_  | \new_[6099]_ ;
  assign \new_[6112]_  = \new_[767]_  | \new_[768]_ ;
  assign \new_[6116]_  = \new_[764]_  | \new_[765]_ ;
  assign \new_[6117]_  = \new_[766]_  | \new_[6116]_ ;
  assign \new_[6118]_  = \new_[6117]_  | \new_[6112]_ ;
  assign \new_[6121]_  = \new_[762]_  | \new_[763]_ ;
  assign \new_[6125]_  = \new_[759]_  | \new_[760]_ ;
  assign \new_[6126]_  = \new_[761]_  | \new_[6125]_ ;
  assign \new_[6127]_  = \new_[6126]_  | \new_[6121]_ ;
  assign \new_[6128]_  = \new_[6127]_  | \new_[6118]_ ;
  assign \new_[6129]_  = \new_[6128]_  | \new_[6109]_ ;
  assign \new_[6130]_  = \new_[6129]_  | \new_[6090]_ ;
  assign \new_[6133]_  = \new_[757]_  | \new_[758]_ ;
  assign \new_[6137]_  = \new_[754]_  | \new_[755]_ ;
  assign \new_[6138]_  = \new_[756]_  | \new_[6137]_ ;
  assign \new_[6139]_  = \new_[6138]_  | \new_[6133]_ ;
  assign \new_[6142]_  = \new_[752]_  | \new_[753]_ ;
  assign \new_[6146]_  = \new_[749]_  | \new_[750]_ ;
  assign \new_[6147]_  = \new_[751]_  | \new_[6146]_ ;
  assign \new_[6148]_  = \new_[6147]_  | \new_[6142]_ ;
  assign \new_[6149]_  = \new_[6148]_  | \new_[6139]_ ;
  assign \new_[6152]_  = \new_[747]_  | \new_[748]_ ;
  assign \new_[6156]_  = \new_[744]_  | \new_[745]_ ;
  assign \new_[6157]_  = \new_[746]_  | \new_[6156]_ ;
  assign \new_[6158]_  = \new_[6157]_  | \new_[6152]_ ;
  assign \new_[6161]_  = \new_[742]_  | \new_[743]_ ;
  assign \new_[6165]_  = \new_[739]_  | \new_[740]_ ;
  assign \new_[6166]_  = \new_[741]_  | \new_[6165]_ ;
  assign \new_[6167]_  = \new_[6166]_  | \new_[6161]_ ;
  assign \new_[6168]_  = \new_[6167]_  | \new_[6158]_ ;
  assign \new_[6169]_  = \new_[6168]_  | \new_[6149]_ ;
  assign \new_[6172]_  = \new_[737]_  | \new_[738]_ ;
  assign \new_[6176]_  = \new_[734]_  | \new_[735]_ ;
  assign \new_[6177]_  = \new_[736]_  | \new_[6176]_ ;
  assign \new_[6178]_  = \new_[6177]_  | \new_[6172]_ ;
  assign \new_[6181]_  = \new_[732]_  | \new_[733]_ ;
  assign \new_[6185]_  = \new_[729]_  | \new_[730]_ ;
  assign \new_[6186]_  = \new_[731]_  | \new_[6185]_ ;
  assign \new_[6187]_  = \new_[6186]_  | \new_[6181]_ ;
  assign \new_[6188]_  = \new_[6187]_  | \new_[6178]_ ;
  assign \new_[6191]_  = \new_[727]_  | \new_[728]_ ;
  assign \new_[6195]_  = \new_[724]_  | \new_[725]_ ;
  assign \new_[6196]_  = \new_[726]_  | \new_[6195]_ ;
  assign \new_[6197]_  = \new_[6196]_  | \new_[6191]_ ;
  assign \new_[6200]_  = \new_[722]_  | \new_[723]_ ;
  assign \new_[6204]_  = \new_[719]_  | \new_[720]_ ;
  assign \new_[6205]_  = \new_[721]_  | \new_[6204]_ ;
  assign \new_[6206]_  = \new_[6205]_  | \new_[6200]_ ;
  assign \new_[6207]_  = \new_[6206]_  | \new_[6197]_ ;
  assign \new_[6208]_  = \new_[6207]_  | \new_[6188]_ ;
  assign \new_[6209]_  = \new_[6208]_  | \new_[6169]_ ;
  assign \new_[6210]_  = \new_[6209]_  | \new_[6130]_ ;
  assign \new_[6213]_  = \new_[717]_  | \new_[718]_ ;
  assign \new_[6217]_  = \new_[714]_  | \new_[715]_ ;
  assign \new_[6218]_  = \new_[716]_  | \new_[6217]_ ;
  assign \new_[6219]_  = \new_[6218]_  | \new_[6213]_ ;
  assign \new_[6222]_  = \new_[712]_  | \new_[713]_ ;
  assign \new_[6226]_  = \new_[709]_  | \new_[710]_ ;
  assign \new_[6227]_  = \new_[711]_  | \new_[6226]_ ;
  assign \new_[6228]_  = \new_[6227]_  | \new_[6222]_ ;
  assign \new_[6229]_  = \new_[6228]_  | \new_[6219]_ ;
  assign \new_[6232]_  = \new_[707]_  | \new_[708]_ ;
  assign \new_[6236]_  = \new_[704]_  | \new_[705]_ ;
  assign \new_[6237]_  = \new_[706]_  | \new_[6236]_ ;
  assign \new_[6238]_  = \new_[6237]_  | \new_[6232]_ ;
  assign \new_[6241]_  = \new_[702]_  | \new_[703]_ ;
  assign \new_[6245]_  = \new_[699]_  | \new_[700]_ ;
  assign \new_[6246]_  = \new_[701]_  | \new_[6245]_ ;
  assign \new_[6247]_  = \new_[6246]_  | \new_[6241]_ ;
  assign \new_[6248]_  = \new_[6247]_  | \new_[6238]_ ;
  assign \new_[6249]_  = \new_[6248]_  | \new_[6229]_ ;
  assign \new_[6252]_  = \new_[697]_  | \new_[698]_ ;
  assign \new_[6256]_  = \new_[694]_  | \new_[695]_ ;
  assign \new_[6257]_  = \new_[696]_  | \new_[6256]_ ;
  assign \new_[6258]_  = \new_[6257]_  | \new_[6252]_ ;
  assign \new_[6261]_  = \new_[692]_  | \new_[693]_ ;
  assign \new_[6265]_  = \new_[689]_  | \new_[690]_ ;
  assign \new_[6266]_  = \new_[691]_  | \new_[6265]_ ;
  assign \new_[6267]_  = \new_[6266]_  | \new_[6261]_ ;
  assign \new_[6268]_  = \new_[6267]_  | \new_[6258]_ ;
  assign \new_[6271]_  = \new_[687]_  | \new_[688]_ ;
  assign \new_[6275]_  = \new_[684]_  | \new_[685]_ ;
  assign \new_[6276]_  = \new_[686]_  | \new_[6275]_ ;
  assign \new_[6277]_  = \new_[6276]_  | \new_[6271]_ ;
  assign \new_[6280]_  = \new_[682]_  | \new_[683]_ ;
  assign \new_[6284]_  = \new_[679]_  | \new_[680]_ ;
  assign \new_[6285]_  = \new_[681]_  | \new_[6284]_ ;
  assign \new_[6286]_  = \new_[6285]_  | \new_[6280]_ ;
  assign \new_[6287]_  = \new_[6286]_  | \new_[6277]_ ;
  assign \new_[6288]_  = \new_[6287]_  | \new_[6268]_ ;
  assign \new_[6289]_  = \new_[6288]_  | \new_[6249]_ ;
  assign \new_[6292]_  = \new_[677]_  | \new_[678]_ ;
  assign \new_[6296]_  = \new_[674]_  | \new_[675]_ ;
  assign \new_[6297]_  = \new_[676]_  | \new_[6296]_ ;
  assign \new_[6298]_  = \new_[6297]_  | \new_[6292]_ ;
  assign \new_[6301]_  = \new_[672]_  | \new_[673]_ ;
  assign \new_[6305]_  = \new_[669]_  | \new_[670]_ ;
  assign \new_[6306]_  = \new_[671]_  | \new_[6305]_ ;
  assign \new_[6307]_  = \new_[6306]_  | \new_[6301]_ ;
  assign \new_[6308]_  = \new_[6307]_  | \new_[6298]_ ;
  assign \new_[6311]_  = \new_[667]_  | \new_[668]_ ;
  assign \new_[6315]_  = \new_[664]_  | \new_[665]_ ;
  assign \new_[6316]_  = \new_[666]_  | \new_[6315]_ ;
  assign \new_[6317]_  = \new_[6316]_  | \new_[6311]_ ;
  assign \new_[6320]_  = \new_[662]_  | \new_[663]_ ;
  assign \new_[6324]_  = \new_[659]_  | \new_[660]_ ;
  assign \new_[6325]_  = \new_[661]_  | \new_[6324]_ ;
  assign \new_[6326]_  = \new_[6325]_  | \new_[6320]_ ;
  assign \new_[6327]_  = \new_[6326]_  | \new_[6317]_ ;
  assign \new_[6328]_  = \new_[6327]_  | \new_[6308]_ ;
  assign \new_[6331]_  = \new_[657]_  | \new_[658]_ ;
  assign \new_[6335]_  = \new_[654]_  | \new_[655]_ ;
  assign \new_[6336]_  = \new_[656]_  | \new_[6335]_ ;
  assign \new_[6337]_  = \new_[6336]_  | \new_[6331]_ ;
  assign \new_[6340]_  = \new_[652]_  | \new_[653]_ ;
  assign \new_[6344]_  = \new_[649]_  | \new_[650]_ ;
  assign \new_[6345]_  = \new_[651]_  | \new_[6344]_ ;
  assign \new_[6346]_  = \new_[6345]_  | \new_[6340]_ ;
  assign \new_[6347]_  = \new_[6346]_  | \new_[6337]_ ;
  assign \new_[6350]_  = \new_[647]_  | \new_[648]_ ;
  assign \new_[6354]_  = \new_[644]_  | \new_[645]_ ;
  assign \new_[6355]_  = \new_[646]_  | \new_[6354]_ ;
  assign \new_[6356]_  = \new_[6355]_  | \new_[6350]_ ;
  assign \new_[6359]_  = \new_[642]_  | \new_[643]_ ;
  assign \new_[6363]_  = \new_[639]_  | \new_[640]_ ;
  assign \new_[6364]_  = \new_[641]_  | \new_[6363]_ ;
  assign \new_[6365]_  = \new_[6364]_  | \new_[6359]_ ;
  assign \new_[6366]_  = \new_[6365]_  | \new_[6356]_ ;
  assign \new_[6367]_  = \new_[6366]_  | \new_[6347]_ ;
  assign \new_[6368]_  = \new_[6367]_  | \new_[6328]_ ;
  assign \new_[6369]_  = \new_[6368]_  | \new_[6289]_ ;
  assign \new_[6370]_  = \new_[6369]_  | \new_[6210]_ ;
  assign \new_[6371]_  = \new_[6370]_  | \new_[6051]_ ;
  assign \new_[6372]_  = \new_[6371]_  | \new_[5734]_ ;
  assign \new_[6375]_  = \new_[637]_  | \new_[638]_ ;
  assign \new_[6378]_  = \new_[635]_  | \new_[636]_ ;
  assign \new_[6379]_  = \new_[6378]_  | \new_[6375]_ ;
  assign \new_[6382]_  = \new_[633]_  | \new_[634]_ ;
  assign \new_[6386]_  = \new_[630]_  | \new_[631]_ ;
  assign \new_[6387]_  = \new_[632]_  | \new_[6386]_ ;
  assign \new_[6388]_  = \new_[6387]_  | \new_[6382]_ ;
  assign \new_[6389]_  = \new_[6388]_  | \new_[6379]_ ;
  assign \new_[6392]_  = \new_[628]_  | \new_[629]_ ;
  assign \new_[6396]_  = \new_[625]_  | \new_[626]_ ;
  assign \new_[6397]_  = \new_[627]_  | \new_[6396]_ ;
  assign \new_[6398]_  = \new_[6397]_  | \new_[6392]_ ;
  assign \new_[6401]_  = \new_[623]_  | \new_[624]_ ;
  assign \new_[6405]_  = \new_[620]_  | \new_[621]_ ;
  assign \new_[6406]_  = \new_[622]_  | \new_[6405]_ ;
  assign \new_[6407]_  = \new_[6406]_  | \new_[6401]_ ;
  assign \new_[6408]_  = \new_[6407]_  | \new_[6398]_ ;
  assign \new_[6409]_  = \new_[6408]_  | \new_[6389]_ ;
  assign \new_[6412]_  = \new_[618]_  | \new_[619]_ ;
  assign \new_[6416]_  = \new_[615]_  | \new_[616]_ ;
  assign \new_[6417]_  = \new_[617]_  | \new_[6416]_ ;
  assign \new_[6418]_  = \new_[6417]_  | \new_[6412]_ ;
  assign \new_[6421]_  = \new_[613]_  | \new_[614]_ ;
  assign \new_[6425]_  = \new_[610]_  | \new_[611]_ ;
  assign \new_[6426]_  = \new_[612]_  | \new_[6425]_ ;
  assign \new_[6427]_  = \new_[6426]_  | \new_[6421]_ ;
  assign \new_[6428]_  = \new_[6427]_  | \new_[6418]_ ;
  assign \new_[6431]_  = \new_[608]_  | \new_[609]_ ;
  assign \new_[6435]_  = \new_[605]_  | \new_[606]_ ;
  assign \new_[6436]_  = \new_[607]_  | \new_[6435]_ ;
  assign \new_[6437]_  = \new_[6436]_  | \new_[6431]_ ;
  assign \new_[6440]_  = \new_[603]_  | \new_[604]_ ;
  assign \new_[6444]_  = \new_[600]_  | \new_[601]_ ;
  assign \new_[6445]_  = \new_[602]_  | \new_[6444]_ ;
  assign \new_[6446]_  = \new_[6445]_  | \new_[6440]_ ;
  assign \new_[6447]_  = \new_[6446]_  | \new_[6437]_ ;
  assign \new_[6448]_  = \new_[6447]_  | \new_[6428]_ ;
  assign \new_[6449]_  = \new_[6448]_  | \new_[6409]_ ;
  assign \new_[6452]_  = \new_[598]_  | \new_[599]_ ;
  assign \new_[6456]_  = \new_[595]_  | \new_[596]_ ;
  assign \new_[6457]_  = \new_[597]_  | \new_[6456]_ ;
  assign \new_[6458]_  = \new_[6457]_  | \new_[6452]_ ;
  assign \new_[6461]_  = \new_[593]_  | \new_[594]_ ;
  assign \new_[6465]_  = \new_[590]_  | \new_[591]_ ;
  assign \new_[6466]_  = \new_[592]_  | \new_[6465]_ ;
  assign \new_[6467]_  = \new_[6466]_  | \new_[6461]_ ;
  assign \new_[6468]_  = \new_[6467]_  | \new_[6458]_ ;
  assign \new_[6471]_  = \new_[588]_  | \new_[589]_ ;
  assign \new_[6475]_  = \new_[585]_  | \new_[586]_ ;
  assign \new_[6476]_  = \new_[587]_  | \new_[6475]_ ;
  assign \new_[6477]_  = \new_[6476]_  | \new_[6471]_ ;
  assign \new_[6480]_  = \new_[583]_  | \new_[584]_ ;
  assign \new_[6484]_  = \new_[580]_  | \new_[581]_ ;
  assign \new_[6485]_  = \new_[582]_  | \new_[6484]_ ;
  assign \new_[6486]_  = \new_[6485]_  | \new_[6480]_ ;
  assign \new_[6487]_  = \new_[6486]_  | \new_[6477]_ ;
  assign \new_[6488]_  = \new_[6487]_  | \new_[6468]_ ;
  assign \new_[6491]_  = \new_[578]_  | \new_[579]_ ;
  assign \new_[6495]_  = \new_[575]_  | \new_[576]_ ;
  assign \new_[6496]_  = \new_[577]_  | \new_[6495]_ ;
  assign \new_[6497]_  = \new_[6496]_  | \new_[6491]_ ;
  assign \new_[6500]_  = \new_[573]_  | \new_[574]_ ;
  assign \new_[6504]_  = \new_[570]_  | \new_[571]_ ;
  assign \new_[6505]_  = \new_[572]_  | \new_[6504]_ ;
  assign \new_[6506]_  = \new_[6505]_  | \new_[6500]_ ;
  assign \new_[6507]_  = \new_[6506]_  | \new_[6497]_ ;
  assign \new_[6510]_  = \new_[568]_  | \new_[569]_ ;
  assign \new_[6514]_  = \new_[565]_  | \new_[566]_ ;
  assign \new_[6515]_  = \new_[567]_  | \new_[6514]_ ;
  assign \new_[6516]_  = \new_[6515]_  | \new_[6510]_ ;
  assign \new_[6519]_  = \new_[563]_  | \new_[564]_ ;
  assign \new_[6523]_  = \new_[560]_  | \new_[561]_ ;
  assign \new_[6524]_  = \new_[562]_  | \new_[6523]_ ;
  assign \new_[6525]_  = \new_[6524]_  | \new_[6519]_ ;
  assign \new_[6526]_  = \new_[6525]_  | \new_[6516]_ ;
  assign \new_[6527]_  = \new_[6526]_  | \new_[6507]_ ;
  assign \new_[6528]_  = \new_[6527]_  | \new_[6488]_ ;
  assign \new_[6529]_  = \new_[6528]_  | \new_[6449]_ ;
  assign \new_[6532]_  = \new_[558]_  | \new_[559]_ ;
  assign \new_[6536]_  = \new_[555]_  | \new_[556]_ ;
  assign \new_[6537]_  = \new_[557]_  | \new_[6536]_ ;
  assign \new_[6538]_  = \new_[6537]_  | \new_[6532]_ ;
  assign \new_[6541]_  = \new_[553]_  | \new_[554]_ ;
  assign \new_[6545]_  = \new_[550]_  | \new_[551]_ ;
  assign \new_[6546]_  = \new_[552]_  | \new_[6545]_ ;
  assign \new_[6547]_  = \new_[6546]_  | \new_[6541]_ ;
  assign \new_[6548]_  = \new_[6547]_  | \new_[6538]_ ;
  assign \new_[6551]_  = \new_[548]_  | \new_[549]_ ;
  assign \new_[6555]_  = \new_[545]_  | \new_[546]_ ;
  assign \new_[6556]_  = \new_[547]_  | \new_[6555]_ ;
  assign \new_[6557]_  = \new_[6556]_  | \new_[6551]_ ;
  assign \new_[6560]_  = \new_[543]_  | \new_[544]_ ;
  assign \new_[6564]_  = \new_[540]_  | \new_[541]_ ;
  assign \new_[6565]_  = \new_[542]_  | \new_[6564]_ ;
  assign \new_[6566]_  = \new_[6565]_  | \new_[6560]_ ;
  assign \new_[6567]_  = \new_[6566]_  | \new_[6557]_ ;
  assign \new_[6568]_  = \new_[6567]_  | \new_[6548]_ ;
  assign \new_[6571]_  = \new_[538]_  | \new_[539]_ ;
  assign \new_[6575]_  = \new_[535]_  | \new_[536]_ ;
  assign \new_[6576]_  = \new_[537]_  | \new_[6575]_ ;
  assign \new_[6577]_  = \new_[6576]_  | \new_[6571]_ ;
  assign \new_[6580]_  = \new_[533]_  | \new_[534]_ ;
  assign \new_[6584]_  = \new_[530]_  | \new_[531]_ ;
  assign \new_[6585]_  = \new_[532]_  | \new_[6584]_ ;
  assign \new_[6586]_  = \new_[6585]_  | \new_[6580]_ ;
  assign \new_[6587]_  = \new_[6586]_  | \new_[6577]_ ;
  assign \new_[6590]_  = \new_[528]_  | \new_[529]_ ;
  assign \new_[6594]_  = \new_[525]_  | \new_[526]_ ;
  assign \new_[6595]_  = \new_[527]_  | \new_[6594]_ ;
  assign \new_[6596]_  = \new_[6595]_  | \new_[6590]_ ;
  assign \new_[6599]_  = \new_[523]_  | \new_[524]_ ;
  assign \new_[6603]_  = \new_[520]_  | \new_[521]_ ;
  assign \new_[6604]_  = \new_[522]_  | \new_[6603]_ ;
  assign \new_[6605]_  = \new_[6604]_  | \new_[6599]_ ;
  assign \new_[6606]_  = \new_[6605]_  | \new_[6596]_ ;
  assign \new_[6607]_  = \new_[6606]_  | \new_[6587]_ ;
  assign \new_[6608]_  = \new_[6607]_  | \new_[6568]_ ;
  assign \new_[6611]_  = \new_[518]_  | \new_[519]_ ;
  assign \new_[6615]_  = \new_[515]_  | \new_[516]_ ;
  assign \new_[6616]_  = \new_[517]_  | \new_[6615]_ ;
  assign \new_[6617]_  = \new_[6616]_  | \new_[6611]_ ;
  assign \new_[6620]_  = \new_[513]_  | \new_[514]_ ;
  assign \new_[6624]_  = \new_[510]_  | \new_[511]_ ;
  assign \new_[6625]_  = \new_[512]_  | \new_[6624]_ ;
  assign \new_[6626]_  = \new_[6625]_  | \new_[6620]_ ;
  assign \new_[6627]_  = \new_[6626]_  | \new_[6617]_ ;
  assign \new_[6630]_  = \new_[508]_  | \new_[509]_ ;
  assign \new_[6634]_  = \new_[505]_  | \new_[506]_ ;
  assign \new_[6635]_  = \new_[507]_  | \new_[6634]_ ;
  assign \new_[6636]_  = \new_[6635]_  | \new_[6630]_ ;
  assign \new_[6639]_  = \new_[503]_  | \new_[504]_ ;
  assign \new_[6643]_  = \new_[500]_  | \new_[501]_ ;
  assign \new_[6644]_  = \new_[502]_  | \new_[6643]_ ;
  assign \new_[6645]_  = \new_[6644]_  | \new_[6639]_ ;
  assign \new_[6646]_  = \new_[6645]_  | \new_[6636]_ ;
  assign \new_[6647]_  = \new_[6646]_  | \new_[6627]_ ;
  assign \new_[6650]_  = \new_[498]_  | \new_[499]_ ;
  assign \new_[6654]_  = \new_[495]_  | \new_[496]_ ;
  assign \new_[6655]_  = \new_[497]_  | \new_[6654]_ ;
  assign \new_[6656]_  = \new_[6655]_  | \new_[6650]_ ;
  assign \new_[6659]_  = \new_[493]_  | \new_[494]_ ;
  assign \new_[6663]_  = \new_[490]_  | \new_[491]_ ;
  assign \new_[6664]_  = \new_[492]_  | \new_[6663]_ ;
  assign \new_[6665]_  = \new_[6664]_  | \new_[6659]_ ;
  assign \new_[6666]_  = \new_[6665]_  | \new_[6656]_ ;
  assign \new_[6669]_  = \new_[488]_  | \new_[489]_ ;
  assign \new_[6673]_  = \new_[485]_  | \new_[486]_ ;
  assign \new_[6674]_  = \new_[487]_  | \new_[6673]_ ;
  assign \new_[6675]_  = \new_[6674]_  | \new_[6669]_ ;
  assign \new_[6678]_  = \new_[483]_  | \new_[484]_ ;
  assign \new_[6682]_  = \new_[480]_  | \new_[481]_ ;
  assign \new_[6683]_  = \new_[482]_  | \new_[6682]_ ;
  assign \new_[6684]_  = \new_[6683]_  | \new_[6678]_ ;
  assign \new_[6685]_  = \new_[6684]_  | \new_[6675]_ ;
  assign \new_[6686]_  = \new_[6685]_  | \new_[6666]_ ;
  assign \new_[6687]_  = \new_[6686]_  | \new_[6647]_ ;
  assign \new_[6688]_  = \new_[6687]_  | \new_[6608]_ ;
  assign \new_[6689]_  = \new_[6688]_  | \new_[6529]_ ;
  assign \new_[6692]_  = \new_[478]_  | \new_[479]_ ;
  assign \new_[6696]_  = \new_[475]_  | \new_[476]_ ;
  assign \new_[6697]_  = \new_[477]_  | \new_[6696]_ ;
  assign \new_[6698]_  = \new_[6697]_  | \new_[6692]_ ;
  assign \new_[6701]_  = \new_[473]_  | \new_[474]_ ;
  assign \new_[6705]_  = \new_[470]_  | \new_[471]_ ;
  assign \new_[6706]_  = \new_[472]_  | \new_[6705]_ ;
  assign \new_[6707]_  = \new_[6706]_  | \new_[6701]_ ;
  assign \new_[6708]_  = \new_[6707]_  | \new_[6698]_ ;
  assign \new_[6711]_  = \new_[468]_  | \new_[469]_ ;
  assign \new_[6715]_  = \new_[465]_  | \new_[466]_ ;
  assign \new_[6716]_  = \new_[467]_  | \new_[6715]_ ;
  assign \new_[6717]_  = \new_[6716]_  | \new_[6711]_ ;
  assign \new_[6720]_  = \new_[463]_  | \new_[464]_ ;
  assign \new_[6724]_  = \new_[460]_  | \new_[461]_ ;
  assign \new_[6725]_  = \new_[462]_  | \new_[6724]_ ;
  assign \new_[6726]_  = \new_[6725]_  | \new_[6720]_ ;
  assign \new_[6727]_  = \new_[6726]_  | \new_[6717]_ ;
  assign \new_[6728]_  = \new_[6727]_  | \new_[6708]_ ;
  assign \new_[6731]_  = \new_[458]_  | \new_[459]_ ;
  assign \new_[6735]_  = \new_[455]_  | \new_[456]_ ;
  assign \new_[6736]_  = \new_[457]_  | \new_[6735]_ ;
  assign \new_[6737]_  = \new_[6736]_  | \new_[6731]_ ;
  assign \new_[6740]_  = \new_[453]_  | \new_[454]_ ;
  assign \new_[6744]_  = \new_[450]_  | \new_[451]_ ;
  assign \new_[6745]_  = \new_[452]_  | \new_[6744]_ ;
  assign \new_[6746]_  = \new_[6745]_  | \new_[6740]_ ;
  assign \new_[6747]_  = \new_[6746]_  | \new_[6737]_ ;
  assign \new_[6750]_  = \new_[448]_  | \new_[449]_ ;
  assign \new_[6754]_  = \new_[445]_  | \new_[446]_ ;
  assign \new_[6755]_  = \new_[447]_  | \new_[6754]_ ;
  assign \new_[6756]_  = \new_[6755]_  | \new_[6750]_ ;
  assign \new_[6759]_  = \new_[443]_  | \new_[444]_ ;
  assign \new_[6763]_  = \new_[440]_  | \new_[441]_ ;
  assign \new_[6764]_  = \new_[442]_  | \new_[6763]_ ;
  assign \new_[6765]_  = \new_[6764]_  | \new_[6759]_ ;
  assign \new_[6766]_  = \new_[6765]_  | \new_[6756]_ ;
  assign \new_[6767]_  = \new_[6766]_  | \new_[6747]_ ;
  assign \new_[6768]_  = \new_[6767]_  | \new_[6728]_ ;
  assign \new_[6771]_  = \new_[438]_  | \new_[439]_ ;
  assign \new_[6775]_  = \new_[435]_  | \new_[436]_ ;
  assign \new_[6776]_  = \new_[437]_  | \new_[6775]_ ;
  assign \new_[6777]_  = \new_[6776]_  | \new_[6771]_ ;
  assign \new_[6780]_  = \new_[433]_  | \new_[434]_ ;
  assign \new_[6784]_  = \new_[430]_  | \new_[431]_ ;
  assign \new_[6785]_  = \new_[432]_  | \new_[6784]_ ;
  assign \new_[6786]_  = \new_[6785]_  | \new_[6780]_ ;
  assign \new_[6787]_  = \new_[6786]_  | \new_[6777]_ ;
  assign \new_[6790]_  = \new_[428]_  | \new_[429]_ ;
  assign \new_[6794]_  = \new_[425]_  | \new_[426]_ ;
  assign \new_[6795]_  = \new_[427]_  | \new_[6794]_ ;
  assign \new_[6796]_  = \new_[6795]_  | \new_[6790]_ ;
  assign \new_[6799]_  = \new_[423]_  | \new_[424]_ ;
  assign \new_[6803]_  = \new_[420]_  | \new_[421]_ ;
  assign \new_[6804]_  = \new_[422]_  | \new_[6803]_ ;
  assign \new_[6805]_  = \new_[6804]_  | \new_[6799]_ ;
  assign \new_[6806]_  = \new_[6805]_  | \new_[6796]_ ;
  assign \new_[6807]_  = \new_[6806]_  | \new_[6787]_ ;
  assign \new_[6810]_  = \new_[418]_  | \new_[419]_ ;
  assign \new_[6814]_  = \new_[415]_  | \new_[416]_ ;
  assign \new_[6815]_  = \new_[417]_  | \new_[6814]_ ;
  assign \new_[6816]_  = \new_[6815]_  | \new_[6810]_ ;
  assign \new_[6819]_  = \new_[413]_  | \new_[414]_ ;
  assign \new_[6823]_  = \new_[410]_  | \new_[411]_ ;
  assign \new_[6824]_  = \new_[412]_  | \new_[6823]_ ;
  assign \new_[6825]_  = \new_[6824]_  | \new_[6819]_ ;
  assign \new_[6826]_  = \new_[6825]_  | \new_[6816]_ ;
  assign \new_[6829]_  = \new_[408]_  | \new_[409]_ ;
  assign \new_[6833]_  = \new_[405]_  | \new_[406]_ ;
  assign \new_[6834]_  = \new_[407]_  | \new_[6833]_ ;
  assign \new_[6835]_  = \new_[6834]_  | \new_[6829]_ ;
  assign \new_[6838]_  = \new_[403]_  | \new_[404]_ ;
  assign \new_[6842]_  = \new_[400]_  | \new_[401]_ ;
  assign \new_[6843]_  = \new_[402]_  | \new_[6842]_ ;
  assign \new_[6844]_  = \new_[6843]_  | \new_[6838]_ ;
  assign \new_[6845]_  = \new_[6844]_  | \new_[6835]_ ;
  assign \new_[6846]_  = \new_[6845]_  | \new_[6826]_ ;
  assign \new_[6847]_  = \new_[6846]_  | \new_[6807]_ ;
  assign \new_[6848]_  = \new_[6847]_  | \new_[6768]_ ;
  assign \new_[6851]_  = \new_[398]_  | \new_[399]_ ;
  assign \new_[6855]_  = \new_[395]_  | \new_[396]_ ;
  assign \new_[6856]_  = \new_[397]_  | \new_[6855]_ ;
  assign \new_[6857]_  = \new_[6856]_  | \new_[6851]_ ;
  assign \new_[6860]_  = \new_[393]_  | \new_[394]_ ;
  assign \new_[6864]_  = \new_[390]_  | \new_[391]_ ;
  assign \new_[6865]_  = \new_[392]_  | \new_[6864]_ ;
  assign \new_[6866]_  = \new_[6865]_  | \new_[6860]_ ;
  assign \new_[6867]_  = \new_[6866]_  | \new_[6857]_ ;
  assign \new_[6870]_  = \new_[388]_  | \new_[389]_ ;
  assign \new_[6874]_  = \new_[385]_  | \new_[386]_ ;
  assign \new_[6875]_  = \new_[387]_  | \new_[6874]_ ;
  assign \new_[6876]_  = \new_[6875]_  | \new_[6870]_ ;
  assign \new_[6879]_  = \new_[383]_  | \new_[384]_ ;
  assign \new_[6883]_  = \new_[380]_  | \new_[381]_ ;
  assign \new_[6884]_  = \new_[382]_  | \new_[6883]_ ;
  assign \new_[6885]_  = \new_[6884]_  | \new_[6879]_ ;
  assign \new_[6886]_  = \new_[6885]_  | \new_[6876]_ ;
  assign \new_[6887]_  = \new_[6886]_  | \new_[6867]_ ;
  assign \new_[6890]_  = \new_[378]_  | \new_[379]_ ;
  assign \new_[6894]_  = \new_[375]_  | \new_[376]_ ;
  assign \new_[6895]_  = \new_[377]_  | \new_[6894]_ ;
  assign \new_[6896]_  = \new_[6895]_  | \new_[6890]_ ;
  assign \new_[6899]_  = \new_[373]_  | \new_[374]_ ;
  assign \new_[6903]_  = \new_[370]_  | \new_[371]_ ;
  assign \new_[6904]_  = \new_[372]_  | \new_[6903]_ ;
  assign \new_[6905]_  = \new_[6904]_  | \new_[6899]_ ;
  assign \new_[6906]_  = \new_[6905]_  | \new_[6896]_ ;
  assign \new_[6909]_  = \new_[368]_  | \new_[369]_ ;
  assign \new_[6913]_  = \new_[365]_  | \new_[366]_ ;
  assign \new_[6914]_  = \new_[367]_  | \new_[6913]_ ;
  assign \new_[6915]_  = \new_[6914]_  | \new_[6909]_ ;
  assign \new_[6918]_  = \new_[363]_  | \new_[364]_ ;
  assign \new_[6922]_  = \new_[360]_  | \new_[361]_ ;
  assign \new_[6923]_  = \new_[362]_  | \new_[6922]_ ;
  assign \new_[6924]_  = \new_[6923]_  | \new_[6918]_ ;
  assign \new_[6925]_  = \new_[6924]_  | \new_[6915]_ ;
  assign \new_[6926]_  = \new_[6925]_  | \new_[6906]_ ;
  assign \new_[6927]_  = \new_[6926]_  | \new_[6887]_ ;
  assign \new_[6930]_  = \new_[358]_  | \new_[359]_ ;
  assign \new_[6934]_  = \new_[355]_  | \new_[356]_ ;
  assign \new_[6935]_  = \new_[357]_  | \new_[6934]_ ;
  assign \new_[6936]_  = \new_[6935]_  | \new_[6930]_ ;
  assign \new_[6939]_  = \new_[353]_  | \new_[354]_ ;
  assign \new_[6943]_  = \new_[350]_  | \new_[351]_ ;
  assign \new_[6944]_  = \new_[352]_  | \new_[6943]_ ;
  assign \new_[6945]_  = \new_[6944]_  | \new_[6939]_ ;
  assign \new_[6946]_  = \new_[6945]_  | \new_[6936]_ ;
  assign \new_[6949]_  = \new_[348]_  | \new_[349]_ ;
  assign \new_[6953]_  = \new_[345]_  | \new_[346]_ ;
  assign \new_[6954]_  = \new_[347]_  | \new_[6953]_ ;
  assign \new_[6955]_  = \new_[6954]_  | \new_[6949]_ ;
  assign \new_[6958]_  = \new_[343]_  | \new_[344]_ ;
  assign \new_[6962]_  = \new_[340]_  | \new_[341]_ ;
  assign \new_[6963]_  = \new_[342]_  | \new_[6962]_ ;
  assign \new_[6964]_  = \new_[6963]_  | \new_[6958]_ ;
  assign \new_[6965]_  = \new_[6964]_  | \new_[6955]_ ;
  assign \new_[6966]_  = \new_[6965]_  | \new_[6946]_ ;
  assign \new_[6969]_  = \new_[338]_  | \new_[339]_ ;
  assign \new_[6973]_  = \new_[335]_  | \new_[336]_ ;
  assign \new_[6974]_  = \new_[337]_  | \new_[6973]_ ;
  assign \new_[6975]_  = \new_[6974]_  | \new_[6969]_ ;
  assign \new_[6978]_  = \new_[333]_  | \new_[334]_ ;
  assign \new_[6982]_  = \new_[330]_  | \new_[331]_ ;
  assign \new_[6983]_  = \new_[332]_  | \new_[6982]_ ;
  assign \new_[6984]_  = \new_[6983]_  | \new_[6978]_ ;
  assign \new_[6985]_  = \new_[6984]_  | \new_[6975]_ ;
  assign \new_[6988]_  = \new_[328]_  | \new_[329]_ ;
  assign \new_[6992]_  = \new_[325]_  | \new_[326]_ ;
  assign \new_[6993]_  = \new_[327]_  | \new_[6992]_ ;
  assign \new_[6994]_  = \new_[6993]_  | \new_[6988]_ ;
  assign \new_[6997]_  = \new_[323]_  | \new_[324]_ ;
  assign \new_[7001]_  = \new_[320]_  | \new_[321]_ ;
  assign \new_[7002]_  = \new_[322]_  | \new_[7001]_ ;
  assign \new_[7003]_  = \new_[7002]_  | \new_[6997]_ ;
  assign \new_[7004]_  = \new_[7003]_  | \new_[6994]_ ;
  assign \new_[7005]_  = \new_[7004]_  | \new_[6985]_ ;
  assign \new_[7006]_  = \new_[7005]_  | \new_[6966]_ ;
  assign \new_[7007]_  = \new_[7006]_  | \new_[6927]_ ;
  assign \new_[7008]_  = \new_[7007]_  | \new_[6848]_ ;
  assign \new_[7009]_  = \new_[7008]_  | \new_[6689]_ ;
  assign \new_[7012]_  = \new_[318]_  | \new_[319]_ ;
  assign \new_[7015]_  = \new_[316]_  | \new_[317]_ ;
  assign \new_[7016]_  = \new_[7015]_  | \new_[7012]_ ;
  assign \new_[7019]_  = \new_[314]_  | \new_[315]_ ;
  assign \new_[7023]_  = \new_[311]_  | \new_[312]_ ;
  assign \new_[7024]_  = \new_[313]_  | \new_[7023]_ ;
  assign \new_[7025]_  = \new_[7024]_  | \new_[7019]_ ;
  assign \new_[7026]_  = \new_[7025]_  | \new_[7016]_ ;
  assign \new_[7029]_  = \new_[309]_  | \new_[310]_ ;
  assign \new_[7033]_  = \new_[306]_  | \new_[307]_ ;
  assign \new_[7034]_  = \new_[308]_  | \new_[7033]_ ;
  assign \new_[7035]_  = \new_[7034]_  | \new_[7029]_ ;
  assign \new_[7038]_  = \new_[304]_  | \new_[305]_ ;
  assign \new_[7042]_  = \new_[301]_  | \new_[302]_ ;
  assign \new_[7043]_  = \new_[303]_  | \new_[7042]_ ;
  assign \new_[7044]_  = \new_[7043]_  | \new_[7038]_ ;
  assign \new_[7045]_  = \new_[7044]_  | \new_[7035]_ ;
  assign \new_[7046]_  = \new_[7045]_  | \new_[7026]_ ;
  assign \new_[7049]_  = \new_[299]_  | \new_[300]_ ;
  assign \new_[7053]_  = \new_[296]_  | \new_[297]_ ;
  assign \new_[7054]_  = \new_[298]_  | \new_[7053]_ ;
  assign \new_[7055]_  = \new_[7054]_  | \new_[7049]_ ;
  assign \new_[7058]_  = \new_[294]_  | \new_[295]_ ;
  assign \new_[7062]_  = \new_[291]_  | \new_[292]_ ;
  assign \new_[7063]_  = \new_[293]_  | \new_[7062]_ ;
  assign \new_[7064]_  = \new_[7063]_  | \new_[7058]_ ;
  assign \new_[7065]_  = \new_[7064]_  | \new_[7055]_ ;
  assign \new_[7068]_  = \new_[289]_  | \new_[290]_ ;
  assign \new_[7072]_  = \new_[286]_  | \new_[287]_ ;
  assign \new_[7073]_  = \new_[288]_  | \new_[7072]_ ;
  assign \new_[7074]_  = \new_[7073]_  | \new_[7068]_ ;
  assign \new_[7077]_  = \new_[284]_  | \new_[285]_ ;
  assign \new_[7081]_  = \new_[281]_  | \new_[282]_ ;
  assign \new_[7082]_  = \new_[283]_  | \new_[7081]_ ;
  assign \new_[7083]_  = \new_[7082]_  | \new_[7077]_ ;
  assign \new_[7084]_  = \new_[7083]_  | \new_[7074]_ ;
  assign \new_[7085]_  = \new_[7084]_  | \new_[7065]_ ;
  assign \new_[7086]_  = \new_[7085]_  | \new_[7046]_ ;
  assign \new_[7089]_  = \new_[279]_  | \new_[280]_ ;
  assign \new_[7093]_  = \new_[276]_  | \new_[277]_ ;
  assign \new_[7094]_  = \new_[278]_  | \new_[7093]_ ;
  assign \new_[7095]_  = \new_[7094]_  | \new_[7089]_ ;
  assign \new_[7098]_  = \new_[274]_  | \new_[275]_ ;
  assign \new_[7102]_  = \new_[271]_  | \new_[272]_ ;
  assign \new_[7103]_  = \new_[273]_  | \new_[7102]_ ;
  assign \new_[7104]_  = \new_[7103]_  | \new_[7098]_ ;
  assign \new_[7105]_  = \new_[7104]_  | \new_[7095]_ ;
  assign \new_[7108]_  = \new_[269]_  | \new_[270]_ ;
  assign \new_[7112]_  = \new_[266]_  | \new_[267]_ ;
  assign \new_[7113]_  = \new_[268]_  | \new_[7112]_ ;
  assign \new_[7114]_  = \new_[7113]_  | \new_[7108]_ ;
  assign \new_[7117]_  = \new_[264]_  | \new_[265]_ ;
  assign \new_[7121]_  = \new_[261]_  | \new_[262]_ ;
  assign \new_[7122]_  = \new_[263]_  | \new_[7121]_ ;
  assign \new_[7123]_  = \new_[7122]_  | \new_[7117]_ ;
  assign \new_[7124]_  = \new_[7123]_  | \new_[7114]_ ;
  assign \new_[7125]_  = \new_[7124]_  | \new_[7105]_ ;
  assign \new_[7128]_  = \new_[259]_  | \new_[260]_ ;
  assign \new_[7132]_  = \new_[256]_  | \new_[257]_ ;
  assign \new_[7133]_  = \new_[258]_  | \new_[7132]_ ;
  assign \new_[7134]_  = \new_[7133]_  | \new_[7128]_ ;
  assign \new_[7137]_  = \new_[254]_  | \new_[255]_ ;
  assign \new_[7141]_  = \new_[251]_  | \new_[252]_ ;
  assign \new_[7142]_  = \new_[253]_  | \new_[7141]_ ;
  assign \new_[7143]_  = \new_[7142]_  | \new_[7137]_ ;
  assign \new_[7144]_  = \new_[7143]_  | \new_[7134]_ ;
  assign \new_[7147]_  = \new_[249]_  | \new_[250]_ ;
  assign \new_[7151]_  = \new_[246]_  | \new_[247]_ ;
  assign \new_[7152]_  = \new_[248]_  | \new_[7151]_ ;
  assign \new_[7153]_  = \new_[7152]_  | \new_[7147]_ ;
  assign \new_[7156]_  = \new_[244]_  | \new_[245]_ ;
  assign \new_[7160]_  = \new_[241]_  | \new_[242]_ ;
  assign \new_[7161]_  = \new_[243]_  | \new_[7160]_ ;
  assign \new_[7162]_  = \new_[7161]_  | \new_[7156]_ ;
  assign \new_[7163]_  = \new_[7162]_  | \new_[7153]_ ;
  assign \new_[7164]_  = \new_[7163]_  | \new_[7144]_ ;
  assign \new_[7165]_  = \new_[7164]_  | \new_[7125]_ ;
  assign \new_[7166]_  = \new_[7165]_  | \new_[7086]_ ;
  assign \new_[7169]_  = \new_[239]_  | \new_[240]_ ;
  assign \new_[7173]_  = \new_[236]_  | \new_[237]_ ;
  assign \new_[7174]_  = \new_[238]_  | \new_[7173]_ ;
  assign \new_[7175]_  = \new_[7174]_  | \new_[7169]_ ;
  assign \new_[7178]_  = \new_[234]_  | \new_[235]_ ;
  assign \new_[7182]_  = \new_[231]_  | \new_[232]_ ;
  assign \new_[7183]_  = \new_[233]_  | \new_[7182]_ ;
  assign \new_[7184]_  = \new_[7183]_  | \new_[7178]_ ;
  assign \new_[7185]_  = \new_[7184]_  | \new_[7175]_ ;
  assign \new_[7188]_  = \new_[229]_  | \new_[230]_ ;
  assign \new_[7192]_  = \new_[226]_  | \new_[227]_ ;
  assign \new_[7193]_  = \new_[228]_  | \new_[7192]_ ;
  assign \new_[7194]_  = \new_[7193]_  | \new_[7188]_ ;
  assign \new_[7197]_  = \new_[224]_  | \new_[225]_ ;
  assign \new_[7201]_  = \new_[221]_  | \new_[222]_ ;
  assign \new_[7202]_  = \new_[223]_  | \new_[7201]_ ;
  assign \new_[7203]_  = \new_[7202]_  | \new_[7197]_ ;
  assign \new_[7204]_  = \new_[7203]_  | \new_[7194]_ ;
  assign \new_[7205]_  = \new_[7204]_  | \new_[7185]_ ;
  assign \new_[7208]_  = \new_[219]_  | \new_[220]_ ;
  assign \new_[7212]_  = \new_[216]_  | \new_[217]_ ;
  assign \new_[7213]_  = \new_[218]_  | \new_[7212]_ ;
  assign \new_[7214]_  = \new_[7213]_  | \new_[7208]_ ;
  assign \new_[7217]_  = \new_[214]_  | \new_[215]_ ;
  assign \new_[7221]_  = \new_[211]_  | \new_[212]_ ;
  assign \new_[7222]_  = \new_[213]_  | \new_[7221]_ ;
  assign \new_[7223]_  = \new_[7222]_  | \new_[7217]_ ;
  assign \new_[7224]_  = \new_[7223]_  | \new_[7214]_ ;
  assign \new_[7227]_  = \new_[209]_  | \new_[210]_ ;
  assign \new_[7231]_  = \new_[206]_  | \new_[207]_ ;
  assign \new_[7232]_  = \new_[208]_  | \new_[7231]_ ;
  assign \new_[7233]_  = \new_[7232]_  | \new_[7227]_ ;
  assign \new_[7236]_  = \new_[204]_  | \new_[205]_ ;
  assign \new_[7240]_  = \new_[201]_  | \new_[202]_ ;
  assign \new_[7241]_  = \new_[203]_  | \new_[7240]_ ;
  assign \new_[7242]_  = \new_[7241]_  | \new_[7236]_ ;
  assign \new_[7243]_  = \new_[7242]_  | \new_[7233]_ ;
  assign \new_[7244]_  = \new_[7243]_  | \new_[7224]_ ;
  assign \new_[7245]_  = \new_[7244]_  | \new_[7205]_ ;
  assign \new_[7248]_  = \new_[199]_  | \new_[200]_ ;
  assign \new_[7252]_  = \new_[196]_  | \new_[197]_ ;
  assign \new_[7253]_  = \new_[198]_  | \new_[7252]_ ;
  assign \new_[7254]_  = \new_[7253]_  | \new_[7248]_ ;
  assign \new_[7257]_  = \new_[194]_  | \new_[195]_ ;
  assign \new_[7261]_  = \new_[191]_  | \new_[192]_ ;
  assign \new_[7262]_  = \new_[193]_  | \new_[7261]_ ;
  assign \new_[7263]_  = \new_[7262]_  | \new_[7257]_ ;
  assign \new_[7264]_  = \new_[7263]_  | \new_[7254]_ ;
  assign \new_[7267]_  = \new_[189]_  | \new_[190]_ ;
  assign \new_[7271]_  = \new_[186]_  | \new_[187]_ ;
  assign \new_[7272]_  = \new_[188]_  | \new_[7271]_ ;
  assign \new_[7273]_  = \new_[7272]_  | \new_[7267]_ ;
  assign \new_[7276]_  = \new_[184]_  | \new_[185]_ ;
  assign \new_[7280]_  = \new_[181]_  | \new_[182]_ ;
  assign \new_[7281]_  = \new_[183]_  | \new_[7280]_ ;
  assign \new_[7282]_  = \new_[7281]_  | \new_[7276]_ ;
  assign \new_[7283]_  = \new_[7282]_  | \new_[7273]_ ;
  assign \new_[7284]_  = \new_[7283]_  | \new_[7264]_ ;
  assign \new_[7287]_  = \new_[179]_  | \new_[180]_ ;
  assign \new_[7291]_  = \new_[176]_  | \new_[177]_ ;
  assign \new_[7292]_  = \new_[178]_  | \new_[7291]_ ;
  assign \new_[7293]_  = \new_[7292]_  | \new_[7287]_ ;
  assign \new_[7296]_  = \new_[174]_  | \new_[175]_ ;
  assign \new_[7300]_  = \new_[171]_  | \new_[172]_ ;
  assign \new_[7301]_  = \new_[173]_  | \new_[7300]_ ;
  assign \new_[7302]_  = \new_[7301]_  | \new_[7296]_ ;
  assign \new_[7303]_  = \new_[7302]_  | \new_[7293]_ ;
  assign \new_[7306]_  = \new_[169]_  | \new_[170]_ ;
  assign \new_[7310]_  = \new_[166]_  | \new_[167]_ ;
  assign \new_[7311]_  = \new_[168]_  | \new_[7310]_ ;
  assign \new_[7312]_  = \new_[7311]_  | \new_[7306]_ ;
  assign \new_[7315]_  = \new_[164]_  | \new_[165]_ ;
  assign \new_[7319]_  = \new_[161]_  | \new_[162]_ ;
  assign \new_[7320]_  = \new_[163]_  | \new_[7319]_ ;
  assign \new_[7321]_  = \new_[7320]_  | \new_[7315]_ ;
  assign \new_[7322]_  = \new_[7321]_  | \new_[7312]_ ;
  assign \new_[7323]_  = \new_[7322]_  | \new_[7303]_ ;
  assign \new_[7324]_  = \new_[7323]_  | \new_[7284]_ ;
  assign \new_[7325]_  = \new_[7324]_  | \new_[7245]_ ;
  assign \new_[7326]_  = \new_[7325]_  | \new_[7166]_ ;
  assign \new_[7329]_  = \new_[159]_  | \new_[160]_ ;
  assign \new_[7333]_  = \new_[156]_  | \new_[157]_ ;
  assign \new_[7334]_  = \new_[158]_  | \new_[7333]_ ;
  assign \new_[7335]_  = \new_[7334]_  | \new_[7329]_ ;
  assign \new_[7338]_  = \new_[154]_  | \new_[155]_ ;
  assign \new_[7342]_  = \new_[151]_  | \new_[152]_ ;
  assign \new_[7343]_  = \new_[153]_  | \new_[7342]_ ;
  assign \new_[7344]_  = \new_[7343]_  | \new_[7338]_ ;
  assign \new_[7345]_  = \new_[7344]_  | \new_[7335]_ ;
  assign \new_[7348]_  = \new_[149]_  | \new_[150]_ ;
  assign \new_[7352]_  = \new_[146]_  | \new_[147]_ ;
  assign \new_[7353]_  = \new_[148]_  | \new_[7352]_ ;
  assign \new_[7354]_  = \new_[7353]_  | \new_[7348]_ ;
  assign \new_[7357]_  = \new_[144]_  | \new_[145]_ ;
  assign \new_[7361]_  = \new_[141]_  | \new_[142]_ ;
  assign \new_[7362]_  = \new_[143]_  | \new_[7361]_ ;
  assign \new_[7363]_  = \new_[7362]_  | \new_[7357]_ ;
  assign \new_[7364]_  = \new_[7363]_  | \new_[7354]_ ;
  assign \new_[7365]_  = \new_[7364]_  | \new_[7345]_ ;
  assign \new_[7368]_  = \new_[139]_  | \new_[140]_ ;
  assign \new_[7372]_  = \new_[136]_  | \new_[137]_ ;
  assign \new_[7373]_  = \new_[138]_  | \new_[7372]_ ;
  assign \new_[7374]_  = \new_[7373]_  | \new_[7368]_ ;
  assign \new_[7377]_  = \new_[134]_  | \new_[135]_ ;
  assign \new_[7381]_  = \new_[131]_  | \new_[132]_ ;
  assign \new_[7382]_  = \new_[133]_  | \new_[7381]_ ;
  assign \new_[7383]_  = \new_[7382]_  | \new_[7377]_ ;
  assign \new_[7384]_  = \new_[7383]_  | \new_[7374]_ ;
  assign \new_[7387]_  = \new_[129]_  | \new_[130]_ ;
  assign \new_[7391]_  = \new_[126]_  | \new_[127]_ ;
  assign \new_[7392]_  = \new_[128]_  | \new_[7391]_ ;
  assign \new_[7393]_  = \new_[7392]_  | \new_[7387]_ ;
  assign \new_[7396]_  = \new_[124]_  | \new_[125]_ ;
  assign \new_[7400]_  = \new_[121]_  | \new_[122]_ ;
  assign \new_[7401]_  = \new_[123]_  | \new_[7400]_ ;
  assign \new_[7402]_  = \new_[7401]_  | \new_[7396]_ ;
  assign \new_[7403]_  = \new_[7402]_  | \new_[7393]_ ;
  assign \new_[7404]_  = \new_[7403]_  | \new_[7384]_ ;
  assign \new_[7405]_  = \new_[7404]_  | \new_[7365]_ ;
  assign \new_[7408]_  = \new_[119]_  | \new_[120]_ ;
  assign \new_[7412]_  = \new_[116]_  | \new_[117]_ ;
  assign \new_[7413]_  = \new_[118]_  | \new_[7412]_ ;
  assign \new_[7414]_  = \new_[7413]_  | \new_[7408]_ ;
  assign \new_[7417]_  = \new_[114]_  | \new_[115]_ ;
  assign \new_[7421]_  = \new_[111]_  | \new_[112]_ ;
  assign \new_[7422]_  = \new_[113]_  | \new_[7421]_ ;
  assign \new_[7423]_  = \new_[7422]_  | \new_[7417]_ ;
  assign \new_[7424]_  = \new_[7423]_  | \new_[7414]_ ;
  assign \new_[7427]_  = \new_[109]_  | \new_[110]_ ;
  assign \new_[7431]_  = \new_[106]_  | \new_[107]_ ;
  assign \new_[7432]_  = \new_[108]_  | \new_[7431]_ ;
  assign \new_[7433]_  = \new_[7432]_  | \new_[7427]_ ;
  assign \new_[7436]_  = \new_[104]_  | \new_[105]_ ;
  assign \new_[7440]_  = \new_[101]_  | \new_[102]_ ;
  assign \new_[7441]_  = \new_[103]_  | \new_[7440]_ ;
  assign \new_[7442]_  = \new_[7441]_  | \new_[7436]_ ;
  assign \new_[7443]_  = \new_[7442]_  | \new_[7433]_ ;
  assign \new_[7444]_  = \new_[7443]_  | \new_[7424]_ ;
  assign \new_[7447]_  = \new_[99]_  | \new_[100]_ ;
  assign \new_[7451]_  = \new_[96]_  | \new_[97]_ ;
  assign \new_[7452]_  = \new_[98]_  | \new_[7451]_ ;
  assign \new_[7453]_  = \new_[7452]_  | \new_[7447]_ ;
  assign \new_[7456]_  = \new_[94]_  | \new_[95]_ ;
  assign \new_[7460]_  = \new_[91]_  | \new_[92]_ ;
  assign \new_[7461]_  = \new_[93]_  | \new_[7460]_ ;
  assign \new_[7462]_  = \new_[7461]_  | \new_[7456]_ ;
  assign \new_[7463]_  = \new_[7462]_  | \new_[7453]_ ;
  assign \new_[7466]_  = \new_[89]_  | \new_[90]_ ;
  assign \new_[7470]_  = \new_[86]_  | \new_[87]_ ;
  assign \new_[7471]_  = \new_[88]_  | \new_[7470]_ ;
  assign \new_[7472]_  = \new_[7471]_  | \new_[7466]_ ;
  assign \new_[7475]_  = \new_[84]_  | \new_[85]_ ;
  assign \new_[7479]_  = \new_[81]_  | \new_[82]_ ;
  assign \new_[7480]_  = \new_[83]_  | \new_[7479]_ ;
  assign \new_[7481]_  = \new_[7480]_  | \new_[7475]_ ;
  assign \new_[7482]_  = \new_[7481]_  | \new_[7472]_ ;
  assign \new_[7483]_  = \new_[7482]_  | \new_[7463]_ ;
  assign \new_[7484]_  = \new_[7483]_  | \new_[7444]_ ;
  assign \new_[7485]_  = \new_[7484]_  | \new_[7405]_ ;
  assign \new_[7488]_  = \new_[79]_  | \new_[80]_ ;
  assign \new_[7492]_  = \new_[76]_  | \new_[77]_ ;
  assign \new_[7493]_  = \new_[78]_  | \new_[7492]_ ;
  assign \new_[7494]_  = \new_[7493]_  | \new_[7488]_ ;
  assign \new_[7497]_  = \new_[74]_  | \new_[75]_ ;
  assign \new_[7501]_  = \new_[71]_  | \new_[72]_ ;
  assign \new_[7502]_  = \new_[73]_  | \new_[7501]_ ;
  assign \new_[7503]_  = \new_[7502]_  | \new_[7497]_ ;
  assign \new_[7504]_  = \new_[7503]_  | \new_[7494]_ ;
  assign \new_[7507]_  = \new_[69]_  | \new_[70]_ ;
  assign \new_[7511]_  = \new_[66]_  | \new_[67]_ ;
  assign \new_[7512]_  = \new_[68]_  | \new_[7511]_ ;
  assign \new_[7513]_  = \new_[7512]_  | \new_[7507]_ ;
  assign \new_[7516]_  = \new_[64]_  | \new_[65]_ ;
  assign \new_[7520]_  = \new_[61]_  | \new_[62]_ ;
  assign \new_[7521]_  = \new_[63]_  | \new_[7520]_ ;
  assign \new_[7522]_  = \new_[7521]_  | \new_[7516]_ ;
  assign \new_[7523]_  = \new_[7522]_  | \new_[7513]_ ;
  assign \new_[7524]_  = \new_[7523]_  | \new_[7504]_ ;
  assign \new_[7527]_  = \new_[59]_  | \new_[60]_ ;
  assign \new_[7531]_  = \new_[56]_  | \new_[57]_ ;
  assign \new_[7532]_  = \new_[58]_  | \new_[7531]_ ;
  assign \new_[7533]_  = \new_[7532]_  | \new_[7527]_ ;
  assign \new_[7536]_  = \new_[54]_  | \new_[55]_ ;
  assign \new_[7540]_  = \new_[51]_  | \new_[52]_ ;
  assign \new_[7541]_  = \new_[53]_  | \new_[7540]_ ;
  assign \new_[7542]_  = \new_[7541]_  | \new_[7536]_ ;
  assign \new_[7543]_  = \new_[7542]_  | \new_[7533]_ ;
  assign \new_[7546]_  = \new_[49]_  | \new_[50]_ ;
  assign \new_[7550]_  = \new_[46]_  | \new_[47]_ ;
  assign \new_[7551]_  = \new_[48]_  | \new_[7550]_ ;
  assign \new_[7552]_  = \new_[7551]_  | \new_[7546]_ ;
  assign \new_[7555]_  = \new_[44]_  | \new_[45]_ ;
  assign \new_[7559]_  = \new_[41]_  | \new_[42]_ ;
  assign \new_[7560]_  = \new_[43]_  | \new_[7559]_ ;
  assign \new_[7561]_  = \new_[7560]_  | \new_[7555]_ ;
  assign \new_[7562]_  = \new_[7561]_  | \new_[7552]_ ;
  assign \new_[7563]_  = \new_[7562]_  | \new_[7543]_ ;
  assign \new_[7564]_  = \new_[7563]_  | \new_[7524]_ ;
  assign \new_[7567]_  = \new_[39]_  | \new_[40]_ ;
  assign \new_[7571]_  = \new_[36]_  | \new_[37]_ ;
  assign \new_[7572]_  = \new_[38]_  | \new_[7571]_ ;
  assign \new_[7573]_  = \new_[7572]_  | \new_[7567]_ ;
  assign \new_[7576]_  = \new_[34]_  | \new_[35]_ ;
  assign \new_[7580]_  = \new_[31]_  | \new_[32]_ ;
  assign \new_[7581]_  = \new_[33]_  | \new_[7580]_ ;
  assign \new_[7582]_  = \new_[7581]_  | \new_[7576]_ ;
  assign \new_[7583]_  = \new_[7582]_  | \new_[7573]_ ;
  assign \new_[7586]_  = \new_[29]_  | \new_[30]_ ;
  assign \new_[7590]_  = \new_[26]_  | \new_[27]_ ;
  assign \new_[7591]_  = \new_[28]_  | \new_[7590]_ ;
  assign \new_[7592]_  = \new_[7591]_  | \new_[7586]_ ;
  assign \new_[7595]_  = \new_[24]_  | \new_[25]_ ;
  assign \new_[7599]_  = \new_[21]_  | \new_[22]_ ;
  assign \new_[7600]_  = \new_[23]_  | \new_[7599]_ ;
  assign \new_[7601]_  = \new_[7600]_  | \new_[7595]_ ;
  assign \new_[7602]_  = \new_[7601]_  | \new_[7592]_ ;
  assign \new_[7603]_  = \new_[7602]_  | \new_[7583]_ ;
  assign \new_[7606]_  = \new_[19]_  | \new_[20]_ ;
  assign \new_[7610]_  = \new_[16]_  | \new_[17]_ ;
  assign \new_[7611]_  = \new_[18]_  | \new_[7610]_ ;
  assign \new_[7612]_  = \new_[7611]_  | \new_[7606]_ ;
  assign \new_[7615]_  = \new_[14]_  | \new_[15]_ ;
  assign \new_[7619]_  = \new_[11]_  | \new_[12]_ ;
  assign \new_[7620]_  = \new_[13]_  | \new_[7619]_ ;
  assign \new_[7621]_  = \new_[7620]_  | \new_[7615]_ ;
  assign \new_[7622]_  = \new_[7621]_  | \new_[7612]_ ;
  assign \new_[7625]_  = \new_[9]_  | \new_[10]_ ;
  assign \new_[7629]_  = \new_[6]_  | \new_[7]_ ;
  assign \new_[7630]_  = \new_[8]_  | \new_[7629]_ ;
  assign \new_[7631]_  = \new_[7630]_  | \new_[7625]_ ;
  assign \new_[7634]_  = \new_[4]_  | \new_[5]_ ;
  assign \new_[7638]_  = \new_[1]_  | \new_[2]_ ;
  assign \new_[7639]_  = \new_[3]_  | \new_[7638]_ ;
  assign \new_[7640]_  = \new_[7639]_  | \new_[7634]_ ;
  assign \new_[7641]_  = \new_[7640]_  | \new_[7631]_ ;
  assign \new_[7642]_  = \new_[7641]_  | \new_[7622]_ ;
  assign \new_[7643]_  = \new_[7642]_  | \new_[7603]_ ;
  assign \new_[7644]_  = \new_[7643]_  | \new_[7564]_ ;
  assign \new_[7645]_  = \new_[7644]_  | \new_[7485]_ ;
  assign \new_[7646]_  = \new_[7645]_  | \new_[7326]_ ;
  assign \new_[7647]_  = \new_[7646]_  | \new_[7009]_ ;
  assign \new_[7648]_  = \new_[7647]_  | \new_[6372]_ ;
  assign \new_[7652]_  = ~A202 & ~A201;
  assign \new_[7653]_  = A169 & \new_[7652]_ ;
  assign \new_[7657]_  = A268 & A235;
  assign \new_[7658]_  = ~A203 & \new_[7657]_ ;
  assign \new_[7662]_  = ~A200 & ~A199;
  assign \new_[7663]_  = A169 & \new_[7662]_ ;
  assign \new_[7667]_  = A268 & A235;
  assign \new_[7668]_  = ~A202 & \new_[7667]_ ;
  assign \new_[7672]_  = ~A166 & ~A167;
  assign \new_[7673]_  = ~A169 & \new_[7672]_ ;
  assign \new_[7677]_  = A268 & A235;
  assign \new_[7678]_  = A202 & \new_[7677]_ ;
  assign \new_[7682]_  = ~A168 & ~A169;
  assign \new_[7683]_  = ~A170 & \new_[7682]_ ;
  assign \new_[7687]_  = A268 & A235;
  assign \new_[7688]_  = A202 & \new_[7687]_ ;
  assign \new_[7692]_  = ~A201 & A166;
  assign \new_[7693]_  = A168 & \new_[7692]_ ;
  assign \new_[7696]_  = ~A203 & ~A202;
  assign \new_[7699]_  = A268 & A235;
  assign \new_[7700]_  = \new_[7699]_  & \new_[7696]_ ;
  assign \new_[7704]_  = ~A199 & A166;
  assign \new_[7705]_  = A168 & \new_[7704]_ ;
  assign \new_[7708]_  = ~A202 & ~A200;
  assign \new_[7711]_  = A268 & A235;
  assign \new_[7712]_  = \new_[7711]_  & \new_[7708]_ ;
  assign \new_[7716]_  = ~A201 & A167;
  assign \new_[7717]_  = A168 & \new_[7716]_ ;
  assign \new_[7720]_  = ~A203 & ~A202;
  assign \new_[7723]_  = A268 & A235;
  assign \new_[7724]_  = \new_[7723]_  & \new_[7720]_ ;
  assign \new_[7728]_  = ~A199 & A167;
  assign \new_[7729]_  = A168 & \new_[7728]_ ;
  assign \new_[7732]_  = ~A202 & ~A200;
  assign \new_[7735]_  = A268 & A235;
  assign \new_[7736]_  = \new_[7735]_  & \new_[7732]_ ;
  assign \new_[7740]_  = ~A202 & ~A201;
  assign \new_[7741]_  = A169 & \new_[7740]_ ;
  assign \new_[7744]_  = A235 & ~A203;
  assign \new_[7747]_  = A267 & A265;
  assign \new_[7748]_  = \new_[7747]_  & \new_[7744]_ ;
  assign \new_[7752]_  = ~A202 & ~A201;
  assign \new_[7753]_  = A169 & \new_[7752]_ ;
  assign \new_[7756]_  = A235 & ~A203;
  assign \new_[7759]_  = A267 & A266;
  assign \new_[7760]_  = \new_[7759]_  & \new_[7756]_ ;
  assign \new_[7764]_  = ~A202 & ~A201;
  assign \new_[7765]_  = A169 & \new_[7764]_ ;
  assign \new_[7768]_  = A232 & ~A203;
  assign \new_[7771]_  = A268 & A234;
  assign \new_[7772]_  = \new_[7771]_  & \new_[7768]_ ;
  assign \new_[7776]_  = ~A202 & ~A201;
  assign \new_[7777]_  = A169 & \new_[7776]_ ;
  assign \new_[7780]_  = A233 & ~A203;
  assign \new_[7783]_  = A268 & A234;
  assign \new_[7784]_  = \new_[7783]_  & \new_[7780]_ ;
  assign \new_[7788]_  = A200 & A199;
  assign \new_[7789]_  = A169 & \new_[7788]_ ;
  assign \new_[7792]_  = ~A202 & ~A201;
  assign \new_[7795]_  = A268 & A235;
  assign \new_[7796]_  = \new_[7795]_  & \new_[7792]_ ;
  assign \new_[7800]_  = ~A200 & ~A199;
  assign \new_[7801]_  = A169 & \new_[7800]_ ;
  assign \new_[7804]_  = A235 & ~A202;
  assign \new_[7807]_  = A267 & A265;
  assign \new_[7808]_  = \new_[7807]_  & \new_[7804]_ ;
  assign \new_[7812]_  = ~A200 & ~A199;
  assign \new_[7813]_  = A169 & \new_[7812]_ ;
  assign \new_[7816]_  = A235 & ~A202;
  assign \new_[7819]_  = A267 & A266;
  assign \new_[7820]_  = \new_[7819]_  & \new_[7816]_ ;
  assign \new_[7824]_  = ~A200 & ~A199;
  assign \new_[7825]_  = A169 & \new_[7824]_ ;
  assign \new_[7828]_  = A232 & ~A202;
  assign \new_[7831]_  = A268 & A234;
  assign \new_[7832]_  = \new_[7831]_  & \new_[7828]_ ;
  assign \new_[7836]_  = ~A200 & ~A199;
  assign \new_[7837]_  = A169 & \new_[7836]_ ;
  assign \new_[7840]_  = A233 & ~A202;
  assign \new_[7843]_  = A268 & A234;
  assign \new_[7844]_  = \new_[7843]_  & \new_[7840]_ ;
  assign \new_[7848]_  = ~A166 & ~A167;
  assign \new_[7849]_  = ~A169 & \new_[7848]_ ;
  assign \new_[7852]_  = A235 & A202;
  assign \new_[7855]_  = A267 & A265;
  assign \new_[7856]_  = \new_[7855]_  & \new_[7852]_ ;
  assign \new_[7860]_  = ~A166 & ~A167;
  assign \new_[7861]_  = ~A169 & \new_[7860]_ ;
  assign \new_[7864]_  = A235 & A202;
  assign \new_[7867]_  = A267 & A266;
  assign \new_[7868]_  = \new_[7867]_  & \new_[7864]_ ;
  assign \new_[7872]_  = ~A166 & ~A167;
  assign \new_[7873]_  = ~A169 & \new_[7872]_ ;
  assign \new_[7876]_  = A232 & A202;
  assign \new_[7879]_  = A268 & A234;
  assign \new_[7880]_  = \new_[7879]_  & \new_[7876]_ ;
  assign \new_[7884]_  = ~A166 & ~A167;
  assign \new_[7885]_  = ~A169 & \new_[7884]_ ;
  assign \new_[7888]_  = A233 & A202;
  assign \new_[7891]_  = A268 & A234;
  assign \new_[7892]_  = \new_[7891]_  & \new_[7888]_ ;
  assign \new_[7896]_  = ~A166 & ~A167;
  assign \new_[7897]_  = ~A169 & \new_[7896]_ ;
  assign \new_[7900]_  = A201 & A199;
  assign \new_[7903]_  = A268 & A235;
  assign \new_[7904]_  = \new_[7903]_  & \new_[7900]_ ;
  assign \new_[7908]_  = ~A166 & ~A167;
  assign \new_[7909]_  = ~A169 & \new_[7908]_ ;
  assign \new_[7912]_  = A201 & A200;
  assign \new_[7915]_  = A268 & A235;
  assign \new_[7916]_  = \new_[7915]_  & \new_[7912]_ ;
  assign \new_[7920]_  = A167 & ~A168;
  assign \new_[7921]_  = ~A169 & \new_[7920]_ ;
  assign \new_[7924]_  = A202 & A166;
  assign \new_[7927]_  = A268 & A235;
  assign \new_[7928]_  = \new_[7927]_  & \new_[7924]_ ;
  assign \new_[7932]_  = ~A168 & ~A169;
  assign \new_[7933]_  = ~A170 & \new_[7932]_ ;
  assign \new_[7936]_  = A235 & A202;
  assign \new_[7939]_  = A267 & A265;
  assign \new_[7940]_  = \new_[7939]_  & \new_[7936]_ ;
  assign \new_[7944]_  = ~A168 & ~A169;
  assign \new_[7945]_  = ~A170 & \new_[7944]_ ;
  assign \new_[7948]_  = A235 & A202;
  assign \new_[7951]_  = A267 & A266;
  assign \new_[7952]_  = \new_[7951]_  & \new_[7948]_ ;
  assign \new_[7956]_  = ~A168 & ~A169;
  assign \new_[7957]_  = ~A170 & \new_[7956]_ ;
  assign \new_[7960]_  = A232 & A202;
  assign \new_[7963]_  = A268 & A234;
  assign \new_[7964]_  = \new_[7963]_  & \new_[7960]_ ;
  assign \new_[7968]_  = ~A168 & ~A169;
  assign \new_[7969]_  = ~A170 & \new_[7968]_ ;
  assign \new_[7972]_  = A233 & A202;
  assign \new_[7975]_  = A268 & A234;
  assign \new_[7976]_  = \new_[7975]_  & \new_[7972]_ ;
  assign \new_[7980]_  = ~A168 & ~A169;
  assign \new_[7981]_  = ~A170 & \new_[7980]_ ;
  assign \new_[7984]_  = A201 & A199;
  assign \new_[7987]_  = A268 & A235;
  assign \new_[7988]_  = \new_[7987]_  & \new_[7984]_ ;
  assign \new_[7992]_  = ~A168 & ~A169;
  assign \new_[7993]_  = ~A170 & \new_[7992]_ ;
  assign \new_[7996]_  = A201 & A200;
  assign \new_[7999]_  = A268 & A235;
  assign \new_[8000]_  = \new_[7999]_  & \new_[7996]_ ;
  assign \new_[8003]_  = A166 & A168;
  assign \new_[8006]_  = ~A202 & ~A201;
  assign \new_[8007]_  = \new_[8006]_  & \new_[8003]_ ;
  assign \new_[8010]_  = A235 & ~A203;
  assign \new_[8013]_  = A267 & A265;
  assign \new_[8014]_  = \new_[8013]_  & \new_[8010]_ ;
  assign \new_[8017]_  = A166 & A168;
  assign \new_[8020]_  = ~A202 & ~A201;
  assign \new_[8021]_  = \new_[8020]_  & \new_[8017]_ ;
  assign \new_[8024]_  = A235 & ~A203;
  assign \new_[8027]_  = A267 & A266;
  assign \new_[8028]_  = \new_[8027]_  & \new_[8024]_ ;
  assign \new_[8031]_  = A166 & A168;
  assign \new_[8034]_  = ~A202 & ~A201;
  assign \new_[8035]_  = \new_[8034]_  & \new_[8031]_ ;
  assign \new_[8038]_  = A232 & ~A203;
  assign \new_[8041]_  = A268 & A234;
  assign \new_[8042]_  = \new_[8041]_  & \new_[8038]_ ;
  assign \new_[8045]_  = A166 & A168;
  assign \new_[8048]_  = ~A202 & ~A201;
  assign \new_[8049]_  = \new_[8048]_  & \new_[8045]_ ;
  assign \new_[8052]_  = A233 & ~A203;
  assign \new_[8055]_  = A268 & A234;
  assign \new_[8056]_  = \new_[8055]_  & \new_[8052]_ ;
  assign \new_[8059]_  = A166 & A168;
  assign \new_[8062]_  = A200 & A199;
  assign \new_[8063]_  = \new_[8062]_  & \new_[8059]_ ;
  assign \new_[8066]_  = ~A202 & ~A201;
  assign \new_[8069]_  = A268 & A235;
  assign \new_[8070]_  = \new_[8069]_  & \new_[8066]_ ;
  assign \new_[8073]_  = A166 & A168;
  assign \new_[8076]_  = ~A200 & ~A199;
  assign \new_[8077]_  = \new_[8076]_  & \new_[8073]_ ;
  assign \new_[8080]_  = A235 & ~A202;
  assign \new_[8083]_  = A267 & A265;
  assign \new_[8084]_  = \new_[8083]_  & \new_[8080]_ ;
  assign \new_[8087]_  = A166 & A168;
  assign \new_[8090]_  = ~A200 & ~A199;
  assign \new_[8091]_  = \new_[8090]_  & \new_[8087]_ ;
  assign \new_[8094]_  = A235 & ~A202;
  assign \new_[8097]_  = A267 & A266;
  assign \new_[8098]_  = \new_[8097]_  & \new_[8094]_ ;
  assign \new_[8101]_  = A166 & A168;
  assign \new_[8104]_  = ~A200 & ~A199;
  assign \new_[8105]_  = \new_[8104]_  & \new_[8101]_ ;
  assign \new_[8108]_  = A232 & ~A202;
  assign \new_[8111]_  = A268 & A234;
  assign \new_[8112]_  = \new_[8111]_  & \new_[8108]_ ;
  assign \new_[8115]_  = A166 & A168;
  assign \new_[8118]_  = ~A200 & ~A199;
  assign \new_[8119]_  = \new_[8118]_  & \new_[8115]_ ;
  assign \new_[8122]_  = A233 & ~A202;
  assign \new_[8125]_  = A268 & A234;
  assign \new_[8126]_  = \new_[8125]_  & \new_[8122]_ ;
  assign \new_[8129]_  = A167 & A168;
  assign \new_[8132]_  = ~A202 & ~A201;
  assign \new_[8133]_  = \new_[8132]_  & \new_[8129]_ ;
  assign \new_[8136]_  = A235 & ~A203;
  assign \new_[8139]_  = A267 & A265;
  assign \new_[8140]_  = \new_[8139]_  & \new_[8136]_ ;
  assign \new_[8143]_  = A167 & A168;
  assign \new_[8146]_  = ~A202 & ~A201;
  assign \new_[8147]_  = \new_[8146]_  & \new_[8143]_ ;
  assign \new_[8150]_  = A235 & ~A203;
  assign \new_[8153]_  = A267 & A266;
  assign \new_[8154]_  = \new_[8153]_  & \new_[8150]_ ;
  assign \new_[8157]_  = A167 & A168;
  assign \new_[8160]_  = ~A202 & ~A201;
  assign \new_[8161]_  = \new_[8160]_  & \new_[8157]_ ;
  assign \new_[8164]_  = A232 & ~A203;
  assign \new_[8167]_  = A268 & A234;
  assign \new_[8168]_  = \new_[8167]_  & \new_[8164]_ ;
  assign \new_[8171]_  = A167 & A168;
  assign \new_[8174]_  = ~A202 & ~A201;
  assign \new_[8175]_  = \new_[8174]_  & \new_[8171]_ ;
  assign \new_[8178]_  = A233 & ~A203;
  assign \new_[8181]_  = A268 & A234;
  assign \new_[8182]_  = \new_[8181]_  & \new_[8178]_ ;
  assign \new_[8185]_  = A167 & A168;
  assign \new_[8188]_  = A200 & A199;
  assign \new_[8189]_  = \new_[8188]_  & \new_[8185]_ ;
  assign \new_[8192]_  = ~A202 & ~A201;
  assign \new_[8195]_  = A268 & A235;
  assign \new_[8196]_  = \new_[8195]_  & \new_[8192]_ ;
  assign \new_[8199]_  = A167 & A168;
  assign \new_[8202]_  = ~A200 & ~A199;
  assign \new_[8203]_  = \new_[8202]_  & \new_[8199]_ ;
  assign \new_[8206]_  = A235 & ~A202;
  assign \new_[8209]_  = A267 & A265;
  assign \new_[8210]_  = \new_[8209]_  & \new_[8206]_ ;
  assign \new_[8213]_  = A167 & A168;
  assign \new_[8216]_  = ~A200 & ~A199;
  assign \new_[8217]_  = \new_[8216]_  & \new_[8213]_ ;
  assign \new_[8220]_  = A235 & ~A202;
  assign \new_[8223]_  = A267 & A266;
  assign \new_[8224]_  = \new_[8223]_  & \new_[8220]_ ;
  assign \new_[8227]_  = A167 & A168;
  assign \new_[8230]_  = ~A200 & ~A199;
  assign \new_[8231]_  = \new_[8230]_  & \new_[8227]_ ;
  assign \new_[8234]_  = A232 & ~A202;
  assign \new_[8237]_  = A268 & A234;
  assign \new_[8238]_  = \new_[8237]_  & \new_[8234]_ ;
  assign \new_[8241]_  = A167 & A168;
  assign \new_[8244]_  = ~A200 & ~A199;
  assign \new_[8245]_  = \new_[8244]_  & \new_[8241]_ ;
  assign \new_[8248]_  = A233 & ~A202;
  assign \new_[8251]_  = A268 & A234;
  assign \new_[8252]_  = \new_[8251]_  & \new_[8248]_ ;
  assign \new_[8255]_  = A167 & A170;
  assign \new_[8258]_  = ~A201 & ~A166;
  assign \new_[8259]_  = \new_[8258]_  & \new_[8255]_ ;
  assign \new_[8262]_  = ~A203 & ~A202;
  assign \new_[8265]_  = A268 & A235;
  assign \new_[8266]_  = \new_[8265]_  & \new_[8262]_ ;
  assign \new_[8269]_  = A167 & A170;
  assign \new_[8272]_  = ~A199 & ~A166;
  assign \new_[8273]_  = \new_[8272]_  & \new_[8269]_ ;
  assign \new_[8276]_  = ~A202 & ~A200;
  assign \new_[8279]_  = A268 & A235;
  assign \new_[8280]_  = \new_[8279]_  & \new_[8276]_ ;
  assign \new_[8283]_  = ~A167 & A170;
  assign \new_[8286]_  = ~A201 & A166;
  assign \new_[8287]_  = \new_[8286]_  & \new_[8283]_ ;
  assign \new_[8290]_  = ~A203 & ~A202;
  assign \new_[8293]_  = A268 & A235;
  assign \new_[8294]_  = \new_[8293]_  & \new_[8290]_ ;
  assign \new_[8297]_  = ~A167 & A170;
  assign \new_[8300]_  = ~A199 & A166;
  assign \new_[8301]_  = \new_[8300]_  & \new_[8297]_ ;
  assign \new_[8304]_  = ~A202 & ~A200;
  assign \new_[8307]_  = A268 & A235;
  assign \new_[8308]_  = \new_[8307]_  & \new_[8304]_ ;
  assign \new_[8311]_  = ~A201 & A169;
  assign \new_[8314]_  = ~A203 & ~A202;
  assign \new_[8315]_  = \new_[8314]_  & \new_[8311]_ ;
  assign \new_[8318]_  = ~A300 & A235;
  assign \new_[8321]_  = ~A302 & ~A301;
  assign \new_[8322]_  = \new_[8321]_  & \new_[8318]_ ;
  assign \new_[8325]_  = ~A201 & A169;
  assign \new_[8328]_  = ~A203 & ~A202;
  assign \new_[8329]_  = \new_[8328]_  & \new_[8325]_ ;
  assign \new_[8332]_  = ~A298 & A235;
  assign \new_[8335]_  = ~A301 & ~A299;
  assign \new_[8336]_  = \new_[8335]_  & \new_[8332]_ ;
  assign \new_[8339]_  = ~A201 & A169;
  assign \new_[8342]_  = ~A203 & ~A202;
  assign \new_[8343]_  = \new_[8342]_  & \new_[8339]_ ;
  assign \new_[8346]_  = ~A265 & A235;
  assign \new_[8349]_  = A269 & A266;
  assign \new_[8350]_  = \new_[8349]_  & \new_[8346]_ ;
  assign \new_[8353]_  = ~A201 & A169;
  assign \new_[8356]_  = ~A203 & ~A202;
  assign \new_[8357]_  = \new_[8356]_  & \new_[8353]_ ;
  assign \new_[8360]_  = A265 & A235;
  assign \new_[8363]_  = A269 & ~A266;
  assign \new_[8364]_  = \new_[8363]_  & \new_[8360]_ ;
  assign \new_[8367]_  = ~A201 & A169;
  assign \new_[8370]_  = ~A203 & ~A202;
  assign \new_[8371]_  = \new_[8370]_  & \new_[8367]_ ;
  assign \new_[8374]_  = A234 & A232;
  assign \new_[8377]_  = A267 & A265;
  assign \new_[8378]_  = \new_[8377]_  & \new_[8374]_ ;
  assign \new_[8381]_  = ~A201 & A169;
  assign \new_[8384]_  = ~A203 & ~A202;
  assign \new_[8385]_  = \new_[8384]_  & \new_[8381]_ ;
  assign \new_[8388]_  = A234 & A232;
  assign \new_[8391]_  = A267 & A266;
  assign \new_[8392]_  = \new_[8391]_  & \new_[8388]_ ;
  assign \new_[8395]_  = ~A201 & A169;
  assign \new_[8398]_  = ~A203 & ~A202;
  assign \new_[8399]_  = \new_[8398]_  & \new_[8395]_ ;
  assign \new_[8402]_  = A234 & A233;
  assign \new_[8405]_  = A267 & A265;
  assign \new_[8406]_  = \new_[8405]_  & \new_[8402]_ ;
  assign \new_[8409]_  = ~A201 & A169;
  assign \new_[8412]_  = ~A203 & ~A202;
  assign \new_[8413]_  = \new_[8412]_  & \new_[8409]_ ;
  assign \new_[8416]_  = A234 & A233;
  assign \new_[8419]_  = A267 & A266;
  assign \new_[8420]_  = \new_[8419]_  & \new_[8416]_ ;
  assign \new_[8423]_  = ~A201 & A169;
  assign \new_[8426]_  = ~A203 & ~A202;
  assign \new_[8427]_  = \new_[8426]_  & \new_[8423]_ ;
  assign \new_[8430]_  = A233 & ~A232;
  assign \new_[8433]_  = A268 & A236;
  assign \new_[8434]_  = \new_[8433]_  & \new_[8430]_ ;
  assign \new_[8437]_  = ~A201 & A169;
  assign \new_[8440]_  = ~A203 & ~A202;
  assign \new_[8441]_  = \new_[8440]_  & \new_[8437]_ ;
  assign \new_[8444]_  = ~A233 & A232;
  assign \new_[8447]_  = A268 & A236;
  assign \new_[8448]_  = \new_[8447]_  & \new_[8444]_ ;
  assign \new_[8451]_  = A199 & A169;
  assign \new_[8454]_  = ~A201 & A200;
  assign \new_[8455]_  = \new_[8454]_  & \new_[8451]_ ;
  assign \new_[8458]_  = A235 & ~A202;
  assign \new_[8461]_  = A267 & A265;
  assign \new_[8462]_  = \new_[8461]_  & \new_[8458]_ ;
  assign \new_[8465]_  = A199 & A169;
  assign \new_[8468]_  = ~A201 & A200;
  assign \new_[8469]_  = \new_[8468]_  & \new_[8465]_ ;
  assign \new_[8472]_  = A235 & ~A202;
  assign \new_[8475]_  = A267 & A266;
  assign \new_[8476]_  = \new_[8475]_  & \new_[8472]_ ;
  assign \new_[8479]_  = A199 & A169;
  assign \new_[8482]_  = ~A201 & A200;
  assign \new_[8483]_  = \new_[8482]_  & \new_[8479]_ ;
  assign \new_[8486]_  = A232 & ~A202;
  assign \new_[8489]_  = A268 & A234;
  assign \new_[8490]_  = \new_[8489]_  & \new_[8486]_ ;
  assign \new_[8493]_  = A199 & A169;
  assign \new_[8496]_  = ~A201 & A200;
  assign \new_[8497]_  = \new_[8496]_  & \new_[8493]_ ;
  assign \new_[8500]_  = A233 & ~A202;
  assign \new_[8503]_  = A268 & A234;
  assign \new_[8504]_  = \new_[8503]_  & \new_[8500]_ ;
  assign \new_[8507]_  = ~A199 & A169;
  assign \new_[8510]_  = ~A202 & ~A200;
  assign \new_[8511]_  = \new_[8510]_  & \new_[8507]_ ;
  assign \new_[8514]_  = ~A300 & A235;
  assign \new_[8517]_  = ~A302 & ~A301;
  assign \new_[8518]_  = \new_[8517]_  & \new_[8514]_ ;
  assign \new_[8521]_  = ~A199 & A169;
  assign \new_[8524]_  = ~A202 & ~A200;
  assign \new_[8525]_  = \new_[8524]_  & \new_[8521]_ ;
  assign \new_[8528]_  = ~A298 & A235;
  assign \new_[8531]_  = ~A301 & ~A299;
  assign \new_[8532]_  = \new_[8531]_  & \new_[8528]_ ;
  assign \new_[8535]_  = ~A199 & A169;
  assign \new_[8538]_  = ~A202 & ~A200;
  assign \new_[8539]_  = \new_[8538]_  & \new_[8535]_ ;
  assign \new_[8542]_  = ~A265 & A235;
  assign \new_[8545]_  = A269 & A266;
  assign \new_[8546]_  = \new_[8545]_  & \new_[8542]_ ;
  assign \new_[8549]_  = ~A199 & A169;
  assign \new_[8552]_  = ~A202 & ~A200;
  assign \new_[8553]_  = \new_[8552]_  & \new_[8549]_ ;
  assign \new_[8556]_  = A265 & A235;
  assign \new_[8559]_  = A269 & ~A266;
  assign \new_[8560]_  = \new_[8559]_  & \new_[8556]_ ;
  assign \new_[8563]_  = ~A199 & A169;
  assign \new_[8566]_  = ~A202 & ~A200;
  assign \new_[8567]_  = \new_[8566]_  & \new_[8563]_ ;
  assign \new_[8570]_  = A234 & A232;
  assign \new_[8573]_  = A267 & A265;
  assign \new_[8574]_  = \new_[8573]_  & \new_[8570]_ ;
  assign \new_[8577]_  = ~A199 & A169;
  assign \new_[8580]_  = ~A202 & ~A200;
  assign \new_[8581]_  = \new_[8580]_  & \new_[8577]_ ;
  assign \new_[8584]_  = A234 & A232;
  assign \new_[8587]_  = A267 & A266;
  assign \new_[8588]_  = \new_[8587]_  & \new_[8584]_ ;
  assign \new_[8591]_  = ~A199 & A169;
  assign \new_[8594]_  = ~A202 & ~A200;
  assign \new_[8595]_  = \new_[8594]_  & \new_[8591]_ ;
  assign \new_[8598]_  = A234 & A233;
  assign \new_[8601]_  = A267 & A265;
  assign \new_[8602]_  = \new_[8601]_  & \new_[8598]_ ;
  assign \new_[8605]_  = ~A199 & A169;
  assign \new_[8608]_  = ~A202 & ~A200;
  assign \new_[8609]_  = \new_[8608]_  & \new_[8605]_ ;
  assign \new_[8612]_  = A234 & A233;
  assign \new_[8615]_  = A267 & A266;
  assign \new_[8616]_  = \new_[8615]_  & \new_[8612]_ ;
  assign \new_[8619]_  = ~A199 & A169;
  assign \new_[8622]_  = ~A202 & ~A200;
  assign \new_[8623]_  = \new_[8622]_  & \new_[8619]_ ;
  assign \new_[8626]_  = A233 & ~A232;
  assign \new_[8629]_  = A268 & A236;
  assign \new_[8630]_  = \new_[8629]_  & \new_[8626]_ ;
  assign \new_[8633]_  = ~A199 & A169;
  assign \new_[8636]_  = ~A202 & ~A200;
  assign \new_[8637]_  = \new_[8636]_  & \new_[8633]_ ;
  assign \new_[8640]_  = ~A233 & A232;
  assign \new_[8643]_  = A268 & A236;
  assign \new_[8644]_  = \new_[8643]_  & \new_[8640]_ ;
  assign \new_[8647]_  = ~A167 & ~A169;
  assign \new_[8650]_  = A202 & ~A166;
  assign \new_[8651]_  = \new_[8650]_  & \new_[8647]_ ;
  assign \new_[8654]_  = ~A300 & A235;
  assign \new_[8657]_  = ~A302 & ~A301;
  assign \new_[8658]_  = \new_[8657]_  & \new_[8654]_ ;
  assign \new_[8661]_  = ~A167 & ~A169;
  assign \new_[8664]_  = A202 & ~A166;
  assign \new_[8665]_  = \new_[8664]_  & \new_[8661]_ ;
  assign \new_[8668]_  = ~A298 & A235;
  assign \new_[8671]_  = ~A301 & ~A299;
  assign \new_[8672]_  = \new_[8671]_  & \new_[8668]_ ;
  assign \new_[8675]_  = ~A167 & ~A169;
  assign \new_[8678]_  = A202 & ~A166;
  assign \new_[8679]_  = \new_[8678]_  & \new_[8675]_ ;
  assign \new_[8682]_  = ~A265 & A235;
  assign \new_[8685]_  = A269 & A266;
  assign \new_[8686]_  = \new_[8685]_  & \new_[8682]_ ;
  assign \new_[8689]_  = ~A167 & ~A169;
  assign \new_[8692]_  = A202 & ~A166;
  assign \new_[8693]_  = \new_[8692]_  & \new_[8689]_ ;
  assign \new_[8696]_  = A265 & A235;
  assign \new_[8699]_  = A269 & ~A266;
  assign \new_[8700]_  = \new_[8699]_  & \new_[8696]_ ;
  assign \new_[8703]_  = ~A167 & ~A169;
  assign \new_[8706]_  = A202 & ~A166;
  assign \new_[8707]_  = \new_[8706]_  & \new_[8703]_ ;
  assign \new_[8710]_  = A234 & A232;
  assign \new_[8713]_  = A267 & A265;
  assign \new_[8714]_  = \new_[8713]_  & \new_[8710]_ ;
  assign \new_[8717]_  = ~A167 & ~A169;
  assign \new_[8720]_  = A202 & ~A166;
  assign \new_[8721]_  = \new_[8720]_  & \new_[8717]_ ;
  assign \new_[8724]_  = A234 & A232;
  assign \new_[8727]_  = A267 & A266;
  assign \new_[8728]_  = \new_[8727]_  & \new_[8724]_ ;
  assign \new_[8731]_  = ~A167 & ~A169;
  assign \new_[8734]_  = A202 & ~A166;
  assign \new_[8735]_  = \new_[8734]_  & \new_[8731]_ ;
  assign \new_[8738]_  = A234 & A233;
  assign \new_[8741]_  = A267 & A265;
  assign \new_[8742]_  = \new_[8741]_  & \new_[8738]_ ;
  assign \new_[8745]_  = ~A167 & ~A169;
  assign \new_[8748]_  = A202 & ~A166;
  assign \new_[8749]_  = \new_[8748]_  & \new_[8745]_ ;
  assign \new_[8752]_  = A234 & A233;
  assign \new_[8755]_  = A267 & A266;
  assign \new_[8756]_  = \new_[8755]_  & \new_[8752]_ ;
  assign \new_[8759]_  = ~A167 & ~A169;
  assign \new_[8762]_  = A202 & ~A166;
  assign \new_[8763]_  = \new_[8762]_  & \new_[8759]_ ;
  assign \new_[8766]_  = A233 & ~A232;
  assign \new_[8769]_  = A268 & A236;
  assign \new_[8770]_  = \new_[8769]_  & \new_[8766]_ ;
  assign \new_[8773]_  = ~A167 & ~A169;
  assign \new_[8776]_  = A202 & ~A166;
  assign \new_[8777]_  = \new_[8776]_  & \new_[8773]_ ;
  assign \new_[8780]_  = ~A233 & A232;
  assign \new_[8783]_  = A268 & A236;
  assign \new_[8784]_  = \new_[8783]_  & \new_[8780]_ ;
  assign \new_[8787]_  = ~A167 & ~A169;
  assign \new_[8790]_  = A199 & ~A166;
  assign \new_[8791]_  = \new_[8790]_  & \new_[8787]_ ;
  assign \new_[8794]_  = A235 & A201;
  assign \new_[8797]_  = A267 & A265;
  assign \new_[8798]_  = \new_[8797]_  & \new_[8794]_ ;
  assign \new_[8801]_  = ~A167 & ~A169;
  assign \new_[8804]_  = A199 & ~A166;
  assign \new_[8805]_  = \new_[8804]_  & \new_[8801]_ ;
  assign \new_[8808]_  = A235 & A201;
  assign \new_[8811]_  = A267 & A266;
  assign \new_[8812]_  = \new_[8811]_  & \new_[8808]_ ;
  assign \new_[8815]_  = ~A167 & ~A169;
  assign \new_[8818]_  = A199 & ~A166;
  assign \new_[8819]_  = \new_[8818]_  & \new_[8815]_ ;
  assign \new_[8822]_  = A232 & A201;
  assign \new_[8825]_  = A268 & A234;
  assign \new_[8826]_  = \new_[8825]_  & \new_[8822]_ ;
  assign \new_[8829]_  = ~A167 & ~A169;
  assign \new_[8832]_  = A199 & ~A166;
  assign \new_[8833]_  = \new_[8832]_  & \new_[8829]_ ;
  assign \new_[8836]_  = A233 & A201;
  assign \new_[8839]_  = A268 & A234;
  assign \new_[8840]_  = \new_[8839]_  & \new_[8836]_ ;
  assign \new_[8843]_  = ~A167 & ~A169;
  assign \new_[8846]_  = A200 & ~A166;
  assign \new_[8847]_  = \new_[8846]_  & \new_[8843]_ ;
  assign \new_[8850]_  = A235 & A201;
  assign \new_[8853]_  = A267 & A265;
  assign \new_[8854]_  = \new_[8853]_  & \new_[8850]_ ;
  assign \new_[8857]_  = ~A167 & ~A169;
  assign \new_[8860]_  = A200 & ~A166;
  assign \new_[8861]_  = \new_[8860]_  & \new_[8857]_ ;
  assign \new_[8864]_  = A235 & A201;
  assign \new_[8867]_  = A267 & A266;
  assign \new_[8868]_  = \new_[8867]_  & \new_[8864]_ ;
  assign \new_[8871]_  = ~A167 & ~A169;
  assign \new_[8874]_  = A200 & ~A166;
  assign \new_[8875]_  = \new_[8874]_  & \new_[8871]_ ;
  assign \new_[8878]_  = A232 & A201;
  assign \new_[8881]_  = A268 & A234;
  assign \new_[8882]_  = \new_[8881]_  & \new_[8878]_ ;
  assign \new_[8885]_  = ~A167 & ~A169;
  assign \new_[8888]_  = A200 & ~A166;
  assign \new_[8889]_  = \new_[8888]_  & \new_[8885]_ ;
  assign \new_[8892]_  = A233 & A201;
  assign \new_[8895]_  = A268 & A234;
  assign \new_[8896]_  = \new_[8895]_  & \new_[8892]_ ;
  assign \new_[8899]_  = ~A167 & ~A169;
  assign \new_[8902]_  = ~A199 & ~A166;
  assign \new_[8903]_  = \new_[8902]_  & \new_[8899]_ ;
  assign \new_[8906]_  = A203 & A200;
  assign \new_[8909]_  = A268 & A235;
  assign \new_[8910]_  = \new_[8909]_  & \new_[8906]_ ;
  assign \new_[8913]_  = ~A167 & ~A169;
  assign \new_[8916]_  = A199 & ~A166;
  assign \new_[8917]_  = \new_[8916]_  & \new_[8913]_ ;
  assign \new_[8920]_  = A203 & ~A200;
  assign \new_[8923]_  = A268 & A235;
  assign \new_[8924]_  = \new_[8923]_  & \new_[8920]_ ;
  assign \new_[8927]_  = ~A168 & ~A169;
  assign \new_[8930]_  = A166 & A167;
  assign \new_[8931]_  = \new_[8930]_  & \new_[8927]_ ;
  assign \new_[8934]_  = A235 & A202;
  assign \new_[8937]_  = A267 & A265;
  assign \new_[8938]_  = \new_[8937]_  & \new_[8934]_ ;
  assign \new_[8941]_  = ~A168 & ~A169;
  assign \new_[8944]_  = A166 & A167;
  assign \new_[8945]_  = \new_[8944]_  & \new_[8941]_ ;
  assign \new_[8948]_  = A235 & A202;
  assign \new_[8951]_  = A267 & A266;
  assign \new_[8952]_  = \new_[8951]_  & \new_[8948]_ ;
  assign \new_[8955]_  = ~A168 & ~A169;
  assign \new_[8958]_  = A166 & A167;
  assign \new_[8959]_  = \new_[8958]_  & \new_[8955]_ ;
  assign \new_[8962]_  = A232 & A202;
  assign \new_[8965]_  = A268 & A234;
  assign \new_[8966]_  = \new_[8965]_  & \new_[8962]_ ;
  assign \new_[8969]_  = ~A168 & ~A169;
  assign \new_[8972]_  = A166 & A167;
  assign \new_[8973]_  = \new_[8972]_  & \new_[8969]_ ;
  assign \new_[8976]_  = A233 & A202;
  assign \new_[8979]_  = A268 & A234;
  assign \new_[8980]_  = \new_[8979]_  & \new_[8976]_ ;
  assign \new_[8983]_  = ~A168 & ~A169;
  assign \new_[8986]_  = A166 & A167;
  assign \new_[8987]_  = \new_[8986]_  & \new_[8983]_ ;
  assign \new_[8990]_  = A201 & A199;
  assign \new_[8993]_  = A268 & A235;
  assign \new_[8994]_  = \new_[8993]_  & \new_[8990]_ ;
  assign \new_[8997]_  = ~A168 & ~A169;
  assign \new_[9000]_  = A166 & A167;
  assign \new_[9001]_  = \new_[9000]_  & \new_[8997]_ ;
  assign \new_[9004]_  = A201 & A200;
  assign \new_[9007]_  = A268 & A235;
  assign \new_[9008]_  = \new_[9007]_  & \new_[9004]_ ;
  assign \new_[9011]_  = ~A169 & ~A170;
  assign \new_[9014]_  = A202 & ~A168;
  assign \new_[9015]_  = \new_[9014]_  & \new_[9011]_ ;
  assign \new_[9018]_  = ~A300 & A235;
  assign \new_[9021]_  = ~A302 & ~A301;
  assign \new_[9022]_  = \new_[9021]_  & \new_[9018]_ ;
  assign \new_[9025]_  = ~A169 & ~A170;
  assign \new_[9028]_  = A202 & ~A168;
  assign \new_[9029]_  = \new_[9028]_  & \new_[9025]_ ;
  assign \new_[9032]_  = ~A298 & A235;
  assign \new_[9035]_  = ~A301 & ~A299;
  assign \new_[9036]_  = \new_[9035]_  & \new_[9032]_ ;
  assign \new_[9039]_  = ~A169 & ~A170;
  assign \new_[9042]_  = A202 & ~A168;
  assign \new_[9043]_  = \new_[9042]_  & \new_[9039]_ ;
  assign \new_[9046]_  = ~A265 & A235;
  assign \new_[9049]_  = A269 & A266;
  assign \new_[9050]_  = \new_[9049]_  & \new_[9046]_ ;
  assign \new_[9053]_  = ~A169 & ~A170;
  assign \new_[9056]_  = A202 & ~A168;
  assign \new_[9057]_  = \new_[9056]_  & \new_[9053]_ ;
  assign \new_[9060]_  = A265 & A235;
  assign \new_[9063]_  = A269 & ~A266;
  assign \new_[9064]_  = \new_[9063]_  & \new_[9060]_ ;
  assign \new_[9067]_  = ~A169 & ~A170;
  assign \new_[9070]_  = A202 & ~A168;
  assign \new_[9071]_  = \new_[9070]_  & \new_[9067]_ ;
  assign \new_[9074]_  = A234 & A232;
  assign \new_[9077]_  = A267 & A265;
  assign \new_[9078]_  = \new_[9077]_  & \new_[9074]_ ;
  assign \new_[9081]_  = ~A169 & ~A170;
  assign \new_[9084]_  = A202 & ~A168;
  assign \new_[9085]_  = \new_[9084]_  & \new_[9081]_ ;
  assign \new_[9088]_  = A234 & A232;
  assign \new_[9091]_  = A267 & A266;
  assign \new_[9092]_  = \new_[9091]_  & \new_[9088]_ ;
  assign \new_[9095]_  = ~A169 & ~A170;
  assign \new_[9098]_  = A202 & ~A168;
  assign \new_[9099]_  = \new_[9098]_  & \new_[9095]_ ;
  assign \new_[9102]_  = A234 & A233;
  assign \new_[9105]_  = A267 & A265;
  assign \new_[9106]_  = \new_[9105]_  & \new_[9102]_ ;
  assign \new_[9109]_  = ~A169 & ~A170;
  assign \new_[9112]_  = A202 & ~A168;
  assign \new_[9113]_  = \new_[9112]_  & \new_[9109]_ ;
  assign \new_[9116]_  = A234 & A233;
  assign \new_[9119]_  = A267 & A266;
  assign \new_[9120]_  = \new_[9119]_  & \new_[9116]_ ;
  assign \new_[9123]_  = ~A169 & ~A170;
  assign \new_[9126]_  = A202 & ~A168;
  assign \new_[9127]_  = \new_[9126]_  & \new_[9123]_ ;
  assign \new_[9130]_  = A233 & ~A232;
  assign \new_[9133]_  = A268 & A236;
  assign \new_[9134]_  = \new_[9133]_  & \new_[9130]_ ;
  assign \new_[9137]_  = ~A169 & ~A170;
  assign \new_[9140]_  = A202 & ~A168;
  assign \new_[9141]_  = \new_[9140]_  & \new_[9137]_ ;
  assign \new_[9144]_  = ~A233 & A232;
  assign \new_[9147]_  = A268 & A236;
  assign \new_[9148]_  = \new_[9147]_  & \new_[9144]_ ;
  assign \new_[9151]_  = ~A169 & ~A170;
  assign \new_[9154]_  = A199 & ~A168;
  assign \new_[9155]_  = \new_[9154]_  & \new_[9151]_ ;
  assign \new_[9158]_  = A235 & A201;
  assign \new_[9161]_  = A267 & A265;
  assign \new_[9162]_  = \new_[9161]_  & \new_[9158]_ ;
  assign \new_[9165]_  = ~A169 & ~A170;
  assign \new_[9168]_  = A199 & ~A168;
  assign \new_[9169]_  = \new_[9168]_  & \new_[9165]_ ;
  assign \new_[9172]_  = A235 & A201;
  assign \new_[9175]_  = A267 & A266;
  assign \new_[9176]_  = \new_[9175]_  & \new_[9172]_ ;
  assign \new_[9179]_  = ~A169 & ~A170;
  assign \new_[9182]_  = A199 & ~A168;
  assign \new_[9183]_  = \new_[9182]_  & \new_[9179]_ ;
  assign \new_[9186]_  = A232 & A201;
  assign \new_[9189]_  = A268 & A234;
  assign \new_[9190]_  = \new_[9189]_  & \new_[9186]_ ;
  assign \new_[9193]_  = ~A169 & ~A170;
  assign \new_[9196]_  = A199 & ~A168;
  assign \new_[9197]_  = \new_[9196]_  & \new_[9193]_ ;
  assign \new_[9200]_  = A233 & A201;
  assign \new_[9203]_  = A268 & A234;
  assign \new_[9204]_  = \new_[9203]_  & \new_[9200]_ ;
  assign \new_[9207]_  = ~A169 & ~A170;
  assign \new_[9210]_  = A200 & ~A168;
  assign \new_[9211]_  = \new_[9210]_  & \new_[9207]_ ;
  assign \new_[9214]_  = A235 & A201;
  assign \new_[9217]_  = A267 & A265;
  assign \new_[9218]_  = \new_[9217]_  & \new_[9214]_ ;
  assign \new_[9221]_  = ~A169 & ~A170;
  assign \new_[9224]_  = A200 & ~A168;
  assign \new_[9225]_  = \new_[9224]_  & \new_[9221]_ ;
  assign \new_[9228]_  = A235 & A201;
  assign \new_[9231]_  = A267 & A266;
  assign \new_[9232]_  = \new_[9231]_  & \new_[9228]_ ;
  assign \new_[9235]_  = ~A169 & ~A170;
  assign \new_[9238]_  = A200 & ~A168;
  assign \new_[9239]_  = \new_[9238]_  & \new_[9235]_ ;
  assign \new_[9242]_  = A232 & A201;
  assign \new_[9245]_  = A268 & A234;
  assign \new_[9246]_  = \new_[9245]_  & \new_[9242]_ ;
  assign \new_[9249]_  = ~A169 & ~A170;
  assign \new_[9252]_  = A200 & ~A168;
  assign \new_[9253]_  = \new_[9252]_  & \new_[9249]_ ;
  assign \new_[9256]_  = A233 & A201;
  assign \new_[9259]_  = A268 & A234;
  assign \new_[9260]_  = \new_[9259]_  & \new_[9256]_ ;
  assign \new_[9263]_  = ~A169 & ~A170;
  assign \new_[9266]_  = ~A199 & ~A168;
  assign \new_[9267]_  = \new_[9266]_  & \new_[9263]_ ;
  assign \new_[9270]_  = A203 & A200;
  assign \new_[9273]_  = A268 & A235;
  assign \new_[9274]_  = \new_[9273]_  & \new_[9270]_ ;
  assign \new_[9277]_  = ~A169 & ~A170;
  assign \new_[9280]_  = A199 & ~A168;
  assign \new_[9281]_  = \new_[9280]_  & \new_[9277]_ ;
  assign \new_[9284]_  = A203 & ~A200;
  assign \new_[9287]_  = A268 & A235;
  assign \new_[9288]_  = \new_[9287]_  & \new_[9284]_ ;
  assign \new_[9291]_  = A166 & A168;
  assign \new_[9294]_  = ~A202 & ~A201;
  assign \new_[9295]_  = \new_[9294]_  & \new_[9291]_ ;
  assign \new_[9298]_  = A235 & ~A203;
  assign \new_[9302]_  = ~A302 & ~A301;
  assign \new_[9303]_  = ~A300 & \new_[9302]_ ;
  assign \new_[9304]_  = \new_[9303]_  & \new_[9298]_ ;
  assign \new_[9307]_  = A166 & A168;
  assign \new_[9310]_  = ~A202 & ~A201;
  assign \new_[9311]_  = \new_[9310]_  & \new_[9307]_ ;
  assign \new_[9314]_  = A235 & ~A203;
  assign \new_[9318]_  = ~A301 & ~A299;
  assign \new_[9319]_  = ~A298 & \new_[9318]_ ;
  assign \new_[9320]_  = \new_[9319]_  & \new_[9314]_ ;
  assign \new_[9323]_  = A166 & A168;
  assign \new_[9326]_  = ~A202 & ~A201;
  assign \new_[9327]_  = \new_[9326]_  & \new_[9323]_ ;
  assign \new_[9330]_  = A235 & ~A203;
  assign \new_[9334]_  = A269 & A266;
  assign \new_[9335]_  = ~A265 & \new_[9334]_ ;
  assign \new_[9336]_  = \new_[9335]_  & \new_[9330]_ ;
  assign \new_[9339]_  = A166 & A168;
  assign \new_[9342]_  = ~A202 & ~A201;
  assign \new_[9343]_  = \new_[9342]_  & \new_[9339]_ ;
  assign \new_[9346]_  = A235 & ~A203;
  assign \new_[9350]_  = A269 & ~A266;
  assign \new_[9351]_  = A265 & \new_[9350]_ ;
  assign \new_[9352]_  = \new_[9351]_  & \new_[9346]_ ;
  assign \new_[9355]_  = A166 & A168;
  assign \new_[9358]_  = ~A202 & ~A201;
  assign \new_[9359]_  = \new_[9358]_  & \new_[9355]_ ;
  assign \new_[9362]_  = A232 & ~A203;
  assign \new_[9366]_  = A267 & A265;
  assign \new_[9367]_  = A234 & \new_[9366]_ ;
  assign \new_[9368]_  = \new_[9367]_  & \new_[9362]_ ;
  assign \new_[9371]_  = A166 & A168;
  assign \new_[9374]_  = ~A202 & ~A201;
  assign \new_[9375]_  = \new_[9374]_  & \new_[9371]_ ;
  assign \new_[9378]_  = A232 & ~A203;
  assign \new_[9382]_  = A267 & A266;
  assign \new_[9383]_  = A234 & \new_[9382]_ ;
  assign \new_[9384]_  = \new_[9383]_  & \new_[9378]_ ;
  assign \new_[9387]_  = A166 & A168;
  assign \new_[9390]_  = ~A202 & ~A201;
  assign \new_[9391]_  = \new_[9390]_  & \new_[9387]_ ;
  assign \new_[9394]_  = A233 & ~A203;
  assign \new_[9398]_  = A267 & A265;
  assign \new_[9399]_  = A234 & \new_[9398]_ ;
  assign \new_[9400]_  = \new_[9399]_  & \new_[9394]_ ;
  assign \new_[9403]_  = A166 & A168;
  assign \new_[9406]_  = ~A202 & ~A201;
  assign \new_[9407]_  = \new_[9406]_  & \new_[9403]_ ;
  assign \new_[9410]_  = A233 & ~A203;
  assign \new_[9414]_  = A267 & A266;
  assign \new_[9415]_  = A234 & \new_[9414]_ ;
  assign \new_[9416]_  = \new_[9415]_  & \new_[9410]_ ;
  assign \new_[9419]_  = A166 & A168;
  assign \new_[9422]_  = ~A202 & ~A201;
  assign \new_[9423]_  = \new_[9422]_  & \new_[9419]_ ;
  assign \new_[9426]_  = ~A232 & ~A203;
  assign \new_[9430]_  = A268 & A236;
  assign \new_[9431]_  = A233 & \new_[9430]_ ;
  assign \new_[9432]_  = \new_[9431]_  & \new_[9426]_ ;
  assign \new_[9435]_  = A166 & A168;
  assign \new_[9438]_  = ~A202 & ~A201;
  assign \new_[9439]_  = \new_[9438]_  & \new_[9435]_ ;
  assign \new_[9442]_  = A232 & ~A203;
  assign \new_[9446]_  = A268 & A236;
  assign \new_[9447]_  = ~A233 & \new_[9446]_ ;
  assign \new_[9448]_  = \new_[9447]_  & \new_[9442]_ ;
  assign \new_[9451]_  = A166 & A168;
  assign \new_[9454]_  = A200 & A199;
  assign \new_[9455]_  = \new_[9454]_  & \new_[9451]_ ;
  assign \new_[9458]_  = ~A202 & ~A201;
  assign \new_[9462]_  = A267 & A265;
  assign \new_[9463]_  = A235 & \new_[9462]_ ;
  assign \new_[9464]_  = \new_[9463]_  & \new_[9458]_ ;
  assign \new_[9467]_  = A166 & A168;
  assign \new_[9470]_  = A200 & A199;
  assign \new_[9471]_  = \new_[9470]_  & \new_[9467]_ ;
  assign \new_[9474]_  = ~A202 & ~A201;
  assign \new_[9478]_  = A267 & A266;
  assign \new_[9479]_  = A235 & \new_[9478]_ ;
  assign \new_[9480]_  = \new_[9479]_  & \new_[9474]_ ;
  assign \new_[9483]_  = A166 & A168;
  assign \new_[9486]_  = A200 & A199;
  assign \new_[9487]_  = \new_[9486]_  & \new_[9483]_ ;
  assign \new_[9490]_  = ~A202 & ~A201;
  assign \new_[9494]_  = A268 & A234;
  assign \new_[9495]_  = A232 & \new_[9494]_ ;
  assign \new_[9496]_  = \new_[9495]_  & \new_[9490]_ ;
  assign \new_[9499]_  = A166 & A168;
  assign \new_[9502]_  = A200 & A199;
  assign \new_[9503]_  = \new_[9502]_  & \new_[9499]_ ;
  assign \new_[9506]_  = ~A202 & ~A201;
  assign \new_[9510]_  = A268 & A234;
  assign \new_[9511]_  = A233 & \new_[9510]_ ;
  assign \new_[9512]_  = \new_[9511]_  & \new_[9506]_ ;
  assign \new_[9515]_  = A166 & A168;
  assign \new_[9518]_  = ~A200 & ~A199;
  assign \new_[9519]_  = \new_[9518]_  & \new_[9515]_ ;
  assign \new_[9522]_  = A235 & ~A202;
  assign \new_[9526]_  = ~A302 & ~A301;
  assign \new_[9527]_  = ~A300 & \new_[9526]_ ;
  assign \new_[9528]_  = \new_[9527]_  & \new_[9522]_ ;
  assign \new_[9531]_  = A166 & A168;
  assign \new_[9534]_  = ~A200 & ~A199;
  assign \new_[9535]_  = \new_[9534]_  & \new_[9531]_ ;
  assign \new_[9538]_  = A235 & ~A202;
  assign \new_[9542]_  = ~A301 & ~A299;
  assign \new_[9543]_  = ~A298 & \new_[9542]_ ;
  assign \new_[9544]_  = \new_[9543]_  & \new_[9538]_ ;
  assign \new_[9547]_  = A166 & A168;
  assign \new_[9550]_  = ~A200 & ~A199;
  assign \new_[9551]_  = \new_[9550]_  & \new_[9547]_ ;
  assign \new_[9554]_  = A235 & ~A202;
  assign \new_[9558]_  = A269 & A266;
  assign \new_[9559]_  = ~A265 & \new_[9558]_ ;
  assign \new_[9560]_  = \new_[9559]_  & \new_[9554]_ ;
  assign \new_[9563]_  = A166 & A168;
  assign \new_[9566]_  = ~A200 & ~A199;
  assign \new_[9567]_  = \new_[9566]_  & \new_[9563]_ ;
  assign \new_[9570]_  = A235 & ~A202;
  assign \new_[9574]_  = A269 & ~A266;
  assign \new_[9575]_  = A265 & \new_[9574]_ ;
  assign \new_[9576]_  = \new_[9575]_  & \new_[9570]_ ;
  assign \new_[9579]_  = A166 & A168;
  assign \new_[9582]_  = ~A200 & ~A199;
  assign \new_[9583]_  = \new_[9582]_  & \new_[9579]_ ;
  assign \new_[9586]_  = A232 & ~A202;
  assign \new_[9590]_  = A267 & A265;
  assign \new_[9591]_  = A234 & \new_[9590]_ ;
  assign \new_[9592]_  = \new_[9591]_  & \new_[9586]_ ;
  assign \new_[9595]_  = A166 & A168;
  assign \new_[9598]_  = ~A200 & ~A199;
  assign \new_[9599]_  = \new_[9598]_  & \new_[9595]_ ;
  assign \new_[9602]_  = A232 & ~A202;
  assign \new_[9606]_  = A267 & A266;
  assign \new_[9607]_  = A234 & \new_[9606]_ ;
  assign \new_[9608]_  = \new_[9607]_  & \new_[9602]_ ;
  assign \new_[9611]_  = A166 & A168;
  assign \new_[9614]_  = ~A200 & ~A199;
  assign \new_[9615]_  = \new_[9614]_  & \new_[9611]_ ;
  assign \new_[9618]_  = A233 & ~A202;
  assign \new_[9622]_  = A267 & A265;
  assign \new_[9623]_  = A234 & \new_[9622]_ ;
  assign \new_[9624]_  = \new_[9623]_  & \new_[9618]_ ;
  assign \new_[9627]_  = A166 & A168;
  assign \new_[9630]_  = ~A200 & ~A199;
  assign \new_[9631]_  = \new_[9630]_  & \new_[9627]_ ;
  assign \new_[9634]_  = A233 & ~A202;
  assign \new_[9638]_  = A267 & A266;
  assign \new_[9639]_  = A234 & \new_[9638]_ ;
  assign \new_[9640]_  = \new_[9639]_  & \new_[9634]_ ;
  assign \new_[9643]_  = A166 & A168;
  assign \new_[9646]_  = ~A200 & ~A199;
  assign \new_[9647]_  = \new_[9646]_  & \new_[9643]_ ;
  assign \new_[9650]_  = ~A232 & ~A202;
  assign \new_[9654]_  = A268 & A236;
  assign \new_[9655]_  = A233 & \new_[9654]_ ;
  assign \new_[9656]_  = \new_[9655]_  & \new_[9650]_ ;
  assign \new_[9659]_  = A166 & A168;
  assign \new_[9662]_  = ~A200 & ~A199;
  assign \new_[9663]_  = \new_[9662]_  & \new_[9659]_ ;
  assign \new_[9666]_  = A232 & ~A202;
  assign \new_[9670]_  = A268 & A236;
  assign \new_[9671]_  = ~A233 & \new_[9670]_ ;
  assign \new_[9672]_  = \new_[9671]_  & \new_[9666]_ ;
  assign \new_[9675]_  = A167 & A168;
  assign \new_[9678]_  = ~A202 & ~A201;
  assign \new_[9679]_  = \new_[9678]_  & \new_[9675]_ ;
  assign \new_[9682]_  = A235 & ~A203;
  assign \new_[9686]_  = ~A302 & ~A301;
  assign \new_[9687]_  = ~A300 & \new_[9686]_ ;
  assign \new_[9688]_  = \new_[9687]_  & \new_[9682]_ ;
  assign \new_[9691]_  = A167 & A168;
  assign \new_[9694]_  = ~A202 & ~A201;
  assign \new_[9695]_  = \new_[9694]_  & \new_[9691]_ ;
  assign \new_[9698]_  = A235 & ~A203;
  assign \new_[9702]_  = ~A301 & ~A299;
  assign \new_[9703]_  = ~A298 & \new_[9702]_ ;
  assign \new_[9704]_  = \new_[9703]_  & \new_[9698]_ ;
  assign \new_[9707]_  = A167 & A168;
  assign \new_[9710]_  = ~A202 & ~A201;
  assign \new_[9711]_  = \new_[9710]_  & \new_[9707]_ ;
  assign \new_[9714]_  = A235 & ~A203;
  assign \new_[9718]_  = A269 & A266;
  assign \new_[9719]_  = ~A265 & \new_[9718]_ ;
  assign \new_[9720]_  = \new_[9719]_  & \new_[9714]_ ;
  assign \new_[9723]_  = A167 & A168;
  assign \new_[9726]_  = ~A202 & ~A201;
  assign \new_[9727]_  = \new_[9726]_  & \new_[9723]_ ;
  assign \new_[9730]_  = A235 & ~A203;
  assign \new_[9734]_  = A269 & ~A266;
  assign \new_[9735]_  = A265 & \new_[9734]_ ;
  assign \new_[9736]_  = \new_[9735]_  & \new_[9730]_ ;
  assign \new_[9739]_  = A167 & A168;
  assign \new_[9742]_  = ~A202 & ~A201;
  assign \new_[9743]_  = \new_[9742]_  & \new_[9739]_ ;
  assign \new_[9746]_  = A232 & ~A203;
  assign \new_[9750]_  = A267 & A265;
  assign \new_[9751]_  = A234 & \new_[9750]_ ;
  assign \new_[9752]_  = \new_[9751]_  & \new_[9746]_ ;
  assign \new_[9755]_  = A167 & A168;
  assign \new_[9758]_  = ~A202 & ~A201;
  assign \new_[9759]_  = \new_[9758]_  & \new_[9755]_ ;
  assign \new_[9762]_  = A232 & ~A203;
  assign \new_[9766]_  = A267 & A266;
  assign \new_[9767]_  = A234 & \new_[9766]_ ;
  assign \new_[9768]_  = \new_[9767]_  & \new_[9762]_ ;
  assign \new_[9771]_  = A167 & A168;
  assign \new_[9774]_  = ~A202 & ~A201;
  assign \new_[9775]_  = \new_[9774]_  & \new_[9771]_ ;
  assign \new_[9778]_  = A233 & ~A203;
  assign \new_[9782]_  = A267 & A265;
  assign \new_[9783]_  = A234 & \new_[9782]_ ;
  assign \new_[9784]_  = \new_[9783]_  & \new_[9778]_ ;
  assign \new_[9787]_  = A167 & A168;
  assign \new_[9790]_  = ~A202 & ~A201;
  assign \new_[9791]_  = \new_[9790]_  & \new_[9787]_ ;
  assign \new_[9794]_  = A233 & ~A203;
  assign \new_[9798]_  = A267 & A266;
  assign \new_[9799]_  = A234 & \new_[9798]_ ;
  assign \new_[9800]_  = \new_[9799]_  & \new_[9794]_ ;
  assign \new_[9803]_  = A167 & A168;
  assign \new_[9806]_  = ~A202 & ~A201;
  assign \new_[9807]_  = \new_[9806]_  & \new_[9803]_ ;
  assign \new_[9810]_  = ~A232 & ~A203;
  assign \new_[9814]_  = A268 & A236;
  assign \new_[9815]_  = A233 & \new_[9814]_ ;
  assign \new_[9816]_  = \new_[9815]_  & \new_[9810]_ ;
  assign \new_[9819]_  = A167 & A168;
  assign \new_[9822]_  = ~A202 & ~A201;
  assign \new_[9823]_  = \new_[9822]_  & \new_[9819]_ ;
  assign \new_[9826]_  = A232 & ~A203;
  assign \new_[9830]_  = A268 & A236;
  assign \new_[9831]_  = ~A233 & \new_[9830]_ ;
  assign \new_[9832]_  = \new_[9831]_  & \new_[9826]_ ;
  assign \new_[9835]_  = A167 & A168;
  assign \new_[9838]_  = A200 & A199;
  assign \new_[9839]_  = \new_[9838]_  & \new_[9835]_ ;
  assign \new_[9842]_  = ~A202 & ~A201;
  assign \new_[9846]_  = A267 & A265;
  assign \new_[9847]_  = A235 & \new_[9846]_ ;
  assign \new_[9848]_  = \new_[9847]_  & \new_[9842]_ ;
  assign \new_[9851]_  = A167 & A168;
  assign \new_[9854]_  = A200 & A199;
  assign \new_[9855]_  = \new_[9854]_  & \new_[9851]_ ;
  assign \new_[9858]_  = ~A202 & ~A201;
  assign \new_[9862]_  = A267 & A266;
  assign \new_[9863]_  = A235 & \new_[9862]_ ;
  assign \new_[9864]_  = \new_[9863]_  & \new_[9858]_ ;
  assign \new_[9867]_  = A167 & A168;
  assign \new_[9870]_  = A200 & A199;
  assign \new_[9871]_  = \new_[9870]_  & \new_[9867]_ ;
  assign \new_[9874]_  = ~A202 & ~A201;
  assign \new_[9878]_  = A268 & A234;
  assign \new_[9879]_  = A232 & \new_[9878]_ ;
  assign \new_[9880]_  = \new_[9879]_  & \new_[9874]_ ;
  assign \new_[9883]_  = A167 & A168;
  assign \new_[9886]_  = A200 & A199;
  assign \new_[9887]_  = \new_[9886]_  & \new_[9883]_ ;
  assign \new_[9890]_  = ~A202 & ~A201;
  assign \new_[9894]_  = A268 & A234;
  assign \new_[9895]_  = A233 & \new_[9894]_ ;
  assign \new_[9896]_  = \new_[9895]_  & \new_[9890]_ ;
  assign \new_[9899]_  = A167 & A168;
  assign \new_[9902]_  = ~A200 & ~A199;
  assign \new_[9903]_  = \new_[9902]_  & \new_[9899]_ ;
  assign \new_[9906]_  = A235 & ~A202;
  assign \new_[9910]_  = ~A302 & ~A301;
  assign \new_[9911]_  = ~A300 & \new_[9910]_ ;
  assign \new_[9912]_  = \new_[9911]_  & \new_[9906]_ ;
  assign \new_[9915]_  = A167 & A168;
  assign \new_[9918]_  = ~A200 & ~A199;
  assign \new_[9919]_  = \new_[9918]_  & \new_[9915]_ ;
  assign \new_[9922]_  = A235 & ~A202;
  assign \new_[9926]_  = ~A301 & ~A299;
  assign \new_[9927]_  = ~A298 & \new_[9926]_ ;
  assign \new_[9928]_  = \new_[9927]_  & \new_[9922]_ ;
  assign \new_[9931]_  = A167 & A168;
  assign \new_[9934]_  = ~A200 & ~A199;
  assign \new_[9935]_  = \new_[9934]_  & \new_[9931]_ ;
  assign \new_[9938]_  = A235 & ~A202;
  assign \new_[9942]_  = A269 & A266;
  assign \new_[9943]_  = ~A265 & \new_[9942]_ ;
  assign \new_[9944]_  = \new_[9943]_  & \new_[9938]_ ;
  assign \new_[9947]_  = A167 & A168;
  assign \new_[9950]_  = ~A200 & ~A199;
  assign \new_[9951]_  = \new_[9950]_  & \new_[9947]_ ;
  assign \new_[9954]_  = A235 & ~A202;
  assign \new_[9958]_  = A269 & ~A266;
  assign \new_[9959]_  = A265 & \new_[9958]_ ;
  assign \new_[9960]_  = \new_[9959]_  & \new_[9954]_ ;
  assign \new_[9963]_  = A167 & A168;
  assign \new_[9966]_  = ~A200 & ~A199;
  assign \new_[9967]_  = \new_[9966]_  & \new_[9963]_ ;
  assign \new_[9970]_  = A232 & ~A202;
  assign \new_[9974]_  = A267 & A265;
  assign \new_[9975]_  = A234 & \new_[9974]_ ;
  assign \new_[9976]_  = \new_[9975]_  & \new_[9970]_ ;
  assign \new_[9979]_  = A167 & A168;
  assign \new_[9982]_  = ~A200 & ~A199;
  assign \new_[9983]_  = \new_[9982]_  & \new_[9979]_ ;
  assign \new_[9986]_  = A232 & ~A202;
  assign \new_[9990]_  = A267 & A266;
  assign \new_[9991]_  = A234 & \new_[9990]_ ;
  assign \new_[9992]_  = \new_[9991]_  & \new_[9986]_ ;
  assign \new_[9995]_  = A167 & A168;
  assign \new_[9998]_  = ~A200 & ~A199;
  assign \new_[9999]_  = \new_[9998]_  & \new_[9995]_ ;
  assign \new_[10002]_  = A233 & ~A202;
  assign \new_[10006]_  = A267 & A265;
  assign \new_[10007]_  = A234 & \new_[10006]_ ;
  assign \new_[10008]_  = \new_[10007]_  & \new_[10002]_ ;
  assign \new_[10011]_  = A167 & A168;
  assign \new_[10014]_  = ~A200 & ~A199;
  assign \new_[10015]_  = \new_[10014]_  & \new_[10011]_ ;
  assign \new_[10018]_  = A233 & ~A202;
  assign \new_[10022]_  = A267 & A266;
  assign \new_[10023]_  = A234 & \new_[10022]_ ;
  assign \new_[10024]_  = \new_[10023]_  & \new_[10018]_ ;
  assign \new_[10027]_  = A167 & A168;
  assign \new_[10030]_  = ~A200 & ~A199;
  assign \new_[10031]_  = \new_[10030]_  & \new_[10027]_ ;
  assign \new_[10034]_  = ~A232 & ~A202;
  assign \new_[10038]_  = A268 & A236;
  assign \new_[10039]_  = A233 & \new_[10038]_ ;
  assign \new_[10040]_  = \new_[10039]_  & \new_[10034]_ ;
  assign \new_[10043]_  = A167 & A168;
  assign \new_[10046]_  = ~A200 & ~A199;
  assign \new_[10047]_  = \new_[10046]_  & \new_[10043]_ ;
  assign \new_[10050]_  = A232 & ~A202;
  assign \new_[10054]_  = A268 & A236;
  assign \new_[10055]_  = ~A233 & \new_[10054]_ ;
  assign \new_[10056]_  = \new_[10055]_  & \new_[10050]_ ;
  assign \new_[10059]_  = A167 & A170;
  assign \new_[10062]_  = ~A201 & ~A166;
  assign \new_[10063]_  = \new_[10062]_  & \new_[10059]_ ;
  assign \new_[10066]_  = ~A203 & ~A202;
  assign \new_[10070]_  = A267 & A265;
  assign \new_[10071]_  = A235 & \new_[10070]_ ;
  assign \new_[10072]_  = \new_[10071]_  & \new_[10066]_ ;
  assign \new_[10075]_  = A167 & A170;
  assign \new_[10078]_  = ~A201 & ~A166;
  assign \new_[10079]_  = \new_[10078]_  & \new_[10075]_ ;
  assign \new_[10082]_  = ~A203 & ~A202;
  assign \new_[10086]_  = A267 & A266;
  assign \new_[10087]_  = A235 & \new_[10086]_ ;
  assign \new_[10088]_  = \new_[10087]_  & \new_[10082]_ ;
  assign \new_[10091]_  = A167 & A170;
  assign \new_[10094]_  = ~A201 & ~A166;
  assign \new_[10095]_  = \new_[10094]_  & \new_[10091]_ ;
  assign \new_[10098]_  = ~A203 & ~A202;
  assign \new_[10102]_  = A268 & A234;
  assign \new_[10103]_  = A232 & \new_[10102]_ ;
  assign \new_[10104]_  = \new_[10103]_  & \new_[10098]_ ;
  assign \new_[10107]_  = A167 & A170;
  assign \new_[10110]_  = ~A201 & ~A166;
  assign \new_[10111]_  = \new_[10110]_  & \new_[10107]_ ;
  assign \new_[10114]_  = ~A203 & ~A202;
  assign \new_[10118]_  = A268 & A234;
  assign \new_[10119]_  = A233 & \new_[10118]_ ;
  assign \new_[10120]_  = \new_[10119]_  & \new_[10114]_ ;
  assign \new_[10123]_  = A167 & A170;
  assign \new_[10126]_  = A199 & ~A166;
  assign \new_[10127]_  = \new_[10126]_  & \new_[10123]_ ;
  assign \new_[10130]_  = ~A201 & A200;
  assign \new_[10134]_  = A268 & A235;
  assign \new_[10135]_  = ~A202 & \new_[10134]_ ;
  assign \new_[10136]_  = \new_[10135]_  & \new_[10130]_ ;
  assign \new_[10139]_  = A167 & A170;
  assign \new_[10142]_  = ~A199 & ~A166;
  assign \new_[10143]_  = \new_[10142]_  & \new_[10139]_ ;
  assign \new_[10146]_  = ~A202 & ~A200;
  assign \new_[10150]_  = A267 & A265;
  assign \new_[10151]_  = A235 & \new_[10150]_ ;
  assign \new_[10152]_  = \new_[10151]_  & \new_[10146]_ ;
  assign \new_[10155]_  = A167 & A170;
  assign \new_[10158]_  = ~A199 & ~A166;
  assign \new_[10159]_  = \new_[10158]_  & \new_[10155]_ ;
  assign \new_[10162]_  = ~A202 & ~A200;
  assign \new_[10166]_  = A267 & A266;
  assign \new_[10167]_  = A235 & \new_[10166]_ ;
  assign \new_[10168]_  = \new_[10167]_  & \new_[10162]_ ;
  assign \new_[10171]_  = A167 & A170;
  assign \new_[10174]_  = ~A199 & ~A166;
  assign \new_[10175]_  = \new_[10174]_  & \new_[10171]_ ;
  assign \new_[10178]_  = ~A202 & ~A200;
  assign \new_[10182]_  = A268 & A234;
  assign \new_[10183]_  = A232 & \new_[10182]_ ;
  assign \new_[10184]_  = \new_[10183]_  & \new_[10178]_ ;
  assign \new_[10187]_  = A167 & A170;
  assign \new_[10190]_  = ~A199 & ~A166;
  assign \new_[10191]_  = \new_[10190]_  & \new_[10187]_ ;
  assign \new_[10194]_  = ~A202 & ~A200;
  assign \new_[10198]_  = A268 & A234;
  assign \new_[10199]_  = A233 & \new_[10198]_ ;
  assign \new_[10200]_  = \new_[10199]_  & \new_[10194]_ ;
  assign \new_[10203]_  = ~A167 & A170;
  assign \new_[10206]_  = ~A201 & A166;
  assign \new_[10207]_  = \new_[10206]_  & \new_[10203]_ ;
  assign \new_[10210]_  = ~A203 & ~A202;
  assign \new_[10214]_  = A267 & A265;
  assign \new_[10215]_  = A235 & \new_[10214]_ ;
  assign \new_[10216]_  = \new_[10215]_  & \new_[10210]_ ;
  assign \new_[10219]_  = ~A167 & A170;
  assign \new_[10222]_  = ~A201 & A166;
  assign \new_[10223]_  = \new_[10222]_  & \new_[10219]_ ;
  assign \new_[10226]_  = ~A203 & ~A202;
  assign \new_[10230]_  = A267 & A266;
  assign \new_[10231]_  = A235 & \new_[10230]_ ;
  assign \new_[10232]_  = \new_[10231]_  & \new_[10226]_ ;
  assign \new_[10235]_  = ~A167 & A170;
  assign \new_[10238]_  = ~A201 & A166;
  assign \new_[10239]_  = \new_[10238]_  & \new_[10235]_ ;
  assign \new_[10242]_  = ~A203 & ~A202;
  assign \new_[10246]_  = A268 & A234;
  assign \new_[10247]_  = A232 & \new_[10246]_ ;
  assign \new_[10248]_  = \new_[10247]_  & \new_[10242]_ ;
  assign \new_[10251]_  = ~A167 & A170;
  assign \new_[10254]_  = ~A201 & A166;
  assign \new_[10255]_  = \new_[10254]_  & \new_[10251]_ ;
  assign \new_[10258]_  = ~A203 & ~A202;
  assign \new_[10262]_  = A268 & A234;
  assign \new_[10263]_  = A233 & \new_[10262]_ ;
  assign \new_[10264]_  = \new_[10263]_  & \new_[10258]_ ;
  assign \new_[10267]_  = ~A167 & A170;
  assign \new_[10270]_  = A199 & A166;
  assign \new_[10271]_  = \new_[10270]_  & \new_[10267]_ ;
  assign \new_[10274]_  = ~A201 & A200;
  assign \new_[10278]_  = A268 & A235;
  assign \new_[10279]_  = ~A202 & \new_[10278]_ ;
  assign \new_[10280]_  = \new_[10279]_  & \new_[10274]_ ;
  assign \new_[10283]_  = ~A167 & A170;
  assign \new_[10286]_  = ~A199 & A166;
  assign \new_[10287]_  = \new_[10286]_  & \new_[10283]_ ;
  assign \new_[10290]_  = ~A202 & ~A200;
  assign \new_[10294]_  = A267 & A265;
  assign \new_[10295]_  = A235 & \new_[10294]_ ;
  assign \new_[10296]_  = \new_[10295]_  & \new_[10290]_ ;
  assign \new_[10299]_  = ~A167 & A170;
  assign \new_[10302]_  = ~A199 & A166;
  assign \new_[10303]_  = \new_[10302]_  & \new_[10299]_ ;
  assign \new_[10306]_  = ~A202 & ~A200;
  assign \new_[10310]_  = A267 & A266;
  assign \new_[10311]_  = A235 & \new_[10310]_ ;
  assign \new_[10312]_  = \new_[10311]_  & \new_[10306]_ ;
  assign \new_[10315]_  = ~A167 & A170;
  assign \new_[10318]_  = ~A199 & A166;
  assign \new_[10319]_  = \new_[10318]_  & \new_[10315]_ ;
  assign \new_[10322]_  = ~A202 & ~A200;
  assign \new_[10326]_  = A268 & A234;
  assign \new_[10327]_  = A232 & \new_[10326]_ ;
  assign \new_[10328]_  = \new_[10327]_  & \new_[10322]_ ;
  assign \new_[10331]_  = ~A167 & A170;
  assign \new_[10334]_  = ~A199 & A166;
  assign \new_[10335]_  = \new_[10334]_  & \new_[10331]_ ;
  assign \new_[10338]_  = ~A202 & ~A200;
  assign \new_[10342]_  = A268 & A234;
  assign \new_[10343]_  = A233 & \new_[10342]_ ;
  assign \new_[10344]_  = \new_[10343]_  & \new_[10338]_ ;
  assign \new_[10347]_  = ~A201 & A169;
  assign \new_[10350]_  = ~A203 & ~A202;
  assign \new_[10351]_  = \new_[10350]_  & \new_[10347]_ ;
  assign \new_[10354]_  = A298 & A235;
  assign \new_[10358]_  = ~A301 & ~A300;
  assign \new_[10359]_  = A299 & \new_[10358]_ ;
  assign \new_[10360]_  = \new_[10359]_  & \new_[10354]_ ;
  assign \new_[10363]_  = ~A201 & A169;
  assign \new_[10366]_  = ~A203 & ~A202;
  assign \new_[10367]_  = \new_[10366]_  & \new_[10363]_ ;
  assign \new_[10370]_  = A234 & A232;
  assign \new_[10374]_  = ~A302 & ~A301;
  assign \new_[10375]_  = ~A300 & \new_[10374]_ ;
  assign \new_[10376]_  = \new_[10375]_  & \new_[10370]_ ;
  assign \new_[10379]_  = ~A201 & A169;
  assign \new_[10382]_  = ~A203 & ~A202;
  assign \new_[10383]_  = \new_[10382]_  & \new_[10379]_ ;
  assign \new_[10386]_  = A234 & A232;
  assign \new_[10390]_  = ~A301 & ~A299;
  assign \new_[10391]_  = ~A298 & \new_[10390]_ ;
  assign \new_[10392]_  = \new_[10391]_  & \new_[10386]_ ;
  assign \new_[10395]_  = ~A201 & A169;
  assign \new_[10398]_  = ~A203 & ~A202;
  assign \new_[10399]_  = \new_[10398]_  & \new_[10395]_ ;
  assign \new_[10402]_  = A234 & A232;
  assign \new_[10406]_  = A269 & A266;
  assign \new_[10407]_  = ~A265 & \new_[10406]_ ;
  assign \new_[10408]_  = \new_[10407]_  & \new_[10402]_ ;
  assign \new_[10411]_  = ~A201 & A169;
  assign \new_[10414]_  = ~A203 & ~A202;
  assign \new_[10415]_  = \new_[10414]_  & \new_[10411]_ ;
  assign \new_[10418]_  = A234 & A232;
  assign \new_[10422]_  = A269 & ~A266;
  assign \new_[10423]_  = A265 & \new_[10422]_ ;
  assign \new_[10424]_  = \new_[10423]_  & \new_[10418]_ ;
  assign \new_[10427]_  = ~A201 & A169;
  assign \new_[10430]_  = ~A203 & ~A202;
  assign \new_[10431]_  = \new_[10430]_  & \new_[10427]_ ;
  assign \new_[10434]_  = A234 & A233;
  assign \new_[10438]_  = ~A302 & ~A301;
  assign \new_[10439]_  = ~A300 & \new_[10438]_ ;
  assign \new_[10440]_  = \new_[10439]_  & \new_[10434]_ ;
  assign \new_[10443]_  = ~A201 & A169;
  assign \new_[10446]_  = ~A203 & ~A202;
  assign \new_[10447]_  = \new_[10446]_  & \new_[10443]_ ;
  assign \new_[10450]_  = A234 & A233;
  assign \new_[10454]_  = ~A301 & ~A299;
  assign \new_[10455]_  = ~A298 & \new_[10454]_ ;
  assign \new_[10456]_  = \new_[10455]_  & \new_[10450]_ ;
  assign \new_[10459]_  = ~A201 & A169;
  assign \new_[10462]_  = ~A203 & ~A202;
  assign \new_[10463]_  = \new_[10462]_  & \new_[10459]_ ;
  assign \new_[10466]_  = A234 & A233;
  assign \new_[10470]_  = A269 & A266;
  assign \new_[10471]_  = ~A265 & \new_[10470]_ ;
  assign \new_[10472]_  = \new_[10471]_  & \new_[10466]_ ;
  assign \new_[10475]_  = ~A201 & A169;
  assign \new_[10478]_  = ~A203 & ~A202;
  assign \new_[10479]_  = \new_[10478]_  & \new_[10475]_ ;
  assign \new_[10482]_  = A234 & A233;
  assign \new_[10486]_  = A269 & ~A266;
  assign \new_[10487]_  = A265 & \new_[10486]_ ;
  assign \new_[10488]_  = \new_[10487]_  & \new_[10482]_ ;
  assign \new_[10491]_  = ~A201 & A169;
  assign \new_[10494]_  = ~A203 & ~A202;
  assign \new_[10495]_  = \new_[10494]_  & \new_[10491]_ ;
  assign \new_[10498]_  = A233 & ~A232;
  assign \new_[10502]_  = A267 & A265;
  assign \new_[10503]_  = A236 & \new_[10502]_ ;
  assign \new_[10504]_  = \new_[10503]_  & \new_[10498]_ ;
  assign \new_[10507]_  = ~A201 & A169;
  assign \new_[10510]_  = ~A203 & ~A202;
  assign \new_[10511]_  = \new_[10510]_  & \new_[10507]_ ;
  assign \new_[10514]_  = A233 & ~A232;
  assign \new_[10518]_  = A267 & A266;
  assign \new_[10519]_  = A236 & \new_[10518]_ ;
  assign \new_[10520]_  = \new_[10519]_  & \new_[10514]_ ;
  assign \new_[10523]_  = ~A201 & A169;
  assign \new_[10526]_  = ~A203 & ~A202;
  assign \new_[10527]_  = \new_[10526]_  & \new_[10523]_ ;
  assign \new_[10530]_  = ~A233 & A232;
  assign \new_[10534]_  = A267 & A265;
  assign \new_[10535]_  = A236 & \new_[10534]_ ;
  assign \new_[10536]_  = \new_[10535]_  & \new_[10530]_ ;
  assign \new_[10539]_  = ~A201 & A169;
  assign \new_[10542]_  = ~A203 & ~A202;
  assign \new_[10543]_  = \new_[10542]_  & \new_[10539]_ ;
  assign \new_[10546]_  = ~A233 & A232;
  assign \new_[10550]_  = A267 & A266;
  assign \new_[10551]_  = A236 & \new_[10550]_ ;
  assign \new_[10552]_  = \new_[10551]_  & \new_[10546]_ ;
  assign \new_[10555]_  = A199 & A169;
  assign \new_[10558]_  = ~A201 & A200;
  assign \new_[10559]_  = \new_[10558]_  & \new_[10555]_ ;
  assign \new_[10562]_  = A235 & ~A202;
  assign \new_[10566]_  = ~A302 & ~A301;
  assign \new_[10567]_  = ~A300 & \new_[10566]_ ;
  assign \new_[10568]_  = \new_[10567]_  & \new_[10562]_ ;
  assign \new_[10571]_  = A199 & A169;
  assign \new_[10574]_  = ~A201 & A200;
  assign \new_[10575]_  = \new_[10574]_  & \new_[10571]_ ;
  assign \new_[10578]_  = A235 & ~A202;
  assign \new_[10582]_  = ~A301 & ~A299;
  assign \new_[10583]_  = ~A298 & \new_[10582]_ ;
  assign \new_[10584]_  = \new_[10583]_  & \new_[10578]_ ;
  assign \new_[10587]_  = A199 & A169;
  assign \new_[10590]_  = ~A201 & A200;
  assign \new_[10591]_  = \new_[10590]_  & \new_[10587]_ ;
  assign \new_[10594]_  = A235 & ~A202;
  assign \new_[10598]_  = A269 & A266;
  assign \new_[10599]_  = ~A265 & \new_[10598]_ ;
  assign \new_[10600]_  = \new_[10599]_  & \new_[10594]_ ;
  assign \new_[10603]_  = A199 & A169;
  assign \new_[10606]_  = ~A201 & A200;
  assign \new_[10607]_  = \new_[10606]_  & \new_[10603]_ ;
  assign \new_[10610]_  = A235 & ~A202;
  assign \new_[10614]_  = A269 & ~A266;
  assign \new_[10615]_  = A265 & \new_[10614]_ ;
  assign \new_[10616]_  = \new_[10615]_  & \new_[10610]_ ;
  assign \new_[10619]_  = A199 & A169;
  assign \new_[10622]_  = ~A201 & A200;
  assign \new_[10623]_  = \new_[10622]_  & \new_[10619]_ ;
  assign \new_[10626]_  = A232 & ~A202;
  assign \new_[10630]_  = A267 & A265;
  assign \new_[10631]_  = A234 & \new_[10630]_ ;
  assign \new_[10632]_  = \new_[10631]_  & \new_[10626]_ ;
  assign \new_[10635]_  = A199 & A169;
  assign \new_[10638]_  = ~A201 & A200;
  assign \new_[10639]_  = \new_[10638]_  & \new_[10635]_ ;
  assign \new_[10642]_  = A232 & ~A202;
  assign \new_[10646]_  = A267 & A266;
  assign \new_[10647]_  = A234 & \new_[10646]_ ;
  assign \new_[10648]_  = \new_[10647]_  & \new_[10642]_ ;
  assign \new_[10651]_  = A199 & A169;
  assign \new_[10654]_  = ~A201 & A200;
  assign \new_[10655]_  = \new_[10654]_  & \new_[10651]_ ;
  assign \new_[10658]_  = A233 & ~A202;
  assign \new_[10662]_  = A267 & A265;
  assign \new_[10663]_  = A234 & \new_[10662]_ ;
  assign \new_[10664]_  = \new_[10663]_  & \new_[10658]_ ;
  assign \new_[10667]_  = A199 & A169;
  assign \new_[10670]_  = ~A201 & A200;
  assign \new_[10671]_  = \new_[10670]_  & \new_[10667]_ ;
  assign \new_[10674]_  = A233 & ~A202;
  assign \new_[10678]_  = A267 & A266;
  assign \new_[10679]_  = A234 & \new_[10678]_ ;
  assign \new_[10680]_  = \new_[10679]_  & \new_[10674]_ ;
  assign \new_[10683]_  = A199 & A169;
  assign \new_[10686]_  = ~A201 & A200;
  assign \new_[10687]_  = \new_[10686]_  & \new_[10683]_ ;
  assign \new_[10690]_  = ~A232 & ~A202;
  assign \new_[10694]_  = A268 & A236;
  assign \new_[10695]_  = A233 & \new_[10694]_ ;
  assign \new_[10696]_  = \new_[10695]_  & \new_[10690]_ ;
  assign \new_[10699]_  = A199 & A169;
  assign \new_[10702]_  = ~A201 & A200;
  assign \new_[10703]_  = \new_[10702]_  & \new_[10699]_ ;
  assign \new_[10706]_  = A232 & ~A202;
  assign \new_[10710]_  = A268 & A236;
  assign \new_[10711]_  = ~A233 & \new_[10710]_ ;
  assign \new_[10712]_  = \new_[10711]_  & \new_[10706]_ ;
  assign \new_[10715]_  = ~A199 & A169;
  assign \new_[10718]_  = ~A202 & ~A200;
  assign \new_[10719]_  = \new_[10718]_  & \new_[10715]_ ;
  assign \new_[10722]_  = A298 & A235;
  assign \new_[10726]_  = ~A301 & ~A300;
  assign \new_[10727]_  = A299 & \new_[10726]_ ;
  assign \new_[10728]_  = \new_[10727]_  & \new_[10722]_ ;
  assign \new_[10731]_  = ~A199 & A169;
  assign \new_[10734]_  = ~A202 & ~A200;
  assign \new_[10735]_  = \new_[10734]_  & \new_[10731]_ ;
  assign \new_[10738]_  = A234 & A232;
  assign \new_[10742]_  = ~A302 & ~A301;
  assign \new_[10743]_  = ~A300 & \new_[10742]_ ;
  assign \new_[10744]_  = \new_[10743]_  & \new_[10738]_ ;
  assign \new_[10747]_  = ~A199 & A169;
  assign \new_[10750]_  = ~A202 & ~A200;
  assign \new_[10751]_  = \new_[10750]_  & \new_[10747]_ ;
  assign \new_[10754]_  = A234 & A232;
  assign \new_[10758]_  = ~A301 & ~A299;
  assign \new_[10759]_  = ~A298 & \new_[10758]_ ;
  assign \new_[10760]_  = \new_[10759]_  & \new_[10754]_ ;
  assign \new_[10763]_  = ~A199 & A169;
  assign \new_[10766]_  = ~A202 & ~A200;
  assign \new_[10767]_  = \new_[10766]_  & \new_[10763]_ ;
  assign \new_[10770]_  = A234 & A232;
  assign \new_[10774]_  = A269 & A266;
  assign \new_[10775]_  = ~A265 & \new_[10774]_ ;
  assign \new_[10776]_  = \new_[10775]_  & \new_[10770]_ ;
  assign \new_[10779]_  = ~A199 & A169;
  assign \new_[10782]_  = ~A202 & ~A200;
  assign \new_[10783]_  = \new_[10782]_  & \new_[10779]_ ;
  assign \new_[10786]_  = A234 & A232;
  assign \new_[10790]_  = A269 & ~A266;
  assign \new_[10791]_  = A265 & \new_[10790]_ ;
  assign \new_[10792]_  = \new_[10791]_  & \new_[10786]_ ;
  assign \new_[10795]_  = ~A199 & A169;
  assign \new_[10798]_  = ~A202 & ~A200;
  assign \new_[10799]_  = \new_[10798]_  & \new_[10795]_ ;
  assign \new_[10802]_  = A234 & A233;
  assign \new_[10806]_  = ~A302 & ~A301;
  assign \new_[10807]_  = ~A300 & \new_[10806]_ ;
  assign \new_[10808]_  = \new_[10807]_  & \new_[10802]_ ;
  assign \new_[10811]_  = ~A199 & A169;
  assign \new_[10814]_  = ~A202 & ~A200;
  assign \new_[10815]_  = \new_[10814]_  & \new_[10811]_ ;
  assign \new_[10818]_  = A234 & A233;
  assign \new_[10822]_  = ~A301 & ~A299;
  assign \new_[10823]_  = ~A298 & \new_[10822]_ ;
  assign \new_[10824]_  = \new_[10823]_  & \new_[10818]_ ;
  assign \new_[10827]_  = ~A199 & A169;
  assign \new_[10830]_  = ~A202 & ~A200;
  assign \new_[10831]_  = \new_[10830]_  & \new_[10827]_ ;
  assign \new_[10834]_  = A234 & A233;
  assign \new_[10838]_  = A269 & A266;
  assign \new_[10839]_  = ~A265 & \new_[10838]_ ;
  assign \new_[10840]_  = \new_[10839]_  & \new_[10834]_ ;
  assign \new_[10843]_  = ~A199 & A169;
  assign \new_[10846]_  = ~A202 & ~A200;
  assign \new_[10847]_  = \new_[10846]_  & \new_[10843]_ ;
  assign \new_[10850]_  = A234 & A233;
  assign \new_[10854]_  = A269 & ~A266;
  assign \new_[10855]_  = A265 & \new_[10854]_ ;
  assign \new_[10856]_  = \new_[10855]_  & \new_[10850]_ ;
  assign \new_[10859]_  = ~A199 & A169;
  assign \new_[10862]_  = ~A202 & ~A200;
  assign \new_[10863]_  = \new_[10862]_  & \new_[10859]_ ;
  assign \new_[10866]_  = A233 & ~A232;
  assign \new_[10870]_  = A267 & A265;
  assign \new_[10871]_  = A236 & \new_[10870]_ ;
  assign \new_[10872]_  = \new_[10871]_  & \new_[10866]_ ;
  assign \new_[10875]_  = ~A199 & A169;
  assign \new_[10878]_  = ~A202 & ~A200;
  assign \new_[10879]_  = \new_[10878]_  & \new_[10875]_ ;
  assign \new_[10882]_  = A233 & ~A232;
  assign \new_[10886]_  = A267 & A266;
  assign \new_[10887]_  = A236 & \new_[10886]_ ;
  assign \new_[10888]_  = \new_[10887]_  & \new_[10882]_ ;
  assign \new_[10891]_  = ~A199 & A169;
  assign \new_[10894]_  = ~A202 & ~A200;
  assign \new_[10895]_  = \new_[10894]_  & \new_[10891]_ ;
  assign \new_[10898]_  = ~A233 & A232;
  assign \new_[10902]_  = A267 & A265;
  assign \new_[10903]_  = A236 & \new_[10902]_ ;
  assign \new_[10904]_  = \new_[10903]_  & \new_[10898]_ ;
  assign \new_[10907]_  = ~A199 & A169;
  assign \new_[10910]_  = ~A202 & ~A200;
  assign \new_[10911]_  = \new_[10910]_  & \new_[10907]_ ;
  assign \new_[10914]_  = ~A233 & A232;
  assign \new_[10918]_  = A267 & A266;
  assign \new_[10919]_  = A236 & \new_[10918]_ ;
  assign \new_[10920]_  = \new_[10919]_  & \new_[10914]_ ;
  assign \new_[10923]_  = ~A167 & ~A169;
  assign \new_[10926]_  = A202 & ~A166;
  assign \new_[10927]_  = \new_[10926]_  & \new_[10923]_ ;
  assign \new_[10930]_  = A298 & A235;
  assign \new_[10934]_  = ~A301 & ~A300;
  assign \new_[10935]_  = A299 & \new_[10934]_ ;
  assign \new_[10936]_  = \new_[10935]_  & \new_[10930]_ ;
  assign \new_[10939]_  = ~A167 & ~A169;
  assign \new_[10942]_  = A202 & ~A166;
  assign \new_[10943]_  = \new_[10942]_  & \new_[10939]_ ;
  assign \new_[10946]_  = A234 & A232;
  assign \new_[10950]_  = ~A302 & ~A301;
  assign \new_[10951]_  = ~A300 & \new_[10950]_ ;
  assign \new_[10952]_  = \new_[10951]_  & \new_[10946]_ ;
  assign \new_[10955]_  = ~A167 & ~A169;
  assign \new_[10958]_  = A202 & ~A166;
  assign \new_[10959]_  = \new_[10958]_  & \new_[10955]_ ;
  assign \new_[10962]_  = A234 & A232;
  assign \new_[10966]_  = ~A301 & ~A299;
  assign \new_[10967]_  = ~A298 & \new_[10966]_ ;
  assign \new_[10968]_  = \new_[10967]_  & \new_[10962]_ ;
  assign \new_[10971]_  = ~A167 & ~A169;
  assign \new_[10974]_  = A202 & ~A166;
  assign \new_[10975]_  = \new_[10974]_  & \new_[10971]_ ;
  assign \new_[10978]_  = A234 & A232;
  assign \new_[10982]_  = A269 & A266;
  assign \new_[10983]_  = ~A265 & \new_[10982]_ ;
  assign \new_[10984]_  = \new_[10983]_  & \new_[10978]_ ;
  assign \new_[10987]_  = ~A167 & ~A169;
  assign \new_[10990]_  = A202 & ~A166;
  assign \new_[10991]_  = \new_[10990]_  & \new_[10987]_ ;
  assign \new_[10994]_  = A234 & A232;
  assign \new_[10998]_  = A269 & ~A266;
  assign \new_[10999]_  = A265 & \new_[10998]_ ;
  assign \new_[11000]_  = \new_[10999]_  & \new_[10994]_ ;
  assign \new_[11003]_  = ~A167 & ~A169;
  assign \new_[11006]_  = A202 & ~A166;
  assign \new_[11007]_  = \new_[11006]_  & \new_[11003]_ ;
  assign \new_[11010]_  = A234 & A233;
  assign \new_[11014]_  = ~A302 & ~A301;
  assign \new_[11015]_  = ~A300 & \new_[11014]_ ;
  assign \new_[11016]_  = \new_[11015]_  & \new_[11010]_ ;
  assign \new_[11019]_  = ~A167 & ~A169;
  assign \new_[11022]_  = A202 & ~A166;
  assign \new_[11023]_  = \new_[11022]_  & \new_[11019]_ ;
  assign \new_[11026]_  = A234 & A233;
  assign \new_[11030]_  = ~A301 & ~A299;
  assign \new_[11031]_  = ~A298 & \new_[11030]_ ;
  assign \new_[11032]_  = \new_[11031]_  & \new_[11026]_ ;
  assign \new_[11035]_  = ~A167 & ~A169;
  assign \new_[11038]_  = A202 & ~A166;
  assign \new_[11039]_  = \new_[11038]_  & \new_[11035]_ ;
  assign \new_[11042]_  = A234 & A233;
  assign \new_[11046]_  = A269 & A266;
  assign \new_[11047]_  = ~A265 & \new_[11046]_ ;
  assign \new_[11048]_  = \new_[11047]_  & \new_[11042]_ ;
  assign \new_[11051]_  = ~A167 & ~A169;
  assign \new_[11054]_  = A202 & ~A166;
  assign \new_[11055]_  = \new_[11054]_  & \new_[11051]_ ;
  assign \new_[11058]_  = A234 & A233;
  assign \new_[11062]_  = A269 & ~A266;
  assign \new_[11063]_  = A265 & \new_[11062]_ ;
  assign \new_[11064]_  = \new_[11063]_  & \new_[11058]_ ;
  assign \new_[11067]_  = ~A167 & ~A169;
  assign \new_[11070]_  = A202 & ~A166;
  assign \new_[11071]_  = \new_[11070]_  & \new_[11067]_ ;
  assign \new_[11074]_  = A233 & ~A232;
  assign \new_[11078]_  = A267 & A265;
  assign \new_[11079]_  = A236 & \new_[11078]_ ;
  assign \new_[11080]_  = \new_[11079]_  & \new_[11074]_ ;
  assign \new_[11083]_  = ~A167 & ~A169;
  assign \new_[11086]_  = A202 & ~A166;
  assign \new_[11087]_  = \new_[11086]_  & \new_[11083]_ ;
  assign \new_[11090]_  = A233 & ~A232;
  assign \new_[11094]_  = A267 & A266;
  assign \new_[11095]_  = A236 & \new_[11094]_ ;
  assign \new_[11096]_  = \new_[11095]_  & \new_[11090]_ ;
  assign \new_[11099]_  = ~A167 & ~A169;
  assign \new_[11102]_  = A202 & ~A166;
  assign \new_[11103]_  = \new_[11102]_  & \new_[11099]_ ;
  assign \new_[11106]_  = ~A233 & A232;
  assign \new_[11110]_  = A267 & A265;
  assign \new_[11111]_  = A236 & \new_[11110]_ ;
  assign \new_[11112]_  = \new_[11111]_  & \new_[11106]_ ;
  assign \new_[11115]_  = ~A167 & ~A169;
  assign \new_[11118]_  = A202 & ~A166;
  assign \new_[11119]_  = \new_[11118]_  & \new_[11115]_ ;
  assign \new_[11122]_  = ~A233 & A232;
  assign \new_[11126]_  = A267 & A266;
  assign \new_[11127]_  = A236 & \new_[11126]_ ;
  assign \new_[11128]_  = \new_[11127]_  & \new_[11122]_ ;
  assign \new_[11131]_  = ~A167 & ~A169;
  assign \new_[11134]_  = A199 & ~A166;
  assign \new_[11135]_  = \new_[11134]_  & \new_[11131]_ ;
  assign \new_[11138]_  = A235 & A201;
  assign \new_[11142]_  = ~A302 & ~A301;
  assign \new_[11143]_  = ~A300 & \new_[11142]_ ;
  assign \new_[11144]_  = \new_[11143]_  & \new_[11138]_ ;
  assign \new_[11147]_  = ~A167 & ~A169;
  assign \new_[11150]_  = A199 & ~A166;
  assign \new_[11151]_  = \new_[11150]_  & \new_[11147]_ ;
  assign \new_[11154]_  = A235 & A201;
  assign \new_[11158]_  = ~A301 & ~A299;
  assign \new_[11159]_  = ~A298 & \new_[11158]_ ;
  assign \new_[11160]_  = \new_[11159]_  & \new_[11154]_ ;
  assign \new_[11163]_  = ~A167 & ~A169;
  assign \new_[11166]_  = A199 & ~A166;
  assign \new_[11167]_  = \new_[11166]_  & \new_[11163]_ ;
  assign \new_[11170]_  = A235 & A201;
  assign \new_[11174]_  = A269 & A266;
  assign \new_[11175]_  = ~A265 & \new_[11174]_ ;
  assign \new_[11176]_  = \new_[11175]_  & \new_[11170]_ ;
  assign \new_[11179]_  = ~A167 & ~A169;
  assign \new_[11182]_  = A199 & ~A166;
  assign \new_[11183]_  = \new_[11182]_  & \new_[11179]_ ;
  assign \new_[11186]_  = A235 & A201;
  assign \new_[11190]_  = A269 & ~A266;
  assign \new_[11191]_  = A265 & \new_[11190]_ ;
  assign \new_[11192]_  = \new_[11191]_  & \new_[11186]_ ;
  assign \new_[11195]_  = ~A167 & ~A169;
  assign \new_[11198]_  = A199 & ~A166;
  assign \new_[11199]_  = \new_[11198]_  & \new_[11195]_ ;
  assign \new_[11202]_  = A232 & A201;
  assign \new_[11206]_  = A267 & A265;
  assign \new_[11207]_  = A234 & \new_[11206]_ ;
  assign \new_[11208]_  = \new_[11207]_  & \new_[11202]_ ;
  assign \new_[11211]_  = ~A167 & ~A169;
  assign \new_[11214]_  = A199 & ~A166;
  assign \new_[11215]_  = \new_[11214]_  & \new_[11211]_ ;
  assign \new_[11218]_  = A232 & A201;
  assign \new_[11222]_  = A267 & A266;
  assign \new_[11223]_  = A234 & \new_[11222]_ ;
  assign \new_[11224]_  = \new_[11223]_  & \new_[11218]_ ;
  assign \new_[11227]_  = ~A167 & ~A169;
  assign \new_[11230]_  = A199 & ~A166;
  assign \new_[11231]_  = \new_[11230]_  & \new_[11227]_ ;
  assign \new_[11234]_  = A233 & A201;
  assign \new_[11238]_  = A267 & A265;
  assign \new_[11239]_  = A234 & \new_[11238]_ ;
  assign \new_[11240]_  = \new_[11239]_  & \new_[11234]_ ;
  assign \new_[11243]_  = ~A167 & ~A169;
  assign \new_[11246]_  = A199 & ~A166;
  assign \new_[11247]_  = \new_[11246]_  & \new_[11243]_ ;
  assign \new_[11250]_  = A233 & A201;
  assign \new_[11254]_  = A267 & A266;
  assign \new_[11255]_  = A234 & \new_[11254]_ ;
  assign \new_[11256]_  = \new_[11255]_  & \new_[11250]_ ;
  assign \new_[11259]_  = ~A167 & ~A169;
  assign \new_[11262]_  = A199 & ~A166;
  assign \new_[11263]_  = \new_[11262]_  & \new_[11259]_ ;
  assign \new_[11266]_  = ~A232 & A201;
  assign \new_[11270]_  = A268 & A236;
  assign \new_[11271]_  = A233 & \new_[11270]_ ;
  assign \new_[11272]_  = \new_[11271]_  & \new_[11266]_ ;
  assign \new_[11275]_  = ~A167 & ~A169;
  assign \new_[11278]_  = A199 & ~A166;
  assign \new_[11279]_  = \new_[11278]_  & \new_[11275]_ ;
  assign \new_[11282]_  = A232 & A201;
  assign \new_[11286]_  = A268 & A236;
  assign \new_[11287]_  = ~A233 & \new_[11286]_ ;
  assign \new_[11288]_  = \new_[11287]_  & \new_[11282]_ ;
  assign \new_[11291]_  = ~A167 & ~A169;
  assign \new_[11294]_  = A200 & ~A166;
  assign \new_[11295]_  = \new_[11294]_  & \new_[11291]_ ;
  assign \new_[11298]_  = A235 & A201;
  assign \new_[11302]_  = ~A302 & ~A301;
  assign \new_[11303]_  = ~A300 & \new_[11302]_ ;
  assign \new_[11304]_  = \new_[11303]_  & \new_[11298]_ ;
  assign \new_[11307]_  = ~A167 & ~A169;
  assign \new_[11310]_  = A200 & ~A166;
  assign \new_[11311]_  = \new_[11310]_  & \new_[11307]_ ;
  assign \new_[11314]_  = A235 & A201;
  assign \new_[11318]_  = ~A301 & ~A299;
  assign \new_[11319]_  = ~A298 & \new_[11318]_ ;
  assign \new_[11320]_  = \new_[11319]_  & \new_[11314]_ ;
  assign \new_[11323]_  = ~A167 & ~A169;
  assign \new_[11326]_  = A200 & ~A166;
  assign \new_[11327]_  = \new_[11326]_  & \new_[11323]_ ;
  assign \new_[11330]_  = A235 & A201;
  assign \new_[11334]_  = A269 & A266;
  assign \new_[11335]_  = ~A265 & \new_[11334]_ ;
  assign \new_[11336]_  = \new_[11335]_  & \new_[11330]_ ;
  assign \new_[11339]_  = ~A167 & ~A169;
  assign \new_[11342]_  = A200 & ~A166;
  assign \new_[11343]_  = \new_[11342]_  & \new_[11339]_ ;
  assign \new_[11346]_  = A235 & A201;
  assign \new_[11350]_  = A269 & ~A266;
  assign \new_[11351]_  = A265 & \new_[11350]_ ;
  assign \new_[11352]_  = \new_[11351]_  & \new_[11346]_ ;
  assign \new_[11355]_  = ~A167 & ~A169;
  assign \new_[11358]_  = A200 & ~A166;
  assign \new_[11359]_  = \new_[11358]_  & \new_[11355]_ ;
  assign \new_[11362]_  = A232 & A201;
  assign \new_[11366]_  = A267 & A265;
  assign \new_[11367]_  = A234 & \new_[11366]_ ;
  assign \new_[11368]_  = \new_[11367]_  & \new_[11362]_ ;
  assign \new_[11371]_  = ~A167 & ~A169;
  assign \new_[11374]_  = A200 & ~A166;
  assign \new_[11375]_  = \new_[11374]_  & \new_[11371]_ ;
  assign \new_[11378]_  = A232 & A201;
  assign \new_[11382]_  = A267 & A266;
  assign \new_[11383]_  = A234 & \new_[11382]_ ;
  assign \new_[11384]_  = \new_[11383]_  & \new_[11378]_ ;
  assign \new_[11387]_  = ~A167 & ~A169;
  assign \new_[11390]_  = A200 & ~A166;
  assign \new_[11391]_  = \new_[11390]_  & \new_[11387]_ ;
  assign \new_[11394]_  = A233 & A201;
  assign \new_[11398]_  = A267 & A265;
  assign \new_[11399]_  = A234 & \new_[11398]_ ;
  assign \new_[11400]_  = \new_[11399]_  & \new_[11394]_ ;
  assign \new_[11403]_  = ~A167 & ~A169;
  assign \new_[11406]_  = A200 & ~A166;
  assign \new_[11407]_  = \new_[11406]_  & \new_[11403]_ ;
  assign \new_[11410]_  = A233 & A201;
  assign \new_[11414]_  = A267 & A266;
  assign \new_[11415]_  = A234 & \new_[11414]_ ;
  assign \new_[11416]_  = \new_[11415]_  & \new_[11410]_ ;
  assign \new_[11419]_  = ~A167 & ~A169;
  assign \new_[11422]_  = A200 & ~A166;
  assign \new_[11423]_  = \new_[11422]_  & \new_[11419]_ ;
  assign \new_[11426]_  = ~A232 & A201;
  assign \new_[11430]_  = A268 & A236;
  assign \new_[11431]_  = A233 & \new_[11430]_ ;
  assign \new_[11432]_  = \new_[11431]_  & \new_[11426]_ ;
  assign \new_[11435]_  = ~A167 & ~A169;
  assign \new_[11438]_  = A200 & ~A166;
  assign \new_[11439]_  = \new_[11438]_  & \new_[11435]_ ;
  assign \new_[11442]_  = A232 & A201;
  assign \new_[11446]_  = A268 & A236;
  assign \new_[11447]_  = ~A233 & \new_[11446]_ ;
  assign \new_[11448]_  = \new_[11447]_  & \new_[11442]_ ;
  assign \new_[11451]_  = ~A167 & ~A169;
  assign \new_[11454]_  = ~A199 & ~A166;
  assign \new_[11455]_  = \new_[11454]_  & \new_[11451]_ ;
  assign \new_[11458]_  = A203 & A200;
  assign \new_[11462]_  = A267 & A265;
  assign \new_[11463]_  = A235 & \new_[11462]_ ;
  assign \new_[11464]_  = \new_[11463]_  & \new_[11458]_ ;
  assign \new_[11467]_  = ~A167 & ~A169;
  assign \new_[11470]_  = ~A199 & ~A166;
  assign \new_[11471]_  = \new_[11470]_  & \new_[11467]_ ;
  assign \new_[11474]_  = A203 & A200;
  assign \new_[11478]_  = A267 & A266;
  assign \new_[11479]_  = A235 & \new_[11478]_ ;
  assign \new_[11480]_  = \new_[11479]_  & \new_[11474]_ ;
  assign \new_[11483]_  = ~A167 & ~A169;
  assign \new_[11486]_  = ~A199 & ~A166;
  assign \new_[11487]_  = \new_[11486]_  & \new_[11483]_ ;
  assign \new_[11490]_  = A203 & A200;
  assign \new_[11494]_  = A268 & A234;
  assign \new_[11495]_  = A232 & \new_[11494]_ ;
  assign \new_[11496]_  = \new_[11495]_  & \new_[11490]_ ;
  assign \new_[11499]_  = ~A167 & ~A169;
  assign \new_[11502]_  = ~A199 & ~A166;
  assign \new_[11503]_  = \new_[11502]_  & \new_[11499]_ ;
  assign \new_[11506]_  = A203 & A200;
  assign \new_[11510]_  = A268 & A234;
  assign \new_[11511]_  = A233 & \new_[11510]_ ;
  assign \new_[11512]_  = \new_[11511]_  & \new_[11506]_ ;
  assign \new_[11515]_  = ~A167 & ~A169;
  assign \new_[11518]_  = A199 & ~A166;
  assign \new_[11519]_  = \new_[11518]_  & \new_[11515]_ ;
  assign \new_[11522]_  = A203 & ~A200;
  assign \new_[11526]_  = A267 & A265;
  assign \new_[11527]_  = A235 & \new_[11526]_ ;
  assign \new_[11528]_  = \new_[11527]_  & \new_[11522]_ ;
  assign \new_[11531]_  = ~A167 & ~A169;
  assign \new_[11534]_  = A199 & ~A166;
  assign \new_[11535]_  = \new_[11534]_  & \new_[11531]_ ;
  assign \new_[11538]_  = A203 & ~A200;
  assign \new_[11542]_  = A267 & A266;
  assign \new_[11543]_  = A235 & \new_[11542]_ ;
  assign \new_[11544]_  = \new_[11543]_  & \new_[11538]_ ;
  assign \new_[11547]_  = ~A167 & ~A169;
  assign \new_[11550]_  = A199 & ~A166;
  assign \new_[11551]_  = \new_[11550]_  & \new_[11547]_ ;
  assign \new_[11554]_  = A203 & ~A200;
  assign \new_[11558]_  = A268 & A234;
  assign \new_[11559]_  = A232 & \new_[11558]_ ;
  assign \new_[11560]_  = \new_[11559]_  & \new_[11554]_ ;
  assign \new_[11563]_  = ~A167 & ~A169;
  assign \new_[11566]_  = A199 & ~A166;
  assign \new_[11567]_  = \new_[11566]_  & \new_[11563]_ ;
  assign \new_[11570]_  = A203 & ~A200;
  assign \new_[11574]_  = A268 & A234;
  assign \new_[11575]_  = A233 & \new_[11574]_ ;
  assign \new_[11576]_  = \new_[11575]_  & \new_[11570]_ ;
  assign \new_[11579]_  = ~A168 & ~A169;
  assign \new_[11582]_  = A166 & A167;
  assign \new_[11583]_  = \new_[11582]_  & \new_[11579]_ ;
  assign \new_[11586]_  = A235 & A202;
  assign \new_[11590]_  = ~A302 & ~A301;
  assign \new_[11591]_  = ~A300 & \new_[11590]_ ;
  assign \new_[11592]_  = \new_[11591]_  & \new_[11586]_ ;
  assign \new_[11595]_  = ~A168 & ~A169;
  assign \new_[11598]_  = A166 & A167;
  assign \new_[11599]_  = \new_[11598]_  & \new_[11595]_ ;
  assign \new_[11602]_  = A235 & A202;
  assign \new_[11606]_  = ~A301 & ~A299;
  assign \new_[11607]_  = ~A298 & \new_[11606]_ ;
  assign \new_[11608]_  = \new_[11607]_  & \new_[11602]_ ;
  assign \new_[11611]_  = ~A168 & ~A169;
  assign \new_[11614]_  = A166 & A167;
  assign \new_[11615]_  = \new_[11614]_  & \new_[11611]_ ;
  assign \new_[11618]_  = A235 & A202;
  assign \new_[11622]_  = A269 & A266;
  assign \new_[11623]_  = ~A265 & \new_[11622]_ ;
  assign \new_[11624]_  = \new_[11623]_  & \new_[11618]_ ;
  assign \new_[11627]_  = ~A168 & ~A169;
  assign \new_[11630]_  = A166 & A167;
  assign \new_[11631]_  = \new_[11630]_  & \new_[11627]_ ;
  assign \new_[11634]_  = A235 & A202;
  assign \new_[11638]_  = A269 & ~A266;
  assign \new_[11639]_  = A265 & \new_[11638]_ ;
  assign \new_[11640]_  = \new_[11639]_  & \new_[11634]_ ;
  assign \new_[11643]_  = ~A168 & ~A169;
  assign \new_[11646]_  = A166 & A167;
  assign \new_[11647]_  = \new_[11646]_  & \new_[11643]_ ;
  assign \new_[11650]_  = A232 & A202;
  assign \new_[11654]_  = A267 & A265;
  assign \new_[11655]_  = A234 & \new_[11654]_ ;
  assign \new_[11656]_  = \new_[11655]_  & \new_[11650]_ ;
  assign \new_[11659]_  = ~A168 & ~A169;
  assign \new_[11662]_  = A166 & A167;
  assign \new_[11663]_  = \new_[11662]_  & \new_[11659]_ ;
  assign \new_[11666]_  = A232 & A202;
  assign \new_[11670]_  = A267 & A266;
  assign \new_[11671]_  = A234 & \new_[11670]_ ;
  assign \new_[11672]_  = \new_[11671]_  & \new_[11666]_ ;
  assign \new_[11675]_  = ~A168 & ~A169;
  assign \new_[11678]_  = A166 & A167;
  assign \new_[11679]_  = \new_[11678]_  & \new_[11675]_ ;
  assign \new_[11682]_  = A233 & A202;
  assign \new_[11686]_  = A267 & A265;
  assign \new_[11687]_  = A234 & \new_[11686]_ ;
  assign \new_[11688]_  = \new_[11687]_  & \new_[11682]_ ;
  assign \new_[11691]_  = ~A168 & ~A169;
  assign \new_[11694]_  = A166 & A167;
  assign \new_[11695]_  = \new_[11694]_  & \new_[11691]_ ;
  assign \new_[11698]_  = A233 & A202;
  assign \new_[11702]_  = A267 & A266;
  assign \new_[11703]_  = A234 & \new_[11702]_ ;
  assign \new_[11704]_  = \new_[11703]_  & \new_[11698]_ ;
  assign \new_[11707]_  = ~A168 & ~A169;
  assign \new_[11710]_  = A166 & A167;
  assign \new_[11711]_  = \new_[11710]_  & \new_[11707]_ ;
  assign \new_[11714]_  = ~A232 & A202;
  assign \new_[11718]_  = A268 & A236;
  assign \new_[11719]_  = A233 & \new_[11718]_ ;
  assign \new_[11720]_  = \new_[11719]_  & \new_[11714]_ ;
  assign \new_[11723]_  = ~A168 & ~A169;
  assign \new_[11726]_  = A166 & A167;
  assign \new_[11727]_  = \new_[11726]_  & \new_[11723]_ ;
  assign \new_[11730]_  = A232 & A202;
  assign \new_[11734]_  = A268 & A236;
  assign \new_[11735]_  = ~A233 & \new_[11734]_ ;
  assign \new_[11736]_  = \new_[11735]_  & \new_[11730]_ ;
  assign \new_[11739]_  = ~A168 & ~A169;
  assign \new_[11742]_  = A166 & A167;
  assign \new_[11743]_  = \new_[11742]_  & \new_[11739]_ ;
  assign \new_[11746]_  = A201 & A199;
  assign \new_[11750]_  = A267 & A265;
  assign \new_[11751]_  = A235 & \new_[11750]_ ;
  assign \new_[11752]_  = \new_[11751]_  & \new_[11746]_ ;
  assign \new_[11755]_  = ~A168 & ~A169;
  assign \new_[11758]_  = A166 & A167;
  assign \new_[11759]_  = \new_[11758]_  & \new_[11755]_ ;
  assign \new_[11762]_  = A201 & A199;
  assign \new_[11766]_  = A267 & A266;
  assign \new_[11767]_  = A235 & \new_[11766]_ ;
  assign \new_[11768]_  = \new_[11767]_  & \new_[11762]_ ;
  assign \new_[11771]_  = ~A168 & ~A169;
  assign \new_[11774]_  = A166 & A167;
  assign \new_[11775]_  = \new_[11774]_  & \new_[11771]_ ;
  assign \new_[11778]_  = A201 & A199;
  assign \new_[11782]_  = A268 & A234;
  assign \new_[11783]_  = A232 & \new_[11782]_ ;
  assign \new_[11784]_  = \new_[11783]_  & \new_[11778]_ ;
  assign \new_[11787]_  = ~A168 & ~A169;
  assign \new_[11790]_  = A166 & A167;
  assign \new_[11791]_  = \new_[11790]_  & \new_[11787]_ ;
  assign \new_[11794]_  = A201 & A199;
  assign \new_[11798]_  = A268 & A234;
  assign \new_[11799]_  = A233 & \new_[11798]_ ;
  assign \new_[11800]_  = \new_[11799]_  & \new_[11794]_ ;
  assign \new_[11803]_  = ~A168 & ~A169;
  assign \new_[11806]_  = A166 & A167;
  assign \new_[11807]_  = \new_[11806]_  & \new_[11803]_ ;
  assign \new_[11810]_  = A201 & A200;
  assign \new_[11814]_  = A267 & A265;
  assign \new_[11815]_  = A235 & \new_[11814]_ ;
  assign \new_[11816]_  = \new_[11815]_  & \new_[11810]_ ;
  assign \new_[11819]_  = ~A168 & ~A169;
  assign \new_[11822]_  = A166 & A167;
  assign \new_[11823]_  = \new_[11822]_  & \new_[11819]_ ;
  assign \new_[11826]_  = A201 & A200;
  assign \new_[11830]_  = A267 & A266;
  assign \new_[11831]_  = A235 & \new_[11830]_ ;
  assign \new_[11832]_  = \new_[11831]_  & \new_[11826]_ ;
  assign \new_[11835]_  = ~A168 & ~A169;
  assign \new_[11838]_  = A166 & A167;
  assign \new_[11839]_  = \new_[11838]_  & \new_[11835]_ ;
  assign \new_[11842]_  = A201 & A200;
  assign \new_[11846]_  = A268 & A234;
  assign \new_[11847]_  = A232 & \new_[11846]_ ;
  assign \new_[11848]_  = \new_[11847]_  & \new_[11842]_ ;
  assign \new_[11851]_  = ~A168 & ~A169;
  assign \new_[11854]_  = A166 & A167;
  assign \new_[11855]_  = \new_[11854]_  & \new_[11851]_ ;
  assign \new_[11858]_  = A201 & A200;
  assign \new_[11862]_  = A268 & A234;
  assign \new_[11863]_  = A233 & \new_[11862]_ ;
  assign \new_[11864]_  = \new_[11863]_  & \new_[11858]_ ;
  assign \new_[11867]_  = ~A168 & ~A169;
  assign \new_[11870]_  = A166 & A167;
  assign \new_[11871]_  = \new_[11870]_  & \new_[11867]_ ;
  assign \new_[11874]_  = A200 & ~A199;
  assign \new_[11878]_  = A268 & A235;
  assign \new_[11879]_  = A203 & \new_[11878]_ ;
  assign \new_[11880]_  = \new_[11879]_  & \new_[11874]_ ;
  assign \new_[11883]_  = ~A168 & ~A169;
  assign \new_[11886]_  = A166 & A167;
  assign \new_[11887]_  = \new_[11886]_  & \new_[11883]_ ;
  assign \new_[11890]_  = ~A200 & A199;
  assign \new_[11894]_  = A268 & A235;
  assign \new_[11895]_  = A203 & \new_[11894]_ ;
  assign \new_[11896]_  = \new_[11895]_  & \new_[11890]_ ;
  assign \new_[11899]_  = ~A169 & ~A170;
  assign \new_[11902]_  = A202 & ~A168;
  assign \new_[11903]_  = \new_[11902]_  & \new_[11899]_ ;
  assign \new_[11906]_  = A298 & A235;
  assign \new_[11910]_  = ~A301 & ~A300;
  assign \new_[11911]_  = A299 & \new_[11910]_ ;
  assign \new_[11912]_  = \new_[11911]_  & \new_[11906]_ ;
  assign \new_[11915]_  = ~A169 & ~A170;
  assign \new_[11918]_  = A202 & ~A168;
  assign \new_[11919]_  = \new_[11918]_  & \new_[11915]_ ;
  assign \new_[11922]_  = A234 & A232;
  assign \new_[11926]_  = ~A302 & ~A301;
  assign \new_[11927]_  = ~A300 & \new_[11926]_ ;
  assign \new_[11928]_  = \new_[11927]_  & \new_[11922]_ ;
  assign \new_[11931]_  = ~A169 & ~A170;
  assign \new_[11934]_  = A202 & ~A168;
  assign \new_[11935]_  = \new_[11934]_  & \new_[11931]_ ;
  assign \new_[11938]_  = A234 & A232;
  assign \new_[11942]_  = ~A301 & ~A299;
  assign \new_[11943]_  = ~A298 & \new_[11942]_ ;
  assign \new_[11944]_  = \new_[11943]_  & \new_[11938]_ ;
  assign \new_[11947]_  = ~A169 & ~A170;
  assign \new_[11950]_  = A202 & ~A168;
  assign \new_[11951]_  = \new_[11950]_  & \new_[11947]_ ;
  assign \new_[11954]_  = A234 & A232;
  assign \new_[11958]_  = A269 & A266;
  assign \new_[11959]_  = ~A265 & \new_[11958]_ ;
  assign \new_[11960]_  = \new_[11959]_  & \new_[11954]_ ;
  assign \new_[11963]_  = ~A169 & ~A170;
  assign \new_[11966]_  = A202 & ~A168;
  assign \new_[11967]_  = \new_[11966]_  & \new_[11963]_ ;
  assign \new_[11970]_  = A234 & A232;
  assign \new_[11974]_  = A269 & ~A266;
  assign \new_[11975]_  = A265 & \new_[11974]_ ;
  assign \new_[11976]_  = \new_[11975]_  & \new_[11970]_ ;
  assign \new_[11979]_  = ~A169 & ~A170;
  assign \new_[11982]_  = A202 & ~A168;
  assign \new_[11983]_  = \new_[11982]_  & \new_[11979]_ ;
  assign \new_[11986]_  = A234 & A233;
  assign \new_[11990]_  = ~A302 & ~A301;
  assign \new_[11991]_  = ~A300 & \new_[11990]_ ;
  assign \new_[11992]_  = \new_[11991]_  & \new_[11986]_ ;
  assign \new_[11995]_  = ~A169 & ~A170;
  assign \new_[11998]_  = A202 & ~A168;
  assign \new_[11999]_  = \new_[11998]_  & \new_[11995]_ ;
  assign \new_[12002]_  = A234 & A233;
  assign \new_[12006]_  = ~A301 & ~A299;
  assign \new_[12007]_  = ~A298 & \new_[12006]_ ;
  assign \new_[12008]_  = \new_[12007]_  & \new_[12002]_ ;
  assign \new_[12011]_  = ~A169 & ~A170;
  assign \new_[12014]_  = A202 & ~A168;
  assign \new_[12015]_  = \new_[12014]_  & \new_[12011]_ ;
  assign \new_[12018]_  = A234 & A233;
  assign \new_[12022]_  = A269 & A266;
  assign \new_[12023]_  = ~A265 & \new_[12022]_ ;
  assign \new_[12024]_  = \new_[12023]_  & \new_[12018]_ ;
  assign \new_[12027]_  = ~A169 & ~A170;
  assign \new_[12030]_  = A202 & ~A168;
  assign \new_[12031]_  = \new_[12030]_  & \new_[12027]_ ;
  assign \new_[12034]_  = A234 & A233;
  assign \new_[12038]_  = A269 & ~A266;
  assign \new_[12039]_  = A265 & \new_[12038]_ ;
  assign \new_[12040]_  = \new_[12039]_  & \new_[12034]_ ;
  assign \new_[12043]_  = ~A169 & ~A170;
  assign \new_[12046]_  = A202 & ~A168;
  assign \new_[12047]_  = \new_[12046]_  & \new_[12043]_ ;
  assign \new_[12050]_  = A233 & ~A232;
  assign \new_[12054]_  = A267 & A265;
  assign \new_[12055]_  = A236 & \new_[12054]_ ;
  assign \new_[12056]_  = \new_[12055]_  & \new_[12050]_ ;
  assign \new_[12059]_  = ~A169 & ~A170;
  assign \new_[12062]_  = A202 & ~A168;
  assign \new_[12063]_  = \new_[12062]_  & \new_[12059]_ ;
  assign \new_[12066]_  = A233 & ~A232;
  assign \new_[12070]_  = A267 & A266;
  assign \new_[12071]_  = A236 & \new_[12070]_ ;
  assign \new_[12072]_  = \new_[12071]_  & \new_[12066]_ ;
  assign \new_[12075]_  = ~A169 & ~A170;
  assign \new_[12078]_  = A202 & ~A168;
  assign \new_[12079]_  = \new_[12078]_  & \new_[12075]_ ;
  assign \new_[12082]_  = ~A233 & A232;
  assign \new_[12086]_  = A267 & A265;
  assign \new_[12087]_  = A236 & \new_[12086]_ ;
  assign \new_[12088]_  = \new_[12087]_  & \new_[12082]_ ;
  assign \new_[12091]_  = ~A169 & ~A170;
  assign \new_[12094]_  = A202 & ~A168;
  assign \new_[12095]_  = \new_[12094]_  & \new_[12091]_ ;
  assign \new_[12098]_  = ~A233 & A232;
  assign \new_[12102]_  = A267 & A266;
  assign \new_[12103]_  = A236 & \new_[12102]_ ;
  assign \new_[12104]_  = \new_[12103]_  & \new_[12098]_ ;
  assign \new_[12107]_  = ~A169 & ~A170;
  assign \new_[12110]_  = A199 & ~A168;
  assign \new_[12111]_  = \new_[12110]_  & \new_[12107]_ ;
  assign \new_[12114]_  = A235 & A201;
  assign \new_[12118]_  = ~A302 & ~A301;
  assign \new_[12119]_  = ~A300 & \new_[12118]_ ;
  assign \new_[12120]_  = \new_[12119]_  & \new_[12114]_ ;
  assign \new_[12123]_  = ~A169 & ~A170;
  assign \new_[12126]_  = A199 & ~A168;
  assign \new_[12127]_  = \new_[12126]_  & \new_[12123]_ ;
  assign \new_[12130]_  = A235 & A201;
  assign \new_[12134]_  = ~A301 & ~A299;
  assign \new_[12135]_  = ~A298 & \new_[12134]_ ;
  assign \new_[12136]_  = \new_[12135]_  & \new_[12130]_ ;
  assign \new_[12139]_  = ~A169 & ~A170;
  assign \new_[12142]_  = A199 & ~A168;
  assign \new_[12143]_  = \new_[12142]_  & \new_[12139]_ ;
  assign \new_[12146]_  = A235 & A201;
  assign \new_[12150]_  = A269 & A266;
  assign \new_[12151]_  = ~A265 & \new_[12150]_ ;
  assign \new_[12152]_  = \new_[12151]_  & \new_[12146]_ ;
  assign \new_[12155]_  = ~A169 & ~A170;
  assign \new_[12158]_  = A199 & ~A168;
  assign \new_[12159]_  = \new_[12158]_  & \new_[12155]_ ;
  assign \new_[12162]_  = A235 & A201;
  assign \new_[12166]_  = A269 & ~A266;
  assign \new_[12167]_  = A265 & \new_[12166]_ ;
  assign \new_[12168]_  = \new_[12167]_  & \new_[12162]_ ;
  assign \new_[12171]_  = ~A169 & ~A170;
  assign \new_[12174]_  = A199 & ~A168;
  assign \new_[12175]_  = \new_[12174]_  & \new_[12171]_ ;
  assign \new_[12178]_  = A232 & A201;
  assign \new_[12182]_  = A267 & A265;
  assign \new_[12183]_  = A234 & \new_[12182]_ ;
  assign \new_[12184]_  = \new_[12183]_  & \new_[12178]_ ;
  assign \new_[12187]_  = ~A169 & ~A170;
  assign \new_[12190]_  = A199 & ~A168;
  assign \new_[12191]_  = \new_[12190]_  & \new_[12187]_ ;
  assign \new_[12194]_  = A232 & A201;
  assign \new_[12198]_  = A267 & A266;
  assign \new_[12199]_  = A234 & \new_[12198]_ ;
  assign \new_[12200]_  = \new_[12199]_  & \new_[12194]_ ;
  assign \new_[12203]_  = ~A169 & ~A170;
  assign \new_[12206]_  = A199 & ~A168;
  assign \new_[12207]_  = \new_[12206]_  & \new_[12203]_ ;
  assign \new_[12210]_  = A233 & A201;
  assign \new_[12214]_  = A267 & A265;
  assign \new_[12215]_  = A234 & \new_[12214]_ ;
  assign \new_[12216]_  = \new_[12215]_  & \new_[12210]_ ;
  assign \new_[12219]_  = ~A169 & ~A170;
  assign \new_[12222]_  = A199 & ~A168;
  assign \new_[12223]_  = \new_[12222]_  & \new_[12219]_ ;
  assign \new_[12226]_  = A233 & A201;
  assign \new_[12230]_  = A267 & A266;
  assign \new_[12231]_  = A234 & \new_[12230]_ ;
  assign \new_[12232]_  = \new_[12231]_  & \new_[12226]_ ;
  assign \new_[12235]_  = ~A169 & ~A170;
  assign \new_[12238]_  = A199 & ~A168;
  assign \new_[12239]_  = \new_[12238]_  & \new_[12235]_ ;
  assign \new_[12242]_  = ~A232 & A201;
  assign \new_[12246]_  = A268 & A236;
  assign \new_[12247]_  = A233 & \new_[12246]_ ;
  assign \new_[12248]_  = \new_[12247]_  & \new_[12242]_ ;
  assign \new_[12251]_  = ~A169 & ~A170;
  assign \new_[12254]_  = A199 & ~A168;
  assign \new_[12255]_  = \new_[12254]_  & \new_[12251]_ ;
  assign \new_[12258]_  = A232 & A201;
  assign \new_[12262]_  = A268 & A236;
  assign \new_[12263]_  = ~A233 & \new_[12262]_ ;
  assign \new_[12264]_  = \new_[12263]_  & \new_[12258]_ ;
  assign \new_[12267]_  = ~A169 & ~A170;
  assign \new_[12270]_  = A200 & ~A168;
  assign \new_[12271]_  = \new_[12270]_  & \new_[12267]_ ;
  assign \new_[12274]_  = A235 & A201;
  assign \new_[12278]_  = ~A302 & ~A301;
  assign \new_[12279]_  = ~A300 & \new_[12278]_ ;
  assign \new_[12280]_  = \new_[12279]_  & \new_[12274]_ ;
  assign \new_[12283]_  = ~A169 & ~A170;
  assign \new_[12286]_  = A200 & ~A168;
  assign \new_[12287]_  = \new_[12286]_  & \new_[12283]_ ;
  assign \new_[12290]_  = A235 & A201;
  assign \new_[12294]_  = ~A301 & ~A299;
  assign \new_[12295]_  = ~A298 & \new_[12294]_ ;
  assign \new_[12296]_  = \new_[12295]_  & \new_[12290]_ ;
  assign \new_[12299]_  = ~A169 & ~A170;
  assign \new_[12302]_  = A200 & ~A168;
  assign \new_[12303]_  = \new_[12302]_  & \new_[12299]_ ;
  assign \new_[12306]_  = A235 & A201;
  assign \new_[12310]_  = A269 & A266;
  assign \new_[12311]_  = ~A265 & \new_[12310]_ ;
  assign \new_[12312]_  = \new_[12311]_  & \new_[12306]_ ;
  assign \new_[12315]_  = ~A169 & ~A170;
  assign \new_[12318]_  = A200 & ~A168;
  assign \new_[12319]_  = \new_[12318]_  & \new_[12315]_ ;
  assign \new_[12322]_  = A235 & A201;
  assign \new_[12326]_  = A269 & ~A266;
  assign \new_[12327]_  = A265 & \new_[12326]_ ;
  assign \new_[12328]_  = \new_[12327]_  & \new_[12322]_ ;
  assign \new_[12331]_  = ~A169 & ~A170;
  assign \new_[12334]_  = A200 & ~A168;
  assign \new_[12335]_  = \new_[12334]_  & \new_[12331]_ ;
  assign \new_[12338]_  = A232 & A201;
  assign \new_[12342]_  = A267 & A265;
  assign \new_[12343]_  = A234 & \new_[12342]_ ;
  assign \new_[12344]_  = \new_[12343]_  & \new_[12338]_ ;
  assign \new_[12347]_  = ~A169 & ~A170;
  assign \new_[12350]_  = A200 & ~A168;
  assign \new_[12351]_  = \new_[12350]_  & \new_[12347]_ ;
  assign \new_[12354]_  = A232 & A201;
  assign \new_[12358]_  = A267 & A266;
  assign \new_[12359]_  = A234 & \new_[12358]_ ;
  assign \new_[12360]_  = \new_[12359]_  & \new_[12354]_ ;
  assign \new_[12363]_  = ~A169 & ~A170;
  assign \new_[12366]_  = A200 & ~A168;
  assign \new_[12367]_  = \new_[12366]_  & \new_[12363]_ ;
  assign \new_[12370]_  = A233 & A201;
  assign \new_[12374]_  = A267 & A265;
  assign \new_[12375]_  = A234 & \new_[12374]_ ;
  assign \new_[12376]_  = \new_[12375]_  & \new_[12370]_ ;
  assign \new_[12379]_  = ~A169 & ~A170;
  assign \new_[12382]_  = A200 & ~A168;
  assign \new_[12383]_  = \new_[12382]_  & \new_[12379]_ ;
  assign \new_[12386]_  = A233 & A201;
  assign \new_[12390]_  = A267 & A266;
  assign \new_[12391]_  = A234 & \new_[12390]_ ;
  assign \new_[12392]_  = \new_[12391]_  & \new_[12386]_ ;
  assign \new_[12395]_  = ~A169 & ~A170;
  assign \new_[12398]_  = A200 & ~A168;
  assign \new_[12399]_  = \new_[12398]_  & \new_[12395]_ ;
  assign \new_[12402]_  = ~A232 & A201;
  assign \new_[12406]_  = A268 & A236;
  assign \new_[12407]_  = A233 & \new_[12406]_ ;
  assign \new_[12408]_  = \new_[12407]_  & \new_[12402]_ ;
  assign \new_[12411]_  = ~A169 & ~A170;
  assign \new_[12414]_  = A200 & ~A168;
  assign \new_[12415]_  = \new_[12414]_  & \new_[12411]_ ;
  assign \new_[12418]_  = A232 & A201;
  assign \new_[12422]_  = A268 & A236;
  assign \new_[12423]_  = ~A233 & \new_[12422]_ ;
  assign \new_[12424]_  = \new_[12423]_  & \new_[12418]_ ;
  assign \new_[12427]_  = ~A169 & ~A170;
  assign \new_[12430]_  = ~A199 & ~A168;
  assign \new_[12431]_  = \new_[12430]_  & \new_[12427]_ ;
  assign \new_[12434]_  = A203 & A200;
  assign \new_[12438]_  = A267 & A265;
  assign \new_[12439]_  = A235 & \new_[12438]_ ;
  assign \new_[12440]_  = \new_[12439]_  & \new_[12434]_ ;
  assign \new_[12443]_  = ~A169 & ~A170;
  assign \new_[12446]_  = ~A199 & ~A168;
  assign \new_[12447]_  = \new_[12446]_  & \new_[12443]_ ;
  assign \new_[12450]_  = A203 & A200;
  assign \new_[12454]_  = A267 & A266;
  assign \new_[12455]_  = A235 & \new_[12454]_ ;
  assign \new_[12456]_  = \new_[12455]_  & \new_[12450]_ ;
  assign \new_[12459]_  = ~A169 & ~A170;
  assign \new_[12462]_  = ~A199 & ~A168;
  assign \new_[12463]_  = \new_[12462]_  & \new_[12459]_ ;
  assign \new_[12466]_  = A203 & A200;
  assign \new_[12470]_  = A268 & A234;
  assign \new_[12471]_  = A232 & \new_[12470]_ ;
  assign \new_[12472]_  = \new_[12471]_  & \new_[12466]_ ;
  assign \new_[12475]_  = ~A169 & ~A170;
  assign \new_[12478]_  = ~A199 & ~A168;
  assign \new_[12479]_  = \new_[12478]_  & \new_[12475]_ ;
  assign \new_[12482]_  = A203 & A200;
  assign \new_[12486]_  = A268 & A234;
  assign \new_[12487]_  = A233 & \new_[12486]_ ;
  assign \new_[12488]_  = \new_[12487]_  & \new_[12482]_ ;
  assign \new_[12491]_  = ~A169 & ~A170;
  assign \new_[12494]_  = A199 & ~A168;
  assign \new_[12495]_  = \new_[12494]_  & \new_[12491]_ ;
  assign \new_[12498]_  = A203 & ~A200;
  assign \new_[12502]_  = A267 & A265;
  assign \new_[12503]_  = A235 & \new_[12502]_ ;
  assign \new_[12504]_  = \new_[12503]_  & \new_[12498]_ ;
  assign \new_[12507]_  = ~A169 & ~A170;
  assign \new_[12510]_  = A199 & ~A168;
  assign \new_[12511]_  = \new_[12510]_  & \new_[12507]_ ;
  assign \new_[12514]_  = A203 & ~A200;
  assign \new_[12518]_  = A267 & A266;
  assign \new_[12519]_  = A235 & \new_[12518]_ ;
  assign \new_[12520]_  = \new_[12519]_  & \new_[12514]_ ;
  assign \new_[12523]_  = ~A169 & ~A170;
  assign \new_[12526]_  = A199 & ~A168;
  assign \new_[12527]_  = \new_[12526]_  & \new_[12523]_ ;
  assign \new_[12530]_  = A203 & ~A200;
  assign \new_[12534]_  = A268 & A234;
  assign \new_[12535]_  = A232 & \new_[12534]_ ;
  assign \new_[12536]_  = \new_[12535]_  & \new_[12530]_ ;
  assign \new_[12539]_  = ~A169 & ~A170;
  assign \new_[12542]_  = A199 & ~A168;
  assign \new_[12543]_  = \new_[12542]_  & \new_[12539]_ ;
  assign \new_[12546]_  = A203 & ~A200;
  assign \new_[12550]_  = A268 & A234;
  assign \new_[12551]_  = A233 & \new_[12550]_ ;
  assign \new_[12552]_  = \new_[12551]_  & \new_[12546]_ ;
  assign \new_[12555]_  = A166 & A168;
  assign \new_[12559]_  = ~A203 & ~A202;
  assign \new_[12560]_  = ~A201 & \new_[12559]_ ;
  assign \new_[12561]_  = \new_[12560]_  & \new_[12555]_ ;
  assign \new_[12564]_  = A298 & A235;
  assign \new_[12568]_  = ~A301 & ~A300;
  assign \new_[12569]_  = A299 & \new_[12568]_ ;
  assign \new_[12570]_  = \new_[12569]_  & \new_[12564]_ ;
  assign \new_[12573]_  = A166 & A168;
  assign \new_[12577]_  = ~A203 & ~A202;
  assign \new_[12578]_  = ~A201 & \new_[12577]_ ;
  assign \new_[12579]_  = \new_[12578]_  & \new_[12573]_ ;
  assign \new_[12582]_  = A234 & A232;
  assign \new_[12586]_  = ~A302 & ~A301;
  assign \new_[12587]_  = ~A300 & \new_[12586]_ ;
  assign \new_[12588]_  = \new_[12587]_  & \new_[12582]_ ;
  assign \new_[12591]_  = A166 & A168;
  assign \new_[12595]_  = ~A203 & ~A202;
  assign \new_[12596]_  = ~A201 & \new_[12595]_ ;
  assign \new_[12597]_  = \new_[12596]_  & \new_[12591]_ ;
  assign \new_[12600]_  = A234 & A232;
  assign \new_[12604]_  = ~A301 & ~A299;
  assign \new_[12605]_  = ~A298 & \new_[12604]_ ;
  assign \new_[12606]_  = \new_[12605]_  & \new_[12600]_ ;
  assign \new_[12609]_  = A166 & A168;
  assign \new_[12613]_  = ~A203 & ~A202;
  assign \new_[12614]_  = ~A201 & \new_[12613]_ ;
  assign \new_[12615]_  = \new_[12614]_  & \new_[12609]_ ;
  assign \new_[12618]_  = A234 & A232;
  assign \new_[12622]_  = A269 & A266;
  assign \new_[12623]_  = ~A265 & \new_[12622]_ ;
  assign \new_[12624]_  = \new_[12623]_  & \new_[12618]_ ;
  assign \new_[12627]_  = A166 & A168;
  assign \new_[12631]_  = ~A203 & ~A202;
  assign \new_[12632]_  = ~A201 & \new_[12631]_ ;
  assign \new_[12633]_  = \new_[12632]_  & \new_[12627]_ ;
  assign \new_[12636]_  = A234 & A232;
  assign \new_[12640]_  = A269 & ~A266;
  assign \new_[12641]_  = A265 & \new_[12640]_ ;
  assign \new_[12642]_  = \new_[12641]_  & \new_[12636]_ ;
  assign \new_[12645]_  = A166 & A168;
  assign \new_[12649]_  = ~A203 & ~A202;
  assign \new_[12650]_  = ~A201 & \new_[12649]_ ;
  assign \new_[12651]_  = \new_[12650]_  & \new_[12645]_ ;
  assign \new_[12654]_  = A234 & A233;
  assign \new_[12658]_  = ~A302 & ~A301;
  assign \new_[12659]_  = ~A300 & \new_[12658]_ ;
  assign \new_[12660]_  = \new_[12659]_  & \new_[12654]_ ;
  assign \new_[12663]_  = A166 & A168;
  assign \new_[12667]_  = ~A203 & ~A202;
  assign \new_[12668]_  = ~A201 & \new_[12667]_ ;
  assign \new_[12669]_  = \new_[12668]_  & \new_[12663]_ ;
  assign \new_[12672]_  = A234 & A233;
  assign \new_[12676]_  = ~A301 & ~A299;
  assign \new_[12677]_  = ~A298 & \new_[12676]_ ;
  assign \new_[12678]_  = \new_[12677]_  & \new_[12672]_ ;
  assign \new_[12681]_  = A166 & A168;
  assign \new_[12685]_  = ~A203 & ~A202;
  assign \new_[12686]_  = ~A201 & \new_[12685]_ ;
  assign \new_[12687]_  = \new_[12686]_  & \new_[12681]_ ;
  assign \new_[12690]_  = A234 & A233;
  assign \new_[12694]_  = A269 & A266;
  assign \new_[12695]_  = ~A265 & \new_[12694]_ ;
  assign \new_[12696]_  = \new_[12695]_  & \new_[12690]_ ;
  assign \new_[12699]_  = A166 & A168;
  assign \new_[12703]_  = ~A203 & ~A202;
  assign \new_[12704]_  = ~A201 & \new_[12703]_ ;
  assign \new_[12705]_  = \new_[12704]_  & \new_[12699]_ ;
  assign \new_[12708]_  = A234 & A233;
  assign \new_[12712]_  = A269 & ~A266;
  assign \new_[12713]_  = A265 & \new_[12712]_ ;
  assign \new_[12714]_  = \new_[12713]_  & \new_[12708]_ ;
  assign \new_[12717]_  = A166 & A168;
  assign \new_[12721]_  = ~A203 & ~A202;
  assign \new_[12722]_  = ~A201 & \new_[12721]_ ;
  assign \new_[12723]_  = \new_[12722]_  & \new_[12717]_ ;
  assign \new_[12726]_  = A233 & ~A232;
  assign \new_[12730]_  = A267 & A265;
  assign \new_[12731]_  = A236 & \new_[12730]_ ;
  assign \new_[12732]_  = \new_[12731]_  & \new_[12726]_ ;
  assign \new_[12735]_  = A166 & A168;
  assign \new_[12739]_  = ~A203 & ~A202;
  assign \new_[12740]_  = ~A201 & \new_[12739]_ ;
  assign \new_[12741]_  = \new_[12740]_  & \new_[12735]_ ;
  assign \new_[12744]_  = A233 & ~A232;
  assign \new_[12748]_  = A267 & A266;
  assign \new_[12749]_  = A236 & \new_[12748]_ ;
  assign \new_[12750]_  = \new_[12749]_  & \new_[12744]_ ;
  assign \new_[12753]_  = A166 & A168;
  assign \new_[12757]_  = ~A203 & ~A202;
  assign \new_[12758]_  = ~A201 & \new_[12757]_ ;
  assign \new_[12759]_  = \new_[12758]_  & \new_[12753]_ ;
  assign \new_[12762]_  = ~A233 & A232;
  assign \new_[12766]_  = A267 & A265;
  assign \new_[12767]_  = A236 & \new_[12766]_ ;
  assign \new_[12768]_  = \new_[12767]_  & \new_[12762]_ ;
  assign \new_[12771]_  = A166 & A168;
  assign \new_[12775]_  = ~A203 & ~A202;
  assign \new_[12776]_  = ~A201 & \new_[12775]_ ;
  assign \new_[12777]_  = \new_[12776]_  & \new_[12771]_ ;
  assign \new_[12780]_  = ~A233 & A232;
  assign \new_[12784]_  = A267 & A266;
  assign \new_[12785]_  = A236 & \new_[12784]_ ;
  assign \new_[12786]_  = \new_[12785]_  & \new_[12780]_ ;
  assign \new_[12789]_  = A166 & A168;
  assign \new_[12793]_  = ~A201 & A200;
  assign \new_[12794]_  = A199 & \new_[12793]_ ;
  assign \new_[12795]_  = \new_[12794]_  & \new_[12789]_ ;
  assign \new_[12798]_  = A235 & ~A202;
  assign \new_[12802]_  = ~A302 & ~A301;
  assign \new_[12803]_  = ~A300 & \new_[12802]_ ;
  assign \new_[12804]_  = \new_[12803]_  & \new_[12798]_ ;
  assign \new_[12807]_  = A166 & A168;
  assign \new_[12811]_  = ~A201 & A200;
  assign \new_[12812]_  = A199 & \new_[12811]_ ;
  assign \new_[12813]_  = \new_[12812]_  & \new_[12807]_ ;
  assign \new_[12816]_  = A235 & ~A202;
  assign \new_[12820]_  = ~A301 & ~A299;
  assign \new_[12821]_  = ~A298 & \new_[12820]_ ;
  assign \new_[12822]_  = \new_[12821]_  & \new_[12816]_ ;
  assign \new_[12825]_  = A166 & A168;
  assign \new_[12829]_  = ~A201 & A200;
  assign \new_[12830]_  = A199 & \new_[12829]_ ;
  assign \new_[12831]_  = \new_[12830]_  & \new_[12825]_ ;
  assign \new_[12834]_  = A235 & ~A202;
  assign \new_[12838]_  = A269 & A266;
  assign \new_[12839]_  = ~A265 & \new_[12838]_ ;
  assign \new_[12840]_  = \new_[12839]_  & \new_[12834]_ ;
  assign \new_[12843]_  = A166 & A168;
  assign \new_[12847]_  = ~A201 & A200;
  assign \new_[12848]_  = A199 & \new_[12847]_ ;
  assign \new_[12849]_  = \new_[12848]_  & \new_[12843]_ ;
  assign \new_[12852]_  = A235 & ~A202;
  assign \new_[12856]_  = A269 & ~A266;
  assign \new_[12857]_  = A265 & \new_[12856]_ ;
  assign \new_[12858]_  = \new_[12857]_  & \new_[12852]_ ;
  assign \new_[12861]_  = A166 & A168;
  assign \new_[12865]_  = ~A201 & A200;
  assign \new_[12866]_  = A199 & \new_[12865]_ ;
  assign \new_[12867]_  = \new_[12866]_  & \new_[12861]_ ;
  assign \new_[12870]_  = A232 & ~A202;
  assign \new_[12874]_  = A267 & A265;
  assign \new_[12875]_  = A234 & \new_[12874]_ ;
  assign \new_[12876]_  = \new_[12875]_  & \new_[12870]_ ;
  assign \new_[12879]_  = A166 & A168;
  assign \new_[12883]_  = ~A201 & A200;
  assign \new_[12884]_  = A199 & \new_[12883]_ ;
  assign \new_[12885]_  = \new_[12884]_  & \new_[12879]_ ;
  assign \new_[12888]_  = A232 & ~A202;
  assign \new_[12892]_  = A267 & A266;
  assign \new_[12893]_  = A234 & \new_[12892]_ ;
  assign \new_[12894]_  = \new_[12893]_  & \new_[12888]_ ;
  assign \new_[12897]_  = A166 & A168;
  assign \new_[12901]_  = ~A201 & A200;
  assign \new_[12902]_  = A199 & \new_[12901]_ ;
  assign \new_[12903]_  = \new_[12902]_  & \new_[12897]_ ;
  assign \new_[12906]_  = A233 & ~A202;
  assign \new_[12910]_  = A267 & A265;
  assign \new_[12911]_  = A234 & \new_[12910]_ ;
  assign \new_[12912]_  = \new_[12911]_  & \new_[12906]_ ;
  assign \new_[12915]_  = A166 & A168;
  assign \new_[12919]_  = ~A201 & A200;
  assign \new_[12920]_  = A199 & \new_[12919]_ ;
  assign \new_[12921]_  = \new_[12920]_  & \new_[12915]_ ;
  assign \new_[12924]_  = A233 & ~A202;
  assign \new_[12928]_  = A267 & A266;
  assign \new_[12929]_  = A234 & \new_[12928]_ ;
  assign \new_[12930]_  = \new_[12929]_  & \new_[12924]_ ;
  assign \new_[12933]_  = A166 & A168;
  assign \new_[12937]_  = ~A201 & A200;
  assign \new_[12938]_  = A199 & \new_[12937]_ ;
  assign \new_[12939]_  = \new_[12938]_  & \new_[12933]_ ;
  assign \new_[12942]_  = ~A232 & ~A202;
  assign \new_[12946]_  = A268 & A236;
  assign \new_[12947]_  = A233 & \new_[12946]_ ;
  assign \new_[12948]_  = \new_[12947]_  & \new_[12942]_ ;
  assign \new_[12951]_  = A166 & A168;
  assign \new_[12955]_  = ~A201 & A200;
  assign \new_[12956]_  = A199 & \new_[12955]_ ;
  assign \new_[12957]_  = \new_[12956]_  & \new_[12951]_ ;
  assign \new_[12960]_  = A232 & ~A202;
  assign \new_[12964]_  = A268 & A236;
  assign \new_[12965]_  = ~A233 & \new_[12964]_ ;
  assign \new_[12966]_  = \new_[12965]_  & \new_[12960]_ ;
  assign \new_[12969]_  = A166 & A168;
  assign \new_[12973]_  = ~A202 & ~A200;
  assign \new_[12974]_  = ~A199 & \new_[12973]_ ;
  assign \new_[12975]_  = \new_[12974]_  & \new_[12969]_ ;
  assign \new_[12978]_  = A298 & A235;
  assign \new_[12982]_  = ~A301 & ~A300;
  assign \new_[12983]_  = A299 & \new_[12982]_ ;
  assign \new_[12984]_  = \new_[12983]_  & \new_[12978]_ ;
  assign \new_[12987]_  = A166 & A168;
  assign \new_[12991]_  = ~A202 & ~A200;
  assign \new_[12992]_  = ~A199 & \new_[12991]_ ;
  assign \new_[12993]_  = \new_[12992]_  & \new_[12987]_ ;
  assign \new_[12996]_  = A234 & A232;
  assign \new_[13000]_  = ~A302 & ~A301;
  assign \new_[13001]_  = ~A300 & \new_[13000]_ ;
  assign \new_[13002]_  = \new_[13001]_  & \new_[12996]_ ;
  assign \new_[13005]_  = A166 & A168;
  assign \new_[13009]_  = ~A202 & ~A200;
  assign \new_[13010]_  = ~A199 & \new_[13009]_ ;
  assign \new_[13011]_  = \new_[13010]_  & \new_[13005]_ ;
  assign \new_[13014]_  = A234 & A232;
  assign \new_[13018]_  = ~A301 & ~A299;
  assign \new_[13019]_  = ~A298 & \new_[13018]_ ;
  assign \new_[13020]_  = \new_[13019]_  & \new_[13014]_ ;
  assign \new_[13023]_  = A166 & A168;
  assign \new_[13027]_  = ~A202 & ~A200;
  assign \new_[13028]_  = ~A199 & \new_[13027]_ ;
  assign \new_[13029]_  = \new_[13028]_  & \new_[13023]_ ;
  assign \new_[13032]_  = A234 & A232;
  assign \new_[13036]_  = A269 & A266;
  assign \new_[13037]_  = ~A265 & \new_[13036]_ ;
  assign \new_[13038]_  = \new_[13037]_  & \new_[13032]_ ;
  assign \new_[13041]_  = A166 & A168;
  assign \new_[13045]_  = ~A202 & ~A200;
  assign \new_[13046]_  = ~A199 & \new_[13045]_ ;
  assign \new_[13047]_  = \new_[13046]_  & \new_[13041]_ ;
  assign \new_[13050]_  = A234 & A232;
  assign \new_[13054]_  = A269 & ~A266;
  assign \new_[13055]_  = A265 & \new_[13054]_ ;
  assign \new_[13056]_  = \new_[13055]_  & \new_[13050]_ ;
  assign \new_[13059]_  = A166 & A168;
  assign \new_[13063]_  = ~A202 & ~A200;
  assign \new_[13064]_  = ~A199 & \new_[13063]_ ;
  assign \new_[13065]_  = \new_[13064]_  & \new_[13059]_ ;
  assign \new_[13068]_  = A234 & A233;
  assign \new_[13072]_  = ~A302 & ~A301;
  assign \new_[13073]_  = ~A300 & \new_[13072]_ ;
  assign \new_[13074]_  = \new_[13073]_  & \new_[13068]_ ;
  assign \new_[13077]_  = A166 & A168;
  assign \new_[13081]_  = ~A202 & ~A200;
  assign \new_[13082]_  = ~A199 & \new_[13081]_ ;
  assign \new_[13083]_  = \new_[13082]_  & \new_[13077]_ ;
  assign \new_[13086]_  = A234 & A233;
  assign \new_[13090]_  = ~A301 & ~A299;
  assign \new_[13091]_  = ~A298 & \new_[13090]_ ;
  assign \new_[13092]_  = \new_[13091]_  & \new_[13086]_ ;
  assign \new_[13095]_  = A166 & A168;
  assign \new_[13099]_  = ~A202 & ~A200;
  assign \new_[13100]_  = ~A199 & \new_[13099]_ ;
  assign \new_[13101]_  = \new_[13100]_  & \new_[13095]_ ;
  assign \new_[13104]_  = A234 & A233;
  assign \new_[13108]_  = A269 & A266;
  assign \new_[13109]_  = ~A265 & \new_[13108]_ ;
  assign \new_[13110]_  = \new_[13109]_  & \new_[13104]_ ;
  assign \new_[13113]_  = A166 & A168;
  assign \new_[13117]_  = ~A202 & ~A200;
  assign \new_[13118]_  = ~A199 & \new_[13117]_ ;
  assign \new_[13119]_  = \new_[13118]_  & \new_[13113]_ ;
  assign \new_[13122]_  = A234 & A233;
  assign \new_[13126]_  = A269 & ~A266;
  assign \new_[13127]_  = A265 & \new_[13126]_ ;
  assign \new_[13128]_  = \new_[13127]_  & \new_[13122]_ ;
  assign \new_[13131]_  = A166 & A168;
  assign \new_[13135]_  = ~A202 & ~A200;
  assign \new_[13136]_  = ~A199 & \new_[13135]_ ;
  assign \new_[13137]_  = \new_[13136]_  & \new_[13131]_ ;
  assign \new_[13140]_  = A233 & ~A232;
  assign \new_[13144]_  = A267 & A265;
  assign \new_[13145]_  = A236 & \new_[13144]_ ;
  assign \new_[13146]_  = \new_[13145]_  & \new_[13140]_ ;
  assign \new_[13149]_  = A166 & A168;
  assign \new_[13153]_  = ~A202 & ~A200;
  assign \new_[13154]_  = ~A199 & \new_[13153]_ ;
  assign \new_[13155]_  = \new_[13154]_  & \new_[13149]_ ;
  assign \new_[13158]_  = A233 & ~A232;
  assign \new_[13162]_  = A267 & A266;
  assign \new_[13163]_  = A236 & \new_[13162]_ ;
  assign \new_[13164]_  = \new_[13163]_  & \new_[13158]_ ;
  assign \new_[13167]_  = A166 & A168;
  assign \new_[13171]_  = ~A202 & ~A200;
  assign \new_[13172]_  = ~A199 & \new_[13171]_ ;
  assign \new_[13173]_  = \new_[13172]_  & \new_[13167]_ ;
  assign \new_[13176]_  = ~A233 & A232;
  assign \new_[13180]_  = A267 & A265;
  assign \new_[13181]_  = A236 & \new_[13180]_ ;
  assign \new_[13182]_  = \new_[13181]_  & \new_[13176]_ ;
  assign \new_[13185]_  = A166 & A168;
  assign \new_[13189]_  = ~A202 & ~A200;
  assign \new_[13190]_  = ~A199 & \new_[13189]_ ;
  assign \new_[13191]_  = \new_[13190]_  & \new_[13185]_ ;
  assign \new_[13194]_  = ~A233 & A232;
  assign \new_[13198]_  = A267 & A266;
  assign \new_[13199]_  = A236 & \new_[13198]_ ;
  assign \new_[13200]_  = \new_[13199]_  & \new_[13194]_ ;
  assign \new_[13203]_  = A167 & A168;
  assign \new_[13207]_  = ~A203 & ~A202;
  assign \new_[13208]_  = ~A201 & \new_[13207]_ ;
  assign \new_[13209]_  = \new_[13208]_  & \new_[13203]_ ;
  assign \new_[13212]_  = A298 & A235;
  assign \new_[13216]_  = ~A301 & ~A300;
  assign \new_[13217]_  = A299 & \new_[13216]_ ;
  assign \new_[13218]_  = \new_[13217]_  & \new_[13212]_ ;
  assign \new_[13221]_  = A167 & A168;
  assign \new_[13225]_  = ~A203 & ~A202;
  assign \new_[13226]_  = ~A201 & \new_[13225]_ ;
  assign \new_[13227]_  = \new_[13226]_  & \new_[13221]_ ;
  assign \new_[13230]_  = A234 & A232;
  assign \new_[13234]_  = ~A302 & ~A301;
  assign \new_[13235]_  = ~A300 & \new_[13234]_ ;
  assign \new_[13236]_  = \new_[13235]_  & \new_[13230]_ ;
  assign \new_[13239]_  = A167 & A168;
  assign \new_[13243]_  = ~A203 & ~A202;
  assign \new_[13244]_  = ~A201 & \new_[13243]_ ;
  assign \new_[13245]_  = \new_[13244]_  & \new_[13239]_ ;
  assign \new_[13248]_  = A234 & A232;
  assign \new_[13252]_  = ~A301 & ~A299;
  assign \new_[13253]_  = ~A298 & \new_[13252]_ ;
  assign \new_[13254]_  = \new_[13253]_  & \new_[13248]_ ;
  assign \new_[13257]_  = A167 & A168;
  assign \new_[13261]_  = ~A203 & ~A202;
  assign \new_[13262]_  = ~A201 & \new_[13261]_ ;
  assign \new_[13263]_  = \new_[13262]_  & \new_[13257]_ ;
  assign \new_[13266]_  = A234 & A232;
  assign \new_[13270]_  = A269 & A266;
  assign \new_[13271]_  = ~A265 & \new_[13270]_ ;
  assign \new_[13272]_  = \new_[13271]_  & \new_[13266]_ ;
  assign \new_[13275]_  = A167 & A168;
  assign \new_[13279]_  = ~A203 & ~A202;
  assign \new_[13280]_  = ~A201 & \new_[13279]_ ;
  assign \new_[13281]_  = \new_[13280]_  & \new_[13275]_ ;
  assign \new_[13284]_  = A234 & A232;
  assign \new_[13288]_  = A269 & ~A266;
  assign \new_[13289]_  = A265 & \new_[13288]_ ;
  assign \new_[13290]_  = \new_[13289]_  & \new_[13284]_ ;
  assign \new_[13293]_  = A167 & A168;
  assign \new_[13297]_  = ~A203 & ~A202;
  assign \new_[13298]_  = ~A201 & \new_[13297]_ ;
  assign \new_[13299]_  = \new_[13298]_  & \new_[13293]_ ;
  assign \new_[13302]_  = A234 & A233;
  assign \new_[13306]_  = ~A302 & ~A301;
  assign \new_[13307]_  = ~A300 & \new_[13306]_ ;
  assign \new_[13308]_  = \new_[13307]_  & \new_[13302]_ ;
  assign \new_[13311]_  = A167 & A168;
  assign \new_[13315]_  = ~A203 & ~A202;
  assign \new_[13316]_  = ~A201 & \new_[13315]_ ;
  assign \new_[13317]_  = \new_[13316]_  & \new_[13311]_ ;
  assign \new_[13320]_  = A234 & A233;
  assign \new_[13324]_  = ~A301 & ~A299;
  assign \new_[13325]_  = ~A298 & \new_[13324]_ ;
  assign \new_[13326]_  = \new_[13325]_  & \new_[13320]_ ;
  assign \new_[13329]_  = A167 & A168;
  assign \new_[13333]_  = ~A203 & ~A202;
  assign \new_[13334]_  = ~A201 & \new_[13333]_ ;
  assign \new_[13335]_  = \new_[13334]_  & \new_[13329]_ ;
  assign \new_[13338]_  = A234 & A233;
  assign \new_[13342]_  = A269 & A266;
  assign \new_[13343]_  = ~A265 & \new_[13342]_ ;
  assign \new_[13344]_  = \new_[13343]_  & \new_[13338]_ ;
  assign \new_[13347]_  = A167 & A168;
  assign \new_[13351]_  = ~A203 & ~A202;
  assign \new_[13352]_  = ~A201 & \new_[13351]_ ;
  assign \new_[13353]_  = \new_[13352]_  & \new_[13347]_ ;
  assign \new_[13356]_  = A234 & A233;
  assign \new_[13360]_  = A269 & ~A266;
  assign \new_[13361]_  = A265 & \new_[13360]_ ;
  assign \new_[13362]_  = \new_[13361]_  & \new_[13356]_ ;
  assign \new_[13365]_  = A167 & A168;
  assign \new_[13369]_  = ~A203 & ~A202;
  assign \new_[13370]_  = ~A201 & \new_[13369]_ ;
  assign \new_[13371]_  = \new_[13370]_  & \new_[13365]_ ;
  assign \new_[13374]_  = A233 & ~A232;
  assign \new_[13378]_  = A267 & A265;
  assign \new_[13379]_  = A236 & \new_[13378]_ ;
  assign \new_[13380]_  = \new_[13379]_  & \new_[13374]_ ;
  assign \new_[13383]_  = A167 & A168;
  assign \new_[13387]_  = ~A203 & ~A202;
  assign \new_[13388]_  = ~A201 & \new_[13387]_ ;
  assign \new_[13389]_  = \new_[13388]_  & \new_[13383]_ ;
  assign \new_[13392]_  = A233 & ~A232;
  assign \new_[13396]_  = A267 & A266;
  assign \new_[13397]_  = A236 & \new_[13396]_ ;
  assign \new_[13398]_  = \new_[13397]_  & \new_[13392]_ ;
  assign \new_[13401]_  = A167 & A168;
  assign \new_[13405]_  = ~A203 & ~A202;
  assign \new_[13406]_  = ~A201 & \new_[13405]_ ;
  assign \new_[13407]_  = \new_[13406]_  & \new_[13401]_ ;
  assign \new_[13410]_  = ~A233 & A232;
  assign \new_[13414]_  = A267 & A265;
  assign \new_[13415]_  = A236 & \new_[13414]_ ;
  assign \new_[13416]_  = \new_[13415]_  & \new_[13410]_ ;
  assign \new_[13419]_  = A167 & A168;
  assign \new_[13423]_  = ~A203 & ~A202;
  assign \new_[13424]_  = ~A201 & \new_[13423]_ ;
  assign \new_[13425]_  = \new_[13424]_  & \new_[13419]_ ;
  assign \new_[13428]_  = ~A233 & A232;
  assign \new_[13432]_  = A267 & A266;
  assign \new_[13433]_  = A236 & \new_[13432]_ ;
  assign \new_[13434]_  = \new_[13433]_  & \new_[13428]_ ;
  assign \new_[13437]_  = A167 & A168;
  assign \new_[13441]_  = ~A201 & A200;
  assign \new_[13442]_  = A199 & \new_[13441]_ ;
  assign \new_[13443]_  = \new_[13442]_  & \new_[13437]_ ;
  assign \new_[13446]_  = A235 & ~A202;
  assign \new_[13450]_  = ~A302 & ~A301;
  assign \new_[13451]_  = ~A300 & \new_[13450]_ ;
  assign \new_[13452]_  = \new_[13451]_  & \new_[13446]_ ;
  assign \new_[13455]_  = A167 & A168;
  assign \new_[13459]_  = ~A201 & A200;
  assign \new_[13460]_  = A199 & \new_[13459]_ ;
  assign \new_[13461]_  = \new_[13460]_  & \new_[13455]_ ;
  assign \new_[13464]_  = A235 & ~A202;
  assign \new_[13468]_  = ~A301 & ~A299;
  assign \new_[13469]_  = ~A298 & \new_[13468]_ ;
  assign \new_[13470]_  = \new_[13469]_  & \new_[13464]_ ;
  assign \new_[13473]_  = A167 & A168;
  assign \new_[13477]_  = ~A201 & A200;
  assign \new_[13478]_  = A199 & \new_[13477]_ ;
  assign \new_[13479]_  = \new_[13478]_  & \new_[13473]_ ;
  assign \new_[13482]_  = A235 & ~A202;
  assign \new_[13486]_  = A269 & A266;
  assign \new_[13487]_  = ~A265 & \new_[13486]_ ;
  assign \new_[13488]_  = \new_[13487]_  & \new_[13482]_ ;
  assign \new_[13491]_  = A167 & A168;
  assign \new_[13495]_  = ~A201 & A200;
  assign \new_[13496]_  = A199 & \new_[13495]_ ;
  assign \new_[13497]_  = \new_[13496]_  & \new_[13491]_ ;
  assign \new_[13500]_  = A235 & ~A202;
  assign \new_[13504]_  = A269 & ~A266;
  assign \new_[13505]_  = A265 & \new_[13504]_ ;
  assign \new_[13506]_  = \new_[13505]_  & \new_[13500]_ ;
  assign \new_[13509]_  = A167 & A168;
  assign \new_[13513]_  = ~A201 & A200;
  assign \new_[13514]_  = A199 & \new_[13513]_ ;
  assign \new_[13515]_  = \new_[13514]_  & \new_[13509]_ ;
  assign \new_[13518]_  = A232 & ~A202;
  assign \new_[13522]_  = A267 & A265;
  assign \new_[13523]_  = A234 & \new_[13522]_ ;
  assign \new_[13524]_  = \new_[13523]_  & \new_[13518]_ ;
  assign \new_[13527]_  = A167 & A168;
  assign \new_[13531]_  = ~A201 & A200;
  assign \new_[13532]_  = A199 & \new_[13531]_ ;
  assign \new_[13533]_  = \new_[13532]_  & \new_[13527]_ ;
  assign \new_[13536]_  = A232 & ~A202;
  assign \new_[13540]_  = A267 & A266;
  assign \new_[13541]_  = A234 & \new_[13540]_ ;
  assign \new_[13542]_  = \new_[13541]_  & \new_[13536]_ ;
  assign \new_[13545]_  = A167 & A168;
  assign \new_[13549]_  = ~A201 & A200;
  assign \new_[13550]_  = A199 & \new_[13549]_ ;
  assign \new_[13551]_  = \new_[13550]_  & \new_[13545]_ ;
  assign \new_[13554]_  = A233 & ~A202;
  assign \new_[13558]_  = A267 & A265;
  assign \new_[13559]_  = A234 & \new_[13558]_ ;
  assign \new_[13560]_  = \new_[13559]_  & \new_[13554]_ ;
  assign \new_[13563]_  = A167 & A168;
  assign \new_[13567]_  = ~A201 & A200;
  assign \new_[13568]_  = A199 & \new_[13567]_ ;
  assign \new_[13569]_  = \new_[13568]_  & \new_[13563]_ ;
  assign \new_[13572]_  = A233 & ~A202;
  assign \new_[13576]_  = A267 & A266;
  assign \new_[13577]_  = A234 & \new_[13576]_ ;
  assign \new_[13578]_  = \new_[13577]_  & \new_[13572]_ ;
  assign \new_[13581]_  = A167 & A168;
  assign \new_[13585]_  = ~A201 & A200;
  assign \new_[13586]_  = A199 & \new_[13585]_ ;
  assign \new_[13587]_  = \new_[13586]_  & \new_[13581]_ ;
  assign \new_[13590]_  = ~A232 & ~A202;
  assign \new_[13594]_  = A268 & A236;
  assign \new_[13595]_  = A233 & \new_[13594]_ ;
  assign \new_[13596]_  = \new_[13595]_  & \new_[13590]_ ;
  assign \new_[13599]_  = A167 & A168;
  assign \new_[13603]_  = ~A201 & A200;
  assign \new_[13604]_  = A199 & \new_[13603]_ ;
  assign \new_[13605]_  = \new_[13604]_  & \new_[13599]_ ;
  assign \new_[13608]_  = A232 & ~A202;
  assign \new_[13612]_  = A268 & A236;
  assign \new_[13613]_  = ~A233 & \new_[13612]_ ;
  assign \new_[13614]_  = \new_[13613]_  & \new_[13608]_ ;
  assign \new_[13617]_  = A167 & A168;
  assign \new_[13621]_  = ~A202 & ~A200;
  assign \new_[13622]_  = ~A199 & \new_[13621]_ ;
  assign \new_[13623]_  = \new_[13622]_  & \new_[13617]_ ;
  assign \new_[13626]_  = A298 & A235;
  assign \new_[13630]_  = ~A301 & ~A300;
  assign \new_[13631]_  = A299 & \new_[13630]_ ;
  assign \new_[13632]_  = \new_[13631]_  & \new_[13626]_ ;
  assign \new_[13635]_  = A167 & A168;
  assign \new_[13639]_  = ~A202 & ~A200;
  assign \new_[13640]_  = ~A199 & \new_[13639]_ ;
  assign \new_[13641]_  = \new_[13640]_  & \new_[13635]_ ;
  assign \new_[13644]_  = A234 & A232;
  assign \new_[13648]_  = ~A302 & ~A301;
  assign \new_[13649]_  = ~A300 & \new_[13648]_ ;
  assign \new_[13650]_  = \new_[13649]_  & \new_[13644]_ ;
  assign \new_[13653]_  = A167 & A168;
  assign \new_[13657]_  = ~A202 & ~A200;
  assign \new_[13658]_  = ~A199 & \new_[13657]_ ;
  assign \new_[13659]_  = \new_[13658]_  & \new_[13653]_ ;
  assign \new_[13662]_  = A234 & A232;
  assign \new_[13666]_  = ~A301 & ~A299;
  assign \new_[13667]_  = ~A298 & \new_[13666]_ ;
  assign \new_[13668]_  = \new_[13667]_  & \new_[13662]_ ;
  assign \new_[13671]_  = A167 & A168;
  assign \new_[13675]_  = ~A202 & ~A200;
  assign \new_[13676]_  = ~A199 & \new_[13675]_ ;
  assign \new_[13677]_  = \new_[13676]_  & \new_[13671]_ ;
  assign \new_[13680]_  = A234 & A232;
  assign \new_[13684]_  = A269 & A266;
  assign \new_[13685]_  = ~A265 & \new_[13684]_ ;
  assign \new_[13686]_  = \new_[13685]_  & \new_[13680]_ ;
  assign \new_[13689]_  = A167 & A168;
  assign \new_[13693]_  = ~A202 & ~A200;
  assign \new_[13694]_  = ~A199 & \new_[13693]_ ;
  assign \new_[13695]_  = \new_[13694]_  & \new_[13689]_ ;
  assign \new_[13698]_  = A234 & A232;
  assign \new_[13702]_  = A269 & ~A266;
  assign \new_[13703]_  = A265 & \new_[13702]_ ;
  assign \new_[13704]_  = \new_[13703]_  & \new_[13698]_ ;
  assign \new_[13707]_  = A167 & A168;
  assign \new_[13711]_  = ~A202 & ~A200;
  assign \new_[13712]_  = ~A199 & \new_[13711]_ ;
  assign \new_[13713]_  = \new_[13712]_  & \new_[13707]_ ;
  assign \new_[13716]_  = A234 & A233;
  assign \new_[13720]_  = ~A302 & ~A301;
  assign \new_[13721]_  = ~A300 & \new_[13720]_ ;
  assign \new_[13722]_  = \new_[13721]_  & \new_[13716]_ ;
  assign \new_[13725]_  = A167 & A168;
  assign \new_[13729]_  = ~A202 & ~A200;
  assign \new_[13730]_  = ~A199 & \new_[13729]_ ;
  assign \new_[13731]_  = \new_[13730]_  & \new_[13725]_ ;
  assign \new_[13734]_  = A234 & A233;
  assign \new_[13738]_  = ~A301 & ~A299;
  assign \new_[13739]_  = ~A298 & \new_[13738]_ ;
  assign \new_[13740]_  = \new_[13739]_  & \new_[13734]_ ;
  assign \new_[13743]_  = A167 & A168;
  assign \new_[13747]_  = ~A202 & ~A200;
  assign \new_[13748]_  = ~A199 & \new_[13747]_ ;
  assign \new_[13749]_  = \new_[13748]_  & \new_[13743]_ ;
  assign \new_[13752]_  = A234 & A233;
  assign \new_[13756]_  = A269 & A266;
  assign \new_[13757]_  = ~A265 & \new_[13756]_ ;
  assign \new_[13758]_  = \new_[13757]_  & \new_[13752]_ ;
  assign \new_[13761]_  = A167 & A168;
  assign \new_[13765]_  = ~A202 & ~A200;
  assign \new_[13766]_  = ~A199 & \new_[13765]_ ;
  assign \new_[13767]_  = \new_[13766]_  & \new_[13761]_ ;
  assign \new_[13770]_  = A234 & A233;
  assign \new_[13774]_  = A269 & ~A266;
  assign \new_[13775]_  = A265 & \new_[13774]_ ;
  assign \new_[13776]_  = \new_[13775]_  & \new_[13770]_ ;
  assign \new_[13779]_  = A167 & A168;
  assign \new_[13783]_  = ~A202 & ~A200;
  assign \new_[13784]_  = ~A199 & \new_[13783]_ ;
  assign \new_[13785]_  = \new_[13784]_  & \new_[13779]_ ;
  assign \new_[13788]_  = A233 & ~A232;
  assign \new_[13792]_  = A267 & A265;
  assign \new_[13793]_  = A236 & \new_[13792]_ ;
  assign \new_[13794]_  = \new_[13793]_  & \new_[13788]_ ;
  assign \new_[13797]_  = A167 & A168;
  assign \new_[13801]_  = ~A202 & ~A200;
  assign \new_[13802]_  = ~A199 & \new_[13801]_ ;
  assign \new_[13803]_  = \new_[13802]_  & \new_[13797]_ ;
  assign \new_[13806]_  = A233 & ~A232;
  assign \new_[13810]_  = A267 & A266;
  assign \new_[13811]_  = A236 & \new_[13810]_ ;
  assign \new_[13812]_  = \new_[13811]_  & \new_[13806]_ ;
  assign \new_[13815]_  = A167 & A168;
  assign \new_[13819]_  = ~A202 & ~A200;
  assign \new_[13820]_  = ~A199 & \new_[13819]_ ;
  assign \new_[13821]_  = \new_[13820]_  & \new_[13815]_ ;
  assign \new_[13824]_  = ~A233 & A232;
  assign \new_[13828]_  = A267 & A265;
  assign \new_[13829]_  = A236 & \new_[13828]_ ;
  assign \new_[13830]_  = \new_[13829]_  & \new_[13824]_ ;
  assign \new_[13833]_  = A167 & A168;
  assign \new_[13837]_  = ~A202 & ~A200;
  assign \new_[13838]_  = ~A199 & \new_[13837]_ ;
  assign \new_[13839]_  = \new_[13838]_  & \new_[13833]_ ;
  assign \new_[13842]_  = ~A233 & A232;
  assign \new_[13846]_  = A267 & A266;
  assign \new_[13847]_  = A236 & \new_[13846]_ ;
  assign \new_[13848]_  = \new_[13847]_  & \new_[13842]_ ;
  assign \new_[13851]_  = A167 & A170;
  assign \new_[13855]_  = ~A202 & ~A201;
  assign \new_[13856]_  = ~A166 & \new_[13855]_ ;
  assign \new_[13857]_  = \new_[13856]_  & \new_[13851]_ ;
  assign \new_[13860]_  = A235 & ~A203;
  assign \new_[13864]_  = ~A302 & ~A301;
  assign \new_[13865]_  = ~A300 & \new_[13864]_ ;
  assign \new_[13866]_  = \new_[13865]_  & \new_[13860]_ ;
  assign \new_[13869]_  = A167 & A170;
  assign \new_[13873]_  = ~A202 & ~A201;
  assign \new_[13874]_  = ~A166 & \new_[13873]_ ;
  assign \new_[13875]_  = \new_[13874]_  & \new_[13869]_ ;
  assign \new_[13878]_  = A235 & ~A203;
  assign \new_[13882]_  = ~A301 & ~A299;
  assign \new_[13883]_  = ~A298 & \new_[13882]_ ;
  assign \new_[13884]_  = \new_[13883]_  & \new_[13878]_ ;
  assign \new_[13887]_  = A167 & A170;
  assign \new_[13891]_  = ~A202 & ~A201;
  assign \new_[13892]_  = ~A166 & \new_[13891]_ ;
  assign \new_[13893]_  = \new_[13892]_  & \new_[13887]_ ;
  assign \new_[13896]_  = A235 & ~A203;
  assign \new_[13900]_  = A269 & A266;
  assign \new_[13901]_  = ~A265 & \new_[13900]_ ;
  assign \new_[13902]_  = \new_[13901]_  & \new_[13896]_ ;
  assign \new_[13905]_  = A167 & A170;
  assign \new_[13909]_  = ~A202 & ~A201;
  assign \new_[13910]_  = ~A166 & \new_[13909]_ ;
  assign \new_[13911]_  = \new_[13910]_  & \new_[13905]_ ;
  assign \new_[13914]_  = A235 & ~A203;
  assign \new_[13918]_  = A269 & ~A266;
  assign \new_[13919]_  = A265 & \new_[13918]_ ;
  assign \new_[13920]_  = \new_[13919]_  & \new_[13914]_ ;
  assign \new_[13923]_  = A167 & A170;
  assign \new_[13927]_  = ~A202 & ~A201;
  assign \new_[13928]_  = ~A166 & \new_[13927]_ ;
  assign \new_[13929]_  = \new_[13928]_  & \new_[13923]_ ;
  assign \new_[13932]_  = A232 & ~A203;
  assign \new_[13936]_  = A267 & A265;
  assign \new_[13937]_  = A234 & \new_[13936]_ ;
  assign \new_[13938]_  = \new_[13937]_  & \new_[13932]_ ;
  assign \new_[13941]_  = A167 & A170;
  assign \new_[13945]_  = ~A202 & ~A201;
  assign \new_[13946]_  = ~A166 & \new_[13945]_ ;
  assign \new_[13947]_  = \new_[13946]_  & \new_[13941]_ ;
  assign \new_[13950]_  = A232 & ~A203;
  assign \new_[13954]_  = A267 & A266;
  assign \new_[13955]_  = A234 & \new_[13954]_ ;
  assign \new_[13956]_  = \new_[13955]_  & \new_[13950]_ ;
  assign \new_[13959]_  = A167 & A170;
  assign \new_[13963]_  = ~A202 & ~A201;
  assign \new_[13964]_  = ~A166 & \new_[13963]_ ;
  assign \new_[13965]_  = \new_[13964]_  & \new_[13959]_ ;
  assign \new_[13968]_  = A233 & ~A203;
  assign \new_[13972]_  = A267 & A265;
  assign \new_[13973]_  = A234 & \new_[13972]_ ;
  assign \new_[13974]_  = \new_[13973]_  & \new_[13968]_ ;
  assign \new_[13977]_  = A167 & A170;
  assign \new_[13981]_  = ~A202 & ~A201;
  assign \new_[13982]_  = ~A166 & \new_[13981]_ ;
  assign \new_[13983]_  = \new_[13982]_  & \new_[13977]_ ;
  assign \new_[13986]_  = A233 & ~A203;
  assign \new_[13990]_  = A267 & A266;
  assign \new_[13991]_  = A234 & \new_[13990]_ ;
  assign \new_[13992]_  = \new_[13991]_  & \new_[13986]_ ;
  assign \new_[13995]_  = A167 & A170;
  assign \new_[13999]_  = ~A202 & ~A201;
  assign \new_[14000]_  = ~A166 & \new_[13999]_ ;
  assign \new_[14001]_  = \new_[14000]_  & \new_[13995]_ ;
  assign \new_[14004]_  = ~A232 & ~A203;
  assign \new_[14008]_  = A268 & A236;
  assign \new_[14009]_  = A233 & \new_[14008]_ ;
  assign \new_[14010]_  = \new_[14009]_  & \new_[14004]_ ;
  assign \new_[14013]_  = A167 & A170;
  assign \new_[14017]_  = ~A202 & ~A201;
  assign \new_[14018]_  = ~A166 & \new_[14017]_ ;
  assign \new_[14019]_  = \new_[14018]_  & \new_[14013]_ ;
  assign \new_[14022]_  = A232 & ~A203;
  assign \new_[14026]_  = A268 & A236;
  assign \new_[14027]_  = ~A233 & \new_[14026]_ ;
  assign \new_[14028]_  = \new_[14027]_  & \new_[14022]_ ;
  assign \new_[14031]_  = A167 & A170;
  assign \new_[14035]_  = A200 & A199;
  assign \new_[14036]_  = ~A166 & \new_[14035]_ ;
  assign \new_[14037]_  = \new_[14036]_  & \new_[14031]_ ;
  assign \new_[14040]_  = ~A202 & ~A201;
  assign \new_[14044]_  = A267 & A265;
  assign \new_[14045]_  = A235 & \new_[14044]_ ;
  assign \new_[14046]_  = \new_[14045]_  & \new_[14040]_ ;
  assign \new_[14049]_  = A167 & A170;
  assign \new_[14053]_  = A200 & A199;
  assign \new_[14054]_  = ~A166 & \new_[14053]_ ;
  assign \new_[14055]_  = \new_[14054]_  & \new_[14049]_ ;
  assign \new_[14058]_  = ~A202 & ~A201;
  assign \new_[14062]_  = A267 & A266;
  assign \new_[14063]_  = A235 & \new_[14062]_ ;
  assign \new_[14064]_  = \new_[14063]_  & \new_[14058]_ ;
  assign \new_[14067]_  = A167 & A170;
  assign \new_[14071]_  = A200 & A199;
  assign \new_[14072]_  = ~A166 & \new_[14071]_ ;
  assign \new_[14073]_  = \new_[14072]_  & \new_[14067]_ ;
  assign \new_[14076]_  = ~A202 & ~A201;
  assign \new_[14080]_  = A268 & A234;
  assign \new_[14081]_  = A232 & \new_[14080]_ ;
  assign \new_[14082]_  = \new_[14081]_  & \new_[14076]_ ;
  assign \new_[14085]_  = A167 & A170;
  assign \new_[14089]_  = A200 & A199;
  assign \new_[14090]_  = ~A166 & \new_[14089]_ ;
  assign \new_[14091]_  = \new_[14090]_  & \new_[14085]_ ;
  assign \new_[14094]_  = ~A202 & ~A201;
  assign \new_[14098]_  = A268 & A234;
  assign \new_[14099]_  = A233 & \new_[14098]_ ;
  assign \new_[14100]_  = \new_[14099]_  & \new_[14094]_ ;
  assign \new_[14103]_  = A167 & A170;
  assign \new_[14107]_  = ~A200 & ~A199;
  assign \new_[14108]_  = ~A166 & \new_[14107]_ ;
  assign \new_[14109]_  = \new_[14108]_  & \new_[14103]_ ;
  assign \new_[14112]_  = A235 & ~A202;
  assign \new_[14116]_  = ~A302 & ~A301;
  assign \new_[14117]_  = ~A300 & \new_[14116]_ ;
  assign \new_[14118]_  = \new_[14117]_  & \new_[14112]_ ;
  assign \new_[14121]_  = A167 & A170;
  assign \new_[14125]_  = ~A200 & ~A199;
  assign \new_[14126]_  = ~A166 & \new_[14125]_ ;
  assign \new_[14127]_  = \new_[14126]_  & \new_[14121]_ ;
  assign \new_[14130]_  = A235 & ~A202;
  assign \new_[14134]_  = ~A301 & ~A299;
  assign \new_[14135]_  = ~A298 & \new_[14134]_ ;
  assign \new_[14136]_  = \new_[14135]_  & \new_[14130]_ ;
  assign \new_[14139]_  = A167 & A170;
  assign \new_[14143]_  = ~A200 & ~A199;
  assign \new_[14144]_  = ~A166 & \new_[14143]_ ;
  assign \new_[14145]_  = \new_[14144]_  & \new_[14139]_ ;
  assign \new_[14148]_  = A235 & ~A202;
  assign \new_[14152]_  = A269 & A266;
  assign \new_[14153]_  = ~A265 & \new_[14152]_ ;
  assign \new_[14154]_  = \new_[14153]_  & \new_[14148]_ ;
  assign \new_[14157]_  = A167 & A170;
  assign \new_[14161]_  = ~A200 & ~A199;
  assign \new_[14162]_  = ~A166 & \new_[14161]_ ;
  assign \new_[14163]_  = \new_[14162]_  & \new_[14157]_ ;
  assign \new_[14166]_  = A235 & ~A202;
  assign \new_[14170]_  = A269 & ~A266;
  assign \new_[14171]_  = A265 & \new_[14170]_ ;
  assign \new_[14172]_  = \new_[14171]_  & \new_[14166]_ ;
  assign \new_[14175]_  = A167 & A170;
  assign \new_[14179]_  = ~A200 & ~A199;
  assign \new_[14180]_  = ~A166 & \new_[14179]_ ;
  assign \new_[14181]_  = \new_[14180]_  & \new_[14175]_ ;
  assign \new_[14184]_  = A232 & ~A202;
  assign \new_[14188]_  = A267 & A265;
  assign \new_[14189]_  = A234 & \new_[14188]_ ;
  assign \new_[14190]_  = \new_[14189]_  & \new_[14184]_ ;
  assign \new_[14193]_  = A167 & A170;
  assign \new_[14197]_  = ~A200 & ~A199;
  assign \new_[14198]_  = ~A166 & \new_[14197]_ ;
  assign \new_[14199]_  = \new_[14198]_  & \new_[14193]_ ;
  assign \new_[14202]_  = A232 & ~A202;
  assign \new_[14206]_  = A267 & A266;
  assign \new_[14207]_  = A234 & \new_[14206]_ ;
  assign \new_[14208]_  = \new_[14207]_  & \new_[14202]_ ;
  assign \new_[14211]_  = A167 & A170;
  assign \new_[14215]_  = ~A200 & ~A199;
  assign \new_[14216]_  = ~A166 & \new_[14215]_ ;
  assign \new_[14217]_  = \new_[14216]_  & \new_[14211]_ ;
  assign \new_[14220]_  = A233 & ~A202;
  assign \new_[14224]_  = A267 & A265;
  assign \new_[14225]_  = A234 & \new_[14224]_ ;
  assign \new_[14226]_  = \new_[14225]_  & \new_[14220]_ ;
  assign \new_[14229]_  = A167 & A170;
  assign \new_[14233]_  = ~A200 & ~A199;
  assign \new_[14234]_  = ~A166 & \new_[14233]_ ;
  assign \new_[14235]_  = \new_[14234]_  & \new_[14229]_ ;
  assign \new_[14238]_  = A233 & ~A202;
  assign \new_[14242]_  = A267 & A266;
  assign \new_[14243]_  = A234 & \new_[14242]_ ;
  assign \new_[14244]_  = \new_[14243]_  & \new_[14238]_ ;
  assign \new_[14247]_  = A167 & A170;
  assign \new_[14251]_  = ~A200 & ~A199;
  assign \new_[14252]_  = ~A166 & \new_[14251]_ ;
  assign \new_[14253]_  = \new_[14252]_  & \new_[14247]_ ;
  assign \new_[14256]_  = ~A232 & ~A202;
  assign \new_[14260]_  = A268 & A236;
  assign \new_[14261]_  = A233 & \new_[14260]_ ;
  assign \new_[14262]_  = \new_[14261]_  & \new_[14256]_ ;
  assign \new_[14265]_  = A167 & A170;
  assign \new_[14269]_  = ~A200 & ~A199;
  assign \new_[14270]_  = ~A166 & \new_[14269]_ ;
  assign \new_[14271]_  = \new_[14270]_  & \new_[14265]_ ;
  assign \new_[14274]_  = A232 & ~A202;
  assign \new_[14278]_  = A268 & A236;
  assign \new_[14279]_  = ~A233 & \new_[14278]_ ;
  assign \new_[14280]_  = \new_[14279]_  & \new_[14274]_ ;
  assign \new_[14283]_  = ~A167 & A170;
  assign \new_[14287]_  = ~A202 & ~A201;
  assign \new_[14288]_  = A166 & \new_[14287]_ ;
  assign \new_[14289]_  = \new_[14288]_  & \new_[14283]_ ;
  assign \new_[14292]_  = A235 & ~A203;
  assign \new_[14296]_  = ~A302 & ~A301;
  assign \new_[14297]_  = ~A300 & \new_[14296]_ ;
  assign \new_[14298]_  = \new_[14297]_  & \new_[14292]_ ;
  assign \new_[14301]_  = ~A167 & A170;
  assign \new_[14305]_  = ~A202 & ~A201;
  assign \new_[14306]_  = A166 & \new_[14305]_ ;
  assign \new_[14307]_  = \new_[14306]_  & \new_[14301]_ ;
  assign \new_[14310]_  = A235 & ~A203;
  assign \new_[14314]_  = ~A301 & ~A299;
  assign \new_[14315]_  = ~A298 & \new_[14314]_ ;
  assign \new_[14316]_  = \new_[14315]_  & \new_[14310]_ ;
  assign \new_[14319]_  = ~A167 & A170;
  assign \new_[14323]_  = ~A202 & ~A201;
  assign \new_[14324]_  = A166 & \new_[14323]_ ;
  assign \new_[14325]_  = \new_[14324]_  & \new_[14319]_ ;
  assign \new_[14328]_  = A235 & ~A203;
  assign \new_[14332]_  = A269 & A266;
  assign \new_[14333]_  = ~A265 & \new_[14332]_ ;
  assign \new_[14334]_  = \new_[14333]_  & \new_[14328]_ ;
  assign \new_[14337]_  = ~A167 & A170;
  assign \new_[14341]_  = ~A202 & ~A201;
  assign \new_[14342]_  = A166 & \new_[14341]_ ;
  assign \new_[14343]_  = \new_[14342]_  & \new_[14337]_ ;
  assign \new_[14346]_  = A235 & ~A203;
  assign \new_[14350]_  = A269 & ~A266;
  assign \new_[14351]_  = A265 & \new_[14350]_ ;
  assign \new_[14352]_  = \new_[14351]_  & \new_[14346]_ ;
  assign \new_[14355]_  = ~A167 & A170;
  assign \new_[14359]_  = ~A202 & ~A201;
  assign \new_[14360]_  = A166 & \new_[14359]_ ;
  assign \new_[14361]_  = \new_[14360]_  & \new_[14355]_ ;
  assign \new_[14364]_  = A232 & ~A203;
  assign \new_[14368]_  = A267 & A265;
  assign \new_[14369]_  = A234 & \new_[14368]_ ;
  assign \new_[14370]_  = \new_[14369]_  & \new_[14364]_ ;
  assign \new_[14373]_  = ~A167 & A170;
  assign \new_[14377]_  = ~A202 & ~A201;
  assign \new_[14378]_  = A166 & \new_[14377]_ ;
  assign \new_[14379]_  = \new_[14378]_  & \new_[14373]_ ;
  assign \new_[14382]_  = A232 & ~A203;
  assign \new_[14386]_  = A267 & A266;
  assign \new_[14387]_  = A234 & \new_[14386]_ ;
  assign \new_[14388]_  = \new_[14387]_  & \new_[14382]_ ;
  assign \new_[14391]_  = ~A167 & A170;
  assign \new_[14395]_  = ~A202 & ~A201;
  assign \new_[14396]_  = A166 & \new_[14395]_ ;
  assign \new_[14397]_  = \new_[14396]_  & \new_[14391]_ ;
  assign \new_[14400]_  = A233 & ~A203;
  assign \new_[14404]_  = A267 & A265;
  assign \new_[14405]_  = A234 & \new_[14404]_ ;
  assign \new_[14406]_  = \new_[14405]_  & \new_[14400]_ ;
  assign \new_[14409]_  = ~A167 & A170;
  assign \new_[14413]_  = ~A202 & ~A201;
  assign \new_[14414]_  = A166 & \new_[14413]_ ;
  assign \new_[14415]_  = \new_[14414]_  & \new_[14409]_ ;
  assign \new_[14418]_  = A233 & ~A203;
  assign \new_[14422]_  = A267 & A266;
  assign \new_[14423]_  = A234 & \new_[14422]_ ;
  assign \new_[14424]_  = \new_[14423]_  & \new_[14418]_ ;
  assign \new_[14427]_  = ~A167 & A170;
  assign \new_[14431]_  = ~A202 & ~A201;
  assign \new_[14432]_  = A166 & \new_[14431]_ ;
  assign \new_[14433]_  = \new_[14432]_  & \new_[14427]_ ;
  assign \new_[14436]_  = ~A232 & ~A203;
  assign \new_[14440]_  = A268 & A236;
  assign \new_[14441]_  = A233 & \new_[14440]_ ;
  assign \new_[14442]_  = \new_[14441]_  & \new_[14436]_ ;
  assign \new_[14445]_  = ~A167 & A170;
  assign \new_[14449]_  = ~A202 & ~A201;
  assign \new_[14450]_  = A166 & \new_[14449]_ ;
  assign \new_[14451]_  = \new_[14450]_  & \new_[14445]_ ;
  assign \new_[14454]_  = A232 & ~A203;
  assign \new_[14458]_  = A268 & A236;
  assign \new_[14459]_  = ~A233 & \new_[14458]_ ;
  assign \new_[14460]_  = \new_[14459]_  & \new_[14454]_ ;
  assign \new_[14463]_  = ~A167 & A170;
  assign \new_[14467]_  = A200 & A199;
  assign \new_[14468]_  = A166 & \new_[14467]_ ;
  assign \new_[14469]_  = \new_[14468]_  & \new_[14463]_ ;
  assign \new_[14472]_  = ~A202 & ~A201;
  assign \new_[14476]_  = A267 & A265;
  assign \new_[14477]_  = A235 & \new_[14476]_ ;
  assign \new_[14478]_  = \new_[14477]_  & \new_[14472]_ ;
  assign \new_[14481]_  = ~A167 & A170;
  assign \new_[14485]_  = A200 & A199;
  assign \new_[14486]_  = A166 & \new_[14485]_ ;
  assign \new_[14487]_  = \new_[14486]_  & \new_[14481]_ ;
  assign \new_[14490]_  = ~A202 & ~A201;
  assign \new_[14494]_  = A267 & A266;
  assign \new_[14495]_  = A235 & \new_[14494]_ ;
  assign \new_[14496]_  = \new_[14495]_  & \new_[14490]_ ;
  assign \new_[14499]_  = ~A167 & A170;
  assign \new_[14503]_  = A200 & A199;
  assign \new_[14504]_  = A166 & \new_[14503]_ ;
  assign \new_[14505]_  = \new_[14504]_  & \new_[14499]_ ;
  assign \new_[14508]_  = ~A202 & ~A201;
  assign \new_[14512]_  = A268 & A234;
  assign \new_[14513]_  = A232 & \new_[14512]_ ;
  assign \new_[14514]_  = \new_[14513]_  & \new_[14508]_ ;
  assign \new_[14517]_  = ~A167 & A170;
  assign \new_[14521]_  = A200 & A199;
  assign \new_[14522]_  = A166 & \new_[14521]_ ;
  assign \new_[14523]_  = \new_[14522]_  & \new_[14517]_ ;
  assign \new_[14526]_  = ~A202 & ~A201;
  assign \new_[14530]_  = A268 & A234;
  assign \new_[14531]_  = A233 & \new_[14530]_ ;
  assign \new_[14532]_  = \new_[14531]_  & \new_[14526]_ ;
  assign \new_[14535]_  = ~A167 & A170;
  assign \new_[14539]_  = ~A200 & ~A199;
  assign \new_[14540]_  = A166 & \new_[14539]_ ;
  assign \new_[14541]_  = \new_[14540]_  & \new_[14535]_ ;
  assign \new_[14544]_  = A235 & ~A202;
  assign \new_[14548]_  = ~A302 & ~A301;
  assign \new_[14549]_  = ~A300 & \new_[14548]_ ;
  assign \new_[14550]_  = \new_[14549]_  & \new_[14544]_ ;
  assign \new_[14553]_  = ~A167 & A170;
  assign \new_[14557]_  = ~A200 & ~A199;
  assign \new_[14558]_  = A166 & \new_[14557]_ ;
  assign \new_[14559]_  = \new_[14558]_  & \new_[14553]_ ;
  assign \new_[14562]_  = A235 & ~A202;
  assign \new_[14566]_  = ~A301 & ~A299;
  assign \new_[14567]_  = ~A298 & \new_[14566]_ ;
  assign \new_[14568]_  = \new_[14567]_  & \new_[14562]_ ;
  assign \new_[14571]_  = ~A167 & A170;
  assign \new_[14575]_  = ~A200 & ~A199;
  assign \new_[14576]_  = A166 & \new_[14575]_ ;
  assign \new_[14577]_  = \new_[14576]_  & \new_[14571]_ ;
  assign \new_[14580]_  = A235 & ~A202;
  assign \new_[14584]_  = A269 & A266;
  assign \new_[14585]_  = ~A265 & \new_[14584]_ ;
  assign \new_[14586]_  = \new_[14585]_  & \new_[14580]_ ;
  assign \new_[14589]_  = ~A167 & A170;
  assign \new_[14593]_  = ~A200 & ~A199;
  assign \new_[14594]_  = A166 & \new_[14593]_ ;
  assign \new_[14595]_  = \new_[14594]_  & \new_[14589]_ ;
  assign \new_[14598]_  = A235 & ~A202;
  assign \new_[14602]_  = A269 & ~A266;
  assign \new_[14603]_  = A265 & \new_[14602]_ ;
  assign \new_[14604]_  = \new_[14603]_  & \new_[14598]_ ;
  assign \new_[14607]_  = ~A167 & A170;
  assign \new_[14611]_  = ~A200 & ~A199;
  assign \new_[14612]_  = A166 & \new_[14611]_ ;
  assign \new_[14613]_  = \new_[14612]_  & \new_[14607]_ ;
  assign \new_[14616]_  = A232 & ~A202;
  assign \new_[14620]_  = A267 & A265;
  assign \new_[14621]_  = A234 & \new_[14620]_ ;
  assign \new_[14622]_  = \new_[14621]_  & \new_[14616]_ ;
  assign \new_[14625]_  = ~A167 & A170;
  assign \new_[14629]_  = ~A200 & ~A199;
  assign \new_[14630]_  = A166 & \new_[14629]_ ;
  assign \new_[14631]_  = \new_[14630]_  & \new_[14625]_ ;
  assign \new_[14634]_  = A232 & ~A202;
  assign \new_[14638]_  = A267 & A266;
  assign \new_[14639]_  = A234 & \new_[14638]_ ;
  assign \new_[14640]_  = \new_[14639]_  & \new_[14634]_ ;
  assign \new_[14643]_  = ~A167 & A170;
  assign \new_[14647]_  = ~A200 & ~A199;
  assign \new_[14648]_  = A166 & \new_[14647]_ ;
  assign \new_[14649]_  = \new_[14648]_  & \new_[14643]_ ;
  assign \new_[14652]_  = A233 & ~A202;
  assign \new_[14656]_  = A267 & A265;
  assign \new_[14657]_  = A234 & \new_[14656]_ ;
  assign \new_[14658]_  = \new_[14657]_  & \new_[14652]_ ;
  assign \new_[14661]_  = ~A167 & A170;
  assign \new_[14665]_  = ~A200 & ~A199;
  assign \new_[14666]_  = A166 & \new_[14665]_ ;
  assign \new_[14667]_  = \new_[14666]_  & \new_[14661]_ ;
  assign \new_[14670]_  = A233 & ~A202;
  assign \new_[14674]_  = A267 & A266;
  assign \new_[14675]_  = A234 & \new_[14674]_ ;
  assign \new_[14676]_  = \new_[14675]_  & \new_[14670]_ ;
  assign \new_[14679]_  = ~A167 & A170;
  assign \new_[14683]_  = ~A200 & ~A199;
  assign \new_[14684]_  = A166 & \new_[14683]_ ;
  assign \new_[14685]_  = \new_[14684]_  & \new_[14679]_ ;
  assign \new_[14688]_  = ~A232 & ~A202;
  assign \new_[14692]_  = A268 & A236;
  assign \new_[14693]_  = A233 & \new_[14692]_ ;
  assign \new_[14694]_  = \new_[14693]_  & \new_[14688]_ ;
  assign \new_[14697]_  = ~A167 & A170;
  assign \new_[14701]_  = ~A200 & ~A199;
  assign \new_[14702]_  = A166 & \new_[14701]_ ;
  assign \new_[14703]_  = \new_[14702]_  & \new_[14697]_ ;
  assign \new_[14706]_  = A232 & ~A202;
  assign \new_[14710]_  = A268 & A236;
  assign \new_[14711]_  = ~A233 & \new_[14710]_ ;
  assign \new_[14712]_  = \new_[14711]_  & \new_[14706]_ ;
  assign \new_[14715]_  = ~A201 & A169;
  assign \new_[14719]_  = A232 & ~A203;
  assign \new_[14720]_  = ~A202 & \new_[14719]_ ;
  assign \new_[14721]_  = \new_[14720]_  & \new_[14715]_ ;
  assign \new_[14724]_  = A298 & A234;
  assign \new_[14728]_  = ~A301 & ~A300;
  assign \new_[14729]_  = A299 & \new_[14728]_ ;
  assign \new_[14730]_  = \new_[14729]_  & \new_[14724]_ ;
  assign \new_[14733]_  = ~A201 & A169;
  assign \new_[14737]_  = A233 & ~A203;
  assign \new_[14738]_  = ~A202 & \new_[14737]_ ;
  assign \new_[14739]_  = \new_[14738]_  & \new_[14733]_ ;
  assign \new_[14742]_  = A298 & A234;
  assign \new_[14746]_  = ~A301 & ~A300;
  assign \new_[14747]_  = A299 & \new_[14746]_ ;
  assign \new_[14748]_  = \new_[14747]_  & \new_[14742]_ ;
  assign \new_[14751]_  = ~A201 & A169;
  assign \new_[14755]_  = ~A232 & ~A203;
  assign \new_[14756]_  = ~A202 & \new_[14755]_ ;
  assign \new_[14757]_  = \new_[14756]_  & \new_[14751]_ ;
  assign \new_[14760]_  = A236 & A233;
  assign \new_[14764]_  = ~A302 & ~A301;
  assign \new_[14765]_  = ~A300 & \new_[14764]_ ;
  assign \new_[14766]_  = \new_[14765]_  & \new_[14760]_ ;
  assign \new_[14769]_  = ~A201 & A169;
  assign \new_[14773]_  = ~A232 & ~A203;
  assign \new_[14774]_  = ~A202 & \new_[14773]_ ;
  assign \new_[14775]_  = \new_[14774]_  & \new_[14769]_ ;
  assign \new_[14778]_  = A236 & A233;
  assign \new_[14782]_  = ~A301 & ~A299;
  assign \new_[14783]_  = ~A298 & \new_[14782]_ ;
  assign \new_[14784]_  = \new_[14783]_  & \new_[14778]_ ;
  assign \new_[14787]_  = ~A201 & A169;
  assign \new_[14791]_  = ~A232 & ~A203;
  assign \new_[14792]_  = ~A202 & \new_[14791]_ ;
  assign \new_[14793]_  = \new_[14792]_  & \new_[14787]_ ;
  assign \new_[14796]_  = A236 & A233;
  assign \new_[14800]_  = A269 & A266;
  assign \new_[14801]_  = ~A265 & \new_[14800]_ ;
  assign \new_[14802]_  = \new_[14801]_  & \new_[14796]_ ;
  assign \new_[14805]_  = ~A201 & A169;
  assign \new_[14809]_  = ~A232 & ~A203;
  assign \new_[14810]_  = ~A202 & \new_[14809]_ ;
  assign \new_[14811]_  = \new_[14810]_  & \new_[14805]_ ;
  assign \new_[14814]_  = A236 & A233;
  assign \new_[14818]_  = A269 & ~A266;
  assign \new_[14819]_  = A265 & \new_[14818]_ ;
  assign \new_[14820]_  = \new_[14819]_  & \new_[14814]_ ;
  assign \new_[14823]_  = ~A201 & A169;
  assign \new_[14827]_  = A232 & ~A203;
  assign \new_[14828]_  = ~A202 & \new_[14827]_ ;
  assign \new_[14829]_  = \new_[14828]_  & \new_[14823]_ ;
  assign \new_[14832]_  = A236 & ~A233;
  assign \new_[14836]_  = ~A302 & ~A301;
  assign \new_[14837]_  = ~A300 & \new_[14836]_ ;
  assign \new_[14838]_  = \new_[14837]_  & \new_[14832]_ ;
  assign \new_[14841]_  = ~A201 & A169;
  assign \new_[14845]_  = A232 & ~A203;
  assign \new_[14846]_  = ~A202 & \new_[14845]_ ;
  assign \new_[14847]_  = \new_[14846]_  & \new_[14841]_ ;
  assign \new_[14850]_  = A236 & ~A233;
  assign \new_[14854]_  = ~A301 & ~A299;
  assign \new_[14855]_  = ~A298 & \new_[14854]_ ;
  assign \new_[14856]_  = \new_[14855]_  & \new_[14850]_ ;
  assign \new_[14859]_  = ~A201 & A169;
  assign \new_[14863]_  = A232 & ~A203;
  assign \new_[14864]_  = ~A202 & \new_[14863]_ ;
  assign \new_[14865]_  = \new_[14864]_  & \new_[14859]_ ;
  assign \new_[14868]_  = A236 & ~A233;
  assign \new_[14872]_  = A269 & A266;
  assign \new_[14873]_  = ~A265 & \new_[14872]_ ;
  assign \new_[14874]_  = \new_[14873]_  & \new_[14868]_ ;
  assign \new_[14877]_  = ~A201 & A169;
  assign \new_[14881]_  = A232 & ~A203;
  assign \new_[14882]_  = ~A202 & \new_[14881]_ ;
  assign \new_[14883]_  = \new_[14882]_  & \new_[14877]_ ;
  assign \new_[14886]_  = A236 & ~A233;
  assign \new_[14890]_  = A269 & ~A266;
  assign \new_[14891]_  = A265 & \new_[14890]_ ;
  assign \new_[14892]_  = \new_[14891]_  & \new_[14886]_ ;
  assign \new_[14895]_  = A199 & A169;
  assign \new_[14899]_  = ~A202 & ~A201;
  assign \new_[14900]_  = A200 & \new_[14899]_ ;
  assign \new_[14901]_  = \new_[14900]_  & \new_[14895]_ ;
  assign \new_[14904]_  = A298 & A235;
  assign \new_[14908]_  = ~A301 & ~A300;
  assign \new_[14909]_  = A299 & \new_[14908]_ ;
  assign \new_[14910]_  = \new_[14909]_  & \new_[14904]_ ;
  assign \new_[14913]_  = A199 & A169;
  assign \new_[14917]_  = ~A202 & ~A201;
  assign \new_[14918]_  = A200 & \new_[14917]_ ;
  assign \new_[14919]_  = \new_[14918]_  & \new_[14913]_ ;
  assign \new_[14922]_  = A234 & A232;
  assign \new_[14926]_  = ~A302 & ~A301;
  assign \new_[14927]_  = ~A300 & \new_[14926]_ ;
  assign \new_[14928]_  = \new_[14927]_  & \new_[14922]_ ;
  assign \new_[14931]_  = A199 & A169;
  assign \new_[14935]_  = ~A202 & ~A201;
  assign \new_[14936]_  = A200 & \new_[14935]_ ;
  assign \new_[14937]_  = \new_[14936]_  & \new_[14931]_ ;
  assign \new_[14940]_  = A234 & A232;
  assign \new_[14944]_  = ~A301 & ~A299;
  assign \new_[14945]_  = ~A298 & \new_[14944]_ ;
  assign \new_[14946]_  = \new_[14945]_  & \new_[14940]_ ;
  assign \new_[14949]_  = A199 & A169;
  assign \new_[14953]_  = ~A202 & ~A201;
  assign \new_[14954]_  = A200 & \new_[14953]_ ;
  assign \new_[14955]_  = \new_[14954]_  & \new_[14949]_ ;
  assign \new_[14958]_  = A234 & A232;
  assign \new_[14962]_  = A269 & A266;
  assign \new_[14963]_  = ~A265 & \new_[14962]_ ;
  assign \new_[14964]_  = \new_[14963]_  & \new_[14958]_ ;
  assign \new_[14967]_  = A199 & A169;
  assign \new_[14971]_  = ~A202 & ~A201;
  assign \new_[14972]_  = A200 & \new_[14971]_ ;
  assign \new_[14973]_  = \new_[14972]_  & \new_[14967]_ ;
  assign \new_[14976]_  = A234 & A232;
  assign \new_[14980]_  = A269 & ~A266;
  assign \new_[14981]_  = A265 & \new_[14980]_ ;
  assign \new_[14982]_  = \new_[14981]_  & \new_[14976]_ ;
  assign \new_[14985]_  = A199 & A169;
  assign \new_[14989]_  = ~A202 & ~A201;
  assign \new_[14990]_  = A200 & \new_[14989]_ ;
  assign \new_[14991]_  = \new_[14990]_  & \new_[14985]_ ;
  assign \new_[14994]_  = A234 & A233;
  assign \new_[14998]_  = ~A302 & ~A301;
  assign \new_[14999]_  = ~A300 & \new_[14998]_ ;
  assign \new_[15000]_  = \new_[14999]_  & \new_[14994]_ ;
  assign \new_[15003]_  = A199 & A169;
  assign \new_[15007]_  = ~A202 & ~A201;
  assign \new_[15008]_  = A200 & \new_[15007]_ ;
  assign \new_[15009]_  = \new_[15008]_  & \new_[15003]_ ;
  assign \new_[15012]_  = A234 & A233;
  assign \new_[15016]_  = ~A301 & ~A299;
  assign \new_[15017]_  = ~A298 & \new_[15016]_ ;
  assign \new_[15018]_  = \new_[15017]_  & \new_[15012]_ ;
  assign \new_[15021]_  = A199 & A169;
  assign \new_[15025]_  = ~A202 & ~A201;
  assign \new_[15026]_  = A200 & \new_[15025]_ ;
  assign \new_[15027]_  = \new_[15026]_  & \new_[15021]_ ;
  assign \new_[15030]_  = A234 & A233;
  assign \new_[15034]_  = A269 & A266;
  assign \new_[15035]_  = ~A265 & \new_[15034]_ ;
  assign \new_[15036]_  = \new_[15035]_  & \new_[15030]_ ;
  assign \new_[15039]_  = A199 & A169;
  assign \new_[15043]_  = ~A202 & ~A201;
  assign \new_[15044]_  = A200 & \new_[15043]_ ;
  assign \new_[15045]_  = \new_[15044]_  & \new_[15039]_ ;
  assign \new_[15048]_  = A234 & A233;
  assign \new_[15052]_  = A269 & ~A266;
  assign \new_[15053]_  = A265 & \new_[15052]_ ;
  assign \new_[15054]_  = \new_[15053]_  & \new_[15048]_ ;
  assign \new_[15057]_  = A199 & A169;
  assign \new_[15061]_  = ~A202 & ~A201;
  assign \new_[15062]_  = A200 & \new_[15061]_ ;
  assign \new_[15063]_  = \new_[15062]_  & \new_[15057]_ ;
  assign \new_[15066]_  = A233 & ~A232;
  assign \new_[15070]_  = A267 & A265;
  assign \new_[15071]_  = A236 & \new_[15070]_ ;
  assign \new_[15072]_  = \new_[15071]_  & \new_[15066]_ ;
  assign \new_[15075]_  = A199 & A169;
  assign \new_[15079]_  = ~A202 & ~A201;
  assign \new_[15080]_  = A200 & \new_[15079]_ ;
  assign \new_[15081]_  = \new_[15080]_  & \new_[15075]_ ;
  assign \new_[15084]_  = A233 & ~A232;
  assign \new_[15088]_  = A267 & A266;
  assign \new_[15089]_  = A236 & \new_[15088]_ ;
  assign \new_[15090]_  = \new_[15089]_  & \new_[15084]_ ;
  assign \new_[15093]_  = A199 & A169;
  assign \new_[15097]_  = ~A202 & ~A201;
  assign \new_[15098]_  = A200 & \new_[15097]_ ;
  assign \new_[15099]_  = \new_[15098]_  & \new_[15093]_ ;
  assign \new_[15102]_  = ~A233 & A232;
  assign \new_[15106]_  = A267 & A265;
  assign \new_[15107]_  = A236 & \new_[15106]_ ;
  assign \new_[15108]_  = \new_[15107]_  & \new_[15102]_ ;
  assign \new_[15111]_  = A199 & A169;
  assign \new_[15115]_  = ~A202 & ~A201;
  assign \new_[15116]_  = A200 & \new_[15115]_ ;
  assign \new_[15117]_  = \new_[15116]_  & \new_[15111]_ ;
  assign \new_[15120]_  = ~A233 & A232;
  assign \new_[15124]_  = A267 & A266;
  assign \new_[15125]_  = A236 & \new_[15124]_ ;
  assign \new_[15126]_  = \new_[15125]_  & \new_[15120]_ ;
  assign \new_[15129]_  = ~A199 & A169;
  assign \new_[15133]_  = A232 & ~A202;
  assign \new_[15134]_  = ~A200 & \new_[15133]_ ;
  assign \new_[15135]_  = \new_[15134]_  & \new_[15129]_ ;
  assign \new_[15138]_  = A298 & A234;
  assign \new_[15142]_  = ~A301 & ~A300;
  assign \new_[15143]_  = A299 & \new_[15142]_ ;
  assign \new_[15144]_  = \new_[15143]_  & \new_[15138]_ ;
  assign \new_[15147]_  = ~A199 & A169;
  assign \new_[15151]_  = A233 & ~A202;
  assign \new_[15152]_  = ~A200 & \new_[15151]_ ;
  assign \new_[15153]_  = \new_[15152]_  & \new_[15147]_ ;
  assign \new_[15156]_  = A298 & A234;
  assign \new_[15160]_  = ~A301 & ~A300;
  assign \new_[15161]_  = A299 & \new_[15160]_ ;
  assign \new_[15162]_  = \new_[15161]_  & \new_[15156]_ ;
  assign \new_[15165]_  = ~A199 & A169;
  assign \new_[15169]_  = ~A232 & ~A202;
  assign \new_[15170]_  = ~A200 & \new_[15169]_ ;
  assign \new_[15171]_  = \new_[15170]_  & \new_[15165]_ ;
  assign \new_[15174]_  = A236 & A233;
  assign \new_[15178]_  = ~A302 & ~A301;
  assign \new_[15179]_  = ~A300 & \new_[15178]_ ;
  assign \new_[15180]_  = \new_[15179]_  & \new_[15174]_ ;
  assign \new_[15183]_  = ~A199 & A169;
  assign \new_[15187]_  = ~A232 & ~A202;
  assign \new_[15188]_  = ~A200 & \new_[15187]_ ;
  assign \new_[15189]_  = \new_[15188]_  & \new_[15183]_ ;
  assign \new_[15192]_  = A236 & A233;
  assign \new_[15196]_  = ~A301 & ~A299;
  assign \new_[15197]_  = ~A298 & \new_[15196]_ ;
  assign \new_[15198]_  = \new_[15197]_  & \new_[15192]_ ;
  assign \new_[15201]_  = ~A199 & A169;
  assign \new_[15205]_  = ~A232 & ~A202;
  assign \new_[15206]_  = ~A200 & \new_[15205]_ ;
  assign \new_[15207]_  = \new_[15206]_  & \new_[15201]_ ;
  assign \new_[15210]_  = A236 & A233;
  assign \new_[15214]_  = A269 & A266;
  assign \new_[15215]_  = ~A265 & \new_[15214]_ ;
  assign \new_[15216]_  = \new_[15215]_  & \new_[15210]_ ;
  assign \new_[15219]_  = ~A199 & A169;
  assign \new_[15223]_  = ~A232 & ~A202;
  assign \new_[15224]_  = ~A200 & \new_[15223]_ ;
  assign \new_[15225]_  = \new_[15224]_  & \new_[15219]_ ;
  assign \new_[15228]_  = A236 & A233;
  assign \new_[15232]_  = A269 & ~A266;
  assign \new_[15233]_  = A265 & \new_[15232]_ ;
  assign \new_[15234]_  = \new_[15233]_  & \new_[15228]_ ;
  assign \new_[15237]_  = ~A199 & A169;
  assign \new_[15241]_  = A232 & ~A202;
  assign \new_[15242]_  = ~A200 & \new_[15241]_ ;
  assign \new_[15243]_  = \new_[15242]_  & \new_[15237]_ ;
  assign \new_[15246]_  = A236 & ~A233;
  assign \new_[15250]_  = ~A302 & ~A301;
  assign \new_[15251]_  = ~A300 & \new_[15250]_ ;
  assign \new_[15252]_  = \new_[15251]_  & \new_[15246]_ ;
  assign \new_[15255]_  = ~A199 & A169;
  assign \new_[15259]_  = A232 & ~A202;
  assign \new_[15260]_  = ~A200 & \new_[15259]_ ;
  assign \new_[15261]_  = \new_[15260]_  & \new_[15255]_ ;
  assign \new_[15264]_  = A236 & ~A233;
  assign \new_[15268]_  = ~A301 & ~A299;
  assign \new_[15269]_  = ~A298 & \new_[15268]_ ;
  assign \new_[15270]_  = \new_[15269]_  & \new_[15264]_ ;
  assign \new_[15273]_  = ~A199 & A169;
  assign \new_[15277]_  = A232 & ~A202;
  assign \new_[15278]_  = ~A200 & \new_[15277]_ ;
  assign \new_[15279]_  = \new_[15278]_  & \new_[15273]_ ;
  assign \new_[15282]_  = A236 & ~A233;
  assign \new_[15286]_  = A269 & A266;
  assign \new_[15287]_  = ~A265 & \new_[15286]_ ;
  assign \new_[15288]_  = \new_[15287]_  & \new_[15282]_ ;
  assign \new_[15291]_  = ~A199 & A169;
  assign \new_[15295]_  = A232 & ~A202;
  assign \new_[15296]_  = ~A200 & \new_[15295]_ ;
  assign \new_[15297]_  = \new_[15296]_  & \new_[15291]_ ;
  assign \new_[15300]_  = A236 & ~A233;
  assign \new_[15304]_  = A269 & ~A266;
  assign \new_[15305]_  = A265 & \new_[15304]_ ;
  assign \new_[15306]_  = \new_[15305]_  & \new_[15300]_ ;
  assign \new_[15309]_  = ~A167 & ~A169;
  assign \new_[15313]_  = A232 & A202;
  assign \new_[15314]_  = ~A166 & \new_[15313]_ ;
  assign \new_[15315]_  = \new_[15314]_  & \new_[15309]_ ;
  assign \new_[15318]_  = A298 & A234;
  assign \new_[15322]_  = ~A301 & ~A300;
  assign \new_[15323]_  = A299 & \new_[15322]_ ;
  assign \new_[15324]_  = \new_[15323]_  & \new_[15318]_ ;
  assign \new_[15327]_  = ~A167 & ~A169;
  assign \new_[15331]_  = A233 & A202;
  assign \new_[15332]_  = ~A166 & \new_[15331]_ ;
  assign \new_[15333]_  = \new_[15332]_  & \new_[15327]_ ;
  assign \new_[15336]_  = A298 & A234;
  assign \new_[15340]_  = ~A301 & ~A300;
  assign \new_[15341]_  = A299 & \new_[15340]_ ;
  assign \new_[15342]_  = \new_[15341]_  & \new_[15336]_ ;
  assign \new_[15345]_  = ~A167 & ~A169;
  assign \new_[15349]_  = ~A232 & A202;
  assign \new_[15350]_  = ~A166 & \new_[15349]_ ;
  assign \new_[15351]_  = \new_[15350]_  & \new_[15345]_ ;
  assign \new_[15354]_  = A236 & A233;
  assign \new_[15358]_  = ~A302 & ~A301;
  assign \new_[15359]_  = ~A300 & \new_[15358]_ ;
  assign \new_[15360]_  = \new_[15359]_  & \new_[15354]_ ;
  assign \new_[15363]_  = ~A167 & ~A169;
  assign \new_[15367]_  = ~A232 & A202;
  assign \new_[15368]_  = ~A166 & \new_[15367]_ ;
  assign \new_[15369]_  = \new_[15368]_  & \new_[15363]_ ;
  assign \new_[15372]_  = A236 & A233;
  assign \new_[15376]_  = ~A301 & ~A299;
  assign \new_[15377]_  = ~A298 & \new_[15376]_ ;
  assign \new_[15378]_  = \new_[15377]_  & \new_[15372]_ ;
  assign \new_[15381]_  = ~A167 & ~A169;
  assign \new_[15385]_  = ~A232 & A202;
  assign \new_[15386]_  = ~A166 & \new_[15385]_ ;
  assign \new_[15387]_  = \new_[15386]_  & \new_[15381]_ ;
  assign \new_[15390]_  = A236 & A233;
  assign \new_[15394]_  = A269 & A266;
  assign \new_[15395]_  = ~A265 & \new_[15394]_ ;
  assign \new_[15396]_  = \new_[15395]_  & \new_[15390]_ ;
  assign \new_[15399]_  = ~A167 & ~A169;
  assign \new_[15403]_  = ~A232 & A202;
  assign \new_[15404]_  = ~A166 & \new_[15403]_ ;
  assign \new_[15405]_  = \new_[15404]_  & \new_[15399]_ ;
  assign \new_[15408]_  = A236 & A233;
  assign \new_[15412]_  = A269 & ~A266;
  assign \new_[15413]_  = A265 & \new_[15412]_ ;
  assign \new_[15414]_  = \new_[15413]_  & \new_[15408]_ ;
  assign \new_[15417]_  = ~A167 & ~A169;
  assign \new_[15421]_  = A232 & A202;
  assign \new_[15422]_  = ~A166 & \new_[15421]_ ;
  assign \new_[15423]_  = \new_[15422]_  & \new_[15417]_ ;
  assign \new_[15426]_  = A236 & ~A233;
  assign \new_[15430]_  = ~A302 & ~A301;
  assign \new_[15431]_  = ~A300 & \new_[15430]_ ;
  assign \new_[15432]_  = \new_[15431]_  & \new_[15426]_ ;
  assign \new_[15435]_  = ~A167 & ~A169;
  assign \new_[15439]_  = A232 & A202;
  assign \new_[15440]_  = ~A166 & \new_[15439]_ ;
  assign \new_[15441]_  = \new_[15440]_  & \new_[15435]_ ;
  assign \new_[15444]_  = A236 & ~A233;
  assign \new_[15448]_  = ~A301 & ~A299;
  assign \new_[15449]_  = ~A298 & \new_[15448]_ ;
  assign \new_[15450]_  = \new_[15449]_  & \new_[15444]_ ;
  assign \new_[15453]_  = ~A167 & ~A169;
  assign \new_[15457]_  = A232 & A202;
  assign \new_[15458]_  = ~A166 & \new_[15457]_ ;
  assign \new_[15459]_  = \new_[15458]_  & \new_[15453]_ ;
  assign \new_[15462]_  = A236 & ~A233;
  assign \new_[15466]_  = A269 & A266;
  assign \new_[15467]_  = ~A265 & \new_[15466]_ ;
  assign \new_[15468]_  = \new_[15467]_  & \new_[15462]_ ;
  assign \new_[15471]_  = ~A167 & ~A169;
  assign \new_[15475]_  = A232 & A202;
  assign \new_[15476]_  = ~A166 & \new_[15475]_ ;
  assign \new_[15477]_  = \new_[15476]_  & \new_[15471]_ ;
  assign \new_[15480]_  = A236 & ~A233;
  assign \new_[15484]_  = A269 & ~A266;
  assign \new_[15485]_  = A265 & \new_[15484]_ ;
  assign \new_[15486]_  = \new_[15485]_  & \new_[15480]_ ;
  assign \new_[15489]_  = ~A167 & ~A169;
  assign \new_[15493]_  = A201 & A199;
  assign \new_[15494]_  = ~A166 & \new_[15493]_ ;
  assign \new_[15495]_  = \new_[15494]_  & \new_[15489]_ ;
  assign \new_[15498]_  = A298 & A235;
  assign \new_[15502]_  = ~A301 & ~A300;
  assign \new_[15503]_  = A299 & \new_[15502]_ ;
  assign \new_[15504]_  = \new_[15503]_  & \new_[15498]_ ;
  assign \new_[15507]_  = ~A167 & ~A169;
  assign \new_[15511]_  = A201 & A199;
  assign \new_[15512]_  = ~A166 & \new_[15511]_ ;
  assign \new_[15513]_  = \new_[15512]_  & \new_[15507]_ ;
  assign \new_[15516]_  = A234 & A232;
  assign \new_[15520]_  = ~A302 & ~A301;
  assign \new_[15521]_  = ~A300 & \new_[15520]_ ;
  assign \new_[15522]_  = \new_[15521]_  & \new_[15516]_ ;
  assign \new_[15525]_  = ~A167 & ~A169;
  assign \new_[15529]_  = A201 & A199;
  assign \new_[15530]_  = ~A166 & \new_[15529]_ ;
  assign \new_[15531]_  = \new_[15530]_  & \new_[15525]_ ;
  assign \new_[15534]_  = A234 & A232;
  assign \new_[15538]_  = ~A301 & ~A299;
  assign \new_[15539]_  = ~A298 & \new_[15538]_ ;
  assign \new_[15540]_  = \new_[15539]_  & \new_[15534]_ ;
  assign \new_[15543]_  = ~A167 & ~A169;
  assign \new_[15547]_  = A201 & A199;
  assign \new_[15548]_  = ~A166 & \new_[15547]_ ;
  assign \new_[15549]_  = \new_[15548]_  & \new_[15543]_ ;
  assign \new_[15552]_  = A234 & A232;
  assign \new_[15556]_  = A269 & A266;
  assign \new_[15557]_  = ~A265 & \new_[15556]_ ;
  assign \new_[15558]_  = \new_[15557]_  & \new_[15552]_ ;
  assign \new_[15561]_  = ~A167 & ~A169;
  assign \new_[15565]_  = A201 & A199;
  assign \new_[15566]_  = ~A166 & \new_[15565]_ ;
  assign \new_[15567]_  = \new_[15566]_  & \new_[15561]_ ;
  assign \new_[15570]_  = A234 & A232;
  assign \new_[15574]_  = A269 & ~A266;
  assign \new_[15575]_  = A265 & \new_[15574]_ ;
  assign \new_[15576]_  = \new_[15575]_  & \new_[15570]_ ;
  assign \new_[15579]_  = ~A167 & ~A169;
  assign \new_[15583]_  = A201 & A199;
  assign \new_[15584]_  = ~A166 & \new_[15583]_ ;
  assign \new_[15585]_  = \new_[15584]_  & \new_[15579]_ ;
  assign \new_[15588]_  = A234 & A233;
  assign \new_[15592]_  = ~A302 & ~A301;
  assign \new_[15593]_  = ~A300 & \new_[15592]_ ;
  assign \new_[15594]_  = \new_[15593]_  & \new_[15588]_ ;
  assign \new_[15597]_  = ~A167 & ~A169;
  assign \new_[15601]_  = A201 & A199;
  assign \new_[15602]_  = ~A166 & \new_[15601]_ ;
  assign \new_[15603]_  = \new_[15602]_  & \new_[15597]_ ;
  assign \new_[15606]_  = A234 & A233;
  assign \new_[15610]_  = ~A301 & ~A299;
  assign \new_[15611]_  = ~A298 & \new_[15610]_ ;
  assign \new_[15612]_  = \new_[15611]_  & \new_[15606]_ ;
  assign \new_[15615]_  = ~A167 & ~A169;
  assign \new_[15619]_  = A201 & A199;
  assign \new_[15620]_  = ~A166 & \new_[15619]_ ;
  assign \new_[15621]_  = \new_[15620]_  & \new_[15615]_ ;
  assign \new_[15624]_  = A234 & A233;
  assign \new_[15628]_  = A269 & A266;
  assign \new_[15629]_  = ~A265 & \new_[15628]_ ;
  assign \new_[15630]_  = \new_[15629]_  & \new_[15624]_ ;
  assign \new_[15633]_  = ~A167 & ~A169;
  assign \new_[15637]_  = A201 & A199;
  assign \new_[15638]_  = ~A166 & \new_[15637]_ ;
  assign \new_[15639]_  = \new_[15638]_  & \new_[15633]_ ;
  assign \new_[15642]_  = A234 & A233;
  assign \new_[15646]_  = A269 & ~A266;
  assign \new_[15647]_  = A265 & \new_[15646]_ ;
  assign \new_[15648]_  = \new_[15647]_  & \new_[15642]_ ;
  assign \new_[15651]_  = ~A167 & ~A169;
  assign \new_[15655]_  = A201 & A199;
  assign \new_[15656]_  = ~A166 & \new_[15655]_ ;
  assign \new_[15657]_  = \new_[15656]_  & \new_[15651]_ ;
  assign \new_[15660]_  = A233 & ~A232;
  assign \new_[15664]_  = A267 & A265;
  assign \new_[15665]_  = A236 & \new_[15664]_ ;
  assign \new_[15666]_  = \new_[15665]_  & \new_[15660]_ ;
  assign \new_[15669]_  = ~A167 & ~A169;
  assign \new_[15673]_  = A201 & A199;
  assign \new_[15674]_  = ~A166 & \new_[15673]_ ;
  assign \new_[15675]_  = \new_[15674]_  & \new_[15669]_ ;
  assign \new_[15678]_  = A233 & ~A232;
  assign \new_[15682]_  = A267 & A266;
  assign \new_[15683]_  = A236 & \new_[15682]_ ;
  assign \new_[15684]_  = \new_[15683]_  & \new_[15678]_ ;
  assign \new_[15687]_  = ~A167 & ~A169;
  assign \new_[15691]_  = A201 & A199;
  assign \new_[15692]_  = ~A166 & \new_[15691]_ ;
  assign \new_[15693]_  = \new_[15692]_  & \new_[15687]_ ;
  assign \new_[15696]_  = ~A233 & A232;
  assign \new_[15700]_  = A267 & A265;
  assign \new_[15701]_  = A236 & \new_[15700]_ ;
  assign \new_[15702]_  = \new_[15701]_  & \new_[15696]_ ;
  assign \new_[15705]_  = ~A167 & ~A169;
  assign \new_[15709]_  = A201 & A199;
  assign \new_[15710]_  = ~A166 & \new_[15709]_ ;
  assign \new_[15711]_  = \new_[15710]_  & \new_[15705]_ ;
  assign \new_[15714]_  = ~A233 & A232;
  assign \new_[15718]_  = A267 & A266;
  assign \new_[15719]_  = A236 & \new_[15718]_ ;
  assign \new_[15720]_  = \new_[15719]_  & \new_[15714]_ ;
  assign \new_[15723]_  = ~A167 & ~A169;
  assign \new_[15727]_  = A201 & A200;
  assign \new_[15728]_  = ~A166 & \new_[15727]_ ;
  assign \new_[15729]_  = \new_[15728]_  & \new_[15723]_ ;
  assign \new_[15732]_  = A298 & A235;
  assign \new_[15736]_  = ~A301 & ~A300;
  assign \new_[15737]_  = A299 & \new_[15736]_ ;
  assign \new_[15738]_  = \new_[15737]_  & \new_[15732]_ ;
  assign \new_[15741]_  = ~A167 & ~A169;
  assign \new_[15745]_  = A201 & A200;
  assign \new_[15746]_  = ~A166 & \new_[15745]_ ;
  assign \new_[15747]_  = \new_[15746]_  & \new_[15741]_ ;
  assign \new_[15750]_  = A234 & A232;
  assign \new_[15754]_  = ~A302 & ~A301;
  assign \new_[15755]_  = ~A300 & \new_[15754]_ ;
  assign \new_[15756]_  = \new_[15755]_  & \new_[15750]_ ;
  assign \new_[15759]_  = ~A167 & ~A169;
  assign \new_[15763]_  = A201 & A200;
  assign \new_[15764]_  = ~A166 & \new_[15763]_ ;
  assign \new_[15765]_  = \new_[15764]_  & \new_[15759]_ ;
  assign \new_[15768]_  = A234 & A232;
  assign \new_[15772]_  = ~A301 & ~A299;
  assign \new_[15773]_  = ~A298 & \new_[15772]_ ;
  assign \new_[15774]_  = \new_[15773]_  & \new_[15768]_ ;
  assign \new_[15777]_  = ~A167 & ~A169;
  assign \new_[15781]_  = A201 & A200;
  assign \new_[15782]_  = ~A166 & \new_[15781]_ ;
  assign \new_[15783]_  = \new_[15782]_  & \new_[15777]_ ;
  assign \new_[15786]_  = A234 & A232;
  assign \new_[15790]_  = A269 & A266;
  assign \new_[15791]_  = ~A265 & \new_[15790]_ ;
  assign \new_[15792]_  = \new_[15791]_  & \new_[15786]_ ;
  assign \new_[15795]_  = ~A167 & ~A169;
  assign \new_[15799]_  = A201 & A200;
  assign \new_[15800]_  = ~A166 & \new_[15799]_ ;
  assign \new_[15801]_  = \new_[15800]_  & \new_[15795]_ ;
  assign \new_[15804]_  = A234 & A232;
  assign \new_[15808]_  = A269 & ~A266;
  assign \new_[15809]_  = A265 & \new_[15808]_ ;
  assign \new_[15810]_  = \new_[15809]_  & \new_[15804]_ ;
  assign \new_[15813]_  = ~A167 & ~A169;
  assign \new_[15817]_  = A201 & A200;
  assign \new_[15818]_  = ~A166 & \new_[15817]_ ;
  assign \new_[15819]_  = \new_[15818]_  & \new_[15813]_ ;
  assign \new_[15822]_  = A234 & A233;
  assign \new_[15826]_  = ~A302 & ~A301;
  assign \new_[15827]_  = ~A300 & \new_[15826]_ ;
  assign \new_[15828]_  = \new_[15827]_  & \new_[15822]_ ;
  assign \new_[15831]_  = ~A167 & ~A169;
  assign \new_[15835]_  = A201 & A200;
  assign \new_[15836]_  = ~A166 & \new_[15835]_ ;
  assign \new_[15837]_  = \new_[15836]_  & \new_[15831]_ ;
  assign \new_[15840]_  = A234 & A233;
  assign \new_[15844]_  = ~A301 & ~A299;
  assign \new_[15845]_  = ~A298 & \new_[15844]_ ;
  assign \new_[15846]_  = \new_[15845]_  & \new_[15840]_ ;
  assign \new_[15849]_  = ~A167 & ~A169;
  assign \new_[15853]_  = A201 & A200;
  assign \new_[15854]_  = ~A166 & \new_[15853]_ ;
  assign \new_[15855]_  = \new_[15854]_  & \new_[15849]_ ;
  assign \new_[15858]_  = A234 & A233;
  assign \new_[15862]_  = A269 & A266;
  assign \new_[15863]_  = ~A265 & \new_[15862]_ ;
  assign \new_[15864]_  = \new_[15863]_  & \new_[15858]_ ;
  assign \new_[15867]_  = ~A167 & ~A169;
  assign \new_[15871]_  = A201 & A200;
  assign \new_[15872]_  = ~A166 & \new_[15871]_ ;
  assign \new_[15873]_  = \new_[15872]_  & \new_[15867]_ ;
  assign \new_[15876]_  = A234 & A233;
  assign \new_[15880]_  = A269 & ~A266;
  assign \new_[15881]_  = A265 & \new_[15880]_ ;
  assign \new_[15882]_  = \new_[15881]_  & \new_[15876]_ ;
  assign \new_[15885]_  = ~A167 & ~A169;
  assign \new_[15889]_  = A201 & A200;
  assign \new_[15890]_  = ~A166 & \new_[15889]_ ;
  assign \new_[15891]_  = \new_[15890]_  & \new_[15885]_ ;
  assign \new_[15894]_  = A233 & ~A232;
  assign \new_[15898]_  = A267 & A265;
  assign \new_[15899]_  = A236 & \new_[15898]_ ;
  assign \new_[15900]_  = \new_[15899]_  & \new_[15894]_ ;
  assign \new_[15903]_  = ~A167 & ~A169;
  assign \new_[15907]_  = A201 & A200;
  assign \new_[15908]_  = ~A166 & \new_[15907]_ ;
  assign \new_[15909]_  = \new_[15908]_  & \new_[15903]_ ;
  assign \new_[15912]_  = A233 & ~A232;
  assign \new_[15916]_  = A267 & A266;
  assign \new_[15917]_  = A236 & \new_[15916]_ ;
  assign \new_[15918]_  = \new_[15917]_  & \new_[15912]_ ;
  assign \new_[15921]_  = ~A167 & ~A169;
  assign \new_[15925]_  = A201 & A200;
  assign \new_[15926]_  = ~A166 & \new_[15925]_ ;
  assign \new_[15927]_  = \new_[15926]_  & \new_[15921]_ ;
  assign \new_[15930]_  = ~A233 & A232;
  assign \new_[15934]_  = A267 & A265;
  assign \new_[15935]_  = A236 & \new_[15934]_ ;
  assign \new_[15936]_  = \new_[15935]_  & \new_[15930]_ ;
  assign \new_[15939]_  = ~A167 & ~A169;
  assign \new_[15943]_  = A201 & A200;
  assign \new_[15944]_  = ~A166 & \new_[15943]_ ;
  assign \new_[15945]_  = \new_[15944]_  & \new_[15939]_ ;
  assign \new_[15948]_  = ~A233 & A232;
  assign \new_[15952]_  = A267 & A266;
  assign \new_[15953]_  = A236 & \new_[15952]_ ;
  assign \new_[15954]_  = \new_[15953]_  & \new_[15948]_ ;
  assign \new_[15957]_  = ~A167 & ~A169;
  assign \new_[15961]_  = A200 & ~A199;
  assign \new_[15962]_  = ~A166 & \new_[15961]_ ;
  assign \new_[15963]_  = \new_[15962]_  & \new_[15957]_ ;
  assign \new_[15966]_  = A235 & A203;
  assign \new_[15970]_  = ~A302 & ~A301;
  assign \new_[15971]_  = ~A300 & \new_[15970]_ ;
  assign \new_[15972]_  = \new_[15971]_  & \new_[15966]_ ;
  assign \new_[15975]_  = ~A167 & ~A169;
  assign \new_[15979]_  = A200 & ~A199;
  assign \new_[15980]_  = ~A166 & \new_[15979]_ ;
  assign \new_[15981]_  = \new_[15980]_  & \new_[15975]_ ;
  assign \new_[15984]_  = A235 & A203;
  assign \new_[15988]_  = ~A301 & ~A299;
  assign \new_[15989]_  = ~A298 & \new_[15988]_ ;
  assign \new_[15990]_  = \new_[15989]_  & \new_[15984]_ ;
  assign \new_[15993]_  = ~A167 & ~A169;
  assign \new_[15997]_  = A200 & ~A199;
  assign \new_[15998]_  = ~A166 & \new_[15997]_ ;
  assign \new_[15999]_  = \new_[15998]_  & \new_[15993]_ ;
  assign \new_[16002]_  = A235 & A203;
  assign \new_[16006]_  = A269 & A266;
  assign \new_[16007]_  = ~A265 & \new_[16006]_ ;
  assign \new_[16008]_  = \new_[16007]_  & \new_[16002]_ ;
  assign \new_[16011]_  = ~A167 & ~A169;
  assign \new_[16015]_  = A200 & ~A199;
  assign \new_[16016]_  = ~A166 & \new_[16015]_ ;
  assign \new_[16017]_  = \new_[16016]_  & \new_[16011]_ ;
  assign \new_[16020]_  = A235 & A203;
  assign \new_[16024]_  = A269 & ~A266;
  assign \new_[16025]_  = A265 & \new_[16024]_ ;
  assign \new_[16026]_  = \new_[16025]_  & \new_[16020]_ ;
  assign \new_[16029]_  = ~A167 & ~A169;
  assign \new_[16033]_  = A200 & ~A199;
  assign \new_[16034]_  = ~A166 & \new_[16033]_ ;
  assign \new_[16035]_  = \new_[16034]_  & \new_[16029]_ ;
  assign \new_[16038]_  = A232 & A203;
  assign \new_[16042]_  = A267 & A265;
  assign \new_[16043]_  = A234 & \new_[16042]_ ;
  assign \new_[16044]_  = \new_[16043]_  & \new_[16038]_ ;
  assign \new_[16047]_  = ~A167 & ~A169;
  assign \new_[16051]_  = A200 & ~A199;
  assign \new_[16052]_  = ~A166 & \new_[16051]_ ;
  assign \new_[16053]_  = \new_[16052]_  & \new_[16047]_ ;
  assign \new_[16056]_  = A232 & A203;
  assign \new_[16060]_  = A267 & A266;
  assign \new_[16061]_  = A234 & \new_[16060]_ ;
  assign \new_[16062]_  = \new_[16061]_  & \new_[16056]_ ;
  assign \new_[16065]_  = ~A167 & ~A169;
  assign \new_[16069]_  = A200 & ~A199;
  assign \new_[16070]_  = ~A166 & \new_[16069]_ ;
  assign \new_[16071]_  = \new_[16070]_  & \new_[16065]_ ;
  assign \new_[16074]_  = A233 & A203;
  assign \new_[16078]_  = A267 & A265;
  assign \new_[16079]_  = A234 & \new_[16078]_ ;
  assign \new_[16080]_  = \new_[16079]_  & \new_[16074]_ ;
  assign \new_[16083]_  = ~A167 & ~A169;
  assign \new_[16087]_  = A200 & ~A199;
  assign \new_[16088]_  = ~A166 & \new_[16087]_ ;
  assign \new_[16089]_  = \new_[16088]_  & \new_[16083]_ ;
  assign \new_[16092]_  = A233 & A203;
  assign \new_[16096]_  = A267 & A266;
  assign \new_[16097]_  = A234 & \new_[16096]_ ;
  assign \new_[16098]_  = \new_[16097]_  & \new_[16092]_ ;
  assign \new_[16101]_  = ~A167 & ~A169;
  assign \new_[16105]_  = A200 & ~A199;
  assign \new_[16106]_  = ~A166 & \new_[16105]_ ;
  assign \new_[16107]_  = \new_[16106]_  & \new_[16101]_ ;
  assign \new_[16110]_  = ~A232 & A203;
  assign \new_[16114]_  = A268 & A236;
  assign \new_[16115]_  = A233 & \new_[16114]_ ;
  assign \new_[16116]_  = \new_[16115]_  & \new_[16110]_ ;
  assign \new_[16119]_  = ~A167 & ~A169;
  assign \new_[16123]_  = A200 & ~A199;
  assign \new_[16124]_  = ~A166 & \new_[16123]_ ;
  assign \new_[16125]_  = \new_[16124]_  & \new_[16119]_ ;
  assign \new_[16128]_  = A232 & A203;
  assign \new_[16132]_  = A268 & A236;
  assign \new_[16133]_  = ~A233 & \new_[16132]_ ;
  assign \new_[16134]_  = \new_[16133]_  & \new_[16128]_ ;
  assign \new_[16137]_  = ~A167 & ~A169;
  assign \new_[16141]_  = ~A200 & A199;
  assign \new_[16142]_  = ~A166 & \new_[16141]_ ;
  assign \new_[16143]_  = \new_[16142]_  & \new_[16137]_ ;
  assign \new_[16146]_  = A235 & A203;
  assign \new_[16150]_  = ~A302 & ~A301;
  assign \new_[16151]_  = ~A300 & \new_[16150]_ ;
  assign \new_[16152]_  = \new_[16151]_  & \new_[16146]_ ;
  assign \new_[16155]_  = ~A167 & ~A169;
  assign \new_[16159]_  = ~A200 & A199;
  assign \new_[16160]_  = ~A166 & \new_[16159]_ ;
  assign \new_[16161]_  = \new_[16160]_  & \new_[16155]_ ;
  assign \new_[16164]_  = A235 & A203;
  assign \new_[16168]_  = ~A301 & ~A299;
  assign \new_[16169]_  = ~A298 & \new_[16168]_ ;
  assign \new_[16170]_  = \new_[16169]_  & \new_[16164]_ ;
  assign \new_[16173]_  = ~A167 & ~A169;
  assign \new_[16177]_  = ~A200 & A199;
  assign \new_[16178]_  = ~A166 & \new_[16177]_ ;
  assign \new_[16179]_  = \new_[16178]_  & \new_[16173]_ ;
  assign \new_[16182]_  = A235 & A203;
  assign \new_[16186]_  = A269 & A266;
  assign \new_[16187]_  = ~A265 & \new_[16186]_ ;
  assign \new_[16188]_  = \new_[16187]_  & \new_[16182]_ ;
  assign \new_[16191]_  = ~A167 & ~A169;
  assign \new_[16195]_  = ~A200 & A199;
  assign \new_[16196]_  = ~A166 & \new_[16195]_ ;
  assign \new_[16197]_  = \new_[16196]_  & \new_[16191]_ ;
  assign \new_[16200]_  = A235 & A203;
  assign \new_[16204]_  = A269 & ~A266;
  assign \new_[16205]_  = A265 & \new_[16204]_ ;
  assign \new_[16206]_  = \new_[16205]_  & \new_[16200]_ ;
  assign \new_[16209]_  = ~A167 & ~A169;
  assign \new_[16213]_  = ~A200 & A199;
  assign \new_[16214]_  = ~A166 & \new_[16213]_ ;
  assign \new_[16215]_  = \new_[16214]_  & \new_[16209]_ ;
  assign \new_[16218]_  = A232 & A203;
  assign \new_[16222]_  = A267 & A265;
  assign \new_[16223]_  = A234 & \new_[16222]_ ;
  assign \new_[16224]_  = \new_[16223]_  & \new_[16218]_ ;
  assign \new_[16227]_  = ~A167 & ~A169;
  assign \new_[16231]_  = ~A200 & A199;
  assign \new_[16232]_  = ~A166 & \new_[16231]_ ;
  assign \new_[16233]_  = \new_[16232]_  & \new_[16227]_ ;
  assign \new_[16236]_  = A232 & A203;
  assign \new_[16240]_  = A267 & A266;
  assign \new_[16241]_  = A234 & \new_[16240]_ ;
  assign \new_[16242]_  = \new_[16241]_  & \new_[16236]_ ;
  assign \new_[16245]_  = ~A167 & ~A169;
  assign \new_[16249]_  = ~A200 & A199;
  assign \new_[16250]_  = ~A166 & \new_[16249]_ ;
  assign \new_[16251]_  = \new_[16250]_  & \new_[16245]_ ;
  assign \new_[16254]_  = A233 & A203;
  assign \new_[16258]_  = A267 & A265;
  assign \new_[16259]_  = A234 & \new_[16258]_ ;
  assign \new_[16260]_  = \new_[16259]_  & \new_[16254]_ ;
  assign \new_[16263]_  = ~A167 & ~A169;
  assign \new_[16267]_  = ~A200 & A199;
  assign \new_[16268]_  = ~A166 & \new_[16267]_ ;
  assign \new_[16269]_  = \new_[16268]_  & \new_[16263]_ ;
  assign \new_[16272]_  = A233 & A203;
  assign \new_[16276]_  = A267 & A266;
  assign \new_[16277]_  = A234 & \new_[16276]_ ;
  assign \new_[16278]_  = \new_[16277]_  & \new_[16272]_ ;
  assign \new_[16281]_  = ~A167 & ~A169;
  assign \new_[16285]_  = ~A200 & A199;
  assign \new_[16286]_  = ~A166 & \new_[16285]_ ;
  assign \new_[16287]_  = \new_[16286]_  & \new_[16281]_ ;
  assign \new_[16290]_  = ~A232 & A203;
  assign \new_[16294]_  = A268 & A236;
  assign \new_[16295]_  = A233 & \new_[16294]_ ;
  assign \new_[16296]_  = \new_[16295]_  & \new_[16290]_ ;
  assign \new_[16299]_  = ~A167 & ~A169;
  assign \new_[16303]_  = ~A200 & A199;
  assign \new_[16304]_  = ~A166 & \new_[16303]_ ;
  assign \new_[16305]_  = \new_[16304]_  & \new_[16299]_ ;
  assign \new_[16308]_  = A232 & A203;
  assign \new_[16312]_  = A268 & A236;
  assign \new_[16313]_  = ~A233 & \new_[16312]_ ;
  assign \new_[16314]_  = \new_[16313]_  & \new_[16308]_ ;
  assign \new_[16317]_  = ~A168 & ~A169;
  assign \new_[16321]_  = A202 & A166;
  assign \new_[16322]_  = A167 & \new_[16321]_ ;
  assign \new_[16323]_  = \new_[16322]_  & \new_[16317]_ ;
  assign \new_[16326]_  = A298 & A235;
  assign \new_[16330]_  = ~A301 & ~A300;
  assign \new_[16331]_  = A299 & \new_[16330]_ ;
  assign \new_[16332]_  = \new_[16331]_  & \new_[16326]_ ;
  assign \new_[16335]_  = ~A168 & ~A169;
  assign \new_[16339]_  = A202 & A166;
  assign \new_[16340]_  = A167 & \new_[16339]_ ;
  assign \new_[16341]_  = \new_[16340]_  & \new_[16335]_ ;
  assign \new_[16344]_  = A234 & A232;
  assign \new_[16348]_  = ~A302 & ~A301;
  assign \new_[16349]_  = ~A300 & \new_[16348]_ ;
  assign \new_[16350]_  = \new_[16349]_  & \new_[16344]_ ;
  assign \new_[16353]_  = ~A168 & ~A169;
  assign \new_[16357]_  = A202 & A166;
  assign \new_[16358]_  = A167 & \new_[16357]_ ;
  assign \new_[16359]_  = \new_[16358]_  & \new_[16353]_ ;
  assign \new_[16362]_  = A234 & A232;
  assign \new_[16366]_  = ~A301 & ~A299;
  assign \new_[16367]_  = ~A298 & \new_[16366]_ ;
  assign \new_[16368]_  = \new_[16367]_  & \new_[16362]_ ;
  assign \new_[16371]_  = ~A168 & ~A169;
  assign \new_[16375]_  = A202 & A166;
  assign \new_[16376]_  = A167 & \new_[16375]_ ;
  assign \new_[16377]_  = \new_[16376]_  & \new_[16371]_ ;
  assign \new_[16380]_  = A234 & A232;
  assign \new_[16384]_  = A269 & A266;
  assign \new_[16385]_  = ~A265 & \new_[16384]_ ;
  assign \new_[16386]_  = \new_[16385]_  & \new_[16380]_ ;
  assign \new_[16389]_  = ~A168 & ~A169;
  assign \new_[16393]_  = A202 & A166;
  assign \new_[16394]_  = A167 & \new_[16393]_ ;
  assign \new_[16395]_  = \new_[16394]_  & \new_[16389]_ ;
  assign \new_[16398]_  = A234 & A232;
  assign \new_[16402]_  = A269 & ~A266;
  assign \new_[16403]_  = A265 & \new_[16402]_ ;
  assign \new_[16404]_  = \new_[16403]_  & \new_[16398]_ ;
  assign \new_[16407]_  = ~A168 & ~A169;
  assign \new_[16411]_  = A202 & A166;
  assign \new_[16412]_  = A167 & \new_[16411]_ ;
  assign \new_[16413]_  = \new_[16412]_  & \new_[16407]_ ;
  assign \new_[16416]_  = A234 & A233;
  assign \new_[16420]_  = ~A302 & ~A301;
  assign \new_[16421]_  = ~A300 & \new_[16420]_ ;
  assign \new_[16422]_  = \new_[16421]_  & \new_[16416]_ ;
  assign \new_[16425]_  = ~A168 & ~A169;
  assign \new_[16429]_  = A202 & A166;
  assign \new_[16430]_  = A167 & \new_[16429]_ ;
  assign \new_[16431]_  = \new_[16430]_  & \new_[16425]_ ;
  assign \new_[16434]_  = A234 & A233;
  assign \new_[16438]_  = ~A301 & ~A299;
  assign \new_[16439]_  = ~A298 & \new_[16438]_ ;
  assign \new_[16440]_  = \new_[16439]_  & \new_[16434]_ ;
  assign \new_[16443]_  = ~A168 & ~A169;
  assign \new_[16447]_  = A202 & A166;
  assign \new_[16448]_  = A167 & \new_[16447]_ ;
  assign \new_[16449]_  = \new_[16448]_  & \new_[16443]_ ;
  assign \new_[16452]_  = A234 & A233;
  assign \new_[16456]_  = A269 & A266;
  assign \new_[16457]_  = ~A265 & \new_[16456]_ ;
  assign \new_[16458]_  = \new_[16457]_  & \new_[16452]_ ;
  assign \new_[16461]_  = ~A168 & ~A169;
  assign \new_[16465]_  = A202 & A166;
  assign \new_[16466]_  = A167 & \new_[16465]_ ;
  assign \new_[16467]_  = \new_[16466]_  & \new_[16461]_ ;
  assign \new_[16470]_  = A234 & A233;
  assign \new_[16474]_  = A269 & ~A266;
  assign \new_[16475]_  = A265 & \new_[16474]_ ;
  assign \new_[16476]_  = \new_[16475]_  & \new_[16470]_ ;
  assign \new_[16479]_  = ~A168 & ~A169;
  assign \new_[16483]_  = A202 & A166;
  assign \new_[16484]_  = A167 & \new_[16483]_ ;
  assign \new_[16485]_  = \new_[16484]_  & \new_[16479]_ ;
  assign \new_[16488]_  = A233 & ~A232;
  assign \new_[16492]_  = A267 & A265;
  assign \new_[16493]_  = A236 & \new_[16492]_ ;
  assign \new_[16494]_  = \new_[16493]_  & \new_[16488]_ ;
  assign \new_[16497]_  = ~A168 & ~A169;
  assign \new_[16501]_  = A202 & A166;
  assign \new_[16502]_  = A167 & \new_[16501]_ ;
  assign \new_[16503]_  = \new_[16502]_  & \new_[16497]_ ;
  assign \new_[16506]_  = A233 & ~A232;
  assign \new_[16510]_  = A267 & A266;
  assign \new_[16511]_  = A236 & \new_[16510]_ ;
  assign \new_[16512]_  = \new_[16511]_  & \new_[16506]_ ;
  assign \new_[16515]_  = ~A168 & ~A169;
  assign \new_[16519]_  = A202 & A166;
  assign \new_[16520]_  = A167 & \new_[16519]_ ;
  assign \new_[16521]_  = \new_[16520]_  & \new_[16515]_ ;
  assign \new_[16524]_  = ~A233 & A232;
  assign \new_[16528]_  = A267 & A265;
  assign \new_[16529]_  = A236 & \new_[16528]_ ;
  assign \new_[16530]_  = \new_[16529]_  & \new_[16524]_ ;
  assign \new_[16533]_  = ~A168 & ~A169;
  assign \new_[16537]_  = A202 & A166;
  assign \new_[16538]_  = A167 & \new_[16537]_ ;
  assign \new_[16539]_  = \new_[16538]_  & \new_[16533]_ ;
  assign \new_[16542]_  = ~A233 & A232;
  assign \new_[16546]_  = A267 & A266;
  assign \new_[16547]_  = A236 & \new_[16546]_ ;
  assign \new_[16548]_  = \new_[16547]_  & \new_[16542]_ ;
  assign \new_[16551]_  = ~A168 & ~A169;
  assign \new_[16555]_  = A199 & A166;
  assign \new_[16556]_  = A167 & \new_[16555]_ ;
  assign \new_[16557]_  = \new_[16556]_  & \new_[16551]_ ;
  assign \new_[16560]_  = A235 & A201;
  assign \new_[16564]_  = ~A302 & ~A301;
  assign \new_[16565]_  = ~A300 & \new_[16564]_ ;
  assign \new_[16566]_  = \new_[16565]_  & \new_[16560]_ ;
  assign \new_[16569]_  = ~A168 & ~A169;
  assign \new_[16573]_  = A199 & A166;
  assign \new_[16574]_  = A167 & \new_[16573]_ ;
  assign \new_[16575]_  = \new_[16574]_  & \new_[16569]_ ;
  assign \new_[16578]_  = A235 & A201;
  assign \new_[16582]_  = ~A301 & ~A299;
  assign \new_[16583]_  = ~A298 & \new_[16582]_ ;
  assign \new_[16584]_  = \new_[16583]_  & \new_[16578]_ ;
  assign \new_[16587]_  = ~A168 & ~A169;
  assign \new_[16591]_  = A199 & A166;
  assign \new_[16592]_  = A167 & \new_[16591]_ ;
  assign \new_[16593]_  = \new_[16592]_  & \new_[16587]_ ;
  assign \new_[16596]_  = A235 & A201;
  assign \new_[16600]_  = A269 & A266;
  assign \new_[16601]_  = ~A265 & \new_[16600]_ ;
  assign \new_[16602]_  = \new_[16601]_  & \new_[16596]_ ;
  assign \new_[16605]_  = ~A168 & ~A169;
  assign \new_[16609]_  = A199 & A166;
  assign \new_[16610]_  = A167 & \new_[16609]_ ;
  assign \new_[16611]_  = \new_[16610]_  & \new_[16605]_ ;
  assign \new_[16614]_  = A235 & A201;
  assign \new_[16618]_  = A269 & ~A266;
  assign \new_[16619]_  = A265 & \new_[16618]_ ;
  assign \new_[16620]_  = \new_[16619]_  & \new_[16614]_ ;
  assign \new_[16623]_  = ~A168 & ~A169;
  assign \new_[16627]_  = A199 & A166;
  assign \new_[16628]_  = A167 & \new_[16627]_ ;
  assign \new_[16629]_  = \new_[16628]_  & \new_[16623]_ ;
  assign \new_[16632]_  = A232 & A201;
  assign \new_[16636]_  = A267 & A265;
  assign \new_[16637]_  = A234 & \new_[16636]_ ;
  assign \new_[16638]_  = \new_[16637]_  & \new_[16632]_ ;
  assign \new_[16641]_  = ~A168 & ~A169;
  assign \new_[16645]_  = A199 & A166;
  assign \new_[16646]_  = A167 & \new_[16645]_ ;
  assign \new_[16647]_  = \new_[16646]_  & \new_[16641]_ ;
  assign \new_[16650]_  = A232 & A201;
  assign \new_[16654]_  = A267 & A266;
  assign \new_[16655]_  = A234 & \new_[16654]_ ;
  assign \new_[16656]_  = \new_[16655]_  & \new_[16650]_ ;
  assign \new_[16659]_  = ~A168 & ~A169;
  assign \new_[16663]_  = A199 & A166;
  assign \new_[16664]_  = A167 & \new_[16663]_ ;
  assign \new_[16665]_  = \new_[16664]_  & \new_[16659]_ ;
  assign \new_[16668]_  = A233 & A201;
  assign \new_[16672]_  = A267 & A265;
  assign \new_[16673]_  = A234 & \new_[16672]_ ;
  assign \new_[16674]_  = \new_[16673]_  & \new_[16668]_ ;
  assign \new_[16677]_  = ~A168 & ~A169;
  assign \new_[16681]_  = A199 & A166;
  assign \new_[16682]_  = A167 & \new_[16681]_ ;
  assign \new_[16683]_  = \new_[16682]_  & \new_[16677]_ ;
  assign \new_[16686]_  = A233 & A201;
  assign \new_[16690]_  = A267 & A266;
  assign \new_[16691]_  = A234 & \new_[16690]_ ;
  assign \new_[16692]_  = \new_[16691]_  & \new_[16686]_ ;
  assign \new_[16695]_  = ~A168 & ~A169;
  assign \new_[16699]_  = A199 & A166;
  assign \new_[16700]_  = A167 & \new_[16699]_ ;
  assign \new_[16701]_  = \new_[16700]_  & \new_[16695]_ ;
  assign \new_[16704]_  = ~A232 & A201;
  assign \new_[16708]_  = A268 & A236;
  assign \new_[16709]_  = A233 & \new_[16708]_ ;
  assign \new_[16710]_  = \new_[16709]_  & \new_[16704]_ ;
  assign \new_[16713]_  = ~A168 & ~A169;
  assign \new_[16717]_  = A199 & A166;
  assign \new_[16718]_  = A167 & \new_[16717]_ ;
  assign \new_[16719]_  = \new_[16718]_  & \new_[16713]_ ;
  assign \new_[16722]_  = A232 & A201;
  assign \new_[16726]_  = A268 & A236;
  assign \new_[16727]_  = ~A233 & \new_[16726]_ ;
  assign \new_[16728]_  = \new_[16727]_  & \new_[16722]_ ;
  assign \new_[16731]_  = ~A168 & ~A169;
  assign \new_[16735]_  = A200 & A166;
  assign \new_[16736]_  = A167 & \new_[16735]_ ;
  assign \new_[16737]_  = \new_[16736]_  & \new_[16731]_ ;
  assign \new_[16740]_  = A235 & A201;
  assign \new_[16744]_  = ~A302 & ~A301;
  assign \new_[16745]_  = ~A300 & \new_[16744]_ ;
  assign \new_[16746]_  = \new_[16745]_  & \new_[16740]_ ;
  assign \new_[16749]_  = ~A168 & ~A169;
  assign \new_[16753]_  = A200 & A166;
  assign \new_[16754]_  = A167 & \new_[16753]_ ;
  assign \new_[16755]_  = \new_[16754]_  & \new_[16749]_ ;
  assign \new_[16758]_  = A235 & A201;
  assign \new_[16762]_  = ~A301 & ~A299;
  assign \new_[16763]_  = ~A298 & \new_[16762]_ ;
  assign \new_[16764]_  = \new_[16763]_  & \new_[16758]_ ;
  assign \new_[16767]_  = ~A168 & ~A169;
  assign \new_[16771]_  = A200 & A166;
  assign \new_[16772]_  = A167 & \new_[16771]_ ;
  assign \new_[16773]_  = \new_[16772]_  & \new_[16767]_ ;
  assign \new_[16776]_  = A235 & A201;
  assign \new_[16780]_  = A269 & A266;
  assign \new_[16781]_  = ~A265 & \new_[16780]_ ;
  assign \new_[16782]_  = \new_[16781]_  & \new_[16776]_ ;
  assign \new_[16785]_  = ~A168 & ~A169;
  assign \new_[16789]_  = A200 & A166;
  assign \new_[16790]_  = A167 & \new_[16789]_ ;
  assign \new_[16791]_  = \new_[16790]_  & \new_[16785]_ ;
  assign \new_[16794]_  = A235 & A201;
  assign \new_[16798]_  = A269 & ~A266;
  assign \new_[16799]_  = A265 & \new_[16798]_ ;
  assign \new_[16800]_  = \new_[16799]_  & \new_[16794]_ ;
  assign \new_[16803]_  = ~A168 & ~A169;
  assign \new_[16807]_  = A200 & A166;
  assign \new_[16808]_  = A167 & \new_[16807]_ ;
  assign \new_[16809]_  = \new_[16808]_  & \new_[16803]_ ;
  assign \new_[16812]_  = A232 & A201;
  assign \new_[16816]_  = A267 & A265;
  assign \new_[16817]_  = A234 & \new_[16816]_ ;
  assign \new_[16818]_  = \new_[16817]_  & \new_[16812]_ ;
  assign \new_[16821]_  = ~A168 & ~A169;
  assign \new_[16825]_  = A200 & A166;
  assign \new_[16826]_  = A167 & \new_[16825]_ ;
  assign \new_[16827]_  = \new_[16826]_  & \new_[16821]_ ;
  assign \new_[16830]_  = A232 & A201;
  assign \new_[16834]_  = A267 & A266;
  assign \new_[16835]_  = A234 & \new_[16834]_ ;
  assign \new_[16836]_  = \new_[16835]_  & \new_[16830]_ ;
  assign \new_[16839]_  = ~A168 & ~A169;
  assign \new_[16843]_  = A200 & A166;
  assign \new_[16844]_  = A167 & \new_[16843]_ ;
  assign \new_[16845]_  = \new_[16844]_  & \new_[16839]_ ;
  assign \new_[16848]_  = A233 & A201;
  assign \new_[16852]_  = A267 & A265;
  assign \new_[16853]_  = A234 & \new_[16852]_ ;
  assign \new_[16854]_  = \new_[16853]_  & \new_[16848]_ ;
  assign \new_[16857]_  = ~A168 & ~A169;
  assign \new_[16861]_  = A200 & A166;
  assign \new_[16862]_  = A167 & \new_[16861]_ ;
  assign \new_[16863]_  = \new_[16862]_  & \new_[16857]_ ;
  assign \new_[16866]_  = A233 & A201;
  assign \new_[16870]_  = A267 & A266;
  assign \new_[16871]_  = A234 & \new_[16870]_ ;
  assign \new_[16872]_  = \new_[16871]_  & \new_[16866]_ ;
  assign \new_[16875]_  = ~A168 & ~A169;
  assign \new_[16879]_  = A200 & A166;
  assign \new_[16880]_  = A167 & \new_[16879]_ ;
  assign \new_[16881]_  = \new_[16880]_  & \new_[16875]_ ;
  assign \new_[16884]_  = ~A232 & A201;
  assign \new_[16888]_  = A268 & A236;
  assign \new_[16889]_  = A233 & \new_[16888]_ ;
  assign \new_[16890]_  = \new_[16889]_  & \new_[16884]_ ;
  assign \new_[16893]_  = ~A168 & ~A169;
  assign \new_[16897]_  = A200 & A166;
  assign \new_[16898]_  = A167 & \new_[16897]_ ;
  assign \new_[16899]_  = \new_[16898]_  & \new_[16893]_ ;
  assign \new_[16902]_  = A232 & A201;
  assign \new_[16906]_  = A268 & A236;
  assign \new_[16907]_  = ~A233 & \new_[16906]_ ;
  assign \new_[16908]_  = \new_[16907]_  & \new_[16902]_ ;
  assign \new_[16911]_  = ~A168 & ~A169;
  assign \new_[16915]_  = ~A199 & A166;
  assign \new_[16916]_  = A167 & \new_[16915]_ ;
  assign \new_[16917]_  = \new_[16916]_  & \new_[16911]_ ;
  assign \new_[16920]_  = A203 & A200;
  assign \new_[16924]_  = A267 & A265;
  assign \new_[16925]_  = A235 & \new_[16924]_ ;
  assign \new_[16926]_  = \new_[16925]_  & \new_[16920]_ ;
  assign \new_[16929]_  = ~A168 & ~A169;
  assign \new_[16933]_  = ~A199 & A166;
  assign \new_[16934]_  = A167 & \new_[16933]_ ;
  assign \new_[16935]_  = \new_[16934]_  & \new_[16929]_ ;
  assign \new_[16938]_  = A203 & A200;
  assign \new_[16942]_  = A267 & A266;
  assign \new_[16943]_  = A235 & \new_[16942]_ ;
  assign \new_[16944]_  = \new_[16943]_  & \new_[16938]_ ;
  assign \new_[16947]_  = ~A168 & ~A169;
  assign \new_[16951]_  = ~A199 & A166;
  assign \new_[16952]_  = A167 & \new_[16951]_ ;
  assign \new_[16953]_  = \new_[16952]_  & \new_[16947]_ ;
  assign \new_[16956]_  = A203 & A200;
  assign \new_[16960]_  = A268 & A234;
  assign \new_[16961]_  = A232 & \new_[16960]_ ;
  assign \new_[16962]_  = \new_[16961]_  & \new_[16956]_ ;
  assign \new_[16965]_  = ~A168 & ~A169;
  assign \new_[16969]_  = ~A199 & A166;
  assign \new_[16970]_  = A167 & \new_[16969]_ ;
  assign \new_[16971]_  = \new_[16970]_  & \new_[16965]_ ;
  assign \new_[16974]_  = A203 & A200;
  assign \new_[16978]_  = A268 & A234;
  assign \new_[16979]_  = A233 & \new_[16978]_ ;
  assign \new_[16980]_  = \new_[16979]_  & \new_[16974]_ ;
  assign \new_[16983]_  = ~A168 & ~A169;
  assign \new_[16987]_  = A199 & A166;
  assign \new_[16988]_  = A167 & \new_[16987]_ ;
  assign \new_[16989]_  = \new_[16988]_  & \new_[16983]_ ;
  assign \new_[16992]_  = A203 & ~A200;
  assign \new_[16996]_  = A267 & A265;
  assign \new_[16997]_  = A235 & \new_[16996]_ ;
  assign \new_[16998]_  = \new_[16997]_  & \new_[16992]_ ;
  assign \new_[17001]_  = ~A168 & ~A169;
  assign \new_[17005]_  = A199 & A166;
  assign \new_[17006]_  = A167 & \new_[17005]_ ;
  assign \new_[17007]_  = \new_[17006]_  & \new_[17001]_ ;
  assign \new_[17010]_  = A203 & ~A200;
  assign \new_[17014]_  = A267 & A266;
  assign \new_[17015]_  = A235 & \new_[17014]_ ;
  assign \new_[17016]_  = \new_[17015]_  & \new_[17010]_ ;
  assign \new_[17019]_  = ~A168 & ~A169;
  assign \new_[17023]_  = A199 & A166;
  assign \new_[17024]_  = A167 & \new_[17023]_ ;
  assign \new_[17025]_  = \new_[17024]_  & \new_[17019]_ ;
  assign \new_[17028]_  = A203 & ~A200;
  assign \new_[17032]_  = A268 & A234;
  assign \new_[17033]_  = A232 & \new_[17032]_ ;
  assign \new_[17034]_  = \new_[17033]_  & \new_[17028]_ ;
  assign \new_[17037]_  = ~A168 & ~A169;
  assign \new_[17041]_  = A199 & A166;
  assign \new_[17042]_  = A167 & \new_[17041]_ ;
  assign \new_[17043]_  = \new_[17042]_  & \new_[17037]_ ;
  assign \new_[17046]_  = A203 & ~A200;
  assign \new_[17050]_  = A268 & A234;
  assign \new_[17051]_  = A233 & \new_[17050]_ ;
  assign \new_[17052]_  = \new_[17051]_  & \new_[17046]_ ;
  assign \new_[17055]_  = ~A169 & ~A170;
  assign \new_[17059]_  = A232 & A202;
  assign \new_[17060]_  = ~A168 & \new_[17059]_ ;
  assign \new_[17061]_  = \new_[17060]_  & \new_[17055]_ ;
  assign \new_[17064]_  = A298 & A234;
  assign \new_[17068]_  = ~A301 & ~A300;
  assign \new_[17069]_  = A299 & \new_[17068]_ ;
  assign \new_[17070]_  = \new_[17069]_  & \new_[17064]_ ;
  assign \new_[17073]_  = ~A169 & ~A170;
  assign \new_[17077]_  = A233 & A202;
  assign \new_[17078]_  = ~A168 & \new_[17077]_ ;
  assign \new_[17079]_  = \new_[17078]_  & \new_[17073]_ ;
  assign \new_[17082]_  = A298 & A234;
  assign \new_[17086]_  = ~A301 & ~A300;
  assign \new_[17087]_  = A299 & \new_[17086]_ ;
  assign \new_[17088]_  = \new_[17087]_  & \new_[17082]_ ;
  assign \new_[17091]_  = ~A169 & ~A170;
  assign \new_[17095]_  = ~A232 & A202;
  assign \new_[17096]_  = ~A168 & \new_[17095]_ ;
  assign \new_[17097]_  = \new_[17096]_  & \new_[17091]_ ;
  assign \new_[17100]_  = A236 & A233;
  assign \new_[17104]_  = ~A302 & ~A301;
  assign \new_[17105]_  = ~A300 & \new_[17104]_ ;
  assign \new_[17106]_  = \new_[17105]_  & \new_[17100]_ ;
  assign \new_[17109]_  = ~A169 & ~A170;
  assign \new_[17113]_  = ~A232 & A202;
  assign \new_[17114]_  = ~A168 & \new_[17113]_ ;
  assign \new_[17115]_  = \new_[17114]_  & \new_[17109]_ ;
  assign \new_[17118]_  = A236 & A233;
  assign \new_[17122]_  = ~A301 & ~A299;
  assign \new_[17123]_  = ~A298 & \new_[17122]_ ;
  assign \new_[17124]_  = \new_[17123]_  & \new_[17118]_ ;
  assign \new_[17127]_  = ~A169 & ~A170;
  assign \new_[17131]_  = ~A232 & A202;
  assign \new_[17132]_  = ~A168 & \new_[17131]_ ;
  assign \new_[17133]_  = \new_[17132]_  & \new_[17127]_ ;
  assign \new_[17136]_  = A236 & A233;
  assign \new_[17140]_  = A269 & A266;
  assign \new_[17141]_  = ~A265 & \new_[17140]_ ;
  assign \new_[17142]_  = \new_[17141]_  & \new_[17136]_ ;
  assign \new_[17145]_  = ~A169 & ~A170;
  assign \new_[17149]_  = ~A232 & A202;
  assign \new_[17150]_  = ~A168 & \new_[17149]_ ;
  assign \new_[17151]_  = \new_[17150]_  & \new_[17145]_ ;
  assign \new_[17154]_  = A236 & A233;
  assign \new_[17158]_  = A269 & ~A266;
  assign \new_[17159]_  = A265 & \new_[17158]_ ;
  assign \new_[17160]_  = \new_[17159]_  & \new_[17154]_ ;
  assign \new_[17163]_  = ~A169 & ~A170;
  assign \new_[17167]_  = A232 & A202;
  assign \new_[17168]_  = ~A168 & \new_[17167]_ ;
  assign \new_[17169]_  = \new_[17168]_  & \new_[17163]_ ;
  assign \new_[17172]_  = A236 & ~A233;
  assign \new_[17176]_  = ~A302 & ~A301;
  assign \new_[17177]_  = ~A300 & \new_[17176]_ ;
  assign \new_[17178]_  = \new_[17177]_  & \new_[17172]_ ;
  assign \new_[17181]_  = ~A169 & ~A170;
  assign \new_[17185]_  = A232 & A202;
  assign \new_[17186]_  = ~A168 & \new_[17185]_ ;
  assign \new_[17187]_  = \new_[17186]_  & \new_[17181]_ ;
  assign \new_[17190]_  = A236 & ~A233;
  assign \new_[17194]_  = ~A301 & ~A299;
  assign \new_[17195]_  = ~A298 & \new_[17194]_ ;
  assign \new_[17196]_  = \new_[17195]_  & \new_[17190]_ ;
  assign \new_[17199]_  = ~A169 & ~A170;
  assign \new_[17203]_  = A232 & A202;
  assign \new_[17204]_  = ~A168 & \new_[17203]_ ;
  assign \new_[17205]_  = \new_[17204]_  & \new_[17199]_ ;
  assign \new_[17208]_  = A236 & ~A233;
  assign \new_[17212]_  = A269 & A266;
  assign \new_[17213]_  = ~A265 & \new_[17212]_ ;
  assign \new_[17214]_  = \new_[17213]_  & \new_[17208]_ ;
  assign \new_[17217]_  = ~A169 & ~A170;
  assign \new_[17221]_  = A232 & A202;
  assign \new_[17222]_  = ~A168 & \new_[17221]_ ;
  assign \new_[17223]_  = \new_[17222]_  & \new_[17217]_ ;
  assign \new_[17226]_  = A236 & ~A233;
  assign \new_[17230]_  = A269 & ~A266;
  assign \new_[17231]_  = A265 & \new_[17230]_ ;
  assign \new_[17232]_  = \new_[17231]_  & \new_[17226]_ ;
  assign \new_[17235]_  = ~A169 & ~A170;
  assign \new_[17239]_  = A201 & A199;
  assign \new_[17240]_  = ~A168 & \new_[17239]_ ;
  assign \new_[17241]_  = \new_[17240]_  & \new_[17235]_ ;
  assign \new_[17244]_  = A298 & A235;
  assign \new_[17248]_  = ~A301 & ~A300;
  assign \new_[17249]_  = A299 & \new_[17248]_ ;
  assign \new_[17250]_  = \new_[17249]_  & \new_[17244]_ ;
  assign \new_[17253]_  = ~A169 & ~A170;
  assign \new_[17257]_  = A201 & A199;
  assign \new_[17258]_  = ~A168 & \new_[17257]_ ;
  assign \new_[17259]_  = \new_[17258]_  & \new_[17253]_ ;
  assign \new_[17262]_  = A234 & A232;
  assign \new_[17266]_  = ~A302 & ~A301;
  assign \new_[17267]_  = ~A300 & \new_[17266]_ ;
  assign \new_[17268]_  = \new_[17267]_  & \new_[17262]_ ;
  assign \new_[17271]_  = ~A169 & ~A170;
  assign \new_[17275]_  = A201 & A199;
  assign \new_[17276]_  = ~A168 & \new_[17275]_ ;
  assign \new_[17277]_  = \new_[17276]_  & \new_[17271]_ ;
  assign \new_[17280]_  = A234 & A232;
  assign \new_[17284]_  = ~A301 & ~A299;
  assign \new_[17285]_  = ~A298 & \new_[17284]_ ;
  assign \new_[17286]_  = \new_[17285]_  & \new_[17280]_ ;
  assign \new_[17289]_  = ~A169 & ~A170;
  assign \new_[17293]_  = A201 & A199;
  assign \new_[17294]_  = ~A168 & \new_[17293]_ ;
  assign \new_[17295]_  = \new_[17294]_  & \new_[17289]_ ;
  assign \new_[17298]_  = A234 & A232;
  assign \new_[17302]_  = A269 & A266;
  assign \new_[17303]_  = ~A265 & \new_[17302]_ ;
  assign \new_[17304]_  = \new_[17303]_  & \new_[17298]_ ;
  assign \new_[17307]_  = ~A169 & ~A170;
  assign \new_[17311]_  = A201 & A199;
  assign \new_[17312]_  = ~A168 & \new_[17311]_ ;
  assign \new_[17313]_  = \new_[17312]_  & \new_[17307]_ ;
  assign \new_[17316]_  = A234 & A232;
  assign \new_[17320]_  = A269 & ~A266;
  assign \new_[17321]_  = A265 & \new_[17320]_ ;
  assign \new_[17322]_  = \new_[17321]_  & \new_[17316]_ ;
  assign \new_[17325]_  = ~A169 & ~A170;
  assign \new_[17329]_  = A201 & A199;
  assign \new_[17330]_  = ~A168 & \new_[17329]_ ;
  assign \new_[17331]_  = \new_[17330]_  & \new_[17325]_ ;
  assign \new_[17334]_  = A234 & A233;
  assign \new_[17338]_  = ~A302 & ~A301;
  assign \new_[17339]_  = ~A300 & \new_[17338]_ ;
  assign \new_[17340]_  = \new_[17339]_  & \new_[17334]_ ;
  assign \new_[17343]_  = ~A169 & ~A170;
  assign \new_[17347]_  = A201 & A199;
  assign \new_[17348]_  = ~A168 & \new_[17347]_ ;
  assign \new_[17349]_  = \new_[17348]_  & \new_[17343]_ ;
  assign \new_[17352]_  = A234 & A233;
  assign \new_[17356]_  = ~A301 & ~A299;
  assign \new_[17357]_  = ~A298 & \new_[17356]_ ;
  assign \new_[17358]_  = \new_[17357]_  & \new_[17352]_ ;
  assign \new_[17361]_  = ~A169 & ~A170;
  assign \new_[17365]_  = A201 & A199;
  assign \new_[17366]_  = ~A168 & \new_[17365]_ ;
  assign \new_[17367]_  = \new_[17366]_  & \new_[17361]_ ;
  assign \new_[17370]_  = A234 & A233;
  assign \new_[17374]_  = A269 & A266;
  assign \new_[17375]_  = ~A265 & \new_[17374]_ ;
  assign \new_[17376]_  = \new_[17375]_  & \new_[17370]_ ;
  assign \new_[17379]_  = ~A169 & ~A170;
  assign \new_[17383]_  = A201 & A199;
  assign \new_[17384]_  = ~A168 & \new_[17383]_ ;
  assign \new_[17385]_  = \new_[17384]_  & \new_[17379]_ ;
  assign \new_[17388]_  = A234 & A233;
  assign \new_[17392]_  = A269 & ~A266;
  assign \new_[17393]_  = A265 & \new_[17392]_ ;
  assign \new_[17394]_  = \new_[17393]_  & \new_[17388]_ ;
  assign \new_[17397]_  = ~A169 & ~A170;
  assign \new_[17401]_  = A201 & A199;
  assign \new_[17402]_  = ~A168 & \new_[17401]_ ;
  assign \new_[17403]_  = \new_[17402]_  & \new_[17397]_ ;
  assign \new_[17406]_  = A233 & ~A232;
  assign \new_[17410]_  = A267 & A265;
  assign \new_[17411]_  = A236 & \new_[17410]_ ;
  assign \new_[17412]_  = \new_[17411]_  & \new_[17406]_ ;
  assign \new_[17415]_  = ~A169 & ~A170;
  assign \new_[17419]_  = A201 & A199;
  assign \new_[17420]_  = ~A168 & \new_[17419]_ ;
  assign \new_[17421]_  = \new_[17420]_  & \new_[17415]_ ;
  assign \new_[17424]_  = A233 & ~A232;
  assign \new_[17428]_  = A267 & A266;
  assign \new_[17429]_  = A236 & \new_[17428]_ ;
  assign \new_[17430]_  = \new_[17429]_  & \new_[17424]_ ;
  assign \new_[17433]_  = ~A169 & ~A170;
  assign \new_[17437]_  = A201 & A199;
  assign \new_[17438]_  = ~A168 & \new_[17437]_ ;
  assign \new_[17439]_  = \new_[17438]_  & \new_[17433]_ ;
  assign \new_[17442]_  = ~A233 & A232;
  assign \new_[17446]_  = A267 & A265;
  assign \new_[17447]_  = A236 & \new_[17446]_ ;
  assign \new_[17448]_  = \new_[17447]_  & \new_[17442]_ ;
  assign \new_[17451]_  = ~A169 & ~A170;
  assign \new_[17455]_  = A201 & A199;
  assign \new_[17456]_  = ~A168 & \new_[17455]_ ;
  assign \new_[17457]_  = \new_[17456]_  & \new_[17451]_ ;
  assign \new_[17460]_  = ~A233 & A232;
  assign \new_[17464]_  = A267 & A266;
  assign \new_[17465]_  = A236 & \new_[17464]_ ;
  assign \new_[17466]_  = \new_[17465]_  & \new_[17460]_ ;
  assign \new_[17469]_  = ~A169 & ~A170;
  assign \new_[17473]_  = A201 & A200;
  assign \new_[17474]_  = ~A168 & \new_[17473]_ ;
  assign \new_[17475]_  = \new_[17474]_  & \new_[17469]_ ;
  assign \new_[17478]_  = A298 & A235;
  assign \new_[17482]_  = ~A301 & ~A300;
  assign \new_[17483]_  = A299 & \new_[17482]_ ;
  assign \new_[17484]_  = \new_[17483]_  & \new_[17478]_ ;
  assign \new_[17487]_  = ~A169 & ~A170;
  assign \new_[17491]_  = A201 & A200;
  assign \new_[17492]_  = ~A168 & \new_[17491]_ ;
  assign \new_[17493]_  = \new_[17492]_  & \new_[17487]_ ;
  assign \new_[17496]_  = A234 & A232;
  assign \new_[17500]_  = ~A302 & ~A301;
  assign \new_[17501]_  = ~A300 & \new_[17500]_ ;
  assign \new_[17502]_  = \new_[17501]_  & \new_[17496]_ ;
  assign \new_[17505]_  = ~A169 & ~A170;
  assign \new_[17509]_  = A201 & A200;
  assign \new_[17510]_  = ~A168 & \new_[17509]_ ;
  assign \new_[17511]_  = \new_[17510]_  & \new_[17505]_ ;
  assign \new_[17514]_  = A234 & A232;
  assign \new_[17518]_  = ~A301 & ~A299;
  assign \new_[17519]_  = ~A298 & \new_[17518]_ ;
  assign \new_[17520]_  = \new_[17519]_  & \new_[17514]_ ;
  assign \new_[17523]_  = ~A169 & ~A170;
  assign \new_[17527]_  = A201 & A200;
  assign \new_[17528]_  = ~A168 & \new_[17527]_ ;
  assign \new_[17529]_  = \new_[17528]_  & \new_[17523]_ ;
  assign \new_[17532]_  = A234 & A232;
  assign \new_[17536]_  = A269 & A266;
  assign \new_[17537]_  = ~A265 & \new_[17536]_ ;
  assign \new_[17538]_  = \new_[17537]_  & \new_[17532]_ ;
  assign \new_[17541]_  = ~A169 & ~A170;
  assign \new_[17545]_  = A201 & A200;
  assign \new_[17546]_  = ~A168 & \new_[17545]_ ;
  assign \new_[17547]_  = \new_[17546]_  & \new_[17541]_ ;
  assign \new_[17550]_  = A234 & A232;
  assign \new_[17554]_  = A269 & ~A266;
  assign \new_[17555]_  = A265 & \new_[17554]_ ;
  assign \new_[17556]_  = \new_[17555]_  & \new_[17550]_ ;
  assign \new_[17559]_  = ~A169 & ~A170;
  assign \new_[17563]_  = A201 & A200;
  assign \new_[17564]_  = ~A168 & \new_[17563]_ ;
  assign \new_[17565]_  = \new_[17564]_  & \new_[17559]_ ;
  assign \new_[17568]_  = A234 & A233;
  assign \new_[17572]_  = ~A302 & ~A301;
  assign \new_[17573]_  = ~A300 & \new_[17572]_ ;
  assign \new_[17574]_  = \new_[17573]_  & \new_[17568]_ ;
  assign \new_[17577]_  = ~A169 & ~A170;
  assign \new_[17581]_  = A201 & A200;
  assign \new_[17582]_  = ~A168 & \new_[17581]_ ;
  assign \new_[17583]_  = \new_[17582]_  & \new_[17577]_ ;
  assign \new_[17586]_  = A234 & A233;
  assign \new_[17590]_  = ~A301 & ~A299;
  assign \new_[17591]_  = ~A298 & \new_[17590]_ ;
  assign \new_[17592]_  = \new_[17591]_  & \new_[17586]_ ;
  assign \new_[17595]_  = ~A169 & ~A170;
  assign \new_[17599]_  = A201 & A200;
  assign \new_[17600]_  = ~A168 & \new_[17599]_ ;
  assign \new_[17601]_  = \new_[17600]_  & \new_[17595]_ ;
  assign \new_[17604]_  = A234 & A233;
  assign \new_[17608]_  = A269 & A266;
  assign \new_[17609]_  = ~A265 & \new_[17608]_ ;
  assign \new_[17610]_  = \new_[17609]_  & \new_[17604]_ ;
  assign \new_[17613]_  = ~A169 & ~A170;
  assign \new_[17617]_  = A201 & A200;
  assign \new_[17618]_  = ~A168 & \new_[17617]_ ;
  assign \new_[17619]_  = \new_[17618]_  & \new_[17613]_ ;
  assign \new_[17622]_  = A234 & A233;
  assign \new_[17626]_  = A269 & ~A266;
  assign \new_[17627]_  = A265 & \new_[17626]_ ;
  assign \new_[17628]_  = \new_[17627]_  & \new_[17622]_ ;
  assign \new_[17631]_  = ~A169 & ~A170;
  assign \new_[17635]_  = A201 & A200;
  assign \new_[17636]_  = ~A168 & \new_[17635]_ ;
  assign \new_[17637]_  = \new_[17636]_  & \new_[17631]_ ;
  assign \new_[17640]_  = A233 & ~A232;
  assign \new_[17644]_  = A267 & A265;
  assign \new_[17645]_  = A236 & \new_[17644]_ ;
  assign \new_[17646]_  = \new_[17645]_  & \new_[17640]_ ;
  assign \new_[17649]_  = ~A169 & ~A170;
  assign \new_[17653]_  = A201 & A200;
  assign \new_[17654]_  = ~A168 & \new_[17653]_ ;
  assign \new_[17655]_  = \new_[17654]_  & \new_[17649]_ ;
  assign \new_[17658]_  = A233 & ~A232;
  assign \new_[17662]_  = A267 & A266;
  assign \new_[17663]_  = A236 & \new_[17662]_ ;
  assign \new_[17664]_  = \new_[17663]_  & \new_[17658]_ ;
  assign \new_[17667]_  = ~A169 & ~A170;
  assign \new_[17671]_  = A201 & A200;
  assign \new_[17672]_  = ~A168 & \new_[17671]_ ;
  assign \new_[17673]_  = \new_[17672]_  & \new_[17667]_ ;
  assign \new_[17676]_  = ~A233 & A232;
  assign \new_[17680]_  = A267 & A265;
  assign \new_[17681]_  = A236 & \new_[17680]_ ;
  assign \new_[17682]_  = \new_[17681]_  & \new_[17676]_ ;
  assign \new_[17685]_  = ~A169 & ~A170;
  assign \new_[17689]_  = A201 & A200;
  assign \new_[17690]_  = ~A168 & \new_[17689]_ ;
  assign \new_[17691]_  = \new_[17690]_  & \new_[17685]_ ;
  assign \new_[17694]_  = ~A233 & A232;
  assign \new_[17698]_  = A267 & A266;
  assign \new_[17699]_  = A236 & \new_[17698]_ ;
  assign \new_[17700]_  = \new_[17699]_  & \new_[17694]_ ;
  assign \new_[17703]_  = ~A169 & ~A170;
  assign \new_[17707]_  = A200 & ~A199;
  assign \new_[17708]_  = ~A168 & \new_[17707]_ ;
  assign \new_[17709]_  = \new_[17708]_  & \new_[17703]_ ;
  assign \new_[17712]_  = A235 & A203;
  assign \new_[17716]_  = ~A302 & ~A301;
  assign \new_[17717]_  = ~A300 & \new_[17716]_ ;
  assign \new_[17718]_  = \new_[17717]_  & \new_[17712]_ ;
  assign \new_[17721]_  = ~A169 & ~A170;
  assign \new_[17725]_  = A200 & ~A199;
  assign \new_[17726]_  = ~A168 & \new_[17725]_ ;
  assign \new_[17727]_  = \new_[17726]_  & \new_[17721]_ ;
  assign \new_[17730]_  = A235 & A203;
  assign \new_[17734]_  = ~A301 & ~A299;
  assign \new_[17735]_  = ~A298 & \new_[17734]_ ;
  assign \new_[17736]_  = \new_[17735]_  & \new_[17730]_ ;
  assign \new_[17739]_  = ~A169 & ~A170;
  assign \new_[17743]_  = A200 & ~A199;
  assign \new_[17744]_  = ~A168 & \new_[17743]_ ;
  assign \new_[17745]_  = \new_[17744]_  & \new_[17739]_ ;
  assign \new_[17748]_  = A235 & A203;
  assign \new_[17752]_  = A269 & A266;
  assign \new_[17753]_  = ~A265 & \new_[17752]_ ;
  assign \new_[17754]_  = \new_[17753]_  & \new_[17748]_ ;
  assign \new_[17757]_  = ~A169 & ~A170;
  assign \new_[17761]_  = A200 & ~A199;
  assign \new_[17762]_  = ~A168 & \new_[17761]_ ;
  assign \new_[17763]_  = \new_[17762]_  & \new_[17757]_ ;
  assign \new_[17766]_  = A235 & A203;
  assign \new_[17770]_  = A269 & ~A266;
  assign \new_[17771]_  = A265 & \new_[17770]_ ;
  assign \new_[17772]_  = \new_[17771]_  & \new_[17766]_ ;
  assign \new_[17775]_  = ~A169 & ~A170;
  assign \new_[17779]_  = A200 & ~A199;
  assign \new_[17780]_  = ~A168 & \new_[17779]_ ;
  assign \new_[17781]_  = \new_[17780]_  & \new_[17775]_ ;
  assign \new_[17784]_  = A232 & A203;
  assign \new_[17788]_  = A267 & A265;
  assign \new_[17789]_  = A234 & \new_[17788]_ ;
  assign \new_[17790]_  = \new_[17789]_  & \new_[17784]_ ;
  assign \new_[17793]_  = ~A169 & ~A170;
  assign \new_[17797]_  = A200 & ~A199;
  assign \new_[17798]_  = ~A168 & \new_[17797]_ ;
  assign \new_[17799]_  = \new_[17798]_  & \new_[17793]_ ;
  assign \new_[17802]_  = A232 & A203;
  assign \new_[17806]_  = A267 & A266;
  assign \new_[17807]_  = A234 & \new_[17806]_ ;
  assign \new_[17808]_  = \new_[17807]_  & \new_[17802]_ ;
  assign \new_[17811]_  = ~A169 & ~A170;
  assign \new_[17815]_  = A200 & ~A199;
  assign \new_[17816]_  = ~A168 & \new_[17815]_ ;
  assign \new_[17817]_  = \new_[17816]_  & \new_[17811]_ ;
  assign \new_[17820]_  = A233 & A203;
  assign \new_[17824]_  = A267 & A265;
  assign \new_[17825]_  = A234 & \new_[17824]_ ;
  assign \new_[17826]_  = \new_[17825]_  & \new_[17820]_ ;
  assign \new_[17829]_  = ~A169 & ~A170;
  assign \new_[17833]_  = A200 & ~A199;
  assign \new_[17834]_  = ~A168 & \new_[17833]_ ;
  assign \new_[17835]_  = \new_[17834]_  & \new_[17829]_ ;
  assign \new_[17838]_  = A233 & A203;
  assign \new_[17842]_  = A267 & A266;
  assign \new_[17843]_  = A234 & \new_[17842]_ ;
  assign \new_[17844]_  = \new_[17843]_  & \new_[17838]_ ;
  assign \new_[17847]_  = ~A169 & ~A170;
  assign \new_[17851]_  = A200 & ~A199;
  assign \new_[17852]_  = ~A168 & \new_[17851]_ ;
  assign \new_[17853]_  = \new_[17852]_  & \new_[17847]_ ;
  assign \new_[17856]_  = ~A232 & A203;
  assign \new_[17860]_  = A268 & A236;
  assign \new_[17861]_  = A233 & \new_[17860]_ ;
  assign \new_[17862]_  = \new_[17861]_  & \new_[17856]_ ;
  assign \new_[17865]_  = ~A169 & ~A170;
  assign \new_[17869]_  = A200 & ~A199;
  assign \new_[17870]_  = ~A168 & \new_[17869]_ ;
  assign \new_[17871]_  = \new_[17870]_  & \new_[17865]_ ;
  assign \new_[17874]_  = A232 & A203;
  assign \new_[17878]_  = A268 & A236;
  assign \new_[17879]_  = ~A233 & \new_[17878]_ ;
  assign \new_[17880]_  = \new_[17879]_  & \new_[17874]_ ;
  assign \new_[17883]_  = ~A169 & ~A170;
  assign \new_[17887]_  = ~A200 & A199;
  assign \new_[17888]_  = ~A168 & \new_[17887]_ ;
  assign \new_[17889]_  = \new_[17888]_  & \new_[17883]_ ;
  assign \new_[17892]_  = A235 & A203;
  assign \new_[17896]_  = ~A302 & ~A301;
  assign \new_[17897]_  = ~A300 & \new_[17896]_ ;
  assign \new_[17898]_  = \new_[17897]_  & \new_[17892]_ ;
  assign \new_[17901]_  = ~A169 & ~A170;
  assign \new_[17905]_  = ~A200 & A199;
  assign \new_[17906]_  = ~A168 & \new_[17905]_ ;
  assign \new_[17907]_  = \new_[17906]_  & \new_[17901]_ ;
  assign \new_[17910]_  = A235 & A203;
  assign \new_[17914]_  = ~A301 & ~A299;
  assign \new_[17915]_  = ~A298 & \new_[17914]_ ;
  assign \new_[17916]_  = \new_[17915]_  & \new_[17910]_ ;
  assign \new_[17919]_  = ~A169 & ~A170;
  assign \new_[17923]_  = ~A200 & A199;
  assign \new_[17924]_  = ~A168 & \new_[17923]_ ;
  assign \new_[17925]_  = \new_[17924]_  & \new_[17919]_ ;
  assign \new_[17928]_  = A235 & A203;
  assign \new_[17932]_  = A269 & A266;
  assign \new_[17933]_  = ~A265 & \new_[17932]_ ;
  assign \new_[17934]_  = \new_[17933]_  & \new_[17928]_ ;
  assign \new_[17937]_  = ~A169 & ~A170;
  assign \new_[17941]_  = ~A200 & A199;
  assign \new_[17942]_  = ~A168 & \new_[17941]_ ;
  assign \new_[17943]_  = \new_[17942]_  & \new_[17937]_ ;
  assign \new_[17946]_  = A235 & A203;
  assign \new_[17950]_  = A269 & ~A266;
  assign \new_[17951]_  = A265 & \new_[17950]_ ;
  assign \new_[17952]_  = \new_[17951]_  & \new_[17946]_ ;
  assign \new_[17955]_  = ~A169 & ~A170;
  assign \new_[17959]_  = ~A200 & A199;
  assign \new_[17960]_  = ~A168 & \new_[17959]_ ;
  assign \new_[17961]_  = \new_[17960]_  & \new_[17955]_ ;
  assign \new_[17964]_  = A232 & A203;
  assign \new_[17968]_  = A267 & A265;
  assign \new_[17969]_  = A234 & \new_[17968]_ ;
  assign \new_[17970]_  = \new_[17969]_  & \new_[17964]_ ;
  assign \new_[17973]_  = ~A169 & ~A170;
  assign \new_[17977]_  = ~A200 & A199;
  assign \new_[17978]_  = ~A168 & \new_[17977]_ ;
  assign \new_[17979]_  = \new_[17978]_  & \new_[17973]_ ;
  assign \new_[17982]_  = A232 & A203;
  assign \new_[17986]_  = A267 & A266;
  assign \new_[17987]_  = A234 & \new_[17986]_ ;
  assign \new_[17988]_  = \new_[17987]_  & \new_[17982]_ ;
  assign \new_[17991]_  = ~A169 & ~A170;
  assign \new_[17995]_  = ~A200 & A199;
  assign \new_[17996]_  = ~A168 & \new_[17995]_ ;
  assign \new_[17997]_  = \new_[17996]_  & \new_[17991]_ ;
  assign \new_[18000]_  = A233 & A203;
  assign \new_[18004]_  = A267 & A265;
  assign \new_[18005]_  = A234 & \new_[18004]_ ;
  assign \new_[18006]_  = \new_[18005]_  & \new_[18000]_ ;
  assign \new_[18009]_  = ~A169 & ~A170;
  assign \new_[18013]_  = ~A200 & A199;
  assign \new_[18014]_  = ~A168 & \new_[18013]_ ;
  assign \new_[18015]_  = \new_[18014]_  & \new_[18009]_ ;
  assign \new_[18018]_  = A233 & A203;
  assign \new_[18022]_  = A267 & A266;
  assign \new_[18023]_  = A234 & \new_[18022]_ ;
  assign \new_[18024]_  = \new_[18023]_  & \new_[18018]_ ;
  assign \new_[18027]_  = ~A169 & ~A170;
  assign \new_[18031]_  = ~A200 & A199;
  assign \new_[18032]_  = ~A168 & \new_[18031]_ ;
  assign \new_[18033]_  = \new_[18032]_  & \new_[18027]_ ;
  assign \new_[18036]_  = ~A232 & A203;
  assign \new_[18040]_  = A268 & A236;
  assign \new_[18041]_  = A233 & \new_[18040]_ ;
  assign \new_[18042]_  = \new_[18041]_  & \new_[18036]_ ;
  assign \new_[18045]_  = ~A169 & ~A170;
  assign \new_[18049]_  = ~A200 & A199;
  assign \new_[18050]_  = ~A168 & \new_[18049]_ ;
  assign \new_[18051]_  = \new_[18050]_  & \new_[18045]_ ;
  assign \new_[18054]_  = A232 & A203;
  assign \new_[18058]_  = A268 & A236;
  assign \new_[18059]_  = ~A233 & \new_[18058]_ ;
  assign \new_[18060]_  = \new_[18059]_  & \new_[18054]_ ;
  assign \new_[18063]_  = A166 & A168;
  assign \new_[18067]_  = ~A203 & ~A202;
  assign \new_[18068]_  = ~A201 & \new_[18067]_ ;
  assign \new_[18069]_  = \new_[18068]_  & \new_[18063]_ ;
  assign \new_[18073]_  = A298 & A234;
  assign \new_[18074]_  = A232 & \new_[18073]_ ;
  assign \new_[18078]_  = ~A301 & ~A300;
  assign \new_[18079]_  = A299 & \new_[18078]_ ;
  assign \new_[18080]_  = \new_[18079]_  & \new_[18074]_ ;
  assign \new_[18083]_  = A166 & A168;
  assign \new_[18087]_  = ~A203 & ~A202;
  assign \new_[18088]_  = ~A201 & \new_[18087]_ ;
  assign \new_[18089]_  = \new_[18088]_  & \new_[18083]_ ;
  assign \new_[18093]_  = A298 & A234;
  assign \new_[18094]_  = A233 & \new_[18093]_ ;
  assign \new_[18098]_  = ~A301 & ~A300;
  assign \new_[18099]_  = A299 & \new_[18098]_ ;
  assign \new_[18100]_  = \new_[18099]_  & \new_[18094]_ ;
  assign \new_[18103]_  = A166 & A168;
  assign \new_[18107]_  = ~A203 & ~A202;
  assign \new_[18108]_  = ~A201 & \new_[18107]_ ;
  assign \new_[18109]_  = \new_[18108]_  & \new_[18103]_ ;
  assign \new_[18113]_  = A236 & A233;
  assign \new_[18114]_  = ~A232 & \new_[18113]_ ;
  assign \new_[18118]_  = ~A302 & ~A301;
  assign \new_[18119]_  = ~A300 & \new_[18118]_ ;
  assign \new_[18120]_  = \new_[18119]_  & \new_[18114]_ ;
  assign \new_[18123]_  = A166 & A168;
  assign \new_[18127]_  = ~A203 & ~A202;
  assign \new_[18128]_  = ~A201 & \new_[18127]_ ;
  assign \new_[18129]_  = \new_[18128]_  & \new_[18123]_ ;
  assign \new_[18133]_  = A236 & A233;
  assign \new_[18134]_  = ~A232 & \new_[18133]_ ;
  assign \new_[18138]_  = ~A301 & ~A299;
  assign \new_[18139]_  = ~A298 & \new_[18138]_ ;
  assign \new_[18140]_  = \new_[18139]_  & \new_[18134]_ ;
  assign \new_[18143]_  = A166 & A168;
  assign \new_[18147]_  = ~A203 & ~A202;
  assign \new_[18148]_  = ~A201 & \new_[18147]_ ;
  assign \new_[18149]_  = \new_[18148]_  & \new_[18143]_ ;
  assign \new_[18153]_  = A236 & A233;
  assign \new_[18154]_  = ~A232 & \new_[18153]_ ;
  assign \new_[18158]_  = A269 & A266;
  assign \new_[18159]_  = ~A265 & \new_[18158]_ ;
  assign \new_[18160]_  = \new_[18159]_  & \new_[18154]_ ;
  assign \new_[18163]_  = A166 & A168;
  assign \new_[18167]_  = ~A203 & ~A202;
  assign \new_[18168]_  = ~A201 & \new_[18167]_ ;
  assign \new_[18169]_  = \new_[18168]_  & \new_[18163]_ ;
  assign \new_[18173]_  = A236 & A233;
  assign \new_[18174]_  = ~A232 & \new_[18173]_ ;
  assign \new_[18178]_  = A269 & ~A266;
  assign \new_[18179]_  = A265 & \new_[18178]_ ;
  assign \new_[18180]_  = \new_[18179]_  & \new_[18174]_ ;
  assign \new_[18183]_  = A166 & A168;
  assign \new_[18187]_  = ~A203 & ~A202;
  assign \new_[18188]_  = ~A201 & \new_[18187]_ ;
  assign \new_[18189]_  = \new_[18188]_  & \new_[18183]_ ;
  assign \new_[18193]_  = A236 & ~A233;
  assign \new_[18194]_  = A232 & \new_[18193]_ ;
  assign \new_[18198]_  = ~A302 & ~A301;
  assign \new_[18199]_  = ~A300 & \new_[18198]_ ;
  assign \new_[18200]_  = \new_[18199]_  & \new_[18194]_ ;
  assign \new_[18203]_  = A166 & A168;
  assign \new_[18207]_  = ~A203 & ~A202;
  assign \new_[18208]_  = ~A201 & \new_[18207]_ ;
  assign \new_[18209]_  = \new_[18208]_  & \new_[18203]_ ;
  assign \new_[18213]_  = A236 & ~A233;
  assign \new_[18214]_  = A232 & \new_[18213]_ ;
  assign \new_[18218]_  = ~A301 & ~A299;
  assign \new_[18219]_  = ~A298 & \new_[18218]_ ;
  assign \new_[18220]_  = \new_[18219]_  & \new_[18214]_ ;
  assign \new_[18223]_  = A166 & A168;
  assign \new_[18227]_  = ~A203 & ~A202;
  assign \new_[18228]_  = ~A201 & \new_[18227]_ ;
  assign \new_[18229]_  = \new_[18228]_  & \new_[18223]_ ;
  assign \new_[18233]_  = A236 & ~A233;
  assign \new_[18234]_  = A232 & \new_[18233]_ ;
  assign \new_[18238]_  = A269 & A266;
  assign \new_[18239]_  = ~A265 & \new_[18238]_ ;
  assign \new_[18240]_  = \new_[18239]_  & \new_[18234]_ ;
  assign \new_[18243]_  = A166 & A168;
  assign \new_[18247]_  = ~A203 & ~A202;
  assign \new_[18248]_  = ~A201 & \new_[18247]_ ;
  assign \new_[18249]_  = \new_[18248]_  & \new_[18243]_ ;
  assign \new_[18253]_  = A236 & ~A233;
  assign \new_[18254]_  = A232 & \new_[18253]_ ;
  assign \new_[18258]_  = A269 & ~A266;
  assign \new_[18259]_  = A265 & \new_[18258]_ ;
  assign \new_[18260]_  = \new_[18259]_  & \new_[18254]_ ;
  assign \new_[18263]_  = A166 & A168;
  assign \new_[18267]_  = ~A201 & A200;
  assign \new_[18268]_  = A199 & \new_[18267]_ ;
  assign \new_[18269]_  = \new_[18268]_  & \new_[18263]_ ;
  assign \new_[18273]_  = A298 & A235;
  assign \new_[18274]_  = ~A202 & \new_[18273]_ ;
  assign \new_[18278]_  = ~A301 & ~A300;
  assign \new_[18279]_  = A299 & \new_[18278]_ ;
  assign \new_[18280]_  = \new_[18279]_  & \new_[18274]_ ;
  assign \new_[18283]_  = A166 & A168;
  assign \new_[18287]_  = ~A201 & A200;
  assign \new_[18288]_  = A199 & \new_[18287]_ ;
  assign \new_[18289]_  = \new_[18288]_  & \new_[18283]_ ;
  assign \new_[18293]_  = A234 & A232;
  assign \new_[18294]_  = ~A202 & \new_[18293]_ ;
  assign \new_[18298]_  = ~A302 & ~A301;
  assign \new_[18299]_  = ~A300 & \new_[18298]_ ;
  assign \new_[18300]_  = \new_[18299]_  & \new_[18294]_ ;
  assign \new_[18303]_  = A166 & A168;
  assign \new_[18307]_  = ~A201 & A200;
  assign \new_[18308]_  = A199 & \new_[18307]_ ;
  assign \new_[18309]_  = \new_[18308]_  & \new_[18303]_ ;
  assign \new_[18313]_  = A234 & A232;
  assign \new_[18314]_  = ~A202 & \new_[18313]_ ;
  assign \new_[18318]_  = ~A301 & ~A299;
  assign \new_[18319]_  = ~A298 & \new_[18318]_ ;
  assign \new_[18320]_  = \new_[18319]_  & \new_[18314]_ ;
  assign \new_[18323]_  = A166 & A168;
  assign \new_[18327]_  = ~A201 & A200;
  assign \new_[18328]_  = A199 & \new_[18327]_ ;
  assign \new_[18329]_  = \new_[18328]_  & \new_[18323]_ ;
  assign \new_[18333]_  = A234 & A232;
  assign \new_[18334]_  = ~A202 & \new_[18333]_ ;
  assign \new_[18338]_  = A269 & A266;
  assign \new_[18339]_  = ~A265 & \new_[18338]_ ;
  assign \new_[18340]_  = \new_[18339]_  & \new_[18334]_ ;
  assign \new_[18343]_  = A166 & A168;
  assign \new_[18347]_  = ~A201 & A200;
  assign \new_[18348]_  = A199 & \new_[18347]_ ;
  assign \new_[18349]_  = \new_[18348]_  & \new_[18343]_ ;
  assign \new_[18353]_  = A234 & A232;
  assign \new_[18354]_  = ~A202 & \new_[18353]_ ;
  assign \new_[18358]_  = A269 & ~A266;
  assign \new_[18359]_  = A265 & \new_[18358]_ ;
  assign \new_[18360]_  = \new_[18359]_  & \new_[18354]_ ;
  assign \new_[18363]_  = A166 & A168;
  assign \new_[18367]_  = ~A201 & A200;
  assign \new_[18368]_  = A199 & \new_[18367]_ ;
  assign \new_[18369]_  = \new_[18368]_  & \new_[18363]_ ;
  assign \new_[18373]_  = A234 & A233;
  assign \new_[18374]_  = ~A202 & \new_[18373]_ ;
  assign \new_[18378]_  = ~A302 & ~A301;
  assign \new_[18379]_  = ~A300 & \new_[18378]_ ;
  assign \new_[18380]_  = \new_[18379]_  & \new_[18374]_ ;
  assign \new_[18383]_  = A166 & A168;
  assign \new_[18387]_  = ~A201 & A200;
  assign \new_[18388]_  = A199 & \new_[18387]_ ;
  assign \new_[18389]_  = \new_[18388]_  & \new_[18383]_ ;
  assign \new_[18393]_  = A234 & A233;
  assign \new_[18394]_  = ~A202 & \new_[18393]_ ;
  assign \new_[18398]_  = ~A301 & ~A299;
  assign \new_[18399]_  = ~A298 & \new_[18398]_ ;
  assign \new_[18400]_  = \new_[18399]_  & \new_[18394]_ ;
  assign \new_[18403]_  = A166 & A168;
  assign \new_[18407]_  = ~A201 & A200;
  assign \new_[18408]_  = A199 & \new_[18407]_ ;
  assign \new_[18409]_  = \new_[18408]_  & \new_[18403]_ ;
  assign \new_[18413]_  = A234 & A233;
  assign \new_[18414]_  = ~A202 & \new_[18413]_ ;
  assign \new_[18418]_  = A269 & A266;
  assign \new_[18419]_  = ~A265 & \new_[18418]_ ;
  assign \new_[18420]_  = \new_[18419]_  & \new_[18414]_ ;
  assign \new_[18423]_  = A166 & A168;
  assign \new_[18427]_  = ~A201 & A200;
  assign \new_[18428]_  = A199 & \new_[18427]_ ;
  assign \new_[18429]_  = \new_[18428]_  & \new_[18423]_ ;
  assign \new_[18433]_  = A234 & A233;
  assign \new_[18434]_  = ~A202 & \new_[18433]_ ;
  assign \new_[18438]_  = A269 & ~A266;
  assign \new_[18439]_  = A265 & \new_[18438]_ ;
  assign \new_[18440]_  = \new_[18439]_  & \new_[18434]_ ;
  assign \new_[18443]_  = A166 & A168;
  assign \new_[18447]_  = ~A201 & A200;
  assign \new_[18448]_  = A199 & \new_[18447]_ ;
  assign \new_[18449]_  = \new_[18448]_  & \new_[18443]_ ;
  assign \new_[18453]_  = A233 & ~A232;
  assign \new_[18454]_  = ~A202 & \new_[18453]_ ;
  assign \new_[18458]_  = A267 & A265;
  assign \new_[18459]_  = A236 & \new_[18458]_ ;
  assign \new_[18460]_  = \new_[18459]_  & \new_[18454]_ ;
  assign \new_[18463]_  = A166 & A168;
  assign \new_[18467]_  = ~A201 & A200;
  assign \new_[18468]_  = A199 & \new_[18467]_ ;
  assign \new_[18469]_  = \new_[18468]_  & \new_[18463]_ ;
  assign \new_[18473]_  = A233 & ~A232;
  assign \new_[18474]_  = ~A202 & \new_[18473]_ ;
  assign \new_[18478]_  = A267 & A266;
  assign \new_[18479]_  = A236 & \new_[18478]_ ;
  assign \new_[18480]_  = \new_[18479]_  & \new_[18474]_ ;
  assign \new_[18483]_  = A166 & A168;
  assign \new_[18487]_  = ~A201 & A200;
  assign \new_[18488]_  = A199 & \new_[18487]_ ;
  assign \new_[18489]_  = \new_[18488]_  & \new_[18483]_ ;
  assign \new_[18493]_  = ~A233 & A232;
  assign \new_[18494]_  = ~A202 & \new_[18493]_ ;
  assign \new_[18498]_  = A267 & A265;
  assign \new_[18499]_  = A236 & \new_[18498]_ ;
  assign \new_[18500]_  = \new_[18499]_  & \new_[18494]_ ;
  assign \new_[18503]_  = A166 & A168;
  assign \new_[18507]_  = ~A201 & A200;
  assign \new_[18508]_  = A199 & \new_[18507]_ ;
  assign \new_[18509]_  = \new_[18508]_  & \new_[18503]_ ;
  assign \new_[18513]_  = ~A233 & A232;
  assign \new_[18514]_  = ~A202 & \new_[18513]_ ;
  assign \new_[18518]_  = A267 & A266;
  assign \new_[18519]_  = A236 & \new_[18518]_ ;
  assign \new_[18520]_  = \new_[18519]_  & \new_[18514]_ ;
  assign \new_[18523]_  = A166 & A168;
  assign \new_[18527]_  = ~A202 & ~A200;
  assign \new_[18528]_  = ~A199 & \new_[18527]_ ;
  assign \new_[18529]_  = \new_[18528]_  & \new_[18523]_ ;
  assign \new_[18533]_  = A298 & A234;
  assign \new_[18534]_  = A232 & \new_[18533]_ ;
  assign \new_[18538]_  = ~A301 & ~A300;
  assign \new_[18539]_  = A299 & \new_[18538]_ ;
  assign \new_[18540]_  = \new_[18539]_  & \new_[18534]_ ;
  assign \new_[18543]_  = A166 & A168;
  assign \new_[18547]_  = ~A202 & ~A200;
  assign \new_[18548]_  = ~A199 & \new_[18547]_ ;
  assign \new_[18549]_  = \new_[18548]_  & \new_[18543]_ ;
  assign \new_[18553]_  = A298 & A234;
  assign \new_[18554]_  = A233 & \new_[18553]_ ;
  assign \new_[18558]_  = ~A301 & ~A300;
  assign \new_[18559]_  = A299 & \new_[18558]_ ;
  assign \new_[18560]_  = \new_[18559]_  & \new_[18554]_ ;
  assign \new_[18563]_  = A166 & A168;
  assign \new_[18567]_  = ~A202 & ~A200;
  assign \new_[18568]_  = ~A199 & \new_[18567]_ ;
  assign \new_[18569]_  = \new_[18568]_  & \new_[18563]_ ;
  assign \new_[18573]_  = A236 & A233;
  assign \new_[18574]_  = ~A232 & \new_[18573]_ ;
  assign \new_[18578]_  = ~A302 & ~A301;
  assign \new_[18579]_  = ~A300 & \new_[18578]_ ;
  assign \new_[18580]_  = \new_[18579]_  & \new_[18574]_ ;
  assign \new_[18583]_  = A166 & A168;
  assign \new_[18587]_  = ~A202 & ~A200;
  assign \new_[18588]_  = ~A199 & \new_[18587]_ ;
  assign \new_[18589]_  = \new_[18588]_  & \new_[18583]_ ;
  assign \new_[18593]_  = A236 & A233;
  assign \new_[18594]_  = ~A232 & \new_[18593]_ ;
  assign \new_[18598]_  = ~A301 & ~A299;
  assign \new_[18599]_  = ~A298 & \new_[18598]_ ;
  assign \new_[18600]_  = \new_[18599]_  & \new_[18594]_ ;
  assign \new_[18603]_  = A166 & A168;
  assign \new_[18607]_  = ~A202 & ~A200;
  assign \new_[18608]_  = ~A199 & \new_[18607]_ ;
  assign \new_[18609]_  = \new_[18608]_  & \new_[18603]_ ;
  assign \new_[18613]_  = A236 & A233;
  assign \new_[18614]_  = ~A232 & \new_[18613]_ ;
  assign \new_[18618]_  = A269 & A266;
  assign \new_[18619]_  = ~A265 & \new_[18618]_ ;
  assign \new_[18620]_  = \new_[18619]_  & \new_[18614]_ ;
  assign \new_[18623]_  = A166 & A168;
  assign \new_[18627]_  = ~A202 & ~A200;
  assign \new_[18628]_  = ~A199 & \new_[18627]_ ;
  assign \new_[18629]_  = \new_[18628]_  & \new_[18623]_ ;
  assign \new_[18633]_  = A236 & A233;
  assign \new_[18634]_  = ~A232 & \new_[18633]_ ;
  assign \new_[18638]_  = A269 & ~A266;
  assign \new_[18639]_  = A265 & \new_[18638]_ ;
  assign \new_[18640]_  = \new_[18639]_  & \new_[18634]_ ;
  assign \new_[18643]_  = A166 & A168;
  assign \new_[18647]_  = ~A202 & ~A200;
  assign \new_[18648]_  = ~A199 & \new_[18647]_ ;
  assign \new_[18649]_  = \new_[18648]_  & \new_[18643]_ ;
  assign \new_[18653]_  = A236 & ~A233;
  assign \new_[18654]_  = A232 & \new_[18653]_ ;
  assign \new_[18658]_  = ~A302 & ~A301;
  assign \new_[18659]_  = ~A300 & \new_[18658]_ ;
  assign \new_[18660]_  = \new_[18659]_  & \new_[18654]_ ;
  assign \new_[18663]_  = A166 & A168;
  assign \new_[18667]_  = ~A202 & ~A200;
  assign \new_[18668]_  = ~A199 & \new_[18667]_ ;
  assign \new_[18669]_  = \new_[18668]_  & \new_[18663]_ ;
  assign \new_[18673]_  = A236 & ~A233;
  assign \new_[18674]_  = A232 & \new_[18673]_ ;
  assign \new_[18678]_  = ~A301 & ~A299;
  assign \new_[18679]_  = ~A298 & \new_[18678]_ ;
  assign \new_[18680]_  = \new_[18679]_  & \new_[18674]_ ;
  assign \new_[18683]_  = A166 & A168;
  assign \new_[18687]_  = ~A202 & ~A200;
  assign \new_[18688]_  = ~A199 & \new_[18687]_ ;
  assign \new_[18689]_  = \new_[18688]_  & \new_[18683]_ ;
  assign \new_[18693]_  = A236 & ~A233;
  assign \new_[18694]_  = A232 & \new_[18693]_ ;
  assign \new_[18698]_  = A269 & A266;
  assign \new_[18699]_  = ~A265 & \new_[18698]_ ;
  assign \new_[18700]_  = \new_[18699]_  & \new_[18694]_ ;
  assign \new_[18703]_  = A166 & A168;
  assign \new_[18707]_  = ~A202 & ~A200;
  assign \new_[18708]_  = ~A199 & \new_[18707]_ ;
  assign \new_[18709]_  = \new_[18708]_  & \new_[18703]_ ;
  assign \new_[18713]_  = A236 & ~A233;
  assign \new_[18714]_  = A232 & \new_[18713]_ ;
  assign \new_[18718]_  = A269 & ~A266;
  assign \new_[18719]_  = A265 & \new_[18718]_ ;
  assign \new_[18720]_  = \new_[18719]_  & \new_[18714]_ ;
  assign \new_[18723]_  = A167 & A168;
  assign \new_[18727]_  = ~A203 & ~A202;
  assign \new_[18728]_  = ~A201 & \new_[18727]_ ;
  assign \new_[18729]_  = \new_[18728]_  & \new_[18723]_ ;
  assign \new_[18733]_  = A298 & A234;
  assign \new_[18734]_  = A232 & \new_[18733]_ ;
  assign \new_[18738]_  = ~A301 & ~A300;
  assign \new_[18739]_  = A299 & \new_[18738]_ ;
  assign \new_[18740]_  = \new_[18739]_  & \new_[18734]_ ;
  assign \new_[18743]_  = A167 & A168;
  assign \new_[18747]_  = ~A203 & ~A202;
  assign \new_[18748]_  = ~A201 & \new_[18747]_ ;
  assign \new_[18749]_  = \new_[18748]_  & \new_[18743]_ ;
  assign \new_[18753]_  = A298 & A234;
  assign \new_[18754]_  = A233 & \new_[18753]_ ;
  assign \new_[18758]_  = ~A301 & ~A300;
  assign \new_[18759]_  = A299 & \new_[18758]_ ;
  assign \new_[18760]_  = \new_[18759]_  & \new_[18754]_ ;
  assign \new_[18763]_  = A167 & A168;
  assign \new_[18767]_  = ~A203 & ~A202;
  assign \new_[18768]_  = ~A201 & \new_[18767]_ ;
  assign \new_[18769]_  = \new_[18768]_  & \new_[18763]_ ;
  assign \new_[18773]_  = A236 & A233;
  assign \new_[18774]_  = ~A232 & \new_[18773]_ ;
  assign \new_[18778]_  = ~A302 & ~A301;
  assign \new_[18779]_  = ~A300 & \new_[18778]_ ;
  assign \new_[18780]_  = \new_[18779]_  & \new_[18774]_ ;
  assign \new_[18783]_  = A167 & A168;
  assign \new_[18787]_  = ~A203 & ~A202;
  assign \new_[18788]_  = ~A201 & \new_[18787]_ ;
  assign \new_[18789]_  = \new_[18788]_  & \new_[18783]_ ;
  assign \new_[18793]_  = A236 & A233;
  assign \new_[18794]_  = ~A232 & \new_[18793]_ ;
  assign \new_[18798]_  = ~A301 & ~A299;
  assign \new_[18799]_  = ~A298 & \new_[18798]_ ;
  assign \new_[18800]_  = \new_[18799]_  & \new_[18794]_ ;
  assign \new_[18803]_  = A167 & A168;
  assign \new_[18807]_  = ~A203 & ~A202;
  assign \new_[18808]_  = ~A201 & \new_[18807]_ ;
  assign \new_[18809]_  = \new_[18808]_  & \new_[18803]_ ;
  assign \new_[18813]_  = A236 & A233;
  assign \new_[18814]_  = ~A232 & \new_[18813]_ ;
  assign \new_[18818]_  = A269 & A266;
  assign \new_[18819]_  = ~A265 & \new_[18818]_ ;
  assign \new_[18820]_  = \new_[18819]_  & \new_[18814]_ ;
  assign \new_[18823]_  = A167 & A168;
  assign \new_[18827]_  = ~A203 & ~A202;
  assign \new_[18828]_  = ~A201 & \new_[18827]_ ;
  assign \new_[18829]_  = \new_[18828]_  & \new_[18823]_ ;
  assign \new_[18833]_  = A236 & A233;
  assign \new_[18834]_  = ~A232 & \new_[18833]_ ;
  assign \new_[18838]_  = A269 & ~A266;
  assign \new_[18839]_  = A265 & \new_[18838]_ ;
  assign \new_[18840]_  = \new_[18839]_  & \new_[18834]_ ;
  assign \new_[18843]_  = A167 & A168;
  assign \new_[18847]_  = ~A203 & ~A202;
  assign \new_[18848]_  = ~A201 & \new_[18847]_ ;
  assign \new_[18849]_  = \new_[18848]_  & \new_[18843]_ ;
  assign \new_[18853]_  = A236 & ~A233;
  assign \new_[18854]_  = A232 & \new_[18853]_ ;
  assign \new_[18858]_  = ~A302 & ~A301;
  assign \new_[18859]_  = ~A300 & \new_[18858]_ ;
  assign \new_[18860]_  = \new_[18859]_  & \new_[18854]_ ;
  assign \new_[18863]_  = A167 & A168;
  assign \new_[18867]_  = ~A203 & ~A202;
  assign \new_[18868]_  = ~A201 & \new_[18867]_ ;
  assign \new_[18869]_  = \new_[18868]_  & \new_[18863]_ ;
  assign \new_[18873]_  = A236 & ~A233;
  assign \new_[18874]_  = A232 & \new_[18873]_ ;
  assign \new_[18878]_  = ~A301 & ~A299;
  assign \new_[18879]_  = ~A298 & \new_[18878]_ ;
  assign \new_[18880]_  = \new_[18879]_  & \new_[18874]_ ;
  assign \new_[18883]_  = A167 & A168;
  assign \new_[18887]_  = ~A203 & ~A202;
  assign \new_[18888]_  = ~A201 & \new_[18887]_ ;
  assign \new_[18889]_  = \new_[18888]_  & \new_[18883]_ ;
  assign \new_[18893]_  = A236 & ~A233;
  assign \new_[18894]_  = A232 & \new_[18893]_ ;
  assign \new_[18898]_  = A269 & A266;
  assign \new_[18899]_  = ~A265 & \new_[18898]_ ;
  assign \new_[18900]_  = \new_[18899]_  & \new_[18894]_ ;
  assign \new_[18903]_  = A167 & A168;
  assign \new_[18907]_  = ~A203 & ~A202;
  assign \new_[18908]_  = ~A201 & \new_[18907]_ ;
  assign \new_[18909]_  = \new_[18908]_  & \new_[18903]_ ;
  assign \new_[18913]_  = A236 & ~A233;
  assign \new_[18914]_  = A232 & \new_[18913]_ ;
  assign \new_[18918]_  = A269 & ~A266;
  assign \new_[18919]_  = A265 & \new_[18918]_ ;
  assign \new_[18920]_  = \new_[18919]_  & \new_[18914]_ ;
  assign \new_[18923]_  = A167 & A168;
  assign \new_[18927]_  = ~A201 & A200;
  assign \new_[18928]_  = A199 & \new_[18927]_ ;
  assign \new_[18929]_  = \new_[18928]_  & \new_[18923]_ ;
  assign \new_[18933]_  = A298 & A235;
  assign \new_[18934]_  = ~A202 & \new_[18933]_ ;
  assign \new_[18938]_  = ~A301 & ~A300;
  assign \new_[18939]_  = A299 & \new_[18938]_ ;
  assign \new_[18940]_  = \new_[18939]_  & \new_[18934]_ ;
  assign \new_[18943]_  = A167 & A168;
  assign \new_[18947]_  = ~A201 & A200;
  assign \new_[18948]_  = A199 & \new_[18947]_ ;
  assign \new_[18949]_  = \new_[18948]_  & \new_[18943]_ ;
  assign \new_[18953]_  = A234 & A232;
  assign \new_[18954]_  = ~A202 & \new_[18953]_ ;
  assign \new_[18958]_  = ~A302 & ~A301;
  assign \new_[18959]_  = ~A300 & \new_[18958]_ ;
  assign \new_[18960]_  = \new_[18959]_  & \new_[18954]_ ;
  assign \new_[18963]_  = A167 & A168;
  assign \new_[18967]_  = ~A201 & A200;
  assign \new_[18968]_  = A199 & \new_[18967]_ ;
  assign \new_[18969]_  = \new_[18968]_  & \new_[18963]_ ;
  assign \new_[18973]_  = A234 & A232;
  assign \new_[18974]_  = ~A202 & \new_[18973]_ ;
  assign \new_[18978]_  = ~A301 & ~A299;
  assign \new_[18979]_  = ~A298 & \new_[18978]_ ;
  assign \new_[18980]_  = \new_[18979]_  & \new_[18974]_ ;
  assign \new_[18983]_  = A167 & A168;
  assign \new_[18987]_  = ~A201 & A200;
  assign \new_[18988]_  = A199 & \new_[18987]_ ;
  assign \new_[18989]_  = \new_[18988]_  & \new_[18983]_ ;
  assign \new_[18993]_  = A234 & A232;
  assign \new_[18994]_  = ~A202 & \new_[18993]_ ;
  assign \new_[18998]_  = A269 & A266;
  assign \new_[18999]_  = ~A265 & \new_[18998]_ ;
  assign \new_[19000]_  = \new_[18999]_  & \new_[18994]_ ;
  assign \new_[19003]_  = A167 & A168;
  assign \new_[19007]_  = ~A201 & A200;
  assign \new_[19008]_  = A199 & \new_[19007]_ ;
  assign \new_[19009]_  = \new_[19008]_  & \new_[19003]_ ;
  assign \new_[19013]_  = A234 & A232;
  assign \new_[19014]_  = ~A202 & \new_[19013]_ ;
  assign \new_[19018]_  = A269 & ~A266;
  assign \new_[19019]_  = A265 & \new_[19018]_ ;
  assign \new_[19020]_  = \new_[19019]_  & \new_[19014]_ ;
  assign \new_[19023]_  = A167 & A168;
  assign \new_[19027]_  = ~A201 & A200;
  assign \new_[19028]_  = A199 & \new_[19027]_ ;
  assign \new_[19029]_  = \new_[19028]_  & \new_[19023]_ ;
  assign \new_[19033]_  = A234 & A233;
  assign \new_[19034]_  = ~A202 & \new_[19033]_ ;
  assign \new_[19038]_  = ~A302 & ~A301;
  assign \new_[19039]_  = ~A300 & \new_[19038]_ ;
  assign \new_[19040]_  = \new_[19039]_  & \new_[19034]_ ;
  assign \new_[19043]_  = A167 & A168;
  assign \new_[19047]_  = ~A201 & A200;
  assign \new_[19048]_  = A199 & \new_[19047]_ ;
  assign \new_[19049]_  = \new_[19048]_  & \new_[19043]_ ;
  assign \new_[19053]_  = A234 & A233;
  assign \new_[19054]_  = ~A202 & \new_[19053]_ ;
  assign \new_[19058]_  = ~A301 & ~A299;
  assign \new_[19059]_  = ~A298 & \new_[19058]_ ;
  assign \new_[19060]_  = \new_[19059]_  & \new_[19054]_ ;
  assign \new_[19063]_  = A167 & A168;
  assign \new_[19067]_  = ~A201 & A200;
  assign \new_[19068]_  = A199 & \new_[19067]_ ;
  assign \new_[19069]_  = \new_[19068]_  & \new_[19063]_ ;
  assign \new_[19073]_  = A234 & A233;
  assign \new_[19074]_  = ~A202 & \new_[19073]_ ;
  assign \new_[19078]_  = A269 & A266;
  assign \new_[19079]_  = ~A265 & \new_[19078]_ ;
  assign \new_[19080]_  = \new_[19079]_  & \new_[19074]_ ;
  assign \new_[19083]_  = A167 & A168;
  assign \new_[19087]_  = ~A201 & A200;
  assign \new_[19088]_  = A199 & \new_[19087]_ ;
  assign \new_[19089]_  = \new_[19088]_  & \new_[19083]_ ;
  assign \new_[19093]_  = A234 & A233;
  assign \new_[19094]_  = ~A202 & \new_[19093]_ ;
  assign \new_[19098]_  = A269 & ~A266;
  assign \new_[19099]_  = A265 & \new_[19098]_ ;
  assign \new_[19100]_  = \new_[19099]_  & \new_[19094]_ ;
  assign \new_[19103]_  = A167 & A168;
  assign \new_[19107]_  = ~A201 & A200;
  assign \new_[19108]_  = A199 & \new_[19107]_ ;
  assign \new_[19109]_  = \new_[19108]_  & \new_[19103]_ ;
  assign \new_[19113]_  = A233 & ~A232;
  assign \new_[19114]_  = ~A202 & \new_[19113]_ ;
  assign \new_[19118]_  = A267 & A265;
  assign \new_[19119]_  = A236 & \new_[19118]_ ;
  assign \new_[19120]_  = \new_[19119]_  & \new_[19114]_ ;
  assign \new_[19123]_  = A167 & A168;
  assign \new_[19127]_  = ~A201 & A200;
  assign \new_[19128]_  = A199 & \new_[19127]_ ;
  assign \new_[19129]_  = \new_[19128]_  & \new_[19123]_ ;
  assign \new_[19133]_  = A233 & ~A232;
  assign \new_[19134]_  = ~A202 & \new_[19133]_ ;
  assign \new_[19138]_  = A267 & A266;
  assign \new_[19139]_  = A236 & \new_[19138]_ ;
  assign \new_[19140]_  = \new_[19139]_  & \new_[19134]_ ;
  assign \new_[19143]_  = A167 & A168;
  assign \new_[19147]_  = ~A201 & A200;
  assign \new_[19148]_  = A199 & \new_[19147]_ ;
  assign \new_[19149]_  = \new_[19148]_  & \new_[19143]_ ;
  assign \new_[19153]_  = ~A233 & A232;
  assign \new_[19154]_  = ~A202 & \new_[19153]_ ;
  assign \new_[19158]_  = A267 & A265;
  assign \new_[19159]_  = A236 & \new_[19158]_ ;
  assign \new_[19160]_  = \new_[19159]_  & \new_[19154]_ ;
  assign \new_[19163]_  = A167 & A168;
  assign \new_[19167]_  = ~A201 & A200;
  assign \new_[19168]_  = A199 & \new_[19167]_ ;
  assign \new_[19169]_  = \new_[19168]_  & \new_[19163]_ ;
  assign \new_[19173]_  = ~A233 & A232;
  assign \new_[19174]_  = ~A202 & \new_[19173]_ ;
  assign \new_[19178]_  = A267 & A266;
  assign \new_[19179]_  = A236 & \new_[19178]_ ;
  assign \new_[19180]_  = \new_[19179]_  & \new_[19174]_ ;
  assign \new_[19183]_  = A167 & A168;
  assign \new_[19187]_  = ~A202 & ~A200;
  assign \new_[19188]_  = ~A199 & \new_[19187]_ ;
  assign \new_[19189]_  = \new_[19188]_  & \new_[19183]_ ;
  assign \new_[19193]_  = A298 & A234;
  assign \new_[19194]_  = A232 & \new_[19193]_ ;
  assign \new_[19198]_  = ~A301 & ~A300;
  assign \new_[19199]_  = A299 & \new_[19198]_ ;
  assign \new_[19200]_  = \new_[19199]_  & \new_[19194]_ ;
  assign \new_[19203]_  = A167 & A168;
  assign \new_[19207]_  = ~A202 & ~A200;
  assign \new_[19208]_  = ~A199 & \new_[19207]_ ;
  assign \new_[19209]_  = \new_[19208]_  & \new_[19203]_ ;
  assign \new_[19213]_  = A298 & A234;
  assign \new_[19214]_  = A233 & \new_[19213]_ ;
  assign \new_[19218]_  = ~A301 & ~A300;
  assign \new_[19219]_  = A299 & \new_[19218]_ ;
  assign \new_[19220]_  = \new_[19219]_  & \new_[19214]_ ;
  assign \new_[19223]_  = A167 & A168;
  assign \new_[19227]_  = ~A202 & ~A200;
  assign \new_[19228]_  = ~A199 & \new_[19227]_ ;
  assign \new_[19229]_  = \new_[19228]_  & \new_[19223]_ ;
  assign \new_[19233]_  = A236 & A233;
  assign \new_[19234]_  = ~A232 & \new_[19233]_ ;
  assign \new_[19238]_  = ~A302 & ~A301;
  assign \new_[19239]_  = ~A300 & \new_[19238]_ ;
  assign \new_[19240]_  = \new_[19239]_  & \new_[19234]_ ;
  assign \new_[19243]_  = A167 & A168;
  assign \new_[19247]_  = ~A202 & ~A200;
  assign \new_[19248]_  = ~A199 & \new_[19247]_ ;
  assign \new_[19249]_  = \new_[19248]_  & \new_[19243]_ ;
  assign \new_[19253]_  = A236 & A233;
  assign \new_[19254]_  = ~A232 & \new_[19253]_ ;
  assign \new_[19258]_  = ~A301 & ~A299;
  assign \new_[19259]_  = ~A298 & \new_[19258]_ ;
  assign \new_[19260]_  = \new_[19259]_  & \new_[19254]_ ;
  assign \new_[19263]_  = A167 & A168;
  assign \new_[19267]_  = ~A202 & ~A200;
  assign \new_[19268]_  = ~A199 & \new_[19267]_ ;
  assign \new_[19269]_  = \new_[19268]_  & \new_[19263]_ ;
  assign \new_[19273]_  = A236 & A233;
  assign \new_[19274]_  = ~A232 & \new_[19273]_ ;
  assign \new_[19278]_  = A269 & A266;
  assign \new_[19279]_  = ~A265 & \new_[19278]_ ;
  assign \new_[19280]_  = \new_[19279]_  & \new_[19274]_ ;
  assign \new_[19283]_  = A167 & A168;
  assign \new_[19287]_  = ~A202 & ~A200;
  assign \new_[19288]_  = ~A199 & \new_[19287]_ ;
  assign \new_[19289]_  = \new_[19288]_  & \new_[19283]_ ;
  assign \new_[19293]_  = A236 & A233;
  assign \new_[19294]_  = ~A232 & \new_[19293]_ ;
  assign \new_[19298]_  = A269 & ~A266;
  assign \new_[19299]_  = A265 & \new_[19298]_ ;
  assign \new_[19300]_  = \new_[19299]_  & \new_[19294]_ ;
  assign \new_[19303]_  = A167 & A168;
  assign \new_[19307]_  = ~A202 & ~A200;
  assign \new_[19308]_  = ~A199 & \new_[19307]_ ;
  assign \new_[19309]_  = \new_[19308]_  & \new_[19303]_ ;
  assign \new_[19313]_  = A236 & ~A233;
  assign \new_[19314]_  = A232 & \new_[19313]_ ;
  assign \new_[19318]_  = ~A302 & ~A301;
  assign \new_[19319]_  = ~A300 & \new_[19318]_ ;
  assign \new_[19320]_  = \new_[19319]_  & \new_[19314]_ ;
  assign \new_[19323]_  = A167 & A168;
  assign \new_[19327]_  = ~A202 & ~A200;
  assign \new_[19328]_  = ~A199 & \new_[19327]_ ;
  assign \new_[19329]_  = \new_[19328]_  & \new_[19323]_ ;
  assign \new_[19333]_  = A236 & ~A233;
  assign \new_[19334]_  = A232 & \new_[19333]_ ;
  assign \new_[19338]_  = ~A301 & ~A299;
  assign \new_[19339]_  = ~A298 & \new_[19338]_ ;
  assign \new_[19340]_  = \new_[19339]_  & \new_[19334]_ ;
  assign \new_[19343]_  = A167 & A168;
  assign \new_[19347]_  = ~A202 & ~A200;
  assign \new_[19348]_  = ~A199 & \new_[19347]_ ;
  assign \new_[19349]_  = \new_[19348]_  & \new_[19343]_ ;
  assign \new_[19353]_  = A236 & ~A233;
  assign \new_[19354]_  = A232 & \new_[19353]_ ;
  assign \new_[19358]_  = A269 & A266;
  assign \new_[19359]_  = ~A265 & \new_[19358]_ ;
  assign \new_[19360]_  = \new_[19359]_  & \new_[19354]_ ;
  assign \new_[19363]_  = A167 & A168;
  assign \new_[19367]_  = ~A202 & ~A200;
  assign \new_[19368]_  = ~A199 & \new_[19367]_ ;
  assign \new_[19369]_  = \new_[19368]_  & \new_[19363]_ ;
  assign \new_[19373]_  = A236 & ~A233;
  assign \new_[19374]_  = A232 & \new_[19373]_ ;
  assign \new_[19378]_  = A269 & ~A266;
  assign \new_[19379]_  = A265 & \new_[19378]_ ;
  assign \new_[19380]_  = \new_[19379]_  & \new_[19374]_ ;
  assign \new_[19383]_  = A167 & A170;
  assign \new_[19387]_  = ~A202 & ~A201;
  assign \new_[19388]_  = ~A166 & \new_[19387]_ ;
  assign \new_[19389]_  = \new_[19388]_  & \new_[19383]_ ;
  assign \new_[19393]_  = A298 & A235;
  assign \new_[19394]_  = ~A203 & \new_[19393]_ ;
  assign \new_[19398]_  = ~A301 & ~A300;
  assign \new_[19399]_  = A299 & \new_[19398]_ ;
  assign \new_[19400]_  = \new_[19399]_  & \new_[19394]_ ;
  assign \new_[19403]_  = A167 & A170;
  assign \new_[19407]_  = ~A202 & ~A201;
  assign \new_[19408]_  = ~A166 & \new_[19407]_ ;
  assign \new_[19409]_  = \new_[19408]_  & \new_[19403]_ ;
  assign \new_[19413]_  = A234 & A232;
  assign \new_[19414]_  = ~A203 & \new_[19413]_ ;
  assign \new_[19418]_  = ~A302 & ~A301;
  assign \new_[19419]_  = ~A300 & \new_[19418]_ ;
  assign \new_[19420]_  = \new_[19419]_  & \new_[19414]_ ;
  assign \new_[19423]_  = A167 & A170;
  assign \new_[19427]_  = ~A202 & ~A201;
  assign \new_[19428]_  = ~A166 & \new_[19427]_ ;
  assign \new_[19429]_  = \new_[19428]_  & \new_[19423]_ ;
  assign \new_[19433]_  = A234 & A232;
  assign \new_[19434]_  = ~A203 & \new_[19433]_ ;
  assign \new_[19438]_  = ~A301 & ~A299;
  assign \new_[19439]_  = ~A298 & \new_[19438]_ ;
  assign \new_[19440]_  = \new_[19439]_  & \new_[19434]_ ;
  assign \new_[19443]_  = A167 & A170;
  assign \new_[19447]_  = ~A202 & ~A201;
  assign \new_[19448]_  = ~A166 & \new_[19447]_ ;
  assign \new_[19449]_  = \new_[19448]_  & \new_[19443]_ ;
  assign \new_[19453]_  = A234 & A232;
  assign \new_[19454]_  = ~A203 & \new_[19453]_ ;
  assign \new_[19458]_  = A269 & A266;
  assign \new_[19459]_  = ~A265 & \new_[19458]_ ;
  assign \new_[19460]_  = \new_[19459]_  & \new_[19454]_ ;
  assign \new_[19463]_  = A167 & A170;
  assign \new_[19467]_  = ~A202 & ~A201;
  assign \new_[19468]_  = ~A166 & \new_[19467]_ ;
  assign \new_[19469]_  = \new_[19468]_  & \new_[19463]_ ;
  assign \new_[19473]_  = A234 & A232;
  assign \new_[19474]_  = ~A203 & \new_[19473]_ ;
  assign \new_[19478]_  = A269 & ~A266;
  assign \new_[19479]_  = A265 & \new_[19478]_ ;
  assign \new_[19480]_  = \new_[19479]_  & \new_[19474]_ ;
  assign \new_[19483]_  = A167 & A170;
  assign \new_[19487]_  = ~A202 & ~A201;
  assign \new_[19488]_  = ~A166 & \new_[19487]_ ;
  assign \new_[19489]_  = \new_[19488]_  & \new_[19483]_ ;
  assign \new_[19493]_  = A234 & A233;
  assign \new_[19494]_  = ~A203 & \new_[19493]_ ;
  assign \new_[19498]_  = ~A302 & ~A301;
  assign \new_[19499]_  = ~A300 & \new_[19498]_ ;
  assign \new_[19500]_  = \new_[19499]_  & \new_[19494]_ ;
  assign \new_[19503]_  = A167 & A170;
  assign \new_[19507]_  = ~A202 & ~A201;
  assign \new_[19508]_  = ~A166 & \new_[19507]_ ;
  assign \new_[19509]_  = \new_[19508]_  & \new_[19503]_ ;
  assign \new_[19513]_  = A234 & A233;
  assign \new_[19514]_  = ~A203 & \new_[19513]_ ;
  assign \new_[19518]_  = ~A301 & ~A299;
  assign \new_[19519]_  = ~A298 & \new_[19518]_ ;
  assign \new_[19520]_  = \new_[19519]_  & \new_[19514]_ ;
  assign \new_[19523]_  = A167 & A170;
  assign \new_[19527]_  = ~A202 & ~A201;
  assign \new_[19528]_  = ~A166 & \new_[19527]_ ;
  assign \new_[19529]_  = \new_[19528]_  & \new_[19523]_ ;
  assign \new_[19533]_  = A234 & A233;
  assign \new_[19534]_  = ~A203 & \new_[19533]_ ;
  assign \new_[19538]_  = A269 & A266;
  assign \new_[19539]_  = ~A265 & \new_[19538]_ ;
  assign \new_[19540]_  = \new_[19539]_  & \new_[19534]_ ;
  assign \new_[19543]_  = A167 & A170;
  assign \new_[19547]_  = ~A202 & ~A201;
  assign \new_[19548]_  = ~A166 & \new_[19547]_ ;
  assign \new_[19549]_  = \new_[19548]_  & \new_[19543]_ ;
  assign \new_[19553]_  = A234 & A233;
  assign \new_[19554]_  = ~A203 & \new_[19553]_ ;
  assign \new_[19558]_  = A269 & ~A266;
  assign \new_[19559]_  = A265 & \new_[19558]_ ;
  assign \new_[19560]_  = \new_[19559]_  & \new_[19554]_ ;
  assign \new_[19563]_  = A167 & A170;
  assign \new_[19567]_  = ~A202 & ~A201;
  assign \new_[19568]_  = ~A166 & \new_[19567]_ ;
  assign \new_[19569]_  = \new_[19568]_  & \new_[19563]_ ;
  assign \new_[19573]_  = A233 & ~A232;
  assign \new_[19574]_  = ~A203 & \new_[19573]_ ;
  assign \new_[19578]_  = A267 & A265;
  assign \new_[19579]_  = A236 & \new_[19578]_ ;
  assign \new_[19580]_  = \new_[19579]_  & \new_[19574]_ ;
  assign \new_[19583]_  = A167 & A170;
  assign \new_[19587]_  = ~A202 & ~A201;
  assign \new_[19588]_  = ~A166 & \new_[19587]_ ;
  assign \new_[19589]_  = \new_[19588]_  & \new_[19583]_ ;
  assign \new_[19593]_  = A233 & ~A232;
  assign \new_[19594]_  = ~A203 & \new_[19593]_ ;
  assign \new_[19598]_  = A267 & A266;
  assign \new_[19599]_  = A236 & \new_[19598]_ ;
  assign \new_[19600]_  = \new_[19599]_  & \new_[19594]_ ;
  assign \new_[19603]_  = A167 & A170;
  assign \new_[19607]_  = ~A202 & ~A201;
  assign \new_[19608]_  = ~A166 & \new_[19607]_ ;
  assign \new_[19609]_  = \new_[19608]_  & \new_[19603]_ ;
  assign \new_[19613]_  = ~A233 & A232;
  assign \new_[19614]_  = ~A203 & \new_[19613]_ ;
  assign \new_[19618]_  = A267 & A265;
  assign \new_[19619]_  = A236 & \new_[19618]_ ;
  assign \new_[19620]_  = \new_[19619]_  & \new_[19614]_ ;
  assign \new_[19623]_  = A167 & A170;
  assign \new_[19627]_  = ~A202 & ~A201;
  assign \new_[19628]_  = ~A166 & \new_[19627]_ ;
  assign \new_[19629]_  = \new_[19628]_  & \new_[19623]_ ;
  assign \new_[19633]_  = ~A233 & A232;
  assign \new_[19634]_  = ~A203 & \new_[19633]_ ;
  assign \new_[19638]_  = A267 & A266;
  assign \new_[19639]_  = A236 & \new_[19638]_ ;
  assign \new_[19640]_  = \new_[19639]_  & \new_[19634]_ ;
  assign \new_[19643]_  = A167 & A170;
  assign \new_[19647]_  = A200 & A199;
  assign \new_[19648]_  = ~A166 & \new_[19647]_ ;
  assign \new_[19649]_  = \new_[19648]_  & \new_[19643]_ ;
  assign \new_[19653]_  = A235 & ~A202;
  assign \new_[19654]_  = ~A201 & \new_[19653]_ ;
  assign \new_[19658]_  = ~A302 & ~A301;
  assign \new_[19659]_  = ~A300 & \new_[19658]_ ;
  assign \new_[19660]_  = \new_[19659]_  & \new_[19654]_ ;
  assign \new_[19663]_  = A167 & A170;
  assign \new_[19667]_  = A200 & A199;
  assign \new_[19668]_  = ~A166 & \new_[19667]_ ;
  assign \new_[19669]_  = \new_[19668]_  & \new_[19663]_ ;
  assign \new_[19673]_  = A235 & ~A202;
  assign \new_[19674]_  = ~A201 & \new_[19673]_ ;
  assign \new_[19678]_  = ~A301 & ~A299;
  assign \new_[19679]_  = ~A298 & \new_[19678]_ ;
  assign \new_[19680]_  = \new_[19679]_  & \new_[19674]_ ;
  assign \new_[19683]_  = A167 & A170;
  assign \new_[19687]_  = A200 & A199;
  assign \new_[19688]_  = ~A166 & \new_[19687]_ ;
  assign \new_[19689]_  = \new_[19688]_  & \new_[19683]_ ;
  assign \new_[19693]_  = A235 & ~A202;
  assign \new_[19694]_  = ~A201 & \new_[19693]_ ;
  assign \new_[19698]_  = A269 & A266;
  assign \new_[19699]_  = ~A265 & \new_[19698]_ ;
  assign \new_[19700]_  = \new_[19699]_  & \new_[19694]_ ;
  assign \new_[19703]_  = A167 & A170;
  assign \new_[19707]_  = A200 & A199;
  assign \new_[19708]_  = ~A166 & \new_[19707]_ ;
  assign \new_[19709]_  = \new_[19708]_  & \new_[19703]_ ;
  assign \new_[19713]_  = A235 & ~A202;
  assign \new_[19714]_  = ~A201 & \new_[19713]_ ;
  assign \new_[19718]_  = A269 & ~A266;
  assign \new_[19719]_  = A265 & \new_[19718]_ ;
  assign \new_[19720]_  = \new_[19719]_  & \new_[19714]_ ;
  assign \new_[19723]_  = A167 & A170;
  assign \new_[19727]_  = A200 & A199;
  assign \new_[19728]_  = ~A166 & \new_[19727]_ ;
  assign \new_[19729]_  = \new_[19728]_  & \new_[19723]_ ;
  assign \new_[19733]_  = A232 & ~A202;
  assign \new_[19734]_  = ~A201 & \new_[19733]_ ;
  assign \new_[19738]_  = A267 & A265;
  assign \new_[19739]_  = A234 & \new_[19738]_ ;
  assign \new_[19740]_  = \new_[19739]_  & \new_[19734]_ ;
  assign \new_[19743]_  = A167 & A170;
  assign \new_[19747]_  = A200 & A199;
  assign \new_[19748]_  = ~A166 & \new_[19747]_ ;
  assign \new_[19749]_  = \new_[19748]_  & \new_[19743]_ ;
  assign \new_[19753]_  = A232 & ~A202;
  assign \new_[19754]_  = ~A201 & \new_[19753]_ ;
  assign \new_[19758]_  = A267 & A266;
  assign \new_[19759]_  = A234 & \new_[19758]_ ;
  assign \new_[19760]_  = \new_[19759]_  & \new_[19754]_ ;
  assign \new_[19763]_  = A167 & A170;
  assign \new_[19767]_  = A200 & A199;
  assign \new_[19768]_  = ~A166 & \new_[19767]_ ;
  assign \new_[19769]_  = \new_[19768]_  & \new_[19763]_ ;
  assign \new_[19773]_  = A233 & ~A202;
  assign \new_[19774]_  = ~A201 & \new_[19773]_ ;
  assign \new_[19778]_  = A267 & A265;
  assign \new_[19779]_  = A234 & \new_[19778]_ ;
  assign \new_[19780]_  = \new_[19779]_  & \new_[19774]_ ;
  assign \new_[19783]_  = A167 & A170;
  assign \new_[19787]_  = A200 & A199;
  assign \new_[19788]_  = ~A166 & \new_[19787]_ ;
  assign \new_[19789]_  = \new_[19788]_  & \new_[19783]_ ;
  assign \new_[19793]_  = A233 & ~A202;
  assign \new_[19794]_  = ~A201 & \new_[19793]_ ;
  assign \new_[19798]_  = A267 & A266;
  assign \new_[19799]_  = A234 & \new_[19798]_ ;
  assign \new_[19800]_  = \new_[19799]_  & \new_[19794]_ ;
  assign \new_[19803]_  = A167 & A170;
  assign \new_[19807]_  = A200 & A199;
  assign \new_[19808]_  = ~A166 & \new_[19807]_ ;
  assign \new_[19809]_  = \new_[19808]_  & \new_[19803]_ ;
  assign \new_[19813]_  = ~A232 & ~A202;
  assign \new_[19814]_  = ~A201 & \new_[19813]_ ;
  assign \new_[19818]_  = A268 & A236;
  assign \new_[19819]_  = A233 & \new_[19818]_ ;
  assign \new_[19820]_  = \new_[19819]_  & \new_[19814]_ ;
  assign \new_[19823]_  = A167 & A170;
  assign \new_[19827]_  = A200 & A199;
  assign \new_[19828]_  = ~A166 & \new_[19827]_ ;
  assign \new_[19829]_  = \new_[19828]_  & \new_[19823]_ ;
  assign \new_[19833]_  = A232 & ~A202;
  assign \new_[19834]_  = ~A201 & \new_[19833]_ ;
  assign \new_[19838]_  = A268 & A236;
  assign \new_[19839]_  = ~A233 & \new_[19838]_ ;
  assign \new_[19840]_  = \new_[19839]_  & \new_[19834]_ ;
  assign \new_[19843]_  = A167 & A170;
  assign \new_[19847]_  = ~A200 & ~A199;
  assign \new_[19848]_  = ~A166 & \new_[19847]_ ;
  assign \new_[19849]_  = \new_[19848]_  & \new_[19843]_ ;
  assign \new_[19853]_  = A298 & A235;
  assign \new_[19854]_  = ~A202 & \new_[19853]_ ;
  assign \new_[19858]_  = ~A301 & ~A300;
  assign \new_[19859]_  = A299 & \new_[19858]_ ;
  assign \new_[19860]_  = \new_[19859]_  & \new_[19854]_ ;
  assign \new_[19863]_  = A167 & A170;
  assign \new_[19867]_  = ~A200 & ~A199;
  assign \new_[19868]_  = ~A166 & \new_[19867]_ ;
  assign \new_[19869]_  = \new_[19868]_  & \new_[19863]_ ;
  assign \new_[19873]_  = A234 & A232;
  assign \new_[19874]_  = ~A202 & \new_[19873]_ ;
  assign \new_[19878]_  = ~A302 & ~A301;
  assign \new_[19879]_  = ~A300 & \new_[19878]_ ;
  assign \new_[19880]_  = \new_[19879]_  & \new_[19874]_ ;
  assign \new_[19883]_  = A167 & A170;
  assign \new_[19887]_  = ~A200 & ~A199;
  assign \new_[19888]_  = ~A166 & \new_[19887]_ ;
  assign \new_[19889]_  = \new_[19888]_  & \new_[19883]_ ;
  assign \new_[19893]_  = A234 & A232;
  assign \new_[19894]_  = ~A202 & \new_[19893]_ ;
  assign \new_[19898]_  = ~A301 & ~A299;
  assign \new_[19899]_  = ~A298 & \new_[19898]_ ;
  assign \new_[19900]_  = \new_[19899]_  & \new_[19894]_ ;
  assign \new_[19903]_  = A167 & A170;
  assign \new_[19907]_  = ~A200 & ~A199;
  assign \new_[19908]_  = ~A166 & \new_[19907]_ ;
  assign \new_[19909]_  = \new_[19908]_  & \new_[19903]_ ;
  assign \new_[19913]_  = A234 & A232;
  assign \new_[19914]_  = ~A202 & \new_[19913]_ ;
  assign \new_[19918]_  = A269 & A266;
  assign \new_[19919]_  = ~A265 & \new_[19918]_ ;
  assign \new_[19920]_  = \new_[19919]_  & \new_[19914]_ ;
  assign \new_[19923]_  = A167 & A170;
  assign \new_[19927]_  = ~A200 & ~A199;
  assign \new_[19928]_  = ~A166 & \new_[19927]_ ;
  assign \new_[19929]_  = \new_[19928]_  & \new_[19923]_ ;
  assign \new_[19933]_  = A234 & A232;
  assign \new_[19934]_  = ~A202 & \new_[19933]_ ;
  assign \new_[19938]_  = A269 & ~A266;
  assign \new_[19939]_  = A265 & \new_[19938]_ ;
  assign \new_[19940]_  = \new_[19939]_  & \new_[19934]_ ;
  assign \new_[19943]_  = A167 & A170;
  assign \new_[19947]_  = ~A200 & ~A199;
  assign \new_[19948]_  = ~A166 & \new_[19947]_ ;
  assign \new_[19949]_  = \new_[19948]_  & \new_[19943]_ ;
  assign \new_[19953]_  = A234 & A233;
  assign \new_[19954]_  = ~A202 & \new_[19953]_ ;
  assign \new_[19958]_  = ~A302 & ~A301;
  assign \new_[19959]_  = ~A300 & \new_[19958]_ ;
  assign \new_[19960]_  = \new_[19959]_  & \new_[19954]_ ;
  assign \new_[19963]_  = A167 & A170;
  assign \new_[19967]_  = ~A200 & ~A199;
  assign \new_[19968]_  = ~A166 & \new_[19967]_ ;
  assign \new_[19969]_  = \new_[19968]_  & \new_[19963]_ ;
  assign \new_[19973]_  = A234 & A233;
  assign \new_[19974]_  = ~A202 & \new_[19973]_ ;
  assign \new_[19978]_  = ~A301 & ~A299;
  assign \new_[19979]_  = ~A298 & \new_[19978]_ ;
  assign \new_[19980]_  = \new_[19979]_  & \new_[19974]_ ;
  assign \new_[19983]_  = A167 & A170;
  assign \new_[19987]_  = ~A200 & ~A199;
  assign \new_[19988]_  = ~A166 & \new_[19987]_ ;
  assign \new_[19989]_  = \new_[19988]_  & \new_[19983]_ ;
  assign \new_[19993]_  = A234 & A233;
  assign \new_[19994]_  = ~A202 & \new_[19993]_ ;
  assign \new_[19998]_  = A269 & A266;
  assign \new_[19999]_  = ~A265 & \new_[19998]_ ;
  assign \new_[20000]_  = \new_[19999]_  & \new_[19994]_ ;
  assign \new_[20003]_  = A167 & A170;
  assign \new_[20007]_  = ~A200 & ~A199;
  assign \new_[20008]_  = ~A166 & \new_[20007]_ ;
  assign \new_[20009]_  = \new_[20008]_  & \new_[20003]_ ;
  assign \new_[20013]_  = A234 & A233;
  assign \new_[20014]_  = ~A202 & \new_[20013]_ ;
  assign \new_[20018]_  = A269 & ~A266;
  assign \new_[20019]_  = A265 & \new_[20018]_ ;
  assign \new_[20020]_  = \new_[20019]_  & \new_[20014]_ ;
  assign \new_[20023]_  = A167 & A170;
  assign \new_[20027]_  = ~A200 & ~A199;
  assign \new_[20028]_  = ~A166 & \new_[20027]_ ;
  assign \new_[20029]_  = \new_[20028]_  & \new_[20023]_ ;
  assign \new_[20033]_  = A233 & ~A232;
  assign \new_[20034]_  = ~A202 & \new_[20033]_ ;
  assign \new_[20038]_  = A267 & A265;
  assign \new_[20039]_  = A236 & \new_[20038]_ ;
  assign \new_[20040]_  = \new_[20039]_  & \new_[20034]_ ;
  assign \new_[20043]_  = A167 & A170;
  assign \new_[20047]_  = ~A200 & ~A199;
  assign \new_[20048]_  = ~A166 & \new_[20047]_ ;
  assign \new_[20049]_  = \new_[20048]_  & \new_[20043]_ ;
  assign \new_[20053]_  = A233 & ~A232;
  assign \new_[20054]_  = ~A202 & \new_[20053]_ ;
  assign \new_[20058]_  = A267 & A266;
  assign \new_[20059]_  = A236 & \new_[20058]_ ;
  assign \new_[20060]_  = \new_[20059]_  & \new_[20054]_ ;
  assign \new_[20063]_  = A167 & A170;
  assign \new_[20067]_  = ~A200 & ~A199;
  assign \new_[20068]_  = ~A166 & \new_[20067]_ ;
  assign \new_[20069]_  = \new_[20068]_  & \new_[20063]_ ;
  assign \new_[20073]_  = ~A233 & A232;
  assign \new_[20074]_  = ~A202 & \new_[20073]_ ;
  assign \new_[20078]_  = A267 & A265;
  assign \new_[20079]_  = A236 & \new_[20078]_ ;
  assign \new_[20080]_  = \new_[20079]_  & \new_[20074]_ ;
  assign \new_[20083]_  = A167 & A170;
  assign \new_[20087]_  = ~A200 & ~A199;
  assign \new_[20088]_  = ~A166 & \new_[20087]_ ;
  assign \new_[20089]_  = \new_[20088]_  & \new_[20083]_ ;
  assign \new_[20093]_  = ~A233 & A232;
  assign \new_[20094]_  = ~A202 & \new_[20093]_ ;
  assign \new_[20098]_  = A267 & A266;
  assign \new_[20099]_  = A236 & \new_[20098]_ ;
  assign \new_[20100]_  = \new_[20099]_  & \new_[20094]_ ;
  assign \new_[20103]_  = ~A167 & A170;
  assign \new_[20107]_  = ~A202 & ~A201;
  assign \new_[20108]_  = A166 & \new_[20107]_ ;
  assign \new_[20109]_  = \new_[20108]_  & \new_[20103]_ ;
  assign \new_[20113]_  = A298 & A235;
  assign \new_[20114]_  = ~A203 & \new_[20113]_ ;
  assign \new_[20118]_  = ~A301 & ~A300;
  assign \new_[20119]_  = A299 & \new_[20118]_ ;
  assign \new_[20120]_  = \new_[20119]_  & \new_[20114]_ ;
  assign \new_[20123]_  = ~A167 & A170;
  assign \new_[20127]_  = ~A202 & ~A201;
  assign \new_[20128]_  = A166 & \new_[20127]_ ;
  assign \new_[20129]_  = \new_[20128]_  & \new_[20123]_ ;
  assign \new_[20133]_  = A234 & A232;
  assign \new_[20134]_  = ~A203 & \new_[20133]_ ;
  assign \new_[20138]_  = ~A302 & ~A301;
  assign \new_[20139]_  = ~A300 & \new_[20138]_ ;
  assign \new_[20140]_  = \new_[20139]_  & \new_[20134]_ ;
  assign \new_[20143]_  = ~A167 & A170;
  assign \new_[20147]_  = ~A202 & ~A201;
  assign \new_[20148]_  = A166 & \new_[20147]_ ;
  assign \new_[20149]_  = \new_[20148]_  & \new_[20143]_ ;
  assign \new_[20153]_  = A234 & A232;
  assign \new_[20154]_  = ~A203 & \new_[20153]_ ;
  assign \new_[20158]_  = ~A301 & ~A299;
  assign \new_[20159]_  = ~A298 & \new_[20158]_ ;
  assign \new_[20160]_  = \new_[20159]_  & \new_[20154]_ ;
  assign \new_[20163]_  = ~A167 & A170;
  assign \new_[20167]_  = ~A202 & ~A201;
  assign \new_[20168]_  = A166 & \new_[20167]_ ;
  assign \new_[20169]_  = \new_[20168]_  & \new_[20163]_ ;
  assign \new_[20173]_  = A234 & A232;
  assign \new_[20174]_  = ~A203 & \new_[20173]_ ;
  assign \new_[20178]_  = A269 & A266;
  assign \new_[20179]_  = ~A265 & \new_[20178]_ ;
  assign \new_[20180]_  = \new_[20179]_  & \new_[20174]_ ;
  assign \new_[20183]_  = ~A167 & A170;
  assign \new_[20187]_  = ~A202 & ~A201;
  assign \new_[20188]_  = A166 & \new_[20187]_ ;
  assign \new_[20189]_  = \new_[20188]_  & \new_[20183]_ ;
  assign \new_[20193]_  = A234 & A232;
  assign \new_[20194]_  = ~A203 & \new_[20193]_ ;
  assign \new_[20198]_  = A269 & ~A266;
  assign \new_[20199]_  = A265 & \new_[20198]_ ;
  assign \new_[20200]_  = \new_[20199]_  & \new_[20194]_ ;
  assign \new_[20203]_  = ~A167 & A170;
  assign \new_[20207]_  = ~A202 & ~A201;
  assign \new_[20208]_  = A166 & \new_[20207]_ ;
  assign \new_[20209]_  = \new_[20208]_  & \new_[20203]_ ;
  assign \new_[20213]_  = A234 & A233;
  assign \new_[20214]_  = ~A203 & \new_[20213]_ ;
  assign \new_[20218]_  = ~A302 & ~A301;
  assign \new_[20219]_  = ~A300 & \new_[20218]_ ;
  assign \new_[20220]_  = \new_[20219]_  & \new_[20214]_ ;
  assign \new_[20223]_  = ~A167 & A170;
  assign \new_[20227]_  = ~A202 & ~A201;
  assign \new_[20228]_  = A166 & \new_[20227]_ ;
  assign \new_[20229]_  = \new_[20228]_  & \new_[20223]_ ;
  assign \new_[20233]_  = A234 & A233;
  assign \new_[20234]_  = ~A203 & \new_[20233]_ ;
  assign \new_[20238]_  = ~A301 & ~A299;
  assign \new_[20239]_  = ~A298 & \new_[20238]_ ;
  assign \new_[20240]_  = \new_[20239]_  & \new_[20234]_ ;
  assign \new_[20243]_  = ~A167 & A170;
  assign \new_[20247]_  = ~A202 & ~A201;
  assign \new_[20248]_  = A166 & \new_[20247]_ ;
  assign \new_[20249]_  = \new_[20248]_  & \new_[20243]_ ;
  assign \new_[20253]_  = A234 & A233;
  assign \new_[20254]_  = ~A203 & \new_[20253]_ ;
  assign \new_[20258]_  = A269 & A266;
  assign \new_[20259]_  = ~A265 & \new_[20258]_ ;
  assign \new_[20260]_  = \new_[20259]_  & \new_[20254]_ ;
  assign \new_[20263]_  = ~A167 & A170;
  assign \new_[20267]_  = ~A202 & ~A201;
  assign \new_[20268]_  = A166 & \new_[20267]_ ;
  assign \new_[20269]_  = \new_[20268]_  & \new_[20263]_ ;
  assign \new_[20273]_  = A234 & A233;
  assign \new_[20274]_  = ~A203 & \new_[20273]_ ;
  assign \new_[20278]_  = A269 & ~A266;
  assign \new_[20279]_  = A265 & \new_[20278]_ ;
  assign \new_[20280]_  = \new_[20279]_  & \new_[20274]_ ;
  assign \new_[20283]_  = ~A167 & A170;
  assign \new_[20287]_  = ~A202 & ~A201;
  assign \new_[20288]_  = A166 & \new_[20287]_ ;
  assign \new_[20289]_  = \new_[20288]_  & \new_[20283]_ ;
  assign \new_[20293]_  = A233 & ~A232;
  assign \new_[20294]_  = ~A203 & \new_[20293]_ ;
  assign \new_[20298]_  = A267 & A265;
  assign \new_[20299]_  = A236 & \new_[20298]_ ;
  assign \new_[20300]_  = \new_[20299]_  & \new_[20294]_ ;
  assign \new_[20303]_  = ~A167 & A170;
  assign \new_[20307]_  = ~A202 & ~A201;
  assign \new_[20308]_  = A166 & \new_[20307]_ ;
  assign \new_[20309]_  = \new_[20308]_  & \new_[20303]_ ;
  assign \new_[20313]_  = A233 & ~A232;
  assign \new_[20314]_  = ~A203 & \new_[20313]_ ;
  assign \new_[20318]_  = A267 & A266;
  assign \new_[20319]_  = A236 & \new_[20318]_ ;
  assign \new_[20320]_  = \new_[20319]_  & \new_[20314]_ ;
  assign \new_[20323]_  = ~A167 & A170;
  assign \new_[20327]_  = ~A202 & ~A201;
  assign \new_[20328]_  = A166 & \new_[20327]_ ;
  assign \new_[20329]_  = \new_[20328]_  & \new_[20323]_ ;
  assign \new_[20333]_  = ~A233 & A232;
  assign \new_[20334]_  = ~A203 & \new_[20333]_ ;
  assign \new_[20338]_  = A267 & A265;
  assign \new_[20339]_  = A236 & \new_[20338]_ ;
  assign \new_[20340]_  = \new_[20339]_  & \new_[20334]_ ;
  assign \new_[20343]_  = ~A167 & A170;
  assign \new_[20347]_  = ~A202 & ~A201;
  assign \new_[20348]_  = A166 & \new_[20347]_ ;
  assign \new_[20349]_  = \new_[20348]_  & \new_[20343]_ ;
  assign \new_[20353]_  = ~A233 & A232;
  assign \new_[20354]_  = ~A203 & \new_[20353]_ ;
  assign \new_[20358]_  = A267 & A266;
  assign \new_[20359]_  = A236 & \new_[20358]_ ;
  assign \new_[20360]_  = \new_[20359]_  & \new_[20354]_ ;
  assign \new_[20363]_  = ~A167 & A170;
  assign \new_[20367]_  = A200 & A199;
  assign \new_[20368]_  = A166 & \new_[20367]_ ;
  assign \new_[20369]_  = \new_[20368]_  & \new_[20363]_ ;
  assign \new_[20373]_  = A235 & ~A202;
  assign \new_[20374]_  = ~A201 & \new_[20373]_ ;
  assign \new_[20378]_  = ~A302 & ~A301;
  assign \new_[20379]_  = ~A300 & \new_[20378]_ ;
  assign \new_[20380]_  = \new_[20379]_  & \new_[20374]_ ;
  assign \new_[20383]_  = ~A167 & A170;
  assign \new_[20387]_  = A200 & A199;
  assign \new_[20388]_  = A166 & \new_[20387]_ ;
  assign \new_[20389]_  = \new_[20388]_  & \new_[20383]_ ;
  assign \new_[20393]_  = A235 & ~A202;
  assign \new_[20394]_  = ~A201 & \new_[20393]_ ;
  assign \new_[20398]_  = ~A301 & ~A299;
  assign \new_[20399]_  = ~A298 & \new_[20398]_ ;
  assign \new_[20400]_  = \new_[20399]_  & \new_[20394]_ ;
  assign \new_[20403]_  = ~A167 & A170;
  assign \new_[20407]_  = A200 & A199;
  assign \new_[20408]_  = A166 & \new_[20407]_ ;
  assign \new_[20409]_  = \new_[20408]_  & \new_[20403]_ ;
  assign \new_[20413]_  = A235 & ~A202;
  assign \new_[20414]_  = ~A201 & \new_[20413]_ ;
  assign \new_[20418]_  = A269 & A266;
  assign \new_[20419]_  = ~A265 & \new_[20418]_ ;
  assign \new_[20420]_  = \new_[20419]_  & \new_[20414]_ ;
  assign \new_[20423]_  = ~A167 & A170;
  assign \new_[20427]_  = A200 & A199;
  assign \new_[20428]_  = A166 & \new_[20427]_ ;
  assign \new_[20429]_  = \new_[20428]_  & \new_[20423]_ ;
  assign \new_[20433]_  = A235 & ~A202;
  assign \new_[20434]_  = ~A201 & \new_[20433]_ ;
  assign \new_[20438]_  = A269 & ~A266;
  assign \new_[20439]_  = A265 & \new_[20438]_ ;
  assign \new_[20440]_  = \new_[20439]_  & \new_[20434]_ ;
  assign \new_[20443]_  = ~A167 & A170;
  assign \new_[20447]_  = A200 & A199;
  assign \new_[20448]_  = A166 & \new_[20447]_ ;
  assign \new_[20449]_  = \new_[20448]_  & \new_[20443]_ ;
  assign \new_[20453]_  = A232 & ~A202;
  assign \new_[20454]_  = ~A201 & \new_[20453]_ ;
  assign \new_[20458]_  = A267 & A265;
  assign \new_[20459]_  = A234 & \new_[20458]_ ;
  assign \new_[20460]_  = \new_[20459]_  & \new_[20454]_ ;
  assign \new_[20463]_  = ~A167 & A170;
  assign \new_[20467]_  = A200 & A199;
  assign \new_[20468]_  = A166 & \new_[20467]_ ;
  assign \new_[20469]_  = \new_[20468]_  & \new_[20463]_ ;
  assign \new_[20473]_  = A232 & ~A202;
  assign \new_[20474]_  = ~A201 & \new_[20473]_ ;
  assign \new_[20478]_  = A267 & A266;
  assign \new_[20479]_  = A234 & \new_[20478]_ ;
  assign \new_[20480]_  = \new_[20479]_  & \new_[20474]_ ;
  assign \new_[20483]_  = ~A167 & A170;
  assign \new_[20487]_  = A200 & A199;
  assign \new_[20488]_  = A166 & \new_[20487]_ ;
  assign \new_[20489]_  = \new_[20488]_  & \new_[20483]_ ;
  assign \new_[20493]_  = A233 & ~A202;
  assign \new_[20494]_  = ~A201 & \new_[20493]_ ;
  assign \new_[20498]_  = A267 & A265;
  assign \new_[20499]_  = A234 & \new_[20498]_ ;
  assign \new_[20500]_  = \new_[20499]_  & \new_[20494]_ ;
  assign \new_[20503]_  = ~A167 & A170;
  assign \new_[20507]_  = A200 & A199;
  assign \new_[20508]_  = A166 & \new_[20507]_ ;
  assign \new_[20509]_  = \new_[20508]_  & \new_[20503]_ ;
  assign \new_[20513]_  = A233 & ~A202;
  assign \new_[20514]_  = ~A201 & \new_[20513]_ ;
  assign \new_[20518]_  = A267 & A266;
  assign \new_[20519]_  = A234 & \new_[20518]_ ;
  assign \new_[20520]_  = \new_[20519]_  & \new_[20514]_ ;
  assign \new_[20523]_  = ~A167 & A170;
  assign \new_[20527]_  = A200 & A199;
  assign \new_[20528]_  = A166 & \new_[20527]_ ;
  assign \new_[20529]_  = \new_[20528]_  & \new_[20523]_ ;
  assign \new_[20533]_  = ~A232 & ~A202;
  assign \new_[20534]_  = ~A201 & \new_[20533]_ ;
  assign \new_[20538]_  = A268 & A236;
  assign \new_[20539]_  = A233 & \new_[20538]_ ;
  assign \new_[20540]_  = \new_[20539]_  & \new_[20534]_ ;
  assign \new_[20543]_  = ~A167 & A170;
  assign \new_[20547]_  = A200 & A199;
  assign \new_[20548]_  = A166 & \new_[20547]_ ;
  assign \new_[20549]_  = \new_[20548]_  & \new_[20543]_ ;
  assign \new_[20553]_  = A232 & ~A202;
  assign \new_[20554]_  = ~A201 & \new_[20553]_ ;
  assign \new_[20558]_  = A268 & A236;
  assign \new_[20559]_  = ~A233 & \new_[20558]_ ;
  assign \new_[20560]_  = \new_[20559]_  & \new_[20554]_ ;
  assign \new_[20563]_  = ~A167 & A170;
  assign \new_[20567]_  = ~A200 & ~A199;
  assign \new_[20568]_  = A166 & \new_[20567]_ ;
  assign \new_[20569]_  = \new_[20568]_  & \new_[20563]_ ;
  assign \new_[20573]_  = A298 & A235;
  assign \new_[20574]_  = ~A202 & \new_[20573]_ ;
  assign \new_[20578]_  = ~A301 & ~A300;
  assign \new_[20579]_  = A299 & \new_[20578]_ ;
  assign \new_[20580]_  = \new_[20579]_  & \new_[20574]_ ;
  assign \new_[20583]_  = ~A167 & A170;
  assign \new_[20587]_  = ~A200 & ~A199;
  assign \new_[20588]_  = A166 & \new_[20587]_ ;
  assign \new_[20589]_  = \new_[20588]_  & \new_[20583]_ ;
  assign \new_[20593]_  = A234 & A232;
  assign \new_[20594]_  = ~A202 & \new_[20593]_ ;
  assign \new_[20598]_  = ~A302 & ~A301;
  assign \new_[20599]_  = ~A300 & \new_[20598]_ ;
  assign \new_[20600]_  = \new_[20599]_  & \new_[20594]_ ;
  assign \new_[20603]_  = ~A167 & A170;
  assign \new_[20607]_  = ~A200 & ~A199;
  assign \new_[20608]_  = A166 & \new_[20607]_ ;
  assign \new_[20609]_  = \new_[20608]_  & \new_[20603]_ ;
  assign \new_[20613]_  = A234 & A232;
  assign \new_[20614]_  = ~A202 & \new_[20613]_ ;
  assign \new_[20618]_  = ~A301 & ~A299;
  assign \new_[20619]_  = ~A298 & \new_[20618]_ ;
  assign \new_[20620]_  = \new_[20619]_  & \new_[20614]_ ;
  assign \new_[20623]_  = ~A167 & A170;
  assign \new_[20627]_  = ~A200 & ~A199;
  assign \new_[20628]_  = A166 & \new_[20627]_ ;
  assign \new_[20629]_  = \new_[20628]_  & \new_[20623]_ ;
  assign \new_[20633]_  = A234 & A232;
  assign \new_[20634]_  = ~A202 & \new_[20633]_ ;
  assign \new_[20638]_  = A269 & A266;
  assign \new_[20639]_  = ~A265 & \new_[20638]_ ;
  assign \new_[20640]_  = \new_[20639]_  & \new_[20634]_ ;
  assign \new_[20643]_  = ~A167 & A170;
  assign \new_[20647]_  = ~A200 & ~A199;
  assign \new_[20648]_  = A166 & \new_[20647]_ ;
  assign \new_[20649]_  = \new_[20648]_  & \new_[20643]_ ;
  assign \new_[20653]_  = A234 & A232;
  assign \new_[20654]_  = ~A202 & \new_[20653]_ ;
  assign \new_[20658]_  = A269 & ~A266;
  assign \new_[20659]_  = A265 & \new_[20658]_ ;
  assign \new_[20660]_  = \new_[20659]_  & \new_[20654]_ ;
  assign \new_[20663]_  = ~A167 & A170;
  assign \new_[20667]_  = ~A200 & ~A199;
  assign \new_[20668]_  = A166 & \new_[20667]_ ;
  assign \new_[20669]_  = \new_[20668]_  & \new_[20663]_ ;
  assign \new_[20673]_  = A234 & A233;
  assign \new_[20674]_  = ~A202 & \new_[20673]_ ;
  assign \new_[20678]_  = ~A302 & ~A301;
  assign \new_[20679]_  = ~A300 & \new_[20678]_ ;
  assign \new_[20680]_  = \new_[20679]_  & \new_[20674]_ ;
  assign \new_[20683]_  = ~A167 & A170;
  assign \new_[20687]_  = ~A200 & ~A199;
  assign \new_[20688]_  = A166 & \new_[20687]_ ;
  assign \new_[20689]_  = \new_[20688]_  & \new_[20683]_ ;
  assign \new_[20693]_  = A234 & A233;
  assign \new_[20694]_  = ~A202 & \new_[20693]_ ;
  assign \new_[20698]_  = ~A301 & ~A299;
  assign \new_[20699]_  = ~A298 & \new_[20698]_ ;
  assign \new_[20700]_  = \new_[20699]_  & \new_[20694]_ ;
  assign \new_[20703]_  = ~A167 & A170;
  assign \new_[20707]_  = ~A200 & ~A199;
  assign \new_[20708]_  = A166 & \new_[20707]_ ;
  assign \new_[20709]_  = \new_[20708]_  & \new_[20703]_ ;
  assign \new_[20713]_  = A234 & A233;
  assign \new_[20714]_  = ~A202 & \new_[20713]_ ;
  assign \new_[20718]_  = A269 & A266;
  assign \new_[20719]_  = ~A265 & \new_[20718]_ ;
  assign \new_[20720]_  = \new_[20719]_  & \new_[20714]_ ;
  assign \new_[20723]_  = ~A167 & A170;
  assign \new_[20727]_  = ~A200 & ~A199;
  assign \new_[20728]_  = A166 & \new_[20727]_ ;
  assign \new_[20729]_  = \new_[20728]_  & \new_[20723]_ ;
  assign \new_[20733]_  = A234 & A233;
  assign \new_[20734]_  = ~A202 & \new_[20733]_ ;
  assign \new_[20738]_  = A269 & ~A266;
  assign \new_[20739]_  = A265 & \new_[20738]_ ;
  assign \new_[20740]_  = \new_[20739]_  & \new_[20734]_ ;
  assign \new_[20743]_  = ~A167 & A170;
  assign \new_[20747]_  = ~A200 & ~A199;
  assign \new_[20748]_  = A166 & \new_[20747]_ ;
  assign \new_[20749]_  = \new_[20748]_  & \new_[20743]_ ;
  assign \new_[20753]_  = A233 & ~A232;
  assign \new_[20754]_  = ~A202 & \new_[20753]_ ;
  assign \new_[20758]_  = A267 & A265;
  assign \new_[20759]_  = A236 & \new_[20758]_ ;
  assign \new_[20760]_  = \new_[20759]_  & \new_[20754]_ ;
  assign \new_[20763]_  = ~A167 & A170;
  assign \new_[20767]_  = ~A200 & ~A199;
  assign \new_[20768]_  = A166 & \new_[20767]_ ;
  assign \new_[20769]_  = \new_[20768]_  & \new_[20763]_ ;
  assign \new_[20773]_  = A233 & ~A232;
  assign \new_[20774]_  = ~A202 & \new_[20773]_ ;
  assign \new_[20778]_  = A267 & A266;
  assign \new_[20779]_  = A236 & \new_[20778]_ ;
  assign \new_[20780]_  = \new_[20779]_  & \new_[20774]_ ;
  assign \new_[20783]_  = ~A167 & A170;
  assign \new_[20787]_  = ~A200 & ~A199;
  assign \new_[20788]_  = A166 & \new_[20787]_ ;
  assign \new_[20789]_  = \new_[20788]_  & \new_[20783]_ ;
  assign \new_[20793]_  = ~A233 & A232;
  assign \new_[20794]_  = ~A202 & \new_[20793]_ ;
  assign \new_[20798]_  = A267 & A265;
  assign \new_[20799]_  = A236 & \new_[20798]_ ;
  assign \new_[20800]_  = \new_[20799]_  & \new_[20794]_ ;
  assign \new_[20803]_  = ~A167 & A170;
  assign \new_[20807]_  = ~A200 & ~A199;
  assign \new_[20808]_  = A166 & \new_[20807]_ ;
  assign \new_[20809]_  = \new_[20808]_  & \new_[20803]_ ;
  assign \new_[20813]_  = ~A233 & A232;
  assign \new_[20814]_  = ~A202 & \new_[20813]_ ;
  assign \new_[20818]_  = A267 & A266;
  assign \new_[20819]_  = A236 & \new_[20818]_ ;
  assign \new_[20820]_  = \new_[20819]_  & \new_[20814]_ ;
  assign \new_[20823]_  = ~A201 & A169;
  assign \new_[20827]_  = ~A234 & ~A203;
  assign \new_[20828]_  = ~A202 & \new_[20827]_ ;
  assign \new_[20829]_  = \new_[20828]_  & \new_[20823]_ ;
  assign \new_[20833]_  = ~A267 & ~A236;
  assign \new_[20834]_  = ~A235 & \new_[20833]_ ;
  assign \new_[20838]_  = A301 & ~A269;
  assign \new_[20839]_  = ~A268 & \new_[20838]_ ;
  assign \new_[20840]_  = \new_[20839]_  & \new_[20834]_ ;
  assign \new_[20843]_  = ~A201 & A169;
  assign \new_[20847]_  = ~A234 & ~A203;
  assign \new_[20848]_  = ~A202 & \new_[20847]_ ;
  assign \new_[20849]_  = \new_[20848]_  & \new_[20843]_ ;
  assign \new_[20853]_  = ~A265 & ~A236;
  assign \new_[20854]_  = ~A235 & \new_[20853]_ ;
  assign \new_[20858]_  = A301 & ~A268;
  assign \new_[20859]_  = ~A266 & \new_[20858]_ ;
  assign \new_[20860]_  = \new_[20859]_  & \new_[20854]_ ;
  assign \new_[20863]_  = ~A201 & A169;
  assign \new_[20867]_  = ~A232 & ~A203;
  assign \new_[20868]_  = ~A202 & \new_[20867]_ ;
  assign \new_[20869]_  = \new_[20868]_  & \new_[20863]_ ;
  assign \new_[20873]_  = A298 & A236;
  assign \new_[20874]_  = A233 & \new_[20873]_ ;
  assign \new_[20878]_  = ~A301 & ~A300;
  assign \new_[20879]_  = A299 & \new_[20878]_ ;
  assign \new_[20880]_  = \new_[20879]_  & \new_[20874]_ ;
  assign \new_[20883]_  = ~A201 & A169;
  assign \new_[20887]_  = A232 & ~A203;
  assign \new_[20888]_  = ~A202 & \new_[20887]_ ;
  assign \new_[20889]_  = \new_[20888]_  & \new_[20883]_ ;
  assign \new_[20893]_  = A298 & A236;
  assign \new_[20894]_  = ~A233 & \new_[20893]_ ;
  assign \new_[20898]_  = ~A301 & ~A300;
  assign \new_[20899]_  = A299 & \new_[20898]_ ;
  assign \new_[20900]_  = \new_[20899]_  & \new_[20894]_ ;
  assign \new_[20903]_  = ~A201 & A169;
  assign \new_[20907]_  = ~A232 & ~A203;
  assign \new_[20908]_  = ~A202 & \new_[20907]_ ;
  assign \new_[20909]_  = \new_[20908]_  & \new_[20903]_ ;
  assign \new_[20913]_  = ~A267 & ~A235;
  assign \new_[20914]_  = ~A233 & \new_[20913]_ ;
  assign \new_[20918]_  = A301 & ~A269;
  assign \new_[20919]_  = ~A268 & \new_[20918]_ ;
  assign \new_[20920]_  = \new_[20919]_  & \new_[20914]_ ;
  assign \new_[20923]_  = ~A201 & A169;
  assign \new_[20927]_  = ~A232 & ~A203;
  assign \new_[20928]_  = ~A202 & \new_[20927]_ ;
  assign \new_[20929]_  = \new_[20928]_  & \new_[20923]_ ;
  assign \new_[20933]_  = ~A265 & ~A235;
  assign \new_[20934]_  = ~A233 & \new_[20933]_ ;
  assign \new_[20938]_  = A301 & ~A268;
  assign \new_[20939]_  = ~A266 & \new_[20938]_ ;
  assign \new_[20940]_  = \new_[20939]_  & \new_[20934]_ ;
  assign \new_[20943]_  = A199 & A169;
  assign \new_[20947]_  = ~A202 & ~A201;
  assign \new_[20948]_  = A200 & \new_[20947]_ ;
  assign \new_[20949]_  = \new_[20948]_  & \new_[20943]_ ;
  assign \new_[20953]_  = A298 & A234;
  assign \new_[20954]_  = A232 & \new_[20953]_ ;
  assign \new_[20958]_  = ~A301 & ~A300;
  assign \new_[20959]_  = A299 & \new_[20958]_ ;
  assign \new_[20960]_  = \new_[20959]_  & \new_[20954]_ ;
  assign \new_[20963]_  = A199 & A169;
  assign \new_[20967]_  = ~A202 & ~A201;
  assign \new_[20968]_  = A200 & \new_[20967]_ ;
  assign \new_[20969]_  = \new_[20968]_  & \new_[20963]_ ;
  assign \new_[20973]_  = A298 & A234;
  assign \new_[20974]_  = A233 & \new_[20973]_ ;
  assign \new_[20978]_  = ~A301 & ~A300;
  assign \new_[20979]_  = A299 & \new_[20978]_ ;
  assign \new_[20980]_  = \new_[20979]_  & \new_[20974]_ ;
  assign \new_[20983]_  = A199 & A169;
  assign \new_[20987]_  = ~A202 & ~A201;
  assign \new_[20988]_  = A200 & \new_[20987]_ ;
  assign \new_[20989]_  = \new_[20988]_  & \new_[20983]_ ;
  assign \new_[20993]_  = A236 & A233;
  assign \new_[20994]_  = ~A232 & \new_[20993]_ ;
  assign \new_[20998]_  = ~A302 & ~A301;
  assign \new_[20999]_  = ~A300 & \new_[20998]_ ;
  assign \new_[21000]_  = \new_[20999]_  & \new_[20994]_ ;
  assign \new_[21003]_  = A199 & A169;
  assign \new_[21007]_  = ~A202 & ~A201;
  assign \new_[21008]_  = A200 & \new_[21007]_ ;
  assign \new_[21009]_  = \new_[21008]_  & \new_[21003]_ ;
  assign \new_[21013]_  = A236 & A233;
  assign \new_[21014]_  = ~A232 & \new_[21013]_ ;
  assign \new_[21018]_  = ~A301 & ~A299;
  assign \new_[21019]_  = ~A298 & \new_[21018]_ ;
  assign \new_[21020]_  = \new_[21019]_  & \new_[21014]_ ;
  assign \new_[21023]_  = A199 & A169;
  assign \new_[21027]_  = ~A202 & ~A201;
  assign \new_[21028]_  = A200 & \new_[21027]_ ;
  assign \new_[21029]_  = \new_[21028]_  & \new_[21023]_ ;
  assign \new_[21033]_  = A236 & A233;
  assign \new_[21034]_  = ~A232 & \new_[21033]_ ;
  assign \new_[21038]_  = A269 & A266;
  assign \new_[21039]_  = ~A265 & \new_[21038]_ ;
  assign \new_[21040]_  = \new_[21039]_  & \new_[21034]_ ;
  assign \new_[21043]_  = A199 & A169;
  assign \new_[21047]_  = ~A202 & ~A201;
  assign \new_[21048]_  = A200 & \new_[21047]_ ;
  assign \new_[21049]_  = \new_[21048]_  & \new_[21043]_ ;
  assign \new_[21053]_  = A236 & A233;
  assign \new_[21054]_  = ~A232 & \new_[21053]_ ;
  assign \new_[21058]_  = A269 & ~A266;
  assign \new_[21059]_  = A265 & \new_[21058]_ ;
  assign \new_[21060]_  = \new_[21059]_  & \new_[21054]_ ;
  assign \new_[21063]_  = A199 & A169;
  assign \new_[21067]_  = ~A202 & ~A201;
  assign \new_[21068]_  = A200 & \new_[21067]_ ;
  assign \new_[21069]_  = \new_[21068]_  & \new_[21063]_ ;
  assign \new_[21073]_  = A236 & ~A233;
  assign \new_[21074]_  = A232 & \new_[21073]_ ;
  assign \new_[21078]_  = ~A302 & ~A301;
  assign \new_[21079]_  = ~A300 & \new_[21078]_ ;
  assign \new_[21080]_  = \new_[21079]_  & \new_[21074]_ ;
  assign \new_[21083]_  = A199 & A169;
  assign \new_[21087]_  = ~A202 & ~A201;
  assign \new_[21088]_  = A200 & \new_[21087]_ ;
  assign \new_[21089]_  = \new_[21088]_  & \new_[21083]_ ;
  assign \new_[21093]_  = A236 & ~A233;
  assign \new_[21094]_  = A232 & \new_[21093]_ ;
  assign \new_[21098]_  = ~A301 & ~A299;
  assign \new_[21099]_  = ~A298 & \new_[21098]_ ;
  assign \new_[21100]_  = \new_[21099]_  & \new_[21094]_ ;
  assign \new_[21103]_  = A199 & A169;
  assign \new_[21107]_  = ~A202 & ~A201;
  assign \new_[21108]_  = A200 & \new_[21107]_ ;
  assign \new_[21109]_  = \new_[21108]_  & \new_[21103]_ ;
  assign \new_[21113]_  = A236 & ~A233;
  assign \new_[21114]_  = A232 & \new_[21113]_ ;
  assign \new_[21118]_  = A269 & A266;
  assign \new_[21119]_  = ~A265 & \new_[21118]_ ;
  assign \new_[21120]_  = \new_[21119]_  & \new_[21114]_ ;
  assign \new_[21123]_  = A199 & A169;
  assign \new_[21127]_  = ~A202 & ~A201;
  assign \new_[21128]_  = A200 & \new_[21127]_ ;
  assign \new_[21129]_  = \new_[21128]_  & \new_[21123]_ ;
  assign \new_[21133]_  = A236 & ~A233;
  assign \new_[21134]_  = A232 & \new_[21133]_ ;
  assign \new_[21138]_  = A269 & ~A266;
  assign \new_[21139]_  = A265 & \new_[21138]_ ;
  assign \new_[21140]_  = \new_[21139]_  & \new_[21134]_ ;
  assign \new_[21143]_  = ~A199 & A169;
  assign \new_[21147]_  = ~A234 & ~A202;
  assign \new_[21148]_  = ~A200 & \new_[21147]_ ;
  assign \new_[21149]_  = \new_[21148]_  & \new_[21143]_ ;
  assign \new_[21153]_  = ~A267 & ~A236;
  assign \new_[21154]_  = ~A235 & \new_[21153]_ ;
  assign \new_[21158]_  = A301 & ~A269;
  assign \new_[21159]_  = ~A268 & \new_[21158]_ ;
  assign \new_[21160]_  = \new_[21159]_  & \new_[21154]_ ;
  assign \new_[21163]_  = ~A199 & A169;
  assign \new_[21167]_  = ~A234 & ~A202;
  assign \new_[21168]_  = ~A200 & \new_[21167]_ ;
  assign \new_[21169]_  = \new_[21168]_  & \new_[21163]_ ;
  assign \new_[21173]_  = ~A265 & ~A236;
  assign \new_[21174]_  = ~A235 & \new_[21173]_ ;
  assign \new_[21178]_  = A301 & ~A268;
  assign \new_[21179]_  = ~A266 & \new_[21178]_ ;
  assign \new_[21180]_  = \new_[21179]_  & \new_[21174]_ ;
  assign \new_[21183]_  = ~A199 & A169;
  assign \new_[21187]_  = ~A232 & ~A202;
  assign \new_[21188]_  = ~A200 & \new_[21187]_ ;
  assign \new_[21189]_  = \new_[21188]_  & \new_[21183]_ ;
  assign \new_[21193]_  = A298 & A236;
  assign \new_[21194]_  = A233 & \new_[21193]_ ;
  assign \new_[21198]_  = ~A301 & ~A300;
  assign \new_[21199]_  = A299 & \new_[21198]_ ;
  assign \new_[21200]_  = \new_[21199]_  & \new_[21194]_ ;
  assign \new_[21203]_  = ~A199 & A169;
  assign \new_[21207]_  = A232 & ~A202;
  assign \new_[21208]_  = ~A200 & \new_[21207]_ ;
  assign \new_[21209]_  = \new_[21208]_  & \new_[21203]_ ;
  assign \new_[21213]_  = A298 & A236;
  assign \new_[21214]_  = ~A233 & \new_[21213]_ ;
  assign \new_[21218]_  = ~A301 & ~A300;
  assign \new_[21219]_  = A299 & \new_[21218]_ ;
  assign \new_[21220]_  = \new_[21219]_  & \new_[21214]_ ;
  assign \new_[21223]_  = ~A199 & A169;
  assign \new_[21227]_  = ~A232 & ~A202;
  assign \new_[21228]_  = ~A200 & \new_[21227]_ ;
  assign \new_[21229]_  = \new_[21228]_  & \new_[21223]_ ;
  assign \new_[21233]_  = ~A267 & ~A235;
  assign \new_[21234]_  = ~A233 & \new_[21233]_ ;
  assign \new_[21238]_  = A301 & ~A269;
  assign \new_[21239]_  = ~A268 & \new_[21238]_ ;
  assign \new_[21240]_  = \new_[21239]_  & \new_[21234]_ ;
  assign \new_[21243]_  = ~A199 & A169;
  assign \new_[21247]_  = ~A232 & ~A202;
  assign \new_[21248]_  = ~A200 & \new_[21247]_ ;
  assign \new_[21249]_  = \new_[21248]_  & \new_[21243]_ ;
  assign \new_[21253]_  = ~A265 & ~A235;
  assign \new_[21254]_  = ~A233 & \new_[21253]_ ;
  assign \new_[21258]_  = A301 & ~A268;
  assign \new_[21259]_  = ~A266 & \new_[21258]_ ;
  assign \new_[21260]_  = \new_[21259]_  & \new_[21254]_ ;
  assign \new_[21263]_  = ~A167 & ~A169;
  assign \new_[21267]_  = ~A234 & A202;
  assign \new_[21268]_  = ~A166 & \new_[21267]_ ;
  assign \new_[21269]_  = \new_[21268]_  & \new_[21263]_ ;
  assign \new_[21273]_  = ~A267 & ~A236;
  assign \new_[21274]_  = ~A235 & \new_[21273]_ ;
  assign \new_[21278]_  = A301 & ~A269;
  assign \new_[21279]_  = ~A268 & \new_[21278]_ ;
  assign \new_[21280]_  = \new_[21279]_  & \new_[21274]_ ;
  assign \new_[21283]_  = ~A167 & ~A169;
  assign \new_[21287]_  = ~A234 & A202;
  assign \new_[21288]_  = ~A166 & \new_[21287]_ ;
  assign \new_[21289]_  = \new_[21288]_  & \new_[21283]_ ;
  assign \new_[21293]_  = ~A265 & ~A236;
  assign \new_[21294]_  = ~A235 & \new_[21293]_ ;
  assign \new_[21298]_  = A301 & ~A268;
  assign \new_[21299]_  = ~A266 & \new_[21298]_ ;
  assign \new_[21300]_  = \new_[21299]_  & \new_[21294]_ ;
  assign \new_[21303]_  = ~A167 & ~A169;
  assign \new_[21307]_  = ~A232 & A202;
  assign \new_[21308]_  = ~A166 & \new_[21307]_ ;
  assign \new_[21309]_  = \new_[21308]_  & \new_[21303]_ ;
  assign \new_[21313]_  = A298 & A236;
  assign \new_[21314]_  = A233 & \new_[21313]_ ;
  assign \new_[21318]_  = ~A301 & ~A300;
  assign \new_[21319]_  = A299 & \new_[21318]_ ;
  assign \new_[21320]_  = \new_[21319]_  & \new_[21314]_ ;
  assign \new_[21323]_  = ~A167 & ~A169;
  assign \new_[21327]_  = A232 & A202;
  assign \new_[21328]_  = ~A166 & \new_[21327]_ ;
  assign \new_[21329]_  = \new_[21328]_  & \new_[21323]_ ;
  assign \new_[21333]_  = A298 & A236;
  assign \new_[21334]_  = ~A233 & \new_[21333]_ ;
  assign \new_[21338]_  = ~A301 & ~A300;
  assign \new_[21339]_  = A299 & \new_[21338]_ ;
  assign \new_[21340]_  = \new_[21339]_  & \new_[21334]_ ;
  assign \new_[21343]_  = ~A167 & ~A169;
  assign \new_[21347]_  = ~A232 & A202;
  assign \new_[21348]_  = ~A166 & \new_[21347]_ ;
  assign \new_[21349]_  = \new_[21348]_  & \new_[21343]_ ;
  assign \new_[21353]_  = ~A267 & ~A235;
  assign \new_[21354]_  = ~A233 & \new_[21353]_ ;
  assign \new_[21358]_  = A301 & ~A269;
  assign \new_[21359]_  = ~A268 & \new_[21358]_ ;
  assign \new_[21360]_  = \new_[21359]_  & \new_[21354]_ ;
  assign \new_[21363]_  = ~A167 & ~A169;
  assign \new_[21367]_  = ~A232 & A202;
  assign \new_[21368]_  = ~A166 & \new_[21367]_ ;
  assign \new_[21369]_  = \new_[21368]_  & \new_[21363]_ ;
  assign \new_[21373]_  = ~A265 & ~A235;
  assign \new_[21374]_  = ~A233 & \new_[21373]_ ;
  assign \new_[21378]_  = A301 & ~A268;
  assign \new_[21379]_  = ~A266 & \new_[21378]_ ;
  assign \new_[21380]_  = \new_[21379]_  & \new_[21374]_ ;
  assign \new_[21383]_  = ~A167 & ~A169;
  assign \new_[21387]_  = A201 & A199;
  assign \new_[21388]_  = ~A166 & \new_[21387]_ ;
  assign \new_[21389]_  = \new_[21388]_  & \new_[21383]_ ;
  assign \new_[21393]_  = A298 & A234;
  assign \new_[21394]_  = A232 & \new_[21393]_ ;
  assign \new_[21398]_  = ~A301 & ~A300;
  assign \new_[21399]_  = A299 & \new_[21398]_ ;
  assign \new_[21400]_  = \new_[21399]_  & \new_[21394]_ ;
  assign \new_[21403]_  = ~A167 & ~A169;
  assign \new_[21407]_  = A201 & A199;
  assign \new_[21408]_  = ~A166 & \new_[21407]_ ;
  assign \new_[21409]_  = \new_[21408]_  & \new_[21403]_ ;
  assign \new_[21413]_  = A298 & A234;
  assign \new_[21414]_  = A233 & \new_[21413]_ ;
  assign \new_[21418]_  = ~A301 & ~A300;
  assign \new_[21419]_  = A299 & \new_[21418]_ ;
  assign \new_[21420]_  = \new_[21419]_  & \new_[21414]_ ;
  assign \new_[21423]_  = ~A167 & ~A169;
  assign \new_[21427]_  = A201 & A199;
  assign \new_[21428]_  = ~A166 & \new_[21427]_ ;
  assign \new_[21429]_  = \new_[21428]_  & \new_[21423]_ ;
  assign \new_[21433]_  = A236 & A233;
  assign \new_[21434]_  = ~A232 & \new_[21433]_ ;
  assign \new_[21438]_  = ~A302 & ~A301;
  assign \new_[21439]_  = ~A300 & \new_[21438]_ ;
  assign \new_[21440]_  = \new_[21439]_  & \new_[21434]_ ;
  assign \new_[21443]_  = ~A167 & ~A169;
  assign \new_[21447]_  = A201 & A199;
  assign \new_[21448]_  = ~A166 & \new_[21447]_ ;
  assign \new_[21449]_  = \new_[21448]_  & \new_[21443]_ ;
  assign \new_[21453]_  = A236 & A233;
  assign \new_[21454]_  = ~A232 & \new_[21453]_ ;
  assign \new_[21458]_  = ~A301 & ~A299;
  assign \new_[21459]_  = ~A298 & \new_[21458]_ ;
  assign \new_[21460]_  = \new_[21459]_  & \new_[21454]_ ;
  assign \new_[21463]_  = ~A167 & ~A169;
  assign \new_[21467]_  = A201 & A199;
  assign \new_[21468]_  = ~A166 & \new_[21467]_ ;
  assign \new_[21469]_  = \new_[21468]_  & \new_[21463]_ ;
  assign \new_[21473]_  = A236 & A233;
  assign \new_[21474]_  = ~A232 & \new_[21473]_ ;
  assign \new_[21478]_  = A269 & A266;
  assign \new_[21479]_  = ~A265 & \new_[21478]_ ;
  assign \new_[21480]_  = \new_[21479]_  & \new_[21474]_ ;
  assign \new_[21483]_  = ~A167 & ~A169;
  assign \new_[21487]_  = A201 & A199;
  assign \new_[21488]_  = ~A166 & \new_[21487]_ ;
  assign \new_[21489]_  = \new_[21488]_  & \new_[21483]_ ;
  assign \new_[21493]_  = A236 & A233;
  assign \new_[21494]_  = ~A232 & \new_[21493]_ ;
  assign \new_[21498]_  = A269 & ~A266;
  assign \new_[21499]_  = A265 & \new_[21498]_ ;
  assign \new_[21500]_  = \new_[21499]_  & \new_[21494]_ ;
  assign \new_[21503]_  = ~A167 & ~A169;
  assign \new_[21507]_  = A201 & A199;
  assign \new_[21508]_  = ~A166 & \new_[21507]_ ;
  assign \new_[21509]_  = \new_[21508]_  & \new_[21503]_ ;
  assign \new_[21513]_  = A236 & ~A233;
  assign \new_[21514]_  = A232 & \new_[21513]_ ;
  assign \new_[21518]_  = ~A302 & ~A301;
  assign \new_[21519]_  = ~A300 & \new_[21518]_ ;
  assign \new_[21520]_  = \new_[21519]_  & \new_[21514]_ ;
  assign \new_[21523]_  = ~A167 & ~A169;
  assign \new_[21527]_  = A201 & A199;
  assign \new_[21528]_  = ~A166 & \new_[21527]_ ;
  assign \new_[21529]_  = \new_[21528]_  & \new_[21523]_ ;
  assign \new_[21533]_  = A236 & ~A233;
  assign \new_[21534]_  = A232 & \new_[21533]_ ;
  assign \new_[21538]_  = ~A301 & ~A299;
  assign \new_[21539]_  = ~A298 & \new_[21538]_ ;
  assign \new_[21540]_  = \new_[21539]_  & \new_[21534]_ ;
  assign \new_[21543]_  = ~A167 & ~A169;
  assign \new_[21547]_  = A201 & A199;
  assign \new_[21548]_  = ~A166 & \new_[21547]_ ;
  assign \new_[21549]_  = \new_[21548]_  & \new_[21543]_ ;
  assign \new_[21553]_  = A236 & ~A233;
  assign \new_[21554]_  = A232 & \new_[21553]_ ;
  assign \new_[21558]_  = A269 & A266;
  assign \new_[21559]_  = ~A265 & \new_[21558]_ ;
  assign \new_[21560]_  = \new_[21559]_  & \new_[21554]_ ;
  assign \new_[21563]_  = ~A167 & ~A169;
  assign \new_[21567]_  = A201 & A199;
  assign \new_[21568]_  = ~A166 & \new_[21567]_ ;
  assign \new_[21569]_  = \new_[21568]_  & \new_[21563]_ ;
  assign \new_[21573]_  = A236 & ~A233;
  assign \new_[21574]_  = A232 & \new_[21573]_ ;
  assign \new_[21578]_  = A269 & ~A266;
  assign \new_[21579]_  = A265 & \new_[21578]_ ;
  assign \new_[21580]_  = \new_[21579]_  & \new_[21574]_ ;
  assign \new_[21583]_  = ~A167 & ~A169;
  assign \new_[21587]_  = A201 & A200;
  assign \new_[21588]_  = ~A166 & \new_[21587]_ ;
  assign \new_[21589]_  = \new_[21588]_  & \new_[21583]_ ;
  assign \new_[21593]_  = A298 & A234;
  assign \new_[21594]_  = A232 & \new_[21593]_ ;
  assign \new_[21598]_  = ~A301 & ~A300;
  assign \new_[21599]_  = A299 & \new_[21598]_ ;
  assign \new_[21600]_  = \new_[21599]_  & \new_[21594]_ ;
  assign \new_[21603]_  = ~A167 & ~A169;
  assign \new_[21607]_  = A201 & A200;
  assign \new_[21608]_  = ~A166 & \new_[21607]_ ;
  assign \new_[21609]_  = \new_[21608]_  & \new_[21603]_ ;
  assign \new_[21613]_  = A298 & A234;
  assign \new_[21614]_  = A233 & \new_[21613]_ ;
  assign \new_[21618]_  = ~A301 & ~A300;
  assign \new_[21619]_  = A299 & \new_[21618]_ ;
  assign \new_[21620]_  = \new_[21619]_  & \new_[21614]_ ;
  assign \new_[21623]_  = ~A167 & ~A169;
  assign \new_[21627]_  = A201 & A200;
  assign \new_[21628]_  = ~A166 & \new_[21627]_ ;
  assign \new_[21629]_  = \new_[21628]_  & \new_[21623]_ ;
  assign \new_[21633]_  = A236 & A233;
  assign \new_[21634]_  = ~A232 & \new_[21633]_ ;
  assign \new_[21638]_  = ~A302 & ~A301;
  assign \new_[21639]_  = ~A300 & \new_[21638]_ ;
  assign \new_[21640]_  = \new_[21639]_  & \new_[21634]_ ;
  assign \new_[21643]_  = ~A167 & ~A169;
  assign \new_[21647]_  = A201 & A200;
  assign \new_[21648]_  = ~A166 & \new_[21647]_ ;
  assign \new_[21649]_  = \new_[21648]_  & \new_[21643]_ ;
  assign \new_[21653]_  = A236 & A233;
  assign \new_[21654]_  = ~A232 & \new_[21653]_ ;
  assign \new_[21658]_  = ~A301 & ~A299;
  assign \new_[21659]_  = ~A298 & \new_[21658]_ ;
  assign \new_[21660]_  = \new_[21659]_  & \new_[21654]_ ;
  assign \new_[21663]_  = ~A167 & ~A169;
  assign \new_[21667]_  = A201 & A200;
  assign \new_[21668]_  = ~A166 & \new_[21667]_ ;
  assign \new_[21669]_  = \new_[21668]_  & \new_[21663]_ ;
  assign \new_[21673]_  = A236 & A233;
  assign \new_[21674]_  = ~A232 & \new_[21673]_ ;
  assign \new_[21678]_  = A269 & A266;
  assign \new_[21679]_  = ~A265 & \new_[21678]_ ;
  assign \new_[21680]_  = \new_[21679]_  & \new_[21674]_ ;
  assign \new_[21683]_  = ~A167 & ~A169;
  assign \new_[21687]_  = A201 & A200;
  assign \new_[21688]_  = ~A166 & \new_[21687]_ ;
  assign \new_[21689]_  = \new_[21688]_  & \new_[21683]_ ;
  assign \new_[21693]_  = A236 & A233;
  assign \new_[21694]_  = ~A232 & \new_[21693]_ ;
  assign \new_[21698]_  = A269 & ~A266;
  assign \new_[21699]_  = A265 & \new_[21698]_ ;
  assign \new_[21700]_  = \new_[21699]_  & \new_[21694]_ ;
  assign \new_[21703]_  = ~A167 & ~A169;
  assign \new_[21707]_  = A201 & A200;
  assign \new_[21708]_  = ~A166 & \new_[21707]_ ;
  assign \new_[21709]_  = \new_[21708]_  & \new_[21703]_ ;
  assign \new_[21713]_  = A236 & ~A233;
  assign \new_[21714]_  = A232 & \new_[21713]_ ;
  assign \new_[21718]_  = ~A302 & ~A301;
  assign \new_[21719]_  = ~A300 & \new_[21718]_ ;
  assign \new_[21720]_  = \new_[21719]_  & \new_[21714]_ ;
  assign \new_[21723]_  = ~A167 & ~A169;
  assign \new_[21727]_  = A201 & A200;
  assign \new_[21728]_  = ~A166 & \new_[21727]_ ;
  assign \new_[21729]_  = \new_[21728]_  & \new_[21723]_ ;
  assign \new_[21733]_  = A236 & ~A233;
  assign \new_[21734]_  = A232 & \new_[21733]_ ;
  assign \new_[21738]_  = ~A301 & ~A299;
  assign \new_[21739]_  = ~A298 & \new_[21738]_ ;
  assign \new_[21740]_  = \new_[21739]_  & \new_[21734]_ ;
  assign \new_[21743]_  = ~A167 & ~A169;
  assign \new_[21747]_  = A201 & A200;
  assign \new_[21748]_  = ~A166 & \new_[21747]_ ;
  assign \new_[21749]_  = \new_[21748]_  & \new_[21743]_ ;
  assign \new_[21753]_  = A236 & ~A233;
  assign \new_[21754]_  = A232 & \new_[21753]_ ;
  assign \new_[21758]_  = A269 & A266;
  assign \new_[21759]_  = ~A265 & \new_[21758]_ ;
  assign \new_[21760]_  = \new_[21759]_  & \new_[21754]_ ;
  assign \new_[21763]_  = ~A167 & ~A169;
  assign \new_[21767]_  = A201 & A200;
  assign \new_[21768]_  = ~A166 & \new_[21767]_ ;
  assign \new_[21769]_  = \new_[21768]_  & \new_[21763]_ ;
  assign \new_[21773]_  = A236 & ~A233;
  assign \new_[21774]_  = A232 & \new_[21773]_ ;
  assign \new_[21778]_  = A269 & ~A266;
  assign \new_[21779]_  = A265 & \new_[21778]_ ;
  assign \new_[21780]_  = \new_[21779]_  & \new_[21774]_ ;
  assign \new_[21783]_  = ~A167 & ~A169;
  assign \new_[21787]_  = A200 & ~A199;
  assign \new_[21788]_  = ~A166 & \new_[21787]_ ;
  assign \new_[21789]_  = \new_[21788]_  & \new_[21783]_ ;
  assign \new_[21793]_  = A298 & A235;
  assign \new_[21794]_  = A203 & \new_[21793]_ ;
  assign \new_[21798]_  = ~A301 & ~A300;
  assign \new_[21799]_  = A299 & \new_[21798]_ ;
  assign \new_[21800]_  = \new_[21799]_  & \new_[21794]_ ;
  assign \new_[21803]_  = ~A167 & ~A169;
  assign \new_[21807]_  = A200 & ~A199;
  assign \new_[21808]_  = ~A166 & \new_[21807]_ ;
  assign \new_[21809]_  = \new_[21808]_  & \new_[21803]_ ;
  assign \new_[21813]_  = A234 & A232;
  assign \new_[21814]_  = A203 & \new_[21813]_ ;
  assign \new_[21818]_  = ~A302 & ~A301;
  assign \new_[21819]_  = ~A300 & \new_[21818]_ ;
  assign \new_[21820]_  = \new_[21819]_  & \new_[21814]_ ;
  assign \new_[21823]_  = ~A167 & ~A169;
  assign \new_[21827]_  = A200 & ~A199;
  assign \new_[21828]_  = ~A166 & \new_[21827]_ ;
  assign \new_[21829]_  = \new_[21828]_  & \new_[21823]_ ;
  assign \new_[21833]_  = A234 & A232;
  assign \new_[21834]_  = A203 & \new_[21833]_ ;
  assign \new_[21838]_  = ~A301 & ~A299;
  assign \new_[21839]_  = ~A298 & \new_[21838]_ ;
  assign \new_[21840]_  = \new_[21839]_  & \new_[21834]_ ;
  assign \new_[21843]_  = ~A167 & ~A169;
  assign \new_[21847]_  = A200 & ~A199;
  assign \new_[21848]_  = ~A166 & \new_[21847]_ ;
  assign \new_[21849]_  = \new_[21848]_  & \new_[21843]_ ;
  assign \new_[21853]_  = A234 & A232;
  assign \new_[21854]_  = A203 & \new_[21853]_ ;
  assign \new_[21858]_  = A269 & A266;
  assign \new_[21859]_  = ~A265 & \new_[21858]_ ;
  assign \new_[21860]_  = \new_[21859]_  & \new_[21854]_ ;
  assign \new_[21863]_  = ~A167 & ~A169;
  assign \new_[21867]_  = A200 & ~A199;
  assign \new_[21868]_  = ~A166 & \new_[21867]_ ;
  assign \new_[21869]_  = \new_[21868]_  & \new_[21863]_ ;
  assign \new_[21873]_  = A234 & A232;
  assign \new_[21874]_  = A203 & \new_[21873]_ ;
  assign \new_[21878]_  = A269 & ~A266;
  assign \new_[21879]_  = A265 & \new_[21878]_ ;
  assign \new_[21880]_  = \new_[21879]_  & \new_[21874]_ ;
  assign \new_[21883]_  = ~A167 & ~A169;
  assign \new_[21887]_  = A200 & ~A199;
  assign \new_[21888]_  = ~A166 & \new_[21887]_ ;
  assign \new_[21889]_  = \new_[21888]_  & \new_[21883]_ ;
  assign \new_[21893]_  = A234 & A233;
  assign \new_[21894]_  = A203 & \new_[21893]_ ;
  assign \new_[21898]_  = ~A302 & ~A301;
  assign \new_[21899]_  = ~A300 & \new_[21898]_ ;
  assign \new_[21900]_  = \new_[21899]_  & \new_[21894]_ ;
  assign \new_[21903]_  = ~A167 & ~A169;
  assign \new_[21907]_  = A200 & ~A199;
  assign \new_[21908]_  = ~A166 & \new_[21907]_ ;
  assign \new_[21909]_  = \new_[21908]_  & \new_[21903]_ ;
  assign \new_[21913]_  = A234 & A233;
  assign \new_[21914]_  = A203 & \new_[21913]_ ;
  assign \new_[21918]_  = ~A301 & ~A299;
  assign \new_[21919]_  = ~A298 & \new_[21918]_ ;
  assign \new_[21920]_  = \new_[21919]_  & \new_[21914]_ ;
  assign \new_[21923]_  = ~A167 & ~A169;
  assign \new_[21927]_  = A200 & ~A199;
  assign \new_[21928]_  = ~A166 & \new_[21927]_ ;
  assign \new_[21929]_  = \new_[21928]_  & \new_[21923]_ ;
  assign \new_[21933]_  = A234 & A233;
  assign \new_[21934]_  = A203 & \new_[21933]_ ;
  assign \new_[21938]_  = A269 & A266;
  assign \new_[21939]_  = ~A265 & \new_[21938]_ ;
  assign \new_[21940]_  = \new_[21939]_  & \new_[21934]_ ;
  assign \new_[21943]_  = ~A167 & ~A169;
  assign \new_[21947]_  = A200 & ~A199;
  assign \new_[21948]_  = ~A166 & \new_[21947]_ ;
  assign \new_[21949]_  = \new_[21948]_  & \new_[21943]_ ;
  assign \new_[21953]_  = A234 & A233;
  assign \new_[21954]_  = A203 & \new_[21953]_ ;
  assign \new_[21958]_  = A269 & ~A266;
  assign \new_[21959]_  = A265 & \new_[21958]_ ;
  assign \new_[21960]_  = \new_[21959]_  & \new_[21954]_ ;
  assign \new_[21963]_  = ~A167 & ~A169;
  assign \new_[21967]_  = A200 & ~A199;
  assign \new_[21968]_  = ~A166 & \new_[21967]_ ;
  assign \new_[21969]_  = \new_[21968]_  & \new_[21963]_ ;
  assign \new_[21973]_  = A233 & ~A232;
  assign \new_[21974]_  = A203 & \new_[21973]_ ;
  assign \new_[21978]_  = A267 & A265;
  assign \new_[21979]_  = A236 & \new_[21978]_ ;
  assign \new_[21980]_  = \new_[21979]_  & \new_[21974]_ ;
  assign \new_[21983]_  = ~A167 & ~A169;
  assign \new_[21987]_  = A200 & ~A199;
  assign \new_[21988]_  = ~A166 & \new_[21987]_ ;
  assign \new_[21989]_  = \new_[21988]_  & \new_[21983]_ ;
  assign \new_[21993]_  = A233 & ~A232;
  assign \new_[21994]_  = A203 & \new_[21993]_ ;
  assign \new_[21998]_  = A267 & A266;
  assign \new_[21999]_  = A236 & \new_[21998]_ ;
  assign \new_[22000]_  = \new_[21999]_  & \new_[21994]_ ;
  assign \new_[22003]_  = ~A167 & ~A169;
  assign \new_[22007]_  = A200 & ~A199;
  assign \new_[22008]_  = ~A166 & \new_[22007]_ ;
  assign \new_[22009]_  = \new_[22008]_  & \new_[22003]_ ;
  assign \new_[22013]_  = ~A233 & A232;
  assign \new_[22014]_  = A203 & \new_[22013]_ ;
  assign \new_[22018]_  = A267 & A265;
  assign \new_[22019]_  = A236 & \new_[22018]_ ;
  assign \new_[22020]_  = \new_[22019]_  & \new_[22014]_ ;
  assign \new_[22023]_  = ~A167 & ~A169;
  assign \new_[22027]_  = A200 & ~A199;
  assign \new_[22028]_  = ~A166 & \new_[22027]_ ;
  assign \new_[22029]_  = \new_[22028]_  & \new_[22023]_ ;
  assign \new_[22033]_  = ~A233 & A232;
  assign \new_[22034]_  = A203 & \new_[22033]_ ;
  assign \new_[22038]_  = A267 & A266;
  assign \new_[22039]_  = A236 & \new_[22038]_ ;
  assign \new_[22040]_  = \new_[22039]_  & \new_[22034]_ ;
  assign \new_[22043]_  = ~A167 & ~A169;
  assign \new_[22047]_  = ~A200 & A199;
  assign \new_[22048]_  = ~A166 & \new_[22047]_ ;
  assign \new_[22049]_  = \new_[22048]_  & \new_[22043]_ ;
  assign \new_[22053]_  = A298 & A235;
  assign \new_[22054]_  = A203 & \new_[22053]_ ;
  assign \new_[22058]_  = ~A301 & ~A300;
  assign \new_[22059]_  = A299 & \new_[22058]_ ;
  assign \new_[22060]_  = \new_[22059]_  & \new_[22054]_ ;
  assign \new_[22063]_  = ~A167 & ~A169;
  assign \new_[22067]_  = ~A200 & A199;
  assign \new_[22068]_  = ~A166 & \new_[22067]_ ;
  assign \new_[22069]_  = \new_[22068]_  & \new_[22063]_ ;
  assign \new_[22073]_  = A234 & A232;
  assign \new_[22074]_  = A203 & \new_[22073]_ ;
  assign \new_[22078]_  = ~A302 & ~A301;
  assign \new_[22079]_  = ~A300 & \new_[22078]_ ;
  assign \new_[22080]_  = \new_[22079]_  & \new_[22074]_ ;
  assign \new_[22083]_  = ~A167 & ~A169;
  assign \new_[22087]_  = ~A200 & A199;
  assign \new_[22088]_  = ~A166 & \new_[22087]_ ;
  assign \new_[22089]_  = \new_[22088]_  & \new_[22083]_ ;
  assign \new_[22093]_  = A234 & A232;
  assign \new_[22094]_  = A203 & \new_[22093]_ ;
  assign \new_[22098]_  = ~A301 & ~A299;
  assign \new_[22099]_  = ~A298 & \new_[22098]_ ;
  assign \new_[22100]_  = \new_[22099]_  & \new_[22094]_ ;
  assign \new_[22103]_  = ~A167 & ~A169;
  assign \new_[22107]_  = ~A200 & A199;
  assign \new_[22108]_  = ~A166 & \new_[22107]_ ;
  assign \new_[22109]_  = \new_[22108]_  & \new_[22103]_ ;
  assign \new_[22113]_  = A234 & A232;
  assign \new_[22114]_  = A203 & \new_[22113]_ ;
  assign \new_[22118]_  = A269 & A266;
  assign \new_[22119]_  = ~A265 & \new_[22118]_ ;
  assign \new_[22120]_  = \new_[22119]_  & \new_[22114]_ ;
  assign \new_[22123]_  = ~A167 & ~A169;
  assign \new_[22127]_  = ~A200 & A199;
  assign \new_[22128]_  = ~A166 & \new_[22127]_ ;
  assign \new_[22129]_  = \new_[22128]_  & \new_[22123]_ ;
  assign \new_[22133]_  = A234 & A232;
  assign \new_[22134]_  = A203 & \new_[22133]_ ;
  assign \new_[22138]_  = A269 & ~A266;
  assign \new_[22139]_  = A265 & \new_[22138]_ ;
  assign \new_[22140]_  = \new_[22139]_  & \new_[22134]_ ;
  assign \new_[22143]_  = ~A167 & ~A169;
  assign \new_[22147]_  = ~A200 & A199;
  assign \new_[22148]_  = ~A166 & \new_[22147]_ ;
  assign \new_[22149]_  = \new_[22148]_  & \new_[22143]_ ;
  assign \new_[22153]_  = A234 & A233;
  assign \new_[22154]_  = A203 & \new_[22153]_ ;
  assign \new_[22158]_  = ~A302 & ~A301;
  assign \new_[22159]_  = ~A300 & \new_[22158]_ ;
  assign \new_[22160]_  = \new_[22159]_  & \new_[22154]_ ;
  assign \new_[22163]_  = ~A167 & ~A169;
  assign \new_[22167]_  = ~A200 & A199;
  assign \new_[22168]_  = ~A166 & \new_[22167]_ ;
  assign \new_[22169]_  = \new_[22168]_  & \new_[22163]_ ;
  assign \new_[22173]_  = A234 & A233;
  assign \new_[22174]_  = A203 & \new_[22173]_ ;
  assign \new_[22178]_  = ~A301 & ~A299;
  assign \new_[22179]_  = ~A298 & \new_[22178]_ ;
  assign \new_[22180]_  = \new_[22179]_  & \new_[22174]_ ;
  assign \new_[22183]_  = ~A167 & ~A169;
  assign \new_[22187]_  = ~A200 & A199;
  assign \new_[22188]_  = ~A166 & \new_[22187]_ ;
  assign \new_[22189]_  = \new_[22188]_  & \new_[22183]_ ;
  assign \new_[22193]_  = A234 & A233;
  assign \new_[22194]_  = A203 & \new_[22193]_ ;
  assign \new_[22198]_  = A269 & A266;
  assign \new_[22199]_  = ~A265 & \new_[22198]_ ;
  assign \new_[22200]_  = \new_[22199]_  & \new_[22194]_ ;
  assign \new_[22203]_  = ~A167 & ~A169;
  assign \new_[22207]_  = ~A200 & A199;
  assign \new_[22208]_  = ~A166 & \new_[22207]_ ;
  assign \new_[22209]_  = \new_[22208]_  & \new_[22203]_ ;
  assign \new_[22213]_  = A234 & A233;
  assign \new_[22214]_  = A203 & \new_[22213]_ ;
  assign \new_[22218]_  = A269 & ~A266;
  assign \new_[22219]_  = A265 & \new_[22218]_ ;
  assign \new_[22220]_  = \new_[22219]_  & \new_[22214]_ ;
  assign \new_[22223]_  = ~A167 & ~A169;
  assign \new_[22227]_  = ~A200 & A199;
  assign \new_[22228]_  = ~A166 & \new_[22227]_ ;
  assign \new_[22229]_  = \new_[22228]_  & \new_[22223]_ ;
  assign \new_[22233]_  = A233 & ~A232;
  assign \new_[22234]_  = A203 & \new_[22233]_ ;
  assign \new_[22238]_  = A267 & A265;
  assign \new_[22239]_  = A236 & \new_[22238]_ ;
  assign \new_[22240]_  = \new_[22239]_  & \new_[22234]_ ;
  assign \new_[22243]_  = ~A167 & ~A169;
  assign \new_[22247]_  = ~A200 & A199;
  assign \new_[22248]_  = ~A166 & \new_[22247]_ ;
  assign \new_[22249]_  = \new_[22248]_  & \new_[22243]_ ;
  assign \new_[22253]_  = A233 & ~A232;
  assign \new_[22254]_  = A203 & \new_[22253]_ ;
  assign \new_[22258]_  = A267 & A266;
  assign \new_[22259]_  = A236 & \new_[22258]_ ;
  assign \new_[22260]_  = \new_[22259]_  & \new_[22254]_ ;
  assign \new_[22263]_  = ~A167 & ~A169;
  assign \new_[22267]_  = ~A200 & A199;
  assign \new_[22268]_  = ~A166 & \new_[22267]_ ;
  assign \new_[22269]_  = \new_[22268]_  & \new_[22263]_ ;
  assign \new_[22273]_  = ~A233 & A232;
  assign \new_[22274]_  = A203 & \new_[22273]_ ;
  assign \new_[22278]_  = A267 & A265;
  assign \new_[22279]_  = A236 & \new_[22278]_ ;
  assign \new_[22280]_  = \new_[22279]_  & \new_[22274]_ ;
  assign \new_[22283]_  = ~A167 & ~A169;
  assign \new_[22287]_  = ~A200 & A199;
  assign \new_[22288]_  = ~A166 & \new_[22287]_ ;
  assign \new_[22289]_  = \new_[22288]_  & \new_[22283]_ ;
  assign \new_[22293]_  = ~A233 & A232;
  assign \new_[22294]_  = A203 & \new_[22293]_ ;
  assign \new_[22298]_  = A267 & A266;
  assign \new_[22299]_  = A236 & \new_[22298]_ ;
  assign \new_[22300]_  = \new_[22299]_  & \new_[22294]_ ;
  assign \new_[22303]_  = ~A168 & ~A169;
  assign \new_[22307]_  = A202 & A166;
  assign \new_[22308]_  = A167 & \new_[22307]_ ;
  assign \new_[22309]_  = \new_[22308]_  & \new_[22303]_ ;
  assign \new_[22313]_  = A298 & A234;
  assign \new_[22314]_  = A232 & \new_[22313]_ ;
  assign \new_[22318]_  = ~A301 & ~A300;
  assign \new_[22319]_  = A299 & \new_[22318]_ ;
  assign \new_[22320]_  = \new_[22319]_  & \new_[22314]_ ;
  assign \new_[22323]_  = ~A168 & ~A169;
  assign \new_[22327]_  = A202 & A166;
  assign \new_[22328]_  = A167 & \new_[22327]_ ;
  assign \new_[22329]_  = \new_[22328]_  & \new_[22323]_ ;
  assign \new_[22333]_  = A298 & A234;
  assign \new_[22334]_  = A233 & \new_[22333]_ ;
  assign \new_[22338]_  = ~A301 & ~A300;
  assign \new_[22339]_  = A299 & \new_[22338]_ ;
  assign \new_[22340]_  = \new_[22339]_  & \new_[22334]_ ;
  assign \new_[22343]_  = ~A168 & ~A169;
  assign \new_[22347]_  = A202 & A166;
  assign \new_[22348]_  = A167 & \new_[22347]_ ;
  assign \new_[22349]_  = \new_[22348]_  & \new_[22343]_ ;
  assign \new_[22353]_  = A236 & A233;
  assign \new_[22354]_  = ~A232 & \new_[22353]_ ;
  assign \new_[22358]_  = ~A302 & ~A301;
  assign \new_[22359]_  = ~A300 & \new_[22358]_ ;
  assign \new_[22360]_  = \new_[22359]_  & \new_[22354]_ ;
  assign \new_[22363]_  = ~A168 & ~A169;
  assign \new_[22367]_  = A202 & A166;
  assign \new_[22368]_  = A167 & \new_[22367]_ ;
  assign \new_[22369]_  = \new_[22368]_  & \new_[22363]_ ;
  assign \new_[22373]_  = A236 & A233;
  assign \new_[22374]_  = ~A232 & \new_[22373]_ ;
  assign \new_[22378]_  = ~A301 & ~A299;
  assign \new_[22379]_  = ~A298 & \new_[22378]_ ;
  assign \new_[22380]_  = \new_[22379]_  & \new_[22374]_ ;
  assign \new_[22383]_  = ~A168 & ~A169;
  assign \new_[22387]_  = A202 & A166;
  assign \new_[22388]_  = A167 & \new_[22387]_ ;
  assign \new_[22389]_  = \new_[22388]_  & \new_[22383]_ ;
  assign \new_[22393]_  = A236 & A233;
  assign \new_[22394]_  = ~A232 & \new_[22393]_ ;
  assign \new_[22398]_  = A269 & A266;
  assign \new_[22399]_  = ~A265 & \new_[22398]_ ;
  assign \new_[22400]_  = \new_[22399]_  & \new_[22394]_ ;
  assign \new_[22403]_  = ~A168 & ~A169;
  assign \new_[22407]_  = A202 & A166;
  assign \new_[22408]_  = A167 & \new_[22407]_ ;
  assign \new_[22409]_  = \new_[22408]_  & \new_[22403]_ ;
  assign \new_[22413]_  = A236 & A233;
  assign \new_[22414]_  = ~A232 & \new_[22413]_ ;
  assign \new_[22418]_  = A269 & ~A266;
  assign \new_[22419]_  = A265 & \new_[22418]_ ;
  assign \new_[22420]_  = \new_[22419]_  & \new_[22414]_ ;
  assign \new_[22423]_  = ~A168 & ~A169;
  assign \new_[22427]_  = A202 & A166;
  assign \new_[22428]_  = A167 & \new_[22427]_ ;
  assign \new_[22429]_  = \new_[22428]_  & \new_[22423]_ ;
  assign \new_[22433]_  = A236 & ~A233;
  assign \new_[22434]_  = A232 & \new_[22433]_ ;
  assign \new_[22438]_  = ~A302 & ~A301;
  assign \new_[22439]_  = ~A300 & \new_[22438]_ ;
  assign \new_[22440]_  = \new_[22439]_  & \new_[22434]_ ;
  assign \new_[22443]_  = ~A168 & ~A169;
  assign \new_[22447]_  = A202 & A166;
  assign \new_[22448]_  = A167 & \new_[22447]_ ;
  assign \new_[22449]_  = \new_[22448]_  & \new_[22443]_ ;
  assign \new_[22453]_  = A236 & ~A233;
  assign \new_[22454]_  = A232 & \new_[22453]_ ;
  assign \new_[22458]_  = ~A301 & ~A299;
  assign \new_[22459]_  = ~A298 & \new_[22458]_ ;
  assign \new_[22460]_  = \new_[22459]_  & \new_[22454]_ ;
  assign \new_[22463]_  = ~A168 & ~A169;
  assign \new_[22467]_  = A202 & A166;
  assign \new_[22468]_  = A167 & \new_[22467]_ ;
  assign \new_[22469]_  = \new_[22468]_  & \new_[22463]_ ;
  assign \new_[22473]_  = A236 & ~A233;
  assign \new_[22474]_  = A232 & \new_[22473]_ ;
  assign \new_[22478]_  = A269 & A266;
  assign \new_[22479]_  = ~A265 & \new_[22478]_ ;
  assign \new_[22480]_  = \new_[22479]_  & \new_[22474]_ ;
  assign \new_[22483]_  = ~A168 & ~A169;
  assign \new_[22487]_  = A202 & A166;
  assign \new_[22488]_  = A167 & \new_[22487]_ ;
  assign \new_[22489]_  = \new_[22488]_  & \new_[22483]_ ;
  assign \new_[22493]_  = A236 & ~A233;
  assign \new_[22494]_  = A232 & \new_[22493]_ ;
  assign \new_[22498]_  = A269 & ~A266;
  assign \new_[22499]_  = A265 & \new_[22498]_ ;
  assign \new_[22500]_  = \new_[22499]_  & \new_[22494]_ ;
  assign \new_[22503]_  = ~A168 & ~A169;
  assign \new_[22507]_  = A199 & A166;
  assign \new_[22508]_  = A167 & \new_[22507]_ ;
  assign \new_[22509]_  = \new_[22508]_  & \new_[22503]_ ;
  assign \new_[22513]_  = A298 & A235;
  assign \new_[22514]_  = A201 & \new_[22513]_ ;
  assign \new_[22518]_  = ~A301 & ~A300;
  assign \new_[22519]_  = A299 & \new_[22518]_ ;
  assign \new_[22520]_  = \new_[22519]_  & \new_[22514]_ ;
  assign \new_[22523]_  = ~A168 & ~A169;
  assign \new_[22527]_  = A199 & A166;
  assign \new_[22528]_  = A167 & \new_[22527]_ ;
  assign \new_[22529]_  = \new_[22528]_  & \new_[22523]_ ;
  assign \new_[22533]_  = A234 & A232;
  assign \new_[22534]_  = A201 & \new_[22533]_ ;
  assign \new_[22538]_  = ~A302 & ~A301;
  assign \new_[22539]_  = ~A300 & \new_[22538]_ ;
  assign \new_[22540]_  = \new_[22539]_  & \new_[22534]_ ;
  assign \new_[22543]_  = ~A168 & ~A169;
  assign \new_[22547]_  = A199 & A166;
  assign \new_[22548]_  = A167 & \new_[22547]_ ;
  assign \new_[22549]_  = \new_[22548]_  & \new_[22543]_ ;
  assign \new_[22553]_  = A234 & A232;
  assign \new_[22554]_  = A201 & \new_[22553]_ ;
  assign \new_[22558]_  = ~A301 & ~A299;
  assign \new_[22559]_  = ~A298 & \new_[22558]_ ;
  assign \new_[22560]_  = \new_[22559]_  & \new_[22554]_ ;
  assign \new_[22563]_  = ~A168 & ~A169;
  assign \new_[22567]_  = A199 & A166;
  assign \new_[22568]_  = A167 & \new_[22567]_ ;
  assign \new_[22569]_  = \new_[22568]_  & \new_[22563]_ ;
  assign \new_[22573]_  = A234 & A232;
  assign \new_[22574]_  = A201 & \new_[22573]_ ;
  assign \new_[22578]_  = A269 & A266;
  assign \new_[22579]_  = ~A265 & \new_[22578]_ ;
  assign \new_[22580]_  = \new_[22579]_  & \new_[22574]_ ;
  assign \new_[22583]_  = ~A168 & ~A169;
  assign \new_[22587]_  = A199 & A166;
  assign \new_[22588]_  = A167 & \new_[22587]_ ;
  assign \new_[22589]_  = \new_[22588]_  & \new_[22583]_ ;
  assign \new_[22593]_  = A234 & A232;
  assign \new_[22594]_  = A201 & \new_[22593]_ ;
  assign \new_[22598]_  = A269 & ~A266;
  assign \new_[22599]_  = A265 & \new_[22598]_ ;
  assign \new_[22600]_  = \new_[22599]_  & \new_[22594]_ ;
  assign \new_[22603]_  = ~A168 & ~A169;
  assign \new_[22607]_  = A199 & A166;
  assign \new_[22608]_  = A167 & \new_[22607]_ ;
  assign \new_[22609]_  = \new_[22608]_  & \new_[22603]_ ;
  assign \new_[22613]_  = A234 & A233;
  assign \new_[22614]_  = A201 & \new_[22613]_ ;
  assign \new_[22618]_  = ~A302 & ~A301;
  assign \new_[22619]_  = ~A300 & \new_[22618]_ ;
  assign \new_[22620]_  = \new_[22619]_  & \new_[22614]_ ;
  assign \new_[22623]_  = ~A168 & ~A169;
  assign \new_[22627]_  = A199 & A166;
  assign \new_[22628]_  = A167 & \new_[22627]_ ;
  assign \new_[22629]_  = \new_[22628]_  & \new_[22623]_ ;
  assign \new_[22633]_  = A234 & A233;
  assign \new_[22634]_  = A201 & \new_[22633]_ ;
  assign \new_[22638]_  = ~A301 & ~A299;
  assign \new_[22639]_  = ~A298 & \new_[22638]_ ;
  assign \new_[22640]_  = \new_[22639]_  & \new_[22634]_ ;
  assign \new_[22643]_  = ~A168 & ~A169;
  assign \new_[22647]_  = A199 & A166;
  assign \new_[22648]_  = A167 & \new_[22647]_ ;
  assign \new_[22649]_  = \new_[22648]_  & \new_[22643]_ ;
  assign \new_[22653]_  = A234 & A233;
  assign \new_[22654]_  = A201 & \new_[22653]_ ;
  assign \new_[22658]_  = A269 & A266;
  assign \new_[22659]_  = ~A265 & \new_[22658]_ ;
  assign \new_[22660]_  = \new_[22659]_  & \new_[22654]_ ;
  assign \new_[22663]_  = ~A168 & ~A169;
  assign \new_[22667]_  = A199 & A166;
  assign \new_[22668]_  = A167 & \new_[22667]_ ;
  assign \new_[22669]_  = \new_[22668]_  & \new_[22663]_ ;
  assign \new_[22673]_  = A234 & A233;
  assign \new_[22674]_  = A201 & \new_[22673]_ ;
  assign \new_[22678]_  = A269 & ~A266;
  assign \new_[22679]_  = A265 & \new_[22678]_ ;
  assign \new_[22680]_  = \new_[22679]_  & \new_[22674]_ ;
  assign \new_[22683]_  = ~A168 & ~A169;
  assign \new_[22687]_  = A199 & A166;
  assign \new_[22688]_  = A167 & \new_[22687]_ ;
  assign \new_[22689]_  = \new_[22688]_  & \new_[22683]_ ;
  assign \new_[22693]_  = A233 & ~A232;
  assign \new_[22694]_  = A201 & \new_[22693]_ ;
  assign \new_[22698]_  = A267 & A265;
  assign \new_[22699]_  = A236 & \new_[22698]_ ;
  assign \new_[22700]_  = \new_[22699]_  & \new_[22694]_ ;
  assign \new_[22703]_  = ~A168 & ~A169;
  assign \new_[22707]_  = A199 & A166;
  assign \new_[22708]_  = A167 & \new_[22707]_ ;
  assign \new_[22709]_  = \new_[22708]_  & \new_[22703]_ ;
  assign \new_[22713]_  = A233 & ~A232;
  assign \new_[22714]_  = A201 & \new_[22713]_ ;
  assign \new_[22718]_  = A267 & A266;
  assign \new_[22719]_  = A236 & \new_[22718]_ ;
  assign \new_[22720]_  = \new_[22719]_  & \new_[22714]_ ;
  assign \new_[22723]_  = ~A168 & ~A169;
  assign \new_[22727]_  = A199 & A166;
  assign \new_[22728]_  = A167 & \new_[22727]_ ;
  assign \new_[22729]_  = \new_[22728]_  & \new_[22723]_ ;
  assign \new_[22733]_  = ~A233 & A232;
  assign \new_[22734]_  = A201 & \new_[22733]_ ;
  assign \new_[22738]_  = A267 & A265;
  assign \new_[22739]_  = A236 & \new_[22738]_ ;
  assign \new_[22740]_  = \new_[22739]_  & \new_[22734]_ ;
  assign \new_[22743]_  = ~A168 & ~A169;
  assign \new_[22747]_  = A199 & A166;
  assign \new_[22748]_  = A167 & \new_[22747]_ ;
  assign \new_[22749]_  = \new_[22748]_  & \new_[22743]_ ;
  assign \new_[22753]_  = ~A233 & A232;
  assign \new_[22754]_  = A201 & \new_[22753]_ ;
  assign \new_[22758]_  = A267 & A266;
  assign \new_[22759]_  = A236 & \new_[22758]_ ;
  assign \new_[22760]_  = \new_[22759]_  & \new_[22754]_ ;
  assign \new_[22763]_  = ~A168 & ~A169;
  assign \new_[22767]_  = A200 & A166;
  assign \new_[22768]_  = A167 & \new_[22767]_ ;
  assign \new_[22769]_  = \new_[22768]_  & \new_[22763]_ ;
  assign \new_[22773]_  = A298 & A235;
  assign \new_[22774]_  = A201 & \new_[22773]_ ;
  assign \new_[22778]_  = ~A301 & ~A300;
  assign \new_[22779]_  = A299 & \new_[22778]_ ;
  assign \new_[22780]_  = \new_[22779]_  & \new_[22774]_ ;
  assign \new_[22783]_  = ~A168 & ~A169;
  assign \new_[22787]_  = A200 & A166;
  assign \new_[22788]_  = A167 & \new_[22787]_ ;
  assign \new_[22789]_  = \new_[22788]_  & \new_[22783]_ ;
  assign \new_[22793]_  = A234 & A232;
  assign \new_[22794]_  = A201 & \new_[22793]_ ;
  assign \new_[22798]_  = ~A302 & ~A301;
  assign \new_[22799]_  = ~A300 & \new_[22798]_ ;
  assign \new_[22800]_  = \new_[22799]_  & \new_[22794]_ ;
  assign \new_[22803]_  = ~A168 & ~A169;
  assign \new_[22807]_  = A200 & A166;
  assign \new_[22808]_  = A167 & \new_[22807]_ ;
  assign \new_[22809]_  = \new_[22808]_  & \new_[22803]_ ;
  assign \new_[22813]_  = A234 & A232;
  assign \new_[22814]_  = A201 & \new_[22813]_ ;
  assign \new_[22818]_  = ~A301 & ~A299;
  assign \new_[22819]_  = ~A298 & \new_[22818]_ ;
  assign \new_[22820]_  = \new_[22819]_  & \new_[22814]_ ;
  assign \new_[22823]_  = ~A168 & ~A169;
  assign \new_[22827]_  = A200 & A166;
  assign \new_[22828]_  = A167 & \new_[22827]_ ;
  assign \new_[22829]_  = \new_[22828]_  & \new_[22823]_ ;
  assign \new_[22833]_  = A234 & A232;
  assign \new_[22834]_  = A201 & \new_[22833]_ ;
  assign \new_[22838]_  = A269 & A266;
  assign \new_[22839]_  = ~A265 & \new_[22838]_ ;
  assign \new_[22840]_  = \new_[22839]_  & \new_[22834]_ ;
  assign \new_[22843]_  = ~A168 & ~A169;
  assign \new_[22847]_  = A200 & A166;
  assign \new_[22848]_  = A167 & \new_[22847]_ ;
  assign \new_[22849]_  = \new_[22848]_  & \new_[22843]_ ;
  assign \new_[22853]_  = A234 & A232;
  assign \new_[22854]_  = A201 & \new_[22853]_ ;
  assign \new_[22858]_  = A269 & ~A266;
  assign \new_[22859]_  = A265 & \new_[22858]_ ;
  assign \new_[22860]_  = \new_[22859]_  & \new_[22854]_ ;
  assign \new_[22863]_  = ~A168 & ~A169;
  assign \new_[22867]_  = A200 & A166;
  assign \new_[22868]_  = A167 & \new_[22867]_ ;
  assign \new_[22869]_  = \new_[22868]_  & \new_[22863]_ ;
  assign \new_[22873]_  = A234 & A233;
  assign \new_[22874]_  = A201 & \new_[22873]_ ;
  assign \new_[22878]_  = ~A302 & ~A301;
  assign \new_[22879]_  = ~A300 & \new_[22878]_ ;
  assign \new_[22880]_  = \new_[22879]_  & \new_[22874]_ ;
  assign \new_[22883]_  = ~A168 & ~A169;
  assign \new_[22887]_  = A200 & A166;
  assign \new_[22888]_  = A167 & \new_[22887]_ ;
  assign \new_[22889]_  = \new_[22888]_  & \new_[22883]_ ;
  assign \new_[22893]_  = A234 & A233;
  assign \new_[22894]_  = A201 & \new_[22893]_ ;
  assign \new_[22898]_  = ~A301 & ~A299;
  assign \new_[22899]_  = ~A298 & \new_[22898]_ ;
  assign \new_[22900]_  = \new_[22899]_  & \new_[22894]_ ;
  assign \new_[22903]_  = ~A168 & ~A169;
  assign \new_[22907]_  = A200 & A166;
  assign \new_[22908]_  = A167 & \new_[22907]_ ;
  assign \new_[22909]_  = \new_[22908]_  & \new_[22903]_ ;
  assign \new_[22913]_  = A234 & A233;
  assign \new_[22914]_  = A201 & \new_[22913]_ ;
  assign \new_[22918]_  = A269 & A266;
  assign \new_[22919]_  = ~A265 & \new_[22918]_ ;
  assign \new_[22920]_  = \new_[22919]_  & \new_[22914]_ ;
  assign \new_[22923]_  = ~A168 & ~A169;
  assign \new_[22927]_  = A200 & A166;
  assign \new_[22928]_  = A167 & \new_[22927]_ ;
  assign \new_[22929]_  = \new_[22928]_  & \new_[22923]_ ;
  assign \new_[22933]_  = A234 & A233;
  assign \new_[22934]_  = A201 & \new_[22933]_ ;
  assign \new_[22938]_  = A269 & ~A266;
  assign \new_[22939]_  = A265 & \new_[22938]_ ;
  assign \new_[22940]_  = \new_[22939]_  & \new_[22934]_ ;
  assign \new_[22943]_  = ~A168 & ~A169;
  assign \new_[22947]_  = A200 & A166;
  assign \new_[22948]_  = A167 & \new_[22947]_ ;
  assign \new_[22949]_  = \new_[22948]_  & \new_[22943]_ ;
  assign \new_[22953]_  = A233 & ~A232;
  assign \new_[22954]_  = A201 & \new_[22953]_ ;
  assign \new_[22958]_  = A267 & A265;
  assign \new_[22959]_  = A236 & \new_[22958]_ ;
  assign \new_[22960]_  = \new_[22959]_  & \new_[22954]_ ;
  assign \new_[22963]_  = ~A168 & ~A169;
  assign \new_[22967]_  = A200 & A166;
  assign \new_[22968]_  = A167 & \new_[22967]_ ;
  assign \new_[22969]_  = \new_[22968]_  & \new_[22963]_ ;
  assign \new_[22973]_  = A233 & ~A232;
  assign \new_[22974]_  = A201 & \new_[22973]_ ;
  assign \new_[22978]_  = A267 & A266;
  assign \new_[22979]_  = A236 & \new_[22978]_ ;
  assign \new_[22980]_  = \new_[22979]_  & \new_[22974]_ ;
  assign \new_[22983]_  = ~A168 & ~A169;
  assign \new_[22987]_  = A200 & A166;
  assign \new_[22988]_  = A167 & \new_[22987]_ ;
  assign \new_[22989]_  = \new_[22988]_  & \new_[22983]_ ;
  assign \new_[22993]_  = ~A233 & A232;
  assign \new_[22994]_  = A201 & \new_[22993]_ ;
  assign \new_[22998]_  = A267 & A265;
  assign \new_[22999]_  = A236 & \new_[22998]_ ;
  assign \new_[23000]_  = \new_[22999]_  & \new_[22994]_ ;
  assign \new_[23003]_  = ~A168 & ~A169;
  assign \new_[23007]_  = A200 & A166;
  assign \new_[23008]_  = A167 & \new_[23007]_ ;
  assign \new_[23009]_  = \new_[23008]_  & \new_[23003]_ ;
  assign \new_[23013]_  = ~A233 & A232;
  assign \new_[23014]_  = A201 & \new_[23013]_ ;
  assign \new_[23018]_  = A267 & A266;
  assign \new_[23019]_  = A236 & \new_[23018]_ ;
  assign \new_[23020]_  = \new_[23019]_  & \new_[23014]_ ;
  assign \new_[23023]_  = ~A168 & ~A169;
  assign \new_[23027]_  = ~A199 & A166;
  assign \new_[23028]_  = A167 & \new_[23027]_ ;
  assign \new_[23029]_  = \new_[23028]_  & \new_[23023]_ ;
  assign \new_[23033]_  = A235 & A203;
  assign \new_[23034]_  = A200 & \new_[23033]_ ;
  assign \new_[23038]_  = ~A302 & ~A301;
  assign \new_[23039]_  = ~A300 & \new_[23038]_ ;
  assign \new_[23040]_  = \new_[23039]_  & \new_[23034]_ ;
  assign \new_[23043]_  = ~A168 & ~A169;
  assign \new_[23047]_  = ~A199 & A166;
  assign \new_[23048]_  = A167 & \new_[23047]_ ;
  assign \new_[23049]_  = \new_[23048]_  & \new_[23043]_ ;
  assign \new_[23053]_  = A235 & A203;
  assign \new_[23054]_  = A200 & \new_[23053]_ ;
  assign \new_[23058]_  = ~A301 & ~A299;
  assign \new_[23059]_  = ~A298 & \new_[23058]_ ;
  assign \new_[23060]_  = \new_[23059]_  & \new_[23054]_ ;
  assign \new_[23063]_  = ~A168 & ~A169;
  assign \new_[23067]_  = ~A199 & A166;
  assign \new_[23068]_  = A167 & \new_[23067]_ ;
  assign \new_[23069]_  = \new_[23068]_  & \new_[23063]_ ;
  assign \new_[23073]_  = A235 & A203;
  assign \new_[23074]_  = A200 & \new_[23073]_ ;
  assign \new_[23078]_  = A269 & A266;
  assign \new_[23079]_  = ~A265 & \new_[23078]_ ;
  assign \new_[23080]_  = \new_[23079]_  & \new_[23074]_ ;
  assign \new_[23083]_  = ~A168 & ~A169;
  assign \new_[23087]_  = ~A199 & A166;
  assign \new_[23088]_  = A167 & \new_[23087]_ ;
  assign \new_[23089]_  = \new_[23088]_  & \new_[23083]_ ;
  assign \new_[23093]_  = A235 & A203;
  assign \new_[23094]_  = A200 & \new_[23093]_ ;
  assign \new_[23098]_  = A269 & ~A266;
  assign \new_[23099]_  = A265 & \new_[23098]_ ;
  assign \new_[23100]_  = \new_[23099]_  & \new_[23094]_ ;
  assign \new_[23103]_  = ~A168 & ~A169;
  assign \new_[23107]_  = ~A199 & A166;
  assign \new_[23108]_  = A167 & \new_[23107]_ ;
  assign \new_[23109]_  = \new_[23108]_  & \new_[23103]_ ;
  assign \new_[23113]_  = A232 & A203;
  assign \new_[23114]_  = A200 & \new_[23113]_ ;
  assign \new_[23118]_  = A267 & A265;
  assign \new_[23119]_  = A234 & \new_[23118]_ ;
  assign \new_[23120]_  = \new_[23119]_  & \new_[23114]_ ;
  assign \new_[23123]_  = ~A168 & ~A169;
  assign \new_[23127]_  = ~A199 & A166;
  assign \new_[23128]_  = A167 & \new_[23127]_ ;
  assign \new_[23129]_  = \new_[23128]_  & \new_[23123]_ ;
  assign \new_[23133]_  = A232 & A203;
  assign \new_[23134]_  = A200 & \new_[23133]_ ;
  assign \new_[23138]_  = A267 & A266;
  assign \new_[23139]_  = A234 & \new_[23138]_ ;
  assign \new_[23140]_  = \new_[23139]_  & \new_[23134]_ ;
  assign \new_[23143]_  = ~A168 & ~A169;
  assign \new_[23147]_  = ~A199 & A166;
  assign \new_[23148]_  = A167 & \new_[23147]_ ;
  assign \new_[23149]_  = \new_[23148]_  & \new_[23143]_ ;
  assign \new_[23153]_  = A233 & A203;
  assign \new_[23154]_  = A200 & \new_[23153]_ ;
  assign \new_[23158]_  = A267 & A265;
  assign \new_[23159]_  = A234 & \new_[23158]_ ;
  assign \new_[23160]_  = \new_[23159]_  & \new_[23154]_ ;
  assign \new_[23163]_  = ~A168 & ~A169;
  assign \new_[23167]_  = ~A199 & A166;
  assign \new_[23168]_  = A167 & \new_[23167]_ ;
  assign \new_[23169]_  = \new_[23168]_  & \new_[23163]_ ;
  assign \new_[23173]_  = A233 & A203;
  assign \new_[23174]_  = A200 & \new_[23173]_ ;
  assign \new_[23178]_  = A267 & A266;
  assign \new_[23179]_  = A234 & \new_[23178]_ ;
  assign \new_[23180]_  = \new_[23179]_  & \new_[23174]_ ;
  assign \new_[23183]_  = ~A168 & ~A169;
  assign \new_[23187]_  = ~A199 & A166;
  assign \new_[23188]_  = A167 & \new_[23187]_ ;
  assign \new_[23189]_  = \new_[23188]_  & \new_[23183]_ ;
  assign \new_[23193]_  = ~A232 & A203;
  assign \new_[23194]_  = A200 & \new_[23193]_ ;
  assign \new_[23198]_  = A268 & A236;
  assign \new_[23199]_  = A233 & \new_[23198]_ ;
  assign \new_[23200]_  = \new_[23199]_  & \new_[23194]_ ;
  assign \new_[23203]_  = ~A168 & ~A169;
  assign \new_[23207]_  = ~A199 & A166;
  assign \new_[23208]_  = A167 & \new_[23207]_ ;
  assign \new_[23209]_  = \new_[23208]_  & \new_[23203]_ ;
  assign \new_[23213]_  = A232 & A203;
  assign \new_[23214]_  = A200 & \new_[23213]_ ;
  assign \new_[23218]_  = A268 & A236;
  assign \new_[23219]_  = ~A233 & \new_[23218]_ ;
  assign \new_[23220]_  = \new_[23219]_  & \new_[23214]_ ;
  assign \new_[23223]_  = ~A168 & ~A169;
  assign \new_[23227]_  = A199 & A166;
  assign \new_[23228]_  = A167 & \new_[23227]_ ;
  assign \new_[23229]_  = \new_[23228]_  & \new_[23223]_ ;
  assign \new_[23233]_  = A235 & A203;
  assign \new_[23234]_  = ~A200 & \new_[23233]_ ;
  assign \new_[23238]_  = ~A302 & ~A301;
  assign \new_[23239]_  = ~A300 & \new_[23238]_ ;
  assign \new_[23240]_  = \new_[23239]_  & \new_[23234]_ ;
  assign \new_[23243]_  = ~A168 & ~A169;
  assign \new_[23247]_  = A199 & A166;
  assign \new_[23248]_  = A167 & \new_[23247]_ ;
  assign \new_[23249]_  = \new_[23248]_  & \new_[23243]_ ;
  assign \new_[23253]_  = A235 & A203;
  assign \new_[23254]_  = ~A200 & \new_[23253]_ ;
  assign \new_[23258]_  = ~A301 & ~A299;
  assign \new_[23259]_  = ~A298 & \new_[23258]_ ;
  assign \new_[23260]_  = \new_[23259]_  & \new_[23254]_ ;
  assign \new_[23263]_  = ~A168 & ~A169;
  assign \new_[23267]_  = A199 & A166;
  assign \new_[23268]_  = A167 & \new_[23267]_ ;
  assign \new_[23269]_  = \new_[23268]_  & \new_[23263]_ ;
  assign \new_[23273]_  = A235 & A203;
  assign \new_[23274]_  = ~A200 & \new_[23273]_ ;
  assign \new_[23278]_  = A269 & A266;
  assign \new_[23279]_  = ~A265 & \new_[23278]_ ;
  assign \new_[23280]_  = \new_[23279]_  & \new_[23274]_ ;
  assign \new_[23283]_  = ~A168 & ~A169;
  assign \new_[23287]_  = A199 & A166;
  assign \new_[23288]_  = A167 & \new_[23287]_ ;
  assign \new_[23289]_  = \new_[23288]_  & \new_[23283]_ ;
  assign \new_[23293]_  = A235 & A203;
  assign \new_[23294]_  = ~A200 & \new_[23293]_ ;
  assign \new_[23298]_  = A269 & ~A266;
  assign \new_[23299]_  = A265 & \new_[23298]_ ;
  assign \new_[23300]_  = \new_[23299]_  & \new_[23294]_ ;
  assign \new_[23303]_  = ~A168 & ~A169;
  assign \new_[23307]_  = A199 & A166;
  assign \new_[23308]_  = A167 & \new_[23307]_ ;
  assign \new_[23309]_  = \new_[23308]_  & \new_[23303]_ ;
  assign \new_[23313]_  = A232 & A203;
  assign \new_[23314]_  = ~A200 & \new_[23313]_ ;
  assign \new_[23318]_  = A267 & A265;
  assign \new_[23319]_  = A234 & \new_[23318]_ ;
  assign \new_[23320]_  = \new_[23319]_  & \new_[23314]_ ;
  assign \new_[23323]_  = ~A168 & ~A169;
  assign \new_[23327]_  = A199 & A166;
  assign \new_[23328]_  = A167 & \new_[23327]_ ;
  assign \new_[23329]_  = \new_[23328]_  & \new_[23323]_ ;
  assign \new_[23333]_  = A232 & A203;
  assign \new_[23334]_  = ~A200 & \new_[23333]_ ;
  assign \new_[23338]_  = A267 & A266;
  assign \new_[23339]_  = A234 & \new_[23338]_ ;
  assign \new_[23340]_  = \new_[23339]_  & \new_[23334]_ ;
  assign \new_[23343]_  = ~A168 & ~A169;
  assign \new_[23347]_  = A199 & A166;
  assign \new_[23348]_  = A167 & \new_[23347]_ ;
  assign \new_[23349]_  = \new_[23348]_  & \new_[23343]_ ;
  assign \new_[23353]_  = A233 & A203;
  assign \new_[23354]_  = ~A200 & \new_[23353]_ ;
  assign \new_[23358]_  = A267 & A265;
  assign \new_[23359]_  = A234 & \new_[23358]_ ;
  assign \new_[23360]_  = \new_[23359]_  & \new_[23354]_ ;
  assign \new_[23363]_  = ~A168 & ~A169;
  assign \new_[23367]_  = A199 & A166;
  assign \new_[23368]_  = A167 & \new_[23367]_ ;
  assign \new_[23369]_  = \new_[23368]_  & \new_[23363]_ ;
  assign \new_[23373]_  = A233 & A203;
  assign \new_[23374]_  = ~A200 & \new_[23373]_ ;
  assign \new_[23378]_  = A267 & A266;
  assign \new_[23379]_  = A234 & \new_[23378]_ ;
  assign \new_[23380]_  = \new_[23379]_  & \new_[23374]_ ;
  assign \new_[23383]_  = ~A168 & ~A169;
  assign \new_[23387]_  = A199 & A166;
  assign \new_[23388]_  = A167 & \new_[23387]_ ;
  assign \new_[23389]_  = \new_[23388]_  & \new_[23383]_ ;
  assign \new_[23393]_  = ~A232 & A203;
  assign \new_[23394]_  = ~A200 & \new_[23393]_ ;
  assign \new_[23398]_  = A268 & A236;
  assign \new_[23399]_  = A233 & \new_[23398]_ ;
  assign \new_[23400]_  = \new_[23399]_  & \new_[23394]_ ;
  assign \new_[23403]_  = ~A168 & ~A169;
  assign \new_[23407]_  = A199 & A166;
  assign \new_[23408]_  = A167 & \new_[23407]_ ;
  assign \new_[23409]_  = \new_[23408]_  & \new_[23403]_ ;
  assign \new_[23413]_  = A232 & A203;
  assign \new_[23414]_  = ~A200 & \new_[23413]_ ;
  assign \new_[23418]_  = A268 & A236;
  assign \new_[23419]_  = ~A233 & \new_[23418]_ ;
  assign \new_[23420]_  = \new_[23419]_  & \new_[23414]_ ;
  assign \new_[23423]_  = ~A169 & ~A170;
  assign \new_[23427]_  = ~A234 & A202;
  assign \new_[23428]_  = ~A168 & \new_[23427]_ ;
  assign \new_[23429]_  = \new_[23428]_  & \new_[23423]_ ;
  assign \new_[23433]_  = ~A267 & ~A236;
  assign \new_[23434]_  = ~A235 & \new_[23433]_ ;
  assign \new_[23438]_  = A301 & ~A269;
  assign \new_[23439]_  = ~A268 & \new_[23438]_ ;
  assign \new_[23440]_  = \new_[23439]_  & \new_[23434]_ ;
  assign \new_[23443]_  = ~A169 & ~A170;
  assign \new_[23447]_  = ~A234 & A202;
  assign \new_[23448]_  = ~A168 & \new_[23447]_ ;
  assign \new_[23449]_  = \new_[23448]_  & \new_[23443]_ ;
  assign \new_[23453]_  = ~A265 & ~A236;
  assign \new_[23454]_  = ~A235 & \new_[23453]_ ;
  assign \new_[23458]_  = A301 & ~A268;
  assign \new_[23459]_  = ~A266 & \new_[23458]_ ;
  assign \new_[23460]_  = \new_[23459]_  & \new_[23454]_ ;
  assign \new_[23463]_  = ~A169 & ~A170;
  assign \new_[23467]_  = ~A232 & A202;
  assign \new_[23468]_  = ~A168 & \new_[23467]_ ;
  assign \new_[23469]_  = \new_[23468]_  & \new_[23463]_ ;
  assign \new_[23473]_  = A298 & A236;
  assign \new_[23474]_  = A233 & \new_[23473]_ ;
  assign \new_[23478]_  = ~A301 & ~A300;
  assign \new_[23479]_  = A299 & \new_[23478]_ ;
  assign \new_[23480]_  = \new_[23479]_  & \new_[23474]_ ;
  assign \new_[23483]_  = ~A169 & ~A170;
  assign \new_[23487]_  = A232 & A202;
  assign \new_[23488]_  = ~A168 & \new_[23487]_ ;
  assign \new_[23489]_  = \new_[23488]_  & \new_[23483]_ ;
  assign \new_[23493]_  = A298 & A236;
  assign \new_[23494]_  = ~A233 & \new_[23493]_ ;
  assign \new_[23498]_  = ~A301 & ~A300;
  assign \new_[23499]_  = A299 & \new_[23498]_ ;
  assign \new_[23500]_  = \new_[23499]_  & \new_[23494]_ ;
  assign \new_[23503]_  = ~A169 & ~A170;
  assign \new_[23507]_  = ~A232 & A202;
  assign \new_[23508]_  = ~A168 & \new_[23507]_ ;
  assign \new_[23509]_  = \new_[23508]_  & \new_[23503]_ ;
  assign \new_[23513]_  = ~A267 & ~A235;
  assign \new_[23514]_  = ~A233 & \new_[23513]_ ;
  assign \new_[23518]_  = A301 & ~A269;
  assign \new_[23519]_  = ~A268 & \new_[23518]_ ;
  assign \new_[23520]_  = \new_[23519]_  & \new_[23514]_ ;
  assign \new_[23523]_  = ~A169 & ~A170;
  assign \new_[23527]_  = ~A232 & A202;
  assign \new_[23528]_  = ~A168 & \new_[23527]_ ;
  assign \new_[23529]_  = \new_[23528]_  & \new_[23523]_ ;
  assign \new_[23533]_  = ~A265 & ~A235;
  assign \new_[23534]_  = ~A233 & \new_[23533]_ ;
  assign \new_[23538]_  = A301 & ~A268;
  assign \new_[23539]_  = ~A266 & \new_[23538]_ ;
  assign \new_[23540]_  = \new_[23539]_  & \new_[23534]_ ;
  assign \new_[23543]_  = ~A169 & ~A170;
  assign \new_[23547]_  = A201 & A199;
  assign \new_[23548]_  = ~A168 & \new_[23547]_ ;
  assign \new_[23549]_  = \new_[23548]_  & \new_[23543]_ ;
  assign \new_[23553]_  = A298 & A234;
  assign \new_[23554]_  = A232 & \new_[23553]_ ;
  assign \new_[23558]_  = ~A301 & ~A300;
  assign \new_[23559]_  = A299 & \new_[23558]_ ;
  assign \new_[23560]_  = \new_[23559]_  & \new_[23554]_ ;
  assign \new_[23563]_  = ~A169 & ~A170;
  assign \new_[23567]_  = A201 & A199;
  assign \new_[23568]_  = ~A168 & \new_[23567]_ ;
  assign \new_[23569]_  = \new_[23568]_  & \new_[23563]_ ;
  assign \new_[23573]_  = A298 & A234;
  assign \new_[23574]_  = A233 & \new_[23573]_ ;
  assign \new_[23578]_  = ~A301 & ~A300;
  assign \new_[23579]_  = A299 & \new_[23578]_ ;
  assign \new_[23580]_  = \new_[23579]_  & \new_[23574]_ ;
  assign \new_[23583]_  = ~A169 & ~A170;
  assign \new_[23587]_  = A201 & A199;
  assign \new_[23588]_  = ~A168 & \new_[23587]_ ;
  assign \new_[23589]_  = \new_[23588]_  & \new_[23583]_ ;
  assign \new_[23593]_  = A236 & A233;
  assign \new_[23594]_  = ~A232 & \new_[23593]_ ;
  assign \new_[23598]_  = ~A302 & ~A301;
  assign \new_[23599]_  = ~A300 & \new_[23598]_ ;
  assign \new_[23600]_  = \new_[23599]_  & \new_[23594]_ ;
  assign \new_[23603]_  = ~A169 & ~A170;
  assign \new_[23607]_  = A201 & A199;
  assign \new_[23608]_  = ~A168 & \new_[23607]_ ;
  assign \new_[23609]_  = \new_[23608]_  & \new_[23603]_ ;
  assign \new_[23613]_  = A236 & A233;
  assign \new_[23614]_  = ~A232 & \new_[23613]_ ;
  assign \new_[23618]_  = ~A301 & ~A299;
  assign \new_[23619]_  = ~A298 & \new_[23618]_ ;
  assign \new_[23620]_  = \new_[23619]_  & \new_[23614]_ ;
  assign \new_[23623]_  = ~A169 & ~A170;
  assign \new_[23627]_  = A201 & A199;
  assign \new_[23628]_  = ~A168 & \new_[23627]_ ;
  assign \new_[23629]_  = \new_[23628]_  & \new_[23623]_ ;
  assign \new_[23633]_  = A236 & A233;
  assign \new_[23634]_  = ~A232 & \new_[23633]_ ;
  assign \new_[23638]_  = A269 & A266;
  assign \new_[23639]_  = ~A265 & \new_[23638]_ ;
  assign \new_[23640]_  = \new_[23639]_  & \new_[23634]_ ;
  assign \new_[23643]_  = ~A169 & ~A170;
  assign \new_[23647]_  = A201 & A199;
  assign \new_[23648]_  = ~A168 & \new_[23647]_ ;
  assign \new_[23649]_  = \new_[23648]_  & \new_[23643]_ ;
  assign \new_[23653]_  = A236 & A233;
  assign \new_[23654]_  = ~A232 & \new_[23653]_ ;
  assign \new_[23658]_  = A269 & ~A266;
  assign \new_[23659]_  = A265 & \new_[23658]_ ;
  assign \new_[23660]_  = \new_[23659]_  & \new_[23654]_ ;
  assign \new_[23663]_  = ~A169 & ~A170;
  assign \new_[23667]_  = A201 & A199;
  assign \new_[23668]_  = ~A168 & \new_[23667]_ ;
  assign \new_[23669]_  = \new_[23668]_  & \new_[23663]_ ;
  assign \new_[23673]_  = A236 & ~A233;
  assign \new_[23674]_  = A232 & \new_[23673]_ ;
  assign \new_[23678]_  = ~A302 & ~A301;
  assign \new_[23679]_  = ~A300 & \new_[23678]_ ;
  assign \new_[23680]_  = \new_[23679]_  & \new_[23674]_ ;
  assign \new_[23683]_  = ~A169 & ~A170;
  assign \new_[23687]_  = A201 & A199;
  assign \new_[23688]_  = ~A168 & \new_[23687]_ ;
  assign \new_[23689]_  = \new_[23688]_  & \new_[23683]_ ;
  assign \new_[23693]_  = A236 & ~A233;
  assign \new_[23694]_  = A232 & \new_[23693]_ ;
  assign \new_[23698]_  = ~A301 & ~A299;
  assign \new_[23699]_  = ~A298 & \new_[23698]_ ;
  assign \new_[23700]_  = \new_[23699]_  & \new_[23694]_ ;
  assign \new_[23703]_  = ~A169 & ~A170;
  assign \new_[23707]_  = A201 & A199;
  assign \new_[23708]_  = ~A168 & \new_[23707]_ ;
  assign \new_[23709]_  = \new_[23708]_  & \new_[23703]_ ;
  assign \new_[23713]_  = A236 & ~A233;
  assign \new_[23714]_  = A232 & \new_[23713]_ ;
  assign \new_[23718]_  = A269 & A266;
  assign \new_[23719]_  = ~A265 & \new_[23718]_ ;
  assign \new_[23720]_  = \new_[23719]_  & \new_[23714]_ ;
  assign \new_[23723]_  = ~A169 & ~A170;
  assign \new_[23727]_  = A201 & A199;
  assign \new_[23728]_  = ~A168 & \new_[23727]_ ;
  assign \new_[23729]_  = \new_[23728]_  & \new_[23723]_ ;
  assign \new_[23733]_  = A236 & ~A233;
  assign \new_[23734]_  = A232 & \new_[23733]_ ;
  assign \new_[23738]_  = A269 & ~A266;
  assign \new_[23739]_  = A265 & \new_[23738]_ ;
  assign \new_[23740]_  = \new_[23739]_  & \new_[23734]_ ;
  assign \new_[23743]_  = ~A169 & ~A170;
  assign \new_[23747]_  = A201 & A200;
  assign \new_[23748]_  = ~A168 & \new_[23747]_ ;
  assign \new_[23749]_  = \new_[23748]_  & \new_[23743]_ ;
  assign \new_[23753]_  = A298 & A234;
  assign \new_[23754]_  = A232 & \new_[23753]_ ;
  assign \new_[23758]_  = ~A301 & ~A300;
  assign \new_[23759]_  = A299 & \new_[23758]_ ;
  assign \new_[23760]_  = \new_[23759]_  & \new_[23754]_ ;
  assign \new_[23763]_  = ~A169 & ~A170;
  assign \new_[23767]_  = A201 & A200;
  assign \new_[23768]_  = ~A168 & \new_[23767]_ ;
  assign \new_[23769]_  = \new_[23768]_  & \new_[23763]_ ;
  assign \new_[23773]_  = A298 & A234;
  assign \new_[23774]_  = A233 & \new_[23773]_ ;
  assign \new_[23778]_  = ~A301 & ~A300;
  assign \new_[23779]_  = A299 & \new_[23778]_ ;
  assign \new_[23780]_  = \new_[23779]_  & \new_[23774]_ ;
  assign \new_[23783]_  = ~A169 & ~A170;
  assign \new_[23787]_  = A201 & A200;
  assign \new_[23788]_  = ~A168 & \new_[23787]_ ;
  assign \new_[23789]_  = \new_[23788]_  & \new_[23783]_ ;
  assign \new_[23793]_  = A236 & A233;
  assign \new_[23794]_  = ~A232 & \new_[23793]_ ;
  assign \new_[23798]_  = ~A302 & ~A301;
  assign \new_[23799]_  = ~A300 & \new_[23798]_ ;
  assign \new_[23800]_  = \new_[23799]_  & \new_[23794]_ ;
  assign \new_[23803]_  = ~A169 & ~A170;
  assign \new_[23807]_  = A201 & A200;
  assign \new_[23808]_  = ~A168 & \new_[23807]_ ;
  assign \new_[23809]_  = \new_[23808]_  & \new_[23803]_ ;
  assign \new_[23813]_  = A236 & A233;
  assign \new_[23814]_  = ~A232 & \new_[23813]_ ;
  assign \new_[23818]_  = ~A301 & ~A299;
  assign \new_[23819]_  = ~A298 & \new_[23818]_ ;
  assign \new_[23820]_  = \new_[23819]_  & \new_[23814]_ ;
  assign \new_[23823]_  = ~A169 & ~A170;
  assign \new_[23827]_  = A201 & A200;
  assign \new_[23828]_  = ~A168 & \new_[23827]_ ;
  assign \new_[23829]_  = \new_[23828]_  & \new_[23823]_ ;
  assign \new_[23833]_  = A236 & A233;
  assign \new_[23834]_  = ~A232 & \new_[23833]_ ;
  assign \new_[23838]_  = A269 & A266;
  assign \new_[23839]_  = ~A265 & \new_[23838]_ ;
  assign \new_[23840]_  = \new_[23839]_  & \new_[23834]_ ;
  assign \new_[23843]_  = ~A169 & ~A170;
  assign \new_[23847]_  = A201 & A200;
  assign \new_[23848]_  = ~A168 & \new_[23847]_ ;
  assign \new_[23849]_  = \new_[23848]_  & \new_[23843]_ ;
  assign \new_[23853]_  = A236 & A233;
  assign \new_[23854]_  = ~A232 & \new_[23853]_ ;
  assign \new_[23858]_  = A269 & ~A266;
  assign \new_[23859]_  = A265 & \new_[23858]_ ;
  assign \new_[23860]_  = \new_[23859]_  & \new_[23854]_ ;
  assign \new_[23863]_  = ~A169 & ~A170;
  assign \new_[23867]_  = A201 & A200;
  assign \new_[23868]_  = ~A168 & \new_[23867]_ ;
  assign \new_[23869]_  = \new_[23868]_  & \new_[23863]_ ;
  assign \new_[23873]_  = A236 & ~A233;
  assign \new_[23874]_  = A232 & \new_[23873]_ ;
  assign \new_[23878]_  = ~A302 & ~A301;
  assign \new_[23879]_  = ~A300 & \new_[23878]_ ;
  assign \new_[23880]_  = \new_[23879]_  & \new_[23874]_ ;
  assign \new_[23883]_  = ~A169 & ~A170;
  assign \new_[23887]_  = A201 & A200;
  assign \new_[23888]_  = ~A168 & \new_[23887]_ ;
  assign \new_[23889]_  = \new_[23888]_  & \new_[23883]_ ;
  assign \new_[23893]_  = A236 & ~A233;
  assign \new_[23894]_  = A232 & \new_[23893]_ ;
  assign \new_[23898]_  = ~A301 & ~A299;
  assign \new_[23899]_  = ~A298 & \new_[23898]_ ;
  assign \new_[23900]_  = \new_[23899]_  & \new_[23894]_ ;
  assign \new_[23903]_  = ~A169 & ~A170;
  assign \new_[23907]_  = A201 & A200;
  assign \new_[23908]_  = ~A168 & \new_[23907]_ ;
  assign \new_[23909]_  = \new_[23908]_  & \new_[23903]_ ;
  assign \new_[23913]_  = A236 & ~A233;
  assign \new_[23914]_  = A232 & \new_[23913]_ ;
  assign \new_[23918]_  = A269 & A266;
  assign \new_[23919]_  = ~A265 & \new_[23918]_ ;
  assign \new_[23920]_  = \new_[23919]_  & \new_[23914]_ ;
  assign \new_[23923]_  = ~A169 & ~A170;
  assign \new_[23927]_  = A201 & A200;
  assign \new_[23928]_  = ~A168 & \new_[23927]_ ;
  assign \new_[23929]_  = \new_[23928]_  & \new_[23923]_ ;
  assign \new_[23933]_  = A236 & ~A233;
  assign \new_[23934]_  = A232 & \new_[23933]_ ;
  assign \new_[23938]_  = A269 & ~A266;
  assign \new_[23939]_  = A265 & \new_[23938]_ ;
  assign \new_[23940]_  = \new_[23939]_  & \new_[23934]_ ;
  assign \new_[23943]_  = ~A169 & ~A170;
  assign \new_[23947]_  = A200 & ~A199;
  assign \new_[23948]_  = ~A168 & \new_[23947]_ ;
  assign \new_[23949]_  = \new_[23948]_  & \new_[23943]_ ;
  assign \new_[23953]_  = A298 & A235;
  assign \new_[23954]_  = A203 & \new_[23953]_ ;
  assign \new_[23958]_  = ~A301 & ~A300;
  assign \new_[23959]_  = A299 & \new_[23958]_ ;
  assign \new_[23960]_  = \new_[23959]_  & \new_[23954]_ ;
  assign \new_[23963]_  = ~A169 & ~A170;
  assign \new_[23967]_  = A200 & ~A199;
  assign \new_[23968]_  = ~A168 & \new_[23967]_ ;
  assign \new_[23969]_  = \new_[23968]_  & \new_[23963]_ ;
  assign \new_[23973]_  = A234 & A232;
  assign \new_[23974]_  = A203 & \new_[23973]_ ;
  assign \new_[23978]_  = ~A302 & ~A301;
  assign \new_[23979]_  = ~A300 & \new_[23978]_ ;
  assign \new_[23980]_  = \new_[23979]_  & \new_[23974]_ ;
  assign \new_[23983]_  = ~A169 & ~A170;
  assign \new_[23987]_  = A200 & ~A199;
  assign \new_[23988]_  = ~A168 & \new_[23987]_ ;
  assign \new_[23989]_  = \new_[23988]_  & \new_[23983]_ ;
  assign \new_[23993]_  = A234 & A232;
  assign \new_[23994]_  = A203 & \new_[23993]_ ;
  assign \new_[23998]_  = ~A301 & ~A299;
  assign \new_[23999]_  = ~A298 & \new_[23998]_ ;
  assign \new_[24000]_  = \new_[23999]_  & \new_[23994]_ ;
  assign \new_[24003]_  = ~A169 & ~A170;
  assign \new_[24007]_  = A200 & ~A199;
  assign \new_[24008]_  = ~A168 & \new_[24007]_ ;
  assign \new_[24009]_  = \new_[24008]_  & \new_[24003]_ ;
  assign \new_[24013]_  = A234 & A232;
  assign \new_[24014]_  = A203 & \new_[24013]_ ;
  assign \new_[24018]_  = A269 & A266;
  assign \new_[24019]_  = ~A265 & \new_[24018]_ ;
  assign \new_[24020]_  = \new_[24019]_  & \new_[24014]_ ;
  assign \new_[24023]_  = ~A169 & ~A170;
  assign \new_[24027]_  = A200 & ~A199;
  assign \new_[24028]_  = ~A168 & \new_[24027]_ ;
  assign \new_[24029]_  = \new_[24028]_  & \new_[24023]_ ;
  assign \new_[24033]_  = A234 & A232;
  assign \new_[24034]_  = A203 & \new_[24033]_ ;
  assign \new_[24038]_  = A269 & ~A266;
  assign \new_[24039]_  = A265 & \new_[24038]_ ;
  assign \new_[24040]_  = \new_[24039]_  & \new_[24034]_ ;
  assign \new_[24043]_  = ~A169 & ~A170;
  assign \new_[24047]_  = A200 & ~A199;
  assign \new_[24048]_  = ~A168 & \new_[24047]_ ;
  assign \new_[24049]_  = \new_[24048]_  & \new_[24043]_ ;
  assign \new_[24053]_  = A234 & A233;
  assign \new_[24054]_  = A203 & \new_[24053]_ ;
  assign \new_[24058]_  = ~A302 & ~A301;
  assign \new_[24059]_  = ~A300 & \new_[24058]_ ;
  assign \new_[24060]_  = \new_[24059]_  & \new_[24054]_ ;
  assign \new_[24063]_  = ~A169 & ~A170;
  assign \new_[24067]_  = A200 & ~A199;
  assign \new_[24068]_  = ~A168 & \new_[24067]_ ;
  assign \new_[24069]_  = \new_[24068]_  & \new_[24063]_ ;
  assign \new_[24073]_  = A234 & A233;
  assign \new_[24074]_  = A203 & \new_[24073]_ ;
  assign \new_[24078]_  = ~A301 & ~A299;
  assign \new_[24079]_  = ~A298 & \new_[24078]_ ;
  assign \new_[24080]_  = \new_[24079]_  & \new_[24074]_ ;
  assign \new_[24083]_  = ~A169 & ~A170;
  assign \new_[24087]_  = A200 & ~A199;
  assign \new_[24088]_  = ~A168 & \new_[24087]_ ;
  assign \new_[24089]_  = \new_[24088]_  & \new_[24083]_ ;
  assign \new_[24093]_  = A234 & A233;
  assign \new_[24094]_  = A203 & \new_[24093]_ ;
  assign \new_[24098]_  = A269 & A266;
  assign \new_[24099]_  = ~A265 & \new_[24098]_ ;
  assign \new_[24100]_  = \new_[24099]_  & \new_[24094]_ ;
  assign \new_[24103]_  = ~A169 & ~A170;
  assign \new_[24107]_  = A200 & ~A199;
  assign \new_[24108]_  = ~A168 & \new_[24107]_ ;
  assign \new_[24109]_  = \new_[24108]_  & \new_[24103]_ ;
  assign \new_[24113]_  = A234 & A233;
  assign \new_[24114]_  = A203 & \new_[24113]_ ;
  assign \new_[24118]_  = A269 & ~A266;
  assign \new_[24119]_  = A265 & \new_[24118]_ ;
  assign \new_[24120]_  = \new_[24119]_  & \new_[24114]_ ;
  assign \new_[24123]_  = ~A169 & ~A170;
  assign \new_[24127]_  = A200 & ~A199;
  assign \new_[24128]_  = ~A168 & \new_[24127]_ ;
  assign \new_[24129]_  = \new_[24128]_  & \new_[24123]_ ;
  assign \new_[24133]_  = A233 & ~A232;
  assign \new_[24134]_  = A203 & \new_[24133]_ ;
  assign \new_[24138]_  = A267 & A265;
  assign \new_[24139]_  = A236 & \new_[24138]_ ;
  assign \new_[24140]_  = \new_[24139]_  & \new_[24134]_ ;
  assign \new_[24143]_  = ~A169 & ~A170;
  assign \new_[24147]_  = A200 & ~A199;
  assign \new_[24148]_  = ~A168 & \new_[24147]_ ;
  assign \new_[24149]_  = \new_[24148]_  & \new_[24143]_ ;
  assign \new_[24153]_  = A233 & ~A232;
  assign \new_[24154]_  = A203 & \new_[24153]_ ;
  assign \new_[24158]_  = A267 & A266;
  assign \new_[24159]_  = A236 & \new_[24158]_ ;
  assign \new_[24160]_  = \new_[24159]_  & \new_[24154]_ ;
  assign \new_[24163]_  = ~A169 & ~A170;
  assign \new_[24167]_  = A200 & ~A199;
  assign \new_[24168]_  = ~A168 & \new_[24167]_ ;
  assign \new_[24169]_  = \new_[24168]_  & \new_[24163]_ ;
  assign \new_[24173]_  = ~A233 & A232;
  assign \new_[24174]_  = A203 & \new_[24173]_ ;
  assign \new_[24178]_  = A267 & A265;
  assign \new_[24179]_  = A236 & \new_[24178]_ ;
  assign \new_[24180]_  = \new_[24179]_  & \new_[24174]_ ;
  assign \new_[24183]_  = ~A169 & ~A170;
  assign \new_[24187]_  = A200 & ~A199;
  assign \new_[24188]_  = ~A168 & \new_[24187]_ ;
  assign \new_[24189]_  = \new_[24188]_  & \new_[24183]_ ;
  assign \new_[24193]_  = ~A233 & A232;
  assign \new_[24194]_  = A203 & \new_[24193]_ ;
  assign \new_[24198]_  = A267 & A266;
  assign \new_[24199]_  = A236 & \new_[24198]_ ;
  assign \new_[24200]_  = \new_[24199]_  & \new_[24194]_ ;
  assign \new_[24203]_  = ~A169 & ~A170;
  assign \new_[24207]_  = ~A200 & A199;
  assign \new_[24208]_  = ~A168 & \new_[24207]_ ;
  assign \new_[24209]_  = \new_[24208]_  & \new_[24203]_ ;
  assign \new_[24213]_  = A298 & A235;
  assign \new_[24214]_  = A203 & \new_[24213]_ ;
  assign \new_[24218]_  = ~A301 & ~A300;
  assign \new_[24219]_  = A299 & \new_[24218]_ ;
  assign \new_[24220]_  = \new_[24219]_  & \new_[24214]_ ;
  assign \new_[24223]_  = ~A169 & ~A170;
  assign \new_[24227]_  = ~A200 & A199;
  assign \new_[24228]_  = ~A168 & \new_[24227]_ ;
  assign \new_[24229]_  = \new_[24228]_  & \new_[24223]_ ;
  assign \new_[24233]_  = A234 & A232;
  assign \new_[24234]_  = A203 & \new_[24233]_ ;
  assign \new_[24238]_  = ~A302 & ~A301;
  assign \new_[24239]_  = ~A300 & \new_[24238]_ ;
  assign \new_[24240]_  = \new_[24239]_  & \new_[24234]_ ;
  assign \new_[24243]_  = ~A169 & ~A170;
  assign \new_[24247]_  = ~A200 & A199;
  assign \new_[24248]_  = ~A168 & \new_[24247]_ ;
  assign \new_[24249]_  = \new_[24248]_  & \new_[24243]_ ;
  assign \new_[24253]_  = A234 & A232;
  assign \new_[24254]_  = A203 & \new_[24253]_ ;
  assign \new_[24258]_  = ~A301 & ~A299;
  assign \new_[24259]_  = ~A298 & \new_[24258]_ ;
  assign \new_[24260]_  = \new_[24259]_  & \new_[24254]_ ;
  assign \new_[24263]_  = ~A169 & ~A170;
  assign \new_[24267]_  = ~A200 & A199;
  assign \new_[24268]_  = ~A168 & \new_[24267]_ ;
  assign \new_[24269]_  = \new_[24268]_  & \new_[24263]_ ;
  assign \new_[24273]_  = A234 & A232;
  assign \new_[24274]_  = A203 & \new_[24273]_ ;
  assign \new_[24278]_  = A269 & A266;
  assign \new_[24279]_  = ~A265 & \new_[24278]_ ;
  assign \new_[24280]_  = \new_[24279]_  & \new_[24274]_ ;
  assign \new_[24283]_  = ~A169 & ~A170;
  assign \new_[24287]_  = ~A200 & A199;
  assign \new_[24288]_  = ~A168 & \new_[24287]_ ;
  assign \new_[24289]_  = \new_[24288]_  & \new_[24283]_ ;
  assign \new_[24293]_  = A234 & A232;
  assign \new_[24294]_  = A203 & \new_[24293]_ ;
  assign \new_[24298]_  = A269 & ~A266;
  assign \new_[24299]_  = A265 & \new_[24298]_ ;
  assign \new_[24300]_  = \new_[24299]_  & \new_[24294]_ ;
  assign \new_[24303]_  = ~A169 & ~A170;
  assign \new_[24307]_  = ~A200 & A199;
  assign \new_[24308]_  = ~A168 & \new_[24307]_ ;
  assign \new_[24309]_  = \new_[24308]_  & \new_[24303]_ ;
  assign \new_[24313]_  = A234 & A233;
  assign \new_[24314]_  = A203 & \new_[24313]_ ;
  assign \new_[24318]_  = ~A302 & ~A301;
  assign \new_[24319]_  = ~A300 & \new_[24318]_ ;
  assign \new_[24320]_  = \new_[24319]_  & \new_[24314]_ ;
  assign \new_[24323]_  = ~A169 & ~A170;
  assign \new_[24327]_  = ~A200 & A199;
  assign \new_[24328]_  = ~A168 & \new_[24327]_ ;
  assign \new_[24329]_  = \new_[24328]_  & \new_[24323]_ ;
  assign \new_[24333]_  = A234 & A233;
  assign \new_[24334]_  = A203 & \new_[24333]_ ;
  assign \new_[24338]_  = ~A301 & ~A299;
  assign \new_[24339]_  = ~A298 & \new_[24338]_ ;
  assign \new_[24340]_  = \new_[24339]_  & \new_[24334]_ ;
  assign \new_[24343]_  = ~A169 & ~A170;
  assign \new_[24347]_  = ~A200 & A199;
  assign \new_[24348]_  = ~A168 & \new_[24347]_ ;
  assign \new_[24349]_  = \new_[24348]_  & \new_[24343]_ ;
  assign \new_[24353]_  = A234 & A233;
  assign \new_[24354]_  = A203 & \new_[24353]_ ;
  assign \new_[24358]_  = A269 & A266;
  assign \new_[24359]_  = ~A265 & \new_[24358]_ ;
  assign \new_[24360]_  = \new_[24359]_  & \new_[24354]_ ;
  assign \new_[24363]_  = ~A169 & ~A170;
  assign \new_[24367]_  = ~A200 & A199;
  assign \new_[24368]_  = ~A168 & \new_[24367]_ ;
  assign \new_[24369]_  = \new_[24368]_  & \new_[24363]_ ;
  assign \new_[24373]_  = A234 & A233;
  assign \new_[24374]_  = A203 & \new_[24373]_ ;
  assign \new_[24378]_  = A269 & ~A266;
  assign \new_[24379]_  = A265 & \new_[24378]_ ;
  assign \new_[24380]_  = \new_[24379]_  & \new_[24374]_ ;
  assign \new_[24383]_  = ~A169 & ~A170;
  assign \new_[24387]_  = ~A200 & A199;
  assign \new_[24388]_  = ~A168 & \new_[24387]_ ;
  assign \new_[24389]_  = \new_[24388]_  & \new_[24383]_ ;
  assign \new_[24393]_  = A233 & ~A232;
  assign \new_[24394]_  = A203 & \new_[24393]_ ;
  assign \new_[24398]_  = A267 & A265;
  assign \new_[24399]_  = A236 & \new_[24398]_ ;
  assign \new_[24400]_  = \new_[24399]_  & \new_[24394]_ ;
  assign \new_[24403]_  = ~A169 & ~A170;
  assign \new_[24407]_  = ~A200 & A199;
  assign \new_[24408]_  = ~A168 & \new_[24407]_ ;
  assign \new_[24409]_  = \new_[24408]_  & \new_[24403]_ ;
  assign \new_[24413]_  = A233 & ~A232;
  assign \new_[24414]_  = A203 & \new_[24413]_ ;
  assign \new_[24418]_  = A267 & A266;
  assign \new_[24419]_  = A236 & \new_[24418]_ ;
  assign \new_[24420]_  = \new_[24419]_  & \new_[24414]_ ;
  assign \new_[24423]_  = ~A169 & ~A170;
  assign \new_[24427]_  = ~A200 & A199;
  assign \new_[24428]_  = ~A168 & \new_[24427]_ ;
  assign \new_[24429]_  = \new_[24428]_  & \new_[24423]_ ;
  assign \new_[24433]_  = ~A233 & A232;
  assign \new_[24434]_  = A203 & \new_[24433]_ ;
  assign \new_[24438]_  = A267 & A265;
  assign \new_[24439]_  = A236 & \new_[24438]_ ;
  assign \new_[24440]_  = \new_[24439]_  & \new_[24434]_ ;
  assign \new_[24443]_  = ~A169 & ~A170;
  assign \new_[24447]_  = ~A200 & A199;
  assign \new_[24448]_  = ~A168 & \new_[24447]_ ;
  assign \new_[24449]_  = \new_[24448]_  & \new_[24443]_ ;
  assign \new_[24453]_  = ~A233 & A232;
  assign \new_[24454]_  = A203 & \new_[24453]_ ;
  assign \new_[24458]_  = A267 & A266;
  assign \new_[24459]_  = A236 & \new_[24458]_ ;
  assign \new_[24460]_  = \new_[24459]_  & \new_[24454]_ ;
  assign \new_[24464]_  = ~A201 & A166;
  assign \new_[24465]_  = A168 & \new_[24464]_ ;
  assign \new_[24469]_  = ~A234 & ~A203;
  assign \new_[24470]_  = ~A202 & \new_[24469]_ ;
  assign \new_[24471]_  = \new_[24470]_  & \new_[24465]_ ;
  assign \new_[24475]_  = ~A267 & ~A236;
  assign \new_[24476]_  = ~A235 & \new_[24475]_ ;
  assign \new_[24480]_  = A301 & ~A269;
  assign \new_[24481]_  = ~A268 & \new_[24480]_ ;
  assign \new_[24482]_  = \new_[24481]_  & \new_[24476]_ ;
  assign \new_[24486]_  = ~A201 & A166;
  assign \new_[24487]_  = A168 & \new_[24486]_ ;
  assign \new_[24491]_  = ~A234 & ~A203;
  assign \new_[24492]_  = ~A202 & \new_[24491]_ ;
  assign \new_[24493]_  = \new_[24492]_  & \new_[24487]_ ;
  assign \new_[24497]_  = ~A265 & ~A236;
  assign \new_[24498]_  = ~A235 & \new_[24497]_ ;
  assign \new_[24502]_  = A301 & ~A268;
  assign \new_[24503]_  = ~A266 & \new_[24502]_ ;
  assign \new_[24504]_  = \new_[24503]_  & \new_[24498]_ ;
  assign \new_[24508]_  = ~A201 & A166;
  assign \new_[24509]_  = A168 & \new_[24508]_ ;
  assign \new_[24513]_  = ~A232 & ~A203;
  assign \new_[24514]_  = ~A202 & \new_[24513]_ ;
  assign \new_[24515]_  = \new_[24514]_  & \new_[24509]_ ;
  assign \new_[24519]_  = A298 & A236;
  assign \new_[24520]_  = A233 & \new_[24519]_ ;
  assign \new_[24524]_  = ~A301 & ~A300;
  assign \new_[24525]_  = A299 & \new_[24524]_ ;
  assign \new_[24526]_  = \new_[24525]_  & \new_[24520]_ ;
  assign \new_[24530]_  = ~A201 & A166;
  assign \new_[24531]_  = A168 & \new_[24530]_ ;
  assign \new_[24535]_  = A232 & ~A203;
  assign \new_[24536]_  = ~A202 & \new_[24535]_ ;
  assign \new_[24537]_  = \new_[24536]_  & \new_[24531]_ ;
  assign \new_[24541]_  = A298 & A236;
  assign \new_[24542]_  = ~A233 & \new_[24541]_ ;
  assign \new_[24546]_  = ~A301 & ~A300;
  assign \new_[24547]_  = A299 & \new_[24546]_ ;
  assign \new_[24548]_  = \new_[24547]_  & \new_[24542]_ ;
  assign \new_[24552]_  = ~A201 & A166;
  assign \new_[24553]_  = A168 & \new_[24552]_ ;
  assign \new_[24557]_  = ~A232 & ~A203;
  assign \new_[24558]_  = ~A202 & \new_[24557]_ ;
  assign \new_[24559]_  = \new_[24558]_  & \new_[24553]_ ;
  assign \new_[24563]_  = ~A267 & ~A235;
  assign \new_[24564]_  = ~A233 & \new_[24563]_ ;
  assign \new_[24568]_  = A301 & ~A269;
  assign \new_[24569]_  = ~A268 & \new_[24568]_ ;
  assign \new_[24570]_  = \new_[24569]_  & \new_[24564]_ ;
  assign \new_[24574]_  = ~A201 & A166;
  assign \new_[24575]_  = A168 & \new_[24574]_ ;
  assign \new_[24579]_  = ~A232 & ~A203;
  assign \new_[24580]_  = ~A202 & \new_[24579]_ ;
  assign \new_[24581]_  = \new_[24580]_  & \new_[24575]_ ;
  assign \new_[24585]_  = ~A265 & ~A235;
  assign \new_[24586]_  = ~A233 & \new_[24585]_ ;
  assign \new_[24590]_  = A301 & ~A268;
  assign \new_[24591]_  = ~A266 & \new_[24590]_ ;
  assign \new_[24592]_  = \new_[24591]_  & \new_[24586]_ ;
  assign \new_[24596]_  = A199 & A166;
  assign \new_[24597]_  = A168 & \new_[24596]_ ;
  assign \new_[24601]_  = ~A202 & ~A201;
  assign \new_[24602]_  = A200 & \new_[24601]_ ;
  assign \new_[24603]_  = \new_[24602]_  & \new_[24597]_ ;
  assign \new_[24607]_  = A298 & A234;
  assign \new_[24608]_  = A232 & \new_[24607]_ ;
  assign \new_[24612]_  = ~A301 & ~A300;
  assign \new_[24613]_  = A299 & \new_[24612]_ ;
  assign \new_[24614]_  = \new_[24613]_  & \new_[24608]_ ;
  assign \new_[24618]_  = A199 & A166;
  assign \new_[24619]_  = A168 & \new_[24618]_ ;
  assign \new_[24623]_  = ~A202 & ~A201;
  assign \new_[24624]_  = A200 & \new_[24623]_ ;
  assign \new_[24625]_  = \new_[24624]_  & \new_[24619]_ ;
  assign \new_[24629]_  = A298 & A234;
  assign \new_[24630]_  = A233 & \new_[24629]_ ;
  assign \new_[24634]_  = ~A301 & ~A300;
  assign \new_[24635]_  = A299 & \new_[24634]_ ;
  assign \new_[24636]_  = \new_[24635]_  & \new_[24630]_ ;
  assign \new_[24640]_  = A199 & A166;
  assign \new_[24641]_  = A168 & \new_[24640]_ ;
  assign \new_[24645]_  = ~A202 & ~A201;
  assign \new_[24646]_  = A200 & \new_[24645]_ ;
  assign \new_[24647]_  = \new_[24646]_  & \new_[24641]_ ;
  assign \new_[24651]_  = A236 & A233;
  assign \new_[24652]_  = ~A232 & \new_[24651]_ ;
  assign \new_[24656]_  = ~A302 & ~A301;
  assign \new_[24657]_  = ~A300 & \new_[24656]_ ;
  assign \new_[24658]_  = \new_[24657]_  & \new_[24652]_ ;
  assign \new_[24662]_  = A199 & A166;
  assign \new_[24663]_  = A168 & \new_[24662]_ ;
  assign \new_[24667]_  = ~A202 & ~A201;
  assign \new_[24668]_  = A200 & \new_[24667]_ ;
  assign \new_[24669]_  = \new_[24668]_  & \new_[24663]_ ;
  assign \new_[24673]_  = A236 & A233;
  assign \new_[24674]_  = ~A232 & \new_[24673]_ ;
  assign \new_[24678]_  = ~A301 & ~A299;
  assign \new_[24679]_  = ~A298 & \new_[24678]_ ;
  assign \new_[24680]_  = \new_[24679]_  & \new_[24674]_ ;
  assign \new_[24684]_  = A199 & A166;
  assign \new_[24685]_  = A168 & \new_[24684]_ ;
  assign \new_[24689]_  = ~A202 & ~A201;
  assign \new_[24690]_  = A200 & \new_[24689]_ ;
  assign \new_[24691]_  = \new_[24690]_  & \new_[24685]_ ;
  assign \new_[24695]_  = A236 & A233;
  assign \new_[24696]_  = ~A232 & \new_[24695]_ ;
  assign \new_[24700]_  = A269 & A266;
  assign \new_[24701]_  = ~A265 & \new_[24700]_ ;
  assign \new_[24702]_  = \new_[24701]_  & \new_[24696]_ ;
  assign \new_[24706]_  = A199 & A166;
  assign \new_[24707]_  = A168 & \new_[24706]_ ;
  assign \new_[24711]_  = ~A202 & ~A201;
  assign \new_[24712]_  = A200 & \new_[24711]_ ;
  assign \new_[24713]_  = \new_[24712]_  & \new_[24707]_ ;
  assign \new_[24717]_  = A236 & A233;
  assign \new_[24718]_  = ~A232 & \new_[24717]_ ;
  assign \new_[24722]_  = A269 & ~A266;
  assign \new_[24723]_  = A265 & \new_[24722]_ ;
  assign \new_[24724]_  = \new_[24723]_  & \new_[24718]_ ;
  assign \new_[24728]_  = A199 & A166;
  assign \new_[24729]_  = A168 & \new_[24728]_ ;
  assign \new_[24733]_  = ~A202 & ~A201;
  assign \new_[24734]_  = A200 & \new_[24733]_ ;
  assign \new_[24735]_  = \new_[24734]_  & \new_[24729]_ ;
  assign \new_[24739]_  = A236 & ~A233;
  assign \new_[24740]_  = A232 & \new_[24739]_ ;
  assign \new_[24744]_  = ~A302 & ~A301;
  assign \new_[24745]_  = ~A300 & \new_[24744]_ ;
  assign \new_[24746]_  = \new_[24745]_  & \new_[24740]_ ;
  assign \new_[24750]_  = A199 & A166;
  assign \new_[24751]_  = A168 & \new_[24750]_ ;
  assign \new_[24755]_  = ~A202 & ~A201;
  assign \new_[24756]_  = A200 & \new_[24755]_ ;
  assign \new_[24757]_  = \new_[24756]_  & \new_[24751]_ ;
  assign \new_[24761]_  = A236 & ~A233;
  assign \new_[24762]_  = A232 & \new_[24761]_ ;
  assign \new_[24766]_  = ~A301 & ~A299;
  assign \new_[24767]_  = ~A298 & \new_[24766]_ ;
  assign \new_[24768]_  = \new_[24767]_  & \new_[24762]_ ;
  assign \new_[24772]_  = A199 & A166;
  assign \new_[24773]_  = A168 & \new_[24772]_ ;
  assign \new_[24777]_  = ~A202 & ~A201;
  assign \new_[24778]_  = A200 & \new_[24777]_ ;
  assign \new_[24779]_  = \new_[24778]_  & \new_[24773]_ ;
  assign \new_[24783]_  = A236 & ~A233;
  assign \new_[24784]_  = A232 & \new_[24783]_ ;
  assign \new_[24788]_  = A269 & A266;
  assign \new_[24789]_  = ~A265 & \new_[24788]_ ;
  assign \new_[24790]_  = \new_[24789]_  & \new_[24784]_ ;
  assign \new_[24794]_  = A199 & A166;
  assign \new_[24795]_  = A168 & \new_[24794]_ ;
  assign \new_[24799]_  = ~A202 & ~A201;
  assign \new_[24800]_  = A200 & \new_[24799]_ ;
  assign \new_[24801]_  = \new_[24800]_  & \new_[24795]_ ;
  assign \new_[24805]_  = A236 & ~A233;
  assign \new_[24806]_  = A232 & \new_[24805]_ ;
  assign \new_[24810]_  = A269 & ~A266;
  assign \new_[24811]_  = A265 & \new_[24810]_ ;
  assign \new_[24812]_  = \new_[24811]_  & \new_[24806]_ ;
  assign \new_[24816]_  = ~A199 & A166;
  assign \new_[24817]_  = A168 & \new_[24816]_ ;
  assign \new_[24821]_  = ~A234 & ~A202;
  assign \new_[24822]_  = ~A200 & \new_[24821]_ ;
  assign \new_[24823]_  = \new_[24822]_  & \new_[24817]_ ;
  assign \new_[24827]_  = ~A267 & ~A236;
  assign \new_[24828]_  = ~A235 & \new_[24827]_ ;
  assign \new_[24832]_  = A301 & ~A269;
  assign \new_[24833]_  = ~A268 & \new_[24832]_ ;
  assign \new_[24834]_  = \new_[24833]_  & \new_[24828]_ ;
  assign \new_[24838]_  = ~A199 & A166;
  assign \new_[24839]_  = A168 & \new_[24838]_ ;
  assign \new_[24843]_  = ~A234 & ~A202;
  assign \new_[24844]_  = ~A200 & \new_[24843]_ ;
  assign \new_[24845]_  = \new_[24844]_  & \new_[24839]_ ;
  assign \new_[24849]_  = ~A265 & ~A236;
  assign \new_[24850]_  = ~A235 & \new_[24849]_ ;
  assign \new_[24854]_  = A301 & ~A268;
  assign \new_[24855]_  = ~A266 & \new_[24854]_ ;
  assign \new_[24856]_  = \new_[24855]_  & \new_[24850]_ ;
  assign \new_[24860]_  = ~A199 & A166;
  assign \new_[24861]_  = A168 & \new_[24860]_ ;
  assign \new_[24865]_  = ~A232 & ~A202;
  assign \new_[24866]_  = ~A200 & \new_[24865]_ ;
  assign \new_[24867]_  = \new_[24866]_  & \new_[24861]_ ;
  assign \new_[24871]_  = A298 & A236;
  assign \new_[24872]_  = A233 & \new_[24871]_ ;
  assign \new_[24876]_  = ~A301 & ~A300;
  assign \new_[24877]_  = A299 & \new_[24876]_ ;
  assign \new_[24878]_  = \new_[24877]_  & \new_[24872]_ ;
  assign \new_[24882]_  = ~A199 & A166;
  assign \new_[24883]_  = A168 & \new_[24882]_ ;
  assign \new_[24887]_  = A232 & ~A202;
  assign \new_[24888]_  = ~A200 & \new_[24887]_ ;
  assign \new_[24889]_  = \new_[24888]_  & \new_[24883]_ ;
  assign \new_[24893]_  = A298 & A236;
  assign \new_[24894]_  = ~A233 & \new_[24893]_ ;
  assign \new_[24898]_  = ~A301 & ~A300;
  assign \new_[24899]_  = A299 & \new_[24898]_ ;
  assign \new_[24900]_  = \new_[24899]_  & \new_[24894]_ ;
  assign \new_[24904]_  = ~A199 & A166;
  assign \new_[24905]_  = A168 & \new_[24904]_ ;
  assign \new_[24909]_  = ~A232 & ~A202;
  assign \new_[24910]_  = ~A200 & \new_[24909]_ ;
  assign \new_[24911]_  = \new_[24910]_  & \new_[24905]_ ;
  assign \new_[24915]_  = ~A267 & ~A235;
  assign \new_[24916]_  = ~A233 & \new_[24915]_ ;
  assign \new_[24920]_  = A301 & ~A269;
  assign \new_[24921]_  = ~A268 & \new_[24920]_ ;
  assign \new_[24922]_  = \new_[24921]_  & \new_[24916]_ ;
  assign \new_[24926]_  = ~A199 & A166;
  assign \new_[24927]_  = A168 & \new_[24926]_ ;
  assign \new_[24931]_  = ~A232 & ~A202;
  assign \new_[24932]_  = ~A200 & \new_[24931]_ ;
  assign \new_[24933]_  = \new_[24932]_  & \new_[24927]_ ;
  assign \new_[24937]_  = ~A265 & ~A235;
  assign \new_[24938]_  = ~A233 & \new_[24937]_ ;
  assign \new_[24942]_  = A301 & ~A268;
  assign \new_[24943]_  = ~A266 & \new_[24942]_ ;
  assign \new_[24944]_  = \new_[24943]_  & \new_[24938]_ ;
  assign \new_[24948]_  = ~A201 & A167;
  assign \new_[24949]_  = A168 & \new_[24948]_ ;
  assign \new_[24953]_  = ~A234 & ~A203;
  assign \new_[24954]_  = ~A202 & \new_[24953]_ ;
  assign \new_[24955]_  = \new_[24954]_  & \new_[24949]_ ;
  assign \new_[24959]_  = ~A267 & ~A236;
  assign \new_[24960]_  = ~A235 & \new_[24959]_ ;
  assign \new_[24964]_  = A301 & ~A269;
  assign \new_[24965]_  = ~A268 & \new_[24964]_ ;
  assign \new_[24966]_  = \new_[24965]_  & \new_[24960]_ ;
  assign \new_[24970]_  = ~A201 & A167;
  assign \new_[24971]_  = A168 & \new_[24970]_ ;
  assign \new_[24975]_  = ~A234 & ~A203;
  assign \new_[24976]_  = ~A202 & \new_[24975]_ ;
  assign \new_[24977]_  = \new_[24976]_  & \new_[24971]_ ;
  assign \new_[24981]_  = ~A265 & ~A236;
  assign \new_[24982]_  = ~A235 & \new_[24981]_ ;
  assign \new_[24986]_  = A301 & ~A268;
  assign \new_[24987]_  = ~A266 & \new_[24986]_ ;
  assign \new_[24988]_  = \new_[24987]_  & \new_[24982]_ ;
  assign \new_[24992]_  = ~A201 & A167;
  assign \new_[24993]_  = A168 & \new_[24992]_ ;
  assign \new_[24997]_  = ~A232 & ~A203;
  assign \new_[24998]_  = ~A202 & \new_[24997]_ ;
  assign \new_[24999]_  = \new_[24998]_  & \new_[24993]_ ;
  assign \new_[25003]_  = A298 & A236;
  assign \new_[25004]_  = A233 & \new_[25003]_ ;
  assign \new_[25008]_  = ~A301 & ~A300;
  assign \new_[25009]_  = A299 & \new_[25008]_ ;
  assign \new_[25010]_  = \new_[25009]_  & \new_[25004]_ ;
  assign \new_[25014]_  = ~A201 & A167;
  assign \new_[25015]_  = A168 & \new_[25014]_ ;
  assign \new_[25019]_  = A232 & ~A203;
  assign \new_[25020]_  = ~A202 & \new_[25019]_ ;
  assign \new_[25021]_  = \new_[25020]_  & \new_[25015]_ ;
  assign \new_[25025]_  = A298 & A236;
  assign \new_[25026]_  = ~A233 & \new_[25025]_ ;
  assign \new_[25030]_  = ~A301 & ~A300;
  assign \new_[25031]_  = A299 & \new_[25030]_ ;
  assign \new_[25032]_  = \new_[25031]_  & \new_[25026]_ ;
  assign \new_[25036]_  = ~A201 & A167;
  assign \new_[25037]_  = A168 & \new_[25036]_ ;
  assign \new_[25041]_  = ~A232 & ~A203;
  assign \new_[25042]_  = ~A202 & \new_[25041]_ ;
  assign \new_[25043]_  = \new_[25042]_  & \new_[25037]_ ;
  assign \new_[25047]_  = ~A267 & ~A235;
  assign \new_[25048]_  = ~A233 & \new_[25047]_ ;
  assign \new_[25052]_  = A301 & ~A269;
  assign \new_[25053]_  = ~A268 & \new_[25052]_ ;
  assign \new_[25054]_  = \new_[25053]_  & \new_[25048]_ ;
  assign \new_[25058]_  = ~A201 & A167;
  assign \new_[25059]_  = A168 & \new_[25058]_ ;
  assign \new_[25063]_  = ~A232 & ~A203;
  assign \new_[25064]_  = ~A202 & \new_[25063]_ ;
  assign \new_[25065]_  = \new_[25064]_  & \new_[25059]_ ;
  assign \new_[25069]_  = ~A265 & ~A235;
  assign \new_[25070]_  = ~A233 & \new_[25069]_ ;
  assign \new_[25074]_  = A301 & ~A268;
  assign \new_[25075]_  = ~A266 & \new_[25074]_ ;
  assign \new_[25076]_  = \new_[25075]_  & \new_[25070]_ ;
  assign \new_[25080]_  = A199 & A167;
  assign \new_[25081]_  = A168 & \new_[25080]_ ;
  assign \new_[25085]_  = ~A202 & ~A201;
  assign \new_[25086]_  = A200 & \new_[25085]_ ;
  assign \new_[25087]_  = \new_[25086]_  & \new_[25081]_ ;
  assign \new_[25091]_  = A298 & A234;
  assign \new_[25092]_  = A232 & \new_[25091]_ ;
  assign \new_[25096]_  = ~A301 & ~A300;
  assign \new_[25097]_  = A299 & \new_[25096]_ ;
  assign \new_[25098]_  = \new_[25097]_  & \new_[25092]_ ;
  assign \new_[25102]_  = A199 & A167;
  assign \new_[25103]_  = A168 & \new_[25102]_ ;
  assign \new_[25107]_  = ~A202 & ~A201;
  assign \new_[25108]_  = A200 & \new_[25107]_ ;
  assign \new_[25109]_  = \new_[25108]_  & \new_[25103]_ ;
  assign \new_[25113]_  = A298 & A234;
  assign \new_[25114]_  = A233 & \new_[25113]_ ;
  assign \new_[25118]_  = ~A301 & ~A300;
  assign \new_[25119]_  = A299 & \new_[25118]_ ;
  assign \new_[25120]_  = \new_[25119]_  & \new_[25114]_ ;
  assign \new_[25124]_  = A199 & A167;
  assign \new_[25125]_  = A168 & \new_[25124]_ ;
  assign \new_[25129]_  = ~A202 & ~A201;
  assign \new_[25130]_  = A200 & \new_[25129]_ ;
  assign \new_[25131]_  = \new_[25130]_  & \new_[25125]_ ;
  assign \new_[25135]_  = A236 & A233;
  assign \new_[25136]_  = ~A232 & \new_[25135]_ ;
  assign \new_[25140]_  = ~A302 & ~A301;
  assign \new_[25141]_  = ~A300 & \new_[25140]_ ;
  assign \new_[25142]_  = \new_[25141]_  & \new_[25136]_ ;
  assign \new_[25146]_  = A199 & A167;
  assign \new_[25147]_  = A168 & \new_[25146]_ ;
  assign \new_[25151]_  = ~A202 & ~A201;
  assign \new_[25152]_  = A200 & \new_[25151]_ ;
  assign \new_[25153]_  = \new_[25152]_  & \new_[25147]_ ;
  assign \new_[25157]_  = A236 & A233;
  assign \new_[25158]_  = ~A232 & \new_[25157]_ ;
  assign \new_[25162]_  = ~A301 & ~A299;
  assign \new_[25163]_  = ~A298 & \new_[25162]_ ;
  assign \new_[25164]_  = \new_[25163]_  & \new_[25158]_ ;
  assign \new_[25168]_  = A199 & A167;
  assign \new_[25169]_  = A168 & \new_[25168]_ ;
  assign \new_[25173]_  = ~A202 & ~A201;
  assign \new_[25174]_  = A200 & \new_[25173]_ ;
  assign \new_[25175]_  = \new_[25174]_  & \new_[25169]_ ;
  assign \new_[25179]_  = A236 & A233;
  assign \new_[25180]_  = ~A232 & \new_[25179]_ ;
  assign \new_[25184]_  = A269 & A266;
  assign \new_[25185]_  = ~A265 & \new_[25184]_ ;
  assign \new_[25186]_  = \new_[25185]_  & \new_[25180]_ ;
  assign \new_[25190]_  = A199 & A167;
  assign \new_[25191]_  = A168 & \new_[25190]_ ;
  assign \new_[25195]_  = ~A202 & ~A201;
  assign \new_[25196]_  = A200 & \new_[25195]_ ;
  assign \new_[25197]_  = \new_[25196]_  & \new_[25191]_ ;
  assign \new_[25201]_  = A236 & A233;
  assign \new_[25202]_  = ~A232 & \new_[25201]_ ;
  assign \new_[25206]_  = A269 & ~A266;
  assign \new_[25207]_  = A265 & \new_[25206]_ ;
  assign \new_[25208]_  = \new_[25207]_  & \new_[25202]_ ;
  assign \new_[25212]_  = A199 & A167;
  assign \new_[25213]_  = A168 & \new_[25212]_ ;
  assign \new_[25217]_  = ~A202 & ~A201;
  assign \new_[25218]_  = A200 & \new_[25217]_ ;
  assign \new_[25219]_  = \new_[25218]_  & \new_[25213]_ ;
  assign \new_[25223]_  = A236 & ~A233;
  assign \new_[25224]_  = A232 & \new_[25223]_ ;
  assign \new_[25228]_  = ~A302 & ~A301;
  assign \new_[25229]_  = ~A300 & \new_[25228]_ ;
  assign \new_[25230]_  = \new_[25229]_  & \new_[25224]_ ;
  assign \new_[25234]_  = A199 & A167;
  assign \new_[25235]_  = A168 & \new_[25234]_ ;
  assign \new_[25239]_  = ~A202 & ~A201;
  assign \new_[25240]_  = A200 & \new_[25239]_ ;
  assign \new_[25241]_  = \new_[25240]_  & \new_[25235]_ ;
  assign \new_[25245]_  = A236 & ~A233;
  assign \new_[25246]_  = A232 & \new_[25245]_ ;
  assign \new_[25250]_  = ~A301 & ~A299;
  assign \new_[25251]_  = ~A298 & \new_[25250]_ ;
  assign \new_[25252]_  = \new_[25251]_  & \new_[25246]_ ;
  assign \new_[25256]_  = A199 & A167;
  assign \new_[25257]_  = A168 & \new_[25256]_ ;
  assign \new_[25261]_  = ~A202 & ~A201;
  assign \new_[25262]_  = A200 & \new_[25261]_ ;
  assign \new_[25263]_  = \new_[25262]_  & \new_[25257]_ ;
  assign \new_[25267]_  = A236 & ~A233;
  assign \new_[25268]_  = A232 & \new_[25267]_ ;
  assign \new_[25272]_  = A269 & A266;
  assign \new_[25273]_  = ~A265 & \new_[25272]_ ;
  assign \new_[25274]_  = \new_[25273]_  & \new_[25268]_ ;
  assign \new_[25278]_  = A199 & A167;
  assign \new_[25279]_  = A168 & \new_[25278]_ ;
  assign \new_[25283]_  = ~A202 & ~A201;
  assign \new_[25284]_  = A200 & \new_[25283]_ ;
  assign \new_[25285]_  = \new_[25284]_  & \new_[25279]_ ;
  assign \new_[25289]_  = A236 & ~A233;
  assign \new_[25290]_  = A232 & \new_[25289]_ ;
  assign \new_[25294]_  = A269 & ~A266;
  assign \new_[25295]_  = A265 & \new_[25294]_ ;
  assign \new_[25296]_  = \new_[25295]_  & \new_[25290]_ ;
  assign \new_[25300]_  = ~A199 & A167;
  assign \new_[25301]_  = A168 & \new_[25300]_ ;
  assign \new_[25305]_  = ~A234 & ~A202;
  assign \new_[25306]_  = ~A200 & \new_[25305]_ ;
  assign \new_[25307]_  = \new_[25306]_  & \new_[25301]_ ;
  assign \new_[25311]_  = ~A267 & ~A236;
  assign \new_[25312]_  = ~A235 & \new_[25311]_ ;
  assign \new_[25316]_  = A301 & ~A269;
  assign \new_[25317]_  = ~A268 & \new_[25316]_ ;
  assign \new_[25318]_  = \new_[25317]_  & \new_[25312]_ ;
  assign \new_[25322]_  = ~A199 & A167;
  assign \new_[25323]_  = A168 & \new_[25322]_ ;
  assign \new_[25327]_  = ~A234 & ~A202;
  assign \new_[25328]_  = ~A200 & \new_[25327]_ ;
  assign \new_[25329]_  = \new_[25328]_  & \new_[25323]_ ;
  assign \new_[25333]_  = ~A265 & ~A236;
  assign \new_[25334]_  = ~A235 & \new_[25333]_ ;
  assign \new_[25338]_  = A301 & ~A268;
  assign \new_[25339]_  = ~A266 & \new_[25338]_ ;
  assign \new_[25340]_  = \new_[25339]_  & \new_[25334]_ ;
  assign \new_[25344]_  = ~A199 & A167;
  assign \new_[25345]_  = A168 & \new_[25344]_ ;
  assign \new_[25349]_  = ~A232 & ~A202;
  assign \new_[25350]_  = ~A200 & \new_[25349]_ ;
  assign \new_[25351]_  = \new_[25350]_  & \new_[25345]_ ;
  assign \new_[25355]_  = A298 & A236;
  assign \new_[25356]_  = A233 & \new_[25355]_ ;
  assign \new_[25360]_  = ~A301 & ~A300;
  assign \new_[25361]_  = A299 & \new_[25360]_ ;
  assign \new_[25362]_  = \new_[25361]_  & \new_[25356]_ ;
  assign \new_[25366]_  = ~A199 & A167;
  assign \new_[25367]_  = A168 & \new_[25366]_ ;
  assign \new_[25371]_  = A232 & ~A202;
  assign \new_[25372]_  = ~A200 & \new_[25371]_ ;
  assign \new_[25373]_  = \new_[25372]_  & \new_[25367]_ ;
  assign \new_[25377]_  = A298 & A236;
  assign \new_[25378]_  = ~A233 & \new_[25377]_ ;
  assign \new_[25382]_  = ~A301 & ~A300;
  assign \new_[25383]_  = A299 & \new_[25382]_ ;
  assign \new_[25384]_  = \new_[25383]_  & \new_[25378]_ ;
  assign \new_[25388]_  = ~A199 & A167;
  assign \new_[25389]_  = A168 & \new_[25388]_ ;
  assign \new_[25393]_  = ~A232 & ~A202;
  assign \new_[25394]_  = ~A200 & \new_[25393]_ ;
  assign \new_[25395]_  = \new_[25394]_  & \new_[25389]_ ;
  assign \new_[25399]_  = ~A267 & ~A235;
  assign \new_[25400]_  = ~A233 & \new_[25399]_ ;
  assign \new_[25404]_  = A301 & ~A269;
  assign \new_[25405]_  = ~A268 & \new_[25404]_ ;
  assign \new_[25406]_  = \new_[25405]_  & \new_[25400]_ ;
  assign \new_[25410]_  = ~A199 & A167;
  assign \new_[25411]_  = A168 & \new_[25410]_ ;
  assign \new_[25415]_  = ~A232 & ~A202;
  assign \new_[25416]_  = ~A200 & \new_[25415]_ ;
  assign \new_[25417]_  = \new_[25416]_  & \new_[25411]_ ;
  assign \new_[25421]_  = ~A265 & ~A235;
  assign \new_[25422]_  = ~A233 & \new_[25421]_ ;
  assign \new_[25426]_  = A301 & ~A268;
  assign \new_[25427]_  = ~A266 & \new_[25426]_ ;
  assign \new_[25428]_  = \new_[25427]_  & \new_[25422]_ ;
  assign \new_[25432]_  = ~A166 & A167;
  assign \new_[25433]_  = A170 & \new_[25432]_ ;
  assign \new_[25437]_  = ~A203 & ~A202;
  assign \new_[25438]_  = ~A201 & \new_[25437]_ ;
  assign \new_[25439]_  = \new_[25438]_  & \new_[25433]_ ;
  assign \new_[25443]_  = A298 & A234;
  assign \new_[25444]_  = A232 & \new_[25443]_ ;
  assign \new_[25448]_  = ~A301 & ~A300;
  assign \new_[25449]_  = A299 & \new_[25448]_ ;
  assign \new_[25450]_  = \new_[25449]_  & \new_[25444]_ ;
  assign \new_[25454]_  = ~A166 & A167;
  assign \new_[25455]_  = A170 & \new_[25454]_ ;
  assign \new_[25459]_  = ~A203 & ~A202;
  assign \new_[25460]_  = ~A201 & \new_[25459]_ ;
  assign \new_[25461]_  = \new_[25460]_  & \new_[25455]_ ;
  assign \new_[25465]_  = A298 & A234;
  assign \new_[25466]_  = A233 & \new_[25465]_ ;
  assign \new_[25470]_  = ~A301 & ~A300;
  assign \new_[25471]_  = A299 & \new_[25470]_ ;
  assign \new_[25472]_  = \new_[25471]_  & \new_[25466]_ ;
  assign \new_[25476]_  = ~A166 & A167;
  assign \new_[25477]_  = A170 & \new_[25476]_ ;
  assign \new_[25481]_  = ~A203 & ~A202;
  assign \new_[25482]_  = ~A201 & \new_[25481]_ ;
  assign \new_[25483]_  = \new_[25482]_  & \new_[25477]_ ;
  assign \new_[25487]_  = A236 & A233;
  assign \new_[25488]_  = ~A232 & \new_[25487]_ ;
  assign \new_[25492]_  = ~A302 & ~A301;
  assign \new_[25493]_  = ~A300 & \new_[25492]_ ;
  assign \new_[25494]_  = \new_[25493]_  & \new_[25488]_ ;
  assign \new_[25498]_  = ~A166 & A167;
  assign \new_[25499]_  = A170 & \new_[25498]_ ;
  assign \new_[25503]_  = ~A203 & ~A202;
  assign \new_[25504]_  = ~A201 & \new_[25503]_ ;
  assign \new_[25505]_  = \new_[25504]_  & \new_[25499]_ ;
  assign \new_[25509]_  = A236 & A233;
  assign \new_[25510]_  = ~A232 & \new_[25509]_ ;
  assign \new_[25514]_  = ~A301 & ~A299;
  assign \new_[25515]_  = ~A298 & \new_[25514]_ ;
  assign \new_[25516]_  = \new_[25515]_  & \new_[25510]_ ;
  assign \new_[25520]_  = ~A166 & A167;
  assign \new_[25521]_  = A170 & \new_[25520]_ ;
  assign \new_[25525]_  = ~A203 & ~A202;
  assign \new_[25526]_  = ~A201 & \new_[25525]_ ;
  assign \new_[25527]_  = \new_[25526]_  & \new_[25521]_ ;
  assign \new_[25531]_  = A236 & A233;
  assign \new_[25532]_  = ~A232 & \new_[25531]_ ;
  assign \new_[25536]_  = A269 & A266;
  assign \new_[25537]_  = ~A265 & \new_[25536]_ ;
  assign \new_[25538]_  = \new_[25537]_  & \new_[25532]_ ;
  assign \new_[25542]_  = ~A166 & A167;
  assign \new_[25543]_  = A170 & \new_[25542]_ ;
  assign \new_[25547]_  = ~A203 & ~A202;
  assign \new_[25548]_  = ~A201 & \new_[25547]_ ;
  assign \new_[25549]_  = \new_[25548]_  & \new_[25543]_ ;
  assign \new_[25553]_  = A236 & A233;
  assign \new_[25554]_  = ~A232 & \new_[25553]_ ;
  assign \new_[25558]_  = A269 & ~A266;
  assign \new_[25559]_  = A265 & \new_[25558]_ ;
  assign \new_[25560]_  = \new_[25559]_  & \new_[25554]_ ;
  assign \new_[25564]_  = ~A166 & A167;
  assign \new_[25565]_  = A170 & \new_[25564]_ ;
  assign \new_[25569]_  = ~A203 & ~A202;
  assign \new_[25570]_  = ~A201 & \new_[25569]_ ;
  assign \new_[25571]_  = \new_[25570]_  & \new_[25565]_ ;
  assign \new_[25575]_  = A236 & ~A233;
  assign \new_[25576]_  = A232 & \new_[25575]_ ;
  assign \new_[25580]_  = ~A302 & ~A301;
  assign \new_[25581]_  = ~A300 & \new_[25580]_ ;
  assign \new_[25582]_  = \new_[25581]_  & \new_[25576]_ ;
  assign \new_[25586]_  = ~A166 & A167;
  assign \new_[25587]_  = A170 & \new_[25586]_ ;
  assign \new_[25591]_  = ~A203 & ~A202;
  assign \new_[25592]_  = ~A201 & \new_[25591]_ ;
  assign \new_[25593]_  = \new_[25592]_  & \new_[25587]_ ;
  assign \new_[25597]_  = A236 & ~A233;
  assign \new_[25598]_  = A232 & \new_[25597]_ ;
  assign \new_[25602]_  = ~A301 & ~A299;
  assign \new_[25603]_  = ~A298 & \new_[25602]_ ;
  assign \new_[25604]_  = \new_[25603]_  & \new_[25598]_ ;
  assign \new_[25608]_  = ~A166 & A167;
  assign \new_[25609]_  = A170 & \new_[25608]_ ;
  assign \new_[25613]_  = ~A203 & ~A202;
  assign \new_[25614]_  = ~A201 & \new_[25613]_ ;
  assign \new_[25615]_  = \new_[25614]_  & \new_[25609]_ ;
  assign \new_[25619]_  = A236 & ~A233;
  assign \new_[25620]_  = A232 & \new_[25619]_ ;
  assign \new_[25624]_  = A269 & A266;
  assign \new_[25625]_  = ~A265 & \new_[25624]_ ;
  assign \new_[25626]_  = \new_[25625]_  & \new_[25620]_ ;
  assign \new_[25630]_  = ~A166 & A167;
  assign \new_[25631]_  = A170 & \new_[25630]_ ;
  assign \new_[25635]_  = ~A203 & ~A202;
  assign \new_[25636]_  = ~A201 & \new_[25635]_ ;
  assign \new_[25637]_  = \new_[25636]_  & \new_[25631]_ ;
  assign \new_[25641]_  = A236 & ~A233;
  assign \new_[25642]_  = A232 & \new_[25641]_ ;
  assign \new_[25646]_  = A269 & ~A266;
  assign \new_[25647]_  = A265 & \new_[25646]_ ;
  assign \new_[25648]_  = \new_[25647]_  & \new_[25642]_ ;
  assign \new_[25652]_  = ~A166 & A167;
  assign \new_[25653]_  = A170 & \new_[25652]_ ;
  assign \new_[25657]_  = ~A201 & A200;
  assign \new_[25658]_  = A199 & \new_[25657]_ ;
  assign \new_[25659]_  = \new_[25658]_  & \new_[25653]_ ;
  assign \new_[25663]_  = A298 & A235;
  assign \new_[25664]_  = ~A202 & \new_[25663]_ ;
  assign \new_[25668]_  = ~A301 & ~A300;
  assign \new_[25669]_  = A299 & \new_[25668]_ ;
  assign \new_[25670]_  = \new_[25669]_  & \new_[25664]_ ;
  assign \new_[25674]_  = ~A166 & A167;
  assign \new_[25675]_  = A170 & \new_[25674]_ ;
  assign \new_[25679]_  = ~A201 & A200;
  assign \new_[25680]_  = A199 & \new_[25679]_ ;
  assign \new_[25681]_  = \new_[25680]_  & \new_[25675]_ ;
  assign \new_[25685]_  = A234 & A232;
  assign \new_[25686]_  = ~A202 & \new_[25685]_ ;
  assign \new_[25690]_  = ~A302 & ~A301;
  assign \new_[25691]_  = ~A300 & \new_[25690]_ ;
  assign \new_[25692]_  = \new_[25691]_  & \new_[25686]_ ;
  assign \new_[25696]_  = ~A166 & A167;
  assign \new_[25697]_  = A170 & \new_[25696]_ ;
  assign \new_[25701]_  = ~A201 & A200;
  assign \new_[25702]_  = A199 & \new_[25701]_ ;
  assign \new_[25703]_  = \new_[25702]_  & \new_[25697]_ ;
  assign \new_[25707]_  = A234 & A232;
  assign \new_[25708]_  = ~A202 & \new_[25707]_ ;
  assign \new_[25712]_  = ~A301 & ~A299;
  assign \new_[25713]_  = ~A298 & \new_[25712]_ ;
  assign \new_[25714]_  = \new_[25713]_  & \new_[25708]_ ;
  assign \new_[25718]_  = ~A166 & A167;
  assign \new_[25719]_  = A170 & \new_[25718]_ ;
  assign \new_[25723]_  = ~A201 & A200;
  assign \new_[25724]_  = A199 & \new_[25723]_ ;
  assign \new_[25725]_  = \new_[25724]_  & \new_[25719]_ ;
  assign \new_[25729]_  = A234 & A232;
  assign \new_[25730]_  = ~A202 & \new_[25729]_ ;
  assign \new_[25734]_  = A269 & A266;
  assign \new_[25735]_  = ~A265 & \new_[25734]_ ;
  assign \new_[25736]_  = \new_[25735]_  & \new_[25730]_ ;
  assign \new_[25740]_  = ~A166 & A167;
  assign \new_[25741]_  = A170 & \new_[25740]_ ;
  assign \new_[25745]_  = ~A201 & A200;
  assign \new_[25746]_  = A199 & \new_[25745]_ ;
  assign \new_[25747]_  = \new_[25746]_  & \new_[25741]_ ;
  assign \new_[25751]_  = A234 & A232;
  assign \new_[25752]_  = ~A202 & \new_[25751]_ ;
  assign \new_[25756]_  = A269 & ~A266;
  assign \new_[25757]_  = A265 & \new_[25756]_ ;
  assign \new_[25758]_  = \new_[25757]_  & \new_[25752]_ ;
  assign \new_[25762]_  = ~A166 & A167;
  assign \new_[25763]_  = A170 & \new_[25762]_ ;
  assign \new_[25767]_  = ~A201 & A200;
  assign \new_[25768]_  = A199 & \new_[25767]_ ;
  assign \new_[25769]_  = \new_[25768]_  & \new_[25763]_ ;
  assign \new_[25773]_  = A234 & A233;
  assign \new_[25774]_  = ~A202 & \new_[25773]_ ;
  assign \new_[25778]_  = ~A302 & ~A301;
  assign \new_[25779]_  = ~A300 & \new_[25778]_ ;
  assign \new_[25780]_  = \new_[25779]_  & \new_[25774]_ ;
  assign \new_[25784]_  = ~A166 & A167;
  assign \new_[25785]_  = A170 & \new_[25784]_ ;
  assign \new_[25789]_  = ~A201 & A200;
  assign \new_[25790]_  = A199 & \new_[25789]_ ;
  assign \new_[25791]_  = \new_[25790]_  & \new_[25785]_ ;
  assign \new_[25795]_  = A234 & A233;
  assign \new_[25796]_  = ~A202 & \new_[25795]_ ;
  assign \new_[25800]_  = ~A301 & ~A299;
  assign \new_[25801]_  = ~A298 & \new_[25800]_ ;
  assign \new_[25802]_  = \new_[25801]_  & \new_[25796]_ ;
  assign \new_[25806]_  = ~A166 & A167;
  assign \new_[25807]_  = A170 & \new_[25806]_ ;
  assign \new_[25811]_  = ~A201 & A200;
  assign \new_[25812]_  = A199 & \new_[25811]_ ;
  assign \new_[25813]_  = \new_[25812]_  & \new_[25807]_ ;
  assign \new_[25817]_  = A234 & A233;
  assign \new_[25818]_  = ~A202 & \new_[25817]_ ;
  assign \new_[25822]_  = A269 & A266;
  assign \new_[25823]_  = ~A265 & \new_[25822]_ ;
  assign \new_[25824]_  = \new_[25823]_  & \new_[25818]_ ;
  assign \new_[25828]_  = ~A166 & A167;
  assign \new_[25829]_  = A170 & \new_[25828]_ ;
  assign \new_[25833]_  = ~A201 & A200;
  assign \new_[25834]_  = A199 & \new_[25833]_ ;
  assign \new_[25835]_  = \new_[25834]_  & \new_[25829]_ ;
  assign \new_[25839]_  = A234 & A233;
  assign \new_[25840]_  = ~A202 & \new_[25839]_ ;
  assign \new_[25844]_  = A269 & ~A266;
  assign \new_[25845]_  = A265 & \new_[25844]_ ;
  assign \new_[25846]_  = \new_[25845]_  & \new_[25840]_ ;
  assign \new_[25850]_  = ~A166 & A167;
  assign \new_[25851]_  = A170 & \new_[25850]_ ;
  assign \new_[25855]_  = ~A201 & A200;
  assign \new_[25856]_  = A199 & \new_[25855]_ ;
  assign \new_[25857]_  = \new_[25856]_  & \new_[25851]_ ;
  assign \new_[25861]_  = A233 & ~A232;
  assign \new_[25862]_  = ~A202 & \new_[25861]_ ;
  assign \new_[25866]_  = A267 & A265;
  assign \new_[25867]_  = A236 & \new_[25866]_ ;
  assign \new_[25868]_  = \new_[25867]_  & \new_[25862]_ ;
  assign \new_[25872]_  = ~A166 & A167;
  assign \new_[25873]_  = A170 & \new_[25872]_ ;
  assign \new_[25877]_  = ~A201 & A200;
  assign \new_[25878]_  = A199 & \new_[25877]_ ;
  assign \new_[25879]_  = \new_[25878]_  & \new_[25873]_ ;
  assign \new_[25883]_  = A233 & ~A232;
  assign \new_[25884]_  = ~A202 & \new_[25883]_ ;
  assign \new_[25888]_  = A267 & A266;
  assign \new_[25889]_  = A236 & \new_[25888]_ ;
  assign \new_[25890]_  = \new_[25889]_  & \new_[25884]_ ;
  assign \new_[25894]_  = ~A166 & A167;
  assign \new_[25895]_  = A170 & \new_[25894]_ ;
  assign \new_[25899]_  = ~A201 & A200;
  assign \new_[25900]_  = A199 & \new_[25899]_ ;
  assign \new_[25901]_  = \new_[25900]_  & \new_[25895]_ ;
  assign \new_[25905]_  = ~A233 & A232;
  assign \new_[25906]_  = ~A202 & \new_[25905]_ ;
  assign \new_[25910]_  = A267 & A265;
  assign \new_[25911]_  = A236 & \new_[25910]_ ;
  assign \new_[25912]_  = \new_[25911]_  & \new_[25906]_ ;
  assign \new_[25916]_  = ~A166 & A167;
  assign \new_[25917]_  = A170 & \new_[25916]_ ;
  assign \new_[25921]_  = ~A201 & A200;
  assign \new_[25922]_  = A199 & \new_[25921]_ ;
  assign \new_[25923]_  = \new_[25922]_  & \new_[25917]_ ;
  assign \new_[25927]_  = ~A233 & A232;
  assign \new_[25928]_  = ~A202 & \new_[25927]_ ;
  assign \new_[25932]_  = A267 & A266;
  assign \new_[25933]_  = A236 & \new_[25932]_ ;
  assign \new_[25934]_  = \new_[25933]_  & \new_[25928]_ ;
  assign \new_[25938]_  = ~A166 & A167;
  assign \new_[25939]_  = A170 & \new_[25938]_ ;
  assign \new_[25943]_  = ~A202 & ~A200;
  assign \new_[25944]_  = ~A199 & \new_[25943]_ ;
  assign \new_[25945]_  = \new_[25944]_  & \new_[25939]_ ;
  assign \new_[25949]_  = A298 & A234;
  assign \new_[25950]_  = A232 & \new_[25949]_ ;
  assign \new_[25954]_  = ~A301 & ~A300;
  assign \new_[25955]_  = A299 & \new_[25954]_ ;
  assign \new_[25956]_  = \new_[25955]_  & \new_[25950]_ ;
  assign \new_[25960]_  = ~A166 & A167;
  assign \new_[25961]_  = A170 & \new_[25960]_ ;
  assign \new_[25965]_  = ~A202 & ~A200;
  assign \new_[25966]_  = ~A199 & \new_[25965]_ ;
  assign \new_[25967]_  = \new_[25966]_  & \new_[25961]_ ;
  assign \new_[25971]_  = A298 & A234;
  assign \new_[25972]_  = A233 & \new_[25971]_ ;
  assign \new_[25976]_  = ~A301 & ~A300;
  assign \new_[25977]_  = A299 & \new_[25976]_ ;
  assign \new_[25978]_  = \new_[25977]_  & \new_[25972]_ ;
  assign \new_[25982]_  = ~A166 & A167;
  assign \new_[25983]_  = A170 & \new_[25982]_ ;
  assign \new_[25987]_  = ~A202 & ~A200;
  assign \new_[25988]_  = ~A199 & \new_[25987]_ ;
  assign \new_[25989]_  = \new_[25988]_  & \new_[25983]_ ;
  assign \new_[25993]_  = A236 & A233;
  assign \new_[25994]_  = ~A232 & \new_[25993]_ ;
  assign \new_[25998]_  = ~A302 & ~A301;
  assign \new_[25999]_  = ~A300 & \new_[25998]_ ;
  assign \new_[26000]_  = \new_[25999]_  & \new_[25994]_ ;
  assign \new_[26004]_  = ~A166 & A167;
  assign \new_[26005]_  = A170 & \new_[26004]_ ;
  assign \new_[26009]_  = ~A202 & ~A200;
  assign \new_[26010]_  = ~A199 & \new_[26009]_ ;
  assign \new_[26011]_  = \new_[26010]_  & \new_[26005]_ ;
  assign \new_[26015]_  = A236 & A233;
  assign \new_[26016]_  = ~A232 & \new_[26015]_ ;
  assign \new_[26020]_  = ~A301 & ~A299;
  assign \new_[26021]_  = ~A298 & \new_[26020]_ ;
  assign \new_[26022]_  = \new_[26021]_  & \new_[26016]_ ;
  assign \new_[26026]_  = ~A166 & A167;
  assign \new_[26027]_  = A170 & \new_[26026]_ ;
  assign \new_[26031]_  = ~A202 & ~A200;
  assign \new_[26032]_  = ~A199 & \new_[26031]_ ;
  assign \new_[26033]_  = \new_[26032]_  & \new_[26027]_ ;
  assign \new_[26037]_  = A236 & A233;
  assign \new_[26038]_  = ~A232 & \new_[26037]_ ;
  assign \new_[26042]_  = A269 & A266;
  assign \new_[26043]_  = ~A265 & \new_[26042]_ ;
  assign \new_[26044]_  = \new_[26043]_  & \new_[26038]_ ;
  assign \new_[26048]_  = ~A166 & A167;
  assign \new_[26049]_  = A170 & \new_[26048]_ ;
  assign \new_[26053]_  = ~A202 & ~A200;
  assign \new_[26054]_  = ~A199 & \new_[26053]_ ;
  assign \new_[26055]_  = \new_[26054]_  & \new_[26049]_ ;
  assign \new_[26059]_  = A236 & A233;
  assign \new_[26060]_  = ~A232 & \new_[26059]_ ;
  assign \new_[26064]_  = A269 & ~A266;
  assign \new_[26065]_  = A265 & \new_[26064]_ ;
  assign \new_[26066]_  = \new_[26065]_  & \new_[26060]_ ;
  assign \new_[26070]_  = ~A166 & A167;
  assign \new_[26071]_  = A170 & \new_[26070]_ ;
  assign \new_[26075]_  = ~A202 & ~A200;
  assign \new_[26076]_  = ~A199 & \new_[26075]_ ;
  assign \new_[26077]_  = \new_[26076]_  & \new_[26071]_ ;
  assign \new_[26081]_  = A236 & ~A233;
  assign \new_[26082]_  = A232 & \new_[26081]_ ;
  assign \new_[26086]_  = ~A302 & ~A301;
  assign \new_[26087]_  = ~A300 & \new_[26086]_ ;
  assign \new_[26088]_  = \new_[26087]_  & \new_[26082]_ ;
  assign \new_[26092]_  = ~A166 & A167;
  assign \new_[26093]_  = A170 & \new_[26092]_ ;
  assign \new_[26097]_  = ~A202 & ~A200;
  assign \new_[26098]_  = ~A199 & \new_[26097]_ ;
  assign \new_[26099]_  = \new_[26098]_  & \new_[26093]_ ;
  assign \new_[26103]_  = A236 & ~A233;
  assign \new_[26104]_  = A232 & \new_[26103]_ ;
  assign \new_[26108]_  = ~A301 & ~A299;
  assign \new_[26109]_  = ~A298 & \new_[26108]_ ;
  assign \new_[26110]_  = \new_[26109]_  & \new_[26104]_ ;
  assign \new_[26114]_  = ~A166 & A167;
  assign \new_[26115]_  = A170 & \new_[26114]_ ;
  assign \new_[26119]_  = ~A202 & ~A200;
  assign \new_[26120]_  = ~A199 & \new_[26119]_ ;
  assign \new_[26121]_  = \new_[26120]_  & \new_[26115]_ ;
  assign \new_[26125]_  = A236 & ~A233;
  assign \new_[26126]_  = A232 & \new_[26125]_ ;
  assign \new_[26130]_  = A269 & A266;
  assign \new_[26131]_  = ~A265 & \new_[26130]_ ;
  assign \new_[26132]_  = \new_[26131]_  & \new_[26126]_ ;
  assign \new_[26136]_  = ~A166 & A167;
  assign \new_[26137]_  = A170 & \new_[26136]_ ;
  assign \new_[26141]_  = ~A202 & ~A200;
  assign \new_[26142]_  = ~A199 & \new_[26141]_ ;
  assign \new_[26143]_  = \new_[26142]_  & \new_[26137]_ ;
  assign \new_[26147]_  = A236 & ~A233;
  assign \new_[26148]_  = A232 & \new_[26147]_ ;
  assign \new_[26152]_  = A269 & ~A266;
  assign \new_[26153]_  = A265 & \new_[26152]_ ;
  assign \new_[26154]_  = \new_[26153]_  & \new_[26148]_ ;
  assign \new_[26158]_  = A166 & ~A167;
  assign \new_[26159]_  = A170 & \new_[26158]_ ;
  assign \new_[26163]_  = ~A203 & ~A202;
  assign \new_[26164]_  = ~A201 & \new_[26163]_ ;
  assign \new_[26165]_  = \new_[26164]_  & \new_[26159]_ ;
  assign \new_[26169]_  = A298 & A234;
  assign \new_[26170]_  = A232 & \new_[26169]_ ;
  assign \new_[26174]_  = ~A301 & ~A300;
  assign \new_[26175]_  = A299 & \new_[26174]_ ;
  assign \new_[26176]_  = \new_[26175]_  & \new_[26170]_ ;
  assign \new_[26180]_  = A166 & ~A167;
  assign \new_[26181]_  = A170 & \new_[26180]_ ;
  assign \new_[26185]_  = ~A203 & ~A202;
  assign \new_[26186]_  = ~A201 & \new_[26185]_ ;
  assign \new_[26187]_  = \new_[26186]_  & \new_[26181]_ ;
  assign \new_[26191]_  = A298 & A234;
  assign \new_[26192]_  = A233 & \new_[26191]_ ;
  assign \new_[26196]_  = ~A301 & ~A300;
  assign \new_[26197]_  = A299 & \new_[26196]_ ;
  assign \new_[26198]_  = \new_[26197]_  & \new_[26192]_ ;
  assign \new_[26202]_  = A166 & ~A167;
  assign \new_[26203]_  = A170 & \new_[26202]_ ;
  assign \new_[26207]_  = ~A203 & ~A202;
  assign \new_[26208]_  = ~A201 & \new_[26207]_ ;
  assign \new_[26209]_  = \new_[26208]_  & \new_[26203]_ ;
  assign \new_[26213]_  = A236 & A233;
  assign \new_[26214]_  = ~A232 & \new_[26213]_ ;
  assign \new_[26218]_  = ~A302 & ~A301;
  assign \new_[26219]_  = ~A300 & \new_[26218]_ ;
  assign \new_[26220]_  = \new_[26219]_  & \new_[26214]_ ;
  assign \new_[26224]_  = A166 & ~A167;
  assign \new_[26225]_  = A170 & \new_[26224]_ ;
  assign \new_[26229]_  = ~A203 & ~A202;
  assign \new_[26230]_  = ~A201 & \new_[26229]_ ;
  assign \new_[26231]_  = \new_[26230]_  & \new_[26225]_ ;
  assign \new_[26235]_  = A236 & A233;
  assign \new_[26236]_  = ~A232 & \new_[26235]_ ;
  assign \new_[26240]_  = ~A301 & ~A299;
  assign \new_[26241]_  = ~A298 & \new_[26240]_ ;
  assign \new_[26242]_  = \new_[26241]_  & \new_[26236]_ ;
  assign \new_[26246]_  = A166 & ~A167;
  assign \new_[26247]_  = A170 & \new_[26246]_ ;
  assign \new_[26251]_  = ~A203 & ~A202;
  assign \new_[26252]_  = ~A201 & \new_[26251]_ ;
  assign \new_[26253]_  = \new_[26252]_  & \new_[26247]_ ;
  assign \new_[26257]_  = A236 & A233;
  assign \new_[26258]_  = ~A232 & \new_[26257]_ ;
  assign \new_[26262]_  = A269 & A266;
  assign \new_[26263]_  = ~A265 & \new_[26262]_ ;
  assign \new_[26264]_  = \new_[26263]_  & \new_[26258]_ ;
  assign \new_[26268]_  = A166 & ~A167;
  assign \new_[26269]_  = A170 & \new_[26268]_ ;
  assign \new_[26273]_  = ~A203 & ~A202;
  assign \new_[26274]_  = ~A201 & \new_[26273]_ ;
  assign \new_[26275]_  = \new_[26274]_  & \new_[26269]_ ;
  assign \new_[26279]_  = A236 & A233;
  assign \new_[26280]_  = ~A232 & \new_[26279]_ ;
  assign \new_[26284]_  = A269 & ~A266;
  assign \new_[26285]_  = A265 & \new_[26284]_ ;
  assign \new_[26286]_  = \new_[26285]_  & \new_[26280]_ ;
  assign \new_[26290]_  = A166 & ~A167;
  assign \new_[26291]_  = A170 & \new_[26290]_ ;
  assign \new_[26295]_  = ~A203 & ~A202;
  assign \new_[26296]_  = ~A201 & \new_[26295]_ ;
  assign \new_[26297]_  = \new_[26296]_  & \new_[26291]_ ;
  assign \new_[26301]_  = A236 & ~A233;
  assign \new_[26302]_  = A232 & \new_[26301]_ ;
  assign \new_[26306]_  = ~A302 & ~A301;
  assign \new_[26307]_  = ~A300 & \new_[26306]_ ;
  assign \new_[26308]_  = \new_[26307]_  & \new_[26302]_ ;
  assign \new_[26312]_  = A166 & ~A167;
  assign \new_[26313]_  = A170 & \new_[26312]_ ;
  assign \new_[26317]_  = ~A203 & ~A202;
  assign \new_[26318]_  = ~A201 & \new_[26317]_ ;
  assign \new_[26319]_  = \new_[26318]_  & \new_[26313]_ ;
  assign \new_[26323]_  = A236 & ~A233;
  assign \new_[26324]_  = A232 & \new_[26323]_ ;
  assign \new_[26328]_  = ~A301 & ~A299;
  assign \new_[26329]_  = ~A298 & \new_[26328]_ ;
  assign \new_[26330]_  = \new_[26329]_  & \new_[26324]_ ;
  assign \new_[26334]_  = A166 & ~A167;
  assign \new_[26335]_  = A170 & \new_[26334]_ ;
  assign \new_[26339]_  = ~A203 & ~A202;
  assign \new_[26340]_  = ~A201 & \new_[26339]_ ;
  assign \new_[26341]_  = \new_[26340]_  & \new_[26335]_ ;
  assign \new_[26345]_  = A236 & ~A233;
  assign \new_[26346]_  = A232 & \new_[26345]_ ;
  assign \new_[26350]_  = A269 & A266;
  assign \new_[26351]_  = ~A265 & \new_[26350]_ ;
  assign \new_[26352]_  = \new_[26351]_  & \new_[26346]_ ;
  assign \new_[26356]_  = A166 & ~A167;
  assign \new_[26357]_  = A170 & \new_[26356]_ ;
  assign \new_[26361]_  = ~A203 & ~A202;
  assign \new_[26362]_  = ~A201 & \new_[26361]_ ;
  assign \new_[26363]_  = \new_[26362]_  & \new_[26357]_ ;
  assign \new_[26367]_  = A236 & ~A233;
  assign \new_[26368]_  = A232 & \new_[26367]_ ;
  assign \new_[26372]_  = A269 & ~A266;
  assign \new_[26373]_  = A265 & \new_[26372]_ ;
  assign \new_[26374]_  = \new_[26373]_  & \new_[26368]_ ;
  assign \new_[26378]_  = A166 & ~A167;
  assign \new_[26379]_  = A170 & \new_[26378]_ ;
  assign \new_[26383]_  = ~A201 & A200;
  assign \new_[26384]_  = A199 & \new_[26383]_ ;
  assign \new_[26385]_  = \new_[26384]_  & \new_[26379]_ ;
  assign \new_[26389]_  = A298 & A235;
  assign \new_[26390]_  = ~A202 & \new_[26389]_ ;
  assign \new_[26394]_  = ~A301 & ~A300;
  assign \new_[26395]_  = A299 & \new_[26394]_ ;
  assign \new_[26396]_  = \new_[26395]_  & \new_[26390]_ ;
  assign \new_[26400]_  = A166 & ~A167;
  assign \new_[26401]_  = A170 & \new_[26400]_ ;
  assign \new_[26405]_  = ~A201 & A200;
  assign \new_[26406]_  = A199 & \new_[26405]_ ;
  assign \new_[26407]_  = \new_[26406]_  & \new_[26401]_ ;
  assign \new_[26411]_  = A234 & A232;
  assign \new_[26412]_  = ~A202 & \new_[26411]_ ;
  assign \new_[26416]_  = ~A302 & ~A301;
  assign \new_[26417]_  = ~A300 & \new_[26416]_ ;
  assign \new_[26418]_  = \new_[26417]_  & \new_[26412]_ ;
  assign \new_[26422]_  = A166 & ~A167;
  assign \new_[26423]_  = A170 & \new_[26422]_ ;
  assign \new_[26427]_  = ~A201 & A200;
  assign \new_[26428]_  = A199 & \new_[26427]_ ;
  assign \new_[26429]_  = \new_[26428]_  & \new_[26423]_ ;
  assign \new_[26433]_  = A234 & A232;
  assign \new_[26434]_  = ~A202 & \new_[26433]_ ;
  assign \new_[26438]_  = ~A301 & ~A299;
  assign \new_[26439]_  = ~A298 & \new_[26438]_ ;
  assign \new_[26440]_  = \new_[26439]_  & \new_[26434]_ ;
  assign \new_[26444]_  = A166 & ~A167;
  assign \new_[26445]_  = A170 & \new_[26444]_ ;
  assign \new_[26449]_  = ~A201 & A200;
  assign \new_[26450]_  = A199 & \new_[26449]_ ;
  assign \new_[26451]_  = \new_[26450]_  & \new_[26445]_ ;
  assign \new_[26455]_  = A234 & A232;
  assign \new_[26456]_  = ~A202 & \new_[26455]_ ;
  assign \new_[26460]_  = A269 & A266;
  assign \new_[26461]_  = ~A265 & \new_[26460]_ ;
  assign \new_[26462]_  = \new_[26461]_  & \new_[26456]_ ;
  assign \new_[26466]_  = A166 & ~A167;
  assign \new_[26467]_  = A170 & \new_[26466]_ ;
  assign \new_[26471]_  = ~A201 & A200;
  assign \new_[26472]_  = A199 & \new_[26471]_ ;
  assign \new_[26473]_  = \new_[26472]_  & \new_[26467]_ ;
  assign \new_[26477]_  = A234 & A232;
  assign \new_[26478]_  = ~A202 & \new_[26477]_ ;
  assign \new_[26482]_  = A269 & ~A266;
  assign \new_[26483]_  = A265 & \new_[26482]_ ;
  assign \new_[26484]_  = \new_[26483]_  & \new_[26478]_ ;
  assign \new_[26488]_  = A166 & ~A167;
  assign \new_[26489]_  = A170 & \new_[26488]_ ;
  assign \new_[26493]_  = ~A201 & A200;
  assign \new_[26494]_  = A199 & \new_[26493]_ ;
  assign \new_[26495]_  = \new_[26494]_  & \new_[26489]_ ;
  assign \new_[26499]_  = A234 & A233;
  assign \new_[26500]_  = ~A202 & \new_[26499]_ ;
  assign \new_[26504]_  = ~A302 & ~A301;
  assign \new_[26505]_  = ~A300 & \new_[26504]_ ;
  assign \new_[26506]_  = \new_[26505]_  & \new_[26500]_ ;
  assign \new_[26510]_  = A166 & ~A167;
  assign \new_[26511]_  = A170 & \new_[26510]_ ;
  assign \new_[26515]_  = ~A201 & A200;
  assign \new_[26516]_  = A199 & \new_[26515]_ ;
  assign \new_[26517]_  = \new_[26516]_  & \new_[26511]_ ;
  assign \new_[26521]_  = A234 & A233;
  assign \new_[26522]_  = ~A202 & \new_[26521]_ ;
  assign \new_[26526]_  = ~A301 & ~A299;
  assign \new_[26527]_  = ~A298 & \new_[26526]_ ;
  assign \new_[26528]_  = \new_[26527]_  & \new_[26522]_ ;
  assign \new_[26532]_  = A166 & ~A167;
  assign \new_[26533]_  = A170 & \new_[26532]_ ;
  assign \new_[26537]_  = ~A201 & A200;
  assign \new_[26538]_  = A199 & \new_[26537]_ ;
  assign \new_[26539]_  = \new_[26538]_  & \new_[26533]_ ;
  assign \new_[26543]_  = A234 & A233;
  assign \new_[26544]_  = ~A202 & \new_[26543]_ ;
  assign \new_[26548]_  = A269 & A266;
  assign \new_[26549]_  = ~A265 & \new_[26548]_ ;
  assign \new_[26550]_  = \new_[26549]_  & \new_[26544]_ ;
  assign \new_[26554]_  = A166 & ~A167;
  assign \new_[26555]_  = A170 & \new_[26554]_ ;
  assign \new_[26559]_  = ~A201 & A200;
  assign \new_[26560]_  = A199 & \new_[26559]_ ;
  assign \new_[26561]_  = \new_[26560]_  & \new_[26555]_ ;
  assign \new_[26565]_  = A234 & A233;
  assign \new_[26566]_  = ~A202 & \new_[26565]_ ;
  assign \new_[26570]_  = A269 & ~A266;
  assign \new_[26571]_  = A265 & \new_[26570]_ ;
  assign \new_[26572]_  = \new_[26571]_  & \new_[26566]_ ;
  assign \new_[26576]_  = A166 & ~A167;
  assign \new_[26577]_  = A170 & \new_[26576]_ ;
  assign \new_[26581]_  = ~A201 & A200;
  assign \new_[26582]_  = A199 & \new_[26581]_ ;
  assign \new_[26583]_  = \new_[26582]_  & \new_[26577]_ ;
  assign \new_[26587]_  = A233 & ~A232;
  assign \new_[26588]_  = ~A202 & \new_[26587]_ ;
  assign \new_[26592]_  = A267 & A265;
  assign \new_[26593]_  = A236 & \new_[26592]_ ;
  assign \new_[26594]_  = \new_[26593]_  & \new_[26588]_ ;
  assign \new_[26598]_  = A166 & ~A167;
  assign \new_[26599]_  = A170 & \new_[26598]_ ;
  assign \new_[26603]_  = ~A201 & A200;
  assign \new_[26604]_  = A199 & \new_[26603]_ ;
  assign \new_[26605]_  = \new_[26604]_  & \new_[26599]_ ;
  assign \new_[26609]_  = A233 & ~A232;
  assign \new_[26610]_  = ~A202 & \new_[26609]_ ;
  assign \new_[26614]_  = A267 & A266;
  assign \new_[26615]_  = A236 & \new_[26614]_ ;
  assign \new_[26616]_  = \new_[26615]_  & \new_[26610]_ ;
  assign \new_[26620]_  = A166 & ~A167;
  assign \new_[26621]_  = A170 & \new_[26620]_ ;
  assign \new_[26625]_  = ~A201 & A200;
  assign \new_[26626]_  = A199 & \new_[26625]_ ;
  assign \new_[26627]_  = \new_[26626]_  & \new_[26621]_ ;
  assign \new_[26631]_  = ~A233 & A232;
  assign \new_[26632]_  = ~A202 & \new_[26631]_ ;
  assign \new_[26636]_  = A267 & A265;
  assign \new_[26637]_  = A236 & \new_[26636]_ ;
  assign \new_[26638]_  = \new_[26637]_  & \new_[26632]_ ;
  assign \new_[26642]_  = A166 & ~A167;
  assign \new_[26643]_  = A170 & \new_[26642]_ ;
  assign \new_[26647]_  = ~A201 & A200;
  assign \new_[26648]_  = A199 & \new_[26647]_ ;
  assign \new_[26649]_  = \new_[26648]_  & \new_[26643]_ ;
  assign \new_[26653]_  = ~A233 & A232;
  assign \new_[26654]_  = ~A202 & \new_[26653]_ ;
  assign \new_[26658]_  = A267 & A266;
  assign \new_[26659]_  = A236 & \new_[26658]_ ;
  assign \new_[26660]_  = \new_[26659]_  & \new_[26654]_ ;
  assign \new_[26664]_  = A166 & ~A167;
  assign \new_[26665]_  = A170 & \new_[26664]_ ;
  assign \new_[26669]_  = ~A202 & ~A200;
  assign \new_[26670]_  = ~A199 & \new_[26669]_ ;
  assign \new_[26671]_  = \new_[26670]_  & \new_[26665]_ ;
  assign \new_[26675]_  = A298 & A234;
  assign \new_[26676]_  = A232 & \new_[26675]_ ;
  assign \new_[26680]_  = ~A301 & ~A300;
  assign \new_[26681]_  = A299 & \new_[26680]_ ;
  assign \new_[26682]_  = \new_[26681]_  & \new_[26676]_ ;
  assign \new_[26686]_  = A166 & ~A167;
  assign \new_[26687]_  = A170 & \new_[26686]_ ;
  assign \new_[26691]_  = ~A202 & ~A200;
  assign \new_[26692]_  = ~A199 & \new_[26691]_ ;
  assign \new_[26693]_  = \new_[26692]_  & \new_[26687]_ ;
  assign \new_[26697]_  = A298 & A234;
  assign \new_[26698]_  = A233 & \new_[26697]_ ;
  assign \new_[26702]_  = ~A301 & ~A300;
  assign \new_[26703]_  = A299 & \new_[26702]_ ;
  assign \new_[26704]_  = \new_[26703]_  & \new_[26698]_ ;
  assign \new_[26708]_  = A166 & ~A167;
  assign \new_[26709]_  = A170 & \new_[26708]_ ;
  assign \new_[26713]_  = ~A202 & ~A200;
  assign \new_[26714]_  = ~A199 & \new_[26713]_ ;
  assign \new_[26715]_  = \new_[26714]_  & \new_[26709]_ ;
  assign \new_[26719]_  = A236 & A233;
  assign \new_[26720]_  = ~A232 & \new_[26719]_ ;
  assign \new_[26724]_  = ~A302 & ~A301;
  assign \new_[26725]_  = ~A300 & \new_[26724]_ ;
  assign \new_[26726]_  = \new_[26725]_  & \new_[26720]_ ;
  assign \new_[26730]_  = A166 & ~A167;
  assign \new_[26731]_  = A170 & \new_[26730]_ ;
  assign \new_[26735]_  = ~A202 & ~A200;
  assign \new_[26736]_  = ~A199 & \new_[26735]_ ;
  assign \new_[26737]_  = \new_[26736]_  & \new_[26731]_ ;
  assign \new_[26741]_  = A236 & A233;
  assign \new_[26742]_  = ~A232 & \new_[26741]_ ;
  assign \new_[26746]_  = ~A301 & ~A299;
  assign \new_[26747]_  = ~A298 & \new_[26746]_ ;
  assign \new_[26748]_  = \new_[26747]_  & \new_[26742]_ ;
  assign \new_[26752]_  = A166 & ~A167;
  assign \new_[26753]_  = A170 & \new_[26752]_ ;
  assign \new_[26757]_  = ~A202 & ~A200;
  assign \new_[26758]_  = ~A199 & \new_[26757]_ ;
  assign \new_[26759]_  = \new_[26758]_  & \new_[26753]_ ;
  assign \new_[26763]_  = A236 & A233;
  assign \new_[26764]_  = ~A232 & \new_[26763]_ ;
  assign \new_[26768]_  = A269 & A266;
  assign \new_[26769]_  = ~A265 & \new_[26768]_ ;
  assign \new_[26770]_  = \new_[26769]_  & \new_[26764]_ ;
  assign \new_[26774]_  = A166 & ~A167;
  assign \new_[26775]_  = A170 & \new_[26774]_ ;
  assign \new_[26779]_  = ~A202 & ~A200;
  assign \new_[26780]_  = ~A199 & \new_[26779]_ ;
  assign \new_[26781]_  = \new_[26780]_  & \new_[26775]_ ;
  assign \new_[26785]_  = A236 & A233;
  assign \new_[26786]_  = ~A232 & \new_[26785]_ ;
  assign \new_[26790]_  = A269 & ~A266;
  assign \new_[26791]_  = A265 & \new_[26790]_ ;
  assign \new_[26792]_  = \new_[26791]_  & \new_[26786]_ ;
  assign \new_[26796]_  = A166 & ~A167;
  assign \new_[26797]_  = A170 & \new_[26796]_ ;
  assign \new_[26801]_  = ~A202 & ~A200;
  assign \new_[26802]_  = ~A199 & \new_[26801]_ ;
  assign \new_[26803]_  = \new_[26802]_  & \new_[26797]_ ;
  assign \new_[26807]_  = A236 & ~A233;
  assign \new_[26808]_  = A232 & \new_[26807]_ ;
  assign \new_[26812]_  = ~A302 & ~A301;
  assign \new_[26813]_  = ~A300 & \new_[26812]_ ;
  assign \new_[26814]_  = \new_[26813]_  & \new_[26808]_ ;
  assign \new_[26818]_  = A166 & ~A167;
  assign \new_[26819]_  = A170 & \new_[26818]_ ;
  assign \new_[26823]_  = ~A202 & ~A200;
  assign \new_[26824]_  = ~A199 & \new_[26823]_ ;
  assign \new_[26825]_  = \new_[26824]_  & \new_[26819]_ ;
  assign \new_[26829]_  = A236 & ~A233;
  assign \new_[26830]_  = A232 & \new_[26829]_ ;
  assign \new_[26834]_  = ~A301 & ~A299;
  assign \new_[26835]_  = ~A298 & \new_[26834]_ ;
  assign \new_[26836]_  = \new_[26835]_  & \new_[26830]_ ;
  assign \new_[26840]_  = A166 & ~A167;
  assign \new_[26841]_  = A170 & \new_[26840]_ ;
  assign \new_[26845]_  = ~A202 & ~A200;
  assign \new_[26846]_  = ~A199 & \new_[26845]_ ;
  assign \new_[26847]_  = \new_[26846]_  & \new_[26841]_ ;
  assign \new_[26851]_  = A236 & ~A233;
  assign \new_[26852]_  = A232 & \new_[26851]_ ;
  assign \new_[26856]_  = A269 & A266;
  assign \new_[26857]_  = ~A265 & \new_[26856]_ ;
  assign \new_[26858]_  = \new_[26857]_  & \new_[26852]_ ;
  assign \new_[26862]_  = A166 & ~A167;
  assign \new_[26863]_  = A170 & \new_[26862]_ ;
  assign \new_[26867]_  = ~A202 & ~A200;
  assign \new_[26868]_  = ~A199 & \new_[26867]_ ;
  assign \new_[26869]_  = \new_[26868]_  & \new_[26863]_ ;
  assign \new_[26873]_  = A236 & ~A233;
  assign \new_[26874]_  = A232 & \new_[26873]_ ;
  assign \new_[26878]_  = A269 & ~A266;
  assign \new_[26879]_  = A265 & \new_[26878]_ ;
  assign \new_[26880]_  = \new_[26879]_  & \new_[26874]_ ;
  assign \new_[26884]_  = ~A202 & ~A201;
  assign \new_[26885]_  = A169 & \new_[26884]_ ;
  assign \new_[26889]_  = ~A235 & ~A234;
  assign \new_[26890]_  = ~A203 & \new_[26889]_ ;
  assign \new_[26891]_  = \new_[26890]_  & \new_[26885]_ ;
  assign \new_[26895]_  = ~A268 & ~A267;
  assign \new_[26896]_  = ~A236 & \new_[26895]_ ;
  assign \new_[26900]_  = A300 & A299;
  assign \new_[26901]_  = ~A269 & \new_[26900]_ ;
  assign \new_[26902]_  = \new_[26901]_  & \new_[26896]_ ;
  assign \new_[26906]_  = ~A202 & ~A201;
  assign \new_[26907]_  = A169 & \new_[26906]_ ;
  assign \new_[26911]_  = ~A235 & ~A234;
  assign \new_[26912]_  = ~A203 & \new_[26911]_ ;
  assign \new_[26913]_  = \new_[26912]_  & \new_[26907]_ ;
  assign \new_[26917]_  = ~A268 & ~A267;
  assign \new_[26918]_  = ~A236 & \new_[26917]_ ;
  assign \new_[26922]_  = A300 & A298;
  assign \new_[26923]_  = ~A269 & \new_[26922]_ ;
  assign \new_[26924]_  = \new_[26923]_  & \new_[26918]_ ;
  assign \new_[26928]_  = ~A202 & ~A201;
  assign \new_[26929]_  = A169 & \new_[26928]_ ;
  assign \new_[26933]_  = ~A235 & ~A234;
  assign \new_[26934]_  = ~A203 & \new_[26933]_ ;
  assign \new_[26935]_  = \new_[26934]_  & \new_[26929]_ ;
  assign \new_[26939]_  = A266 & A265;
  assign \new_[26940]_  = ~A236 & \new_[26939]_ ;
  assign \new_[26944]_  = A301 & ~A268;
  assign \new_[26945]_  = ~A267 & \new_[26944]_ ;
  assign \new_[26946]_  = \new_[26945]_  & \new_[26940]_ ;
  assign \new_[26950]_  = ~A202 & ~A201;
  assign \new_[26951]_  = A169 & \new_[26950]_ ;
  assign \new_[26955]_  = ~A235 & ~A234;
  assign \new_[26956]_  = ~A203 & \new_[26955]_ ;
  assign \new_[26957]_  = \new_[26956]_  & \new_[26951]_ ;
  assign \new_[26961]_  = ~A266 & ~A265;
  assign \new_[26962]_  = ~A236 & \new_[26961]_ ;
  assign \new_[26966]_  = A300 & A299;
  assign \new_[26967]_  = ~A268 & \new_[26966]_ ;
  assign \new_[26968]_  = \new_[26967]_  & \new_[26962]_ ;
  assign \new_[26972]_  = ~A202 & ~A201;
  assign \new_[26973]_  = A169 & \new_[26972]_ ;
  assign \new_[26977]_  = ~A235 & ~A234;
  assign \new_[26978]_  = ~A203 & \new_[26977]_ ;
  assign \new_[26979]_  = \new_[26978]_  & \new_[26973]_ ;
  assign \new_[26983]_  = ~A266 & ~A265;
  assign \new_[26984]_  = ~A236 & \new_[26983]_ ;
  assign \new_[26988]_  = A300 & A298;
  assign \new_[26989]_  = ~A268 & \new_[26988]_ ;
  assign \new_[26990]_  = \new_[26989]_  & \new_[26984]_ ;
  assign \new_[26994]_  = ~A202 & ~A201;
  assign \new_[26995]_  = A169 & \new_[26994]_ ;
  assign \new_[26999]_  = A233 & A232;
  assign \new_[27000]_  = ~A203 & \new_[26999]_ ;
  assign \new_[27001]_  = \new_[27000]_  & \new_[26995]_ ;
  assign \new_[27005]_  = ~A267 & ~A235;
  assign \new_[27006]_  = ~A234 & \new_[27005]_ ;
  assign \new_[27010]_  = A301 & ~A269;
  assign \new_[27011]_  = ~A268 & \new_[27010]_ ;
  assign \new_[27012]_  = \new_[27011]_  & \new_[27006]_ ;
  assign \new_[27016]_  = ~A202 & ~A201;
  assign \new_[27017]_  = A169 & \new_[27016]_ ;
  assign \new_[27021]_  = A233 & A232;
  assign \new_[27022]_  = ~A203 & \new_[27021]_ ;
  assign \new_[27023]_  = \new_[27022]_  & \new_[27017]_ ;
  assign \new_[27027]_  = ~A265 & ~A235;
  assign \new_[27028]_  = ~A234 & \new_[27027]_ ;
  assign \new_[27032]_  = A301 & ~A268;
  assign \new_[27033]_  = ~A266 & \new_[27032]_ ;
  assign \new_[27034]_  = \new_[27033]_  & \new_[27028]_ ;
  assign \new_[27038]_  = ~A202 & ~A201;
  assign \new_[27039]_  = A169 & \new_[27038]_ ;
  assign \new_[27043]_  = ~A233 & ~A232;
  assign \new_[27044]_  = ~A203 & \new_[27043]_ ;
  assign \new_[27045]_  = \new_[27044]_  & \new_[27039]_ ;
  assign \new_[27049]_  = ~A268 & ~A267;
  assign \new_[27050]_  = ~A235 & \new_[27049]_ ;
  assign \new_[27054]_  = A300 & A299;
  assign \new_[27055]_  = ~A269 & \new_[27054]_ ;
  assign \new_[27056]_  = \new_[27055]_  & \new_[27050]_ ;
  assign \new_[27060]_  = ~A202 & ~A201;
  assign \new_[27061]_  = A169 & \new_[27060]_ ;
  assign \new_[27065]_  = ~A233 & ~A232;
  assign \new_[27066]_  = ~A203 & \new_[27065]_ ;
  assign \new_[27067]_  = \new_[27066]_  & \new_[27061]_ ;
  assign \new_[27071]_  = ~A268 & ~A267;
  assign \new_[27072]_  = ~A235 & \new_[27071]_ ;
  assign \new_[27076]_  = A300 & A298;
  assign \new_[27077]_  = ~A269 & \new_[27076]_ ;
  assign \new_[27078]_  = \new_[27077]_  & \new_[27072]_ ;
  assign \new_[27082]_  = ~A202 & ~A201;
  assign \new_[27083]_  = A169 & \new_[27082]_ ;
  assign \new_[27087]_  = ~A233 & ~A232;
  assign \new_[27088]_  = ~A203 & \new_[27087]_ ;
  assign \new_[27089]_  = \new_[27088]_  & \new_[27083]_ ;
  assign \new_[27093]_  = A266 & A265;
  assign \new_[27094]_  = ~A235 & \new_[27093]_ ;
  assign \new_[27098]_  = A301 & ~A268;
  assign \new_[27099]_  = ~A267 & \new_[27098]_ ;
  assign \new_[27100]_  = \new_[27099]_  & \new_[27094]_ ;
  assign \new_[27104]_  = ~A202 & ~A201;
  assign \new_[27105]_  = A169 & \new_[27104]_ ;
  assign \new_[27109]_  = ~A233 & ~A232;
  assign \new_[27110]_  = ~A203 & \new_[27109]_ ;
  assign \new_[27111]_  = \new_[27110]_  & \new_[27105]_ ;
  assign \new_[27115]_  = ~A266 & ~A265;
  assign \new_[27116]_  = ~A235 & \new_[27115]_ ;
  assign \new_[27120]_  = A300 & A299;
  assign \new_[27121]_  = ~A268 & \new_[27120]_ ;
  assign \new_[27122]_  = \new_[27121]_  & \new_[27116]_ ;
  assign \new_[27126]_  = ~A202 & ~A201;
  assign \new_[27127]_  = A169 & \new_[27126]_ ;
  assign \new_[27131]_  = ~A233 & ~A232;
  assign \new_[27132]_  = ~A203 & \new_[27131]_ ;
  assign \new_[27133]_  = \new_[27132]_  & \new_[27127]_ ;
  assign \new_[27137]_  = ~A266 & ~A265;
  assign \new_[27138]_  = ~A235 & \new_[27137]_ ;
  assign \new_[27142]_  = A300 & A298;
  assign \new_[27143]_  = ~A268 & \new_[27142]_ ;
  assign \new_[27144]_  = \new_[27143]_  & \new_[27138]_ ;
  assign \new_[27148]_  = A200 & A199;
  assign \new_[27149]_  = A169 & \new_[27148]_ ;
  assign \new_[27153]_  = ~A234 & ~A202;
  assign \new_[27154]_  = ~A201 & \new_[27153]_ ;
  assign \new_[27155]_  = \new_[27154]_  & \new_[27149]_ ;
  assign \new_[27159]_  = ~A267 & ~A236;
  assign \new_[27160]_  = ~A235 & \new_[27159]_ ;
  assign \new_[27164]_  = A301 & ~A269;
  assign \new_[27165]_  = ~A268 & \new_[27164]_ ;
  assign \new_[27166]_  = \new_[27165]_  & \new_[27160]_ ;
  assign \new_[27170]_  = A200 & A199;
  assign \new_[27171]_  = A169 & \new_[27170]_ ;
  assign \new_[27175]_  = ~A234 & ~A202;
  assign \new_[27176]_  = ~A201 & \new_[27175]_ ;
  assign \new_[27177]_  = \new_[27176]_  & \new_[27171]_ ;
  assign \new_[27181]_  = ~A265 & ~A236;
  assign \new_[27182]_  = ~A235 & \new_[27181]_ ;
  assign \new_[27186]_  = A301 & ~A268;
  assign \new_[27187]_  = ~A266 & \new_[27186]_ ;
  assign \new_[27188]_  = \new_[27187]_  & \new_[27182]_ ;
  assign \new_[27192]_  = A200 & A199;
  assign \new_[27193]_  = A169 & \new_[27192]_ ;
  assign \new_[27197]_  = ~A232 & ~A202;
  assign \new_[27198]_  = ~A201 & \new_[27197]_ ;
  assign \new_[27199]_  = \new_[27198]_  & \new_[27193]_ ;
  assign \new_[27203]_  = A298 & A236;
  assign \new_[27204]_  = A233 & \new_[27203]_ ;
  assign \new_[27208]_  = ~A301 & ~A300;
  assign \new_[27209]_  = A299 & \new_[27208]_ ;
  assign \new_[27210]_  = \new_[27209]_  & \new_[27204]_ ;
  assign \new_[27214]_  = A200 & A199;
  assign \new_[27215]_  = A169 & \new_[27214]_ ;
  assign \new_[27219]_  = A232 & ~A202;
  assign \new_[27220]_  = ~A201 & \new_[27219]_ ;
  assign \new_[27221]_  = \new_[27220]_  & \new_[27215]_ ;
  assign \new_[27225]_  = A298 & A236;
  assign \new_[27226]_  = ~A233 & \new_[27225]_ ;
  assign \new_[27230]_  = ~A301 & ~A300;
  assign \new_[27231]_  = A299 & \new_[27230]_ ;
  assign \new_[27232]_  = \new_[27231]_  & \new_[27226]_ ;
  assign \new_[27236]_  = A200 & A199;
  assign \new_[27237]_  = A169 & \new_[27236]_ ;
  assign \new_[27241]_  = ~A232 & ~A202;
  assign \new_[27242]_  = ~A201 & \new_[27241]_ ;
  assign \new_[27243]_  = \new_[27242]_  & \new_[27237]_ ;
  assign \new_[27247]_  = ~A267 & ~A235;
  assign \new_[27248]_  = ~A233 & \new_[27247]_ ;
  assign \new_[27252]_  = A301 & ~A269;
  assign \new_[27253]_  = ~A268 & \new_[27252]_ ;
  assign \new_[27254]_  = \new_[27253]_  & \new_[27248]_ ;
  assign \new_[27258]_  = A200 & A199;
  assign \new_[27259]_  = A169 & \new_[27258]_ ;
  assign \new_[27263]_  = ~A232 & ~A202;
  assign \new_[27264]_  = ~A201 & \new_[27263]_ ;
  assign \new_[27265]_  = \new_[27264]_  & \new_[27259]_ ;
  assign \new_[27269]_  = ~A265 & ~A235;
  assign \new_[27270]_  = ~A233 & \new_[27269]_ ;
  assign \new_[27274]_  = A301 & ~A268;
  assign \new_[27275]_  = ~A266 & \new_[27274]_ ;
  assign \new_[27276]_  = \new_[27275]_  & \new_[27270]_ ;
  assign \new_[27280]_  = ~A200 & ~A199;
  assign \new_[27281]_  = A169 & \new_[27280]_ ;
  assign \new_[27285]_  = ~A235 & ~A234;
  assign \new_[27286]_  = ~A202 & \new_[27285]_ ;
  assign \new_[27287]_  = \new_[27286]_  & \new_[27281]_ ;
  assign \new_[27291]_  = ~A268 & ~A267;
  assign \new_[27292]_  = ~A236 & \new_[27291]_ ;
  assign \new_[27296]_  = A300 & A299;
  assign \new_[27297]_  = ~A269 & \new_[27296]_ ;
  assign \new_[27298]_  = \new_[27297]_  & \new_[27292]_ ;
  assign \new_[27302]_  = ~A200 & ~A199;
  assign \new_[27303]_  = A169 & \new_[27302]_ ;
  assign \new_[27307]_  = ~A235 & ~A234;
  assign \new_[27308]_  = ~A202 & \new_[27307]_ ;
  assign \new_[27309]_  = \new_[27308]_  & \new_[27303]_ ;
  assign \new_[27313]_  = ~A268 & ~A267;
  assign \new_[27314]_  = ~A236 & \new_[27313]_ ;
  assign \new_[27318]_  = A300 & A298;
  assign \new_[27319]_  = ~A269 & \new_[27318]_ ;
  assign \new_[27320]_  = \new_[27319]_  & \new_[27314]_ ;
  assign \new_[27324]_  = ~A200 & ~A199;
  assign \new_[27325]_  = A169 & \new_[27324]_ ;
  assign \new_[27329]_  = ~A235 & ~A234;
  assign \new_[27330]_  = ~A202 & \new_[27329]_ ;
  assign \new_[27331]_  = \new_[27330]_  & \new_[27325]_ ;
  assign \new_[27335]_  = A266 & A265;
  assign \new_[27336]_  = ~A236 & \new_[27335]_ ;
  assign \new_[27340]_  = A301 & ~A268;
  assign \new_[27341]_  = ~A267 & \new_[27340]_ ;
  assign \new_[27342]_  = \new_[27341]_  & \new_[27336]_ ;
  assign \new_[27346]_  = ~A200 & ~A199;
  assign \new_[27347]_  = A169 & \new_[27346]_ ;
  assign \new_[27351]_  = ~A235 & ~A234;
  assign \new_[27352]_  = ~A202 & \new_[27351]_ ;
  assign \new_[27353]_  = \new_[27352]_  & \new_[27347]_ ;
  assign \new_[27357]_  = ~A266 & ~A265;
  assign \new_[27358]_  = ~A236 & \new_[27357]_ ;
  assign \new_[27362]_  = A300 & A299;
  assign \new_[27363]_  = ~A268 & \new_[27362]_ ;
  assign \new_[27364]_  = \new_[27363]_  & \new_[27358]_ ;
  assign \new_[27368]_  = ~A200 & ~A199;
  assign \new_[27369]_  = A169 & \new_[27368]_ ;
  assign \new_[27373]_  = ~A235 & ~A234;
  assign \new_[27374]_  = ~A202 & \new_[27373]_ ;
  assign \new_[27375]_  = \new_[27374]_  & \new_[27369]_ ;
  assign \new_[27379]_  = ~A266 & ~A265;
  assign \new_[27380]_  = ~A236 & \new_[27379]_ ;
  assign \new_[27384]_  = A300 & A298;
  assign \new_[27385]_  = ~A268 & \new_[27384]_ ;
  assign \new_[27386]_  = \new_[27385]_  & \new_[27380]_ ;
  assign \new_[27390]_  = ~A200 & ~A199;
  assign \new_[27391]_  = A169 & \new_[27390]_ ;
  assign \new_[27395]_  = A233 & A232;
  assign \new_[27396]_  = ~A202 & \new_[27395]_ ;
  assign \new_[27397]_  = \new_[27396]_  & \new_[27391]_ ;
  assign \new_[27401]_  = ~A267 & ~A235;
  assign \new_[27402]_  = ~A234 & \new_[27401]_ ;
  assign \new_[27406]_  = A301 & ~A269;
  assign \new_[27407]_  = ~A268 & \new_[27406]_ ;
  assign \new_[27408]_  = \new_[27407]_  & \new_[27402]_ ;
  assign \new_[27412]_  = ~A200 & ~A199;
  assign \new_[27413]_  = A169 & \new_[27412]_ ;
  assign \new_[27417]_  = A233 & A232;
  assign \new_[27418]_  = ~A202 & \new_[27417]_ ;
  assign \new_[27419]_  = \new_[27418]_  & \new_[27413]_ ;
  assign \new_[27423]_  = ~A265 & ~A235;
  assign \new_[27424]_  = ~A234 & \new_[27423]_ ;
  assign \new_[27428]_  = A301 & ~A268;
  assign \new_[27429]_  = ~A266 & \new_[27428]_ ;
  assign \new_[27430]_  = \new_[27429]_  & \new_[27424]_ ;
  assign \new_[27434]_  = ~A200 & ~A199;
  assign \new_[27435]_  = A169 & \new_[27434]_ ;
  assign \new_[27439]_  = ~A233 & ~A232;
  assign \new_[27440]_  = ~A202 & \new_[27439]_ ;
  assign \new_[27441]_  = \new_[27440]_  & \new_[27435]_ ;
  assign \new_[27445]_  = ~A268 & ~A267;
  assign \new_[27446]_  = ~A235 & \new_[27445]_ ;
  assign \new_[27450]_  = A300 & A299;
  assign \new_[27451]_  = ~A269 & \new_[27450]_ ;
  assign \new_[27452]_  = \new_[27451]_  & \new_[27446]_ ;
  assign \new_[27456]_  = ~A200 & ~A199;
  assign \new_[27457]_  = A169 & \new_[27456]_ ;
  assign \new_[27461]_  = ~A233 & ~A232;
  assign \new_[27462]_  = ~A202 & \new_[27461]_ ;
  assign \new_[27463]_  = \new_[27462]_  & \new_[27457]_ ;
  assign \new_[27467]_  = ~A268 & ~A267;
  assign \new_[27468]_  = ~A235 & \new_[27467]_ ;
  assign \new_[27472]_  = A300 & A298;
  assign \new_[27473]_  = ~A269 & \new_[27472]_ ;
  assign \new_[27474]_  = \new_[27473]_  & \new_[27468]_ ;
  assign \new_[27478]_  = ~A200 & ~A199;
  assign \new_[27479]_  = A169 & \new_[27478]_ ;
  assign \new_[27483]_  = ~A233 & ~A232;
  assign \new_[27484]_  = ~A202 & \new_[27483]_ ;
  assign \new_[27485]_  = \new_[27484]_  & \new_[27479]_ ;
  assign \new_[27489]_  = A266 & A265;
  assign \new_[27490]_  = ~A235 & \new_[27489]_ ;
  assign \new_[27494]_  = A301 & ~A268;
  assign \new_[27495]_  = ~A267 & \new_[27494]_ ;
  assign \new_[27496]_  = \new_[27495]_  & \new_[27490]_ ;
  assign \new_[27500]_  = ~A200 & ~A199;
  assign \new_[27501]_  = A169 & \new_[27500]_ ;
  assign \new_[27505]_  = ~A233 & ~A232;
  assign \new_[27506]_  = ~A202 & \new_[27505]_ ;
  assign \new_[27507]_  = \new_[27506]_  & \new_[27501]_ ;
  assign \new_[27511]_  = ~A266 & ~A265;
  assign \new_[27512]_  = ~A235 & \new_[27511]_ ;
  assign \new_[27516]_  = A300 & A299;
  assign \new_[27517]_  = ~A268 & \new_[27516]_ ;
  assign \new_[27518]_  = \new_[27517]_  & \new_[27512]_ ;
  assign \new_[27522]_  = ~A200 & ~A199;
  assign \new_[27523]_  = A169 & \new_[27522]_ ;
  assign \new_[27527]_  = ~A233 & ~A232;
  assign \new_[27528]_  = ~A202 & \new_[27527]_ ;
  assign \new_[27529]_  = \new_[27528]_  & \new_[27523]_ ;
  assign \new_[27533]_  = ~A266 & ~A265;
  assign \new_[27534]_  = ~A235 & \new_[27533]_ ;
  assign \new_[27538]_  = A300 & A298;
  assign \new_[27539]_  = ~A268 & \new_[27538]_ ;
  assign \new_[27540]_  = \new_[27539]_  & \new_[27534]_ ;
  assign \new_[27544]_  = ~A166 & ~A167;
  assign \new_[27545]_  = ~A169 & \new_[27544]_ ;
  assign \new_[27549]_  = ~A235 & ~A234;
  assign \new_[27550]_  = A202 & \new_[27549]_ ;
  assign \new_[27551]_  = \new_[27550]_  & \new_[27545]_ ;
  assign \new_[27555]_  = ~A268 & ~A267;
  assign \new_[27556]_  = ~A236 & \new_[27555]_ ;
  assign \new_[27560]_  = A300 & A299;
  assign \new_[27561]_  = ~A269 & \new_[27560]_ ;
  assign \new_[27562]_  = \new_[27561]_  & \new_[27556]_ ;
  assign \new_[27566]_  = ~A166 & ~A167;
  assign \new_[27567]_  = ~A169 & \new_[27566]_ ;
  assign \new_[27571]_  = ~A235 & ~A234;
  assign \new_[27572]_  = A202 & \new_[27571]_ ;
  assign \new_[27573]_  = \new_[27572]_  & \new_[27567]_ ;
  assign \new_[27577]_  = ~A268 & ~A267;
  assign \new_[27578]_  = ~A236 & \new_[27577]_ ;
  assign \new_[27582]_  = A300 & A298;
  assign \new_[27583]_  = ~A269 & \new_[27582]_ ;
  assign \new_[27584]_  = \new_[27583]_  & \new_[27578]_ ;
  assign \new_[27588]_  = ~A166 & ~A167;
  assign \new_[27589]_  = ~A169 & \new_[27588]_ ;
  assign \new_[27593]_  = ~A235 & ~A234;
  assign \new_[27594]_  = A202 & \new_[27593]_ ;
  assign \new_[27595]_  = \new_[27594]_  & \new_[27589]_ ;
  assign \new_[27599]_  = A266 & A265;
  assign \new_[27600]_  = ~A236 & \new_[27599]_ ;
  assign \new_[27604]_  = A301 & ~A268;
  assign \new_[27605]_  = ~A267 & \new_[27604]_ ;
  assign \new_[27606]_  = \new_[27605]_  & \new_[27600]_ ;
  assign \new_[27610]_  = ~A166 & ~A167;
  assign \new_[27611]_  = ~A169 & \new_[27610]_ ;
  assign \new_[27615]_  = ~A235 & ~A234;
  assign \new_[27616]_  = A202 & \new_[27615]_ ;
  assign \new_[27617]_  = \new_[27616]_  & \new_[27611]_ ;
  assign \new_[27621]_  = ~A266 & ~A265;
  assign \new_[27622]_  = ~A236 & \new_[27621]_ ;
  assign \new_[27626]_  = A300 & A299;
  assign \new_[27627]_  = ~A268 & \new_[27626]_ ;
  assign \new_[27628]_  = \new_[27627]_  & \new_[27622]_ ;
  assign \new_[27632]_  = ~A166 & ~A167;
  assign \new_[27633]_  = ~A169 & \new_[27632]_ ;
  assign \new_[27637]_  = ~A235 & ~A234;
  assign \new_[27638]_  = A202 & \new_[27637]_ ;
  assign \new_[27639]_  = \new_[27638]_  & \new_[27633]_ ;
  assign \new_[27643]_  = ~A266 & ~A265;
  assign \new_[27644]_  = ~A236 & \new_[27643]_ ;
  assign \new_[27648]_  = A300 & A298;
  assign \new_[27649]_  = ~A268 & \new_[27648]_ ;
  assign \new_[27650]_  = \new_[27649]_  & \new_[27644]_ ;
  assign \new_[27654]_  = ~A166 & ~A167;
  assign \new_[27655]_  = ~A169 & \new_[27654]_ ;
  assign \new_[27659]_  = A233 & A232;
  assign \new_[27660]_  = A202 & \new_[27659]_ ;
  assign \new_[27661]_  = \new_[27660]_  & \new_[27655]_ ;
  assign \new_[27665]_  = ~A267 & ~A235;
  assign \new_[27666]_  = ~A234 & \new_[27665]_ ;
  assign \new_[27670]_  = A301 & ~A269;
  assign \new_[27671]_  = ~A268 & \new_[27670]_ ;
  assign \new_[27672]_  = \new_[27671]_  & \new_[27666]_ ;
  assign \new_[27676]_  = ~A166 & ~A167;
  assign \new_[27677]_  = ~A169 & \new_[27676]_ ;
  assign \new_[27681]_  = A233 & A232;
  assign \new_[27682]_  = A202 & \new_[27681]_ ;
  assign \new_[27683]_  = \new_[27682]_  & \new_[27677]_ ;
  assign \new_[27687]_  = ~A265 & ~A235;
  assign \new_[27688]_  = ~A234 & \new_[27687]_ ;
  assign \new_[27692]_  = A301 & ~A268;
  assign \new_[27693]_  = ~A266 & \new_[27692]_ ;
  assign \new_[27694]_  = \new_[27693]_  & \new_[27688]_ ;
  assign \new_[27698]_  = ~A166 & ~A167;
  assign \new_[27699]_  = ~A169 & \new_[27698]_ ;
  assign \new_[27703]_  = ~A233 & ~A232;
  assign \new_[27704]_  = A202 & \new_[27703]_ ;
  assign \new_[27705]_  = \new_[27704]_  & \new_[27699]_ ;
  assign \new_[27709]_  = ~A268 & ~A267;
  assign \new_[27710]_  = ~A235 & \new_[27709]_ ;
  assign \new_[27714]_  = A300 & A299;
  assign \new_[27715]_  = ~A269 & \new_[27714]_ ;
  assign \new_[27716]_  = \new_[27715]_  & \new_[27710]_ ;
  assign \new_[27720]_  = ~A166 & ~A167;
  assign \new_[27721]_  = ~A169 & \new_[27720]_ ;
  assign \new_[27725]_  = ~A233 & ~A232;
  assign \new_[27726]_  = A202 & \new_[27725]_ ;
  assign \new_[27727]_  = \new_[27726]_  & \new_[27721]_ ;
  assign \new_[27731]_  = ~A268 & ~A267;
  assign \new_[27732]_  = ~A235 & \new_[27731]_ ;
  assign \new_[27736]_  = A300 & A298;
  assign \new_[27737]_  = ~A269 & \new_[27736]_ ;
  assign \new_[27738]_  = \new_[27737]_  & \new_[27732]_ ;
  assign \new_[27742]_  = ~A166 & ~A167;
  assign \new_[27743]_  = ~A169 & \new_[27742]_ ;
  assign \new_[27747]_  = ~A233 & ~A232;
  assign \new_[27748]_  = A202 & \new_[27747]_ ;
  assign \new_[27749]_  = \new_[27748]_  & \new_[27743]_ ;
  assign \new_[27753]_  = A266 & A265;
  assign \new_[27754]_  = ~A235 & \new_[27753]_ ;
  assign \new_[27758]_  = A301 & ~A268;
  assign \new_[27759]_  = ~A267 & \new_[27758]_ ;
  assign \new_[27760]_  = \new_[27759]_  & \new_[27754]_ ;
  assign \new_[27764]_  = ~A166 & ~A167;
  assign \new_[27765]_  = ~A169 & \new_[27764]_ ;
  assign \new_[27769]_  = ~A233 & ~A232;
  assign \new_[27770]_  = A202 & \new_[27769]_ ;
  assign \new_[27771]_  = \new_[27770]_  & \new_[27765]_ ;
  assign \new_[27775]_  = ~A266 & ~A265;
  assign \new_[27776]_  = ~A235 & \new_[27775]_ ;
  assign \new_[27780]_  = A300 & A299;
  assign \new_[27781]_  = ~A268 & \new_[27780]_ ;
  assign \new_[27782]_  = \new_[27781]_  & \new_[27776]_ ;
  assign \new_[27786]_  = ~A166 & ~A167;
  assign \new_[27787]_  = ~A169 & \new_[27786]_ ;
  assign \new_[27791]_  = ~A233 & ~A232;
  assign \new_[27792]_  = A202 & \new_[27791]_ ;
  assign \new_[27793]_  = \new_[27792]_  & \new_[27787]_ ;
  assign \new_[27797]_  = ~A266 & ~A265;
  assign \new_[27798]_  = ~A235 & \new_[27797]_ ;
  assign \new_[27802]_  = A300 & A298;
  assign \new_[27803]_  = ~A268 & \new_[27802]_ ;
  assign \new_[27804]_  = \new_[27803]_  & \new_[27798]_ ;
  assign \new_[27808]_  = ~A166 & ~A167;
  assign \new_[27809]_  = ~A169 & \new_[27808]_ ;
  assign \new_[27813]_  = ~A234 & A201;
  assign \new_[27814]_  = A199 & \new_[27813]_ ;
  assign \new_[27815]_  = \new_[27814]_  & \new_[27809]_ ;
  assign \new_[27819]_  = ~A267 & ~A236;
  assign \new_[27820]_  = ~A235 & \new_[27819]_ ;
  assign \new_[27824]_  = A301 & ~A269;
  assign \new_[27825]_  = ~A268 & \new_[27824]_ ;
  assign \new_[27826]_  = \new_[27825]_  & \new_[27820]_ ;
  assign \new_[27830]_  = ~A166 & ~A167;
  assign \new_[27831]_  = ~A169 & \new_[27830]_ ;
  assign \new_[27835]_  = ~A234 & A201;
  assign \new_[27836]_  = A199 & \new_[27835]_ ;
  assign \new_[27837]_  = \new_[27836]_  & \new_[27831]_ ;
  assign \new_[27841]_  = ~A265 & ~A236;
  assign \new_[27842]_  = ~A235 & \new_[27841]_ ;
  assign \new_[27846]_  = A301 & ~A268;
  assign \new_[27847]_  = ~A266 & \new_[27846]_ ;
  assign \new_[27848]_  = \new_[27847]_  & \new_[27842]_ ;
  assign \new_[27852]_  = ~A166 & ~A167;
  assign \new_[27853]_  = ~A169 & \new_[27852]_ ;
  assign \new_[27857]_  = ~A232 & A201;
  assign \new_[27858]_  = A199 & \new_[27857]_ ;
  assign \new_[27859]_  = \new_[27858]_  & \new_[27853]_ ;
  assign \new_[27863]_  = A298 & A236;
  assign \new_[27864]_  = A233 & \new_[27863]_ ;
  assign \new_[27868]_  = ~A301 & ~A300;
  assign \new_[27869]_  = A299 & \new_[27868]_ ;
  assign \new_[27870]_  = \new_[27869]_  & \new_[27864]_ ;
  assign \new_[27874]_  = ~A166 & ~A167;
  assign \new_[27875]_  = ~A169 & \new_[27874]_ ;
  assign \new_[27879]_  = A232 & A201;
  assign \new_[27880]_  = A199 & \new_[27879]_ ;
  assign \new_[27881]_  = \new_[27880]_  & \new_[27875]_ ;
  assign \new_[27885]_  = A298 & A236;
  assign \new_[27886]_  = ~A233 & \new_[27885]_ ;
  assign \new_[27890]_  = ~A301 & ~A300;
  assign \new_[27891]_  = A299 & \new_[27890]_ ;
  assign \new_[27892]_  = \new_[27891]_  & \new_[27886]_ ;
  assign \new_[27896]_  = ~A166 & ~A167;
  assign \new_[27897]_  = ~A169 & \new_[27896]_ ;
  assign \new_[27901]_  = ~A232 & A201;
  assign \new_[27902]_  = A199 & \new_[27901]_ ;
  assign \new_[27903]_  = \new_[27902]_  & \new_[27897]_ ;
  assign \new_[27907]_  = ~A267 & ~A235;
  assign \new_[27908]_  = ~A233 & \new_[27907]_ ;
  assign \new_[27912]_  = A301 & ~A269;
  assign \new_[27913]_  = ~A268 & \new_[27912]_ ;
  assign \new_[27914]_  = \new_[27913]_  & \new_[27908]_ ;
  assign \new_[27918]_  = ~A166 & ~A167;
  assign \new_[27919]_  = ~A169 & \new_[27918]_ ;
  assign \new_[27923]_  = ~A232 & A201;
  assign \new_[27924]_  = A199 & \new_[27923]_ ;
  assign \new_[27925]_  = \new_[27924]_  & \new_[27919]_ ;
  assign \new_[27929]_  = ~A265 & ~A235;
  assign \new_[27930]_  = ~A233 & \new_[27929]_ ;
  assign \new_[27934]_  = A301 & ~A268;
  assign \new_[27935]_  = ~A266 & \new_[27934]_ ;
  assign \new_[27936]_  = \new_[27935]_  & \new_[27930]_ ;
  assign \new_[27940]_  = ~A166 & ~A167;
  assign \new_[27941]_  = ~A169 & \new_[27940]_ ;
  assign \new_[27945]_  = ~A234 & A201;
  assign \new_[27946]_  = A200 & \new_[27945]_ ;
  assign \new_[27947]_  = \new_[27946]_  & \new_[27941]_ ;
  assign \new_[27951]_  = ~A267 & ~A236;
  assign \new_[27952]_  = ~A235 & \new_[27951]_ ;
  assign \new_[27956]_  = A301 & ~A269;
  assign \new_[27957]_  = ~A268 & \new_[27956]_ ;
  assign \new_[27958]_  = \new_[27957]_  & \new_[27952]_ ;
  assign \new_[27962]_  = ~A166 & ~A167;
  assign \new_[27963]_  = ~A169 & \new_[27962]_ ;
  assign \new_[27967]_  = ~A234 & A201;
  assign \new_[27968]_  = A200 & \new_[27967]_ ;
  assign \new_[27969]_  = \new_[27968]_  & \new_[27963]_ ;
  assign \new_[27973]_  = ~A265 & ~A236;
  assign \new_[27974]_  = ~A235 & \new_[27973]_ ;
  assign \new_[27978]_  = A301 & ~A268;
  assign \new_[27979]_  = ~A266 & \new_[27978]_ ;
  assign \new_[27980]_  = \new_[27979]_  & \new_[27974]_ ;
  assign \new_[27984]_  = ~A166 & ~A167;
  assign \new_[27985]_  = ~A169 & \new_[27984]_ ;
  assign \new_[27989]_  = ~A232 & A201;
  assign \new_[27990]_  = A200 & \new_[27989]_ ;
  assign \new_[27991]_  = \new_[27990]_  & \new_[27985]_ ;
  assign \new_[27995]_  = A298 & A236;
  assign \new_[27996]_  = A233 & \new_[27995]_ ;
  assign \new_[28000]_  = ~A301 & ~A300;
  assign \new_[28001]_  = A299 & \new_[28000]_ ;
  assign \new_[28002]_  = \new_[28001]_  & \new_[27996]_ ;
  assign \new_[28006]_  = ~A166 & ~A167;
  assign \new_[28007]_  = ~A169 & \new_[28006]_ ;
  assign \new_[28011]_  = A232 & A201;
  assign \new_[28012]_  = A200 & \new_[28011]_ ;
  assign \new_[28013]_  = \new_[28012]_  & \new_[28007]_ ;
  assign \new_[28017]_  = A298 & A236;
  assign \new_[28018]_  = ~A233 & \new_[28017]_ ;
  assign \new_[28022]_  = ~A301 & ~A300;
  assign \new_[28023]_  = A299 & \new_[28022]_ ;
  assign \new_[28024]_  = \new_[28023]_  & \new_[28018]_ ;
  assign \new_[28028]_  = ~A166 & ~A167;
  assign \new_[28029]_  = ~A169 & \new_[28028]_ ;
  assign \new_[28033]_  = ~A232 & A201;
  assign \new_[28034]_  = A200 & \new_[28033]_ ;
  assign \new_[28035]_  = \new_[28034]_  & \new_[28029]_ ;
  assign \new_[28039]_  = ~A267 & ~A235;
  assign \new_[28040]_  = ~A233 & \new_[28039]_ ;
  assign \new_[28044]_  = A301 & ~A269;
  assign \new_[28045]_  = ~A268 & \new_[28044]_ ;
  assign \new_[28046]_  = \new_[28045]_  & \new_[28040]_ ;
  assign \new_[28050]_  = ~A166 & ~A167;
  assign \new_[28051]_  = ~A169 & \new_[28050]_ ;
  assign \new_[28055]_  = ~A232 & A201;
  assign \new_[28056]_  = A200 & \new_[28055]_ ;
  assign \new_[28057]_  = \new_[28056]_  & \new_[28051]_ ;
  assign \new_[28061]_  = ~A265 & ~A235;
  assign \new_[28062]_  = ~A233 & \new_[28061]_ ;
  assign \new_[28066]_  = A301 & ~A268;
  assign \new_[28067]_  = ~A266 & \new_[28066]_ ;
  assign \new_[28068]_  = \new_[28067]_  & \new_[28062]_ ;
  assign \new_[28072]_  = ~A166 & ~A167;
  assign \new_[28073]_  = ~A169 & \new_[28072]_ ;
  assign \new_[28077]_  = A203 & A200;
  assign \new_[28078]_  = ~A199 & \new_[28077]_ ;
  assign \new_[28079]_  = \new_[28078]_  & \new_[28073]_ ;
  assign \new_[28083]_  = A298 & A234;
  assign \new_[28084]_  = A232 & \new_[28083]_ ;
  assign \new_[28088]_  = ~A301 & ~A300;
  assign \new_[28089]_  = A299 & \new_[28088]_ ;
  assign \new_[28090]_  = \new_[28089]_  & \new_[28084]_ ;
  assign \new_[28094]_  = ~A166 & ~A167;
  assign \new_[28095]_  = ~A169 & \new_[28094]_ ;
  assign \new_[28099]_  = A203 & A200;
  assign \new_[28100]_  = ~A199 & \new_[28099]_ ;
  assign \new_[28101]_  = \new_[28100]_  & \new_[28095]_ ;
  assign \new_[28105]_  = A298 & A234;
  assign \new_[28106]_  = A233 & \new_[28105]_ ;
  assign \new_[28110]_  = ~A301 & ~A300;
  assign \new_[28111]_  = A299 & \new_[28110]_ ;
  assign \new_[28112]_  = \new_[28111]_  & \new_[28106]_ ;
  assign \new_[28116]_  = ~A166 & ~A167;
  assign \new_[28117]_  = ~A169 & \new_[28116]_ ;
  assign \new_[28121]_  = A203 & A200;
  assign \new_[28122]_  = ~A199 & \new_[28121]_ ;
  assign \new_[28123]_  = \new_[28122]_  & \new_[28117]_ ;
  assign \new_[28127]_  = A236 & A233;
  assign \new_[28128]_  = ~A232 & \new_[28127]_ ;
  assign \new_[28132]_  = ~A302 & ~A301;
  assign \new_[28133]_  = ~A300 & \new_[28132]_ ;
  assign \new_[28134]_  = \new_[28133]_  & \new_[28128]_ ;
  assign \new_[28138]_  = ~A166 & ~A167;
  assign \new_[28139]_  = ~A169 & \new_[28138]_ ;
  assign \new_[28143]_  = A203 & A200;
  assign \new_[28144]_  = ~A199 & \new_[28143]_ ;
  assign \new_[28145]_  = \new_[28144]_  & \new_[28139]_ ;
  assign \new_[28149]_  = A236 & A233;
  assign \new_[28150]_  = ~A232 & \new_[28149]_ ;
  assign \new_[28154]_  = ~A301 & ~A299;
  assign \new_[28155]_  = ~A298 & \new_[28154]_ ;
  assign \new_[28156]_  = \new_[28155]_  & \new_[28150]_ ;
  assign \new_[28160]_  = ~A166 & ~A167;
  assign \new_[28161]_  = ~A169 & \new_[28160]_ ;
  assign \new_[28165]_  = A203 & A200;
  assign \new_[28166]_  = ~A199 & \new_[28165]_ ;
  assign \new_[28167]_  = \new_[28166]_  & \new_[28161]_ ;
  assign \new_[28171]_  = A236 & A233;
  assign \new_[28172]_  = ~A232 & \new_[28171]_ ;
  assign \new_[28176]_  = A269 & A266;
  assign \new_[28177]_  = ~A265 & \new_[28176]_ ;
  assign \new_[28178]_  = \new_[28177]_  & \new_[28172]_ ;
  assign \new_[28182]_  = ~A166 & ~A167;
  assign \new_[28183]_  = ~A169 & \new_[28182]_ ;
  assign \new_[28187]_  = A203 & A200;
  assign \new_[28188]_  = ~A199 & \new_[28187]_ ;
  assign \new_[28189]_  = \new_[28188]_  & \new_[28183]_ ;
  assign \new_[28193]_  = A236 & A233;
  assign \new_[28194]_  = ~A232 & \new_[28193]_ ;
  assign \new_[28198]_  = A269 & ~A266;
  assign \new_[28199]_  = A265 & \new_[28198]_ ;
  assign \new_[28200]_  = \new_[28199]_  & \new_[28194]_ ;
  assign \new_[28204]_  = ~A166 & ~A167;
  assign \new_[28205]_  = ~A169 & \new_[28204]_ ;
  assign \new_[28209]_  = A203 & A200;
  assign \new_[28210]_  = ~A199 & \new_[28209]_ ;
  assign \new_[28211]_  = \new_[28210]_  & \new_[28205]_ ;
  assign \new_[28215]_  = A236 & ~A233;
  assign \new_[28216]_  = A232 & \new_[28215]_ ;
  assign \new_[28220]_  = ~A302 & ~A301;
  assign \new_[28221]_  = ~A300 & \new_[28220]_ ;
  assign \new_[28222]_  = \new_[28221]_  & \new_[28216]_ ;
  assign \new_[28226]_  = ~A166 & ~A167;
  assign \new_[28227]_  = ~A169 & \new_[28226]_ ;
  assign \new_[28231]_  = A203 & A200;
  assign \new_[28232]_  = ~A199 & \new_[28231]_ ;
  assign \new_[28233]_  = \new_[28232]_  & \new_[28227]_ ;
  assign \new_[28237]_  = A236 & ~A233;
  assign \new_[28238]_  = A232 & \new_[28237]_ ;
  assign \new_[28242]_  = ~A301 & ~A299;
  assign \new_[28243]_  = ~A298 & \new_[28242]_ ;
  assign \new_[28244]_  = \new_[28243]_  & \new_[28238]_ ;
  assign \new_[28248]_  = ~A166 & ~A167;
  assign \new_[28249]_  = ~A169 & \new_[28248]_ ;
  assign \new_[28253]_  = A203 & A200;
  assign \new_[28254]_  = ~A199 & \new_[28253]_ ;
  assign \new_[28255]_  = \new_[28254]_  & \new_[28249]_ ;
  assign \new_[28259]_  = A236 & ~A233;
  assign \new_[28260]_  = A232 & \new_[28259]_ ;
  assign \new_[28264]_  = A269 & A266;
  assign \new_[28265]_  = ~A265 & \new_[28264]_ ;
  assign \new_[28266]_  = \new_[28265]_  & \new_[28260]_ ;
  assign \new_[28270]_  = ~A166 & ~A167;
  assign \new_[28271]_  = ~A169 & \new_[28270]_ ;
  assign \new_[28275]_  = A203 & A200;
  assign \new_[28276]_  = ~A199 & \new_[28275]_ ;
  assign \new_[28277]_  = \new_[28276]_  & \new_[28271]_ ;
  assign \new_[28281]_  = A236 & ~A233;
  assign \new_[28282]_  = A232 & \new_[28281]_ ;
  assign \new_[28286]_  = A269 & ~A266;
  assign \new_[28287]_  = A265 & \new_[28286]_ ;
  assign \new_[28288]_  = \new_[28287]_  & \new_[28282]_ ;
  assign \new_[28292]_  = ~A166 & ~A167;
  assign \new_[28293]_  = ~A169 & \new_[28292]_ ;
  assign \new_[28297]_  = A203 & ~A200;
  assign \new_[28298]_  = A199 & \new_[28297]_ ;
  assign \new_[28299]_  = \new_[28298]_  & \new_[28293]_ ;
  assign \new_[28303]_  = A298 & A234;
  assign \new_[28304]_  = A232 & \new_[28303]_ ;
  assign \new_[28308]_  = ~A301 & ~A300;
  assign \new_[28309]_  = A299 & \new_[28308]_ ;
  assign \new_[28310]_  = \new_[28309]_  & \new_[28304]_ ;
  assign \new_[28314]_  = ~A166 & ~A167;
  assign \new_[28315]_  = ~A169 & \new_[28314]_ ;
  assign \new_[28319]_  = A203 & ~A200;
  assign \new_[28320]_  = A199 & \new_[28319]_ ;
  assign \new_[28321]_  = \new_[28320]_  & \new_[28315]_ ;
  assign \new_[28325]_  = A298 & A234;
  assign \new_[28326]_  = A233 & \new_[28325]_ ;
  assign \new_[28330]_  = ~A301 & ~A300;
  assign \new_[28331]_  = A299 & \new_[28330]_ ;
  assign \new_[28332]_  = \new_[28331]_  & \new_[28326]_ ;
  assign \new_[28336]_  = ~A166 & ~A167;
  assign \new_[28337]_  = ~A169 & \new_[28336]_ ;
  assign \new_[28341]_  = A203 & ~A200;
  assign \new_[28342]_  = A199 & \new_[28341]_ ;
  assign \new_[28343]_  = \new_[28342]_  & \new_[28337]_ ;
  assign \new_[28347]_  = A236 & A233;
  assign \new_[28348]_  = ~A232 & \new_[28347]_ ;
  assign \new_[28352]_  = ~A302 & ~A301;
  assign \new_[28353]_  = ~A300 & \new_[28352]_ ;
  assign \new_[28354]_  = \new_[28353]_  & \new_[28348]_ ;
  assign \new_[28358]_  = ~A166 & ~A167;
  assign \new_[28359]_  = ~A169 & \new_[28358]_ ;
  assign \new_[28363]_  = A203 & ~A200;
  assign \new_[28364]_  = A199 & \new_[28363]_ ;
  assign \new_[28365]_  = \new_[28364]_  & \new_[28359]_ ;
  assign \new_[28369]_  = A236 & A233;
  assign \new_[28370]_  = ~A232 & \new_[28369]_ ;
  assign \new_[28374]_  = ~A301 & ~A299;
  assign \new_[28375]_  = ~A298 & \new_[28374]_ ;
  assign \new_[28376]_  = \new_[28375]_  & \new_[28370]_ ;
  assign \new_[28380]_  = ~A166 & ~A167;
  assign \new_[28381]_  = ~A169 & \new_[28380]_ ;
  assign \new_[28385]_  = A203 & ~A200;
  assign \new_[28386]_  = A199 & \new_[28385]_ ;
  assign \new_[28387]_  = \new_[28386]_  & \new_[28381]_ ;
  assign \new_[28391]_  = A236 & A233;
  assign \new_[28392]_  = ~A232 & \new_[28391]_ ;
  assign \new_[28396]_  = A269 & A266;
  assign \new_[28397]_  = ~A265 & \new_[28396]_ ;
  assign \new_[28398]_  = \new_[28397]_  & \new_[28392]_ ;
  assign \new_[28402]_  = ~A166 & ~A167;
  assign \new_[28403]_  = ~A169 & \new_[28402]_ ;
  assign \new_[28407]_  = A203 & ~A200;
  assign \new_[28408]_  = A199 & \new_[28407]_ ;
  assign \new_[28409]_  = \new_[28408]_  & \new_[28403]_ ;
  assign \new_[28413]_  = A236 & A233;
  assign \new_[28414]_  = ~A232 & \new_[28413]_ ;
  assign \new_[28418]_  = A269 & ~A266;
  assign \new_[28419]_  = A265 & \new_[28418]_ ;
  assign \new_[28420]_  = \new_[28419]_  & \new_[28414]_ ;
  assign \new_[28424]_  = ~A166 & ~A167;
  assign \new_[28425]_  = ~A169 & \new_[28424]_ ;
  assign \new_[28429]_  = A203 & ~A200;
  assign \new_[28430]_  = A199 & \new_[28429]_ ;
  assign \new_[28431]_  = \new_[28430]_  & \new_[28425]_ ;
  assign \new_[28435]_  = A236 & ~A233;
  assign \new_[28436]_  = A232 & \new_[28435]_ ;
  assign \new_[28440]_  = ~A302 & ~A301;
  assign \new_[28441]_  = ~A300 & \new_[28440]_ ;
  assign \new_[28442]_  = \new_[28441]_  & \new_[28436]_ ;
  assign \new_[28446]_  = ~A166 & ~A167;
  assign \new_[28447]_  = ~A169 & \new_[28446]_ ;
  assign \new_[28451]_  = A203 & ~A200;
  assign \new_[28452]_  = A199 & \new_[28451]_ ;
  assign \new_[28453]_  = \new_[28452]_  & \new_[28447]_ ;
  assign \new_[28457]_  = A236 & ~A233;
  assign \new_[28458]_  = A232 & \new_[28457]_ ;
  assign \new_[28462]_  = ~A301 & ~A299;
  assign \new_[28463]_  = ~A298 & \new_[28462]_ ;
  assign \new_[28464]_  = \new_[28463]_  & \new_[28458]_ ;
  assign \new_[28468]_  = ~A166 & ~A167;
  assign \new_[28469]_  = ~A169 & \new_[28468]_ ;
  assign \new_[28473]_  = A203 & ~A200;
  assign \new_[28474]_  = A199 & \new_[28473]_ ;
  assign \new_[28475]_  = \new_[28474]_  & \new_[28469]_ ;
  assign \new_[28479]_  = A236 & ~A233;
  assign \new_[28480]_  = A232 & \new_[28479]_ ;
  assign \new_[28484]_  = A269 & A266;
  assign \new_[28485]_  = ~A265 & \new_[28484]_ ;
  assign \new_[28486]_  = \new_[28485]_  & \new_[28480]_ ;
  assign \new_[28490]_  = ~A166 & ~A167;
  assign \new_[28491]_  = ~A169 & \new_[28490]_ ;
  assign \new_[28495]_  = A203 & ~A200;
  assign \new_[28496]_  = A199 & \new_[28495]_ ;
  assign \new_[28497]_  = \new_[28496]_  & \new_[28491]_ ;
  assign \new_[28501]_  = A236 & ~A233;
  assign \new_[28502]_  = A232 & \new_[28501]_ ;
  assign \new_[28506]_  = A269 & ~A266;
  assign \new_[28507]_  = A265 & \new_[28506]_ ;
  assign \new_[28508]_  = \new_[28507]_  & \new_[28502]_ ;
  assign \new_[28512]_  = A167 & ~A168;
  assign \new_[28513]_  = ~A169 & \new_[28512]_ ;
  assign \new_[28517]_  = ~A234 & A202;
  assign \new_[28518]_  = A166 & \new_[28517]_ ;
  assign \new_[28519]_  = \new_[28518]_  & \new_[28513]_ ;
  assign \new_[28523]_  = ~A267 & ~A236;
  assign \new_[28524]_  = ~A235 & \new_[28523]_ ;
  assign \new_[28528]_  = A301 & ~A269;
  assign \new_[28529]_  = ~A268 & \new_[28528]_ ;
  assign \new_[28530]_  = \new_[28529]_  & \new_[28524]_ ;
  assign \new_[28534]_  = A167 & ~A168;
  assign \new_[28535]_  = ~A169 & \new_[28534]_ ;
  assign \new_[28539]_  = ~A234 & A202;
  assign \new_[28540]_  = A166 & \new_[28539]_ ;
  assign \new_[28541]_  = \new_[28540]_  & \new_[28535]_ ;
  assign \new_[28545]_  = ~A265 & ~A236;
  assign \new_[28546]_  = ~A235 & \new_[28545]_ ;
  assign \new_[28550]_  = A301 & ~A268;
  assign \new_[28551]_  = ~A266 & \new_[28550]_ ;
  assign \new_[28552]_  = \new_[28551]_  & \new_[28546]_ ;
  assign \new_[28556]_  = A167 & ~A168;
  assign \new_[28557]_  = ~A169 & \new_[28556]_ ;
  assign \new_[28561]_  = ~A232 & A202;
  assign \new_[28562]_  = A166 & \new_[28561]_ ;
  assign \new_[28563]_  = \new_[28562]_  & \new_[28557]_ ;
  assign \new_[28567]_  = A298 & A236;
  assign \new_[28568]_  = A233 & \new_[28567]_ ;
  assign \new_[28572]_  = ~A301 & ~A300;
  assign \new_[28573]_  = A299 & \new_[28572]_ ;
  assign \new_[28574]_  = \new_[28573]_  & \new_[28568]_ ;
  assign \new_[28578]_  = A167 & ~A168;
  assign \new_[28579]_  = ~A169 & \new_[28578]_ ;
  assign \new_[28583]_  = A232 & A202;
  assign \new_[28584]_  = A166 & \new_[28583]_ ;
  assign \new_[28585]_  = \new_[28584]_  & \new_[28579]_ ;
  assign \new_[28589]_  = A298 & A236;
  assign \new_[28590]_  = ~A233 & \new_[28589]_ ;
  assign \new_[28594]_  = ~A301 & ~A300;
  assign \new_[28595]_  = A299 & \new_[28594]_ ;
  assign \new_[28596]_  = \new_[28595]_  & \new_[28590]_ ;
  assign \new_[28600]_  = A167 & ~A168;
  assign \new_[28601]_  = ~A169 & \new_[28600]_ ;
  assign \new_[28605]_  = ~A232 & A202;
  assign \new_[28606]_  = A166 & \new_[28605]_ ;
  assign \new_[28607]_  = \new_[28606]_  & \new_[28601]_ ;
  assign \new_[28611]_  = ~A267 & ~A235;
  assign \new_[28612]_  = ~A233 & \new_[28611]_ ;
  assign \new_[28616]_  = A301 & ~A269;
  assign \new_[28617]_  = ~A268 & \new_[28616]_ ;
  assign \new_[28618]_  = \new_[28617]_  & \new_[28612]_ ;
  assign \new_[28622]_  = A167 & ~A168;
  assign \new_[28623]_  = ~A169 & \new_[28622]_ ;
  assign \new_[28627]_  = ~A232 & A202;
  assign \new_[28628]_  = A166 & \new_[28627]_ ;
  assign \new_[28629]_  = \new_[28628]_  & \new_[28623]_ ;
  assign \new_[28633]_  = ~A265 & ~A235;
  assign \new_[28634]_  = ~A233 & \new_[28633]_ ;
  assign \new_[28638]_  = A301 & ~A268;
  assign \new_[28639]_  = ~A266 & \new_[28638]_ ;
  assign \new_[28640]_  = \new_[28639]_  & \new_[28634]_ ;
  assign \new_[28644]_  = A167 & ~A168;
  assign \new_[28645]_  = ~A169 & \new_[28644]_ ;
  assign \new_[28649]_  = A201 & A199;
  assign \new_[28650]_  = A166 & \new_[28649]_ ;
  assign \new_[28651]_  = \new_[28650]_  & \new_[28645]_ ;
  assign \new_[28655]_  = A298 & A234;
  assign \new_[28656]_  = A232 & \new_[28655]_ ;
  assign \new_[28660]_  = ~A301 & ~A300;
  assign \new_[28661]_  = A299 & \new_[28660]_ ;
  assign \new_[28662]_  = \new_[28661]_  & \new_[28656]_ ;
  assign \new_[28666]_  = A167 & ~A168;
  assign \new_[28667]_  = ~A169 & \new_[28666]_ ;
  assign \new_[28671]_  = A201 & A199;
  assign \new_[28672]_  = A166 & \new_[28671]_ ;
  assign \new_[28673]_  = \new_[28672]_  & \new_[28667]_ ;
  assign \new_[28677]_  = A298 & A234;
  assign \new_[28678]_  = A233 & \new_[28677]_ ;
  assign \new_[28682]_  = ~A301 & ~A300;
  assign \new_[28683]_  = A299 & \new_[28682]_ ;
  assign \new_[28684]_  = \new_[28683]_  & \new_[28678]_ ;
  assign \new_[28688]_  = A167 & ~A168;
  assign \new_[28689]_  = ~A169 & \new_[28688]_ ;
  assign \new_[28693]_  = A201 & A199;
  assign \new_[28694]_  = A166 & \new_[28693]_ ;
  assign \new_[28695]_  = \new_[28694]_  & \new_[28689]_ ;
  assign \new_[28699]_  = A236 & A233;
  assign \new_[28700]_  = ~A232 & \new_[28699]_ ;
  assign \new_[28704]_  = ~A302 & ~A301;
  assign \new_[28705]_  = ~A300 & \new_[28704]_ ;
  assign \new_[28706]_  = \new_[28705]_  & \new_[28700]_ ;
  assign \new_[28710]_  = A167 & ~A168;
  assign \new_[28711]_  = ~A169 & \new_[28710]_ ;
  assign \new_[28715]_  = A201 & A199;
  assign \new_[28716]_  = A166 & \new_[28715]_ ;
  assign \new_[28717]_  = \new_[28716]_  & \new_[28711]_ ;
  assign \new_[28721]_  = A236 & A233;
  assign \new_[28722]_  = ~A232 & \new_[28721]_ ;
  assign \new_[28726]_  = ~A301 & ~A299;
  assign \new_[28727]_  = ~A298 & \new_[28726]_ ;
  assign \new_[28728]_  = \new_[28727]_  & \new_[28722]_ ;
  assign \new_[28732]_  = A167 & ~A168;
  assign \new_[28733]_  = ~A169 & \new_[28732]_ ;
  assign \new_[28737]_  = A201 & A199;
  assign \new_[28738]_  = A166 & \new_[28737]_ ;
  assign \new_[28739]_  = \new_[28738]_  & \new_[28733]_ ;
  assign \new_[28743]_  = A236 & A233;
  assign \new_[28744]_  = ~A232 & \new_[28743]_ ;
  assign \new_[28748]_  = A269 & A266;
  assign \new_[28749]_  = ~A265 & \new_[28748]_ ;
  assign \new_[28750]_  = \new_[28749]_  & \new_[28744]_ ;
  assign \new_[28754]_  = A167 & ~A168;
  assign \new_[28755]_  = ~A169 & \new_[28754]_ ;
  assign \new_[28759]_  = A201 & A199;
  assign \new_[28760]_  = A166 & \new_[28759]_ ;
  assign \new_[28761]_  = \new_[28760]_  & \new_[28755]_ ;
  assign \new_[28765]_  = A236 & A233;
  assign \new_[28766]_  = ~A232 & \new_[28765]_ ;
  assign \new_[28770]_  = A269 & ~A266;
  assign \new_[28771]_  = A265 & \new_[28770]_ ;
  assign \new_[28772]_  = \new_[28771]_  & \new_[28766]_ ;
  assign \new_[28776]_  = A167 & ~A168;
  assign \new_[28777]_  = ~A169 & \new_[28776]_ ;
  assign \new_[28781]_  = A201 & A199;
  assign \new_[28782]_  = A166 & \new_[28781]_ ;
  assign \new_[28783]_  = \new_[28782]_  & \new_[28777]_ ;
  assign \new_[28787]_  = A236 & ~A233;
  assign \new_[28788]_  = A232 & \new_[28787]_ ;
  assign \new_[28792]_  = ~A302 & ~A301;
  assign \new_[28793]_  = ~A300 & \new_[28792]_ ;
  assign \new_[28794]_  = \new_[28793]_  & \new_[28788]_ ;
  assign \new_[28798]_  = A167 & ~A168;
  assign \new_[28799]_  = ~A169 & \new_[28798]_ ;
  assign \new_[28803]_  = A201 & A199;
  assign \new_[28804]_  = A166 & \new_[28803]_ ;
  assign \new_[28805]_  = \new_[28804]_  & \new_[28799]_ ;
  assign \new_[28809]_  = A236 & ~A233;
  assign \new_[28810]_  = A232 & \new_[28809]_ ;
  assign \new_[28814]_  = ~A301 & ~A299;
  assign \new_[28815]_  = ~A298 & \new_[28814]_ ;
  assign \new_[28816]_  = \new_[28815]_  & \new_[28810]_ ;
  assign \new_[28820]_  = A167 & ~A168;
  assign \new_[28821]_  = ~A169 & \new_[28820]_ ;
  assign \new_[28825]_  = A201 & A199;
  assign \new_[28826]_  = A166 & \new_[28825]_ ;
  assign \new_[28827]_  = \new_[28826]_  & \new_[28821]_ ;
  assign \new_[28831]_  = A236 & ~A233;
  assign \new_[28832]_  = A232 & \new_[28831]_ ;
  assign \new_[28836]_  = A269 & A266;
  assign \new_[28837]_  = ~A265 & \new_[28836]_ ;
  assign \new_[28838]_  = \new_[28837]_  & \new_[28832]_ ;
  assign \new_[28842]_  = A167 & ~A168;
  assign \new_[28843]_  = ~A169 & \new_[28842]_ ;
  assign \new_[28847]_  = A201 & A199;
  assign \new_[28848]_  = A166 & \new_[28847]_ ;
  assign \new_[28849]_  = \new_[28848]_  & \new_[28843]_ ;
  assign \new_[28853]_  = A236 & ~A233;
  assign \new_[28854]_  = A232 & \new_[28853]_ ;
  assign \new_[28858]_  = A269 & ~A266;
  assign \new_[28859]_  = A265 & \new_[28858]_ ;
  assign \new_[28860]_  = \new_[28859]_  & \new_[28854]_ ;
  assign \new_[28864]_  = A167 & ~A168;
  assign \new_[28865]_  = ~A169 & \new_[28864]_ ;
  assign \new_[28869]_  = A201 & A200;
  assign \new_[28870]_  = A166 & \new_[28869]_ ;
  assign \new_[28871]_  = \new_[28870]_  & \new_[28865]_ ;
  assign \new_[28875]_  = A298 & A234;
  assign \new_[28876]_  = A232 & \new_[28875]_ ;
  assign \new_[28880]_  = ~A301 & ~A300;
  assign \new_[28881]_  = A299 & \new_[28880]_ ;
  assign \new_[28882]_  = \new_[28881]_  & \new_[28876]_ ;
  assign \new_[28886]_  = A167 & ~A168;
  assign \new_[28887]_  = ~A169 & \new_[28886]_ ;
  assign \new_[28891]_  = A201 & A200;
  assign \new_[28892]_  = A166 & \new_[28891]_ ;
  assign \new_[28893]_  = \new_[28892]_  & \new_[28887]_ ;
  assign \new_[28897]_  = A298 & A234;
  assign \new_[28898]_  = A233 & \new_[28897]_ ;
  assign \new_[28902]_  = ~A301 & ~A300;
  assign \new_[28903]_  = A299 & \new_[28902]_ ;
  assign \new_[28904]_  = \new_[28903]_  & \new_[28898]_ ;
  assign \new_[28908]_  = A167 & ~A168;
  assign \new_[28909]_  = ~A169 & \new_[28908]_ ;
  assign \new_[28913]_  = A201 & A200;
  assign \new_[28914]_  = A166 & \new_[28913]_ ;
  assign \new_[28915]_  = \new_[28914]_  & \new_[28909]_ ;
  assign \new_[28919]_  = A236 & A233;
  assign \new_[28920]_  = ~A232 & \new_[28919]_ ;
  assign \new_[28924]_  = ~A302 & ~A301;
  assign \new_[28925]_  = ~A300 & \new_[28924]_ ;
  assign \new_[28926]_  = \new_[28925]_  & \new_[28920]_ ;
  assign \new_[28930]_  = A167 & ~A168;
  assign \new_[28931]_  = ~A169 & \new_[28930]_ ;
  assign \new_[28935]_  = A201 & A200;
  assign \new_[28936]_  = A166 & \new_[28935]_ ;
  assign \new_[28937]_  = \new_[28936]_  & \new_[28931]_ ;
  assign \new_[28941]_  = A236 & A233;
  assign \new_[28942]_  = ~A232 & \new_[28941]_ ;
  assign \new_[28946]_  = ~A301 & ~A299;
  assign \new_[28947]_  = ~A298 & \new_[28946]_ ;
  assign \new_[28948]_  = \new_[28947]_  & \new_[28942]_ ;
  assign \new_[28952]_  = A167 & ~A168;
  assign \new_[28953]_  = ~A169 & \new_[28952]_ ;
  assign \new_[28957]_  = A201 & A200;
  assign \new_[28958]_  = A166 & \new_[28957]_ ;
  assign \new_[28959]_  = \new_[28958]_  & \new_[28953]_ ;
  assign \new_[28963]_  = A236 & A233;
  assign \new_[28964]_  = ~A232 & \new_[28963]_ ;
  assign \new_[28968]_  = A269 & A266;
  assign \new_[28969]_  = ~A265 & \new_[28968]_ ;
  assign \new_[28970]_  = \new_[28969]_  & \new_[28964]_ ;
  assign \new_[28974]_  = A167 & ~A168;
  assign \new_[28975]_  = ~A169 & \new_[28974]_ ;
  assign \new_[28979]_  = A201 & A200;
  assign \new_[28980]_  = A166 & \new_[28979]_ ;
  assign \new_[28981]_  = \new_[28980]_  & \new_[28975]_ ;
  assign \new_[28985]_  = A236 & A233;
  assign \new_[28986]_  = ~A232 & \new_[28985]_ ;
  assign \new_[28990]_  = A269 & ~A266;
  assign \new_[28991]_  = A265 & \new_[28990]_ ;
  assign \new_[28992]_  = \new_[28991]_  & \new_[28986]_ ;
  assign \new_[28996]_  = A167 & ~A168;
  assign \new_[28997]_  = ~A169 & \new_[28996]_ ;
  assign \new_[29001]_  = A201 & A200;
  assign \new_[29002]_  = A166 & \new_[29001]_ ;
  assign \new_[29003]_  = \new_[29002]_  & \new_[28997]_ ;
  assign \new_[29007]_  = A236 & ~A233;
  assign \new_[29008]_  = A232 & \new_[29007]_ ;
  assign \new_[29012]_  = ~A302 & ~A301;
  assign \new_[29013]_  = ~A300 & \new_[29012]_ ;
  assign \new_[29014]_  = \new_[29013]_  & \new_[29008]_ ;
  assign \new_[29018]_  = A167 & ~A168;
  assign \new_[29019]_  = ~A169 & \new_[29018]_ ;
  assign \new_[29023]_  = A201 & A200;
  assign \new_[29024]_  = A166 & \new_[29023]_ ;
  assign \new_[29025]_  = \new_[29024]_  & \new_[29019]_ ;
  assign \new_[29029]_  = A236 & ~A233;
  assign \new_[29030]_  = A232 & \new_[29029]_ ;
  assign \new_[29034]_  = ~A301 & ~A299;
  assign \new_[29035]_  = ~A298 & \new_[29034]_ ;
  assign \new_[29036]_  = \new_[29035]_  & \new_[29030]_ ;
  assign \new_[29040]_  = A167 & ~A168;
  assign \new_[29041]_  = ~A169 & \new_[29040]_ ;
  assign \new_[29045]_  = A201 & A200;
  assign \new_[29046]_  = A166 & \new_[29045]_ ;
  assign \new_[29047]_  = \new_[29046]_  & \new_[29041]_ ;
  assign \new_[29051]_  = A236 & ~A233;
  assign \new_[29052]_  = A232 & \new_[29051]_ ;
  assign \new_[29056]_  = A269 & A266;
  assign \new_[29057]_  = ~A265 & \new_[29056]_ ;
  assign \new_[29058]_  = \new_[29057]_  & \new_[29052]_ ;
  assign \new_[29062]_  = A167 & ~A168;
  assign \new_[29063]_  = ~A169 & \new_[29062]_ ;
  assign \new_[29067]_  = A201 & A200;
  assign \new_[29068]_  = A166 & \new_[29067]_ ;
  assign \new_[29069]_  = \new_[29068]_  & \new_[29063]_ ;
  assign \new_[29073]_  = A236 & ~A233;
  assign \new_[29074]_  = A232 & \new_[29073]_ ;
  assign \new_[29078]_  = A269 & ~A266;
  assign \new_[29079]_  = A265 & \new_[29078]_ ;
  assign \new_[29080]_  = \new_[29079]_  & \new_[29074]_ ;
  assign \new_[29084]_  = A167 & ~A168;
  assign \new_[29085]_  = ~A169 & \new_[29084]_ ;
  assign \new_[29089]_  = A200 & ~A199;
  assign \new_[29090]_  = A166 & \new_[29089]_ ;
  assign \new_[29091]_  = \new_[29090]_  & \new_[29085]_ ;
  assign \new_[29095]_  = A298 & A235;
  assign \new_[29096]_  = A203 & \new_[29095]_ ;
  assign \new_[29100]_  = ~A301 & ~A300;
  assign \new_[29101]_  = A299 & \new_[29100]_ ;
  assign \new_[29102]_  = \new_[29101]_  & \new_[29096]_ ;
  assign \new_[29106]_  = A167 & ~A168;
  assign \new_[29107]_  = ~A169 & \new_[29106]_ ;
  assign \new_[29111]_  = A200 & ~A199;
  assign \new_[29112]_  = A166 & \new_[29111]_ ;
  assign \new_[29113]_  = \new_[29112]_  & \new_[29107]_ ;
  assign \new_[29117]_  = A234 & A232;
  assign \new_[29118]_  = A203 & \new_[29117]_ ;
  assign \new_[29122]_  = ~A302 & ~A301;
  assign \new_[29123]_  = ~A300 & \new_[29122]_ ;
  assign \new_[29124]_  = \new_[29123]_  & \new_[29118]_ ;
  assign \new_[29128]_  = A167 & ~A168;
  assign \new_[29129]_  = ~A169 & \new_[29128]_ ;
  assign \new_[29133]_  = A200 & ~A199;
  assign \new_[29134]_  = A166 & \new_[29133]_ ;
  assign \new_[29135]_  = \new_[29134]_  & \new_[29129]_ ;
  assign \new_[29139]_  = A234 & A232;
  assign \new_[29140]_  = A203 & \new_[29139]_ ;
  assign \new_[29144]_  = ~A301 & ~A299;
  assign \new_[29145]_  = ~A298 & \new_[29144]_ ;
  assign \new_[29146]_  = \new_[29145]_  & \new_[29140]_ ;
  assign \new_[29150]_  = A167 & ~A168;
  assign \new_[29151]_  = ~A169 & \new_[29150]_ ;
  assign \new_[29155]_  = A200 & ~A199;
  assign \new_[29156]_  = A166 & \new_[29155]_ ;
  assign \new_[29157]_  = \new_[29156]_  & \new_[29151]_ ;
  assign \new_[29161]_  = A234 & A232;
  assign \new_[29162]_  = A203 & \new_[29161]_ ;
  assign \new_[29166]_  = A269 & A266;
  assign \new_[29167]_  = ~A265 & \new_[29166]_ ;
  assign \new_[29168]_  = \new_[29167]_  & \new_[29162]_ ;
  assign \new_[29172]_  = A167 & ~A168;
  assign \new_[29173]_  = ~A169 & \new_[29172]_ ;
  assign \new_[29177]_  = A200 & ~A199;
  assign \new_[29178]_  = A166 & \new_[29177]_ ;
  assign \new_[29179]_  = \new_[29178]_  & \new_[29173]_ ;
  assign \new_[29183]_  = A234 & A232;
  assign \new_[29184]_  = A203 & \new_[29183]_ ;
  assign \new_[29188]_  = A269 & ~A266;
  assign \new_[29189]_  = A265 & \new_[29188]_ ;
  assign \new_[29190]_  = \new_[29189]_  & \new_[29184]_ ;
  assign \new_[29194]_  = A167 & ~A168;
  assign \new_[29195]_  = ~A169 & \new_[29194]_ ;
  assign \new_[29199]_  = A200 & ~A199;
  assign \new_[29200]_  = A166 & \new_[29199]_ ;
  assign \new_[29201]_  = \new_[29200]_  & \new_[29195]_ ;
  assign \new_[29205]_  = A234 & A233;
  assign \new_[29206]_  = A203 & \new_[29205]_ ;
  assign \new_[29210]_  = ~A302 & ~A301;
  assign \new_[29211]_  = ~A300 & \new_[29210]_ ;
  assign \new_[29212]_  = \new_[29211]_  & \new_[29206]_ ;
  assign \new_[29216]_  = A167 & ~A168;
  assign \new_[29217]_  = ~A169 & \new_[29216]_ ;
  assign \new_[29221]_  = A200 & ~A199;
  assign \new_[29222]_  = A166 & \new_[29221]_ ;
  assign \new_[29223]_  = \new_[29222]_  & \new_[29217]_ ;
  assign \new_[29227]_  = A234 & A233;
  assign \new_[29228]_  = A203 & \new_[29227]_ ;
  assign \new_[29232]_  = ~A301 & ~A299;
  assign \new_[29233]_  = ~A298 & \new_[29232]_ ;
  assign \new_[29234]_  = \new_[29233]_  & \new_[29228]_ ;
  assign \new_[29238]_  = A167 & ~A168;
  assign \new_[29239]_  = ~A169 & \new_[29238]_ ;
  assign \new_[29243]_  = A200 & ~A199;
  assign \new_[29244]_  = A166 & \new_[29243]_ ;
  assign \new_[29245]_  = \new_[29244]_  & \new_[29239]_ ;
  assign \new_[29249]_  = A234 & A233;
  assign \new_[29250]_  = A203 & \new_[29249]_ ;
  assign \new_[29254]_  = A269 & A266;
  assign \new_[29255]_  = ~A265 & \new_[29254]_ ;
  assign \new_[29256]_  = \new_[29255]_  & \new_[29250]_ ;
  assign \new_[29260]_  = A167 & ~A168;
  assign \new_[29261]_  = ~A169 & \new_[29260]_ ;
  assign \new_[29265]_  = A200 & ~A199;
  assign \new_[29266]_  = A166 & \new_[29265]_ ;
  assign \new_[29267]_  = \new_[29266]_  & \new_[29261]_ ;
  assign \new_[29271]_  = A234 & A233;
  assign \new_[29272]_  = A203 & \new_[29271]_ ;
  assign \new_[29276]_  = A269 & ~A266;
  assign \new_[29277]_  = A265 & \new_[29276]_ ;
  assign \new_[29278]_  = \new_[29277]_  & \new_[29272]_ ;
  assign \new_[29282]_  = A167 & ~A168;
  assign \new_[29283]_  = ~A169 & \new_[29282]_ ;
  assign \new_[29287]_  = A200 & ~A199;
  assign \new_[29288]_  = A166 & \new_[29287]_ ;
  assign \new_[29289]_  = \new_[29288]_  & \new_[29283]_ ;
  assign \new_[29293]_  = A233 & ~A232;
  assign \new_[29294]_  = A203 & \new_[29293]_ ;
  assign \new_[29298]_  = A267 & A265;
  assign \new_[29299]_  = A236 & \new_[29298]_ ;
  assign \new_[29300]_  = \new_[29299]_  & \new_[29294]_ ;
  assign \new_[29304]_  = A167 & ~A168;
  assign \new_[29305]_  = ~A169 & \new_[29304]_ ;
  assign \new_[29309]_  = A200 & ~A199;
  assign \new_[29310]_  = A166 & \new_[29309]_ ;
  assign \new_[29311]_  = \new_[29310]_  & \new_[29305]_ ;
  assign \new_[29315]_  = A233 & ~A232;
  assign \new_[29316]_  = A203 & \new_[29315]_ ;
  assign \new_[29320]_  = A267 & A266;
  assign \new_[29321]_  = A236 & \new_[29320]_ ;
  assign \new_[29322]_  = \new_[29321]_  & \new_[29316]_ ;
  assign \new_[29326]_  = A167 & ~A168;
  assign \new_[29327]_  = ~A169 & \new_[29326]_ ;
  assign \new_[29331]_  = A200 & ~A199;
  assign \new_[29332]_  = A166 & \new_[29331]_ ;
  assign \new_[29333]_  = \new_[29332]_  & \new_[29327]_ ;
  assign \new_[29337]_  = ~A233 & A232;
  assign \new_[29338]_  = A203 & \new_[29337]_ ;
  assign \new_[29342]_  = A267 & A265;
  assign \new_[29343]_  = A236 & \new_[29342]_ ;
  assign \new_[29344]_  = \new_[29343]_  & \new_[29338]_ ;
  assign \new_[29348]_  = A167 & ~A168;
  assign \new_[29349]_  = ~A169 & \new_[29348]_ ;
  assign \new_[29353]_  = A200 & ~A199;
  assign \new_[29354]_  = A166 & \new_[29353]_ ;
  assign \new_[29355]_  = \new_[29354]_  & \new_[29349]_ ;
  assign \new_[29359]_  = ~A233 & A232;
  assign \new_[29360]_  = A203 & \new_[29359]_ ;
  assign \new_[29364]_  = A267 & A266;
  assign \new_[29365]_  = A236 & \new_[29364]_ ;
  assign \new_[29366]_  = \new_[29365]_  & \new_[29360]_ ;
  assign \new_[29370]_  = A167 & ~A168;
  assign \new_[29371]_  = ~A169 & \new_[29370]_ ;
  assign \new_[29375]_  = ~A200 & A199;
  assign \new_[29376]_  = A166 & \new_[29375]_ ;
  assign \new_[29377]_  = \new_[29376]_  & \new_[29371]_ ;
  assign \new_[29381]_  = A298 & A235;
  assign \new_[29382]_  = A203 & \new_[29381]_ ;
  assign \new_[29386]_  = ~A301 & ~A300;
  assign \new_[29387]_  = A299 & \new_[29386]_ ;
  assign \new_[29388]_  = \new_[29387]_  & \new_[29382]_ ;
  assign \new_[29392]_  = A167 & ~A168;
  assign \new_[29393]_  = ~A169 & \new_[29392]_ ;
  assign \new_[29397]_  = ~A200 & A199;
  assign \new_[29398]_  = A166 & \new_[29397]_ ;
  assign \new_[29399]_  = \new_[29398]_  & \new_[29393]_ ;
  assign \new_[29403]_  = A234 & A232;
  assign \new_[29404]_  = A203 & \new_[29403]_ ;
  assign \new_[29408]_  = ~A302 & ~A301;
  assign \new_[29409]_  = ~A300 & \new_[29408]_ ;
  assign \new_[29410]_  = \new_[29409]_  & \new_[29404]_ ;
  assign \new_[29414]_  = A167 & ~A168;
  assign \new_[29415]_  = ~A169 & \new_[29414]_ ;
  assign \new_[29419]_  = ~A200 & A199;
  assign \new_[29420]_  = A166 & \new_[29419]_ ;
  assign \new_[29421]_  = \new_[29420]_  & \new_[29415]_ ;
  assign \new_[29425]_  = A234 & A232;
  assign \new_[29426]_  = A203 & \new_[29425]_ ;
  assign \new_[29430]_  = ~A301 & ~A299;
  assign \new_[29431]_  = ~A298 & \new_[29430]_ ;
  assign \new_[29432]_  = \new_[29431]_  & \new_[29426]_ ;
  assign \new_[29436]_  = A167 & ~A168;
  assign \new_[29437]_  = ~A169 & \new_[29436]_ ;
  assign \new_[29441]_  = ~A200 & A199;
  assign \new_[29442]_  = A166 & \new_[29441]_ ;
  assign \new_[29443]_  = \new_[29442]_  & \new_[29437]_ ;
  assign \new_[29447]_  = A234 & A232;
  assign \new_[29448]_  = A203 & \new_[29447]_ ;
  assign \new_[29452]_  = A269 & A266;
  assign \new_[29453]_  = ~A265 & \new_[29452]_ ;
  assign \new_[29454]_  = \new_[29453]_  & \new_[29448]_ ;
  assign \new_[29458]_  = A167 & ~A168;
  assign \new_[29459]_  = ~A169 & \new_[29458]_ ;
  assign \new_[29463]_  = ~A200 & A199;
  assign \new_[29464]_  = A166 & \new_[29463]_ ;
  assign \new_[29465]_  = \new_[29464]_  & \new_[29459]_ ;
  assign \new_[29469]_  = A234 & A232;
  assign \new_[29470]_  = A203 & \new_[29469]_ ;
  assign \new_[29474]_  = A269 & ~A266;
  assign \new_[29475]_  = A265 & \new_[29474]_ ;
  assign \new_[29476]_  = \new_[29475]_  & \new_[29470]_ ;
  assign \new_[29480]_  = A167 & ~A168;
  assign \new_[29481]_  = ~A169 & \new_[29480]_ ;
  assign \new_[29485]_  = ~A200 & A199;
  assign \new_[29486]_  = A166 & \new_[29485]_ ;
  assign \new_[29487]_  = \new_[29486]_  & \new_[29481]_ ;
  assign \new_[29491]_  = A234 & A233;
  assign \new_[29492]_  = A203 & \new_[29491]_ ;
  assign \new_[29496]_  = ~A302 & ~A301;
  assign \new_[29497]_  = ~A300 & \new_[29496]_ ;
  assign \new_[29498]_  = \new_[29497]_  & \new_[29492]_ ;
  assign \new_[29502]_  = A167 & ~A168;
  assign \new_[29503]_  = ~A169 & \new_[29502]_ ;
  assign \new_[29507]_  = ~A200 & A199;
  assign \new_[29508]_  = A166 & \new_[29507]_ ;
  assign \new_[29509]_  = \new_[29508]_  & \new_[29503]_ ;
  assign \new_[29513]_  = A234 & A233;
  assign \new_[29514]_  = A203 & \new_[29513]_ ;
  assign \new_[29518]_  = ~A301 & ~A299;
  assign \new_[29519]_  = ~A298 & \new_[29518]_ ;
  assign \new_[29520]_  = \new_[29519]_  & \new_[29514]_ ;
  assign \new_[29524]_  = A167 & ~A168;
  assign \new_[29525]_  = ~A169 & \new_[29524]_ ;
  assign \new_[29529]_  = ~A200 & A199;
  assign \new_[29530]_  = A166 & \new_[29529]_ ;
  assign \new_[29531]_  = \new_[29530]_  & \new_[29525]_ ;
  assign \new_[29535]_  = A234 & A233;
  assign \new_[29536]_  = A203 & \new_[29535]_ ;
  assign \new_[29540]_  = A269 & A266;
  assign \new_[29541]_  = ~A265 & \new_[29540]_ ;
  assign \new_[29542]_  = \new_[29541]_  & \new_[29536]_ ;
  assign \new_[29546]_  = A167 & ~A168;
  assign \new_[29547]_  = ~A169 & \new_[29546]_ ;
  assign \new_[29551]_  = ~A200 & A199;
  assign \new_[29552]_  = A166 & \new_[29551]_ ;
  assign \new_[29553]_  = \new_[29552]_  & \new_[29547]_ ;
  assign \new_[29557]_  = A234 & A233;
  assign \new_[29558]_  = A203 & \new_[29557]_ ;
  assign \new_[29562]_  = A269 & ~A266;
  assign \new_[29563]_  = A265 & \new_[29562]_ ;
  assign \new_[29564]_  = \new_[29563]_  & \new_[29558]_ ;
  assign \new_[29568]_  = A167 & ~A168;
  assign \new_[29569]_  = ~A169 & \new_[29568]_ ;
  assign \new_[29573]_  = ~A200 & A199;
  assign \new_[29574]_  = A166 & \new_[29573]_ ;
  assign \new_[29575]_  = \new_[29574]_  & \new_[29569]_ ;
  assign \new_[29579]_  = A233 & ~A232;
  assign \new_[29580]_  = A203 & \new_[29579]_ ;
  assign \new_[29584]_  = A267 & A265;
  assign \new_[29585]_  = A236 & \new_[29584]_ ;
  assign \new_[29586]_  = \new_[29585]_  & \new_[29580]_ ;
  assign \new_[29590]_  = A167 & ~A168;
  assign \new_[29591]_  = ~A169 & \new_[29590]_ ;
  assign \new_[29595]_  = ~A200 & A199;
  assign \new_[29596]_  = A166 & \new_[29595]_ ;
  assign \new_[29597]_  = \new_[29596]_  & \new_[29591]_ ;
  assign \new_[29601]_  = A233 & ~A232;
  assign \new_[29602]_  = A203 & \new_[29601]_ ;
  assign \new_[29606]_  = A267 & A266;
  assign \new_[29607]_  = A236 & \new_[29606]_ ;
  assign \new_[29608]_  = \new_[29607]_  & \new_[29602]_ ;
  assign \new_[29612]_  = A167 & ~A168;
  assign \new_[29613]_  = ~A169 & \new_[29612]_ ;
  assign \new_[29617]_  = ~A200 & A199;
  assign \new_[29618]_  = A166 & \new_[29617]_ ;
  assign \new_[29619]_  = \new_[29618]_  & \new_[29613]_ ;
  assign \new_[29623]_  = ~A233 & A232;
  assign \new_[29624]_  = A203 & \new_[29623]_ ;
  assign \new_[29628]_  = A267 & A265;
  assign \new_[29629]_  = A236 & \new_[29628]_ ;
  assign \new_[29630]_  = \new_[29629]_  & \new_[29624]_ ;
  assign \new_[29634]_  = A167 & ~A168;
  assign \new_[29635]_  = ~A169 & \new_[29634]_ ;
  assign \new_[29639]_  = ~A200 & A199;
  assign \new_[29640]_  = A166 & \new_[29639]_ ;
  assign \new_[29641]_  = \new_[29640]_  & \new_[29635]_ ;
  assign \new_[29645]_  = ~A233 & A232;
  assign \new_[29646]_  = A203 & \new_[29645]_ ;
  assign \new_[29650]_  = A267 & A266;
  assign \new_[29651]_  = A236 & \new_[29650]_ ;
  assign \new_[29652]_  = \new_[29651]_  & \new_[29646]_ ;
  assign \new_[29656]_  = ~A168 & ~A169;
  assign \new_[29657]_  = ~A170 & \new_[29656]_ ;
  assign \new_[29661]_  = ~A235 & ~A234;
  assign \new_[29662]_  = A202 & \new_[29661]_ ;
  assign \new_[29663]_  = \new_[29662]_  & \new_[29657]_ ;
  assign \new_[29667]_  = ~A268 & ~A267;
  assign \new_[29668]_  = ~A236 & \new_[29667]_ ;
  assign \new_[29672]_  = A300 & A299;
  assign \new_[29673]_  = ~A269 & \new_[29672]_ ;
  assign \new_[29674]_  = \new_[29673]_  & \new_[29668]_ ;
  assign \new_[29678]_  = ~A168 & ~A169;
  assign \new_[29679]_  = ~A170 & \new_[29678]_ ;
  assign \new_[29683]_  = ~A235 & ~A234;
  assign \new_[29684]_  = A202 & \new_[29683]_ ;
  assign \new_[29685]_  = \new_[29684]_  & \new_[29679]_ ;
  assign \new_[29689]_  = ~A268 & ~A267;
  assign \new_[29690]_  = ~A236 & \new_[29689]_ ;
  assign \new_[29694]_  = A300 & A298;
  assign \new_[29695]_  = ~A269 & \new_[29694]_ ;
  assign \new_[29696]_  = \new_[29695]_  & \new_[29690]_ ;
  assign \new_[29700]_  = ~A168 & ~A169;
  assign \new_[29701]_  = ~A170 & \new_[29700]_ ;
  assign \new_[29705]_  = ~A235 & ~A234;
  assign \new_[29706]_  = A202 & \new_[29705]_ ;
  assign \new_[29707]_  = \new_[29706]_  & \new_[29701]_ ;
  assign \new_[29711]_  = A266 & A265;
  assign \new_[29712]_  = ~A236 & \new_[29711]_ ;
  assign \new_[29716]_  = A301 & ~A268;
  assign \new_[29717]_  = ~A267 & \new_[29716]_ ;
  assign \new_[29718]_  = \new_[29717]_  & \new_[29712]_ ;
  assign \new_[29722]_  = ~A168 & ~A169;
  assign \new_[29723]_  = ~A170 & \new_[29722]_ ;
  assign \new_[29727]_  = ~A235 & ~A234;
  assign \new_[29728]_  = A202 & \new_[29727]_ ;
  assign \new_[29729]_  = \new_[29728]_  & \new_[29723]_ ;
  assign \new_[29733]_  = ~A266 & ~A265;
  assign \new_[29734]_  = ~A236 & \new_[29733]_ ;
  assign \new_[29738]_  = A300 & A299;
  assign \new_[29739]_  = ~A268 & \new_[29738]_ ;
  assign \new_[29740]_  = \new_[29739]_  & \new_[29734]_ ;
  assign \new_[29744]_  = ~A168 & ~A169;
  assign \new_[29745]_  = ~A170 & \new_[29744]_ ;
  assign \new_[29749]_  = ~A235 & ~A234;
  assign \new_[29750]_  = A202 & \new_[29749]_ ;
  assign \new_[29751]_  = \new_[29750]_  & \new_[29745]_ ;
  assign \new_[29755]_  = ~A266 & ~A265;
  assign \new_[29756]_  = ~A236 & \new_[29755]_ ;
  assign \new_[29760]_  = A300 & A298;
  assign \new_[29761]_  = ~A268 & \new_[29760]_ ;
  assign \new_[29762]_  = \new_[29761]_  & \new_[29756]_ ;
  assign \new_[29766]_  = ~A168 & ~A169;
  assign \new_[29767]_  = ~A170 & \new_[29766]_ ;
  assign \new_[29771]_  = A233 & A232;
  assign \new_[29772]_  = A202 & \new_[29771]_ ;
  assign \new_[29773]_  = \new_[29772]_  & \new_[29767]_ ;
  assign \new_[29777]_  = ~A267 & ~A235;
  assign \new_[29778]_  = ~A234 & \new_[29777]_ ;
  assign \new_[29782]_  = A301 & ~A269;
  assign \new_[29783]_  = ~A268 & \new_[29782]_ ;
  assign \new_[29784]_  = \new_[29783]_  & \new_[29778]_ ;
  assign \new_[29788]_  = ~A168 & ~A169;
  assign \new_[29789]_  = ~A170 & \new_[29788]_ ;
  assign \new_[29793]_  = A233 & A232;
  assign \new_[29794]_  = A202 & \new_[29793]_ ;
  assign \new_[29795]_  = \new_[29794]_  & \new_[29789]_ ;
  assign \new_[29799]_  = ~A265 & ~A235;
  assign \new_[29800]_  = ~A234 & \new_[29799]_ ;
  assign \new_[29804]_  = A301 & ~A268;
  assign \new_[29805]_  = ~A266 & \new_[29804]_ ;
  assign \new_[29806]_  = \new_[29805]_  & \new_[29800]_ ;
  assign \new_[29810]_  = ~A168 & ~A169;
  assign \new_[29811]_  = ~A170 & \new_[29810]_ ;
  assign \new_[29815]_  = ~A233 & ~A232;
  assign \new_[29816]_  = A202 & \new_[29815]_ ;
  assign \new_[29817]_  = \new_[29816]_  & \new_[29811]_ ;
  assign \new_[29821]_  = ~A268 & ~A267;
  assign \new_[29822]_  = ~A235 & \new_[29821]_ ;
  assign \new_[29826]_  = A300 & A299;
  assign \new_[29827]_  = ~A269 & \new_[29826]_ ;
  assign \new_[29828]_  = \new_[29827]_  & \new_[29822]_ ;
  assign \new_[29832]_  = ~A168 & ~A169;
  assign \new_[29833]_  = ~A170 & \new_[29832]_ ;
  assign \new_[29837]_  = ~A233 & ~A232;
  assign \new_[29838]_  = A202 & \new_[29837]_ ;
  assign \new_[29839]_  = \new_[29838]_  & \new_[29833]_ ;
  assign \new_[29843]_  = ~A268 & ~A267;
  assign \new_[29844]_  = ~A235 & \new_[29843]_ ;
  assign \new_[29848]_  = A300 & A298;
  assign \new_[29849]_  = ~A269 & \new_[29848]_ ;
  assign \new_[29850]_  = \new_[29849]_  & \new_[29844]_ ;
  assign \new_[29854]_  = ~A168 & ~A169;
  assign \new_[29855]_  = ~A170 & \new_[29854]_ ;
  assign \new_[29859]_  = ~A233 & ~A232;
  assign \new_[29860]_  = A202 & \new_[29859]_ ;
  assign \new_[29861]_  = \new_[29860]_  & \new_[29855]_ ;
  assign \new_[29865]_  = A266 & A265;
  assign \new_[29866]_  = ~A235 & \new_[29865]_ ;
  assign \new_[29870]_  = A301 & ~A268;
  assign \new_[29871]_  = ~A267 & \new_[29870]_ ;
  assign \new_[29872]_  = \new_[29871]_  & \new_[29866]_ ;
  assign \new_[29876]_  = ~A168 & ~A169;
  assign \new_[29877]_  = ~A170 & \new_[29876]_ ;
  assign \new_[29881]_  = ~A233 & ~A232;
  assign \new_[29882]_  = A202 & \new_[29881]_ ;
  assign \new_[29883]_  = \new_[29882]_  & \new_[29877]_ ;
  assign \new_[29887]_  = ~A266 & ~A265;
  assign \new_[29888]_  = ~A235 & \new_[29887]_ ;
  assign \new_[29892]_  = A300 & A299;
  assign \new_[29893]_  = ~A268 & \new_[29892]_ ;
  assign \new_[29894]_  = \new_[29893]_  & \new_[29888]_ ;
  assign \new_[29898]_  = ~A168 & ~A169;
  assign \new_[29899]_  = ~A170 & \new_[29898]_ ;
  assign \new_[29903]_  = ~A233 & ~A232;
  assign \new_[29904]_  = A202 & \new_[29903]_ ;
  assign \new_[29905]_  = \new_[29904]_  & \new_[29899]_ ;
  assign \new_[29909]_  = ~A266 & ~A265;
  assign \new_[29910]_  = ~A235 & \new_[29909]_ ;
  assign \new_[29914]_  = A300 & A298;
  assign \new_[29915]_  = ~A268 & \new_[29914]_ ;
  assign \new_[29916]_  = \new_[29915]_  & \new_[29910]_ ;
  assign \new_[29920]_  = ~A168 & ~A169;
  assign \new_[29921]_  = ~A170 & \new_[29920]_ ;
  assign \new_[29925]_  = ~A234 & A201;
  assign \new_[29926]_  = A199 & \new_[29925]_ ;
  assign \new_[29927]_  = \new_[29926]_  & \new_[29921]_ ;
  assign \new_[29931]_  = ~A267 & ~A236;
  assign \new_[29932]_  = ~A235 & \new_[29931]_ ;
  assign \new_[29936]_  = A301 & ~A269;
  assign \new_[29937]_  = ~A268 & \new_[29936]_ ;
  assign \new_[29938]_  = \new_[29937]_  & \new_[29932]_ ;
  assign \new_[29942]_  = ~A168 & ~A169;
  assign \new_[29943]_  = ~A170 & \new_[29942]_ ;
  assign \new_[29947]_  = ~A234 & A201;
  assign \new_[29948]_  = A199 & \new_[29947]_ ;
  assign \new_[29949]_  = \new_[29948]_  & \new_[29943]_ ;
  assign \new_[29953]_  = ~A265 & ~A236;
  assign \new_[29954]_  = ~A235 & \new_[29953]_ ;
  assign \new_[29958]_  = A301 & ~A268;
  assign \new_[29959]_  = ~A266 & \new_[29958]_ ;
  assign \new_[29960]_  = \new_[29959]_  & \new_[29954]_ ;
  assign \new_[29964]_  = ~A168 & ~A169;
  assign \new_[29965]_  = ~A170 & \new_[29964]_ ;
  assign \new_[29969]_  = ~A232 & A201;
  assign \new_[29970]_  = A199 & \new_[29969]_ ;
  assign \new_[29971]_  = \new_[29970]_  & \new_[29965]_ ;
  assign \new_[29975]_  = A298 & A236;
  assign \new_[29976]_  = A233 & \new_[29975]_ ;
  assign \new_[29980]_  = ~A301 & ~A300;
  assign \new_[29981]_  = A299 & \new_[29980]_ ;
  assign \new_[29982]_  = \new_[29981]_  & \new_[29976]_ ;
  assign \new_[29986]_  = ~A168 & ~A169;
  assign \new_[29987]_  = ~A170 & \new_[29986]_ ;
  assign \new_[29991]_  = A232 & A201;
  assign \new_[29992]_  = A199 & \new_[29991]_ ;
  assign \new_[29993]_  = \new_[29992]_  & \new_[29987]_ ;
  assign \new_[29997]_  = A298 & A236;
  assign \new_[29998]_  = ~A233 & \new_[29997]_ ;
  assign \new_[30002]_  = ~A301 & ~A300;
  assign \new_[30003]_  = A299 & \new_[30002]_ ;
  assign \new_[30004]_  = \new_[30003]_  & \new_[29998]_ ;
  assign \new_[30008]_  = ~A168 & ~A169;
  assign \new_[30009]_  = ~A170 & \new_[30008]_ ;
  assign \new_[30013]_  = ~A232 & A201;
  assign \new_[30014]_  = A199 & \new_[30013]_ ;
  assign \new_[30015]_  = \new_[30014]_  & \new_[30009]_ ;
  assign \new_[30019]_  = ~A267 & ~A235;
  assign \new_[30020]_  = ~A233 & \new_[30019]_ ;
  assign \new_[30024]_  = A301 & ~A269;
  assign \new_[30025]_  = ~A268 & \new_[30024]_ ;
  assign \new_[30026]_  = \new_[30025]_  & \new_[30020]_ ;
  assign \new_[30030]_  = ~A168 & ~A169;
  assign \new_[30031]_  = ~A170 & \new_[30030]_ ;
  assign \new_[30035]_  = ~A232 & A201;
  assign \new_[30036]_  = A199 & \new_[30035]_ ;
  assign \new_[30037]_  = \new_[30036]_  & \new_[30031]_ ;
  assign \new_[30041]_  = ~A265 & ~A235;
  assign \new_[30042]_  = ~A233 & \new_[30041]_ ;
  assign \new_[30046]_  = A301 & ~A268;
  assign \new_[30047]_  = ~A266 & \new_[30046]_ ;
  assign \new_[30048]_  = \new_[30047]_  & \new_[30042]_ ;
  assign \new_[30052]_  = ~A168 & ~A169;
  assign \new_[30053]_  = ~A170 & \new_[30052]_ ;
  assign \new_[30057]_  = ~A234 & A201;
  assign \new_[30058]_  = A200 & \new_[30057]_ ;
  assign \new_[30059]_  = \new_[30058]_  & \new_[30053]_ ;
  assign \new_[30063]_  = ~A267 & ~A236;
  assign \new_[30064]_  = ~A235 & \new_[30063]_ ;
  assign \new_[30068]_  = A301 & ~A269;
  assign \new_[30069]_  = ~A268 & \new_[30068]_ ;
  assign \new_[30070]_  = \new_[30069]_  & \new_[30064]_ ;
  assign \new_[30074]_  = ~A168 & ~A169;
  assign \new_[30075]_  = ~A170 & \new_[30074]_ ;
  assign \new_[30079]_  = ~A234 & A201;
  assign \new_[30080]_  = A200 & \new_[30079]_ ;
  assign \new_[30081]_  = \new_[30080]_  & \new_[30075]_ ;
  assign \new_[30085]_  = ~A265 & ~A236;
  assign \new_[30086]_  = ~A235 & \new_[30085]_ ;
  assign \new_[30090]_  = A301 & ~A268;
  assign \new_[30091]_  = ~A266 & \new_[30090]_ ;
  assign \new_[30092]_  = \new_[30091]_  & \new_[30086]_ ;
  assign \new_[30096]_  = ~A168 & ~A169;
  assign \new_[30097]_  = ~A170 & \new_[30096]_ ;
  assign \new_[30101]_  = ~A232 & A201;
  assign \new_[30102]_  = A200 & \new_[30101]_ ;
  assign \new_[30103]_  = \new_[30102]_  & \new_[30097]_ ;
  assign \new_[30107]_  = A298 & A236;
  assign \new_[30108]_  = A233 & \new_[30107]_ ;
  assign \new_[30112]_  = ~A301 & ~A300;
  assign \new_[30113]_  = A299 & \new_[30112]_ ;
  assign \new_[30114]_  = \new_[30113]_  & \new_[30108]_ ;
  assign \new_[30118]_  = ~A168 & ~A169;
  assign \new_[30119]_  = ~A170 & \new_[30118]_ ;
  assign \new_[30123]_  = A232 & A201;
  assign \new_[30124]_  = A200 & \new_[30123]_ ;
  assign \new_[30125]_  = \new_[30124]_  & \new_[30119]_ ;
  assign \new_[30129]_  = A298 & A236;
  assign \new_[30130]_  = ~A233 & \new_[30129]_ ;
  assign \new_[30134]_  = ~A301 & ~A300;
  assign \new_[30135]_  = A299 & \new_[30134]_ ;
  assign \new_[30136]_  = \new_[30135]_  & \new_[30130]_ ;
  assign \new_[30140]_  = ~A168 & ~A169;
  assign \new_[30141]_  = ~A170 & \new_[30140]_ ;
  assign \new_[30145]_  = ~A232 & A201;
  assign \new_[30146]_  = A200 & \new_[30145]_ ;
  assign \new_[30147]_  = \new_[30146]_  & \new_[30141]_ ;
  assign \new_[30151]_  = ~A267 & ~A235;
  assign \new_[30152]_  = ~A233 & \new_[30151]_ ;
  assign \new_[30156]_  = A301 & ~A269;
  assign \new_[30157]_  = ~A268 & \new_[30156]_ ;
  assign \new_[30158]_  = \new_[30157]_  & \new_[30152]_ ;
  assign \new_[30162]_  = ~A168 & ~A169;
  assign \new_[30163]_  = ~A170 & \new_[30162]_ ;
  assign \new_[30167]_  = ~A232 & A201;
  assign \new_[30168]_  = A200 & \new_[30167]_ ;
  assign \new_[30169]_  = \new_[30168]_  & \new_[30163]_ ;
  assign \new_[30173]_  = ~A265 & ~A235;
  assign \new_[30174]_  = ~A233 & \new_[30173]_ ;
  assign \new_[30178]_  = A301 & ~A268;
  assign \new_[30179]_  = ~A266 & \new_[30178]_ ;
  assign \new_[30180]_  = \new_[30179]_  & \new_[30174]_ ;
  assign \new_[30184]_  = ~A168 & ~A169;
  assign \new_[30185]_  = ~A170 & \new_[30184]_ ;
  assign \new_[30189]_  = A203 & A200;
  assign \new_[30190]_  = ~A199 & \new_[30189]_ ;
  assign \new_[30191]_  = \new_[30190]_  & \new_[30185]_ ;
  assign \new_[30195]_  = A298 & A234;
  assign \new_[30196]_  = A232 & \new_[30195]_ ;
  assign \new_[30200]_  = ~A301 & ~A300;
  assign \new_[30201]_  = A299 & \new_[30200]_ ;
  assign \new_[30202]_  = \new_[30201]_  & \new_[30196]_ ;
  assign \new_[30206]_  = ~A168 & ~A169;
  assign \new_[30207]_  = ~A170 & \new_[30206]_ ;
  assign \new_[30211]_  = A203 & A200;
  assign \new_[30212]_  = ~A199 & \new_[30211]_ ;
  assign \new_[30213]_  = \new_[30212]_  & \new_[30207]_ ;
  assign \new_[30217]_  = A298 & A234;
  assign \new_[30218]_  = A233 & \new_[30217]_ ;
  assign \new_[30222]_  = ~A301 & ~A300;
  assign \new_[30223]_  = A299 & \new_[30222]_ ;
  assign \new_[30224]_  = \new_[30223]_  & \new_[30218]_ ;
  assign \new_[30228]_  = ~A168 & ~A169;
  assign \new_[30229]_  = ~A170 & \new_[30228]_ ;
  assign \new_[30233]_  = A203 & A200;
  assign \new_[30234]_  = ~A199 & \new_[30233]_ ;
  assign \new_[30235]_  = \new_[30234]_  & \new_[30229]_ ;
  assign \new_[30239]_  = A236 & A233;
  assign \new_[30240]_  = ~A232 & \new_[30239]_ ;
  assign \new_[30244]_  = ~A302 & ~A301;
  assign \new_[30245]_  = ~A300 & \new_[30244]_ ;
  assign \new_[30246]_  = \new_[30245]_  & \new_[30240]_ ;
  assign \new_[30250]_  = ~A168 & ~A169;
  assign \new_[30251]_  = ~A170 & \new_[30250]_ ;
  assign \new_[30255]_  = A203 & A200;
  assign \new_[30256]_  = ~A199 & \new_[30255]_ ;
  assign \new_[30257]_  = \new_[30256]_  & \new_[30251]_ ;
  assign \new_[30261]_  = A236 & A233;
  assign \new_[30262]_  = ~A232 & \new_[30261]_ ;
  assign \new_[30266]_  = ~A301 & ~A299;
  assign \new_[30267]_  = ~A298 & \new_[30266]_ ;
  assign \new_[30268]_  = \new_[30267]_  & \new_[30262]_ ;
  assign \new_[30272]_  = ~A168 & ~A169;
  assign \new_[30273]_  = ~A170 & \new_[30272]_ ;
  assign \new_[30277]_  = A203 & A200;
  assign \new_[30278]_  = ~A199 & \new_[30277]_ ;
  assign \new_[30279]_  = \new_[30278]_  & \new_[30273]_ ;
  assign \new_[30283]_  = A236 & A233;
  assign \new_[30284]_  = ~A232 & \new_[30283]_ ;
  assign \new_[30288]_  = A269 & A266;
  assign \new_[30289]_  = ~A265 & \new_[30288]_ ;
  assign \new_[30290]_  = \new_[30289]_  & \new_[30284]_ ;
  assign \new_[30294]_  = ~A168 & ~A169;
  assign \new_[30295]_  = ~A170 & \new_[30294]_ ;
  assign \new_[30299]_  = A203 & A200;
  assign \new_[30300]_  = ~A199 & \new_[30299]_ ;
  assign \new_[30301]_  = \new_[30300]_  & \new_[30295]_ ;
  assign \new_[30305]_  = A236 & A233;
  assign \new_[30306]_  = ~A232 & \new_[30305]_ ;
  assign \new_[30310]_  = A269 & ~A266;
  assign \new_[30311]_  = A265 & \new_[30310]_ ;
  assign \new_[30312]_  = \new_[30311]_  & \new_[30306]_ ;
  assign \new_[30316]_  = ~A168 & ~A169;
  assign \new_[30317]_  = ~A170 & \new_[30316]_ ;
  assign \new_[30321]_  = A203 & A200;
  assign \new_[30322]_  = ~A199 & \new_[30321]_ ;
  assign \new_[30323]_  = \new_[30322]_  & \new_[30317]_ ;
  assign \new_[30327]_  = A236 & ~A233;
  assign \new_[30328]_  = A232 & \new_[30327]_ ;
  assign \new_[30332]_  = ~A302 & ~A301;
  assign \new_[30333]_  = ~A300 & \new_[30332]_ ;
  assign \new_[30334]_  = \new_[30333]_  & \new_[30328]_ ;
  assign \new_[30338]_  = ~A168 & ~A169;
  assign \new_[30339]_  = ~A170 & \new_[30338]_ ;
  assign \new_[30343]_  = A203 & A200;
  assign \new_[30344]_  = ~A199 & \new_[30343]_ ;
  assign \new_[30345]_  = \new_[30344]_  & \new_[30339]_ ;
  assign \new_[30349]_  = A236 & ~A233;
  assign \new_[30350]_  = A232 & \new_[30349]_ ;
  assign \new_[30354]_  = ~A301 & ~A299;
  assign \new_[30355]_  = ~A298 & \new_[30354]_ ;
  assign \new_[30356]_  = \new_[30355]_  & \new_[30350]_ ;
  assign \new_[30360]_  = ~A168 & ~A169;
  assign \new_[30361]_  = ~A170 & \new_[30360]_ ;
  assign \new_[30365]_  = A203 & A200;
  assign \new_[30366]_  = ~A199 & \new_[30365]_ ;
  assign \new_[30367]_  = \new_[30366]_  & \new_[30361]_ ;
  assign \new_[30371]_  = A236 & ~A233;
  assign \new_[30372]_  = A232 & \new_[30371]_ ;
  assign \new_[30376]_  = A269 & A266;
  assign \new_[30377]_  = ~A265 & \new_[30376]_ ;
  assign \new_[30378]_  = \new_[30377]_  & \new_[30372]_ ;
  assign \new_[30382]_  = ~A168 & ~A169;
  assign \new_[30383]_  = ~A170 & \new_[30382]_ ;
  assign \new_[30387]_  = A203 & A200;
  assign \new_[30388]_  = ~A199 & \new_[30387]_ ;
  assign \new_[30389]_  = \new_[30388]_  & \new_[30383]_ ;
  assign \new_[30393]_  = A236 & ~A233;
  assign \new_[30394]_  = A232 & \new_[30393]_ ;
  assign \new_[30398]_  = A269 & ~A266;
  assign \new_[30399]_  = A265 & \new_[30398]_ ;
  assign \new_[30400]_  = \new_[30399]_  & \new_[30394]_ ;
  assign \new_[30404]_  = ~A168 & ~A169;
  assign \new_[30405]_  = ~A170 & \new_[30404]_ ;
  assign \new_[30409]_  = A203 & ~A200;
  assign \new_[30410]_  = A199 & \new_[30409]_ ;
  assign \new_[30411]_  = \new_[30410]_  & \new_[30405]_ ;
  assign \new_[30415]_  = A298 & A234;
  assign \new_[30416]_  = A232 & \new_[30415]_ ;
  assign \new_[30420]_  = ~A301 & ~A300;
  assign \new_[30421]_  = A299 & \new_[30420]_ ;
  assign \new_[30422]_  = \new_[30421]_  & \new_[30416]_ ;
  assign \new_[30426]_  = ~A168 & ~A169;
  assign \new_[30427]_  = ~A170 & \new_[30426]_ ;
  assign \new_[30431]_  = A203 & ~A200;
  assign \new_[30432]_  = A199 & \new_[30431]_ ;
  assign \new_[30433]_  = \new_[30432]_  & \new_[30427]_ ;
  assign \new_[30437]_  = A298 & A234;
  assign \new_[30438]_  = A233 & \new_[30437]_ ;
  assign \new_[30442]_  = ~A301 & ~A300;
  assign \new_[30443]_  = A299 & \new_[30442]_ ;
  assign \new_[30444]_  = \new_[30443]_  & \new_[30438]_ ;
  assign \new_[30448]_  = ~A168 & ~A169;
  assign \new_[30449]_  = ~A170 & \new_[30448]_ ;
  assign \new_[30453]_  = A203 & ~A200;
  assign \new_[30454]_  = A199 & \new_[30453]_ ;
  assign \new_[30455]_  = \new_[30454]_  & \new_[30449]_ ;
  assign \new_[30459]_  = A236 & A233;
  assign \new_[30460]_  = ~A232 & \new_[30459]_ ;
  assign \new_[30464]_  = ~A302 & ~A301;
  assign \new_[30465]_  = ~A300 & \new_[30464]_ ;
  assign \new_[30466]_  = \new_[30465]_  & \new_[30460]_ ;
  assign \new_[30470]_  = ~A168 & ~A169;
  assign \new_[30471]_  = ~A170 & \new_[30470]_ ;
  assign \new_[30475]_  = A203 & ~A200;
  assign \new_[30476]_  = A199 & \new_[30475]_ ;
  assign \new_[30477]_  = \new_[30476]_  & \new_[30471]_ ;
  assign \new_[30481]_  = A236 & A233;
  assign \new_[30482]_  = ~A232 & \new_[30481]_ ;
  assign \new_[30486]_  = ~A301 & ~A299;
  assign \new_[30487]_  = ~A298 & \new_[30486]_ ;
  assign \new_[30488]_  = \new_[30487]_  & \new_[30482]_ ;
  assign \new_[30492]_  = ~A168 & ~A169;
  assign \new_[30493]_  = ~A170 & \new_[30492]_ ;
  assign \new_[30497]_  = A203 & ~A200;
  assign \new_[30498]_  = A199 & \new_[30497]_ ;
  assign \new_[30499]_  = \new_[30498]_  & \new_[30493]_ ;
  assign \new_[30503]_  = A236 & A233;
  assign \new_[30504]_  = ~A232 & \new_[30503]_ ;
  assign \new_[30508]_  = A269 & A266;
  assign \new_[30509]_  = ~A265 & \new_[30508]_ ;
  assign \new_[30510]_  = \new_[30509]_  & \new_[30504]_ ;
  assign \new_[30514]_  = ~A168 & ~A169;
  assign \new_[30515]_  = ~A170 & \new_[30514]_ ;
  assign \new_[30519]_  = A203 & ~A200;
  assign \new_[30520]_  = A199 & \new_[30519]_ ;
  assign \new_[30521]_  = \new_[30520]_  & \new_[30515]_ ;
  assign \new_[30525]_  = A236 & A233;
  assign \new_[30526]_  = ~A232 & \new_[30525]_ ;
  assign \new_[30530]_  = A269 & ~A266;
  assign \new_[30531]_  = A265 & \new_[30530]_ ;
  assign \new_[30532]_  = \new_[30531]_  & \new_[30526]_ ;
  assign \new_[30536]_  = ~A168 & ~A169;
  assign \new_[30537]_  = ~A170 & \new_[30536]_ ;
  assign \new_[30541]_  = A203 & ~A200;
  assign \new_[30542]_  = A199 & \new_[30541]_ ;
  assign \new_[30543]_  = \new_[30542]_  & \new_[30537]_ ;
  assign \new_[30547]_  = A236 & ~A233;
  assign \new_[30548]_  = A232 & \new_[30547]_ ;
  assign \new_[30552]_  = ~A302 & ~A301;
  assign \new_[30553]_  = ~A300 & \new_[30552]_ ;
  assign \new_[30554]_  = \new_[30553]_  & \new_[30548]_ ;
  assign \new_[30558]_  = ~A168 & ~A169;
  assign \new_[30559]_  = ~A170 & \new_[30558]_ ;
  assign \new_[30563]_  = A203 & ~A200;
  assign \new_[30564]_  = A199 & \new_[30563]_ ;
  assign \new_[30565]_  = \new_[30564]_  & \new_[30559]_ ;
  assign \new_[30569]_  = A236 & ~A233;
  assign \new_[30570]_  = A232 & \new_[30569]_ ;
  assign \new_[30574]_  = ~A301 & ~A299;
  assign \new_[30575]_  = ~A298 & \new_[30574]_ ;
  assign \new_[30576]_  = \new_[30575]_  & \new_[30570]_ ;
  assign \new_[30580]_  = ~A168 & ~A169;
  assign \new_[30581]_  = ~A170 & \new_[30580]_ ;
  assign \new_[30585]_  = A203 & ~A200;
  assign \new_[30586]_  = A199 & \new_[30585]_ ;
  assign \new_[30587]_  = \new_[30586]_  & \new_[30581]_ ;
  assign \new_[30591]_  = A236 & ~A233;
  assign \new_[30592]_  = A232 & \new_[30591]_ ;
  assign \new_[30596]_  = A269 & A266;
  assign \new_[30597]_  = ~A265 & \new_[30596]_ ;
  assign \new_[30598]_  = \new_[30597]_  & \new_[30592]_ ;
  assign \new_[30602]_  = ~A168 & ~A169;
  assign \new_[30603]_  = ~A170 & \new_[30602]_ ;
  assign \new_[30607]_  = A203 & ~A200;
  assign \new_[30608]_  = A199 & \new_[30607]_ ;
  assign \new_[30609]_  = \new_[30608]_  & \new_[30603]_ ;
  assign \new_[30613]_  = A236 & ~A233;
  assign \new_[30614]_  = A232 & \new_[30613]_ ;
  assign \new_[30618]_  = A269 & ~A266;
  assign \new_[30619]_  = A265 & \new_[30618]_ ;
  assign \new_[30620]_  = \new_[30619]_  & \new_[30614]_ ;
  assign \new_[30624]_  = ~A201 & A166;
  assign \new_[30625]_  = A168 & \new_[30624]_ ;
  assign \new_[30629]_  = ~A234 & ~A203;
  assign \new_[30630]_  = ~A202 & \new_[30629]_ ;
  assign \new_[30631]_  = \new_[30630]_  & \new_[30625]_ ;
  assign \new_[30635]_  = ~A267 & ~A236;
  assign \new_[30636]_  = ~A235 & \new_[30635]_ ;
  assign \new_[30639]_  = ~A269 & ~A268;
  assign \new_[30642]_  = A300 & A299;
  assign \new_[30643]_  = \new_[30642]_  & \new_[30639]_ ;
  assign \new_[30644]_  = \new_[30643]_  & \new_[30636]_ ;
  assign \new_[30648]_  = ~A201 & A166;
  assign \new_[30649]_  = A168 & \new_[30648]_ ;
  assign \new_[30653]_  = ~A234 & ~A203;
  assign \new_[30654]_  = ~A202 & \new_[30653]_ ;
  assign \new_[30655]_  = \new_[30654]_  & \new_[30649]_ ;
  assign \new_[30659]_  = ~A267 & ~A236;
  assign \new_[30660]_  = ~A235 & \new_[30659]_ ;
  assign \new_[30663]_  = ~A269 & ~A268;
  assign \new_[30666]_  = A300 & A298;
  assign \new_[30667]_  = \new_[30666]_  & \new_[30663]_ ;
  assign \new_[30668]_  = \new_[30667]_  & \new_[30660]_ ;
  assign \new_[30672]_  = ~A201 & A166;
  assign \new_[30673]_  = A168 & \new_[30672]_ ;
  assign \new_[30677]_  = ~A234 & ~A203;
  assign \new_[30678]_  = ~A202 & \new_[30677]_ ;
  assign \new_[30679]_  = \new_[30678]_  & \new_[30673]_ ;
  assign \new_[30683]_  = A265 & ~A236;
  assign \new_[30684]_  = ~A235 & \new_[30683]_ ;
  assign \new_[30687]_  = ~A267 & A266;
  assign \new_[30690]_  = A301 & ~A268;
  assign \new_[30691]_  = \new_[30690]_  & \new_[30687]_ ;
  assign \new_[30692]_  = \new_[30691]_  & \new_[30684]_ ;
  assign \new_[30696]_  = ~A201 & A166;
  assign \new_[30697]_  = A168 & \new_[30696]_ ;
  assign \new_[30701]_  = ~A234 & ~A203;
  assign \new_[30702]_  = ~A202 & \new_[30701]_ ;
  assign \new_[30703]_  = \new_[30702]_  & \new_[30697]_ ;
  assign \new_[30707]_  = ~A265 & ~A236;
  assign \new_[30708]_  = ~A235 & \new_[30707]_ ;
  assign \new_[30711]_  = ~A268 & ~A266;
  assign \new_[30714]_  = A300 & A299;
  assign \new_[30715]_  = \new_[30714]_  & \new_[30711]_ ;
  assign \new_[30716]_  = \new_[30715]_  & \new_[30708]_ ;
  assign \new_[30720]_  = ~A201 & A166;
  assign \new_[30721]_  = A168 & \new_[30720]_ ;
  assign \new_[30725]_  = ~A234 & ~A203;
  assign \new_[30726]_  = ~A202 & \new_[30725]_ ;
  assign \new_[30727]_  = \new_[30726]_  & \new_[30721]_ ;
  assign \new_[30731]_  = ~A265 & ~A236;
  assign \new_[30732]_  = ~A235 & \new_[30731]_ ;
  assign \new_[30735]_  = ~A268 & ~A266;
  assign \new_[30738]_  = A300 & A298;
  assign \new_[30739]_  = \new_[30738]_  & \new_[30735]_ ;
  assign \new_[30740]_  = \new_[30739]_  & \new_[30732]_ ;
  assign \new_[30744]_  = ~A201 & A166;
  assign \new_[30745]_  = A168 & \new_[30744]_ ;
  assign \new_[30749]_  = A232 & ~A203;
  assign \new_[30750]_  = ~A202 & \new_[30749]_ ;
  assign \new_[30751]_  = \new_[30750]_  & \new_[30745]_ ;
  assign \new_[30755]_  = ~A235 & ~A234;
  assign \new_[30756]_  = A233 & \new_[30755]_ ;
  assign \new_[30759]_  = ~A268 & ~A267;
  assign \new_[30762]_  = A301 & ~A269;
  assign \new_[30763]_  = \new_[30762]_  & \new_[30759]_ ;
  assign \new_[30764]_  = \new_[30763]_  & \new_[30756]_ ;
  assign \new_[30768]_  = ~A201 & A166;
  assign \new_[30769]_  = A168 & \new_[30768]_ ;
  assign \new_[30773]_  = A232 & ~A203;
  assign \new_[30774]_  = ~A202 & \new_[30773]_ ;
  assign \new_[30775]_  = \new_[30774]_  & \new_[30769]_ ;
  assign \new_[30779]_  = ~A235 & ~A234;
  assign \new_[30780]_  = A233 & \new_[30779]_ ;
  assign \new_[30783]_  = ~A266 & ~A265;
  assign \new_[30786]_  = A301 & ~A268;
  assign \new_[30787]_  = \new_[30786]_  & \new_[30783]_ ;
  assign \new_[30788]_  = \new_[30787]_  & \new_[30780]_ ;
  assign \new_[30792]_  = ~A201 & A166;
  assign \new_[30793]_  = A168 & \new_[30792]_ ;
  assign \new_[30797]_  = ~A232 & ~A203;
  assign \new_[30798]_  = ~A202 & \new_[30797]_ ;
  assign \new_[30799]_  = \new_[30798]_  & \new_[30793]_ ;
  assign \new_[30803]_  = ~A267 & ~A235;
  assign \new_[30804]_  = ~A233 & \new_[30803]_ ;
  assign \new_[30807]_  = ~A269 & ~A268;
  assign \new_[30810]_  = A300 & A299;
  assign \new_[30811]_  = \new_[30810]_  & \new_[30807]_ ;
  assign \new_[30812]_  = \new_[30811]_  & \new_[30804]_ ;
  assign \new_[30816]_  = ~A201 & A166;
  assign \new_[30817]_  = A168 & \new_[30816]_ ;
  assign \new_[30821]_  = ~A232 & ~A203;
  assign \new_[30822]_  = ~A202 & \new_[30821]_ ;
  assign \new_[30823]_  = \new_[30822]_  & \new_[30817]_ ;
  assign \new_[30827]_  = ~A267 & ~A235;
  assign \new_[30828]_  = ~A233 & \new_[30827]_ ;
  assign \new_[30831]_  = ~A269 & ~A268;
  assign \new_[30834]_  = A300 & A298;
  assign \new_[30835]_  = \new_[30834]_  & \new_[30831]_ ;
  assign \new_[30836]_  = \new_[30835]_  & \new_[30828]_ ;
  assign \new_[30840]_  = ~A201 & A166;
  assign \new_[30841]_  = A168 & \new_[30840]_ ;
  assign \new_[30845]_  = ~A232 & ~A203;
  assign \new_[30846]_  = ~A202 & \new_[30845]_ ;
  assign \new_[30847]_  = \new_[30846]_  & \new_[30841]_ ;
  assign \new_[30851]_  = A265 & ~A235;
  assign \new_[30852]_  = ~A233 & \new_[30851]_ ;
  assign \new_[30855]_  = ~A267 & A266;
  assign \new_[30858]_  = A301 & ~A268;
  assign \new_[30859]_  = \new_[30858]_  & \new_[30855]_ ;
  assign \new_[30860]_  = \new_[30859]_  & \new_[30852]_ ;
  assign \new_[30864]_  = ~A201 & A166;
  assign \new_[30865]_  = A168 & \new_[30864]_ ;
  assign \new_[30869]_  = ~A232 & ~A203;
  assign \new_[30870]_  = ~A202 & \new_[30869]_ ;
  assign \new_[30871]_  = \new_[30870]_  & \new_[30865]_ ;
  assign \new_[30875]_  = ~A265 & ~A235;
  assign \new_[30876]_  = ~A233 & \new_[30875]_ ;
  assign \new_[30879]_  = ~A268 & ~A266;
  assign \new_[30882]_  = A300 & A299;
  assign \new_[30883]_  = \new_[30882]_  & \new_[30879]_ ;
  assign \new_[30884]_  = \new_[30883]_  & \new_[30876]_ ;
  assign \new_[30888]_  = ~A201 & A166;
  assign \new_[30889]_  = A168 & \new_[30888]_ ;
  assign \new_[30893]_  = ~A232 & ~A203;
  assign \new_[30894]_  = ~A202 & \new_[30893]_ ;
  assign \new_[30895]_  = \new_[30894]_  & \new_[30889]_ ;
  assign \new_[30899]_  = ~A265 & ~A235;
  assign \new_[30900]_  = ~A233 & \new_[30899]_ ;
  assign \new_[30903]_  = ~A268 & ~A266;
  assign \new_[30906]_  = A300 & A298;
  assign \new_[30907]_  = \new_[30906]_  & \new_[30903]_ ;
  assign \new_[30908]_  = \new_[30907]_  & \new_[30900]_ ;
  assign \new_[30912]_  = A199 & A166;
  assign \new_[30913]_  = A168 & \new_[30912]_ ;
  assign \new_[30917]_  = ~A202 & ~A201;
  assign \new_[30918]_  = A200 & \new_[30917]_ ;
  assign \new_[30919]_  = \new_[30918]_  & \new_[30913]_ ;
  assign \new_[30923]_  = ~A236 & ~A235;
  assign \new_[30924]_  = ~A234 & \new_[30923]_ ;
  assign \new_[30927]_  = ~A268 & ~A267;
  assign \new_[30930]_  = A301 & ~A269;
  assign \new_[30931]_  = \new_[30930]_  & \new_[30927]_ ;
  assign \new_[30932]_  = \new_[30931]_  & \new_[30924]_ ;
  assign \new_[30936]_  = A199 & A166;
  assign \new_[30937]_  = A168 & \new_[30936]_ ;
  assign \new_[30941]_  = ~A202 & ~A201;
  assign \new_[30942]_  = A200 & \new_[30941]_ ;
  assign \new_[30943]_  = \new_[30942]_  & \new_[30937]_ ;
  assign \new_[30947]_  = ~A236 & ~A235;
  assign \new_[30948]_  = ~A234 & \new_[30947]_ ;
  assign \new_[30951]_  = ~A266 & ~A265;
  assign \new_[30954]_  = A301 & ~A268;
  assign \new_[30955]_  = \new_[30954]_  & \new_[30951]_ ;
  assign \new_[30956]_  = \new_[30955]_  & \new_[30948]_ ;
  assign \new_[30960]_  = A199 & A166;
  assign \new_[30961]_  = A168 & \new_[30960]_ ;
  assign \new_[30965]_  = ~A202 & ~A201;
  assign \new_[30966]_  = A200 & \new_[30965]_ ;
  assign \new_[30967]_  = \new_[30966]_  & \new_[30961]_ ;
  assign \new_[30971]_  = A236 & A233;
  assign \new_[30972]_  = ~A232 & \new_[30971]_ ;
  assign \new_[30975]_  = A299 & A298;
  assign \new_[30978]_  = ~A301 & ~A300;
  assign \new_[30979]_  = \new_[30978]_  & \new_[30975]_ ;
  assign \new_[30980]_  = \new_[30979]_  & \new_[30972]_ ;
  assign \new_[30984]_  = A199 & A166;
  assign \new_[30985]_  = A168 & \new_[30984]_ ;
  assign \new_[30989]_  = ~A202 & ~A201;
  assign \new_[30990]_  = A200 & \new_[30989]_ ;
  assign \new_[30991]_  = \new_[30990]_  & \new_[30985]_ ;
  assign \new_[30995]_  = A236 & ~A233;
  assign \new_[30996]_  = A232 & \new_[30995]_ ;
  assign \new_[30999]_  = A299 & A298;
  assign \new_[31002]_  = ~A301 & ~A300;
  assign \new_[31003]_  = \new_[31002]_  & \new_[30999]_ ;
  assign \new_[31004]_  = \new_[31003]_  & \new_[30996]_ ;
  assign \new_[31008]_  = A199 & A166;
  assign \new_[31009]_  = A168 & \new_[31008]_ ;
  assign \new_[31013]_  = ~A202 & ~A201;
  assign \new_[31014]_  = A200 & \new_[31013]_ ;
  assign \new_[31015]_  = \new_[31014]_  & \new_[31009]_ ;
  assign \new_[31019]_  = ~A235 & ~A233;
  assign \new_[31020]_  = ~A232 & \new_[31019]_ ;
  assign \new_[31023]_  = ~A268 & ~A267;
  assign \new_[31026]_  = A301 & ~A269;
  assign \new_[31027]_  = \new_[31026]_  & \new_[31023]_ ;
  assign \new_[31028]_  = \new_[31027]_  & \new_[31020]_ ;
  assign \new_[31032]_  = A199 & A166;
  assign \new_[31033]_  = A168 & \new_[31032]_ ;
  assign \new_[31037]_  = ~A202 & ~A201;
  assign \new_[31038]_  = A200 & \new_[31037]_ ;
  assign \new_[31039]_  = \new_[31038]_  & \new_[31033]_ ;
  assign \new_[31043]_  = ~A235 & ~A233;
  assign \new_[31044]_  = ~A232 & \new_[31043]_ ;
  assign \new_[31047]_  = ~A266 & ~A265;
  assign \new_[31050]_  = A301 & ~A268;
  assign \new_[31051]_  = \new_[31050]_  & \new_[31047]_ ;
  assign \new_[31052]_  = \new_[31051]_  & \new_[31044]_ ;
  assign \new_[31056]_  = ~A199 & A166;
  assign \new_[31057]_  = A168 & \new_[31056]_ ;
  assign \new_[31061]_  = ~A234 & ~A202;
  assign \new_[31062]_  = ~A200 & \new_[31061]_ ;
  assign \new_[31063]_  = \new_[31062]_  & \new_[31057]_ ;
  assign \new_[31067]_  = ~A267 & ~A236;
  assign \new_[31068]_  = ~A235 & \new_[31067]_ ;
  assign \new_[31071]_  = ~A269 & ~A268;
  assign \new_[31074]_  = A300 & A299;
  assign \new_[31075]_  = \new_[31074]_  & \new_[31071]_ ;
  assign \new_[31076]_  = \new_[31075]_  & \new_[31068]_ ;
  assign \new_[31080]_  = ~A199 & A166;
  assign \new_[31081]_  = A168 & \new_[31080]_ ;
  assign \new_[31085]_  = ~A234 & ~A202;
  assign \new_[31086]_  = ~A200 & \new_[31085]_ ;
  assign \new_[31087]_  = \new_[31086]_  & \new_[31081]_ ;
  assign \new_[31091]_  = ~A267 & ~A236;
  assign \new_[31092]_  = ~A235 & \new_[31091]_ ;
  assign \new_[31095]_  = ~A269 & ~A268;
  assign \new_[31098]_  = A300 & A298;
  assign \new_[31099]_  = \new_[31098]_  & \new_[31095]_ ;
  assign \new_[31100]_  = \new_[31099]_  & \new_[31092]_ ;
  assign \new_[31104]_  = ~A199 & A166;
  assign \new_[31105]_  = A168 & \new_[31104]_ ;
  assign \new_[31109]_  = ~A234 & ~A202;
  assign \new_[31110]_  = ~A200 & \new_[31109]_ ;
  assign \new_[31111]_  = \new_[31110]_  & \new_[31105]_ ;
  assign \new_[31115]_  = A265 & ~A236;
  assign \new_[31116]_  = ~A235 & \new_[31115]_ ;
  assign \new_[31119]_  = ~A267 & A266;
  assign \new_[31122]_  = A301 & ~A268;
  assign \new_[31123]_  = \new_[31122]_  & \new_[31119]_ ;
  assign \new_[31124]_  = \new_[31123]_  & \new_[31116]_ ;
  assign \new_[31128]_  = ~A199 & A166;
  assign \new_[31129]_  = A168 & \new_[31128]_ ;
  assign \new_[31133]_  = ~A234 & ~A202;
  assign \new_[31134]_  = ~A200 & \new_[31133]_ ;
  assign \new_[31135]_  = \new_[31134]_  & \new_[31129]_ ;
  assign \new_[31139]_  = ~A265 & ~A236;
  assign \new_[31140]_  = ~A235 & \new_[31139]_ ;
  assign \new_[31143]_  = ~A268 & ~A266;
  assign \new_[31146]_  = A300 & A299;
  assign \new_[31147]_  = \new_[31146]_  & \new_[31143]_ ;
  assign \new_[31148]_  = \new_[31147]_  & \new_[31140]_ ;
  assign \new_[31152]_  = ~A199 & A166;
  assign \new_[31153]_  = A168 & \new_[31152]_ ;
  assign \new_[31157]_  = ~A234 & ~A202;
  assign \new_[31158]_  = ~A200 & \new_[31157]_ ;
  assign \new_[31159]_  = \new_[31158]_  & \new_[31153]_ ;
  assign \new_[31163]_  = ~A265 & ~A236;
  assign \new_[31164]_  = ~A235 & \new_[31163]_ ;
  assign \new_[31167]_  = ~A268 & ~A266;
  assign \new_[31170]_  = A300 & A298;
  assign \new_[31171]_  = \new_[31170]_  & \new_[31167]_ ;
  assign \new_[31172]_  = \new_[31171]_  & \new_[31164]_ ;
  assign \new_[31176]_  = ~A199 & A166;
  assign \new_[31177]_  = A168 & \new_[31176]_ ;
  assign \new_[31181]_  = A232 & ~A202;
  assign \new_[31182]_  = ~A200 & \new_[31181]_ ;
  assign \new_[31183]_  = \new_[31182]_  & \new_[31177]_ ;
  assign \new_[31187]_  = ~A235 & ~A234;
  assign \new_[31188]_  = A233 & \new_[31187]_ ;
  assign \new_[31191]_  = ~A268 & ~A267;
  assign \new_[31194]_  = A301 & ~A269;
  assign \new_[31195]_  = \new_[31194]_  & \new_[31191]_ ;
  assign \new_[31196]_  = \new_[31195]_  & \new_[31188]_ ;
  assign \new_[31200]_  = ~A199 & A166;
  assign \new_[31201]_  = A168 & \new_[31200]_ ;
  assign \new_[31205]_  = A232 & ~A202;
  assign \new_[31206]_  = ~A200 & \new_[31205]_ ;
  assign \new_[31207]_  = \new_[31206]_  & \new_[31201]_ ;
  assign \new_[31211]_  = ~A235 & ~A234;
  assign \new_[31212]_  = A233 & \new_[31211]_ ;
  assign \new_[31215]_  = ~A266 & ~A265;
  assign \new_[31218]_  = A301 & ~A268;
  assign \new_[31219]_  = \new_[31218]_  & \new_[31215]_ ;
  assign \new_[31220]_  = \new_[31219]_  & \new_[31212]_ ;
  assign \new_[31224]_  = ~A199 & A166;
  assign \new_[31225]_  = A168 & \new_[31224]_ ;
  assign \new_[31229]_  = ~A232 & ~A202;
  assign \new_[31230]_  = ~A200 & \new_[31229]_ ;
  assign \new_[31231]_  = \new_[31230]_  & \new_[31225]_ ;
  assign \new_[31235]_  = ~A267 & ~A235;
  assign \new_[31236]_  = ~A233 & \new_[31235]_ ;
  assign \new_[31239]_  = ~A269 & ~A268;
  assign \new_[31242]_  = A300 & A299;
  assign \new_[31243]_  = \new_[31242]_  & \new_[31239]_ ;
  assign \new_[31244]_  = \new_[31243]_  & \new_[31236]_ ;
  assign \new_[31248]_  = ~A199 & A166;
  assign \new_[31249]_  = A168 & \new_[31248]_ ;
  assign \new_[31253]_  = ~A232 & ~A202;
  assign \new_[31254]_  = ~A200 & \new_[31253]_ ;
  assign \new_[31255]_  = \new_[31254]_  & \new_[31249]_ ;
  assign \new_[31259]_  = ~A267 & ~A235;
  assign \new_[31260]_  = ~A233 & \new_[31259]_ ;
  assign \new_[31263]_  = ~A269 & ~A268;
  assign \new_[31266]_  = A300 & A298;
  assign \new_[31267]_  = \new_[31266]_  & \new_[31263]_ ;
  assign \new_[31268]_  = \new_[31267]_  & \new_[31260]_ ;
  assign \new_[31272]_  = ~A199 & A166;
  assign \new_[31273]_  = A168 & \new_[31272]_ ;
  assign \new_[31277]_  = ~A232 & ~A202;
  assign \new_[31278]_  = ~A200 & \new_[31277]_ ;
  assign \new_[31279]_  = \new_[31278]_  & \new_[31273]_ ;
  assign \new_[31283]_  = A265 & ~A235;
  assign \new_[31284]_  = ~A233 & \new_[31283]_ ;
  assign \new_[31287]_  = ~A267 & A266;
  assign \new_[31290]_  = A301 & ~A268;
  assign \new_[31291]_  = \new_[31290]_  & \new_[31287]_ ;
  assign \new_[31292]_  = \new_[31291]_  & \new_[31284]_ ;
  assign \new_[31296]_  = ~A199 & A166;
  assign \new_[31297]_  = A168 & \new_[31296]_ ;
  assign \new_[31301]_  = ~A232 & ~A202;
  assign \new_[31302]_  = ~A200 & \new_[31301]_ ;
  assign \new_[31303]_  = \new_[31302]_  & \new_[31297]_ ;
  assign \new_[31307]_  = ~A265 & ~A235;
  assign \new_[31308]_  = ~A233 & \new_[31307]_ ;
  assign \new_[31311]_  = ~A268 & ~A266;
  assign \new_[31314]_  = A300 & A299;
  assign \new_[31315]_  = \new_[31314]_  & \new_[31311]_ ;
  assign \new_[31316]_  = \new_[31315]_  & \new_[31308]_ ;
  assign \new_[31320]_  = ~A199 & A166;
  assign \new_[31321]_  = A168 & \new_[31320]_ ;
  assign \new_[31325]_  = ~A232 & ~A202;
  assign \new_[31326]_  = ~A200 & \new_[31325]_ ;
  assign \new_[31327]_  = \new_[31326]_  & \new_[31321]_ ;
  assign \new_[31331]_  = ~A265 & ~A235;
  assign \new_[31332]_  = ~A233 & \new_[31331]_ ;
  assign \new_[31335]_  = ~A268 & ~A266;
  assign \new_[31338]_  = A300 & A298;
  assign \new_[31339]_  = \new_[31338]_  & \new_[31335]_ ;
  assign \new_[31340]_  = \new_[31339]_  & \new_[31332]_ ;
  assign \new_[31344]_  = ~A201 & A167;
  assign \new_[31345]_  = A168 & \new_[31344]_ ;
  assign \new_[31349]_  = ~A234 & ~A203;
  assign \new_[31350]_  = ~A202 & \new_[31349]_ ;
  assign \new_[31351]_  = \new_[31350]_  & \new_[31345]_ ;
  assign \new_[31355]_  = ~A267 & ~A236;
  assign \new_[31356]_  = ~A235 & \new_[31355]_ ;
  assign \new_[31359]_  = ~A269 & ~A268;
  assign \new_[31362]_  = A300 & A299;
  assign \new_[31363]_  = \new_[31362]_  & \new_[31359]_ ;
  assign \new_[31364]_  = \new_[31363]_  & \new_[31356]_ ;
  assign \new_[31368]_  = ~A201 & A167;
  assign \new_[31369]_  = A168 & \new_[31368]_ ;
  assign \new_[31373]_  = ~A234 & ~A203;
  assign \new_[31374]_  = ~A202 & \new_[31373]_ ;
  assign \new_[31375]_  = \new_[31374]_  & \new_[31369]_ ;
  assign \new_[31379]_  = ~A267 & ~A236;
  assign \new_[31380]_  = ~A235 & \new_[31379]_ ;
  assign \new_[31383]_  = ~A269 & ~A268;
  assign \new_[31386]_  = A300 & A298;
  assign \new_[31387]_  = \new_[31386]_  & \new_[31383]_ ;
  assign \new_[31388]_  = \new_[31387]_  & \new_[31380]_ ;
  assign \new_[31392]_  = ~A201 & A167;
  assign \new_[31393]_  = A168 & \new_[31392]_ ;
  assign \new_[31397]_  = ~A234 & ~A203;
  assign \new_[31398]_  = ~A202 & \new_[31397]_ ;
  assign \new_[31399]_  = \new_[31398]_  & \new_[31393]_ ;
  assign \new_[31403]_  = A265 & ~A236;
  assign \new_[31404]_  = ~A235 & \new_[31403]_ ;
  assign \new_[31407]_  = ~A267 & A266;
  assign \new_[31410]_  = A301 & ~A268;
  assign \new_[31411]_  = \new_[31410]_  & \new_[31407]_ ;
  assign \new_[31412]_  = \new_[31411]_  & \new_[31404]_ ;
  assign \new_[31416]_  = ~A201 & A167;
  assign \new_[31417]_  = A168 & \new_[31416]_ ;
  assign \new_[31421]_  = ~A234 & ~A203;
  assign \new_[31422]_  = ~A202 & \new_[31421]_ ;
  assign \new_[31423]_  = \new_[31422]_  & \new_[31417]_ ;
  assign \new_[31427]_  = ~A265 & ~A236;
  assign \new_[31428]_  = ~A235 & \new_[31427]_ ;
  assign \new_[31431]_  = ~A268 & ~A266;
  assign \new_[31434]_  = A300 & A299;
  assign \new_[31435]_  = \new_[31434]_  & \new_[31431]_ ;
  assign \new_[31436]_  = \new_[31435]_  & \new_[31428]_ ;
  assign \new_[31440]_  = ~A201 & A167;
  assign \new_[31441]_  = A168 & \new_[31440]_ ;
  assign \new_[31445]_  = ~A234 & ~A203;
  assign \new_[31446]_  = ~A202 & \new_[31445]_ ;
  assign \new_[31447]_  = \new_[31446]_  & \new_[31441]_ ;
  assign \new_[31451]_  = ~A265 & ~A236;
  assign \new_[31452]_  = ~A235 & \new_[31451]_ ;
  assign \new_[31455]_  = ~A268 & ~A266;
  assign \new_[31458]_  = A300 & A298;
  assign \new_[31459]_  = \new_[31458]_  & \new_[31455]_ ;
  assign \new_[31460]_  = \new_[31459]_  & \new_[31452]_ ;
  assign \new_[31464]_  = ~A201 & A167;
  assign \new_[31465]_  = A168 & \new_[31464]_ ;
  assign \new_[31469]_  = A232 & ~A203;
  assign \new_[31470]_  = ~A202 & \new_[31469]_ ;
  assign \new_[31471]_  = \new_[31470]_  & \new_[31465]_ ;
  assign \new_[31475]_  = ~A235 & ~A234;
  assign \new_[31476]_  = A233 & \new_[31475]_ ;
  assign \new_[31479]_  = ~A268 & ~A267;
  assign \new_[31482]_  = A301 & ~A269;
  assign \new_[31483]_  = \new_[31482]_  & \new_[31479]_ ;
  assign \new_[31484]_  = \new_[31483]_  & \new_[31476]_ ;
  assign \new_[31488]_  = ~A201 & A167;
  assign \new_[31489]_  = A168 & \new_[31488]_ ;
  assign \new_[31493]_  = A232 & ~A203;
  assign \new_[31494]_  = ~A202 & \new_[31493]_ ;
  assign \new_[31495]_  = \new_[31494]_  & \new_[31489]_ ;
  assign \new_[31499]_  = ~A235 & ~A234;
  assign \new_[31500]_  = A233 & \new_[31499]_ ;
  assign \new_[31503]_  = ~A266 & ~A265;
  assign \new_[31506]_  = A301 & ~A268;
  assign \new_[31507]_  = \new_[31506]_  & \new_[31503]_ ;
  assign \new_[31508]_  = \new_[31507]_  & \new_[31500]_ ;
  assign \new_[31512]_  = ~A201 & A167;
  assign \new_[31513]_  = A168 & \new_[31512]_ ;
  assign \new_[31517]_  = ~A232 & ~A203;
  assign \new_[31518]_  = ~A202 & \new_[31517]_ ;
  assign \new_[31519]_  = \new_[31518]_  & \new_[31513]_ ;
  assign \new_[31523]_  = ~A267 & ~A235;
  assign \new_[31524]_  = ~A233 & \new_[31523]_ ;
  assign \new_[31527]_  = ~A269 & ~A268;
  assign \new_[31530]_  = A300 & A299;
  assign \new_[31531]_  = \new_[31530]_  & \new_[31527]_ ;
  assign \new_[31532]_  = \new_[31531]_  & \new_[31524]_ ;
  assign \new_[31536]_  = ~A201 & A167;
  assign \new_[31537]_  = A168 & \new_[31536]_ ;
  assign \new_[31541]_  = ~A232 & ~A203;
  assign \new_[31542]_  = ~A202 & \new_[31541]_ ;
  assign \new_[31543]_  = \new_[31542]_  & \new_[31537]_ ;
  assign \new_[31547]_  = ~A267 & ~A235;
  assign \new_[31548]_  = ~A233 & \new_[31547]_ ;
  assign \new_[31551]_  = ~A269 & ~A268;
  assign \new_[31554]_  = A300 & A298;
  assign \new_[31555]_  = \new_[31554]_  & \new_[31551]_ ;
  assign \new_[31556]_  = \new_[31555]_  & \new_[31548]_ ;
  assign \new_[31560]_  = ~A201 & A167;
  assign \new_[31561]_  = A168 & \new_[31560]_ ;
  assign \new_[31565]_  = ~A232 & ~A203;
  assign \new_[31566]_  = ~A202 & \new_[31565]_ ;
  assign \new_[31567]_  = \new_[31566]_  & \new_[31561]_ ;
  assign \new_[31571]_  = A265 & ~A235;
  assign \new_[31572]_  = ~A233 & \new_[31571]_ ;
  assign \new_[31575]_  = ~A267 & A266;
  assign \new_[31578]_  = A301 & ~A268;
  assign \new_[31579]_  = \new_[31578]_  & \new_[31575]_ ;
  assign \new_[31580]_  = \new_[31579]_  & \new_[31572]_ ;
  assign \new_[31584]_  = ~A201 & A167;
  assign \new_[31585]_  = A168 & \new_[31584]_ ;
  assign \new_[31589]_  = ~A232 & ~A203;
  assign \new_[31590]_  = ~A202 & \new_[31589]_ ;
  assign \new_[31591]_  = \new_[31590]_  & \new_[31585]_ ;
  assign \new_[31595]_  = ~A265 & ~A235;
  assign \new_[31596]_  = ~A233 & \new_[31595]_ ;
  assign \new_[31599]_  = ~A268 & ~A266;
  assign \new_[31602]_  = A300 & A299;
  assign \new_[31603]_  = \new_[31602]_  & \new_[31599]_ ;
  assign \new_[31604]_  = \new_[31603]_  & \new_[31596]_ ;
  assign \new_[31608]_  = ~A201 & A167;
  assign \new_[31609]_  = A168 & \new_[31608]_ ;
  assign \new_[31613]_  = ~A232 & ~A203;
  assign \new_[31614]_  = ~A202 & \new_[31613]_ ;
  assign \new_[31615]_  = \new_[31614]_  & \new_[31609]_ ;
  assign \new_[31619]_  = ~A265 & ~A235;
  assign \new_[31620]_  = ~A233 & \new_[31619]_ ;
  assign \new_[31623]_  = ~A268 & ~A266;
  assign \new_[31626]_  = A300 & A298;
  assign \new_[31627]_  = \new_[31626]_  & \new_[31623]_ ;
  assign \new_[31628]_  = \new_[31627]_  & \new_[31620]_ ;
  assign \new_[31632]_  = A199 & A167;
  assign \new_[31633]_  = A168 & \new_[31632]_ ;
  assign \new_[31637]_  = ~A202 & ~A201;
  assign \new_[31638]_  = A200 & \new_[31637]_ ;
  assign \new_[31639]_  = \new_[31638]_  & \new_[31633]_ ;
  assign \new_[31643]_  = ~A236 & ~A235;
  assign \new_[31644]_  = ~A234 & \new_[31643]_ ;
  assign \new_[31647]_  = ~A268 & ~A267;
  assign \new_[31650]_  = A301 & ~A269;
  assign \new_[31651]_  = \new_[31650]_  & \new_[31647]_ ;
  assign \new_[31652]_  = \new_[31651]_  & \new_[31644]_ ;
  assign \new_[31656]_  = A199 & A167;
  assign \new_[31657]_  = A168 & \new_[31656]_ ;
  assign \new_[31661]_  = ~A202 & ~A201;
  assign \new_[31662]_  = A200 & \new_[31661]_ ;
  assign \new_[31663]_  = \new_[31662]_  & \new_[31657]_ ;
  assign \new_[31667]_  = ~A236 & ~A235;
  assign \new_[31668]_  = ~A234 & \new_[31667]_ ;
  assign \new_[31671]_  = ~A266 & ~A265;
  assign \new_[31674]_  = A301 & ~A268;
  assign \new_[31675]_  = \new_[31674]_  & \new_[31671]_ ;
  assign \new_[31676]_  = \new_[31675]_  & \new_[31668]_ ;
  assign \new_[31680]_  = A199 & A167;
  assign \new_[31681]_  = A168 & \new_[31680]_ ;
  assign \new_[31685]_  = ~A202 & ~A201;
  assign \new_[31686]_  = A200 & \new_[31685]_ ;
  assign \new_[31687]_  = \new_[31686]_  & \new_[31681]_ ;
  assign \new_[31691]_  = A236 & A233;
  assign \new_[31692]_  = ~A232 & \new_[31691]_ ;
  assign \new_[31695]_  = A299 & A298;
  assign \new_[31698]_  = ~A301 & ~A300;
  assign \new_[31699]_  = \new_[31698]_  & \new_[31695]_ ;
  assign \new_[31700]_  = \new_[31699]_  & \new_[31692]_ ;
  assign \new_[31704]_  = A199 & A167;
  assign \new_[31705]_  = A168 & \new_[31704]_ ;
  assign \new_[31709]_  = ~A202 & ~A201;
  assign \new_[31710]_  = A200 & \new_[31709]_ ;
  assign \new_[31711]_  = \new_[31710]_  & \new_[31705]_ ;
  assign \new_[31715]_  = A236 & ~A233;
  assign \new_[31716]_  = A232 & \new_[31715]_ ;
  assign \new_[31719]_  = A299 & A298;
  assign \new_[31722]_  = ~A301 & ~A300;
  assign \new_[31723]_  = \new_[31722]_  & \new_[31719]_ ;
  assign \new_[31724]_  = \new_[31723]_  & \new_[31716]_ ;
  assign \new_[31728]_  = A199 & A167;
  assign \new_[31729]_  = A168 & \new_[31728]_ ;
  assign \new_[31733]_  = ~A202 & ~A201;
  assign \new_[31734]_  = A200 & \new_[31733]_ ;
  assign \new_[31735]_  = \new_[31734]_  & \new_[31729]_ ;
  assign \new_[31739]_  = ~A235 & ~A233;
  assign \new_[31740]_  = ~A232 & \new_[31739]_ ;
  assign \new_[31743]_  = ~A268 & ~A267;
  assign \new_[31746]_  = A301 & ~A269;
  assign \new_[31747]_  = \new_[31746]_  & \new_[31743]_ ;
  assign \new_[31748]_  = \new_[31747]_  & \new_[31740]_ ;
  assign \new_[31752]_  = A199 & A167;
  assign \new_[31753]_  = A168 & \new_[31752]_ ;
  assign \new_[31757]_  = ~A202 & ~A201;
  assign \new_[31758]_  = A200 & \new_[31757]_ ;
  assign \new_[31759]_  = \new_[31758]_  & \new_[31753]_ ;
  assign \new_[31763]_  = ~A235 & ~A233;
  assign \new_[31764]_  = ~A232 & \new_[31763]_ ;
  assign \new_[31767]_  = ~A266 & ~A265;
  assign \new_[31770]_  = A301 & ~A268;
  assign \new_[31771]_  = \new_[31770]_  & \new_[31767]_ ;
  assign \new_[31772]_  = \new_[31771]_  & \new_[31764]_ ;
  assign \new_[31776]_  = ~A199 & A167;
  assign \new_[31777]_  = A168 & \new_[31776]_ ;
  assign \new_[31781]_  = ~A234 & ~A202;
  assign \new_[31782]_  = ~A200 & \new_[31781]_ ;
  assign \new_[31783]_  = \new_[31782]_  & \new_[31777]_ ;
  assign \new_[31787]_  = ~A267 & ~A236;
  assign \new_[31788]_  = ~A235 & \new_[31787]_ ;
  assign \new_[31791]_  = ~A269 & ~A268;
  assign \new_[31794]_  = A300 & A299;
  assign \new_[31795]_  = \new_[31794]_  & \new_[31791]_ ;
  assign \new_[31796]_  = \new_[31795]_  & \new_[31788]_ ;
  assign \new_[31800]_  = ~A199 & A167;
  assign \new_[31801]_  = A168 & \new_[31800]_ ;
  assign \new_[31805]_  = ~A234 & ~A202;
  assign \new_[31806]_  = ~A200 & \new_[31805]_ ;
  assign \new_[31807]_  = \new_[31806]_  & \new_[31801]_ ;
  assign \new_[31811]_  = ~A267 & ~A236;
  assign \new_[31812]_  = ~A235 & \new_[31811]_ ;
  assign \new_[31815]_  = ~A269 & ~A268;
  assign \new_[31818]_  = A300 & A298;
  assign \new_[31819]_  = \new_[31818]_  & \new_[31815]_ ;
  assign \new_[31820]_  = \new_[31819]_  & \new_[31812]_ ;
  assign \new_[31824]_  = ~A199 & A167;
  assign \new_[31825]_  = A168 & \new_[31824]_ ;
  assign \new_[31829]_  = ~A234 & ~A202;
  assign \new_[31830]_  = ~A200 & \new_[31829]_ ;
  assign \new_[31831]_  = \new_[31830]_  & \new_[31825]_ ;
  assign \new_[31835]_  = A265 & ~A236;
  assign \new_[31836]_  = ~A235 & \new_[31835]_ ;
  assign \new_[31839]_  = ~A267 & A266;
  assign \new_[31842]_  = A301 & ~A268;
  assign \new_[31843]_  = \new_[31842]_  & \new_[31839]_ ;
  assign \new_[31844]_  = \new_[31843]_  & \new_[31836]_ ;
  assign \new_[31848]_  = ~A199 & A167;
  assign \new_[31849]_  = A168 & \new_[31848]_ ;
  assign \new_[31853]_  = ~A234 & ~A202;
  assign \new_[31854]_  = ~A200 & \new_[31853]_ ;
  assign \new_[31855]_  = \new_[31854]_  & \new_[31849]_ ;
  assign \new_[31859]_  = ~A265 & ~A236;
  assign \new_[31860]_  = ~A235 & \new_[31859]_ ;
  assign \new_[31863]_  = ~A268 & ~A266;
  assign \new_[31866]_  = A300 & A299;
  assign \new_[31867]_  = \new_[31866]_  & \new_[31863]_ ;
  assign \new_[31868]_  = \new_[31867]_  & \new_[31860]_ ;
  assign \new_[31872]_  = ~A199 & A167;
  assign \new_[31873]_  = A168 & \new_[31872]_ ;
  assign \new_[31877]_  = ~A234 & ~A202;
  assign \new_[31878]_  = ~A200 & \new_[31877]_ ;
  assign \new_[31879]_  = \new_[31878]_  & \new_[31873]_ ;
  assign \new_[31883]_  = ~A265 & ~A236;
  assign \new_[31884]_  = ~A235 & \new_[31883]_ ;
  assign \new_[31887]_  = ~A268 & ~A266;
  assign \new_[31890]_  = A300 & A298;
  assign \new_[31891]_  = \new_[31890]_  & \new_[31887]_ ;
  assign \new_[31892]_  = \new_[31891]_  & \new_[31884]_ ;
  assign \new_[31896]_  = ~A199 & A167;
  assign \new_[31897]_  = A168 & \new_[31896]_ ;
  assign \new_[31901]_  = A232 & ~A202;
  assign \new_[31902]_  = ~A200 & \new_[31901]_ ;
  assign \new_[31903]_  = \new_[31902]_  & \new_[31897]_ ;
  assign \new_[31907]_  = ~A235 & ~A234;
  assign \new_[31908]_  = A233 & \new_[31907]_ ;
  assign \new_[31911]_  = ~A268 & ~A267;
  assign \new_[31914]_  = A301 & ~A269;
  assign \new_[31915]_  = \new_[31914]_  & \new_[31911]_ ;
  assign \new_[31916]_  = \new_[31915]_  & \new_[31908]_ ;
  assign \new_[31920]_  = ~A199 & A167;
  assign \new_[31921]_  = A168 & \new_[31920]_ ;
  assign \new_[31925]_  = A232 & ~A202;
  assign \new_[31926]_  = ~A200 & \new_[31925]_ ;
  assign \new_[31927]_  = \new_[31926]_  & \new_[31921]_ ;
  assign \new_[31931]_  = ~A235 & ~A234;
  assign \new_[31932]_  = A233 & \new_[31931]_ ;
  assign \new_[31935]_  = ~A266 & ~A265;
  assign \new_[31938]_  = A301 & ~A268;
  assign \new_[31939]_  = \new_[31938]_  & \new_[31935]_ ;
  assign \new_[31940]_  = \new_[31939]_  & \new_[31932]_ ;
  assign \new_[31944]_  = ~A199 & A167;
  assign \new_[31945]_  = A168 & \new_[31944]_ ;
  assign \new_[31949]_  = ~A232 & ~A202;
  assign \new_[31950]_  = ~A200 & \new_[31949]_ ;
  assign \new_[31951]_  = \new_[31950]_  & \new_[31945]_ ;
  assign \new_[31955]_  = ~A267 & ~A235;
  assign \new_[31956]_  = ~A233 & \new_[31955]_ ;
  assign \new_[31959]_  = ~A269 & ~A268;
  assign \new_[31962]_  = A300 & A299;
  assign \new_[31963]_  = \new_[31962]_  & \new_[31959]_ ;
  assign \new_[31964]_  = \new_[31963]_  & \new_[31956]_ ;
  assign \new_[31968]_  = ~A199 & A167;
  assign \new_[31969]_  = A168 & \new_[31968]_ ;
  assign \new_[31973]_  = ~A232 & ~A202;
  assign \new_[31974]_  = ~A200 & \new_[31973]_ ;
  assign \new_[31975]_  = \new_[31974]_  & \new_[31969]_ ;
  assign \new_[31979]_  = ~A267 & ~A235;
  assign \new_[31980]_  = ~A233 & \new_[31979]_ ;
  assign \new_[31983]_  = ~A269 & ~A268;
  assign \new_[31986]_  = A300 & A298;
  assign \new_[31987]_  = \new_[31986]_  & \new_[31983]_ ;
  assign \new_[31988]_  = \new_[31987]_  & \new_[31980]_ ;
  assign \new_[31992]_  = ~A199 & A167;
  assign \new_[31993]_  = A168 & \new_[31992]_ ;
  assign \new_[31997]_  = ~A232 & ~A202;
  assign \new_[31998]_  = ~A200 & \new_[31997]_ ;
  assign \new_[31999]_  = \new_[31998]_  & \new_[31993]_ ;
  assign \new_[32003]_  = A265 & ~A235;
  assign \new_[32004]_  = ~A233 & \new_[32003]_ ;
  assign \new_[32007]_  = ~A267 & A266;
  assign \new_[32010]_  = A301 & ~A268;
  assign \new_[32011]_  = \new_[32010]_  & \new_[32007]_ ;
  assign \new_[32012]_  = \new_[32011]_  & \new_[32004]_ ;
  assign \new_[32016]_  = ~A199 & A167;
  assign \new_[32017]_  = A168 & \new_[32016]_ ;
  assign \new_[32021]_  = ~A232 & ~A202;
  assign \new_[32022]_  = ~A200 & \new_[32021]_ ;
  assign \new_[32023]_  = \new_[32022]_  & \new_[32017]_ ;
  assign \new_[32027]_  = ~A265 & ~A235;
  assign \new_[32028]_  = ~A233 & \new_[32027]_ ;
  assign \new_[32031]_  = ~A268 & ~A266;
  assign \new_[32034]_  = A300 & A299;
  assign \new_[32035]_  = \new_[32034]_  & \new_[32031]_ ;
  assign \new_[32036]_  = \new_[32035]_  & \new_[32028]_ ;
  assign \new_[32040]_  = ~A199 & A167;
  assign \new_[32041]_  = A168 & \new_[32040]_ ;
  assign \new_[32045]_  = ~A232 & ~A202;
  assign \new_[32046]_  = ~A200 & \new_[32045]_ ;
  assign \new_[32047]_  = \new_[32046]_  & \new_[32041]_ ;
  assign \new_[32051]_  = ~A265 & ~A235;
  assign \new_[32052]_  = ~A233 & \new_[32051]_ ;
  assign \new_[32055]_  = ~A268 & ~A266;
  assign \new_[32058]_  = A300 & A298;
  assign \new_[32059]_  = \new_[32058]_  & \new_[32055]_ ;
  assign \new_[32060]_  = \new_[32059]_  & \new_[32052]_ ;
  assign \new_[32064]_  = ~A166 & A167;
  assign \new_[32065]_  = A170 & \new_[32064]_ ;
  assign \new_[32069]_  = ~A203 & ~A202;
  assign \new_[32070]_  = ~A201 & \new_[32069]_ ;
  assign \new_[32071]_  = \new_[32070]_  & \new_[32065]_ ;
  assign \new_[32075]_  = ~A236 & ~A235;
  assign \new_[32076]_  = ~A234 & \new_[32075]_ ;
  assign \new_[32079]_  = ~A268 & ~A267;
  assign \new_[32082]_  = A301 & ~A269;
  assign \new_[32083]_  = \new_[32082]_  & \new_[32079]_ ;
  assign \new_[32084]_  = \new_[32083]_  & \new_[32076]_ ;
  assign \new_[32088]_  = ~A166 & A167;
  assign \new_[32089]_  = A170 & \new_[32088]_ ;
  assign \new_[32093]_  = ~A203 & ~A202;
  assign \new_[32094]_  = ~A201 & \new_[32093]_ ;
  assign \new_[32095]_  = \new_[32094]_  & \new_[32089]_ ;
  assign \new_[32099]_  = ~A236 & ~A235;
  assign \new_[32100]_  = ~A234 & \new_[32099]_ ;
  assign \new_[32103]_  = ~A266 & ~A265;
  assign \new_[32106]_  = A301 & ~A268;
  assign \new_[32107]_  = \new_[32106]_  & \new_[32103]_ ;
  assign \new_[32108]_  = \new_[32107]_  & \new_[32100]_ ;
  assign \new_[32112]_  = ~A166 & A167;
  assign \new_[32113]_  = A170 & \new_[32112]_ ;
  assign \new_[32117]_  = ~A203 & ~A202;
  assign \new_[32118]_  = ~A201 & \new_[32117]_ ;
  assign \new_[32119]_  = \new_[32118]_  & \new_[32113]_ ;
  assign \new_[32123]_  = A236 & A233;
  assign \new_[32124]_  = ~A232 & \new_[32123]_ ;
  assign \new_[32127]_  = A299 & A298;
  assign \new_[32130]_  = ~A301 & ~A300;
  assign \new_[32131]_  = \new_[32130]_  & \new_[32127]_ ;
  assign \new_[32132]_  = \new_[32131]_  & \new_[32124]_ ;
  assign \new_[32136]_  = ~A166 & A167;
  assign \new_[32137]_  = A170 & \new_[32136]_ ;
  assign \new_[32141]_  = ~A203 & ~A202;
  assign \new_[32142]_  = ~A201 & \new_[32141]_ ;
  assign \new_[32143]_  = \new_[32142]_  & \new_[32137]_ ;
  assign \new_[32147]_  = A236 & ~A233;
  assign \new_[32148]_  = A232 & \new_[32147]_ ;
  assign \new_[32151]_  = A299 & A298;
  assign \new_[32154]_  = ~A301 & ~A300;
  assign \new_[32155]_  = \new_[32154]_  & \new_[32151]_ ;
  assign \new_[32156]_  = \new_[32155]_  & \new_[32148]_ ;
  assign \new_[32160]_  = ~A166 & A167;
  assign \new_[32161]_  = A170 & \new_[32160]_ ;
  assign \new_[32165]_  = ~A203 & ~A202;
  assign \new_[32166]_  = ~A201 & \new_[32165]_ ;
  assign \new_[32167]_  = \new_[32166]_  & \new_[32161]_ ;
  assign \new_[32171]_  = ~A235 & ~A233;
  assign \new_[32172]_  = ~A232 & \new_[32171]_ ;
  assign \new_[32175]_  = ~A268 & ~A267;
  assign \new_[32178]_  = A301 & ~A269;
  assign \new_[32179]_  = \new_[32178]_  & \new_[32175]_ ;
  assign \new_[32180]_  = \new_[32179]_  & \new_[32172]_ ;
  assign \new_[32184]_  = ~A166 & A167;
  assign \new_[32185]_  = A170 & \new_[32184]_ ;
  assign \new_[32189]_  = ~A203 & ~A202;
  assign \new_[32190]_  = ~A201 & \new_[32189]_ ;
  assign \new_[32191]_  = \new_[32190]_  & \new_[32185]_ ;
  assign \new_[32195]_  = ~A235 & ~A233;
  assign \new_[32196]_  = ~A232 & \new_[32195]_ ;
  assign \new_[32199]_  = ~A266 & ~A265;
  assign \new_[32202]_  = A301 & ~A268;
  assign \new_[32203]_  = \new_[32202]_  & \new_[32199]_ ;
  assign \new_[32204]_  = \new_[32203]_  & \new_[32196]_ ;
  assign \new_[32208]_  = ~A166 & A167;
  assign \new_[32209]_  = A170 & \new_[32208]_ ;
  assign \new_[32213]_  = ~A201 & A200;
  assign \new_[32214]_  = A199 & \new_[32213]_ ;
  assign \new_[32215]_  = \new_[32214]_  & \new_[32209]_ ;
  assign \new_[32219]_  = A234 & A232;
  assign \new_[32220]_  = ~A202 & \new_[32219]_ ;
  assign \new_[32223]_  = A299 & A298;
  assign \new_[32226]_  = ~A301 & ~A300;
  assign \new_[32227]_  = \new_[32226]_  & \new_[32223]_ ;
  assign \new_[32228]_  = \new_[32227]_  & \new_[32220]_ ;
  assign \new_[32232]_  = ~A166 & A167;
  assign \new_[32233]_  = A170 & \new_[32232]_ ;
  assign \new_[32237]_  = ~A201 & A200;
  assign \new_[32238]_  = A199 & \new_[32237]_ ;
  assign \new_[32239]_  = \new_[32238]_  & \new_[32233]_ ;
  assign \new_[32243]_  = A234 & A233;
  assign \new_[32244]_  = ~A202 & \new_[32243]_ ;
  assign \new_[32247]_  = A299 & A298;
  assign \new_[32250]_  = ~A301 & ~A300;
  assign \new_[32251]_  = \new_[32250]_  & \new_[32247]_ ;
  assign \new_[32252]_  = \new_[32251]_  & \new_[32244]_ ;
  assign \new_[32256]_  = ~A166 & A167;
  assign \new_[32257]_  = A170 & \new_[32256]_ ;
  assign \new_[32261]_  = ~A201 & A200;
  assign \new_[32262]_  = A199 & \new_[32261]_ ;
  assign \new_[32263]_  = \new_[32262]_  & \new_[32257]_ ;
  assign \new_[32267]_  = A233 & ~A232;
  assign \new_[32268]_  = ~A202 & \new_[32267]_ ;
  assign \new_[32271]_  = ~A300 & A236;
  assign \new_[32274]_  = ~A302 & ~A301;
  assign \new_[32275]_  = \new_[32274]_  & \new_[32271]_ ;
  assign \new_[32276]_  = \new_[32275]_  & \new_[32268]_ ;
  assign \new_[32280]_  = ~A166 & A167;
  assign \new_[32281]_  = A170 & \new_[32280]_ ;
  assign \new_[32285]_  = ~A201 & A200;
  assign \new_[32286]_  = A199 & \new_[32285]_ ;
  assign \new_[32287]_  = \new_[32286]_  & \new_[32281]_ ;
  assign \new_[32291]_  = A233 & ~A232;
  assign \new_[32292]_  = ~A202 & \new_[32291]_ ;
  assign \new_[32295]_  = ~A298 & A236;
  assign \new_[32298]_  = ~A301 & ~A299;
  assign \new_[32299]_  = \new_[32298]_  & \new_[32295]_ ;
  assign \new_[32300]_  = \new_[32299]_  & \new_[32292]_ ;
  assign \new_[32304]_  = ~A166 & A167;
  assign \new_[32305]_  = A170 & \new_[32304]_ ;
  assign \new_[32309]_  = ~A201 & A200;
  assign \new_[32310]_  = A199 & \new_[32309]_ ;
  assign \new_[32311]_  = \new_[32310]_  & \new_[32305]_ ;
  assign \new_[32315]_  = A233 & ~A232;
  assign \new_[32316]_  = ~A202 & \new_[32315]_ ;
  assign \new_[32319]_  = ~A265 & A236;
  assign \new_[32322]_  = A269 & A266;
  assign \new_[32323]_  = \new_[32322]_  & \new_[32319]_ ;
  assign \new_[32324]_  = \new_[32323]_  & \new_[32316]_ ;
  assign \new_[32328]_  = ~A166 & A167;
  assign \new_[32329]_  = A170 & \new_[32328]_ ;
  assign \new_[32333]_  = ~A201 & A200;
  assign \new_[32334]_  = A199 & \new_[32333]_ ;
  assign \new_[32335]_  = \new_[32334]_  & \new_[32329]_ ;
  assign \new_[32339]_  = A233 & ~A232;
  assign \new_[32340]_  = ~A202 & \new_[32339]_ ;
  assign \new_[32343]_  = A265 & A236;
  assign \new_[32346]_  = A269 & ~A266;
  assign \new_[32347]_  = \new_[32346]_  & \new_[32343]_ ;
  assign \new_[32348]_  = \new_[32347]_  & \new_[32340]_ ;
  assign \new_[32352]_  = ~A166 & A167;
  assign \new_[32353]_  = A170 & \new_[32352]_ ;
  assign \new_[32357]_  = ~A201 & A200;
  assign \new_[32358]_  = A199 & \new_[32357]_ ;
  assign \new_[32359]_  = \new_[32358]_  & \new_[32353]_ ;
  assign \new_[32363]_  = ~A233 & A232;
  assign \new_[32364]_  = ~A202 & \new_[32363]_ ;
  assign \new_[32367]_  = ~A300 & A236;
  assign \new_[32370]_  = ~A302 & ~A301;
  assign \new_[32371]_  = \new_[32370]_  & \new_[32367]_ ;
  assign \new_[32372]_  = \new_[32371]_  & \new_[32364]_ ;
  assign \new_[32376]_  = ~A166 & A167;
  assign \new_[32377]_  = A170 & \new_[32376]_ ;
  assign \new_[32381]_  = ~A201 & A200;
  assign \new_[32382]_  = A199 & \new_[32381]_ ;
  assign \new_[32383]_  = \new_[32382]_  & \new_[32377]_ ;
  assign \new_[32387]_  = ~A233 & A232;
  assign \new_[32388]_  = ~A202 & \new_[32387]_ ;
  assign \new_[32391]_  = ~A298 & A236;
  assign \new_[32394]_  = ~A301 & ~A299;
  assign \new_[32395]_  = \new_[32394]_  & \new_[32391]_ ;
  assign \new_[32396]_  = \new_[32395]_  & \new_[32388]_ ;
  assign \new_[32400]_  = ~A166 & A167;
  assign \new_[32401]_  = A170 & \new_[32400]_ ;
  assign \new_[32405]_  = ~A201 & A200;
  assign \new_[32406]_  = A199 & \new_[32405]_ ;
  assign \new_[32407]_  = \new_[32406]_  & \new_[32401]_ ;
  assign \new_[32411]_  = ~A233 & A232;
  assign \new_[32412]_  = ~A202 & \new_[32411]_ ;
  assign \new_[32415]_  = ~A265 & A236;
  assign \new_[32418]_  = A269 & A266;
  assign \new_[32419]_  = \new_[32418]_  & \new_[32415]_ ;
  assign \new_[32420]_  = \new_[32419]_  & \new_[32412]_ ;
  assign \new_[32424]_  = ~A166 & A167;
  assign \new_[32425]_  = A170 & \new_[32424]_ ;
  assign \new_[32429]_  = ~A201 & A200;
  assign \new_[32430]_  = A199 & \new_[32429]_ ;
  assign \new_[32431]_  = \new_[32430]_  & \new_[32425]_ ;
  assign \new_[32435]_  = ~A233 & A232;
  assign \new_[32436]_  = ~A202 & \new_[32435]_ ;
  assign \new_[32439]_  = A265 & A236;
  assign \new_[32442]_  = A269 & ~A266;
  assign \new_[32443]_  = \new_[32442]_  & \new_[32439]_ ;
  assign \new_[32444]_  = \new_[32443]_  & \new_[32436]_ ;
  assign \new_[32448]_  = ~A166 & A167;
  assign \new_[32449]_  = A170 & \new_[32448]_ ;
  assign \new_[32453]_  = ~A202 & ~A200;
  assign \new_[32454]_  = ~A199 & \new_[32453]_ ;
  assign \new_[32455]_  = \new_[32454]_  & \new_[32449]_ ;
  assign \new_[32459]_  = ~A236 & ~A235;
  assign \new_[32460]_  = ~A234 & \new_[32459]_ ;
  assign \new_[32463]_  = ~A268 & ~A267;
  assign \new_[32466]_  = A301 & ~A269;
  assign \new_[32467]_  = \new_[32466]_  & \new_[32463]_ ;
  assign \new_[32468]_  = \new_[32467]_  & \new_[32460]_ ;
  assign \new_[32472]_  = ~A166 & A167;
  assign \new_[32473]_  = A170 & \new_[32472]_ ;
  assign \new_[32477]_  = ~A202 & ~A200;
  assign \new_[32478]_  = ~A199 & \new_[32477]_ ;
  assign \new_[32479]_  = \new_[32478]_  & \new_[32473]_ ;
  assign \new_[32483]_  = ~A236 & ~A235;
  assign \new_[32484]_  = ~A234 & \new_[32483]_ ;
  assign \new_[32487]_  = ~A266 & ~A265;
  assign \new_[32490]_  = A301 & ~A268;
  assign \new_[32491]_  = \new_[32490]_  & \new_[32487]_ ;
  assign \new_[32492]_  = \new_[32491]_  & \new_[32484]_ ;
  assign \new_[32496]_  = ~A166 & A167;
  assign \new_[32497]_  = A170 & \new_[32496]_ ;
  assign \new_[32501]_  = ~A202 & ~A200;
  assign \new_[32502]_  = ~A199 & \new_[32501]_ ;
  assign \new_[32503]_  = \new_[32502]_  & \new_[32497]_ ;
  assign \new_[32507]_  = A236 & A233;
  assign \new_[32508]_  = ~A232 & \new_[32507]_ ;
  assign \new_[32511]_  = A299 & A298;
  assign \new_[32514]_  = ~A301 & ~A300;
  assign \new_[32515]_  = \new_[32514]_  & \new_[32511]_ ;
  assign \new_[32516]_  = \new_[32515]_  & \new_[32508]_ ;
  assign \new_[32520]_  = ~A166 & A167;
  assign \new_[32521]_  = A170 & \new_[32520]_ ;
  assign \new_[32525]_  = ~A202 & ~A200;
  assign \new_[32526]_  = ~A199 & \new_[32525]_ ;
  assign \new_[32527]_  = \new_[32526]_  & \new_[32521]_ ;
  assign \new_[32531]_  = A236 & ~A233;
  assign \new_[32532]_  = A232 & \new_[32531]_ ;
  assign \new_[32535]_  = A299 & A298;
  assign \new_[32538]_  = ~A301 & ~A300;
  assign \new_[32539]_  = \new_[32538]_  & \new_[32535]_ ;
  assign \new_[32540]_  = \new_[32539]_  & \new_[32532]_ ;
  assign \new_[32544]_  = ~A166 & A167;
  assign \new_[32545]_  = A170 & \new_[32544]_ ;
  assign \new_[32549]_  = ~A202 & ~A200;
  assign \new_[32550]_  = ~A199 & \new_[32549]_ ;
  assign \new_[32551]_  = \new_[32550]_  & \new_[32545]_ ;
  assign \new_[32555]_  = ~A235 & ~A233;
  assign \new_[32556]_  = ~A232 & \new_[32555]_ ;
  assign \new_[32559]_  = ~A268 & ~A267;
  assign \new_[32562]_  = A301 & ~A269;
  assign \new_[32563]_  = \new_[32562]_  & \new_[32559]_ ;
  assign \new_[32564]_  = \new_[32563]_  & \new_[32556]_ ;
  assign \new_[32568]_  = ~A166 & A167;
  assign \new_[32569]_  = A170 & \new_[32568]_ ;
  assign \new_[32573]_  = ~A202 & ~A200;
  assign \new_[32574]_  = ~A199 & \new_[32573]_ ;
  assign \new_[32575]_  = \new_[32574]_  & \new_[32569]_ ;
  assign \new_[32579]_  = ~A235 & ~A233;
  assign \new_[32580]_  = ~A232 & \new_[32579]_ ;
  assign \new_[32583]_  = ~A266 & ~A265;
  assign \new_[32586]_  = A301 & ~A268;
  assign \new_[32587]_  = \new_[32586]_  & \new_[32583]_ ;
  assign \new_[32588]_  = \new_[32587]_  & \new_[32580]_ ;
  assign \new_[32592]_  = A166 & ~A167;
  assign \new_[32593]_  = A170 & \new_[32592]_ ;
  assign \new_[32597]_  = ~A203 & ~A202;
  assign \new_[32598]_  = ~A201 & \new_[32597]_ ;
  assign \new_[32599]_  = \new_[32598]_  & \new_[32593]_ ;
  assign \new_[32603]_  = ~A236 & ~A235;
  assign \new_[32604]_  = ~A234 & \new_[32603]_ ;
  assign \new_[32607]_  = ~A268 & ~A267;
  assign \new_[32610]_  = A301 & ~A269;
  assign \new_[32611]_  = \new_[32610]_  & \new_[32607]_ ;
  assign \new_[32612]_  = \new_[32611]_  & \new_[32604]_ ;
  assign \new_[32616]_  = A166 & ~A167;
  assign \new_[32617]_  = A170 & \new_[32616]_ ;
  assign \new_[32621]_  = ~A203 & ~A202;
  assign \new_[32622]_  = ~A201 & \new_[32621]_ ;
  assign \new_[32623]_  = \new_[32622]_  & \new_[32617]_ ;
  assign \new_[32627]_  = ~A236 & ~A235;
  assign \new_[32628]_  = ~A234 & \new_[32627]_ ;
  assign \new_[32631]_  = ~A266 & ~A265;
  assign \new_[32634]_  = A301 & ~A268;
  assign \new_[32635]_  = \new_[32634]_  & \new_[32631]_ ;
  assign \new_[32636]_  = \new_[32635]_  & \new_[32628]_ ;
  assign \new_[32640]_  = A166 & ~A167;
  assign \new_[32641]_  = A170 & \new_[32640]_ ;
  assign \new_[32645]_  = ~A203 & ~A202;
  assign \new_[32646]_  = ~A201 & \new_[32645]_ ;
  assign \new_[32647]_  = \new_[32646]_  & \new_[32641]_ ;
  assign \new_[32651]_  = A236 & A233;
  assign \new_[32652]_  = ~A232 & \new_[32651]_ ;
  assign \new_[32655]_  = A299 & A298;
  assign \new_[32658]_  = ~A301 & ~A300;
  assign \new_[32659]_  = \new_[32658]_  & \new_[32655]_ ;
  assign \new_[32660]_  = \new_[32659]_  & \new_[32652]_ ;
  assign \new_[32664]_  = A166 & ~A167;
  assign \new_[32665]_  = A170 & \new_[32664]_ ;
  assign \new_[32669]_  = ~A203 & ~A202;
  assign \new_[32670]_  = ~A201 & \new_[32669]_ ;
  assign \new_[32671]_  = \new_[32670]_  & \new_[32665]_ ;
  assign \new_[32675]_  = A236 & ~A233;
  assign \new_[32676]_  = A232 & \new_[32675]_ ;
  assign \new_[32679]_  = A299 & A298;
  assign \new_[32682]_  = ~A301 & ~A300;
  assign \new_[32683]_  = \new_[32682]_  & \new_[32679]_ ;
  assign \new_[32684]_  = \new_[32683]_  & \new_[32676]_ ;
  assign \new_[32688]_  = A166 & ~A167;
  assign \new_[32689]_  = A170 & \new_[32688]_ ;
  assign \new_[32693]_  = ~A203 & ~A202;
  assign \new_[32694]_  = ~A201 & \new_[32693]_ ;
  assign \new_[32695]_  = \new_[32694]_  & \new_[32689]_ ;
  assign \new_[32699]_  = ~A235 & ~A233;
  assign \new_[32700]_  = ~A232 & \new_[32699]_ ;
  assign \new_[32703]_  = ~A268 & ~A267;
  assign \new_[32706]_  = A301 & ~A269;
  assign \new_[32707]_  = \new_[32706]_  & \new_[32703]_ ;
  assign \new_[32708]_  = \new_[32707]_  & \new_[32700]_ ;
  assign \new_[32712]_  = A166 & ~A167;
  assign \new_[32713]_  = A170 & \new_[32712]_ ;
  assign \new_[32717]_  = ~A203 & ~A202;
  assign \new_[32718]_  = ~A201 & \new_[32717]_ ;
  assign \new_[32719]_  = \new_[32718]_  & \new_[32713]_ ;
  assign \new_[32723]_  = ~A235 & ~A233;
  assign \new_[32724]_  = ~A232 & \new_[32723]_ ;
  assign \new_[32727]_  = ~A266 & ~A265;
  assign \new_[32730]_  = A301 & ~A268;
  assign \new_[32731]_  = \new_[32730]_  & \new_[32727]_ ;
  assign \new_[32732]_  = \new_[32731]_  & \new_[32724]_ ;
  assign \new_[32736]_  = A166 & ~A167;
  assign \new_[32737]_  = A170 & \new_[32736]_ ;
  assign \new_[32741]_  = ~A201 & A200;
  assign \new_[32742]_  = A199 & \new_[32741]_ ;
  assign \new_[32743]_  = \new_[32742]_  & \new_[32737]_ ;
  assign \new_[32747]_  = A234 & A232;
  assign \new_[32748]_  = ~A202 & \new_[32747]_ ;
  assign \new_[32751]_  = A299 & A298;
  assign \new_[32754]_  = ~A301 & ~A300;
  assign \new_[32755]_  = \new_[32754]_  & \new_[32751]_ ;
  assign \new_[32756]_  = \new_[32755]_  & \new_[32748]_ ;
  assign \new_[32760]_  = A166 & ~A167;
  assign \new_[32761]_  = A170 & \new_[32760]_ ;
  assign \new_[32765]_  = ~A201 & A200;
  assign \new_[32766]_  = A199 & \new_[32765]_ ;
  assign \new_[32767]_  = \new_[32766]_  & \new_[32761]_ ;
  assign \new_[32771]_  = A234 & A233;
  assign \new_[32772]_  = ~A202 & \new_[32771]_ ;
  assign \new_[32775]_  = A299 & A298;
  assign \new_[32778]_  = ~A301 & ~A300;
  assign \new_[32779]_  = \new_[32778]_  & \new_[32775]_ ;
  assign \new_[32780]_  = \new_[32779]_  & \new_[32772]_ ;
  assign \new_[32784]_  = A166 & ~A167;
  assign \new_[32785]_  = A170 & \new_[32784]_ ;
  assign \new_[32789]_  = ~A201 & A200;
  assign \new_[32790]_  = A199 & \new_[32789]_ ;
  assign \new_[32791]_  = \new_[32790]_  & \new_[32785]_ ;
  assign \new_[32795]_  = A233 & ~A232;
  assign \new_[32796]_  = ~A202 & \new_[32795]_ ;
  assign \new_[32799]_  = ~A300 & A236;
  assign \new_[32802]_  = ~A302 & ~A301;
  assign \new_[32803]_  = \new_[32802]_  & \new_[32799]_ ;
  assign \new_[32804]_  = \new_[32803]_  & \new_[32796]_ ;
  assign \new_[32808]_  = A166 & ~A167;
  assign \new_[32809]_  = A170 & \new_[32808]_ ;
  assign \new_[32813]_  = ~A201 & A200;
  assign \new_[32814]_  = A199 & \new_[32813]_ ;
  assign \new_[32815]_  = \new_[32814]_  & \new_[32809]_ ;
  assign \new_[32819]_  = A233 & ~A232;
  assign \new_[32820]_  = ~A202 & \new_[32819]_ ;
  assign \new_[32823]_  = ~A298 & A236;
  assign \new_[32826]_  = ~A301 & ~A299;
  assign \new_[32827]_  = \new_[32826]_  & \new_[32823]_ ;
  assign \new_[32828]_  = \new_[32827]_  & \new_[32820]_ ;
  assign \new_[32832]_  = A166 & ~A167;
  assign \new_[32833]_  = A170 & \new_[32832]_ ;
  assign \new_[32837]_  = ~A201 & A200;
  assign \new_[32838]_  = A199 & \new_[32837]_ ;
  assign \new_[32839]_  = \new_[32838]_  & \new_[32833]_ ;
  assign \new_[32843]_  = A233 & ~A232;
  assign \new_[32844]_  = ~A202 & \new_[32843]_ ;
  assign \new_[32847]_  = ~A265 & A236;
  assign \new_[32850]_  = A269 & A266;
  assign \new_[32851]_  = \new_[32850]_  & \new_[32847]_ ;
  assign \new_[32852]_  = \new_[32851]_  & \new_[32844]_ ;
  assign \new_[32856]_  = A166 & ~A167;
  assign \new_[32857]_  = A170 & \new_[32856]_ ;
  assign \new_[32861]_  = ~A201 & A200;
  assign \new_[32862]_  = A199 & \new_[32861]_ ;
  assign \new_[32863]_  = \new_[32862]_  & \new_[32857]_ ;
  assign \new_[32867]_  = A233 & ~A232;
  assign \new_[32868]_  = ~A202 & \new_[32867]_ ;
  assign \new_[32871]_  = A265 & A236;
  assign \new_[32874]_  = A269 & ~A266;
  assign \new_[32875]_  = \new_[32874]_  & \new_[32871]_ ;
  assign \new_[32876]_  = \new_[32875]_  & \new_[32868]_ ;
  assign \new_[32880]_  = A166 & ~A167;
  assign \new_[32881]_  = A170 & \new_[32880]_ ;
  assign \new_[32885]_  = ~A201 & A200;
  assign \new_[32886]_  = A199 & \new_[32885]_ ;
  assign \new_[32887]_  = \new_[32886]_  & \new_[32881]_ ;
  assign \new_[32891]_  = ~A233 & A232;
  assign \new_[32892]_  = ~A202 & \new_[32891]_ ;
  assign \new_[32895]_  = ~A300 & A236;
  assign \new_[32898]_  = ~A302 & ~A301;
  assign \new_[32899]_  = \new_[32898]_  & \new_[32895]_ ;
  assign \new_[32900]_  = \new_[32899]_  & \new_[32892]_ ;
  assign \new_[32904]_  = A166 & ~A167;
  assign \new_[32905]_  = A170 & \new_[32904]_ ;
  assign \new_[32909]_  = ~A201 & A200;
  assign \new_[32910]_  = A199 & \new_[32909]_ ;
  assign \new_[32911]_  = \new_[32910]_  & \new_[32905]_ ;
  assign \new_[32915]_  = ~A233 & A232;
  assign \new_[32916]_  = ~A202 & \new_[32915]_ ;
  assign \new_[32919]_  = ~A298 & A236;
  assign \new_[32922]_  = ~A301 & ~A299;
  assign \new_[32923]_  = \new_[32922]_  & \new_[32919]_ ;
  assign \new_[32924]_  = \new_[32923]_  & \new_[32916]_ ;
  assign \new_[32928]_  = A166 & ~A167;
  assign \new_[32929]_  = A170 & \new_[32928]_ ;
  assign \new_[32933]_  = ~A201 & A200;
  assign \new_[32934]_  = A199 & \new_[32933]_ ;
  assign \new_[32935]_  = \new_[32934]_  & \new_[32929]_ ;
  assign \new_[32939]_  = ~A233 & A232;
  assign \new_[32940]_  = ~A202 & \new_[32939]_ ;
  assign \new_[32943]_  = ~A265 & A236;
  assign \new_[32946]_  = A269 & A266;
  assign \new_[32947]_  = \new_[32946]_  & \new_[32943]_ ;
  assign \new_[32948]_  = \new_[32947]_  & \new_[32940]_ ;
  assign \new_[32952]_  = A166 & ~A167;
  assign \new_[32953]_  = A170 & \new_[32952]_ ;
  assign \new_[32957]_  = ~A201 & A200;
  assign \new_[32958]_  = A199 & \new_[32957]_ ;
  assign \new_[32959]_  = \new_[32958]_  & \new_[32953]_ ;
  assign \new_[32963]_  = ~A233 & A232;
  assign \new_[32964]_  = ~A202 & \new_[32963]_ ;
  assign \new_[32967]_  = A265 & A236;
  assign \new_[32970]_  = A269 & ~A266;
  assign \new_[32971]_  = \new_[32970]_  & \new_[32967]_ ;
  assign \new_[32972]_  = \new_[32971]_  & \new_[32964]_ ;
  assign \new_[32976]_  = A166 & ~A167;
  assign \new_[32977]_  = A170 & \new_[32976]_ ;
  assign \new_[32981]_  = ~A202 & ~A200;
  assign \new_[32982]_  = ~A199 & \new_[32981]_ ;
  assign \new_[32983]_  = \new_[32982]_  & \new_[32977]_ ;
  assign \new_[32987]_  = ~A236 & ~A235;
  assign \new_[32988]_  = ~A234 & \new_[32987]_ ;
  assign \new_[32991]_  = ~A268 & ~A267;
  assign \new_[32994]_  = A301 & ~A269;
  assign \new_[32995]_  = \new_[32994]_  & \new_[32991]_ ;
  assign \new_[32996]_  = \new_[32995]_  & \new_[32988]_ ;
  assign \new_[33000]_  = A166 & ~A167;
  assign \new_[33001]_  = A170 & \new_[33000]_ ;
  assign \new_[33005]_  = ~A202 & ~A200;
  assign \new_[33006]_  = ~A199 & \new_[33005]_ ;
  assign \new_[33007]_  = \new_[33006]_  & \new_[33001]_ ;
  assign \new_[33011]_  = ~A236 & ~A235;
  assign \new_[33012]_  = ~A234 & \new_[33011]_ ;
  assign \new_[33015]_  = ~A266 & ~A265;
  assign \new_[33018]_  = A301 & ~A268;
  assign \new_[33019]_  = \new_[33018]_  & \new_[33015]_ ;
  assign \new_[33020]_  = \new_[33019]_  & \new_[33012]_ ;
  assign \new_[33024]_  = A166 & ~A167;
  assign \new_[33025]_  = A170 & \new_[33024]_ ;
  assign \new_[33029]_  = ~A202 & ~A200;
  assign \new_[33030]_  = ~A199 & \new_[33029]_ ;
  assign \new_[33031]_  = \new_[33030]_  & \new_[33025]_ ;
  assign \new_[33035]_  = A236 & A233;
  assign \new_[33036]_  = ~A232 & \new_[33035]_ ;
  assign \new_[33039]_  = A299 & A298;
  assign \new_[33042]_  = ~A301 & ~A300;
  assign \new_[33043]_  = \new_[33042]_  & \new_[33039]_ ;
  assign \new_[33044]_  = \new_[33043]_  & \new_[33036]_ ;
  assign \new_[33048]_  = A166 & ~A167;
  assign \new_[33049]_  = A170 & \new_[33048]_ ;
  assign \new_[33053]_  = ~A202 & ~A200;
  assign \new_[33054]_  = ~A199 & \new_[33053]_ ;
  assign \new_[33055]_  = \new_[33054]_  & \new_[33049]_ ;
  assign \new_[33059]_  = A236 & ~A233;
  assign \new_[33060]_  = A232 & \new_[33059]_ ;
  assign \new_[33063]_  = A299 & A298;
  assign \new_[33066]_  = ~A301 & ~A300;
  assign \new_[33067]_  = \new_[33066]_  & \new_[33063]_ ;
  assign \new_[33068]_  = \new_[33067]_  & \new_[33060]_ ;
  assign \new_[33072]_  = A166 & ~A167;
  assign \new_[33073]_  = A170 & \new_[33072]_ ;
  assign \new_[33077]_  = ~A202 & ~A200;
  assign \new_[33078]_  = ~A199 & \new_[33077]_ ;
  assign \new_[33079]_  = \new_[33078]_  & \new_[33073]_ ;
  assign \new_[33083]_  = ~A235 & ~A233;
  assign \new_[33084]_  = ~A232 & \new_[33083]_ ;
  assign \new_[33087]_  = ~A268 & ~A267;
  assign \new_[33090]_  = A301 & ~A269;
  assign \new_[33091]_  = \new_[33090]_  & \new_[33087]_ ;
  assign \new_[33092]_  = \new_[33091]_  & \new_[33084]_ ;
  assign \new_[33096]_  = A166 & ~A167;
  assign \new_[33097]_  = A170 & \new_[33096]_ ;
  assign \new_[33101]_  = ~A202 & ~A200;
  assign \new_[33102]_  = ~A199 & \new_[33101]_ ;
  assign \new_[33103]_  = \new_[33102]_  & \new_[33097]_ ;
  assign \new_[33107]_  = ~A235 & ~A233;
  assign \new_[33108]_  = ~A232 & \new_[33107]_ ;
  assign \new_[33111]_  = ~A266 & ~A265;
  assign \new_[33114]_  = A301 & ~A268;
  assign \new_[33115]_  = \new_[33114]_  & \new_[33111]_ ;
  assign \new_[33116]_  = \new_[33115]_  & \new_[33108]_ ;
  assign \new_[33120]_  = ~A202 & ~A201;
  assign \new_[33121]_  = A169 & \new_[33120]_ ;
  assign \new_[33125]_  = ~A235 & ~A234;
  assign \new_[33126]_  = ~A203 & \new_[33125]_ ;
  assign \new_[33127]_  = \new_[33126]_  & \new_[33121]_ ;
  assign \new_[33131]_  = ~A268 & ~A267;
  assign \new_[33132]_  = ~A236 & \new_[33131]_ ;
  assign \new_[33135]_  = A298 & ~A269;
  assign \new_[33138]_  = A302 & ~A299;
  assign \new_[33139]_  = \new_[33138]_  & \new_[33135]_ ;
  assign \new_[33140]_  = \new_[33139]_  & \new_[33132]_ ;
  assign \new_[33144]_  = ~A202 & ~A201;
  assign \new_[33145]_  = A169 & \new_[33144]_ ;
  assign \new_[33149]_  = ~A235 & ~A234;
  assign \new_[33150]_  = ~A203 & \new_[33149]_ ;
  assign \new_[33151]_  = \new_[33150]_  & \new_[33145]_ ;
  assign \new_[33155]_  = ~A268 & ~A267;
  assign \new_[33156]_  = ~A236 & \new_[33155]_ ;
  assign \new_[33159]_  = ~A298 & ~A269;
  assign \new_[33162]_  = A302 & A299;
  assign \new_[33163]_  = \new_[33162]_  & \new_[33159]_ ;
  assign \new_[33164]_  = \new_[33163]_  & \new_[33156]_ ;
  assign \new_[33168]_  = ~A202 & ~A201;
  assign \new_[33169]_  = A169 & \new_[33168]_ ;
  assign \new_[33173]_  = ~A235 & ~A234;
  assign \new_[33174]_  = ~A203 & \new_[33173]_ ;
  assign \new_[33175]_  = \new_[33174]_  & \new_[33169]_ ;
  assign \new_[33179]_  = A266 & A265;
  assign \new_[33180]_  = ~A236 & \new_[33179]_ ;
  assign \new_[33183]_  = ~A268 & ~A267;
  assign \new_[33186]_  = A300 & A299;
  assign \new_[33187]_  = \new_[33186]_  & \new_[33183]_ ;
  assign \new_[33188]_  = \new_[33187]_  & \new_[33180]_ ;
  assign \new_[33192]_  = ~A202 & ~A201;
  assign \new_[33193]_  = A169 & \new_[33192]_ ;
  assign \new_[33197]_  = ~A235 & ~A234;
  assign \new_[33198]_  = ~A203 & \new_[33197]_ ;
  assign \new_[33199]_  = \new_[33198]_  & \new_[33193]_ ;
  assign \new_[33203]_  = A266 & A265;
  assign \new_[33204]_  = ~A236 & \new_[33203]_ ;
  assign \new_[33207]_  = ~A268 & ~A267;
  assign \new_[33210]_  = A300 & A298;
  assign \new_[33211]_  = \new_[33210]_  & \new_[33207]_ ;
  assign \new_[33212]_  = \new_[33211]_  & \new_[33204]_ ;
  assign \new_[33216]_  = ~A202 & ~A201;
  assign \new_[33217]_  = A169 & \new_[33216]_ ;
  assign \new_[33221]_  = ~A235 & ~A234;
  assign \new_[33222]_  = ~A203 & \new_[33221]_ ;
  assign \new_[33223]_  = \new_[33222]_  & \new_[33217]_ ;
  assign \new_[33227]_  = ~A266 & ~A265;
  assign \new_[33228]_  = ~A236 & \new_[33227]_ ;
  assign \new_[33231]_  = A298 & ~A268;
  assign \new_[33234]_  = A302 & ~A299;
  assign \new_[33235]_  = \new_[33234]_  & \new_[33231]_ ;
  assign \new_[33236]_  = \new_[33235]_  & \new_[33228]_ ;
  assign \new_[33240]_  = ~A202 & ~A201;
  assign \new_[33241]_  = A169 & \new_[33240]_ ;
  assign \new_[33245]_  = ~A235 & ~A234;
  assign \new_[33246]_  = ~A203 & \new_[33245]_ ;
  assign \new_[33247]_  = \new_[33246]_  & \new_[33241]_ ;
  assign \new_[33251]_  = ~A266 & ~A265;
  assign \new_[33252]_  = ~A236 & \new_[33251]_ ;
  assign \new_[33255]_  = ~A298 & ~A268;
  assign \new_[33258]_  = A302 & A299;
  assign \new_[33259]_  = \new_[33258]_  & \new_[33255]_ ;
  assign \new_[33260]_  = \new_[33259]_  & \new_[33252]_ ;
  assign \new_[33264]_  = ~A202 & ~A201;
  assign \new_[33265]_  = A169 & \new_[33264]_ ;
  assign \new_[33269]_  = A233 & A232;
  assign \new_[33270]_  = ~A203 & \new_[33269]_ ;
  assign \new_[33271]_  = \new_[33270]_  & \new_[33265]_ ;
  assign \new_[33275]_  = ~A267 & ~A235;
  assign \new_[33276]_  = ~A234 & \new_[33275]_ ;
  assign \new_[33279]_  = ~A269 & ~A268;
  assign \new_[33282]_  = A300 & A299;
  assign \new_[33283]_  = \new_[33282]_  & \new_[33279]_ ;
  assign \new_[33284]_  = \new_[33283]_  & \new_[33276]_ ;
  assign \new_[33288]_  = ~A202 & ~A201;
  assign \new_[33289]_  = A169 & \new_[33288]_ ;
  assign \new_[33293]_  = A233 & A232;
  assign \new_[33294]_  = ~A203 & \new_[33293]_ ;
  assign \new_[33295]_  = \new_[33294]_  & \new_[33289]_ ;
  assign \new_[33299]_  = ~A267 & ~A235;
  assign \new_[33300]_  = ~A234 & \new_[33299]_ ;
  assign \new_[33303]_  = ~A269 & ~A268;
  assign \new_[33306]_  = A300 & A298;
  assign \new_[33307]_  = \new_[33306]_  & \new_[33303]_ ;
  assign \new_[33308]_  = \new_[33307]_  & \new_[33300]_ ;
  assign \new_[33312]_  = ~A202 & ~A201;
  assign \new_[33313]_  = A169 & \new_[33312]_ ;
  assign \new_[33317]_  = A233 & A232;
  assign \new_[33318]_  = ~A203 & \new_[33317]_ ;
  assign \new_[33319]_  = \new_[33318]_  & \new_[33313]_ ;
  assign \new_[33323]_  = A265 & ~A235;
  assign \new_[33324]_  = ~A234 & \new_[33323]_ ;
  assign \new_[33327]_  = ~A267 & A266;
  assign \new_[33330]_  = A301 & ~A268;
  assign \new_[33331]_  = \new_[33330]_  & \new_[33327]_ ;
  assign \new_[33332]_  = \new_[33331]_  & \new_[33324]_ ;
  assign \new_[33336]_  = ~A202 & ~A201;
  assign \new_[33337]_  = A169 & \new_[33336]_ ;
  assign \new_[33341]_  = A233 & A232;
  assign \new_[33342]_  = ~A203 & \new_[33341]_ ;
  assign \new_[33343]_  = \new_[33342]_  & \new_[33337]_ ;
  assign \new_[33347]_  = ~A265 & ~A235;
  assign \new_[33348]_  = ~A234 & \new_[33347]_ ;
  assign \new_[33351]_  = ~A268 & ~A266;
  assign \new_[33354]_  = A300 & A299;
  assign \new_[33355]_  = \new_[33354]_  & \new_[33351]_ ;
  assign \new_[33356]_  = \new_[33355]_  & \new_[33348]_ ;
  assign \new_[33360]_  = ~A202 & ~A201;
  assign \new_[33361]_  = A169 & \new_[33360]_ ;
  assign \new_[33365]_  = A233 & A232;
  assign \new_[33366]_  = ~A203 & \new_[33365]_ ;
  assign \new_[33367]_  = \new_[33366]_  & \new_[33361]_ ;
  assign \new_[33371]_  = ~A265 & ~A235;
  assign \new_[33372]_  = ~A234 & \new_[33371]_ ;
  assign \new_[33375]_  = ~A268 & ~A266;
  assign \new_[33378]_  = A300 & A298;
  assign \new_[33379]_  = \new_[33378]_  & \new_[33375]_ ;
  assign \new_[33380]_  = \new_[33379]_  & \new_[33372]_ ;
  assign \new_[33384]_  = ~A202 & ~A201;
  assign \new_[33385]_  = A169 & \new_[33384]_ ;
  assign \new_[33389]_  = ~A233 & ~A232;
  assign \new_[33390]_  = ~A203 & \new_[33389]_ ;
  assign \new_[33391]_  = \new_[33390]_  & \new_[33385]_ ;
  assign \new_[33395]_  = ~A268 & ~A267;
  assign \new_[33396]_  = ~A235 & \new_[33395]_ ;
  assign \new_[33399]_  = A298 & ~A269;
  assign \new_[33402]_  = A302 & ~A299;
  assign \new_[33403]_  = \new_[33402]_  & \new_[33399]_ ;
  assign \new_[33404]_  = \new_[33403]_  & \new_[33396]_ ;
  assign \new_[33408]_  = ~A202 & ~A201;
  assign \new_[33409]_  = A169 & \new_[33408]_ ;
  assign \new_[33413]_  = ~A233 & ~A232;
  assign \new_[33414]_  = ~A203 & \new_[33413]_ ;
  assign \new_[33415]_  = \new_[33414]_  & \new_[33409]_ ;
  assign \new_[33419]_  = ~A268 & ~A267;
  assign \new_[33420]_  = ~A235 & \new_[33419]_ ;
  assign \new_[33423]_  = ~A298 & ~A269;
  assign \new_[33426]_  = A302 & A299;
  assign \new_[33427]_  = \new_[33426]_  & \new_[33423]_ ;
  assign \new_[33428]_  = \new_[33427]_  & \new_[33420]_ ;
  assign \new_[33432]_  = ~A202 & ~A201;
  assign \new_[33433]_  = A169 & \new_[33432]_ ;
  assign \new_[33437]_  = ~A233 & ~A232;
  assign \new_[33438]_  = ~A203 & \new_[33437]_ ;
  assign \new_[33439]_  = \new_[33438]_  & \new_[33433]_ ;
  assign \new_[33443]_  = A266 & A265;
  assign \new_[33444]_  = ~A235 & \new_[33443]_ ;
  assign \new_[33447]_  = ~A268 & ~A267;
  assign \new_[33450]_  = A300 & A299;
  assign \new_[33451]_  = \new_[33450]_  & \new_[33447]_ ;
  assign \new_[33452]_  = \new_[33451]_  & \new_[33444]_ ;
  assign \new_[33456]_  = ~A202 & ~A201;
  assign \new_[33457]_  = A169 & \new_[33456]_ ;
  assign \new_[33461]_  = ~A233 & ~A232;
  assign \new_[33462]_  = ~A203 & \new_[33461]_ ;
  assign \new_[33463]_  = \new_[33462]_  & \new_[33457]_ ;
  assign \new_[33467]_  = A266 & A265;
  assign \new_[33468]_  = ~A235 & \new_[33467]_ ;
  assign \new_[33471]_  = ~A268 & ~A267;
  assign \new_[33474]_  = A300 & A298;
  assign \new_[33475]_  = \new_[33474]_  & \new_[33471]_ ;
  assign \new_[33476]_  = \new_[33475]_  & \new_[33468]_ ;
  assign \new_[33480]_  = ~A202 & ~A201;
  assign \new_[33481]_  = A169 & \new_[33480]_ ;
  assign \new_[33485]_  = ~A233 & ~A232;
  assign \new_[33486]_  = ~A203 & \new_[33485]_ ;
  assign \new_[33487]_  = \new_[33486]_  & \new_[33481]_ ;
  assign \new_[33491]_  = ~A266 & ~A265;
  assign \new_[33492]_  = ~A235 & \new_[33491]_ ;
  assign \new_[33495]_  = A298 & ~A268;
  assign \new_[33498]_  = A302 & ~A299;
  assign \new_[33499]_  = \new_[33498]_  & \new_[33495]_ ;
  assign \new_[33500]_  = \new_[33499]_  & \new_[33492]_ ;
  assign \new_[33504]_  = ~A202 & ~A201;
  assign \new_[33505]_  = A169 & \new_[33504]_ ;
  assign \new_[33509]_  = ~A233 & ~A232;
  assign \new_[33510]_  = ~A203 & \new_[33509]_ ;
  assign \new_[33511]_  = \new_[33510]_  & \new_[33505]_ ;
  assign \new_[33515]_  = ~A266 & ~A265;
  assign \new_[33516]_  = ~A235 & \new_[33515]_ ;
  assign \new_[33519]_  = ~A298 & ~A268;
  assign \new_[33522]_  = A302 & A299;
  assign \new_[33523]_  = \new_[33522]_  & \new_[33519]_ ;
  assign \new_[33524]_  = \new_[33523]_  & \new_[33516]_ ;
  assign \new_[33528]_  = A200 & A199;
  assign \new_[33529]_  = A169 & \new_[33528]_ ;
  assign \new_[33533]_  = ~A234 & ~A202;
  assign \new_[33534]_  = ~A201 & \new_[33533]_ ;
  assign \new_[33535]_  = \new_[33534]_  & \new_[33529]_ ;
  assign \new_[33539]_  = ~A267 & ~A236;
  assign \new_[33540]_  = ~A235 & \new_[33539]_ ;
  assign \new_[33543]_  = ~A269 & ~A268;
  assign \new_[33546]_  = A300 & A299;
  assign \new_[33547]_  = \new_[33546]_  & \new_[33543]_ ;
  assign \new_[33548]_  = \new_[33547]_  & \new_[33540]_ ;
  assign \new_[33552]_  = A200 & A199;
  assign \new_[33553]_  = A169 & \new_[33552]_ ;
  assign \new_[33557]_  = ~A234 & ~A202;
  assign \new_[33558]_  = ~A201 & \new_[33557]_ ;
  assign \new_[33559]_  = \new_[33558]_  & \new_[33553]_ ;
  assign \new_[33563]_  = ~A267 & ~A236;
  assign \new_[33564]_  = ~A235 & \new_[33563]_ ;
  assign \new_[33567]_  = ~A269 & ~A268;
  assign \new_[33570]_  = A300 & A298;
  assign \new_[33571]_  = \new_[33570]_  & \new_[33567]_ ;
  assign \new_[33572]_  = \new_[33571]_  & \new_[33564]_ ;
  assign \new_[33576]_  = A200 & A199;
  assign \new_[33577]_  = A169 & \new_[33576]_ ;
  assign \new_[33581]_  = ~A234 & ~A202;
  assign \new_[33582]_  = ~A201 & \new_[33581]_ ;
  assign \new_[33583]_  = \new_[33582]_  & \new_[33577]_ ;
  assign \new_[33587]_  = A265 & ~A236;
  assign \new_[33588]_  = ~A235 & \new_[33587]_ ;
  assign \new_[33591]_  = ~A267 & A266;
  assign \new_[33594]_  = A301 & ~A268;
  assign \new_[33595]_  = \new_[33594]_  & \new_[33591]_ ;
  assign \new_[33596]_  = \new_[33595]_  & \new_[33588]_ ;
  assign \new_[33600]_  = A200 & A199;
  assign \new_[33601]_  = A169 & \new_[33600]_ ;
  assign \new_[33605]_  = ~A234 & ~A202;
  assign \new_[33606]_  = ~A201 & \new_[33605]_ ;
  assign \new_[33607]_  = \new_[33606]_  & \new_[33601]_ ;
  assign \new_[33611]_  = ~A265 & ~A236;
  assign \new_[33612]_  = ~A235 & \new_[33611]_ ;
  assign \new_[33615]_  = ~A268 & ~A266;
  assign \new_[33618]_  = A300 & A299;
  assign \new_[33619]_  = \new_[33618]_  & \new_[33615]_ ;
  assign \new_[33620]_  = \new_[33619]_  & \new_[33612]_ ;
  assign \new_[33624]_  = A200 & A199;
  assign \new_[33625]_  = A169 & \new_[33624]_ ;
  assign \new_[33629]_  = ~A234 & ~A202;
  assign \new_[33630]_  = ~A201 & \new_[33629]_ ;
  assign \new_[33631]_  = \new_[33630]_  & \new_[33625]_ ;
  assign \new_[33635]_  = ~A265 & ~A236;
  assign \new_[33636]_  = ~A235 & \new_[33635]_ ;
  assign \new_[33639]_  = ~A268 & ~A266;
  assign \new_[33642]_  = A300 & A298;
  assign \new_[33643]_  = \new_[33642]_  & \new_[33639]_ ;
  assign \new_[33644]_  = \new_[33643]_  & \new_[33636]_ ;
  assign \new_[33648]_  = A200 & A199;
  assign \new_[33649]_  = A169 & \new_[33648]_ ;
  assign \new_[33653]_  = A232 & ~A202;
  assign \new_[33654]_  = ~A201 & \new_[33653]_ ;
  assign \new_[33655]_  = \new_[33654]_  & \new_[33649]_ ;
  assign \new_[33659]_  = ~A235 & ~A234;
  assign \new_[33660]_  = A233 & \new_[33659]_ ;
  assign \new_[33663]_  = ~A268 & ~A267;
  assign \new_[33666]_  = A301 & ~A269;
  assign \new_[33667]_  = \new_[33666]_  & \new_[33663]_ ;
  assign \new_[33668]_  = \new_[33667]_  & \new_[33660]_ ;
  assign \new_[33672]_  = A200 & A199;
  assign \new_[33673]_  = A169 & \new_[33672]_ ;
  assign \new_[33677]_  = A232 & ~A202;
  assign \new_[33678]_  = ~A201 & \new_[33677]_ ;
  assign \new_[33679]_  = \new_[33678]_  & \new_[33673]_ ;
  assign \new_[33683]_  = ~A235 & ~A234;
  assign \new_[33684]_  = A233 & \new_[33683]_ ;
  assign \new_[33687]_  = ~A266 & ~A265;
  assign \new_[33690]_  = A301 & ~A268;
  assign \new_[33691]_  = \new_[33690]_  & \new_[33687]_ ;
  assign \new_[33692]_  = \new_[33691]_  & \new_[33684]_ ;
  assign \new_[33696]_  = A200 & A199;
  assign \new_[33697]_  = A169 & \new_[33696]_ ;
  assign \new_[33701]_  = ~A232 & ~A202;
  assign \new_[33702]_  = ~A201 & \new_[33701]_ ;
  assign \new_[33703]_  = \new_[33702]_  & \new_[33697]_ ;
  assign \new_[33707]_  = ~A267 & ~A235;
  assign \new_[33708]_  = ~A233 & \new_[33707]_ ;
  assign \new_[33711]_  = ~A269 & ~A268;
  assign \new_[33714]_  = A300 & A299;
  assign \new_[33715]_  = \new_[33714]_  & \new_[33711]_ ;
  assign \new_[33716]_  = \new_[33715]_  & \new_[33708]_ ;
  assign \new_[33720]_  = A200 & A199;
  assign \new_[33721]_  = A169 & \new_[33720]_ ;
  assign \new_[33725]_  = ~A232 & ~A202;
  assign \new_[33726]_  = ~A201 & \new_[33725]_ ;
  assign \new_[33727]_  = \new_[33726]_  & \new_[33721]_ ;
  assign \new_[33731]_  = ~A267 & ~A235;
  assign \new_[33732]_  = ~A233 & \new_[33731]_ ;
  assign \new_[33735]_  = ~A269 & ~A268;
  assign \new_[33738]_  = A300 & A298;
  assign \new_[33739]_  = \new_[33738]_  & \new_[33735]_ ;
  assign \new_[33740]_  = \new_[33739]_  & \new_[33732]_ ;
  assign \new_[33744]_  = A200 & A199;
  assign \new_[33745]_  = A169 & \new_[33744]_ ;
  assign \new_[33749]_  = ~A232 & ~A202;
  assign \new_[33750]_  = ~A201 & \new_[33749]_ ;
  assign \new_[33751]_  = \new_[33750]_  & \new_[33745]_ ;
  assign \new_[33755]_  = A265 & ~A235;
  assign \new_[33756]_  = ~A233 & \new_[33755]_ ;
  assign \new_[33759]_  = ~A267 & A266;
  assign \new_[33762]_  = A301 & ~A268;
  assign \new_[33763]_  = \new_[33762]_  & \new_[33759]_ ;
  assign \new_[33764]_  = \new_[33763]_  & \new_[33756]_ ;
  assign \new_[33768]_  = A200 & A199;
  assign \new_[33769]_  = A169 & \new_[33768]_ ;
  assign \new_[33773]_  = ~A232 & ~A202;
  assign \new_[33774]_  = ~A201 & \new_[33773]_ ;
  assign \new_[33775]_  = \new_[33774]_  & \new_[33769]_ ;
  assign \new_[33779]_  = ~A265 & ~A235;
  assign \new_[33780]_  = ~A233 & \new_[33779]_ ;
  assign \new_[33783]_  = ~A268 & ~A266;
  assign \new_[33786]_  = A300 & A299;
  assign \new_[33787]_  = \new_[33786]_  & \new_[33783]_ ;
  assign \new_[33788]_  = \new_[33787]_  & \new_[33780]_ ;
  assign \new_[33792]_  = A200 & A199;
  assign \new_[33793]_  = A169 & \new_[33792]_ ;
  assign \new_[33797]_  = ~A232 & ~A202;
  assign \new_[33798]_  = ~A201 & \new_[33797]_ ;
  assign \new_[33799]_  = \new_[33798]_  & \new_[33793]_ ;
  assign \new_[33803]_  = ~A265 & ~A235;
  assign \new_[33804]_  = ~A233 & \new_[33803]_ ;
  assign \new_[33807]_  = ~A268 & ~A266;
  assign \new_[33810]_  = A300 & A298;
  assign \new_[33811]_  = \new_[33810]_  & \new_[33807]_ ;
  assign \new_[33812]_  = \new_[33811]_  & \new_[33804]_ ;
  assign \new_[33816]_  = ~A200 & ~A199;
  assign \new_[33817]_  = A169 & \new_[33816]_ ;
  assign \new_[33821]_  = ~A235 & ~A234;
  assign \new_[33822]_  = ~A202 & \new_[33821]_ ;
  assign \new_[33823]_  = \new_[33822]_  & \new_[33817]_ ;
  assign \new_[33827]_  = ~A268 & ~A267;
  assign \new_[33828]_  = ~A236 & \new_[33827]_ ;
  assign \new_[33831]_  = A298 & ~A269;
  assign \new_[33834]_  = A302 & ~A299;
  assign \new_[33835]_  = \new_[33834]_  & \new_[33831]_ ;
  assign \new_[33836]_  = \new_[33835]_  & \new_[33828]_ ;
  assign \new_[33840]_  = ~A200 & ~A199;
  assign \new_[33841]_  = A169 & \new_[33840]_ ;
  assign \new_[33845]_  = ~A235 & ~A234;
  assign \new_[33846]_  = ~A202 & \new_[33845]_ ;
  assign \new_[33847]_  = \new_[33846]_  & \new_[33841]_ ;
  assign \new_[33851]_  = ~A268 & ~A267;
  assign \new_[33852]_  = ~A236 & \new_[33851]_ ;
  assign \new_[33855]_  = ~A298 & ~A269;
  assign \new_[33858]_  = A302 & A299;
  assign \new_[33859]_  = \new_[33858]_  & \new_[33855]_ ;
  assign \new_[33860]_  = \new_[33859]_  & \new_[33852]_ ;
  assign \new_[33864]_  = ~A200 & ~A199;
  assign \new_[33865]_  = A169 & \new_[33864]_ ;
  assign \new_[33869]_  = ~A235 & ~A234;
  assign \new_[33870]_  = ~A202 & \new_[33869]_ ;
  assign \new_[33871]_  = \new_[33870]_  & \new_[33865]_ ;
  assign \new_[33875]_  = A266 & A265;
  assign \new_[33876]_  = ~A236 & \new_[33875]_ ;
  assign \new_[33879]_  = ~A268 & ~A267;
  assign \new_[33882]_  = A300 & A299;
  assign \new_[33883]_  = \new_[33882]_  & \new_[33879]_ ;
  assign \new_[33884]_  = \new_[33883]_  & \new_[33876]_ ;
  assign \new_[33888]_  = ~A200 & ~A199;
  assign \new_[33889]_  = A169 & \new_[33888]_ ;
  assign \new_[33893]_  = ~A235 & ~A234;
  assign \new_[33894]_  = ~A202 & \new_[33893]_ ;
  assign \new_[33895]_  = \new_[33894]_  & \new_[33889]_ ;
  assign \new_[33899]_  = A266 & A265;
  assign \new_[33900]_  = ~A236 & \new_[33899]_ ;
  assign \new_[33903]_  = ~A268 & ~A267;
  assign \new_[33906]_  = A300 & A298;
  assign \new_[33907]_  = \new_[33906]_  & \new_[33903]_ ;
  assign \new_[33908]_  = \new_[33907]_  & \new_[33900]_ ;
  assign \new_[33912]_  = ~A200 & ~A199;
  assign \new_[33913]_  = A169 & \new_[33912]_ ;
  assign \new_[33917]_  = ~A235 & ~A234;
  assign \new_[33918]_  = ~A202 & \new_[33917]_ ;
  assign \new_[33919]_  = \new_[33918]_  & \new_[33913]_ ;
  assign \new_[33923]_  = ~A266 & ~A265;
  assign \new_[33924]_  = ~A236 & \new_[33923]_ ;
  assign \new_[33927]_  = A298 & ~A268;
  assign \new_[33930]_  = A302 & ~A299;
  assign \new_[33931]_  = \new_[33930]_  & \new_[33927]_ ;
  assign \new_[33932]_  = \new_[33931]_  & \new_[33924]_ ;
  assign \new_[33936]_  = ~A200 & ~A199;
  assign \new_[33937]_  = A169 & \new_[33936]_ ;
  assign \new_[33941]_  = ~A235 & ~A234;
  assign \new_[33942]_  = ~A202 & \new_[33941]_ ;
  assign \new_[33943]_  = \new_[33942]_  & \new_[33937]_ ;
  assign \new_[33947]_  = ~A266 & ~A265;
  assign \new_[33948]_  = ~A236 & \new_[33947]_ ;
  assign \new_[33951]_  = ~A298 & ~A268;
  assign \new_[33954]_  = A302 & A299;
  assign \new_[33955]_  = \new_[33954]_  & \new_[33951]_ ;
  assign \new_[33956]_  = \new_[33955]_  & \new_[33948]_ ;
  assign \new_[33960]_  = ~A200 & ~A199;
  assign \new_[33961]_  = A169 & \new_[33960]_ ;
  assign \new_[33965]_  = A233 & A232;
  assign \new_[33966]_  = ~A202 & \new_[33965]_ ;
  assign \new_[33967]_  = \new_[33966]_  & \new_[33961]_ ;
  assign \new_[33971]_  = ~A267 & ~A235;
  assign \new_[33972]_  = ~A234 & \new_[33971]_ ;
  assign \new_[33975]_  = ~A269 & ~A268;
  assign \new_[33978]_  = A300 & A299;
  assign \new_[33979]_  = \new_[33978]_  & \new_[33975]_ ;
  assign \new_[33980]_  = \new_[33979]_  & \new_[33972]_ ;
  assign \new_[33984]_  = ~A200 & ~A199;
  assign \new_[33985]_  = A169 & \new_[33984]_ ;
  assign \new_[33989]_  = A233 & A232;
  assign \new_[33990]_  = ~A202 & \new_[33989]_ ;
  assign \new_[33991]_  = \new_[33990]_  & \new_[33985]_ ;
  assign \new_[33995]_  = ~A267 & ~A235;
  assign \new_[33996]_  = ~A234 & \new_[33995]_ ;
  assign \new_[33999]_  = ~A269 & ~A268;
  assign \new_[34002]_  = A300 & A298;
  assign \new_[34003]_  = \new_[34002]_  & \new_[33999]_ ;
  assign \new_[34004]_  = \new_[34003]_  & \new_[33996]_ ;
  assign \new_[34008]_  = ~A200 & ~A199;
  assign \new_[34009]_  = A169 & \new_[34008]_ ;
  assign \new_[34013]_  = A233 & A232;
  assign \new_[34014]_  = ~A202 & \new_[34013]_ ;
  assign \new_[34015]_  = \new_[34014]_  & \new_[34009]_ ;
  assign \new_[34019]_  = A265 & ~A235;
  assign \new_[34020]_  = ~A234 & \new_[34019]_ ;
  assign \new_[34023]_  = ~A267 & A266;
  assign \new_[34026]_  = A301 & ~A268;
  assign \new_[34027]_  = \new_[34026]_  & \new_[34023]_ ;
  assign \new_[34028]_  = \new_[34027]_  & \new_[34020]_ ;
  assign \new_[34032]_  = ~A200 & ~A199;
  assign \new_[34033]_  = A169 & \new_[34032]_ ;
  assign \new_[34037]_  = A233 & A232;
  assign \new_[34038]_  = ~A202 & \new_[34037]_ ;
  assign \new_[34039]_  = \new_[34038]_  & \new_[34033]_ ;
  assign \new_[34043]_  = ~A265 & ~A235;
  assign \new_[34044]_  = ~A234 & \new_[34043]_ ;
  assign \new_[34047]_  = ~A268 & ~A266;
  assign \new_[34050]_  = A300 & A299;
  assign \new_[34051]_  = \new_[34050]_  & \new_[34047]_ ;
  assign \new_[34052]_  = \new_[34051]_  & \new_[34044]_ ;
  assign \new_[34056]_  = ~A200 & ~A199;
  assign \new_[34057]_  = A169 & \new_[34056]_ ;
  assign \new_[34061]_  = A233 & A232;
  assign \new_[34062]_  = ~A202 & \new_[34061]_ ;
  assign \new_[34063]_  = \new_[34062]_  & \new_[34057]_ ;
  assign \new_[34067]_  = ~A265 & ~A235;
  assign \new_[34068]_  = ~A234 & \new_[34067]_ ;
  assign \new_[34071]_  = ~A268 & ~A266;
  assign \new_[34074]_  = A300 & A298;
  assign \new_[34075]_  = \new_[34074]_  & \new_[34071]_ ;
  assign \new_[34076]_  = \new_[34075]_  & \new_[34068]_ ;
  assign \new_[34080]_  = ~A200 & ~A199;
  assign \new_[34081]_  = A169 & \new_[34080]_ ;
  assign \new_[34085]_  = ~A233 & ~A232;
  assign \new_[34086]_  = ~A202 & \new_[34085]_ ;
  assign \new_[34087]_  = \new_[34086]_  & \new_[34081]_ ;
  assign \new_[34091]_  = ~A268 & ~A267;
  assign \new_[34092]_  = ~A235 & \new_[34091]_ ;
  assign \new_[34095]_  = A298 & ~A269;
  assign \new_[34098]_  = A302 & ~A299;
  assign \new_[34099]_  = \new_[34098]_  & \new_[34095]_ ;
  assign \new_[34100]_  = \new_[34099]_  & \new_[34092]_ ;
  assign \new_[34104]_  = ~A200 & ~A199;
  assign \new_[34105]_  = A169 & \new_[34104]_ ;
  assign \new_[34109]_  = ~A233 & ~A232;
  assign \new_[34110]_  = ~A202 & \new_[34109]_ ;
  assign \new_[34111]_  = \new_[34110]_  & \new_[34105]_ ;
  assign \new_[34115]_  = ~A268 & ~A267;
  assign \new_[34116]_  = ~A235 & \new_[34115]_ ;
  assign \new_[34119]_  = ~A298 & ~A269;
  assign \new_[34122]_  = A302 & A299;
  assign \new_[34123]_  = \new_[34122]_  & \new_[34119]_ ;
  assign \new_[34124]_  = \new_[34123]_  & \new_[34116]_ ;
  assign \new_[34128]_  = ~A200 & ~A199;
  assign \new_[34129]_  = A169 & \new_[34128]_ ;
  assign \new_[34133]_  = ~A233 & ~A232;
  assign \new_[34134]_  = ~A202 & \new_[34133]_ ;
  assign \new_[34135]_  = \new_[34134]_  & \new_[34129]_ ;
  assign \new_[34139]_  = A266 & A265;
  assign \new_[34140]_  = ~A235 & \new_[34139]_ ;
  assign \new_[34143]_  = ~A268 & ~A267;
  assign \new_[34146]_  = A300 & A299;
  assign \new_[34147]_  = \new_[34146]_  & \new_[34143]_ ;
  assign \new_[34148]_  = \new_[34147]_  & \new_[34140]_ ;
  assign \new_[34152]_  = ~A200 & ~A199;
  assign \new_[34153]_  = A169 & \new_[34152]_ ;
  assign \new_[34157]_  = ~A233 & ~A232;
  assign \new_[34158]_  = ~A202 & \new_[34157]_ ;
  assign \new_[34159]_  = \new_[34158]_  & \new_[34153]_ ;
  assign \new_[34163]_  = A266 & A265;
  assign \new_[34164]_  = ~A235 & \new_[34163]_ ;
  assign \new_[34167]_  = ~A268 & ~A267;
  assign \new_[34170]_  = A300 & A298;
  assign \new_[34171]_  = \new_[34170]_  & \new_[34167]_ ;
  assign \new_[34172]_  = \new_[34171]_  & \new_[34164]_ ;
  assign \new_[34176]_  = ~A200 & ~A199;
  assign \new_[34177]_  = A169 & \new_[34176]_ ;
  assign \new_[34181]_  = ~A233 & ~A232;
  assign \new_[34182]_  = ~A202 & \new_[34181]_ ;
  assign \new_[34183]_  = \new_[34182]_  & \new_[34177]_ ;
  assign \new_[34187]_  = ~A266 & ~A265;
  assign \new_[34188]_  = ~A235 & \new_[34187]_ ;
  assign \new_[34191]_  = A298 & ~A268;
  assign \new_[34194]_  = A302 & ~A299;
  assign \new_[34195]_  = \new_[34194]_  & \new_[34191]_ ;
  assign \new_[34196]_  = \new_[34195]_  & \new_[34188]_ ;
  assign \new_[34200]_  = ~A200 & ~A199;
  assign \new_[34201]_  = A169 & \new_[34200]_ ;
  assign \new_[34205]_  = ~A233 & ~A232;
  assign \new_[34206]_  = ~A202 & \new_[34205]_ ;
  assign \new_[34207]_  = \new_[34206]_  & \new_[34201]_ ;
  assign \new_[34211]_  = ~A266 & ~A265;
  assign \new_[34212]_  = ~A235 & \new_[34211]_ ;
  assign \new_[34215]_  = ~A298 & ~A268;
  assign \new_[34218]_  = A302 & A299;
  assign \new_[34219]_  = \new_[34218]_  & \new_[34215]_ ;
  assign \new_[34220]_  = \new_[34219]_  & \new_[34212]_ ;
  assign \new_[34224]_  = ~A166 & ~A167;
  assign \new_[34225]_  = ~A169 & \new_[34224]_ ;
  assign \new_[34229]_  = ~A235 & ~A234;
  assign \new_[34230]_  = A202 & \new_[34229]_ ;
  assign \new_[34231]_  = \new_[34230]_  & \new_[34225]_ ;
  assign \new_[34235]_  = ~A268 & ~A267;
  assign \new_[34236]_  = ~A236 & \new_[34235]_ ;
  assign \new_[34239]_  = A298 & ~A269;
  assign \new_[34242]_  = A302 & ~A299;
  assign \new_[34243]_  = \new_[34242]_  & \new_[34239]_ ;
  assign \new_[34244]_  = \new_[34243]_  & \new_[34236]_ ;
  assign \new_[34248]_  = ~A166 & ~A167;
  assign \new_[34249]_  = ~A169 & \new_[34248]_ ;
  assign \new_[34253]_  = ~A235 & ~A234;
  assign \new_[34254]_  = A202 & \new_[34253]_ ;
  assign \new_[34255]_  = \new_[34254]_  & \new_[34249]_ ;
  assign \new_[34259]_  = ~A268 & ~A267;
  assign \new_[34260]_  = ~A236 & \new_[34259]_ ;
  assign \new_[34263]_  = ~A298 & ~A269;
  assign \new_[34266]_  = A302 & A299;
  assign \new_[34267]_  = \new_[34266]_  & \new_[34263]_ ;
  assign \new_[34268]_  = \new_[34267]_  & \new_[34260]_ ;
  assign \new_[34272]_  = ~A166 & ~A167;
  assign \new_[34273]_  = ~A169 & \new_[34272]_ ;
  assign \new_[34277]_  = ~A235 & ~A234;
  assign \new_[34278]_  = A202 & \new_[34277]_ ;
  assign \new_[34279]_  = \new_[34278]_  & \new_[34273]_ ;
  assign \new_[34283]_  = A266 & A265;
  assign \new_[34284]_  = ~A236 & \new_[34283]_ ;
  assign \new_[34287]_  = ~A268 & ~A267;
  assign \new_[34290]_  = A300 & A299;
  assign \new_[34291]_  = \new_[34290]_  & \new_[34287]_ ;
  assign \new_[34292]_  = \new_[34291]_  & \new_[34284]_ ;
  assign \new_[34296]_  = ~A166 & ~A167;
  assign \new_[34297]_  = ~A169 & \new_[34296]_ ;
  assign \new_[34301]_  = ~A235 & ~A234;
  assign \new_[34302]_  = A202 & \new_[34301]_ ;
  assign \new_[34303]_  = \new_[34302]_  & \new_[34297]_ ;
  assign \new_[34307]_  = A266 & A265;
  assign \new_[34308]_  = ~A236 & \new_[34307]_ ;
  assign \new_[34311]_  = ~A268 & ~A267;
  assign \new_[34314]_  = A300 & A298;
  assign \new_[34315]_  = \new_[34314]_  & \new_[34311]_ ;
  assign \new_[34316]_  = \new_[34315]_  & \new_[34308]_ ;
  assign \new_[34320]_  = ~A166 & ~A167;
  assign \new_[34321]_  = ~A169 & \new_[34320]_ ;
  assign \new_[34325]_  = ~A235 & ~A234;
  assign \new_[34326]_  = A202 & \new_[34325]_ ;
  assign \new_[34327]_  = \new_[34326]_  & \new_[34321]_ ;
  assign \new_[34331]_  = ~A266 & ~A265;
  assign \new_[34332]_  = ~A236 & \new_[34331]_ ;
  assign \new_[34335]_  = A298 & ~A268;
  assign \new_[34338]_  = A302 & ~A299;
  assign \new_[34339]_  = \new_[34338]_  & \new_[34335]_ ;
  assign \new_[34340]_  = \new_[34339]_  & \new_[34332]_ ;
  assign \new_[34344]_  = ~A166 & ~A167;
  assign \new_[34345]_  = ~A169 & \new_[34344]_ ;
  assign \new_[34349]_  = ~A235 & ~A234;
  assign \new_[34350]_  = A202 & \new_[34349]_ ;
  assign \new_[34351]_  = \new_[34350]_  & \new_[34345]_ ;
  assign \new_[34355]_  = ~A266 & ~A265;
  assign \new_[34356]_  = ~A236 & \new_[34355]_ ;
  assign \new_[34359]_  = ~A298 & ~A268;
  assign \new_[34362]_  = A302 & A299;
  assign \new_[34363]_  = \new_[34362]_  & \new_[34359]_ ;
  assign \new_[34364]_  = \new_[34363]_  & \new_[34356]_ ;
  assign \new_[34368]_  = ~A166 & ~A167;
  assign \new_[34369]_  = ~A169 & \new_[34368]_ ;
  assign \new_[34373]_  = A233 & A232;
  assign \new_[34374]_  = A202 & \new_[34373]_ ;
  assign \new_[34375]_  = \new_[34374]_  & \new_[34369]_ ;
  assign \new_[34379]_  = ~A267 & ~A235;
  assign \new_[34380]_  = ~A234 & \new_[34379]_ ;
  assign \new_[34383]_  = ~A269 & ~A268;
  assign \new_[34386]_  = A300 & A299;
  assign \new_[34387]_  = \new_[34386]_  & \new_[34383]_ ;
  assign \new_[34388]_  = \new_[34387]_  & \new_[34380]_ ;
  assign \new_[34392]_  = ~A166 & ~A167;
  assign \new_[34393]_  = ~A169 & \new_[34392]_ ;
  assign \new_[34397]_  = A233 & A232;
  assign \new_[34398]_  = A202 & \new_[34397]_ ;
  assign \new_[34399]_  = \new_[34398]_  & \new_[34393]_ ;
  assign \new_[34403]_  = ~A267 & ~A235;
  assign \new_[34404]_  = ~A234 & \new_[34403]_ ;
  assign \new_[34407]_  = ~A269 & ~A268;
  assign \new_[34410]_  = A300 & A298;
  assign \new_[34411]_  = \new_[34410]_  & \new_[34407]_ ;
  assign \new_[34412]_  = \new_[34411]_  & \new_[34404]_ ;
  assign \new_[34416]_  = ~A166 & ~A167;
  assign \new_[34417]_  = ~A169 & \new_[34416]_ ;
  assign \new_[34421]_  = A233 & A232;
  assign \new_[34422]_  = A202 & \new_[34421]_ ;
  assign \new_[34423]_  = \new_[34422]_  & \new_[34417]_ ;
  assign \new_[34427]_  = A265 & ~A235;
  assign \new_[34428]_  = ~A234 & \new_[34427]_ ;
  assign \new_[34431]_  = ~A267 & A266;
  assign \new_[34434]_  = A301 & ~A268;
  assign \new_[34435]_  = \new_[34434]_  & \new_[34431]_ ;
  assign \new_[34436]_  = \new_[34435]_  & \new_[34428]_ ;
  assign \new_[34440]_  = ~A166 & ~A167;
  assign \new_[34441]_  = ~A169 & \new_[34440]_ ;
  assign \new_[34445]_  = A233 & A232;
  assign \new_[34446]_  = A202 & \new_[34445]_ ;
  assign \new_[34447]_  = \new_[34446]_  & \new_[34441]_ ;
  assign \new_[34451]_  = ~A265 & ~A235;
  assign \new_[34452]_  = ~A234 & \new_[34451]_ ;
  assign \new_[34455]_  = ~A268 & ~A266;
  assign \new_[34458]_  = A300 & A299;
  assign \new_[34459]_  = \new_[34458]_  & \new_[34455]_ ;
  assign \new_[34460]_  = \new_[34459]_  & \new_[34452]_ ;
  assign \new_[34464]_  = ~A166 & ~A167;
  assign \new_[34465]_  = ~A169 & \new_[34464]_ ;
  assign \new_[34469]_  = A233 & A232;
  assign \new_[34470]_  = A202 & \new_[34469]_ ;
  assign \new_[34471]_  = \new_[34470]_  & \new_[34465]_ ;
  assign \new_[34475]_  = ~A265 & ~A235;
  assign \new_[34476]_  = ~A234 & \new_[34475]_ ;
  assign \new_[34479]_  = ~A268 & ~A266;
  assign \new_[34482]_  = A300 & A298;
  assign \new_[34483]_  = \new_[34482]_  & \new_[34479]_ ;
  assign \new_[34484]_  = \new_[34483]_  & \new_[34476]_ ;
  assign \new_[34488]_  = ~A166 & ~A167;
  assign \new_[34489]_  = ~A169 & \new_[34488]_ ;
  assign \new_[34493]_  = ~A233 & ~A232;
  assign \new_[34494]_  = A202 & \new_[34493]_ ;
  assign \new_[34495]_  = \new_[34494]_  & \new_[34489]_ ;
  assign \new_[34499]_  = ~A268 & ~A267;
  assign \new_[34500]_  = ~A235 & \new_[34499]_ ;
  assign \new_[34503]_  = A298 & ~A269;
  assign \new_[34506]_  = A302 & ~A299;
  assign \new_[34507]_  = \new_[34506]_  & \new_[34503]_ ;
  assign \new_[34508]_  = \new_[34507]_  & \new_[34500]_ ;
  assign \new_[34512]_  = ~A166 & ~A167;
  assign \new_[34513]_  = ~A169 & \new_[34512]_ ;
  assign \new_[34517]_  = ~A233 & ~A232;
  assign \new_[34518]_  = A202 & \new_[34517]_ ;
  assign \new_[34519]_  = \new_[34518]_  & \new_[34513]_ ;
  assign \new_[34523]_  = ~A268 & ~A267;
  assign \new_[34524]_  = ~A235 & \new_[34523]_ ;
  assign \new_[34527]_  = ~A298 & ~A269;
  assign \new_[34530]_  = A302 & A299;
  assign \new_[34531]_  = \new_[34530]_  & \new_[34527]_ ;
  assign \new_[34532]_  = \new_[34531]_  & \new_[34524]_ ;
  assign \new_[34536]_  = ~A166 & ~A167;
  assign \new_[34537]_  = ~A169 & \new_[34536]_ ;
  assign \new_[34541]_  = ~A233 & ~A232;
  assign \new_[34542]_  = A202 & \new_[34541]_ ;
  assign \new_[34543]_  = \new_[34542]_  & \new_[34537]_ ;
  assign \new_[34547]_  = A266 & A265;
  assign \new_[34548]_  = ~A235 & \new_[34547]_ ;
  assign \new_[34551]_  = ~A268 & ~A267;
  assign \new_[34554]_  = A300 & A299;
  assign \new_[34555]_  = \new_[34554]_  & \new_[34551]_ ;
  assign \new_[34556]_  = \new_[34555]_  & \new_[34548]_ ;
  assign \new_[34560]_  = ~A166 & ~A167;
  assign \new_[34561]_  = ~A169 & \new_[34560]_ ;
  assign \new_[34565]_  = ~A233 & ~A232;
  assign \new_[34566]_  = A202 & \new_[34565]_ ;
  assign \new_[34567]_  = \new_[34566]_  & \new_[34561]_ ;
  assign \new_[34571]_  = A266 & A265;
  assign \new_[34572]_  = ~A235 & \new_[34571]_ ;
  assign \new_[34575]_  = ~A268 & ~A267;
  assign \new_[34578]_  = A300 & A298;
  assign \new_[34579]_  = \new_[34578]_  & \new_[34575]_ ;
  assign \new_[34580]_  = \new_[34579]_  & \new_[34572]_ ;
  assign \new_[34584]_  = ~A166 & ~A167;
  assign \new_[34585]_  = ~A169 & \new_[34584]_ ;
  assign \new_[34589]_  = ~A233 & ~A232;
  assign \new_[34590]_  = A202 & \new_[34589]_ ;
  assign \new_[34591]_  = \new_[34590]_  & \new_[34585]_ ;
  assign \new_[34595]_  = ~A266 & ~A265;
  assign \new_[34596]_  = ~A235 & \new_[34595]_ ;
  assign \new_[34599]_  = A298 & ~A268;
  assign \new_[34602]_  = A302 & ~A299;
  assign \new_[34603]_  = \new_[34602]_  & \new_[34599]_ ;
  assign \new_[34604]_  = \new_[34603]_  & \new_[34596]_ ;
  assign \new_[34608]_  = ~A166 & ~A167;
  assign \new_[34609]_  = ~A169 & \new_[34608]_ ;
  assign \new_[34613]_  = ~A233 & ~A232;
  assign \new_[34614]_  = A202 & \new_[34613]_ ;
  assign \new_[34615]_  = \new_[34614]_  & \new_[34609]_ ;
  assign \new_[34619]_  = ~A266 & ~A265;
  assign \new_[34620]_  = ~A235 & \new_[34619]_ ;
  assign \new_[34623]_  = ~A298 & ~A268;
  assign \new_[34626]_  = A302 & A299;
  assign \new_[34627]_  = \new_[34626]_  & \new_[34623]_ ;
  assign \new_[34628]_  = \new_[34627]_  & \new_[34620]_ ;
  assign \new_[34632]_  = ~A166 & ~A167;
  assign \new_[34633]_  = ~A169 & \new_[34632]_ ;
  assign \new_[34637]_  = ~A234 & A201;
  assign \new_[34638]_  = A199 & \new_[34637]_ ;
  assign \new_[34639]_  = \new_[34638]_  & \new_[34633]_ ;
  assign \new_[34643]_  = ~A267 & ~A236;
  assign \new_[34644]_  = ~A235 & \new_[34643]_ ;
  assign \new_[34647]_  = ~A269 & ~A268;
  assign \new_[34650]_  = A300 & A299;
  assign \new_[34651]_  = \new_[34650]_  & \new_[34647]_ ;
  assign \new_[34652]_  = \new_[34651]_  & \new_[34644]_ ;
  assign \new_[34656]_  = ~A166 & ~A167;
  assign \new_[34657]_  = ~A169 & \new_[34656]_ ;
  assign \new_[34661]_  = ~A234 & A201;
  assign \new_[34662]_  = A199 & \new_[34661]_ ;
  assign \new_[34663]_  = \new_[34662]_  & \new_[34657]_ ;
  assign \new_[34667]_  = ~A267 & ~A236;
  assign \new_[34668]_  = ~A235 & \new_[34667]_ ;
  assign \new_[34671]_  = ~A269 & ~A268;
  assign \new_[34674]_  = A300 & A298;
  assign \new_[34675]_  = \new_[34674]_  & \new_[34671]_ ;
  assign \new_[34676]_  = \new_[34675]_  & \new_[34668]_ ;
  assign \new_[34680]_  = ~A166 & ~A167;
  assign \new_[34681]_  = ~A169 & \new_[34680]_ ;
  assign \new_[34685]_  = ~A234 & A201;
  assign \new_[34686]_  = A199 & \new_[34685]_ ;
  assign \new_[34687]_  = \new_[34686]_  & \new_[34681]_ ;
  assign \new_[34691]_  = A265 & ~A236;
  assign \new_[34692]_  = ~A235 & \new_[34691]_ ;
  assign \new_[34695]_  = ~A267 & A266;
  assign \new_[34698]_  = A301 & ~A268;
  assign \new_[34699]_  = \new_[34698]_  & \new_[34695]_ ;
  assign \new_[34700]_  = \new_[34699]_  & \new_[34692]_ ;
  assign \new_[34704]_  = ~A166 & ~A167;
  assign \new_[34705]_  = ~A169 & \new_[34704]_ ;
  assign \new_[34709]_  = ~A234 & A201;
  assign \new_[34710]_  = A199 & \new_[34709]_ ;
  assign \new_[34711]_  = \new_[34710]_  & \new_[34705]_ ;
  assign \new_[34715]_  = ~A265 & ~A236;
  assign \new_[34716]_  = ~A235 & \new_[34715]_ ;
  assign \new_[34719]_  = ~A268 & ~A266;
  assign \new_[34722]_  = A300 & A299;
  assign \new_[34723]_  = \new_[34722]_  & \new_[34719]_ ;
  assign \new_[34724]_  = \new_[34723]_  & \new_[34716]_ ;
  assign \new_[34728]_  = ~A166 & ~A167;
  assign \new_[34729]_  = ~A169 & \new_[34728]_ ;
  assign \new_[34733]_  = ~A234 & A201;
  assign \new_[34734]_  = A199 & \new_[34733]_ ;
  assign \new_[34735]_  = \new_[34734]_  & \new_[34729]_ ;
  assign \new_[34739]_  = ~A265 & ~A236;
  assign \new_[34740]_  = ~A235 & \new_[34739]_ ;
  assign \new_[34743]_  = ~A268 & ~A266;
  assign \new_[34746]_  = A300 & A298;
  assign \new_[34747]_  = \new_[34746]_  & \new_[34743]_ ;
  assign \new_[34748]_  = \new_[34747]_  & \new_[34740]_ ;
  assign \new_[34752]_  = ~A166 & ~A167;
  assign \new_[34753]_  = ~A169 & \new_[34752]_ ;
  assign \new_[34757]_  = A232 & A201;
  assign \new_[34758]_  = A199 & \new_[34757]_ ;
  assign \new_[34759]_  = \new_[34758]_  & \new_[34753]_ ;
  assign \new_[34763]_  = ~A235 & ~A234;
  assign \new_[34764]_  = A233 & \new_[34763]_ ;
  assign \new_[34767]_  = ~A268 & ~A267;
  assign \new_[34770]_  = A301 & ~A269;
  assign \new_[34771]_  = \new_[34770]_  & \new_[34767]_ ;
  assign \new_[34772]_  = \new_[34771]_  & \new_[34764]_ ;
  assign \new_[34776]_  = ~A166 & ~A167;
  assign \new_[34777]_  = ~A169 & \new_[34776]_ ;
  assign \new_[34781]_  = A232 & A201;
  assign \new_[34782]_  = A199 & \new_[34781]_ ;
  assign \new_[34783]_  = \new_[34782]_  & \new_[34777]_ ;
  assign \new_[34787]_  = ~A235 & ~A234;
  assign \new_[34788]_  = A233 & \new_[34787]_ ;
  assign \new_[34791]_  = ~A266 & ~A265;
  assign \new_[34794]_  = A301 & ~A268;
  assign \new_[34795]_  = \new_[34794]_  & \new_[34791]_ ;
  assign \new_[34796]_  = \new_[34795]_  & \new_[34788]_ ;
  assign \new_[34800]_  = ~A166 & ~A167;
  assign \new_[34801]_  = ~A169 & \new_[34800]_ ;
  assign \new_[34805]_  = ~A232 & A201;
  assign \new_[34806]_  = A199 & \new_[34805]_ ;
  assign \new_[34807]_  = \new_[34806]_  & \new_[34801]_ ;
  assign \new_[34811]_  = ~A267 & ~A235;
  assign \new_[34812]_  = ~A233 & \new_[34811]_ ;
  assign \new_[34815]_  = ~A269 & ~A268;
  assign \new_[34818]_  = A300 & A299;
  assign \new_[34819]_  = \new_[34818]_  & \new_[34815]_ ;
  assign \new_[34820]_  = \new_[34819]_  & \new_[34812]_ ;
  assign \new_[34824]_  = ~A166 & ~A167;
  assign \new_[34825]_  = ~A169 & \new_[34824]_ ;
  assign \new_[34829]_  = ~A232 & A201;
  assign \new_[34830]_  = A199 & \new_[34829]_ ;
  assign \new_[34831]_  = \new_[34830]_  & \new_[34825]_ ;
  assign \new_[34835]_  = ~A267 & ~A235;
  assign \new_[34836]_  = ~A233 & \new_[34835]_ ;
  assign \new_[34839]_  = ~A269 & ~A268;
  assign \new_[34842]_  = A300 & A298;
  assign \new_[34843]_  = \new_[34842]_  & \new_[34839]_ ;
  assign \new_[34844]_  = \new_[34843]_  & \new_[34836]_ ;
  assign \new_[34848]_  = ~A166 & ~A167;
  assign \new_[34849]_  = ~A169 & \new_[34848]_ ;
  assign \new_[34853]_  = ~A232 & A201;
  assign \new_[34854]_  = A199 & \new_[34853]_ ;
  assign \new_[34855]_  = \new_[34854]_  & \new_[34849]_ ;
  assign \new_[34859]_  = A265 & ~A235;
  assign \new_[34860]_  = ~A233 & \new_[34859]_ ;
  assign \new_[34863]_  = ~A267 & A266;
  assign \new_[34866]_  = A301 & ~A268;
  assign \new_[34867]_  = \new_[34866]_  & \new_[34863]_ ;
  assign \new_[34868]_  = \new_[34867]_  & \new_[34860]_ ;
  assign \new_[34872]_  = ~A166 & ~A167;
  assign \new_[34873]_  = ~A169 & \new_[34872]_ ;
  assign \new_[34877]_  = ~A232 & A201;
  assign \new_[34878]_  = A199 & \new_[34877]_ ;
  assign \new_[34879]_  = \new_[34878]_  & \new_[34873]_ ;
  assign \new_[34883]_  = ~A265 & ~A235;
  assign \new_[34884]_  = ~A233 & \new_[34883]_ ;
  assign \new_[34887]_  = ~A268 & ~A266;
  assign \new_[34890]_  = A300 & A299;
  assign \new_[34891]_  = \new_[34890]_  & \new_[34887]_ ;
  assign \new_[34892]_  = \new_[34891]_  & \new_[34884]_ ;
  assign \new_[34896]_  = ~A166 & ~A167;
  assign \new_[34897]_  = ~A169 & \new_[34896]_ ;
  assign \new_[34901]_  = ~A232 & A201;
  assign \new_[34902]_  = A199 & \new_[34901]_ ;
  assign \new_[34903]_  = \new_[34902]_  & \new_[34897]_ ;
  assign \new_[34907]_  = ~A265 & ~A235;
  assign \new_[34908]_  = ~A233 & \new_[34907]_ ;
  assign \new_[34911]_  = ~A268 & ~A266;
  assign \new_[34914]_  = A300 & A298;
  assign \new_[34915]_  = \new_[34914]_  & \new_[34911]_ ;
  assign \new_[34916]_  = \new_[34915]_  & \new_[34908]_ ;
  assign \new_[34920]_  = ~A166 & ~A167;
  assign \new_[34921]_  = ~A169 & \new_[34920]_ ;
  assign \new_[34925]_  = ~A234 & A201;
  assign \new_[34926]_  = A200 & \new_[34925]_ ;
  assign \new_[34927]_  = \new_[34926]_  & \new_[34921]_ ;
  assign \new_[34931]_  = ~A267 & ~A236;
  assign \new_[34932]_  = ~A235 & \new_[34931]_ ;
  assign \new_[34935]_  = ~A269 & ~A268;
  assign \new_[34938]_  = A300 & A299;
  assign \new_[34939]_  = \new_[34938]_  & \new_[34935]_ ;
  assign \new_[34940]_  = \new_[34939]_  & \new_[34932]_ ;
  assign \new_[34944]_  = ~A166 & ~A167;
  assign \new_[34945]_  = ~A169 & \new_[34944]_ ;
  assign \new_[34949]_  = ~A234 & A201;
  assign \new_[34950]_  = A200 & \new_[34949]_ ;
  assign \new_[34951]_  = \new_[34950]_  & \new_[34945]_ ;
  assign \new_[34955]_  = ~A267 & ~A236;
  assign \new_[34956]_  = ~A235 & \new_[34955]_ ;
  assign \new_[34959]_  = ~A269 & ~A268;
  assign \new_[34962]_  = A300 & A298;
  assign \new_[34963]_  = \new_[34962]_  & \new_[34959]_ ;
  assign \new_[34964]_  = \new_[34963]_  & \new_[34956]_ ;
  assign \new_[34968]_  = ~A166 & ~A167;
  assign \new_[34969]_  = ~A169 & \new_[34968]_ ;
  assign \new_[34973]_  = ~A234 & A201;
  assign \new_[34974]_  = A200 & \new_[34973]_ ;
  assign \new_[34975]_  = \new_[34974]_  & \new_[34969]_ ;
  assign \new_[34979]_  = A265 & ~A236;
  assign \new_[34980]_  = ~A235 & \new_[34979]_ ;
  assign \new_[34983]_  = ~A267 & A266;
  assign \new_[34986]_  = A301 & ~A268;
  assign \new_[34987]_  = \new_[34986]_  & \new_[34983]_ ;
  assign \new_[34988]_  = \new_[34987]_  & \new_[34980]_ ;
  assign \new_[34992]_  = ~A166 & ~A167;
  assign \new_[34993]_  = ~A169 & \new_[34992]_ ;
  assign \new_[34997]_  = ~A234 & A201;
  assign \new_[34998]_  = A200 & \new_[34997]_ ;
  assign \new_[34999]_  = \new_[34998]_  & \new_[34993]_ ;
  assign \new_[35003]_  = ~A265 & ~A236;
  assign \new_[35004]_  = ~A235 & \new_[35003]_ ;
  assign \new_[35007]_  = ~A268 & ~A266;
  assign \new_[35010]_  = A300 & A299;
  assign \new_[35011]_  = \new_[35010]_  & \new_[35007]_ ;
  assign \new_[35012]_  = \new_[35011]_  & \new_[35004]_ ;
  assign \new_[35016]_  = ~A166 & ~A167;
  assign \new_[35017]_  = ~A169 & \new_[35016]_ ;
  assign \new_[35021]_  = ~A234 & A201;
  assign \new_[35022]_  = A200 & \new_[35021]_ ;
  assign \new_[35023]_  = \new_[35022]_  & \new_[35017]_ ;
  assign \new_[35027]_  = ~A265 & ~A236;
  assign \new_[35028]_  = ~A235 & \new_[35027]_ ;
  assign \new_[35031]_  = ~A268 & ~A266;
  assign \new_[35034]_  = A300 & A298;
  assign \new_[35035]_  = \new_[35034]_  & \new_[35031]_ ;
  assign \new_[35036]_  = \new_[35035]_  & \new_[35028]_ ;
  assign \new_[35040]_  = ~A166 & ~A167;
  assign \new_[35041]_  = ~A169 & \new_[35040]_ ;
  assign \new_[35045]_  = A232 & A201;
  assign \new_[35046]_  = A200 & \new_[35045]_ ;
  assign \new_[35047]_  = \new_[35046]_  & \new_[35041]_ ;
  assign \new_[35051]_  = ~A235 & ~A234;
  assign \new_[35052]_  = A233 & \new_[35051]_ ;
  assign \new_[35055]_  = ~A268 & ~A267;
  assign \new_[35058]_  = A301 & ~A269;
  assign \new_[35059]_  = \new_[35058]_  & \new_[35055]_ ;
  assign \new_[35060]_  = \new_[35059]_  & \new_[35052]_ ;
  assign \new_[35064]_  = ~A166 & ~A167;
  assign \new_[35065]_  = ~A169 & \new_[35064]_ ;
  assign \new_[35069]_  = A232 & A201;
  assign \new_[35070]_  = A200 & \new_[35069]_ ;
  assign \new_[35071]_  = \new_[35070]_  & \new_[35065]_ ;
  assign \new_[35075]_  = ~A235 & ~A234;
  assign \new_[35076]_  = A233 & \new_[35075]_ ;
  assign \new_[35079]_  = ~A266 & ~A265;
  assign \new_[35082]_  = A301 & ~A268;
  assign \new_[35083]_  = \new_[35082]_  & \new_[35079]_ ;
  assign \new_[35084]_  = \new_[35083]_  & \new_[35076]_ ;
  assign \new_[35088]_  = ~A166 & ~A167;
  assign \new_[35089]_  = ~A169 & \new_[35088]_ ;
  assign \new_[35093]_  = ~A232 & A201;
  assign \new_[35094]_  = A200 & \new_[35093]_ ;
  assign \new_[35095]_  = \new_[35094]_  & \new_[35089]_ ;
  assign \new_[35099]_  = ~A267 & ~A235;
  assign \new_[35100]_  = ~A233 & \new_[35099]_ ;
  assign \new_[35103]_  = ~A269 & ~A268;
  assign \new_[35106]_  = A300 & A299;
  assign \new_[35107]_  = \new_[35106]_  & \new_[35103]_ ;
  assign \new_[35108]_  = \new_[35107]_  & \new_[35100]_ ;
  assign \new_[35112]_  = ~A166 & ~A167;
  assign \new_[35113]_  = ~A169 & \new_[35112]_ ;
  assign \new_[35117]_  = ~A232 & A201;
  assign \new_[35118]_  = A200 & \new_[35117]_ ;
  assign \new_[35119]_  = \new_[35118]_  & \new_[35113]_ ;
  assign \new_[35123]_  = ~A267 & ~A235;
  assign \new_[35124]_  = ~A233 & \new_[35123]_ ;
  assign \new_[35127]_  = ~A269 & ~A268;
  assign \new_[35130]_  = A300 & A298;
  assign \new_[35131]_  = \new_[35130]_  & \new_[35127]_ ;
  assign \new_[35132]_  = \new_[35131]_  & \new_[35124]_ ;
  assign \new_[35136]_  = ~A166 & ~A167;
  assign \new_[35137]_  = ~A169 & \new_[35136]_ ;
  assign \new_[35141]_  = ~A232 & A201;
  assign \new_[35142]_  = A200 & \new_[35141]_ ;
  assign \new_[35143]_  = \new_[35142]_  & \new_[35137]_ ;
  assign \new_[35147]_  = A265 & ~A235;
  assign \new_[35148]_  = ~A233 & \new_[35147]_ ;
  assign \new_[35151]_  = ~A267 & A266;
  assign \new_[35154]_  = A301 & ~A268;
  assign \new_[35155]_  = \new_[35154]_  & \new_[35151]_ ;
  assign \new_[35156]_  = \new_[35155]_  & \new_[35148]_ ;
  assign \new_[35160]_  = ~A166 & ~A167;
  assign \new_[35161]_  = ~A169 & \new_[35160]_ ;
  assign \new_[35165]_  = ~A232 & A201;
  assign \new_[35166]_  = A200 & \new_[35165]_ ;
  assign \new_[35167]_  = \new_[35166]_  & \new_[35161]_ ;
  assign \new_[35171]_  = ~A265 & ~A235;
  assign \new_[35172]_  = ~A233 & \new_[35171]_ ;
  assign \new_[35175]_  = ~A268 & ~A266;
  assign \new_[35178]_  = A300 & A299;
  assign \new_[35179]_  = \new_[35178]_  & \new_[35175]_ ;
  assign \new_[35180]_  = \new_[35179]_  & \new_[35172]_ ;
  assign \new_[35184]_  = ~A166 & ~A167;
  assign \new_[35185]_  = ~A169 & \new_[35184]_ ;
  assign \new_[35189]_  = ~A232 & A201;
  assign \new_[35190]_  = A200 & \new_[35189]_ ;
  assign \new_[35191]_  = \new_[35190]_  & \new_[35185]_ ;
  assign \new_[35195]_  = ~A265 & ~A235;
  assign \new_[35196]_  = ~A233 & \new_[35195]_ ;
  assign \new_[35199]_  = ~A268 & ~A266;
  assign \new_[35202]_  = A300 & A298;
  assign \new_[35203]_  = \new_[35202]_  & \new_[35199]_ ;
  assign \new_[35204]_  = \new_[35203]_  & \new_[35196]_ ;
  assign \new_[35208]_  = ~A166 & ~A167;
  assign \new_[35209]_  = ~A169 & \new_[35208]_ ;
  assign \new_[35213]_  = A203 & A200;
  assign \new_[35214]_  = ~A199 & \new_[35213]_ ;
  assign \new_[35215]_  = \new_[35214]_  & \new_[35209]_ ;
  assign \new_[35219]_  = ~A236 & ~A235;
  assign \new_[35220]_  = ~A234 & \new_[35219]_ ;
  assign \new_[35223]_  = ~A268 & ~A267;
  assign \new_[35226]_  = A301 & ~A269;
  assign \new_[35227]_  = \new_[35226]_  & \new_[35223]_ ;
  assign \new_[35228]_  = \new_[35227]_  & \new_[35220]_ ;
  assign \new_[35232]_  = ~A166 & ~A167;
  assign \new_[35233]_  = ~A169 & \new_[35232]_ ;
  assign \new_[35237]_  = A203 & A200;
  assign \new_[35238]_  = ~A199 & \new_[35237]_ ;
  assign \new_[35239]_  = \new_[35238]_  & \new_[35233]_ ;
  assign \new_[35243]_  = ~A236 & ~A235;
  assign \new_[35244]_  = ~A234 & \new_[35243]_ ;
  assign \new_[35247]_  = ~A266 & ~A265;
  assign \new_[35250]_  = A301 & ~A268;
  assign \new_[35251]_  = \new_[35250]_  & \new_[35247]_ ;
  assign \new_[35252]_  = \new_[35251]_  & \new_[35244]_ ;
  assign \new_[35256]_  = ~A166 & ~A167;
  assign \new_[35257]_  = ~A169 & \new_[35256]_ ;
  assign \new_[35261]_  = A203 & A200;
  assign \new_[35262]_  = ~A199 & \new_[35261]_ ;
  assign \new_[35263]_  = \new_[35262]_  & \new_[35257]_ ;
  assign \new_[35267]_  = A236 & A233;
  assign \new_[35268]_  = ~A232 & \new_[35267]_ ;
  assign \new_[35271]_  = A299 & A298;
  assign \new_[35274]_  = ~A301 & ~A300;
  assign \new_[35275]_  = \new_[35274]_  & \new_[35271]_ ;
  assign \new_[35276]_  = \new_[35275]_  & \new_[35268]_ ;
  assign \new_[35280]_  = ~A166 & ~A167;
  assign \new_[35281]_  = ~A169 & \new_[35280]_ ;
  assign \new_[35285]_  = A203 & A200;
  assign \new_[35286]_  = ~A199 & \new_[35285]_ ;
  assign \new_[35287]_  = \new_[35286]_  & \new_[35281]_ ;
  assign \new_[35291]_  = A236 & ~A233;
  assign \new_[35292]_  = A232 & \new_[35291]_ ;
  assign \new_[35295]_  = A299 & A298;
  assign \new_[35298]_  = ~A301 & ~A300;
  assign \new_[35299]_  = \new_[35298]_  & \new_[35295]_ ;
  assign \new_[35300]_  = \new_[35299]_  & \new_[35292]_ ;
  assign \new_[35304]_  = ~A166 & ~A167;
  assign \new_[35305]_  = ~A169 & \new_[35304]_ ;
  assign \new_[35309]_  = A203 & A200;
  assign \new_[35310]_  = ~A199 & \new_[35309]_ ;
  assign \new_[35311]_  = \new_[35310]_  & \new_[35305]_ ;
  assign \new_[35315]_  = ~A235 & ~A233;
  assign \new_[35316]_  = ~A232 & \new_[35315]_ ;
  assign \new_[35319]_  = ~A268 & ~A267;
  assign \new_[35322]_  = A301 & ~A269;
  assign \new_[35323]_  = \new_[35322]_  & \new_[35319]_ ;
  assign \new_[35324]_  = \new_[35323]_  & \new_[35316]_ ;
  assign \new_[35328]_  = ~A166 & ~A167;
  assign \new_[35329]_  = ~A169 & \new_[35328]_ ;
  assign \new_[35333]_  = A203 & A200;
  assign \new_[35334]_  = ~A199 & \new_[35333]_ ;
  assign \new_[35335]_  = \new_[35334]_  & \new_[35329]_ ;
  assign \new_[35339]_  = ~A235 & ~A233;
  assign \new_[35340]_  = ~A232 & \new_[35339]_ ;
  assign \new_[35343]_  = ~A266 & ~A265;
  assign \new_[35346]_  = A301 & ~A268;
  assign \new_[35347]_  = \new_[35346]_  & \new_[35343]_ ;
  assign \new_[35348]_  = \new_[35347]_  & \new_[35340]_ ;
  assign \new_[35352]_  = ~A166 & ~A167;
  assign \new_[35353]_  = ~A169 & \new_[35352]_ ;
  assign \new_[35357]_  = A203 & ~A200;
  assign \new_[35358]_  = A199 & \new_[35357]_ ;
  assign \new_[35359]_  = \new_[35358]_  & \new_[35353]_ ;
  assign \new_[35363]_  = ~A236 & ~A235;
  assign \new_[35364]_  = ~A234 & \new_[35363]_ ;
  assign \new_[35367]_  = ~A268 & ~A267;
  assign \new_[35370]_  = A301 & ~A269;
  assign \new_[35371]_  = \new_[35370]_  & \new_[35367]_ ;
  assign \new_[35372]_  = \new_[35371]_  & \new_[35364]_ ;
  assign \new_[35376]_  = ~A166 & ~A167;
  assign \new_[35377]_  = ~A169 & \new_[35376]_ ;
  assign \new_[35381]_  = A203 & ~A200;
  assign \new_[35382]_  = A199 & \new_[35381]_ ;
  assign \new_[35383]_  = \new_[35382]_  & \new_[35377]_ ;
  assign \new_[35387]_  = ~A236 & ~A235;
  assign \new_[35388]_  = ~A234 & \new_[35387]_ ;
  assign \new_[35391]_  = ~A266 & ~A265;
  assign \new_[35394]_  = A301 & ~A268;
  assign \new_[35395]_  = \new_[35394]_  & \new_[35391]_ ;
  assign \new_[35396]_  = \new_[35395]_  & \new_[35388]_ ;
  assign \new_[35400]_  = ~A166 & ~A167;
  assign \new_[35401]_  = ~A169 & \new_[35400]_ ;
  assign \new_[35405]_  = A203 & ~A200;
  assign \new_[35406]_  = A199 & \new_[35405]_ ;
  assign \new_[35407]_  = \new_[35406]_  & \new_[35401]_ ;
  assign \new_[35411]_  = A236 & A233;
  assign \new_[35412]_  = ~A232 & \new_[35411]_ ;
  assign \new_[35415]_  = A299 & A298;
  assign \new_[35418]_  = ~A301 & ~A300;
  assign \new_[35419]_  = \new_[35418]_  & \new_[35415]_ ;
  assign \new_[35420]_  = \new_[35419]_  & \new_[35412]_ ;
  assign \new_[35424]_  = ~A166 & ~A167;
  assign \new_[35425]_  = ~A169 & \new_[35424]_ ;
  assign \new_[35429]_  = A203 & ~A200;
  assign \new_[35430]_  = A199 & \new_[35429]_ ;
  assign \new_[35431]_  = \new_[35430]_  & \new_[35425]_ ;
  assign \new_[35435]_  = A236 & ~A233;
  assign \new_[35436]_  = A232 & \new_[35435]_ ;
  assign \new_[35439]_  = A299 & A298;
  assign \new_[35442]_  = ~A301 & ~A300;
  assign \new_[35443]_  = \new_[35442]_  & \new_[35439]_ ;
  assign \new_[35444]_  = \new_[35443]_  & \new_[35436]_ ;
  assign \new_[35448]_  = ~A166 & ~A167;
  assign \new_[35449]_  = ~A169 & \new_[35448]_ ;
  assign \new_[35453]_  = A203 & ~A200;
  assign \new_[35454]_  = A199 & \new_[35453]_ ;
  assign \new_[35455]_  = \new_[35454]_  & \new_[35449]_ ;
  assign \new_[35459]_  = ~A235 & ~A233;
  assign \new_[35460]_  = ~A232 & \new_[35459]_ ;
  assign \new_[35463]_  = ~A268 & ~A267;
  assign \new_[35466]_  = A301 & ~A269;
  assign \new_[35467]_  = \new_[35466]_  & \new_[35463]_ ;
  assign \new_[35468]_  = \new_[35467]_  & \new_[35460]_ ;
  assign \new_[35472]_  = ~A166 & ~A167;
  assign \new_[35473]_  = ~A169 & \new_[35472]_ ;
  assign \new_[35477]_  = A203 & ~A200;
  assign \new_[35478]_  = A199 & \new_[35477]_ ;
  assign \new_[35479]_  = \new_[35478]_  & \new_[35473]_ ;
  assign \new_[35483]_  = ~A235 & ~A233;
  assign \new_[35484]_  = ~A232 & \new_[35483]_ ;
  assign \new_[35487]_  = ~A266 & ~A265;
  assign \new_[35490]_  = A301 & ~A268;
  assign \new_[35491]_  = \new_[35490]_  & \new_[35487]_ ;
  assign \new_[35492]_  = \new_[35491]_  & \new_[35484]_ ;
  assign \new_[35496]_  = A167 & ~A168;
  assign \new_[35497]_  = ~A169 & \new_[35496]_ ;
  assign \new_[35501]_  = ~A234 & A202;
  assign \new_[35502]_  = A166 & \new_[35501]_ ;
  assign \new_[35503]_  = \new_[35502]_  & \new_[35497]_ ;
  assign \new_[35507]_  = ~A267 & ~A236;
  assign \new_[35508]_  = ~A235 & \new_[35507]_ ;
  assign \new_[35511]_  = ~A269 & ~A268;
  assign \new_[35514]_  = A300 & A299;
  assign \new_[35515]_  = \new_[35514]_  & \new_[35511]_ ;
  assign \new_[35516]_  = \new_[35515]_  & \new_[35508]_ ;
  assign \new_[35520]_  = A167 & ~A168;
  assign \new_[35521]_  = ~A169 & \new_[35520]_ ;
  assign \new_[35525]_  = ~A234 & A202;
  assign \new_[35526]_  = A166 & \new_[35525]_ ;
  assign \new_[35527]_  = \new_[35526]_  & \new_[35521]_ ;
  assign \new_[35531]_  = ~A267 & ~A236;
  assign \new_[35532]_  = ~A235 & \new_[35531]_ ;
  assign \new_[35535]_  = ~A269 & ~A268;
  assign \new_[35538]_  = A300 & A298;
  assign \new_[35539]_  = \new_[35538]_  & \new_[35535]_ ;
  assign \new_[35540]_  = \new_[35539]_  & \new_[35532]_ ;
  assign \new_[35544]_  = A167 & ~A168;
  assign \new_[35545]_  = ~A169 & \new_[35544]_ ;
  assign \new_[35549]_  = ~A234 & A202;
  assign \new_[35550]_  = A166 & \new_[35549]_ ;
  assign \new_[35551]_  = \new_[35550]_  & \new_[35545]_ ;
  assign \new_[35555]_  = A265 & ~A236;
  assign \new_[35556]_  = ~A235 & \new_[35555]_ ;
  assign \new_[35559]_  = ~A267 & A266;
  assign \new_[35562]_  = A301 & ~A268;
  assign \new_[35563]_  = \new_[35562]_  & \new_[35559]_ ;
  assign \new_[35564]_  = \new_[35563]_  & \new_[35556]_ ;
  assign \new_[35568]_  = A167 & ~A168;
  assign \new_[35569]_  = ~A169 & \new_[35568]_ ;
  assign \new_[35573]_  = ~A234 & A202;
  assign \new_[35574]_  = A166 & \new_[35573]_ ;
  assign \new_[35575]_  = \new_[35574]_  & \new_[35569]_ ;
  assign \new_[35579]_  = ~A265 & ~A236;
  assign \new_[35580]_  = ~A235 & \new_[35579]_ ;
  assign \new_[35583]_  = ~A268 & ~A266;
  assign \new_[35586]_  = A300 & A299;
  assign \new_[35587]_  = \new_[35586]_  & \new_[35583]_ ;
  assign \new_[35588]_  = \new_[35587]_  & \new_[35580]_ ;
  assign \new_[35592]_  = A167 & ~A168;
  assign \new_[35593]_  = ~A169 & \new_[35592]_ ;
  assign \new_[35597]_  = ~A234 & A202;
  assign \new_[35598]_  = A166 & \new_[35597]_ ;
  assign \new_[35599]_  = \new_[35598]_  & \new_[35593]_ ;
  assign \new_[35603]_  = ~A265 & ~A236;
  assign \new_[35604]_  = ~A235 & \new_[35603]_ ;
  assign \new_[35607]_  = ~A268 & ~A266;
  assign \new_[35610]_  = A300 & A298;
  assign \new_[35611]_  = \new_[35610]_  & \new_[35607]_ ;
  assign \new_[35612]_  = \new_[35611]_  & \new_[35604]_ ;
  assign \new_[35616]_  = A167 & ~A168;
  assign \new_[35617]_  = ~A169 & \new_[35616]_ ;
  assign \new_[35621]_  = A232 & A202;
  assign \new_[35622]_  = A166 & \new_[35621]_ ;
  assign \new_[35623]_  = \new_[35622]_  & \new_[35617]_ ;
  assign \new_[35627]_  = ~A235 & ~A234;
  assign \new_[35628]_  = A233 & \new_[35627]_ ;
  assign \new_[35631]_  = ~A268 & ~A267;
  assign \new_[35634]_  = A301 & ~A269;
  assign \new_[35635]_  = \new_[35634]_  & \new_[35631]_ ;
  assign \new_[35636]_  = \new_[35635]_  & \new_[35628]_ ;
  assign \new_[35640]_  = A167 & ~A168;
  assign \new_[35641]_  = ~A169 & \new_[35640]_ ;
  assign \new_[35645]_  = A232 & A202;
  assign \new_[35646]_  = A166 & \new_[35645]_ ;
  assign \new_[35647]_  = \new_[35646]_  & \new_[35641]_ ;
  assign \new_[35651]_  = ~A235 & ~A234;
  assign \new_[35652]_  = A233 & \new_[35651]_ ;
  assign \new_[35655]_  = ~A266 & ~A265;
  assign \new_[35658]_  = A301 & ~A268;
  assign \new_[35659]_  = \new_[35658]_  & \new_[35655]_ ;
  assign \new_[35660]_  = \new_[35659]_  & \new_[35652]_ ;
  assign \new_[35664]_  = A167 & ~A168;
  assign \new_[35665]_  = ~A169 & \new_[35664]_ ;
  assign \new_[35669]_  = ~A232 & A202;
  assign \new_[35670]_  = A166 & \new_[35669]_ ;
  assign \new_[35671]_  = \new_[35670]_  & \new_[35665]_ ;
  assign \new_[35675]_  = ~A267 & ~A235;
  assign \new_[35676]_  = ~A233 & \new_[35675]_ ;
  assign \new_[35679]_  = ~A269 & ~A268;
  assign \new_[35682]_  = A300 & A299;
  assign \new_[35683]_  = \new_[35682]_  & \new_[35679]_ ;
  assign \new_[35684]_  = \new_[35683]_  & \new_[35676]_ ;
  assign \new_[35688]_  = A167 & ~A168;
  assign \new_[35689]_  = ~A169 & \new_[35688]_ ;
  assign \new_[35693]_  = ~A232 & A202;
  assign \new_[35694]_  = A166 & \new_[35693]_ ;
  assign \new_[35695]_  = \new_[35694]_  & \new_[35689]_ ;
  assign \new_[35699]_  = ~A267 & ~A235;
  assign \new_[35700]_  = ~A233 & \new_[35699]_ ;
  assign \new_[35703]_  = ~A269 & ~A268;
  assign \new_[35706]_  = A300 & A298;
  assign \new_[35707]_  = \new_[35706]_  & \new_[35703]_ ;
  assign \new_[35708]_  = \new_[35707]_  & \new_[35700]_ ;
  assign \new_[35712]_  = A167 & ~A168;
  assign \new_[35713]_  = ~A169 & \new_[35712]_ ;
  assign \new_[35717]_  = ~A232 & A202;
  assign \new_[35718]_  = A166 & \new_[35717]_ ;
  assign \new_[35719]_  = \new_[35718]_  & \new_[35713]_ ;
  assign \new_[35723]_  = A265 & ~A235;
  assign \new_[35724]_  = ~A233 & \new_[35723]_ ;
  assign \new_[35727]_  = ~A267 & A266;
  assign \new_[35730]_  = A301 & ~A268;
  assign \new_[35731]_  = \new_[35730]_  & \new_[35727]_ ;
  assign \new_[35732]_  = \new_[35731]_  & \new_[35724]_ ;
  assign \new_[35736]_  = A167 & ~A168;
  assign \new_[35737]_  = ~A169 & \new_[35736]_ ;
  assign \new_[35741]_  = ~A232 & A202;
  assign \new_[35742]_  = A166 & \new_[35741]_ ;
  assign \new_[35743]_  = \new_[35742]_  & \new_[35737]_ ;
  assign \new_[35747]_  = ~A265 & ~A235;
  assign \new_[35748]_  = ~A233 & \new_[35747]_ ;
  assign \new_[35751]_  = ~A268 & ~A266;
  assign \new_[35754]_  = A300 & A299;
  assign \new_[35755]_  = \new_[35754]_  & \new_[35751]_ ;
  assign \new_[35756]_  = \new_[35755]_  & \new_[35748]_ ;
  assign \new_[35760]_  = A167 & ~A168;
  assign \new_[35761]_  = ~A169 & \new_[35760]_ ;
  assign \new_[35765]_  = ~A232 & A202;
  assign \new_[35766]_  = A166 & \new_[35765]_ ;
  assign \new_[35767]_  = \new_[35766]_  & \new_[35761]_ ;
  assign \new_[35771]_  = ~A265 & ~A235;
  assign \new_[35772]_  = ~A233 & \new_[35771]_ ;
  assign \new_[35775]_  = ~A268 & ~A266;
  assign \new_[35778]_  = A300 & A298;
  assign \new_[35779]_  = \new_[35778]_  & \new_[35775]_ ;
  assign \new_[35780]_  = \new_[35779]_  & \new_[35772]_ ;
  assign \new_[35784]_  = A167 & ~A168;
  assign \new_[35785]_  = ~A169 & \new_[35784]_ ;
  assign \new_[35789]_  = A201 & A199;
  assign \new_[35790]_  = A166 & \new_[35789]_ ;
  assign \new_[35791]_  = \new_[35790]_  & \new_[35785]_ ;
  assign \new_[35795]_  = ~A236 & ~A235;
  assign \new_[35796]_  = ~A234 & \new_[35795]_ ;
  assign \new_[35799]_  = ~A268 & ~A267;
  assign \new_[35802]_  = A301 & ~A269;
  assign \new_[35803]_  = \new_[35802]_  & \new_[35799]_ ;
  assign \new_[35804]_  = \new_[35803]_  & \new_[35796]_ ;
  assign \new_[35808]_  = A167 & ~A168;
  assign \new_[35809]_  = ~A169 & \new_[35808]_ ;
  assign \new_[35813]_  = A201 & A199;
  assign \new_[35814]_  = A166 & \new_[35813]_ ;
  assign \new_[35815]_  = \new_[35814]_  & \new_[35809]_ ;
  assign \new_[35819]_  = ~A236 & ~A235;
  assign \new_[35820]_  = ~A234 & \new_[35819]_ ;
  assign \new_[35823]_  = ~A266 & ~A265;
  assign \new_[35826]_  = A301 & ~A268;
  assign \new_[35827]_  = \new_[35826]_  & \new_[35823]_ ;
  assign \new_[35828]_  = \new_[35827]_  & \new_[35820]_ ;
  assign \new_[35832]_  = A167 & ~A168;
  assign \new_[35833]_  = ~A169 & \new_[35832]_ ;
  assign \new_[35837]_  = A201 & A199;
  assign \new_[35838]_  = A166 & \new_[35837]_ ;
  assign \new_[35839]_  = \new_[35838]_  & \new_[35833]_ ;
  assign \new_[35843]_  = A236 & A233;
  assign \new_[35844]_  = ~A232 & \new_[35843]_ ;
  assign \new_[35847]_  = A299 & A298;
  assign \new_[35850]_  = ~A301 & ~A300;
  assign \new_[35851]_  = \new_[35850]_  & \new_[35847]_ ;
  assign \new_[35852]_  = \new_[35851]_  & \new_[35844]_ ;
  assign \new_[35856]_  = A167 & ~A168;
  assign \new_[35857]_  = ~A169 & \new_[35856]_ ;
  assign \new_[35861]_  = A201 & A199;
  assign \new_[35862]_  = A166 & \new_[35861]_ ;
  assign \new_[35863]_  = \new_[35862]_  & \new_[35857]_ ;
  assign \new_[35867]_  = A236 & ~A233;
  assign \new_[35868]_  = A232 & \new_[35867]_ ;
  assign \new_[35871]_  = A299 & A298;
  assign \new_[35874]_  = ~A301 & ~A300;
  assign \new_[35875]_  = \new_[35874]_  & \new_[35871]_ ;
  assign \new_[35876]_  = \new_[35875]_  & \new_[35868]_ ;
  assign \new_[35880]_  = A167 & ~A168;
  assign \new_[35881]_  = ~A169 & \new_[35880]_ ;
  assign \new_[35885]_  = A201 & A199;
  assign \new_[35886]_  = A166 & \new_[35885]_ ;
  assign \new_[35887]_  = \new_[35886]_  & \new_[35881]_ ;
  assign \new_[35891]_  = ~A235 & ~A233;
  assign \new_[35892]_  = ~A232 & \new_[35891]_ ;
  assign \new_[35895]_  = ~A268 & ~A267;
  assign \new_[35898]_  = A301 & ~A269;
  assign \new_[35899]_  = \new_[35898]_  & \new_[35895]_ ;
  assign \new_[35900]_  = \new_[35899]_  & \new_[35892]_ ;
  assign \new_[35904]_  = A167 & ~A168;
  assign \new_[35905]_  = ~A169 & \new_[35904]_ ;
  assign \new_[35909]_  = A201 & A199;
  assign \new_[35910]_  = A166 & \new_[35909]_ ;
  assign \new_[35911]_  = \new_[35910]_  & \new_[35905]_ ;
  assign \new_[35915]_  = ~A235 & ~A233;
  assign \new_[35916]_  = ~A232 & \new_[35915]_ ;
  assign \new_[35919]_  = ~A266 & ~A265;
  assign \new_[35922]_  = A301 & ~A268;
  assign \new_[35923]_  = \new_[35922]_  & \new_[35919]_ ;
  assign \new_[35924]_  = \new_[35923]_  & \new_[35916]_ ;
  assign \new_[35928]_  = A167 & ~A168;
  assign \new_[35929]_  = ~A169 & \new_[35928]_ ;
  assign \new_[35933]_  = A201 & A200;
  assign \new_[35934]_  = A166 & \new_[35933]_ ;
  assign \new_[35935]_  = \new_[35934]_  & \new_[35929]_ ;
  assign \new_[35939]_  = ~A236 & ~A235;
  assign \new_[35940]_  = ~A234 & \new_[35939]_ ;
  assign \new_[35943]_  = ~A268 & ~A267;
  assign \new_[35946]_  = A301 & ~A269;
  assign \new_[35947]_  = \new_[35946]_  & \new_[35943]_ ;
  assign \new_[35948]_  = \new_[35947]_  & \new_[35940]_ ;
  assign \new_[35952]_  = A167 & ~A168;
  assign \new_[35953]_  = ~A169 & \new_[35952]_ ;
  assign \new_[35957]_  = A201 & A200;
  assign \new_[35958]_  = A166 & \new_[35957]_ ;
  assign \new_[35959]_  = \new_[35958]_  & \new_[35953]_ ;
  assign \new_[35963]_  = ~A236 & ~A235;
  assign \new_[35964]_  = ~A234 & \new_[35963]_ ;
  assign \new_[35967]_  = ~A266 & ~A265;
  assign \new_[35970]_  = A301 & ~A268;
  assign \new_[35971]_  = \new_[35970]_  & \new_[35967]_ ;
  assign \new_[35972]_  = \new_[35971]_  & \new_[35964]_ ;
  assign \new_[35976]_  = A167 & ~A168;
  assign \new_[35977]_  = ~A169 & \new_[35976]_ ;
  assign \new_[35981]_  = A201 & A200;
  assign \new_[35982]_  = A166 & \new_[35981]_ ;
  assign \new_[35983]_  = \new_[35982]_  & \new_[35977]_ ;
  assign \new_[35987]_  = A236 & A233;
  assign \new_[35988]_  = ~A232 & \new_[35987]_ ;
  assign \new_[35991]_  = A299 & A298;
  assign \new_[35994]_  = ~A301 & ~A300;
  assign \new_[35995]_  = \new_[35994]_  & \new_[35991]_ ;
  assign \new_[35996]_  = \new_[35995]_  & \new_[35988]_ ;
  assign \new_[36000]_  = A167 & ~A168;
  assign \new_[36001]_  = ~A169 & \new_[36000]_ ;
  assign \new_[36005]_  = A201 & A200;
  assign \new_[36006]_  = A166 & \new_[36005]_ ;
  assign \new_[36007]_  = \new_[36006]_  & \new_[36001]_ ;
  assign \new_[36011]_  = A236 & ~A233;
  assign \new_[36012]_  = A232 & \new_[36011]_ ;
  assign \new_[36015]_  = A299 & A298;
  assign \new_[36018]_  = ~A301 & ~A300;
  assign \new_[36019]_  = \new_[36018]_  & \new_[36015]_ ;
  assign \new_[36020]_  = \new_[36019]_  & \new_[36012]_ ;
  assign \new_[36024]_  = A167 & ~A168;
  assign \new_[36025]_  = ~A169 & \new_[36024]_ ;
  assign \new_[36029]_  = A201 & A200;
  assign \new_[36030]_  = A166 & \new_[36029]_ ;
  assign \new_[36031]_  = \new_[36030]_  & \new_[36025]_ ;
  assign \new_[36035]_  = ~A235 & ~A233;
  assign \new_[36036]_  = ~A232 & \new_[36035]_ ;
  assign \new_[36039]_  = ~A268 & ~A267;
  assign \new_[36042]_  = A301 & ~A269;
  assign \new_[36043]_  = \new_[36042]_  & \new_[36039]_ ;
  assign \new_[36044]_  = \new_[36043]_  & \new_[36036]_ ;
  assign \new_[36048]_  = A167 & ~A168;
  assign \new_[36049]_  = ~A169 & \new_[36048]_ ;
  assign \new_[36053]_  = A201 & A200;
  assign \new_[36054]_  = A166 & \new_[36053]_ ;
  assign \new_[36055]_  = \new_[36054]_  & \new_[36049]_ ;
  assign \new_[36059]_  = ~A235 & ~A233;
  assign \new_[36060]_  = ~A232 & \new_[36059]_ ;
  assign \new_[36063]_  = ~A266 & ~A265;
  assign \new_[36066]_  = A301 & ~A268;
  assign \new_[36067]_  = \new_[36066]_  & \new_[36063]_ ;
  assign \new_[36068]_  = \new_[36067]_  & \new_[36060]_ ;
  assign \new_[36072]_  = A167 & ~A168;
  assign \new_[36073]_  = ~A169 & \new_[36072]_ ;
  assign \new_[36077]_  = A200 & ~A199;
  assign \new_[36078]_  = A166 & \new_[36077]_ ;
  assign \new_[36079]_  = \new_[36078]_  & \new_[36073]_ ;
  assign \new_[36083]_  = A234 & A232;
  assign \new_[36084]_  = A203 & \new_[36083]_ ;
  assign \new_[36087]_  = A299 & A298;
  assign \new_[36090]_  = ~A301 & ~A300;
  assign \new_[36091]_  = \new_[36090]_  & \new_[36087]_ ;
  assign \new_[36092]_  = \new_[36091]_  & \new_[36084]_ ;
  assign \new_[36096]_  = A167 & ~A168;
  assign \new_[36097]_  = ~A169 & \new_[36096]_ ;
  assign \new_[36101]_  = A200 & ~A199;
  assign \new_[36102]_  = A166 & \new_[36101]_ ;
  assign \new_[36103]_  = \new_[36102]_  & \new_[36097]_ ;
  assign \new_[36107]_  = A234 & A233;
  assign \new_[36108]_  = A203 & \new_[36107]_ ;
  assign \new_[36111]_  = A299 & A298;
  assign \new_[36114]_  = ~A301 & ~A300;
  assign \new_[36115]_  = \new_[36114]_  & \new_[36111]_ ;
  assign \new_[36116]_  = \new_[36115]_  & \new_[36108]_ ;
  assign \new_[36120]_  = A167 & ~A168;
  assign \new_[36121]_  = ~A169 & \new_[36120]_ ;
  assign \new_[36125]_  = A200 & ~A199;
  assign \new_[36126]_  = A166 & \new_[36125]_ ;
  assign \new_[36127]_  = \new_[36126]_  & \new_[36121]_ ;
  assign \new_[36131]_  = A233 & ~A232;
  assign \new_[36132]_  = A203 & \new_[36131]_ ;
  assign \new_[36135]_  = ~A300 & A236;
  assign \new_[36138]_  = ~A302 & ~A301;
  assign \new_[36139]_  = \new_[36138]_  & \new_[36135]_ ;
  assign \new_[36140]_  = \new_[36139]_  & \new_[36132]_ ;
  assign \new_[36144]_  = A167 & ~A168;
  assign \new_[36145]_  = ~A169 & \new_[36144]_ ;
  assign \new_[36149]_  = A200 & ~A199;
  assign \new_[36150]_  = A166 & \new_[36149]_ ;
  assign \new_[36151]_  = \new_[36150]_  & \new_[36145]_ ;
  assign \new_[36155]_  = A233 & ~A232;
  assign \new_[36156]_  = A203 & \new_[36155]_ ;
  assign \new_[36159]_  = ~A298 & A236;
  assign \new_[36162]_  = ~A301 & ~A299;
  assign \new_[36163]_  = \new_[36162]_  & \new_[36159]_ ;
  assign \new_[36164]_  = \new_[36163]_  & \new_[36156]_ ;
  assign \new_[36168]_  = A167 & ~A168;
  assign \new_[36169]_  = ~A169 & \new_[36168]_ ;
  assign \new_[36173]_  = A200 & ~A199;
  assign \new_[36174]_  = A166 & \new_[36173]_ ;
  assign \new_[36175]_  = \new_[36174]_  & \new_[36169]_ ;
  assign \new_[36179]_  = A233 & ~A232;
  assign \new_[36180]_  = A203 & \new_[36179]_ ;
  assign \new_[36183]_  = ~A265 & A236;
  assign \new_[36186]_  = A269 & A266;
  assign \new_[36187]_  = \new_[36186]_  & \new_[36183]_ ;
  assign \new_[36188]_  = \new_[36187]_  & \new_[36180]_ ;
  assign \new_[36192]_  = A167 & ~A168;
  assign \new_[36193]_  = ~A169 & \new_[36192]_ ;
  assign \new_[36197]_  = A200 & ~A199;
  assign \new_[36198]_  = A166 & \new_[36197]_ ;
  assign \new_[36199]_  = \new_[36198]_  & \new_[36193]_ ;
  assign \new_[36203]_  = A233 & ~A232;
  assign \new_[36204]_  = A203 & \new_[36203]_ ;
  assign \new_[36207]_  = A265 & A236;
  assign \new_[36210]_  = A269 & ~A266;
  assign \new_[36211]_  = \new_[36210]_  & \new_[36207]_ ;
  assign \new_[36212]_  = \new_[36211]_  & \new_[36204]_ ;
  assign \new_[36216]_  = A167 & ~A168;
  assign \new_[36217]_  = ~A169 & \new_[36216]_ ;
  assign \new_[36221]_  = A200 & ~A199;
  assign \new_[36222]_  = A166 & \new_[36221]_ ;
  assign \new_[36223]_  = \new_[36222]_  & \new_[36217]_ ;
  assign \new_[36227]_  = ~A233 & A232;
  assign \new_[36228]_  = A203 & \new_[36227]_ ;
  assign \new_[36231]_  = ~A300 & A236;
  assign \new_[36234]_  = ~A302 & ~A301;
  assign \new_[36235]_  = \new_[36234]_  & \new_[36231]_ ;
  assign \new_[36236]_  = \new_[36235]_  & \new_[36228]_ ;
  assign \new_[36240]_  = A167 & ~A168;
  assign \new_[36241]_  = ~A169 & \new_[36240]_ ;
  assign \new_[36245]_  = A200 & ~A199;
  assign \new_[36246]_  = A166 & \new_[36245]_ ;
  assign \new_[36247]_  = \new_[36246]_  & \new_[36241]_ ;
  assign \new_[36251]_  = ~A233 & A232;
  assign \new_[36252]_  = A203 & \new_[36251]_ ;
  assign \new_[36255]_  = ~A298 & A236;
  assign \new_[36258]_  = ~A301 & ~A299;
  assign \new_[36259]_  = \new_[36258]_  & \new_[36255]_ ;
  assign \new_[36260]_  = \new_[36259]_  & \new_[36252]_ ;
  assign \new_[36264]_  = A167 & ~A168;
  assign \new_[36265]_  = ~A169 & \new_[36264]_ ;
  assign \new_[36269]_  = A200 & ~A199;
  assign \new_[36270]_  = A166 & \new_[36269]_ ;
  assign \new_[36271]_  = \new_[36270]_  & \new_[36265]_ ;
  assign \new_[36275]_  = ~A233 & A232;
  assign \new_[36276]_  = A203 & \new_[36275]_ ;
  assign \new_[36279]_  = ~A265 & A236;
  assign \new_[36282]_  = A269 & A266;
  assign \new_[36283]_  = \new_[36282]_  & \new_[36279]_ ;
  assign \new_[36284]_  = \new_[36283]_  & \new_[36276]_ ;
  assign \new_[36288]_  = A167 & ~A168;
  assign \new_[36289]_  = ~A169 & \new_[36288]_ ;
  assign \new_[36293]_  = A200 & ~A199;
  assign \new_[36294]_  = A166 & \new_[36293]_ ;
  assign \new_[36295]_  = \new_[36294]_  & \new_[36289]_ ;
  assign \new_[36299]_  = ~A233 & A232;
  assign \new_[36300]_  = A203 & \new_[36299]_ ;
  assign \new_[36303]_  = A265 & A236;
  assign \new_[36306]_  = A269 & ~A266;
  assign \new_[36307]_  = \new_[36306]_  & \new_[36303]_ ;
  assign \new_[36308]_  = \new_[36307]_  & \new_[36300]_ ;
  assign \new_[36312]_  = A167 & ~A168;
  assign \new_[36313]_  = ~A169 & \new_[36312]_ ;
  assign \new_[36317]_  = ~A200 & A199;
  assign \new_[36318]_  = A166 & \new_[36317]_ ;
  assign \new_[36319]_  = \new_[36318]_  & \new_[36313]_ ;
  assign \new_[36323]_  = A234 & A232;
  assign \new_[36324]_  = A203 & \new_[36323]_ ;
  assign \new_[36327]_  = A299 & A298;
  assign \new_[36330]_  = ~A301 & ~A300;
  assign \new_[36331]_  = \new_[36330]_  & \new_[36327]_ ;
  assign \new_[36332]_  = \new_[36331]_  & \new_[36324]_ ;
  assign \new_[36336]_  = A167 & ~A168;
  assign \new_[36337]_  = ~A169 & \new_[36336]_ ;
  assign \new_[36341]_  = ~A200 & A199;
  assign \new_[36342]_  = A166 & \new_[36341]_ ;
  assign \new_[36343]_  = \new_[36342]_  & \new_[36337]_ ;
  assign \new_[36347]_  = A234 & A233;
  assign \new_[36348]_  = A203 & \new_[36347]_ ;
  assign \new_[36351]_  = A299 & A298;
  assign \new_[36354]_  = ~A301 & ~A300;
  assign \new_[36355]_  = \new_[36354]_  & \new_[36351]_ ;
  assign \new_[36356]_  = \new_[36355]_  & \new_[36348]_ ;
  assign \new_[36360]_  = A167 & ~A168;
  assign \new_[36361]_  = ~A169 & \new_[36360]_ ;
  assign \new_[36365]_  = ~A200 & A199;
  assign \new_[36366]_  = A166 & \new_[36365]_ ;
  assign \new_[36367]_  = \new_[36366]_  & \new_[36361]_ ;
  assign \new_[36371]_  = A233 & ~A232;
  assign \new_[36372]_  = A203 & \new_[36371]_ ;
  assign \new_[36375]_  = ~A300 & A236;
  assign \new_[36378]_  = ~A302 & ~A301;
  assign \new_[36379]_  = \new_[36378]_  & \new_[36375]_ ;
  assign \new_[36380]_  = \new_[36379]_  & \new_[36372]_ ;
  assign \new_[36384]_  = A167 & ~A168;
  assign \new_[36385]_  = ~A169 & \new_[36384]_ ;
  assign \new_[36389]_  = ~A200 & A199;
  assign \new_[36390]_  = A166 & \new_[36389]_ ;
  assign \new_[36391]_  = \new_[36390]_  & \new_[36385]_ ;
  assign \new_[36395]_  = A233 & ~A232;
  assign \new_[36396]_  = A203 & \new_[36395]_ ;
  assign \new_[36399]_  = ~A298 & A236;
  assign \new_[36402]_  = ~A301 & ~A299;
  assign \new_[36403]_  = \new_[36402]_  & \new_[36399]_ ;
  assign \new_[36404]_  = \new_[36403]_  & \new_[36396]_ ;
  assign \new_[36408]_  = A167 & ~A168;
  assign \new_[36409]_  = ~A169 & \new_[36408]_ ;
  assign \new_[36413]_  = ~A200 & A199;
  assign \new_[36414]_  = A166 & \new_[36413]_ ;
  assign \new_[36415]_  = \new_[36414]_  & \new_[36409]_ ;
  assign \new_[36419]_  = A233 & ~A232;
  assign \new_[36420]_  = A203 & \new_[36419]_ ;
  assign \new_[36423]_  = ~A265 & A236;
  assign \new_[36426]_  = A269 & A266;
  assign \new_[36427]_  = \new_[36426]_  & \new_[36423]_ ;
  assign \new_[36428]_  = \new_[36427]_  & \new_[36420]_ ;
  assign \new_[36432]_  = A167 & ~A168;
  assign \new_[36433]_  = ~A169 & \new_[36432]_ ;
  assign \new_[36437]_  = ~A200 & A199;
  assign \new_[36438]_  = A166 & \new_[36437]_ ;
  assign \new_[36439]_  = \new_[36438]_  & \new_[36433]_ ;
  assign \new_[36443]_  = A233 & ~A232;
  assign \new_[36444]_  = A203 & \new_[36443]_ ;
  assign \new_[36447]_  = A265 & A236;
  assign \new_[36450]_  = A269 & ~A266;
  assign \new_[36451]_  = \new_[36450]_  & \new_[36447]_ ;
  assign \new_[36452]_  = \new_[36451]_  & \new_[36444]_ ;
  assign \new_[36456]_  = A167 & ~A168;
  assign \new_[36457]_  = ~A169 & \new_[36456]_ ;
  assign \new_[36461]_  = ~A200 & A199;
  assign \new_[36462]_  = A166 & \new_[36461]_ ;
  assign \new_[36463]_  = \new_[36462]_  & \new_[36457]_ ;
  assign \new_[36467]_  = ~A233 & A232;
  assign \new_[36468]_  = A203 & \new_[36467]_ ;
  assign \new_[36471]_  = ~A300 & A236;
  assign \new_[36474]_  = ~A302 & ~A301;
  assign \new_[36475]_  = \new_[36474]_  & \new_[36471]_ ;
  assign \new_[36476]_  = \new_[36475]_  & \new_[36468]_ ;
  assign \new_[36480]_  = A167 & ~A168;
  assign \new_[36481]_  = ~A169 & \new_[36480]_ ;
  assign \new_[36485]_  = ~A200 & A199;
  assign \new_[36486]_  = A166 & \new_[36485]_ ;
  assign \new_[36487]_  = \new_[36486]_  & \new_[36481]_ ;
  assign \new_[36491]_  = ~A233 & A232;
  assign \new_[36492]_  = A203 & \new_[36491]_ ;
  assign \new_[36495]_  = ~A298 & A236;
  assign \new_[36498]_  = ~A301 & ~A299;
  assign \new_[36499]_  = \new_[36498]_  & \new_[36495]_ ;
  assign \new_[36500]_  = \new_[36499]_  & \new_[36492]_ ;
  assign \new_[36504]_  = A167 & ~A168;
  assign \new_[36505]_  = ~A169 & \new_[36504]_ ;
  assign \new_[36509]_  = ~A200 & A199;
  assign \new_[36510]_  = A166 & \new_[36509]_ ;
  assign \new_[36511]_  = \new_[36510]_  & \new_[36505]_ ;
  assign \new_[36515]_  = ~A233 & A232;
  assign \new_[36516]_  = A203 & \new_[36515]_ ;
  assign \new_[36519]_  = ~A265 & A236;
  assign \new_[36522]_  = A269 & A266;
  assign \new_[36523]_  = \new_[36522]_  & \new_[36519]_ ;
  assign \new_[36524]_  = \new_[36523]_  & \new_[36516]_ ;
  assign \new_[36528]_  = A167 & ~A168;
  assign \new_[36529]_  = ~A169 & \new_[36528]_ ;
  assign \new_[36533]_  = ~A200 & A199;
  assign \new_[36534]_  = A166 & \new_[36533]_ ;
  assign \new_[36535]_  = \new_[36534]_  & \new_[36529]_ ;
  assign \new_[36539]_  = ~A233 & A232;
  assign \new_[36540]_  = A203 & \new_[36539]_ ;
  assign \new_[36543]_  = A265 & A236;
  assign \new_[36546]_  = A269 & ~A266;
  assign \new_[36547]_  = \new_[36546]_  & \new_[36543]_ ;
  assign \new_[36548]_  = \new_[36547]_  & \new_[36540]_ ;
  assign \new_[36552]_  = ~A168 & ~A169;
  assign \new_[36553]_  = ~A170 & \new_[36552]_ ;
  assign \new_[36557]_  = ~A235 & ~A234;
  assign \new_[36558]_  = A202 & \new_[36557]_ ;
  assign \new_[36559]_  = \new_[36558]_  & \new_[36553]_ ;
  assign \new_[36563]_  = ~A268 & ~A267;
  assign \new_[36564]_  = ~A236 & \new_[36563]_ ;
  assign \new_[36567]_  = A298 & ~A269;
  assign \new_[36570]_  = A302 & ~A299;
  assign \new_[36571]_  = \new_[36570]_  & \new_[36567]_ ;
  assign \new_[36572]_  = \new_[36571]_  & \new_[36564]_ ;
  assign \new_[36576]_  = ~A168 & ~A169;
  assign \new_[36577]_  = ~A170 & \new_[36576]_ ;
  assign \new_[36581]_  = ~A235 & ~A234;
  assign \new_[36582]_  = A202 & \new_[36581]_ ;
  assign \new_[36583]_  = \new_[36582]_  & \new_[36577]_ ;
  assign \new_[36587]_  = ~A268 & ~A267;
  assign \new_[36588]_  = ~A236 & \new_[36587]_ ;
  assign \new_[36591]_  = ~A298 & ~A269;
  assign \new_[36594]_  = A302 & A299;
  assign \new_[36595]_  = \new_[36594]_  & \new_[36591]_ ;
  assign \new_[36596]_  = \new_[36595]_  & \new_[36588]_ ;
  assign \new_[36600]_  = ~A168 & ~A169;
  assign \new_[36601]_  = ~A170 & \new_[36600]_ ;
  assign \new_[36605]_  = ~A235 & ~A234;
  assign \new_[36606]_  = A202 & \new_[36605]_ ;
  assign \new_[36607]_  = \new_[36606]_  & \new_[36601]_ ;
  assign \new_[36611]_  = A266 & A265;
  assign \new_[36612]_  = ~A236 & \new_[36611]_ ;
  assign \new_[36615]_  = ~A268 & ~A267;
  assign \new_[36618]_  = A300 & A299;
  assign \new_[36619]_  = \new_[36618]_  & \new_[36615]_ ;
  assign \new_[36620]_  = \new_[36619]_  & \new_[36612]_ ;
  assign \new_[36624]_  = ~A168 & ~A169;
  assign \new_[36625]_  = ~A170 & \new_[36624]_ ;
  assign \new_[36629]_  = ~A235 & ~A234;
  assign \new_[36630]_  = A202 & \new_[36629]_ ;
  assign \new_[36631]_  = \new_[36630]_  & \new_[36625]_ ;
  assign \new_[36635]_  = A266 & A265;
  assign \new_[36636]_  = ~A236 & \new_[36635]_ ;
  assign \new_[36639]_  = ~A268 & ~A267;
  assign \new_[36642]_  = A300 & A298;
  assign \new_[36643]_  = \new_[36642]_  & \new_[36639]_ ;
  assign \new_[36644]_  = \new_[36643]_  & \new_[36636]_ ;
  assign \new_[36648]_  = ~A168 & ~A169;
  assign \new_[36649]_  = ~A170 & \new_[36648]_ ;
  assign \new_[36653]_  = ~A235 & ~A234;
  assign \new_[36654]_  = A202 & \new_[36653]_ ;
  assign \new_[36655]_  = \new_[36654]_  & \new_[36649]_ ;
  assign \new_[36659]_  = ~A266 & ~A265;
  assign \new_[36660]_  = ~A236 & \new_[36659]_ ;
  assign \new_[36663]_  = A298 & ~A268;
  assign \new_[36666]_  = A302 & ~A299;
  assign \new_[36667]_  = \new_[36666]_  & \new_[36663]_ ;
  assign \new_[36668]_  = \new_[36667]_  & \new_[36660]_ ;
  assign \new_[36672]_  = ~A168 & ~A169;
  assign \new_[36673]_  = ~A170 & \new_[36672]_ ;
  assign \new_[36677]_  = ~A235 & ~A234;
  assign \new_[36678]_  = A202 & \new_[36677]_ ;
  assign \new_[36679]_  = \new_[36678]_  & \new_[36673]_ ;
  assign \new_[36683]_  = ~A266 & ~A265;
  assign \new_[36684]_  = ~A236 & \new_[36683]_ ;
  assign \new_[36687]_  = ~A298 & ~A268;
  assign \new_[36690]_  = A302 & A299;
  assign \new_[36691]_  = \new_[36690]_  & \new_[36687]_ ;
  assign \new_[36692]_  = \new_[36691]_  & \new_[36684]_ ;
  assign \new_[36696]_  = ~A168 & ~A169;
  assign \new_[36697]_  = ~A170 & \new_[36696]_ ;
  assign \new_[36701]_  = A233 & A232;
  assign \new_[36702]_  = A202 & \new_[36701]_ ;
  assign \new_[36703]_  = \new_[36702]_  & \new_[36697]_ ;
  assign \new_[36707]_  = ~A267 & ~A235;
  assign \new_[36708]_  = ~A234 & \new_[36707]_ ;
  assign \new_[36711]_  = ~A269 & ~A268;
  assign \new_[36714]_  = A300 & A299;
  assign \new_[36715]_  = \new_[36714]_  & \new_[36711]_ ;
  assign \new_[36716]_  = \new_[36715]_  & \new_[36708]_ ;
  assign \new_[36720]_  = ~A168 & ~A169;
  assign \new_[36721]_  = ~A170 & \new_[36720]_ ;
  assign \new_[36725]_  = A233 & A232;
  assign \new_[36726]_  = A202 & \new_[36725]_ ;
  assign \new_[36727]_  = \new_[36726]_  & \new_[36721]_ ;
  assign \new_[36731]_  = ~A267 & ~A235;
  assign \new_[36732]_  = ~A234 & \new_[36731]_ ;
  assign \new_[36735]_  = ~A269 & ~A268;
  assign \new_[36738]_  = A300 & A298;
  assign \new_[36739]_  = \new_[36738]_  & \new_[36735]_ ;
  assign \new_[36740]_  = \new_[36739]_  & \new_[36732]_ ;
  assign \new_[36744]_  = ~A168 & ~A169;
  assign \new_[36745]_  = ~A170 & \new_[36744]_ ;
  assign \new_[36749]_  = A233 & A232;
  assign \new_[36750]_  = A202 & \new_[36749]_ ;
  assign \new_[36751]_  = \new_[36750]_  & \new_[36745]_ ;
  assign \new_[36755]_  = A265 & ~A235;
  assign \new_[36756]_  = ~A234 & \new_[36755]_ ;
  assign \new_[36759]_  = ~A267 & A266;
  assign \new_[36762]_  = A301 & ~A268;
  assign \new_[36763]_  = \new_[36762]_  & \new_[36759]_ ;
  assign \new_[36764]_  = \new_[36763]_  & \new_[36756]_ ;
  assign \new_[36768]_  = ~A168 & ~A169;
  assign \new_[36769]_  = ~A170 & \new_[36768]_ ;
  assign \new_[36773]_  = A233 & A232;
  assign \new_[36774]_  = A202 & \new_[36773]_ ;
  assign \new_[36775]_  = \new_[36774]_  & \new_[36769]_ ;
  assign \new_[36779]_  = ~A265 & ~A235;
  assign \new_[36780]_  = ~A234 & \new_[36779]_ ;
  assign \new_[36783]_  = ~A268 & ~A266;
  assign \new_[36786]_  = A300 & A299;
  assign \new_[36787]_  = \new_[36786]_  & \new_[36783]_ ;
  assign \new_[36788]_  = \new_[36787]_  & \new_[36780]_ ;
  assign \new_[36792]_  = ~A168 & ~A169;
  assign \new_[36793]_  = ~A170 & \new_[36792]_ ;
  assign \new_[36797]_  = A233 & A232;
  assign \new_[36798]_  = A202 & \new_[36797]_ ;
  assign \new_[36799]_  = \new_[36798]_  & \new_[36793]_ ;
  assign \new_[36803]_  = ~A265 & ~A235;
  assign \new_[36804]_  = ~A234 & \new_[36803]_ ;
  assign \new_[36807]_  = ~A268 & ~A266;
  assign \new_[36810]_  = A300 & A298;
  assign \new_[36811]_  = \new_[36810]_  & \new_[36807]_ ;
  assign \new_[36812]_  = \new_[36811]_  & \new_[36804]_ ;
  assign \new_[36816]_  = ~A168 & ~A169;
  assign \new_[36817]_  = ~A170 & \new_[36816]_ ;
  assign \new_[36821]_  = ~A233 & ~A232;
  assign \new_[36822]_  = A202 & \new_[36821]_ ;
  assign \new_[36823]_  = \new_[36822]_  & \new_[36817]_ ;
  assign \new_[36827]_  = ~A268 & ~A267;
  assign \new_[36828]_  = ~A235 & \new_[36827]_ ;
  assign \new_[36831]_  = A298 & ~A269;
  assign \new_[36834]_  = A302 & ~A299;
  assign \new_[36835]_  = \new_[36834]_  & \new_[36831]_ ;
  assign \new_[36836]_  = \new_[36835]_  & \new_[36828]_ ;
  assign \new_[36840]_  = ~A168 & ~A169;
  assign \new_[36841]_  = ~A170 & \new_[36840]_ ;
  assign \new_[36845]_  = ~A233 & ~A232;
  assign \new_[36846]_  = A202 & \new_[36845]_ ;
  assign \new_[36847]_  = \new_[36846]_  & \new_[36841]_ ;
  assign \new_[36851]_  = ~A268 & ~A267;
  assign \new_[36852]_  = ~A235 & \new_[36851]_ ;
  assign \new_[36855]_  = ~A298 & ~A269;
  assign \new_[36858]_  = A302 & A299;
  assign \new_[36859]_  = \new_[36858]_  & \new_[36855]_ ;
  assign \new_[36860]_  = \new_[36859]_  & \new_[36852]_ ;
  assign \new_[36864]_  = ~A168 & ~A169;
  assign \new_[36865]_  = ~A170 & \new_[36864]_ ;
  assign \new_[36869]_  = ~A233 & ~A232;
  assign \new_[36870]_  = A202 & \new_[36869]_ ;
  assign \new_[36871]_  = \new_[36870]_  & \new_[36865]_ ;
  assign \new_[36875]_  = A266 & A265;
  assign \new_[36876]_  = ~A235 & \new_[36875]_ ;
  assign \new_[36879]_  = ~A268 & ~A267;
  assign \new_[36882]_  = A300 & A299;
  assign \new_[36883]_  = \new_[36882]_  & \new_[36879]_ ;
  assign \new_[36884]_  = \new_[36883]_  & \new_[36876]_ ;
  assign \new_[36888]_  = ~A168 & ~A169;
  assign \new_[36889]_  = ~A170 & \new_[36888]_ ;
  assign \new_[36893]_  = ~A233 & ~A232;
  assign \new_[36894]_  = A202 & \new_[36893]_ ;
  assign \new_[36895]_  = \new_[36894]_  & \new_[36889]_ ;
  assign \new_[36899]_  = A266 & A265;
  assign \new_[36900]_  = ~A235 & \new_[36899]_ ;
  assign \new_[36903]_  = ~A268 & ~A267;
  assign \new_[36906]_  = A300 & A298;
  assign \new_[36907]_  = \new_[36906]_  & \new_[36903]_ ;
  assign \new_[36908]_  = \new_[36907]_  & \new_[36900]_ ;
  assign \new_[36912]_  = ~A168 & ~A169;
  assign \new_[36913]_  = ~A170 & \new_[36912]_ ;
  assign \new_[36917]_  = ~A233 & ~A232;
  assign \new_[36918]_  = A202 & \new_[36917]_ ;
  assign \new_[36919]_  = \new_[36918]_  & \new_[36913]_ ;
  assign \new_[36923]_  = ~A266 & ~A265;
  assign \new_[36924]_  = ~A235 & \new_[36923]_ ;
  assign \new_[36927]_  = A298 & ~A268;
  assign \new_[36930]_  = A302 & ~A299;
  assign \new_[36931]_  = \new_[36930]_  & \new_[36927]_ ;
  assign \new_[36932]_  = \new_[36931]_  & \new_[36924]_ ;
  assign \new_[36936]_  = ~A168 & ~A169;
  assign \new_[36937]_  = ~A170 & \new_[36936]_ ;
  assign \new_[36941]_  = ~A233 & ~A232;
  assign \new_[36942]_  = A202 & \new_[36941]_ ;
  assign \new_[36943]_  = \new_[36942]_  & \new_[36937]_ ;
  assign \new_[36947]_  = ~A266 & ~A265;
  assign \new_[36948]_  = ~A235 & \new_[36947]_ ;
  assign \new_[36951]_  = ~A298 & ~A268;
  assign \new_[36954]_  = A302 & A299;
  assign \new_[36955]_  = \new_[36954]_  & \new_[36951]_ ;
  assign \new_[36956]_  = \new_[36955]_  & \new_[36948]_ ;
  assign \new_[36960]_  = ~A168 & ~A169;
  assign \new_[36961]_  = ~A170 & \new_[36960]_ ;
  assign \new_[36965]_  = ~A234 & A201;
  assign \new_[36966]_  = A199 & \new_[36965]_ ;
  assign \new_[36967]_  = \new_[36966]_  & \new_[36961]_ ;
  assign \new_[36971]_  = ~A267 & ~A236;
  assign \new_[36972]_  = ~A235 & \new_[36971]_ ;
  assign \new_[36975]_  = ~A269 & ~A268;
  assign \new_[36978]_  = A300 & A299;
  assign \new_[36979]_  = \new_[36978]_  & \new_[36975]_ ;
  assign \new_[36980]_  = \new_[36979]_  & \new_[36972]_ ;
  assign \new_[36984]_  = ~A168 & ~A169;
  assign \new_[36985]_  = ~A170 & \new_[36984]_ ;
  assign \new_[36989]_  = ~A234 & A201;
  assign \new_[36990]_  = A199 & \new_[36989]_ ;
  assign \new_[36991]_  = \new_[36990]_  & \new_[36985]_ ;
  assign \new_[36995]_  = ~A267 & ~A236;
  assign \new_[36996]_  = ~A235 & \new_[36995]_ ;
  assign \new_[36999]_  = ~A269 & ~A268;
  assign \new_[37002]_  = A300 & A298;
  assign \new_[37003]_  = \new_[37002]_  & \new_[36999]_ ;
  assign \new_[37004]_  = \new_[37003]_  & \new_[36996]_ ;
  assign \new_[37008]_  = ~A168 & ~A169;
  assign \new_[37009]_  = ~A170 & \new_[37008]_ ;
  assign \new_[37013]_  = ~A234 & A201;
  assign \new_[37014]_  = A199 & \new_[37013]_ ;
  assign \new_[37015]_  = \new_[37014]_  & \new_[37009]_ ;
  assign \new_[37019]_  = A265 & ~A236;
  assign \new_[37020]_  = ~A235 & \new_[37019]_ ;
  assign \new_[37023]_  = ~A267 & A266;
  assign \new_[37026]_  = A301 & ~A268;
  assign \new_[37027]_  = \new_[37026]_  & \new_[37023]_ ;
  assign \new_[37028]_  = \new_[37027]_  & \new_[37020]_ ;
  assign \new_[37032]_  = ~A168 & ~A169;
  assign \new_[37033]_  = ~A170 & \new_[37032]_ ;
  assign \new_[37037]_  = ~A234 & A201;
  assign \new_[37038]_  = A199 & \new_[37037]_ ;
  assign \new_[37039]_  = \new_[37038]_  & \new_[37033]_ ;
  assign \new_[37043]_  = ~A265 & ~A236;
  assign \new_[37044]_  = ~A235 & \new_[37043]_ ;
  assign \new_[37047]_  = ~A268 & ~A266;
  assign \new_[37050]_  = A300 & A299;
  assign \new_[37051]_  = \new_[37050]_  & \new_[37047]_ ;
  assign \new_[37052]_  = \new_[37051]_  & \new_[37044]_ ;
  assign \new_[37056]_  = ~A168 & ~A169;
  assign \new_[37057]_  = ~A170 & \new_[37056]_ ;
  assign \new_[37061]_  = ~A234 & A201;
  assign \new_[37062]_  = A199 & \new_[37061]_ ;
  assign \new_[37063]_  = \new_[37062]_  & \new_[37057]_ ;
  assign \new_[37067]_  = ~A265 & ~A236;
  assign \new_[37068]_  = ~A235 & \new_[37067]_ ;
  assign \new_[37071]_  = ~A268 & ~A266;
  assign \new_[37074]_  = A300 & A298;
  assign \new_[37075]_  = \new_[37074]_  & \new_[37071]_ ;
  assign \new_[37076]_  = \new_[37075]_  & \new_[37068]_ ;
  assign \new_[37080]_  = ~A168 & ~A169;
  assign \new_[37081]_  = ~A170 & \new_[37080]_ ;
  assign \new_[37085]_  = A232 & A201;
  assign \new_[37086]_  = A199 & \new_[37085]_ ;
  assign \new_[37087]_  = \new_[37086]_  & \new_[37081]_ ;
  assign \new_[37091]_  = ~A235 & ~A234;
  assign \new_[37092]_  = A233 & \new_[37091]_ ;
  assign \new_[37095]_  = ~A268 & ~A267;
  assign \new_[37098]_  = A301 & ~A269;
  assign \new_[37099]_  = \new_[37098]_  & \new_[37095]_ ;
  assign \new_[37100]_  = \new_[37099]_  & \new_[37092]_ ;
  assign \new_[37104]_  = ~A168 & ~A169;
  assign \new_[37105]_  = ~A170 & \new_[37104]_ ;
  assign \new_[37109]_  = A232 & A201;
  assign \new_[37110]_  = A199 & \new_[37109]_ ;
  assign \new_[37111]_  = \new_[37110]_  & \new_[37105]_ ;
  assign \new_[37115]_  = ~A235 & ~A234;
  assign \new_[37116]_  = A233 & \new_[37115]_ ;
  assign \new_[37119]_  = ~A266 & ~A265;
  assign \new_[37122]_  = A301 & ~A268;
  assign \new_[37123]_  = \new_[37122]_  & \new_[37119]_ ;
  assign \new_[37124]_  = \new_[37123]_  & \new_[37116]_ ;
  assign \new_[37128]_  = ~A168 & ~A169;
  assign \new_[37129]_  = ~A170 & \new_[37128]_ ;
  assign \new_[37133]_  = ~A232 & A201;
  assign \new_[37134]_  = A199 & \new_[37133]_ ;
  assign \new_[37135]_  = \new_[37134]_  & \new_[37129]_ ;
  assign \new_[37139]_  = ~A267 & ~A235;
  assign \new_[37140]_  = ~A233 & \new_[37139]_ ;
  assign \new_[37143]_  = ~A269 & ~A268;
  assign \new_[37146]_  = A300 & A299;
  assign \new_[37147]_  = \new_[37146]_  & \new_[37143]_ ;
  assign \new_[37148]_  = \new_[37147]_  & \new_[37140]_ ;
  assign \new_[37152]_  = ~A168 & ~A169;
  assign \new_[37153]_  = ~A170 & \new_[37152]_ ;
  assign \new_[37157]_  = ~A232 & A201;
  assign \new_[37158]_  = A199 & \new_[37157]_ ;
  assign \new_[37159]_  = \new_[37158]_  & \new_[37153]_ ;
  assign \new_[37163]_  = ~A267 & ~A235;
  assign \new_[37164]_  = ~A233 & \new_[37163]_ ;
  assign \new_[37167]_  = ~A269 & ~A268;
  assign \new_[37170]_  = A300 & A298;
  assign \new_[37171]_  = \new_[37170]_  & \new_[37167]_ ;
  assign \new_[37172]_  = \new_[37171]_  & \new_[37164]_ ;
  assign \new_[37176]_  = ~A168 & ~A169;
  assign \new_[37177]_  = ~A170 & \new_[37176]_ ;
  assign \new_[37181]_  = ~A232 & A201;
  assign \new_[37182]_  = A199 & \new_[37181]_ ;
  assign \new_[37183]_  = \new_[37182]_  & \new_[37177]_ ;
  assign \new_[37187]_  = A265 & ~A235;
  assign \new_[37188]_  = ~A233 & \new_[37187]_ ;
  assign \new_[37191]_  = ~A267 & A266;
  assign \new_[37194]_  = A301 & ~A268;
  assign \new_[37195]_  = \new_[37194]_  & \new_[37191]_ ;
  assign \new_[37196]_  = \new_[37195]_  & \new_[37188]_ ;
  assign \new_[37200]_  = ~A168 & ~A169;
  assign \new_[37201]_  = ~A170 & \new_[37200]_ ;
  assign \new_[37205]_  = ~A232 & A201;
  assign \new_[37206]_  = A199 & \new_[37205]_ ;
  assign \new_[37207]_  = \new_[37206]_  & \new_[37201]_ ;
  assign \new_[37211]_  = ~A265 & ~A235;
  assign \new_[37212]_  = ~A233 & \new_[37211]_ ;
  assign \new_[37215]_  = ~A268 & ~A266;
  assign \new_[37218]_  = A300 & A299;
  assign \new_[37219]_  = \new_[37218]_  & \new_[37215]_ ;
  assign \new_[37220]_  = \new_[37219]_  & \new_[37212]_ ;
  assign \new_[37224]_  = ~A168 & ~A169;
  assign \new_[37225]_  = ~A170 & \new_[37224]_ ;
  assign \new_[37229]_  = ~A232 & A201;
  assign \new_[37230]_  = A199 & \new_[37229]_ ;
  assign \new_[37231]_  = \new_[37230]_  & \new_[37225]_ ;
  assign \new_[37235]_  = ~A265 & ~A235;
  assign \new_[37236]_  = ~A233 & \new_[37235]_ ;
  assign \new_[37239]_  = ~A268 & ~A266;
  assign \new_[37242]_  = A300 & A298;
  assign \new_[37243]_  = \new_[37242]_  & \new_[37239]_ ;
  assign \new_[37244]_  = \new_[37243]_  & \new_[37236]_ ;
  assign \new_[37248]_  = ~A168 & ~A169;
  assign \new_[37249]_  = ~A170 & \new_[37248]_ ;
  assign \new_[37253]_  = ~A234 & A201;
  assign \new_[37254]_  = A200 & \new_[37253]_ ;
  assign \new_[37255]_  = \new_[37254]_  & \new_[37249]_ ;
  assign \new_[37259]_  = ~A267 & ~A236;
  assign \new_[37260]_  = ~A235 & \new_[37259]_ ;
  assign \new_[37263]_  = ~A269 & ~A268;
  assign \new_[37266]_  = A300 & A299;
  assign \new_[37267]_  = \new_[37266]_  & \new_[37263]_ ;
  assign \new_[37268]_  = \new_[37267]_  & \new_[37260]_ ;
  assign \new_[37272]_  = ~A168 & ~A169;
  assign \new_[37273]_  = ~A170 & \new_[37272]_ ;
  assign \new_[37277]_  = ~A234 & A201;
  assign \new_[37278]_  = A200 & \new_[37277]_ ;
  assign \new_[37279]_  = \new_[37278]_  & \new_[37273]_ ;
  assign \new_[37283]_  = ~A267 & ~A236;
  assign \new_[37284]_  = ~A235 & \new_[37283]_ ;
  assign \new_[37287]_  = ~A269 & ~A268;
  assign \new_[37290]_  = A300 & A298;
  assign \new_[37291]_  = \new_[37290]_  & \new_[37287]_ ;
  assign \new_[37292]_  = \new_[37291]_  & \new_[37284]_ ;
  assign \new_[37296]_  = ~A168 & ~A169;
  assign \new_[37297]_  = ~A170 & \new_[37296]_ ;
  assign \new_[37301]_  = ~A234 & A201;
  assign \new_[37302]_  = A200 & \new_[37301]_ ;
  assign \new_[37303]_  = \new_[37302]_  & \new_[37297]_ ;
  assign \new_[37307]_  = A265 & ~A236;
  assign \new_[37308]_  = ~A235 & \new_[37307]_ ;
  assign \new_[37311]_  = ~A267 & A266;
  assign \new_[37314]_  = A301 & ~A268;
  assign \new_[37315]_  = \new_[37314]_  & \new_[37311]_ ;
  assign \new_[37316]_  = \new_[37315]_  & \new_[37308]_ ;
  assign \new_[37320]_  = ~A168 & ~A169;
  assign \new_[37321]_  = ~A170 & \new_[37320]_ ;
  assign \new_[37325]_  = ~A234 & A201;
  assign \new_[37326]_  = A200 & \new_[37325]_ ;
  assign \new_[37327]_  = \new_[37326]_  & \new_[37321]_ ;
  assign \new_[37331]_  = ~A265 & ~A236;
  assign \new_[37332]_  = ~A235 & \new_[37331]_ ;
  assign \new_[37335]_  = ~A268 & ~A266;
  assign \new_[37338]_  = A300 & A299;
  assign \new_[37339]_  = \new_[37338]_  & \new_[37335]_ ;
  assign \new_[37340]_  = \new_[37339]_  & \new_[37332]_ ;
  assign \new_[37344]_  = ~A168 & ~A169;
  assign \new_[37345]_  = ~A170 & \new_[37344]_ ;
  assign \new_[37349]_  = ~A234 & A201;
  assign \new_[37350]_  = A200 & \new_[37349]_ ;
  assign \new_[37351]_  = \new_[37350]_  & \new_[37345]_ ;
  assign \new_[37355]_  = ~A265 & ~A236;
  assign \new_[37356]_  = ~A235 & \new_[37355]_ ;
  assign \new_[37359]_  = ~A268 & ~A266;
  assign \new_[37362]_  = A300 & A298;
  assign \new_[37363]_  = \new_[37362]_  & \new_[37359]_ ;
  assign \new_[37364]_  = \new_[37363]_  & \new_[37356]_ ;
  assign \new_[37368]_  = ~A168 & ~A169;
  assign \new_[37369]_  = ~A170 & \new_[37368]_ ;
  assign \new_[37373]_  = A232 & A201;
  assign \new_[37374]_  = A200 & \new_[37373]_ ;
  assign \new_[37375]_  = \new_[37374]_  & \new_[37369]_ ;
  assign \new_[37379]_  = ~A235 & ~A234;
  assign \new_[37380]_  = A233 & \new_[37379]_ ;
  assign \new_[37383]_  = ~A268 & ~A267;
  assign \new_[37386]_  = A301 & ~A269;
  assign \new_[37387]_  = \new_[37386]_  & \new_[37383]_ ;
  assign \new_[37388]_  = \new_[37387]_  & \new_[37380]_ ;
  assign \new_[37392]_  = ~A168 & ~A169;
  assign \new_[37393]_  = ~A170 & \new_[37392]_ ;
  assign \new_[37397]_  = A232 & A201;
  assign \new_[37398]_  = A200 & \new_[37397]_ ;
  assign \new_[37399]_  = \new_[37398]_  & \new_[37393]_ ;
  assign \new_[37403]_  = ~A235 & ~A234;
  assign \new_[37404]_  = A233 & \new_[37403]_ ;
  assign \new_[37407]_  = ~A266 & ~A265;
  assign \new_[37410]_  = A301 & ~A268;
  assign \new_[37411]_  = \new_[37410]_  & \new_[37407]_ ;
  assign \new_[37412]_  = \new_[37411]_  & \new_[37404]_ ;
  assign \new_[37416]_  = ~A168 & ~A169;
  assign \new_[37417]_  = ~A170 & \new_[37416]_ ;
  assign \new_[37421]_  = ~A232 & A201;
  assign \new_[37422]_  = A200 & \new_[37421]_ ;
  assign \new_[37423]_  = \new_[37422]_  & \new_[37417]_ ;
  assign \new_[37427]_  = ~A267 & ~A235;
  assign \new_[37428]_  = ~A233 & \new_[37427]_ ;
  assign \new_[37431]_  = ~A269 & ~A268;
  assign \new_[37434]_  = A300 & A299;
  assign \new_[37435]_  = \new_[37434]_  & \new_[37431]_ ;
  assign \new_[37436]_  = \new_[37435]_  & \new_[37428]_ ;
  assign \new_[37440]_  = ~A168 & ~A169;
  assign \new_[37441]_  = ~A170 & \new_[37440]_ ;
  assign \new_[37445]_  = ~A232 & A201;
  assign \new_[37446]_  = A200 & \new_[37445]_ ;
  assign \new_[37447]_  = \new_[37446]_  & \new_[37441]_ ;
  assign \new_[37451]_  = ~A267 & ~A235;
  assign \new_[37452]_  = ~A233 & \new_[37451]_ ;
  assign \new_[37455]_  = ~A269 & ~A268;
  assign \new_[37458]_  = A300 & A298;
  assign \new_[37459]_  = \new_[37458]_  & \new_[37455]_ ;
  assign \new_[37460]_  = \new_[37459]_  & \new_[37452]_ ;
  assign \new_[37464]_  = ~A168 & ~A169;
  assign \new_[37465]_  = ~A170 & \new_[37464]_ ;
  assign \new_[37469]_  = ~A232 & A201;
  assign \new_[37470]_  = A200 & \new_[37469]_ ;
  assign \new_[37471]_  = \new_[37470]_  & \new_[37465]_ ;
  assign \new_[37475]_  = A265 & ~A235;
  assign \new_[37476]_  = ~A233 & \new_[37475]_ ;
  assign \new_[37479]_  = ~A267 & A266;
  assign \new_[37482]_  = A301 & ~A268;
  assign \new_[37483]_  = \new_[37482]_  & \new_[37479]_ ;
  assign \new_[37484]_  = \new_[37483]_  & \new_[37476]_ ;
  assign \new_[37488]_  = ~A168 & ~A169;
  assign \new_[37489]_  = ~A170 & \new_[37488]_ ;
  assign \new_[37493]_  = ~A232 & A201;
  assign \new_[37494]_  = A200 & \new_[37493]_ ;
  assign \new_[37495]_  = \new_[37494]_  & \new_[37489]_ ;
  assign \new_[37499]_  = ~A265 & ~A235;
  assign \new_[37500]_  = ~A233 & \new_[37499]_ ;
  assign \new_[37503]_  = ~A268 & ~A266;
  assign \new_[37506]_  = A300 & A299;
  assign \new_[37507]_  = \new_[37506]_  & \new_[37503]_ ;
  assign \new_[37508]_  = \new_[37507]_  & \new_[37500]_ ;
  assign \new_[37512]_  = ~A168 & ~A169;
  assign \new_[37513]_  = ~A170 & \new_[37512]_ ;
  assign \new_[37517]_  = ~A232 & A201;
  assign \new_[37518]_  = A200 & \new_[37517]_ ;
  assign \new_[37519]_  = \new_[37518]_  & \new_[37513]_ ;
  assign \new_[37523]_  = ~A265 & ~A235;
  assign \new_[37524]_  = ~A233 & \new_[37523]_ ;
  assign \new_[37527]_  = ~A268 & ~A266;
  assign \new_[37530]_  = A300 & A298;
  assign \new_[37531]_  = \new_[37530]_  & \new_[37527]_ ;
  assign \new_[37532]_  = \new_[37531]_  & \new_[37524]_ ;
  assign \new_[37536]_  = ~A168 & ~A169;
  assign \new_[37537]_  = ~A170 & \new_[37536]_ ;
  assign \new_[37541]_  = A203 & A200;
  assign \new_[37542]_  = ~A199 & \new_[37541]_ ;
  assign \new_[37543]_  = \new_[37542]_  & \new_[37537]_ ;
  assign \new_[37547]_  = ~A236 & ~A235;
  assign \new_[37548]_  = ~A234 & \new_[37547]_ ;
  assign \new_[37551]_  = ~A268 & ~A267;
  assign \new_[37554]_  = A301 & ~A269;
  assign \new_[37555]_  = \new_[37554]_  & \new_[37551]_ ;
  assign \new_[37556]_  = \new_[37555]_  & \new_[37548]_ ;
  assign \new_[37560]_  = ~A168 & ~A169;
  assign \new_[37561]_  = ~A170 & \new_[37560]_ ;
  assign \new_[37565]_  = A203 & A200;
  assign \new_[37566]_  = ~A199 & \new_[37565]_ ;
  assign \new_[37567]_  = \new_[37566]_  & \new_[37561]_ ;
  assign \new_[37571]_  = ~A236 & ~A235;
  assign \new_[37572]_  = ~A234 & \new_[37571]_ ;
  assign \new_[37575]_  = ~A266 & ~A265;
  assign \new_[37578]_  = A301 & ~A268;
  assign \new_[37579]_  = \new_[37578]_  & \new_[37575]_ ;
  assign \new_[37580]_  = \new_[37579]_  & \new_[37572]_ ;
  assign \new_[37584]_  = ~A168 & ~A169;
  assign \new_[37585]_  = ~A170 & \new_[37584]_ ;
  assign \new_[37589]_  = A203 & A200;
  assign \new_[37590]_  = ~A199 & \new_[37589]_ ;
  assign \new_[37591]_  = \new_[37590]_  & \new_[37585]_ ;
  assign \new_[37595]_  = A236 & A233;
  assign \new_[37596]_  = ~A232 & \new_[37595]_ ;
  assign \new_[37599]_  = A299 & A298;
  assign \new_[37602]_  = ~A301 & ~A300;
  assign \new_[37603]_  = \new_[37602]_  & \new_[37599]_ ;
  assign \new_[37604]_  = \new_[37603]_  & \new_[37596]_ ;
  assign \new_[37608]_  = ~A168 & ~A169;
  assign \new_[37609]_  = ~A170 & \new_[37608]_ ;
  assign \new_[37613]_  = A203 & A200;
  assign \new_[37614]_  = ~A199 & \new_[37613]_ ;
  assign \new_[37615]_  = \new_[37614]_  & \new_[37609]_ ;
  assign \new_[37619]_  = A236 & ~A233;
  assign \new_[37620]_  = A232 & \new_[37619]_ ;
  assign \new_[37623]_  = A299 & A298;
  assign \new_[37626]_  = ~A301 & ~A300;
  assign \new_[37627]_  = \new_[37626]_  & \new_[37623]_ ;
  assign \new_[37628]_  = \new_[37627]_  & \new_[37620]_ ;
  assign \new_[37632]_  = ~A168 & ~A169;
  assign \new_[37633]_  = ~A170 & \new_[37632]_ ;
  assign \new_[37637]_  = A203 & A200;
  assign \new_[37638]_  = ~A199 & \new_[37637]_ ;
  assign \new_[37639]_  = \new_[37638]_  & \new_[37633]_ ;
  assign \new_[37643]_  = ~A235 & ~A233;
  assign \new_[37644]_  = ~A232 & \new_[37643]_ ;
  assign \new_[37647]_  = ~A268 & ~A267;
  assign \new_[37650]_  = A301 & ~A269;
  assign \new_[37651]_  = \new_[37650]_  & \new_[37647]_ ;
  assign \new_[37652]_  = \new_[37651]_  & \new_[37644]_ ;
  assign \new_[37656]_  = ~A168 & ~A169;
  assign \new_[37657]_  = ~A170 & \new_[37656]_ ;
  assign \new_[37661]_  = A203 & A200;
  assign \new_[37662]_  = ~A199 & \new_[37661]_ ;
  assign \new_[37663]_  = \new_[37662]_  & \new_[37657]_ ;
  assign \new_[37667]_  = ~A235 & ~A233;
  assign \new_[37668]_  = ~A232 & \new_[37667]_ ;
  assign \new_[37671]_  = ~A266 & ~A265;
  assign \new_[37674]_  = A301 & ~A268;
  assign \new_[37675]_  = \new_[37674]_  & \new_[37671]_ ;
  assign \new_[37676]_  = \new_[37675]_  & \new_[37668]_ ;
  assign \new_[37680]_  = ~A168 & ~A169;
  assign \new_[37681]_  = ~A170 & \new_[37680]_ ;
  assign \new_[37685]_  = A203 & ~A200;
  assign \new_[37686]_  = A199 & \new_[37685]_ ;
  assign \new_[37687]_  = \new_[37686]_  & \new_[37681]_ ;
  assign \new_[37691]_  = ~A236 & ~A235;
  assign \new_[37692]_  = ~A234 & \new_[37691]_ ;
  assign \new_[37695]_  = ~A268 & ~A267;
  assign \new_[37698]_  = A301 & ~A269;
  assign \new_[37699]_  = \new_[37698]_  & \new_[37695]_ ;
  assign \new_[37700]_  = \new_[37699]_  & \new_[37692]_ ;
  assign \new_[37704]_  = ~A168 & ~A169;
  assign \new_[37705]_  = ~A170 & \new_[37704]_ ;
  assign \new_[37709]_  = A203 & ~A200;
  assign \new_[37710]_  = A199 & \new_[37709]_ ;
  assign \new_[37711]_  = \new_[37710]_  & \new_[37705]_ ;
  assign \new_[37715]_  = ~A236 & ~A235;
  assign \new_[37716]_  = ~A234 & \new_[37715]_ ;
  assign \new_[37719]_  = ~A266 & ~A265;
  assign \new_[37722]_  = A301 & ~A268;
  assign \new_[37723]_  = \new_[37722]_  & \new_[37719]_ ;
  assign \new_[37724]_  = \new_[37723]_  & \new_[37716]_ ;
  assign \new_[37728]_  = ~A168 & ~A169;
  assign \new_[37729]_  = ~A170 & \new_[37728]_ ;
  assign \new_[37733]_  = A203 & ~A200;
  assign \new_[37734]_  = A199 & \new_[37733]_ ;
  assign \new_[37735]_  = \new_[37734]_  & \new_[37729]_ ;
  assign \new_[37739]_  = A236 & A233;
  assign \new_[37740]_  = ~A232 & \new_[37739]_ ;
  assign \new_[37743]_  = A299 & A298;
  assign \new_[37746]_  = ~A301 & ~A300;
  assign \new_[37747]_  = \new_[37746]_  & \new_[37743]_ ;
  assign \new_[37748]_  = \new_[37747]_  & \new_[37740]_ ;
  assign \new_[37752]_  = ~A168 & ~A169;
  assign \new_[37753]_  = ~A170 & \new_[37752]_ ;
  assign \new_[37757]_  = A203 & ~A200;
  assign \new_[37758]_  = A199 & \new_[37757]_ ;
  assign \new_[37759]_  = \new_[37758]_  & \new_[37753]_ ;
  assign \new_[37763]_  = A236 & ~A233;
  assign \new_[37764]_  = A232 & \new_[37763]_ ;
  assign \new_[37767]_  = A299 & A298;
  assign \new_[37770]_  = ~A301 & ~A300;
  assign \new_[37771]_  = \new_[37770]_  & \new_[37767]_ ;
  assign \new_[37772]_  = \new_[37771]_  & \new_[37764]_ ;
  assign \new_[37776]_  = ~A168 & ~A169;
  assign \new_[37777]_  = ~A170 & \new_[37776]_ ;
  assign \new_[37781]_  = A203 & ~A200;
  assign \new_[37782]_  = A199 & \new_[37781]_ ;
  assign \new_[37783]_  = \new_[37782]_  & \new_[37777]_ ;
  assign \new_[37787]_  = ~A235 & ~A233;
  assign \new_[37788]_  = ~A232 & \new_[37787]_ ;
  assign \new_[37791]_  = ~A268 & ~A267;
  assign \new_[37794]_  = A301 & ~A269;
  assign \new_[37795]_  = \new_[37794]_  & \new_[37791]_ ;
  assign \new_[37796]_  = \new_[37795]_  & \new_[37788]_ ;
  assign \new_[37800]_  = ~A168 & ~A169;
  assign \new_[37801]_  = ~A170 & \new_[37800]_ ;
  assign \new_[37805]_  = A203 & ~A200;
  assign \new_[37806]_  = A199 & \new_[37805]_ ;
  assign \new_[37807]_  = \new_[37806]_  & \new_[37801]_ ;
  assign \new_[37811]_  = ~A235 & ~A233;
  assign \new_[37812]_  = ~A232 & \new_[37811]_ ;
  assign \new_[37815]_  = ~A266 & ~A265;
  assign \new_[37818]_  = A301 & ~A268;
  assign \new_[37819]_  = \new_[37818]_  & \new_[37815]_ ;
  assign \new_[37820]_  = \new_[37819]_  & \new_[37812]_ ;
  assign \new_[37824]_  = ~A201 & A166;
  assign \new_[37825]_  = A168 & \new_[37824]_ ;
  assign \new_[37828]_  = ~A203 & ~A202;
  assign \new_[37831]_  = ~A235 & ~A234;
  assign \new_[37832]_  = \new_[37831]_  & \new_[37828]_ ;
  assign \new_[37833]_  = \new_[37832]_  & \new_[37825]_ ;
  assign \new_[37837]_  = ~A268 & ~A267;
  assign \new_[37838]_  = ~A236 & \new_[37837]_ ;
  assign \new_[37841]_  = A298 & ~A269;
  assign \new_[37844]_  = A302 & ~A299;
  assign \new_[37845]_  = \new_[37844]_  & \new_[37841]_ ;
  assign \new_[37846]_  = \new_[37845]_  & \new_[37838]_ ;
  assign \new_[37850]_  = ~A201 & A166;
  assign \new_[37851]_  = A168 & \new_[37850]_ ;
  assign \new_[37854]_  = ~A203 & ~A202;
  assign \new_[37857]_  = ~A235 & ~A234;
  assign \new_[37858]_  = \new_[37857]_  & \new_[37854]_ ;
  assign \new_[37859]_  = \new_[37858]_  & \new_[37851]_ ;
  assign \new_[37863]_  = ~A268 & ~A267;
  assign \new_[37864]_  = ~A236 & \new_[37863]_ ;
  assign \new_[37867]_  = ~A298 & ~A269;
  assign \new_[37870]_  = A302 & A299;
  assign \new_[37871]_  = \new_[37870]_  & \new_[37867]_ ;
  assign \new_[37872]_  = \new_[37871]_  & \new_[37864]_ ;
  assign \new_[37876]_  = ~A201 & A166;
  assign \new_[37877]_  = A168 & \new_[37876]_ ;
  assign \new_[37880]_  = ~A203 & ~A202;
  assign \new_[37883]_  = ~A235 & ~A234;
  assign \new_[37884]_  = \new_[37883]_  & \new_[37880]_ ;
  assign \new_[37885]_  = \new_[37884]_  & \new_[37877]_ ;
  assign \new_[37889]_  = A266 & A265;
  assign \new_[37890]_  = ~A236 & \new_[37889]_ ;
  assign \new_[37893]_  = ~A268 & ~A267;
  assign \new_[37896]_  = A300 & A299;
  assign \new_[37897]_  = \new_[37896]_  & \new_[37893]_ ;
  assign \new_[37898]_  = \new_[37897]_  & \new_[37890]_ ;
  assign \new_[37902]_  = ~A201 & A166;
  assign \new_[37903]_  = A168 & \new_[37902]_ ;
  assign \new_[37906]_  = ~A203 & ~A202;
  assign \new_[37909]_  = ~A235 & ~A234;
  assign \new_[37910]_  = \new_[37909]_  & \new_[37906]_ ;
  assign \new_[37911]_  = \new_[37910]_  & \new_[37903]_ ;
  assign \new_[37915]_  = A266 & A265;
  assign \new_[37916]_  = ~A236 & \new_[37915]_ ;
  assign \new_[37919]_  = ~A268 & ~A267;
  assign \new_[37922]_  = A300 & A298;
  assign \new_[37923]_  = \new_[37922]_  & \new_[37919]_ ;
  assign \new_[37924]_  = \new_[37923]_  & \new_[37916]_ ;
  assign \new_[37928]_  = ~A201 & A166;
  assign \new_[37929]_  = A168 & \new_[37928]_ ;
  assign \new_[37932]_  = ~A203 & ~A202;
  assign \new_[37935]_  = ~A235 & ~A234;
  assign \new_[37936]_  = \new_[37935]_  & \new_[37932]_ ;
  assign \new_[37937]_  = \new_[37936]_  & \new_[37929]_ ;
  assign \new_[37941]_  = ~A266 & ~A265;
  assign \new_[37942]_  = ~A236 & \new_[37941]_ ;
  assign \new_[37945]_  = A298 & ~A268;
  assign \new_[37948]_  = A302 & ~A299;
  assign \new_[37949]_  = \new_[37948]_  & \new_[37945]_ ;
  assign \new_[37950]_  = \new_[37949]_  & \new_[37942]_ ;
  assign \new_[37954]_  = ~A201 & A166;
  assign \new_[37955]_  = A168 & \new_[37954]_ ;
  assign \new_[37958]_  = ~A203 & ~A202;
  assign \new_[37961]_  = ~A235 & ~A234;
  assign \new_[37962]_  = \new_[37961]_  & \new_[37958]_ ;
  assign \new_[37963]_  = \new_[37962]_  & \new_[37955]_ ;
  assign \new_[37967]_  = ~A266 & ~A265;
  assign \new_[37968]_  = ~A236 & \new_[37967]_ ;
  assign \new_[37971]_  = ~A298 & ~A268;
  assign \new_[37974]_  = A302 & A299;
  assign \new_[37975]_  = \new_[37974]_  & \new_[37971]_ ;
  assign \new_[37976]_  = \new_[37975]_  & \new_[37968]_ ;
  assign \new_[37980]_  = ~A201 & A166;
  assign \new_[37981]_  = A168 & \new_[37980]_ ;
  assign \new_[37984]_  = ~A203 & ~A202;
  assign \new_[37987]_  = A233 & A232;
  assign \new_[37988]_  = \new_[37987]_  & \new_[37984]_ ;
  assign \new_[37989]_  = \new_[37988]_  & \new_[37981]_ ;
  assign \new_[37993]_  = ~A267 & ~A235;
  assign \new_[37994]_  = ~A234 & \new_[37993]_ ;
  assign \new_[37997]_  = ~A269 & ~A268;
  assign \new_[38000]_  = A300 & A299;
  assign \new_[38001]_  = \new_[38000]_  & \new_[37997]_ ;
  assign \new_[38002]_  = \new_[38001]_  & \new_[37994]_ ;
  assign \new_[38006]_  = ~A201 & A166;
  assign \new_[38007]_  = A168 & \new_[38006]_ ;
  assign \new_[38010]_  = ~A203 & ~A202;
  assign \new_[38013]_  = A233 & A232;
  assign \new_[38014]_  = \new_[38013]_  & \new_[38010]_ ;
  assign \new_[38015]_  = \new_[38014]_  & \new_[38007]_ ;
  assign \new_[38019]_  = ~A267 & ~A235;
  assign \new_[38020]_  = ~A234 & \new_[38019]_ ;
  assign \new_[38023]_  = ~A269 & ~A268;
  assign \new_[38026]_  = A300 & A298;
  assign \new_[38027]_  = \new_[38026]_  & \new_[38023]_ ;
  assign \new_[38028]_  = \new_[38027]_  & \new_[38020]_ ;
  assign \new_[38032]_  = ~A201 & A166;
  assign \new_[38033]_  = A168 & \new_[38032]_ ;
  assign \new_[38036]_  = ~A203 & ~A202;
  assign \new_[38039]_  = A233 & A232;
  assign \new_[38040]_  = \new_[38039]_  & \new_[38036]_ ;
  assign \new_[38041]_  = \new_[38040]_  & \new_[38033]_ ;
  assign \new_[38045]_  = A265 & ~A235;
  assign \new_[38046]_  = ~A234 & \new_[38045]_ ;
  assign \new_[38049]_  = ~A267 & A266;
  assign \new_[38052]_  = A301 & ~A268;
  assign \new_[38053]_  = \new_[38052]_  & \new_[38049]_ ;
  assign \new_[38054]_  = \new_[38053]_  & \new_[38046]_ ;
  assign \new_[38058]_  = ~A201 & A166;
  assign \new_[38059]_  = A168 & \new_[38058]_ ;
  assign \new_[38062]_  = ~A203 & ~A202;
  assign \new_[38065]_  = A233 & A232;
  assign \new_[38066]_  = \new_[38065]_  & \new_[38062]_ ;
  assign \new_[38067]_  = \new_[38066]_  & \new_[38059]_ ;
  assign \new_[38071]_  = ~A265 & ~A235;
  assign \new_[38072]_  = ~A234 & \new_[38071]_ ;
  assign \new_[38075]_  = ~A268 & ~A266;
  assign \new_[38078]_  = A300 & A299;
  assign \new_[38079]_  = \new_[38078]_  & \new_[38075]_ ;
  assign \new_[38080]_  = \new_[38079]_  & \new_[38072]_ ;
  assign \new_[38084]_  = ~A201 & A166;
  assign \new_[38085]_  = A168 & \new_[38084]_ ;
  assign \new_[38088]_  = ~A203 & ~A202;
  assign \new_[38091]_  = A233 & A232;
  assign \new_[38092]_  = \new_[38091]_  & \new_[38088]_ ;
  assign \new_[38093]_  = \new_[38092]_  & \new_[38085]_ ;
  assign \new_[38097]_  = ~A265 & ~A235;
  assign \new_[38098]_  = ~A234 & \new_[38097]_ ;
  assign \new_[38101]_  = ~A268 & ~A266;
  assign \new_[38104]_  = A300 & A298;
  assign \new_[38105]_  = \new_[38104]_  & \new_[38101]_ ;
  assign \new_[38106]_  = \new_[38105]_  & \new_[38098]_ ;
  assign \new_[38110]_  = ~A201 & A166;
  assign \new_[38111]_  = A168 & \new_[38110]_ ;
  assign \new_[38114]_  = ~A203 & ~A202;
  assign \new_[38117]_  = ~A233 & ~A232;
  assign \new_[38118]_  = \new_[38117]_  & \new_[38114]_ ;
  assign \new_[38119]_  = \new_[38118]_  & \new_[38111]_ ;
  assign \new_[38123]_  = ~A268 & ~A267;
  assign \new_[38124]_  = ~A235 & \new_[38123]_ ;
  assign \new_[38127]_  = A298 & ~A269;
  assign \new_[38130]_  = A302 & ~A299;
  assign \new_[38131]_  = \new_[38130]_  & \new_[38127]_ ;
  assign \new_[38132]_  = \new_[38131]_  & \new_[38124]_ ;
  assign \new_[38136]_  = ~A201 & A166;
  assign \new_[38137]_  = A168 & \new_[38136]_ ;
  assign \new_[38140]_  = ~A203 & ~A202;
  assign \new_[38143]_  = ~A233 & ~A232;
  assign \new_[38144]_  = \new_[38143]_  & \new_[38140]_ ;
  assign \new_[38145]_  = \new_[38144]_  & \new_[38137]_ ;
  assign \new_[38149]_  = ~A268 & ~A267;
  assign \new_[38150]_  = ~A235 & \new_[38149]_ ;
  assign \new_[38153]_  = ~A298 & ~A269;
  assign \new_[38156]_  = A302 & A299;
  assign \new_[38157]_  = \new_[38156]_  & \new_[38153]_ ;
  assign \new_[38158]_  = \new_[38157]_  & \new_[38150]_ ;
  assign \new_[38162]_  = ~A201 & A166;
  assign \new_[38163]_  = A168 & \new_[38162]_ ;
  assign \new_[38166]_  = ~A203 & ~A202;
  assign \new_[38169]_  = ~A233 & ~A232;
  assign \new_[38170]_  = \new_[38169]_  & \new_[38166]_ ;
  assign \new_[38171]_  = \new_[38170]_  & \new_[38163]_ ;
  assign \new_[38175]_  = A266 & A265;
  assign \new_[38176]_  = ~A235 & \new_[38175]_ ;
  assign \new_[38179]_  = ~A268 & ~A267;
  assign \new_[38182]_  = A300 & A299;
  assign \new_[38183]_  = \new_[38182]_  & \new_[38179]_ ;
  assign \new_[38184]_  = \new_[38183]_  & \new_[38176]_ ;
  assign \new_[38188]_  = ~A201 & A166;
  assign \new_[38189]_  = A168 & \new_[38188]_ ;
  assign \new_[38192]_  = ~A203 & ~A202;
  assign \new_[38195]_  = ~A233 & ~A232;
  assign \new_[38196]_  = \new_[38195]_  & \new_[38192]_ ;
  assign \new_[38197]_  = \new_[38196]_  & \new_[38189]_ ;
  assign \new_[38201]_  = A266 & A265;
  assign \new_[38202]_  = ~A235 & \new_[38201]_ ;
  assign \new_[38205]_  = ~A268 & ~A267;
  assign \new_[38208]_  = A300 & A298;
  assign \new_[38209]_  = \new_[38208]_  & \new_[38205]_ ;
  assign \new_[38210]_  = \new_[38209]_  & \new_[38202]_ ;
  assign \new_[38214]_  = ~A201 & A166;
  assign \new_[38215]_  = A168 & \new_[38214]_ ;
  assign \new_[38218]_  = ~A203 & ~A202;
  assign \new_[38221]_  = ~A233 & ~A232;
  assign \new_[38222]_  = \new_[38221]_  & \new_[38218]_ ;
  assign \new_[38223]_  = \new_[38222]_  & \new_[38215]_ ;
  assign \new_[38227]_  = ~A266 & ~A265;
  assign \new_[38228]_  = ~A235 & \new_[38227]_ ;
  assign \new_[38231]_  = A298 & ~A268;
  assign \new_[38234]_  = A302 & ~A299;
  assign \new_[38235]_  = \new_[38234]_  & \new_[38231]_ ;
  assign \new_[38236]_  = \new_[38235]_  & \new_[38228]_ ;
  assign \new_[38240]_  = ~A201 & A166;
  assign \new_[38241]_  = A168 & \new_[38240]_ ;
  assign \new_[38244]_  = ~A203 & ~A202;
  assign \new_[38247]_  = ~A233 & ~A232;
  assign \new_[38248]_  = \new_[38247]_  & \new_[38244]_ ;
  assign \new_[38249]_  = \new_[38248]_  & \new_[38241]_ ;
  assign \new_[38253]_  = ~A266 & ~A265;
  assign \new_[38254]_  = ~A235 & \new_[38253]_ ;
  assign \new_[38257]_  = ~A298 & ~A268;
  assign \new_[38260]_  = A302 & A299;
  assign \new_[38261]_  = \new_[38260]_  & \new_[38257]_ ;
  assign \new_[38262]_  = \new_[38261]_  & \new_[38254]_ ;
  assign \new_[38266]_  = A199 & A166;
  assign \new_[38267]_  = A168 & \new_[38266]_ ;
  assign \new_[38270]_  = ~A201 & A200;
  assign \new_[38273]_  = ~A234 & ~A202;
  assign \new_[38274]_  = \new_[38273]_  & \new_[38270]_ ;
  assign \new_[38275]_  = \new_[38274]_  & \new_[38267]_ ;
  assign \new_[38279]_  = ~A267 & ~A236;
  assign \new_[38280]_  = ~A235 & \new_[38279]_ ;
  assign \new_[38283]_  = ~A269 & ~A268;
  assign \new_[38286]_  = A300 & A299;
  assign \new_[38287]_  = \new_[38286]_  & \new_[38283]_ ;
  assign \new_[38288]_  = \new_[38287]_  & \new_[38280]_ ;
  assign \new_[38292]_  = A199 & A166;
  assign \new_[38293]_  = A168 & \new_[38292]_ ;
  assign \new_[38296]_  = ~A201 & A200;
  assign \new_[38299]_  = ~A234 & ~A202;
  assign \new_[38300]_  = \new_[38299]_  & \new_[38296]_ ;
  assign \new_[38301]_  = \new_[38300]_  & \new_[38293]_ ;
  assign \new_[38305]_  = ~A267 & ~A236;
  assign \new_[38306]_  = ~A235 & \new_[38305]_ ;
  assign \new_[38309]_  = ~A269 & ~A268;
  assign \new_[38312]_  = A300 & A298;
  assign \new_[38313]_  = \new_[38312]_  & \new_[38309]_ ;
  assign \new_[38314]_  = \new_[38313]_  & \new_[38306]_ ;
  assign \new_[38318]_  = A199 & A166;
  assign \new_[38319]_  = A168 & \new_[38318]_ ;
  assign \new_[38322]_  = ~A201 & A200;
  assign \new_[38325]_  = ~A234 & ~A202;
  assign \new_[38326]_  = \new_[38325]_  & \new_[38322]_ ;
  assign \new_[38327]_  = \new_[38326]_  & \new_[38319]_ ;
  assign \new_[38331]_  = A265 & ~A236;
  assign \new_[38332]_  = ~A235 & \new_[38331]_ ;
  assign \new_[38335]_  = ~A267 & A266;
  assign \new_[38338]_  = A301 & ~A268;
  assign \new_[38339]_  = \new_[38338]_  & \new_[38335]_ ;
  assign \new_[38340]_  = \new_[38339]_  & \new_[38332]_ ;
  assign \new_[38344]_  = A199 & A166;
  assign \new_[38345]_  = A168 & \new_[38344]_ ;
  assign \new_[38348]_  = ~A201 & A200;
  assign \new_[38351]_  = ~A234 & ~A202;
  assign \new_[38352]_  = \new_[38351]_  & \new_[38348]_ ;
  assign \new_[38353]_  = \new_[38352]_  & \new_[38345]_ ;
  assign \new_[38357]_  = ~A265 & ~A236;
  assign \new_[38358]_  = ~A235 & \new_[38357]_ ;
  assign \new_[38361]_  = ~A268 & ~A266;
  assign \new_[38364]_  = A300 & A299;
  assign \new_[38365]_  = \new_[38364]_  & \new_[38361]_ ;
  assign \new_[38366]_  = \new_[38365]_  & \new_[38358]_ ;
  assign \new_[38370]_  = A199 & A166;
  assign \new_[38371]_  = A168 & \new_[38370]_ ;
  assign \new_[38374]_  = ~A201 & A200;
  assign \new_[38377]_  = ~A234 & ~A202;
  assign \new_[38378]_  = \new_[38377]_  & \new_[38374]_ ;
  assign \new_[38379]_  = \new_[38378]_  & \new_[38371]_ ;
  assign \new_[38383]_  = ~A265 & ~A236;
  assign \new_[38384]_  = ~A235 & \new_[38383]_ ;
  assign \new_[38387]_  = ~A268 & ~A266;
  assign \new_[38390]_  = A300 & A298;
  assign \new_[38391]_  = \new_[38390]_  & \new_[38387]_ ;
  assign \new_[38392]_  = \new_[38391]_  & \new_[38384]_ ;
  assign \new_[38396]_  = A199 & A166;
  assign \new_[38397]_  = A168 & \new_[38396]_ ;
  assign \new_[38400]_  = ~A201 & A200;
  assign \new_[38403]_  = A232 & ~A202;
  assign \new_[38404]_  = \new_[38403]_  & \new_[38400]_ ;
  assign \new_[38405]_  = \new_[38404]_  & \new_[38397]_ ;
  assign \new_[38409]_  = ~A235 & ~A234;
  assign \new_[38410]_  = A233 & \new_[38409]_ ;
  assign \new_[38413]_  = ~A268 & ~A267;
  assign \new_[38416]_  = A301 & ~A269;
  assign \new_[38417]_  = \new_[38416]_  & \new_[38413]_ ;
  assign \new_[38418]_  = \new_[38417]_  & \new_[38410]_ ;
  assign \new_[38422]_  = A199 & A166;
  assign \new_[38423]_  = A168 & \new_[38422]_ ;
  assign \new_[38426]_  = ~A201 & A200;
  assign \new_[38429]_  = A232 & ~A202;
  assign \new_[38430]_  = \new_[38429]_  & \new_[38426]_ ;
  assign \new_[38431]_  = \new_[38430]_  & \new_[38423]_ ;
  assign \new_[38435]_  = ~A235 & ~A234;
  assign \new_[38436]_  = A233 & \new_[38435]_ ;
  assign \new_[38439]_  = ~A266 & ~A265;
  assign \new_[38442]_  = A301 & ~A268;
  assign \new_[38443]_  = \new_[38442]_  & \new_[38439]_ ;
  assign \new_[38444]_  = \new_[38443]_  & \new_[38436]_ ;
  assign \new_[38448]_  = A199 & A166;
  assign \new_[38449]_  = A168 & \new_[38448]_ ;
  assign \new_[38452]_  = ~A201 & A200;
  assign \new_[38455]_  = ~A232 & ~A202;
  assign \new_[38456]_  = \new_[38455]_  & \new_[38452]_ ;
  assign \new_[38457]_  = \new_[38456]_  & \new_[38449]_ ;
  assign \new_[38461]_  = ~A267 & ~A235;
  assign \new_[38462]_  = ~A233 & \new_[38461]_ ;
  assign \new_[38465]_  = ~A269 & ~A268;
  assign \new_[38468]_  = A300 & A299;
  assign \new_[38469]_  = \new_[38468]_  & \new_[38465]_ ;
  assign \new_[38470]_  = \new_[38469]_  & \new_[38462]_ ;
  assign \new_[38474]_  = A199 & A166;
  assign \new_[38475]_  = A168 & \new_[38474]_ ;
  assign \new_[38478]_  = ~A201 & A200;
  assign \new_[38481]_  = ~A232 & ~A202;
  assign \new_[38482]_  = \new_[38481]_  & \new_[38478]_ ;
  assign \new_[38483]_  = \new_[38482]_  & \new_[38475]_ ;
  assign \new_[38487]_  = ~A267 & ~A235;
  assign \new_[38488]_  = ~A233 & \new_[38487]_ ;
  assign \new_[38491]_  = ~A269 & ~A268;
  assign \new_[38494]_  = A300 & A298;
  assign \new_[38495]_  = \new_[38494]_  & \new_[38491]_ ;
  assign \new_[38496]_  = \new_[38495]_  & \new_[38488]_ ;
  assign \new_[38500]_  = A199 & A166;
  assign \new_[38501]_  = A168 & \new_[38500]_ ;
  assign \new_[38504]_  = ~A201 & A200;
  assign \new_[38507]_  = ~A232 & ~A202;
  assign \new_[38508]_  = \new_[38507]_  & \new_[38504]_ ;
  assign \new_[38509]_  = \new_[38508]_  & \new_[38501]_ ;
  assign \new_[38513]_  = A265 & ~A235;
  assign \new_[38514]_  = ~A233 & \new_[38513]_ ;
  assign \new_[38517]_  = ~A267 & A266;
  assign \new_[38520]_  = A301 & ~A268;
  assign \new_[38521]_  = \new_[38520]_  & \new_[38517]_ ;
  assign \new_[38522]_  = \new_[38521]_  & \new_[38514]_ ;
  assign \new_[38526]_  = A199 & A166;
  assign \new_[38527]_  = A168 & \new_[38526]_ ;
  assign \new_[38530]_  = ~A201 & A200;
  assign \new_[38533]_  = ~A232 & ~A202;
  assign \new_[38534]_  = \new_[38533]_  & \new_[38530]_ ;
  assign \new_[38535]_  = \new_[38534]_  & \new_[38527]_ ;
  assign \new_[38539]_  = ~A265 & ~A235;
  assign \new_[38540]_  = ~A233 & \new_[38539]_ ;
  assign \new_[38543]_  = ~A268 & ~A266;
  assign \new_[38546]_  = A300 & A299;
  assign \new_[38547]_  = \new_[38546]_  & \new_[38543]_ ;
  assign \new_[38548]_  = \new_[38547]_  & \new_[38540]_ ;
  assign \new_[38552]_  = A199 & A166;
  assign \new_[38553]_  = A168 & \new_[38552]_ ;
  assign \new_[38556]_  = ~A201 & A200;
  assign \new_[38559]_  = ~A232 & ~A202;
  assign \new_[38560]_  = \new_[38559]_  & \new_[38556]_ ;
  assign \new_[38561]_  = \new_[38560]_  & \new_[38553]_ ;
  assign \new_[38565]_  = ~A265 & ~A235;
  assign \new_[38566]_  = ~A233 & \new_[38565]_ ;
  assign \new_[38569]_  = ~A268 & ~A266;
  assign \new_[38572]_  = A300 & A298;
  assign \new_[38573]_  = \new_[38572]_  & \new_[38569]_ ;
  assign \new_[38574]_  = \new_[38573]_  & \new_[38566]_ ;
  assign \new_[38578]_  = ~A199 & A166;
  assign \new_[38579]_  = A168 & \new_[38578]_ ;
  assign \new_[38582]_  = ~A202 & ~A200;
  assign \new_[38585]_  = ~A235 & ~A234;
  assign \new_[38586]_  = \new_[38585]_  & \new_[38582]_ ;
  assign \new_[38587]_  = \new_[38586]_  & \new_[38579]_ ;
  assign \new_[38591]_  = ~A268 & ~A267;
  assign \new_[38592]_  = ~A236 & \new_[38591]_ ;
  assign \new_[38595]_  = A298 & ~A269;
  assign \new_[38598]_  = A302 & ~A299;
  assign \new_[38599]_  = \new_[38598]_  & \new_[38595]_ ;
  assign \new_[38600]_  = \new_[38599]_  & \new_[38592]_ ;
  assign \new_[38604]_  = ~A199 & A166;
  assign \new_[38605]_  = A168 & \new_[38604]_ ;
  assign \new_[38608]_  = ~A202 & ~A200;
  assign \new_[38611]_  = ~A235 & ~A234;
  assign \new_[38612]_  = \new_[38611]_  & \new_[38608]_ ;
  assign \new_[38613]_  = \new_[38612]_  & \new_[38605]_ ;
  assign \new_[38617]_  = ~A268 & ~A267;
  assign \new_[38618]_  = ~A236 & \new_[38617]_ ;
  assign \new_[38621]_  = ~A298 & ~A269;
  assign \new_[38624]_  = A302 & A299;
  assign \new_[38625]_  = \new_[38624]_  & \new_[38621]_ ;
  assign \new_[38626]_  = \new_[38625]_  & \new_[38618]_ ;
  assign \new_[38630]_  = ~A199 & A166;
  assign \new_[38631]_  = A168 & \new_[38630]_ ;
  assign \new_[38634]_  = ~A202 & ~A200;
  assign \new_[38637]_  = ~A235 & ~A234;
  assign \new_[38638]_  = \new_[38637]_  & \new_[38634]_ ;
  assign \new_[38639]_  = \new_[38638]_  & \new_[38631]_ ;
  assign \new_[38643]_  = A266 & A265;
  assign \new_[38644]_  = ~A236 & \new_[38643]_ ;
  assign \new_[38647]_  = ~A268 & ~A267;
  assign \new_[38650]_  = A300 & A299;
  assign \new_[38651]_  = \new_[38650]_  & \new_[38647]_ ;
  assign \new_[38652]_  = \new_[38651]_  & \new_[38644]_ ;
  assign \new_[38656]_  = ~A199 & A166;
  assign \new_[38657]_  = A168 & \new_[38656]_ ;
  assign \new_[38660]_  = ~A202 & ~A200;
  assign \new_[38663]_  = ~A235 & ~A234;
  assign \new_[38664]_  = \new_[38663]_  & \new_[38660]_ ;
  assign \new_[38665]_  = \new_[38664]_  & \new_[38657]_ ;
  assign \new_[38669]_  = A266 & A265;
  assign \new_[38670]_  = ~A236 & \new_[38669]_ ;
  assign \new_[38673]_  = ~A268 & ~A267;
  assign \new_[38676]_  = A300 & A298;
  assign \new_[38677]_  = \new_[38676]_  & \new_[38673]_ ;
  assign \new_[38678]_  = \new_[38677]_  & \new_[38670]_ ;
  assign \new_[38682]_  = ~A199 & A166;
  assign \new_[38683]_  = A168 & \new_[38682]_ ;
  assign \new_[38686]_  = ~A202 & ~A200;
  assign \new_[38689]_  = ~A235 & ~A234;
  assign \new_[38690]_  = \new_[38689]_  & \new_[38686]_ ;
  assign \new_[38691]_  = \new_[38690]_  & \new_[38683]_ ;
  assign \new_[38695]_  = ~A266 & ~A265;
  assign \new_[38696]_  = ~A236 & \new_[38695]_ ;
  assign \new_[38699]_  = A298 & ~A268;
  assign \new_[38702]_  = A302 & ~A299;
  assign \new_[38703]_  = \new_[38702]_  & \new_[38699]_ ;
  assign \new_[38704]_  = \new_[38703]_  & \new_[38696]_ ;
  assign \new_[38708]_  = ~A199 & A166;
  assign \new_[38709]_  = A168 & \new_[38708]_ ;
  assign \new_[38712]_  = ~A202 & ~A200;
  assign \new_[38715]_  = ~A235 & ~A234;
  assign \new_[38716]_  = \new_[38715]_  & \new_[38712]_ ;
  assign \new_[38717]_  = \new_[38716]_  & \new_[38709]_ ;
  assign \new_[38721]_  = ~A266 & ~A265;
  assign \new_[38722]_  = ~A236 & \new_[38721]_ ;
  assign \new_[38725]_  = ~A298 & ~A268;
  assign \new_[38728]_  = A302 & A299;
  assign \new_[38729]_  = \new_[38728]_  & \new_[38725]_ ;
  assign \new_[38730]_  = \new_[38729]_  & \new_[38722]_ ;
  assign \new_[38734]_  = ~A199 & A166;
  assign \new_[38735]_  = A168 & \new_[38734]_ ;
  assign \new_[38738]_  = ~A202 & ~A200;
  assign \new_[38741]_  = A233 & A232;
  assign \new_[38742]_  = \new_[38741]_  & \new_[38738]_ ;
  assign \new_[38743]_  = \new_[38742]_  & \new_[38735]_ ;
  assign \new_[38747]_  = ~A267 & ~A235;
  assign \new_[38748]_  = ~A234 & \new_[38747]_ ;
  assign \new_[38751]_  = ~A269 & ~A268;
  assign \new_[38754]_  = A300 & A299;
  assign \new_[38755]_  = \new_[38754]_  & \new_[38751]_ ;
  assign \new_[38756]_  = \new_[38755]_  & \new_[38748]_ ;
  assign \new_[38760]_  = ~A199 & A166;
  assign \new_[38761]_  = A168 & \new_[38760]_ ;
  assign \new_[38764]_  = ~A202 & ~A200;
  assign \new_[38767]_  = A233 & A232;
  assign \new_[38768]_  = \new_[38767]_  & \new_[38764]_ ;
  assign \new_[38769]_  = \new_[38768]_  & \new_[38761]_ ;
  assign \new_[38773]_  = ~A267 & ~A235;
  assign \new_[38774]_  = ~A234 & \new_[38773]_ ;
  assign \new_[38777]_  = ~A269 & ~A268;
  assign \new_[38780]_  = A300 & A298;
  assign \new_[38781]_  = \new_[38780]_  & \new_[38777]_ ;
  assign \new_[38782]_  = \new_[38781]_  & \new_[38774]_ ;
  assign \new_[38786]_  = ~A199 & A166;
  assign \new_[38787]_  = A168 & \new_[38786]_ ;
  assign \new_[38790]_  = ~A202 & ~A200;
  assign \new_[38793]_  = A233 & A232;
  assign \new_[38794]_  = \new_[38793]_  & \new_[38790]_ ;
  assign \new_[38795]_  = \new_[38794]_  & \new_[38787]_ ;
  assign \new_[38799]_  = A265 & ~A235;
  assign \new_[38800]_  = ~A234 & \new_[38799]_ ;
  assign \new_[38803]_  = ~A267 & A266;
  assign \new_[38806]_  = A301 & ~A268;
  assign \new_[38807]_  = \new_[38806]_  & \new_[38803]_ ;
  assign \new_[38808]_  = \new_[38807]_  & \new_[38800]_ ;
  assign \new_[38812]_  = ~A199 & A166;
  assign \new_[38813]_  = A168 & \new_[38812]_ ;
  assign \new_[38816]_  = ~A202 & ~A200;
  assign \new_[38819]_  = A233 & A232;
  assign \new_[38820]_  = \new_[38819]_  & \new_[38816]_ ;
  assign \new_[38821]_  = \new_[38820]_  & \new_[38813]_ ;
  assign \new_[38825]_  = ~A265 & ~A235;
  assign \new_[38826]_  = ~A234 & \new_[38825]_ ;
  assign \new_[38829]_  = ~A268 & ~A266;
  assign \new_[38832]_  = A300 & A299;
  assign \new_[38833]_  = \new_[38832]_  & \new_[38829]_ ;
  assign \new_[38834]_  = \new_[38833]_  & \new_[38826]_ ;
  assign \new_[38838]_  = ~A199 & A166;
  assign \new_[38839]_  = A168 & \new_[38838]_ ;
  assign \new_[38842]_  = ~A202 & ~A200;
  assign \new_[38845]_  = A233 & A232;
  assign \new_[38846]_  = \new_[38845]_  & \new_[38842]_ ;
  assign \new_[38847]_  = \new_[38846]_  & \new_[38839]_ ;
  assign \new_[38851]_  = ~A265 & ~A235;
  assign \new_[38852]_  = ~A234 & \new_[38851]_ ;
  assign \new_[38855]_  = ~A268 & ~A266;
  assign \new_[38858]_  = A300 & A298;
  assign \new_[38859]_  = \new_[38858]_  & \new_[38855]_ ;
  assign \new_[38860]_  = \new_[38859]_  & \new_[38852]_ ;
  assign \new_[38864]_  = ~A199 & A166;
  assign \new_[38865]_  = A168 & \new_[38864]_ ;
  assign \new_[38868]_  = ~A202 & ~A200;
  assign \new_[38871]_  = ~A233 & ~A232;
  assign \new_[38872]_  = \new_[38871]_  & \new_[38868]_ ;
  assign \new_[38873]_  = \new_[38872]_  & \new_[38865]_ ;
  assign \new_[38877]_  = ~A268 & ~A267;
  assign \new_[38878]_  = ~A235 & \new_[38877]_ ;
  assign \new_[38881]_  = A298 & ~A269;
  assign \new_[38884]_  = A302 & ~A299;
  assign \new_[38885]_  = \new_[38884]_  & \new_[38881]_ ;
  assign \new_[38886]_  = \new_[38885]_  & \new_[38878]_ ;
  assign \new_[38890]_  = ~A199 & A166;
  assign \new_[38891]_  = A168 & \new_[38890]_ ;
  assign \new_[38894]_  = ~A202 & ~A200;
  assign \new_[38897]_  = ~A233 & ~A232;
  assign \new_[38898]_  = \new_[38897]_  & \new_[38894]_ ;
  assign \new_[38899]_  = \new_[38898]_  & \new_[38891]_ ;
  assign \new_[38903]_  = ~A268 & ~A267;
  assign \new_[38904]_  = ~A235 & \new_[38903]_ ;
  assign \new_[38907]_  = ~A298 & ~A269;
  assign \new_[38910]_  = A302 & A299;
  assign \new_[38911]_  = \new_[38910]_  & \new_[38907]_ ;
  assign \new_[38912]_  = \new_[38911]_  & \new_[38904]_ ;
  assign \new_[38916]_  = ~A199 & A166;
  assign \new_[38917]_  = A168 & \new_[38916]_ ;
  assign \new_[38920]_  = ~A202 & ~A200;
  assign \new_[38923]_  = ~A233 & ~A232;
  assign \new_[38924]_  = \new_[38923]_  & \new_[38920]_ ;
  assign \new_[38925]_  = \new_[38924]_  & \new_[38917]_ ;
  assign \new_[38929]_  = A266 & A265;
  assign \new_[38930]_  = ~A235 & \new_[38929]_ ;
  assign \new_[38933]_  = ~A268 & ~A267;
  assign \new_[38936]_  = A300 & A299;
  assign \new_[38937]_  = \new_[38936]_  & \new_[38933]_ ;
  assign \new_[38938]_  = \new_[38937]_  & \new_[38930]_ ;
  assign \new_[38942]_  = ~A199 & A166;
  assign \new_[38943]_  = A168 & \new_[38942]_ ;
  assign \new_[38946]_  = ~A202 & ~A200;
  assign \new_[38949]_  = ~A233 & ~A232;
  assign \new_[38950]_  = \new_[38949]_  & \new_[38946]_ ;
  assign \new_[38951]_  = \new_[38950]_  & \new_[38943]_ ;
  assign \new_[38955]_  = A266 & A265;
  assign \new_[38956]_  = ~A235 & \new_[38955]_ ;
  assign \new_[38959]_  = ~A268 & ~A267;
  assign \new_[38962]_  = A300 & A298;
  assign \new_[38963]_  = \new_[38962]_  & \new_[38959]_ ;
  assign \new_[38964]_  = \new_[38963]_  & \new_[38956]_ ;
  assign \new_[38968]_  = ~A199 & A166;
  assign \new_[38969]_  = A168 & \new_[38968]_ ;
  assign \new_[38972]_  = ~A202 & ~A200;
  assign \new_[38975]_  = ~A233 & ~A232;
  assign \new_[38976]_  = \new_[38975]_  & \new_[38972]_ ;
  assign \new_[38977]_  = \new_[38976]_  & \new_[38969]_ ;
  assign \new_[38981]_  = ~A266 & ~A265;
  assign \new_[38982]_  = ~A235 & \new_[38981]_ ;
  assign \new_[38985]_  = A298 & ~A268;
  assign \new_[38988]_  = A302 & ~A299;
  assign \new_[38989]_  = \new_[38988]_  & \new_[38985]_ ;
  assign \new_[38990]_  = \new_[38989]_  & \new_[38982]_ ;
  assign \new_[38994]_  = ~A199 & A166;
  assign \new_[38995]_  = A168 & \new_[38994]_ ;
  assign \new_[38998]_  = ~A202 & ~A200;
  assign \new_[39001]_  = ~A233 & ~A232;
  assign \new_[39002]_  = \new_[39001]_  & \new_[38998]_ ;
  assign \new_[39003]_  = \new_[39002]_  & \new_[38995]_ ;
  assign \new_[39007]_  = ~A266 & ~A265;
  assign \new_[39008]_  = ~A235 & \new_[39007]_ ;
  assign \new_[39011]_  = ~A298 & ~A268;
  assign \new_[39014]_  = A302 & A299;
  assign \new_[39015]_  = \new_[39014]_  & \new_[39011]_ ;
  assign \new_[39016]_  = \new_[39015]_  & \new_[39008]_ ;
  assign \new_[39020]_  = ~A201 & A167;
  assign \new_[39021]_  = A168 & \new_[39020]_ ;
  assign \new_[39024]_  = ~A203 & ~A202;
  assign \new_[39027]_  = ~A235 & ~A234;
  assign \new_[39028]_  = \new_[39027]_  & \new_[39024]_ ;
  assign \new_[39029]_  = \new_[39028]_  & \new_[39021]_ ;
  assign \new_[39033]_  = ~A268 & ~A267;
  assign \new_[39034]_  = ~A236 & \new_[39033]_ ;
  assign \new_[39037]_  = A298 & ~A269;
  assign \new_[39040]_  = A302 & ~A299;
  assign \new_[39041]_  = \new_[39040]_  & \new_[39037]_ ;
  assign \new_[39042]_  = \new_[39041]_  & \new_[39034]_ ;
  assign \new_[39046]_  = ~A201 & A167;
  assign \new_[39047]_  = A168 & \new_[39046]_ ;
  assign \new_[39050]_  = ~A203 & ~A202;
  assign \new_[39053]_  = ~A235 & ~A234;
  assign \new_[39054]_  = \new_[39053]_  & \new_[39050]_ ;
  assign \new_[39055]_  = \new_[39054]_  & \new_[39047]_ ;
  assign \new_[39059]_  = ~A268 & ~A267;
  assign \new_[39060]_  = ~A236 & \new_[39059]_ ;
  assign \new_[39063]_  = ~A298 & ~A269;
  assign \new_[39066]_  = A302 & A299;
  assign \new_[39067]_  = \new_[39066]_  & \new_[39063]_ ;
  assign \new_[39068]_  = \new_[39067]_  & \new_[39060]_ ;
  assign \new_[39072]_  = ~A201 & A167;
  assign \new_[39073]_  = A168 & \new_[39072]_ ;
  assign \new_[39076]_  = ~A203 & ~A202;
  assign \new_[39079]_  = ~A235 & ~A234;
  assign \new_[39080]_  = \new_[39079]_  & \new_[39076]_ ;
  assign \new_[39081]_  = \new_[39080]_  & \new_[39073]_ ;
  assign \new_[39085]_  = A266 & A265;
  assign \new_[39086]_  = ~A236 & \new_[39085]_ ;
  assign \new_[39089]_  = ~A268 & ~A267;
  assign \new_[39092]_  = A300 & A299;
  assign \new_[39093]_  = \new_[39092]_  & \new_[39089]_ ;
  assign \new_[39094]_  = \new_[39093]_  & \new_[39086]_ ;
  assign \new_[39098]_  = ~A201 & A167;
  assign \new_[39099]_  = A168 & \new_[39098]_ ;
  assign \new_[39102]_  = ~A203 & ~A202;
  assign \new_[39105]_  = ~A235 & ~A234;
  assign \new_[39106]_  = \new_[39105]_  & \new_[39102]_ ;
  assign \new_[39107]_  = \new_[39106]_  & \new_[39099]_ ;
  assign \new_[39111]_  = A266 & A265;
  assign \new_[39112]_  = ~A236 & \new_[39111]_ ;
  assign \new_[39115]_  = ~A268 & ~A267;
  assign \new_[39118]_  = A300 & A298;
  assign \new_[39119]_  = \new_[39118]_  & \new_[39115]_ ;
  assign \new_[39120]_  = \new_[39119]_  & \new_[39112]_ ;
  assign \new_[39124]_  = ~A201 & A167;
  assign \new_[39125]_  = A168 & \new_[39124]_ ;
  assign \new_[39128]_  = ~A203 & ~A202;
  assign \new_[39131]_  = ~A235 & ~A234;
  assign \new_[39132]_  = \new_[39131]_  & \new_[39128]_ ;
  assign \new_[39133]_  = \new_[39132]_  & \new_[39125]_ ;
  assign \new_[39137]_  = ~A266 & ~A265;
  assign \new_[39138]_  = ~A236 & \new_[39137]_ ;
  assign \new_[39141]_  = A298 & ~A268;
  assign \new_[39144]_  = A302 & ~A299;
  assign \new_[39145]_  = \new_[39144]_  & \new_[39141]_ ;
  assign \new_[39146]_  = \new_[39145]_  & \new_[39138]_ ;
  assign \new_[39150]_  = ~A201 & A167;
  assign \new_[39151]_  = A168 & \new_[39150]_ ;
  assign \new_[39154]_  = ~A203 & ~A202;
  assign \new_[39157]_  = ~A235 & ~A234;
  assign \new_[39158]_  = \new_[39157]_  & \new_[39154]_ ;
  assign \new_[39159]_  = \new_[39158]_  & \new_[39151]_ ;
  assign \new_[39163]_  = ~A266 & ~A265;
  assign \new_[39164]_  = ~A236 & \new_[39163]_ ;
  assign \new_[39167]_  = ~A298 & ~A268;
  assign \new_[39170]_  = A302 & A299;
  assign \new_[39171]_  = \new_[39170]_  & \new_[39167]_ ;
  assign \new_[39172]_  = \new_[39171]_  & \new_[39164]_ ;
  assign \new_[39176]_  = ~A201 & A167;
  assign \new_[39177]_  = A168 & \new_[39176]_ ;
  assign \new_[39180]_  = ~A203 & ~A202;
  assign \new_[39183]_  = A233 & A232;
  assign \new_[39184]_  = \new_[39183]_  & \new_[39180]_ ;
  assign \new_[39185]_  = \new_[39184]_  & \new_[39177]_ ;
  assign \new_[39189]_  = ~A267 & ~A235;
  assign \new_[39190]_  = ~A234 & \new_[39189]_ ;
  assign \new_[39193]_  = ~A269 & ~A268;
  assign \new_[39196]_  = A300 & A299;
  assign \new_[39197]_  = \new_[39196]_  & \new_[39193]_ ;
  assign \new_[39198]_  = \new_[39197]_  & \new_[39190]_ ;
  assign \new_[39202]_  = ~A201 & A167;
  assign \new_[39203]_  = A168 & \new_[39202]_ ;
  assign \new_[39206]_  = ~A203 & ~A202;
  assign \new_[39209]_  = A233 & A232;
  assign \new_[39210]_  = \new_[39209]_  & \new_[39206]_ ;
  assign \new_[39211]_  = \new_[39210]_  & \new_[39203]_ ;
  assign \new_[39215]_  = ~A267 & ~A235;
  assign \new_[39216]_  = ~A234 & \new_[39215]_ ;
  assign \new_[39219]_  = ~A269 & ~A268;
  assign \new_[39222]_  = A300 & A298;
  assign \new_[39223]_  = \new_[39222]_  & \new_[39219]_ ;
  assign \new_[39224]_  = \new_[39223]_  & \new_[39216]_ ;
  assign \new_[39228]_  = ~A201 & A167;
  assign \new_[39229]_  = A168 & \new_[39228]_ ;
  assign \new_[39232]_  = ~A203 & ~A202;
  assign \new_[39235]_  = A233 & A232;
  assign \new_[39236]_  = \new_[39235]_  & \new_[39232]_ ;
  assign \new_[39237]_  = \new_[39236]_  & \new_[39229]_ ;
  assign \new_[39241]_  = A265 & ~A235;
  assign \new_[39242]_  = ~A234 & \new_[39241]_ ;
  assign \new_[39245]_  = ~A267 & A266;
  assign \new_[39248]_  = A301 & ~A268;
  assign \new_[39249]_  = \new_[39248]_  & \new_[39245]_ ;
  assign \new_[39250]_  = \new_[39249]_  & \new_[39242]_ ;
  assign \new_[39254]_  = ~A201 & A167;
  assign \new_[39255]_  = A168 & \new_[39254]_ ;
  assign \new_[39258]_  = ~A203 & ~A202;
  assign \new_[39261]_  = A233 & A232;
  assign \new_[39262]_  = \new_[39261]_  & \new_[39258]_ ;
  assign \new_[39263]_  = \new_[39262]_  & \new_[39255]_ ;
  assign \new_[39267]_  = ~A265 & ~A235;
  assign \new_[39268]_  = ~A234 & \new_[39267]_ ;
  assign \new_[39271]_  = ~A268 & ~A266;
  assign \new_[39274]_  = A300 & A299;
  assign \new_[39275]_  = \new_[39274]_  & \new_[39271]_ ;
  assign \new_[39276]_  = \new_[39275]_  & \new_[39268]_ ;
  assign \new_[39280]_  = ~A201 & A167;
  assign \new_[39281]_  = A168 & \new_[39280]_ ;
  assign \new_[39284]_  = ~A203 & ~A202;
  assign \new_[39287]_  = A233 & A232;
  assign \new_[39288]_  = \new_[39287]_  & \new_[39284]_ ;
  assign \new_[39289]_  = \new_[39288]_  & \new_[39281]_ ;
  assign \new_[39293]_  = ~A265 & ~A235;
  assign \new_[39294]_  = ~A234 & \new_[39293]_ ;
  assign \new_[39297]_  = ~A268 & ~A266;
  assign \new_[39300]_  = A300 & A298;
  assign \new_[39301]_  = \new_[39300]_  & \new_[39297]_ ;
  assign \new_[39302]_  = \new_[39301]_  & \new_[39294]_ ;
  assign \new_[39306]_  = ~A201 & A167;
  assign \new_[39307]_  = A168 & \new_[39306]_ ;
  assign \new_[39310]_  = ~A203 & ~A202;
  assign \new_[39313]_  = ~A233 & ~A232;
  assign \new_[39314]_  = \new_[39313]_  & \new_[39310]_ ;
  assign \new_[39315]_  = \new_[39314]_  & \new_[39307]_ ;
  assign \new_[39319]_  = ~A268 & ~A267;
  assign \new_[39320]_  = ~A235 & \new_[39319]_ ;
  assign \new_[39323]_  = A298 & ~A269;
  assign \new_[39326]_  = A302 & ~A299;
  assign \new_[39327]_  = \new_[39326]_  & \new_[39323]_ ;
  assign \new_[39328]_  = \new_[39327]_  & \new_[39320]_ ;
  assign \new_[39332]_  = ~A201 & A167;
  assign \new_[39333]_  = A168 & \new_[39332]_ ;
  assign \new_[39336]_  = ~A203 & ~A202;
  assign \new_[39339]_  = ~A233 & ~A232;
  assign \new_[39340]_  = \new_[39339]_  & \new_[39336]_ ;
  assign \new_[39341]_  = \new_[39340]_  & \new_[39333]_ ;
  assign \new_[39345]_  = ~A268 & ~A267;
  assign \new_[39346]_  = ~A235 & \new_[39345]_ ;
  assign \new_[39349]_  = ~A298 & ~A269;
  assign \new_[39352]_  = A302 & A299;
  assign \new_[39353]_  = \new_[39352]_  & \new_[39349]_ ;
  assign \new_[39354]_  = \new_[39353]_  & \new_[39346]_ ;
  assign \new_[39358]_  = ~A201 & A167;
  assign \new_[39359]_  = A168 & \new_[39358]_ ;
  assign \new_[39362]_  = ~A203 & ~A202;
  assign \new_[39365]_  = ~A233 & ~A232;
  assign \new_[39366]_  = \new_[39365]_  & \new_[39362]_ ;
  assign \new_[39367]_  = \new_[39366]_  & \new_[39359]_ ;
  assign \new_[39371]_  = A266 & A265;
  assign \new_[39372]_  = ~A235 & \new_[39371]_ ;
  assign \new_[39375]_  = ~A268 & ~A267;
  assign \new_[39378]_  = A300 & A299;
  assign \new_[39379]_  = \new_[39378]_  & \new_[39375]_ ;
  assign \new_[39380]_  = \new_[39379]_  & \new_[39372]_ ;
  assign \new_[39384]_  = ~A201 & A167;
  assign \new_[39385]_  = A168 & \new_[39384]_ ;
  assign \new_[39388]_  = ~A203 & ~A202;
  assign \new_[39391]_  = ~A233 & ~A232;
  assign \new_[39392]_  = \new_[39391]_  & \new_[39388]_ ;
  assign \new_[39393]_  = \new_[39392]_  & \new_[39385]_ ;
  assign \new_[39397]_  = A266 & A265;
  assign \new_[39398]_  = ~A235 & \new_[39397]_ ;
  assign \new_[39401]_  = ~A268 & ~A267;
  assign \new_[39404]_  = A300 & A298;
  assign \new_[39405]_  = \new_[39404]_  & \new_[39401]_ ;
  assign \new_[39406]_  = \new_[39405]_  & \new_[39398]_ ;
  assign \new_[39410]_  = ~A201 & A167;
  assign \new_[39411]_  = A168 & \new_[39410]_ ;
  assign \new_[39414]_  = ~A203 & ~A202;
  assign \new_[39417]_  = ~A233 & ~A232;
  assign \new_[39418]_  = \new_[39417]_  & \new_[39414]_ ;
  assign \new_[39419]_  = \new_[39418]_  & \new_[39411]_ ;
  assign \new_[39423]_  = ~A266 & ~A265;
  assign \new_[39424]_  = ~A235 & \new_[39423]_ ;
  assign \new_[39427]_  = A298 & ~A268;
  assign \new_[39430]_  = A302 & ~A299;
  assign \new_[39431]_  = \new_[39430]_  & \new_[39427]_ ;
  assign \new_[39432]_  = \new_[39431]_  & \new_[39424]_ ;
  assign \new_[39436]_  = ~A201 & A167;
  assign \new_[39437]_  = A168 & \new_[39436]_ ;
  assign \new_[39440]_  = ~A203 & ~A202;
  assign \new_[39443]_  = ~A233 & ~A232;
  assign \new_[39444]_  = \new_[39443]_  & \new_[39440]_ ;
  assign \new_[39445]_  = \new_[39444]_  & \new_[39437]_ ;
  assign \new_[39449]_  = ~A266 & ~A265;
  assign \new_[39450]_  = ~A235 & \new_[39449]_ ;
  assign \new_[39453]_  = ~A298 & ~A268;
  assign \new_[39456]_  = A302 & A299;
  assign \new_[39457]_  = \new_[39456]_  & \new_[39453]_ ;
  assign \new_[39458]_  = \new_[39457]_  & \new_[39450]_ ;
  assign \new_[39462]_  = A199 & A167;
  assign \new_[39463]_  = A168 & \new_[39462]_ ;
  assign \new_[39466]_  = ~A201 & A200;
  assign \new_[39469]_  = ~A234 & ~A202;
  assign \new_[39470]_  = \new_[39469]_  & \new_[39466]_ ;
  assign \new_[39471]_  = \new_[39470]_  & \new_[39463]_ ;
  assign \new_[39475]_  = ~A267 & ~A236;
  assign \new_[39476]_  = ~A235 & \new_[39475]_ ;
  assign \new_[39479]_  = ~A269 & ~A268;
  assign \new_[39482]_  = A300 & A299;
  assign \new_[39483]_  = \new_[39482]_  & \new_[39479]_ ;
  assign \new_[39484]_  = \new_[39483]_  & \new_[39476]_ ;
  assign \new_[39488]_  = A199 & A167;
  assign \new_[39489]_  = A168 & \new_[39488]_ ;
  assign \new_[39492]_  = ~A201 & A200;
  assign \new_[39495]_  = ~A234 & ~A202;
  assign \new_[39496]_  = \new_[39495]_  & \new_[39492]_ ;
  assign \new_[39497]_  = \new_[39496]_  & \new_[39489]_ ;
  assign \new_[39501]_  = ~A267 & ~A236;
  assign \new_[39502]_  = ~A235 & \new_[39501]_ ;
  assign \new_[39505]_  = ~A269 & ~A268;
  assign \new_[39508]_  = A300 & A298;
  assign \new_[39509]_  = \new_[39508]_  & \new_[39505]_ ;
  assign \new_[39510]_  = \new_[39509]_  & \new_[39502]_ ;
  assign \new_[39514]_  = A199 & A167;
  assign \new_[39515]_  = A168 & \new_[39514]_ ;
  assign \new_[39518]_  = ~A201 & A200;
  assign \new_[39521]_  = ~A234 & ~A202;
  assign \new_[39522]_  = \new_[39521]_  & \new_[39518]_ ;
  assign \new_[39523]_  = \new_[39522]_  & \new_[39515]_ ;
  assign \new_[39527]_  = A265 & ~A236;
  assign \new_[39528]_  = ~A235 & \new_[39527]_ ;
  assign \new_[39531]_  = ~A267 & A266;
  assign \new_[39534]_  = A301 & ~A268;
  assign \new_[39535]_  = \new_[39534]_  & \new_[39531]_ ;
  assign \new_[39536]_  = \new_[39535]_  & \new_[39528]_ ;
  assign \new_[39540]_  = A199 & A167;
  assign \new_[39541]_  = A168 & \new_[39540]_ ;
  assign \new_[39544]_  = ~A201 & A200;
  assign \new_[39547]_  = ~A234 & ~A202;
  assign \new_[39548]_  = \new_[39547]_  & \new_[39544]_ ;
  assign \new_[39549]_  = \new_[39548]_  & \new_[39541]_ ;
  assign \new_[39553]_  = ~A265 & ~A236;
  assign \new_[39554]_  = ~A235 & \new_[39553]_ ;
  assign \new_[39557]_  = ~A268 & ~A266;
  assign \new_[39560]_  = A300 & A299;
  assign \new_[39561]_  = \new_[39560]_  & \new_[39557]_ ;
  assign \new_[39562]_  = \new_[39561]_  & \new_[39554]_ ;
  assign \new_[39566]_  = A199 & A167;
  assign \new_[39567]_  = A168 & \new_[39566]_ ;
  assign \new_[39570]_  = ~A201 & A200;
  assign \new_[39573]_  = ~A234 & ~A202;
  assign \new_[39574]_  = \new_[39573]_  & \new_[39570]_ ;
  assign \new_[39575]_  = \new_[39574]_  & \new_[39567]_ ;
  assign \new_[39579]_  = ~A265 & ~A236;
  assign \new_[39580]_  = ~A235 & \new_[39579]_ ;
  assign \new_[39583]_  = ~A268 & ~A266;
  assign \new_[39586]_  = A300 & A298;
  assign \new_[39587]_  = \new_[39586]_  & \new_[39583]_ ;
  assign \new_[39588]_  = \new_[39587]_  & \new_[39580]_ ;
  assign \new_[39592]_  = A199 & A167;
  assign \new_[39593]_  = A168 & \new_[39592]_ ;
  assign \new_[39596]_  = ~A201 & A200;
  assign \new_[39599]_  = A232 & ~A202;
  assign \new_[39600]_  = \new_[39599]_  & \new_[39596]_ ;
  assign \new_[39601]_  = \new_[39600]_  & \new_[39593]_ ;
  assign \new_[39605]_  = ~A235 & ~A234;
  assign \new_[39606]_  = A233 & \new_[39605]_ ;
  assign \new_[39609]_  = ~A268 & ~A267;
  assign \new_[39612]_  = A301 & ~A269;
  assign \new_[39613]_  = \new_[39612]_  & \new_[39609]_ ;
  assign \new_[39614]_  = \new_[39613]_  & \new_[39606]_ ;
  assign \new_[39618]_  = A199 & A167;
  assign \new_[39619]_  = A168 & \new_[39618]_ ;
  assign \new_[39622]_  = ~A201 & A200;
  assign \new_[39625]_  = A232 & ~A202;
  assign \new_[39626]_  = \new_[39625]_  & \new_[39622]_ ;
  assign \new_[39627]_  = \new_[39626]_  & \new_[39619]_ ;
  assign \new_[39631]_  = ~A235 & ~A234;
  assign \new_[39632]_  = A233 & \new_[39631]_ ;
  assign \new_[39635]_  = ~A266 & ~A265;
  assign \new_[39638]_  = A301 & ~A268;
  assign \new_[39639]_  = \new_[39638]_  & \new_[39635]_ ;
  assign \new_[39640]_  = \new_[39639]_  & \new_[39632]_ ;
  assign \new_[39644]_  = A199 & A167;
  assign \new_[39645]_  = A168 & \new_[39644]_ ;
  assign \new_[39648]_  = ~A201 & A200;
  assign \new_[39651]_  = ~A232 & ~A202;
  assign \new_[39652]_  = \new_[39651]_  & \new_[39648]_ ;
  assign \new_[39653]_  = \new_[39652]_  & \new_[39645]_ ;
  assign \new_[39657]_  = ~A267 & ~A235;
  assign \new_[39658]_  = ~A233 & \new_[39657]_ ;
  assign \new_[39661]_  = ~A269 & ~A268;
  assign \new_[39664]_  = A300 & A299;
  assign \new_[39665]_  = \new_[39664]_  & \new_[39661]_ ;
  assign \new_[39666]_  = \new_[39665]_  & \new_[39658]_ ;
  assign \new_[39670]_  = A199 & A167;
  assign \new_[39671]_  = A168 & \new_[39670]_ ;
  assign \new_[39674]_  = ~A201 & A200;
  assign \new_[39677]_  = ~A232 & ~A202;
  assign \new_[39678]_  = \new_[39677]_  & \new_[39674]_ ;
  assign \new_[39679]_  = \new_[39678]_  & \new_[39671]_ ;
  assign \new_[39683]_  = ~A267 & ~A235;
  assign \new_[39684]_  = ~A233 & \new_[39683]_ ;
  assign \new_[39687]_  = ~A269 & ~A268;
  assign \new_[39690]_  = A300 & A298;
  assign \new_[39691]_  = \new_[39690]_  & \new_[39687]_ ;
  assign \new_[39692]_  = \new_[39691]_  & \new_[39684]_ ;
  assign \new_[39696]_  = A199 & A167;
  assign \new_[39697]_  = A168 & \new_[39696]_ ;
  assign \new_[39700]_  = ~A201 & A200;
  assign \new_[39703]_  = ~A232 & ~A202;
  assign \new_[39704]_  = \new_[39703]_  & \new_[39700]_ ;
  assign \new_[39705]_  = \new_[39704]_  & \new_[39697]_ ;
  assign \new_[39709]_  = A265 & ~A235;
  assign \new_[39710]_  = ~A233 & \new_[39709]_ ;
  assign \new_[39713]_  = ~A267 & A266;
  assign \new_[39716]_  = A301 & ~A268;
  assign \new_[39717]_  = \new_[39716]_  & \new_[39713]_ ;
  assign \new_[39718]_  = \new_[39717]_  & \new_[39710]_ ;
  assign \new_[39722]_  = A199 & A167;
  assign \new_[39723]_  = A168 & \new_[39722]_ ;
  assign \new_[39726]_  = ~A201 & A200;
  assign \new_[39729]_  = ~A232 & ~A202;
  assign \new_[39730]_  = \new_[39729]_  & \new_[39726]_ ;
  assign \new_[39731]_  = \new_[39730]_  & \new_[39723]_ ;
  assign \new_[39735]_  = ~A265 & ~A235;
  assign \new_[39736]_  = ~A233 & \new_[39735]_ ;
  assign \new_[39739]_  = ~A268 & ~A266;
  assign \new_[39742]_  = A300 & A299;
  assign \new_[39743]_  = \new_[39742]_  & \new_[39739]_ ;
  assign \new_[39744]_  = \new_[39743]_  & \new_[39736]_ ;
  assign \new_[39748]_  = A199 & A167;
  assign \new_[39749]_  = A168 & \new_[39748]_ ;
  assign \new_[39752]_  = ~A201 & A200;
  assign \new_[39755]_  = ~A232 & ~A202;
  assign \new_[39756]_  = \new_[39755]_  & \new_[39752]_ ;
  assign \new_[39757]_  = \new_[39756]_  & \new_[39749]_ ;
  assign \new_[39761]_  = ~A265 & ~A235;
  assign \new_[39762]_  = ~A233 & \new_[39761]_ ;
  assign \new_[39765]_  = ~A268 & ~A266;
  assign \new_[39768]_  = A300 & A298;
  assign \new_[39769]_  = \new_[39768]_  & \new_[39765]_ ;
  assign \new_[39770]_  = \new_[39769]_  & \new_[39762]_ ;
  assign \new_[39774]_  = ~A199 & A167;
  assign \new_[39775]_  = A168 & \new_[39774]_ ;
  assign \new_[39778]_  = ~A202 & ~A200;
  assign \new_[39781]_  = ~A235 & ~A234;
  assign \new_[39782]_  = \new_[39781]_  & \new_[39778]_ ;
  assign \new_[39783]_  = \new_[39782]_  & \new_[39775]_ ;
  assign \new_[39787]_  = ~A268 & ~A267;
  assign \new_[39788]_  = ~A236 & \new_[39787]_ ;
  assign \new_[39791]_  = A298 & ~A269;
  assign \new_[39794]_  = A302 & ~A299;
  assign \new_[39795]_  = \new_[39794]_  & \new_[39791]_ ;
  assign \new_[39796]_  = \new_[39795]_  & \new_[39788]_ ;
  assign \new_[39800]_  = ~A199 & A167;
  assign \new_[39801]_  = A168 & \new_[39800]_ ;
  assign \new_[39804]_  = ~A202 & ~A200;
  assign \new_[39807]_  = ~A235 & ~A234;
  assign \new_[39808]_  = \new_[39807]_  & \new_[39804]_ ;
  assign \new_[39809]_  = \new_[39808]_  & \new_[39801]_ ;
  assign \new_[39813]_  = ~A268 & ~A267;
  assign \new_[39814]_  = ~A236 & \new_[39813]_ ;
  assign \new_[39817]_  = ~A298 & ~A269;
  assign \new_[39820]_  = A302 & A299;
  assign \new_[39821]_  = \new_[39820]_  & \new_[39817]_ ;
  assign \new_[39822]_  = \new_[39821]_  & \new_[39814]_ ;
  assign \new_[39826]_  = ~A199 & A167;
  assign \new_[39827]_  = A168 & \new_[39826]_ ;
  assign \new_[39830]_  = ~A202 & ~A200;
  assign \new_[39833]_  = ~A235 & ~A234;
  assign \new_[39834]_  = \new_[39833]_  & \new_[39830]_ ;
  assign \new_[39835]_  = \new_[39834]_  & \new_[39827]_ ;
  assign \new_[39839]_  = A266 & A265;
  assign \new_[39840]_  = ~A236 & \new_[39839]_ ;
  assign \new_[39843]_  = ~A268 & ~A267;
  assign \new_[39846]_  = A300 & A299;
  assign \new_[39847]_  = \new_[39846]_  & \new_[39843]_ ;
  assign \new_[39848]_  = \new_[39847]_  & \new_[39840]_ ;
  assign \new_[39852]_  = ~A199 & A167;
  assign \new_[39853]_  = A168 & \new_[39852]_ ;
  assign \new_[39856]_  = ~A202 & ~A200;
  assign \new_[39859]_  = ~A235 & ~A234;
  assign \new_[39860]_  = \new_[39859]_  & \new_[39856]_ ;
  assign \new_[39861]_  = \new_[39860]_  & \new_[39853]_ ;
  assign \new_[39865]_  = A266 & A265;
  assign \new_[39866]_  = ~A236 & \new_[39865]_ ;
  assign \new_[39869]_  = ~A268 & ~A267;
  assign \new_[39872]_  = A300 & A298;
  assign \new_[39873]_  = \new_[39872]_  & \new_[39869]_ ;
  assign \new_[39874]_  = \new_[39873]_  & \new_[39866]_ ;
  assign \new_[39878]_  = ~A199 & A167;
  assign \new_[39879]_  = A168 & \new_[39878]_ ;
  assign \new_[39882]_  = ~A202 & ~A200;
  assign \new_[39885]_  = ~A235 & ~A234;
  assign \new_[39886]_  = \new_[39885]_  & \new_[39882]_ ;
  assign \new_[39887]_  = \new_[39886]_  & \new_[39879]_ ;
  assign \new_[39891]_  = ~A266 & ~A265;
  assign \new_[39892]_  = ~A236 & \new_[39891]_ ;
  assign \new_[39895]_  = A298 & ~A268;
  assign \new_[39898]_  = A302 & ~A299;
  assign \new_[39899]_  = \new_[39898]_  & \new_[39895]_ ;
  assign \new_[39900]_  = \new_[39899]_  & \new_[39892]_ ;
  assign \new_[39904]_  = ~A199 & A167;
  assign \new_[39905]_  = A168 & \new_[39904]_ ;
  assign \new_[39908]_  = ~A202 & ~A200;
  assign \new_[39911]_  = ~A235 & ~A234;
  assign \new_[39912]_  = \new_[39911]_  & \new_[39908]_ ;
  assign \new_[39913]_  = \new_[39912]_  & \new_[39905]_ ;
  assign \new_[39917]_  = ~A266 & ~A265;
  assign \new_[39918]_  = ~A236 & \new_[39917]_ ;
  assign \new_[39921]_  = ~A298 & ~A268;
  assign \new_[39924]_  = A302 & A299;
  assign \new_[39925]_  = \new_[39924]_  & \new_[39921]_ ;
  assign \new_[39926]_  = \new_[39925]_  & \new_[39918]_ ;
  assign \new_[39930]_  = ~A199 & A167;
  assign \new_[39931]_  = A168 & \new_[39930]_ ;
  assign \new_[39934]_  = ~A202 & ~A200;
  assign \new_[39937]_  = A233 & A232;
  assign \new_[39938]_  = \new_[39937]_  & \new_[39934]_ ;
  assign \new_[39939]_  = \new_[39938]_  & \new_[39931]_ ;
  assign \new_[39943]_  = ~A267 & ~A235;
  assign \new_[39944]_  = ~A234 & \new_[39943]_ ;
  assign \new_[39947]_  = ~A269 & ~A268;
  assign \new_[39950]_  = A300 & A299;
  assign \new_[39951]_  = \new_[39950]_  & \new_[39947]_ ;
  assign \new_[39952]_  = \new_[39951]_  & \new_[39944]_ ;
  assign \new_[39956]_  = ~A199 & A167;
  assign \new_[39957]_  = A168 & \new_[39956]_ ;
  assign \new_[39960]_  = ~A202 & ~A200;
  assign \new_[39963]_  = A233 & A232;
  assign \new_[39964]_  = \new_[39963]_  & \new_[39960]_ ;
  assign \new_[39965]_  = \new_[39964]_  & \new_[39957]_ ;
  assign \new_[39969]_  = ~A267 & ~A235;
  assign \new_[39970]_  = ~A234 & \new_[39969]_ ;
  assign \new_[39973]_  = ~A269 & ~A268;
  assign \new_[39976]_  = A300 & A298;
  assign \new_[39977]_  = \new_[39976]_  & \new_[39973]_ ;
  assign \new_[39978]_  = \new_[39977]_  & \new_[39970]_ ;
  assign \new_[39982]_  = ~A199 & A167;
  assign \new_[39983]_  = A168 & \new_[39982]_ ;
  assign \new_[39986]_  = ~A202 & ~A200;
  assign \new_[39989]_  = A233 & A232;
  assign \new_[39990]_  = \new_[39989]_  & \new_[39986]_ ;
  assign \new_[39991]_  = \new_[39990]_  & \new_[39983]_ ;
  assign \new_[39995]_  = A265 & ~A235;
  assign \new_[39996]_  = ~A234 & \new_[39995]_ ;
  assign \new_[39999]_  = ~A267 & A266;
  assign \new_[40002]_  = A301 & ~A268;
  assign \new_[40003]_  = \new_[40002]_  & \new_[39999]_ ;
  assign \new_[40004]_  = \new_[40003]_  & \new_[39996]_ ;
  assign \new_[40008]_  = ~A199 & A167;
  assign \new_[40009]_  = A168 & \new_[40008]_ ;
  assign \new_[40012]_  = ~A202 & ~A200;
  assign \new_[40015]_  = A233 & A232;
  assign \new_[40016]_  = \new_[40015]_  & \new_[40012]_ ;
  assign \new_[40017]_  = \new_[40016]_  & \new_[40009]_ ;
  assign \new_[40021]_  = ~A265 & ~A235;
  assign \new_[40022]_  = ~A234 & \new_[40021]_ ;
  assign \new_[40025]_  = ~A268 & ~A266;
  assign \new_[40028]_  = A300 & A299;
  assign \new_[40029]_  = \new_[40028]_  & \new_[40025]_ ;
  assign \new_[40030]_  = \new_[40029]_  & \new_[40022]_ ;
  assign \new_[40034]_  = ~A199 & A167;
  assign \new_[40035]_  = A168 & \new_[40034]_ ;
  assign \new_[40038]_  = ~A202 & ~A200;
  assign \new_[40041]_  = A233 & A232;
  assign \new_[40042]_  = \new_[40041]_  & \new_[40038]_ ;
  assign \new_[40043]_  = \new_[40042]_  & \new_[40035]_ ;
  assign \new_[40047]_  = ~A265 & ~A235;
  assign \new_[40048]_  = ~A234 & \new_[40047]_ ;
  assign \new_[40051]_  = ~A268 & ~A266;
  assign \new_[40054]_  = A300 & A298;
  assign \new_[40055]_  = \new_[40054]_  & \new_[40051]_ ;
  assign \new_[40056]_  = \new_[40055]_  & \new_[40048]_ ;
  assign \new_[40060]_  = ~A199 & A167;
  assign \new_[40061]_  = A168 & \new_[40060]_ ;
  assign \new_[40064]_  = ~A202 & ~A200;
  assign \new_[40067]_  = ~A233 & ~A232;
  assign \new_[40068]_  = \new_[40067]_  & \new_[40064]_ ;
  assign \new_[40069]_  = \new_[40068]_  & \new_[40061]_ ;
  assign \new_[40073]_  = ~A268 & ~A267;
  assign \new_[40074]_  = ~A235 & \new_[40073]_ ;
  assign \new_[40077]_  = A298 & ~A269;
  assign \new_[40080]_  = A302 & ~A299;
  assign \new_[40081]_  = \new_[40080]_  & \new_[40077]_ ;
  assign \new_[40082]_  = \new_[40081]_  & \new_[40074]_ ;
  assign \new_[40086]_  = ~A199 & A167;
  assign \new_[40087]_  = A168 & \new_[40086]_ ;
  assign \new_[40090]_  = ~A202 & ~A200;
  assign \new_[40093]_  = ~A233 & ~A232;
  assign \new_[40094]_  = \new_[40093]_  & \new_[40090]_ ;
  assign \new_[40095]_  = \new_[40094]_  & \new_[40087]_ ;
  assign \new_[40099]_  = ~A268 & ~A267;
  assign \new_[40100]_  = ~A235 & \new_[40099]_ ;
  assign \new_[40103]_  = ~A298 & ~A269;
  assign \new_[40106]_  = A302 & A299;
  assign \new_[40107]_  = \new_[40106]_  & \new_[40103]_ ;
  assign \new_[40108]_  = \new_[40107]_  & \new_[40100]_ ;
  assign \new_[40112]_  = ~A199 & A167;
  assign \new_[40113]_  = A168 & \new_[40112]_ ;
  assign \new_[40116]_  = ~A202 & ~A200;
  assign \new_[40119]_  = ~A233 & ~A232;
  assign \new_[40120]_  = \new_[40119]_  & \new_[40116]_ ;
  assign \new_[40121]_  = \new_[40120]_  & \new_[40113]_ ;
  assign \new_[40125]_  = A266 & A265;
  assign \new_[40126]_  = ~A235 & \new_[40125]_ ;
  assign \new_[40129]_  = ~A268 & ~A267;
  assign \new_[40132]_  = A300 & A299;
  assign \new_[40133]_  = \new_[40132]_  & \new_[40129]_ ;
  assign \new_[40134]_  = \new_[40133]_  & \new_[40126]_ ;
  assign \new_[40138]_  = ~A199 & A167;
  assign \new_[40139]_  = A168 & \new_[40138]_ ;
  assign \new_[40142]_  = ~A202 & ~A200;
  assign \new_[40145]_  = ~A233 & ~A232;
  assign \new_[40146]_  = \new_[40145]_  & \new_[40142]_ ;
  assign \new_[40147]_  = \new_[40146]_  & \new_[40139]_ ;
  assign \new_[40151]_  = A266 & A265;
  assign \new_[40152]_  = ~A235 & \new_[40151]_ ;
  assign \new_[40155]_  = ~A268 & ~A267;
  assign \new_[40158]_  = A300 & A298;
  assign \new_[40159]_  = \new_[40158]_  & \new_[40155]_ ;
  assign \new_[40160]_  = \new_[40159]_  & \new_[40152]_ ;
  assign \new_[40164]_  = ~A199 & A167;
  assign \new_[40165]_  = A168 & \new_[40164]_ ;
  assign \new_[40168]_  = ~A202 & ~A200;
  assign \new_[40171]_  = ~A233 & ~A232;
  assign \new_[40172]_  = \new_[40171]_  & \new_[40168]_ ;
  assign \new_[40173]_  = \new_[40172]_  & \new_[40165]_ ;
  assign \new_[40177]_  = ~A266 & ~A265;
  assign \new_[40178]_  = ~A235 & \new_[40177]_ ;
  assign \new_[40181]_  = A298 & ~A268;
  assign \new_[40184]_  = A302 & ~A299;
  assign \new_[40185]_  = \new_[40184]_  & \new_[40181]_ ;
  assign \new_[40186]_  = \new_[40185]_  & \new_[40178]_ ;
  assign \new_[40190]_  = ~A199 & A167;
  assign \new_[40191]_  = A168 & \new_[40190]_ ;
  assign \new_[40194]_  = ~A202 & ~A200;
  assign \new_[40197]_  = ~A233 & ~A232;
  assign \new_[40198]_  = \new_[40197]_  & \new_[40194]_ ;
  assign \new_[40199]_  = \new_[40198]_  & \new_[40191]_ ;
  assign \new_[40203]_  = ~A266 & ~A265;
  assign \new_[40204]_  = ~A235 & \new_[40203]_ ;
  assign \new_[40207]_  = ~A298 & ~A268;
  assign \new_[40210]_  = A302 & A299;
  assign \new_[40211]_  = \new_[40210]_  & \new_[40207]_ ;
  assign \new_[40212]_  = \new_[40211]_  & \new_[40204]_ ;
  assign \new_[40216]_  = ~A166 & A167;
  assign \new_[40217]_  = A170 & \new_[40216]_ ;
  assign \new_[40220]_  = ~A202 & ~A201;
  assign \new_[40223]_  = ~A234 & ~A203;
  assign \new_[40224]_  = \new_[40223]_  & \new_[40220]_ ;
  assign \new_[40225]_  = \new_[40224]_  & \new_[40217]_ ;
  assign \new_[40229]_  = ~A267 & ~A236;
  assign \new_[40230]_  = ~A235 & \new_[40229]_ ;
  assign \new_[40233]_  = ~A269 & ~A268;
  assign \new_[40236]_  = A300 & A299;
  assign \new_[40237]_  = \new_[40236]_  & \new_[40233]_ ;
  assign \new_[40238]_  = \new_[40237]_  & \new_[40230]_ ;
  assign \new_[40242]_  = ~A166 & A167;
  assign \new_[40243]_  = A170 & \new_[40242]_ ;
  assign \new_[40246]_  = ~A202 & ~A201;
  assign \new_[40249]_  = ~A234 & ~A203;
  assign \new_[40250]_  = \new_[40249]_  & \new_[40246]_ ;
  assign \new_[40251]_  = \new_[40250]_  & \new_[40243]_ ;
  assign \new_[40255]_  = ~A267 & ~A236;
  assign \new_[40256]_  = ~A235 & \new_[40255]_ ;
  assign \new_[40259]_  = ~A269 & ~A268;
  assign \new_[40262]_  = A300 & A298;
  assign \new_[40263]_  = \new_[40262]_  & \new_[40259]_ ;
  assign \new_[40264]_  = \new_[40263]_  & \new_[40256]_ ;
  assign \new_[40268]_  = ~A166 & A167;
  assign \new_[40269]_  = A170 & \new_[40268]_ ;
  assign \new_[40272]_  = ~A202 & ~A201;
  assign \new_[40275]_  = ~A234 & ~A203;
  assign \new_[40276]_  = \new_[40275]_  & \new_[40272]_ ;
  assign \new_[40277]_  = \new_[40276]_  & \new_[40269]_ ;
  assign \new_[40281]_  = A265 & ~A236;
  assign \new_[40282]_  = ~A235 & \new_[40281]_ ;
  assign \new_[40285]_  = ~A267 & A266;
  assign \new_[40288]_  = A301 & ~A268;
  assign \new_[40289]_  = \new_[40288]_  & \new_[40285]_ ;
  assign \new_[40290]_  = \new_[40289]_  & \new_[40282]_ ;
  assign \new_[40294]_  = ~A166 & A167;
  assign \new_[40295]_  = A170 & \new_[40294]_ ;
  assign \new_[40298]_  = ~A202 & ~A201;
  assign \new_[40301]_  = ~A234 & ~A203;
  assign \new_[40302]_  = \new_[40301]_  & \new_[40298]_ ;
  assign \new_[40303]_  = \new_[40302]_  & \new_[40295]_ ;
  assign \new_[40307]_  = ~A265 & ~A236;
  assign \new_[40308]_  = ~A235 & \new_[40307]_ ;
  assign \new_[40311]_  = ~A268 & ~A266;
  assign \new_[40314]_  = A300 & A299;
  assign \new_[40315]_  = \new_[40314]_  & \new_[40311]_ ;
  assign \new_[40316]_  = \new_[40315]_  & \new_[40308]_ ;
  assign \new_[40320]_  = ~A166 & A167;
  assign \new_[40321]_  = A170 & \new_[40320]_ ;
  assign \new_[40324]_  = ~A202 & ~A201;
  assign \new_[40327]_  = ~A234 & ~A203;
  assign \new_[40328]_  = \new_[40327]_  & \new_[40324]_ ;
  assign \new_[40329]_  = \new_[40328]_  & \new_[40321]_ ;
  assign \new_[40333]_  = ~A265 & ~A236;
  assign \new_[40334]_  = ~A235 & \new_[40333]_ ;
  assign \new_[40337]_  = ~A268 & ~A266;
  assign \new_[40340]_  = A300 & A298;
  assign \new_[40341]_  = \new_[40340]_  & \new_[40337]_ ;
  assign \new_[40342]_  = \new_[40341]_  & \new_[40334]_ ;
  assign \new_[40346]_  = ~A166 & A167;
  assign \new_[40347]_  = A170 & \new_[40346]_ ;
  assign \new_[40350]_  = ~A202 & ~A201;
  assign \new_[40353]_  = A232 & ~A203;
  assign \new_[40354]_  = \new_[40353]_  & \new_[40350]_ ;
  assign \new_[40355]_  = \new_[40354]_  & \new_[40347]_ ;
  assign \new_[40359]_  = ~A235 & ~A234;
  assign \new_[40360]_  = A233 & \new_[40359]_ ;
  assign \new_[40363]_  = ~A268 & ~A267;
  assign \new_[40366]_  = A301 & ~A269;
  assign \new_[40367]_  = \new_[40366]_  & \new_[40363]_ ;
  assign \new_[40368]_  = \new_[40367]_  & \new_[40360]_ ;
  assign \new_[40372]_  = ~A166 & A167;
  assign \new_[40373]_  = A170 & \new_[40372]_ ;
  assign \new_[40376]_  = ~A202 & ~A201;
  assign \new_[40379]_  = A232 & ~A203;
  assign \new_[40380]_  = \new_[40379]_  & \new_[40376]_ ;
  assign \new_[40381]_  = \new_[40380]_  & \new_[40373]_ ;
  assign \new_[40385]_  = ~A235 & ~A234;
  assign \new_[40386]_  = A233 & \new_[40385]_ ;
  assign \new_[40389]_  = ~A266 & ~A265;
  assign \new_[40392]_  = A301 & ~A268;
  assign \new_[40393]_  = \new_[40392]_  & \new_[40389]_ ;
  assign \new_[40394]_  = \new_[40393]_  & \new_[40386]_ ;
  assign \new_[40398]_  = ~A166 & A167;
  assign \new_[40399]_  = A170 & \new_[40398]_ ;
  assign \new_[40402]_  = ~A202 & ~A201;
  assign \new_[40405]_  = ~A232 & ~A203;
  assign \new_[40406]_  = \new_[40405]_  & \new_[40402]_ ;
  assign \new_[40407]_  = \new_[40406]_  & \new_[40399]_ ;
  assign \new_[40411]_  = ~A267 & ~A235;
  assign \new_[40412]_  = ~A233 & \new_[40411]_ ;
  assign \new_[40415]_  = ~A269 & ~A268;
  assign \new_[40418]_  = A300 & A299;
  assign \new_[40419]_  = \new_[40418]_  & \new_[40415]_ ;
  assign \new_[40420]_  = \new_[40419]_  & \new_[40412]_ ;
  assign \new_[40424]_  = ~A166 & A167;
  assign \new_[40425]_  = A170 & \new_[40424]_ ;
  assign \new_[40428]_  = ~A202 & ~A201;
  assign \new_[40431]_  = ~A232 & ~A203;
  assign \new_[40432]_  = \new_[40431]_  & \new_[40428]_ ;
  assign \new_[40433]_  = \new_[40432]_  & \new_[40425]_ ;
  assign \new_[40437]_  = ~A267 & ~A235;
  assign \new_[40438]_  = ~A233 & \new_[40437]_ ;
  assign \new_[40441]_  = ~A269 & ~A268;
  assign \new_[40444]_  = A300 & A298;
  assign \new_[40445]_  = \new_[40444]_  & \new_[40441]_ ;
  assign \new_[40446]_  = \new_[40445]_  & \new_[40438]_ ;
  assign \new_[40450]_  = ~A166 & A167;
  assign \new_[40451]_  = A170 & \new_[40450]_ ;
  assign \new_[40454]_  = ~A202 & ~A201;
  assign \new_[40457]_  = ~A232 & ~A203;
  assign \new_[40458]_  = \new_[40457]_  & \new_[40454]_ ;
  assign \new_[40459]_  = \new_[40458]_  & \new_[40451]_ ;
  assign \new_[40463]_  = A265 & ~A235;
  assign \new_[40464]_  = ~A233 & \new_[40463]_ ;
  assign \new_[40467]_  = ~A267 & A266;
  assign \new_[40470]_  = A301 & ~A268;
  assign \new_[40471]_  = \new_[40470]_  & \new_[40467]_ ;
  assign \new_[40472]_  = \new_[40471]_  & \new_[40464]_ ;
  assign \new_[40476]_  = ~A166 & A167;
  assign \new_[40477]_  = A170 & \new_[40476]_ ;
  assign \new_[40480]_  = ~A202 & ~A201;
  assign \new_[40483]_  = ~A232 & ~A203;
  assign \new_[40484]_  = \new_[40483]_  & \new_[40480]_ ;
  assign \new_[40485]_  = \new_[40484]_  & \new_[40477]_ ;
  assign \new_[40489]_  = ~A265 & ~A235;
  assign \new_[40490]_  = ~A233 & \new_[40489]_ ;
  assign \new_[40493]_  = ~A268 & ~A266;
  assign \new_[40496]_  = A300 & A299;
  assign \new_[40497]_  = \new_[40496]_  & \new_[40493]_ ;
  assign \new_[40498]_  = \new_[40497]_  & \new_[40490]_ ;
  assign \new_[40502]_  = ~A166 & A167;
  assign \new_[40503]_  = A170 & \new_[40502]_ ;
  assign \new_[40506]_  = ~A202 & ~A201;
  assign \new_[40509]_  = ~A232 & ~A203;
  assign \new_[40510]_  = \new_[40509]_  & \new_[40506]_ ;
  assign \new_[40511]_  = \new_[40510]_  & \new_[40503]_ ;
  assign \new_[40515]_  = ~A265 & ~A235;
  assign \new_[40516]_  = ~A233 & \new_[40515]_ ;
  assign \new_[40519]_  = ~A268 & ~A266;
  assign \new_[40522]_  = A300 & A298;
  assign \new_[40523]_  = \new_[40522]_  & \new_[40519]_ ;
  assign \new_[40524]_  = \new_[40523]_  & \new_[40516]_ ;
  assign \new_[40528]_  = ~A166 & A167;
  assign \new_[40529]_  = A170 & \new_[40528]_ ;
  assign \new_[40532]_  = A200 & A199;
  assign \new_[40535]_  = ~A202 & ~A201;
  assign \new_[40536]_  = \new_[40535]_  & \new_[40532]_ ;
  assign \new_[40537]_  = \new_[40536]_  & \new_[40529]_ ;
  assign \new_[40541]_  = ~A236 & ~A235;
  assign \new_[40542]_  = ~A234 & \new_[40541]_ ;
  assign \new_[40545]_  = ~A268 & ~A267;
  assign \new_[40548]_  = A301 & ~A269;
  assign \new_[40549]_  = \new_[40548]_  & \new_[40545]_ ;
  assign \new_[40550]_  = \new_[40549]_  & \new_[40542]_ ;
  assign \new_[40554]_  = ~A166 & A167;
  assign \new_[40555]_  = A170 & \new_[40554]_ ;
  assign \new_[40558]_  = A200 & A199;
  assign \new_[40561]_  = ~A202 & ~A201;
  assign \new_[40562]_  = \new_[40561]_  & \new_[40558]_ ;
  assign \new_[40563]_  = \new_[40562]_  & \new_[40555]_ ;
  assign \new_[40567]_  = ~A236 & ~A235;
  assign \new_[40568]_  = ~A234 & \new_[40567]_ ;
  assign \new_[40571]_  = ~A266 & ~A265;
  assign \new_[40574]_  = A301 & ~A268;
  assign \new_[40575]_  = \new_[40574]_  & \new_[40571]_ ;
  assign \new_[40576]_  = \new_[40575]_  & \new_[40568]_ ;
  assign \new_[40580]_  = ~A166 & A167;
  assign \new_[40581]_  = A170 & \new_[40580]_ ;
  assign \new_[40584]_  = A200 & A199;
  assign \new_[40587]_  = ~A202 & ~A201;
  assign \new_[40588]_  = \new_[40587]_  & \new_[40584]_ ;
  assign \new_[40589]_  = \new_[40588]_  & \new_[40581]_ ;
  assign \new_[40593]_  = A236 & A233;
  assign \new_[40594]_  = ~A232 & \new_[40593]_ ;
  assign \new_[40597]_  = A299 & A298;
  assign \new_[40600]_  = ~A301 & ~A300;
  assign \new_[40601]_  = \new_[40600]_  & \new_[40597]_ ;
  assign \new_[40602]_  = \new_[40601]_  & \new_[40594]_ ;
  assign \new_[40606]_  = ~A166 & A167;
  assign \new_[40607]_  = A170 & \new_[40606]_ ;
  assign \new_[40610]_  = A200 & A199;
  assign \new_[40613]_  = ~A202 & ~A201;
  assign \new_[40614]_  = \new_[40613]_  & \new_[40610]_ ;
  assign \new_[40615]_  = \new_[40614]_  & \new_[40607]_ ;
  assign \new_[40619]_  = A236 & ~A233;
  assign \new_[40620]_  = A232 & \new_[40619]_ ;
  assign \new_[40623]_  = A299 & A298;
  assign \new_[40626]_  = ~A301 & ~A300;
  assign \new_[40627]_  = \new_[40626]_  & \new_[40623]_ ;
  assign \new_[40628]_  = \new_[40627]_  & \new_[40620]_ ;
  assign \new_[40632]_  = ~A166 & A167;
  assign \new_[40633]_  = A170 & \new_[40632]_ ;
  assign \new_[40636]_  = A200 & A199;
  assign \new_[40639]_  = ~A202 & ~A201;
  assign \new_[40640]_  = \new_[40639]_  & \new_[40636]_ ;
  assign \new_[40641]_  = \new_[40640]_  & \new_[40633]_ ;
  assign \new_[40645]_  = ~A235 & ~A233;
  assign \new_[40646]_  = ~A232 & \new_[40645]_ ;
  assign \new_[40649]_  = ~A268 & ~A267;
  assign \new_[40652]_  = A301 & ~A269;
  assign \new_[40653]_  = \new_[40652]_  & \new_[40649]_ ;
  assign \new_[40654]_  = \new_[40653]_  & \new_[40646]_ ;
  assign \new_[40658]_  = ~A166 & A167;
  assign \new_[40659]_  = A170 & \new_[40658]_ ;
  assign \new_[40662]_  = A200 & A199;
  assign \new_[40665]_  = ~A202 & ~A201;
  assign \new_[40666]_  = \new_[40665]_  & \new_[40662]_ ;
  assign \new_[40667]_  = \new_[40666]_  & \new_[40659]_ ;
  assign \new_[40671]_  = ~A235 & ~A233;
  assign \new_[40672]_  = ~A232 & \new_[40671]_ ;
  assign \new_[40675]_  = ~A266 & ~A265;
  assign \new_[40678]_  = A301 & ~A268;
  assign \new_[40679]_  = \new_[40678]_  & \new_[40675]_ ;
  assign \new_[40680]_  = \new_[40679]_  & \new_[40672]_ ;
  assign \new_[40684]_  = ~A166 & A167;
  assign \new_[40685]_  = A170 & \new_[40684]_ ;
  assign \new_[40688]_  = ~A200 & ~A199;
  assign \new_[40691]_  = ~A234 & ~A202;
  assign \new_[40692]_  = \new_[40691]_  & \new_[40688]_ ;
  assign \new_[40693]_  = \new_[40692]_  & \new_[40685]_ ;
  assign \new_[40697]_  = ~A267 & ~A236;
  assign \new_[40698]_  = ~A235 & \new_[40697]_ ;
  assign \new_[40701]_  = ~A269 & ~A268;
  assign \new_[40704]_  = A300 & A299;
  assign \new_[40705]_  = \new_[40704]_  & \new_[40701]_ ;
  assign \new_[40706]_  = \new_[40705]_  & \new_[40698]_ ;
  assign \new_[40710]_  = ~A166 & A167;
  assign \new_[40711]_  = A170 & \new_[40710]_ ;
  assign \new_[40714]_  = ~A200 & ~A199;
  assign \new_[40717]_  = ~A234 & ~A202;
  assign \new_[40718]_  = \new_[40717]_  & \new_[40714]_ ;
  assign \new_[40719]_  = \new_[40718]_  & \new_[40711]_ ;
  assign \new_[40723]_  = ~A267 & ~A236;
  assign \new_[40724]_  = ~A235 & \new_[40723]_ ;
  assign \new_[40727]_  = ~A269 & ~A268;
  assign \new_[40730]_  = A300 & A298;
  assign \new_[40731]_  = \new_[40730]_  & \new_[40727]_ ;
  assign \new_[40732]_  = \new_[40731]_  & \new_[40724]_ ;
  assign \new_[40736]_  = ~A166 & A167;
  assign \new_[40737]_  = A170 & \new_[40736]_ ;
  assign \new_[40740]_  = ~A200 & ~A199;
  assign \new_[40743]_  = ~A234 & ~A202;
  assign \new_[40744]_  = \new_[40743]_  & \new_[40740]_ ;
  assign \new_[40745]_  = \new_[40744]_  & \new_[40737]_ ;
  assign \new_[40749]_  = A265 & ~A236;
  assign \new_[40750]_  = ~A235 & \new_[40749]_ ;
  assign \new_[40753]_  = ~A267 & A266;
  assign \new_[40756]_  = A301 & ~A268;
  assign \new_[40757]_  = \new_[40756]_  & \new_[40753]_ ;
  assign \new_[40758]_  = \new_[40757]_  & \new_[40750]_ ;
  assign \new_[40762]_  = ~A166 & A167;
  assign \new_[40763]_  = A170 & \new_[40762]_ ;
  assign \new_[40766]_  = ~A200 & ~A199;
  assign \new_[40769]_  = ~A234 & ~A202;
  assign \new_[40770]_  = \new_[40769]_  & \new_[40766]_ ;
  assign \new_[40771]_  = \new_[40770]_  & \new_[40763]_ ;
  assign \new_[40775]_  = ~A265 & ~A236;
  assign \new_[40776]_  = ~A235 & \new_[40775]_ ;
  assign \new_[40779]_  = ~A268 & ~A266;
  assign \new_[40782]_  = A300 & A299;
  assign \new_[40783]_  = \new_[40782]_  & \new_[40779]_ ;
  assign \new_[40784]_  = \new_[40783]_  & \new_[40776]_ ;
  assign \new_[40788]_  = ~A166 & A167;
  assign \new_[40789]_  = A170 & \new_[40788]_ ;
  assign \new_[40792]_  = ~A200 & ~A199;
  assign \new_[40795]_  = ~A234 & ~A202;
  assign \new_[40796]_  = \new_[40795]_  & \new_[40792]_ ;
  assign \new_[40797]_  = \new_[40796]_  & \new_[40789]_ ;
  assign \new_[40801]_  = ~A265 & ~A236;
  assign \new_[40802]_  = ~A235 & \new_[40801]_ ;
  assign \new_[40805]_  = ~A268 & ~A266;
  assign \new_[40808]_  = A300 & A298;
  assign \new_[40809]_  = \new_[40808]_  & \new_[40805]_ ;
  assign \new_[40810]_  = \new_[40809]_  & \new_[40802]_ ;
  assign \new_[40814]_  = ~A166 & A167;
  assign \new_[40815]_  = A170 & \new_[40814]_ ;
  assign \new_[40818]_  = ~A200 & ~A199;
  assign \new_[40821]_  = A232 & ~A202;
  assign \new_[40822]_  = \new_[40821]_  & \new_[40818]_ ;
  assign \new_[40823]_  = \new_[40822]_  & \new_[40815]_ ;
  assign \new_[40827]_  = ~A235 & ~A234;
  assign \new_[40828]_  = A233 & \new_[40827]_ ;
  assign \new_[40831]_  = ~A268 & ~A267;
  assign \new_[40834]_  = A301 & ~A269;
  assign \new_[40835]_  = \new_[40834]_  & \new_[40831]_ ;
  assign \new_[40836]_  = \new_[40835]_  & \new_[40828]_ ;
  assign \new_[40840]_  = ~A166 & A167;
  assign \new_[40841]_  = A170 & \new_[40840]_ ;
  assign \new_[40844]_  = ~A200 & ~A199;
  assign \new_[40847]_  = A232 & ~A202;
  assign \new_[40848]_  = \new_[40847]_  & \new_[40844]_ ;
  assign \new_[40849]_  = \new_[40848]_  & \new_[40841]_ ;
  assign \new_[40853]_  = ~A235 & ~A234;
  assign \new_[40854]_  = A233 & \new_[40853]_ ;
  assign \new_[40857]_  = ~A266 & ~A265;
  assign \new_[40860]_  = A301 & ~A268;
  assign \new_[40861]_  = \new_[40860]_  & \new_[40857]_ ;
  assign \new_[40862]_  = \new_[40861]_  & \new_[40854]_ ;
  assign \new_[40866]_  = ~A166 & A167;
  assign \new_[40867]_  = A170 & \new_[40866]_ ;
  assign \new_[40870]_  = ~A200 & ~A199;
  assign \new_[40873]_  = ~A232 & ~A202;
  assign \new_[40874]_  = \new_[40873]_  & \new_[40870]_ ;
  assign \new_[40875]_  = \new_[40874]_  & \new_[40867]_ ;
  assign \new_[40879]_  = ~A267 & ~A235;
  assign \new_[40880]_  = ~A233 & \new_[40879]_ ;
  assign \new_[40883]_  = ~A269 & ~A268;
  assign \new_[40886]_  = A300 & A299;
  assign \new_[40887]_  = \new_[40886]_  & \new_[40883]_ ;
  assign \new_[40888]_  = \new_[40887]_  & \new_[40880]_ ;
  assign \new_[40892]_  = ~A166 & A167;
  assign \new_[40893]_  = A170 & \new_[40892]_ ;
  assign \new_[40896]_  = ~A200 & ~A199;
  assign \new_[40899]_  = ~A232 & ~A202;
  assign \new_[40900]_  = \new_[40899]_  & \new_[40896]_ ;
  assign \new_[40901]_  = \new_[40900]_  & \new_[40893]_ ;
  assign \new_[40905]_  = ~A267 & ~A235;
  assign \new_[40906]_  = ~A233 & \new_[40905]_ ;
  assign \new_[40909]_  = ~A269 & ~A268;
  assign \new_[40912]_  = A300 & A298;
  assign \new_[40913]_  = \new_[40912]_  & \new_[40909]_ ;
  assign \new_[40914]_  = \new_[40913]_  & \new_[40906]_ ;
  assign \new_[40918]_  = ~A166 & A167;
  assign \new_[40919]_  = A170 & \new_[40918]_ ;
  assign \new_[40922]_  = ~A200 & ~A199;
  assign \new_[40925]_  = ~A232 & ~A202;
  assign \new_[40926]_  = \new_[40925]_  & \new_[40922]_ ;
  assign \new_[40927]_  = \new_[40926]_  & \new_[40919]_ ;
  assign \new_[40931]_  = A265 & ~A235;
  assign \new_[40932]_  = ~A233 & \new_[40931]_ ;
  assign \new_[40935]_  = ~A267 & A266;
  assign \new_[40938]_  = A301 & ~A268;
  assign \new_[40939]_  = \new_[40938]_  & \new_[40935]_ ;
  assign \new_[40940]_  = \new_[40939]_  & \new_[40932]_ ;
  assign \new_[40944]_  = ~A166 & A167;
  assign \new_[40945]_  = A170 & \new_[40944]_ ;
  assign \new_[40948]_  = ~A200 & ~A199;
  assign \new_[40951]_  = ~A232 & ~A202;
  assign \new_[40952]_  = \new_[40951]_  & \new_[40948]_ ;
  assign \new_[40953]_  = \new_[40952]_  & \new_[40945]_ ;
  assign \new_[40957]_  = ~A265 & ~A235;
  assign \new_[40958]_  = ~A233 & \new_[40957]_ ;
  assign \new_[40961]_  = ~A268 & ~A266;
  assign \new_[40964]_  = A300 & A299;
  assign \new_[40965]_  = \new_[40964]_  & \new_[40961]_ ;
  assign \new_[40966]_  = \new_[40965]_  & \new_[40958]_ ;
  assign \new_[40970]_  = ~A166 & A167;
  assign \new_[40971]_  = A170 & \new_[40970]_ ;
  assign \new_[40974]_  = ~A200 & ~A199;
  assign \new_[40977]_  = ~A232 & ~A202;
  assign \new_[40978]_  = \new_[40977]_  & \new_[40974]_ ;
  assign \new_[40979]_  = \new_[40978]_  & \new_[40971]_ ;
  assign \new_[40983]_  = ~A265 & ~A235;
  assign \new_[40984]_  = ~A233 & \new_[40983]_ ;
  assign \new_[40987]_  = ~A268 & ~A266;
  assign \new_[40990]_  = A300 & A298;
  assign \new_[40991]_  = \new_[40990]_  & \new_[40987]_ ;
  assign \new_[40992]_  = \new_[40991]_  & \new_[40984]_ ;
  assign \new_[40996]_  = A166 & ~A167;
  assign \new_[40997]_  = A170 & \new_[40996]_ ;
  assign \new_[41000]_  = ~A202 & ~A201;
  assign \new_[41003]_  = ~A234 & ~A203;
  assign \new_[41004]_  = \new_[41003]_  & \new_[41000]_ ;
  assign \new_[41005]_  = \new_[41004]_  & \new_[40997]_ ;
  assign \new_[41009]_  = ~A267 & ~A236;
  assign \new_[41010]_  = ~A235 & \new_[41009]_ ;
  assign \new_[41013]_  = ~A269 & ~A268;
  assign \new_[41016]_  = A300 & A299;
  assign \new_[41017]_  = \new_[41016]_  & \new_[41013]_ ;
  assign \new_[41018]_  = \new_[41017]_  & \new_[41010]_ ;
  assign \new_[41022]_  = A166 & ~A167;
  assign \new_[41023]_  = A170 & \new_[41022]_ ;
  assign \new_[41026]_  = ~A202 & ~A201;
  assign \new_[41029]_  = ~A234 & ~A203;
  assign \new_[41030]_  = \new_[41029]_  & \new_[41026]_ ;
  assign \new_[41031]_  = \new_[41030]_  & \new_[41023]_ ;
  assign \new_[41035]_  = ~A267 & ~A236;
  assign \new_[41036]_  = ~A235 & \new_[41035]_ ;
  assign \new_[41039]_  = ~A269 & ~A268;
  assign \new_[41042]_  = A300 & A298;
  assign \new_[41043]_  = \new_[41042]_  & \new_[41039]_ ;
  assign \new_[41044]_  = \new_[41043]_  & \new_[41036]_ ;
  assign \new_[41048]_  = A166 & ~A167;
  assign \new_[41049]_  = A170 & \new_[41048]_ ;
  assign \new_[41052]_  = ~A202 & ~A201;
  assign \new_[41055]_  = ~A234 & ~A203;
  assign \new_[41056]_  = \new_[41055]_  & \new_[41052]_ ;
  assign \new_[41057]_  = \new_[41056]_  & \new_[41049]_ ;
  assign \new_[41061]_  = A265 & ~A236;
  assign \new_[41062]_  = ~A235 & \new_[41061]_ ;
  assign \new_[41065]_  = ~A267 & A266;
  assign \new_[41068]_  = A301 & ~A268;
  assign \new_[41069]_  = \new_[41068]_  & \new_[41065]_ ;
  assign \new_[41070]_  = \new_[41069]_  & \new_[41062]_ ;
  assign \new_[41074]_  = A166 & ~A167;
  assign \new_[41075]_  = A170 & \new_[41074]_ ;
  assign \new_[41078]_  = ~A202 & ~A201;
  assign \new_[41081]_  = ~A234 & ~A203;
  assign \new_[41082]_  = \new_[41081]_  & \new_[41078]_ ;
  assign \new_[41083]_  = \new_[41082]_  & \new_[41075]_ ;
  assign \new_[41087]_  = ~A265 & ~A236;
  assign \new_[41088]_  = ~A235 & \new_[41087]_ ;
  assign \new_[41091]_  = ~A268 & ~A266;
  assign \new_[41094]_  = A300 & A299;
  assign \new_[41095]_  = \new_[41094]_  & \new_[41091]_ ;
  assign \new_[41096]_  = \new_[41095]_  & \new_[41088]_ ;
  assign \new_[41100]_  = A166 & ~A167;
  assign \new_[41101]_  = A170 & \new_[41100]_ ;
  assign \new_[41104]_  = ~A202 & ~A201;
  assign \new_[41107]_  = ~A234 & ~A203;
  assign \new_[41108]_  = \new_[41107]_  & \new_[41104]_ ;
  assign \new_[41109]_  = \new_[41108]_  & \new_[41101]_ ;
  assign \new_[41113]_  = ~A265 & ~A236;
  assign \new_[41114]_  = ~A235 & \new_[41113]_ ;
  assign \new_[41117]_  = ~A268 & ~A266;
  assign \new_[41120]_  = A300 & A298;
  assign \new_[41121]_  = \new_[41120]_  & \new_[41117]_ ;
  assign \new_[41122]_  = \new_[41121]_  & \new_[41114]_ ;
  assign \new_[41126]_  = A166 & ~A167;
  assign \new_[41127]_  = A170 & \new_[41126]_ ;
  assign \new_[41130]_  = ~A202 & ~A201;
  assign \new_[41133]_  = A232 & ~A203;
  assign \new_[41134]_  = \new_[41133]_  & \new_[41130]_ ;
  assign \new_[41135]_  = \new_[41134]_  & \new_[41127]_ ;
  assign \new_[41139]_  = ~A235 & ~A234;
  assign \new_[41140]_  = A233 & \new_[41139]_ ;
  assign \new_[41143]_  = ~A268 & ~A267;
  assign \new_[41146]_  = A301 & ~A269;
  assign \new_[41147]_  = \new_[41146]_  & \new_[41143]_ ;
  assign \new_[41148]_  = \new_[41147]_  & \new_[41140]_ ;
  assign \new_[41152]_  = A166 & ~A167;
  assign \new_[41153]_  = A170 & \new_[41152]_ ;
  assign \new_[41156]_  = ~A202 & ~A201;
  assign \new_[41159]_  = A232 & ~A203;
  assign \new_[41160]_  = \new_[41159]_  & \new_[41156]_ ;
  assign \new_[41161]_  = \new_[41160]_  & \new_[41153]_ ;
  assign \new_[41165]_  = ~A235 & ~A234;
  assign \new_[41166]_  = A233 & \new_[41165]_ ;
  assign \new_[41169]_  = ~A266 & ~A265;
  assign \new_[41172]_  = A301 & ~A268;
  assign \new_[41173]_  = \new_[41172]_  & \new_[41169]_ ;
  assign \new_[41174]_  = \new_[41173]_  & \new_[41166]_ ;
  assign \new_[41178]_  = A166 & ~A167;
  assign \new_[41179]_  = A170 & \new_[41178]_ ;
  assign \new_[41182]_  = ~A202 & ~A201;
  assign \new_[41185]_  = ~A232 & ~A203;
  assign \new_[41186]_  = \new_[41185]_  & \new_[41182]_ ;
  assign \new_[41187]_  = \new_[41186]_  & \new_[41179]_ ;
  assign \new_[41191]_  = ~A267 & ~A235;
  assign \new_[41192]_  = ~A233 & \new_[41191]_ ;
  assign \new_[41195]_  = ~A269 & ~A268;
  assign \new_[41198]_  = A300 & A299;
  assign \new_[41199]_  = \new_[41198]_  & \new_[41195]_ ;
  assign \new_[41200]_  = \new_[41199]_  & \new_[41192]_ ;
  assign \new_[41204]_  = A166 & ~A167;
  assign \new_[41205]_  = A170 & \new_[41204]_ ;
  assign \new_[41208]_  = ~A202 & ~A201;
  assign \new_[41211]_  = ~A232 & ~A203;
  assign \new_[41212]_  = \new_[41211]_  & \new_[41208]_ ;
  assign \new_[41213]_  = \new_[41212]_  & \new_[41205]_ ;
  assign \new_[41217]_  = ~A267 & ~A235;
  assign \new_[41218]_  = ~A233 & \new_[41217]_ ;
  assign \new_[41221]_  = ~A269 & ~A268;
  assign \new_[41224]_  = A300 & A298;
  assign \new_[41225]_  = \new_[41224]_  & \new_[41221]_ ;
  assign \new_[41226]_  = \new_[41225]_  & \new_[41218]_ ;
  assign \new_[41230]_  = A166 & ~A167;
  assign \new_[41231]_  = A170 & \new_[41230]_ ;
  assign \new_[41234]_  = ~A202 & ~A201;
  assign \new_[41237]_  = ~A232 & ~A203;
  assign \new_[41238]_  = \new_[41237]_  & \new_[41234]_ ;
  assign \new_[41239]_  = \new_[41238]_  & \new_[41231]_ ;
  assign \new_[41243]_  = A265 & ~A235;
  assign \new_[41244]_  = ~A233 & \new_[41243]_ ;
  assign \new_[41247]_  = ~A267 & A266;
  assign \new_[41250]_  = A301 & ~A268;
  assign \new_[41251]_  = \new_[41250]_  & \new_[41247]_ ;
  assign \new_[41252]_  = \new_[41251]_  & \new_[41244]_ ;
  assign \new_[41256]_  = A166 & ~A167;
  assign \new_[41257]_  = A170 & \new_[41256]_ ;
  assign \new_[41260]_  = ~A202 & ~A201;
  assign \new_[41263]_  = ~A232 & ~A203;
  assign \new_[41264]_  = \new_[41263]_  & \new_[41260]_ ;
  assign \new_[41265]_  = \new_[41264]_  & \new_[41257]_ ;
  assign \new_[41269]_  = ~A265 & ~A235;
  assign \new_[41270]_  = ~A233 & \new_[41269]_ ;
  assign \new_[41273]_  = ~A268 & ~A266;
  assign \new_[41276]_  = A300 & A299;
  assign \new_[41277]_  = \new_[41276]_  & \new_[41273]_ ;
  assign \new_[41278]_  = \new_[41277]_  & \new_[41270]_ ;
  assign \new_[41282]_  = A166 & ~A167;
  assign \new_[41283]_  = A170 & \new_[41282]_ ;
  assign \new_[41286]_  = ~A202 & ~A201;
  assign \new_[41289]_  = ~A232 & ~A203;
  assign \new_[41290]_  = \new_[41289]_  & \new_[41286]_ ;
  assign \new_[41291]_  = \new_[41290]_  & \new_[41283]_ ;
  assign \new_[41295]_  = ~A265 & ~A235;
  assign \new_[41296]_  = ~A233 & \new_[41295]_ ;
  assign \new_[41299]_  = ~A268 & ~A266;
  assign \new_[41302]_  = A300 & A298;
  assign \new_[41303]_  = \new_[41302]_  & \new_[41299]_ ;
  assign \new_[41304]_  = \new_[41303]_  & \new_[41296]_ ;
  assign \new_[41308]_  = A166 & ~A167;
  assign \new_[41309]_  = A170 & \new_[41308]_ ;
  assign \new_[41312]_  = A200 & A199;
  assign \new_[41315]_  = ~A202 & ~A201;
  assign \new_[41316]_  = \new_[41315]_  & \new_[41312]_ ;
  assign \new_[41317]_  = \new_[41316]_  & \new_[41309]_ ;
  assign \new_[41321]_  = ~A236 & ~A235;
  assign \new_[41322]_  = ~A234 & \new_[41321]_ ;
  assign \new_[41325]_  = ~A268 & ~A267;
  assign \new_[41328]_  = A301 & ~A269;
  assign \new_[41329]_  = \new_[41328]_  & \new_[41325]_ ;
  assign \new_[41330]_  = \new_[41329]_  & \new_[41322]_ ;
  assign \new_[41334]_  = A166 & ~A167;
  assign \new_[41335]_  = A170 & \new_[41334]_ ;
  assign \new_[41338]_  = A200 & A199;
  assign \new_[41341]_  = ~A202 & ~A201;
  assign \new_[41342]_  = \new_[41341]_  & \new_[41338]_ ;
  assign \new_[41343]_  = \new_[41342]_  & \new_[41335]_ ;
  assign \new_[41347]_  = ~A236 & ~A235;
  assign \new_[41348]_  = ~A234 & \new_[41347]_ ;
  assign \new_[41351]_  = ~A266 & ~A265;
  assign \new_[41354]_  = A301 & ~A268;
  assign \new_[41355]_  = \new_[41354]_  & \new_[41351]_ ;
  assign \new_[41356]_  = \new_[41355]_  & \new_[41348]_ ;
  assign \new_[41360]_  = A166 & ~A167;
  assign \new_[41361]_  = A170 & \new_[41360]_ ;
  assign \new_[41364]_  = A200 & A199;
  assign \new_[41367]_  = ~A202 & ~A201;
  assign \new_[41368]_  = \new_[41367]_  & \new_[41364]_ ;
  assign \new_[41369]_  = \new_[41368]_  & \new_[41361]_ ;
  assign \new_[41373]_  = A236 & A233;
  assign \new_[41374]_  = ~A232 & \new_[41373]_ ;
  assign \new_[41377]_  = A299 & A298;
  assign \new_[41380]_  = ~A301 & ~A300;
  assign \new_[41381]_  = \new_[41380]_  & \new_[41377]_ ;
  assign \new_[41382]_  = \new_[41381]_  & \new_[41374]_ ;
  assign \new_[41386]_  = A166 & ~A167;
  assign \new_[41387]_  = A170 & \new_[41386]_ ;
  assign \new_[41390]_  = A200 & A199;
  assign \new_[41393]_  = ~A202 & ~A201;
  assign \new_[41394]_  = \new_[41393]_  & \new_[41390]_ ;
  assign \new_[41395]_  = \new_[41394]_  & \new_[41387]_ ;
  assign \new_[41399]_  = A236 & ~A233;
  assign \new_[41400]_  = A232 & \new_[41399]_ ;
  assign \new_[41403]_  = A299 & A298;
  assign \new_[41406]_  = ~A301 & ~A300;
  assign \new_[41407]_  = \new_[41406]_  & \new_[41403]_ ;
  assign \new_[41408]_  = \new_[41407]_  & \new_[41400]_ ;
  assign \new_[41412]_  = A166 & ~A167;
  assign \new_[41413]_  = A170 & \new_[41412]_ ;
  assign \new_[41416]_  = A200 & A199;
  assign \new_[41419]_  = ~A202 & ~A201;
  assign \new_[41420]_  = \new_[41419]_  & \new_[41416]_ ;
  assign \new_[41421]_  = \new_[41420]_  & \new_[41413]_ ;
  assign \new_[41425]_  = ~A235 & ~A233;
  assign \new_[41426]_  = ~A232 & \new_[41425]_ ;
  assign \new_[41429]_  = ~A268 & ~A267;
  assign \new_[41432]_  = A301 & ~A269;
  assign \new_[41433]_  = \new_[41432]_  & \new_[41429]_ ;
  assign \new_[41434]_  = \new_[41433]_  & \new_[41426]_ ;
  assign \new_[41438]_  = A166 & ~A167;
  assign \new_[41439]_  = A170 & \new_[41438]_ ;
  assign \new_[41442]_  = A200 & A199;
  assign \new_[41445]_  = ~A202 & ~A201;
  assign \new_[41446]_  = \new_[41445]_  & \new_[41442]_ ;
  assign \new_[41447]_  = \new_[41446]_  & \new_[41439]_ ;
  assign \new_[41451]_  = ~A235 & ~A233;
  assign \new_[41452]_  = ~A232 & \new_[41451]_ ;
  assign \new_[41455]_  = ~A266 & ~A265;
  assign \new_[41458]_  = A301 & ~A268;
  assign \new_[41459]_  = \new_[41458]_  & \new_[41455]_ ;
  assign \new_[41460]_  = \new_[41459]_  & \new_[41452]_ ;
  assign \new_[41464]_  = A166 & ~A167;
  assign \new_[41465]_  = A170 & \new_[41464]_ ;
  assign \new_[41468]_  = ~A200 & ~A199;
  assign \new_[41471]_  = ~A234 & ~A202;
  assign \new_[41472]_  = \new_[41471]_  & \new_[41468]_ ;
  assign \new_[41473]_  = \new_[41472]_  & \new_[41465]_ ;
  assign \new_[41477]_  = ~A267 & ~A236;
  assign \new_[41478]_  = ~A235 & \new_[41477]_ ;
  assign \new_[41481]_  = ~A269 & ~A268;
  assign \new_[41484]_  = A300 & A299;
  assign \new_[41485]_  = \new_[41484]_  & \new_[41481]_ ;
  assign \new_[41486]_  = \new_[41485]_  & \new_[41478]_ ;
  assign \new_[41490]_  = A166 & ~A167;
  assign \new_[41491]_  = A170 & \new_[41490]_ ;
  assign \new_[41494]_  = ~A200 & ~A199;
  assign \new_[41497]_  = ~A234 & ~A202;
  assign \new_[41498]_  = \new_[41497]_  & \new_[41494]_ ;
  assign \new_[41499]_  = \new_[41498]_  & \new_[41491]_ ;
  assign \new_[41503]_  = ~A267 & ~A236;
  assign \new_[41504]_  = ~A235 & \new_[41503]_ ;
  assign \new_[41507]_  = ~A269 & ~A268;
  assign \new_[41510]_  = A300 & A298;
  assign \new_[41511]_  = \new_[41510]_  & \new_[41507]_ ;
  assign \new_[41512]_  = \new_[41511]_  & \new_[41504]_ ;
  assign \new_[41516]_  = A166 & ~A167;
  assign \new_[41517]_  = A170 & \new_[41516]_ ;
  assign \new_[41520]_  = ~A200 & ~A199;
  assign \new_[41523]_  = ~A234 & ~A202;
  assign \new_[41524]_  = \new_[41523]_  & \new_[41520]_ ;
  assign \new_[41525]_  = \new_[41524]_  & \new_[41517]_ ;
  assign \new_[41529]_  = A265 & ~A236;
  assign \new_[41530]_  = ~A235 & \new_[41529]_ ;
  assign \new_[41533]_  = ~A267 & A266;
  assign \new_[41536]_  = A301 & ~A268;
  assign \new_[41537]_  = \new_[41536]_  & \new_[41533]_ ;
  assign \new_[41538]_  = \new_[41537]_  & \new_[41530]_ ;
  assign \new_[41542]_  = A166 & ~A167;
  assign \new_[41543]_  = A170 & \new_[41542]_ ;
  assign \new_[41546]_  = ~A200 & ~A199;
  assign \new_[41549]_  = ~A234 & ~A202;
  assign \new_[41550]_  = \new_[41549]_  & \new_[41546]_ ;
  assign \new_[41551]_  = \new_[41550]_  & \new_[41543]_ ;
  assign \new_[41555]_  = ~A265 & ~A236;
  assign \new_[41556]_  = ~A235 & \new_[41555]_ ;
  assign \new_[41559]_  = ~A268 & ~A266;
  assign \new_[41562]_  = A300 & A299;
  assign \new_[41563]_  = \new_[41562]_  & \new_[41559]_ ;
  assign \new_[41564]_  = \new_[41563]_  & \new_[41556]_ ;
  assign \new_[41568]_  = A166 & ~A167;
  assign \new_[41569]_  = A170 & \new_[41568]_ ;
  assign \new_[41572]_  = ~A200 & ~A199;
  assign \new_[41575]_  = ~A234 & ~A202;
  assign \new_[41576]_  = \new_[41575]_  & \new_[41572]_ ;
  assign \new_[41577]_  = \new_[41576]_  & \new_[41569]_ ;
  assign \new_[41581]_  = ~A265 & ~A236;
  assign \new_[41582]_  = ~A235 & \new_[41581]_ ;
  assign \new_[41585]_  = ~A268 & ~A266;
  assign \new_[41588]_  = A300 & A298;
  assign \new_[41589]_  = \new_[41588]_  & \new_[41585]_ ;
  assign \new_[41590]_  = \new_[41589]_  & \new_[41582]_ ;
  assign \new_[41594]_  = A166 & ~A167;
  assign \new_[41595]_  = A170 & \new_[41594]_ ;
  assign \new_[41598]_  = ~A200 & ~A199;
  assign \new_[41601]_  = A232 & ~A202;
  assign \new_[41602]_  = \new_[41601]_  & \new_[41598]_ ;
  assign \new_[41603]_  = \new_[41602]_  & \new_[41595]_ ;
  assign \new_[41607]_  = ~A235 & ~A234;
  assign \new_[41608]_  = A233 & \new_[41607]_ ;
  assign \new_[41611]_  = ~A268 & ~A267;
  assign \new_[41614]_  = A301 & ~A269;
  assign \new_[41615]_  = \new_[41614]_  & \new_[41611]_ ;
  assign \new_[41616]_  = \new_[41615]_  & \new_[41608]_ ;
  assign \new_[41620]_  = A166 & ~A167;
  assign \new_[41621]_  = A170 & \new_[41620]_ ;
  assign \new_[41624]_  = ~A200 & ~A199;
  assign \new_[41627]_  = A232 & ~A202;
  assign \new_[41628]_  = \new_[41627]_  & \new_[41624]_ ;
  assign \new_[41629]_  = \new_[41628]_  & \new_[41621]_ ;
  assign \new_[41633]_  = ~A235 & ~A234;
  assign \new_[41634]_  = A233 & \new_[41633]_ ;
  assign \new_[41637]_  = ~A266 & ~A265;
  assign \new_[41640]_  = A301 & ~A268;
  assign \new_[41641]_  = \new_[41640]_  & \new_[41637]_ ;
  assign \new_[41642]_  = \new_[41641]_  & \new_[41634]_ ;
  assign \new_[41646]_  = A166 & ~A167;
  assign \new_[41647]_  = A170 & \new_[41646]_ ;
  assign \new_[41650]_  = ~A200 & ~A199;
  assign \new_[41653]_  = ~A232 & ~A202;
  assign \new_[41654]_  = \new_[41653]_  & \new_[41650]_ ;
  assign \new_[41655]_  = \new_[41654]_  & \new_[41647]_ ;
  assign \new_[41659]_  = ~A267 & ~A235;
  assign \new_[41660]_  = ~A233 & \new_[41659]_ ;
  assign \new_[41663]_  = ~A269 & ~A268;
  assign \new_[41666]_  = A300 & A299;
  assign \new_[41667]_  = \new_[41666]_  & \new_[41663]_ ;
  assign \new_[41668]_  = \new_[41667]_  & \new_[41660]_ ;
  assign \new_[41672]_  = A166 & ~A167;
  assign \new_[41673]_  = A170 & \new_[41672]_ ;
  assign \new_[41676]_  = ~A200 & ~A199;
  assign \new_[41679]_  = ~A232 & ~A202;
  assign \new_[41680]_  = \new_[41679]_  & \new_[41676]_ ;
  assign \new_[41681]_  = \new_[41680]_  & \new_[41673]_ ;
  assign \new_[41685]_  = ~A267 & ~A235;
  assign \new_[41686]_  = ~A233 & \new_[41685]_ ;
  assign \new_[41689]_  = ~A269 & ~A268;
  assign \new_[41692]_  = A300 & A298;
  assign \new_[41693]_  = \new_[41692]_  & \new_[41689]_ ;
  assign \new_[41694]_  = \new_[41693]_  & \new_[41686]_ ;
  assign \new_[41698]_  = A166 & ~A167;
  assign \new_[41699]_  = A170 & \new_[41698]_ ;
  assign \new_[41702]_  = ~A200 & ~A199;
  assign \new_[41705]_  = ~A232 & ~A202;
  assign \new_[41706]_  = \new_[41705]_  & \new_[41702]_ ;
  assign \new_[41707]_  = \new_[41706]_  & \new_[41699]_ ;
  assign \new_[41711]_  = A265 & ~A235;
  assign \new_[41712]_  = ~A233 & \new_[41711]_ ;
  assign \new_[41715]_  = ~A267 & A266;
  assign \new_[41718]_  = A301 & ~A268;
  assign \new_[41719]_  = \new_[41718]_  & \new_[41715]_ ;
  assign \new_[41720]_  = \new_[41719]_  & \new_[41712]_ ;
  assign \new_[41724]_  = A166 & ~A167;
  assign \new_[41725]_  = A170 & \new_[41724]_ ;
  assign \new_[41728]_  = ~A200 & ~A199;
  assign \new_[41731]_  = ~A232 & ~A202;
  assign \new_[41732]_  = \new_[41731]_  & \new_[41728]_ ;
  assign \new_[41733]_  = \new_[41732]_  & \new_[41725]_ ;
  assign \new_[41737]_  = ~A265 & ~A235;
  assign \new_[41738]_  = ~A233 & \new_[41737]_ ;
  assign \new_[41741]_  = ~A268 & ~A266;
  assign \new_[41744]_  = A300 & A299;
  assign \new_[41745]_  = \new_[41744]_  & \new_[41741]_ ;
  assign \new_[41746]_  = \new_[41745]_  & \new_[41738]_ ;
  assign \new_[41750]_  = A166 & ~A167;
  assign \new_[41751]_  = A170 & \new_[41750]_ ;
  assign \new_[41754]_  = ~A200 & ~A199;
  assign \new_[41757]_  = ~A232 & ~A202;
  assign \new_[41758]_  = \new_[41757]_  & \new_[41754]_ ;
  assign \new_[41759]_  = \new_[41758]_  & \new_[41751]_ ;
  assign \new_[41763]_  = ~A265 & ~A235;
  assign \new_[41764]_  = ~A233 & \new_[41763]_ ;
  assign \new_[41767]_  = ~A268 & ~A266;
  assign \new_[41770]_  = A300 & A298;
  assign \new_[41771]_  = \new_[41770]_  & \new_[41767]_ ;
  assign \new_[41772]_  = \new_[41771]_  & \new_[41764]_ ;
  assign \new_[41776]_  = ~A202 & ~A201;
  assign \new_[41777]_  = A169 & \new_[41776]_ ;
  assign \new_[41780]_  = ~A234 & ~A203;
  assign \new_[41783]_  = ~A236 & ~A235;
  assign \new_[41784]_  = \new_[41783]_  & \new_[41780]_ ;
  assign \new_[41785]_  = \new_[41784]_  & \new_[41777]_ ;
  assign \new_[41789]_  = ~A267 & A266;
  assign \new_[41790]_  = A265 & \new_[41789]_ ;
  assign \new_[41793]_  = A298 & ~A268;
  assign \new_[41796]_  = A302 & ~A299;
  assign \new_[41797]_  = \new_[41796]_  & \new_[41793]_ ;
  assign \new_[41798]_  = \new_[41797]_  & \new_[41790]_ ;
  assign \new_[41802]_  = ~A202 & ~A201;
  assign \new_[41803]_  = A169 & \new_[41802]_ ;
  assign \new_[41806]_  = ~A234 & ~A203;
  assign \new_[41809]_  = ~A236 & ~A235;
  assign \new_[41810]_  = \new_[41809]_  & \new_[41806]_ ;
  assign \new_[41811]_  = \new_[41810]_  & \new_[41803]_ ;
  assign \new_[41815]_  = ~A267 & A266;
  assign \new_[41816]_  = A265 & \new_[41815]_ ;
  assign \new_[41819]_  = ~A298 & ~A268;
  assign \new_[41822]_  = A302 & A299;
  assign \new_[41823]_  = \new_[41822]_  & \new_[41819]_ ;
  assign \new_[41824]_  = \new_[41823]_  & \new_[41816]_ ;
  assign \new_[41828]_  = ~A202 & ~A201;
  assign \new_[41829]_  = A169 & \new_[41828]_ ;
  assign \new_[41832]_  = A232 & ~A203;
  assign \new_[41835]_  = ~A234 & A233;
  assign \new_[41836]_  = \new_[41835]_  & \new_[41832]_ ;
  assign \new_[41837]_  = \new_[41836]_  & \new_[41829]_ ;
  assign \new_[41841]_  = ~A268 & ~A267;
  assign \new_[41842]_  = ~A235 & \new_[41841]_ ;
  assign \new_[41845]_  = A298 & ~A269;
  assign \new_[41848]_  = A302 & ~A299;
  assign \new_[41849]_  = \new_[41848]_  & \new_[41845]_ ;
  assign \new_[41850]_  = \new_[41849]_  & \new_[41842]_ ;
  assign \new_[41854]_  = ~A202 & ~A201;
  assign \new_[41855]_  = A169 & \new_[41854]_ ;
  assign \new_[41858]_  = A232 & ~A203;
  assign \new_[41861]_  = ~A234 & A233;
  assign \new_[41862]_  = \new_[41861]_  & \new_[41858]_ ;
  assign \new_[41863]_  = \new_[41862]_  & \new_[41855]_ ;
  assign \new_[41867]_  = ~A268 & ~A267;
  assign \new_[41868]_  = ~A235 & \new_[41867]_ ;
  assign \new_[41871]_  = ~A298 & ~A269;
  assign \new_[41874]_  = A302 & A299;
  assign \new_[41875]_  = \new_[41874]_  & \new_[41871]_ ;
  assign \new_[41876]_  = \new_[41875]_  & \new_[41868]_ ;
  assign \new_[41880]_  = ~A202 & ~A201;
  assign \new_[41881]_  = A169 & \new_[41880]_ ;
  assign \new_[41884]_  = A232 & ~A203;
  assign \new_[41887]_  = ~A234 & A233;
  assign \new_[41888]_  = \new_[41887]_  & \new_[41884]_ ;
  assign \new_[41889]_  = \new_[41888]_  & \new_[41881]_ ;
  assign \new_[41893]_  = A266 & A265;
  assign \new_[41894]_  = ~A235 & \new_[41893]_ ;
  assign \new_[41897]_  = ~A268 & ~A267;
  assign \new_[41900]_  = A300 & A299;
  assign \new_[41901]_  = \new_[41900]_  & \new_[41897]_ ;
  assign \new_[41902]_  = \new_[41901]_  & \new_[41894]_ ;
  assign \new_[41906]_  = ~A202 & ~A201;
  assign \new_[41907]_  = A169 & \new_[41906]_ ;
  assign \new_[41910]_  = A232 & ~A203;
  assign \new_[41913]_  = ~A234 & A233;
  assign \new_[41914]_  = \new_[41913]_  & \new_[41910]_ ;
  assign \new_[41915]_  = \new_[41914]_  & \new_[41907]_ ;
  assign \new_[41919]_  = A266 & A265;
  assign \new_[41920]_  = ~A235 & \new_[41919]_ ;
  assign \new_[41923]_  = ~A268 & ~A267;
  assign \new_[41926]_  = A300 & A298;
  assign \new_[41927]_  = \new_[41926]_  & \new_[41923]_ ;
  assign \new_[41928]_  = \new_[41927]_  & \new_[41920]_ ;
  assign \new_[41932]_  = ~A202 & ~A201;
  assign \new_[41933]_  = A169 & \new_[41932]_ ;
  assign \new_[41936]_  = A232 & ~A203;
  assign \new_[41939]_  = ~A234 & A233;
  assign \new_[41940]_  = \new_[41939]_  & \new_[41936]_ ;
  assign \new_[41941]_  = \new_[41940]_  & \new_[41933]_ ;
  assign \new_[41945]_  = ~A266 & ~A265;
  assign \new_[41946]_  = ~A235 & \new_[41945]_ ;
  assign \new_[41949]_  = A298 & ~A268;
  assign \new_[41952]_  = A302 & ~A299;
  assign \new_[41953]_  = \new_[41952]_  & \new_[41949]_ ;
  assign \new_[41954]_  = \new_[41953]_  & \new_[41946]_ ;
  assign \new_[41958]_  = ~A202 & ~A201;
  assign \new_[41959]_  = A169 & \new_[41958]_ ;
  assign \new_[41962]_  = A232 & ~A203;
  assign \new_[41965]_  = ~A234 & A233;
  assign \new_[41966]_  = \new_[41965]_  & \new_[41962]_ ;
  assign \new_[41967]_  = \new_[41966]_  & \new_[41959]_ ;
  assign \new_[41971]_  = ~A266 & ~A265;
  assign \new_[41972]_  = ~A235 & \new_[41971]_ ;
  assign \new_[41975]_  = ~A298 & ~A268;
  assign \new_[41978]_  = A302 & A299;
  assign \new_[41979]_  = \new_[41978]_  & \new_[41975]_ ;
  assign \new_[41980]_  = \new_[41979]_  & \new_[41972]_ ;
  assign \new_[41984]_  = ~A202 & ~A201;
  assign \new_[41985]_  = A169 & \new_[41984]_ ;
  assign \new_[41988]_  = ~A232 & ~A203;
  assign \new_[41991]_  = ~A235 & ~A233;
  assign \new_[41992]_  = \new_[41991]_  & \new_[41988]_ ;
  assign \new_[41993]_  = \new_[41992]_  & \new_[41985]_ ;
  assign \new_[41997]_  = ~A267 & A266;
  assign \new_[41998]_  = A265 & \new_[41997]_ ;
  assign \new_[42001]_  = A298 & ~A268;
  assign \new_[42004]_  = A302 & ~A299;
  assign \new_[42005]_  = \new_[42004]_  & \new_[42001]_ ;
  assign \new_[42006]_  = \new_[42005]_  & \new_[41998]_ ;
  assign \new_[42010]_  = ~A202 & ~A201;
  assign \new_[42011]_  = A169 & \new_[42010]_ ;
  assign \new_[42014]_  = ~A232 & ~A203;
  assign \new_[42017]_  = ~A235 & ~A233;
  assign \new_[42018]_  = \new_[42017]_  & \new_[42014]_ ;
  assign \new_[42019]_  = \new_[42018]_  & \new_[42011]_ ;
  assign \new_[42023]_  = ~A267 & A266;
  assign \new_[42024]_  = A265 & \new_[42023]_ ;
  assign \new_[42027]_  = ~A298 & ~A268;
  assign \new_[42030]_  = A302 & A299;
  assign \new_[42031]_  = \new_[42030]_  & \new_[42027]_ ;
  assign \new_[42032]_  = \new_[42031]_  & \new_[42024]_ ;
  assign \new_[42036]_  = A200 & A199;
  assign \new_[42037]_  = A169 & \new_[42036]_ ;
  assign \new_[42040]_  = ~A202 & ~A201;
  assign \new_[42043]_  = ~A235 & ~A234;
  assign \new_[42044]_  = \new_[42043]_  & \new_[42040]_ ;
  assign \new_[42045]_  = \new_[42044]_  & \new_[42037]_ ;
  assign \new_[42049]_  = ~A268 & ~A267;
  assign \new_[42050]_  = ~A236 & \new_[42049]_ ;
  assign \new_[42053]_  = A298 & ~A269;
  assign \new_[42056]_  = A302 & ~A299;
  assign \new_[42057]_  = \new_[42056]_  & \new_[42053]_ ;
  assign \new_[42058]_  = \new_[42057]_  & \new_[42050]_ ;
  assign \new_[42062]_  = A200 & A199;
  assign \new_[42063]_  = A169 & \new_[42062]_ ;
  assign \new_[42066]_  = ~A202 & ~A201;
  assign \new_[42069]_  = ~A235 & ~A234;
  assign \new_[42070]_  = \new_[42069]_  & \new_[42066]_ ;
  assign \new_[42071]_  = \new_[42070]_  & \new_[42063]_ ;
  assign \new_[42075]_  = ~A268 & ~A267;
  assign \new_[42076]_  = ~A236 & \new_[42075]_ ;
  assign \new_[42079]_  = ~A298 & ~A269;
  assign \new_[42082]_  = A302 & A299;
  assign \new_[42083]_  = \new_[42082]_  & \new_[42079]_ ;
  assign \new_[42084]_  = \new_[42083]_  & \new_[42076]_ ;
  assign \new_[42088]_  = A200 & A199;
  assign \new_[42089]_  = A169 & \new_[42088]_ ;
  assign \new_[42092]_  = ~A202 & ~A201;
  assign \new_[42095]_  = ~A235 & ~A234;
  assign \new_[42096]_  = \new_[42095]_  & \new_[42092]_ ;
  assign \new_[42097]_  = \new_[42096]_  & \new_[42089]_ ;
  assign \new_[42101]_  = A266 & A265;
  assign \new_[42102]_  = ~A236 & \new_[42101]_ ;
  assign \new_[42105]_  = ~A268 & ~A267;
  assign \new_[42108]_  = A300 & A299;
  assign \new_[42109]_  = \new_[42108]_  & \new_[42105]_ ;
  assign \new_[42110]_  = \new_[42109]_  & \new_[42102]_ ;
  assign \new_[42114]_  = A200 & A199;
  assign \new_[42115]_  = A169 & \new_[42114]_ ;
  assign \new_[42118]_  = ~A202 & ~A201;
  assign \new_[42121]_  = ~A235 & ~A234;
  assign \new_[42122]_  = \new_[42121]_  & \new_[42118]_ ;
  assign \new_[42123]_  = \new_[42122]_  & \new_[42115]_ ;
  assign \new_[42127]_  = A266 & A265;
  assign \new_[42128]_  = ~A236 & \new_[42127]_ ;
  assign \new_[42131]_  = ~A268 & ~A267;
  assign \new_[42134]_  = A300 & A298;
  assign \new_[42135]_  = \new_[42134]_  & \new_[42131]_ ;
  assign \new_[42136]_  = \new_[42135]_  & \new_[42128]_ ;
  assign \new_[42140]_  = A200 & A199;
  assign \new_[42141]_  = A169 & \new_[42140]_ ;
  assign \new_[42144]_  = ~A202 & ~A201;
  assign \new_[42147]_  = ~A235 & ~A234;
  assign \new_[42148]_  = \new_[42147]_  & \new_[42144]_ ;
  assign \new_[42149]_  = \new_[42148]_  & \new_[42141]_ ;
  assign \new_[42153]_  = ~A266 & ~A265;
  assign \new_[42154]_  = ~A236 & \new_[42153]_ ;
  assign \new_[42157]_  = A298 & ~A268;
  assign \new_[42160]_  = A302 & ~A299;
  assign \new_[42161]_  = \new_[42160]_  & \new_[42157]_ ;
  assign \new_[42162]_  = \new_[42161]_  & \new_[42154]_ ;
  assign \new_[42166]_  = A200 & A199;
  assign \new_[42167]_  = A169 & \new_[42166]_ ;
  assign \new_[42170]_  = ~A202 & ~A201;
  assign \new_[42173]_  = ~A235 & ~A234;
  assign \new_[42174]_  = \new_[42173]_  & \new_[42170]_ ;
  assign \new_[42175]_  = \new_[42174]_  & \new_[42167]_ ;
  assign \new_[42179]_  = ~A266 & ~A265;
  assign \new_[42180]_  = ~A236 & \new_[42179]_ ;
  assign \new_[42183]_  = ~A298 & ~A268;
  assign \new_[42186]_  = A302 & A299;
  assign \new_[42187]_  = \new_[42186]_  & \new_[42183]_ ;
  assign \new_[42188]_  = \new_[42187]_  & \new_[42180]_ ;
  assign \new_[42192]_  = A200 & A199;
  assign \new_[42193]_  = A169 & \new_[42192]_ ;
  assign \new_[42196]_  = ~A202 & ~A201;
  assign \new_[42199]_  = A233 & A232;
  assign \new_[42200]_  = \new_[42199]_  & \new_[42196]_ ;
  assign \new_[42201]_  = \new_[42200]_  & \new_[42193]_ ;
  assign \new_[42205]_  = ~A267 & ~A235;
  assign \new_[42206]_  = ~A234 & \new_[42205]_ ;
  assign \new_[42209]_  = ~A269 & ~A268;
  assign \new_[42212]_  = A300 & A299;
  assign \new_[42213]_  = \new_[42212]_  & \new_[42209]_ ;
  assign \new_[42214]_  = \new_[42213]_  & \new_[42206]_ ;
  assign \new_[42218]_  = A200 & A199;
  assign \new_[42219]_  = A169 & \new_[42218]_ ;
  assign \new_[42222]_  = ~A202 & ~A201;
  assign \new_[42225]_  = A233 & A232;
  assign \new_[42226]_  = \new_[42225]_  & \new_[42222]_ ;
  assign \new_[42227]_  = \new_[42226]_  & \new_[42219]_ ;
  assign \new_[42231]_  = ~A267 & ~A235;
  assign \new_[42232]_  = ~A234 & \new_[42231]_ ;
  assign \new_[42235]_  = ~A269 & ~A268;
  assign \new_[42238]_  = A300 & A298;
  assign \new_[42239]_  = \new_[42238]_  & \new_[42235]_ ;
  assign \new_[42240]_  = \new_[42239]_  & \new_[42232]_ ;
  assign \new_[42244]_  = A200 & A199;
  assign \new_[42245]_  = A169 & \new_[42244]_ ;
  assign \new_[42248]_  = ~A202 & ~A201;
  assign \new_[42251]_  = A233 & A232;
  assign \new_[42252]_  = \new_[42251]_  & \new_[42248]_ ;
  assign \new_[42253]_  = \new_[42252]_  & \new_[42245]_ ;
  assign \new_[42257]_  = A265 & ~A235;
  assign \new_[42258]_  = ~A234 & \new_[42257]_ ;
  assign \new_[42261]_  = ~A267 & A266;
  assign \new_[42264]_  = A301 & ~A268;
  assign \new_[42265]_  = \new_[42264]_  & \new_[42261]_ ;
  assign \new_[42266]_  = \new_[42265]_  & \new_[42258]_ ;
  assign \new_[42270]_  = A200 & A199;
  assign \new_[42271]_  = A169 & \new_[42270]_ ;
  assign \new_[42274]_  = ~A202 & ~A201;
  assign \new_[42277]_  = A233 & A232;
  assign \new_[42278]_  = \new_[42277]_  & \new_[42274]_ ;
  assign \new_[42279]_  = \new_[42278]_  & \new_[42271]_ ;
  assign \new_[42283]_  = ~A265 & ~A235;
  assign \new_[42284]_  = ~A234 & \new_[42283]_ ;
  assign \new_[42287]_  = ~A268 & ~A266;
  assign \new_[42290]_  = A300 & A299;
  assign \new_[42291]_  = \new_[42290]_  & \new_[42287]_ ;
  assign \new_[42292]_  = \new_[42291]_  & \new_[42284]_ ;
  assign \new_[42296]_  = A200 & A199;
  assign \new_[42297]_  = A169 & \new_[42296]_ ;
  assign \new_[42300]_  = ~A202 & ~A201;
  assign \new_[42303]_  = A233 & A232;
  assign \new_[42304]_  = \new_[42303]_  & \new_[42300]_ ;
  assign \new_[42305]_  = \new_[42304]_  & \new_[42297]_ ;
  assign \new_[42309]_  = ~A265 & ~A235;
  assign \new_[42310]_  = ~A234 & \new_[42309]_ ;
  assign \new_[42313]_  = ~A268 & ~A266;
  assign \new_[42316]_  = A300 & A298;
  assign \new_[42317]_  = \new_[42316]_  & \new_[42313]_ ;
  assign \new_[42318]_  = \new_[42317]_  & \new_[42310]_ ;
  assign \new_[42322]_  = A200 & A199;
  assign \new_[42323]_  = A169 & \new_[42322]_ ;
  assign \new_[42326]_  = ~A202 & ~A201;
  assign \new_[42329]_  = ~A233 & ~A232;
  assign \new_[42330]_  = \new_[42329]_  & \new_[42326]_ ;
  assign \new_[42331]_  = \new_[42330]_  & \new_[42323]_ ;
  assign \new_[42335]_  = ~A268 & ~A267;
  assign \new_[42336]_  = ~A235 & \new_[42335]_ ;
  assign \new_[42339]_  = A298 & ~A269;
  assign \new_[42342]_  = A302 & ~A299;
  assign \new_[42343]_  = \new_[42342]_  & \new_[42339]_ ;
  assign \new_[42344]_  = \new_[42343]_  & \new_[42336]_ ;
  assign \new_[42348]_  = A200 & A199;
  assign \new_[42349]_  = A169 & \new_[42348]_ ;
  assign \new_[42352]_  = ~A202 & ~A201;
  assign \new_[42355]_  = ~A233 & ~A232;
  assign \new_[42356]_  = \new_[42355]_  & \new_[42352]_ ;
  assign \new_[42357]_  = \new_[42356]_  & \new_[42349]_ ;
  assign \new_[42361]_  = ~A268 & ~A267;
  assign \new_[42362]_  = ~A235 & \new_[42361]_ ;
  assign \new_[42365]_  = ~A298 & ~A269;
  assign \new_[42368]_  = A302 & A299;
  assign \new_[42369]_  = \new_[42368]_  & \new_[42365]_ ;
  assign \new_[42370]_  = \new_[42369]_  & \new_[42362]_ ;
  assign \new_[42374]_  = A200 & A199;
  assign \new_[42375]_  = A169 & \new_[42374]_ ;
  assign \new_[42378]_  = ~A202 & ~A201;
  assign \new_[42381]_  = ~A233 & ~A232;
  assign \new_[42382]_  = \new_[42381]_  & \new_[42378]_ ;
  assign \new_[42383]_  = \new_[42382]_  & \new_[42375]_ ;
  assign \new_[42387]_  = A266 & A265;
  assign \new_[42388]_  = ~A235 & \new_[42387]_ ;
  assign \new_[42391]_  = ~A268 & ~A267;
  assign \new_[42394]_  = A300 & A299;
  assign \new_[42395]_  = \new_[42394]_  & \new_[42391]_ ;
  assign \new_[42396]_  = \new_[42395]_  & \new_[42388]_ ;
  assign \new_[42400]_  = A200 & A199;
  assign \new_[42401]_  = A169 & \new_[42400]_ ;
  assign \new_[42404]_  = ~A202 & ~A201;
  assign \new_[42407]_  = ~A233 & ~A232;
  assign \new_[42408]_  = \new_[42407]_  & \new_[42404]_ ;
  assign \new_[42409]_  = \new_[42408]_  & \new_[42401]_ ;
  assign \new_[42413]_  = A266 & A265;
  assign \new_[42414]_  = ~A235 & \new_[42413]_ ;
  assign \new_[42417]_  = ~A268 & ~A267;
  assign \new_[42420]_  = A300 & A298;
  assign \new_[42421]_  = \new_[42420]_  & \new_[42417]_ ;
  assign \new_[42422]_  = \new_[42421]_  & \new_[42414]_ ;
  assign \new_[42426]_  = A200 & A199;
  assign \new_[42427]_  = A169 & \new_[42426]_ ;
  assign \new_[42430]_  = ~A202 & ~A201;
  assign \new_[42433]_  = ~A233 & ~A232;
  assign \new_[42434]_  = \new_[42433]_  & \new_[42430]_ ;
  assign \new_[42435]_  = \new_[42434]_  & \new_[42427]_ ;
  assign \new_[42439]_  = ~A266 & ~A265;
  assign \new_[42440]_  = ~A235 & \new_[42439]_ ;
  assign \new_[42443]_  = A298 & ~A268;
  assign \new_[42446]_  = A302 & ~A299;
  assign \new_[42447]_  = \new_[42446]_  & \new_[42443]_ ;
  assign \new_[42448]_  = \new_[42447]_  & \new_[42440]_ ;
  assign \new_[42452]_  = A200 & A199;
  assign \new_[42453]_  = A169 & \new_[42452]_ ;
  assign \new_[42456]_  = ~A202 & ~A201;
  assign \new_[42459]_  = ~A233 & ~A232;
  assign \new_[42460]_  = \new_[42459]_  & \new_[42456]_ ;
  assign \new_[42461]_  = \new_[42460]_  & \new_[42453]_ ;
  assign \new_[42465]_  = ~A266 & ~A265;
  assign \new_[42466]_  = ~A235 & \new_[42465]_ ;
  assign \new_[42469]_  = ~A298 & ~A268;
  assign \new_[42472]_  = A302 & A299;
  assign \new_[42473]_  = \new_[42472]_  & \new_[42469]_ ;
  assign \new_[42474]_  = \new_[42473]_  & \new_[42466]_ ;
  assign \new_[42478]_  = ~A200 & ~A199;
  assign \new_[42479]_  = A169 & \new_[42478]_ ;
  assign \new_[42482]_  = ~A234 & ~A202;
  assign \new_[42485]_  = ~A236 & ~A235;
  assign \new_[42486]_  = \new_[42485]_  & \new_[42482]_ ;
  assign \new_[42487]_  = \new_[42486]_  & \new_[42479]_ ;
  assign \new_[42491]_  = ~A267 & A266;
  assign \new_[42492]_  = A265 & \new_[42491]_ ;
  assign \new_[42495]_  = A298 & ~A268;
  assign \new_[42498]_  = A302 & ~A299;
  assign \new_[42499]_  = \new_[42498]_  & \new_[42495]_ ;
  assign \new_[42500]_  = \new_[42499]_  & \new_[42492]_ ;
  assign \new_[42504]_  = ~A200 & ~A199;
  assign \new_[42505]_  = A169 & \new_[42504]_ ;
  assign \new_[42508]_  = ~A234 & ~A202;
  assign \new_[42511]_  = ~A236 & ~A235;
  assign \new_[42512]_  = \new_[42511]_  & \new_[42508]_ ;
  assign \new_[42513]_  = \new_[42512]_  & \new_[42505]_ ;
  assign \new_[42517]_  = ~A267 & A266;
  assign \new_[42518]_  = A265 & \new_[42517]_ ;
  assign \new_[42521]_  = ~A298 & ~A268;
  assign \new_[42524]_  = A302 & A299;
  assign \new_[42525]_  = \new_[42524]_  & \new_[42521]_ ;
  assign \new_[42526]_  = \new_[42525]_  & \new_[42518]_ ;
  assign \new_[42530]_  = ~A200 & ~A199;
  assign \new_[42531]_  = A169 & \new_[42530]_ ;
  assign \new_[42534]_  = A232 & ~A202;
  assign \new_[42537]_  = ~A234 & A233;
  assign \new_[42538]_  = \new_[42537]_  & \new_[42534]_ ;
  assign \new_[42539]_  = \new_[42538]_  & \new_[42531]_ ;
  assign \new_[42543]_  = ~A268 & ~A267;
  assign \new_[42544]_  = ~A235 & \new_[42543]_ ;
  assign \new_[42547]_  = A298 & ~A269;
  assign \new_[42550]_  = A302 & ~A299;
  assign \new_[42551]_  = \new_[42550]_  & \new_[42547]_ ;
  assign \new_[42552]_  = \new_[42551]_  & \new_[42544]_ ;
  assign \new_[42556]_  = ~A200 & ~A199;
  assign \new_[42557]_  = A169 & \new_[42556]_ ;
  assign \new_[42560]_  = A232 & ~A202;
  assign \new_[42563]_  = ~A234 & A233;
  assign \new_[42564]_  = \new_[42563]_  & \new_[42560]_ ;
  assign \new_[42565]_  = \new_[42564]_  & \new_[42557]_ ;
  assign \new_[42569]_  = ~A268 & ~A267;
  assign \new_[42570]_  = ~A235 & \new_[42569]_ ;
  assign \new_[42573]_  = ~A298 & ~A269;
  assign \new_[42576]_  = A302 & A299;
  assign \new_[42577]_  = \new_[42576]_  & \new_[42573]_ ;
  assign \new_[42578]_  = \new_[42577]_  & \new_[42570]_ ;
  assign \new_[42582]_  = ~A200 & ~A199;
  assign \new_[42583]_  = A169 & \new_[42582]_ ;
  assign \new_[42586]_  = A232 & ~A202;
  assign \new_[42589]_  = ~A234 & A233;
  assign \new_[42590]_  = \new_[42589]_  & \new_[42586]_ ;
  assign \new_[42591]_  = \new_[42590]_  & \new_[42583]_ ;
  assign \new_[42595]_  = A266 & A265;
  assign \new_[42596]_  = ~A235 & \new_[42595]_ ;
  assign \new_[42599]_  = ~A268 & ~A267;
  assign \new_[42602]_  = A300 & A299;
  assign \new_[42603]_  = \new_[42602]_  & \new_[42599]_ ;
  assign \new_[42604]_  = \new_[42603]_  & \new_[42596]_ ;
  assign \new_[42608]_  = ~A200 & ~A199;
  assign \new_[42609]_  = A169 & \new_[42608]_ ;
  assign \new_[42612]_  = A232 & ~A202;
  assign \new_[42615]_  = ~A234 & A233;
  assign \new_[42616]_  = \new_[42615]_  & \new_[42612]_ ;
  assign \new_[42617]_  = \new_[42616]_  & \new_[42609]_ ;
  assign \new_[42621]_  = A266 & A265;
  assign \new_[42622]_  = ~A235 & \new_[42621]_ ;
  assign \new_[42625]_  = ~A268 & ~A267;
  assign \new_[42628]_  = A300 & A298;
  assign \new_[42629]_  = \new_[42628]_  & \new_[42625]_ ;
  assign \new_[42630]_  = \new_[42629]_  & \new_[42622]_ ;
  assign \new_[42634]_  = ~A200 & ~A199;
  assign \new_[42635]_  = A169 & \new_[42634]_ ;
  assign \new_[42638]_  = A232 & ~A202;
  assign \new_[42641]_  = ~A234 & A233;
  assign \new_[42642]_  = \new_[42641]_  & \new_[42638]_ ;
  assign \new_[42643]_  = \new_[42642]_  & \new_[42635]_ ;
  assign \new_[42647]_  = ~A266 & ~A265;
  assign \new_[42648]_  = ~A235 & \new_[42647]_ ;
  assign \new_[42651]_  = A298 & ~A268;
  assign \new_[42654]_  = A302 & ~A299;
  assign \new_[42655]_  = \new_[42654]_  & \new_[42651]_ ;
  assign \new_[42656]_  = \new_[42655]_  & \new_[42648]_ ;
  assign \new_[42660]_  = ~A200 & ~A199;
  assign \new_[42661]_  = A169 & \new_[42660]_ ;
  assign \new_[42664]_  = A232 & ~A202;
  assign \new_[42667]_  = ~A234 & A233;
  assign \new_[42668]_  = \new_[42667]_  & \new_[42664]_ ;
  assign \new_[42669]_  = \new_[42668]_  & \new_[42661]_ ;
  assign \new_[42673]_  = ~A266 & ~A265;
  assign \new_[42674]_  = ~A235 & \new_[42673]_ ;
  assign \new_[42677]_  = ~A298 & ~A268;
  assign \new_[42680]_  = A302 & A299;
  assign \new_[42681]_  = \new_[42680]_  & \new_[42677]_ ;
  assign \new_[42682]_  = \new_[42681]_  & \new_[42674]_ ;
  assign \new_[42686]_  = ~A200 & ~A199;
  assign \new_[42687]_  = A169 & \new_[42686]_ ;
  assign \new_[42690]_  = ~A232 & ~A202;
  assign \new_[42693]_  = ~A235 & ~A233;
  assign \new_[42694]_  = \new_[42693]_  & \new_[42690]_ ;
  assign \new_[42695]_  = \new_[42694]_  & \new_[42687]_ ;
  assign \new_[42699]_  = ~A267 & A266;
  assign \new_[42700]_  = A265 & \new_[42699]_ ;
  assign \new_[42703]_  = A298 & ~A268;
  assign \new_[42706]_  = A302 & ~A299;
  assign \new_[42707]_  = \new_[42706]_  & \new_[42703]_ ;
  assign \new_[42708]_  = \new_[42707]_  & \new_[42700]_ ;
  assign \new_[42712]_  = ~A200 & ~A199;
  assign \new_[42713]_  = A169 & \new_[42712]_ ;
  assign \new_[42716]_  = ~A232 & ~A202;
  assign \new_[42719]_  = ~A235 & ~A233;
  assign \new_[42720]_  = \new_[42719]_  & \new_[42716]_ ;
  assign \new_[42721]_  = \new_[42720]_  & \new_[42713]_ ;
  assign \new_[42725]_  = ~A267 & A266;
  assign \new_[42726]_  = A265 & \new_[42725]_ ;
  assign \new_[42729]_  = ~A298 & ~A268;
  assign \new_[42732]_  = A302 & A299;
  assign \new_[42733]_  = \new_[42732]_  & \new_[42729]_ ;
  assign \new_[42734]_  = \new_[42733]_  & \new_[42726]_ ;
  assign \new_[42738]_  = ~A166 & ~A167;
  assign \new_[42739]_  = ~A169 & \new_[42738]_ ;
  assign \new_[42742]_  = ~A234 & A202;
  assign \new_[42745]_  = ~A236 & ~A235;
  assign \new_[42746]_  = \new_[42745]_  & \new_[42742]_ ;
  assign \new_[42747]_  = \new_[42746]_  & \new_[42739]_ ;
  assign \new_[42751]_  = ~A267 & A266;
  assign \new_[42752]_  = A265 & \new_[42751]_ ;
  assign \new_[42755]_  = A298 & ~A268;
  assign \new_[42758]_  = A302 & ~A299;
  assign \new_[42759]_  = \new_[42758]_  & \new_[42755]_ ;
  assign \new_[42760]_  = \new_[42759]_  & \new_[42752]_ ;
  assign \new_[42764]_  = ~A166 & ~A167;
  assign \new_[42765]_  = ~A169 & \new_[42764]_ ;
  assign \new_[42768]_  = ~A234 & A202;
  assign \new_[42771]_  = ~A236 & ~A235;
  assign \new_[42772]_  = \new_[42771]_  & \new_[42768]_ ;
  assign \new_[42773]_  = \new_[42772]_  & \new_[42765]_ ;
  assign \new_[42777]_  = ~A267 & A266;
  assign \new_[42778]_  = A265 & \new_[42777]_ ;
  assign \new_[42781]_  = ~A298 & ~A268;
  assign \new_[42784]_  = A302 & A299;
  assign \new_[42785]_  = \new_[42784]_  & \new_[42781]_ ;
  assign \new_[42786]_  = \new_[42785]_  & \new_[42778]_ ;
  assign \new_[42790]_  = ~A166 & ~A167;
  assign \new_[42791]_  = ~A169 & \new_[42790]_ ;
  assign \new_[42794]_  = A232 & A202;
  assign \new_[42797]_  = ~A234 & A233;
  assign \new_[42798]_  = \new_[42797]_  & \new_[42794]_ ;
  assign \new_[42799]_  = \new_[42798]_  & \new_[42791]_ ;
  assign \new_[42803]_  = ~A268 & ~A267;
  assign \new_[42804]_  = ~A235 & \new_[42803]_ ;
  assign \new_[42807]_  = A298 & ~A269;
  assign \new_[42810]_  = A302 & ~A299;
  assign \new_[42811]_  = \new_[42810]_  & \new_[42807]_ ;
  assign \new_[42812]_  = \new_[42811]_  & \new_[42804]_ ;
  assign \new_[42816]_  = ~A166 & ~A167;
  assign \new_[42817]_  = ~A169 & \new_[42816]_ ;
  assign \new_[42820]_  = A232 & A202;
  assign \new_[42823]_  = ~A234 & A233;
  assign \new_[42824]_  = \new_[42823]_  & \new_[42820]_ ;
  assign \new_[42825]_  = \new_[42824]_  & \new_[42817]_ ;
  assign \new_[42829]_  = ~A268 & ~A267;
  assign \new_[42830]_  = ~A235 & \new_[42829]_ ;
  assign \new_[42833]_  = ~A298 & ~A269;
  assign \new_[42836]_  = A302 & A299;
  assign \new_[42837]_  = \new_[42836]_  & \new_[42833]_ ;
  assign \new_[42838]_  = \new_[42837]_  & \new_[42830]_ ;
  assign \new_[42842]_  = ~A166 & ~A167;
  assign \new_[42843]_  = ~A169 & \new_[42842]_ ;
  assign \new_[42846]_  = A232 & A202;
  assign \new_[42849]_  = ~A234 & A233;
  assign \new_[42850]_  = \new_[42849]_  & \new_[42846]_ ;
  assign \new_[42851]_  = \new_[42850]_  & \new_[42843]_ ;
  assign \new_[42855]_  = A266 & A265;
  assign \new_[42856]_  = ~A235 & \new_[42855]_ ;
  assign \new_[42859]_  = ~A268 & ~A267;
  assign \new_[42862]_  = A300 & A299;
  assign \new_[42863]_  = \new_[42862]_  & \new_[42859]_ ;
  assign \new_[42864]_  = \new_[42863]_  & \new_[42856]_ ;
  assign \new_[42868]_  = ~A166 & ~A167;
  assign \new_[42869]_  = ~A169 & \new_[42868]_ ;
  assign \new_[42872]_  = A232 & A202;
  assign \new_[42875]_  = ~A234 & A233;
  assign \new_[42876]_  = \new_[42875]_  & \new_[42872]_ ;
  assign \new_[42877]_  = \new_[42876]_  & \new_[42869]_ ;
  assign \new_[42881]_  = A266 & A265;
  assign \new_[42882]_  = ~A235 & \new_[42881]_ ;
  assign \new_[42885]_  = ~A268 & ~A267;
  assign \new_[42888]_  = A300 & A298;
  assign \new_[42889]_  = \new_[42888]_  & \new_[42885]_ ;
  assign \new_[42890]_  = \new_[42889]_  & \new_[42882]_ ;
  assign \new_[42894]_  = ~A166 & ~A167;
  assign \new_[42895]_  = ~A169 & \new_[42894]_ ;
  assign \new_[42898]_  = A232 & A202;
  assign \new_[42901]_  = ~A234 & A233;
  assign \new_[42902]_  = \new_[42901]_  & \new_[42898]_ ;
  assign \new_[42903]_  = \new_[42902]_  & \new_[42895]_ ;
  assign \new_[42907]_  = ~A266 & ~A265;
  assign \new_[42908]_  = ~A235 & \new_[42907]_ ;
  assign \new_[42911]_  = A298 & ~A268;
  assign \new_[42914]_  = A302 & ~A299;
  assign \new_[42915]_  = \new_[42914]_  & \new_[42911]_ ;
  assign \new_[42916]_  = \new_[42915]_  & \new_[42908]_ ;
  assign \new_[42920]_  = ~A166 & ~A167;
  assign \new_[42921]_  = ~A169 & \new_[42920]_ ;
  assign \new_[42924]_  = A232 & A202;
  assign \new_[42927]_  = ~A234 & A233;
  assign \new_[42928]_  = \new_[42927]_  & \new_[42924]_ ;
  assign \new_[42929]_  = \new_[42928]_  & \new_[42921]_ ;
  assign \new_[42933]_  = ~A266 & ~A265;
  assign \new_[42934]_  = ~A235 & \new_[42933]_ ;
  assign \new_[42937]_  = ~A298 & ~A268;
  assign \new_[42940]_  = A302 & A299;
  assign \new_[42941]_  = \new_[42940]_  & \new_[42937]_ ;
  assign \new_[42942]_  = \new_[42941]_  & \new_[42934]_ ;
  assign \new_[42946]_  = ~A166 & ~A167;
  assign \new_[42947]_  = ~A169 & \new_[42946]_ ;
  assign \new_[42950]_  = ~A232 & A202;
  assign \new_[42953]_  = ~A235 & ~A233;
  assign \new_[42954]_  = \new_[42953]_  & \new_[42950]_ ;
  assign \new_[42955]_  = \new_[42954]_  & \new_[42947]_ ;
  assign \new_[42959]_  = ~A267 & A266;
  assign \new_[42960]_  = A265 & \new_[42959]_ ;
  assign \new_[42963]_  = A298 & ~A268;
  assign \new_[42966]_  = A302 & ~A299;
  assign \new_[42967]_  = \new_[42966]_  & \new_[42963]_ ;
  assign \new_[42968]_  = \new_[42967]_  & \new_[42960]_ ;
  assign \new_[42972]_  = ~A166 & ~A167;
  assign \new_[42973]_  = ~A169 & \new_[42972]_ ;
  assign \new_[42976]_  = ~A232 & A202;
  assign \new_[42979]_  = ~A235 & ~A233;
  assign \new_[42980]_  = \new_[42979]_  & \new_[42976]_ ;
  assign \new_[42981]_  = \new_[42980]_  & \new_[42973]_ ;
  assign \new_[42985]_  = ~A267 & A266;
  assign \new_[42986]_  = A265 & \new_[42985]_ ;
  assign \new_[42989]_  = ~A298 & ~A268;
  assign \new_[42992]_  = A302 & A299;
  assign \new_[42993]_  = \new_[42992]_  & \new_[42989]_ ;
  assign \new_[42994]_  = \new_[42993]_  & \new_[42986]_ ;
  assign \new_[42998]_  = ~A166 & ~A167;
  assign \new_[42999]_  = ~A169 & \new_[42998]_ ;
  assign \new_[43002]_  = A201 & A199;
  assign \new_[43005]_  = ~A235 & ~A234;
  assign \new_[43006]_  = \new_[43005]_  & \new_[43002]_ ;
  assign \new_[43007]_  = \new_[43006]_  & \new_[42999]_ ;
  assign \new_[43011]_  = ~A268 & ~A267;
  assign \new_[43012]_  = ~A236 & \new_[43011]_ ;
  assign \new_[43015]_  = A298 & ~A269;
  assign \new_[43018]_  = A302 & ~A299;
  assign \new_[43019]_  = \new_[43018]_  & \new_[43015]_ ;
  assign \new_[43020]_  = \new_[43019]_  & \new_[43012]_ ;
  assign \new_[43024]_  = ~A166 & ~A167;
  assign \new_[43025]_  = ~A169 & \new_[43024]_ ;
  assign \new_[43028]_  = A201 & A199;
  assign \new_[43031]_  = ~A235 & ~A234;
  assign \new_[43032]_  = \new_[43031]_  & \new_[43028]_ ;
  assign \new_[43033]_  = \new_[43032]_  & \new_[43025]_ ;
  assign \new_[43037]_  = ~A268 & ~A267;
  assign \new_[43038]_  = ~A236 & \new_[43037]_ ;
  assign \new_[43041]_  = ~A298 & ~A269;
  assign \new_[43044]_  = A302 & A299;
  assign \new_[43045]_  = \new_[43044]_  & \new_[43041]_ ;
  assign \new_[43046]_  = \new_[43045]_  & \new_[43038]_ ;
  assign \new_[43050]_  = ~A166 & ~A167;
  assign \new_[43051]_  = ~A169 & \new_[43050]_ ;
  assign \new_[43054]_  = A201 & A199;
  assign \new_[43057]_  = ~A235 & ~A234;
  assign \new_[43058]_  = \new_[43057]_  & \new_[43054]_ ;
  assign \new_[43059]_  = \new_[43058]_  & \new_[43051]_ ;
  assign \new_[43063]_  = A266 & A265;
  assign \new_[43064]_  = ~A236 & \new_[43063]_ ;
  assign \new_[43067]_  = ~A268 & ~A267;
  assign \new_[43070]_  = A300 & A299;
  assign \new_[43071]_  = \new_[43070]_  & \new_[43067]_ ;
  assign \new_[43072]_  = \new_[43071]_  & \new_[43064]_ ;
  assign \new_[43076]_  = ~A166 & ~A167;
  assign \new_[43077]_  = ~A169 & \new_[43076]_ ;
  assign \new_[43080]_  = A201 & A199;
  assign \new_[43083]_  = ~A235 & ~A234;
  assign \new_[43084]_  = \new_[43083]_  & \new_[43080]_ ;
  assign \new_[43085]_  = \new_[43084]_  & \new_[43077]_ ;
  assign \new_[43089]_  = A266 & A265;
  assign \new_[43090]_  = ~A236 & \new_[43089]_ ;
  assign \new_[43093]_  = ~A268 & ~A267;
  assign \new_[43096]_  = A300 & A298;
  assign \new_[43097]_  = \new_[43096]_  & \new_[43093]_ ;
  assign \new_[43098]_  = \new_[43097]_  & \new_[43090]_ ;
  assign \new_[43102]_  = ~A166 & ~A167;
  assign \new_[43103]_  = ~A169 & \new_[43102]_ ;
  assign \new_[43106]_  = A201 & A199;
  assign \new_[43109]_  = ~A235 & ~A234;
  assign \new_[43110]_  = \new_[43109]_  & \new_[43106]_ ;
  assign \new_[43111]_  = \new_[43110]_  & \new_[43103]_ ;
  assign \new_[43115]_  = ~A266 & ~A265;
  assign \new_[43116]_  = ~A236 & \new_[43115]_ ;
  assign \new_[43119]_  = A298 & ~A268;
  assign \new_[43122]_  = A302 & ~A299;
  assign \new_[43123]_  = \new_[43122]_  & \new_[43119]_ ;
  assign \new_[43124]_  = \new_[43123]_  & \new_[43116]_ ;
  assign \new_[43128]_  = ~A166 & ~A167;
  assign \new_[43129]_  = ~A169 & \new_[43128]_ ;
  assign \new_[43132]_  = A201 & A199;
  assign \new_[43135]_  = ~A235 & ~A234;
  assign \new_[43136]_  = \new_[43135]_  & \new_[43132]_ ;
  assign \new_[43137]_  = \new_[43136]_  & \new_[43129]_ ;
  assign \new_[43141]_  = ~A266 & ~A265;
  assign \new_[43142]_  = ~A236 & \new_[43141]_ ;
  assign \new_[43145]_  = ~A298 & ~A268;
  assign \new_[43148]_  = A302 & A299;
  assign \new_[43149]_  = \new_[43148]_  & \new_[43145]_ ;
  assign \new_[43150]_  = \new_[43149]_  & \new_[43142]_ ;
  assign \new_[43154]_  = ~A166 & ~A167;
  assign \new_[43155]_  = ~A169 & \new_[43154]_ ;
  assign \new_[43158]_  = A201 & A199;
  assign \new_[43161]_  = A233 & A232;
  assign \new_[43162]_  = \new_[43161]_  & \new_[43158]_ ;
  assign \new_[43163]_  = \new_[43162]_  & \new_[43155]_ ;
  assign \new_[43167]_  = ~A267 & ~A235;
  assign \new_[43168]_  = ~A234 & \new_[43167]_ ;
  assign \new_[43171]_  = ~A269 & ~A268;
  assign \new_[43174]_  = A300 & A299;
  assign \new_[43175]_  = \new_[43174]_  & \new_[43171]_ ;
  assign \new_[43176]_  = \new_[43175]_  & \new_[43168]_ ;
  assign \new_[43180]_  = ~A166 & ~A167;
  assign \new_[43181]_  = ~A169 & \new_[43180]_ ;
  assign \new_[43184]_  = A201 & A199;
  assign \new_[43187]_  = A233 & A232;
  assign \new_[43188]_  = \new_[43187]_  & \new_[43184]_ ;
  assign \new_[43189]_  = \new_[43188]_  & \new_[43181]_ ;
  assign \new_[43193]_  = ~A267 & ~A235;
  assign \new_[43194]_  = ~A234 & \new_[43193]_ ;
  assign \new_[43197]_  = ~A269 & ~A268;
  assign \new_[43200]_  = A300 & A298;
  assign \new_[43201]_  = \new_[43200]_  & \new_[43197]_ ;
  assign \new_[43202]_  = \new_[43201]_  & \new_[43194]_ ;
  assign \new_[43206]_  = ~A166 & ~A167;
  assign \new_[43207]_  = ~A169 & \new_[43206]_ ;
  assign \new_[43210]_  = A201 & A199;
  assign \new_[43213]_  = A233 & A232;
  assign \new_[43214]_  = \new_[43213]_  & \new_[43210]_ ;
  assign \new_[43215]_  = \new_[43214]_  & \new_[43207]_ ;
  assign \new_[43219]_  = A265 & ~A235;
  assign \new_[43220]_  = ~A234 & \new_[43219]_ ;
  assign \new_[43223]_  = ~A267 & A266;
  assign \new_[43226]_  = A301 & ~A268;
  assign \new_[43227]_  = \new_[43226]_  & \new_[43223]_ ;
  assign \new_[43228]_  = \new_[43227]_  & \new_[43220]_ ;
  assign \new_[43232]_  = ~A166 & ~A167;
  assign \new_[43233]_  = ~A169 & \new_[43232]_ ;
  assign \new_[43236]_  = A201 & A199;
  assign \new_[43239]_  = A233 & A232;
  assign \new_[43240]_  = \new_[43239]_  & \new_[43236]_ ;
  assign \new_[43241]_  = \new_[43240]_  & \new_[43233]_ ;
  assign \new_[43245]_  = ~A265 & ~A235;
  assign \new_[43246]_  = ~A234 & \new_[43245]_ ;
  assign \new_[43249]_  = ~A268 & ~A266;
  assign \new_[43252]_  = A300 & A299;
  assign \new_[43253]_  = \new_[43252]_  & \new_[43249]_ ;
  assign \new_[43254]_  = \new_[43253]_  & \new_[43246]_ ;
  assign \new_[43258]_  = ~A166 & ~A167;
  assign \new_[43259]_  = ~A169 & \new_[43258]_ ;
  assign \new_[43262]_  = A201 & A199;
  assign \new_[43265]_  = A233 & A232;
  assign \new_[43266]_  = \new_[43265]_  & \new_[43262]_ ;
  assign \new_[43267]_  = \new_[43266]_  & \new_[43259]_ ;
  assign \new_[43271]_  = ~A265 & ~A235;
  assign \new_[43272]_  = ~A234 & \new_[43271]_ ;
  assign \new_[43275]_  = ~A268 & ~A266;
  assign \new_[43278]_  = A300 & A298;
  assign \new_[43279]_  = \new_[43278]_  & \new_[43275]_ ;
  assign \new_[43280]_  = \new_[43279]_  & \new_[43272]_ ;
  assign \new_[43284]_  = ~A166 & ~A167;
  assign \new_[43285]_  = ~A169 & \new_[43284]_ ;
  assign \new_[43288]_  = A201 & A199;
  assign \new_[43291]_  = ~A233 & ~A232;
  assign \new_[43292]_  = \new_[43291]_  & \new_[43288]_ ;
  assign \new_[43293]_  = \new_[43292]_  & \new_[43285]_ ;
  assign \new_[43297]_  = ~A268 & ~A267;
  assign \new_[43298]_  = ~A235 & \new_[43297]_ ;
  assign \new_[43301]_  = A298 & ~A269;
  assign \new_[43304]_  = A302 & ~A299;
  assign \new_[43305]_  = \new_[43304]_  & \new_[43301]_ ;
  assign \new_[43306]_  = \new_[43305]_  & \new_[43298]_ ;
  assign \new_[43310]_  = ~A166 & ~A167;
  assign \new_[43311]_  = ~A169 & \new_[43310]_ ;
  assign \new_[43314]_  = A201 & A199;
  assign \new_[43317]_  = ~A233 & ~A232;
  assign \new_[43318]_  = \new_[43317]_  & \new_[43314]_ ;
  assign \new_[43319]_  = \new_[43318]_  & \new_[43311]_ ;
  assign \new_[43323]_  = ~A268 & ~A267;
  assign \new_[43324]_  = ~A235 & \new_[43323]_ ;
  assign \new_[43327]_  = ~A298 & ~A269;
  assign \new_[43330]_  = A302 & A299;
  assign \new_[43331]_  = \new_[43330]_  & \new_[43327]_ ;
  assign \new_[43332]_  = \new_[43331]_  & \new_[43324]_ ;
  assign \new_[43336]_  = ~A166 & ~A167;
  assign \new_[43337]_  = ~A169 & \new_[43336]_ ;
  assign \new_[43340]_  = A201 & A199;
  assign \new_[43343]_  = ~A233 & ~A232;
  assign \new_[43344]_  = \new_[43343]_  & \new_[43340]_ ;
  assign \new_[43345]_  = \new_[43344]_  & \new_[43337]_ ;
  assign \new_[43349]_  = A266 & A265;
  assign \new_[43350]_  = ~A235 & \new_[43349]_ ;
  assign \new_[43353]_  = ~A268 & ~A267;
  assign \new_[43356]_  = A300 & A299;
  assign \new_[43357]_  = \new_[43356]_  & \new_[43353]_ ;
  assign \new_[43358]_  = \new_[43357]_  & \new_[43350]_ ;
  assign \new_[43362]_  = ~A166 & ~A167;
  assign \new_[43363]_  = ~A169 & \new_[43362]_ ;
  assign \new_[43366]_  = A201 & A199;
  assign \new_[43369]_  = ~A233 & ~A232;
  assign \new_[43370]_  = \new_[43369]_  & \new_[43366]_ ;
  assign \new_[43371]_  = \new_[43370]_  & \new_[43363]_ ;
  assign \new_[43375]_  = A266 & A265;
  assign \new_[43376]_  = ~A235 & \new_[43375]_ ;
  assign \new_[43379]_  = ~A268 & ~A267;
  assign \new_[43382]_  = A300 & A298;
  assign \new_[43383]_  = \new_[43382]_  & \new_[43379]_ ;
  assign \new_[43384]_  = \new_[43383]_  & \new_[43376]_ ;
  assign \new_[43388]_  = ~A166 & ~A167;
  assign \new_[43389]_  = ~A169 & \new_[43388]_ ;
  assign \new_[43392]_  = A201 & A199;
  assign \new_[43395]_  = ~A233 & ~A232;
  assign \new_[43396]_  = \new_[43395]_  & \new_[43392]_ ;
  assign \new_[43397]_  = \new_[43396]_  & \new_[43389]_ ;
  assign \new_[43401]_  = ~A266 & ~A265;
  assign \new_[43402]_  = ~A235 & \new_[43401]_ ;
  assign \new_[43405]_  = A298 & ~A268;
  assign \new_[43408]_  = A302 & ~A299;
  assign \new_[43409]_  = \new_[43408]_  & \new_[43405]_ ;
  assign \new_[43410]_  = \new_[43409]_  & \new_[43402]_ ;
  assign \new_[43414]_  = ~A166 & ~A167;
  assign \new_[43415]_  = ~A169 & \new_[43414]_ ;
  assign \new_[43418]_  = A201 & A199;
  assign \new_[43421]_  = ~A233 & ~A232;
  assign \new_[43422]_  = \new_[43421]_  & \new_[43418]_ ;
  assign \new_[43423]_  = \new_[43422]_  & \new_[43415]_ ;
  assign \new_[43427]_  = ~A266 & ~A265;
  assign \new_[43428]_  = ~A235 & \new_[43427]_ ;
  assign \new_[43431]_  = ~A298 & ~A268;
  assign \new_[43434]_  = A302 & A299;
  assign \new_[43435]_  = \new_[43434]_  & \new_[43431]_ ;
  assign \new_[43436]_  = \new_[43435]_  & \new_[43428]_ ;
  assign \new_[43440]_  = ~A166 & ~A167;
  assign \new_[43441]_  = ~A169 & \new_[43440]_ ;
  assign \new_[43444]_  = A201 & A200;
  assign \new_[43447]_  = ~A235 & ~A234;
  assign \new_[43448]_  = \new_[43447]_  & \new_[43444]_ ;
  assign \new_[43449]_  = \new_[43448]_  & \new_[43441]_ ;
  assign \new_[43453]_  = ~A268 & ~A267;
  assign \new_[43454]_  = ~A236 & \new_[43453]_ ;
  assign \new_[43457]_  = A298 & ~A269;
  assign \new_[43460]_  = A302 & ~A299;
  assign \new_[43461]_  = \new_[43460]_  & \new_[43457]_ ;
  assign \new_[43462]_  = \new_[43461]_  & \new_[43454]_ ;
  assign \new_[43466]_  = ~A166 & ~A167;
  assign \new_[43467]_  = ~A169 & \new_[43466]_ ;
  assign \new_[43470]_  = A201 & A200;
  assign \new_[43473]_  = ~A235 & ~A234;
  assign \new_[43474]_  = \new_[43473]_  & \new_[43470]_ ;
  assign \new_[43475]_  = \new_[43474]_  & \new_[43467]_ ;
  assign \new_[43479]_  = ~A268 & ~A267;
  assign \new_[43480]_  = ~A236 & \new_[43479]_ ;
  assign \new_[43483]_  = ~A298 & ~A269;
  assign \new_[43486]_  = A302 & A299;
  assign \new_[43487]_  = \new_[43486]_  & \new_[43483]_ ;
  assign \new_[43488]_  = \new_[43487]_  & \new_[43480]_ ;
  assign \new_[43492]_  = ~A166 & ~A167;
  assign \new_[43493]_  = ~A169 & \new_[43492]_ ;
  assign \new_[43496]_  = A201 & A200;
  assign \new_[43499]_  = ~A235 & ~A234;
  assign \new_[43500]_  = \new_[43499]_  & \new_[43496]_ ;
  assign \new_[43501]_  = \new_[43500]_  & \new_[43493]_ ;
  assign \new_[43505]_  = A266 & A265;
  assign \new_[43506]_  = ~A236 & \new_[43505]_ ;
  assign \new_[43509]_  = ~A268 & ~A267;
  assign \new_[43512]_  = A300 & A299;
  assign \new_[43513]_  = \new_[43512]_  & \new_[43509]_ ;
  assign \new_[43514]_  = \new_[43513]_  & \new_[43506]_ ;
  assign \new_[43518]_  = ~A166 & ~A167;
  assign \new_[43519]_  = ~A169 & \new_[43518]_ ;
  assign \new_[43522]_  = A201 & A200;
  assign \new_[43525]_  = ~A235 & ~A234;
  assign \new_[43526]_  = \new_[43525]_  & \new_[43522]_ ;
  assign \new_[43527]_  = \new_[43526]_  & \new_[43519]_ ;
  assign \new_[43531]_  = A266 & A265;
  assign \new_[43532]_  = ~A236 & \new_[43531]_ ;
  assign \new_[43535]_  = ~A268 & ~A267;
  assign \new_[43538]_  = A300 & A298;
  assign \new_[43539]_  = \new_[43538]_  & \new_[43535]_ ;
  assign \new_[43540]_  = \new_[43539]_  & \new_[43532]_ ;
  assign \new_[43544]_  = ~A166 & ~A167;
  assign \new_[43545]_  = ~A169 & \new_[43544]_ ;
  assign \new_[43548]_  = A201 & A200;
  assign \new_[43551]_  = ~A235 & ~A234;
  assign \new_[43552]_  = \new_[43551]_  & \new_[43548]_ ;
  assign \new_[43553]_  = \new_[43552]_  & \new_[43545]_ ;
  assign \new_[43557]_  = ~A266 & ~A265;
  assign \new_[43558]_  = ~A236 & \new_[43557]_ ;
  assign \new_[43561]_  = A298 & ~A268;
  assign \new_[43564]_  = A302 & ~A299;
  assign \new_[43565]_  = \new_[43564]_  & \new_[43561]_ ;
  assign \new_[43566]_  = \new_[43565]_  & \new_[43558]_ ;
  assign \new_[43570]_  = ~A166 & ~A167;
  assign \new_[43571]_  = ~A169 & \new_[43570]_ ;
  assign \new_[43574]_  = A201 & A200;
  assign \new_[43577]_  = ~A235 & ~A234;
  assign \new_[43578]_  = \new_[43577]_  & \new_[43574]_ ;
  assign \new_[43579]_  = \new_[43578]_  & \new_[43571]_ ;
  assign \new_[43583]_  = ~A266 & ~A265;
  assign \new_[43584]_  = ~A236 & \new_[43583]_ ;
  assign \new_[43587]_  = ~A298 & ~A268;
  assign \new_[43590]_  = A302 & A299;
  assign \new_[43591]_  = \new_[43590]_  & \new_[43587]_ ;
  assign \new_[43592]_  = \new_[43591]_  & \new_[43584]_ ;
  assign \new_[43596]_  = ~A166 & ~A167;
  assign \new_[43597]_  = ~A169 & \new_[43596]_ ;
  assign \new_[43600]_  = A201 & A200;
  assign \new_[43603]_  = A233 & A232;
  assign \new_[43604]_  = \new_[43603]_  & \new_[43600]_ ;
  assign \new_[43605]_  = \new_[43604]_  & \new_[43597]_ ;
  assign \new_[43609]_  = ~A267 & ~A235;
  assign \new_[43610]_  = ~A234 & \new_[43609]_ ;
  assign \new_[43613]_  = ~A269 & ~A268;
  assign \new_[43616]_  = A300 & A299;
  assign \new_[43617]_  = \new_[43616]_  & \new_[43613]_ ;
  assign \new_[43618]_  = \new_[43617]_  & \new_[43610]_ ;
  assign \new_[43622]_  = ~A166 & ~A167;
  assign \new_[43623]_  = ~A169 & \new_[43622]_ ;
  assign \new_[43626]_  = A201 & A200;
  assign \new_[43629]_  = A233 & A232;
  assign \new_[43630]_  = \new_[43629]_  & \new_[43626]_ ;
  assign \new_[43631]_  = \new_[43630]_  & \new_[43623]_ ;
  assign \new_[43635]_  = ~A267 & ~A235;
  assign \new_[43636]_  = ~A234 & \new_[43635]_ ;
  assign \new_[43639]_  = ~A269 & ~A268;
  assign \new_[43642]_  = A300 & A298;
  assign \new_[43643]_  = \new_[43642]_  & \new_[43639]_ ;
  assign \new_[43644]_  = \new_[43643]_  & \new_[43636]_ ;
  assign \new_[43648]_  = ~A166 & ~A167;
  assign \new_[43649]_  = ~A169 & \new_[43648]_ ;
  assign \new_[43652]_  = A201 & A200;
  assign \new_[43655]_  = A233 & A232;
  assign \new_[43656]_  = \new_[43655]_  & \new_[43652]_ ;
  assign \new_[43657]_  = \new_[43656]_  & \new_[43649]_ ;
  assign \new_[43661]_  = A265 & ~A235;
  assign \new_[43662]_  = ~A234 & \new_[43661]_ ;
  assign \new_[43665]_  = ~A267 & A266;
  assign \new_[43668]_  = A301 & ~A268;
  assign \new_[43669]_  = \new_[43668]_  & \new_[43665]_ ;
  assign \new_[43670]_  = \new_[43669]_  & \new_[43662]_ ;
  assign \new_[43674]_  = ~A166 & ~A167;
  assign \new_[43675]_  = ~A169 & \new_[43674]_ ;
  assign \new_[43678]_  = A201 & A200;
  assign \new_[43681]_  = A233 & A232;
  assign \new_[43682]_  = \new_[43681]_  & \new_[43678]_ ;
  assign \new_[43683]_  = \new_[43682]_  & \new_[43675]_ ;
  assign \new_[43687]_  = ~A265 & ~A235;
  assign \new_[43688]_  = ~A234 & \new_[43687]_ ;
  assign \new_[43691]_  = ~A268 & ~A266;
  assign \new_[43694]_  = A300 & A299;
  assign \new_[43695]_  = \new_[43694]_  & \new_[43691]_ ;
  assign \new_[43696]_  = \new_[43695]_  & \new_[43688]_ ;
  assign \new_[43700]_  = ~A166 & ~A167;
  assign \new_[43701]_  = ~A169 & \new_[43700]_ ;
  assign \new_[43704]_  = A201 & A200;
  assign \new_[43707]_  = A233 & A232;
  assign \new_[43708]_  = \new_[43707]_  & \new_[43704]_ ;
  assign \new_[43709]_  = \new_[43708]_  & \new_[43701]_ ;
  assign \new_[43713]_  = ~A265 & ~A235;
  assign \new_[43714]_  = ~A234 & \new_[43713]_ ;
  assign \new_[43717]_  = ~A268 & ~A266;
  assign \new_[43720]_  = A300 & A298;
  assign \new_[43721]_  = \new_[43720]_  & \new_[43717]_ ;
  assign \new_[43722]_  = \new_[43721]_  & \new_[43714]_ ;
  assign \new_[43726]_  = ~A166 & ~A167;
  assign \new_[43727]_  = ~A169 & \new_[43726]_ ;
  assign \new_[43730]_  = A201 & A200;
  assign \new_[43733]_  = ~A233 & ~A232;
  assign \new_[43734]_  = \new_[43733]_  & \new_[43730]_ ;
  assign \new_[43735]_  = \new_[43734]_  & \new_[43727]_ ;
  assign \new_[43739]_  = ~A268 & ~A267;
  assign \new_[43740]_  = ~A235 & \new_[43739]_ ;
  assign \new_[43743]_  = A298 & ~A269;
  assign \new_[43746]_  = A302 & ~A299;
  assign \new_[43747]_  = \new_[43746]_  & \new_[43743]_ ;
  assign \new_[43748]_  = \new_[43747]_  & \new_[43740]_ ;
  assign \new_[43752]_  = ~A166 & ~A167;
  assign \new_[43753]_  = ~A169 & \new_[43752]_ ;
  assign \new_[43756]_  = A201 & A200;
  assign \new_[43759]_  = ~A233 & ~A232;
  assign \new_[43760]_  = \new_[43759]_  & \new_[43756]_ ;
  assign \new_[43761]_  = \new_[43760]_  & \new_[43753]_ ;
  assign \new_[43765]_  = ~A268 & ~A267;
  assign \new_[43766]_  = ~A235 & \new_[43765]_ ;
  assign \new_[43769]_  = ~A298 & ~A269;
  assign \new_[43772]_  = A302 & A299;
  assign \new_[43773]_  = \new_[43772]_  & \new_[43769]_ ;
  assign \new_[43774]_  = \new_[43773]_  & \new_[43766]_ ;
  assign \new_[43778]_  = ~A166 & ~A167;
  assign \new_[43779]_  = ~A169 & \new_[43778]_ ;
  assign \new_[43782]_  = A201 & A200;
  assign \new_[43785]_  = ~A233 & ~A232;
  assign \new_[43786]_  = \new_[43785]_  & \new_[43782]_ ;
  assign \new_[43787]_  = \new_[43786]_  & \new_[43779]_ ;
  assign \new_[43791]_  = A266 & A265;
  assign \new_[43792]_  = ~A235 & \new_[43791]_ ;
  assign \new_[43795]_  = ~A268 & ~A267;
  assign \new_[43798]_  = A300 & A299;
  assign \new_[43799]_  = \new_[43798]_  & \new_[43795]_ ;
  assign \new_[43800]_  = \new_[43799]_  & \new_[43792]_ ;
  assign \new_[43804]_  = ~A166 & ~A167;
  assign \new_[43805]_  = ~A169 & \new_[43804]_ ;
  assign \new_[43808]_  = A201 & A200;
  assign \new_[43811]_  = ~A233 & ~A232;
  assign \new_[43812]_  = \new_[43811]_  & \new_[43808]_ ;
  assign \new_[43813]_  = \new_[43812]_  & \new_[43805]_ ;
  assign \new_[43817]_  = A266 & A265;
  assign \new_[43818]_  = ~A235 & \new_[43817]_ ;
  assign \new_[43821]_  = ~A268 & ~A267;
  assign \new_[43824]_  = A300 & A298;
  assign \new_[43825]_  = \new_[43824]_  & \new_[43821]_ ;
  assign \new_[43826]_  = \new_[43825]_  & \new_[43818]_ ;
  assign \new_[43830]_  = ~A166 & ~A167;
  assign \new_[43831]_  = ~A169 & \new_[43830]_ ;
  assign \new_[43834]_  = A201 & A200;
  assign \new_[43837]_  = ~A233 & ~A232;
  assign \new_[43838]_  = \new_[43837]_  & \new_[43834]_ ;
  assign \new_[43839]_  = \new_[43838]_  & \new_[43831]_ ;
  assign \new_[43843]_  = ~A266 & ~A265;
  assign \new_[43844]_  = ~A235 & \new_[43843]_ ;
  assign \new_[43847]_  = A298 & ~A268;
  assign \new_[43850]_  = A302 & ~A299;
  assign \new_[43851]_  = \new_[43850]_  & \new_[43847]_ ;
  assign \new_[43852]_  = \new_[43851]_  & \new_[43844]_ ;
  assign \new_[43856]_  = ~A166 & ~A167;
  assign \new_[43857]_  = ~A169 & \new_[43856]_ ;
  assign \new_[43860]_  = A201 & A200;
  assign \new_[43863]_  = ~A233 & ~A232;
  assign \new_[43864]_  = \new_[43863]_  & \new_[43860]_ ;
  assign \new_[43865]_  = \new_[43864]_  & \new_[43857]_ ;
  assign \new_[43869]_  = ~A266 & ~A265;
  assign \new_[43870]_  = ~A235 & \new_[43869]_ ;
  assign \new_[43873]_  = ~A298 & ~A268;
  assign \new_[43876]_  = A302 & A299;
  assign \new_[43877]_  = \new_[43876]_  & \new_[43873]_ ;
  assign \new_[43878]_  = \new_[43877]_  & \new_[43870]_ ;
  assign \new_[43882]_  = ~A166 & ~A167;
  assign \new_[43883]_  = ~A169 & \new_[43882]_ ;
  assign \new_[43886]_  = A200 & ~A199;
  assign \new_[43889]_  = ~A234 & A203;
  assign \new_[43890]_  = \new_[43889]_  & \new_[43886]_ ;
  assign \new_[43891]_  = \new_[43890]_  & \new_[43883]_ ;
  assign \new_[43895]_  = ~A267 & ~A236;
  assign \new_[43896]_  = ~A235 & \new_[43895]_ ;
  assign \new_[43899]_  = ~A269 & ~A268;
  assign \new_[43902]_  = A300 & A299;
  assign \new_[43903]_  = \new_[43902]_  & \new_[43899]_ ;
  assign \new_[43904]_  = \new_[43903]_  & \new_[43896]_ ;
  assign \new_[43908]_  = ~A166 & ~A167;
  assign \new_[43909]_  = ~A169 & \new_[43908]_ ;
  assign \new_[43912]_  = A200 & ~A199;
  assign \new_[43915]_  = ~A234 & A203;
  assign \new_[43916]_  = \new_[43915]_  & \new_[43912]_ ;
  assign \new_[43917]_  = \new_[43916]_  & \new_[43909]_ ;
  assign \new_[43921]_  = ~A267 & ~A236;
  assign \new_[43922]_  = ~A235 & \new_[43921]_ ;
  assign \new_[43925]_  = ~A269 & ~A268;
  assign \new_[43928]_  = A300 & A298;
  assign \new_[43929]_  = \new_[43928]_  & \new_[43925]_ ;
  assign \new_[43930]_  = \new_[43929]_  & \new_[43922]_ ;
  assign \new_[43934]_  = ~A166 & ~A167;
  assign \new_[43935]_  = ~A169 & \new_[43934]_ ;
  assign \new_[43938]_  = A200 & ~A199;
  assign \new_[43941]_  = ~A234 & A203;
  assign \new_[43942]_  = \new_[43941]_  & \new_[43938]_ ;
  assign \new_[43943]_  = \new_[43942]_  & \new_[43935]_ ;
  assign \new_[43947]_  = A265 & ~A236;
  assign \new_[43948]_  = ~A235 & \new_[43947]_ ;
  assign \new_[43951]_  = ~A267 & A266;
  assign \new_[43954]_  = A301 & ~A268;
  assign \new_[43955]_  = \new_[43954]_  & \new_[43951]_ ;
  assign \new_[43956]_  = \new_[43955]_  & \new_[43948]_ ;
  assign \new_[43960]_  = ~A166 & ~A167;
  assign \new_[43961]_  = ~A169 & \new_[43960]_ ;
  assign \new_[43964]_  = A200 & ~A199;
  assign \new_[43967]_  = ~A234 & A203;
  assign \new_[43968]_  = \new_[43967]_  & \new_[43964]_ ;
  assign \new_[43969]_  = \new_[43968]_  & \new_[43961]_ ;
  assign \new_[43973]_  = ~A265 & ~A236;
  assign \new_[43974]_  = ~A235 & \new_[43973]_ ;
  assign \new_[43977]_  = ~A268 & ~A266;
  assign \new_[43980]_  = A300 & A299;
  assign \new_[43981]_  = \new_[43980]_  & \new_[43977]_ ;
  assign \new_[43982]_  = \new_[43981]_  & \new_[43974]_ ;
  assign \new_[43986]_  = ~A166 & ~A167;
  assign \new_[43987]_  = ~A169 & \new_[43986]_ ;
  assign \new_[43990]_  = A200 & ~A199;
  assign \new_[43993]_  = ~A234 & A203;
  assign \new_[43994]_  = \new_[43993]_  & \new_[43990]_ ;
  assign \new_[43995]_  = \new_[43994]_  & \new_[43987]_ ;
  assign \new_[43999]_  = ~A265 & ~A236;
  assign \new_[44000]_  = ~A235 & \new_[43999]_ ;
  assign \new_[44003]_  = ~A268 & ~A266;
  assign \new_[44006]_  = A300 & A298;
  assign \new_[44007]_  = \new_[44006]_  & \new_[44003]_ ;
  assign \new_[44008]_  = \new_[44007]_  & \new_[44000]_ ;
  assign \new_[44012]_  = ~A166 & ~A167;
  assign \new_[44013]_  = ~A169 & \new_[44012]_ ;
  assign \new_[44016]_  = A200 & ~A199;
  assign \new_[44019]_  = A232 & A203;
  assign \new_[44020]_  = \new_[44019]_  & \new_[44016]_ ;
  assign \new_[44021]_  = \new_[44020]_  & \new_[44013]_ ;
  assign \new_[44025]_  = ~A235 & ~A234;
  assign \new_[44026]_  = A233 & \new_[44025]_ ;
  assign \new_[44029]_  = ~A268 & ~A267;
  assign \new_[44032]_  = A301 & ~A269;
  assign \new_[44033]_  = \new_[44032]_  & \new_[44029]_ ;
  assign \new_[44034]_  = \new_[44033]_  & \new_[44026]_ ;
  assign \new_[44038]_  = ~A166 & ~A167;
  assign \new_[44039]_  = ~A169 & \new_[44038]_ ;
  assign \new_[44042]_  = A200 & ~A199;
  assign \new_[44045]_  = A232 & A203;
  assign \new_[44046]_  = \new_[44045]_  & \new_[44042]_ ;
  assign \new_[44047]_  = \new_[44046]_  & \new_[44039]_ ;
  assign \new_[44051]_  = ~A235 & ~A234;
  assign \new_[44052]_  = A233 & \new_[44051]_ ;
  assign \new_[44055]_  = ~A266 & ~A265;
  assign \new_[44058]_  = A301 & ~A268;
  assign \new_[44059]_  = \new_[44058]_  & \new_[44055]_ ;
  assign \new_[44060]_  = \new_[44059]_  & \new_[44052]_ ;
  assign \new_[44064]_  = ~A166 & ~A167;
  assign \new_[44065]_  = ~A169 & \new_[44064]_ ;
  assign \new_[44068]_  = A200 & ~A199;
  assign \new_[44071]_  = ~A232 & A203;
  assign \new_[44072]_  = \new_[44071]_  & \new_[44068]_ ;
  assign \new_[44073]_  = \new_[44072]_  & \new_[44065]_ ;
  assign \new_[44077]_  = ~A267 & ~A235;
  assign \new_[44078]_  = ~A233 & \new_[44077]_ ;
  assign \new_[44081]_  = ~A269 & ~A268;
  assign \new_[44084]_  = A300 & A299;
  assign \new_[44085]_  = \new_[44084]_  & \new_[44081]_ ;
  assign \new_[44086]_  = \new_[44085]_  & \new_[44078]_ ;
  assign \new_[44090]_  = ~A166 & ~A167;
  assign \new_[44091]_  = ~A169 & \new_[44090]_ ;
  assign \new_[44094]_  = A200 & ~A199;
  assign \new_[44097]_  = ~A232 & A203;
  assign \new_[44098]_  = \new_[44097]_  & \new_[44094]_ ;
  assign \new_[44099]_  = \new_[44098]_  & \new_[44091]_ ;
  assign \new_[44103]_  = ~A267 & ~A235;
  assign \new_[44104]_  = ~A233 & \new_[44103]_ ;
  assign \new_[44107]_  = ~A269 & ~A268;
  assign \new_[44110]_  = A300 & A298;
  assign \new_[44111]_  = \new_[44110]_  & \new_[44107]_ ;
  assign \new_[44112]_  = \new_[44111]_  & \new_[44104]_ ;
  assign \new_[44116]_  = ~A166 & ~A167;
  assign \new_[44117]_  = ~A169 & \new_[44116]_ ;
  assign \new_[44120]_  = A200 & ~A199;
  assign \new_[44123]_  = ~A232 & A203;
  assign \new_[44124]_  = \new_[44123]_  & \new_[44120]_ ;
  assign \new_[44125]_  = \new_[44124]_  & \new_[44117]_ ;
  assign \new_[44129]_  = A265 & ~A235;
  assign \new_[44130]_  = ~A233 & \new_[44129]_ ;
  assign \new_[44133]_  = ~A267 & A266;
  assign \new_[44136]_  = A301 & ~A268;
  assign \new_[44137]_  = \new_[44136]_  & \new_[44133]_ ;
  assign \new_[44138]_  = \new_[44137]_  & \new_[44130]_ ;
  assign \new_[44142]_  = ~A166 & ~A167;
  assign \new_[44143]_  = ~A169 & \new_[44142]_ ;
  assign \new_[44146]_  = A200 & ~A199;
  assign \new_[44149]_  = ~A232 & A203;
  assign \new_[44150]_  = \new_[44149]_  & \new_[44146]_ ;
  assign \new_[44151]_  = \new_[44150]_  & \new_[44143]_ ;
  assign \new_[44155]_  = ~A265 & ~A235;
  assign \new_[44156]_  = ~A233 & \new_[44155]_ ;
  assign \new_[44159]_  = ~A268 & ~A266;
  assign \new_[44162]_  = A300 & A299;
  assign \new_[44163]_  = \new_[44162]_  & \new_[44159]_ ;
  assign \new_[44164]_  = \new_[44163]_  & \new_[44156]_ ;
  assign \new_[44168]_  = ~A166 & ~A167;
  assign \new_[44169]_  = ~A169 & \new_[44168]_ ;
  assign \new_[44172]_  = A200 & ~A199;
  assign \new_[44175]_  = ~A232 & A203;
  assign \new_[44176]_  = \new_[44175]_  & \new_[44172]_ ;
  assign \new_[44177]_  = \new_[44176]_  & \new_[44169]_ ;
  assign \new_[44181]_  = ~A265 & ~A235;
  assign \new_[44182]_  = ~A233 & \new_[44181]_ ;
  assign \new_[44185]_  = ~A268 & ~A266;
  assign \new_[44188]_  = A300 & A298;
  assign \new_[44189]_  = \new_[44188]_  & \new_[44185]_ ;
  assign \new_[44190]_  = \new_[44189]_  & \new_[44182]_ ;
  assign \new_[44194]_  = ~A166 & ~A167;
  assign \new_[44195]_  = ~A169 & \new_[44194]_ ;
  assign \new_[44198]_  = ~A200 & A199;
  assign \new_[44201]_  = ~A234 & A203;
  assign \new_[44202]_  = \new_[44201]_  & \new_[44198]_ ;
  assign \new_[44203]_  = \new_[44202]_  & \new_[44195]_ ;
  assign \new_[44207]_  = ~A267 & ~A236;
  assign \new_[44208]_  = ~A235 & \new_[44207]_ ;
  assign \new_[44211]_  = ~A269 & ~A268;
  assign \new_[44214]_  = A300 & A299;
  assign \new_[44215]_  = \new_[44214]_  & \new_[44211]_ ;
  assign \new_[44216]_  = \new_[44215]_  & \new_[44208]_ ;
  assign \new_[44220]_  = ~A166 & ~A167;
  assign \new_[44221]_  = ~A169 & \new_[44220]_ ;
  assign \new_[44224]_  = ~A200 & A199;
  assign \new_[44227]_  = ~A234 & A203;
  assign \new_[44228]_  = \new_[44227]_  & \new_[44224]_ ;
  assign \new_[44229]_  = \new_[44228]_  & \new_[44221]_ ;
  assign \new_[44233]_  = ~A267 & ~A236;
  assign \new_[44234]_  = ~A235 & \new_[44233]_ ;
  assign \new_[44237]_  = ~A269 & ~A268;
  assign \new_[44240]_  = A300 & A298;
  assign \new_[44241]_  = \new_[44240]_  & \new_[44237]_ ;
  assign \new_[44242]_  = \new_[44241]_  & \new_[44234]_ ;
  assign \new_[44246]_  = ~A166 & ~A167;
  assign \new_[44247]_  = ~A169 & \new_[44246]_ ;
  assign \new_[44250]_  = ~A200 & A199;
  assign \new_[44253]_  = ~A234 & A203;
  assign \new_[44254]_  = \new_[44253]_  & \new_[44250]_ ;
  assign \new_[44255]_  = \new_[44254]_  & \new_[44247]_ ;
  assign \new_[44259]_  = A265 & ~A236;
  assign \new_[44260]_  = ~A235 & \new_[44259]_ ;
  assign \new_[44263]_  = ~A267 & A266;
  assign \new_[44266]_  = A301 & ~A268;
  assign \new_[44267]_  = \new_[44266]_  & \new_[44263]_ ;
  assign \new_[44268]_  = \new_[44267]_  & \new_[44260]_ ;
  assign \new_[44272]_  = ~A166 & ~A167;
  assign \new_[44273]_  = ~A169 & \new_[44272]_ ;
  assign \new_[44276]_  = ~A200 & A199;
  assign \new_[44279]_  = ~A234 & A203;
  assign \new_[44280]_  = \new_[44279]_  & \new_[44276]_ ;
  assign \new_[44281]_  = \new_[44280]_  & \new_[44273]_ ;
  assign \new_[44285]_  = ~A265 & ~A236;
  assign \new_[44286]_  = ~A235 & \new_[44285]_ ;
  assign \new_[44289]_  = ~A268 & ~A266;
  assign \new_[44292]_  = A300 & A299;
  assign \new_[44293]_  = \new_[44292]_  & \new_[44289]_ ;
  assign \new_[44294]_  = \new_[44293]_  & \new_[44286]_ ;
  assign \new_[44298]_  = ~A166 & ~A167;
  assign \new_[44299]_  = ~A169 & \new_[44298]_ ;
  assign \new_[44302]_  = ~A200 & A199;
  assign \new_[44305]_  = ~A234 & A203;
  assign \new_[44306]_  = \new_[44305]_  & \new_[44302]_ ;
  assign \new_[44307]_  = \new_[44306]_  & \new_[44299]_ ;
  assign \new_[44311]_  = ~A265 & ~A236;
  assign \new_[44312]_  = ~A235 & \new_[44311]_ ;
  assign \new_[44315]_  = ~A268 & ~A266;
  assign \new_[44318]_  = A300 & A298;
  assign \new_[44319]_  = \new_[44318]_  & \new_[44315]_ ;
  assign \new_[44320]_  = \new_[44319]_  & \new_[44312]_ ;
  assign \new_[44324]_  = ~A166 & ~A167;
  assign \new_[44325]_  = ~A169 & \new_[44324]_ ;
  assign \new_[44328]_  = ~A200 & A199;
  assign \new_[44331]_  = A232 & A203;
  assign \new_[44332]_  = \new_[44331]_  & \new_[44328]_ ;
  assign \new_[44333]_  = \new_[44332]_  & \new_[44325]_ ;
  assign \new_[44337]_  = ~A235 & ~A234;
  assign \new_[44338]_  = A233 & \new_[44337]_ ;
  assign \new_[44341]_  = ~A268 & ~A267;
  assign \new_[44344]_  = A301 & ~A269;
  assign \new_[44345]_  = \new_[44344]_  & \new_[44341]_ ;
  assign \new_[44346]_  = \new_[44345]_  & \new_[44338]_ ;
  assign \new_[44350]_  = ~A166 & ~A167;
  assign \new_[44351]_  = ~A169 & \new_[44350]_ ;
  assign \new_[44354]_  = ~A200 & A199;
  assign \new_[44357]_  = A232 & A203;
  assign \new_[44358]_  = \new_[44357]_  & \new_[44354]_ ;
  assign \new_[44359]_  = \new_[44358]_  & \new_[44351]_ ;
  assign \new_[44363]_  = ~A235 & ~A234;
  assign \new_[44364]_  = A233 & \new_[44363]_ ;
  assign \new_[44367]_  = ~A266 & ~A265;
  assign \new_[44370]_  = A301 & ~A268;
  assign \new_[44371]_  = \new_[44370]_  & \new_[44367]_ ;
  assign \new_[44372]_  = \new_[44371]_  & \new_[44364]_ ;
  assign \new_[44376]_  = ~A166 & ~A167;
  assign \new_[44377]_  = ~A169 & \new_[44376]_ ;
  assign \new_[44380]_  = ~A200 & A199;
  assign \new_[44383]_  = ~A232 & A203;
  assign \new_[44384]_  = \new_[44383]_  & \new_[44380]_ ;
  assign \new_[44385]_  = \new_[44384]_  & \new_[44377]_ ;
  assign \new_[44389]_  = ~A267 & ~A235;
  assign \new_[44390]_  = ~A233 & \new_[44389]_ ;
  assign \new_[44393]_  = ~A269 & ~A268;
  assign \new_[44396]_  = A300 & A299;
  assign \new_[44397]_  = \new_[44396]_  & \new_[44393]_ ;
  assign \new_[44398]_  = \new_[44397]_  & \new_[44390]_ ;
  assign \new_[44402]_  = ~A166 & ~A167;
  assign \new_[44403]_  = ~A169 & \new_[44402]_ ;
  assign \new_[44406]_  = ~A200 & A199;
  assign \new_[44409]_  = ~A232 & A203;
  assign \new_[44410]_  = \new_[44409]_  & \new_[44406]_ ;
  assign \new_[44411]_  = \new_[44410]_  & \new_[44403]_ ;
  assign \new_[44415]_  = ~A267 & ~A235;
  assign \new_[44416]_  = ~A233 & \new_[44415]_ ;
  assign \new_[44419]_  = ~A269 & ~A268;
  assign \new_[44422]_  = A300 & A298;
  assign \new_[44423]_  = \new_[44422]_  & \new_[44419]_ ;
  assign \new_[44424]_  = \new_[44423]_  & \new_[44416]_ ;
  assign \new_[44428]_  = ~A166 & ~A167;
  assign \new_[44429]_  = ~A169 & \new_[44428]_ ;
  assign \new_[44432]_  = ~A200 & A199;
  assign \new_[44435]_  = ~A232 & A203;
  assign \new_[44436]_  = \new_[44435]_  & \new_[44432]_ ;
  assign \new_[44437]_  = \new_[44436]_  & \new_[44429]_ ;
  assign \new_[44441]_  = A265 & ~A235;
  assign \new_[44442]_  = ~A233 & \new_[44441]_ ;
  assign \new_[44445]_  = ~A267 & A266;
  assign \new_[44448]_  = A301 & ~A268;
  assign \new_[44449]_  = \new_[44448]_  & \new_[44445]_ ;
  assign \new_[44450]_  = \new_[44449]_  & \new_[44442]_ ;
  assign \new_[44454]_  = ~A166 & ~A167;
  assign \new_[44455]_  = ~A169 & \new_[44454]_ ;
  assign \new_[44458]_  = ~A200 & A199;
  assign \new_[44461]_  = ~A232 & A203;
  assign \new_[44462]_  = \new_[44461]_  & \new_[44458]_ ;
  assign \new_[44463]_  = \new_[44462]_  & \new_[44455]_ ;
  assign \new_[44467]_  = ~A265 & ~A235;
  assign \new_[44468]_  = ~A233 & \new_[44467]_ ;
  assign \new_[44471]_  = ~A268 & ~A266;
  assign \new_[44474]_  = A300 & A299;
  assign \new_[44475]_  = \new_[44474]_  & \new_[44471]_ ;
  assign \new_[44476]_  = \new_[44475]_  & \new_[44468]_ ;
  assign \new_[44480]_  = ~A166 & ~A167;
  assign \new_[44481]_  = ~A169 & \new_[44480]_ ;
  assign \new_[44484]_  = ~A200 & A199;
  assign \new_[44487]_  = ~A232 & A203;
  assign \new_[44488]_  = \new_[44487]_  & \new_[44484]_ ;
  assign \new_[44489]_  = \new_[44488]_  & \new_[44481]_ ;
  assign \new_[44493]_  = ~A265 & ~A235;
  assign \new_[44494]_  = ~A233 & \new_[44493]_ ;
  assign \new_[44497]_  = ~A268 & ~A266;
  assign \new_[44500]_  = A300 & A298;
  assign \new_[44501]_  = \new_[44500]_  & \new_[44497]_ ;
  assign \new_[44502]_  = \new_[44501]_  & \new_[44494]_ ;
  assign \new_[44506]_  = A167 & ~A168;
  assign \new_[44507]_  = ~A169 & \new_[44506]_ ;
  assign \new_[44510]_  = A202 & A166;
  assign \new_[44513]_  = ~A235 & ~A234;
  assign \new_[44514]_  = \new_[44513]_  & \new_[44510]_ ;
  assign \new_[44515]_  = \new_[44514]_  & \new_[44507]_ ;
  assign \new_[44519]_  = ~A268 & ~A267;
  assign \new_[44520]_  = ~A236 & \new_[44519]_ ;
  assign \new_[44523]_  = A298 & ~A269;
  assign \new_[44526]_  = A302 & ~A299;
  assign \new_[44527]_  = \new_[44526]_  & \new_[44523]_ ;
  assign \new_[44528]_  = \new_[44527]_  & \new_[44520]_ ;
  assign \new_[44532]_  = A167 & ~A168;
  assign \new_[44533]_  = ~A169 & \new_[44532]_ ;
  assign \new_[44536]_  = A202 & A166;
  assign \new_[44539]_  = ~A235 & ~A234;
  assign \new_[44540]_  = \new_[44539]_  & \new_[44536]_ ;
  assign \new_[44541]_  = \new_[44540]_  & \new_[44533]_ ;
  assign \new_[44545]_  = ~A268 & ~A267;
  assign \new_[44546]_  = ~A236 & \new_[44545]_ ;
  assign \new_[44549]_  = ~A298 & ~A269;
  assign \new_[44552]_  = A302 & A299;
  assign \new_[44553]_  = \new_[44552]_  & \new_[44549]_ ;
  assign \new_[44554]_  = \new_[44553]_  & \new_[44546]_ ;
  assign \new_[44558]_  = A167 & ~A168;
  assign \new_[44559]_  = ~A169 & \new_[44558]_ ;
  assign \new_[44562]_  = A202 & A166;
  assign \new_[44565]_  = ~A235 & ~A234;
  assign \new_[44566]_  = \new_[44565]_  & \new_[44562]_ ;
  assign \new_[44567]_  = \new_[44566]_  & \new_[44559]_ ;
  assign \new_[44571]_  = A266 & A265;
  assign \new_[44572]_  = ~A236 & \new_[44571]_ ;
  assign \new_[44575]_  = ~A268 & ~A267;
  assign \new_[44578]_  = A300 & A299;
  assign \new_[44579]_  = \new_[44578]_  & \new_[44575]_ ;
  assign \new_[44580]_  = \new_[44579]_  & \new_[44572]_ ;
  assign \new_[44584]_  = A167 & ~A168;
  assign \new_[44585]_  = ~A169 & \new_[44584]_ ;
  assign \new_[44588]_  = A202 & A166;
  assign \new_[44591]_  = ~A235 & ~A234;
  assign \new_[44592]_  = \new_[44591]_  & \new_[44588]_ ;
  assign \new_[44593]_  = \new_[44592]_  & \new_[44585]_ ;
  assign \new_[44597]_  = A266 & A265;
  assign \new_[44598]_  = ~A236 & \new_[44597]_ ;
  assign \new_[44601]_  = ~A268 & ~A267;
  assign \new_[44604]_  = A300 & A298;
  assign \new_[44605]_  = \new_[44604]_  & \new_[44601]_ ;
  assign \new_[44606]_  = \new_[44605]_  & \new_[44598]_ ;
  assign \new_[44610]_  = A167 & ~A168;
  assign \new_[44611]_  = ~A169 & \new_[44610]_ ;
  assign \new_[44614]_  = A202 & A166;
  assign \new_[44617]_  = ~A235 & ~A234;
  assign \new_[44618]_  = \new_[44617]_  & \new_[44614]_ ;
  assign \new_[44619]_  = \new_[44618]_  & \new_[44611]_ ;
  assign \new_[44623]_  = ~A266 & ~A265;
  assign \new_[44624]_  = ~A236 & \new_[44623]_ ;
  assign \new_[44627]_  = A298 & ~A268;
  assign \new_[44630]_  = A302 & ~A299;
  assign \new_[44631]_  = \new_[44630]_  & \new_[44627]_ ;
  assign \new_[44632]_  = \new_[44631]_  & \new_[44624]_ ;
  assign \new_[44636]_  = A167 & ~A168;
  assign \new_[44637]_  = ~A169 & \new_[44636]_ ;
  assign \new_[44640]_  = A202 & A166;
  assign \new_[44643]_  = ~A235 & ~A234;
  assign \new_[44644]_  = \new_[44643]_  & \new_[44640]_ ;
  assign \new_[44645]_  = \new_[44644]_  & \new_[44637]_ ;
  assign \new_[44649]_  = ~A266 & ~A265;
  assign \new_[44650]_  = ~A236 & \new_[44649]_ ;
  assign \new_[44653]_  = ~A298 & ~A268;
  assign \new_[44656]_  = A302 & A299;
  assign \new_[44657]_  = \new_[44656]_  & \new_[44653]_ ;
  assign \new_[44658]_  = \new_[44657]_  & \new_[44650]_ ;
  assign \new_[44662]_  = A167 & ~A168;
  assign \new_[44663]_  = ~A169 & \new_[44662]_ ;
  assign \new_[44666]_  = A202 & A166;
  assign \new_[44669]_  = A233 & A232;
  assign \new_[44670]_  = \new_[44669]_  & \new_[44666]_ ;
  assign \new_[44671]_  = \new_[44670]_  & \new_[44663]_ ;
  assign \new_[44675]_  = ~A267 & ~A235;
  assign \new_[44676]_  = ~A234 & \new_[44675]_ ;
  assign \new_[44679]_  = ~A269 & ~A268;
  assign \new_[44682]_  = A300 & A299;
  assign \new_[44683]_  = \new_[44682]_  & \new_[44679]_ ;
  assign \new_[44684]_  = \new_[44683]_  & \new_[44676]_ ;
  assign \new_[44688]_  = A167 & ~A168;
  assign \new_[44689]_  = ~A169 & \new_[44688]_ ;
  assign \new_[44692]_  = A202 & A166;
  assign \new_[44695]_  = A233 & A232;
  assign \new_[44696]_  = \new_[44695]_  & \new_[44692]_ ;
  assign \new_[44697]_  = \new_[44696]_  & \new_[44689]_ ;
  assign \new_[44701]_  = ~A267 & ~A235;
  assign \new_[44702]_  = ~A234 & \new_[44701]_ ;
  assign \new_[44705]_  = ~A269 & ~A268;
  assign \new_[44708]_  = A300 & A298;
  assign \new_[44709]_  = \new_[44708]_  & \new_[44705]_ ;
  assign \new_[44710]_  = \new_[44709]_  & \new_[44702]_ ;
  assign \new_[44714]_  = A167 & ~A168;
  assign \new_[44715]_  = ~A169 & \new_[44714]_ ;
  assign \new_[44718]_  = A202 & A166;
  assign \new_[44721]_  = A233 & A232;
  assign \new_[44722]_  = \new_[44721]_  & \new_[44718]_ ;
  assign \new_[44723]_  = \new_[44722]_  & \new_[44715]_ ;
  assign \new_[44727]_  = A265 & ~A235;
  assign \new_[44728]_  = ~A234 & \new_[44727]_ ;
  assign \new_[44731]_  = ~A267 & A266;
  assign \new_[44734]_  = A301 & ~A268;
  assign \new_[44735]_  = \new_[44734]_  & \new_[44731]_ ;
  assign \new_[44736]_  = \new_[44735]_  & \new_[44728]_ ;
  assign \new_[44740]_  = A167 & ~A168;
  assign \new_[44741]_  = ~A169 & \new_[44740]_ ;
  assign \new_[44744]_  = A202 & A166;
  assign \new_[44747]_  = A233 & A232;
  assign \new_[44748]_  = \new_[44747]_  & \new_[44744]_ ;
  assign \new_[44749]_  = \new_[44748]_  & \new_[44741]_ ;
  assign \new_[44753]_  = ~A265 & ~A235;
  assign \new_[44754]_  = ~A234 & \new_[44753]_ ;
  assign \new_[44757]_  = ~A268 & ~A266;
  assign \new_[44760]_  = A300 & A299;
  assign \new_[44761]_  = \new_[44760]_  & \new_[44757]_ ;
  assign \new_[44762]_  = \new_[44761]_  & \new_[44754]_ ;
  assign \new_[44766]_  = A167 & ~A168;
  assign \new_[44767]_  = ~A169 & \new_[44766]_ ;
  assign \new_[44770]_  = A202 & A166;
  assign \new_[44773]_  = A233 & A232;
  assign \new_[44774]_  = \new_[44773]_  & \new_[44770]_ ;
  assign \new_[44775]_  = \new_[44774]_  & \new_[44767]_ ;
  assign \new_[44779]_  = ~A265 & ~A235;
  assign \new_[44780]_  = ~A234 & \new_[44779]_ ;
  assign \new_[44783]_  = ~A268 & ~A266;
  assign \new_[44786]_  = A300 & A298;
  assign \new_[44787]_  = \new_[44786]_  & \new_[44783]_ ;
  assign \new_[44788]_  = \new_[44787]_  & \new_[44780]_ ;
  assign \new_[44792]_  = A167 & ~A168;
  assign \new_[44793]_  = ~A169 & \new_[44792]_ ;
  assign \new_[44796]_  = A202 & A166;
  assign \new_[44799]_  = ~A233 & ~A232;
  assign \new_[44800]_  = \new_[44799]_  & \new_[44796]_ ;
  assign \new_[44801]_  = \new_[44800]_  & \new_[44793]_ ;
  assign \new_[44805]_  = ~A268 & ~A267;
  assign \new_[44806]_  = ~A235 & \new_[44805]_ ;
  assign \new_[44809]_  = A298 & ~A269;
  assign \new_[44812]_  = A302 & ~A299;
  assign \new_[44813]_  = \new_[44812]_  & \new_[44809]_ ;
  assign \new_[44814]_  = \new_[44813]_  & \new_[44806]_ ;
  assign \new_[44818]_  = A167 & ~A168;
  assign \new_[44819]_  = ~A169 & \new_[44818]_ ;
  assign \new_[44822]_  = A202 & A166;
  assign \new_[44825]_  = ~A233 & ~A232;
  assign \new_[44826]_  = \new_[44825]_  & \new_[44822]_ ;
  assign \new_[44827]_  = \new_[44826]_  & \new_[44819]_ ;
  assign \new_[44831]_  = ~A268 & ~A267;
  assign \new_[44832]_  = ~A235 & \new_[44831]_ ;
  assign \new_[44835]_  = ~A298 & ~A269;
  assign \new_[44838]_  = A302 & A299;
  assign \new_[44839]_  = \new_[44838]_  & \new_[44835]_ ;
  assign \new_[44840]_  = \new_[44839]_  & \new_[44832]_ ;
  assign \new_[44844]_  = A167 & ~A168;
  assign \new_[44845]_  = ~A169 & \new_[44844]_ ;
  assign \new_[44848]_  = A202 & A166;
  assign \new_[44851]_  = ~A233 & ~A232;
  assign \new_[44852]_  = \new_[44851]_  & \new_[44848]_ ;
  assign \new_[44853]_  = \new_[44852]_  & \new_[44845]_ ;
  assign \new_[44857]_  = A266 & A265;
  assign \new_[44858]_  = ~A235 & \new_[44857]_ ;
  assign \new_[44861]_  = ~A268 & ~A267;
  assign \new_[44864]_  = A300 & A299;
  assign \new_[44865]_  = \new_[44864]_  & \new_[44861]_ ;
  assign \new_[44866]_  = \new_[44865]_  & \new_[44858]_ ;
  assign \new_[44870]_  = A167 & ~A168;
  assign \new_[44871]_  = ~A169 & \new_[44870]_ ;
  assign \new_[44874]_  = A202 & A166;
  assign \new_[44877]_  = ~A233 & ~A232;
  assign \new_[44878]_  = \new_[44877]_  & \new_[44874]_ ;
  assign \new_[44879]_  = \new_[44878]_  & \new_[44871]_ ;
  assign \new_[44883]_  = A266 & A265;
  assign \new_[44884]_  = ~A235 & \new_[44883]_ ;
  assign \new_[44887]_  = ~A268 & ~A267;
  assign \new_[44890]_  = A300 & A298;
  assign \new_[44891]_  = \new_[44890]_  & \new_[44887]_ ;
  assign \new_[44892]_  = \new_[44891]_  & \new_[44884]_ ;
  assign \new_[44896]_  = A167 & ~A168;
  assign \new_[44897]_  = ~A169 & \new_[44896]_ ;
  assign \new_[44900]_  = A202 & A166;
  assign \new_[44903]_  = ~A233 & ~A232;
  assign \new_[44904]_  = \new_[44903]_  & \new_[44900]_ ;
  assign \new_[44905]_  = \new_[44904]_  & \new_[44897]_ ;
  assign \new_[44909]_  = ~A266 & ~A265;
  assign \new_[44910]_  = ~A235 & \new_[44909]_ ;
  assign \new_[44913]_  = A298 & ~A268;
  assign \new_[44916]_  = A302 & ~A299;
  assign \new_[44917]_  = \new_[44916]_  & \new_[44913]_ ;
  assign \new_[44918]_  = \new_[44917]_  & \new_[44910]_ ;
  assign \new_[44922]_  = A167 & ~A168;
  assign \new_[44923]_  = ~A169 & \new_[44922]_ ;
  assign \new_[44926]_  = A202 & A166;
  assign \new_[44929]_  = ~A233 & ~A232;
  assign \new_[44930]_  = \new_[44929]_  & \new_[44926]_ ;
  assign \new_[44931]_  = \new_[44930]_  & \new_[44923]_ ;
  assign \new_[44935]_  = ~A266 & ~A265;
  assign \new_[44936]_  = ~A235 & \new_[44935]_ ;
  assign \new_[44939]_  = ~A298 & ~A268;
  assign \new_[44942]_  = A302 & A299;
  assign \new_[44943]_  = \new_[44942]_  & \new_[44939]_ ;
  assign \new_[44944]_  = \new_[44943]_  & \new_[44936]_ ;
  assign \new_[44948]_  = A167 & ~A168;
  assign \new_[44949]_  = ~A169 & \new_[44948]_ ;
  assign \new_[44952]_  = A199 & A166;
  assign \new_[44955]_  = ~A234 & A201;
  assign \new_[44956]_  = \new_[44955]_  & \new_[44952]_ ;
  assign \new_[44957]_  = \new_[44956]_  & \new_[44949]_ ;
  assign \new_[44961]_  = ~A267 & ~A236;
  assign \new_[44962]_  = ~A235 & \new_[44961]_ ;
  assign \new_[44965]_  = ~A269 & ~A268;
  assign \new_[44968]_  = A300 & A299;
  assign \new_[44969]_  = \new_[44968]_  & \new_[44965]_ ;
  assign \new_[44970]_  = \new_[44969]_  & \new_[44962]_ ;
  assign \new_[44974]_  = A167 & ~A168;
  assign \new_[44975]_  = ~A169 & \new_[44974]_ ;
  assign \new_[44978]_  = A199 & A166;
  assign \new_[44981]_  = ~A234 & A201;
  assign \new_[44982]_  = \new_[44981]_  & \new_[44978]_ ;
  assign \new_[44983]_  = \new_[44982]_  & \new_[44975]_ ;
  assign \new_[44987]_  = ~A267 & ~A236;
  assign \new_[44988]_  = ~A235 & \new_[44987]_ ;
  assign \new_[44991]_  = ~A269 & ~A268;
  assign \new_[44994]_  = A300 & A298;
  assign \new_[44995]_  = \new_[44994]_  & \new_[44991]_ ;
  assign \new_[44996]_  = \new_[44995]_  & \new_[44988]_ ;
  assign \new_[45000]_  = A167 & ~A168;
  assign \new_[45001]_  = ~A169 & \new_[45000]_ ;
  assign \new_[45004]_  = A199 & A166;
  assign \new_[45007]_  = ~A234 & A201;
  assign \new_[45008]_  = \new_[45007]_  & \new_[45004]_ ;
  assign \new_[45009]_  = \new_[45008]_  & \new_[45001]_ ;
  assign \new_[45013]_  = A265 & ~A236;
  assign \new_[45014]_  = ~A235 & \new_[45013]_ ;
  assign \new_[45017]_  = ~A267 & A266;
  assign \new_[45020]_  = A301 & ~A268;
  assign \new_[45021]_  = \new_[45020]_  & \new_[45017]_ ;
  assign \new_[45022]_  = \new_[45021]_  & \new_[45014]_ ;
  assign \new_[45026]_  = A167 & ~A168;
  assign \new_[45027]_  = ~A169 & \new_[45026]_ ;
  assign \new_[45030]_  = A199 & A166;
  assign \new_[45033]_  = ~A234 & A201;
  assign \new_[45034]_  = \new_[45033]_  & \new_[45030]_ ;
  assign \new_[45035]_  = \new_[45034]_  & \new_[45027]_ ;
  assign \new_[45039]_  = ~A265 & ~A236;
  assign \new_[45040]_  = ~A235 & \new_[45039]_ ;
  assign \new_[45043]_  = ~A268 & ~A266;
  assign \new_[45046]_  = A300 & A299;
  assign \new_[45047]_  = \new_[45046]_  & \new_[45043]_ ;
  assign \new_[45048]_  = \new_[45047]_  & \new_[45040]_ ;
  assign \new_[45052]_  = A167 & ~A168;
  assign \new_[45053]_  = ~A169 & \new_[45052]_ ;
  assign \new_[45056]_  = A199 & A166;
  assign \new_[45059]_  = ~A234 & A201;
  assign \new_[45060]_  = \new_[45059]_  & \new_[45056]_ ;
  assign \new_[45061]_  = \new_[45060]_  & \new_[45053]_ ;
  assign \new_[45065]_  = ~A265 & ~A236;
  assign \new_[45066]_  = ~A235 & \new_[45065]_ ;
  assign \new_[45069]_  = ~A268 & ~A266;
  assign \new_[45072]_  = A300 & A298;
  assign \new_[45073]_  = \new_[45072]_  & \new_[45069]_ ;
  assign \new_[45074]_  = \new_[45073]_  & \new_[45066]_ ;
  assign \new_[45078]_  = A167 & ~A168;
  assign \new_[45079]_  = ~A169 & \new_[45078]_ ;
  assign \new_[45082]_  = A199 & A166;
  assign \new_[45085]_  = A232 & A201;
  assign \new_[45086]_  = \new_[45085]_  & \new_[45082]_ ;
  assign \new_[45087]_  = \new_[45086]_  & \new_[45079]_ ;
  assign \new_[45091]_  = ~A235 & ~A234;
  assign \new_[45092]_  = A233 & \new_[45091]_ ;
  assign \new_[45095]_  = ~A268 & ~A267;
  assign \new_[45098]_  = A301 & ~A269;
  assign \new_[45099]_  = \new_[45098]_  & \new_[45095]_ ;
  assign \new_[45100]_  = \new_[45099]_  & \new_[45092]_ ;
  assign \new_[45104]_  = A167 & ~A168;
  assign \new_[45105]_  = ~A169 & \new_[45104]_ ;
  assign \new_[45108]_  = A199 & A166;
  assign \new_[45111]_  = A232 & A201;
  assign \new_[45112]_  = \new_[45111]_  & \new_[45108]_ ;
  assign \new_[45113]_  = \new_[45112]_  & \new_[45105]_ ;
  assign \new_[45117]_  = ~A235 & ~A234;
  assign \new_[45118]_  = A233 & \new_[45117]_ ;
  assign \new_[45121]_  = ~A266 & ~A265;
  assign \new_[45124]_  = A301 & ~A268;
  assign \new_[45125]_  = \new_[45124]_  & \new_[45121]_ ;
  assign \new_[45126]_  = \new_[45125]_  & \new_[45118]_ ;
  assign \new_[45130]_  = A167 & ~A168;
  assign \new_[45131]_  = ~A169 & \new_[45130]_ ;
  assign \new_[45134]_  = A199 & A166;
  assign \new_[45137]_  = ~A232 & A201;
  assign \new_[45138]_  = \new_[45137]_  & \new_[45134]_ ;
  assign \new_[45139]_  = \new_[45138]_  & \new_[45131]_ ;
  assign \new_[45143]_  = ~A267 & ~A235;
  assign \new_[45144]_  = ~A233 & \new_[45143]_ ;
  assign \new_[45147]_  = ~A269 & ~A268;
  assign \new_[45150]_  = A300 & A299;
  assign \new_[45151]_  = \new_[45150]_  & \new_[45147]_ ;
  assign \new_[45152]_  = \new_[45151]_  & \new_[45144]_ ;
  assign \new_[45156]_  = A167 & ~A168;
  assign \new_[45157]_  = ~A169 & \new_[45156]_ ;
  assign \new_[45160]_  = A199 & A166;
  assign \new_[45163]_  = ~A232 & A201;
  assign \new_[45164]_  = \new_[45163]_  & \new_[45160]_ ;
  assign \new_[45165]_  = \new_[45164]_  & \new_[45157]_ ;
  assign \new_[45169]_  = ~A267 & ~A235;
  assign \new_[45170]_  = ~A233 & \new_[45169]_ ;
  assign \new_[45173]_  = ~A269 & ~A268;
  assign \new_[45176]_  = A300 & A298;
  assign \new_[45177]_  = \new_[45176]_  & \new_[45173]_ ;
  assign \new_[45178]_  = \new_[45177]_  & \new_[45170]_ ;
  assign \new_[45182]_  = A167 & ~A168;
  assign \new_[45183]_  = ~A169 & \new_[45182]_ ;
  assign \new_[45186]_  = A199 & A166;
  assign \new_[45189]_  = ~A232 & A201;
  assign \new_[45190]_  = \new_[45189]_  & \new_[45186]_ ;
  assign \new_[45191]_  = \new_[45190]_  & \new_[45183]_ ;
  assign \new_[45195]_  = A265 & ~A235;
  assign \new_[45196]_  = ~A233 & \new_[45195]_ ;
  assign \new_[45199]_  = ~A267 & A266;
  assign \new_[45202]_  = A301 & ~A268;
  assign \new_[45203]_  = \new_[45202]_  & \new_[45199]_ ;
  assign \new_[45204]_  = \new_[45203]_  & \new_[45196]_ ;
  assign \new_[45208]_  = A167 & ~A168;
  assign \new_[45209]_  = ~A169 & \new_[45208]_ ;
  assign \new_[45212]_  = A199 & A166;
  assign \new_[45215]_  = ~A232 & A201;
  assign \new_[45216]_  = \new_[45215]_  & \new_[45212]_ ;
  assign \new_[45217]_  = \new_[45216]_  & \new_[45209]_ ;
  assign \new_[45221]_  = ~A265 & ~A235;
  assign \new_[45222]_  = ~A233 & \new_[45221]_ ;
  assign \new_[45225]_  = ~A268 & ~A266;
  assign \new_[45228]_  = A300 & A299;
  assign \new_[45229]_  = \new_[45228]_  & \new_[45225]_ ;
  assign \new_[45230]_  = \new_[45229]_  & \new_[45222]_ ;
  assign \new_[45234]_  = A167 & ~A168;
  assign \new_[45235]_  = ~A169 & \new_[45234]_ ;
  assign \new_[45238]_  = A199 & A166;
  assign \new_[45241]_  = ~A232 & A201;
  assign \new_[45242]_  = \new_[45241]_  & \new_[45238]_ ;
  assign \new_[45243]_  = \new_[45242]_  & \new_[45235]_ ;
  assign \new_[45247]_  = ~A265 & ~A235;
  assign \new_[45248]_  = ~A233 & \new_[45247]_ ;
  assign \new_[45251]_  = ~A268 & ~A266;
  assign \new_[45254]_  = A300 & A298;
  assign \new_[45255]_  = \new_[45254]_  & \new_[45251]_ ;
  assign \new_[45256]_  = \new_[45255]_  & \new_[45248]_ ;
  assign \new_[45260]_  = A167 & ~A168;
  assign \new_[45261]_  = ~A169 & \new_[45260]_ ;
  assign \new_[45264]_  = A200 & A166;
  assign \new_[45267]_  = ~A234 & A201;
  assign \new_[45268]_  = \new_[45267]_  & \new_[45264]_ ;
  assign \new_[45269]_  = \new_[45268]_  & \new_[45261]_ ;
  assign \new_[45273]_  = ~A267 & ~A236;
  assign \new_[45274]_  = ~A235 & \new_[45273]_ ;
  assign \new_[45277]_  = ~A269 & ~A268;
  assign \new_[45280]_  = A300 & A299;
  assign \new_[45281]_  = \new_[45280]_  & \new_[45277]_ ;
  assign \new_[45282]_  = \new_[45281]_  & \new_[45274]_ ;
  assign \new_[45286]_  = A167 & ~A168;
  assign \new_[45287]_  = ~A169 & \new_[45286]_ ;
  assign \new_[45290]_  = A200 & A166;
  assign \new_[45293]_  = ~A234 & A201;
  assign \new_[45294]_  = \new_[45293]_  & \new_[45290]_ ;
  assign \new_[45295]_  = \new_[45294]_  & \new_[45287]_ ;
  assign \new_[45299]_  = ~A267 & ~A236;
  assign \new_[45300]_  = ~A235 & \new_[45299]_ ;
  assign \new_[45303]_  = ~A269 & ~A268;
  assign \new_[45306]_  = A300 & A298;
  assign \new_[45307]_  = \new_[45306]_  & \new_[45303]_ ;
  assign \new_[45308]_  = \new_[45307]_  & \new_[45300]_ ;
  assign \new_[45312]_  = A167 & ~A168;
  assign \new_[45313]_  = ~A169 & \new_[45312]_ ;
  assign \new_[45316]_  = A200 & A166;
  assign \new_[45319]_  = ~A234 & A201;
  assign \new_[45320]_  = \new_[45319]_  & \new_[45316]_ ;
  assign \new_[45321]_  = \new_[45320]_  & \new_[45313]_ ;
  assign \new_[45325]_  = A265 & ~A236;
  assign \new_[45326]_  = ~A235 & \new_[45325]_ ;
  assign \new_[45329]_  = ~A267 & A266;
  assign \new_[45332]_  = A301 & ~A268;
  assign \new_[45333]_  = \new_[45332]_  & \new_[45329]_ ;
  assign \new_[45334]_  = \new_[45333]_  & \new_[45326]_ ;
  assign \new_[45338]_  = A167 & ~A168;
  assign \new_[45339]_  = ~A169 & \new_[45338]_ ;
  assign \new_[45342]_  = A200 & A166;
  assign \new_[45345]_  = ~A234 & A201;
  assign \new_[45346]_  = \new_[45345]_  & \new_[45342]_ ;
  assign \new_[45347]_  = \new_[45346]_  & \new_[45339]_ ;
  assign \new_[45351]_  = ~A265 & ~A236;
  assign \new_[45352]_  = ~A235 & \new_[45351]_ ;
  assign \new_[45355]_  = ~A268 & ~A266;
  assign \new_[45358]_  = A300 & A299;
  assign \new_[45359]_  = \new_[45358]_  & \new_[45355]_ ;
  assign \new_[45360]_  = \new_[45359]_  & \new_[45352]_ ;
  assign \new_[45364]_  = A167 & ~A168;
  assign \new_[45365]_  = ~A169 & \new_[45364]_ ;
  assign \new_[45368]_  = A200 & A166;
  assign \new_[45371]_  = ~A234 & A201;
  assign \new_[45372]_  = \new_[45371]_  & \new_[45368]_ ;
  assign \new_[45373]_  = \new_[45372]_  & \new_[45365]_ ;
  assign \new_[45377]_  = ~A265 & ~A236;
  assign \new_[45378]_  = ~A235 & \new_[45377]_ ;
  assign \new_[45381]_  = ~A268 & ~A266;
  assign \new_[45384]_  = A300 & A298;
  assign \new_[45385]_  = \new_[45384]_  & \new_[45381]_ ;
  assign \new_[45386]_  = \new_[45385]_  & \new_[45378]_ ;
  assign \new_[45390]_  = A167 & ~A168;
  assign \new_[45391]_  = ~A169 & \new_[45390]_ ;
  assign \new_[45394]_  = A200 & A166;
  assign \new_[45397]_  = A232 & A201;
  assign \new_[45398]_  = \new_[45397]_  & \new_[45394]_ ;
  assign \new_[45399]_  = \new_[45398]_  & \new_[45391]_ ;
  assign \new_[45403]_  = ~A235 & ~A234;
  assign \new_[45404]_  = A233 & \new_[45403]_ ;
  assign \new_[45407]_  = ~A268 & ~A267;
  assign \new_[45410]_  = A301 & ~A269;
  assign \new_[45411]_  = \new_[45410]_  & \new_[45407]_ ;
  assign \new_[45412]_  = \new_[45411]_  & \new_[45404]_ ;
  assign \new_[45416]_  = A167 & ~A168;
  assign \new_[45417]_  = ~A169 & \new_[45416]_ ;
  assign \new_[45420]_  = A200 & A166;
  assign \new_[45423]_  = A232 & A201;
  assign \new_[45424]_  = \new_[45423]_  & \new_[45420]_ ;
  assign \new_[45425]_  = \new_[45424]_  & \new_[45417]_ ;
  assign \new_[45429]_  = ~A235 & ~A234;
  assign \new_[45430]_  = A233 & \new_[45429]_ ;
  assign \new_[45433]_  = ~A266 & ~A265;
  assign \new_[45436]_  = A301 & ~A268;
  assign \new_[45437]_  = \new_[45436]_  & \new_[45433]_ ;
  assign \new_[45438]_  = \new_[45437]_  & \new_[45430]_ ;
  assign \new_[45442]_  = A167 & ~A168;
  assign \new_[45443]_  = ~A169 & \new_[45442]_ ;
  assign \new_[45446]_  = A200 & A166;
  assign \new_[45449]_  = ~A232 & A201;
  assign \new_[45450]_  = \new_[45449]_  & \new_[45446]_ ;
  assign \new_[45451]_  = \new_[45450]_  & \new_[45443]_ ;
  assign \new_[45455]_  = ~A267 & ~A235;
  assign \new_[45456]_  = ~A233 & \new_[45455]_ ;
  assign \new_[45459]_  = ~A269 & ~A268;
  assign \new_[45462]_  = A300 & A299;
  assign \new_[45463]_  = \new_[45462]_  & \new_[45459]_ ;
  assign \new_[45464]_  = \new_[45463]_  & \new_[45456]_ ;
  assign \new_[45468]_  = A167 & ~A168;
  assign \new_[45469]_  = ~A169 & \new_[45468]_ ;
  assign \new_[45472]_  = A200 & A166;
  assign \new_[45475]_  = ~A232 & A201;
  assign \new_[45476]_  = \new_[45475]_  & \new_[45472]_ ;
  assign \new_[45477]_  = \new_[45476]_  & \new_[45469]_ ;
  assign \new_[45481]_  = ~A267 & ~A235;
  assign \new_[45482]_  = ~A233 & \new_[45481]_ ;
  assign \new_[45485]_  = ~A269 & ~A268;
  assign \new_[45488]_  = A300 & A298;
  assign \new_[45489]_  = \new_[45488]_  & \new_[45485]_ ;
  assign \new_[45490]_  = \new_[45489]_  & \new_[45482]_ ;
  assign \new_[45494]_  = A167 & ~A168;
  assign \new_[45495]_  = ~A169 & \new_[45494]_ ;
  assign \new_[45498]_  = A200 & A166;
  assign \new_[45501]_  = ~A232 & A201;
  assign \new_[45502]_  = \new_[45501]_  & \new_[45498]_ ;
  assign \new_[45503]_  = \new_[45502]_  & \new_[45495]_ ;
  assign \new_[45507]_  = A265 & ~A235;
  assign \new_[45508]_  = ~A233 & \new_[45507]_ ;
  assign \new_[45511]_  = ~A267 & A266;
  assign \new_[45514]_  = A301 & ~A268;
  assign \new_[45515]_  = \new_[45514]_  & \new_[45511]_ ;
  assign \new_[45516]_  = \new_[45515]_  & \new_[45508]_ ;
  assign \new_[45520]_  = A167 & ~A168;
  assign \new_[45521]_  = ~A169 & \new_[45520]_ ;
  assign \new_[45524]_  = A200 & A166;
  assign \new_[45527]_  = ~A232 & A201;
  assign \new_[45528]_  = \new_[45527]_  & \new_[45524]_ ;
  assign \new_[45529]_  = \new_[45528]_  & \new_[45521]_ ;
  assign \new_[45533]_  = ~A265 & ~A235;
  assign \new_[45534]_  = ~A233 & \new_[45533]_ ;
  assign \new_[45537]_  = ~A268 & ~A266;
  assign \new_[45540]_  = A300 & A299;
  assign \new_[45541]_  = \new_[45540]_  & \new_[45537]_ ;
  assign \new_[45542]_  = \new_[45541]_  & \new_[45534]_ ;
  assign \new_[45546]_  = A167 & ~A168;
  assign \new_[45547]_  = ~A169 & \new_[45546]_ ;
  assign \new_[45550]_  = A200 & A166;
  assign \new_[45553]_  = ~A232 & A201;
  assign \new_[45554]_  = \new_[45553]_  & \new_[45550]_ ;
  assign \new_[45555]_  = \new_[45554]_  & \new_[45547]_ ;
  assign \new_[45559]_  = ~A265 & ~A235;
  assign \new_[45560]_  = ~A233 & \new_[45559]_ ;
  assign \new_[45563]_  = ~A268 & ~A266;
  assign \new_[45566]_  = A300 & A298;
  assign \new_[45567]_  = \new_[45566]_  & \new_[45563]_ ;
  assign \new_[45568]_  = \new_[45567]_  & \new_[45560]_ ;
  assign \new_[45572]_  = A167 & ~A168;
  assign \new_[45573]_  = ~A169 & \new_[45572]_ ;
  assign \new_[45576]_  = ~A199 & A166;
  assign \new_[45579]_  = A203 & A200;
  assign \new_[45580]_  = \new_[45579]_  & \new_[45576]_ ;
  assign \new_[45581]_  = \new_[45580]_  & \new_[45573]_ ;
  assign \new_[45585]_  = ~A236 & ~A235;
  assign \new_[45586]_  = ~A234 & \new_[45585]_ ;
  assign \new_[45589]_  = ~A268 & ~A267;
  assign \new_[45592]_  = A301 & ~A269;
  assign \new_[45593]_  = \new_[45592]_  & \new_[45589]_ ;
  assign \new_[45594]_  = \new_[45593]_  & \new_[45586]_ ;
  assign \new_[45598]_  = A167 & ~A168;
  assign \new_[45599]_  = ~A169 & \new_[45598]_ ;
  assign \new_[45602]_  = ~A199 & A166;
  assign \new_[45605]_  = A203 & A200;
  assign \new_[45606]_  = \new_[45605]_  & \new_[45602]_ ;
  assign \new_[45607]_  = \new_[45606]_  & \new_[45599]_ ;
  assign \new_[45611]_  = ~A236 & ~A235;
  assign \new_[45612]_  = ~A234 & \new_[45611]_ ;
  assign \new_[45615]_  = ~A266 & ~A265;
  assign \new_[45618]_  = A301 & ~A268;
  assign \new_[45619]_  = \new_[45618]_  & \new_[45615]_ ;
  assign \new_[45620]_  = \new_[45619]_  & \new_[45612]_ ;
  assign \new_[45624]_  = A167 & ~A168;
  assign \new_[45625]_  = ~A169 & \new_[45624]_ ;
  assign \new_[45628]_  = ~A199 & A166;
  assign \new_[45631]_  = A203 & A200;
  assign \new_[45632]_  = \new_[45631]_  & \new_[45628]_ ;
  assign \new_[45633]_  = \new_[45632]_  & \new_[45625]_ ;
  assign \new_[45637]_  = A236 & A233;
  assign \new_[45638]_  = ~A232 & \new_[45637]_ ;
  assign \new_[45641]_  = A299 & A298;
  assign \new_[45644]_  = ~A301 & ~A300;
  assign \new_[45645]_  = \new_[45644]_  & \new_[45641]_ ;
  assign \new_[45646]_  = \new_[45645]_  & \new_[45638]_ ;
  assign \new_[45650]_  = A167 & ~A168;
  assign \new_[45651]_  = ~A169 & \new_[45650]_ ;
  assign \new_[45654]_  = ~A199 & A166;
  assign \new_[45657]_  = A203 & A200;
  assign \new_[45658]_  = \new_[45657]_  & \new_[45654]_ ;
  assign \new_[45659]_  = \new_[45658]_  & \new_[45651]_ ;
  assign \new_[45663]_  = A236 & ~A233;
  assign \new_[45664]_  = A232 & \new_[45663]_ ;
  assign \new_[45667]_  = A299 & A298;
  assign \new_[45670]_  = ~A301 & ~A300;
  assign \new_[45671]_  = \new_[45670]_  & \new_[45667]_ ;
  assign \new_[45672]_  = \new_[45671]_  & \new_[45664]_ ;
  assign \new_[45676]_  = A167 & ~A168;
  assign \new_[45677]_  = ~A169 & \new_[45676]_ ;
  assign \new_[45680]_  = ~A199 & A166;
  assign \new_[45683]_  = A203 & A200;
  assign \new_[45684]_  = \new_[45683]_  & \new_[45680]_ ;
  assign \new_[45685]_  = \new_[45684]_  & \new_[45677]_ ;
  assign \new_[45689]_  = ~A235 & ~A233;
  assign \new_[45690]_  = ~A232 & \new_[45689]_ ;
  assign \new_[45693]_  = ~A268 & ~A267;
  assign \new_[45696]_  = A301 & ~A269;
  assign \new_[45697]_  = \new_[45696]_  & \new_[45693]_ ;
  assign \new_[45698]_  = \new_[45697]_  & \new_[45690]_ ;
  assign \new_[45702]_  = A167 & ~A168;
  assign \new_[45703]_  = ~A169 & \new_[45702]_ ;
  assign \new_[45706]_  = ~A199 & A166;
  assign \new_[45709]_  = A203 & A200;
  assign \new_[45710]_  = \new_[45709]_  & \new_[45706]_ ;
  assign \new_[45711]_  = \new_[45710]_  & \new_[45703]_ ;
  assign \new_[45715]_  = ~A235 & ~A233;
  assign \new_[45716]_  = ~A232 & \new_[45715]_ ;
  assign \new_[45719]_  = ~A266 & ~A265;
  assign \new_[45722]_  = A301 & ~A268;
  assign \new_[45723]_  = \new_[45722]_  & \new_[45719]_ ;
  assign \new_[45724]_  = \new_[45723]_  & \new_[45716]_ ;
  assign \new_[45728]_  = A167 & ~A168;
  assign \new_[45729]_  = ~A169 & \new_[45728]_ ;
  assign \new_[45732]_  = A199 & A166;
  assign \new_[45735]_  = A203 & ~A200;
  assign \new_[45736]_  = \new_[45735]_  & \new_[45732]_ ;
  assign \new_[45737]_  = \new_[45736]_  & \new_[45729]_ ;
  assign \new_[45741]_  = ~A236 & ~A235;
  assign \new_[45742]_  = ~A234 & \new_[45741]_ ;
  assign \new_[45745]_  = ~A268 & ~A267;
  assign \new_[45748]_  = A301 & ~A269;
  assign \new_[45749]_  = \new_[45748]_  & \new_[45745]_ ;
  assign \new_[45750]_  = \new_[45749]_  & \new_[45742]_ ;
  assign \new_[45754]_  = A167 & ~A168;
  assign \new_[45755]_  = ~A169 & \new_[45754]_ ;
  assign \new_[45758]_  = A199 & A166;
  assign \new_[45761]_  = A203 & ~A200;
  assign \new_[45762]_  = \new_[45761]_  & \new_[45758]_ ;
  assign \new_[45763]_  = \new_[45762]_  & \new_[45755]_ ;
  assign \new_[45767]_  = ~A236 & ~A235;
  assign \new_[45768]_  = ~A234 & \new_[45767]_ ;
  assign \new_[45771]_  = ~A266 & ~A265;
  assign \new_[45774]_  = A301 & ~A268;
  assign \new_[45775]_  = \new_[45774]_  & \new_[45771]_ ;
  assign \new_[45776]_  = \new_[45775]_  & \new_[45768]_ ;
  assign \new_[45780]_  = A167 & ~A168;
  assign \new_[45781]_  = ~A169 & \new_[45780]_ ;
  assign \new_[45784]_  = A199 & A166;
  assign \new_[45787]_  = A203 & ~A200;
  assign \new_[45788]_  = \new_[45787]_  & \new_[45784]_ ;
  assign \new_[45789]_  = \new_[45788]_  & \new_[45781]_ ;
  assign \new_[45793]_  = A236 & A233;
  assign \new_[45794]_  = ~A232 & \new_[45793]_ ;
  assign \new_[45797]_  = A299 & A298;
  assign \new_[45800]_  = ~A301 & ~A300;
  assign \new_[45801]_  = \new_[45800]_  & \new_[45797]_ ;
  assign \new_[45802]_  = \new_[45801]_  & \new_[45794]_ ;
  assign \new_[45806]_  = A167 & ~A168;
  assign \new_[45807]_  = ~A169 & \new_[45806]_ ;
  assign \new_[45810]_  = A199 & A166;
  assign \new_[45813]_  = A203 & ~A200;
  assign \new_[45814]_  = \new_[45813]_  & \new_[45810]_ ;
  assign \new_[45815]_  = \new_[45814]_  & \new_[45807]_ ;
  assign \new_[45819]_  = A236 & ~A233;
  assign \new_[45820]_  = A232 & \new_[45819]_ ;
  assign \new_[45823]_  = A299 & A298;
  assign \new_[45826]_  = ~A301 & ~A300;
  assign \new_[45827]_  = \new_[45826]_  & \new_[45823]_ ;
  assign \new_[45828]_  = \new_[45827]_  & \new_[45820]_ ;
  assign \new_[45832]_  = A167 & ~A168;
  assign \new_[45833]_  = ~A169 & \new_[45832]_ ;
  assign \new_[45836]_  = A199 & A166;
  assign \new_[45839]_  = A203 & ~A200;
  assign \new_[45840]_  = \new_[45839]_  & \new_[45836]_ ;
  assign \new_[45841]_  = \new_[45840]_  & \new_[45833]_ ;
  assign \new_[45845]_  = ~A235 & ~A233;
  assign \new_[45846]_  = ~A232 & \new_[45845]_ ;
  assign \new_[45849]_  = ~A268 & ~A267;
  assign \new_[45852]_  = A301 & ~A269;
  assign \new_[45853]_  = \new_[45852]_  & \new_[45849]_ ;
  assign \new_[45854]_  = \new_[45853]_  & \new_[45846]_ ;
  assign \new_[45858]_  = A167 & ~A168;
  assign \new_[45859]_  = ~A169 & \new_[45858]_ ;
  assign \new_[45862]_  = A199 & A166;
  assign \new_[45865]_  = A203 & ~A200;
  assign \new_[45866]_  = \new_[45865]_  & \new_[45862]_ ;
  assign \new_[45867]_  = \new_[45866]_  & \new_[45859]_ ;
  assign \new_[45871]_  = ~A235 & ~A233;
  assign \new_[45872]_  = ~A232 & \new_[45871]_ ;
  assign \new_[45875]_  = ~A266 & ~A265;
  assign \new_[45878]_  = A301 & ~A268;
  assign \new_[45879]_  = \new_[45878]_  & \new_[45875]_ ;
  assign \new_[45880]_  = \new_[45879]_  & \new_[45872]_ ;
  assign \new_[45884]_  = ~A168 & ~A169;
  assign \new_[45885]_  = ~A170 & \new_[45884]_ ;
  assign \new_[45888]_  = ~A234 & A202;
  assign \new_[45891]_  = ~A236 & ~A235;
  assign \new_[45892]_  = \new_[45891]_  & \new_[45888]_ ;
  assign \new_[45893]_  = \new_[45892]_  & \new_[45885]_ ;
  assign \new_[45897]_  = ~A267 & A266;
  assign \new_[45898]_  = A265 & \new_[45897]_ ;
  assign \new_[45901]_  = A298 & ~A268;
  assign \new_[45904]_  = A302 & ~A299;
  assign \new_[45905]_  = \new_[45904]_  & \new_[45901]_ ;
  assign \new_[45906]_  = \new_[45905]_  & \new_[45898]_ ;
  assign \new_[45910]_  = ~A168 & ~A169;
  assign \new_[45911]_  = ~A170 & \new_[45910]_ ;
  assign \new_[45914]_  = ~A234 & A202;
  assign \new_[45917]_  = ~A236 & ~A235;
  assign \new_[45918]_  = \new_[45917]_  & \new_[45914]_ ;
  assign \new_[45919]_  = \new_[45918]_  & \new_[45911]_ ;
  assign \new_[45923]_  = ~A267 & A266;
  assign \new_[45924]_  = A265 & \new_[45923]_ ;
  assign \new_[45927]_  = ~A298 & ~A268;
  assign \new_[45930]_  = A302 & A299;
  assign \new_[45931]_  = \new_[45930]_  & \new_[45927]_ ;
  assign \new_[45932]_  = \new_[45931]_  & \new_[45924]_ ;
  assign \new_[45936]_  = ~A168 & ~A169;
  assign \new_[45937]_  = ~A170 & \new_[45936]_ ;
  assign \new_[45940]_  = A232 & A202;
  assign \new_[45943]_  = ~A234 & A233;
  assign \new_[45944]_  = \new_[45943]_  & \new_[45940]_ ;
  assign \new_[45945]_  = \new_[45944]_  & \new_[45937]_ ;
  assign \new_[45949]_  = ~A268 & ~A267;
  assign \new_[45950]_  = ~A235 & \new_[45949]_ ;
  assign \new_[45953]_  = A298 & ~A269;
  assign \new_[45956]_  = A302 & ~A299;
  assign \new_[45957]_  = \new_[45956]_  & \new_[45953]_ ;
  assign \new_[45958]_  = \new_[45957]_  & \new_[45950]_ ;
  assign \new_[45962]_  = ~A168 & ~A169;
  assign \new_[45963]_  = ~A170 & \new_[45962]_ ;
  assign \new_[45966]_  = A232 & A202;
  assign \new_[45969]_  = ~A234 & A233;
  assign \new_[45970]_  = \new_[45969]_  & \new_[45966]_ ;
  assign \new_[45971]_  = \new_[45970]_  & \new_[45963]_ ;
  assign \new_[45975]_  = ~A268 & ~A267;
  assign \new_[45976]_  = ~A235 & \new_[45975]_ ;
  assign \new_[45979]_  = ~A298 & ~A269;
  assign \new_[45982]_  = A302 & A299;
  assign \new_[45983]_  = \new_[45982]_  & \new_[45979]_ ;
  assign \new_[45984]_  = \new_[45983]_  & \new_[45976]_ ;
  assign \new_[45988]_  = ~A168 & ~A169;
  assign \new_[45989]_  = ~A170 & \new_[45988]_ ;
  assign \new_[45992]_  = A232 & A202;
  assign \new_[45995]_  = ~A234 & A233;
  assign \new_[45996]_  = \new_[45995]_  & \new_[45992]_ ;
  assign \new_[45997]_  = \new_[45996]_  & \new_[45989]_ ;
  assign \new_[46001]_  = A266 & A265;
  assign \new_[46002]_  = ~A235 & \new_[46001]_ ;
  assign \new_[46005]_  = ~A268 & ~A267;
  assign \new_[46008]_  = A300 & A299;
  assign \new_[46009]_  = \new_[46008]_  & \new_[46005]_ ;
  assign \new_[46010]_  = \new_[46009]_  & \new_[46002]_ ;
  assign \new_[46014]_  = ~A168 & ~A169;
  assign \new_[46015]_  = ~A170 & \new_[46014]_ ;
  assign \new_[46018]_  = A232 & A202;
  assign \new_[46021]_  = ~A234 & A233;
  assign \new_[46022]_  = \new_[46021]_  & \new_[46018]_ ;
  assign \new_[46023]_  = \new_[46022]_  & \new_[46015]_ ;
  assign \new_[46027]_  = A266 & A265;
  assign \new_[46028]_  = ~A235 & \new_[46027]_ ;
  assign \new_[46031]_  = ~A268 & ~A267;
  assign \new_[46034]_  = A300 & A298;
  assign \new_[46035]_  = \new_[46034]_  & \new_[46031]_ ;
  assign \new_[46036]_  = \new_[46035]_  & \new_[46028]_ ;
  assign \new_[46040]_  = ~A168 & ~A169;
  assign \new_[46041]_  = ~A170 & \new_[46040]_ ;
  assign \new_[46044]_  = A232 & A202;
  assign \new_[46047]_  = ~A234 & A233;
  assign \new_[46048]_  = \new_[46047]_  & \new_[46044]_ ;
  assign \new_[46049]_  = \new_[46048]_  & \new_[46041]_ ;
  assign \new_[46053]_  = ~A266 & ~A265;
  assign \new_[46054]_  = ~A235 & \new_[46053]_ ;
  assign \new_[46057]_  = A298 & ~A268;
  assign \new_[46060]_  = A302 & ~A299;
  assign \new_[46061]_  = \new_[46060]_  & \new_[46057]_ ;
  assign \new_[46062]_  = \new_[46061]_  & \new_[46054]_ ;
  assign \new_[46066]_  = ~A168 & ~A169;
  assign \new_[46067]_  = ~A170 & \new_[46066]_ ;
  assign \new_[46070]_  = A232 & A202;
  assign \new_[46073]_  = ~A234 & A233;
  assign \new_[46074]_  = \new_[46073]_  & \new_[46070]_ ;
  assign \new_[46075]_  = \new_[46074]_  & \new_[46067]_ ;
  assign \new_[46079]_  = ~A266 & ~A265;
  assign \new_[46080]_  = ~A235 & \new_[46079]_ ;
  assign \new_[46083]_  = ~A298 & ~A268;
  assign \new_[46086]_  = A302 & A299;
  assign \new_[46087]_  = \new_[46086]_  & \new_[46083]_ ;
  assign \new_[46088]_  = \new_[46087]_  & \new_[46080]_ ;
  assign \new_[46092]_  = ~A168 & ~A169;
  assign \new_[46093]_  = ~A170 & \new_[46092]_ ;
  assign \new_[46096]_  = ~A232 & A202;
  assign \new_[46099]_  = ~A235 & ~A233;
  assign \new_[46100]_  = \new_[46099]_  & \new_[46096]_ ;
  assign \new_[46101]_  = \new_[46100]_  & \new_[46093]_ ;
  assign \new_[46105]_  = ~A267 & A266;
  assign \new_[46106]_  = A265 & \new_[46105]_ ;
  assign \new_[46109]_  = A298 & ~A268;
  assign \new_[46112]_  = A302 & ~A299;
  assign \new_[46113]_  = \new_[46112]_  & \new_[46109]_ ;
  assign \new_[46114]_  = \new_[46113]_  & \new_[46106]_ ;
  assign \new_[46118]_  = ~A168 & ~A169;
  assign \new_[46119]_  = ~A170 & \new_[46118]_ ;
  assign \new_[46122]_  = ~A232 & A202;
  assign \new_[46125]_  = ~A235 & ~A233;
  assign \new_[46126]_  = \new_[46125]_  & \new_[46122]_ ;
  assign \new_[46127]_  = \new_[46126]_  & \new_[46119]_ ;
  assign \new_[46131]_  = ~A267 & A266;
  assign \new_[46132]_  = A265 & \new_[46131]_ ;
  assign \new_[46135]_  = ~A298 & ~A268;
  assign \new_[46138]_  = A302 & A299;
  assign \new_[46139]_  = \new_[46138]_  & \new_[46135]_ ;
  assign \new_[46140]_  = \new_[46139]_  & \new_[46132]_ ;
  assign \new_[46144]_  = ~A168 & ~A169;
  assign \new_[46145]_  = ~A170 & \new_[46144]_ ;
  assign \new_[46148]_  = A201 & A199;
  assign \new_[46151]_  = ~A235 & ~A234;
  assign \new_[46152]_  = \new_[46151]_  & \new_[46148]_ ;
  assign \new_[46153]_  = \new_[46152]_  & \new_[46145]_ ;
  assign \new_[46157]_  = ~A268 & ~A267;
  assign \new_[46158]_  = ~A236 & \new_[46157]_ ;
  assign \new_[46161]_  = A298 & ~A269;
  assign \new_[46164]_  = A302 & ~A299;
  assign \new_[46165]_  = \new_[46164]_  & \new_[46161]_ ;
  assign \new_[46166]_  = \new_[46165]_  & \new_[46158]_ ;
  assign \new_[46170]_  = ~A168 & ~A169;
  assign \new_[46171]_  = ~A170 & \new_[46170]_ ;
  assign \new_[46174]_  = A201 & A199;
  assign \new_[46177]_  = ~A235 & ~A234;
  assign \new_[46178]_  = \new_[46177]_  & \new_[46174]_ ;
  assign \new_[46179]_  = \new_[46178]_  & \new_[46171]_ ;
  assign \new_[46183]_  = ~A268 & ~A267;
  assign \new_[46184]_  = ~A236 & \new_[46183]_ ;
  assign \new_[46187]_  = ~A298 & ~A269;
  assign \new_[46190]_  = A302 & A299;
  assign \new_[46191]_  = \new_[46190]_  & \new_[46187]_ ;
  assign \new_[46192]_  = \new_[46191]_  & \new_[46184]_ ;
  assign \new_[46196]_  = ~A168 & ~A169;
  assign \new_[46197]_  = ~A170 & \new_[46196]_ ;
  assign \new_[46200]_  = A201 & A199;
  assign \new_[46203]_  = ~A235 & ~A234;
  assign \new_[46204]_  = \new_[46203]_  & \new_[46200]_ ;
  assign \new_[46205]_  = \new_[46204]_  & \new_[46197]_ ;
  assign \new_[46209]_  = A266 & A265;
  assign \new_[46210]_  = ~A236 & \new_[46209]_ ;
  assign \new_[46213]_  = ~A268 & ~A267;
  assign \new_[46216]_  = A300 & A299;
  assign \new_[46217]_  = \new_[46216]_  & \new_[46213]_ ;
  assign \new_[46218]_  = \new_[46217]_  & \new_[46210]_ ;
  assign \new_[46222]_  = ~A168 & ~A169;
  assign \new_[46223]_  = ~A170 & \new_[46222]_ ;
  assign \new_[46226]_  = A201 & A199;
  assign \new_[46229]_  = ~A235 & ~A234;
  assign \new_[46230]_  = \new_[46229]_  & \new_[46226]_ ;
  assign \new_[46231]_  = \new_[46230]_  & \new_[46223]_ ;
  assign \new_[46235]_  = A266 & A265;
  assign \new_[46236]_  = ~A236 & \new_[46235]_ ;
  assign \new_[46239]_  = ~A268 & ~A267;
  assign \new_[46242]_  = A300 & A298;
  assign \new_[46243]_  = \new_[46242]_  & \new_[46239]_ ;
  assign \new_[46244]_  = \new_[46243]_  & \new_[46236]_ ;
  assign \new_[46248]_  = ~A168 & ~A169;
  assign \new_[46249]_  = ~A170 & \new_[46248]_ ;
  assign \new_[46252]_  = A201 & A199;
  assign \new_[46255]_  = ~A235 & ~A234;
  assign \new_[46256]_  = \new_[46255]_  & \new_[46252]_ ;
  assign \new_[46257]_  = \new_[46256]_  & \new_[46249]_ ;
  assign \new_[46261]_  = ~A266 & ~A265;
  assign \new_[46262]_  = ~A236 & \new_[46261]_ ;
  assign \new_[46265]_  = A298 & ~A268;
  assign \new_[46268]_  = A302 & ~A299;
  assign \new_[46269]_  = \new_[46268]_  & \new_[46265]_ ;
  assign \new_[46270]_  = \new_[46269]_  & \new_[46262]_ ;
  assign \new_[46274]_  = ~A168 & ~A169;
  assign \new_[46275]_  = ~A170 & \new_[46274]_ ;
  assign \new_[46278]_  = A201 & A199;
  assign \new_[46281]_  = ~A235 & ~A234;
  assign \new_[46282]_  = \new_[46281]_  & \new_[46278]_ ;
  assign \new_[46283]_  = \new_[46282]_  & \new_[46275]_ ;
  assign \new_[46287]_  = ~A266 & ~A265;
  assign \new_[46288]_  = ~A236 & \new_[46287]_ ;
  assign \new_[46291]_  = ~A298 & ~A268;
  assign \new_[46294]_  = A302 & A299;
  assign \new_[46295]_  = \new_[46294]_  & \new_[46291]_ ;
  assign \new_[46296]_  = \new_[46295]_  & \new_[46288]_ ;
  assign \new_[46300]_  = ~A168 & ~A169;
  assign \new_[46301]_  = ~A170 & \new_[46300]_ ;
  assign \new_[46304]_  = A201 & A199;
  assign \new_[46307]_  = A233 & A232;
  assign \new_[46308]_  = \new_[46307]_  & \new_[46304]_ ;
  assign \new_[46309]_  = \new_[46308]_  & \new_[46301]_ ;
  assign \new_[46313]_  = ~A267 & ~A235;
  assign \new_[46314]_  = ~A234 & \new_[46313]_ ;
  assign \new_[46317]_  = ~A269 & ~A268;
  assign \new_[46320]_  = A300 & A299;
  assign \new_[46321]_  = \new_[46320]_  & \new_[46317]_ ;
  assign \new_[46322]_  = \new_[46321]_  & \new_[46314]_ ;
  assign \new_[46326]_  = ~A168 & ~A169;
  assign \new_[46327]_  = ~A170 & \new_[46326]_ ;
  assign \new_[46330]_  = A201 & A199;
  assign \new_[46333]_  = A233 & A232;
  assign \new_[46334]_  = \new_[46333]_  & \new_[46330]_ ;
  assign \new_[46335]_  = \new_[46334]_  & \new_[46327]_ ;
  assign \new_[46339]_  = ~A267 & ~A235;
  assign \new_[46340]_  = ~A234 & \new_[46339]_ ;
  assign \new_[46343]_  = ~A269 & ~A268;
  assign \new_[46346]_  = A300 & A298;
  assign \new_[46347]_  = \new_[46346]_  & \new_[46343]_ ;
  assign \new_[46348]_  = \new_[46347]_  & \new_[46340]_ ;
  assign \new_[46352]_  = ~A168 & ~A169;
  assign \new_[46353]_  = ~A170 & \new_[46352]_ ;
  assign \new_[46356]_  = A201 & A199;
  assign \new_[46359]_  = A233 & A232;
  assign \new_[46360]_  = \new_[46359]_  & \new_[46356]_ ;
  assign \new_[46361]_  = \new_[46360]_  & \new_[46353]_ ;
  assign \new_[46365]_  = A265 & ~A235;
  assign \new_[46366]_  = ~A234 & \new_[46365]_ ;
  assign \new_[46369]_  = ~A267 & A266;
  assign \new_[46372]_  = A301 & ~A268;
  assign \new_[46373]_  = \new_[46372]_  & \new_[46369]_ ;
  assign \new_[46374]_  = \new_[46373]_  & \new_[46366]_ ;
  assign \new_[46378]_  = ~A168 & ~A169;
  assign \new_[46379]_  = ~A170 & \new_[46378]_ ;
  assign \new_[46382]_  = A201 & A199;
  assign \new_[46385]_  = A233 & A232;
  assign \new_[46386]_  = \new_[46385]_  & \new_[46382]_ ;
  assign \new_[46387]_  = \new_[46386]_  & \new_[46379]_ ;
  assign \new_[46391]_  = ~A265 & ~A235;
  assign \new_[46392]_  = ~A234 & \new_[46391]_ ;
  assign \new_[46395]_  = ~A268 & ~A266;
  assign \new_[46398]_  = A300 & A299;
  assign \new_[46399]_  = \new_[46398]_  & \new_[46395]_ ;
  assign \new_[46400]_  = \new_[46399]_  & \new_[46392]_ ;
  assign \new_[46404]_  = ~A168 & ~A169;
  assign \new_[46405]_  = ~A170 & \new_[46404]_ ;
  assign \new_[46408]_  = A201 & A199;
  assign \new_[46411]_  = A233 & A232;
  assign \new_[46412]_  = \new_[46411]_  & \new_[46408]_ ;
  assign \new_[46413]_  = \new_[46412]_  & \new_[46405]_ ;
  assign \new_[46417]_  = ~A265 & ~A235;
  assign \new_[46418]_  = ~A234 & \new_[46417]_ ;
  assign \new_[46421]_  = ~A268 & ~A266;
  assign \new_[46424]_  = A300 & A298;
  assign \new_[46425]_  = \new_[46424]_  & \new_[46421]_ ;
  assign \new_[46426]_  = \new_[46425]_  & \new_[46418]_ ;
  assign \new_[46430]_  = ~A168 & ~A169;
  assign \new_[46431]_  = ~A170 & \new_[46430]_ ;
  assign \new_[46434]_  = A201 & A199;
  assign \new_[46437]_  = ~A233 & ~A232;
  assign \new_[46438]_  = \new_[46437]_  & \new_[46434]_ ;
  assign \new_[46439]_  = \new_[46438]_  & \new_[46431]_ ;
  assign \new_[46443]_  = ~A268 & ~A267;
  assign \new_[46444]_  = ~A235 & \new_[46443]_ ;
  assign \new_[46447]_  = A298 & ~A269;
  assign \new_[46450]_  = A302 & ~A299;
  assign \new_[46451]_  = \new_[46450]_  & \new_[46447]_ ;
  assign \new_[46452]_  = \new_[46451]_  & \new_[46444]_ ;
  assign \new_[46456]_  = ~A168 & ~A169;
  assign \new_[46457]_  = ~A170 & \new_[46456]_ ;
  assign \new_[46460]_  = A201 & A199;
  assign \new_[46463]_  = ~A233 & ~A232;
  assign \new_[46464]_  = \new_[46463]_  & \new_[46460]_ ;
  assign \new_[46465]_  = \new_[46464]_  & \new_[46457]_ ;
  assign \new_[46469]_  = ~A268 & ~A267;
  assign \new_[46470]_  = ~A235 & \new_[46469]_ ;
  assign \new_[46473]_  = ~A298 & ~A269;
  assign \new_[46476]_  = A302 & A299;
  assign \new_[46477]_  = \new_[46476]_  & \new_[46473]_ ;
  assign \new_[46478]_  = \new_[46477]_  & \new_[46470]_ ;
  assign \new_[46482]_  = ~A168 & ~A169;
  assign \new_[46483]_  = ~A170 & \new_[46482]_ ;
  assign \new_[46486]_  = A201 & A199;
  assign \new_[46489]_  = ~A233 & ~A232;
  assign \new_[46490]_  = \new_[46489]_  & \new_[46486]_ ;
  assign \new_[46491]_  = \new_[46490]_  & \new_[46483]_ ;
  assign \new_[46495]_  = A266 & A265;
  assign \new_[46496]_  = ~A235 & \new_[46495]_ ;
  assign \new_[46499]_  = ~A268 & ~A267;
  assign \new_[46502]_  = A300 & A299;
  assign \new_[46503]_  = \new_[46502]_  & \new_[46499]_ ;
  assign \new_[46504]_  = \new_[46503]_  & \new_[46496]_ ;
  assign \new_[46508]_  = ~A168 & ~A169;
  assign \new_[46509]_  = ~A170 & \new_[46508]_ ;
  assign \new_[46512]_  = A201 & A199;
  assign \new_[46515]_  = ~A233 & ~A232;
  assign \new_[46516]_  = \new_[46515]_  & \new_[46512]_ ;
  assign \new_[46517]_  = \new_[46516]_  & \new_[46509]_ ;
  assign \new_[46521]_  = A266 & A265;
  assign \new_[46522]_  = ~A235 & \new_[46521]_ ;
  assign \new_[46525]_  = ~A268 & ~A267;
  assign \new_[46528]_  = A300 & A298;
  assign \new_[46529]_  = \new_[46528]_  & \new_[46525]_ ;
  assign \new_[46530]_  = \new_[46529]_  & \new_[46522]_ ;
  assign \new_[46534]_  = ~A168 & ~A169;
  assign \new_[46535]_  = ~A170 & \new_[46534]_ ;
  assign \new_[46538]_  = A201 & A199;
  assign \new_[46541]_  = ~A233 & ~A232;
  assign \new_[46542]_  = \new_[46541]_  & \new_[46538]_ ;
  assign \new_[46543]_  = \new_[46542]_  & \new_[46535]_ ;
  assign \new_[46547]_  = ~A266 & ~A265;
  assign \new_[46548]_  = ~A235 & \new_[46547]_ ;
  assign \new_[46551]_  = A298 & ~A268;
  assign \new_[46554]_  = A302 & ~A299;
  assign \new_[46555]_  = \new_[46554]_  & \new_[46551]_ ;
  assign \new_[46556]_  = \new_[46555]_  & \new_[46548]_ ;
  assign \new_[46560]_  = ~A168 & ~A169;
  assign \new_[46561]_  = ~A170 & \new_[46560]_ ;
  assign \new_[46564]_  = A201 & A199;
  assign \new_[46567]_  = ~A233 & ~A232;
  assign \new_[46568]_  = \new_[46567]_  & \new_[46564]_ ;
  assign \new_[46569]_  = \new_[46568]_  & \new_[46561]_ ;
  assign \new_[46573]_  = ~A266 & ~A265;
  assign \new_[46574]_  = ~A235 & \new_[46573]_ ;
  assign \new_[46577]_  = ~A298 & ~A268;
  assign \new_[46580]_  = A302 & A299;
  assign \new_[46581]_  = \new_[46580]_  & \new_[46577]_ ;
  assign \new_[46582]_  = \new_[46581]_  & \new_[46574]_ ;
  assign \new_[46586]_  = ~A168 & ~A169;
  assign \new_[46587]_  = ~A170 & \new_[46586]_ ;
  assign \new_[46590]_  = A201 & A200;
  assign \new_[46593]_  = ~A235 & ~A234;
  assign \new_[46594]_  = \new_[46593]_  & \new_[46590]_ ;
  assign \new_[46595]_  = \new_[46594]_  & \new_[46587]_ ;
  assign \new_[46599]_  = ~A268 & ~A267;
  assign \new_[46600]_  = ~A236 & \new_[46599]_ ;
  assign \new_[46603]_  = A298 & ~A269;
  assign \new_[46606]_  = A302 & ~A299;
  assign \new_[46607]_  = \new_[46606]_  & \new_[46603]_ ;
  assign \new_[46608]_  = \new_[46607]_  & \new_[46600]_ ;
  assign \new_[46612]_  = ~A168 & ~A169;
  assign \new_[46613]_  = ~A170 & \new_[46612]_ ;
  assign \new_[46616]_  = A201 & A200;
  assign \new_[46619]_  = ~A235 & ~A234;
  assign \new_[46620]_  = \new_[46619]_  & \new_[46616]_ ;
  assign \new_[46621]_  = \new_[46620]_  & \new_[46613]_ ;
  assign \new_[46625]_  = ~A268 & ~A267;
  assign \new_[46626]_  = ~A236 & \new_[46625]_ ;
  assign \new_[46629]_  = ~A298 & ~A269;
  assign \new_[46632]_  = A302 & A299;
  assign \new_[46633]_  = \new_[46632]_  & \new_[46629]_ ;
  assign \new_[46634]_  = \new_[46633]_  & \new_[46626]_ ;
  assign \new_[46638]_  = ~A168 & ~A169;
  assign \new_[46639]_  = ~A170 & \new_[46638]_ ;
  assign \new_[46642]_  = A201 & A200;
  assign \new_[46645]_  = ~A235 & ~A234;
  assign \new_[46646]_  = \new_[46645]_  & \new_[46642]_ ;
  assign \new_[46647]_  = \new_[46646]_  & \new_[46639]_ ;
  assign \new_[46651]_  = A266 & A265;
  assign \new_[46652]_  = ~A236 & \new_[46651]_ ;
  assign \new_[46655]_  = ~A268 & ~A267;
  assign \new_[46658]_  = A300 & A299;
  assign \new_[46659]_  = \new_[46658]_  & \new_[46655]_ ;
  assign \new_[46660]_  = \new_[46659]_  & \new_[46652]_ ;
  assign \new_[46664]_  = ~A168 & ~A169;
  assign \new_[46665]_  = ~A170 & \new_[46664]_ ;
  assign \new_[46668]_  = A201 & A200;
  assign \new_[46671]_  = ~A235 & ~A234;
  assign \new_[46672]_  = \new_[46671]_  & \new_[46668]_ ;
  assign \new_[46673]_  = \new_[46672]_  & \new_[46665]_ ;
  assign \new_[46677]_  = A266 & A265;
  assign \new_[46678]_  = ~A236 & \new_[46677]_ ;
  assign \new_[46681]_  = ~A268 & ~A267;
  assign \new_[46684]_  = A300 & A298;
  assign \new_[46685]_  = \new_[46684]_  & \new_[46681]_ ;
  assign \new_[46686]_  = \new_[46685]_  & \new_[46678]_ ;
  assign \new_[46690]_  = ~A168 & ~A169;
  assign \new_[46691]_  = ~A170 & \new_[46690]_ ;
  assign \new_[46694]_  = A201 & A200;
  assign \new_[46697]_  = ~A235 & ~A234;
  assign \new_[46698]_  = \new_[46697]_  & \new_[46694]_ ;
  assign \new_[46699]_  = \new_[46698]_  & \new_[46691]_ ;
  assign \new_[46703]_  = ~A266 & ~A265;
  assign \new_[46704]_  = ~A236 & \new_[46703]_ ;
  assign \new_[46707]_  = A298 & ~A268;
  assign \new_[46710]_  = A302 & ~A299;
  assign \new_[46711]_  = \new_[46710]_  & \new_[46707]_ ;
  assign \new_[46712]_  = \new_[46711]_  & \new_[46704]_ ;
  assign \new_[46716]_  = ~A168 & ~A169;
  assign \new_[46717]_  = ~A170 & \new_[46716]_ ;
  assign \new_[46720]_  = A201 & A200;
  assign \new_[46723]_  = ~A235 & ~A234;
  assign \new_[46724]_  = \new_[46723]_  & \new_[46720]_ ;
  assign \new_[46725]_  = \new_[46724]_  & \new_[46717]_ ;
  assign \new_[46729]_  = ~A266 & ~A265;
  assign \new_[46730]_  = ~A236 & \new_[46729]_ ;
  assign \new_[46733]_  = ~A298 & ~A268;
  assign \new_[46736]_  = A302 & A299;
  assign \new_[46737]_  = \new_[46736]_  & \new_[46733]_ ;
  assign \new_[46738]_  = \new_[46737]_  & \new_[46730]_ ;
  assign \new_[46742]_  = ~A168 & ~A169;
  assign \new_[46743]_  = ~A170 & \new_[46742]_ ;
  assign \new_[46746]_  = A201 & A200;
  assign \new_[46749]_  = A233 & A232;
  assign \new_[46750]_  = \new_[46749]_  & \new_[46746]_ ;
  assign \new_[46751]_  = \new_[46750]_  & \new_[46743]_ ;
  assign \new_[46755]_  = ~A267 & ~A235;
  assign \new_[46756]_  = ~A234 & \new_[46755]_ ;
  assign \new_[46759]_  = ~A269 & ~A268;
  assign \new_[46762]_  = A300 & A299;
  assign \new_[46763]_  = \new_[46762]_  & \new_[46759]_ ;
  assign \new_[46764]_  = \new_[46763]_  & \new_[46756]_ ;
  assign \new_[46768]_  = ~A168 & ~A169;
  assign \new_[46769]_  = ~A170 & \new_[46768]_ ;
  assign \new_[46772]_  = A201 & A200;
  assign \new_[46775]_  = A233 & A232;
  assign \new_[46776]_  = \new_[46775]_  & \new_[46772]_ ;
  assign \new_[46777]_  = \new_[46776]_  & \new_[46769]_ ;
  assign \new_[46781]_  = ~A267 & ~A235;
  assign \new_[46782]_  = ~A234 & \new_[46781]_ ;
  assign \new_[46785]_  = ~A269 & ~A268;
  assign \new_[46788]_  = A300 & A298;
  assign \new_[46789]_  = \new_[46788]_  & \new_[46785]_ ;
  assign \new_[46790]_  = \new_[46789]_  & \new_[46782]_ ;
  assign \new_[46794]_  = ~A168 & ~A169;
  assign \new_[46795]_  = ~A170 & \new_[46794]_ ;
  assign \new_[46798]_  = A201 & A200;
  assign \new_[46801]_  = A233 & A232;
  assign \new_[46802]_  = \new_[46801]_  & \new_[46798]_ ;
  assign \new_[46803]_  = \new_[46802]_  & \new_[46795]_ ;
  assign \new_[46807]_  = A265 & ~A235;
  assign \new_[46808]_  = ~A234 & \new_[46807]_ ;
  assign \new_[46811]_  = ~A267 & A266;
  assign \new_[46814]_  = A301 & ~A268;
  assign \new_[46815]_  = \new_[46814]_  & \new_[46811]_ ;
  assign \new_[46816]_  = \new_[46815]_  & \new_[46808]_ ;
  assign \new_[46820]_  = ~A168 & ~A169;
  assign \new_[46821]_  = ~A170 & \new_[46820]_ ;
  assign \new_[46824]_  = A201 & A200;
  assign \new_[46827]_  = A233 & A232;
  assign \new_[46828]_  = \new_[46827]_  & \new_[46824]_ ;
  assign \new_[46829]_  = \new_[46828]_  & \new_[46821]_ ;
  assign \new_[46833]_  = ~A265 & ~A235;
  assign \new_[46834]_  = ~A234 & \new_[46833]_ ;
  assign \new_[46837]_  = ~A268 & ~A266;
  assign \new_[46840]_  = A300 & A299;
  assign \new_[46841]_  = \new_[46840]_  & \new_[46837]_ ;
  assign \new_[46842]_  = \new_[46841]_  & \new_[46834]_ ;
  assign \new_[46846]_  = ~A168 & ~A169;
  assign \new_[46847]_  = ~A170 & \new_[46846]_ ;
  assign \new_[46850]_  = A201 & A200;
  assign \new_[46853]_  = A233 & A232;
  assign \new_[46854]_  = \new_[46853]_  & \new_[46850]_ ;
  assign \new_[46855]_  = \new_[46854]_  & \new_[46847]_ ;
  assign \new_[46859]_  = ~A265 & ~A235;
  assign \new_[46860]_  = ~A234 & \new_[46859]_ ;
  assign \new_[46863]_  = ~A268 & ~A266;
  assign \new_[46866]_  = A300 & A298;
  assign \new_[46867]_  = \new_[46866]_  & \new_[46863]_ ;
  assign \new_[46868]_  = \new_[46867]_  & \new_[46860]_ ;
  assign \new_[46872]_  = ~A168 & ~A169;
  assign \new_[46873]_  = ~A170 & \new_[46872]_ ;
  assign \new_[46876]_  = A201 & A200;
  assign \new_[46879]_  = ~A233 & ~A232;
  assign \new_[46880]_  = \new_[46879]_  & \new_[46876]_ ;
  assign \new_[46881]_  = \new_[46880]_  & \new_[46873]_ ;
  assign \new_[46885]_  = ~A268 & ~A267;
  assign \new_[46886]_  = ~A235 & \new_[46885]_ ;
  assign \new_[46889]_  = A298 & ~A269;
  assign \new_[46892]_  = A302 & ~A299;
  assign \new_[46893]_  = \new_[46892]_  & \new_[46889]_ ;
  assign \new_[46894]_  = \new_[46893]_  & \new_[46886]_ ;
  assign \new_[46898]_  = ~A168 & ~A169;
  assign \new_[46899]_  = ~A170 & \new_[46898]_ ;
  assign \new_[46902]_  = A201 & A200;
  assign \new_[46905]_  = ~A233 & ~A232;
  assign \new_[46906]_  = \new_[46905]_  & \new_[46902]_ ;
  assign \new_[46907]_  = \new_[46906]_  & \new_[46899]_ ;
  assign \new_[46911]_  = ~A268 & ~A267;
  assign \new_[46912]_  = ~A235 & \new_[46911]_ ;
  assign \new_[46915]_  = ~A298 & ~A269;
  assign \new_[46918]_  = A302 & A299;
  assign \new_[46919]_  = \new_[46918]_  & \new_[46915]_ ;
  assign \new_[46920]_  = \new_[46919]_  & \new_[46912]_ ;
  assign \new_[46924]_  = ~A168 & ~A169;
  assign \new_[46925]_  = ~A170 & \new_[46924]_ ;
  assign \new_[46928]_  = A201 & A200;
  assign \new_[46931]_  = ~A233 & ~A232;
  assign \new_[46932]_  = \new_[46931]_  & \new_[46928]_ ;
  assign \new_[46933]_  = \new_[46932]_  & \new_[46925]_ ;
  assign \new_[46937]_  = A266 & A265;
  assign \new_[46938]_  = ~A235 & \new_[46937]_ ;
  assign \new_[46941]_  = ~A268 & ~A267;
  assign \new_[46944]_  = A300 & A299;
  assign \new_[46945]_  = \new_[46944]_  & \new_[46941]_ ;
  assign \new_[46946]_  = \new_[46945]_  & \new_[46938]_ ;
  assign \new_[46950]_  = ~A168 & ~A169;
  assign \new_[46951]_  = ~A170 & \new_[46950]_ ;
  assign \new_[46954]_  = A201 & A200;
  assign \new_[46957]_  = ~A233 & ~A232;
  assign \new_[46958]_  = \new_[46957]_  & \new_[46954]_ ;
  assign \new_[46959]_  = \new_[46958]_  & \new_[46951]_ ;
  assign \new_[46963]_  = A266 & A265;
  assign \new_[46964]_  = ~A235 & \new_[46963]_ ;
  assign \new_[46967]_  = ~A268 & ~A267;
  assign \new_[46970]_  = A300 & A298;
  assign \new_[46971]_  = \new_[46970]_  & \new_[46967]_ ;
  assign \new_[46972]_  = \new_[46971]_  & \new_[46964]_ ;
  assign \new_[46976]_  = ~A168 & ~A169;
  assign \new_[46977]_  = ~A170 & \new_[46976]_ ;
  assign \new_[46980]_  = A201 & A200;
  assign \new_[46983]_  = ~A233 & ~A232;
  assign \new_[46984]_  = \new_[46983]_  & \new_[46980]_ ;
  assign \new_[46985]_  = \new_[46984]_  & \new_[46977]_ ;
  assign \new_[46989]_  = ~A266 & ~A265;
  assign \new_[46990]_  = ~A235 & \new_[46989]_ ;
  assign \new_[46993]_  = A298 & ~A268;
  assign \new_[46996]_  = A302 & ~A299;
  assign \new_[46997]_  = \new_[46996]_  & \new_[46993]_ ;
  assign \new_[46998]_  = \new_[46997]_  & \new_[46990]_ ;
  assign \new_[47002]_  = ~A168 & ~A169;
  assign \new_[47003]_  = ~A170 & \new_[47002]_ ;
  assign \new_[47006]_  = A201 & A200;
  assign \new_[47009]_  = ~A233 & ~A232;
  assign \new_[47010]_  = \new_[47009]_  & \new_[47006]_ ;
  assign \new_[47011]_  = \new_[47010]_  & \new_[47003]_ ;
  assign \new_[47015]_  = ~A266 & ~A265;
  assign \new_[47016]_  = ~A235 & \new_[47015]_ ;
  assign \new_[47019]_  = ~A298 & ~A268;
  assign \new_[47022]_  = A302 & A299;
  assign \new_[47023]_  = \new_[47022]_  & \new_[47019]_ ;
  assign \new_[47024]_  = \new_[47023]_  & \new_[47016]_ ;
  assign \new_[47028]_  = ~A168 & ~A169;
  assign \new_[47029]_  = ~A170 & \new_[47028]_ ;
  assign \new_[47032]_  = A200 & ~A199;
  assign \new_[47035]_  = ~A234 & A203;
  assign \new_[47036]_  = \new_[47035]_  & \new_[47032]_ ;
  assign \new_[47037]_  = \new_[47036]_  & \new_[47029]_ ;
  assign \new_[47041]_  = ~A267 & ~A236;
  assign \new_[47042]_  = ~A235 & \new_[47041]_ ;
  assign \new_[47045]_  = ~A269 & ~A268;
  assign \new_[47048]_  = A300 & A299;
  assign \new_[47049]_  = \new_[47048]_  & \new_[47045]_ ;
  assign \new_[47050]_  = \new_[47049]_  & \new_[47042]_ ;
  assign \new_[47054]_  = ~A168 & ~A169;
  assign \new_[47055]_  = ~A170 & \new_[47054]_ ;
  assign \new_[47058]_  = A200 & ~A199;
  assign \new_[47061]_  = ~A234 & A203;
  assign \new_[47062]_  = \new_[47061]_  & \new_[47058]_ ;
  assign \new_[47063]_  = \new_[47062]_  & \new_[47055]_ ;
  assign \new_[47067]_  = ~A267 & ~A236;
  assign \new_[47068]_  = ~A235 & \new_[47067]_ ;
  assign \new_[47071]_  = ~A269 & ~A268;
  assign \new_[47074]_  = A300 & A298;
  assign \new_[47075]_  = \new_[47074]_  & \new_[47071]_ ;
  assign \new_[47076]_  = \new_[47075]_  & \new_[47068]_ ;
  assign \new_[47080]_  = ~A168 & ~A169;
  assign \new_[47081]_  = ~A170 & \new_[47080]_ ;
  assign \new_[47084]_  = A200 & ~A199;
  assign \new_[47087]_  = ~A234 & A203;
  assign \new_[47088]_  = \new_[47087]_  & \new_[47084]_ ;
  assign \new_[47089]_  = \new_[47088]_  & \new_[47081]_ ;
  assign \new_[47093]_  = A265 & ~A236;
  assign \new_[47094]_  = ~A235 & \new_[47093]_ ;
  assign \new_[47097]_  = ~A267 & A266;
  assign \new_[47100]_  = A301 & ~A268;
  assign \new_[47101]_  = \new_[47100]_  & \new_[47097]_ ;
  assign \new_[47102]_  = \new_[47101]_  & \new_[47094]_ ;
  assign \new_[47106]_  = ~A168 & ~A169;
  assign \new_[47107]_  = ~A170 & \new_[47106]_ ;
  assign \new_[47110]_  = A200 & ~A199;
  assign \new_[47113]_  = ~A234 & A203;
  assign \new_[47114]_  = \new_[47113]_  & \new_[47110]_ ;
  assign \new_[47115]_  = \new_[47114]_  & \new_[47107]_ ;
  assign \new_[47119]_  = ~A265 & ~A236;
  assign \new_[47120]_  = ~A235 & \new_[47119]_ ;
  assign \new_[47123]_  = ~A268 & ~A266;
  assign \new_[47126]_  = A300 & A299;
  assign \new_[47127]_  = \new_[47126]_  & \new_[47123]_ ;
  assign \new_[47128]_  = \new_[47127]_  & \new_[47120]_ ;
  assign \new_[47132]_  = ~A168 & ~A169;
  assign \new_[47133]_  = ~A170 & \new_[47132]_ ;
  assign \new_[47136]_  = A200 & ~A199;
  assign \new_[47139]_  = ~A234 & A203;
  assign \new_[47140]_  = \new_[47139]_  & \new_[47136]_ ;
  assign \new_[47141]_  = \new_[47140]_  & \new_[47133]_ ;
  assign \new_[47145]_  = ~A265 & ~A236;
  assign \new_[47146]_  = ~A235 & \new_[47145]_ ;
  assign \new_[47149]_  = ~A268 & ~A266;
  assign \new_[47152]_  = A300 & A298;
  assign \new_[47153]_  = \new_[47152]_  & \new_[47149]_ ;
  assign \new_[47154]_  = \new_[47153]_  & \new_[47146]_ ;
  assign \new_[47158]_  = ~A168 & ~A169;
  assign \new_[47159]_  = ~A170 & \new_[47158]_ ;
  assign \new_[47162]_  = A200 & ~A199;
  assign \new_[47165]_  = A232 & A203;
  assign \new_[47166]_  = \new_[47165]_  & \new_[47162]_ ;
  assign \new_[47167]_  = \new_[47166]_  & \new_[47159]_ ;
  assign \new_[47171]_  = ~A235 & ~A234;
  assign \new_[47172]_  = A233 & \new_[47171]_ ;
  assign \new_[47175]_  = ~A268 & ~A267;
  assign \new_[47178]_  = A301 & ~A269;
  assign \new_[47179]_  = \new_[47178]_  & \new_[47175]_ ;
  assign \new_[47180]_  = \new_[47179]_  & \new_[47172]_ ;
  assign \new_[47184]_  = ~A168 & ~A169;
  assign \new_[47185]_  = ~A170 & \new_[47184]_ ;
  assign \new_[47188]_  = A200 & ~A199;
  assign \new_[47191]_  = A232 & A203;
  assign \new_[47192]_  = \new_[47191]_  & \new_[47188]_ ;
  assign \new_[47193]_  = \new_[47192]_  & \new_[47185]_ ;
  assign \new_[47197]_  = ~A235 & ~A234;
  assign \new_[47198]_  = A233 & \new_[47197]_ ;
  assign \new_[47201]_  = ~A266 & ~A265;
  assign \new_[47204]_  = A301 & ~A268;
  assign \new_[47205]_  = \new_[47204]_  & \new_[47201]_ ;
  assign \new_[47206]_  = \new_[47205]_  & \new_[47198]_ ;
  assign \new_[47210]_  = ~A168 & ~A169;
  assign \new_[47211]_  = ~A170 & \new_[47210]_ ;
  assign \new_[47214]_  = A200 & ~A199;
  assign \new_[47217]_  = ~A232 & A203;
  assign \new_[47218]_  = \new_[47217]_  & \new_[47214]_ ;
  assign \new_[47219]_  = \new_[47218]_  & \new_[47211]_ ;
  assign \new_[47223]_  = ~A267 & ~A235;
  assign \new_[47224]_  = ~A233 & \new_[47223]_ ;
  assign \new_[47227]_  = ~A269 & ~A268;
  assign \new_[47230]_  = A300 & A299;
  assign \new_[47231]_  = \new_[47230]_  & \new_[47227]_ ;
  assign \new_[47232]_  = \new_[47231]_  & \new_[47224]_ ;
  assign \new_[47236]_  = ~A168 & ~A169;
  assign \new_[47237]_  = ~A170 & \new_[47236]_ ;
  assign \new_[47240]_  = A200 & ~A199;
  assign \new_[47243]_  = ~A232 & A203;
  assign \new_[47244]_  = \new_[47243]_  & \new_[47240]_ ;
  assign \new_[47245]_  = \new_[47244]_  & \new_[47237]_ ;
  assign \new_[47249]_  = ~A267 & ~A235;
  assign \new_[47250]_  = ~A233 & \new_[47249]_ ;
  assign \new_[47253]_  = ~A269 & ~A268;
  assign \new_[47256]_  = A300 & A298;
  assign \new_[47257]_  = \new_[47256]_  & \new_[47253]_ ;
  assign \new_[47258]_  = \new_[47257]_  & \new_[47250]_ ;
  assign \new_[47262]_  = ~A168 & ~A169;
  assign \new_[47263]_  = ~A170 & \new_[47262]_ ;
  assign \new_[47266]_  = A200 & ~A199;
  assign \new_[47269]_  = ~A232 & A203;
  assign \new_[47270]_  = \new_[47269]_  & \new_[47266]_ ;
  assign \new_[47271]_  = \new_[47270]_  & \new_[47263]_ ;
  assign \new_[47275]_  = A265 & ~A235;
  assign \new_[47276]_  = ~A233 & \new_[47275]_ ;
  assign \new_[47279]_  = ~A267 & A266;
  assign \new_[47282]_  = A301 & ~A268;
  assign \new_[47283]_  = \new_[47282]_  & \new_[47279]_ ;
  assign \new_[47284]_  = \new_[47283]_  & \new_[47276]_ ;
  assign \new_[47288]_  = ~A168 & ~A169;
  assign \new_[47289]_  = ~A170 & \new_[47288]_ ;
  assign \new_[47292]_  = A200 & ~A199;
  assign \new_[47295]_  = ~A232 & A203;
  assign \new_[47296]_  = \new_[47295]_  & \new_[47292]_ ;
  assign \new_[47297]_  = \new_[47296]_  & \new_[47289]_ ;
  assign \new_[47301]_  = ~A265 & ~A235;
  assign \new_[47302]_  = ~A233 & \new_[47301]_ ;
  assign \new_[47305]_  = ~A268 & ~A266;
  assign \new_[47308]_  = A300 & A299;
  assign \new_[47309]_  = \new_[47308]_  & \new_[47305]_ ;
  assign \new_[47310]_  = \new_[47309]_  & \new_[47302]_ ;
  assign \new_[47314]_  = ~A168 & ~A169;
  assign \new_[47315]_  = ~A170 & \new_[47314]_ ;
  assign \new_[47318]_  = A200 & ~A199;
  assign \new_[47321]_  = ~A232 & A203;
  assign \new_[47322]_  = \new_[47321]_  & \new_[47318]_ ;
  assign \new_[47323]_  = \new_[47322]_  & \new_[47315]_ ;
  assign \new_[47327]_  = ~A265 & ~A235;
  assign \new_[47328]_  = ~A233 & \new_[47327]_ ;
  assign \new_[47331]_  = ~A268 & ~A266;
  assign \new_[47334]_  = A300 & A298;
  assign \new_[47335]_  = \new_[47334]_  & \new_[47331]_ ;
  assign \new_[47336]_  = \new_[47335]_  & \new_[47328]_ ;
  assign \new_[47340]_  = ~A168 & ~A169;
  assign \new_[47341]_  = ~A170 & \new_[47340]_ ;
  assign \new_[47344]_  = ~A200 & A199;
  assign \new_[47347]_  = ~A234 & A203;
  assign \new_[47348]_  = \new_[47347]_  & \new_[47344]_ ;
  assign \new_[47349]_  = \new_[47348]_  & \new_[47341]_ ;
  assign \new_[47353]_  = ~A267 & ~A236;
  assign \new_[47354]_  = ~A235 & \new_[47353]_ ;
  assign \new_[47357]_  = ~A269 & ~A268;
  assign \new_[47360]_  = A300 & A299;
  assign \new_[47361]_  = \new_[47360]_  & \new_[47357]_ ;
  assign \new_[47362]_  = \new_[47361]_  & \new_[47354]_ ;
  assign \new_[47366]_  = ~A168 & ~A169;
  assign \new_[47367]_  = ~A170 & \new_[47366]_ ;
  assign \new_[47370]_  = ~A200 & A199;
  assign \new_[47373]_  = ~A234 & A203;
  assign \new_[47374]_  = \new_[47373]_  & \new_[47370]_ ;
  assign \new_[47375]_  = \new_[47374]_  & \new_[47367]_ ;
  assign \new_[47379]_  = ~A267 & ~A236;
  assign \new_[47380]_  = ~A235 & \new_[47379]_ ;
  assign \new_[47383]_  = ~A269 & ~A268;
  assign \new_[47386]_  = A300 & A298;
  assign \new_[47387]_  = \new_[47386]_  & \new_[47383]_ ;
  assign \new_[47388]_  = \new_[47387]_  & \new_[47380]_ ;
  assign \new_[47392]_  = ~A168 & ~A169;
  assign \new_[47393]_  = ~A170 & \new_[47392]_ ;
  assign \new_[47396]_  = ~A200 & A199;
  assign \new_[47399]_  = ~A234 & A203;
  assign \new_[47400]_  = \new_[47399]_  & \new_[47396]_ ;
  assign \new_[47401]_  = \new_[47400]_  & \new_[47393]_ ;
  assign \new_[47405]_  = A265 & ~A236;
  assign \new_[47406]_  = ~A235 & \new_[47405]_ ;
  assign \new_[47409]_  = ~A267 & A266;
  assign \new_[47412]_  = A301 & ~A268;
  assign \new_[47413]_  = \new_[47412]_  & \new_[47409]_ ;
  assign \new_[47414]_  = \new_[47413]_  & \new_[47406]_ ;
  assign \new_[47418]_  = ~A168 & ~A169;
  assign \new_[47419]_  = ~A170 & \new_[47418]_ ;
  assign \new_[47422]_  = ~A200 & A199;
  assign \new_[47425]_  = ~A234 & A203;
  assign \new_[47426]_  = \new_[47425]_  & \new_[47422]_ ;
  assign \new_[47427]_  = \new_[47426]_  & \new_[47419]_ ;
  assign \new_[47431]_  = ~A265 & ~A236;
  assign \new_[47432]_  = ~A235 & \new_[47431]_ ;
  assign \new_[47435]_  = ~A268 & ~A266;
  assign \new_[47438]_  = A300 & A299;
  assign \new_[47439]_  = \new_[47438]_  & \new_[47435]_ ;
  assign \new_[47440]_  = \new_[47439]_  & \new_[47432]_ ;
  assign \new_[47444]_  = ~A168 & ~A169;
  assign \new_[47445]_  = ~A170 & \new_[47444]_ ;
  assign \new_[47448]_  = ~A200 & A199;
  assign \new_[47451]_  = ~A234 & A203;
  assign \new_[47452]_  = \new_[47451]_  & \new_[47448]_ ;
  assign \new_[47453]_  = \new_[47452]_  & \new_[47445]_ ;
  assign \new_[47457]_  = ~A265 & ~A236;
  assign \new_[47458]_  = ~A235 & \new_[47457]_ ;
  assign \new_[47461]_  = ~A268 & ~A266;
  assign \new_[47464]_  = A300 & A298;
  assign \new_[47465]_  = \new_[47464]_  & \new_[47461]_ ;
  assign \new_[47466]_  = \new_[47465]_  & \new_[47458]_ ;
  assign \new_[47470]_  = ~A168 & ~A169;
  assign \new_[47471]_  = ~A170 & \new_[47470]_ ;
  assign \new_[47474]_  = ~A200 & A199;
  assign \new_[47477]_  = A232 & A203;
  assign \new_[47478]_  = \new_[47477]_  & \new_[47474]_ ;
  assign \new_[47479]_  = \new_[47478]_  & \new_[47471]_ ;
  assign \new_[47483]_  = ~A235 & ~A234;
  assign \new_[47484]_  = A233 & \new_[47483]_ ;
  assign \new_[47487]_  = ~A268 & ~A267;
  assign \new_[47490]_  = A301 & ~A269;
  assign \new_[47491]_  = \new_[47490]_  & \new_[47487]_ ;
  assign \new_[47492]_  = \new_[47491]_  & \new_[47484]_ ;
  assign \new_[47496]_  = ~A168 & ~A169;
  assign \new_[47497]_  = ~A170 & \new_[47496]_ ;
  assign \new_[47500]_  = ~A200 & A199;
  assign \new_[47503]_  = A232 & A203;
  assign \new_[47504]_  = \new_[47503]_  & \new_[47500]_ ;
  assign \new_[47505]_  = \new_[47504]_  & \new_[47497]_ ;
  assign \new_[47509]_  = ~A235 & ~A234;
  assign \new_[47510]_  = A233 & \new_[47509]_ ;
  assign \new_[47513]_  = ~A266 & ~A265;
  assign \new_[47516]_  = A301 & ~A268;
  assign \new_[47517]_  = \new_[47516]_  & \new_[47513]_ ;
  assign \new_[47518]_  = \new_[47517]_  & \new_[47510]_ ;
  assign \new_[47522]_  = ~A168 & ~A169;
  assign \new_[47523]_  = ~A170 & \new_[47522]_ ;
  assign \new_[47526]_  = ~A200 & A199;
  assign \new_[47529]_  = ~A232 & A203;
  assign \new_[47530]_  = \new_[47529]_  & \new_[47526]_ ;
  assign \new_[47531]_  = \new_[47530]_  & \new_[47523]_ ;
  assign \new_[47535]_  = ~A267 & ~A235;
  assign \new_[47536]_  = ~A233 & \new_[47535]_ ;
  assign \new_[47539]_  = ~A269 & ~A268;
  assign \new_[47542]_  = A300 & A299;
  assign \new_[47543]_  = \new_[47542]_  & \new_[47539]_ ;
  assign \new_[47544]_  = \new_[47543]_  & \new_[47536]_ ;
  assign \new_[47548]_  = ~A168 & ~A169;
  assign \new_[47549]_  = ~A170 & \new_[47548]_ ;
  assign \new_[47552]_  = ~A200 & A199;
  assign \new_[47555]_  = ~A232 & A203;
  assign \new_[47556]_  = \new_[47555]_  & \new_[47552]_ ;
  assign \new_[47557]_  = \new_[47556]_  & \new_[47549]_ ;
  assign \new_[47561]_  = ~A267 & ~A235;
  assign \new_[47562]_  = ~A233 & \new_[47561]_ ;
  assign \new_[47565]_  = ~A269 & ~A268;
  assign \new_[47568]_  = A300 & A298;
  assign \new_[47569]_  = \new_[47568]_  & \new_[47565]_ ;
  assign \new_[47570]_  = \new_[47569]_  & \new_[47562]_ ;
  assign \new_[47574]_  = ~A168 & ~A169;
  assign \new_[47575]_  = ~A170 & \new_[47574]_ ;
  assign \new_[47578]_  = ~A200 & A199;
  assign \new_[47581]_  = ~A232 & A203;
  assign \new_[47582]_  = \new_[47581]_  & \new_[47578]_ ;
  assign \new_[47583]_  = \new_[47582]_  & \new_[47575]_ ;
  assign \new_[47587]_  = A265 & ~A235;
  assign \new_[47588]_  = ~A233 & \new_[47587]_ ;
  assign \new_[47591]_  = ~A267 & A266;
  assign \new_[47594]_  = A301 & ~A268;
  assign \new_[47595]_  = \new_[47594]_  & \new_[47591]_ ;
  assign \new_[47596]_  = \new_[47595]_  & \new_[47588]_ ;
  assign \new_[47600]_  = ~A168 & ~A169;
  assign \new_[47601]_  = ~A170 & \new_[47600]_ ;
  assign \new_[47604]_  = ~A200 & A199;
  assign \new_[47607]_  = ~A232 & A203;
  assign \new_[47608]_  = \new_[47607]_  & \new_[47604]_ ;
  assign \new_[47609]_  = \new_[47608]_  & \new_[47601]_ ;
  assign \new_[47613]_  = ~A265 & ~A235;
  assign \new_[47614]_  = ~A233 & \new_[47613]_ ;
  assign \new_[47617]_  = ~A268 & ~A266;
  assign \new_[47620]_  = A300 & A299;
  assign \new_[47621]_  = \new_[47620]_  & \new_[47617]_ ;
  assign \new_[47622]_  = \new_[47621]_  & \new_[47614]_ ;
  assign \new_[47626]_  = ~A168 & ~A169;
  assign \new_[47627]_  = ~A170 & \new_[47626]_ ;
  assign \new_[47630]_  = ~A200 & A199;
  assign \new_[47633]_  = ~A232 & A203;
  assign \new_[47634]_  = \new_[47633]_  & \new_[47630]_ ;
  assign \new_[47635]_  = \new_[47634]_  & \new_[47627]_ ;
  assign \new_[47639]_  = ~A265 & ~A235;
  assign \new_[47640]_  = ~A233 & \new_[47639]_ ;
  assign \new_[47643]_  = ~A268 & ~A266;
  assign \new_[47646]_  = A300 & A298;
  assign \new_[47647]_  = \new_[47646]_  & \new_[47643]_ ;
  assign \new_[47648]_  = \new_[47647]_  & \new_[47640]_ ;
  assign \new_[47652]_  = ~A201 & A166;
  assign \new_[47653]_  = A168 & \new_[47652]_ ;
  assign \new_[47656]_  = ~A203 & ~A202;
  assign \new_[47659]_  = ~A235 & ~A234;
  assign \new_[47660]_  = \new_[47659]_  & \new_[47656]_ ;
  assign \new_[47661]_  = \new_[47660]_  & \new_[47653]_ ;
  assign \new_[47664]_  = A265 & ~A236;
  assign \new_[47667]_  = ~A267 & A266;
  assign \new_[47668]_  = \new_[47667]_  & \new_[47664]_ ;
  assign \new_[47671]_  = A298 & ~A268;
  assign \new_[47674]_  = A302 & ~A299;
  assign \new_[47675]_  = \new_[47674]_  & \new_[47671]_ ;
  assign \new_[47676]_  = \new_[47675]_  & \new_[47668]_ ;
  assign \new_[47680]_  = ~A201 & A166;
  assign \new_[47681]_  = A168 & \new_[47680]_ ;
  assign \new_[47684]_  = ~A203 & ~A202;
  assign \new_[47687]_  = ~A235 & ~A234;
  assign \new_[47688]_  = \new_[47687]_  & \new_[47684]_ ;
  assign \new_[47689]_  = \new_[47688]_  & \new_[47681]_ ;
  assign \new_[47692]_  = A265 & ~A236;
  assign \new_[47695]_  = ~A267 & A266;
  assign \new_[47696]_  = \new_[47695]_  & \new_[47692]_ ;
  assign \new_[47699]_  = ~A298 & ~A268;
  assign \new_[47702]_  = A302 & A299;
  assign \new_[47703]_  = \new_[47702]_  & \new_[47699]_ ;
  assign \new_[47704]_  = \new_[47703]_  & \new_[47696]_ ;
  assign \new_[47708]_  = ~A201 & A166;
  assign \new_[47709]_  = A168 & \new_[47708]_ ;
  assign \new_[47712]_  = ~A203 & ~A202;
  assign \new_[47715]_  = A233 & A232;
  assign \new_[47716]_  = \new_[47715]_  & \new_[47712]_ ;
  assign \new_[47717]_  = \new_[47716]_  & \new_[47709]_ ;
  assign \new_[47720]_  = ~A235 & ~A234;
  assign \new_[47723]_  = ~A268 & ~A267;
  assign \new_[47724]_  = \new_[47723]_  & \new_[47720]_ ;
  assign \new_[47727]_  = A298 & ~A269;
  assign \new_[47730]_  = A302 & ~A299;
  assign \new_[47731]_  = \new_[47730]_  & \new_[47727]_ ;
  assign \new_[47732]_  = \new_[47731]_  & \new_[47724]_ ;
  assign \new_[47736]_  = ~A201 & A166;
  assign \new_[47737]_  = A168 & \new_[47736]_ ;
  assign \new_[47740]_  = ~A203 & ~A202;
  assign \new_[47743]_  = A233 & A232;
  assign \new_[47744]_  = \new_[47743]_  & \new_[47740]_ ;
  assign \new_[47745]_  = \new_[47744]_  & \new_[47737]_ ;
  assign \new_[47748]_  = ~A235 & ~A234;
  assign \new_[47751]_  = ~A268 & ~A267;
  assign \new_[47752]_  = \new_[47751]_  & \new_[47748]_ ;
  assign \new_[47755]_  = ~A298 & ~A269;
  assign \new_[47758]_  = A302 & A299;
  assign \new_[47759]_  = \new_[47758]_  & \new_[47755]_ ;
  assign \new_[47760]_  = \new_[47759]_  & \new_[47752]_ ;
  assign \new_[47764]_  = ~A201 & A166;
  assign \new_[47765]_  = A168 & \new_[47764]_ ;
  assign \new_[47768]_  = ~A203 & ~A202;
  assign \new_[47771]_  = A233 & A232;
  assign \new_[47772]_  = \new_[47771]_  & \new_[47768]_ ;
  assign \new_[47773]_  = \new_[47772]_  & \new_[47765]_ ;
  assign \new_[47776]_  = ~A235 & ~A234;
  assign \new_[47779]_  = A266 & A265;
  assign \new_[47780]_  = \new_[47779]_  & \new_[47776]_ ;
  assign \new_[47783]_  = ~A268 & ~A267;
  assign \new_[47786]_  = A300 & A299;
  assign \new_[47787]_  = \new_[47786]_  & \new_[47783]_ ;
  assign \new_[47788]_  = \new_[47787]_  & \new_[47780]_ ;
  assign \new_[47792]_  = ~A201 & A166;
  assign \new_[47793]_  = A168 & \new_[47792]_ ;
  assign \new_[47796]_  = ~A203 & ~A202;
  assign \new_[47799]_  = A233 & A232;
  assign \new_[47800]_  = \new_[47799]_  & \new_[47796]_ ;
  assign \new_[47801]_  = \new_[47800]_  & \new_[47793]_ ;
  assign \new_[47804]_  = ~A235 & ~A234;
  assign \new_[47807]_  = A266 & A265;
  assign \new_[47808]_  = \new_[47807]_  & \new_[47804]_ ;
  assign \new_[47811]_  = ~A268 & ~A267;
  assign \new_[47814]_  = A300 & A298;
  assign \new_[47815]_  = \new_[47814]_  & \new_[47811]_ ;
  assign \new_[47816]_  = \new_[47815]_  & \new_[47808]_ ;
  assign \new_[47820]_  = ~A201 & A166;
  assign \new_[47821]_  = A168 & \new_[47820]_ ;
  assign \new_[47824]_  = ~A203 & ~A202;
  assign \new_[47827]_  = A233 & A232;
  assign \new_[47828]_  = \new_[47827]_  & \new_[47824]_ ;
  assign \new_[47829]_  = \new_[47828]_  & \new_[47821]_ ;
  assign \new_[47832]_  = ~A235 & ~A234;
  assign \new_[47835]_  = ~A266 & ~A265;
  assign \new_[47836]_  = \new_[47835]_  & \new_[47832]_ ;
  assign \new_[47839]_  = A298 & ~A268;
  assign \new_[47842]_  = A302 & ~A299;
  assign \new_[47843]_  = \new_[47842]_  & \new_[47839]_ ;
  assign \new_[47844]_  = \new_[47843]_  & \new_[47836]_ ;
  assign \new_[47848]_  = ~A201 & A166;
  assign \new_[47849]_  = A168 & \new_[47848]_ ;
  assign \new_[47852]_  = ~A203 & ~A202;
  assign \new_[47855]_  = A233 & A232;
  assign \new_[47856]_  = \new_[47855]_  & \new_[47852]_ ;
  assign \new_[47857]_  = \new_[47856]_  & \new_[47849]_ ;
  assign \new_[47860]_  = ~A235 & ~A234;
  assign \new_[47863]_  = ~A266 & ~A265;
  assign \new_[47864]_  = \new_[47863]_  & \new_[47860]_ ;
  assign \new_[47867]_  = ~A298 & ~A268;
  assign \new_[47870]_  = A302 & A299;
  assign \new_[47871]_  = \new_[47870]_  & \new_[47867]_ ;
  assign \new_[47872]_  = \new_[47871]_  & \new_[47864]_ ;
  assign \new_[47876]_  = ~A201 & A166;
  assign \new_[47877]_  = A168 & \new_[47876]_ ;
  assign \new_[47880]_  = ~A203 & ~A202;
  assign \new_[47883]_  = ~A233 & ~A232;
  assign \new_[47884]_  = \new_[47883]_  & \new_[47880]_ ;
  assign \new_[47885]_  = \new_[47884]_  & \new_[47877]_ ;
  assign \new_[47888]_  = A265 & ~A235;
  assign \new_[47891]_  = ~A267 & A266;
  assign \new_[47892]_  = \new_[47891]_  & \new_[47888]_ ;
  assign \new_[47895]_  = A298 & ~A268;
  assign \new_[47898]_  = A302 & ~A299;
  assign \new_[47899]_  = \new_[47898]_  & \new_[47895]_ ;
  assign \new_[47900]_  = \new_[47899]_  & \new_[47892]_ ;
  assign \new_[47904]_  = ~A201 & A166;
  assign \new_[47905]_  = A168 & \new_[47904]_ ;
  assign \new_[47908]_  = ~A203 & ~A202;
  assign \new_[47911]_  = ~A233 & ~A232;
  assign \new_[47912]_  = \new_[47911]_  & \new_[47908]_ ;
  assign \new_[47913]_  = \new_[47912]_  & \new_[47905]_ ;
  assign \new_[47916]_  = A265 & ~A235;
  assign \new_[47919]_  = ~A267 & A266;
  assign \new_[47920]_  = \new_[47919]_  & \new_[47916]_ ;
  assign \new_[47923]_  = ~A298 & ~A268;
  assign \new_[47926]_  = A302 & A299;
  assign \new_[47927]_  = \new_[47926]_  & \new_[47923]_ ;
  assign \new_[47928]_  = \new_[47927]_  & \new_[47920]_ ;
  assign \new_[47932]_  = A199 & A166;
  assign \new_[47933]_  = A168 & \new_[47932]_ ;
  assign \new_[47936]_  = ~A201 & A200;
  assign \new_[47939]_  = ~A234 & ~A202;
  assign \new_[47940]_  = \new_[47939]_  & \new_[47936]_ ;
  assign \new_[47941]_  = \new_[47940]_  & \new_[47933]_ ;
  assign \new_[47944]_  = ~A236 & ~A235;
  assign \new_[47947]_  = ~A268 & ~A267;
  assign \new_[47948]_  = \new_[47947]_  & \new_[47944]_ ;
  assign \new_[47951]_  = A298 & ~A269;
  assign \new_[47954]_  = A302 & ~A299;
  assign \new_[47955]_  = \new_[47954]_  & \new_[47951]_ ;
  assign \new_[47956]_  = \new_[47955]_  & \new_[47948]_ ;
  assign \new_[47960]_  = A199 & A166;
  assign \new_[47961]_  = A168 & \new_[47960]_ ;
  assign \new_[47964]_  = ~A201 & A200;
  assign \new_[47967]_  = ~A234 & ~A202;
  assign \new_[47968]_  = \new_[47967]_  & \new_[47964]_ ;
  assign \new_[47969]_  = \new_[47968]_  & \new_[47961]_ ;
  assign \new_[47972]_  = ~A236 & ~A235;
  assign \new_[47975]_  = ~A268 & ~A267;
  assign \new_[47976]_  = \new_[47975]_  & \new_[47972]_ ;
  assign \new_[47979]_  = ~A298 & ~A269;
  assign \new_[47982]_  = A302 & A299;
  assign \new_[47983]_  = \new_[47982]_  & \new_[47979]_ ;
  assign \new_[47984]_  = \new_[47983]_  & \new_[47976]_ ;
  assign \new_[47988]_  = A199 & A166;
  assign \new_[47989]_  = A168 & \new_[47988]_ ;
  assign \new_[47992]_  = ~A201 & A200;
  assign \new_[47995]_  = ~A234 & ~A202;
  assign \new_[47996]_  = \new_[47995]_  & \new_[47992]_ ;
  assign \new_[47997]_  = \new_[47996]_  & \new_[47989]_ ;
  assign \new_[48000]_  = ~A236 & ~A235;
  assign \new_[48003]_  = A266 & A265;
  assign \new_[48004]_  = \new_[48003]_  & \new_[48000]_ ;
  assign \new_[48007]_  = ~A268 & ~A267;
  assign \new_[48010]_  = A300 & A299;
  assign \new_[48011]_  = \new_[48010]_  & \new_[48007]_ ;
  assign \new_[48012]_  = \new_[48011]_  & \new_[48004]_ ;
  assign \new_[48016]_  = A199 & A166;
  assign \new_[48017]_  = A168 & \new_[48016]_ ;
  assign \new_[48020]_  = ~A201 & A200;
  assign \new_[48023]_  = ~A234 & ~A202;
  assign \new_[48024]_  = \new_[48023]_  & \new_[48020]_ ;
  assign \new_[48025]_  = \new_[48024]_  & \new_[48017]_ ;
  assign \new_[48028]_  = ~A236 & ~A235;
  assign \new_[48031]_  = A266 & A265;
  assign \new_[48032]_  = \new_[48031]_  & \new_[48028]_ ;
  assign \new_[48035]_  = ~A268 & ~A267;
  assign \new_[48038]_  = A300 & A298;
  assign \new_[48039]_  = \new_[48038]_  & \new_[48035]_ ;
  assign \new_[48040]_  = \new_[48039]_  & \new_[48032]_ ;
  assign \new_[48044]_  = A199 & A166;
  assign \new_[48045]_  = A168 & \new_[48044]_ ;
  assign \new_[48048]_  = ~A201 & A200;
  assign \new_[48051]_  = ~A234 & ~A202;
  assign \new_[48052]_  = \new_[48051]_  & \new_[48048]_ ;
  assign \new_[48053]_  = \new_[48052]_  & \new_[48045]_ ;
  assign \new_[48056]_  = ~A236 & ~A235;
  assign \new_[48059]_  = ~A266 & ~A265;
  assign \new_[48060]_  = \new_[48059]_  & \new_[48056]_ ;
  assign \new_[48063]_  = A298 & ~A268;
  assign \new_[48066]_  = A302 & ~A299;
  assign \new_[48067]_  = \new_[48066]_  & \new_[48063]_ ;
  assign \new_[48068]_  = \new_[48067]_  & \new_[48060]_ ;
  assign \new_[48072]_  = A199 & A166;
  assign \new_[48073]_  = A168 & \new_[48072]_ ;
  assign \new_[48076]_  = ~A201 & A200;
  assign \new_[48079]_  = ~A234 & ~A202;
  assign \new_[48080]_  = \new_[48079]_  & \new_[48076]_ ;
  assign \new_[48081]_  = \new_[48080]_  & \new_[48073]_ ;
  assign \new_[48084]_  = ~A236 & ~A235;
  assign \new_[48087]_  = ~A266 & ~A265;
  assign \new_[48088]_  = \new_[48087]_  & \new_[48084]_ ;
  assign \new_[48091]_  = ~A298 & ~A268;
  assign \new_[48094]_  = A302 & A299;
  assign \new_[48095]_  = \new_[48094]_  & \new_[48091]_ ;
  assign \new_[48096]_  = \new_[48095]_  & \new_[48088]_ ;
  assign \new_[48100]_  = A199 & A166;
  assign \new_[48101]_  = A168 & \new_[48100]_ ;
  assign \new_[48104]_  = ~A201 & A200;
  assign \new_[48107]_  = A232 & ~A202;
  assign \new_[48108]_  = \new_[48107]_  & \new_[48104]_ ;
  assign \new_[48109]_  = \new_[48108]_  & \new_[48101]_ ;
  assign \new_[48112]_  = ~A234 & A233;
  assign \new_[48115]_  = ~A267 & ~A235;
  assign \new_[48116]_  = \new_[48115]_  & \new_[48112]_ ;
  assign \new_[48119]_  = ~A269 & ~A268;
  assign \new_[48122]_  = A300 & A299;
  assign \new_[48123]_  = \new_[48122]_  & \new_[48119]_ ;
  assign \new_[48124]_  = \new_[48123]_  & \new_[48116]_ ;
  assign \new_[48128]_  = A199 & A166;
  assign \new_[48129]_  = A168 & \new_[48128]_ ;
  assign \new_[48132]_  = ~A201 & A200;
  assign \new_[48135]_  = A232 & ~A202;
  assign \new_[48136]_  = \new_[48135]_  & \new_[48132]_ ;
  assign \new_[48137]_  = \new_[48136]_  & \new_[48129]_ ;
  assign \new_[48140]_  = ~A234 & A233;
  assign \new_[48143]_  = ~A267 & ~A235;
  assign \new_[48144]_  = \new_[48143]_  & \new_[48140]_ ;
  assign \new_[48147]_  = ~A269 & ~A268;
  assign \new_[48150]_  = A300 & A298;
  assign \new_[48151]_  = \new_[48150]_  & \new_[48147]_ ;
  assign \new_[48152]_  = \new_[48151]_  & \new_[48144]_ ;
  assign \new_[48156]_  = A199 & A166;
  assign \new_[48157]_  = A168 & \new_[48156]_ ;
  assign \new_[48160]_  = ~A201 & A200;
  assign \new_[48163]_  = A232 & ~A202;
  assign \new_[48164]_  = \new_[48163]_  & \new_[48160]_ ;
  assign \new_[48165]_  = \new_[48164]_  & \new_[48157]_ ;
  assign \new_[48168]_  = ~A234 & A233;
  assign \new_[48171]_  = A265 & ~A235;
  assign \new_[48172]_  = \new_[48171]_  & \new_[48168]_ ;
  assign \new_[48175]_  = ~A267 & A266;
  assign \new_[48178]_  = A301 & ~A268;
  assign \new_[48179]_  = \new_[48178]_  & \new_[48175]_ ;
  assign \new_[48180]_  = \new_[48179]_  & \new_[48172]_ ;
  assign \new_[48184]_  = A199 & A166;
  assign \new_[48185]_  = A168 & \new_[48184]_ ;
  assign \new_[48188]_  = ~A201 & A200;
  assign \new_[48191]_  = A232 & ~A202;
  assign \new_[48192]_  = \new_[48191]_  & \new_[48188]_ ;
  assign \new_[48193]_  = \new_[48192]_  & \new_[48185]_ ;
  assign \new_[48196]_  = ~A234 & A233;
  assign \new_[48199]_  = ~A265 & ~A235;
  assign \new_[48200]_  = \new_[48199]_  & \new_[48196]_ ;
  assign \new_[48203]_  = ~A268 & ~A266;
  assign \new_[48206]_  = A300 & A299;
  assign \new_[48207]_  = \new_[48206]_  & \new_[48203]_ ;
  assign \new_[48208]_  = \new_[48207]_  & \new_[48200]_ ;
  assign \new_[48212]_  = A199 & A166;
  assign \new_[48213]_  = A168 & \new_[48212]_ ;
  assign \new_[48216]_  = ~A201 & A200;
  assign \new_[48219]_  = A232 & ~A202;
  assign \new_[48220]_  = \new_[48219]_  & \new_[48216]_ ;
  assign \new_[48221]_  = \new_[48220]_  & \new_[48213]_ ;
  assign \new_[48224]_  = ~A234 & A233;
  assign \new_[48227]_  = ~A265 & ~A235;
  assign \new_[48228]_  = \new_[48227]_  & \new_[48224]_ ;
  assign \new_[48231]_  = ~A268 & ~A266;
  assign \new_[48234]_  = A300 & A298;
  assign \new_[48235]_  = \new_[48234]_  & \new_[48231]_ ;
  assign \new_[48236]_  = \new_[48235]_  & \new_[48228]_ ;
  assign \new_[48240]_  = A199 & A166;
  assign \new_[48241]_  = A168 & \new_[48240]_ ;
  assign \new_[48244]_  = ~A201 & A200;
  assign \new_[48247]_  = ~A232 & ~A202;
  assign \new_[48248]_  = \new_[48247]_  & \new_[48244]_ ;
  assign \new_[48249]_  = \new_[48248]_  & \new_[48241]_ ;
  assign \new_[48252]_  = ~A235 & ~A233;
  assign \new_[48255]_  = ~A268 & ~A267;
  assign \new_[48256]_  = \new_[48255]_  & \new_[48252]_ ;
  assign \new_[48259]_  = A298 & ~A269;
  assign \new_[48262]_  = A302 & ~A299;
  assign \new_[48263]_  = \new_[48262]_  & \new_[48259]_ ;
  assign \new_[48264]_  = \new_[48263]_  & \new_[48256]_ ;
  assign \new_[48268]_  = A199 & A166;
  assign \new_[48269]_  = A168 & \new_[48268]_ ;
  assign \new_[48272]_  = ~A201 & A200;
  assign \new_[48275]_  = ~A232 & ~A202;
  assign \new_[48276]_  = \new_[48275]_  & \new_[48272]_ ;
  assign \new_[48277]_  = \new_[48276]_  & \new_[48269]_ ;
  assign \new_[48280]_  = ~A235 & ~A233;
  assign \new_[48283]_  = ~A268 & ~A267;
  assign \new_[48284]_  = \new_[48283]_  & \new_[48280]_ ;
  assign \new_[48287]_  = ~A298 & ~A269;
  assign \new_[48290]_  = A302 & A299;
  assign \new_[48291]_  = \new_[48290]_  & \new_[48287]_ ;
  assign \new_[48292]_  = \new_[48291]_  & \new_[48284]_ ;
  assign \new_[48296]_  = A199 & A166;
  assign \new_[48297]_  = A168 & \new_[48296]_ ;
  assign \new_[48300]_  = ~A201 & A200;
  assign \new_[48303]_  = ~A232 & ~A202;
  assign \new_[48304]_  = \new_[48303]_  & \new_[48300]_ ;
  assign \new_[48305]_  = \new_[48304]_  & \new_[48297]_ ;
  assign \new_[48308]_  = ~A235 & ~A233;
  assign \new_[48311]_  = A266 & A265;
  assign \new_[48312]_  = \new_[48311]_  & \new_[48308]_ ;
  assign \new_[48315]_  = ~A268 & ~A267;
  assign \new_[48318]_  = A300 & A299;
  assign \new_[48319]_  = \new_[48318]_  & \new_[48315]_ ;
  assign \new_[48320]_  = \new_[48319]_  & \new_[48312]_ ;
  assign \new_[48324]_  = A199 & A166;
  assign \new_[48325]_  = A168 & \new_[48324]_ ;
  assign \new_[48328]_  = ~A201 & A200;
  assign \new_[48331]_  = ~A232 & ~A202;
  assign \new_[48332]_  = \new_[48331]_  & \new_[48328]_ ;
  assign \new_[48333]_  = \new_[48332]_  & \new_[48325]_ ;
  assign \new_[48336]_  = ~A235 & ~A233;
  assign \new_[48339]_  = A266 & A265;
  assign \new_[48340]_  = \new_[48339]_  & \new_[48336]_ ;
  assign \new_[48343]_  = ~A268 & ~A267;
  assign \new_[48346]_  = A300 & A298;
  assign \new_[48347]_  = \new_[48346]_  & \new_[48343]_ ;
  assign \new_[48348]_  = \new_[48347]_  & \new_[48340]_ ;
  assign \new_[48352]_  = A199 & A166;
  assign \new_[48353]_  = A168 & \new_[48352]_ ;
  assign \new_[48356]_  = ~A201 & A200;
  assign \new_[48359]_  = ~A232 & ~A202;
  assign \new_[48360]_  = \new_[48359]_  & \new_[48356]_ ;
  assign \new_[48361]_  = \new_[48360]_  & \new_[48353]_ ;
  assign \new_[48364]_  = ~A235 & ~A233;
  assign \new_[48367]_  = ~A266 & ~A265;
  assign \new_[48368]_  = \new_[48367]_  & \new_[48364]_ ;
  assign \new_[48371]_  = A298 & ~A268;
  assign \new_[48374]_  = A302 & ~A299;
  assign \new_[48375]_  = \new_[48374]_  & \new_[48371]_ ;
  assign \new_[48376]_  = \new_[48375]_  & \new_[48368]_ ;
  assign \new_[48380]_  = A199 & A166;
  assign \new_[48381]_  = A168 & \new_[48380]_ ;
  assign \new_[48384]_  = ~A201 & A200;
  assign \new_[48387]_  = ~A232 & ~A202;
  assign \new_[48388]_  = \new_[48387]_  & \new_[48384]_ ;
  assign \new_[48389]_  = \new_[48388]_  & \new_[48381]_ ;
  assign \new_[48392]_  = ~A235 & ~A233;
  assign \new_[48395]_  = ~A266 & ~A265;
  assign \new_[48396]_  = \new_[48395]_  & \new_[48392]_ ;
  assign \new_[48399]_  = ~A298 & ~A268;
  assign \new_[48402]_  = A302 & A299;
  assign \new_[48403]_  = \new_[48402]_  & \new_[48399]_ ;
  assign \new_[48404]_  = \new_[48403]_  & \new_[48396]_ ;
  assign \new_[48408]_  = ~A199 & A166;
  assign \new_[48409]_  = A168 & \new_[48408]_ ;
  assign \new_[48412]_  = ~A202 & ~A200;
  assign \new_[48415]_  = ~A235 & ~A234;
  assign \new_[48416]_  = \new_[48415]_  & \new_[48412]_ ;
  assign \new_[48417]_  = \new_[48416]_  & \new_[48409]_ ;
  assign \new_[48420]_  = A265 & ~A236;
  assign \new_[48423]_  = ~A267 & A266;
  assign \new_[48424]_  = \new_[48423]_  & \new_[48420]_ ;
  assign \new_[48427]_  = A298 & ~A268;
  assign \new_[48430]_  = A302 & ~A299;
  assign \new_[48431]_  = \new_[48430]_  & \new_[48427]_ ;
  assign \new_[48432]_  = \new_[48431]_  & \new_[48424]_ ;
  assign \new_[48436]_  = ~A199 & A166;
  assign \new_[48437]_  = A168 & \new_[48436]_ ;
  assign \new_[48440]_  = ~A202 & ~A200;
  assign \new_[48443]_  = ~A235 & ~A234;
  assign \new_[48444]_  = \new_[48443]_  & \new_[48440]_ ;
  assign \new_[48445]_  = \new_[48444]_  & \new_[48437]_ ;
  assign \new_[48448]_  = A265 & ~A236;
  assign \new_[48451]_  = ~A267 & A266;
  assign \new_[48452]_  = \new_[48451]_  & \new_[48448]_ ;
  assign \new_[48455]_  = ~A298 & ~A268;
  assign \new_[48458]_  = A302 & A299;
  assign \new_[48459]_  = \new_[48458]_  & \new_[48455]_ ;
  assign \new_[48460]_  = \new_[48459]_  & \new_[48452]_ ;
  assign \new_[48464]_  = ~A199 & A166;
  assign \new_[48465]_  = A168 & \new_[48464]_ ;
  assign \new_[48468]_  = ~A202 & ~A200;
  assign \new_[48471]_  = A233 & A232;
  assign \new_[48472]_  = \new_[48471]_  & \new_[48468]_ ;
  assign \new_[48473]_  = \new_[48472]_  & \new_[48465]_ ;
  assign \new_[48476]_  = ~A235 & ~A234;
  assign \new_[48479]_  = ~A268 & ~A267;
  assign \new_[48480]_  = \new_[48479]_  & \new_[48476]_ ;
  assign \new_[48483]_  = A298 & ~A269;
  assign \new_[48486]_  = A302 & ~A299;
  assign \new_[48487]_  = \new_[48486]_  & \new_[48483]_ ;
  assign \new_[48488]_  = \new_[48487]_  & \new_[48480]_ ;
  assign \new_[48492]_  = ~A199 & A166;
  assign \new_[48493]_  = A168 & \new_[48492]_ ;
  assign \new_[48496]_  = ~A202 & ~A200;
  assign \new_[48499]_  = A233 & A232;
  assign \new_[48500]_  = \new_[48499]_  & \new_[48496]_ ;
  assign \new_[48501]_  = \new_[48500]_  & \new_[48493]_ ;
  assign \new_[48504]_  = ~A235 & ~A234;
  assign \new_[48507]_  = ~A268 & ~A267;
  assign \new_[48508]_  = \new_[48507]_  & \new_[48504]_ ;
  assign \new_[48511]_  = ~A298 & ~A269;
  assign \new_[48514]_  = A302 & A299;
  assign \new_[48515]_  = \new_[48514]_  & \new_[48511]_ ;
  assign \new_[48516]_  = \new_[48515]_  & \new_[48508]_ ;
  assign \new_[48520]_  = ~A199 & A166;
  assign \new_[48521]_  = A168 & \new_[48520]_ ;
  assign \new_[48524]_  = ~A202 & ~A200;
  assign \new_[48527]_  = A233 & A232;
  assign \new_[48528]_  = \new_[48527]_  & \new_[48524]_ ;
  assign \new_[48529]_  = \new_[48528]_  & \new_[48521]_ ;
  assign \new_[48532]_  = ~A235 & ~A234;
  assign \new_[48535]_  = A266 & A265;
  assign \new_[48536]_  = \new_[48535]_  & \new_[48532]_ ;
  assign \new_[48539]_  = ~A268 & ~A267;
  assign \new_[48542]_  = A300 & A299;
  assign \new_[48543]_  = \new_[48542]_  & \new_[48539]_ ;
  assign \new_[48544]_  = \new_[48543]_  & \new_[48536]_ ;
  assign \new_[48548]_  = ~A199 & A166;
  assign \new_[48549]_  = A168 & \new_[48548]_ ;
  assign \new_[48552]_  = ~A202 & ~A200;
  assign \new_[48555]_  = A233 & A232;
  assign \new_[48556]_  = \new_[48555]_  & \new_[48552]_ ;
  assign \new_[48557]_  = \new_[48556]_  & \new_[48549]_ ;
  assign \new_[48560]_  = ~A235 & ~A234;
  assign \new_[48563]_  = A266 & A265;
  assign \new_[48564]_  = \new_[48563]_  & \new_[48560]_ ;
  assign \new_[48567]_  = ~A268 & ~A267;
  assign \new_[48570]_  = A300 & A298;
  assign \new_[48571]_  = \new_[48570]_  & \new_[48567]_ ;
  assign \new_[48572]_  = \new_[48571]_  & \new_[48564]_ ;
  assign \new_[48576]_  = ~A199 & A166;
  assign \new_[48577]_  = A168 & \new_[48576]_ ;
  assign \new_[48580]_  = ~A202 & ~A200;
  assign \new_[48583]_  = A233 & A232;
  assign \new_[48584]_  = \new_[48583]_  & \new_[48580]_ ;
  assign \new_[48585]_  = \new_[48584]_  & \new_[48577]_ ;
  assign \new_[48588]_  = ~A235 & ~A234;
  assign \new_[48591]_  = ~A266 & ~A265;
  assign \new_[48592]_  = \new_[48591]_  & \new_[48588]_ ;
  assign \new_[48595]_  = A298 & ~A268;
  assign \new_[48598]_  = A302 & ~A299;
  assign \new_[48599]_  = \new_[48598]_  & \new_[48595]_ ;
  assign \new_[48600]_  = \new_[48599]_  & \new_[48592]_ ;
  assign \new_[48604]_  = ~A199 & A166;
  assign \new_[48605]_  = A168 & \new_[48604]_ ;
  assign \new_[48608]_  = ~A202 & ~A200;
  assign \new_[48611]_  = A233 & A232;
  assign \new_[48612]_  = \new_[48611]_  & \new_[48608]_ ;
  assign \new_[48613]_  = \new_[48612]_  & \new_[48605]_ ;
  assign \new_[48616]_  = ~A235 & ~A234;
  assign \new_[48619]_  = ~A266 & ~A265;
  assign \new_[48620]_  = \new_[48619]_  & \new_[48616]_ ;
  assign \new_[48623]_  = ~A298 & ~A268;
  assign \new_[48626]_  = A302 & A299;
  assign \new_[48627]_  = \new_[48626]_  & \new_[48623]_ ;
  assign \new_[48628]_  = \new_[48627]_  & \new_[48620]_ ;
  assign \new_[48632]_  = ~A199 & A166;
  assign \new_[48633]_  = A168 & \new_[48632]_ ;
  assign \new_[48636]_  = ~A202 & ~A200;
  assign \new_[48639]_  = ~A233 & ~A232;
  assign \new_[48640]_  = \new_[48639]_  & \new_[48636]_ ;
  assign \new_[48641]_  = \new_[48640]_  & \new_[48633]_ ;
  assign \new_[48644]_  = A265 & ~A235;
  assign \new_[48647]_  = ~A267 & A266;
  assign \new_[48648]_  = \new_[48647]_  & \new_[48644]_ ;
  assign \new_[48651]_  = A298 & ~A268;
  assign \new_[48654]_  = A302 & ~A299;
  assign \new_[48655]_  = \new_[48654]_  & \new_[48651]_ ;
  assign \new_[48656]_  = \new_[48655]_  & \new_[48648]_ ;
  assign \new_[48660]_  = ~A199 & A166;
  assign \new_[48661]_  = A168 & \new_[48660]_ ;
  assign \new_[48664]_  = ~A202 & ~A200;
  assign \new_[48667]_  = ~A233 & ~A232;
  assign \new_[48668]_  = \new_[48667]_  & \new_[48664]_ ;
  assign \new_[48669]_  = \new_[48668]_  & \new_[48661]_ ;
  assign \new_[48672]_  = A265 & ~A235;
  assign \new_[48675]_  = ~A267 & A266;
  assign \new_[48676]_  = \new_[48675]_  & \new_[48672]_ ;
  assign \new_[48679]_  = ~A298 & ~A268;
  assign \new_[48682]_  = A302 & A299;
  assign \new_[48683]_  = \new_[48682]_  & \new_[48679]_ ;
  assign \new_[48684]_  = \new_[48683]_  & \new_[48676]_ ;
  assign \new_[48688]_  = ~A201 & A167;
  assign \new_[48689]_  = A168 & \new_[48688]_ ;
  assign \new_[48692]_  = ~A203 & ~A202;
  assign \new_[48695]_  = ~A235 & ~A234;
  assign \new_[48696]_  = \new_[48695]_  & \new_[48692]_ ;
  assign \new_[48697]_  = \new_[48696]_  & \new_[48689]_ ;
  assign \new_[48700]_  = A265 & ~A236;
  assign \new_[48703]_  = ~A267 & A266;
  assign \new_[48704]_  = \new_[48703]_  & \new_[48700]_ ;
  assign \new_[48707]_  = A298 & ~A268;
  assign \new_[48710]_  = A302 & ~A299;
  assign \new_[48711]_  = \new_[48710]_  & \new_[48707]_ ;
  assign \new_[48712]_  = \new_[48711]_  & \new_[48704]_ ;
  assign \new_[48716]_  = ~A201 & A167;
  assign \new_[48717]_  = A168 & \new_[48716]_ ;
  assign \new_[48720]_  = ~A203 & ~A202;
  assign \new_[48723]_  = ~A235 & ~A234;
  assign \new_[48724]_  = \new_[48723]_  & \new_[48720]_ ;
  assign \new_[48725]_  = \new_[48724]_  & \new_[48717]_ ;
  assign \new_[48728]_  = A265 & ~A236;
  assign \new_[48731]_  = ~A267 & A266;
  assign \new_[48732]_  = \new_[48731]_  & \new_[48728]_ ;
  assign \new_[48735]_  = ~A298 & ~A268;
  assign \new_[48738]_  = A302 & A299;
  assign \new_[48739]_  = \new_[48738]_  & \new_[48735]_ ;
  assign \new_[48740]_  = \new_[48739]_  & \new_[48732]_ ;
  assign \new_[48744]_  = ~A201 & A167;
  assign \new_[48745]_  = A168 & \new_[48744]_ ;
  assign \new_[48748]_  = ~A203 & ~A202;
  assign \new_[48751]_  = A233 & A232;
  assign \new_[48752]_  = \new_[48751]_  & \new_[48748]_ ;
  assign \new_[48753]_  = \new_[48752]_  & \new_[48745]_ ;
  assign \new_[48756]_  = ~A235 & ~A234;
  assign \new_[48759]_  = ~A268 & ~A267;
  assign \new_[48760]_  = \new_[48759]_  & \new_[48756]_ ;
  assign \new_[48763]_  = A298 & ~A269;
  assign \new_[48766]_  = A302 & ~A299;
  assign \new_[48767]_  = \new_[48766]_  & \new_[48763]_ ;
  assign \new_[48768]_  = \new_[48767]_  & \new_[48760]_ ;
  assign \new_[48772]_  = ~A201 & A167;
  assign \new_[48773]_  = A168 & \new_[48772]_ ;
  assign \new_[48776]_  = ~A203 & ~A202;
  assign \new_[48779]_  = A233 & A232;
  assign \new_[48780]_  = \new_[48779]_  & \new_[48776]_ ;
  assign \new_[48781]_  = \new_[48780]_  & \new_[48773]_ ;
  assign \new_[48784]_  = ~A235 & ~A234;
  assign \new_[48787]_  = ~A268 & ~A267;
  assign \new_[48788]_  = \new_[48787]_  & \new_[48784]_ ;
  assign \new_[48791]_  = ~A298 & ~A269;
  assign \new_[48794]_  = A302 & A299;
  assign \new_[48795]_  = \new_[48794]_  & \new_[48791]_ ;
  assign \new_[48796]_  = \new_[48795]_  & \new_[48788]_ ;
  assign \new_[48800]_  = ~A201 & A167;
  assign \new_[48801]_  = A168 & \new_[48800]_ ;
  assign \new_[48804]_  = ~A203 & ~A202;
  assign \new_[48807]_  = A233 & A232;
  assign \new_[48808]_  = \new_[48807]_  & \new_[48804]_ ;
  assign \new_[48809]_  = \new_[48808]_  & \new_[48801]_ ;
  assign \new_[48812]_  = ~A235 & ~A234;
  assign \new_[48815]_  = A266 & A265;
  assign \new_[48816]_  = \new_[48815]_  & \new_[48812]_ ;
  assign \new_[48819]_  = ~A268 & ~A267;
  assign \new_[48822]_  = A300 & A299;
  assign \new_[48823]_  = \new_[48822]_  & \new_[48819]_ ;
  assign \new_[48824]_  = \new_[48823]_  & \new_[48816]_ ;
  assign \new_[48828]_  = ~A201 & A167;
  assign \new_[48829]_  = A168 & \new_[48828]_ ;
  assign \new_[48832]_  = ~A203 & ~A202;
  assign \new_[48835]_  = A233 & A232;
  assign \new_[48836]_  = \new_[48835]_  & \new_[48832]_ ;
  assign \new_[48837]_  = \new_[48836]_  & \new_[48829]_ ;
  assign \new_[48840]_  = ~A235 & ~A234;
  assign \new_[48843]_  = A266 & A265;
  assign \new_[48844]_  = \new_[48843]_  & \new_[48840]_ ;
  assign \new_[48847]_  = ~A268 & ~A267;
  assign \new_[48850]_  = A300 & A298;
  assign \new_[48851]_  = \new_[48850]_  & \new_[48847]_ ;
  assign \new_[48852]_  = \new_[48851]_  & \new_[48844]_ ;
  assign \new_[48856]_  = ~A201 & A167;
  assign \new_[48857]_  = A168 & \new_[48856]_ ;
  assign \new_[48860]_  = ~A203 & ~A202;
  assign \new_[48863]_  = A233 & A232;
  assign \new_[48864]_  = \new_[48863]_  & \new_[48860]_ ;
  assign \new_[48865]_  = \new_[48864]_  & \new_[48857]_ ;
  assign \new_[48868]_  = ~A235 & ~A234;
  assign \new_[48871]_  = ~A266 & ~A265;
  assign \new_[48872]_  = \new_[48871]_  & \new_[48868]_ ;
  assign \new_[48875]_  = A298 & ~A268;
  assign \new_[48878]_  = A302 & ~A299;
  assign \new_[48879]_  = \new_[48878]_  & \new_[48875]_ ;
  assign \new_[48880]_  = \new_[48879]_  & \new_[48872]_ ;
  assign \new_[48884]_  = ~A201 & A167;
  assign \new_[48885]_  = A168 & \new_[48884]_ ;
  assign \new_[48888]_  = ~A203 & ~A202;
  assign \new_[48891]_  = A233 & A232;
  assign \new_[48892]_  = \new_[48891]_  & \new_[48888]_ ;
  assign \new_[48893]_  = \new_[48892]_  & \new_[48885]_ ;
  assign \new_[48896]_  = ~A235 & ~A234;
  assign \new_[48899]_  = ~A266 & ~A265;
  assign \new_[48900]_  = \new_[48899]_  & \new_[48896]_ ;
  assign \new_[48903]_  = ~A298 & ~A268;
  assign \new_[48906]_  = A302 & A299;
  assign \new_[48907]_  = \new_[48906]_  & \new_[48903]_ ;
  assign \new_[48908]_  = \new_[48907]_  & \new_[48900]_ ;
  assign \new_[48912]_  = ~A201 & A167;
  assign \new_[48913]_  = A168 & \new_[48912]_ ;
  assign \new_[48916]_  = ~A203 & ~A202;
  assign \new_[48919]_  = ~A233 & ~A232;
  assign \new_[48920]_  = \new_[48919]_  & \new_[48916]_ ;
  assign \new_[48921]_  = \new_[48920]_  & \new_[48913]_ ;
  assign \new_[48924]_  = A265 & ~A235;
  assign \new_[48927]_  = ~A267 & A266;
  assign \new_[48928]_  = \new_[48927]_  & \new_[48924]_ ;
  assign \new_[48931]_  = A298 & ~A268;
  assign \new_[48934]_  = A302 & ~A299;
  assign \new_[48935]_  = \new_[48934]_  & \new_[48931]_ ;
  assign \new_[48936]_  = \new_[48935]_  & \new_[48928]_ ;
  assign \new_[48940]_  = ~A201 & A167;
  assign \new_[48941]_  = A168 & \new_[48940]_ ;
  assign \new_[48944]_  = ~A203 & ~A202;
  assign \new_[48947]_  = ~A233 & ~A232;
  assign \new_[48948]_  = \new_[48947]_  & \new_[48944]_ ;
  assign \new_[48949]_  = \new_[48948]_  & \new_[48941]_ ;
  assign \new_[48952]_  = A265 & ~A235;
  assign \new_[48955]_  = ~A267 & A266;
  assign \new_[48956]_  = \new_[48955]_  & \new_[48952]_ ;
  assign \new_[48959]_  = ~A298 & ~A268;
  assign \new_[48962]_  = A302 & A299;
  assign \new_[48963]_  = \new_[48962]_  & \new_[48959]_ ;
  assign \new_[48964]_  = \new_[48963]_  & \new_[48956]_ ;
  assign \new_[48968]_  = A199 & A167;
  assign \new_[48969]_  = A168 & \new_[48968]_ ;
  assign \new_[48972]_  = ~A201 & A200;
  assign \new_[48975]_  = ~A234 & ~A202;
  assign \new_[48976]_  = \new_[48975]_  & \new_[48972]_ ;
  assign \new_[48977]_  = \new_[48976]_  & \new_[48969]_ ;
  assign \new_[48980]_  = ~A236 & ~A235;
  assign \new_[48983]_  = ~A268 & ~A267;
  assign \new_[48984]_  = \new_[48983]_  & \new_[48980]_ ;
  assign \new_[48987]_  = A298 & ~A269;
  assign \new_[48990]_  = A302 & ~A299;
  assign \new_[48991]_  = \new_[48990]_  & \new_[48987]_ ;
  assign \new_[48992]_  = \new_[48991]_  & \new_[48984]_ ;
  assign \new_[48996]_  = A199 & A167;
  assign \new_[48997]_  = A168 & \new_[48996]_ ;
  assign \new_[49000]_  = ~A201 & A200;
  assign \new_[49003]_  = ~A234 & ~A202;
  assign \new_[49004]_  = \new_[49003]_  & \new_[49000]_ ;
  assign \new_[49005]_  = \new_[49004]_  & \new_[48997]_ ;
  assign \new_[49008]_  = ~A236 & ~A235;
  assign \new_[49011]_  = ~A268 & ~A267;
  assign \new_[49012]_  = \new_[49011]_  & \new_[49008]_ ;
  assign \new_[49015]_  = ~A298 & ~A269;
  assign \new_[49018]_  = A302 & A299;
  assign \new_[49019]_  = \new_[49018]_  & \new_[49015]_ ;
  assign \new_[49020]_  = \new_[49019]_  & \new_[49012]_ ;
  assign \new_[49024]_  = A199 & A167;
  assign \new_[49025]_  = A168 & \new_[49024]_ ;
  assign \new_[49028]_  = ~A201 & A200;
  assign \new_[49031]_  = ~A234 & ~A202;
  assign \new_[49032]_  = \new_[49031]_  & \new_[49028]_ ;
  assign \new_[49033]_  = \new_[49032]_  & \new_[49025]_ ;
  assign \new_[49036]_  = ~A236 & ~A235;
  assign \new_[49039]_  = A266 & A265;
  assign \new_[49040]_  = \new_[49039]_  & \new_[49036]_ ;
  assign \new_[49043]_  = ~A268 & ~A267;
  assign \new_[49046]_  = A300 & A299;
  assign \new_[49047]_  = \new_[49046]_  & \new_[49043]_ ;
  assign \new_[49048]_  = \new_[49047]_  & \new_[49040]_ ;
  assign \new_[49052]_  = A199 & A167;
  assign \new_[49053]_  = A168 & \new_[49052]_ ;
  assign \new_[49056]_  = ~A201 & A200;
  assign \new_[49059]_  = ~A234 & ~A202;
  assign \new_[49060]_  = \new_[49059]_  & \new_[49056]_ ;
  assign \new_[49061]_  = \new_[49060]_  & \new_[49053]_ ;
  assign \new_[49064]_  = ~A236 & ~A235;
  assign \new_[49067]_  = A266 & A265;
  assign \new_[49068]_  = \new_[49067]_  & \new_[49064]_ ;
  assign \new_[49071]_  = ~A268 & ~A267;
  assign \new_[49074]_  = A300 & A298;
  assign \new_[49075]_  = \new_[49074]_  & \new_[49071]_ ;
  assign \new_[49076]_  = \new_[49075]_  & \new_[49068]_ ;
  assign \new_[49080]_  = A199 & A167;
  assign \new_[49081]_  = A168 & \new_[49080]_ ;
  assign \new_[49084]_  = ~A201 & A200;
  assign \new_[49087]_  = ~A234 & ~A202;
  assign \new_[49088]_  = \new_[49087]_  & \new_[49084]_ ;
  assign \new_[49089]_  = \new_[49088]_  & \new_[49081]_ ;
  assign \new_[49092]_  = ~A236 & ~A235;
  assign \new_[49095]_  = ~A266 & ~A265;
  assign \new_[49096]_  = \new_[49095]_  & \new_[49092]_ ;
  assign \new_[49099]_  = A298 & ~A268;
  assign \new_[49102]_  = A302 & ~A299;
  assign \new_[49103]_  = \new_[49102]_  & \new_[49099]_ ;
  assign \new_[49104]_  = \new_[49103]_  & \new_[49096]_ ;
  assign \new_[49108]_  = A199 & A167;
  assign \new_[49109]_  = A168 & \new_[49108]_ ;
  assign \new_[49112]_  = ~A201 & A200;
  assign \new_[49115]_  = ~A234 & ~A202;
  assign \new_[49116]_  = \new_[49115]_  & \new_[49112]_ ;
  assign \new_[49117]_  = \new_[49116]_  & \new_[49109]_ ;
  assign \new_[49120]_  = ~A236 & ~A235;
  assign \new_[49123]_  = ~A266 & ~A265;
  assign \new_[49124]_  = \new_[49123]_  & \new_[49120]_ ;
  assign \new_[49127]_  = ~A298 & ~A268;
  assign \new_[49130]_  = A302 & A299;
  assign \new_[49131]_  = \new_[49130]_  & \new_[49127]_ ;
  assign \new_[49132]_  = \new_[49131]_  & \new_[49124]_ ;
  assign \new_[49136]_  = A199 & A167;
  assign \new_[49137]_  = A168 & \new_[49136]_ ;
  assign \new_[49140]_  = ~A201 & A200;
  assign \new_[49143]_  = A232 & ~A202;
  assign \new_[49144]_  = \new_[49143]_  & \new_[49140]_ ;
  assign \new_[49145]_  = \new_[49144]_  & \new_[49137]_ ;
  assign \new_[49148]_  = ~A234 & A233;
  assign \new_[49151]_  = ~A267 & ~A235;
  assign \new_[49152]_  = \new_[49151]_  & \new_[49148]_ ;
  assign \new_[49155]_  = ~A269 & ~A268;
  assign \new_[49158]_  = A300 & A299;
  assign \new_[49159]_  = \new_[49158]_  & \new_[49155]_ ;
  assign \new_[49160]_  = \new_[49159]_  & \new_[49152]_ ;
  assign \new_[49164]_  = A199 & A167;
  assign \new_[49165]_  = A168 & \new_[49164]_ ;
  assign \new_[49168]_  = ~A201 & A200;
  assign \new_[49171]_  = A232 & ~A202;
  assign \new_[49172]_  = \new_[49171]_  & \new_[49168]_ ;
  assign \new_[49173]_  = \new_[49172]_  & \new_[49165]_ ;
  assign \new_[49176]_  = ~A234 & A233;
  assign \new_[49179]_  = ~A267 & ~A235;
  assign \new_[49180]_  = \new_[49179]_  & \new_[49176]_ ;
  assign \new_[49183]_  = ~A269 & ~A268;
  assign \new_[49186]_  = A300 & A298;
  assign \new_[49187]_  = \new_[49186]_  & \new_[49183]_ ;
  assign \new_[49188]_  = \new_[49187]_  & \new_[49180]_ ;
  assign \new_[49192]_  = A199 & A167;
  assign \new_[49193]_  = A168 & \new_[49192]_ ;
  assign \new_[49196]_  = ~A201 & A200;
  assign \new_[49199]_  = A232 & ~A202;
  assign \new_[49200]_  = \new_[49199]_  & \new_[49196]_ ;
  assign \new_[49201]_  = \new_[49200]_  & \new_[49193]_ ;
  assign \new_[49204]_  = ~A234 & A233;
  assign \new_[49207]_  = A265 & ~A235;
  assign \new_[49208]_  = \new_[49207]_  & \new_[49204]_ ;
  assign \new_[49211]_  = ~A267 & A266;
  assign \new_[49214]_  = A301 & ~A268;
  assign \new_[49215]_  = \new_[49214]_  & \new_[49211]_ ;
  assign \new_[49216]_  = \new_[49215]_  & \new_[49208]_ ;
  assign \new_[49220]_  = A199 & A167;
  assign \new_[49221]_  = A168 & \new_[49220]_ ;
  assign \new_[49224]_  = ~A201 & A200;
  assign \new_[49227]_  = A232 & ~A202;
  assign \new_[49228]_  = \new_[49227]_  & \new_[49224]_ ;
  assign \new_[49229]_  = \new_[49228]_  & \new_[49221]_ ;
  assign \new_[49232]_  = ~A234 & A233;
  assign \new_[49235]_  = ~A265 & ~A235;
  assign \new_[49236]_  = \new_[49235]_  & \new_[49232]_ ;
  assign \new_[49239]_  = ~A268 & ~A266;
  assign \new_[49242]_  = A300 & A299;
  assign \new_[49243]_  = \new_[49242]_  & \new_[49239]_ ;
  assign \new_[49244]_  = \new_[49243]_  & \new_[49236]_ ;
  assign \new_[49248]_  = A199 & A167;
  assign \new_[49249]_  = A168 & \new_[49248]_ ;
  assign \new_[49252]_  = ~A201 & A200;
  assign \new_[49255]_  = A232 & ~A202;
  assign \new_[49256]_  = \new_[49255]_  & \new_[49252]_ ;
  assign \new_[49257]_  = \new_[49256]_  & \new_[49249]_ ;
  assign \new_[49260]_  = ~A234 & A233;
  assign \new_[49263]_  = ~A265 & ~A235;
  assign \new_[49264]_  = \new_[49263]_  & \new_[49260]_ ;
  assign \new_[49267]_  = ~A268 & ~A266;
  assign \new_[49270]_  = A300 & A298;
  assign \new_[49271]_  = \new_[49270]_  & \new_[49267]_ ;
  assign \new_[49272]_  = \new_[49271]_  & \new_[49264]_ ;
  assign \new_[49276]_  = A199 & A167;
  assign \new_[49277]_  = A168 & \new_[49276]_ ;
  assign \new_[49280]_  = ~A201 & A200;
  assign \new_[49283]_  = ~A232 & ~A202;
  assign \new_[49284]_  = \new_[49283]_  & \new_[49280]_ ;
  assign \new_[49285]_  = \new_[49284]_  & \new_[49277]_ ;
  assign \new_[49288]_  = ~A235 & ~A233;
  assign \new_[49291]_  = ~A268 & ~A267;
  assign \new_[49292]_  = \new_[49291]_  & \new_[49288]_ ;
  assign \new_[49295]_  = A298 & ~A269;
  assign \new_[49298]_  = A302 & ~A299;
  assign \new_[49299]_  = \new_[49298]_  & \new_[49295]_ ;
  assign \new_[49300]_  = \new_[49299]_  & \new_[49292]_ ;
  assign \new_[49304]_  = A199 & A167;
  assign \new_[49305]_  = A168 & \new_[49304]_ ;
  assign \new_[49308]_  = ~A201 & A200;
  assign \new_[49311]_  = ~A232 & ~A202;
  assign \new_[49312]_  = \new_[49311]_  & \new_[49308]_ ;
  assign \new_[49313]_  = \new_[49312]_  & \new_[49305]_ ;
  assign \new_[49316]_  = ~A235 & ~A233;
  assign \new_[49319]_  = ~A268 & ~A267;
  assign \new_[49320]_  = \new_[49319]_  & \new_[49316]_ ;
  assign \new_[49323]_  = ~A298 & ~A269;
  assign \new_[49326]_  = A302 & A299;
  assign \new_[49327]_  = \new_[49326]_  & \new_[49323]_ ;
  assign \new_[49328]_  = \new_[49327]_  & \new_[49320]_ ;
  assign \new_[49332]_  = A199 & A167;
  assign \new_[49333]_  = A168 & \new_[49332]_ ;
  assign \new_[49336]_  = ~A201 & A200;
  assign \new_[49339]_  = ~A232 & ~A202;
  assign \new_[49340]_  = \new_[49339]_  & \new_[49336]_ ;
  assign \new_[49341]_  = \new_[49340]_  & \new_[49333]_ ;
  assign \new_[49344]_  = ~A235 & ~A233;
  assign \new_[49347]_  = A266 & A265;
  assign \new_[49348]_  = \new_[49347]_  & \new_[49344]_ ;
  assign \new_[49351]_  = ~A268 & ~A267;
  assign \new_[49354]_  = A300 & A299;
  assign \new_[49355]_  = \new_[49354]_  & \new_[49351]_ ;
  assign \new_[49356]_  = \new_[49355]_  & \new_[49348]_ ;
  assign \new_[49360]_  = A199 & A167;
  assign \new_[49361]_  = A168 & \new_[49360]_ ;
  assign \new_[49364]_  = ~A201 & A200;
  assign \new_[49367]_  = ~A232 & ~A202;
  assign \new_[49368]_  = \new_[49367]_  & \new_[49364]_ ;
  assign \new_[49369]_  = \new_[49368]_  & \new_[49361]_ ;
  assign \new_[49372]_  = ~A235 & ~A233;
  assign \new_[49375]_  = A266 & A265;
  assign \new_[49376]_  = \new_[49375]_  & \new_[49372]_ ;
  assign \new_[49379]_  = ~A268 & ~A267;
  assign \new_[49382]_  = A300 & A298;
  assign \new_[49383]_  = \new_[49382]_  & \new_[49379]_ ;
  assign \new_[49384]_  = \new_[49383]_  & \new_[49376]_ ;
  assign \new_[49388]_  = A199 & A167;
  assign \new_[49389]_  = A168 & \new_[49388]_ ;
  assign \new_[49392]_  = ~A201 & A200;
  assign \new_[49395]_  = ~A232 & ~A202;
  assign \new_[49396]_  = \new_[49395]_  & \new_[49392]_ ;
  assign \new_[49397]_  = \new_[49396]_  & \new_[49389]_ ;
  assign \new_[49400]_  = ~A235 & ~A233;
  assign \new_[49403]_  = ~A266 & ~A265;
  assign \new_[49404]_  = \new_[49403]_  & \new_[49400]_ ;
  assign \new_[49407]_  = A298 & ~A268;
  assign \new_[49410]_  = A302 & ~A299;
  assign \new_[49411]_  = \new_[49410]_  & \new_[49407]_ ;
  assign \new_[49412]_  = \new_[49411]_  & \new_[49404]_ ;
  assign \new_[49416]_  = A199 & A167;
  assign \new_[49417]_  = A168 & \new_[49416]_ ;
  assign \new_[49420]_  = ~A201 & A200;
  assign \new_[49423]_  = ~A232 & ~A202;
  assign \new_[49424]_  = \new_[49423]_  & \new_[49420]_ ;
  assign \new_[49425]_  = \new_[49424]_  & \new_[49417]_ ;
  assign \new_[49428]_  = ~A235 & ~A233;
  assign \new_[49431]_  = ~A266 & ~A265;
  assign \new_[49432]_  = \new_[49431]_  & \new_[49428]_ ;
  assign \new_[49435]_  = ~A298 & ~A268;
  assign \new_[49438]_  = A302 & A299;
  assign \new_[49439]_  = \new_[49438]_  & \new_[49435]_ ;
  assign \new_[49440]_  = \new_[49439]_  & \new_[49432]_ ;
  assign \new_[49444]_  = ~A199 & A167;
  assign \new_[49445]_  = A168 & \new_[49444]_ ;
  assign \new_[49448]_  = ~A202 & ~A200;
  assign \new_[49451]_  = ~A235 & ~A234;
  assign \new_[49452]_  = \new_[49451]_  & \new_[49448]_ ;
  assign \new_[49453]_  = \new_[49452]_  & \new_[49445]_ ;
  assign \new_[49456]_  = A265 & ~A236;
  assign \new_[49459]_  = ~A267 & A266;
  assign \new_[49460]_  = \new_[49459]_  & \new_[49456]_ ;
  assign \new_[49463]_  = A298 & ~A268;
  assign \new_[49466]_  = A302 & ~A299;
  assign \new_[49467]_  = \new_[49466]_  & \new_[49463]_ ;
  assign \new_[49468]_  = \new_[49467]_  & \new_[49460]_ ;
  assign \new_[49472]_  = ~A199 & A167;
  assign \new_[49473]_  = A168 & \new_[49472]_ ;
  assign \new_[49476]_  = ~A202 & ~A200;
  assign \new_[49479]_  = ~A235 & ~A234;
  assign \new_[49480]_  = \new_[49479]_  & \new_[49476]_ ;
  assign \new_[49481]_  = \new_[49480]_  & \new_[49473]_ ;
  assign \new_[49484]_  = A265 & ~A236;
  assign \new_[49487]_  = ~A267 & A266;
  assign \new_[49488]_  = \new_[49487]_  & \new_[49484]_ ;
  assign \new_[49491]_  = ~A298 & ~A268;
  assign \new_[49494]_  = A302 & A299;
  assign \new_[49495]_  = \new_[49494]_  & \new_[49491]_ ;
  assign \new_[49496]_  = \new_[49495]_  & \new_[49488]_ ;
  assign \new_[49500]_  = ~A199 & A167;
  assign \new_[49501]_  = A168 & \new_[49500]_ ;
  assign \new_[49504]_  = ~A202 & ~A200;
  assign \new_[49507]_  = A233 & A232;
  assign \new_[49508]_  = \new_[49507]_  & \new_[49504]_ ;
  assign \new_[49509]_  = \new_[49508]_  & \new_[49501]_ ;
  assign \new_[49512]_  = ~A235 & ~A234;
  assign \new_[49515]_  = ~A268 & ~A267;
  assign \new_[49516]_  = \new_[49515]_  & \new_[49512]_ ;
  assign \new_[49519]_  = A298 & ~A269;
  assign \new_[49522]_  = A302 & ~A299;
  assign \new_[49523]_  = \new_[49522]_  & \new_[49519]_ ;
  assign \new_[49524]_  = \new_[49523]_  & \new_[49516]_ ;
  assign \new_[49528]_  = ~A199 & A167;
  assign \new_[49529]_  = A168 & \new_[49528]_ ;
  assign \new_[49532]_  = ~A202 & ~A200;
  assign \new_[49535]_  = A233 & A232;
  assign \new_[49536]_  = \new_[49535]_  & \new_[49532]_ ;
  assign \new_[49537]_  = \new_[49536]_  & \new_[49529]_ ;
  assign \new_[49540]_  = ~A235 & ~A234;
  assign \new_[49543]_  = ~A268 & ~A267;
  assign \new_[49544]_  = \new_[49543]_  & \new_[49540]_ ;
  assign \new_[49547]_  = ~A298 & ~A269;
  assign \new_[49550]_  = A302 & A299;
  assign \new_[49551]_  = \new_[49550]_  & \new_[49547]_ ;
  assign \new_[49552]_  = \new_[49551]_  & \new_[49544]_ ;
  assign \new_[49556]_  = ~A199 & A167;
  assign \new_[49557]_  = A168 & \new_[49556]_ ;
  assign \new_[49560]_  = ~A202 & ~A200;
  assign \new_[49563]_  = A233 & A232;
  assign \new_[49564]_  = \new_[49563]_  & \new_[49560]_ ;
  assign \new_[49565]_  = \new_[49564]_  & \new_[49557]_ ;
  assign \new_[49568]_  = ~A235 & ~A234;
  assign \new_[49571]_  = A266 & A265;
  assign \new_[49572]_  = \new_[49571]_  & \new_[49568]_ ;
  assign \new_[49575]_  = ~A268 & ~A267;
  assign \new_[49578]_  = A300 & A299;
  assign \new_[49579]_  = \new_[49578]_  & \new_[49575]_ ;
  assign \new_[49580]_  = \new_[49579]_  & \new_[49572]_ ;
  assign \new_[49584]_  = ~A199 & A167;
  assign \new_[49585]_  = A168 & \new_[49584]_ ;
  assign \new_[49588]_  = ~A202 & ~A200;
  assign \new_[49591]_  = A233 & A232;
  assign \new_[49592]_  = \new_[49591]_  & \new_[49588]_ ;
  assign \new_[49593]_  = \new_[49592]_  & \new_[49585]_ ;
  assign \new_[49596]_  = ~A235 & ~A234;
  assign \new_[49599]_  = A266 & A265;
  assign \new_[49600]_  = \new_[49599]_  & \new_[49596]_ ;
  assign \new_[49603]_  = ~A268 & ~A267;
  assign \new_[49606]_  = A300 & A298;
  assign \new_[49607]_  = \new_[49606]_  & \new_[49603]_ ;
  assign \new_[49608]_  = \new_[49607]_  & \new_[49600]_ ;
  assign \new_[49612]_  = ~A199 & A167;
  assign \new_[49613]_  = A168 & \new_[49612]_ ;
  assign \new_[49616]_  = ~A202 & ~A200;
  assign \new_[49619]_  = A233 & A232;
  assign \new_[49620]_  = \new_[49619]_  & \new_[49616]_ ;
  assign \new_[49621]_  = \new_[49620]_  & \new_[49613]_ ;
  assign \new_[49624]_  = ~A235 & ~A234;
  assign \new_[49627]_  = ~A266 & ~A265;
  assign \new_[49628]_  = \new_[49627]_  & \new_[49624]_ ;
  assign \new_[49631]_  = A298 & ~A268;
  assign \new_[49634]_  = A302 & ~A299;
  assign \new_[49635]_  = \new_[49634]_  & \new_[49631]_ ;
  assign \new_[49636]_  = \new_[49635]_  & \new_[49628]_ ;
  assign \new_[49640]_  = ~A199 & A167;
  assign \new_[49641]_  = A168 & \new_[49640]_ ;
  assign \new_[49644]_  = ~A202 & ~A200;
  assign \new_[49647]_  = A233 & A232;
  assign \new_[49648]_  = \new_[49647]_  & \new_[49644]_ ;
  assign \new_[49649]_  = \new_[49648]_  & \new_[49641]_ ;
  assign \new_[49652]_  = ~A235 & ~A234;
  assign \new_[49655]_  = ~A266 & ~A265;
  assign \new_[49656]_  = \new_[49655]_  & \new_[49652]_ ;
  assign \new_[49659]_  = ~A298 & ~A268;
  assign \new_[49662]_  = A302 & A299;
  assign \new_[49663]_  = \new_[49662]_  & \new_[49659]_ ;
  assign \new_[49664]_  = \new_[49663]_  & \new_[49656]_ ;
  assign \new_[49668]_  = ~A199 & A167;
  assign \new_[49669]_  = A168 & \new_[49668]_ ;
  assign \new_[49672]_  = ~A202 & ~A200;
  assign \new_[49675]_  = ~A233 & ~A232;
  assign \new_[49676]_  = \new_[49675]_  & \new_[49672]_ ;
  assign \new_[49677]_  = \new_[49676]_  & \new_[49669]_ ;
  assign \new_[49680]_  = A265 & ~A235;
  assign \new_[49683]_  = ~A267 & A266;
  assign \new_[49684]_  = \new_[49683]_  & \new_[49680]_ ;
  assign \new_[49687]_  = A298 & ~A268;
  assign \new_[49690]_  = A302 & ~A299;
  assign \new_[49691]_  = \new_[49690]_  & \new_[49687]_ ;
  assign \new_[49692]_  = \new_[49691]_  & \new_[49684]_ ;
  assign \new_[49696]_  = ~A199 & A167;
  assign \new_[49697]_  = A168 & \new_[49696]_ ;
  assign \new_[49700]_  = ~A202 & ~A200;
  assign \new_[49703]_  = ~A233 & ~A232;
  assign \new_[49704]_  = \new_[49703]_  & \new_[49700]_ ;
  assign \new_[49705]_  = \new_[49704]_  & \new_[49697]_ ;
  assign \new_[49708]_  = A265 & ~A235;
  assign \new_[49711]_  = ~A267 & A266;
  assign \new_[49712]_  = \new_[49711]_  & \new_[49708]_ ;
  assign \new_[49715]_  = ~A298 & ~A268;
  assign \new_[49718]_  = A302 & A299;
  assign \new_[49719]_  = \new_[49718]_  & \new_[49715]_ ;
  assign \new_[49720]_  = \new_[49719]_  & \new_[49712]_ ;
  assign \new_[49724]_  = ~A166 & A167;
  assign \new_[49725]_  = A170 & \new_[49724]_ ;
  assign \new_[49728]_  = ~A202 & ~A201;
  assign \new_[49731]_  = ~A234 & ~A203;
  assign \new_[49732]_  = \new_[49731]_  & \new_[49728]_ ;
  assign \new_[49733]_  = \new_[49732]_  & \new_[49725]_ ;
  assign \new_[49736]_  = ~A236 & ~A235;
  assign \new_[49739]_  = ~A268 & ~A267;
  assign \new_[49740]_  = \new_[49739]_  & \new_[49736]_ ;
  assign \new_[49743]_  = A298 & ~A269;
  assign \new_[49746]_  = A302 & ~A299;
  assign \new_[49747]_  = \new_[49746]_  & \new_[49743]_ ;
  assign \new_[49748]_  = \new_[49747]_  & \new_[49740]_ ;
  assign \new_[49752]_  = ~A166 & A167;
  assign \new_[49753]_  = A170 & \new_[49752]_ ;
  assign \new_[49756]_  = ~A202 & ~A201;
  assign \new_[49759]_  = ~A234 & ~A203;
  assign \new_[49760]_  = \new_[49759]_  & \new_[49756]_ ;
  assign \new_[49761]_  = \new_[49760]_  & \new_[49753]_ ;
  assign \new_[49764]_  = ~A236 & ~A235;
  assign \new_[49767]_  = ~A268 & ~A267;
  assign \new_[49768]_  = \new_[49767]_  & \new_[49764]_ ;
  assign \new_[49771]_  = ~A298 & ~A269;
  assign \new_[49774]_  = A302 & A299;
  assign \new_[49775]_  = \new_[49774]_  & \new_[49771]_ ;
  assign \new_[49776]_  = \new_[49775]_  & \new_[49768]_ ;
  assign \new_[49780]_  = ~A166 & A167;
  assign \new_[49781]_  = A170 & \new_[49780]_ ;
  assign \new_[49784]_  = ~A202 & ~A201;
  assign \new_[49787]_  = ~A234 & ~A203;
  assign \new_[49788]_  = \new_[49787]_  & \new_[49784]_ ;
  assign \new_[49789]_  = \new_[49788]_  & \new_[49781]_ ;
  assign \new_[49792]_  = ~A236 & ~A235;
  assign \new_[49795]_  = A266 & A265;
  assign \new_[49796]_  = \new_[49795]_  & \new_[49792]_ ;
  assign \new_[49799]_  = ~A268 & ~A267;
  assign \new_[49802]_  = A300 & A299;
  assign \new_[49803]_  = \new_[49802]_  & \new_[49799]_ ;
  assign \new_[49804]_  = \new_[49803]_  & \new_[49796]_ ;
  assign \new_[49808]_  = ~A166 & A167;
  assign \new_[49809]_  = A170 & \new_[49808]_ ;
  assign \new_[49812]_  = ~A202 & ~A201;
  assign \new_[49815]_  = ~A234 & ~A203;
  assign \new_[49816]_  = \new_[49815]_  & \new_[49812]_ ;
  assign \new_[49817]_  = \new_[49816]_  & \new_[49809]_ ;
  assign \new_[49820]_  = ~A236 & ~A235;
  assign \new_[49823]_  = A266 & A265;
  assign \new_[49824]_  = \new_[49823]_  & \new_[49820]_ ;
  assign \new_[49827]_  = ~A268 & ~A267;
  assign \new_[49830]_  = A300 & A298;
  assign \new_[49831]_  = \new_[49830]_  & \new_[49827]_ ;
  assign \new_[49832]_  = \new_[49831]_  & \new_[49824]_ ;
  assign \new_[49836]_  = ~A166 & A167;
  assign \new_[49837]_  = A170 & \new_[49836]_ ;
  assign \new_[49840]_  = ~A202 & ~A201;
  assign \new_[49843]_  = ~A234 & ~A203;
  assign \new_[49844]_  = \new_[49843]_  & \new_[49840]_ ;
  assign \new_[49845]_  = \new_[49844]_  & \new_[49837]_ ;
  assign \new_[49848]_  = ~A236 & ~A235;
  assign \new_[49851]_  = ~A266 & ~A265;
  assign \new_[49852]_  = \new_[49851]_  & \new_[49848]_ ;
  assign \new_[49855]_  = A298 & ~A268;
  assign \new_[49858]_  = A302 & ~A299;
  assign \new_[49859]_  = \new_[49858]_  & \new_[49855]_ ;
  assign \new_[49860]_  = \new_[49859]_  & \new_[49852]_ ;
  assign \new_[49864]_  = ~A166 & A167;
  assign \new_[49865]_  = A170 & \new_[49864]_ ;
  assign \new_[49868]_  = ~A202 & ~A201;
  assign \new_[49871]_  = ~A234 & ~A203;
  assign \new_[49872]_  = \new_[49871]_  & \new_[49868]_ ;
  assign \new_[49873]_  = \new_[49872]_  & \new_[49865]_ ;
  assign \new_[49876]_  = ~A236 & ~A235;
  assign \new_[49879]_  = ~A266 & ~A265;
  assign \new_[49880]_  = \new_[49879]_  & \new_[49876]_ ;
  assign \new_[49883]_  = ~A298 & ~A268;
  assign \new_[49886]_  = A302 & A299;
  assign \new_[49887]_  = \new_[49886]_  & \new_[49883]_ ;
  assign \new_[49888]_  = \new_[49887]_  & \new_[49880]_ ;
  assign \new_[49892]_  = ~A166 & A167;
  assign \new_[49893]_  = A170 & \new_[49892]_ ;
  assign \new_[49896]_  = ~A202 & ~A201;
  assign \new_[49899]_  = A232 & ~A203;
  assign \new_[49900]_  = \new_[49899]_  & \new_[49896]_ ;
  assign \new_[49901]_  = \new_[49900]_  & \new_[49893]_ ;
  assign \new_[49904]_  = ~A234 & A233;
  assign \new_[49907]_  = ~A267 & ~A235;
  assign \new_[49908]_  = \new_[49907]_  & \new_[49904]_ ;
  assign \new_[49911]_  = ~A269 & ~A268;
  assign \new_[49914]_  = A300 & A299;
  assign \new_[49915]_  = \new_[49914]_  & \new_[49911]_ ;
  assign \new_[49916]_  = \new_[49915]_  & \new_[49908]_ ;
  assign \new_[49920]_  = ~A166 & A167;
  assign \new_[49921]_  = A170 & \new_[49920]_ ;
  assign \new_[49924]_  = ~A202 & ~A201;
  assign \new_[49927]_  = A232 & ~A203;
  assign \new_[49928]_  = \new_[49927]_  & \new_[49924]_ ;
  assign \new_[49929]_  = \new_[49928]_  & \new_[49921]_ ;
  assign \new_[49932]_  = ~A234 & A233;
  assign \new_[49935]_  = ~A267 & ~A235;
  assign \new_[49936]_  = \new_[49935]_  & \new_[49932]_ ;
  assign \new_[49939]_  = ~A269 & ~A268;
  assign \new_[49942]_  = A300 & A298;
  assign \new_[49943]_  = \new_[49942]_  & \new_[49939]_ ;
  assign \new_[49944]_  = \new_[49943]_  & \new_[49936]_ ;
  assign \new_[49948]_  = ~A166 & A167;
  assign \new_[49949]_  = A170 & \new_[49948]_ ;
  assign \new_[49952]_  = ~A202 & ~A201;
  assign \new_[49955]_  = A232 & ~A203;
  assign \new_[49956]_  = \new_[49955]_  & \new_[49952]_ ;
  assign \new_[49957]_  = \new_[49956]_  & \new_[49949]_ ;
  assign \new_[49960]_  = ~A234 & A233;
  assign \new_[49963]_  = A265 & ~A235;
  assign \new_[49964]_  = \new_[49963]_  & \new_[49960]_ ;
  assign \new_[49967]_  = ~A267 & A266;
  assign \new_[49970]_  = A301 & ~A268;
  assign \new_[49971]_  = \new_[49970]_  & \new_[49967]_ ;
  assign \new_[49972]_  = \new_[49971]_  & \new_[49964]_ ;
  assign \new_[49976]_  = ~A166 & A167;
  assign \new_[49977]_  = A170 & \new_[49976]_ ;
  assign \new_[49980]_  = ~A202 & ~A201;
  assign \new_[49983]_  = A232 & ~A203;
  assign \new_[49984]_  = \new_[49983]_  & \new_[49980]_ ;
  assign \new_[49985]_  = \new_[49984]_  & \new_[49977]_ ;
  assign \new_[49988]_  = ~A234 & A233;
  assign \new_[49991]_  = ~A265 & ~A235;
  assign \new_[49992]_  = \new_[49991]_  & \new_[49988]_ ;
  assign \new_[49995]_  = ~A268 & ~A266;
  assign \new_[49998]_  = A300 & A299;
  assign \new_[49999]_  = \new_[49998]_  & \new_[49995]_ ;
  assign \new_[50000]_  = \new_[49999]_  & \new_[49992]_ ;
  assign \new_[50004]_  = ~A166 & A167;
  assign \new_[50005]_  = A170 & \new_[50004]_ ;
  assign \new_[50008]_  = ~A202 & ~A201;
  assign \new_[50011]_  = A232 & ~A203;
  assign \new_[50012]_  = \new_[50011]_  & \new_[50008]_ ;
  assign \new_[50013]_  = \new_[50012]_  & \new_[50005]_ ;
  assign \new_[50016]_  = ~A234 & A233;
  assign \new_[50019]_  = ~A265 & ~A235;
  assign \new_[50020]_  = \new_[50019]_  & \new_[50016]_ ;
  assign \new_[50023]_  = ~A268 & ~A266;
  assign \new_[50026]_  = A300 & A298;
  assign \new_[50027]_  = \new_[50026]_  & \new_[50023]_ ;
  assign \new_[50028]_  = \new_[50027]_  & \new_[50020]_ ;
  assign \new_[50032]_  = ~A166 & A167;
  assign \new_[50033]_  = A170 & \new_[50032]_ ;
  assign \new_[50036]_  = ~A202 & ~A201;
  assign \new_[50039]_  = ~A232 & ~A203;
  assign \new_[50040]_  = \new_[50039]_  & \new_[50036]_ ;
  assign \new_[50041]_  = \new_[50040]_  & \new_[50033]_ ;
  assign \new_[50044]_  = ~A235 & ~A233;
  assign \new_[50047]_  = ~A268 & ~A267;
  assign \new_[50048]_  = \new_[50047]_  & \new_[50044]_ ;
  assign \new_[50051]_  = A298 & ~A269;
  assign \new_[50054]_  = A302 & ~A299;
  assign \new_[50055]_  = \new_[50054]_  & \new_[50051]_ ;
  assign \new_[50056]_  = \new_[50055]_  & \new_[50048]_ ;
  assign \new_[50060]_  = ~A166 & A167;
  assign \new_[50061]_  = A170 & \new_[50060]_ ;
  assign \new_[50064]_  = ~A202 & ~A201;
  assign \new_[50067]_  = ~A232 & ~A203;
  assign \new_[50068]_  = \new_[50067]_  & \new_[50064]_ ;
  assign \new_[50069]_  = \new_[50068]_  & \new_[50061]_ ;
  assign \new_[50072]_  = ~A235 & ~A233;
  assign \new_[50075]_  = ~A268 & ~A267;
  assign \new_[50076]_  = \new_[50075]_  & \new_[50072]_ ;
  assign \new_[50079]_  = ~A298 & ~A269;
  assign \new_[50082]_  = A302 & A299;
  assign \new_[50083]_  = \new_[50082]_  & \new_[50079]_ ;
  assign \new_[50084]_  = \new_[50083]_  & \new_[50076]_ ;
  assign \new_[50088]_  = ~A166 & A167;
  assign \new_[50089]_  = A170 & \new_[50088]_ ;
  assign \new_[50092]_  = ~A202 & ~A201;
  assign \new_[50095]_  = ~A232 & ~A203;
  assign \new_[50096]_  = \new_[50095]_  & \new_[50092]_ ;
  assign \new_[50097]_  = \new_[50096]_  & \new_[50089]_ ;
  assign \new_[50100]_  = ~A235 & ~A233;
  assign \new_[50103]_  = A266 & A265;
  assign \new_[50104]_  = \new_[50103]_  & \new_[50100]_ ;
  assign \new_[50107]_  = ~A268 & ~A267;
  assign \new_[50110]_  = A300 & A299;
  assign \new_[50111]_  = \new_[50110]_  & \new_[50107]_ ;
  assign \new_[50112]_  = \new_[50111]_  & \new_[50104]_ ;
  assign \new_[50116]_  = ~A166 & A167;
  assign \new_[50117]_  = A170 & \new_[50116]_ ;
  assign \new_[50120]_  = ~A202 & ~A201;
  assign \new_[50123]_  = ~A232 & ~A203;
  assign \new_[50124]_  = \new_[50123]_  & \new_[50120]_ ;
  assign \new_[50125]_  = \new_[50124]_  & \new_[50117]_ ;
  assign \new_[50128]_  = ~A235 & ~A233;
  assign \new_[50131]_  = A266 & A265;
  assign \new_[50132]_  = \new_[50131]_  & \new_[50128]_ ;
  assign \new_[50135]_  = ~A268 & ~A267;
  assign \new_[50138]_  = A300 & A298;
  assign \new_[50139]_  = \new_[50138]_  & \new_[50135]_ ;
  assign \new_[50140]_  = \new_[50139]_  & \new_[50132]_ ;
  assign \new_[50144]_  = ~A166 & A167;
  assign \new_[50145]_  = A170 & \new_[50144]_ ;
  assign \new_[50148]_  = ~A202 & ~A201;
  assign \new_[50151]_  = ~A232 & ~A203;
  assign \new_[50152]_  = \new_[50151]_  & \new_[50148]_ ;
  assign \new_[50153]_  = \new_[50152]_  & \new_[50145]_ ;
  assign \new_[50156]_  = ~A235 & ~A233;
  assign \new_[50159]_  = ~A266 & ~A265;
  assign \new_[50160]_  = \new_[50159]_  & \new_[50156]_ ;
  assign \new_[50163]_  = A298 & ~A268;
  assign \new_[50166]_  = A302 & ~A299;
  assign \new_[50167]_  = \new_[50166]_  & \new_[50163]_ ;
  assign \new_[50168]_  = \new_[50167]_  & \new_[50160]_ ;
  assign \new_[50172]_  = ~A166 & A167;
  assign \new_[50173]_  = A170 & \new_[50172]_ ;
  assign \new_[50176]_  = ~A202 & ~A201;
  assign \new_[50179]_  = ~A232 & ~A203;
  assign \new_[50180]_  = \new_[50179]_  & \new_[50176]_ ;
  assign \new_[50181]_  = \new_[50180]_  & \new_[50173]_ ;
  assign \new_[50184]_  = ~A235 & ~A233;
  assign \new_[50187]_  = ~A266 & ~A265;
  assign \new_[50188]_  = \new_[50187]_  & \new_[50184]_ ;
  assign \new_[50191]_  = ~A298 & ~A268;
  assign \new_[50194]_  = A302 & A299;
  assign \new_[50195]_  = \new_[50194]_  & \new_[50191]_ ;
  assign \new_[50196]_  = \new_[50195]_  & \new_[50188]_ ;
  assign \new_[50200]_  = ~A166 & A167;
  assign \new_[50201]_  = A170 & \new_[50200]_ ;
  assign \new_[50204]_  = A200 & A199;
  assign \new_[50207]_  = ~A202 & ~A201;
  assign \new_[50208]_  = \new_[50207]_  & \new_[50204]_ ;
  assign \new_[50209]_  = \new_[50208]_  & \new_[50201]_ ;
  assign \new_[50212]_  = ~A235 & ~A234;
  assign \new_[50215]_  = ~A267 & ~A236;
  assign \new_[50216]_  = \new_[50215]_  & \new_[50212]_ ;
  assign \new_[50219]_  = ~A269 & ~A268;
  assign \new_[50222]_  = A300 & A299;
  assign \new_[50223]_  = \new_[50222]_  & \new_[50219]_ ;
  assign \new_[50224]_  = \new_[50223]_  & \new_[50216]_ ;
  assign \new_[50228]_  = ~A166 & A167;
  assign \new_[50229]_  = A170 & \new_[50228]_ ;
  assign \new_[50232]_  = A200 & A199;
  assign \new_[50235]_  = ~A202 & ~A201;
  assign \new_[50236]_  = \new_[50235]_  & \new_[50232]_ ;
  assign \new_[50237]_  = \new_[50236]_  & \new_[50229]_ ;
  assign \new_[50240]_  = ~A235 & ~A234;
  assign \new_[50243]_  = ~A267 & ~A236;
  assign \new_[50244]_  = \new_[50243]_  & \new_[50240]_ ;
  assign \new_[50247]_  = ~A269 & ~A268;
  assign \new_[50250]_  = A300 & A298;
  assign \new_[50251]_  = \new_[50250]_  & \new_[50247]_ ;
  assign \new_[50252]_  = \new_[50251]_  & \new_[50244]_ ;
  assign \new_[50256]_  = ~A166 & A167;
  assign \new_[50257]_  = A170 & \new_[50256]_ ;
  assign \new_[50260]_  = A200 & A199;
  assign \new_[50263]_  = ~A202 & ~A201;
  assign \new_[50264]_  = \new_[50263]_  & \new_[50260]_ ;
  assign \new_[50265]_  = \new_[50264]_  & \new_[50257]_ ;
  assign \new_[50268]_  = ~A235 & ~A234;
  assign \new_[50271]_  = A265 & ~A236;
  assign \new_[50272]_  = \new_[50271]_  & \new_[50268]_ ;
  assign \new_[50275]_  = ~A267 & A266;
  assign \new_[50278]_  = A301 & ~A268;
  assign \new_[50279]_  = \new_[50278]_  & \new_[50275]_ ;
  assign \new_[50280]_  = \new_[50279]_  & \new_[50272]_ ;
  assign \new_[50284]_  = ~A166 & A167;
  assign \new_[50285]_  = A170 & \new_[50284]_ ;
  assign \new_[50288]_  = A200 & A199;
  assign \new_[50291]_  = ~A202 & ~A201;
  assign \new_[50292]_  = \new_[50291]_  & \new_[50288]_ ;
  assign \new_[50293]_  = \new_[50292]_  & \new_[50285]_ ;
  assign \new_[50296]_  = ~A235 & ~A234;
  assign \new_[50299]_  = ~A265 & ~A236;
  assign \new_[50300]_  = \new_[50299]_  & \new_[50296]_ ;
  assign \new_[50303]_  = ~A268 & ~A266;
  assign \new_[50306]_  = A300 & A299;
  assign \new_[50307]_  = \new_[50306]_  & \new_[50303]_ ;
  assign \new_[50308]_  = \new_[50307]_  & \new_[50300]_ ;
  assign \new_[50312]_  = ~A166 & A167;
  assign \new_[50313]_  = A170 & \new_[50312]_ ;
  assign \new_[50316]_  = A200 & A199;
  assign \new_[50319]_  = ~A202 & ~A201;
  assign \new_[50320]_  = \new_[50319]_  & \new_[50316]_ ;
  assign \new_[50321]_  = \new_[50320]_  & \new_[50313]_ ;
  assign \new_[50324]_  = ~A235 & ~A234;
  assign \new_[50327]_  = ~A265 & ~A236;
  assign \new_[50328]_  = \new_[50327]_  & \new_[50324]_ ;
  assign \new_[50331]_  = ~A268 & ~A266;
  assign \new_[50334]_  = A300 & A298;
  assign \new_[50335]_  = \new_[50334]_  & \new_[50331]_ ;
  assign \new_[50336]_  = \new_[50335]_  & \new_[50328]_ ;
  assign \new_[50340]_  = ~A166 & A167;
  assign \new_[50341]_  = A170 & \new_[50340]_ ;
  assign \new_[50344]_  = A200 & A199;
  assign \new_[50347]_  = ~A202 & ~A201;
  assign \new_[50348]_  = \new_[50347]_  & \new_[50344]_ ;
  assign \new_[50349]_  = \new_[50348]_  & \new_[50341]_ ;
  assign \new_[50352]_  = A233 & A232;
  assign \new_[50355]_  = ~A235 & ~A234;
  assign \new_[50356]_  = \new_[50355]_  & \new_[50352]_ ;
  assign \new_[50359]_  = ~A268 & ~A267;
  assign \new_[50362]_  = A301 & ~A269;
  assign \new_[50363]_  = \new_[50362]_  & \new_[50359]_ ;
  assign \new_[50364]_  = \new_[50363]_  & \new_[50356]_ ;
  assign \new_[50368]_  = ~A166 & A167;
  assign \new_[50369]_  = A170 & \new_[50368]_ ;
  assign \new_[50372]_  = A200 & A199;
  assign \new_[50375]_  = ~A202 & ~A201;
  assign \new_[50376]_  = \new_[50375]_  & \new_[50372]_ ;
  assign \new_[50377]_  = \new_[50376]_  & \new_[50369]_ ;
  assign \new_[50380]_  = A233 & A232;
  assign \new_[50383]_  = ~A235 & ~A234;
  assign \new_[50384]_  = \new_[50383]_  & \new_[50380]_ ;
  assign \new_[50387]_  = ~A266 & ~A265;
  assign \new_[50390]_  = A301 & ~A268;
  assign \new_[50391]_  = \new_[50390]_  & \new_[50387]_ ;
  assign \new_[50392]_  = \new_[50391]_  & \new_[50384]_ ;
  assign \new_[50396]_  = ~A166 & A167;
  assign \new_[50397]_  = A170 & \new_[50396]_ ;
  assign \new_[50400]_  = A200 & A199;
  assign \new_[50403]_  = ~A202 & ~A201;
  assign \new_[50404]_  = \new_[50403]_  & \new_[50400]_ ;
  assign \new_[50405]_  = \new_[50404]_  & \new_[50397]_ ;
  assign \new_[50408]_  = ~A233 & ~A232;
  assign \new_[50411]_  = ~A267 & ~A235;
  assign \new_[50412]_  = \new_[50411]_  & \new_[50408]_ ;
  assign \new_[50415]_  = ~A269 & ~A268;
  assign \new_[50418]_  = A300 & A299;
  assign \new_[50419]_  = \new_[50418]_  & \new_[50415]_ ;
  assign \new_[50420]_  = \new_[50419]_  & \new_[50412]_ ;
  assign \new_[50424]_  = ~A166 & A167;
  assign \new_[50425]_  = A170 & \new_[50424]_ ;
  assign \new_[50428]_  = A200 & A199;
  assign \new_[50431]_  = ~A202 & ~A201;
  assign \new_[50432]_  = \new_[50431]_  & \new_[50428]_ ;
  assign \new_[50433]_  = \new_[50432]_  & \new_[50425]_ ;
  assign \new_[50436]_  = ~A233 & ~A232;
  assign \new_[50439]_  = ~A267 & ~A235;
  assign \new_[50440]_  = \new_[50439]_  & \new_[50436]_ ;
  assign \new_[50443]_  = ~A269 & ~A268;
  assign \new_[50446]_  = A300 & A298;
  assign \new_[50447]_  = \new_[50446]_  & \new_[50443]_ ;
  assign \new_[50448]_  = \new_[50447]_  & \new_[50440]_ ;
  assign \new_[50452]_  = ~A166 & A167;
  assign \new_[50453]_  = A170 & \new_[50452]_ ;
  assign \new_[50456]_  = A200 & A199;
  assign \new_[50459]_  = ~A202 & ~A201;
  assign \new_[50460]_  = \new_[50459]_  & \new_[50456]_ ;
  assign \new_[50461]_  = \new_[50460]_  & \new_[50453]_ ;
  assign \new_[50464]_  = ~A233 & ~A232;
  assign \new_[50467]_  = A265 & ~A235;
  assign \new_[50468]_  = \new_[50467]_  & \new_[50464]_ ;
  assign \new_[50471]_  = ~A267 & A266;
  assign \new_[50474]_  = A301 & ~A268;
  assign \new_[50475]_  = \new_[50474]_  & \new_[50471]_ ;
  assign \new_[50476]_  = \new_[50475]_  & \new_[50468]_ ;
  assign \new_[50480]_  = ~A166 & A167;
  assign \new_[50481]_  = A170 & \new_[50480]_ ;
  assign \new_[50484]_  = A200 & A199;
  assign \new_[50487]_  = ~A202 & ~A201;
  assign \new_[50488]_  = \new_[50487]_  & \new_[50484]_ ;
  assign \new_[50489]_  = \new_[50488]_  & \new_[50481]_ ;
  assign \new_[50492]_  = ~A233 & ~A232;
  assign \new_[50495]_  = ~A265 & ~A235;
  assign \new_[50496]_  = \new_[50495]_  & \new_[50492]_ ;
  assign \new_[50499]_  = ~A268 & ~A266;
  assign \new_[50502]_  = A300 & A299;
  assign \new_[50503]_  = \new_[50502]_  & \new_[50499]_ ;
  assign \new_[50504]_  = \new_[50503]_  & \new_[50496]_ ;
  assign \new_[50508]_  = ~A166 & A167;
  assign \new_[50509]_  = A170 & \new_[50508]_ ;
  assign \new_[50512]_  = A200 & A199;
  assign \new_[50515]_  = ~A202 & ~A201;
  assign \new_[50516]_  = \new_[50515]_  & \new_[50512]_ ;
  assign \new_[50517]_  = \new_[50516]_  & \new_[50509]_ ;
  assign \new_[50520]_  = ~A233 & ~A232;
  assign \new_[50523]_  = ~A265 & ~A235;
  assign \new_[50524]_  = \new_[50523]_  & \new_[50520]_ ;
  assign \new_[50527]_  = ~A268 & ~A266;
  assign \new_[50530]_  = A300 & A298;
  assign \new_[50531]_  = \new_[50530]_  & \new_[50527]_ ;
  assign \new_[50532]_  = \new_[50531]_  & \new_[50524]_ ;
  assign \new_[50536]_  = ~A166 & A167;
  assign \new_[50537]_  = A170 & \new_[50536]_ ;
  assign \new_[50540]_  = ~A200 & ~A199;
  assign \new_[50543]_  = ~A234 & ~A202;
  assign \new_[50544]_  = \new_[50543]_  & \new_[50540]_ ;
  assign \new_[50545]_  = \new_[50544]_  & \new_[50537]_ ;
  assign \new_[50548]_  = ~A236 & ~A235;
  assign \new_[50551]_  = ~A268 & ~A267;
  assign \new_[50552]_  = \new_[50551]_  & \new_[50548]_ ;
  assign \new_[50555]_  = A298 & ~A269;
  assign \new_[50558]_  = A302 & ~A299;
  assign \new_[50559]_  = \new_[50558]_  & \new_[50555]_ ;
  assign \new_[50560]_  = \new_[50559]_  & \new_[50552]_ ;
  assign \new_[50564]_  = ~A166 & A167;
  assign \new_[50565]_  = A170 & \new_[50564]_ ;
  assign \new_[50568]_  = ~A200 & ~A199;
  assign \new_[50571]_  = ~A234 & ~A202;
  assign \new_[50572]_  = \new_[50571]_  & \new_[50568]_ ;
  assign \new_[50573]_  = \new_[50572]_  & \new_[50565]_ ;
  assign \new_[50576]_  = ~A236 & ~A235;
  assign \new_[50579]_  = ~A268 & ~A267;
  assign \new_[50580]_  = \new_[50579]_  & \new_[50576]_ ;
  assign \new_[50583]_  = ~A298 & ~A269;
  assign \new_[50586]_  = A302 & A299;
  assign \new_[50587]_  = \new_[50586]_  & \new_[50583]_ ;
  assign \new_[50588]_  = \new_[50587]_  & \new_[50580]_ ;
  assign \new_[50592]_  = ~A166 & A167;
  assign \new_[50593]_  = A170 & \new_[50592]_ ;
  assign \new_[50596]_  = ~A200 & ~A199;
  assign \new_[50599]_  = ~A234 & ~A202;
  assign \new_[50600]_  = \new_[50599]_  & \new_[50596]_ ;
  assign \new_[50601]_  = \new_[50600]_  & \new_[50593]_ ;
  assign \new_[50604]_  = ~A236 & ~A235;
  assign \new_[50607]_  = A266 & A265;
  assign \new_[50608]_  = \new_[50607]_  & \new_[50604]_ ;
  assign \new_[50611]_  = ~A268 & ~A267;
  assign \new_[50614]_  = A300 & A299;
  assign \new_[50615]_  = \new_[50614]_  & \new_[50611]_ ;
  assign \new_[50616]_  = \new_[50615]_  & \new_[50608]_ ;
  assign \new_[50620]_  = ~A166 & A167;
  assign \new_[50621]_  = A170 & \new_[50620]_ ;
  assign \new_[50624]_  = ~A200 & ~A199;
  assign \new_[50627]_  = ~A234 & ~A202;
  assign \new_[50628]_  = \new_[50627]_  & \new_[50624]_ ;
  assign \new_[50629]_  = \new_[50628]_  & \new_[50621]_ ;
  assign \new_[50632]_  = ~A236 & ~A235;
  assign \new_[50635]_  = A266 & A265;
  assign \new_[50636]_  = \new_[50635]_  & \new_[50632]_ ;
  assign \new_[50639]_  = ~A268 & ~A267;
  assign \new_[50642]_  = A300 & A298;
  assign \new_[50643]_  = \new_[50642]_  & \new_[50639]_ ;
  assign \new_[50644]_  = \new_[50643]_  & \new_[50636]_ ;
  assign \new_[50648]_  = ~A166 & A167;
  assign \new_[50649]_  = A170 & \new_[50648]_ ;
  assign \new_[50652]_  = ~A200 & ~A199;
  assign \new_[50655]_  = ~A234 & ~A202;
  assign \new_[50656]_  = \new_[50655]_  & \new_[50652]_ ;
  assign \new_[50657]_  = \new_[50656]_  & \new_[50649]_ ;
  assign \new_[50660]_  = ~A236 & ~A235;
  assign \new_[50663]_  = ~A266 & ~A265;
  assign \new_[50664]_  = \new_[50663]_  & \new_[50660]_ ;
  assign \new_[50667]_  = A298 & ~A268;
  assign \new_[50670]_  = A302 & ~A299;
  assign \new_[50671]_  = \new_[50670]_  & \new_[50667]_ ;
  assign \new_[50672]_  = \new_[50671]_  & \new_[50664]_ ;
  assign \new_[50676]_  = ~A166 & A167;
  assign \new_[50677]_  = A170 & \new_[50676]_ ;
  assign \new_[50680]_  = ~A200 & ~A199;
  assign \new_[50683]_  = ~A234 & ~A202;
  assign \new_[50684]_  = \new_[50683]_  & \new_[50680]_ ;
  assign \new_[50685]_  = \new_[50684]_  & \new_[50677]_ ;
  assign \new_[50688]_  = ~A236 & ~A235;
  assign \new_[50691]_  = ~A266 & ~A265;
  assign \new_[50692]_  = \new_[50691]_  & \new_[50688]_ ;
  assign \new_[50695]_  = ~A298 & ~A268;
  assign \new_[50698]_  = A302 & A299;
  assign \new_[50699]_  = \new_[50698]_  & \new_[50695]_ ;
  assign \new_[50700]_  = \new_[50699]_  & \new_[50692]_ ;
  assign \new_[50704]_  = ~A166 & A167;
  assign \new_[50705]_  = A170 & \new_[50704]_ ;
  assign \new_[50708]_  = ~A200 & ~A199;
  assign \new_[50711]_  = A232 & ~A202;
  assign \new_[50712]_  = \new_[50711]_  & \new_[50708]_ ;
  assign \new_[50713]_  = \new_[50712]_  & \new_[50705]_ ;
  assign \new_[50716]_  = ~A234 & A233;
  assign \new_[50719]_  = ~A267 & ~A235;
  assign \new_[50720]_  = \new_[50719]_  & \new_[50716]_ ;
  assign \new_[50723]_  = ~A269 & ~A268;
  assign \new_[50726]_  = A300 & A299;
  assign \new_[50727]_  = \new_[50726]_  & \new_[50723]_ ;
  assign \new_[50728]_  = \new_[50727]_  & \new_[50720]_ ;
  assign \new_[50732]_  = ~A166 & A167;
  assign \new_[50733]_  = A170 & \new_[50732]_ ;
  assign \new_[50736]_  = ~A200 & ~A199;
  assign \new_[50739]_  = A232 & ~A202;
  assign \new_[50740]_  = \new_[50739]_  & \new_[50736]_ ;
  assign \new_[50741]_  = \new_[50740]_  & \new_[50733]_ ;
  assign \new_[50744]_  = ~A234 & A233;
  assign \new_[50747]_  = ~A267 & ~A235;
  assign \new_[50748]_  = \new_[50747]_  & \new_[50744]_ ;
  assign \new_[50751]_  = ~A269 & ~A268;
  assign \new_[50754]_  = A300 & A298;
  assign \new_[50755]_  = \new_[50754]_  & \new_[50751]_ ;
  assign \new_[50756]_  = \new_[50755]_  & \new_[50748]_ ;
  assign \new_[50760]_  = ~A166 & A167;
  assign \new_[50761]_  = A170 & \new_[50760]_ ;
  assign \new_[50764]_  = ~A200 & ~A199;
  assign \new_[50767]_  = A232 & ~A202;
  assign \new_[50768]_  = \new_[50767]_  & \new_[50764]_ ;
  assign \new_[50769]_  = \new_[50768]_  & \new_[50761]_ ;
  assign \new_[50772]_  = ~A234 & A233;
  assign \new_[50775]_  = A265 & ~A235;
  assign \new_[50776]_  = \new_[50775]_  & \new_[50772]_ ;
  assign \new_[50779]_  = ~A267 & A266;
  assign \new_[50782]_  = A301 & ~A268;
  assign \new_[50783]_  = \new_[50782]_  & \new_[50779]_ ;
  assign \new_[50784]_  = \new_[50783]_  & \new_[50776]_ ;
  assign \new_[50788]_  = ~A166 & A167;
  assign \new_[50789]_  = A170 & \new_[50788]_ ;
  assign \new_[50792]_  = ~A200 & ~A199;
  assign \new_[50795]_  = A232 & ~A202;
  assign \new_[50796]_  = \new_[50795]_  & \new_[50792]_ ;
  assign \new_[50797]_  = \new_[50796]_  & \new_[50789]_ ;
  assign \new_[50800]_  = ~A234 & A233;
  assign \new_[50803]_  = ~A265 & ~A235;
  assign \new_[50804]_  = \new_[50803]_  & \new_[50800]_ ;
  assign \new_[50807]_  = ~A268 & ~A266;
  assign \new_[50810]_  = A300 & A299;
  assign \new_[50811]_  = \new_[50810]_  & \new_[50807]_ ;
  assign \new_[50812]_  = \new_[50811]_  & \new_[50804]_ ;
  assign \new_[50816]_  = ~A166 & A167;
  assign \new_[50817]_  = A170 & \new_[50816]_ ;
  assign \new_[50820]_  = ~A200 & ~A199;
  assign \new_[50823]_  = A232 & ~A202;
  assign \new_[50824]_  = \new_[50823]_  & \new_[50820]_ ;
  assign \new_[50825]_  = \new_[50824]_  & \new_[50817]_ ;
  assign \new_[50828]_  = ~A234 & A233;
  assign \new_[50831]_  = ~A265 & ~A235;
  assign \new_[50832]_  = \new_[50831]_  & \new_[50828]_ ;
  assign \new_[50835]_  = ~A268 & ~A266;
  assign \new_[50838]_  = A300 & A298;
  assign \new_[50839]_  = \new_[50838]_  & \new_[50835]_ ;
  assign \new_[50840]_  = \new_[50839]_  & \new_[50832]_ ;
  assign \new_[50844]_  = ~A166 & A167;
  assign \new_[50845]_  = A170 & \new_[50844]_ ;
  assign \new_[50848]_  = ~A200 & ~A199;
  assign \new_[50851]_  = ~A232 & ~A202;
  assign \new_[50852]_  = \new_[50851]_  & \new_[50848]_ ;
  assign \new_[50853]_  = \new_[50852]_  & \new_[50845]_ ;
  assign \new_[50856]_  = ~A235 & ~A233;
  assign \new_[50859]_  = ~A268 & ~A267;
  assign \new_[50860]_  = \new_[50859]_  & \new_[50856]_ ;
  assign \new_[50863]_  = A298 & ~A269;
  assign \new_[50866]_  = A302 & ~A299;
  assign \new_[50867]_  = \new_[50866]_  & \new_[50863]_ ;
  assign \new_[50868]_  = \new_[50867]_  & \new_[50860]_ ;
  assign \new_[50872]_  = ~A166 & A167;
  assign \new_[50873]_  = A170 & \new_[50872]_ ;
  assign \new_[50876]_  = ~A200 & ~A199;
  assign \new_[50879]_  = ~A232 & ~A202;
  assign \new_[50880]_  = \new_[50879]_  & \new_[50876]_ ;
  assign \new_[50881]_  = \new_[50880]_  & \new_[50873]_ ;
  assign \new_[50884]_  = ~A235 & ~A233;
  assign \new_[50887]_  = ~A268 & ~A267;
  assign \new_[50888]_  = \new_[50887]_  & \new_[50884]_ ;
  assign \new_[50891]_  = ~A298 & ~A269;
  assign \new_[50894]_  = A302 & A299;
  assign \new_[50895]_  = \new_[50894]_  & \new_[50891]_ ;
  assign \new_[50896]_  = \new_[50895]_  & \new_[50888]_ ;
  assign \new_[50900]_  = ~A166 & A167;
  assign \new_[50901]_  = A170 & \new_[50900]_ ;
  assign \new_[50904]_  = ~A200 & ~A199;
  assign \new_[50907]_  = ~A232 & ~A202;
  assign \new_[50908]_  = \new_[50907]_  & \new_[50904]_ ;
  assign \new_[50909]_  = \new_[50908]_  & \new_[50901]_ ;
  assign \new_[50912]_  = ~A235 & ~A233;
  assign \new_[50915]_  = A266 & A265;
  assign \new_[50916]_  = \new_[50915]_  & \new_[50912]_ ;
  assign \new_[50919]_  = ~A268 & ~A267;
  assign \new_[50922]_  = A300 & A299;
  assign \new_[50923]_  = \new_[50922]_  & \new_[50919]_ ;
  assign \new_[50924]_  = \new_[50923]_  & \new_[50916]_ ;
  assign \new_[50928]_  = ~A166 & A167;
  assign \new_[50929]_  = A170 & \new_[50928]_ ;
  assign \new_[50932]_  = ~A200 & ~A199;
  assign \new_[50935]_  = ~A232 & ~A202;
  assign \new_[50936]_  = \new_[50935]_  & \new_[50932]_ ;
  assign \new_[50937]_  = \new_[50936]_  & \new_[50929]_ ;
  assign \new_[50940]_  = ~A235 & ~A233;
  assign \new_[50943]_  = A266 & A265;
  assign \new_[50944]_  = \new_[50943]_  & \new_[50940]_ ;
  assign \new_[50947]_  = ~A268 & ~A267;
  assign \new_[50950]_  = A300 & A298;
  assign \new_[50951]_  = \new_[50950]_  & \new_[50947]_ ;
  assign \new_[50952]_  = \new_[50951]_  & \new_[50944]_ ;
  assign \new_[50956]_  = ~A166 & A167;
  assign \new_[50957]_  = A170 & \new_[50956]_ ;
  assign \new_[50960]_  = ~A200 & ~A199;
  assign \new_[50963]_  = ~A232 & ~A202;
  assign \new_[50964]_  = \new_[50963]_  & \new_[50960]_ ;
  assign \new_[50965]_  = \new_[50964]_  & \new_[50957]_ ;
  assign \new_[50968]_  = ~A235 & ~A233;
  assign \new_[50971]_  = ~A266 & ~A265;
  assign \new_[50972]_  = \new_[50971]_  & \new_[50968]_ ;
  assign \new_[50975]_  = A298 & ~A268;
  assign \new_[50978]_  = A302 & ~A299;
  assign \new_[50979]_  = \new_[50978]_  & \new_[50975]_ ;
  assign \new_[50980]_  = \new_[50979]_  & \new_[50972]_ ;
  assign \new_[50984]_  = ~A166 & A167;
  assign \new_[50985]_  = A170 & \new_[50984]_ ;
  assign \new_[50988]_  = ~A200 & ~A199;
  assign \new_[50991]_  = ~A232 & ~A202;
  assign \new_[50992]_  = \new_[50991]_  & \new_[50988]_ ;
  assign \new_[50993]_  = \new_[50992]_  & \new_[50985]_ ;
  assign \new_[50996]_  = ~A235 & ~A233;
  assign \new_[50999]_  = ~A266 & ~A265;
  assign \new_[51000]_  = \new_[50999]_  & \new_[50996]_ ;
  assign \new_[51003]_  = ~A298 & ~A268;
  assign \new_[51006]_  = A302 & A299;
  assign \new_[51007]_  = \new_[51006]_  & \new_[51003]_ ;
  assign \new_[51008]_  = \new_[51007]_  & \new_[51000]_ ;
  assign \new_[51012]_  = A166 & ~A167;
  assign \new_[51013]_  = A170 & \new_[51012]_ ;
  assign \new_[51016]_  = ~A202 & ~A201;
  assign \new_[51019]_  = ~A234 & ~A203;
  assign \new_[51020]_  = \new_[51019]_  & \new_[51016]_ ;
  assign \new_[51021]_  = \new_[51020]_  & \new_[51013]_ ;
  assign \new_[51024]_  = ~A236 & ~A235;
  assign \new_[51027]_  = ~A268 & ~A267;
  assign \new_[51028]_  = \new_[51027]_  & \new_[51024]_ ;
  assign \new_[51031]_  = A298 & ~A269;
  assign \new_[51034]_  = A302 & ~A299;
  assign \new_[51035]_  = \new_[51034]_  & \new_[51031]_ ;
  assign \new_[51036]_  = \new_[51035]_  & \new_[51028]_ ;
  assign \new_[51040]_  = A166 & ~A167;
  assign \new_[51041]_  = A170 & \new_[51040]_ ;
  assign \new_[51044]_  = ~A202 & ~A201;
  assign \new_[51047]_  = ~A234 & ~A203;
  assign \new_[51048]_  = \new_[51047]_  & \new_[51044]_ ;
  assign \new_[51049]_  = \new_[51048]_  & \new_[51041]_ ;
  assign \new_[51052]_  = ~A236 & ~A235;
  assign \new_[51055]_  = ~A268 & ~A267;
  assign \new_[51056]_  = \new_[51055]_  & \new_[51052]_ ;
  assign \new_[51059]_  = ~A298 & ~A269;
  assign \new_[51062]_  = A302 & A299;
  assign \new_[51063]_  = \new_[51062]_  & \new_[51059]_ ;
  assign \new_[51064]_  = \new_[51063]_  & \new_[51056]_ ;
  assign \new_[51068]_  = A166 & ~A167;
  assign \new_[51069]_  = A170 & \new_[51068]_ ;
  assign \new_[51072]_  = ~A202 & ~A201;
  assign \new_[51075]_  = ~A234 & ~A203;
  assign \new_[51076]_  = \new_[51075]_  & \new_[51072]_ ;
  assign \new_[51077]_  = \new_[51076]_  & \new_[51069]_ ;
  assign \new_[51080]_  = ~A236 & ~A235;
  assign \new_[51083]_  = A266 & A265;
  assign \new_[51084]_  = \new_[51083]_  & \new_[51080]_ ;
  assign \new_[51087]_  = ~A268 & ~A267;
  assign \new_[51090]_  = A300 & A299;
  assign \new_[51091]_  = \new_[51090]_  & \new_[51087]_ ;
  assign \new_[51092]_  = \new_[51091]_  & \new_[51084]_ ;
  assign \new_[51096]_  = A166 & ~A167;
  assign \new_[51097]_  = A170 & \new_[51096]_ ;
  assign \new_[51100]_  = ~A202 & ~A201;
  assign \new_[51103]_  = ~A234 & ~A203;
  assign \new_[51104]_  = \new_[51103]_  & \new_[51100]_ ;
  assign \new_[51105]_  = \new_[51104]_  & \new_[51097]_ ;
  assign \new_[51108]_  = ~A236 & ~A235;
  assign \new_[51111]_  = A266 & A265;
  assign \new_[51112]_  = \new_[51111]_  & \new_[51108]_ ;
  assign \new_[51115]_  = ~A268 & ~A267;
  assign \new_[51118]_  = A300 & A298;
  assign \new_[51119]_  = \new_[51118]_  & \new_[51115]_ ;
  assign \new_[51120]_  = \new_[51119]_  & \new_[51112]_ ;
  assign \new_[51124]_  = A166 & ~A167;
  assign \new_[51125]_  = A170 & \new_[51124]_ ;
  assign \new_[51128]_  = ~A202 & ~A201;
  assign \new_[51131]_  = ~A234 & ~A203;
  assign \new_[51132]_  = \new_[51131]_  & \new_[51128]_ ;
  assign \new_[51133]_  = \new_[51132]_  & \new_[51125]_ ;
  assign \new_[51136]_  = ~A236 & ~A235;
  assign \new_[51139]_  = ~A266 & ~A265;
  assign \new_[51140]_  = \new_[51139]_  & \new_[51136]_ ;
  assign \new_[51143]_  = A298 & ~A268;
  assign \new_[51146]_  = A302 & ~A299;
  assign \new_[51147]_  = \new_[51146]_  & \new_[51143]_ ;
  assign \new_[51148]_  = \new_[51147]_  & \new_[51140]_ ;
  assign \new_[51152]_  = A166 & ~A167;
  assign \new_[51153]_  = A170 & \new_[51152]_ ;
  assign \new_[51156]_  = ~A202 & ~A201;
  assign \new_[51159]_  = ~A234 & ~A203;
  assign \new_[51160]_  = \new_[51159]_  & \new_[51156]_ ;
  assign \new_[51161]_  = \new_[51160]_  & \new_[51153]_ ;
  assign \new_[51164]_  = ~A236 & ~A235;
  assign \new_[51167]_  = ~A266 & ~A265;
  assign \new_[51168]_  = \new_[51167]_  & \new_[51164]_ ;
  assign \new_[51171]_  = ~A298 & ~A268;
  assign \new_[51174]_  = A302 & A299;
  assign \new_[51175]_  = \new_[51174]_  & \new_[51171]_ ;
  assign \new_[51176]_  = \new_[51175]_  & \new_[51168]_ ;
  assign \new_[51180]_  = A166 & ~A167;
  assign \new_[51181]_  = A170 & \new_[51180]_ ;
  assign \new_[51184]_  = ~A202 & ~A201;
  assign \new_[51187]_  = A232 & ~A203;
  assign \new_[51188]_  = \new_[51187]_  & \new_[51184]_ ;
  assign \new_[51189]_  = \new_[51188]_  & \new_[51181]_ ;
  assign \new_[51192]_  = ~A234 & A233;
  assign \new_[51195]_  = ~A267 & ~A235;
  assign \new_[51196]_  = \new_[51195]_  & \new_[51192]_ ;
  assign \new_[51199]_  = ~A269 & ~A268;
  assign \new_[51202]_  = A300 & A299;
  assign \new_[51203]_  = \new_[51202]_  & \new_[51199]_ ;
  assign \new_[51204]_  = \new_[51203]_  & \new_[51196]_ ;
  assign \new_[51208]_  = A166 & ~A167;
  assign \new_[51209]_  = A170 & \new_[51208]_ ;
  assign \new_[51212]_  = ~A202 & ~A201;
  assign \new_[51215]_  = A232 & ~A203;
  assign \new_[51216]_  = \new_[51215]_  & \new_[51212]_ ;
  assign \new_[51217]_  = \new_[51216]_  & \new_[51209]_ ;
  assign \new_[51220]_  = ~A234 & A233;
  assign \new_[51223]_  = ~A267 & ~A235;
  assign \new_[51224]_  = \new_[51223]_  & \new_[51220]_ ;
  assign \new_[51227]_  = ~A269 & ~A268;
  assign \new_[51230]_  = A300 & A298;
  assign \new_[51231]_  = \new_[51230]_  & \new_[51227]_ ;
  assign \new_[51232]_  = \new_[51231]_  & \new_[51224]_ ;
  assign \new_[51236]_  = A166 & ~A167;
  assign \new_[51237]_  = A170 & \new_[51236]_ ;
  assign \new_[51240]_  = ~A202 & ~A201;
  assign \new_[51243]_  = A232 & ~A203;
  assign \new_[51244]_  = \new_[51243]_  & \new_[51240]_ ;
  assign \new_[51245]_  = \new_[51244]_  & \new_[51237]_ ;
  assign \new_[51248]_  = ~A234 & A233;
  assign \new_[51251]_  = A265 & ~A235;
  assign \new_[51252]_  = \new_[51251]_  & \new_[51248]_ ;
  assign \new_[51255]_  = ~A267 & A266;
  assign \new_[51258]_  = A301 & ~A268;
  assign \new_[51259]_  = \new_[51258]_  & \new_[51255]_ ;
  assign \new_[51260]_  = \new_[51259]_  & \new_[51252]_ ;
  assign \new_[51264]_  = A166 & ~A167;
  assign \new_[51265]_  = A170 & \new_[51264]_ ;
  assign \new_[51268]_  = ~A202 & ~A201;
  assign \new_[51271]_  = A232 & ~A203;
  assign \new_[51272]_  = \new_[51271]_  & \new_[51268]_ ;
  assign \new_[51273]_  = \new_[51272]_  & \new_[51265]_ ;
  assign \new_[51276]_  = ~A234 & A233;
  assign \new_[51279]_  = ~A265 & ~A235;
  assign \new_[51280]_  = \new_[51279]_  & \new_[51276]_ ;
  assign \new_[51283]_  = ~A268 & ~A266;
  assign \new_[51286]_  = A300 & A299;
  assign \new_[51287]_  = \new_[51286]_  & \new_[51283]_ ;
  assign \new_[51288]_  = \new_[51287]_  & \new_[51280]_ ;
  assign \new_[51292]_  = A166 & ~A167;
  assign \new_[51293]_  = A170 & \new_[51292]_ ;
  assign \new_[51296]_  = ~A202 & ~A201;
  assign \new_[51299]_  = A232 & ~A203;
  assign \new_[51300]_  = \new_[51299]_  & \new_[51296]_ ;
  assign \new_[51301]_  = \new_[51300]_  & \new_[51293]_ ;
  assign \new_[51304]_  = ~A234 & A233;
  assign \new_[51307]_  = ~A265 & ~A235;
  assign \new_[51308]_  = \new_[51307]_  & \new_[51304]_ ;
  assign \new_[51311]_  = ~A268 & ~A266;
  assign \new_[51314]_  = A300 & A298;
  assign \new_[51315]_  = \new_[51314]_  & \new_[51311]_ ;
  assign \new_[51316]_  = \new_[51315]_  & \new_[51308]_ ;
  assign \new_[51320]_  = A166 & ~A167;
  assign \new_[51321]_  = A170 & \new_[51320]_ ;
  assign \new_[51324]_  = ~A202 & ~A201;
  assign \new_[51327]_  = ~A232 & ~A203;
  assign \new_[51328]_  = \new_[51327]_  & \new_[51324]_ ;
  assign \new_[51329]_  = \new_[51328]_  & \new_[51321]_ ;
  assign \new_[51332]_  = ~A235 & ~A233;
  assign \new_[51335]_  = ~A268 & ~A267;
  assign \new_[51336]_  = \new_[51335]_  & \new_[51332]_ ;
  assign \new_[51339]_  = A298 & ~A269;
  assign \new_[51342]_  = A302 & ~A299;
  assign \new_[51343]_  = \new_[51342]_  & \new_[51339]_ ;
  assign \new_[51344]_  = \new_[51343]_  & \new_[51336]_ ;
  assign \new_[51348]_  = A166 & ~A167;
  assign \new_[51349]_  = A170 & \new_[51348]_ ;
  assign \new_[51352]_  = ~A202 & ~A201;
  assign \new_[51355]_  = ~A232 & ~A203;
  assign \new_[51356]_  = \new_[51355]_  & \new_[51352]_ ;
  assign \new_[51357]_  = \new_[51356]_  & \new_[51349]_ ;
  assign \new_[51360]_  = ~A235 & ~A233;
  assign \new_[51363]_  = ~A268 & ~A267;
  assign \new_[51364]_  = \new_[51363]_  & \new_[51360]_ ;
  assign \new_[51367]_  = ~A298 & ~A269;
  assign \new_[51370]_  = A302 & A299;
  assign \new_[51371]_  = \new_[51370]_  & \new_[51367]_ ;
  assign \new_[51372]_  = \new_[51371]_  & \new_[51364]_ ;
  assign \new_[51376]_  = A166 & ~A167;
  assign \new_[51377]_  = A170 & \new_[51376]_ ;
  assign \new_[51380]_  = ~A202 & ~A201;
  assign \new_[51383]_  = ~A232 & ~A203;
  assign \new_[51384]_  = \new_[51383]_  & \new_[51380]_ ;
  assign \new_[51385]_  = \new_[51384]_  & \new_[51377]_ ;
  assign \new_[51388]_  = ~A235 & ~A233;
  assign \new_[51391]_  = A266 & A265;
  assign \new_[51392]_  = \new_[51391]_  & \new_[51388]_ ;
  assign \new_[51395]_  = ~A268 & ~A267;
  assign \new_[51398]_  = A300 & A299;
  assign \new_[51399]_  = \new_[51398]_  & \new_[51395]_ ;
  assign \new_[51400]_  = \new_[51399]_  & \new_[51392]_ ;
  assign \new_[51404]_  = A166 & ~A167;
  assign \new_[51405]_  = A170 & \new_[51404]_ ;
  assign \new_[51408]_  = ~A202 & ~A201;
  assign \new_[51411]_  = ~A232 & ~A203;
  assign \new_[51412]_  = \new_[51411]_  & \new_[51408]_ ;
  assign \new_[51413]_  = \new_[51412]_  & \new_[51405]_ ;
  assign \new_[51416]_  = ~A235 & ~A233;
  assign \new_[51419]_  = A266 & A265;
  assign \new_[51420]_  = \new_[51419]_  & \new_[51416]_ ;
  assign \new_[51423]_  = ~A268 & ~A267;
  assign \new_[51426]_  = A300 & A298;
  assign \new_[51427]_  = \new_[51426]_  & \new_[51423]_ ;
  assign \new_[51428]_  = \new_[51427]_  & \new_[51420]_ ;
  assign \new_[51432]_  = A166 & ~A167;
  assign \new_[51433]_  = A170 & \new_[51432]_ ;
  assign \new_[51436]_  = ~A202 & ~A201;
  assign \new_[51439]_  = ~A232 & ~A203;
  assign \new_[51440]_  = \new_[51439]_  & \new_[51436]_ ;
  assign \new_[51441]_  = \new_[51440]_  & \new_[51433]_ ;
  assign \new_[51444]_  = ~A235 & ~A233;
  assign \new_[51447]_  = ~A266 & ~A265;
  assign \new_[51448]_  = \new_[51447]_  & \new_[51444]_ ;
  assign \new_[51451]_  = A298 & ~A268;
  assign \new_[51454]_  = A302 & ~A299;
  assign \new_[51455]_  = \new_[51454]_  & \new_[51451]_ ;
  assign \new_[51456]_  = \new_[51455]_  & \new_[51448]_ ;
  assign \new_[51460]_  = A166 & ~A167;
  assign \new_[51461]_  = A170 & \new_[51460]_ ;
  assign \new_[51464]_  = ~A202 & ~A201;
  assign \new_[51467]_  = ~A232 & ~A203;
  assign \new_[51468]_  = \new_[51467]_  & \new_[51464]_ ;
  assign \new_[51469]_  = \new_[51468]_  & \new_[51461]_ ;
  assign \new_[51472]_  = ~A235 & ~A233;
  assign \new_[51475]_  = ~A266 & ~A265;
  assign \new_[51476]_  = \new_[51475]_  & \new_[51472]_ ;
  assign \new_[51479]_  = ~A298 & ~A268;
  assign \new_[51482]_  = A302 & A299;
  assign \new_[51483]_  = \new_[51482]_  & \new_[51479]_ ;
  assign \new_[51484]_  = \new_[51483]_  & \new_[51476]_ ;
  assign \new_[51488]_  = A166 & ~A167;
  assign \new_[51489]_  = A170 & \new_[51488]_ ;
  assign \new_[51492]_  = A200 & A199;
  assign \new_[51495]_  = ~A202 & ~A201;
  assign \new_[51496]_  = \new_[51495]_  & \new_[51492]_ ;
  assign \new_[51497]_  = \new_[51496]_  & \new_[51489]_ ;
  assign \new_[51500]_  = ~A235 & ~A234;
  assign \new_[51503]_  = ~A267 & ~A236;
  assign \new_[51504]_  = \new_[51503]_  & \new_[51500]_ ;
  assign \new_[51507]_  = ~A269 & ~A268;
  assign \new_[51510]_  = A300 & A299;
  assign \new_[51511]_  = \new_[51510]_  & \new_[51507]_ ;
  assign \new_[51512]_  = \new_[51511]_  & \new_[51504]_ ;
  assign \new_[51516]_  = A166 & ~A167;
  assign \new_[51517]_  = A170 & \new_[51516]_ ;
  assign \new_[51520]_  = A200 & A199;
  assign \new_[51523]_  = ~A202 & ~A201;
  assign \new_[51524]_  = \new_[51523]_  & \new_[51520]_ ;
  assign \new_[51525]_  = \new_[51524]_  & \new_[51517]_ ;
  assign \new_[51528]_  = ~A235 & ~A234;
  assign \new_[51531]_  = ~A267 & ~A236;
  assign \new_[51532]_  = \new_[51531]_  & \new_[51528]_ ;
  assign \new_[51535]_  = ~A269 & ~A268;
  assign \new_[51538]_  = A300 & A298;
  assign \new_[51539]_  = \new_[51538]_  & \new_[51535]_ ;
  assign \new_[51540]_  = \new_[51539]_  & \new_[51532]_ ;
  assign \new_[51544]_  = A166 & ~A167;
  assign \new_[51545]_  = A170 & \new_[51544]_ ;
  assign \new_[51548]_  = A200 & A199;
  assign \new_[51551]_  = ~A202 & ~A201;
  assign \new_[51552]_  = \new_[51551]_  & \new_[51548]_ ;
  assign \new_[51553]_  = \new_[51552]_  & \new_[51545]_ ;
  assign \new_[51556]_  = ~A235 & ~A234;
  assign \new_[51559]_  = A265 & ~A236;
  assign \new_[51560]_  = \new_[51559]_  & \new_[51556]_ ;
  assign \new_[51563]_  = ~A267 & A266;
  assign \new_[51566]_  = A301 & ~A268;
  assign \new_[51567]_  = \new_[51566]_  & \new_[51563]_ ;
  assign \new_[51568]_  = \new_[51567]_  & \new_[51560]_ ;
  assign \new_[51572]_  = A166 & ~A167;
  assign \new_[51573]_  = A170 & \new_[51572]_ ;
  assign \new_[51576]_  = A200 & A199;
  assign \new_[51579]_  = ~A202 & ~A201;
  assign \new_[51580]_  = \new_[51579]_  & \new_[51576]_ ;
  assign \new_[51581]_  = \new_[51580]_  & \new_[51573]_ ;
  assign \new_[51584]_  = ~A235 & ~A234;
  assign \new_[51587]_  = ~A265 & ~A236;
  assign \new_[51588]_  = \new_[51587]_  & \new_[51584]_ ;
  assign \new_[51591]_  = ~A268 & ~A266;
  assign \new_[51594]_  = A300 & A299;
  assign \new_[51595]_  = \new_[51594]_  & \new_[51591]_ ;
  assign \new_[51596]_  = \new_[51595]_  & \new_[51588]_ ;
  assign \new_[51600]_  = A166 & ~A167;
  assign \new_[51601]_  = A170 & \new_[51600]_ ;
  assign \new_[51604]_  = A200 & A199;
  assign \new_[51607]_  = ~A202 & ~A201;
  assign \new_[51608]_  = \new_[51607]_  & \new_[51604]_ ;
  assign \new_[51609]_  = \new_[51608]_  & \new_[51601]_ ;
  assign \new_[51612]_  = ~A235 & ~A234;
  assign \new_[51615]_  = ~A265 & ~A236;
  assign \new_[51616]_  = \new_[51615]_  & \new_[51612]_ ;
  assign \new_[51619]_  = ~A268 & ~A266;
  assign \new_[51622]_  = A300 & A298;
  assign \new_[51623]_  = \new_[51622]_  & \new_[51619]_ ;
  assign \new_[51624]_  = \new_[51623]_  & \new_[51616]_ ;
  assign \new_[51628]_  = A166 & ~A167;
  assign \new_[51629]_  = A170 & \new_[51628]_ ;
  assign \new_[51632]_  = A200 & A199;
  assign \new_[51635]_  = ~A202 & ~A201;
  assign \new_[51636]_  = \new_[51635]_  & \new_[51632]_ ;
  assign \new_[51637]_  = \new_[51636]_  & \new_[51629]_ ;
  assign \new_[51640]_  = A233 & A232;
  assign \new_[51643]_  = ~A235 & ~A234;
  assign \new_[51644]_  = \new_[51643]_  & \new_[51640]_ ;
  assign \new_[51647]_  = ~A268 & ~A267;
  assign \new_[51650]_  = A301 & ~A269;
  assign \new_[51651]_  = \new_[51650]_  & \new_[51647]_ ;
  assign \new_[51652]_  = \new_[51651]_  & \new_[51644]_ ;
  assign \new_[51656]_  = A166 & ~A167;
  assign \new_[51657]_  = A170 & \new_[51656]_ ;
  assign \new_[51660]_  = A200 & A199;
  assign \new_[51663]_  = ~A202 & ~A201;
  assign \new_[51664]_  = \new_[51663]_  & \new_[51660]_ ;
  assign \new_[51665]_  = \new_[51664]_  & \new_[51657]_ ;
  assign \new_[51668]_  = A233 & A232;
  assign \new_[51671]_  = ~A235 & ~A234;
  assign \new_[51672]_  = \new_[51671]_  & \new_[51668]_ ;
  assign \new_[51675]_  = ~A266 & ~A265;
  assign \new_[51678]_  = A301 & ~A268;
  assign \new_[51679]_  = \new_[51678]_  & \new_[51675]_ ;
  assign \new_[51680]_  = \new_[51679]_  & \new_[51672]_ ;
  assign \new_[51684]_  = A166 & ~A167;
  assign \new_[51685]_  = A170 & \new_[51684]_ ;
  assign \new_[51688]_  = A200 & A199;
  assign \new_[51691]_  = ~A202 & ~A201;
  assign \new_[51692]_  = \new_[51691]_  & \new_[51688]_ ;
  assign \new_[51693]_  = \new_[51692]_  & \new_[51685]_ ;
  assign \new_[51696]_  = ~A233 & ~A232;
  assign \new_[51699]_  = ~A267 & ~A235;
  assign \new_[51700]_  = \new_[51699]_  & \new_[51696]_ ;
  assign \new_[51703]_  = ~A269 & ~A268;
  assign \new_[51706]_  = A300 & A299;
  assign \new_[51707]_  = \new_[51706]_  & \new_[51703]_ ;
  assign \new_[51708]_  = \new_[51707]_  & \new_[51700]_ ;
  assign \new_[51712]_  = A166 & ~A167;
  assign \new_[51713]_  = A170 & \new_[51712]_ ;
  assign \new_[51716]_  = A200 & A199;
  assign \new_[51719]_  = ~A202 & ~A201;
  assign \new_[51720]_  = \new_[51719]_  & \new_[51716]_ ;
  assign \new_[51721]_  = \new_[51720]_  & \new_[51713]_ ;
  assign \new_[51724]_  = ~A233 & ~A232;
  assign \new_[51727]_  = ~A267 & ~A235;
  assign \new_[51728]_  = \new_[51727]_  & \new_[51724]_ ;
  assign \new_[51731]_  = ~A269 & ~A268;
  assign \new_[51734]_  = A300 & A298;
  assign \new_[51735]_  = \new_[51734]_  & \new_[51731]_ ;
  assign \new_[51736]_  = \new_[51735]_  & \new_[51728]_ ;
  assign \new_[51740]_  = A166 & ~A167;
  assign \new_[51741]_  = A170 & \new_[51740]_ ;
  assign \new_[51744]_  = A200 & A199;
  assign \new_[51747]_  = ~A202 & ~A201;
  assign \new_[51748]_  = \new_[51747]_  & \new_[51744]_ ;
  assign \new_[51749]_  = \new_[51748]_  & \new_[51741]_ ;
  assign \new_[51752]_  = ~A233 & ~A232;
  assign \new_[51755]_  = A265 & ~A235;
  assign \new_[51756]_  = \new_[51755]_  & \new_[51752]_ ;
  assign \new_[51759]_  = ~A267 & A266;
  assign \new_[51762]_  = A301 & ~A268;
  assign \new_[51763]_  = \new_[51762]_  & \new_[51759]_ ;
  assign \new_[51764]_  = \new_[51763]_  & \new_[51756]_ ;
  assign \new_[51768]_  = A166 & ~A167;
  assign \new_[51769]_  = A170 & \new_[51768]_ ;
  assign \new_[51772]_  = A200 & A199;
  assign \new_[51775]_  = ~A202 & ~A201;
  assign \new_[51776]_  = \new_[51775]_  & \new_[51772]_ ;
  assign \new_[51777]_  = \new_[51776]_  & \new_[51769]_ ;
  assign \new_[51780]_  = ~A233 & ~A232;
  assign \new_[51783]_  = ~A265 & ~A235;
  assign \new_[51784]_  = \new_[51783]_  & \new_[51780]_ ;
  assign \new_[51787]_  = ~A268 & ~A266;
  assign \new_[51790]_  = A300 & A299;
  assign \new_[51791]_  = \new_[51790]_  & \new_[51787]_ ;
  assign \new_[51792]_  = \new_[51791]_  & \new_[51784]_ ;
  assign \new_[51796]_  = A166 & ~A167;
  assign \new_[51797]_  = A170 & \new_[51796]_ ;
  assign \new_[51800]_  = A200 & A199;
  assign \new_[51803]_  = ~A202 & ~A201;
  assign \new_[51804]_  = \new_[51803]_  & \new_[51800]_ ;
  assign \new_[51805]_  = \new_[51804]_  & \new_[51797]_ ;
  assign \new_[51808]_  = ~A233 & ~A232;
  assign \new_[51811]_  = ~A265 & ~A235;
  assign \new_[51812]_  = \new_[51811]_  & \new_[51808]_ ;
  assign \new_[51815]_  = ~A268 & ~A266;
  assign \new_[51818]_  = A300 & A298;
  assign \new_[51819]_  = \new_[51818]_  & \new_[51815]_ ;
  assign \new_[51820]_  = \new_[51819]_  & \new_[51812]_ ;
  assign \new_[51824]_  = A166 & ~A167;
  assign \new_[51825]_  = A170 & \new_[51824]_ ;
  assign \new_[51828]_  = ~A200 & ~A199;
  assign \new_[51831]_  = ~A234 & ~A202;
  assign \new_[51832]_  = \new_[51831]_  & \new_[51828]_ ;
  assign \new_[51833]_  = \new_[51832]_  & \new_[51825]_ ;
  assign \new_[51836]_  = ~A236 & ~A235;
  assign \new_[51839]_  = ~A268 & ~A267;
  assign \new_[51840]_  = \new_[51839]_  & \new_[51836]_ ;
  assign \new_[51843]_  = A298 & ~A269;
  assign \new_[51846]_  = A302 & ~A299;
  assign \new_[51847]_  = \new_[51846]_  & \new_[51843]_ ;
  assign \new_[51848]_  = \new_[51847]_  & \new_[51840]_ ;
  assign \new_[51852]_  = A166 & ~A167;
  assign \new_[51853]_  = A170 & \new_[51852]_ ;
  assign \new_[51856]_  = ~A200 & ~A199;
  assign \new_[51859]_  = ~A234 & ~A202;
  assign \new_[51860]_  = \new_[51859]_  & \new_[51856]_ ;
  assign \new_[51861]_  = \new_[51860]_  & \new_[51853]_ ;
  assign \new_[51864]_  = ~A236 & ~A235;
  assign \new_[51867]_  = ~A268 & ~A267;
  assign \new_[51868]_  = \new_[51867]_  & \new_[51864]_ ;
  assign \new_[51871]_  = ~A298 & ~A269;
  assign \new_[51874]_  = A302 & A299;
  assign \new_[51875]_  = \new_[51874]_  & \new_[51871]_ ;
  assign \new_[51876]_  = \new_[51875]_  & \new_[51868]_ ;
  assign \new_[51880]_  = A166 & ~A167;
  assign \new_[51881]_  = A170 & \new_[51880]_ ;
  assign \new_[51884]_  = ~A200 & ~A199;
  assign \new_[51887]_  = ~A234 & ~A202;
  assign \new_[51888]_  = \new_[51887]_  & \new_[51884]_ ;
  assign \new_[51889]_  = \new_[51888]_  & \new_[51881]_ ;
  assign \new_[51892]_  = ~A236 & ~A235;
  assign \new_[51895]_  = A266 & A265;
  assign \new_[51896]_  = \new_[51895]_  & \new_[51892]_ ;
  assign \new_[51899]_  = ~A268 & ~A267;
  assign \new_[51902]_  = A300 & A299;
  assign \new_[51903]_  = \new_[51902]_  & \new_[51899]_ ;
  assign \new_[51904]_  = \new_[51903]_  & \new_[51896]_ ;
  assign \new_[51908]_  = A166 & ~A167;
  assign \new_[51909]_  = A170 & \new_[51908]_ ;
  assign \new_[51912]_  = ~A200 & ~A199;
  assign \new_[51915]_  = ~A234 & ~A202;
  assign \new_[51916]_  = \new_[51915]_  & \new_[51912]_ ;
  assign \new_[51917]_  = \new_[51916]_  & \new_[51909]_ ;
  assign \new_[51920]_  = ~A236 & ~A235;
  assign \new_[51923]_  = A266 & A265;
  assign \new_[51924]_  = \new_[51923]_  & \new_[51920]_ ;
  assign \new_[51927]_  = ~A268 & ~A267;
  assign \new_[51930]_  = A300 & A298;
  assign \new_[51931]_  = \new_[51930]_  & \new_[51927]_ ;
  assign \new_[51932]_  = \new_[51931]_  & \new_[51924]_ ;
  assign \new_[51936]_  = A166 & ~A167;
  assign \new_[51937]_  = A170 & \new_[51936]_ ;
  assign \new_[51940]_  = ~A200 & ~A199;
  assign \new_[51943]_  = ~A234 & ~A202;
  assign \new_[51944]_  = \new_[51943]_  & \new_[51940]_ ;
  assign \new_[51945]_  = \new_[51944]_  & \new_[51937]_ ;
  assign \new_[51948]_  = ~A236 & ~A235;
  assign \new_[51951]_  = ~A266 & ~A265;
  assign \new_[51952]_  = \new_[51951]_  & \new_[51948]_ ;
  assign \new_[51955]_  = A298 & ~A268;
  assign \new_[51958]_  = A302 & ~A299;
  assign \new_[51959]_  = \new_[51958]_  & \new_[51955]_ ;
  assign \new_[51960]_  = \new_[51959]_  & \new_[51952]_ ;
  assign \new_[51964]_  = A166 & ~A167;
  assign \new_[51965]_  = A170 & \new_[51964]_ ;
  assign \new_[51968]_  = ~A200 & ~A199;
  assign \new_[51971]_  = ~A234 & ~A202;
  assign \new_[51972]_  = \new_[51971]_  & \new_[51968]_ ;
  assign \new_[51973]_  = \new_[51972]_  & \new_[51965]_ ;
  assign \new_[51976]_  = ~A236 & ~A235;
  assign \new_[51979]_  = ~A266 & ~A265;
  assign \new_[51980]_  = \new_[51979]_  & \new_[51976]_ ;
  assign \new_[51983]_  = ~A298 & ~A268;
  assign \new_[51986]_  = A302 & A299;
  assign \new_[51987]_  = \new_[51986]_  & \new_[51983]_ ;
  assign \new_[51988]_  = \new_[51987]_  & \new_[51980]_ ;
  assign \new_[51992]_  = A166 & ~A167;
  assign \new_[51993]_  = A170 & \new_[51992]_ ;
  assign \new_[51996]_  = ~A200 & ~A199;
  assign \new_[51999]_  = A232 & ~A202;
  assign \new_[52000]_  = \new_[51999]_  & \new_[51996]_ ;
  assign \new_[52001]_  = \new_[52000]_  & \new_[51993]_ ;
  assign \new_[52004]_  = ~A234 & A233;
  assign \new_[52007]_  = ~A267 & ~A235;
  assign \new_[52008]_  = \new_[52007]_  & \new_[52004]_ ;
  assign \new_[52011]_  = ~A269 & ~A268;
  assign \new_[52014]_  = A300 & A299;
  assign \new_[52015]_  = \new_[52014]_  & \new_[52011]_ ;
  assign \new_[52016]_  = \new_[52015]_  & \new_[52008]_ ;
  assign \new_[52020]_  = A166 & ~A167;
  assign \new_[52021]_  = A170 & \new_[52020]_ ;
  assign \new_[52024]_  = ~A200 & ~A199;
  assign \new_[52027]_  = A232 & ~A202;
  assign \new_[52028]_  = \new_[52027]_  & \new_[52024]_ ;
  assign \new_[52029]_  = \new_[52028]_  & \new_[52021]_ ;
  assign \new_[52032]_  = ~A234 & A233;
  assign \new_[52035]_  = ~A267 & ~A235;
  assign \new_[52036]_  = \new_[52035]_  & \new_[52032]_ ;
  assign \new_[52039]_  = ~A269 & ~A268;
  assign \new_[52042]_  = A300 & A298;
  assign \new_[52043]_  = \new_[52042]_  & \new_[52039]_ ;
  assign \new_[52044]_  = \new_[52043]_  & \new_[52036]_ ;
  assign \new_[52048]_  = A166 & ~A167;
  assign \new_[52049]_  = A170 & \new_[52048]_ ;
  assign \new_[52052]_  = ~A200 & ~A199;
  assign \new_[52055]_  = A232 & ~A202;
  assign \new_[52056]_  = \new_[52055]_  & \new_[52052]_ ;
  assign \new_[52057]_  = \new_[52056]_  & \new_[52049]_ ;
  assign \new_[52060]_  = ~A234 & A233;
  assign \new_[52063]_  = A265 & ~A235;
  assign \new_[52064]_  = \new_[52063]_  & \new_[52060]_ ;
  assign \new_[52067]_  = ~A267 & A266;
  assign \new_[52070]_  = A301 & ~A268;
  assign \new_[52071]_  = \new_[52070]_  & \new_[52067]_ ;
  assign \new_[52072]_  = \new_[52071]_  & \new_[52064]_ ;
  assign \new_[52076]_  = A166 & ~A167;
  assign \new_[52077]_  = A170 & \new_[52076]_ ;
  assign \new_[52080]_  = ~A200 & ~A199;
  assign \new_[52083]_  = A232 & ~A202;
  assign \new_[52084]_  = \new_[52083]_  & \new_[52080]_ ;
  assign \new_[52085]_  = \new_[52084]_  & \new_[52077]_ ;
  assign \new_[52088]_  = ~A234 & A233;
  assign \new_[52091]_  = ~A265 & ~A235;
  assign \new_[52092]_  = \new_[52091]_  & \new_[52088]_ ;
  assign \new_[52095]_  = ~A268 & ~A266;
  assign \new_[52098]_  = A300 & A299;
  assign \new_[52099]_  = \new_[52098]_  & \new_[52095]_ ;
  assign \new_[52100]_  = \new_[52099]_  & \new_[52092]_ ;
  assign \new_[52104]_  = A166 & ~A167;
  assign \new_[52105]_  = A170 & \new_[52104]_ ;
  assign \new_[52108]_  = ~A200 & ~A199;
  assign \new_[52111]_  = A232 & ~A202;
  assign \new_[52112]_  = \new_[52111]_  & \new_[52108]_ ;
  assign \new_[52113]_  = \new_[52112]_  & \new_[52105]_ ;
  assign \new_[52116]_  = ~A234 & A233;
  assign \new_[52119]_  = ~A265 & ~A235;
  assign \new_[52120]_  = \new_[52119]_  & \new_[52116]_ ;
  assign \new_[52123]_  = ~A268 & ~A266;
  assign \new_[52126]_  = A300 & A298;
  assign \new_[52127]_  = \new_[52126]_  & \new_[52123]_ ;
  assign \new_[52128]_  = \new_[52127]_  & \new_[52120]_ ;
  assign \new_[52132]_  = A166 & ~A167;
  assign \new_[52133]_  = A170 & \new_[52132]_ ;
  assign \new_[52136]_  = ~A200 & ~A199;
  assign \new_[52139]_  = ~A232 & ~A202;
  assign \new_[52140]_  = \new_[52139]_  & \new_[52136]_ ;
  assign \new_[52141]_  = \new_[52140]_  & \new_[52133]_ ;
  assign \new_[52144]_  = ~A235 & ~A233;
  assign \new_[52147]_  = ~A268 & ~A267;
  assign \new_[52148]_  = \new_[52147]_  & \new_[52144]_ ;
  assign \new_[52151]_  = A298 & ~A269;
  assign \new_[52154]_  = A302 & ~A299;
  assign \new_[52155]_  = \new_[52154]_  & \new_[52151]_ ;
  assign \new_[52156]_  = \new_[52155]_  & \new_[52148]_ ;
  assign \new_[52160]_  = A166 & ~A167;
  assign \new_[52161]_  = A170 & \new_[52160]_ ;
  assign \new_[52164]_  = ~A200 & ~A199;
  assign \new_[52167]_  = ~A232 & ~A202;
  assign \new_[52168]_  = \new_[52167]_  & \new_[52164]_ ;
  assign \new_[52169]_  = \new_[52168]_  & \new_[52161]_ ;
  assign \new_[52172]_  = ~A235 & ~A233;
  assign \new_[52175]_  = ~A268 & ~A267;
  assign \new_[52176]_  = \new_[52175]_  & \new_[52172]_ ;
  assign \new_[52179]_  = ~A298 & ~A269;
  assign \new_[52182]_  = A302 & A299;
  assign \new_[52183]_  = \new_[52182]_  & \new_[52179]_ ;
  assign \new_[52184]_  = \new_[52183]_  & \new_[52176]_ ;
  assign \new_[52188]_  = A166 & ~A167;
  assign \new_[52189]_  = A170 & \new_[52188]_ ;
  assign \new_[52192]_  = ~A200 & ~A199;
  assign \new_[52195]_  = ~A232 & ~A202;
  assign \new_[52196]_  = \new_[52195]_  & \new_[52192]_ ;
  assign \new_[52197]_  = \new_[52196]_  & \new_[52189]_ ;
  assign \new_[52200]_  = ~A235 & ~A233;
  assign \new_[52203]_  = A266 & A265;
  assign \new_[52204]_  = \new_[52203]_  & \new_[52200]_ ;
  assign \new_[52207]_  = ~A268 & ~A267;
  assign \new_[52210]_  = A300 & A299;
  assign \new_[52211]_  = \new_[52210]_  & \new_[52207]_ ;
  assign \new_[52212]_  = \new_[52211]_  & \new_[52204]_ ;
  assign \new_[52216]_  = A166 & ~A167;
  assign \new_[52217]_  = A170 & \new_[52216]_ ;
  assign \new_[52220]_  = ~A200 & ~A199;
  assign \new_[52223]_  = ~A232 & ~A202;
  assign \new_[52224]_  = \new_[52223]_  & \new_[52220]_ ;
  assign \new_[52225]_  = \new_[52224]_  & \new_[52217]_ ;
  assign \new_[52228]_  = ~A235 & ~A233;
  assign \new_[52231]_  = A266 & A265;
  assign \new_[52232]_  = \new_[52231]_  & \new_[52228]_ ;
  assign \new_[52235]_  = ~A268 & ~A267;
  assign \new_[52238]_  = A300 & A298;
  assign \new_[52239]_  = \new_[52238]_  & \new_[52235]_ ;
  assign \new_[52240]_  = \new_[52239]_  & \new_[52232]_ ;
  assign \new_[52244]_  = A166 & ~A167;
  assign \new_[52245]_  = A170 & \new_[52244]_ ;
  assign \new_[52248]_  = ~A200 & ~A199;
  assign \new_[52251]_  = ~A232 & ~A202;
  assign \new_[52252]_  = \new_[52251]_  & \new_[52248]_ ;
  assign \new_[52253]_  = \new_[52252]_  & \new_[52245]_ ;
  assign \new_[52256]_  = ~A235 & ~A233;
  assign \new_[52259]_  = ~A266 & ~A265;
  assign \new_[52260]_  = \new_[52259]_  & \new_[52256]_ ;
  assign \new_[52263]_  = A298 & ~A268;
  assign \new_[52266]_  = A302 & ~A299;
  assign \new_[52267]_  = \new_[52266]_  & \new_[52263]_ ;
  assign \new_[52268]_  = \new_[52267]_  & \new_[52260]_ ;
  assign \new_[52272]_  = A166 & ~A167;
  assign \new_[52273]_  = A170 & \new_[52272]_ ;
  assign \new_[52276]_  = ~A200 & ~A199;
  assign \new_[52279]_  = ~A232 & ~A202;
  assign \new_[52280]_  = \new_[52279]_  & \new_[52276]_ ;
  assign \new_[52281]_  = \new_[52280]_  & \new_[52273]_ ;
  assign \new_[52284]_  = ~A235 & ~A233;
  assign \new_[52287]_  = ~A266 & ~A265;
  assign \new_[52288]_  = \new_[52287]_  & \new_[52284]_ ;
  assign \new_[52291]_  = ~A298 & ~A268;
  assign \new_[52294]_  = A302 & A299;
  assign \new_[52295]_  = \new_[52294]_  & \new_[52291]_ ;
  assign \new_[52296]_  = \new_[52295]_  & \new_[52288]_ ;
  assign \new_[52300]_  = ~A202 & ~A201;
  assign \new_[52301]_  = A169 & \new_[52300]_ ;
  assign \new_[52304]_  = A232 & ~A203;
  assign \new_[52307]_  = ~A234 & A233;
  assign \new_[52308]_  = \new_[52307]_  & \new_[52304]_ ;
  assign \new_[52309]_  = \new_[52308]_  & \new_[52301]_ ;
  assign \new_[52312]_  = A265 & ~A235;
  assign \new_[52315]_  = ~A267 & A266;
  assign \new_[52316]_  = \new_[52315]_  & \new_[52312]_ ;
  assign \new_[52319]_  = A298 & ~A268;
  assign \new_[52322]_  = A302 & ~A299;
  assign \new_[52323]_  = \new_[52322]_  & \new_[52319]_ ;
  assign \new_[52324]_  = \new_[52323]_  & \new_[52316]_ ;
  assign \new_[52328]_  = ~A202 & ~A201;
  assign \new_[52329]_  = A169 & \new_[52328]_ ;
  assign \new_[52332]_  = A232 & ~A203;
  assign \new_[52335]_  = ~A234 & A233;
  assign \new_[52336]_  = \new_[52335]_  & \new_[52332]_ ;
  assign \new_[52337]_  = \new_[52336]_  & \new_[52329]_ ;
  assign \new_[52340]_  = A265 & ~A235;
  assign \new_[52343]_  = ~A267 & A266;
  assign \new_[52344]_  = \new_[52343]_  & \new_[52340]_ ;
  assign \new_[52347]_  = ~A298 & ~A268;
  assign \new_[52350]_  = A302 & A299;
  assign \new_[52351]_  = \new_[52350]_  & \new_[52347]_ ;
  assign \new_[52352]_  = \new_[52351]_  & \new_[52344]_ ;
  assign \new_[52356]_  = A200 & A199;
  assign \new_[52357]_  = A169 & \new_[52356]_ ;
  assign \new_[52360]_  = ~A202 & ~A201;
  assign \new_[52363]_  = ~A235 & ~A234;
  assign \new_[52364]_  = \new_[52363]_  & \new_[52360]_ ;
  assign \new_[52365]_  = \new_[52364]_  & \new_[52357]_ ;
  assign \new_[52368]_  = A265 & ~A236;
  assign \new_[52371]_  = ~A267 & A266;
  assign \new_[52372]_  = \new_[52371]_  & \new_[52368]_ ;
  assign \new_[52375]_  = A298 & ~A268;
  assign \new_[52378]_  = A302 & ~A299;
  assign \new_[52379]_  = \new_[52378]_  & \new_[52375]_ ;
  assign \new_[52380]_  = \new_[52379]_  & \new_[52372]_ ;
  assign \new_[52384]_  = A200 & A199;
  assign \new_[52385]_  = A169 & \new_[52384]_ ;
  assign \new_[52388]_  = ~A202 & ~A201;
  assign \new_[52391]_  = ~A235 & ~A234;
  assign \new_[52392]_  = \new_[52391]_  & \new_[52388]_ ;
  assign \new_[52393]_  = \new_[52392]_  & \new_[52385]_ ;
  assign \new_[52396]_  = A265 & ~A236;
  assign \new_[52399]_  = ~A267 & A266;
  assign \new_[52400]_  = \new_[52399]_  & \new_[52396]_ ;
  assign \new_[52403]_  = ~A298 & ~A268;
  assign \new_[52406]_  = A302 & A299;
  assign \new_[52407]_  = \new_[52406]_  & \new_[52403]_ ;
  assign \new_[52408]_  = \new_[52407]_  & \new_[52400]_ ;
  assign \new_[52412]_  = A200 & A199;
  assign \new_[52413]_  = A169 & \new_[52412]_ ;
  assign \new_[52416]_  = ~A202 & ~A201;
  assign \new_[52419]_  = A233 & A232;
  assign \new_[52420]_  = \new_[52419]_  & \new_[52416]_ ;
  assign \new_[52421]_  = \new_[52420]_  & \new_[52413]_ ;
  assign \new_[52424]_  = ~A235 & ~A234;
  assign \new_[52427]_  = ~A268 & ~A267;
  assign \new_[52428]_  = \new_[52427]_  & \new_[52424]_ ;
  assign \new_[52431]_  = A298 & ~A269;
  assign \new_[52434]_  = A302 & ~A299;
  assign \new_[52435]_  = \new_[52434]_  & \new_[52431]_ ;
  assign \new_[52436]_  = \new_[52435]_  & \new_[52428]_ ;
  assign \new_[52440]_  = A200 & A199;
  assign \new_[52441]_  = A169 & \new_[52440]_ ;
  assign \new_[52444]_  = ~A202 & ~A201;
  assign \new_[52447]_  = A233 & A232;
  assign \new_[52448]_  = \new_[52447]_  & \new_[52444]_ ;
  assign \new_[52449]_  = \new_[52448]_  & \new_[52441]_ ;
  assign \new_[52452]_  = ~A235 & ~A234;
  assign \new_[52455]_  = ~A268 & ~A267;
  assign \new_[52456]_  = \new_[52455]_  & \new_[52452]_ ;
  assign \new_[52459]_  = ~A298 & ~A269;
  assign \new_[52462]_  = A302 & A299;
  assign \new_[52463]_  = \new_[52462]_  & \new_[52459]_ ;
  assign \new_[52464]_  = \new_[52463]_  & \new_[52456]_ ;
  assign \new_[52468]_  = A200 & A199;
  assign \new_[52469]_  = A169 & \new_[52468]_ ;
  assign \new_[52472]_  = ~A202 & ~A201;
  assign \new_[52475]_  = A233 & A232;
  assign \new_[52476]_  = \new_[52475]_  & \new_[52472]_ ;
  assign \new_[52477]_  = \new_[52476]_  & \new_[52469]_ ;
  assign \new_[52480]_  = ~A235 & ~A234;
  assign \new_[52483]_  = A266 & A265;
  assign \new_[52484]_  = \new_[52483]_  & \new_[52480]_ ;
  assign \new_[52487]_  = ~A268 & ~A267;
  assign \new_[52490]_  = A300 & A299;
  assign \new_[52491]_  = \new_[52490]_  & \new_[52487]_ ;
  assign \new_[52492]_  = \new_[52491]_  & \new_[52484]_ ;
  assign \new_[52496]_  = A200 & A199;
  assign \new_[52497]_  = A169 & \new_[52496]_ ;
  assign \new_[52500]_  = ~A202 & ~A201;
  assign \new_[52503]_  = A233 & A232;
  assign \new_[52504]_  = \new_[52503]_  & \new_[52500]_ ;
  assign \new_[52505]_  = \new_[52504]_  & \new_[52497]_ ;
  assign \new_[52508]_  = ~A235 & ~A234;
  assign \new_[52511]_  = A266 & A265;
  assign \new_[52512]_  = \new_[52511]_  & \new_[52508]_ ;
  assign \new_[52515]_  = ~A268 & ~A267;
  assign \new_[52518]_  = A300 & A298;
  assign \new_[52519]_  = \new_[52518]_  & \new_[52515]_ ;
  assign \new_[52520]_  = \new_[52519]_  & \new_[52512]_ ;
  assign \new_[52524]_  = A200 & A199;
  assign \new_[52525]_  = A169 & \new_[52524]_ ;
  assign \new_[52528]_  = ~A202 & ~A201;
  assign \new_[52531]_  = A233 & A232;
  assign \new_[52532]_  = \new_[52531]_  & \new_[52528]_ ;
  assign \new_[52533]_  = \new_[52532]_  & \new_[52525]_ ;
  assign \new_[52536]_  = ~A235 & ~A234;
  assign \new_[52539]_  = ~A266 & ~A265;
  assign \new_[52540]_  = \new_[52539]_  & \new_[52536]_ ;
  assign \new_[52543]_  = A298 & ~A268;
  assign \new_[52546]_  = A302 & ~A299;
  assign \new_[52547]_  = \new_[52546]_  & \new_[52543]_ ;
  assign \new_[52548]_  = \new_[52547]_  & \new_[52540]_ ;
  assign \new_[52552]_  = A200 & A199;
  assign \new_[52553]_  = A169 & \new_[52552]_ ;
  assign \new_[52556]_  = ~A202 & ~A201;
  assign \new_[52559]_  = A233 & A232;
  assign \new_[52560]_  = \new_[52559]_  & \new_[52556]_ ;
  assign \new_[52561]_  = \new_[52560]_  & \new_[52553]_ ;
  assign \new_[52564]_  = ~A235 & ~A234;
  assign \new_[52567]_  = ~A266 & ~A265;
  assign \new_[52568]_  = \new_[52567]_  & \new_[52564]_ ;
  assign \new_[52571]_  = ~A298 & ~A268;
  assign \new_[52574]_  = A302 & A299;
  assign \new_[52575]_  = \new_[52574]_  & \new_[52571]_ ;
  assign \new_[52576]_  = \new_[52575]_  & \new_[52568]_ ;
  assign \new_[52580]_  = A200 & A199;
  assign \new_[52581]_  = A169 & \new_[52580]_ ;
  assign \new_[52584]_  = ~A202 & ~A201;
  assign \new_[52587]_  = ~A233 & ~A232;
  assign \new_[52588]_  = \new_[52587]_  & \new_[52584]_ ;
  assign \new_[52589]_  = \new_[52588]_  & \new_[52581]_ ;
  assign \new_[52592]_  = A265 & ~A235;
  assign \new_[52595]_  = ~A267 & A266;
  assign \new_[52596]_  = \new_[52595]_  & \new_[52592]_ ;
  assign \new_[52599]_  = A298 & ~A268;
  assign \new_[52602]_  = A302 & ~A299;
  assign \new_[52603]_  = \new_[52602]_  & \new_[52599]_ ;
  assign \new_[52604]_  = \new_[52603]_  & \new_[52596]_ ;
  assign \new_[52608]_  = A200 & A199;
  assign \new_[52609]_  = A169 & \new_[52608]_ ;
  assign \new_[52612]_  = ~A202 & ~A201;
  assign \new_[52615]_  = ~A233 & ~A232;
  assign \new_[52616]_  = \new_[52615]_  & \new_[52612]_ ;
  assign \new_[52617]_  = \new_[52616]_  & \new_[52609]_ ;
  assign \new_[52620]_  = A265 & ~A235;
  assign \new_[52623]_  = ~A267 & A266;
  assign \new_[52624]_  = \new_[52623]_  & \new_[52620]_ ;
  assign \new_[52627]_  = ~A298 & ~A268;
  assign \new_[52630]_  = A302 & A299;
  assign \new_[52631]_  = \new_[52630]_  & \new_[52627]_ ;
  assign \new_[52632]_  = \new_[52631]_  & \new_[52624]_ ;
  assign \new_[52636]_  = ~A200 & ~A199;
  assign \new_[52637]_  = A169 & \new_[52636]_ ;
  assign \new_[52640]_  = A232 & ~A202;
  assign \new_[52643]_  = ~A234 & A233;
  assign \new_[52644]_  = \new_[52643]_  & \new_[52640]_ ;
  assign \new_[52645]_  = \new_[52644]_  & \new_[52637]_ ;
  assign \new_[52648]_  = A265 & ~A235;
  assign \new_[52651]_  = ~A267 & A266;
  assign \new_[52652]_  = \new_[52651]_  & \new_[52648]_ ;
  assign \new_[52655]_  = A298 & ~A268;
  assign \new_[52658]_  = A302 & ~A299;
  assign \new_[52659]_  = \new_[52658]_  & \new_[52655]_ ;
  assign \new_[52660]_  = \new_[52659]_  & \new_[52652]_ ;
  assign \new_[52664]_  = ~A200 & ~A199;
  assign \new_[52665]_  = A169 & \new_[52664]_ ;
  assign \new_[52668]_  = A232 & ~A202;
  assign \new_[52671]_  = ~A234 & A233;
  assign \new_[52672]_  = \new_[52671]_  & \new_[52668]_ ;
  assign \new_[52673]_  = \new_[52672]_  & \new_[52665]_ ;
  assign \new_[52676]_  = A265 & ~A235;
  assign \new_[52679]_  = ~A267 & A266;
  assign \new_[52680]_  = \new_[52679]_  & \new_[52676]_ ;
  assign \new_[52683]_  = ~A298 & ~A268;
  assign \new_[52686]_  = A302 & A299;
  assign \new_[52687]_  = \new_[52686]_  & \new_[52683]_ ;
  assign \new_[52688]_  = \new_[52687]_  & \new_[52680]_ ;
  assign \new_[52692]_  = ~A166 & ~A167;
  assign \new_[52693]_  = ~A169 & \new_[52692]_ ;
  assign \new_[52696]_  = A232 & A202;
  assign \new_[52699]_  = ~A234 & A233;
  assign \new_[52700]_  = \new_[52699]_  & \new_[52696]_ ;
  assign \new_[52701]_  = \new_[52700]_  & \new_[52693]_ ;
  assign \new_[52704]_  = A265 & ~A235;
  assign \new_[52707]_  = ~A267 & A266;
  assign \new_[52708]_  = \new_[52707]_  & \new_[52704]_ ;
  assign \new_[52711]_  = A298 & ~A268;
  assign \new_[52714]_  = A302 & ~A299;
  assign \new_[52715]_  = \new_[52714]_  & \new_[52711]_ ;
  assign \new_[52716]_  = \new_[52715]_  & \new_[52708]_ ;
  assign \new_[52720]_  = ~A166 & ~A167;
  assign \new_[52721]_  = ~A169 & \new_[52720]_ ;
  assign \new_[52724]_  = A232 & A202;
  assign \new_[52727]_  = ~A234 & A233;
  assign \new_[52728]_  = \new_[52727]_  & \new_[52724]_ ;
  assign \new_[52729]_  = \new_[52728]_  & \new_[52721]_ ;
  assign \new_[52732]_  = A265 & ~A235;
  assign \new_[52735]_  = ~A267 & A266;
  assign \new_[52736]_  = \new_[52735]_  & \new_[52732]_ ;
  assign \new_[52739]_  = ~A298 & ~A268;
  assign \new_[52742]_  = A302 & A299;
  assign \new_[52743]_  = \new_[52742]_  & \new_[52739]_ ;
  assign \new_[52744]_  = \new_[52743]_  & \new_[52736]_ ;
  assign \new_[52748]_  = ~A166 & ~A167;
  assign \new_[52749]_  = ~A169 & \new_[52748]_ ;
  assign \new_[52752]_  = A201 & A199;
  assign \new_[52755]_  = ~A235 & ~A234;
  assign \new_[52756]_  = \new_[52755]_  & \new_[52752]_ ;
  assign \new_[52757]_  = \new_[52756]_  & \new_[52749]_ ;
  assign \new_[52760]_  = A265 & ~A236;
  assign \new_[52763]_  = ~A267 & A266;
  assign \new_[52764]_  = \new_[52763]_  & \new_[52760]_ ;
  assign \new_[52767]_  = A298 & ~A268;
  assign \new_[52770]_  = A302 & ~A299;
  assign \new_[52771]_  = \new_[52770]_  & \new_[52767]_ ;
  assign \new_[52772]_  = \new_[52771]_  & \new_[52764]_ ;
  assign \new_[52776]_  = ~A166 & ~A167;
  assign \new_[52777]_  = ~A169 & \new_[52776]_ ;
  assign \new_[52780]_  = A201 & A199;
  assign \new_[52783]_  = ~A235 & ~A234;
  assign \new_[52784]_  = \new_[52783]_  & \new_[52780]_ ;
  assign \new_[52785]_  = \new_[52784]_  & \new_[52777]_ ;
  assign \new_[52788]_  = A265 & ~A236;
  assign \new_[52791]_  = ~A267 & A266;
  assign \new_[52792]_  = \new_[52791]_  & \new_[52788]_ ;
  assign \new_[52795]_  = ~A298 & ~A268;
  assign \new_[52798]_  = A302 & A299;
  assign \new_[52799]_  = \new_[52798]_  & \new_[52795]_ ;
  assign \new_[52800]_  = \new_[52799]_  & \new_[52792]_ ;
  assign \new_[52804]_  = ~A166 & ~A167;
  assign \new_[52805]_  = ~A169 & \new_[52804]_ ;
  assign \new_[52808]_  = A201 & A199;
  assign \new_[52811]_  = A233 & A232;
  assign \new_[52812]_  = \new_[52811]_  & \new_[52808]_ ;
  assign \new_[52813]_  = \new_[52812]_  & \new_[52805]_ ;
  assign \new_[52816]_  = ~A235 & ~A234;
  assign \new_[52819]_  = ~A268 & ~A267;
  assign \new_[52820]_  = \new_[52819]_  & \new_[52816]_ ;
  assign \new_[52823]_  = A298 & ~A269;
  assign \new_[52826]_  = A302 & ~A299;
  assign \new_[52827]_  = \new_[52826]_  & \new_[52823]_ ;
  assign \new_[52828]_  = \new_[52827]_  & \new_[52820]_ ;
  assign \new_[52832]_  = ~A166 & ~A167;
  assign \new_[52833]_  = ~A169 & \new_[52832]_ ;
  assign \new_[52836]_  = A201 & A199;
  assign \new_[52839]_  = A233 & A232;
  assign \new_[52840]_  = \new_[52839]_  & \new_[52836]_ ;
  assign \new_[52841]_  = \new_[52840]_  & \new_[52833]_ ;
  assign \new_[52844]_  = ~A235 & ~A234;
  assign \new_[52847]_  = ~A268 & ~A267;
  assign \new_[52848]_  = \new_[52847]_  & \new_[52844]_ ;
  assign \new_[52851]_  = ~A298 & ~A269;
  assign \new_[52854]_  = A302 & A299;
  assign \new_[52855]_  = \new_[52854]_  & \new_[52851]_ ;
  assign \new_[52856]_  = \new_[52855]_  & \new_[52848]_ ;
  assign \new_[52860]_  = ~A166 & ~A167;
  assign \new_[52861]_  = ~A169 & \new_[52860]_ ;
  assign \new_[52864]_  = A201 & A199;
  assign \new_[52867]_  = A233 & A232;
  assign \new_[52868]_  = \new_[52867]_  & \new_[52864]_ ;
  assign \new_[52869]_  = \new_[52868]_  & \new_[52861]_ ;
  assign \new_[52872]_  = ~A235 & ~A234;
  assign \new_[52875]_  = A266 & A265;
  assign \new_[52876]_  = \new_[52875]_  & \new_[52872]_ ;
  assign \new_[52879]_  = ~A268 & ~A267;
  assign \new_[52882]_  = A300 & A299;
  assign \new_[52883]_  = \new_[52882]_  & \new_[52879]_ ;
  assign \new_[52884]_  = \new_[52883]_  & \new_[52876]_ ;
  assign \new_[52888]_  = ~A166 & ~A167;
  assign \new_[52889]_  = ~A169 & \new_[52888]_ ;
  assign \new_[52892]_  = A201 & A199;
  assign \new_[52895]_  = A233 & A232;
  assign \new_[52896]_  = \new_[52895]_  & \new_[52892]_ ;
  assign \new_[52897]_  = \new_[52896]_  & \new_[52889]_ ;
  assign \new_[52900]_  = ~A235 & ~A234;
  assign \new_[52903]_  = A266 & A265;
  assign \new_[52904]_  = \new_[52903]_  & \new_[52900]_ ;
  assign \new_[52907]_  = ~A268 & ~A267;
  assign \new_[52910]_  = A300 & A298;
  assign \new_[52911]_  = \new_[52910]_  & \new_[52907]_ ;
  assign \new_[52912]_  = \new_[52911]_  & \new_[52904]_ ;
  assign \new_[52916]_  = ~A166 & ~A167;
  assign \new_[52917]_  = ~A169 & \new_[52916]_ ;
  assign \new_[52920]_  = A201 & A199;
  assign \new_[52923]_  = A233 & A232;
  assign \new_[52924]_  = \new_[52923]_  & \new_[52920]_ ;
  assign \new_[52925]_  = \new_[52924]_  & \new_[52917]_ ;
  assign \new_[52928]_  = ~A235 & ~A234;
  assign \new_[52931]_  = ~A266 & ~A265;
  assign \new_[52932]_  = \new_[52931]_  & \new_[52928]_ ;
  assign \new_[52935]_  = A298 & ~A268;
  assign \new_[52938]_  = A302 & ~A299;
  assign \new_[52939]_  = \new_[52938]_  & \new_[52935]_ ;
  assign \new_[52940]_  = \new_[52939]_  & \new_[52932]_ ;
  assign \new_[52944]_  = ~A166 & ~A167;
  assign \new_[52945]_  = ~A169 & \new_[52944]_ ;
  assign \new_[52948]_  = A201 & A199;
  assign \new_[52951]_  = A233 & A232;
  assign \new_[52952]_  = \new_[52951]_  & \new_[52948]_ ;
  assign \new_[52953]_  = \new_[52952]_  & \new_[52945]_ ;
  assign \new_[52956]_  = ~A235 & ~A234;
  assign \new_[52959]_  = ~A266 & ~A265;
  assign \new_[52960]_  = \new_[52959]_  & \new_[52956]_ ;
  assign \new_[52963]_  = ~A298 & ~A268;
  assign \new_[52966]_  = A302 & A299;
  assign \new_[52967]_  = \new_[52966]_  & \new_[52963]_ ;
  assign \new_[52968]_  = \new_[52967]_  & \new_[52960]_ ;
  assign \new_[52972]_  = ~A166 & ~A167;
  assign \new_[52973]_  = ~A169 & \new_[52972]_ ;
  assign \new_[52976]_  = A201 & A199;
  assign \new_[52979]_  = ~A233 & ~A232;
  assign \new_[52980]_  = \new_[52979]_  & \new_[52976]_ ;
  assign \new_[52981]_  = \new_[52980]_  & \new_[52973]_ ;
  assign \new_[52984]_  = A265 & ~A235;
  assign \new_[52987]_  = ~A267 & A266;
  assign \new_[52988]_  = \new_[52987]_  & \new_[52984]_ ;
  assign \new_[52991]_  = A298 & ~A268;
  assign \new_[52994]_  = A302 & ~A299;
  assign \new_[52995]_  = \new_[52994]_  & \new_[52991]_ ;
  assign \new_[52996]_  = \new_[52995]_  & \new_[52988]_ ;
  assign \new_[53000]_  = ~A166 & ~A167;
  assign \new_[53001]_  = ~A169 & \new_[53000]_ ;
  assign \new_[53004]_  = A201 & A199;
  assign \new_[53007]_  = ~A233 & ~A232;
  assign \new_[53008]_  = \new_[53007]_  & \new_[53004]_ ;
  assign \new_[53009]_  = \new_[53008]_  & \new_[53001]_ ;
  assign \new_[53012]_  = A265 & ~A235;
  assign \new_[53015]_  = ~A267 & A266;
  assign \new_[53016]_  = \new_[53015]_  & \new_[53012]_ ;
  assign \new_[53019]_  = ~A298 & ~A268;
  assign \new_[53022]_  = A302 & A299;
  assign \new_[53023]_  = \new_[53022]_  & \new_[53019]_ ;
  assign \new_[53024]_  = \new_[53023]_  & \new_[53016]_ ;
  assign \new_[53028]_  = ~A166 & ~A167;
  assign \new_[53029]_  = ~A169 & \new_[53028]_ ;
  assign \new_[53032]_  = A201 & A200;
  assign \new_[53035]_  = ~A235 & ~A234;
  assign \new_[53036]_  = \new_[53035]_  & \new_[53032]_ ;
  assign \new_[53037]_  = \new_[53036]_  & \new_[53029]_ ;
  assign \new_[53040]_  = A265 & ~A236;
  assign \new_[53043]_  = ~A267 & A266;
  assign \new_[53044]_  = \new_[53043]_  & \new_[53040]_ ;
  assign \new_[53047]_  = A298 & ~A268;
  assign \new_[53050]_  = A302 & ~A299;
  assign \new_[53051]_  = \new_[53050]_  & \new_[53047]_ ;
  assign \new_[53052]_  = \new_[53051]_  & \new_[53044]_ ;
  assign \new_[53056]_  = ~A166 & ~A167;
  assign \new_[53057]_  = ~A169 & \new_[53056]_ ;
  assign \new_[53060]_  = A201 & A200;
  assign \new_[53063]_  = ~A235 & ~A234;
  assign \new_[53064]_  = \new_[53063]_  & \new_[53060]_ ;
  assign \new_[53065]_  = \new_[53064]_  & \new_[53057]_ ;
  assign \new_[53068]_  = A265 & ~A236;
  assign \new_[53071]_  = ~A267 & A266;
  assign \new_[53072]_  = \new_[53071]_  & \new_[53068]_ ;
  assign \new_[53075]_  = ~A298 & ~A268;
  assign \new_[53078]_  = A302 & A299;
  assign \new_[53079]_  = \new_[53078]_  & \new_[53075]_ ;
  assign \new_[53080]_  = \new_[53079]_  & \new_[53072]_ ;
  assign \new_[53084]_  = ~A166 & ~A167;
  assign \new_[53085]_  = ~A169 & \new_[53084]_ ;
  assign \new_[53088]_  = A201 & A200;
  assign \new_[53091]_  = A233 & A232;
  assign \new_[53092]_  = \new_[53091]_  & \new_[53088]_ ;
  assign \new_[53093]_  = \new_[53092]_  & \new_[53085]_ ;
  assign \new_[53096]_  = ~A235 & ~A234;
  assign \new_[53099]_  = ~A268 & ~A267;
  assign \new_[53100]_  = \new_[53099]_  & \new_[53096]_ ;
  assign \new_[53103]_  = A298 & ~A269;
  assign \new_[53106]_  = A302 & ~A299;
  assign \new_[53107]_  = \new_[53106]_  & \new_[53103]_ ;
  assign \new_[53108]_  = \new_[53107]_  & \new_[53100]_ ;
  assign \new_[53112]_  = ~A166 & ~A167;
  assign \new_[53113]_  = ~A169 & \new_[53112]_ ;
  assign \new_[53116]_  = A201 & A200;
  assign \new_[53119]_  = A233 & A232;
  assign \new_[53120]_  = \new_[53119]_  & \new_[53116]_ ;
  assign \new_[53121]_  = \new_[53120]_  & \new_[53113]_ ;
  assign \new_[53124]_  = ~A235 & ~A234;
  assign \new_[53127]_  = ~A268 & ~A267;
  assign \new_[53128]_  = \new_[53127]_  & \new_[53124]_ ;
  assign \new_[53131]_  = ~A298 & ~A269;
  assign \new_[53134]_  = A302 & A299;
  assign \new_[53135]_  = \new_[53134]_  & \new_[53131]_ ;
  assign \new_[53136]_  = \new_[53135]_  & \new_[53128]_ ;
  assign \new_[53140]_  = ~A166 & ~A167;
  assign \new_[53141]_  = ~A169 & \new_[53140]_ ;
  assign \new_[53144]_  = A201 & A200;
  assign \new_[53147]_  = A233 & A232;
  assign \new_[53148]_  = \new_[53147]_  & \new_[53144]_ ;
  assign \new_[53149]_  = \new_[53148]_  & \new_[53141]_ ;
  assign \new_[53152]_  = ~A235 & ~A234;
  assign \new_[53155]_  = A266 & A265;
  assign \new_[53156]_  = \new_[53155]_  & \new_[53152]_ ;
  assign \new_[53159]_  = ~A268 & ~A267;
  assign \new_[53162]_  = A300 & A299;
  assign \new_[53163]_  = \new_[53162]_  & \new_[53159]_ ;
  assign \new_[53164]_  = \new_[53163]_  & \new_[53156]_ ;
  assign \new_[53168]_  = ~A166 & ~A167;
  assign \new_[53169]_  = ~A169 & \new_[53168]_ ;
  assign \new_[53172]_  = A201 & A200;
  assign \new_[53175]_  = A233 & A232;
  assign \new_[53176]_  = \new_[53175]_  & \new_[53172]_ ;
  assign \new_[53177]_  = \new_[53176]_  & \new_[53169]_ ;
  assign \new_[53180]_  = ~A235 & ~A234;
  assign \new_[53183]_  = A266 & A265;
  assign \new_[53184]_  = \new_[53183]_  & \new_[53180]_ ;
  assign \new_[53187]_  = ~A268 & ~A267;
  assign \new_[53190]_  = A300 & A298;
  assign \new_[53191]_  = \new_[53190]_  & \new_[53187]_ ;
  assign \new_[53192]_  = \new_[53191]_  & \new_[53184]_ ;
  assign \new_[53196]_  = ~A166 & ~A167;
  assign \new_[53197]_  = ~A169 & \new_[53196]_ ;
  assign \new_[53200]_  = A201 & A200;
  assign \new_[53203]_  = A233 & A232;
  assign \new_[53204]_  = \new_[53203]_  & \new_[53200]_ ;
  assign \new_[53205]_  = \new_[53204]_  & \new_[53197]_ ;
  assign \new_[53208]_  = ~A235 & ~A234;
  assign \new_[53211]_  = ~A266 & ~A265;
  assign \new_[53212]_  = \new_[53211]_  & \new_[53208]_ ;
  assign \new_[53215]_  = A298 & ~A268;
  assign \new_[53218]_  = A302 & ~A299;
  assign \new_[53219]_  = \new_[53218]_  & \new_[53215]_ ;
  assign \new_[53220]_  = \new_[53219]_  & \new_[53212]_ ;
  assign \new_[53224]_  = ~A166 & ~A167;
  assign \new_[53225]_  = ~A169 & \new_[53224]_ ;
  assign \new_[53228]_  = A201 & A200;
  assign \new_[53231]_  = A233 & A232;
  assign \new_[53232]_  = \new_[53231]_  & \new_[53228]_ ;
  assign \new_[53233]_  = \new_[53232]_  & \new_[53225]_ ;
  assign \new_[53236]_  = ~A235 & ~A234;
  assign \new_[53239]_  = ~A266 & ~A265;
  assign \new_[53240]_  = \new_[53239]_  & \new_[53236]_ ;
  assign \new_[53243]_  = ~A298 & ~A268;
  assign \new_[53246]_  = A302 & A299;
  assign \new_[53247]_  = \new_[53246]_  & \new_[53243]_ ;
  assign \new_[53248]_  = \new_[53247]_  & \new_[53240]_ ;
  assign \new_[53252]_  = ~A166 & ~A167;
  assign \new_[53253]_  = ~A169 & \new_[53252]_ ;
  assign \new_[53256]_  = A201 & A200;
  assign \new_[53259]_  = ~A233 & ~A232;
  assign \new_[53260]_  = \new_[53259]_  & \new_[53256]_ ;
  assign \new_[53261]_  = \new_[53260]_  & \new_[53253]_ ;
  assign \new_[53264]_  = A265 & ~A235;
  assign \new_[53267]_  = ~A267 & A266;
  assign \new_[53268]_  = \new_[53267]_  & \new_[53264]_ ;
  assign \new_[53271]_  = A298 & ~A268;
  assign \new_[53274]_  = A302 & ~A299;
  assign \new_[53275]_  = \new_[53274]_  & \new_[53271]_ ;
  assign \new_[53276]_  = \new_[53275]_  & \new_[53268]_ ;
  assign \new_[53280]_  = ~A166 & ~A167;
  assign \new_[53281]_  = ~A169 & \new_[53280]_ ;
  assign \new_[53284]_  = A201 & A200;
  assign \new_[53287]_  = ~A233 & ~A232;
  assign \new_[53288]_  = \new_[53287]_  & \new_[53284]_ ;
  assign \new_[53289]_  = \new_[53288]_  & \new_[53281]_ ;
  assign \new_[53292]_  = A265 & ~A235;
  assign \new_[53295]_  = ~A267 & A266;
  assign \new_[53296]_  = \new_[53295]_  & \new_[53292]_ ;
  assign \new_[53299]_  = ~A298 & ~A268;
  assign \new_[53302]_  = A302 & A299;
  assign \new_[53303]_  = \new_[53302]_  & \new_[53299]_ ;
  assign \new_[53304]_  = \new_[53303]_  & \new_[53296]_ ;
  assign \new_[53308]_  = ~A166 & ~A167;
  assign \new_[53309]_  = ~A169 & \new_[53308]_ ;
  assign \new_[53312]_  = A200 & ~A199;
  assign \new_[53315]_  = ~A234 & A203;
  assign \new_[53316]_  = \new_[53315]_  & \new_[53312]_ ;
  assign \new_[53317]_  = \new_[53316]_  & \new_[53309]_ ;
  assign \new_[53320]_  = ~A236 & ~A235;
  assign \new_[53323]_  = ~A268 & ~A267;
  assign \new_[53324]_  = \new_[53323]_  & \new_[53320]_ ;
  assign \new_[53327]_  = A298 & ~A269;
  assign \new_[53330]_  = A302 & ~A299;
  assign \new_[53331]_  = \new_[53330]_  & \new_[53327]_ ;
  assign \new_[53332]_  = \new_[53331]_  & \new_[53324]_ ;
  assign \new_[53336]_  = ~A166 & ~A167;
  assign \new_[53337]_  = ~A169 & \new_[53336]_ ;
  assign \new_[53340]_  = A200 & ~A199;
  assign \new_[53343]_  = ~A234 & A203;
  assign \new_[53344]_  = \new_[53343]_  & \new_[53340]_ ;
  assign \new_[53345]_  = \new_[53344]_  & \new_[53337]_ ;
  assign \new_[53348]_  = ~A236 & ~A235;
  assign \new_[53351]_  = ~A268 & ~A267;
  assign \new_[53352]_  = \new_[53351]_  & \new_[53348]_ ;
  assign \new_[53355]_  = ~A298 & ~A269;
  assign \new_[53358]_  = A302 & A299;
  assign \new_[53359]_  = \new_[53358]_  & \new_[53355]_ ;
  assign \new_[53360]_  = \new_[53359]_  & \new_[53352]_ ;
  assign \new_[53364]_  = ~A166 & ~A167;
  assign \new_[53365]_  = ~A169 & \new_[53364]_ ;
  assign \new_[53368]_  = A200 & ~A199;
  assign \new_[53371]_  = ~A234 & A203;
  assign \new_[53372]_  = \new_[53371]_  & \new_[53368]_ ;
  assign \new_[53373]_  = \new_[53372]_  & \new_[53365]_ ;
  assign \new_[53376]_  = ~A236 & ~A235;
  assign \new_[53379]_  = A266 & A265;
  assign \new_[53380]_  = \new_[53379]_  & \new_[53376]_ ;
  assign \new_[53383]_  = ~A268 & ~A267;
  assign \new_[53386]_  = A300 & A299;
  assign \new_[53387]_  = \new_[53386]_  & \new_[53383]_ ;
  assign \new_[53388]_  = \new_[53387]_  & \new_[53380]_ ;
  assign \new_[53392]_  = ~A166 & ~A167;
  assign \new_[53393]_  = ~A169 & \new_[53392]_ ;
  assign \new_[53396]_  = A200 & ~A199;
  assign \new_[53399]_  = ~A234 & A203;
  assign \new_[53400]_  = \new_[53399]_  & \new_[53396]_ ;
  assign \new_[53401]_  = \new_[53400]_  & \new_[53393]_ ;
  assign \new_[53404]_  = ~A236 & ~A235;
  assign \new_[53407]_  = A266 & A265;
  assign \new_[53408]_  = \new_[53407]_  & \new_[53404]_ ;
  assign \new_[53411]_  = ~A268 & ~A267;
  assign \new_[53414]_  = A300 & A298;
  assign \new_[53415]_  = \new_[53414]_  & \new_[53411]_ ;
  assign \new_[53416]_  = \new_[53415]_  & \new_[53408]_ ;
  assign \new_[53420]_  = ~A166 & ~A167;
  assign \new_[53421]_  = ~A169 & \new_[53420]_ ;
  assign \new_[53424]_  = A200 & ~A199;
  assign \new_[53427]_  = ~A234 & A203;
  assign \new_[53428]_  = \new_[53427]_  & \new_[53424]_ ;
  assign \new_[53429]_  = \new_[53428]_  & \new_[53421]_ ;
  assign \new_[53432]_  = ~A236 & ~A235;
  assign \new_[53435]_  = ~A266 & ~A265;
  assign \new_[53436]_  = \new_[53435]_  & \new_[53432]_ ;
  assign \new_[53439]_  = A298 & ~A268;
  assign \new_[53442]_  = A302 & ~A299;
  assign \new_[53443]_  = \new_[53442]_  & \new_[53439]_ ;
  assign \new_[53444]_  = \new_[53443]_  & \new_[53436]_ ;
  assign \new_[53448]_  = ~A166 & ~A167;
  assign \new_[53449]_  = ~A169 & \new_[53448]_ ;
  assign \new_[53452]_  = A200 & ~A199;
  assign \new_[53455]_  = ~A234 & A203;
  assign \new_[53456]_  = \new_[53455]_  & \new_[53452]_ ;
  assign \new_[53457]_  = \new_[53456]_  & \new_[53449]_ ;
  assign \new_[53460]_  = ~A236 & ~A235;
  assign \new_[53463]_  = ~A266 & ~A265;
  assign \new_[53464]_  = \new_[53463]_  & \new_[53460]_ ;
  assign \new_[53467]_  = ~A298 & ~A268;
  assign \new_[53470]_  = A302 & A299;
  assign \new_[53471]_  = \new_[53470]_  & \new_[53467]_ ;
  assign \new_[53472]_  = \new_[53471]_  & \new_[53464]_ ;
  assign \new_[53476]_  = ~A166 & ~A167;
  assign \new_[53477]_  = ~A169 & \new_[53476]_ ;
  assign \new_[53480]_  = A200 & ~A199;
  assign \new_[53483]_  = A232 & A203;
  assign \new_[53484]_  = \new_[53483]_  & \new_[53480]_ ;
  assign \new_[53485]_  = \new_[53484]_  & \new_[53477]_ ;
  assign \new_[53488]_  = ~A234 & A233;
  assign \new_[53491]_  = ~A267 & ~A235;
  assign \new_[53492]_  = \new_[53491]_  & \new_[53488]_ ;
  assign \new_[53495]_  = ~A269 & ~A268;
  assign \new_[53498]_  = A300 & A299;
  assign \new_[53499]_  = \new_[53498]_  & \new_[53495]_ ;
  assign \new_[53500]_  = \new_[53499]_  & \new_[53492]_ ;
  assign \new_[53504]_  = ~A166 & ~A167;
  assign \new_[53505]_  = ~A169 & \new_[53504]_ ;
  assign \new_[53508]_  = A200 & ~A199;
  assign \new_[53511]_  = A232 & A203;
  assign \new_[53512]_  = \new_[53511]_  & \new_[53508]_ ;
  assign \new_[53513]_  = \new_[53512]_  & \new_[53505]_ ;
  assign \new_[53516]_  = ~A234 & A233;
  assign \new_[53519]_  = ~A267 & ~A235;
  assign \new_[53520]_  = \new_[53519]_  & \new_[53516]_ ;
  assign \new_[53523]_  = ~A269 & ~A268;
  assign \new_[53526]_  = A300 & A298;
  assign \new_[53527]_  = \new_[53526]_  & \new_[53523]_ ;
  assign \new_[53528]_  = \new_[53527]_  & \new_[53520]_ ;
  assign \new_[53532]_  = ~A166 & ~A167;
  assign \new_[53533]_  = ~A169 & \new_[53532]_ ;
  assign \new_[53536]_  = A200 & ~A199;
  assign \new_[53539]_  = A232 & A203;
  assign \new_[53540]_  = \new_[53539]_  & \new_[53536]_ ;
  assign \new_[53541]_  = \new_[53540]_  & \new_[53533]_ ;
  assign \new_[53544]_  = ~A234 & A233;
  assign \new_[53547]_  = A265 & ~A235;
  assign \new_[53548]_  = \new_[53547]_  & \new_[53544]_ ;
  assign \new_[53551]_  = ~A267 & A266;
  assign \new_[53554]_  = A301 & ~A268;
  assign \new_[53555]_  = \new_[53554]_  & \new_[53551]_ ;
  assign \new_[53556]_  = \new_[53555]_  & \new_[53548]_ ;
  assign \new_[53560]_  = ~A166 & ~A167;
  assign \new_[53561]_  = ~A169 & \new_[53560]_ ;
  assign \new_[53564]_  = A200 & ~A199;
  assign \new_[53567]_  = A232 & A203;
  assign \new_[53568]_  = \new_[53567]_  & \new_[53564]_ ;
  assign \new_[53569]_  = \new_[53568]_  & \new_[53561]_ ;
  assign \new_[53572]_  = ~A234 & A233;
  assign \new_[53575]_  = ~A265 & ~A235;
  assign \new_[53576]_  = \new_[53575]_  & \new_[53572]_ ;
  assign \new_[53579]_  = ~A268 & ~A266;
  assign \new_[53582]_  = A300 & A299;
  assign \new_[53583]_  = \new_[53582]_  & \new_[53579]_ ;
  assign \new_[53584]_  = \new_[53583]_  & \new_[53576]_ ;
  assign \new_[53588]_  = ~A166 & ~A167;
  assign \new_[53589]_  = ~A169 & \new_[53588]_ ;
  assign \new_[53592]_  = A200 & ~A199;
  assign \new_[53595]_  = A232 & A203;
  assign \new_[53596]_  = \new_[53595]_  & \new_[53592]_ ;
  assign \new_[53597]_  = \new_[53596]_  & \new_[53589]_ ;
  assign \new_[53600]_  = ~A234 & A233;
  assign \new_[53603]_  = ~A265 & ~A235;
  assign \new_[53604]_  = \new_[53603]_  & \new_[53600]_ ;
  assign \new_[53607]_  = ~A268 & ~A266;
  assign \new_[53610]_  = A300 & A298;
  assign \new_[53611]_  = \new_[53610]_  & \new_[53607]_ ;
  assign \new_[53612]_  = \new_[53611]_  & \new_[53604]_ ;
  assign \new_[53616]_  = ~A166 & ~A167;
  assign \new_[53617]_  = ~A169 & \new_[53616]_ ;
  assign \new_[53620]_  = A200 & ~A199;
  assign \new_[53623]_  = ~A232 & A203;
  assign \new_[53624]_  = \new_[53623]_  & \new_[53620]_ ;
  assign \new_[53625]_  = \new_[53624]_  & \new_[53617]_ ;
  assign \new_[53628]_  = ~A235 & ~A233;
  assign \new_[53631]_  = ~A268 & ~A267;
  assign \new_[53632]_  = \new_[53631]_  & \new_[53628]_ ;
  assign \new_[53635]_  = A298 & ~A269;
  assign \new_[53638]_  = A302 & ~A299;
  assign \new_[53639]_  = \new_[53638]_  & \new_[53635]_ ;
  assign \new_[53640]_  = \new_[53639]_  & \new_[53632]_ ;
  assign \new_[53644]_  = ~A166 & ~A167;
  assign \new_[53645]_  = ~A169 & \new_[53644]_ ;
  assign \new_[53648]_  = A200 & ~A199;
  assign \new_[53651]_  = ~A232 & A203;
  assign \new_[53652]_  = \new_[53651]_  & \new_[53648]_ ;
  assign \new_[53653]_  = \new_[53652]_  & \new_[53645]_ ;
  assign \new_[53656]_  = ~A235 & ~A233;
  assign \new_[53659]_  = ~A268 & ~A267;
  assign \new_[53660]_  = \new_[53659]_  & \new_[53656]_ ;
  assign \new_[53663]_  = ~A298 & ~A269;
  assign \new_[53666]_  = A302 & A299;
  assign \new_[53667]_  = \new_[53666]_  & \new_[53663]_ ;
  assign \new_[53668]_  = \new_[53667]_  & \new_[53660]_ ;
  assign \new_[53672]_  = ~A166 & ~A167;
  assign \new_[53673]_  = ~A169 & \new_[53672]_ ;
  assign \new_[53676]_  = A200 & ~A199;
  assign \new_[53679]_  = ~A232 & A203;
  assign \new_[53680]_  = \new_[53679]_  & \new_[53676]_ ;
  assign \new_[53681]_  = \new_[53680]_  & \new_[53673]_ ;
  assign \new_[53684]_  = ~A235 & ~A233;
  assign \new_[53687]_  = A266 & A265;
  assign \new_[53688]_  = \new_[53687]_  & \new_[53684]_ ;
  assign \new_[53691]_  = ~A268 & ~A267;
  assign \new_[53694]_  = A300 & A299;
  assign \new_[53695]_  = \new_[53694]_  & \new_[53691]_ ;
  assign \new_[53696]_  = \new_[53695]_  & \new_[53688]_ ;
  assign \new_[53700]_  = ~A166 & ~A167;
  assign \new_[53701]_  = ~A169 & \new_[53700]_ ;
  assign \new_[53704]_  = A200 & ~A199;
  assign \new_[53707]_  = ~A232 & A203;
  assign \new_[53708]_  = \new_[53707]_  & \new_[53704]_ ;
  assign \new_[53709]_  = \new_[53708]_  & \new_[53701]_ ;
  assign \new_[53712]_  = ~A235 & ~A233;
  assign \new_[53715]_  = A266 & A265;
  assign \new_[53716]_  = \new_[53715]_  & \new_[53712]_ ;
  assign \new_[53719]_  = ~A268 & ~A267;
  assign \new_[53722]_  = A300 & A298;
  assign \new_[53723]_  = \new_[53722]_  & \new_[53719]_ ;
  assign \new_[53724]_  = \new_[53723]_  & \new_[53716]_ ;
  assign \new_[53728]_  = ~A166 & ~A167;
  assign \new_[53729]_  = ~A169 & \new_[53728]_ ;
  assign \new_[53732]_  = A200 & ~A199;
  assign \new_[53735]_  = ~A232 & A203;
  assign \new_[53736]_  = \new_[53735]_  & \new_[53732]_ ;
  assign \new_[53737]_  = \new_[53736]_  & \new_[53729]_ ;
  assign \new_[53740]_  = ~A235 & ~A233;
  assign \new_[53743]_  = ~A266 & ~A265;
  assign \new_[53744]_  = \new_[53743]_  & \new_[53740]_ ;
  assign \new_[53747]_  = A298 & ~A268;
  assign \new_[53750]_  = A302 & ~A299;
  assign \new_[53751]_  = \new_[53750]_  & \new_[53747]_ ;
  assign \new_[53752]_  = \new_[53751]_  & \new_[53744]_ ;
  assign \new_[53756]_  = ~A166 & ~A167;
  assign \new_[53757]_  = ~A169 & \new_[53756]_ ;
  assign \new_[53760]_  = A200 & ~A199;
  assign \new_[53763]_  = ~A232 & A203;
  assign \new_[53764]_  = \new_[53763]_  & \new_[53760]_ ;
  assign \new_[53765]_  = \new_[53764]_  & \new_[53757]_ ;
  assign \new_[53768]_  = ~A235 & ~A233;
  assign \new_[53771]_  = ~A266 & ~A265;
  assign \new_[53772]_  = \new_[53771]_  & \new_[53768]_ ;
  assign \new_[53775]_  = ~A298 & ~A268;
  assign \new_[53778]_  = A302 & A299;
  assign \new_[53779]_  = \new_[53778]_  & \new_[53775]_ ;
  assign \new_[53780]_  = \new_[53779]_  & \new_[53772]_ ;
  assign \new_[53784]_  = ~A166 & ~A167;
  assign \new_[53785]_  = ~A169 & \new_[53784]_ ;
  assign \new_[53788]_  = ~A200 & A199;
  assign \new_[53791]_  = ~A234 & A203;
  assign \new_[53792]_  = \new_[53791]_  & \new_[53788]_ ;
  assign \new_[53793]_  = \new_[53792]_  & \new_[53785]_ ;
  assign \new_[53796]_  = ~A236 & ~A235;
  assign \new_[53799]_  = ~A268 & ~A267;
  assign \new_[53800]_  = \new_[53799]_  & \new_[53796]_ ;
  assign \new_[53803]_  = A298 & ~A269;
  assign \new_[53806]_  = A302 & ~A299;
  assign \new_[53807]_  = \new_[53806]_  & \new_[53803]_ ;
  assign \new_[53808]_  = \new_[53807]_  & \new_[53800]_ ;
  assign \new_[53812]_  = ~A166 & ~A167;
  assign \new_[53813]_  = ~A169 & \new_[53812]_ ;
  assign \new_[53816]_  = ~A200 & A199;
  assign \new_[53819]_  = ~A234 & A203;
  assign \new_[53820]_  = \new_[53819]_  & \new_[53816]_ ;
  assign \new_[53821]_  = \new_[53820]_  & \new_[53813]_ ;
  assign \new_[53824]_  = ~A236 & ~A235;
  assign \new_[53827]_  = ~A268 & ~A267;
  assign \new_[53828]_  = \new_[53827]_  & \new_[53824]_ ;
  assign \new_[53831]_  = ~A298 & ~A269;
  assign \new_[53834]_  = A302 & A299;
  assign \new_[53835]_  = \new_[53834]_  & \new_[53831]_ ;
  assign \new_[53836]_  = \new_[53835]_  & \new_[53828]_ ;
  assign \new_[53840]_  = ~A166 & ~A167;
  assign \new_[53841]_  = ~A169 & \new_[53840]_ ;
  assign \new_[53844]_  = ~A200 & A199;
  assign \new_[53847]_  = ~A234 & A203;
  assign \new_[53848]_  = \new_[53847]_  & \new_[53844]_ ;
  assign \new_[53849]_  = \new_[53848]_  & \new_[53841]_ ;
  assign \new_[53852]_  = ~A236 & ~A235;
  assign \new_[53855]_  = A266 & A265;
  assign \new_[53856]_  = \new_[53855]_  & \new_[53852]_ ;
  assign \new_[53859]_  = ~A268 & ~A267;
  assign \new_[53862]_  = A300 & A299;
  assign \new_[53863]_  = \new_[53862]_  & \new_[53859]_ ;
  assign \new_[53864]_  = \new_[53863]_  & \new_[53856]_ ;
  assign \new_[53868]_  = ~A166 & ~A167;
  assign \new_[53869]_  = ~A169 & \new_[53868]_ ;
  assign \new_[53872]_  = ~A200 & A199;
  assign \new_[53875]_  = ~A234 & A203;
  assign \new_[53876]_  = \new_[53875]_  & \new_[53872]_ ;
  assign \new_[53877]_  = \new_[53876]_  & \new_[53869]_ ;
  assign \new_[53880]_  = ~A236 & ~A235;
  assign \new_[53883]_  = A266 & A265;
  assign \new_[53884]_  = \new_[53883]_  & \new_[53880]_ ;
  assign \new_[53887]_  = ~A268 & ~A267;
  assign \new_[53890]_  = A300 & A298;
  assign \new_[53891]_  = \new_[53890]_  & \new_[53887]_ ;
  assign \new_[53892]_  = \new_[53891]_  & \new_[53884]_ ;
  assign \new_[53896]_  = ~A166 & ~A167;
  assign \new_[53897]_  = ~A169 & \new_[53896]_ ;
  assign \new_[53900]_  = ~A200 & A199;
  assign \new_[53903]_  = ~A234 & A203;
  assign \new_[53904]_  = \new_[53903]_  & \new_[53900]_ ;
  assign \new_[53905]_  = \new_[53904]_  & \new_[53897]_ ;
  assign \new_[53908]_  = ~A236 & ~A235;
  assign \new_[53911]_  = ~A266 & ~A265;
  assign \new_[53912]_  = \new_[53911]_  & \new_[53908]_ ;
  assign \new_[53915]_  = A298 & ~A268;
  assign \new_[53918]_  = A302 & ~A299;
  assign \new_[53919]_  = \new_[53918]_  & \new_[53915]_ ;
  assign \new_[53920]_  = \new_[53919]_  & \new_[53912]_ ;
  assign \new_[53924]_  = ~A166 & ~A167;
  assign \new_[53925]_  = ~A169 & \new_[53924]_ ;
  assign \new_[53928]_  = ~A200 & A199;
  assign \new_[53931]_  = ~A234 & A203;
  assign \new_[53932]_  = \new_[53931]_  & \new_[53928]_ ;
  assign \new_[53933]_  = \new_[53932]_  & \new_[53925]_ ;
  assign \new_[53936]_  = ~A236 & ~A235;
  assign \new_[53939]_  = ~A266 & ~A265;
  assign \new_[53940]_  = \new_[53939]_  & \new_[53936]_ ;
  assign \new_[53943]_  = ~A298 & ~A268;
  assign \new_[53946]_  = A302 & A299;
  assign \new_[53947]_  = \new_[53946]_  & \new_[53943]_ ;
  assign \new_[53948]_  = \new_[53947]_  & \new_[53940]_ ;
  assign \new_[53952]_  = ~A166 & ~A167;
  assign \new_[53953]_  = ~A169 & \new_[53952]_ ;
  assign \new_[53956]_  = ~A200 & A199;
  assign \new_[53959]_  = A232 & A203;
  assign \new_[53960]_  = \new_[53959]_  & \new_[53956]_ ;
  assign \new_[53961]_  = \new_[53960]_  & \new_[53953]_ ;
  assign \new_[53964]_  = ~A234 & A233;
  assign \new_[53967]_  = ~A267 & ~A235;
  assign \new_[53968]_  = \new_[53967]_  & \new_[53964]_ ;
  assign \new_[53971]_  = ~A269 & ~A268;
  assign \new_[53974]_  = A300 & A299;
  assign \new_[53975]_  = \new_[53974]_  & \new_[53971]_ ;
  assign \new_[53976]_  = \new_[53975]_  & \new_[53968]_ ;
  assign \new_[53980]_  = ~A166 & ~A167;
  assign \new_[53981]_  = ~A169 & \new_[53980]_ ;
  assign \new_[53984]_  = ~A200 & A199;
  assign \new_[53987]_  = A232 & A203;
  assign \new_[53988]_  = \new_[53987]_  & \new_[53984]_ ;
  assign \new_[53989]_  = \new_[53988]_  & \new_[53981]_ ;
  assign \new_[53992]_  = ~A234 & A233;
  assign \new_[53995]_  = ~A267 & ~A235;
  assign \new_[53996]_  = \new_[53995]_  & \new_[53992]_ ;
  assign \new_[53999]_  = ~A269 & ~A268;
  assign \new_[54002]_  = A300 & A298;
  assign \new_[54003]_  = \new_[54002]_  & \new_[53999]_ ;
  assign \new_[54004]_  = \new_[54003]_  & \new_[53996]_ ;
  assign \new_[54008]_  = ~A166 & ~A167;
  assign \new_[54009]_  = ~A169 & \new_[54008]_ ;
  assign \new_[54012]_  = ~A200 & A199;
  assign \new_[54015]_  = A232 & A203;
  assign \new_[54016]_  = \new_[54015]_  & \new_[54012]_ ;
  assign \new_[54017]_  = \new_[54016]_  & \new_[54009]_ ;
  assign \new_[54020]_  = ~A234 & A233;
  assign \new_[54023]_  = A265 & ~A235;
  assign \new_[54024]_  = \new_[54023]_  & \new_[54020]_ ;
  assign \new_[54027]_  = ~A267 & A266;
  assign \new_[54030]_  = A301 & ~A268;
  assign \new_[54031]_  = \new_[54030]_  & \new_[54027]_ ;
  assign \new_[54032]_  = \new_[54031]_  & \new_[54024]_ ;
  assign \new_[54036]_  = ~A166 & ~A167;
  assign \new_[54037]_  = ~A169 & \new_[54036]_ ;
  assign \new_[54040]_  = ~A200 & A199;
  assign \new_[54043]_  = A232 & A203;
  assign \new_[54044]_  = \new_[54043]_  & \new_[54040]_ ;
  assign \new_[54045]_  = \new_[54044]_  & \new_[54037]_ ;
  assign \new_[54048]_  = ~A234 & A233;
  assign \new_[54051]_  = ~A265 & ~A235;
  assign \new_[54052]_  = \new_[54051]_  & \new_[54048]_ ;
  assign \new_[54055]_  = ~A268 & ~A266;
  assign \new_[54058]_  = A300 & A299;
  assign \new_[54059]_  = \new_[54058]_  & \new_[54055]_ ;
  assign \new_[54060]_  = \new_[54059]_  & \new_[54052]_ ;
  assign \new_[54064]_  = ~A166 & ~A167;
  assign \new_[54065]_  = ~A169 & \new_[54064]_ ;
  assign \new_[54068]_  = ~A200 & A199;
  assign \new_[54071]_  = A232 & A203;
  assign \new_[54072]_  = \new_[54071]_  & \new_[54068]_ ;
  assign \new_[54073]_  = \new_[54072]_  & \new_[54065]_ ;
  assign \new_[54076]_  = ~A234 & A233;
  assign \new_[54079]_  = ~A265 & ~A235;
  assign \new_[54080]_  = \new_[54079]_  & \new_[54076]_ ;
  assign \new_[54083]_  = ~A268 & ~A266;
  assign \new_[54086]_  = A300 & A298;
  assign \new_[54087]_  = \new_[54086]_  & \new_[54083]_ ;
  assign \new_[54088]_  = \new_[54087]_  & \new_[54080]_ ;
  assign \new_[54092]_  = ~A166 & ~A167;
  assign \new_[54093]_  = ~A169 & \new_[54092]_ ;
  assign \new_[54096]_  = ~A200 & A199;
  assign \new_[54099]_  = ~A232 & A203;
  assign \new_[54100]_  = \new_[54099]_  & \new_[54096]_ ;
  assign \new_[54101]_  = \new_[54100]_  & \new_[54093]_ ;
  assign \new_[54104]_  = ~A235 & ~A233;
  assign \new_[54107]_  = ~A268 & ~A267;
  assign \new_[54108]_  = \new_[54107]_  & \new_[54104]_ ;
  assign \new_[54111]_  = A298 & ~A269;
  assign \new_[54114]_  = A302 & ~A299;
  assign \new_[54115]_  = \new_[54114]_  & \new_[54111]_ ;
  assign \new_[54116]_  = \new_[54115]_  & \new_[54108]_ ;
  assign \new_[54120]_  = ~A166 & ~A167;
  assign \new_[54121]_  = ~A169 & \new_[54120]_ ;
  assign \new_[54124]_  = ~A200 & A199;
  assign \new_[54127]_  = ~A232 & A203;
  assign \new_[54128]_  = \new_[54127]_  & \new_[54124]_ ;
  assign \new_[54129]_  = \new_[54128]_  & \new_[54121]_ ;
  assign \new_[54132]_  = ~A235 & ~A233;
  assign \new_[54135]_  = ~A268 & ~A267;
  assign \new_[54136]_  = \new_[54135]_  & \new_[54132]_ ;
  assign \new_[54139]_  = ~A298 & ~A269;
  assign \new_[54142]_  = A302 & A299;
  assign \new_[54143]_  = \new_[54142]_  & \new_[54139]_ ;
  assign \new_[54144]_  = \new_[54143]_  & \new_[54136]_ ;
  assign \new_[54148]_  = ~A166 & ~A167;
  assign \new_[54149]_  = ~A169 & \new_[54148]_ ;
  assign \new_[54152]_  = ~A200 & A199;
  assign \new_[54155]_  = ~A232 & A203;
  assign \new_[54156]_  = \new_[54155]_  & \new_[54152]_ ;
  assign \new_[54157]_  = \new_[54156]_  & \new_[54149]_ ;
  assign \new_[54160]_  = ~A235 & ~A233;
  assign \new_[54163]_  = A266 & A265;
  assign \new_[54164]_  = \new_[54163]_  & \new_[54160]_ ;
  assign \new_[54167]_  = ~A268 & ~A267;
  assign \new_[54170]_  = A300 & A299;
  assign \new_[54171]_  = \new_[54170]_  & \new_[54167]_ ;
  assign \new_[54172]_  = \new_[54171]_  & \new_[54164]_ ;
  assign \new_[54176]_  = ~A166 & ~A167;
  assign \new_[54177]_  = ~A169 & \new_[54176]_ ;
  assign \new_[54180]_  = ~A200 & A199;
  assign \new_[54183]_  = ~A232 & A203;
  assign \new_[54184]_  = \new_[54183]_  & \new_[54180]_ ;
  assign \new_[54185]_  = \new_[54184]_  & \new_[54177]_ ;
  assign \new_[54188]_  = ~A235 & ~A233;
  assign \new_[54191]_  = A266 & A265;
  assign \new_[54192]_  = \new_[54191]_  & \new_[54188]_ ;
  assign \new_[54195]_  = ~A268 & ~A267;
  assign \new_[54198]_  = A300 & A298;
  assign \new_[54199]_  = \new_[54198]_  & \new_[54195]_ ;
  assign \new_[54200]_  = \new_[54199]_  & \new_[54192]_ ;
  assign \new_[54204]_  = ~A166 & ~A167;
  assign \new_[54205]_  = ~A169 & \new_[54204]_ ;
  assign \new_[54208]_  = ~A200 & A199;
  assign \new_[54211]_  = ~A232 & A203;
  assign \new_[54212]_  = \new_[54211]_  & \new_[54208]_ ;
  assign \new_[54213]_  = \new_[54212]_  & \new_[54205]_ ;
  assign \new_[54216]_  = ~A235 & ~A233;
  assign \new_[54219]_  = ~A266 & ~A265;
  assign \new_[54220]_  = \new_[54219]_  & \new_[54216]_ ;
  assign \new_[54223]_  = A298 & ~A268;
  assign \new_[54226]_  = A302 & ~A299;
  assign \new_[54227]_  = \new_[54226]_  & \new_[54223]_ ;
  assign \new_[54228]_  = \new_[54227]_  & \new_[54220]_ ;
  assign \new_[54232]_  = ~A166 & ~A167;
  assign \new_[54233]_  = ~A169 & \new_[54232]_ ;
  assign \new_[54236]_  = ~A200 & A199;
  assign \new_[54239]_  = ~A232 & A203;
  assign \new_[54240]_  = \new_[54239]_  & \new_[54236]_ ;
  assign \new_[54241]_  = \new_[54240]_  & \new_[54233]_ ;
  assign \new_[54244]_  = ~A235 & ~A233;
  assign \new_[54247]_  = ~A266 & ~A265;
  assign \new_[54248]_  = \new_[54247]_  & \new_[54244]_ ;
  assign \new_[54251]_  = ~A298 & ~A268;
  assign \new_[54254]_  = A302 & A299;
  assign \new_[54255]_  = \new_[54254]_  & \new_[54251]_ ;
  assign \new_[54256]_  = \new_[54255]_  & \new_[54248]_ ;
  assign \new_[54260]_  = A167 & ~A168;
  assign \new_[54261]_  = ~A169 & \new_[54260]_ ;
  assign \new_[54264]_  = A202 & A166;
  assign \new_[54267]_  = ~A235 & ~A234;
  assign \new_[54268]_  = \new_[54267]_  & \new_[54264]_ ;
  assign \new_[54269]_  = \new_[54268]_  & \new_[54261]_ ;
  assign \new_[54272]_  = A265 & ~A236;
  assign \new_[54275]_  = ~A267 & A266;
  assign \new_[54276]_  = \new_[54275]_  & \new_[54272]_ ;
  assign \new_[54279]_  = A298 & ~A268;
  assign \new_[54282]_  = A302 & ~A299;
  assign \new_[54283]_  = \new_[54282]_  & \new_[54279]_ ;
  assign \new_[54284]_  = \new_[54283]_  & \new_[54276]_ ;
  assign \new_[54288]_  = A167 & ~A168;
  assign \new_[54289]_  = ~A169 & \new_[54288]_ ;
  assign \new_[54292]_  = A202 & A166;
  assign \new_[54295]_  = ~A235 & ~A234;
  assign \new_[54296]_  = \new_[54295]_  & \new_[54292]_ ;
  assign \new_[54297]_  = \new_[54296]_  & \new_[54289]_ ;
  assign \new_[54300]_  = A265 & ~A236;
  assign \new_[54303]_  = ~A267 & A266;
  assign \new_[54304]_  = \new_[54303]_  & \new_[54300]_ ;
  assign \new_[54307]_  = ~A298 & ~A268;
  assign \new_[54310]_  = A302 & A299;
  assign \new_[54311]_  = \new_[54310]_  & \new_[54307]_ ;
  assign \new_[54312]_  = \new_[54311]_  & \new_[54304]_ ;
  assign \new_[54316]_  = A167 & ~A168;
  assign \new_[54317]_  = ~A169 & \new_[54316]_ ;
  assign \new_[54320]_  = A202 & A166;
  assign \new_[54323]_  = A233 & A232;
  assign \new_[54324]_  = \new_[54323]_  & \new_[54320]_ ;
  assign \new_[54325]_  = \new_[54324]_  & \new_[54317]_ ;
  assign \new_[54328]_  = ~A235 & ~A234;
  assign \new_[54331]_  = ~A268 & ~A267;
  assign \new_[54332]_  = \new_[54331]_  & \new_[54328]_ ;
  assign \new_[54335]_  = A298 & ~A269;
  assign \new_[54338]_  = A302 & ~A299;
  assign \new_[54339]_  = \new_[54338]_  & \new_[54335]_ ;
  assign \new_[54340]_  = \new_[54339]_  & \new_[54332]_ ;
  assign \new_[54344]_  = A167 & ~A168;
  assign \new_[54345]_  = ~A169 & \new_[54344]_ ;
  assign \new_[54348]_  = A202 & A166;
  assign \new_[54351]_  = A233 & A232;
  assign \new_[54352]_  = \new_[54351]_  & \new_[54348]_ ;
  assign \new_[54353]_  = \new_[54352]_  & \new_[54345]_ ;
  assign \new_[54356]_  = ~A235 & ~A234;
  assign \new_[54359]_  = ~A268 & ~A267;
  assign \new_[54360]_  = \new_[54359]_  & \new_[54356]_ ;
  assign \new_[54363]_  = ~A298 & ~A269;
  assign \new_[54366]_  = A302 & A299;
  assign \new_[54367]_  = \new_[54366]_  & \new_[54363]_ ;
  assign \new_[54368]_  = \new_[54367]_  & \new_[54360]_ ;
  assign \new_[54372]_  = A167 & ~A168;
  assign \new_[54373]_  = ~A169 & \new_[54372]_ ;
  assign \new_[54376]_  = A202 & A166;
  assign \new_[54379]_  = A233 & A232;
  assign \new_[54380]_  = \new_[54379]_  & \new_[54376]_ ;
  assign \new_[54381]_  = \new_[54380]_  & \new_[54373]_ ;
  assign \new_[54384]_  = ~A235 & ~A234;
  assign \new_[54387]_  = A266 & A265;
  assign \new_[54388]_  = \new_[54387]_  & \new_[54384]_ ;
  assign \new_[54391]_  = ~A268 & ~A267;
  assign \new_[54394]_  = A300 & A299;
  assign \new_[54395]_  = \new_[54394]_  & \new_[54391]_ ;
  assign \new_[54396]_  = \new_[54395]_  & \new_[54388]_ ;
  assign \new_[54400]_  = A167 & ~A168;
  assign \new_[54401]_  = ~A169 & \new_[54400]_ ;
  assign \new_[54404]_  = A202 & A166;
  assign \new_[54407]_  = A233 & A232;
  assign \new_[54408]_  = \new_[54407]_  & \new_[54404]_ ;
  assign \new_[54409]_  = \new_[54408]_  & \new_[54401]_ ;
  assign \new_[54412]_  = ~A235 & ~A234;
  assign \new_[54415]_  = A266 & A265;
  assign \new_[54416]_  = \new_[54415]_  & \new_[54412]_ ;
  assign \new_[54419]_  = ~A268 & ~A267;
  assign \new_[54422]_  = A300 & A298;
  assign \new_[54423]_  = \new_[54422]_  & \new_[54419]_ ;
  assign \new_[54424]_  = \new_[54423]_  & \new_[54416]_ ;
  assign \new_[54428]_  = A167 & ~A168;
  assign \new_[54429]_  = ~A169 & \new_[54428]_ ;
  assign \new_[54432]_  = A202 & A166;
  assign \new_[54435]_  = A233 & A232;
  assign \new_[54436]_  = \new_[54435]_  & \new_[54432]_ ;
  assign \new_[54437]_  = \new_[54436]_  & \new_[54429]_ ;
  assign \new_[54440]_  = ~A235 & ~A234;
  assign \new_[54443]_  = ~A266 & ~A265;
  assign \new_[54444]_  = \new_[54443]_  & \new_[54440]_ ;
  assign \new_[54447]_  = A298 & ~A268;
  assign \new_[54450]_  = A302 & ~A299;
  assign \new_[54451]_  = \new_[54450]_  & \new_[54447]_ ;
  assign \new_[54452]_  = \new_[54451]_  & \new_[54444]_ ;
  assign \new_[54456]_  = A167 & ~A168;
  assign \new_[54457]_  = ~A169 & \new_[54456]_ ;
  assign \new_[54460]_  = A202 & A166;
  assign \new_[54463]_  = A233 & A232;
  assign \new_[54464]_  = \new_[54463]_  & \new_[54460]_ ;
  assign \new_[54465]_  = \new_[54464]_  & \new_[54457]_ ;
  assign \new_[54468]_  = ~A235 & ~A234;
  assign \new_[54471]_  = ~A266 & ~A265;
  assign \new_[54472]_  = \new_[54471]_  & \new_[54468]_ ;
  assign \new_[54475]_  = ~A298 & ~A268;
  assign \new_[54478]_  = A302 & A299;
  assign \new_[54479]_  = \new_[54478]_  & \new_[54475]_ ;
  assign \new_[54480]_  = \new_[54479]_  & \new_[54472]_ ;
  assign \new_[54484]_  = A167 & ~A168;
  assign \new_[54485]_  = ~A169 & \new_[54484]_ ;
  assign \new_[54488]_  = A202 & A166;
  assign \new_[54491]_  = ~A233 & ~A232;
  assign \new_[54492]_  = \new_[54491]_  & \new_[54488]_ ;
  assign \new_[54493]_  = \new_[54492]_  & \new_[54485]_ ;
  assign \new_[54496]_  = A265 & ~A235;
  assign \new_[54499]_  = ~A267 & A266;
  assign \new_[54500]_  = \new_[54499]_  & \new_[54496]_ ;
  assign \new_[54503]_  = A298 & ~A268;
  assign \new_[54506]_  = A302 & ~A299;
  assign \new_[54507]_  = \new_[54506]_  & \new_[54503]_ ;
  assign \new_[54508]_  = \new_[54507]_  & \new_[54500]_ ;
  assign \new_[54512]_  = A167 & ~A168;
  assign \new_[54513]_  = ~A169 & \new_[54512]_ ;
  assign \new_[54516]_  = A202 & A166;
  assign \new_[54519]_  = ~A233 & ~A232;
  assign \new_[54520]_  = \new_[54519]_  & \new_[54516]_ ;
  assign \new_[54521]_  = \new_[54520]_  & \new_[54513]_ ;
  assign \new_[54524]_  = A265 & ~A235;
  assign \new_[54527]_  = ~A267 & A266;
  assign \new_[54528]_  = \new_[54527]_  & \new_[54524]_ ;
  assign \new_[54531]_  = ~A298 & ~A268;
  assign \new_[54534]_  = A302 & A299;
  assign \new_[54535]_  = \new_[54534]_  & \new_[54531]_ ;
  assign \new_[54536]_  = \new_[54535]_  & \new_[54528]_ ;
  assign \new_[54540]_  = A167 & ~A168;
  assign \new_[54541]_  = ~A169 & \new_[54540]_ ;
  assign \new_[54544]_  = A199 & A166;
  assign \new_[54547]_  = ~A234 & A201;
  assign \new_[54548]_  = \new_[54547]_  & \new_[54544]_ ;
  assign \new_[54549]_  = \new_[54548]_  & \new_[54541]_ ;
  assign \new_[54552]_  = ~A236 & ~A235;
  assign \new_[54555]_  = ~A268 & ~A267;
  assign \new_[54556]_  = \new_[54555]_  & \new_[54552]_ ;
  assign \new_[54559]_  = A298 & ~A269;
  assign \new_[54562]_  = A302 & ~A299;
  assign \new_[54563]_  = \new_[54562]_  & \new_[54559]_ ;
  assign \new_[54564]_  = \new_[54563]_  & \new_[54556]_ ;
  assign \new_[54568]_  = A167 & ~A168;
  assign \new_[54569]_  = ~A169 & \new_[54568]_ ;
  assign \new_[54572]_  = A199 & A166;
  assign \new_[54575]_  = ~A234 & A201;
  assign \new_[54576]_  = \new_[54575]_  & \new_[54572]_ ;
  assign \new_[54577]_  = \new_[54576]_  & \new_[54569]_ ;
  assign \new_[54580]_  = ~A236 & ~A235;
  assign \new_[54583]_  = ~A268 & ~A267;
  assign \new_[54584]_  = \new_[54583]_  & \new_[54580]_ ;
  assign \new_[54587]_  = ~A298 & ~A269;
  assign \new_[54590]_  = A302 & A299;
  assign \new_[54591]_  = \new_[54590]_  & \new_[54587]_ ;
  assign \new_[54592]_  = \new_[54591]_  & \new_[54584]_ ;
  assign \new_[54596]_  = A167 & ~A168;
  assign \new_[54597]_  = ~A169 & \new_[54596]_ ;
  assign \new_[54600]_  = A199 & A166;
  assign \new_[54603]_  = ~A234 & A201;
  assign \new_[54604]_  = \new_[54603]_  & \new_[54600]_ ;
  assign \new_[54605]_  = \new_[54604]_  & \new_[54597]_ ;
  assign \new_[54608]_  = ~A236 & ~A235;
  assign \new_[54611]_  = A266 & A265;
  assign \new_[54612]_  = \new_[54611]_  & \new_[54608]_ ;
  assign \new_[54615]_  = ~A268 & ~A267;
  assign \new_[54618]_  = A300 & A299;
  assign \new_[54619]_  = \new_[54618]_  & \new_[54615]_ ;
  assign \new_[54620]_  = \new_[54619]_  & \new_[54612]_ ;
  assign \new_[54624]_  = A167 & ~A168;
  assign \new_[54625]_  = ~A169 & \new_[54624]_ ;
  assign \new_[54628]_  = A199 & A166;
  assign \new_[54631]_  = ~A234 & A201;
  assign \new_[54632]_  = \new_[54631]_  & \new_[54628]_ ;
  assign \new_[54633]_  = \new_[54632]_  & \new_[54625]_ ;
  assign \new_[54636]_  = ~A236 & ~A235;
  assign \new_[54639]_  = A266 & A265;
  assign \new_[54640]_  = \new_[54639]_  & \new_[54636]_ ;
  assign \new_[54643]_  = ~A268 & ~A267;
  assign \new_[54646]_  = A300 & A298;
  assign \new_[54647]_  = \new_[54646]_  & \new_[54643]_ ;
  assign \new_[54648]_  = \new_[54647]_  & \new_[54640]_ ;
  assign \new_[54652]_  = A167 & ~A168;
  assign \new_[54653]_  = ~A169 & \new_[54652]_ ;
  assign \new_[54656]_  = A199 & A166;
  assign \new_[54659]_  = ~A234 & A201;
  assign \new_[54660]_  = \new_[54659]_  & \new_[54656]_ ;
  assign \new_[54661]_  = \new_[54660]_  & \new_[54653]_ ;
  assign \new_[54664]_  = ~A236 & ~A235;
  assign \new_[54667]_  = ~A266 & ~A265;
  assign \new_[54668]_  = \new_[54667]_  & \new_[54664]_ ;
  assign \new_[54671]_  = A298 & ~A268;
  assign \new_[54674]_  = A302 & ~A299;
  assign \new_[54675]_  = \new_[54674]_  & \new_[54671]_ ;
  assign \new_[54676]_  = \new_[54675]_  & \new_[54668]_ ;
  assign \new_[54680]_  = A167 & ~A168;
  assign \new_[54681]_  = ~A169 & \new_[54680]_ ;
  assign \new_[54684]_  = A199 & A166;
  assign \new_[54687]_  = ~A234 & A201;
  assign \new_[54688]_  = \new_[54687]_  & \new_[54684]_ ;
  assign \new_[54689]_  = \new_[54688]_  & \new_[54681]_ ;
  assign \new_[54692]_  = ~A236 & ~A235;
  assign \new_[54695]_  = ~A266 & ~A265;
  assign \new_[54696]_  = \new_[54695]_  & \new_[54692]_ ;
  assign \new_[54699]_  = ~A298 & ~A268;
  assign \new_[54702]_  = A302 & A299;
  assign \new_[54703]_  = \new_[54702]_  & \new_[54699]_ ;
  assign \new_[54704]_  = \new_[54703]_  & \new_[54696]_ ;
  assign \new_[54708]_  = A167 & ~A168;
  assign \new_[54709]_  = ~A169 & \new_[54708]_ ;
  assign \new_[54712]_  = A199 & A166;
  assign \new_[54715]_  = A232 & A201;
  assign \new_[54716]_  = \new_[54715]_  & \new_[54712]_ ;
  assign \new_[54717]_  = \new_[54716]_  & \new_[54709]_ ;
  assign \new_[54720]_  = ~A234 & A233;
  assign \new_[54723]_  = ~A267 & ~A235;
  assign \new_[54724]_  = \new_[54723]_  & \new_[54720]_ ;
  assign \new_[54727]_  = ~A269 & ~A268;
  assign \new_[54730]_  = A300 & A299;
  assign \new_[54731]_  = \new_[54730]_  & \new_[54727]_ ;
  assign \new_[54732]_  = \new_[54731]_  & \new_[54724]_ ;
  assign \new_[54736]_  = A167 & ~A168;
  assign \new_[54737]_  = ~A169 & \new_[54736]_ ;
  assign \new_[54740]_  = A199 & A166;
  assign \new_[54743]_  = A232 & A201;
  assign \new_[54744]_  = \new_[54743]_  & \new_[54740]_ ;
  assign \new_[54745]_  = \new_[54744]_  & \new_[54737]_ ;
  assign \new_[54748]_  = ~A234 & A233;
  assign \new_[54751]_  = ~A267 & ~A235;
  assign \new_[54752]_  = \new_[54751]_  & \new_[54748]_ ;
  assign \new_[54755]_  = ~A269 & ~A268;
  assign \new_[54758]_  = A300 & A298;
  assign \new_[54759]_  = \new_[54758]_  & \new_[54755]_ ;
  assign \new_[54760]_  = \new_[54759]_  & \new_[54752]_ ;
  assign \new_[54764]_  = A167 & ~A168;
  assign \new_[54765]_  = ~A169 & \new_[54764]_ ;
  assign \new_[54768]_  = A199 & A166;
  assign \new_[54771]_  = A232 & A201;
  assign \new_[54772]_  = \new_[54771]_  & \new_[54768]_ ;
  assign \new_[54773]_  = \new_[54772]_  & \new_[54765]_ ;
  assign \new_[54776]_  = ~A234 & A233;
  assign \new_[54779]_  = A265 & ~A235;
  assign \new_[54780]_  = \new_[54779]_  & \new_[54776]_ ;
  assign \new_[54783]_  = ~A267 & A266;
  assign \new_[54786]_  = A301 & ~A268;
  assign \new_[54787]_  = \new_[54786]_  & \new_[54783]_ ;
  assign \new_[54788]_  = \new_[54787]_  & \new_[54780]_ ;
  assign \new_[54792]_  = A167 & ~A168;
  assign \new_[54793]_  = ~A169 & \new_[54792]_ ;
  assign \new_[54796]_  = A199 & A166;
  assign \new_[54799]_  = A232 & A201;
  assign \new_[54800]_  = \new_[54799]_  & \new_[54796]_ ;
  assign \new_[54801]_  = \new_[54800]_  & \new_[54793]_ ;
  assign \new_[54804]_  = ~A234 & A233;
  assign \new_[54807]_  = ~A265 & ~A235;
  assign \new_[54808]_  = \new_[54807]_  & \new_[54804]_ ;
  assign \new_[54811]_  = ~A268 & ~A266;
  assign \new_[54814]_  = A300 & A299;
  assign \new_[54815]_  = \new_[54814]_  & \new_[54811]_ ;
  assign \new_[54816]_  = \new_[54815]_  & \new_[54808]_ ;
  assign \new_[54820]_  = A167 & ~A168;
  assign \new_[54821]_  = ~A169 & \new_[54820]_ ;
  assign \new_[54824]_  = A199 & A166;
  assign \new_[54827]_  = A232 & A201;
  assign \new_[54828]_  = \new_[54827]_  & \new_[54824]_ ;
  assign \new_[54829]_  = \new_[54828]_  & \new_[54821]_ ;
  assign \new_[54832]_  = ~A234 & A233;
  assign \new_[54835]_  = ~A265 & ~A235;
  assign \new_[54836]_  = \new_[54835]_  & \new_[54832]_ ;
  assign \new_[54839]_  = ~A268 & ~A266;
  assign \new_[54842]_  = A300 & A298;
  assign \new_[54843]_  = \new_[54842]_  & \new_[54839]_ ;
  assign \new_[54844]_  = \new_[54843]_  & \new_[54836]_ ;
  assign \new_[54848]_  = A167 & ~A168;
  assign \new_[54849]_  = ~A169 & \new_[54848]_ ;
  assign \new_[54852]_  = A199 & A166;
  assign \new_[54855]_  = ~A232 & A201;
  assign \new_[54856]_  = \new_[54855]_  & \new_[54852]_ ;
  assign \new_[54857]_  = \new_[54856]_  & \new_[54849]_ ;
  assign \new_[54860]_  = ~A235 & ~A233;
  assign \new_[54863]_  = ~A268 & ~A267;
  assign \new_[54864]_  = \new_[54863]_  & \new_[54860]_ ;
  assign \new_[54867]_  = A298 & ~A269;
  assign \new_[54870]_  = A302 & ~A299;
  assign \new_[54871]_  = \new_[54870]_  & \new_[54867]_ ;
  assign \new_[54872]_  = \new_[54871]_  & \new_[54864]_ ;
  assign \new_[54876]_  = A167 & ~A168;
  assign \new_[54877]_  = ~A169 & \new_[54876]_ ;
  assign \new_[54880]_  = A199 & A166;
  assign \new_[54883]_  = ~A232 & A201;
  assign \new_[54884]_  = \new_[54883]_  & \new_[54880]_ ;
  assign \new_[54885]_  = \new_[54884]_  & \new_[54877]_ ;
  assign \new_[54888]_  = ~A235 & ~A233;
  assign \new_[54891]_  = ~A268 & ~A267;
  assign \new_[54892]_  = \new_[54891]_  & \new_[54888]_ ;
  assign \new_[54895]_  = ~A298 & ~A269;
  assign \new_[54898]_  = A302 & A299;
  assign \new_[54899]_  = \new_[54898]_  & \new_[54895]_ ;
  assign \new_[54900]_  = \new_[54899]_  & \new_[54892]_ ;
  assign \new_[54904]_  = A167 & ~A168;
  assign \new_[54905]_  = ~A169 & \new_[54904]_ ;
  assign \new_[54908]_  = A199 & A166;
  assign \new_[54911]_  = ~A232 & A201;
  assign \new_[54912]_  = \new_[54911]_  & \new_[54908]_ ;
  assign \new_[54913]_  = \new_[54912]_  & \new_[54905]_ ;
  assign \new_[54916]_  = ~A235 & ~A233;
  assign \new_[54919]_  = A266 & A265;
  assign \new_[54920]_  = \new_[54919]_  & \new_[54916]_ ;
  assign \new_[54923]_  = ~A268 & ~A267;
  assign \new_[54926]_  = A300 & A299;
  assign \new_[54927]_  = \new_[54926]_  & \new_[54923]_ ;
  assign \new_[54928]_  = \new_[54927]_  & \new_[54920]_ ;
  assign \new_[54932]_  = A167 & ~A168;
  assign \new_[54933]_  = ~A169 & \new_[54932]_ ;
  assign \new_[54936]_  = A199 & A166;
  assign \new_[54939]_  = ~A232 & A201;
  assign \new_[54940]_  = \new_[54939]_  & \new_[54936]_ ;
  assign \new_[54941]_  = \new_[54940]_  & \new_[54933]_ ;
  assign \new_[54944]_  = ~A235 & ~A233;
  assign \new_[54947]_  = A266 & A265;
  assign \new_[54948]_  = \new_[54947]_  & \new_[54944]_ ;
  assign \new_[54951]_  = ~A268 & ~A267;
  assign \new_[54954]_  = A300 & A298;
  assign \new_[54955]_  = \new_[54954]_  & \new_[54951]_ ;
  assign \new_[54956]_  = \new_[54955]_  & \new_[54948]_ ;
  assign \new_[54960]_  = A167 & ~A168;
  assign \new_[54961]_  = ~A169 & \new_[54960]_ ;
  assign \new_[54964]_  = A199 & A166;
  assign \new_[54967]_  = ~A232 & A201;
  assign \new_[54968]_  = \new_[54967]_  & \new_[54964]_ ;
  assign \new_[54969]_  = \new_[54968]_  & \new_[54961]_ ;
  assign \new_[54972]_  = ~A235 & ~A233;
  assign \new_[54975]_  = ~A266 & ~A265;
  assign \new_[54976]_  = \new_[54975]_  & \new_[54972]_ ;
  assign \new_[54979]_  = A298 & ~A268;
  assign \new_[54982]_  = A302 & ~A299;
  assign \new_[54983]_  = \new_[54982]_  & \new_[54979]_ ;
  assign \new_[54984]_  = \new_[54983]_  & \new_[54976]_ ;
  assign \new_[54988]_  = A167 & ~A168;
  assign \new_[54989]_  = ~A169 & \new_[54988]_ ;
  assign \new_[54992]_  = A199 & A166;
  assign \new_[54995]_  = ~A232 & A201;
  assign \new_[54996]_  = \new_[54995]_  & \new_[54992]_ ;
  assign \new_[54997]_  = \new_[54996]_  & \new_[54989]_ ;
  assign \new_[55000]_  = ~A235 & ~A233;
  assign \new_[55003]_  = ~A266 & ~A265;
  assign \new_[55004]_  = \new_[55003]_  & \new_[55000]_ ;
  assign \new_[55007]_  = ~A298 & ~A268;
  assign \new_[55010]_  = A302 & A299;
  assign \new_[55011]_  = \new_[55010]_  & \new_[55007]_ ;
  assign \new_[55012]_  = \new_[55011]_  & \new_[55004]_ ;
  assign \new_[55016]_  = A167 & ~A168;
  assign \new_[55017]_  = ~A169 & \new_[55016]_ ;
  assign \new_[55020]_  = A200 & A166;
  assign \new_[55023]_  = ~A234 & A201;
  assign \new_[55024]_  = \new_[55023]_  & \new_[55020]_ ;
  assign \new_[55025]_  = \new_[55024]_  & \new_[55017]_ ;
  assign \new_[55028]_  = ~A236 & ~A235;
  assign \new_[55031]_  = ~A268 & ~A267;
  assign \new_[55032]_  = \new_[55031]_  & \new_[55028]_ ;
  assign \new_[55035]_  = A298 & ~A269;
  assign \new_[55038]_  = A302 & ~A299;
  assign \new_[55039]_  = \new_[55038]_  & \new_[55035]_ ;
  assign \new_[55040]_  = \new_[55039]_  & \new_[55032]_ ;
  assign \new_[55044]_  = A167 & ~A168;
  assign \new_[55045]_  = ~A169 & \new_[55044]_ ;
  assign \new_[55048]_  = A200 & A166;
  assign \new_[55051]_  = ~A234 & A201;
  assign \new_[55052]_  = \new_[55051]_  & \new_[55048]_ ;
  assign \new_[55053]_  = \new_[55052]_  & \new_[55045]_ ;
  assign \new_[55056]_  = ~A236 & ~A235;
  assign \new_[55059]_  = ~A268 & ~A267;
  assign \new_[55060]_  = \new_[55059]_  & \new_[55056]_ ;
  assign \new_[55063]_  = ~A298 & ~A269;
  assign \new_[55066]_  = A302 & A299;
  assign \new_[55067]_  = \new_[55066]_  & \new_[55063]_ ;
  assign \new_[55068]_  = \new_[55067]_  & \new_[55060]_ ;
  assign \new_[55072]_  = A167 & ~A168;
  assign \new_[55073]_  = ~A169 & \new_[55072]_ ;
  assign \new_[55076]_  = A200 & A166;
  assign \new_[55079]_  = ~A234 & A201;
  assign \new_[55080]_  = \new_[55079]_  & \new_[55076]_ ;
  assign \new_[55081]_  = \new_[55080]_  & \new_[55073]_ ;
  assign \new_[55084]_  = ~A236 & ~A235;
  assign \new_[55087]_  = A266 & A265;
  assign \new_[55088]_  = \new_[55087]_  & \new_[55084]_ ;
  assign \new_[55091]_  = ~A268 & ~A267;
  assign \new_[55094]_  = A300 & A299;
  assign \new_[55095]_  = \new_[55094]_  & \new_[55091]_ ;
  assign \new_[55096]_  = \new_[55095]_  & \new_[55088]_ ;
  assign \new_[55100]_  = A167 & ~A168;
  assign \new_[55101]_  = ~A169 & \new_[55100]_ ;
  assign \new_[55104]_  = A200 & A166;
  assign \new_[55107]_  = ~A234 & A201;
  assign \new_[55108]_  = \new_[55107]_  & \new_[55104]_ ;
  assign \new_[55109]_  = \new_[55108]_  & \new_[55101]_ ;
  assign \new_[55112]_  = ~A236 & ~A235;
  assign \new_[55115]_  = A266 & A265;
  assign \new_[55116]_  = \new_[55115]_  & \new_[55112]_ ;
  assign \new_[55119]_  = ~A268 & ~A267;
  assign \new_[55122]_  = A300 & A298;
  assign \new_[55123]_  = \new_[55122]_  & \new_[55119]_ ;
  assign \new_[55124]_  = \new_[55123]_  & \new_[55116]_ ;
  assign \new_[55128]_  = A167 & ~A168;
  assign \new_[55129]_  = ~A169 & \new_[55128]_ ;
  assign \new_[55132]_  = A200 & A166;
  assign \new_[55135]_  = ~A234 & A201;
  assign \new_[55136]_  = \new_[55135]_  & \new_[55132]_ ;
  assign \new_[55137]_  = \new_[55136]_  & \new_[55129]_ ;
  assign \new_[55140]_  = ~A236 & ~A235;
  assign \new_[55143]_  = ~A266 & ~A265;
  assign \new_[55144]_  = \new_[55143]_  & \new_[55140]_ ;
  assign \new_[55147]_  = A298 & ~A268;
  assign \new_[55150]_  = A302 & ~A299;
  assign \new_[55151]_  = \new_[55150]_  & \new_[55147]_ ;
  assign \new_[55152]_  = \new_[55151]_  & \new_[55144]_ ;
  assign \new_[55156]_  = A167 & ~A168;
  assign \new_[55157]_  = ~A169 & \new_[55156]_ ;
  assign \new_[55160]_  = A200 & A166;
  assign \new_[55163]_  = ~A234 & A201;
  assign \new_[55164]_  = \new_[55163]_  & \new_[55160]_ ;
  assign \new_[55165]_  = \new_[55164]_  & \new_[55157]_ ;
  assign \new_[55168]_  = ~A236 & ~A235;
  assign \new_[55171]_  = ~A266 & ~A265;
  assign \new_[55172]_  = \new_[55171]_  & \new_[55168]_ ;
  assign \new_[55175]_  = ~A298 & ~A268;
  assign \new_[55178]_  = A302 & A299;
  assign \new_[55179]_  = \new_[55178]_  & \new_[55175]_ ;
  assign \new_[55180]_  = \new_[55179]_  & \new_[55172]_ ;
  assign \new_[55184]_  = A167 & ~A168;
  assign \new_[55185]_  = ~A169 & \new_[55184]_ ;
  assign \new_[55188]_  = A200 & A166;
  assign \new_[55191]_  = A232 & A201;
  assign \new_[55192]_  = \new_[55191]_  & \new_[55188]_ ;
  assign \new_[55193]_  = \new_[55192]_  & \new_[55185]_ ;
  assign \new_[55196]_  = ~A234 & A233;
  assign \new_[55199]_  = ~A267 & ~A235;
  assign \new_[55200]_  = \new_[55199]_  & \new_[55196]_ ;
  assign \new_[55203]_  = ~A269 & ~A268;
  assign \new_[55206]_  = A300 & A299;
  assign \new_[55207]_  = \new_[55206]_  & \new_[55203]_ ;
  assign \new_[55208]_  = \new_[55207]_  & \new_[55200]_ ;
  assign \new_[55212]_  = A167 & ~A168;
  assign \new_[55213]_  = ~A169 & \new_[55212]_ ;
  assign \new_[55216]_  = A200 & A166;
  assign \new_[55219]_  = A232 & A201;
  assign \new_[55220]_  = \new_[55219]_  & \new_[55216]_ ;
  assign \new_[55221]_  = \new_[55220]_  & \new_[55213]_ ;
  assign \new_[55224]_  = ~A234 & A233;
  assign \new_[55227]_  = ~A267 & ~A235;
  assign \new_[55228]_  = \new_[55227]_  & \new_[55224]_ ;
  assign \new_[55231]_  = ~A269 & ~A268;
  assign \new_[55234]_  = A300 & A298;
  assign \new_[55235]_  = \new_[55234]_  & \new_[55231]_ ;
  assign \new_[55236]_  = \new_[55235]_  & \new_[55228]_ ;
  assign \new_[55240]_  = A167 & ~A168;
  assign \new_[55241]_  = ~A169 & \new_[55240]_ ;
  assign \new_[55244]_  = A200 & A166;
  assign \new_[55247]_  = A232 & A201;
  assign \new_[55248]_  = \new_[55247]_  & \new_[55244]_ ;
  assign \new_[55249]_  = \new_[55248]_  & \new_[55241]_ ;
  assign \new_[55252]_  = ~A234 & A233;
  assign \new_[55255]_  = A265 & ~A235;
  assign \new_[55256]_  = \new_[55255]_  & \new_[55252]_ ;
  assign \new_[55259]_  = ~A267 & A266;
  assign \new_[55262]_  = A301 & ~A268;
  assign \new_[55263]_  = \new_[55262]_  & \new_[55259]_ ;
  assign \new_[55264]_  = \new_[55263]_  & \new_[55256]_ ;
  assign \new_[55268]_  = A167 & ~A168;
  assign \new_[55269]_  = ~A169 & \new_[55268]_ ;
  assign \new_[55272]_  = A200 & A166;
  assign \new_[55275]_  = A232 & A201;
  assign \new_[55276]_  = \new_[55275]_  & \new_[55272]_ ;
  assign \new_[55277]_  = \new_[55276]_  & \new_[55269]_ ;
  assign \new_[55280]_  = ~A234 & A233;
  assign \new_[55283]_  = ~A265 & ~A235;
  assign \new_[55284]_  = \new_[55283]_  & \new_[55280]_ ;
  assign \new_[55287]_  = ~A268 & ~A266;
  assign \new_[55290]_  = A300 & A299;
  assign \new_[55291]_  = \new_[55290]_  & \new_[55287]_ ;
  assign \new_[55292]_  = \new_[55291]_  & \new_[55284]_ ;
  assign \new_[55296]_  = A167 & ~A168;
  assign \new_[55297]_  = ~A169 & \new_[55296]_ ;
  assign \new_[55300]_  = A200 & A166;
  assign \new_[55303]_  = A232 & A201;
  assign \new_[55304]_  = \new_[55303]_  & \new_[55300]_ ;
  assign \new_[55305]_  = \new_[55304]_  & \new_[55297]_ ;
  assign \new_[55308]_  = ~A234 & A233;
  assign \new_[55311]_  = ~A265 & ~A235;
  assign \new_[55312]_  = \new_[55311]_  & \new_[55308]_ ;
  assign \new_[55315]_  = ~A268 & ~A266;
  assign \new_[55318]_  = A300 & A298;
  assign \new_[55319]_  = \new_[55318]_  & \new_[55315]_ ;
  assign \new_[55320]_  = \new_[55319]_  & \new_[55312]_ ;
  assign \new_[55324]_  = A167 & ~A168;
  assign \new_[55325]_  = ~A169 & \new_[55324]_ ;
  assign \new_[55328]_  = A200 & A166;
  assign \new_[55331]_  = ~A232 & A201;
  assign \new_[55332]_  = \new_[55331]_  & \new_[55328]_ ;
  assign \new_[55333]_  = \new_[55332]_  & \new_[55325]_ ;
  assign \new_[55336]_  = ~A235 & ~A233;
  assign \new_[55339]_  = ~A268 & ~A267;
  assign \new_[55340]_  = \new_[55339]_  & \new_[55336]_ ;
  assign \new_[55343]_  = A298 & ~A269;
  assign \new_[55346]_  = A302 & ~A299;
  assign \new_[55347]_  = \new_[55346]_  & \new_[55343]_ ;
  assign \new_[55348]_  = \new_[55347]_  & \new_[55340]_ ;
  assign \new_[55352]_  = A167 & ~A168;
  assign \new_[55353]_  = ~A169 & \new_[55352]_ ;
  assign \new_[55356]_  = A200 & A166;
  assign \new_[55359]_  = ~A232 & A201;
  assign \new_[55360]_  = \new_[55359]_  & \new_[55356]_ ;
  assign \new_[55361]_  = \new_[55360]_  & \new_[55353]_ ;
  assign \new_[55364]_  = ~A235 & ~A233;
  assign \new_[55367]_  = ~A268 & ~A267;
  assign \new_[55368]_  = \new_[55367]_  & \new_[55364]_ ;
  assign \new_[55371]_  = ~A298 & ~A269;
  assign \new_[55374]_  = A302 & A299;
  assign \new_[55375]_  = \new_[55374]_  & \new_[55371]_ ;
  assign \new_[55376]_  = \new_[55375]_  & \new_[55368]_ ;
  assign \new_[55380]_  = A167 & ~A168;
  assign \new_[55381]_  = ~A169 & \new_[55380]_ ;
  assign \new_[55384]_  = A200 & A166;
  assign \new_[55387]_  = ~A232 & A201;
  assign \new_[55388]_  = \new_[55387]_  & \new_[55384]_ ;
  assign \new_[55389]_  = \new_[55388]_  & \new_[55381]_ ;
  assign \new_[55392]_  = ~A235 & ~A233;
  assign \new_[55395]_  = A266 & A265;
  assign \new_[55396]_  = \new_[55395]_  & \new_[55392]_ ;
  assign \new_[55399]_  = ~A268 & ~A267;
  assign \new_[55402]_  = A300 & A299;
  assign \new_[55403]_  = \new_[55402]_  & \new_[55399]_ ;
  assign \new_[55404]_  = \new_[55403]_  & \new_[55396]_ ;
  assign \new_[55408]_  = A167 & ~A168;
  assign \new_[55409]_  = ~A169 & \new_[55408]_ ;
  assign \new_[55412]_  = A200 & A166;
  assign \new_[55415]_  = ~A232 & A201;
  assign \new_[55416]_  = \new_[55415]_  & \new_[55412]_ ;
  assign \new_[55417]_  = \new_[55416]_  & \new_[55409]_ ;
  assign \new_[55420]_  = ~A235 & ~A233;
  assign \new_[55423]_  = A266 & A265;
  assign \new_[55424]_  = \new_[55423]_  & \new_[55420]_ ;
  assign \new_[55427]_  = ~A268 & ~A267;
  assign \new_[55430]_  = A300 & A298;
  assign \new_[55431]_  = \new_[55430]_  & \new_[55427]_ ;
  assign \new_[55432]_  = \new_[55431]_  & \new_[55424]_ ;
  assign \new_[55436]_  = A167 & ~A168;
  assign \new_[55437]_  = ~A169 & \new_[55436]_ ;
  assign \new_[55440]_  = A200 & A166;
  assign \new_[55443]_  = ~A232 & A201;
  assign \new_[55444]_  = \new_[55443]_  & \new_[55440]_ ;
  assign \new_[55445]_  = \new_[55444]_  & \new_[55437]_ ;
  assign \new_[55448]_  = ~A235 & ~A233;
  assign \new_[55451]_  = ~A266 & ~A265;
  assign \new_[55452]_  = \new_[55451]_  & \new_[55448]_ ;
  assign \new_[55455]_  = A298 & ~A268;
  assign \new_[55458]_  = A302 & ~A299;
  assign \new_[55459]_  = \new_[55458]_  & \new_[55455]_ ;
  assign \new_[55460]_  = \new_[55459]_  & \new_[55452]_ ;
  assign \new_[55464]_  = A167 & ~A168;
  assign \new_[55465]_  = ~A169 & \new_[55464]_ ;
  assign \new_[55468]_  = A200 & A166;
  assign \new_[55471]_  = ~A232 & A201;
  assign \new_[55472]_  = \new_[55471]_  & \new_[55468]_ ;
  assign \new_[55473]_  = \new_[55472]_  & \new_[55465]_ ;
  assign \new_[55476]_  = ~A235 & ~A233;
  assign \new_[55479]_  = ~A266 & ~A265;
  assign \new_[55480]_  = \new_[55479]_  & \new_[55476]_ ;
  assign \new_[55483]_  = ~A298 & ~A268;
  assign \new_[55486]_  = A302 & A299;
  assign \new_[55487]_  = \new_[55486]_  & \new_[55483]_ ;
  assign \new_[55488]_  = \new_[55487]_  & \new_[55480]_ ;
  assign \new_[55492]_  = A167 & ~A168;
  assign \new_[55493]_  = ~A169 & \new_[55492]_ ;
  assign \new_[55496]_  = ~A199 & A166;
  assign \new_[55499]_  = A203 & A200;
  assign \new_[55500]_  = \new_[55499]_  & \new_[55496]_ ;
  assign \new_[55501]_  = \new_[55500]_  & \new_[55493]_ ;
  assign \new_[55504]_  = ~A235 & ~A234;
  assign \new_[55507]_  = ~A267 & ~A236;
  assign \new_[55508]_  = \new_[55507]_  & \new_[55504]_ ;
  assign \new_[55511]_  = ~A269 & ~A268;
  assign \new_[55514]_  = A300 & A299;
  assign \new_[55515]_  = \new_[55514]_  & \new_[55511]_ ;
  assign \new_[55516]_  = \new_[55515]_  & \new_[55508]_ ;
  assign \new_[55520]_  = A167 & ~A168;
  assign \new_[55521]_  = ~A169 & \new_[55520]_ ;
  assign \new_[55524]_  = ~A199 & A166;
  assign \new_[55527]_  = A203 & A200;
  assign \new_[55528]_  = \new_[55527]_  & \new_[55524]_ ;
  assign \new_[55529]_  = \new_[55528]_  & \new_[55521]_ ;
  assign \new_[55532]_  = ~A235 & ~A234;
  assign \new_[55535]_  = ~A267 & ~A236;
  assign \new_[55536]_  = \new_[55535]_  & \new_[55532]_ ;
  assign \new_[55539]_  = ~A269 & ~A268;
  assign \new_[55542]_  = A300 & A298;
  assign \new_[55543]_  = \new_[55542]_  & \new_[55539]_ ;
  assign \new_[55544]_  = \new_[55543]_  & \new_[55536]_ ;
  assign \new_[55548]_  = A167 & ~A168;
  assign \new_[55549]_  = ~A169 & \new_[55548]_ ;
  assign \new_[55552]_  = ~A199 & A166;
  assign \new_[55555]_  = A203 & A200;
  assign \new_[55556]_  = \new_[55555]_  & \new_[55552]_ ;
  assign \new_[55557]_  = \new_[55556]_  & \new_[55549]_ ;
  assign \new_[55560]_  = ~A235 & ~A234;
  assign \new_[55563]_  = A265 & ~A236;
  assign \new_[55564]_  = \new_[55563]_  & \new_[55560]_ ;
  assign \new_[55567]_  = ~A267 & A266;
  assign \new_[55570]_  = A301 & ~A268;
  assign \new_[55571]_  = \new_[55570]_  & \new_[55567]_ ;
  assign \new_[55572]_  = \new_[55571]_  & \new_[55564]_ ;
  assign \new_[55576]_  = A167 & ~A168;
  assign \new_[55577]_  = ~A169 & \new_[55576]_ ;
  assign \new_[55580]_  = ~A199 & A166;
  assign \new_[55583]_  = A203 & A200;
  assign \new_[55584]_  = \new_[55583]_  & \new_[55580]_ ;
  assign \new_[55585]_  = \new_[55584]_  & \new_[55577]_ ;
  assign \new_[55588]_  = ~A235 & ~A234;
  assign \new_[55591]_  = ~A265 & ~A236;
  assign \new_[55592]_  = \new_[55591]_  & \new_[55588]_ ;
  assign \new_[55595]_  = ~A268 & ~A266;
  assign \new_[55598]_  = A300 & A299;
  assign \new_[55599]_  = \new_[55598]_  & \new_[55595]_ ;
  assign \new_[55600]_  = \new_[55599]_  & \new_[55592]_ ;
  assign \new_[55604]_  = A167 & ~A168;
  assign \new_[55605]_  = ~A169 & \new_[55604]_ ;
  assign \new_[55608]_  = ~A199 & A166;
  assign \new_[55611]_  = A203 & A200;
  assign \new_[55612]_  = \new_[55611]_  & \new_[55608]_ ;
  assign \new_[55613]_  = \new_[55612]_  & \new_[55605]_ ;
  assign \new_[55616]_  = ~A235 & ~A234;
  assign \new_[55619]_  = ~A265 & ~A236;
  assign \new_[55620]_  = \new_[55619]_  & \new_[55616]_ ;
  assign \new_[55623]_  = ~A268 & ~A266;
  assign \new_[55626]_  = A300 & A298;
  assign \new_[55627]_  = \new_[55626]_  & \new_[55623]_ ;
  assign \new_[55628]_  = \new_[55627]_  & \new_[55620]_ ;
  assign \new_[55632]_  = A167 & ~A168;
  assign \new_[55633]_  = ~A169 & \new_[55632]_ ;
  assign \new_[55636]_  = ~A199 & A166;
  assign \new_[55639]_  = A203 & A200;
  assign \new_[55640]_  = \new_[55639]_  & \new_[55636]_ ;
  assign \new_[55641]_  = \new_[55640]_  & \new_[55633]_ ;
  assign \new_[55644]_  = A233 & A232;
  assign \new_[55647]_  = ~A235 & ~A234;
  assign \new_[55648]_  = \new_[55647]_  & \new_[55644]_ ;
  assign \new_[55651]_  = ~A268 & ~A267;
  assign \new_[55654]_  = A301 & ~A269;
  assign \new_[55655]_  = \new_[55654]_  & \new_[55651]_ ;
  assign \new_[55656]_  = \new_[55655]_  & \new_[55648]_ ;
  assign \new_[55660]_  = A167 & ~A168;
  assign \new_[55661]_  = ~A169 & \new_[55660]_ ;
  assign \new_[55664]_  = ~A199 & A166;
  assign \new_[55667]_  = A203 & A200;
  assign \new_[55668]_  = \new_[55667]_  & \new_[55664]_ ;
  assign \new_[55669]_  = \new_[55668]_  & \new_[55661]_ ;
  assign \new_[55672]_  = A233 & A232;
  assign \new_[55675]_  = ~A235 & ~A234;
  assign \new_[55676]_  = \new_[55675]_  & \new_[55672]_ ;
  assign \new_[55679]_  = ~A266 & ~A265;
  assign \new_[55682]_  = A301 & ~A268;
  assign \new_[55683]_  = \new_[55682]_  & \new_[55679]_ ;
  assign \new_[55684]_  = \new_[55683]_  & \new_[55676]_ ;
  assign \new_[55688]_  = A167 & ~A168;
  assign \new_[55689]_  = ~A169 & \new_[55688]_ ;
  assign \new_[55692]_  = ~A199 & A166;
  assign \new_[55695]_  = A203 & A200;
  assign \new_[55696]_  = \new_[55695]_  & \new_[55692]_ ;
  assign \new_[55697]_  = \new_[55696]_  & \new_[55689]_ ;
  assign \new_[55700]_  = ~A233 & ~A232;
  assign \new_[55703]_  = ~A267 & ~A235;
  assign \new_[55704]_  = \new_[55703]_  & \new_[55700]_ ;
  assign \new_[55707]_  = ~A269 & ~A268;
  assign \new_[55710]_  = A300 & A299;
  assign \new_[55711]_  = \new_[55710]_  & \new_[55707]_ ;
  assign \new_[55712]_  = \new_[55711]_  & \new_[55704]_ ;
  assign \new_[55716]_  = A167 & ~A168;
  assign \new_[55717]_  = ~A169 & \new_[55716]_ ;
  assign \new_[55720]_  = ~A199 & A166;
  assign \new_[55723]_  = A203 & A200;
  assign \new_[55724]_  = \new_[55723]_  & \new_[55720]_ ;
  assign \new_[55725]_  = \new_[55724]_  & \new_[55717]_ ;
  assign \new_[55728]_  = ~A233 & ~A232;
  assign \new_[55731]_  = ~A267 & ~A235;
  assign \new_[55732]_  = \new_[55731]_  & \new_[55728]_ ;
  assign \new_[55735]_  = ~A269 & ~A268;
  assign \new_[55738]_  = A300 & A298;
  assign \new_[55739]_  = \new_[55738]_  & \new_[55735]_ ;
  assign \new_[55740]_  = \new_[55739]_  & \new_[55732]_ ;
  assign \new_[55744]_  = A167 & ~A168;
  assign \new_[55745]_  = ~A169 & \new_[55744]_ ;
  assign \new_[55748]_  = ~A199 & A166;
  assign \new_[55751]_  = A203 & A200;
  assign \new_[55752]_  = \new_[55751]_  & \new_[55748]_ ;
  assign \new_[55753]_  = \new_[55752]_  & \new_[55745]_ ;
  assign \new_[55756]_  = ~A233 & ~A232;
  assign \new_[55759]_  = A265 & ~A235;
  assign \new_[55760]_  = \new_[55759]_  & \new_[55756]_ ;
  assign \new_[55763]_  = ~A267 & A266;
  assign \new_[55766]_  = A301 & ~A268;
  assign \new_[55767]_  = \new_[55766]_  & \new_[55763]_ ;
  assign \new_[55768]_  = \new_[55767]_  & \new_[55760]_ ;
  assign \new_[55772]_  = A167 & ~A168;
  assign \new_[55773]_  = ~A169 & \new_[55772]_ ;
  assign \new_[55776]_  = ~A199 & A166;
  assign \new_[55779]_  = A203 & A200;
  assign \new_[55780]_  = \new_[55779]_  & \new_[55776]_ ;
  assign \new_[55781]_  = \new_[55780]_  & \new_[55773]_ ;
  assign \new_[55784]_  = ~A233 & ~A232;
  assign \new_[55787]_  = ~A265 & ~A235;
  assign \new_[55788]_  = \new_[55787]_  & \new_[55784]_ ;
  assign \new_[55791]_  = ~A268 & ~A266;
  assign \new_[55794]_  = A300 & A299;
  assign \new_[55795]_  = \new_[55794]_  & \new_[55791]_ ;
  assign \new_[55796]_  = \new_[55795]_  & \new_[55788]_ ;
  assign \new_[55800]_  = A167 & ~A168;
  assign \new_[55801]_  = ~A169 & \new_[55800]_ ;
  assign \new_[55804]_  = ~A199 & A166;
  assign \new_[55807]_  = A203 & A200;
  assign \new_[55808]_  = \new_[55807]_  & \new_[55804]_ ;
  assign \new_[55809]_  = \new_[55808]_  & \new_[55801]_ ;
  assign \new_[55812]_  = ~A233 & ~A232;
  assign \new_[55815]_  = ~A265 & ~A235;
  assign \new_[55816]_  = \new_[55815]_  & \new_[55812]_ ;
  assign \new_[55819]_  = ~A268 & ~A266;
  assign \new_[55822]_  = A300 & A298;
  assign \new_[55823]_  = \new_[55822]_  & \new_[55819]_ ;
  assign \new_[55824]_  = \new_[55823]_  & \new_[55816]_ ;
  assign \new_[55828]_  = A167 & ~A168;
  assign \new_[55829]_  = ~A169 & \new_[55828]_ ;
  assign \new_[55832]_  = A199 & A166;
  assign \new_[55835]_  = A203 & ~A200;
  assign \new_[55836]_  = \new_[55835]_  & \new_[55832]_ ;
  assign \new_[55837]_  = \new_[55836]_  & \new_[55829]_ ;
  assign \new_[55840]_  = ~A235 & ~A234;
  assign \new_[55843]_  = ~A267 & ~A236;
  assign \new_[55844]_  = \new_[55843]_  & \new_[55840]_ ;
  assign \new_[55847]_  = ~A269 & ~A268;
  assign \new_[55850]_  = A300 & A299;
  assign \new_[55851]_  = \new_[55850]_  & \new_[55847]_ ;
  assign \new_[55852]_  = \new_[55851]_  & \new_[55844]_ ;
  assign \new_[55856]_  = A167 & ~A168;
  assign \new_[55857]_  = ~A169 & \new_[55856]_ ;
  assign \new_[55860]_  = A199 & A166;
  assign \new_[55863]_  = A203 & ~A200;
  assign \new_[55864]_  = \new_[55863]_  & \new_[55860]_ ;
  assign \new_[55865]_  = \new_[55864]_  & \new_[55857]_ ;
  assign \new_[55868]_  = ~A235 & ~A234;
  assign \new_[55871]_  = ~A267 & ~A236;
  assign \new_[55872]_  = \new_[55871]_  & \new_[55868]_ ;
  assign \new_[55875]_  = ~A269 & ~A268;
  assign \new_[55878]_  = A300 & A298;
  assign \new_[55879]_  = \new_[55878]_  & \new_[55875]_ ;
  assign \new_[55880]_  = \new_[55879]_  & \new_[55872]_ ;
  assign \new_[55884]_  = A167 & ~A168;
  assign \new_[55885]_  = ~A169 & \new_[55884]_ ;
  assign \new_[55888]_  = A199 & A166;
  assign \new_[55891]_  = A203 & ~A200;
  assign \new_[55892]_  = \new_[55891]_  & \new_[55888]_ ;
  assign \new_[55893]_  = \new_[55892]_  & \new_[55885]_ ;
  assign \new_[55896]_  = ~A235 & ~A234;
  assign \new_[55899]_  = A265 & ~A236;
  assign \new_[55900]_  = \new_[55899]_  & \new_[55896]_ ;
  assign \new_[55903]_  = ~A267 & A266;
  assign \new_[55906]_  = A301 & ~A268;
  assign \new_[55907]_  = \new_[55906]_  & \new_[55903]_ ;
  assign \new_[55908]_  = \new_[55907]_  & \new_[55900]_ ;
  assign \new_[55912]_  = A167 & ~A168;
  assign \new_[55913]_  = ~A169 & \new_[55912]_ ;
  assign \new_[55916]_  = A199 & A166;
  assign \new_[55919]_  = A203 & ~A200;
  assign \new_[55920]_  = \new_[55919]_  & \new_[55916]_ ;
  assign \new_[55921]_  = \new_[55920]_  & \new_[55913]_ ;
  assign \new_[55924]_  = ~A235 & ~A234;
  assign \new_[55927]_  = ~A265 & ~A236;
  assign \new_[55928]_  = \new_[55927]_  & \new_[55924]_ ;
  assign \new_[55931]_  = ~A268 & ~A266;
  assign \new_[55934]_  = A300 & A299;
  assign \new_[55935]_  = \new_[55934]_  & \new_[55931]_ ;
  assign \new_[55936]_  = \new_[55935]_  & \new_[55928]_ ;
  assign \new_[55940]_  = A167 & ~A168;
  assign \new_[55941]_  = ~A169 & \new_[55940]_ ;
  assign \new_[55944]_  = A199 & A166;
  assign \new_[55947]_  = A203 & ~A200;
  assign \new_[55948]_  = \new_[55947]_  & \new_[55944]_ ;
  assign \new_[55949]_  = \new_[55948]_  & \new_[55941]_ ;
  assign \new_[55952]_  = ~A235 & ~A234;
  assign \new_[55955]_  = ~A265 & ~A236;
  assign \new_[55956]_  = \new_[55955]_  & \new_[55952]_ ;
  assign \new_[55959]_  = ~A268 & ~A266;
  assign \new_[55962]_  = A300 & A298;
  assign \new_[55963]_  = \new_[55962]_  & \new_[55959]_ ;
  assign \new_[55964]_  = \new_[55963]_  & \new_[55956]_ ;
  assign \new_[55968]_  = A167 & ~A168;
  assign \new_[55969]_  = ~A169 & \new_[55968]_ ;
  assign \new_[55972]_  = A199 & A166;
  assign \new_[55975]_  = A203 & ~A200;
  assign \new_[55976]_  = \new_[55975]_  & \new_[55972]_ ;
  assign \new_[55977]_  = \new_[55976]_  & \new_[55969]_ ;
  assign \new_[55980]_  = A233 & A232;
  assign \new_[55983]_  = ~A235 & ~A234;
  assign \new_[55984]_  = \new_[55983]_  & \new_[55980]_ ;
  assign \new_[55987]_  = ~A268 & ~A267;
  assign \new_[55990]_  = A301 & ~A269;
  assign \new_[55991]_  = \new_[55990]_  & \new_[55987]_ ;
  assign \new_[55992]_  = \new_[55991]_  & \new_[55984]_ ;
  assign \new_[55996]_  = A167 & ~A168;
  assign \new_[55997]_  = ~A169 & \new_[55996]_ ;
  assign \new_[56000]_  = A199 & A166;
  assign \new_[56003]_  = A203 & ~A200;
  assign \new_[56004]_  = \new_[56003]_  & \new_[56000]_ ;
  assign \new_[56005]_  = \new_[56004]_  & \new_[55997]_ ;
  assign \new_[56008]_  = A233 & A232;
  assign \new_[56011]_  = ~A235 & ~A234;
  assign \new_[56012]_  = \new_[56011]_  & \new_[56008]_ ;
  assign \new_[56015]_  = ~A266 & ~A265;
  assign \new_[56018]_  = A301 & ~A268;
  assign \new_[56019]_  = \new_[56018]_  & \new_[56015]_ ;
  assign \new_[56020]_  = \new_[56019]_  & \new_[56012]_ ;
  assign \new_[56024]_  = A167 & ~A168;
  assign \new_[56025]_  = ~A169 & \new_[56024]_ ;
  assign \new_[56028]_  = A199 & A166;
  assign \new_[56031]_  = A203 & ~A200;
  assign \new_[56032]_  = \new_[56031]_  & \new_[56028]_ ;
  assign \new_[56033]_  = \new_[56032]_  & \new_[56025]_ ;
  assign \new_[56036]_  = ~A233 & ~A232;
  assign \new_[56039]_  = ~A267 & ~A235;
  assign \new_[56040]_  = \new_[56039]_  & \new_[56036]_ ;
  assign \new_[56043]_  = ~A269 & ~A268;
  assign \new_[56046]_  = A300 & A299;
  assign \new_[56047]_  = \new_[56046]_  & \new_[56043]_ ;
  assign \new_[56048]_  = \new_[56047]_  & \new_[56040]_ ;
  assign \new_[56052]_  = A167 & ~A168;
  assign \new_[56053]_  = ~A169 & \new_[56052]_ ;
  assign \new_[56056]_  = A199 & A166;
  assign \new_[56059]_  = A203 & ~A200;
  assign \new_[56060]_  = \new_[56059]_  & \new_[56056]_ ;
  assign \new_[56061]_  = \new_[56060]_  & \new_[56053]_ ;
  assign \new_[56064]_  = ~A233 & ~A232;
  assign \new_[56067]_  = ~A267 & ~A235;
  assign \new_[56068]_  = \new_[56067]_  & \new_[56064]_ ;
  assign \new_[56071]_  = ~A269 & ~A268;
  assign \new_[56074]_  = A300 & A298;
  assign \new_[56075]_  = \new_[56074]_  & \new_[56071]_ ;
  assign \new_[56076]_  = \new_[56075]_  & \new_[56068]_ ;
  assign \new_[56080]_  = A167 & ~A168;
  assign \new_[56081]_  = ~A169 & \new_[56080]_ ;
  assign \new_[56084]_  = A199 & A166;
  assign \new_[56087]_  = A203 & ~A200;
  assign \new_[56088]_  = \new_[56087]_  & \new_[56084]_ ;
  assign \new_[56089]_  = \new_[56088]_  & \new_[56081]_ ;
  assign \new_[56092]_  = ~A233 & ~A232;
  assign \new_[56095]_  = A265 & ~A235;
  assign \new_[56096]_  = \new_[56095]_  & \new_[56092]_ ;
  assign \new_[56099]_  = ~A267 & A266;
  assign \new_[56102]_  = A301 & ~A268;
  assign \new_[56103]_  = \new_[56102]_  & \new_[56099]_ ;
  assign \new_[56104]_  = \new_[56103]_  & \new_[56096]_ ;
  assign \new_[56108]_  = A167 & ~A168;
  assign \new_[56109]_  = ~A169 & \new_[56108]_ ;
  assign \new_[56112]_  = A199 & A166;
  assign \new_[56115]_  = A203 & ~A200;
  assign \new_[56116]_  = \new_[56115]_  & \new_[56112]_ ;
  assign \new_[56117]_  = \new_[56116]_  & \new_[56109]_ ;
  assign \new_[56120]_  = ~A233 & ~A232;
  assign \new_[56123]_  = ~A265 & ~A235;
  assign \new_[56124]_  = \new_[56123]_  & \new_[56120]_ ;
  assign \new_[56127]_  = ~A268 & ~A266;
  assign \new_[56130]_  = A300 & A299;
  assign \new_[56131]_  = \new_[56130]_  & \new_[56127]_ ;
  assign \new_[56132]_  = \new_[56131]_  & \new_[56124]_ ;
  assign \new_[56136]_  = A167 & ~A168;
  assign \new_[56137]_  = ~A169 & \new_[56136]_ ;
  assign \new_[56140]_  = A199 & A166;
  assign \new_[56143]_  = A203 & ~A200;
  assign \new_[56144]_  = \new_[56143]_  & \new_[56140]_ ;
  assign \new_[56145]_  = \new_[56144]_  & \new_[56137]_ ;
  assign \new_[56148]_  = ~A233 & ~A232;
  assign \new_[56151]_  = ~A265 & ~A235;
  assign \new_[56152]_  = \new_[56151]_  & \new_[56148]_ ;
  assign \new_[56155]_  = ~A268 & ~A266;
  assign \new_[56158]_  = A300 & A298;
  assign \new_[56159]_  = \new_[56158]_  & \new_[56155]_ ;
  assign \new_[56160]_  = \new_[56159]_  & \new_[56152]_ ;
  assign \new_[56164]_  = ~A168 & ~A169;
  assign \new_[56165]_  = ~A170 & \new_[56164]_ ;
  assign \new_[56168]_  = A232 & A202;
  assign \new_[56171]_  = ~A234 & A233;
  assign \new_[56172]_  = \new_[56171]_  & \new_[56168]_ ;
  assign \new_[56173]_  = \new_[56172]_  & \new_[56165]_ ;
  assign \new_[56176]_  = A265 & ~A235;
  assign \new_[56179]_  = ~A267 & A266;
  assign \new_[56180]_  = \new_[56179]_  & \new_[56176]_ ;
  assign \new_[56183]_  = A298 & ~A268;
  assign \new_[56186]_  = A302 & ~A299;
  assign \new_[56187]_  = \new_[56186]_  & \new_[56183]_ ;
  assign \new_[56188]_  = \new_[56187]_  & \new_[56180]_ ;
  assign \new_[56192]_  = ~A168 & ~A169;
  assign \new_[56193]_  = ~A170 & \new_[56192]_ ;
  assign \new_[56196]_  = A232 & A202;
  assign \new_[56199]_  = ~A234 & A233;
  assign \new_[56200]_  = \new_[56199]_  & \new_[56196]_ ;
  assign \new_[56201]_  = \new_[56200]_  & \new_[56193]_ ;
  assign \new_[56204]_  = A265 & ~A235;
  assign \new_[56207]_  = ~A267 & A266;
  assign \new_[56208]_  = \new_[56207]_  & \new_[56204]_ ;
  assign \new_[56211]_  = ~A298 & ~A268;
  assign \new_[56214]_  = A302 & A299;
  assign \new_[56215]_  = \new_[56214]_  & \new_[56211]_ ;
  assign \new_[56216]_  = \new_[56215]_  & \new_[56208]_ ;
  assign \new_[56220]_  = ~A168 & ~A169;
  assign \new_[56221]_  = ~A170 & \new_[56220]_ ;
  assign \new_[56224]_  = A201 & A199;
  assign \new_[56227]_  = ~A235 & ~A234;
  assign \new_[56228]_  = \new_[56227]_  & \new_[56224]_ ;
  assign \new_[56229]_  = \new_[56228]_  & \new_[56221]_ ;
  assign \new_[56232]_  = A265 & ~A236;
  assign \new_[56235]_  = ~A267 & A266;
  assign \new_[56236]_  = \new_[56235]_  & \new_[56232]_ ;
  assign \new_[56239]_  = A298 & ~A268;
  assign \new_[56242]_  = A302 & ~A299;
  assign \new_[56243]_  = \new_[56242]_  & \new_[56239]_ ;
  assign \new_[56244]_  = \new_[56243]_  & \new_[56236]_ ;
  assign \new_[56248]_  = ~A168 & ~A169;
  assign \new_[56249]_  = ~A170 & \new_[56248]_ ;
  assign \new_[56252]_  = A201 & A199;
  assign \new_[56255]_  = ~A235 & ~A234;
  assign \new_[56256]_  = \new_[56255]_  & \new_[56252]_ ;
  assign \new_[56257]_  = \new_[56256]_  & \new_[56249]_ ;
  assign \new_[56260]_  = A265 & ~A236;
  assign \new_[56263]_  = ~A267 & A266;
  assign \new_[56264]_  = \new_[56263]_  & \new_[56260]_ ;
  assign \new_[56267]_  = ~A298 & ~A268;
  assign \new_[56270]_  = A302 & A299;
  assign \new_[56271]_  = \new_[56270]_  & \new_[56267]_ ;
  assign \new_[56272]_  = \new_[56271]_  & \new_[56264]_ ;
  assign \new_[56276]_  = ~A168 & ~A169;
  assign \new_[56277]_  = ~A170 & \new_[56276]_ ;
  assign \new_[56280]_  = A201 & A199;
  assign \new_[56283]_  = A233 & A232;
  assign \new_[56284]_  = \new_[56283]_  & \new_[56280]_ ;
  assign \new_[56285]_  = \new_[56284]_  & \new_[56277]_ ;
  assign \new_[56288]_  = ~A235 & ~A234;
  assign \new_[56291]_  = ~A268 & ~A267;
  assign \new_[56292]_  = \new_[56291]_  & \new_[56288]_ ;
  assign \new_[56295]_  = A298 & ~A269;
  assign \new_[56298]_  = A302 & ~A299;
  assign \new_[56299]_  = \new_[56298]_  & \new_[56295]_ ;
  assign \new_[56300]_  = \new_[56299]_  & \new_[56292]_ ;
  assign \new_[56304]_  = ~A168 & ~A169;
  assign \new_[56305]_  = ~A170 & \new_[56304]_ ;
  assign \new_[56308]_  = A201 & A199;
  assign \new_[56311]_  = A233 & A232;
  assign \new_[56312]_  = \new_[56311]_  & \new_[56308]_ ;
  assign \new_[56313]_  = \new_[56312]_  & \new_[56305]_ ;
  assign \new_[56316]_  = ~A235 & ~A234;
  assign \new_[56319]_  = ~A268 & ~A267;
  assign \new_[56320]_  = \new_[56319]_  & \new_[56316]_ ;
  assign \new_[56323]_  = ~A298 & ~A269;
  assign \new_[56326]_  = A302 & A299;
  assign \new_[56327]_  = \new_[56326]_  & \new_[56323]_ ;
  assign \new_[56328]_  = \new_[56327]_  & \new_[56320]_ ;
  assign \new_[56332]_  = ~A168 & ~A169;
  assign \new_[56333]_  = ~A170 & \new_[56332]_ ;
  assign \new_[56336]_  = A201 & A199;
  assign \new_[56339]_  = A233 & A232;
  assign \new_[56340]_  = \new_[56339]_  & \new_[56336]_ ;
  assign \new_[56341]_  = \new_[56340]_  & \new_[56333]_ ;
  assign \new_[56344]_  = ~A235 & ~A234;
  assign \new_[56347]_  = A266 & A265;
  assign \new_[56348]_  = \new_[56347]_  & \new_[56344]_ ;
  assign \new_[56351]_  = ~A268 & ~A267;
  assign \new_[56354]_  = A300 & A299;
  assign \new_[56355]_  = \new_[56354]_  & \new_[56351]_ ;
  assign \new_[56356]_  = \new_[56355]_  & \new_[56348]_ ;
  assign \new_[56360]_  = ~A168 & ~A169;
  assign \new_[56361]_  = ~A170 & \new_[56360]_ ;
  assign \new_[56364]_  = A201 & A199;
  assign \new_[56367]_  = A233 & A232;
  assign \new_[56368]_  = \new_[56367]_  & \new_[56364]_ ;
  assign \new_[56369]_  = \new_[56368]_  & \new_[56361]_ ;
  assign \new_[56372]_  = ~A235 & ~A234;
  assign \new_[56375]_  = A266 & A265;
  assign \new_[56376]_  = \new_[56375]_  & \new_[56372]_ ;
  assign \new_[56379]_  = ~A268 & ~A267;
  assign \new_[56382]_  = A300 & A298;
  assign \new_[56383]_  = \new_[56382]_  & \new_[56379]_ ;
  assign \new_[56384]_  = \new_[56383]_  & \new_[56376]_ ;
  assign \new_[56388]_  = ~A168 & ~A169;
  assign \new_[56389]_  = ~A170 & \new_[56388]_ ;
  assign \new_[56392]_  = A201 & A199;
  assign \new_[56395]_  = A233 & A232;
  assign \new_[56396]_  = \new_[56395]_  & \new_[56392]_ ;
  assign \new_[56397]_  = \new_[56396]_  & \new_[56389]_ ;
  assign \new_[56400]_  = ~A235 & ~A234;
  assign \new_[56403]_  = ~A266 & ~A265;
  assign \new_[56404]_  = \new_[56403]_  & \new_[56400]_ ;
  assign \new_[56407]_  = A298 & ~A268;
  assign \new_[56410]_  = A302 & ~A299;
  assign \new_[56411]_  = \new_[56410]_  & \new_[56407]_ ;
  assign \new_[56412]_  = \new_[56411]_  & \new_[56404]_ ;
  assign \new_[56416]_  = ~A168 & ~A169;
  assign \new_[56417]_  = ~A170 & \new_[56416]_ ;
  assign \new_[56420]_  = A201 & A199;
  assign \new_[56423]_  = A233 & A232;
  assign \new_[56424]_  = \new_[56423]_  & \new_[56420]_ ;
  assign \new_[56425]_  = \new_[56424]_  & \new_[56417]_ ;
  assign \new_[56428]_  = ~A235 & ~A234;
  assign \new_[56431]_  = ~A266 & ~A265;
  assign \new_[56432]_  = \new_[56431]_  & \new_[56428]_ ;
  assign \new_[56435]_  = ~A298 & ~A268;
  assign \new_[56438]_  = A302 & A299;
  assign \new_[56439]_  = \new_[56438]_  & \new_[56435]_ ;
  assign \new_[56440]_  = \new_[56439]_  & \new_[56432]_ ;
  assign \new_[56444]_  = ~A168 & ~A169;
  assign \new_[56445]_  = ~A170 & \new_[56444]_ ;
  assign \new_[56448]_  = A201 & A199;
  assign \new_[56451]_  = ~A233 & ~A232;
  assign \new_[56452]_  = \new_[56451]_  & \new_[56448]_ ;
  assign \new_[56453]_  = \new_[56452]_  & \new_[56445]_ ;
  assign \new_[56456]_  = A265 & ~A235;
  assign \new_[56459]_  = ~A267 & A266;
  assign \new_[56460]_  = \new_[56459]_  & \new_[56456]_ ;
  assign \new_[56463]_  = A298 & ~A268;
  assign \new_[56466]_  = A302 & ~A299;
  assign \new_[56467]_  = \new_[56466]_  & \new_[56463]_ ;
  assign \new_[56468]_  = \new_[56467]_  & \new_[56460]_ ;
  assign \new_[56472]_  = ~A168 & ~A169;
  assign \new_[56473]_  = ~A170 & \new_[56472]_ ;
  assign \new_[56476]_  = A201 & A199;
  assign \new_[56479]_  = ~A233 & ~A232;
  assign \new_[56480]_  = \new_[56479]_  & \new_[56476]_ ;
  assign \new_[56481]_  = \new_[56480]_  & \new_[56473]_ ;
  assign \new_[56484]_  = A265 & ~A235;
  assign \new_[56487]_  = ~A267 & A266;
  assign \new_[56488]_  = \new_[56487]_  & \new_[56484]_ ;
  assign \new_[56491]_  = ~A298 & ~A268;
  assign \new_[56494]_  = A302 & A299;
  assign \new_[56495]_  = \new_[56494]_  & \new_[56491]_ ;
  assign \new_[56496]_  = \new_[56495]_  & \new_[56488]_ ;
  assign \new_[56500]_  = ~A168 & ~A169;
  assign \new_[56501]_  = ~A170 & \new_[56500]_ ;
  assign \new_[56504]_  = A201 & A200;
  assign \new_[56507]_  = ~A235 & ~A234;
  assign \new_[56508]_  = \new_[56507]_  & \new_[56504]_ ;
  assign \new_[56509]_  = \new_[56508]_  & \new_[56501]_ ;
  assign \new_[56512]_  = A265 & ~A236;
  assign \new_[56515]_  = ~A267 & A266;
  assign \new_[56516]_  = \new_[56515]_  & \new_[56512]_ ;
  assign \new_[56519]_  = A298 & ~A268;
  assign \new_[56522]_  = A302 & ~A299;
  assign \new_[56523]_  = \new_[56522]_  & \new_[56519]_ ;
  assign \new_[56524]_  = \new_[56523]_  & \new_[56516]_ ;
  assign \new_[56528]_  = ~A168 & ~A169;
  assign \new_[56529]_  = ~A170 & \new_[56528]_ ;
  assign \new_[56532]_  = A201 & A200;
  assign \new_[56535]_  = ~A235 & ~A234;
  assign \new_[56536]_  = \new_[56535]_  & \new_[56532]_ ;
  assign \new_[56537]_  = \new_[56536]_  & \new_[56529]_ ;
  assign \new_[56540]_  = A265 & ~A236;
  assign \new_[56543]_  = ~A267 & A266;
  assign \new_[56544]_  = \new_[56543]_  & \new_[56540]_ ;
  assign \new_[56547]_  = ~A298 & ~A268;
  assign \new_[56550]_  = A302 & A299;
  assign \new_[56551]_  = \new_[56550]_  & \new_[56547]_ ;
  assign \new_[56552]_  = \new_[56551]_  & \new_[56544]_ ;
  assign \new_[56556]_  = ~A168 & ~A169;
  assign \new_[56557]_  = ~A170 & \new_[56556]_ ;
  assign \new_[56560]_  = A201 & A200;
  assign \new_[56563]_  = A233 & A232;
  assign \new_[56564]_  = \new_[56563]_  & \new_[56560]_ ;
  assign \new_[56565]_  = \new_[56564]_  & \new_[56557]_ ;
  assign \new_[56568]_  = ~A235 & ~A234;
  assign \new_[56571]_  = ~A268 & ~A267;
  assign \new_[56572]_  = \new_[56571]_  & \new_[56568]_ ;
  assign \new_[56575]_  = A298 & ~A269;
  assign \new_[56578]_  = A302 & ~A299;
  assign \new_[56579]_  = \new_[56578]_  & \new_[56575]_ ;
  assign \new_[56580]_  = \new_[56579]_  & \new_[56572]_ ;
  assign \new_[56584]_  = ~A168 & ~A169;
  assign \new_[56585]_  = ~A170 & \new_[56584]_ ;
  assign \new_[56588]_  = A201 & A200;
  assign \new_[56591]_  = A233 & A232;
  assign \new_[56592]_  = \new_[56591]_  & \new_[56588]_ ;
  assign \new_[56593]_  = \new_[56592]_  & \new_[56585]_ ;
  assign \new_[56596]_  = ~A235 & ~A234;
  assign \new_[56599]_  = ~A268 & ~A267;
  assign \new_[56600]_  = \new_[56599]_  & \new_[56596]_ ;
  assign \new_[56603]_  = ~A298 & ~A269;
  assign \new_[56606]_  = A302 & A299;
  assign \new_[56607]_  = \new_[56606]_  & \new_[56603]_ ;
  assign \new_[56608]_  = \new_[56607]_  & \new_[56600]_ ;
  assign \new_[56612]_  = ~A168 & ~A169;
  assign \new_[56613]_  = ~A170 & \new_[56612]_ ;
  assign \new_[56616]_  = A201 & A200;
  assign \new_[56619]_  = A233 & A232;
  assign \new_[56620]_  = \new_[56619]_  & \new_[56616]_ ;
  assign \new_[56621]_  = \new_[56620]_  & \new_[56613]_ ;
  assign \new_[56624]_  = ~A235 & ~A234;
  assign \new_[56627]_  = A266 & A265;
  assign \new_[56628]_  = \new_[56627]_  & \new_[56624]_ ;
  assign \new_[56631]_  = ~A268 & ~A267;
  assign \new_[56634]_  = A300 & A299;
  assign \new_[56635]_  = \new_[56634]_  & \new_[56631]_ ;
  assign \new_[56636]_  = \new_[56635]_  & \new_[56628]_ ;
  assign \new_[56640]_  = ~A168 & ~A169;
  assign \new_[56641]_  = ~A170 & \new_[56640]_ ;
  assign \new_[56644]_  = A201 & A200;
  assign \new_[56647]_  = A233 & A232;
  assign \new_[56648]_  = \new_[56647]_  & \new_[56644]_ ;
  assign \new_[56649]_  = \new_[56648]_  & \new_[56641]_ ;
  assign \new_[56652]_  = ~A235 & ~A234;
  assign \new_[56655]_  = A266 & A265;
  assign \new_[56656]_  = \new_[56655]_  & \new_[56652]_ ;
  assign \new_[56659]_  = ~A268 & ~A267;
  assign \new_[56662]_  = A300 & A298;
  assign \new_[56663]_  = \new_[56662]_  & \new_[56659]_ ;
  assign \new_[56664]_  = \new_[56663]_  & \new_[56656]_ ;
  assign \new_[56668]_  = ~A168 & ~A169;
  assign \new_[56669]_  = ~A170 & \new_[56668]_ ;
  assign \new_[56672]_  = A201 & A200;
  assign \new_[56675]_  = A233 & A232;
  assign \new_[56676]_  = \new_[56675]_  & \new_[56672]_ ;
  assign \new_[56677]_  = \new_[56676]_  & \new_[56669]_ ;
  assign \new_[56680]_  = ~A235 & ~A234;
  assign \new_[56683]_  = ~A266 & ~A265;
  assign \new_[56684]_  = \new_[56683]_  & \new_[56680]_ ;
  assign \new_[56687]_  = A298 & ~A268;
  assign \new_[56690]_  = A302 & ~A299;
  assign \new_[56691]_  = \new_[56690]_  & \new_[56687]_ ;
  assign \new_[56692]_  = \new_[56691]_  & \new_[56684]_ ;
  assign \new_[56696]_  = ~A168 & ~A169;
  assign \new_[56697]_  = ~A170 & \new_[56696]_ ;
  assign \new_[56700]_  = A201 & A200;
  assign \new_[56703]_  = A233 & A232;
  assign \new_[56704]_  = \new_[56703]_  & \new_[56700]_ ;
  assign \new_[56705]_  = \new_[56704]_  & \new_[56697]_ ;
  assign \new_[56708]_  = ~A235 & ~A234;
  assign \new_[56711]_  = ~A266 & ~A265;
  assign \new_[56712]_  = \new_[56711]_  & \new_[56708]_ ;
  assign \new_[56715]_  = ~A298 & ~A268;
  assign \new_[56718]_  = A302 & A299;
  assign \new_[56719]_  = \new_[56718]_  & \new_[56715]_ ;
  assign \new_[56720]_  = \new_[56719]_  & \new_[56712]_ ;
  assign \new_[56724]_  = ~A168 & ~A169;
  assign \new_[56725]_  = ~A170 & \new_[56724]_ ;
  assign \new_[56728]_  = A201 & A200;
  assign \new_[56731]_  = ~A233 & ~A232;
  assign \new_[56732]_  = \new_[56731]_  & \new_[56728]_ ;
  assign \new_[56733]_  = \new_[56732]_  & \new_[56725]_ ;
  assign \new_[56736]_  = A265 & ~A235;
  assign \new_[56739]_  = ~A267 & A266;
  assign \new_[56740]_  = \new_[56739]_  & \new_[56736]_ ;
  assign \new_[56743]_  = A298 & ~A268;
  assign \new_[56746]_  = A302 & ~A299;
  assign \new_[56747]_  = \new_[56746]_  & \new_[56743]_ ;
  assign \new_[56748]_  = \new_[56747]_  & \new_[56740]_ ;
  assign \new_[56752]_  = ~A168 & ~A169;
  assign \new_[56753]_  = ~A170 & \new_[56752]_ ;
  assign \new_[56756]_  = A201 & A200;
  assign \new_[56759]_  = ~A233 & ~A232;
  assign \new_[56760]_  = \new_[56759]_  & \new_[56756]_ ;
  assign \new_[56761]_  = \new_[56760]_  & \new_[56753]_ ;
  assign \new_[56764]_  = A265 & ~A235;
  assign \new_[56767]_  = ~A267 & A266;
  assign \new_[56768]_  = \new_[56767]_  & \new_[56764]_ ;
  assign \new_[56771]_  = ~A298 & ~A268;
  assign \new_[56774]_  = A302 & A299;
  assign \new_[56775]_  = \new_[56774]_  & \new_[56771]_ ;
  assign \new_[56776]_  = \new_[56775]_  & \new_[56768]_ ;
  assign \new_[56780]_  = ~A168 & ~A169;
  assign \new_[56781]_  = ~A170 & \new_[56780]_ ;
  assign \new_[56784]_  = A200 & ~A199;
  assign \new_[56787]_  = ~A234 & A203;
  assign \new_[56788]_  = \new_[56787]_  & \new_[56784]_ ;
  assign \new_[56789]_  = \new_[56788]_  & \new_[56781]_ ;
  assign \new_[56792]_  = ~A236 & ~A235;
  assign \new_[56795]_  = ~A268 & ~A267;
  assign \new_[56796]_  = \new_[56795]_  & \new_[56792]_ ;
  assign \new_[56799]_  = A298 & ~A269;
  assign \new_[56802]_  = A302 & ~A299;
  assign \new_[56803]_  = \new_[56802]_  & \new_[56799]_ ;
  assign \new_[56804]_  = \new_[56803]_  & \new_[56796]_ ;
  assign \new_[56808]_  = ~A168 & ~A169;
  assign \new_[56809]_  = ~A170 & \new_[56808]_ ;
  assign \new_[56812]_  = A200 & ~A199;
  assign \new_[56815]_  = ~A234 & A203;
  assign \new_[56816]_  = \new_[56815]_  & \new_[56812]_ ;
  assign \new_[56817]_  = \new_[56816]_  & \new_[56809]_ ;
  assign \new_[56820]_  = ~A236 & ~A235;
  assign \new_[56823]_  = ~A268 & ~A267;
  assign \new_[56824]_  = \new_[56823]_  & \new_[56820]_ ;
  assign \new_[56827]_  = ~A298 & ~A269;
  assign \new_[56830]_  = A302 & A299;
  assign \new_[56831]_  = \new_[56830]_  & \new_[56827]_ ;
  assign \new_[56832]_  = \new_[56831]_  & \new_[56824]_ ;
  assign \new_[56836]_  = ~A168 & ~A169;
  assign \new_[56837]_  = ~A170 & \new_[56836]_ ;
  assign \new_[56840]_  = A200 & ~A199;
  assign \new_[56843]_  = ~A234 & A203;
  assign \new_[56844]_  = \new_[56843]_  & \new_[56840]_ ;
  assign \new_[56845]_  = \new_[56844]_  & \new_[56837]_ ;
  assign \new_[56848]_  = ~A236 & ~A235;
  assign \new_[56851]_  = A266 & A265;
  assign \new_[56852]_  = \new_[56851]_  & \new_[56848]_ ;
  assign \new_[56855]_  = ~A268 & ~A267;
  assign \new_[56858]_  = A300 & A299;
  assign \new_[56859]_  = \new_[56858]_  & \new_[56855]_ ;
  assign \new_[56860]_  = \new_[56859]_  & \new_[56852]_ ;
  assign \new_[56864]_  = ~A168 & ~A169;
  assign \new_[56865]_  = ~A170 & \new_[56864]_ ;
  assign \new_[56868]_  = A200 & ~A199;
  assign \new_[56871]_  = ~A234 & A203;
  assign \new_[56872]_  = \new_[56871]_  & \new_[56868]_ ;
  assign \new_[56873]_  = \new_[56872]_  & \new_[56865]_ ;
  assign \new_[56876]_  = ~A236 & ~A235;
  assign \new_[56879]_  = A266 & A265;
  assign \new_[56880]_  = \new_[56879]_  & \new_[56876]_ ;
  assign \new_[56883]_  = ~A268 & ~A267;
  assign \new_[56886]_  = A300 & A298;
  assign \new_[56887]_  = \new_[56886]_  & \new_[56883]_ ;
  assign \new_[56888]_  = \new_[56887]_  & \new_[56880]_ ;
  assign \new_[56892]_  = ~A168 & ~A169;
  assign \new_[56893]_  = ~A170 & \new_[56892]_ ;
  assign \new_[56896]_  = A200 & ~A199;
  assign \new_[56899]_  = ~A234 & A203;
  assign \new_[56900]_  = \new_[56899]_  & \new_[56896]_ ;
  assign \new_[56901]_  = \new_[56900]_  & \new_[56893]_ ;
  assign \new_[56904]_  = ~A236 & ~A235;
  assign \new_[56907]_  = ~A266 & ~A265;
  assign \new_[56908]_  = \new_[56907]_  & \new_[56904]_ ;
  assign \new_[56911]_  = A298 & ~A268;
  assign \new_[56914]_  = A302 & ~A299;
  assign \new_[56915]_  = \new_[56914]_  & \new_[56911]_ ;
  assign \new_[56916]_  = \new_[56915]_  & \new_[56908]_ ;
  assign \new_[56920]_  = ~A168 & ~A169;
  assign \new_[56921]_  = ~A170 & \new_[56920]_ ;
  assign \new_[56924]_  = A200 & ~A199;
  assign \new_[56927]_  = ~A234 & A203;
  assign \new_[56928]_  = \new_[56927]_  & \new_[56924]_ ;
  assign \new_[56929]_  = \new_[56928]_  & \new_[56921]_ ;
  assign \new_[56932]_  = ~A236 & ~A235;
  assign \new_[56935]_  = ~A266 & ~A265;
  assign \new_[56936]_  = \new_[56935]_  & \new_[56932]_ ;
  assign \new_[56939]_  = ~A298 & ~A268;
  assign \new_[56942]_  = A302 & A299;
  assign \new_[56943]_  = \new_[56942]_  & \new_[56939]_ ;
  assign \new_[56944]_  = \new_[56943]_  & \new_[56936]_ ;
  assign \new_[56948]_  = ~A168 & ~A169;
  assign \new_[56949]_  = ~A170 & \new_[56948]_ ;
  assign \new_[56952]_  = A200 & ~A199;
  assign \new_[56955]_  = A232 & A203;
  assign \new_[56956]_  = \new_[56955]_  & \new_[56952]_ ;
  assign \new_[56957]_  = \new_[56956]_  & \new_[56949]_ ;
  assign \new_[56960]_  = ~A234 & A233;
  assign \new_[56963]_  = ~A267 & ~A235;
  assign \new_[56964]_  = \new_[56963]_  & \new_[56960]_ ;
  assign \new_[56967]_  = ~A269 & ~A268;
  assign \new_[56970]_  = A300 & A299;
  assign \new_[56971]_  = \new_[56970]_  & \new_[56967]_ ;
  assign \new_[56972]_  = \new_[56971]_  & \new_[56964]_ ;
  assign \new_[56976]_  = ~A168 & ~A169;
  assign \new_[56977]_  = ~A170 & \new_[56976]_ ;
  assign \new_[56980]_  = A200 & ~A199;
  assign \new_[56983]_  = A232 & A203;
  assign \new_[56984]_  = \new_[56983]_  & \new_[56980]_ ;
  assign \new_[56985]_  = \new_[56984]_  & \new_[56977]_ ;
  assign \new_[56988]_  = ~A234 & A233;
  assign \new_[56991]_  = ~A267 & ~A235;
  assign \new_[56992]_  = \new_[56991]_  & \new_[56988]_ ;
  assign \new_[56995]_  = ~A269 & ~A268;
  assign \new_[56998]_  = A300 & A298;
  assign \new_[56999]_  = \new_[56998]_  & \new_[56995]_ ;
  assign \new_[57000]_  = \new_[56999]_  & \new_[56992]_ ;
  assign \new_[57004]_  = ~A168 & ~A169;
  assign \new_[57005]_  = ~A170 & \new_[57004]_ ;
  assign \new_[57008]_  = A200 & ~A199;
  assign \new_[57011]_  = A232 & A203;
  assign \new_[57012]_  = \new_[57011]_  & \new_[57008]_ ;
  assign \new_[57013]_  = \new_[57012]_  & \new_[57005]_ ;
  assign \new_[57016]_  = ~A234 & A233;
  assign \new_[57019]_  = A265 & ~A235;
  assign \new_[57020]_  = \new_[57019]_  & \new_[57016]_ ;
  assign \new_[57023]_  = ~A267 & A266;
  assign \new_[57026]_  = A301 & ~A268;
  assign \new_[57027]_  = \new_[57026]_  & \new_[57023]_ ;
  assign \new_[57028]_  = \new_[57027]_  & \new_[57020]_ ;
  assign \new_[57032]_  = ~A168 & ~A169;
  assign \new_[57033]_  = ~A170 & \new_[57032]_ ;
  assign \new_[57036]_  = A200 & ~A199;
  assign \new_[57039]_  = A232 & A203;
  assign \new_[57040]_  = \new_[57039]_  & \new_[57036]_ ;
  assign \new_[57041]_  = \new_[57040]_  & \new_[57033]_ ;
  assign \new_[57044]_  = ~A234 & A233;
  assign \new_[57047]_  = ~A265 & ~A235;
  assign \new_[57048]_  = \new_[57047]_  & \new_[57044]_ ;
  assign \new_[57051]_  = ~A268 & ~A266;
  assign \new_[57054]_  = A300 & A299;
  assign \new_[57055]_  = \new_[57054]_  & \new_[57051]_ ;
  assign \new_[57056]_  = \new_[57055]_  & \new_[57048]_ ;
  assign \new_[57060]_  = ~A168 & ~A169;
  assign \new_[57061]_  = ~A170 & \new_[57060]_ ;
  assign \new_[57064]_  = A200 & ~A199;
  assign \new_[57067]_  = A232 & A203;
  assign \new_[57068]_  = \new_[57067]_  & \new_[57064]_ ;
  assign \new_[57069]_  = \new_[57068]_  & \new_[57061]_ ;
  assign \new_[57072]_  = ~A234 & A233;
  assign \new_[57075]_  = ~A265 & ~A235;
  assign \new_[57076]_  = \new_[57075]_  & \new_[57072]_ ;
  assign \new_[57079]_  = ~A268 & ~A266;
  assign \new_[57082]_  = A300 & A298;
  assign \new_[57083]_  = \new_[57082]_  & \new_[57079]_ ;
  assign \new_[57084]_  = \new_[57083]_  & \new_[57076]_ ;
  assign \new_[57088]_  = ~A168 & ~A169;
  assign \new_[57089]_  = ~A170 & \new_[57088]_ ;
  assign \new_[57092]_  = A200 & ~A199;
  assign \new_[57095]_  = ~A232 & A203;
  assign \new_[57096]_  = \new_[57095]_  & \new_[57092]_ ;
  assign \new_[57097]_  = \new_[57096]_  & \new_[57089]_ ;
  assign \new_[57100]_  = ~A235 & ~A233;
  assign \new_[57103]_  = ~A268 & ~A267;
  assign \new_[57104]_  = \new_[57103]_  & \new_[57100]_ ;
  assign \new_[57107]_  = A298 & ~A269;
  assign \new_[57110]_  = A302 & ~A299;
  assign \new_[57111]_  = \new_[57110]_  & \new_[57107]_ ;
  assign \new_[57112]_  = \new_[57111]_  & \new_[57104]_ ;
  assign \new_[57116]_  = ~A168 & ~A169;
  assign \new_[57117]_  = ~A170 & \new_[57116]_ ;
  assign \new_[57120]_  = A200 & ~A199;
  assign \new_[57123]_  = ~A232 & A203;
  assign \new_[57124]_  = \new_[57123]_  & \new_[57120]_ ;
  assign \new_[57125]_  = \new_[57124]_  & \new_[57117]_ ;
  assign \new_[57128]_  = ~A235 & ~A233;
  assign \new_[57131]_  = ~A268 & ~A267;
  assign \new_[57132]_  = \new_[57131]_  & \new_[57128]_ ;
  assign \new_[57135]_  = ~A298 & ~A269;
  assign \new_[57138]_  = A302 & A299;
  assign \new_[57139]_  = \new_[57138]_  & \new_[57135]_ ;
  assign \new_[57140]_  = \new_[57139]_  & \new_[57132]_ ;
  assign \new_[57144]_  = ~A168 & ~A169;
  assign \new_[57145]_  = ~A170 & \new_[57144]_ ;
  assign \new_[57148]_  = A200 & ~A199;
  assign \new_[57151]_  = ~A232 & A203;
  assign \new_[57152]_  = \new_[57151]_  & \new_[57148]_ ;
  assign \new_[57153]_  = \new_[57152]_  & \new_[57145]_ ;
  assign \new_[57156]_  = ~A235 & ~A233;
  assign \new_[57159]_  = A266 & A265;
  assign \new_[57160]_  = \new_[57159]_  & \new_[57156]_ ;
  assign \new_[57163]_  = ~A268 & ~A267;
  assign \new_[57166]_  = A300 & A299;
  assign \new_[57167]_  = \new_[57166]_  & \new_[57163]_ ;
  assign \new_[57168]_  = \new_[57167]_  & \new_[57160]_ ;
  assign \new_[57172]_  = ~A168 & ~A169;
  assign \new_[57173]_  = ~A170 & \new_[57172]_ ;
  assign \new_[57176]_  = A200 & ~A199;
  assign \new_[57179]_  = ~A232 & A203;
  assign \new_[57180]_  = \new_[57179]_  & \new_[57176]_ ;
  assign \new_[57181]_  = \new_[57180]_  & \new_[57173]_ ;
  assign \new_[57184]_  = ~A235 & ~A233;
  assign \new_[57187]_  = A266 & A265;
  assign \new_[57188]_  = \new_[57187]_  & \new_[57184]_ ;
  assign \new_[57191]_  = ~A268 & ~A267;
  assign \new_[57194]_  = A300 & A298;
  assign \new_[57195]_  = \new_[57194]_  & \new_[57191]_ ;
  assign \new_[57196]_  = \new_[57195]_  & \new_[57188]_ ;
  assign \new_[57200]_  = ~A168 & ~A169;
  assign \new_[57201]_  = ~A170 & \new_[57200]_ ;
  assign \new_[57204]_  = A200 & ~A199;
  assign \new_[57207]_  = ~A232 & A203;
  assign \new_[57208]_  = \new_[57207]_  & \new_[57204]_ ;
  assign \new_[57209]_  = \new_[57208]_  & \new_[57201]_ ;
  assign \new_[57212]_  = ~A235 & ~A233;
  assign \new_[57215]_  = ~A266 & ~A265;
  assign \new_[57216]_  = \new_[57215]_  & \new_[57212]_ ;
  assign \new_[57219]_  = A298 & ~A268;
  assign \new_[57222]_  = A302 & ~A299;
  assign \new_[57223]_  = \new_[57222]_  & \new_[57219]_ ;
  assign \new_[57224]_  = \new_[57223]_  & \new_[57216]_ ;
  assign \new_[57228]_  = ~A168 & ~A169;
  assign \new_[57229]_  = ~A170 & \new_[57228]_ ;
  assign \new_[57232]_  = A200 & ~A199;
  assign \new_[57235]_  = ~A232 & A203;
  assign \new_[57236]_  = \new_[57235]_  & \new_[57232]_ ;
  assign \new_[57237]_  = \new_[57236]_  & \new_[57229]_ ;
  assign \new_[57240]_  = ~A235 & ~A233;
  assign \new_[57243]_  = ~A266 & ~A265;
  assign \new_[57244]_  = \new_[57243]_  & \new_[57240]_ ;
  assign \new_[57247]_  = ~A298 & ~A268;
  assign \new_[57250]_  = A302 & A299;
  assign \new_[57251]_  = \new_[57250]_  & \new_[57247]_ ;
  assign \new_[57252]_  = \new_[57251]_  & \new_[57244]_ ;
  assign \new_[57256]_  = ~A168 & ~A169;
  assign \new_[57257]_  = ~A170 & \new_[57256]_ ;
  assign \new_[57260]_  = ~A200 & A199;
  assign \new_[57263]_  = ~A234 & A203;
  assign \new_[57264]_  = \new_[57263]_  & \new_[57260]_ ;
  assign \new_[57265]_  = \new_[57264]_  & \new_[57257]_ ;
  assign \new_[57268]_  = ~A236 & ~A235;
  assign \new_[57271]_  = ~A268 & ~A267;
  assign \new_[57272]_  = \new_[57271]_  & \new_[57268]_ ;
  assign \new_[57275]_  = A298 & ~A269;
  assign \new_[57278]_  = A302 & ~A299;
  assign \new_[57279]_  = \new_[57278]_  & \new_[57275]_ ;
  assign \new_[57280]_  = \new_[57279]_  & \new_[57272]_ ;
  assign \new_[57284]_  = ~A168 & ~A169;
  assign \new_[57285]_  = ~A170 & \new_[57284]_ ;
  assign \new_[57288]_  = ~A200 & A199;
  assign \new_[57291]_  = ~A234 & A203;
  assign \new_[57292]_  = \new_[57291]_  & \new_[57288]_ ;
  assign \new_[57293]_  = \new_[57292]_  & \new_[57285]_ ;
  assign \new_[57296]_  = ~A236 & ~A235;
  assign \new_[57299]_  = ~A268 & ~A267;
  assign \new_[57300]_  = \new_[57299]_  & \new_[57296]_ ;
  assign \new_[57303]_  = ~A298 & ~A269;
  assign \new_[57306]_  = A302 & A299;
  assign \new_[57307]_  = \new_[57306]_  & \new_[57303]_ ;
  assign \new_[57308]_  = \new_[57307]_  & \new_[57300]_ ;
  assign \new_[57312]_  = ~A168 & ~A169;
  assign \new_[57313]_  = ~A170 & \new_[57312]_ ;
  assign \new_[57316]_  = ~A200 & A199;
  assign \new_[57319]_  = ~A234 & A203;
  assign \new_[57320]_  = \new_[57319]_  & \new_[57316]_ ;
  assign \new_[57321]_  = \new_[57320]_  & \new_[57313]_ ;
  assign \new_[57324]_  = ~A236 & ~A235;
  assign \new_[57327]_  = A266 & A265;
  assign \new_[57328]_  = \new_[57327]_  & \new_[57324]_ ;
  assign \new_[57331]_  = ~A268 & ~A267;
  assign \new_[57334]_  = A300 & A299;
  assign \new_[57335]_  = \new_[57334]_  & \new_[57331]_ ;
  assign \new_[57336]_  = \new_[57335]_  & \new_[57328]_ ;
  assign \new_[57340]_  = ~A168 & ~A169;
  assign \new_[57341]_  = ~A170 & \new_[57340]_ ;
  assign \new_[57344]_  = ~A200 & A199;
  assign \new_[57347]_  = ~A234 & A203;
  assign \new_[57348]_  = \new_[57347]_  & \new_[57344]_ ;
  assign \new_[57349]_  = \new_[57348]_  & \new_[57341]_ ;
  assign \new_[57352]_  = ~A236 & ~A235;
  assign \new_[57355]_  = A266 & A265;
  assign \new_[57356]_  = \new_[57355]_  & \new_[57352]_ ;
  assign \new_[57359]_  = ~A268 & ~A267;
  assign \new_[57362]_  = A300 & A298;
  assign \new_[57363]_  = \new_[57362]_  & \new_[57359]_ ;
  assign \new_[57364]_  = \new_[57363]_  & \new_[57356]_ ;
  assign \new_[57368]_  = ~A168 & ~A169;
  assign \new_[57369]_  = ~A170 & \new_[57368]_ ;
  assign \new_[57372]_  = ~A200 & A199;
  assign \new_[57375]_  = ~A234 & A203;
  assign \new_[57376]_  = \new_[57375]_  & \new_[57372]_ ;
  assign \new_[57377]_  = \new_[57376]_  & \new_[57369]_ ;
  assign \new_[57380]_  = ~A236 & ~A235;
  assign \new_[57383]_  = ~A266 & ~A265;
  assign \new_[57384]_  = \new_[57383]_  & \new_[57380]_ ;
  assign \new_[57387]_  = A298 & ~A268;
  assign \new_[57390]_  = A302 & ~A299;
  assign \new_[57391]_  = \new_[57390]_  & \new_[57387]_ ;
  assign \new_[57392]_  = \new_[57391]_  & \new_[57384]_ ;
  assign \new_[57396]_  = ~A168 & ~A169;
  assign \new_[57397]_  = ~A170 & \new_[57396]_ ;
  assign \new_[57400]_  = ~A200 & A199;
  assign \new_[57403]_  = ~A234 & A203;
  assign \new_[57404]_  = \new_[57403]_  & \new_[57400]_ ;
  assign \new_[57405]_  = \new_[57404]_  & \new_[57397]_ ;
  assign \new_[57408]_  = ~A236 & ~A235;
  assign \new_[57411]_  = ~A266 & ~A265;
  assign \new_[57412]_  = \new_[57411]_  & \new_[57408]_ ;
  assign \new_[57415]_  = ~A298 & ~A268;
  assign \new_[57418]_  = A302 & A299;
  assign \new_[57419]_  = \new_[57418]_  & \new_[57415]_ ;
  assign \new_[57420]_  = \new_[57419]_  & \new_[57412]_ ;
  assign \new_[57424]_  = ~A168 & ~A169;
  assign \new_[57425]_  = ~A170 & \new_[57424]_ ;
  assign \new_[57428]_  = ~A200 & A199;
  assign \new_[57431]_  = A232 & A203;
  assign \new_[57432]_  = \new_[57431]_  & \new_[57428]_ ;
  assign \new_[57433]_  = \new_[57432]_  & \new_[57425]_ ;
  assign \new_[57436]_  = ~A234 & A233;
  assign \new_[57439]_  = ~A267 & ~A235;
  assign \new_[57440]_  = \new_[57439]_  & \new_[57436]_ ;
  assign \new_[57443]_  = ~A269 & ~A268;
  assign \new_[57446]_  = A300 & A299;
  assign \new_[57447]_  = \new_[57446]_  & \new_[57443]_ ;
  assign \new_[57448]_  = \new_[57447]_  & \new_[57440]_ ;
  assign \new_[57452]_  = ~A168 & ~A169;
  assign \new_[57453]_  = ~A170 & \new_[57452]_ ;
  assign \new_[57456]_  = ~A200 & A199;
  assign \new_[57459]_  = A232 & A203;
  assign \new_[57460]_  = \new_[57459]_  & \new_[57456]_ ;
  assign \new_[57461]_  = \new_[57460]_  & \new_[57453]_ ;
  assign \new_[57464]_  = ~A234 & A233;
  assign \new_[57467]_  = ~A267 & ~A235;
  assign \new_[57468]_  = \new_[57467]_  & \new_[57464]_ ;
  assign \new_[57471]_  = ~A269 & ~A268;
  assign \new_[57474]_  = A300 & A298;
  assign \new_[57475]_  = \new_[57474]_  & \new_[57471]_ ;
  assign \new_[57476]_  = \new_[57475]_  & \new_[57468]_ ;
  assign \new_[57480]_  = ~A168 & ~A169;
  assign \new_[57481]_  = ~A170 & \new_[57480]_ ;
  assign \new_[57484]_  = ~A200 & A199;
  assign \new_[57487]_  = A232 & A203;
  assign \new_[57488]_  = \new_[57487]_  & \new_[57484]_ ;
  assign \new_[57489]_  = \new_[57488]_  & \new_[57481]_ ;
  assign \new_[57492]_  = ~A234 & A233;
  assign \new_[57495]_  = A265 & ~A235;
  assign \new_[57496]_  = \new_[57495]_  & \new_[57492]_ ;
  assign \new_[57499]_  = ~A267 & A266;
  assign \new_[57502]_  = A301 & ~A268;
  assign \new_[57503]_  = \new_[57502]_  & \new_[57499]_ ;
  assign \new_[57504]_  = \new_[57503]_  & \new_[57496]_ ;
  assign \new_[57508]_  = ~A168 & ~A169;
  assign \new_[57509]_  = ~A170 & \new_[57508]_ ;
  assign \new_[57512]_  = ~A200 & A199;
  assign \new_[57515]_  = A232 & A203;
  assign \new_[57516]_  = \new_[57515]_  & \new_[57512]_ ;
  assign \new_[57517]_  = \new_[57516]_  & \new_[57509]_ ;
  assign \new_[57520]_  = ~A234 & A233;
  assign \new_[57523]_  = ~A265 & ~A235;
  assign \new_[57524]_  = \new_[57523]_  & \new_[57520]_ ;
  assign \new_[57527]_  = ~A268 & ~A266;
  assign \new_[57530]_  = A300 & A299;
  assign \new_[57531]_  = \new_[57530]_  & \new_[57527]_ ;
  assign \new_[57532]_  = \new_[57531]_  & \new_[57524]_ ;
  assign \new_[57536]_  = ~A168 & ~A169;
  assign \new_[57537]_  = ~A170 & \new_[57536]_ ;
  assign \new_[57540]_  = ~A200 & A199;
  assign \new_[57543]_  = A232 & A203;
  assign \new_[57544]_  = \new_[57543]_  & \new_[57540]_ ;
  assign \new_[57545]_  = \new_[57544]_  & \new_[57537]_ ;
  assign \new_[57548]_  = ~A234 & A233;
  assign \new_[57551]_  = ~A265 & ~A235;
  assign \new_[57552]_  = \new_[57551]_  & \new_[57548]_ ;
  assign \new_[57555]_  = ~A268 & ~A266;
  assign \new_[57558]_  = A300 & A298;
  assign \new_[57559]_  = \new_[57558]_  & \new_[57555]_ ;
  assign \new_[57560]_  = \new_[57559]_  & \new_[57552]_ ;
  assign \new_[57564]_  = ~A168 & ~A169;
  assign \new_[57565]_  = ~A170 & \new_[57564]_ ;
  assign \new_[57568]_  = ~A200 & A199;
  assign \new_[57571]_  = ~A232 & A203;
  assign \new_[57572]_  = \new_[57571]_  & \new_[57568]_ ;
  assign \new_[57573]_  = \new_[57572]_  & \new_[57565]_ ;
  assign \new_[57576]_  = ~A235 & ~A233;
  assign \new_[57579]_  = ~A268 & ~A267;
  assign \new_[57580]_  = \new_[57579]_  & \new_[57576]_ ;
  assign \new_[57583]_  = A298 & ~A269;
  assign \new_[57586]_  = A302 & ~A299;
  assign \new_[57587]_  = \new_[57586]_  & \new_[57583]_ ;
  assign \new_[57588]_  = \new_[57587]_  & \new_[57580]_ ;
  assign \new_[57592]_  = ~A168 & ~A169;
  assign \new_[57593]_  = ~A170 & \new_[57592]_ ;
  assign \new_[57596]_  = ~A200 & A199;
  assign \new_[57599]_  = ~A232 & A203;
  assign \new_[57600]_  = \new_[57599]_  & \new_[57596]_ ;
  assign \new_[57601]_  = \new_[57600]_  & \new_[57593]_ ;
  assign \new_[57604]_  = ~A235 & ~A233;
  assign \new_[57607]_  = ~A268 & ~A267;
  assign \new_[57608]_  = \new_[57607]_  & \new_[57604]_ ;
  assign \new_[57611]_  = ~A298 & ~A269;
  assign \new_[57614]_  = A302 & A299;
  assign \new_[57615]_  = \new_[57614]_  & \new_[57611]_ ;
  assign \new_[57616]_  = \new_[57615]_  & \new_[57608]_ ;
  assign \new_[57620]_  = ~A168 & ~A169;
  assign \new_[57621]_  = ~A170 & \new_[57620]_ ;
  assign \new_[57624]_  = ~A200 & A199;
  assign \new_[57627]_  = ~A232 & A203;
  assign \new_[57628]_  = \new_[57627]_  & \new_[57624]_ ;
  assign \new_[57629]_  = \new_[57628]_  & \new_[57621]_ ;
  assign \new_[57632]_  = ~A235 & ~A233;
  assign \new_[57635]_  = A266 & A265;
  assign \new_[57636]_  = \new_[57635]_  & \new_[57632]_ ;
  assign \new_[57639]_  = ~A268 & ~A267;
  assign \new_[57642]_  = A300 & A299;
  assign \new_[57643]_  = \new_[57642]_  & \new_[57639]_ ;
  assign \new_[57644]_  = \new_[57643]_  & \new_[57636]_ ;
  assign \new_[57648]_  = ~A168 & ~A169;
  assign \new_[57649]_  = ~A170 & \new_[57648]_ ;
  assign \new_[57652]_  = ~A200 & A199;
  assign \new_[57655]_  = ~A232 & A203;
  assign \new_[57656]_  = \new_[57655]_  & \new_[57652]_ ;
  assign \new_[57657]_  = \new_[57656]_  & \new_[57649]_ ;
  assign \new_[57660]_  = ~A235 & ~A233;
  assign \new_[57663]_  = A266 & A265;
  assign \new_[57664]_  = \new_[57663]_  & \new_[57660]_ ;
  assign \new_[57667]_  = ~A268 & ~A267;
  assign \new_[57670]_  = A300 & A298;
  assign \new_[57671]_  = \new_[57670]_  & \new_[57667]_ ;
  assign \new_[57672]_  = \new_[57671]_  & \new_[57664]_ ;
  assign \new_[57676]_  = ~A168 & ~A169;
  assign \new_[57677]_  = ~A170 & \new_[57676]_ ;
  assign \new_[57680]_  = ~A200 & A199;
  assign \new_[57683]_  = ~A232 & A203;
  assign \new_[57684]_  = \new_[57683]_  & \new_[57680]_ ;
  assign \new_[57685]_  = \new_[57684]_  & \new_[57677]_ ;
  assign \new_[57688]_  = ~A235 & ~A233;
  assign \new_[57691]_  = ~A266 & ~A265;
  assign \new_[57692]_  = \new_[57691]_  & \new_[57688]_ ;
  assign \new_[57695]_  = A298 & ~A268;
  assign \new_[57698]_  = A302 & ~A299;
  assign \new_[57699]_  = \new_[57698]_  & \new_[57695]_ ;
  assign \new_[57700]_  = \new_[57699]_  & \new_[57692]_ ;
  assign \new_[57704]_  = ~A168 & ~A169;
  assign \new_[57705]_  = ~A170 & \new_[57704]_ ;
  assign \new_[57708]_  = ~A200 & A199;
  assign \new_[57711]_  = ~A232 & A203;
  assign \new_[57712]_  = \new_[57711]_  & \new_[57708]_ ;
  assign \new_[57713]_  = \new_[57712]_  & \new_[57705]_ ;
  assign \new_[57716]_  = ~A235 & ~A233;
  assign \new_[57719]_  = ~A266 & ~A265;
  assign \new_[57720]_  = \new_[57719]_  & \new_[57716]_ ;
  assign \new_[57723]_  = ~A298 & ~A268;
  assign \new_[57726]_  = A302 & A299;
  assign \new_[57727]_  = \new_[57726]_  & \new_[57723]_ ;
  assign \new_[57728]_  = \new_[57727]_  & \new_[57720]_ ;
  assign \new_[57731]_  = A166 & A168;
  assign \new_[57734]_  = ~A202 & ~A201;
  assign \new_[57735]_  = \new_[57734]_  & \new_[57731]_ ;
  assign \new_[57738]_  = A232 & ~A203;
  assign \new_[57741]_  = ~A234 & A233;
  assign \new_[57742]_  = \new_[57741]_  & \new_[57738]_ ;
  assign \new_[57743]_  = \new_[57742]_  & \new_[57735]_ ;
  assign \new_[57746]_  = A265 & ~A235;
  assign \new_[57749]_  = ~A267 & A266;
  assign \new_[57750]_  = \new_[57749]_  & \new_[57746]_ ;
  assign \new_[57753]_  = A298 & ~A268;
  assign \new_[57756]_  = A302 & ~A299;
  assign \new_[57757]_  = \new_[57756]_  & \new_[57753]_ ;
  assign \new_[57758]_  = \new_[57757]_  & \new_[57750]_ ;
  assign \new_[57761]_  = A166 & A168;
  assign \new_[57764]_  = ~A202 & ~A201;
  assign \new_[57765]_  = \new_[57764]_  & \new_[57761]_ ;
  assign \new_[57768]_  = A232 & ~A203;
  assign \new_[57771]_  = ~A234 & A233;
  assign \new_[57772]_  = \new_[57771]_  & \new_[57768]_ ;
  assign \new_[57773]_  = \new_[57772]_  & \new_[57765]_ ;
  assign \new_[57776]_  = A265 & ~A235;
  assign \new_[57779]_  = ~A267 & A266;
  assign \new_[57780]_  = \new_[57779]_  & \new_[57776]_ ;
  assign \new_[57783]_  = ~A298 & ~A268;
  assign \new_[57786]_  = A302 & A299;
  assign \new_[57787]_  = \new_[57786]_  & \new_[57783]_ ;
  assign \new_[57788]_  = \new_[57787]_  & \new_[57780]_ ;
  assign \new_[57791]_  = A166 & A168;
  assign \new_[57794]_  = A200 & A199;
  assign \new_[57795]_  = \new_[57794]_  & \new_[57791]_ ;
  assign \new_[57798]_  = ~A202 & ~A201;
  assign \new_[57801]_  = ~A235 & ~A234;
  assign \new_[57802]_  = \new_[57801]_  & \new_[57798]_ ;
  assign \new_[57803]_  = \new_[57802]_  & \new_[57795]_ ;
  assign \new_[57806]_  = A265 & ~A236;
  assign \new_[57809]_  = ~A267 & A266;
  assign \new_[57810]_  = \new_[57809]_  & \new_[57806]_ ;
  assign \new_[57813]_  = A298 & ~A268;
  assign \new_[57816]_  = A302 & ~A299;
  assign \new_[57817]_  = \new_[57816]_  & \new_[57813]_ ;
  assign \new_[57818]_  = \new_[57817]_  & \new_[57810]_ ;
  assign \new_[57821]_  = A166 & A168;
  assign \new_[57824]_  = A200 & A199;
  assign \new_[57825]_  = \new_[57824]_  & \new_[57821]_ ;
  assign \new_[57828]_  = ~A202 & ~A201;
  assign \new_[57831]_  = ~A235 & ~A234;
  assign \new_[57832]_  = \new_[57831]_  & \new_[57828]_ ;
  assign \new_[57833]_  = \new_[57832]_  & \new_[57825]_ ;
  assign \new_[57836]_  = A265 & ~A236;
  assign \new_[57839]_  = ~A267 & A266;
  assign \new_[57840]_  = \new_[57839]_  & \new_[57836]_ ;
  assign \new_[57843]_  = ~A298 & ~A268;
  assign \new_[57846]_  = A302 & A299;
  assign \new_[57847]_  = \new_[57846]_  & \new_[57843]_ ;
  assign \new_[57848]_  = \new_[57847]_  & \new_[57840]_ ;
  assign \new_[57851]_  = A166 & A168;
  assign \new_[57854]_  = A200 & A199;
  assign \new_[57855]_  = \new_[57854]_  & \new_[57851]_ ;
  assign \new_[57858]_  = ~A202 & ~A201;
  assign \new_[57861]_  = A233 & A232;
  assign \new_[57862]_  = \new_[57861]_  & \new_[57858]_ ;
  assign \new_[57863]_  = \new_[57862]_  & \new_[57855]_ ;
  assign \new_[57866]_  = ~A235 & ~A234;
  assign \new_[57869]_  = ~A268 & ~A267;
  assign \new_[57870]_  = \new_[57869]_  & \new_[57866]_ ;
  assign \new_[57873]_  = A298 & ~A269;
  assign \new_[57876]_  = A302 & ~A299;
  assign \new_[57877]_  = \new_[57876]_  & \new_[57873]_ ;
  assign \new_[57878]_  = \new_[57877]_  & \new_[57870]_ ;
  assign \new_[57881]_  = A166 & A168;
  assign \new_[57884]_  = A200 & A199;
  assign \new_[57885]_  = \new_[57884]_  & \new_[57881]_ ;
  assign \new_[57888]_  = ~A202 & ~A201;
  assign \new_[57891]_  = A233 & A232;
  assign \new_[57892]_  = \new_[57891]_  & \new_[57888]_ ;
  assign \new_[57893]_  = \new_[57892]_  & \new_[57885]_ ;
  assign \new_[57896]_  = ~A235 & ~A234;
  assign \new_[57899]_  = ~A268 & ~A267;
  assign \new_[57900]_  = \new_[57899]_  & \new_[57896]_ ;
  assign \new_[57903]_  = ~A298 & ~A269;
  assign \new_[57906]_  = A302 & A299;
  assign \new_[57907]_  = \new_[57906]_  & \new_[57903]_ ;
  assign \new_[57908]_  = \new_[57907]_  & \new_[57900]_ ;
  assign \new_[57911]_  = A166 & A168;
  assign \new_[57914]_  = A200 & A199;
  assign \new_[57915]_  = \new_[57914]_  & \new_[57911]_ ;
  assign \new_[57918]_  = ~A202 & ~A201;
  assign \new_[57921]_  = A233 & A232;
  assign \new_[57922]_  = \new_[57921]_  & \new_[57918]_ ;
  assign \new_[57923]_  = \new_[57922]_  & \new_[57915]_ ;
  assign \new_[57926]_  = ~A235 & ~A234;
  assign \new_[57929]_  = A266 & A265;
  assign \new_[57930]_  = \new_[57929]_  & \new_[57926]_ ;
  assign \new_[57933]_  = ~A268 & ~A267;
  assign \new_[57936]_  = A300 & A299;
  assign \new_[57937]_  = \new_[57936]_  & \new_[57933]_ ;
  assign \new_[57938]_  = \new_[57937]_  & \new_[57930]_ ;
  assign \new_[57941]_  = A166 & A168;
  assign \new_[57944]_  = A200 & A199;
  assign \new_[57945]_  = \new_[57944]_  & \new_[57941]_ ;
  assign \new_[57948]_  = ~A202 & ~A201;
  assign \new_[57951]_  = A233 & A232;
  assign \new_[57952]_  = \new_[57951]_  & \new_[57948]_ ;
  assign \new_[57953]_  = \new_[57952]_  & \new_[57945]_ ;
  assign \new_[57956]_  = ~A235 & ~A234;
  assign \new_[57959]_  = A266 & A265;
  assign \new_[57960]_  = \new_[57959]_  & \new_[57956]_ ;
  assign \new_[57963]_  = ~A268 & ~A267;
  assign \new_[57966]_  = A300 & A298;
  assign \new_[57967]_  = \new_[57966]_  & \new_[57963]_ ;
  assign \new_[57968]_  = \new_[57967]_  & \new_[57960]_ ;
  assign \new_[57971]_  = A166 & A168;
  assign \new_[57974]_  = A200 & A199;
  assign \new_[57975]_  = \new_[57974]_  & \new_[57971]_ ;
  assign \new_[57978]_  = ~A202 & ~A201;
  assign \new_[57981]_  = A233 & A232;
  assign \new_[57982]_  = \new_[57981]_  & \new_[57978]_ ;
  assign \new_[57983]_  = \new_[57982]_  & \new_[57975]_ ;
  assign \new_[57986]_  = ~A235 & ~A234;
  assign \new_[57989]_  = ~A266 & ~A265;
  assign \new_[57990]_  = \new_[57989]_  & \new_[57986]_ ;
  assign \new_[57993]_  = A298 & ~A268;
  assign \new_[57996]_  = A302 & ~A299;
  assign \new_[57997]_  = \new_[57996]_  & \new_[57993]_ ;
  assign \new_[57998]_  = \new_[57997]_  & \new_[57990]_ ;
  assign \new_[58001]_  = A166 & A168;
  assign \new_[58004]_  = A200 & A199;
  assign \new_[58005]_  = \new_[58004]_  & \new_[58001]_ ;
  assign \new_[58008]_  = ~A202 & ~A201;
  assign \new_[58011]_  = A233 & A232;
  assign \new_[58012]_  = \new_[58011]_  & \new_[58008]_ ;
  assign \new_[58013]_  = \new_[58012]_  & \new_[58005]_ ;
  assign \new_[58016]_  = ~A235 & ~A234;
  assign \new_[58019]_  = ~A266 & ~A265;
  assign \new_[58020]_  = \new_[58019]_  & \new_[58016]_ ;
  assign \new_[58023]_  = ~A298 & ~A268;
  assign \new_[58026]_  = A302 & A299;
  assign \new_[58027]_  = \new_[58026]_  & \new_[58023]_ ;
  assign \new_[58028]_  = \new_[58027]_  & \new_[58020]_ ;
  assign \new_[58031]_  = A166 & A168;
  assign \new_[58034]_  = A200 & A199;
  assign \new_[58035]_  = \new_[58034]_  & \new_[58031]_ ;
  assign \new_[58038]_  = ~A202 & ~A201;
  assign \new_[58041]_  = ~A233 & ~A232;
  assign \new_[58042]_  = \new_[58041]_  & \new_[58038]_ ;
  assign \new_[58043]_  = \new_[58042]_  & \new_[58035]_ ;
  assign \new_[58046]_  = A265 & ~A235;
  assign \new_[58049]_  = ~A267 & A266;
  assign \new_[58050]_  = \new_[58049]_  & \new_[58046]_ ;
  assign \new_[58053]_  = A298 & ~A268;
  assign \new_[58056]_  = A302 & ~A299;
  assign \new_[58057]_  = \new_[58056]_  & \new_[58053]_ ;
  assign \new_[58058]_  = \new_[58057]_  & \new_[58050]_ ;
  assign \new_[58061]_  = A166 & A168;
  assign \new_[58064]_  = A200 & A199;
  assign \new_[58065]_  = \new_[58064]_  & \new_[58061]_ ;
  assign \new_[58068]_  = ~A202 & ~A201;
  assign \new_[58071]_  = ~A233 & ~A232;
  assign \new_[58072]_  = \new_[58071]_  & \new_[58068]_ ;
  assign \new_[58073]_  = \new_[58072]_  & \new_[58065]_ ;
  assign \new_[58076]_  = A265 & ~A235;
  assign \new_[58079]_  = ~A267 & A266;
  assign \new_[58080]_  = \new_[58079]_  & \new_[58076]_ ;
  assign \new_[58083]_  = ~A298 & ~A268;
  assign \new_[58086]_  = A302 & A299;
  assign \new_[58087]_  = \new_[58086]_  & \new_[58083]_ ;
  assign \new_[58088]_  = \new_[58087]_  & \new_[58080]_ ;
  assign \new_[58091]_  = A166 & A168;
  assign \new_[58094]_  = ~A200 & ~A199;
  assign \new_[58095]_  = \new_[58094]_  & \new_[58091]_ ;
  assign \new_[58098]_  = A232 & ~A202;
  assign \new_[58101]_  = ~A234 & A233;
  assign \new_[58102]_  = \new_[58101]_  & \new_[58098]_ ;
  assign \new_[58103]_  = \new_[58102]_  & \new_[58095]_ ;
  assign \new_[58106]_  = A265 & ~A235;
  assign \new_[58109]_  = ~A267 & A266;
  assign \new_[58110]_  = \new_[58109]_  & \new_[58106]_ ;
  assign \new_[58113]_  = A298 & ~A268;
  assign \new_[58116]_  = A302 & ~A299;
  assign \new_[58117]_  = \new_[58116]_  & \new_[58113]_ ;
  assign \new_[58118]_  = \new_[58117]_  & \new_[58110]_ ;
  assign \new_[58121]_  = A166 & A168;
  assign \new_[58124]_  = ~A200 & ~A199;
  assign \new_[58125]_  = \new_[58124]_  & \new_[58121]_ ;
  assign \new_[58128]_  = A232 & ~A202;
  assign \new_[58131]_  = ~A234 & A233;
  assign \new_[58132]_  = \new_[58131]_  & \new_[58128]_ ;
  assign \new_[58133]_  = \new_[58132]_  & \new_[58125]_ ;
  assign \new_[58136]_  = A265 & ~A235;
  assign \new_[58139]_  = ~A267 & A266;
  assign \new_[58140]_  = \new_[58139]_  & \new_[58136]_ ;
  assign \new_[58143]_  = ~A298 & ~A268;
  assign \new_[58146]_  = A302 & A299;
  assign \new_[58147]_  = \new_[58146]_  & \new_[58143]_ ;
  assign \new_[58148]_  = \new_[58147]_  & \new_[58140]_ ;
  assign \new_[58151]_  = A167 & A168;
  assign \new_[58154]_  = ~A202 & ~A201;
  assign \new_[58155]_  = \new_[58154]_  & \new_[58151]_ ;
  assign \new_[58158]_  = A232 & ~A203;
  assign \new_[58161]_  = ~A234 & A233;
  assign \new_[58162]_  = \new_[58161]_  & \new_[58158]_ ;
  assign \new_[58163]_  = \new_[58162]_  & \new_[58155]_ ;
  assign \new_[58166]_  = A265 & ~A235;
  assign \new_[58169]_  = ~A267 & A266;
  assign \new_[58170]_  = \new_[58169]_  & \new_[58166]_ ;
  assign \new_[58173]_  = A298 & ~A268;
  assign \new_[58176]_  = A302 & ~A299;
  assign \new_[58177]_  = \new_[58176]_  & \new_[58173]_ ;
  assign \new_[58178]_  = \new_[58177]_  & \new_[58170]_ ;
  assign \new_[58181]_  = A167 & A168;
  assign \new_[58184]_  = ~A202 & ~A201;
  assign \new_[58185]_  = \new_[58184]_  & \new_[58181]_ ;
  assign \new_[58188]_  = A232 & ~A203;
  assign \new_[58191]_  = ~A234 & A233;
  assign \new_[58192]_  = \new_[58191]_  & \new_[58188]_ ;
  assign \new_[58193]_  = \new_[58192]_  & \new_[58185]_ ;
  assign \new_[58196]_  = A265 & ~A235;
  assign \new_[58199]_  = ~A267 & A266;
  assign \new_[58200]_  = \new_[58199]_  & \new_[58196]_ ;
  assign \new_[58203]_  = ~A298 & ~A268;
  assign \new_[58206]_  = A302 & A299;
  assign \new_[58207]_  = \new_[58206]_  & \new_[58203]_ ;
  assign \new_[58208]_  = \new_[58207]_  & \new_[58200]_ ;
  assign \new_[58211]_  = A167 & A168;
  assign \new_[58214]_  = A200 & A199;
  assign \new_[58215]_  = \new_[58214]_  & \new_[58211]_ ;
  assign \new_[58218]_  = ~A202 & ~A201;
  assign \new_[58221]_  = ~A235 & ~A234;
  assign \new_[58222]_  = \new_[58221]_  & \new_[58218]_ ;
  assign \new_[58223]_  = \new_[58222]_  & \new_[58215]_ ;
  assign \new_[58226]_  = A265 & ~A236;
  assign \new_[58229]_  = ~A267 & A266;
  assign \new_[58230]_  = \new_[58229]_  & \new_[58226]_ ;
  assign \new_[58233]_  = A298 & ~A268;
  assign \new_[58236]_  = A302 & ~A299;
  assign \new_[58237]_  = \new_[58236]_  & \new_[58233]_ ;
  assign \new_[58238]_  = \new_[58237]_  & \new_[58230]_ ;
  assign \new_[58241]_  = A167 & A168;
  assign \new_[58244]_  = A200 & A199;
  assign \new_[58245]_  = \new_[58244]_  & \new_[58241]_ ;
  assign \new_[58248]_  = ~A202 & ~A201;
  assign \new_[58251]_  = ~A235 & ~A234;
  assign \new_[58252]_  = \new_[58251]_  & \new_[58248]_ ;
  assign \new_[58253]_  = \new_[58252]_  & \new_[58245]_ ;
  assign \new_[58256]_  = A265 & ~A236;
  assign \new_[58259]_  = ~A267 & A266;
  assign \new_[58260]_  = \new_[58259]_  & \new_[58256]_ ;
  assign \new_[58263]_  = ~A298 & ~A268;
  assign \new_[58266]_  = A302 & A299;
  assign \new_[58267]_  = \new_[58266]_  & \new_[58263]_ ;
  assign \new_[58268]_  = \new_[58267]_  & \new_[58260]_ ;
  assign \new_[58271]_  = A167 & A168;
  assign \new_[58274]_  = A200 & A199;
  assign \new_[58275]_  = \new_[58274]_  & \new_[58271]_ ;
  assign \new_[58278]_  = ~A202 & ~A201;
  assign \new_[58281]_  = A233 & A232;
  assign \new_[58282]_  = \new_[58281]_  & \new_[58278]_ ;
  assign \new_[58283]_  = \new_[58282]_  & \new_[58275]_ ;
  assign \new_[58286]_  = ~A235 & ~A234;
  assign \new_[58289]_  = ~A268 & ~A267;
  assign \new_[58290]_  = \new_[58289]_  & \new_[58286]_ ;
  assign \new_[58293]_  = A298 & ~A269;
  assign \new_[58296]_  = A302 & ~A299;
  assign \new_[58297]_  = \new_[58296]_  & \new_[58293]_ ;
  assign \new_[58298]_  = \new_[58297]_  & \new_[58290]_ ;
  assign \new_[58301]_  = A167 & A168;
  assign \new_[58304]_  = A200 & A199;
  assign \new_[58305]_  = \new_[58304]_  & \new_[58301]_ ;
  assign \new_[58308]_  = ~A202 & ~A201;
  assign \new_[58311]_  = A233 & A232;
  assign \new_[58312]_  = \new_[58311]_  & \new_[58308]_ ;
  assign \new_[58313]_  = \new_[58312]_  & \new_[58305]_ ;
  assign \new_[58316]_  = ~A235 & ~A234;
  assign \new_[58319]_  = ~A268 & ~A267;
  assign \new_[58320]_  = \new_[58319]_  & \new_[58316]_ ;
  assign \new_[58323]_  = ~A298 & ~A269;
  assign \new_[58326]_  = A302 & A299;
  assign \new_[58327]_  = \new_[58326]_  & \new_[58323]_ ;
  assign \new_[58328]_  = \new_[58327]_  & \new_[58320]_ ;
  assign \new_[58331]_  = A167 & A168;
  assign \new_[58334]_  = A200 & A199;
  assign \new_[58335]_  = \new_[58334]_  & \new_[58331]_ ;
  assign \new_[58338]_  = ~A202 & ~A201;
  assign \new_[58341]_  = A233 & A232;
  assign \new_[58342]_  = \new_[58341]_  & \new_[58338]_ ;
  assign \new_[58343]_  = \new_[58342]_  & \new_[58335]_ ;
  assign \new_[58346]_  = ~A235 & ~A234;
  assign \new_[58349]_  = A266 & A265;
  assign \new_[58350]_  = \new_[58349]_  & \new_[58346]_ ;
  assign \new_[58353]_  = ~A268 & ~A267;
  assign \new_[58356]_  = A300 & A299;
  assign \new_[58357]_  = \new_[58356]_  & \new_[58353]_ ;
  assign \new_[58358]_  = \new_[58357]_  & \new_[58350]_ ;
  assign \new_[58361]_  = A167 & A168;
  assign \new_[58364]_  = A200 & A199;
  assign \new_[58365]_  = \new_[58364]_  & \new_[58361]_ ;
  assign \new_[58368]_  = ~A202 & ~A201;
  assign \new_[58371]_  = A233 & A232;
  assign \new_[58372]_  = \new_[58371]_  & \new_[58368]_ ;
  assign \new_[58373]_  = \new_[58372]_  & \new_[58365]_ ;
  assign \new_[58376]_  = ~A235 & ~A234;
  assign \new_[58379]_  = A266 & A265;
  assign \new_[58380]_  = \new_[58379]_  & \new_[58376]_ ;
  assign \new_[58383]_  = ~A268 & ~A267;
  assign \new_[58386]_  = A300 & A298;
  assign \new_[58387]_  = \new_[58386]_  & \new_[58383]_ ;
  assign \new_[58388]_  = \new_[58387]_  & \new_[58380]_ ;
  assign \new_[58391]_  = A167 & A168;
  assign \new_[58394]_  = A200 & A199;
  assign \new_[58395]_  = \new_[58394]_  & \new_[58391]_ ;
  assign \new_[58398]_  = ~A202 & ~A201;
  assign \new_[58401]_  = A233 & A232;
  assign \new_[58402]_  = \new_[58401]_  & \new_[58398]_ ;
  assign \new_[58403]_  = \new_[58402]_  & \new_[58395]_ ;
  assign \new_[58406]_  = ~A235 & ~A234;
  assign \new_[58409]_  = ~A266 & ~A265;
  assign \new_[58410]_  = \new_[58409]_  & \new_[58406]_ ;
  assign \new_[58413]_  = A298 & ~A268;
  assign \new_[58416]_  = A302 & ~A299;
  assign \new_[58417]_  = \new_[58416]_  & \new_[58413]_ ;
  assign \new_[58418]_  = \new_[58417]_  & \new_[58410]_ ;
  assign \new_[58421]_  = A167 & A168;
  assign \new_[58424]_  = A200 & A199;
  assign \new_[58425]_  = \new_[58424]_  & \new_[58421]_ ;
  assign \new_[58428]_  = ~A202 & ~A201;
  assign \new_[58431]_  = A233 & A232;
  assign \new_[58432]_  = \new_[58431]_  & \new_[58428]_ ;
  assign \new_[58433]_  = \new_[58432]_  & \new_[58425]_ ;
  assign \new_[58436]_  = ~A235 & ~A234;
  assign \new_[58439]_  = ~A266 & ~A265;
  assign \new_[58440]_  = \new_[58439]_  & \new_[58436]_ ;
  assign \new_[58443]_  = ~A298 & ~A268;
  assign \new_[58446]_  = A302 & A299;
  assign \new_[58447]_  = \new_[58446]_  & \new_[58443]_ ;
  assign \new_[58448]_  = \new_[58447]_  & \new_[58440]_ ;
  assign \new_[58451]_  = A167 & A168;
  assign \new_[58454]_  = A200 & A199;
  assign \new_[58455]_  = \new_[58454]_  & \new_[58451]_ ;
  assign \new_[58458]_  = ~A202 & ~A201;
  assign \new_[58461]_  = ~A233 & ~A232;
  assign \new_[58462]_  = \new_[58461]_  & \new_[58458]_ ;
  assign \new_[58463]_  = \new_[58462]_  & \new_[58455]_ ;
  assign \new_[58466]_  = A265 & ~A235;
  assign \new_[58469]_  = ~A267 & A266;
  assign \new_[58470]_  = \new_[58469]_  & \new_[58466]_ ;
  assign \new_[58473]_  = A298 & ~A268;
  assign \new_[58476]_  = A302 & ~A299;
  assign \new_[58477]_  = \new_[58476]_  & \new_[58473]_ ;
  assign \new_[58478]_  = \new_[58477]_  & \new_[58470]_ ;
  assign \new_[58481]_  = A167 & A168;
  assign \new_[58484]_  = A200 & A199;
  assign \new_[58485]_  = \new_[58484]_  & \new_[58481]_ ;
  assign \new_[58488]_  = ~A202 & ~A201;
  assign \new_[58491]_  = ~A233 & ~A232;
  assign \new_[58492]_  = \new_[58491]_  & \new_[58488]_ ;
  assign \new_[58493]_  = \new_[58492]_  & \new_[58485]_ ;
  assign \new_[58496]_  = A265 & ~A235;
  assign \new_[58499]_  = ~A267 & A266;
  assign \new_[58500]_  = \new_[58499]_  & \new_[58496]_ ;
  assign \new_[58503]_  = ~A298 & ~A268;
  assign \new_[58506]_  = A302 & A299;
  assign \new_[58507]_  = \new_[58506]_  & \new_[58503]_ ;
  assign \new_[58508]_  = \new_[58507]_  & \new_[58500]_ ;
  assign \new_[58511]_  = A167 & A168;
  assign \new_[58514]_  = ~A200 & ~A199;
  assign \new_[58515]_  = \new_[58514]_  & \new_[58511]_ ;
  assign \new_[58518]_  = A232 & ~A202;
  assign \new_[58521]_  = ~A234 & A233;
  assign \new_[58522]_  = \new_[58521]_  & \new_[58518]_ ;
  assign \new_[58523]_  = \new_[58522]_  & \new_[58515]_ ;
  assign \new_[58526]_  = A265 & ~A235;
  assign \new_[58529]_  = ~A267 & A266;
  assign \new_[58530]_  = \new_[58529]_  & \new_[58526]_ ;
  assign \new_[58533]_  = A298 & ~A268;
  assign \new_[58536]_  = A302 & ~A299;
  assign \new_[58537]_  = \new_[58536]_  & \new_[58533]_ ;
  assign \new_[58538]_  = \new_[58537]_  & \new_[58530]_ ;
  assign \new_[58541]_  = A167 & A168;
  assign \new_[58544]_  = ~A200 & ~A199;
  assign \new_[58545]_  = \new_[58544]_  & \new_[58541]_ ;
  assign \new_[58548]_  = A232 & ~A202;
  assign \new_[58551]_  = ~A234 & A233;
  assign \new_[58552]_  = \new_[58551]_  & \new_[58548]_ ;
  assign \new_[58553]_  = \new_[58552]_  & \new_[58545]_ ;
  assign \new_[58556]_  = A265 & ~A235;
  assign \new_[58559]_  = ~A267 & A266;
  assign \new_[58560]_  = \new_[58559]_  & \new_[58556]_ ;
  assign \new_[58563]_  = ~A298 & ~A268;
  assign \new_[58566]_  = A302 & A299;
  assign \new_[58567]_  = \new_[58566]_  & \new_[58563]_ ;
  assign \new_[58568]_  = \new_[58567]_  & \new_[58560]_ ;
  assign \new_[58571]_  = A167 & A170;
  assign \new_[58574]_  = ~A201 & ~A166;
  assign \new_[58575]_  = \new_[58574]_  & \new_[58571]_ ;
  assign \new_[58578]_  = ~A203 & ~A202;
  assign \new_[58581]_  = ~A235 & ~A234;
  assign \new_[58582]_  = \new_[58581]_  & \new_[58578]_ ;
  assign \new_[58583]_  = \new_[58582]_  & \new_[58575]_ ;
  assign \new_[58586]_  = A265 & ~A236;
  assign \new_[58589]_  = ~A267 & A266;
  assign \new_[58590]_  = \new_[58589]_  & \new_[58586]_ ;
  assign \new_[58593]_  = A298 & ~A268;
  assign \new_[58596]_  = A302 & ~A299;
  assign \new_[58597]_  = \new_[58596]_  & \new_[58593]_ ;
  assign \new_[58598]_  = \new_[58597]_  & \new_[58590]_ ;
  assign \new_[58601]_  = A167 & A170;
  assign \new_[58604]_  = ~A201 & ~A166;
  assign \new_[58605]_  = \new_[58604]_  & \new_[58601]_ ;
  assign \new_[58608]_  = ~A203 & ~A202;
  assign \new_[58611]_  = ~A235 & ~A234;
  assign \new_[58612]_  = \new_[58611]_  & \new_[58608]_ ;
  assign \new_[58613]_  = \new_[58612]_  & \new_[58605]_ ;
  assign \new_[58616]_  = A265 & ~A236;
  assign \new_[58619]_  = ~A267 & A266;
  assign \new_[58620]_  = \new_[58619]_  & \new_[58616]_ ;
  assign \new_[58623]_  = ~A298 & ~A268;
  assign \new_[58626]_  = A302 & A299;
  assign \new_[58627]_  = \new_[58626]_  & \new_[58623]_ ;
  assign \new_[58628]_  = \new_[58627]_  & \new_[58620]_ ;
  assign \new_[58631]_  = A167 & A170;
  assign \new_[58634]_  = ~A201 & ~A166;
  assign \new_[58635]_  = \new_[58634]_  & \new_[58631]_ ;
  assign \new_[58638]_  = ~A203 & ~A202;
  assign \new_[58641]_  = A233 & A232;
  assign \new_[58642]_  = \new_[58641]_  & \new_[58638]_ ;
  assign \new_[58643]_  = \new_[58642]_  & \new_[58635]_ ;
  assign \new_[58646]_  = ~A235 & ~A234;
  assign \new_[58649]_  = ~A268 & ~A267;
  assign \new_[58650]_  = \new_[58649]_  & \new_[58646]_ ;
  assign \new_[58653]_  = A298 & ~A269;
  assign \new_[58656]_  = A302 & ~A299;
  assign \new_[58657]_  = \new_[58656]_  & \new_[58653]_ ;
  assign \new_[58658]_  = \new_[58657]_  & \new_[58650]_ ;
  assign \new_[58661]_  = A167 & A170;
  assign \new_[58664]_  = ~A201 & ~A166;
  assign \new_[58665]_  = \new_[58664]_  & \new_[58661]_ ;
  assign \new_[58668]_  = ~A203 & ~A202;
  assign \new_[58671]_  = A233 & A232;
  assign \new_[58672]_  = \new_[58671]_  & \new_[58668]_ ;
  assign \new_[58673]_  = \new_[58672]_  & \new_[58665]_ ;
  assign \new_[58676]_  = ~A235 & ~A234;
  assign \new_[58679]_  = ~A268 & ~A267;
  assign \new_[58680]_  = \new_[58679]_  & \new_[58676]_ ;
  assign \new_[58683]_  = ~A298 & ~A269;
  assign \new_[58686]_  = A302 & A299;
  assign \new_[58687]_  = \new_[58686]_  & \new_[58683]_ ;
  assign \new_[58688]_  = \new_[58687]_  & \new_[58680]_ ;
  assign \new_[58691]_  = A167 & A170;
  assign \new_[58694]_  = ~A201 & ~A166;
  assign \new_[58695]_  = \new_[58694]_  & \new_[58691]_ ;
  assign \new_[58698]_  = ~A203 & ~A202;
  assign \new_[58701]_  = A233 & A232;
  assign \new_[58702]_  = \new_[58701]_  & \new_[58698]_ ;
  assign \new_[58703]_  = \new_[58702]_  & \new_[58695]_ ;
  assign \new_[58706]_  = ~A235 & ~A234;
  assign \new_[58709]_  = A266 & A265;
  assign \new_[58710]_  = \new_[58709]_  & \new_[58706]_ ;
  assign \new_[58713]_  = ~A268 & ~A267;
  assign \new_[58716]_  = A300 & A299;
  assign \new_[58717]_  = \new_[58716]_  & \new_[58713]_ ;
  assign \new_[58718]_  = \new_[58717]_  & \new_[58710]_ ;
  assign \new_[58721]_  = A167 & A170;
  assign \new_[58724]_  = ~A201 & ~A166;
  assign \new_[58725]_  = \new_[58724]_  & \new_[58721]_ ;
  assign \new_[58728]_  = ~A203 & ~A202;
  assign \new_[58731]_  = A233 & A232;
  assign \new_[58732]_  = \new_[58731]_  & \new_[58728]_ ;
  assign \new_[58733]_  = \new_[58732]_  & \new_[58725]_ ;
  assign \new_[58736]_  = ~A235 & ~A234;
  assign \new_[58739]_  = A266 & A265;
  assign \new_[58740]_  = \new_[58739]_  & \new_[58736]_ ;
  assign \new_[58743]_  = ~A268 & ~A267;
  assign \new_[58746]_  = A300 & A298;
  assign \new_[58747]_  = \new_[58746]_  & \new_[58743]_ ;
  assign \new_[58748]_  = \new_[58747]_  & \new_[58740]_ ;
  assign \new_[58751]_  = A167 & A170;
  assign \new_[58754]_  = ~A201 & ~A166;
  assign \new_[58755]_  = \new_[58754]_  & \new_[58751]_ ;
  assign \new_[58758]_  = ~A203 & ~A202;
  assign \new_[58761]_  = A233 & A232;
  assign \new_[58762]_  = \new_[58761]_  & \new_[58758]_ ;
  assign \new_[58763]_  = \new_[58762]_  & \new_[58755]_ ;
  assign \new_[58766]_  = ~A235 & ~A234;
  assign \new_[58769]_  = ~A266 & ~A265;
  assign \new_[58770]_  = \new_[58769]_  & \new_[58766]_ ;
  assign \new_[58773]_  = A298 & ~A268;
  assign \new_[58776]_  = A302 & ~A299;
  assign \new_[58777]_  = \new_[58776]_  & \new_[58773]_ ;
  assign \new_[58778]_  = \new_[58777]_  & \new_[58770]_ ;
  assign \new_[58781]_  = A167 & A170;
  assign \new_[58784]_  = ~A201 & ~A166;
  assign \new_[58785]_  = \new_[58784]_  & \new_[58781]_ ;
  assign \new_[58788]_  = ~A203 & ~A202;
  assign \new_[58791]_  = A233 & A232;
  assign \new_[58792]_  = \new_[58791]_  & \new_[58788]_ ;
  assign \new_[58793]_  = \new_[58792]_  & \new_[58785]_ ;
  assign \new_[58796]_  = ~A235 & ~A234;
  assign \new_[58799]_  = ~A266 & ~A265;
  assign \new_[58800]_  = \new_[58799]_  & \new_[58796]_ ;
  assign \new_[58803]_  = ~A298 & ~A268;
  assign \new_[58806]_  = A302 & A299;
  assign \new_[58807]_  = \new_[58806]_  & \new_[58803]_ ;
  assign \new_[58808]_  = \new_[58807]_  & \new_[58800]_ ;
  assign \new_[58811]_  = A167 & A170;
  assign \new_[58814]_  = ~A201 & ~A166;
  assign \new_[58815]_  = \new_[58814]_  & \new_[58811]_ ;
  assign \new_[58818]_  = ~A203 & ~A202;
  assign \new_[58821]_  = ~A233 & ~A232;
  assign \new_[58822]_  = \new_[58821]_  & \new_[58818]_ ;
  assign \new_[58823]_  = \new_[58822]_  & \new_[58815]_ ;
  assign \new_[58826]_  = A265 & ~A235;
  assign \new_[58829]_  = ~A267 & A266;
  assign \new_[58830]_  = \new_[58829]_  & \new_[58826]_ ;
  assign \new_[58833]_  = A298 & ~A268;
  assign \new_[58836]_  = A302 & ~A299;
  assign \new_[58837]_  = \new_[58836]_  & \new_[58833]_ ;
  assign \new_[58838]_  = \new_[58837]_  & \new_[58830]_ ;
  assign \new_[58841]_  = A167 & A170;
  assign \new_[58844]_  = ~A201 & ~A166;
  assign \new_[58845]_  = \new_[58844]_  & \new_[58841]_ ;
  assign \new_[58848]_  = ~A203 & ~A202;
  assign \new_[58851]_  = ~A233 & ~A232;
  assign \new_[58852]_  = \new_[58851]_  & \new_[58848]_ ;
  assign \new_[58853]_  = \new_[58852]_  & \new_[58845]_ ;
  assign \new_[58856]_  = A265 & ~A235;
  assign \new_[58859]_  = ~A267 & A266;
  assign \new_[58860]_  = \new_[58859]_  & \new_[58856]_ ;
  assign \new_[58863]_  = ~A298 & ~A268;
  assign \new_[58866]_  = A302 & A299;
  assign \new_[58867]_  = \new_[58866]_  & \new_[58863]_ ;
  assign \new_[58868]_  = \new_[58867]_  & \new_[58860]_ ;
  assign \new_[58871]_  = A167 & A170;
  assign \new_[58874]_  = A199 & ~A166;
  assign \new_[58875]_  = \new_[58874]_  & \new_[58871]_ ;
  assign \new_[58878]_  = ~A201 & A200;
  assign \new_[58881]_  = ~A234 & ~A202;
  assign \new_[58882]_  = \new_[58881]_  & \new_[58878]_ ;
  assign \new_[58883]_  = \new_[58882]_  & \new_[58875]_ ;
  assign \new_[58886]_  = ~A236 & ~A235;
  assign \new_[58889]_  = ~A268 & ~A267;
  assign \new_[58890]_  = \new_[58889]_  & \new_[58886]_ ;
  assign \new_[58893]_  = A298 & ~A269;
  assign \new_[58896]_  = A302 & ~A299;
  assign \new_[58897]_  = \new_[58896]_  & \new_[58893]_ ;
  assign \new_[58898]_  = \new_[58897]_  & \new_[58890]_ ;
  assign \new_[58901]_  = A167 & A170;
  assign \new_[58904]_  = A199 & ~A166;
  assign \new_[58905]_  = \new_[58904]_  & \new_[58901]_ ;
  assign \new_[58908]_  = ~A201 & A200;
  assign \new_[58911]_  = ~A234 & ~A202;
  assign \new_[58912]_  = \new_[58911]_  & \new_[58908]_ ;
  assign \new_[58913]_  = \new_[58912]_  & \new_[58905]_ ;
  assign \new_[58916]_  = ~A236 & ~A235;
  assign \new_[58919]_  = ~A268 & ~A267;
  assign \new_[58920]_  = \new_[58919]_  & \new_[58916]_ ;
  assign \new_[58923]_  = ~A298 & ~A269;
  assign \new_[58926]_  = A302 & A299;
  assign \new_[58927]_  = \new_[58926]_  & \new_[58923]_ ;
  assign \new_[58928]_  = \new_[58927]_  & \new_[58920]_ ;
  assign \new_[58931]_  = A167 & A170;
  assign \new_[58934]_  = A199 & ~A166;
  assign \new_[58935]_  = \new_[58934]_  & \new_[58931]_ ;
  assign \new_[58938]_  = ~A201 & A200;
  assign \new_[58941]_  = ~A234 & ~A202;
  assign \new_[58942]_  = \new_[58941]_  & \new_[58938]_ ;
  assign \new_[58943]_  = \new_[58942]_  & \new_[58935]_ ;
  assign \new_[58946]_  = ~A236 & ~A235;
  assign \new_[58949]_  = A266 & A265;
  assign \new_[58950]_  = \new_[58949]_  & \new_[58946]_ ;
  assign \new_[58953]_  = ~A268 & ~A267;
  assign \new_[58956]_  = A300 & A299;
  assign \new_[58957]_  = \new_[58956]_  & \new_[58953]_ ;
  assign \new_[58958]_  = \new_[58957]_  & \new_[58950]_ ;
  assign \new_[58961]_  = A167 & A170;
  assign \new_[58964]_  = A199 & ~A166;
  assign \new_[58965]_  = \new_[58964]_  & \new_[58961]_ ;
  assign \new_[58968]_  = ~A201 & A200;
  assign \new_[58971]_  = ~A234 & ~A202;
  assign \new_[58972]_  = \new_[58971]_  & \new_[58968]_ ;
  assign \new_[58973]_  = \new_[58972]_  & \new_[58965]_ ;
  assign \new_[58976]_  = ~A236 & ~A235;
  assign \new_[58979]_  = A266 & A265;
  assign \new_[58980]_  = \new_[58979]_  & \new_[58976]_ ;
  assign \new_[58983]_  = ~A268 & ~A267;
  assign \new_[58986]_  = A300 & A298;
  assign \new_[58987]_  = \new_[58986]_  & \new_[58983]_ ;
  assign \new_[58988]_  = \new_[58987]_  & \new_[58980]_ ;
  assign \new_[58991]_  = A167 & A170;
  assign \new_[58994]_  = A199 & ~A166;
  assign \new_[58995]_  = \new_[58994]_  & \new_[58991]_ ;
  assign \new_[58998]_  = ~A201 & A200;
  assign \new_[59001]_  = ~A234 & ~A202;
  assign \new_[59002]_  = \new_[59001]_  & \new_[58998]_ ;
  assign \new_[59003]_  = \new_[59002]_  & \new_[58995]_ ;
  assign \new_[59006]_  = ~A236 & ~A235;
  assign \new_[59009]_  = ~A266 & ~A265;
  assign \new_[59010]_  = \new_[59009]_  & \new_[59006]_ ;
  assign \new_[59013]_  = A298 & ~A268;
  assign \new_[59016]_  = A302 & ~A299;
  assign \new_[59017]_  = \new_[59016]_  & \new_[59013]_ ;
  assign \new_[59018]_  = \new_[59017]_  & \new_[59010]_ ;
  assign \new_[59021]_  = A167 & A170;
  assign \new_[59024]_  = A199 & ~A166;
  assign \new_[59025]_  = \new_[59024]_  & \new_[59021]_ ;
  assign \new_[59028]_  = ~A201 & A200;
  assign \new_[59031]_  = ~A234 & ~A202;
  assign \new_[59032]_  = \new_[59031]_  & \new_[59028]_ ;
  assign \new_[59033]_  = \new_[59032]_  & \new_[59025]_ ;
  assign \new_[59036]_  = ~A236 & ~A235;
  assign \new_[59039]_  = ~A266 & ~A265;
  assign \new_[59040]_  = \new_[59039]_  & \new_[59036]_ ;
  assign \new_[59043]_  = ~A298 & ~A268;
  assign \new_[59046]_  = A302 & A299;
  assign \new_[59047]_  = \new_[59046]_  & \new_[59043]_ ;
  assign \new_[59048]_  = \new_[59047]_  & \new_[59040]_ ;
  assign \new_[59051]_  = A167 & A170;
  assign \new_[59054]_  = A199 & ~A166;
  assign \new_[59055]_  = \new_[59054]_  & \new_[59051]_ ;
  assign \new_[59058]_  = ~A201 & A200;
  assign \new_[59061]_  = A232 & ~A202;
  assign \new_[59062]_  = \new_[59061]_  & \new_[59058]_ ;
  assign \new_[59063]_  = \new_[59062]_  & \new_[59055]_ ;
  assign \new_[59066]_  = ~A234 & A233;
  assign \new_[59069]_  = ~A267 & ~A235;
  assign \new_[59070]_  = \new_[59069]_  & \new_[59066]_ ;
  assign \new_[59073]_  = ~A269 & ~A268;
  assign \new_[59076]_  = A300 & A299;
  assign \new_[59077]_  = \new_[59076]_  & \new_[59073]_ ;
  assign \new_[59078]_  = \new_[59077]_  & \new_[59070]_ ;
  assign \new_[59081]_  = A167 & A170;
  assign \new_[59084]_  = A199 & ~A166;
  assign \new_[59085]_  = \new_[59084]_  & \new_[59081]_ ;
  assign \new_[59088]_  = ~A201 & A200;
  assign \new_[59091]_  = A232 & ~A202;
  assign \new_[59092]_  = \new_[59091]_  & \new_[59088]_ ;
  assign \new_[59093]_  = \new_[59092]_  & \new_[59085]_ ;
  assign \new_[59096]_  = ~A234 & A233;
  assign \new_[59099]_  = ~A267 & ~A235;
  assign \new_[59100]_  = \new_[59099]_  & \new_[59096]_ ;
  assign \new_[59103]_  = ~A269 & ~A268;
  assign \new_[59106]_  = A300 & A298;
  assign \new_[59107]_  = \new_[59106]_  & \new_[59103]_ ;
  assign \new_[59108]_  = \new_[59107]_  & \new_[59100]_ ;
  assign \new_[59111]_  = A167 & A170;
  assign \new_[59114]_  = A199 & ~A166;
  assign \new_[59115]_  = \new_[59114]_  & \new_[59111]_ ;
  assign \new_[59118]_  = ~A201 & A200;
  assign \new_[59121]_  = A232 & ~A202;
  assign \new_[59122]_  = \new_[59121]_  & \new_[59118]_ ;
  assign \new_[59123]_  = \new_[59122]_  & \new_[59115]_ ;
  assign \new_[59126]_  = ~A234 & A233;
  assign \new_[59129]_  = A265 & ~A235;
  assign \new_[59130]_  = \new_[59129]_  & \new_[59126]_ ;
  assign \new_[59133]_  = ~A267 & A266;
  assign \new_[59136]_  = A301 & ~A268;
  assign \new_[59137]_  = \new_[59136]_  & \new_[59133]_ ;
  assign \new_[59138]_  = \new_[59137]_  & \new_[59130]_ ;
  assign \new_[59141]_  = A167 & A170;
  assign \new_[59144]_  = A199 & ~A166;
  assign \new_[59145]_  = \new_[59144]_  & \new_[59141]_ ;
  assign \new_[59148]_  = ~A201 & A200;
  assign \new_[59151]_  = A232 & ~A202;
  assign \new_[59152]_  = \new_[59151]_  & \new_[59148]_ ;
  assign \new_[59153]_  = \new_[59152]_  & \new_[59145]_ ;
  assign \new_[59156]_  = ~A234 & A233;
  assign \new_[59159]_  = ~A265 & ~A235;
  assign \new_[59160]_  = \new_[59159]_  & \new_[59156]_ ;
  assign \new_[59163]_  = ~A268 & ~A266;
  assign \new_[59166]_  = A300 & A299;
  assign \new_[59167]_  = \new_[59166]_  & \new_[59163]_ ;
  assign \new_[59168]_  = \new_[59167]_  & \new_[59160]_ ;
  assign \new_[59171]_  = A167 & A170;
  assign \new_[59174]_  = A199 & ~A166;
  assign \new_[59175]_  = \new_[59174]_  & \new_[59171]_ ;
  assign \new_[59178]_  = ~A201 & A200;
  assign \new_[59181]_  = A232 & ~A202;
  assign \new_[59182]_  = \new_[59181]_  & \new_[59178]_ ;
  assign \new_[59183]_  = \new_[59182]_  & \new_[59175]_ ;
  assign \new_[59186]_  = ~A234 & A233;
  assign \new_[59189]_  = ~A265 & ~A235;
  assign \new_[59190]_  = \new_[59189]_  & \new_[59186]_ ;
  assign \new_[59193]_  = ~A268 & ~A266;
  assign \new_[59196]_  = A300 & A298;
  assign \new_[59197]_  = \new_[59196]_  & \new_[59193]_ ;
  assign \new_[59198]_  = \new_[59197]_  & \new_[59190]_ ;
  assign \new_[59201]_  = A167 & A170;
  assign \new_[59204]_  = A199 & ~A166;
  assign \new_[59205]_  = \new_[59204]_  & \new_[59201]_ ;
  assign \new_[59208]_  = ~A201 & A200;
  assign \new_[59211]_  = ~A232 & ~A202;
  assign \new_[59212]_  = \new_[59211]_  & \new_[59208]_ ;
  assign \new_[59213]_  = \new_[59212]_  & \new_[59205]_ ;
  assign \new_[59216]_  = ~A235 & ~A233;
  assign \new_[59219]_  = ~A268 & ~A267;
  assign \new_[59220]_  = \new_[59219]_  & \new_[59216]_ ;
  assign \new_[59223]_  = A298 & ~A269;
  assign \new_[59226]_  = A302 & ~A299;
  assign \new_[59227]_  = \new_[59226]_  & \new_[59223]_ ;
  assign \new_[59228]_  = \new_[59227]_  & \new_[59220]_ ;
  assign \new_[59231]_  = A167 & A170;
  assign \new_[59234]_  = A199 & ~A166;
  assign \new_[59235]_  = \new_[59234]_  & \new_[59231]_ ;
  assign \new_[59238]_  = ~A201 & A200;
  assign \new_[59241]_  = ~A232 & ~A202;
  assign \new_[59242]_  = \new_[59241]_  & \new_[59238]_ ;
  assign \new_[59243]_  = \new_[59242]_  & \new_[59235]_ ;
  assign \new_[59246]_  = ~A235 & ~A233;
  assign \new_[59249]_  = ~A268 & ~A267;
  assign \new_[59250]_  = \new_[59249]_  & \new_[59246]_ ;
  assign \new_[59253]_  = ~A298 & ~A269;
  assign \new_[59256]_  = A302 & A299;
  assign \new_[59257]_  = \new_[59256]_  & \new_[59253]_ ;
  assign \new_[59258]_  = \new_[59257]_  & \new_[59250]_ ;
  assign \new_[59261]_  = A167 & A170;
  assign \new_[59264]_  = A199 & ~A166;
  assign \new_[59265]_  = \new_[59264]_  & \new_[59261]_ ;
  assign \new_[59268]_  = ~A201 & A200;
  assign \new_[59271]_  = ~A232 & ~A202;
  assign \new_[59272]_  = \new_[59271]_  & \new_[59268]_ ;
  assign \new_[59273]_  = \new_[59272]_  & \new_[59265]_ ;
  assign \new_[59276]_  = ~A235 & ~A233;
  assign \new_[59279]_  = A266 & A265;
  assign \new_[59280]_  = \new_[59279]_  & \new_[59276]_ ;
  assign \new_[59283]_  = ~A268 & ~A267;
  assign \new_[59286]_  = A300 & A299;
  assign \new_[59287]_  = \new_[59286]_  & \new_[59283]_ ;
  assign \new_[59288]_  = \new_[59287]_  & \new_[59280]_ ;
  assign \new_[59291]_  = A167 & A170;
  assign \new_[59294]_  = A199 & ~A166;
  assign \new_[59295]_  = \new_[59294]_  & \new_[59291]_ ;
  assign \new_[59298]_  = ~A201 & A200;
  assign \new_[59301]_  = ~A232 & ~A202;
  assign \new_[59302]_  = \new_[59301]_  & \new_[59298]_ ;
  assign \new_[59303]_  = \new_[59302]_  & \new_[59295]_ ;
  assign \new_[59306]_  = ~A235 & ~A233;
  assign \new_[59309]_  = A266 & A265;
  assign \new_[59310]_  = \new_[59309]_  & \new_[59306]_ ;
  assign \new_[59313]_  = ~A268 & ~A267;
  assign \new_[59316]_  = A300 & A298;
  assign \new_[59317]_  = \new_[59316]_  & \new_[59313]_ ;
  assign \new_[59318]_  = \new_[59317]_  & \new_[59310]_ ;
  assign \new_[59321]_  = A167 & A170;
  assign \new_[59324]_  = A199 & ~A166;
  assign \new_[59325]_  = \new_[59324]_  & \new_[59321]_ ;
  assign \new_[59328]_  = ~A201 & A200;
  assign \new_[59331]_  = ~A232 & ~A202;
  assign \new_[59332]_  = \new_[59331]_  & \new_[59328]_ ;
  assign \new_[59333]_  = \new_[59332]_  & \new_[59325]_ ;
  assign \new_[59336]_  = ~A235 & ~A233;
  assign \new_[59339]_  = ~A266 & ~A265;
  assign \new_[59340]_  = \new_[59339]_  & \new_[59336]_ ;
  assign \new_[59343]_  = A298 & ~A268;
  assign \new_[59346]_  = A302 & ~A299;
  assign \new_[59347]_  = \new_[59346]_  & \new_[59343]_ ;
  assign \new_[59348]_  = \new_[59347]_  & \new_[59340]_ ;
  assign \new_[59351]_  = A167 & A170;
  assign \new_[59354]_  = A199 & ~A166;
  assign \new_[59355]_  = \new_[59354]_  & \new_[59351]_ ;
  assign \new_[59358]_  = ~A201 & A200;
  assign \new_[59361]_  = ~A232 & ~A202;
  assign \new_[59362]_  = \new_[59361]_  & \new_[59358]_ ;
  assign \new_[59363]_  = \new_[59362]_  & \new_[59355]_ ;
  assign \new_[59366]_  = ~A235 & ~A233;
  assign \new_[59369]_  = ~A266 & ~A265;
  assign \new_[59370]_  = \new_[59369]_  & \new_[59366]_ ;
  assign \new_[59373]_  = ~A298 & ~A268;
  assign \new_[59376]_  = A302 & A299;
  assign \new_[59377]_  = \new_[59376]_  & \new_[59373]_ ;
  assign \new_[59378]_  = \new_[59377]_  & \new_[59370]_ ;
  assign \new_[59381]_  = A167 & A170;
  assign \new_[59384]_  = ~A199 & ~A166;
  assign \new_[59385]_  = \new_[59384]_  & \new_[59381]_ ;
  assign \new_[59388]_  = ~A202 & ~A200;
  assign \new_[59391]_  = ~A235 & ~A234;
  assign \new_[59392]_  = \new_[59391]_  & \new_[59388]_ ;
  assign \new_[59393]_  = \new_[59392]_  & \new_[59385]_ ;
  assign \new_[59396]_  = A265 & ~A236;
  assign \new_[59399]_  = ~A267 & A266;
  assign \new_[59400]_  = \new_[59399]_  & \new_[59396]_ ;
  assign \new_[59403]_  = A298 & ~A268;
  assign \new_[59406]_  = A302 & ~A299;
  assign \new_[59407]_  = \new_[59406]_  & \new_[59403]_ ;
  assign \new_[59408]_  = \new_[59407]_  & \new_[59400]_ ;
  assign \new_[59411]_  = A167 & A170;
  assign \new_[59414]_  = ~A199 & ~A166;
  assign \new_[59415]_  = \new_[59414]_  & \new_[59411]_ ;
  assign \new_[59418]_  = ~A202 & ~A200;
  assign \new_[59421]_  = ~A235 & ~A234;
  assign \new_[59422]_  = \new_[59421]_  & \new_[59418]_ ;
  assign \new_[59423]_  = \new_[59422]_  & \new_[59415]_ ;
  assign \new_[59426]_  = A265 & ~A236;
  assign \new_[59429]_  = ~A267 & A266;
  assign \new_[59430]_  = \new_[59429]_  & \new_[59426]_ ;
  assign \new_[59433]_  = ~A298 & ~A268;
  assign \new_[59436]_  = A302 & A299;
  assign \new_[59437]_  = \new_[59436]_  & \new_[59433]_ ;
  assign \new_[59438]_  = \new_[59437]_  & \new_[59430]_ ;
  assign \new_[59441]_  = A167 & A170;
  assign \new_[59444]_  = ~A199 & ~A166;
  assign \new_[59445]_  = \new_[59444]_  & \new_[59441]_ ;
  assign \new_[59448]_  = ~A202 & ~A200;
  assign \new_[59451]_  = A233 & A232;
  assign \new_[59452]_  = \new_[59451]_  & \new_[59448]_ ;
  assign \new_[59453]_  = \new_[59452]_  & \new_[59445]_ ;
  assign \new_[59456]_  = ~A235 & ~A234;
  assign \new_[59459]_  = ~A268 & ~A267;
  assign \new_[59460]_  = \new_[59459]_  & \new_[59456]_ ;
  assign \new_[59463]_  = A298 & ~A269;
  assign \new_[59466]_  = A302 & ~A299;
  assign \new_[59467]_  = \new_[59466]_  & \new_[59463]_ ;
  assign \new_[59468]_  = \new_[59467]_  & \new_[59460]_ ;
  assign \new_[59471]_  = A167 & A170;
  assign \new_[59474]_  = ~A199 & ~A166;
  assign \new_[59475]_  = \new_[59474]_  & \new_[59471]_ ;
  assign \new_[59478]_  = ~A202 & ~A200;
  assign \new_[59481]_  = A233 & A232;
  assign \new_[59482]_  = \new_[59481]_  & \new_[59478]_ ;
  assign \new_[59483]_  = \new_[59482]_  & \new_[59475]_ ;
  assign \new_[59486]_  = ~A235 & ~A234;
  assign \new_[59489]_  = ~A268 & ~A267;
  assign \new_[59490]_  = \new_[59489]_  & \new_[59486]_ ;
  assign \new_[59493]_  = ~A298 & ~A269;
  assign \new_[59496]_  = A302 & A299;
  assign \new_[59497]_  = \new_[59496]_  & \new_[59493]_ ;
  assign \new_[59498]_  = \new_[59497]_  & \new_[59490]_ ;
  assign \new_[59501]_  = A167 & A170;
  assign \new_[59504]_  = ~A199 & ~A166;
  assign \new_[59505]_  = \new_[59504]_  & \new_[59501]_ ;
  assign \new_[59508]_  = ~A202 & ~A200;
  assign \new_[59511]_  = A233 & A232;
  assign \new_[59512]_  = \new_[59511]_  & \new_[59508]_ ;
  assign \new_[59513]_  = \new_[59512]_  & \new_[59505]_ ;
  assign \new_[59516]_  = ~A235 & ~A234;
  assign \new_[59519]_  = A266 & A265;
  assign \new_[59520]_  = \new_[59519]_  & \new_[59516]_ ;
  assign \new_[59523]_  = ~A268 & ~A267;
  assign \new_[59526]_  = A300 & A299;
  assign \new_[59527]_  = \new_[59526]_  & \new_[59523]_ ;
  assign \new_[59528]_  = \new_[59527]_  & \new_[59520]_ ;
  assign \new_[59531]_  = A167 & A170;
  assign \new_[59534]_  = ~A199 & ~A166;
  assign \new_[59535]_  = \new_[59534]_  & \new_[59531]_ ;
  assign \new_[59538]_  = ~A202 & ~A200;
  assign \new_[59541]_  = A233 & A232;
  assign \new_[59542]_  = \new_[59541]_  & \new_[59538]_ ;
  assign \new_[59543]_  = \new_[59542]_  & \new_[59535]_ ;
  assign \new_[59546]_  = ~A235 & ~A234;
  assign \new_[59549]_  = A266 & A265;
  assign \new_[59550]_  = \new_[59549]_  & \new_[59546]_ ;
  assign \new_[59553]_  = ~A268 & ~A267;
  assign \new_[59556]_  = A300 & A298;
  assign \new_[59557]_  = \new_[59556]_  & \new_[59553]_ ;
  assign \new_[59558]_  = \new_[59557]_  & \new_[59550]_ ;
  assign \new_[59561]_  = A167 & A170;
  assign \new_[59564]_  = ~A199 & ~A166;
  assign \new_[59565]_  = \new_[59564]_  & \new_[59561]_ ;
  assign \new_[59568]_  = ~A202 & ~A200;
  assign \new_[59571]_  = A233 & A232;
  assign \new_[59572]_  = \new_[59571]_  & \new_[59568]_ ;
  assign \new_[59573]_  = \new_[59572]_  & \new_[59565]_ ;
  assign \new_[59576]_  = ~A235 & ~A234;
  assign \new_[59579]_  = ~A266 & ~A265;
  assign \new_[59580]_  = \new_[59579]_  & \new_[59576]_ ;
  assign \new_[59583]_  = A298 & ~A268;
  assign \new_[59586]_  = A302 & ~A299;
  assign \new_[59587]_  = \new_[59586]_  & \new_[59583]_ ;
  assign \new_[59588]_  = \new_[59587]_  & \new_[59580]_ ;
  assign \new_[59591]_  = A167 & A170;
  assign \new_[59594]_  = ~A199 & ~A166;
  assign \new_[59595]_  = \new_[59594]_  & \new_[59591]_ ;
  assign \new_[59598]_  = ~A202 & ~A200;
  assign \new_[59601]_  = A233 & A232;
  assign \new_[59602]_  = \new_[59601]_  & \new_[59598]_ ;
  assign \new_[59603]_  = \new_[59602]_  & \new_[59595]_ ;
  assign \new_[59606]_  = ~A235 & ~A234;
  assign \new_[59609]_  = ~A266 & ~A265;
  assign \new_[59610]_  = \new_[59609]_  & \new_[59606]_ ;
  assign \new_[59613]_  = ~A298 & ~A268;
  assign \new_[59616]_  = A302 & A299;
  assign \new_[59617]_  = \new_[59616]_  & \new_[59613]_ ;
  assign \new_[59618]_  = \new_[59617]_  & \new_[59610]_ ;
  assign \new_[59621]_  = A167 & A170;
  assign \new_[59624]_  = ~A199 & ~A166;
  assign \new_[59625]_  = \new_[59624]_  & \new_[59621]_ ;
  assign \new_[59628]_  = ~A202 & ~A200;
  assign \new_[59631]_  = ~A233 & ~A232;
  assign \new_[59632]_  = \new_[59631]_  & \new_[59628]_ ;
  assign \new_[59633]_  = \new_[59632]_  & \new_[59625]_ ;
  assign \new_[59636]_  = A265 & ~A235;
  assign \new_[59639]_  = ~A267 & A266;
  assign \new_[59640]_  = \new_[59639]_  & \new_[59636]_ ;
  assign \new_[59643]_  = A298 & ~A268;
  assign \new_[59646]_  = A302 & ~A299;
  assign \new_[59647]_  = \new_[59646]_  & \new_[59643]_ ;
  assign \new_[59648]_  = \new_[59647]_  & \new_[59640]_ ;
  assign \new_[59651]_  = A167 & A170;
  assign \new_[59654]_  = ~A199 & ~A166;
  assign \new_[59655]_  = \new_[59654]_  & \new_[59651]_ ;
  assign \new_[59658]_  = ~A202 & ~A200;
  assign \new_[59661]_  = ~A233 & ~A232;
  assign \new_[59662]_  = \new_[59661]_  & \new_[59658]_ ;
  assign \new_[59663]_  = \new_[59662]_  & \new_[59655]_ ;
  assign \new_[59666]_  = A265 & ~A235;
  assign \new_[59669]_  = ~A267 & A266;
  assign \new_[59670]_  = \new_[59669]_  & \new_[59666]_ ;
  assign \new_[59673]_  = ~A298 & ~A268;
  assign \new_[59676]_  = A302 & A299;
  assign \new_[59677]_  = \new_[59676]_  & \new_[59673]_ ;
  assign \new_[59678]_  = \new_[59677]_  & \new_[59670]_ ;
  assign \new_[59681]_  = ~A167 & A170;
  assign \new_[59684]_  = ~A201 & A166;
  assign \new_[59685]_  = \new_[59684]_  & \new_[59681]_ ;
  assign \new_[59688]_  = ~A203 & ~A202;
  assign \new_[59691]_  = ~A235 & ~A234;
  assign \new_[59692]_  = \new_[59691]_  & \new_[59688]_ ;
  assign \new_[59693]_  = \new_[59692]_  & \new_[59685]_ ;
  assign \new_[59696]_  = A265 & ~A236;
  assign \new_[59699]_  = ~A267 & A266;
  assign \new_[59700]_  = \new_[59699]_  & \new_[59696]_ ;
  assign \new_[59703]_  = A298 & ~A268;
  assign \new_[59706]_  = A302 & ~A299;
  assign \new_[59707]_  = \new_[59706]_  & \new_[59703]_ ;
  assign \new_[59708]_  = \new_[59707]_  & \new_[59700]_ ;
  assign \new_[59711]_  = ~A167 & A170;
  assign \new_[59714]_  = ~A201 & A166;
  assign \new_[59715]_  = \new_[59714]_  & \new_[59711]_ ;
  assign \new_[59718]_  = ~A203 & ~A202;
  assign \new_[59721]_  = ~A235 & ~A234;
  assign \new_[59722]_  = \new_[59721]_  & \new_[59718]_ ;
  assign \new_[59723]_  = \new_[59722]_  & \new_[59715]_ ;
  assign \new_[59726]_  = A265 & ~A236;
  assign \new_[59729]_  = ~A267 & A266;
  assign \new_[59730]_  = \new_[59729]_  & \new_[59726]_ ;
  assign \new_[59733]_  = ~A298 & ~A268;
  assign \new_[59736]_  = A302 & A299;
  assign \new_[59737]_  = \new_[59736]_  & \new_[59733]_ ;
  assign \new_[59738]_  = \new_[59737]_  & \new_[59730]_ ;
  assign \new_[59741]_  = ~A167 & A170;
  assign \new_[59744]_  = ~A201 & A166;
  assign \new_[59745]_  = \new_[59744]_  & \new_[59741]_ ;
  assign \new_[59748]_  = ~A203 & ~A202;
  assign \new_[59751]_  = A233 & A232;
  assign \new_[59752]_  = \new_[59751]_  & \new_[59748]_ ;
  assign \new_[59753]_  = \new_[59752]_  & \new_[59745]_ ;
  assign \new_[59756]_  = ~A235 & ~A234;
  assign \new_[59759]_  = ~A268 & ~A267;
  assign \new_[59760]_  = \new_[59759]_  & \new_[59756]_ ;
  assign \new_[59763]_  = A298 & ~A269;
  assign \new_[59766]_  = A302 & ~A299;
  assign \new_[59767]_  = \new_[59766]_  & \new_[59763]_ ;
  assign \new_[59768]_  = \new_[59767]_  & \new_[59760]_ ;
  assign \new_[59771]_  = ~A167 & A170;
  assign \new_[59774]_  = ~A201 & A166;
  assign \new_[59775]_  = \new_[59774]_  & \new_[59771]_ ;
  assign \new_[59778]_  = ~A203 & ~A202;
  assign \new_[59781]_  = A233 & A232;
  assign \new_[59782]_  = \new_[59781]_  & \new_[59778]_ ;
  assign \new_[59783]_  = \new_[59782]_  & \new_[59775]_ ;
  assign \new_[59786]_  = ~A235 & ~A234;
  assign \new_[59789]_  = ~A268 & ~A267;
  assign \new_[59790]_  = \new_[59789]_  & \new_[59786]_ ;
  assign \new_[59793]_  = ~A298 & ~A269;
  assign \new_[59796]_  = A302 & A299;
  assign \new_[59797]_  = \new_[59796]_  & \new_[59793]_ ;
  assign \new_[59798]_  = \new_[59797]_  & \new_[59790]_ ;
  assign \new_[59801]_  = ~A167 & A170;
  assign \new_[59804]_  = ~A201 & A166;
  assign \new_[59805]_  = \new_[59804]_  & \new_[59801]_ ;
  assign \new_[59808]_  = ~A203 & ~A202;
  assign \new_[59811]_  = A233 & A232;
  assign \new_[59812]_  = \new_[59811]_  & \new_[59808]_ ;
  assign \new_[59813]_  = \new_[59812]_  & \new_[59805]_ ;
  assign \new_[59816]_  = ~A235 & ~A234;
  assign \new_[59819]_  = A266 & A265;
  assign \new_[59820]_  = \new_[59819]_  & \new_[59816]_ ;
  assign \new_[59823]_  = ~A268 & ~A267;
  assign \new_[59826]_  = A300 & A299;
  assign \new_[59827]_  = \new_[59826]_  & \new_[59823]_ ;
  assign \new_[59828]_  = \new_[59827]_  & \new_[59820]_ ;
  assign \new_[59831]_  = ~A167 & A170;
  assign \new_[59834]_  = ~A201 & A166;
  assign \new_[59835]_  = \new_[59834]_  & \new_[59831]_ ;
  assign \new_[59838]_  = ~A203 & ~A202;
  assign \new_[59841]_  = A233 & A232;
  assign \new_[59842]_  = \new_[59841]_  & \new_[59838]_ ;
  assign \new_[59843]_  = \new_[59842]_  & \new_[59835]_ ;
  assign \new_[59846]_  = ~A235 & ~A234;
  assign \new_[59849]_  = A266 & A265;
  assign \new_[59850]_  = \new_[59849]_  & \new_[59846]_ ;
  assign \new_[59853]_  = ~A268 & ~A267;
  assign \new_[59856]_  = A300 & A298;
  assign \new_[59857]_  = \new_[59856]_  & \new_[59853]_ ;
  assign \new_[59858]_  = \new_[59857]_  & \new_[59850]_ ;
  assign \new_[59861]_  = ~A167 & A170;
  assign \new_[59864]_  = ~A201 & A166;
  assign \new_[59865]_  = \new_[59864]_  & \new_[59861]_ ;
  assign \new_[59868]_  = ~A203 & ~A202;
  assign \new_[59871]_  = A233 & A232;
  assign \new_[59872]_  = \new_[59871]_  & \new_[59868]_ ;
  assign \new_[59873]_  = \new_[59872]_  & \new_[59865]_ ;
  assign \new_[59876]_  = ~A235 & ~A234;
  assign \new_[59879]_  = ~A266 & ~A265;
  assign \new_[59880]_  = \new_[59879]_  & \new_[59876]_ ;
  assign \new_[59883]_  = A298 & ~A268;
  assign \new_[59886]_  = A302 & ~A299;
  assign \new_[59887]_  = \new_[59886]_  & \new_[59883]_ ;
  assign \new_[59888]_  = \new_[59887]_  & \new_[59880]_ ;
  assign \new_[59891]_  = ~A167 & A170;
  assign \new_[59894]_  = ~A201 & A166;
  assign \new_[59895]_  = \new_[59894]_  & \new_[59891]_ ;
  assign \new_[59898]_  = ~A203 & ~A202;
  assign \new_[59901]_  = A233 & A232;
  assign \new_[59902]_  = \new_[59901]_  & \new_[59898]_ ;
  assign \new_[59903]_  = \new_[59902]_  & \new_[59895]_ ;
  assign \new_[59906]_  = ~A235 & ~A234;
  assign \new_[59909]_  = ~A266 & ~A265;
  assign \new_[59910]_  = \new_[59909]_  & \new_[59906]_ ;
  assign \new_[59913]_  = ~A298 & ~A268;
  assign \new_[59916]_  = A302 & A299;
  assign \new_[59917]_  = \new_[59916]_  & \new_[59913]_ ;
  assign \new_[59918]_  = \new_[59917]_  & \new_[59910]_ ;
  assign \new_[59921]_  = ~A167 & A170;
  assign \new_[59924]_  = ~A201 & A166;
  assign \new_[59925]_  = \new_[59924]_  & \new_[59921]_ ;
  assign \new_[59928]_  = ~A203 & ~A202;
  assign \new_[59931]_  = ~A233 & ~A232;
  assign \new_[59932]_  = \new_[59931]_  & \new_[59928]_ ;
  assign \new_[59933]_  = \new_[59932]_  & \new_[59925]_ ;
  assign \new_[59936]_  = A265 & ~A235;
  assign \new_[59939]_  = ~A267 & A266;
  assign \new_[59940]_  = \new_[59939]_  & \new_[59936]_ ;
  assign \new_[59943]_  = A298 & ~A268;
  assign \new_[59946]_  = A302 & ~A299;
  assign \new_[59947]_  = \new_[59946]_  & \new_[59943]_ ;
  assign \new_[59948]_  = \new_[59947]_  & \new_[59940]_ ;
  assign \new_[59951]_  = ~A167 & A170;
  assign \new_[59954]_  = ~A201 & A166;
  assign \new_[59955]_  = \new_[59954]_  & \new_[59951]_ ;
  assign \new_[59958]_  = ~A203 & ~A202;
  assign \new_[59961]_  = ~A233 & ~A232;
  assign \new_[59962]_  = \new_[59961]_  & \new_[59958]_ ;
  assign \new_[59963]_  = \new_[59962]_  & \new_[59955]_ ;
  assign \new_[59966]_  = A265 & ~A235;
  assign \new_[59969]_  = ~A267 & A266;
  assign \new_[59970]_  = \new_[59969]_  & \new_[59966]_ ;
  assign \new_[59973]_  = ~A298 & ~A268;
  assign \new_[59976]_  = A302 & A299;
  assign \new_[59977]_  = \new_[59976]_  & \new_[59973]_ ;
  assign \new_[59978]_  = \new_[59977]_  & \new_[59970]_ ;
  assign \new_[59981]_  = ~A167 & A170;
  assign \new_[59984]_  = A199 & A166;
  assign \new_[59985]_  = \new_[59984]_  & \new_[59981]_ ;
  assign \new_[59988]_  = ~A201 & A200;
  assign \new_[59991]_  = ~A234 & ~A202;
  assign \new_[59992]_  = \new_[59991]_  & \new_[59988]_ ;
  assign \new_[59993]_  = \new_[59992]_  & \new_[59985]_ ;
  assign \new_[59996]_  = ~A236 & ~A235;
  assign \new_[59999]_  = ~A268 & ~A267;
  assign \new_[60000]_  = \new_[59999]_  & \new_[59996]_ ;
  assign \new_[60003]_  = A298 & ~A269;
  assign \new_[60006]_  = A302 & ~A299;
  assign \new_[60007]_  = \new_[60006]_  & \new_[60003]_ ;
  assign \new_[60008]_  = \new_[60007]_  & \new_[60000]_ ;
  assign \new_[60011]_  = ~A167 & A170;
  assign \new_[60014]_  = A199 & A166;
  assign \new_[60015]_  = \new_[60014]_  & \new_[60011]_ ;
  assign \new_[60018]_  = ~A201 & A200;
  assign \new_[60021]_  = ~A234 & ~A202;
  assign \new_[60022]_  = \new_[60021]_  & \new_[60018]_ ;
  assign \new_[60023]_  = \new_[60022]_  & \new_[60015]_ ;
  assign \new_[60026]_  = ~A236 & ~A235;
  assign \new_[60029]_  = ~A268 & ~A267;
  assign \new_[60030]_  = \new_[60029]_  & \new_[60026]_ ;
  assign \new_[60033]_  = ~A298 & ~A269;
  assign \new_[60036]_  = A302 & A299;
  assign \new_[60037]_  = \new_[60036]_  & \new_[60033]_ ;
  assign \new_[60038]_  = \new_[60037]_  & \new_[60030]_ ;
  assign \new_[60041]_  = ~A167 & A170;
  assign \new_[60044]_  = A199 & A166;
  assign \new_[60045]_  = \new_[60044]_  & \new_[60041]_ ;
  assign \new_[60048]_  = ~A201 & A200;
  assign \new_[60051]_  = ~A234 & ~A202;
  assign \new_[60052]_  = \new_[60051]_  & \new_[60048]_ ;
  assign \new_[60053]_  = \new_[60052]_  & \new_[60045]_ ;
  assign \new_[60056]_  = ~A236 & ~A235;
  assign \new_[60059]_  = A266 & A265;
  assign \new_[60060]_  = \new_[60059]_  & \new_[60056]_ ;
  assign \new_[60063]_  = ~A268 & ~A267;
  assign \new_[60066]_  = A300 & A299;
  assign \new_[60067]_  = \new_[60066]_  & \new_[60063]_ ;
  assign \new_[60068]_  = \new_[60067]_  & \new_[60060]_ ;
  assign \new_[60071]_  = ~A167 & A170;
  assign \new_[60074]_  = A199 & A166;
  assign \new_[60075]_  = \new_[60074]_  & \new_[60071]_ ;
  assign \new_[60078]_  = ~A201 & A200;
  assign \new_[60081]_  = ~A234 & ~A202;
  assign \new_[60082]_  = \new_[60081]_  & \new_[60078]_ ;
  assign \new_[60083]_  = \new_[60082]_  & \new_[60075]_ ;
  assign \new_[60086]_  = ~A236 & ~A235;
  assign \new_[60089]_  = A266 & A265;
  assign \new_[60090]_  = \new_[60089]_  & \new_[60086]_ ;
  assign \new_[60093]_  = ~A268 & ~A267;
  assign \new_[60096]_  = A300 & A298;
  assign \new_[60097]_  = \new_[60096]_  & \new_[60093]_ ;
  assign \new_[60098]_  = \new_[60097]_  & \new_[60090]_ ;
  assign \new_[60101]_  = ~A167 & A170;
  assign \new_[60104]_  = A199 & A166;
  assign \new_[60105]_  = \new_[60104]_  & \new_[60101]_ ;
  assign \new_[60108]_  = ~A201 & A200;
  assign \new_[60111]_  = ~A234 & ~A202;
  assign \new_[60112]_  = \new_[60111]_  & \new_[60108]_ ;
  assign \new_[60113]_  = \new_[60112]_  & \new_[60105]_ ;
  assign \new_[60116]_  = ~A236 & ~A235;
  assign \new_[60119]_  = ~A266 & ~A265;
  assign \new_[60120]_  = \new_[60119]_  & \new_[60116]_ ;
  assign \new_[60123]_  = A298 & ~A268;
  assign \new_[60126]_  = A302 & ~A299;
  assign \new_[60127]_  = \new_[60126]_  & \new_[60123]_ ;
  assign \new_[60128]_  = \new_[60127]_  & \new_[60120]_ ;
  assign \new_[60131]_  = ~A167 & A170;
  assign \new_[60134]_  = A199 & A166;
  assign \new_[60135]_  = \new_[60134]_  & \new_[60131]_ ;
  assign \new_[60138]_  = ~A201 & A200;
  assign \new_[60141]_  = ~A234 & ~A202;
  assign \new_[60142]_  = \new_[60141]_  & \new_[60138]_ ;
  assign \new_[60143]_  = \new_[60142]_  & \new_[60135]_ ;
  assign \new_[60146]_  = ~A236 & ~A235;
  assign \new_[60149]_  = ~A266 & ~A265;
  assign \new_[60150]_  = \new_[60149]_  & \new_[60146]_ ;
  assign \new_[60153]_  = ~A298 & ~A268;
  assign \new_[60156]_  = A302 & A299;
  assign \new_[60157]_  = \new_[60156]_  & \new_[60153]_ ;
  assign \new_[60158]_  = \new_[60157]_  & \new_[60150]_ ;
  assign \new_[60161]_  = ~A167 & A170;
  assign \new_[60164]_  = A199 & A166;
  assign \new_[60165]_  = \new_[60164]_  & \new_[60161]_ ;
  assign \new_[60168]_  = ~A201 & A200;
  assign \new_[60171]_  = A232 & ~A202;
  assign \new_[60172]_  = \new_[60171]_  & \new_[60168]_ ;
  assign \new_[60173]_  = \new_[60172]_  & \new_[60165]_ ;
  assign \new_[60176]_  = ~A234 & A233;
  assign \new_[60179]_  = ~A267 & ~A235;
  assign \new_[60180]_  = \new_[60179]_  & \new_[60176]_ ;
  assign \new_[60183]_  = ~A269 & ~A268;
  assign \new_[60186]_  = A300 & A299;
  assign \new_[60187]_  = \new_[60186]_  & \new_[60183]_ ;
  assign \new_[60188]_  = \new_[60187]_  & \new_[60180]_ ;
  assign \new_[60191]_  = ~A167 & A170;
  assign \new_[60194]_  = A199 & A166;
  assign \new_[60195]_  = \new_[60194]_  & \new_[60191]_ ;
  assign \new_[60198]_  = ~A201 & A200;
  assign \new_[60201]_  = A232 & ~A202;
  assign \new_[60202]_  = \new_[60201]_  & \new_[60198]_ ;
  assign \new_[60203]_  = \new_[60202]_  & \new_[60195]_ ;
  assign \new_[60206]_  = ~A234 & A233;
  assign \new_[60209]_  = ~A267 & ~A235;
  assign \new_[60210]_  = \new_[60209]_  & \new_[60206]_ ;
  assign \new_[60213]_  = ~A269 & ~A268;
  assign \new_[60216]_  = A300 & A298;
  assign \new_[60217]_  = \new_[60216]_  & \new_[60213]_ ;
  assign \new_[60218]_  = \new_[60217]_  & \new_[60210]_ ;
  assign \new_[60221]_  = ~A167 & A170;
  assign \new_[60224]_  = A199 & A166;
  assign \new_[60225]_  = \new_[60224]_  & \new_[60221]_ ;
  assign \new_[60228]_  = ~A201 & A200;
  assign \new_[60231]_  = A232 & ~A202;
  assign \new_[60232]_  = \new_[60231]_  & \new_[60228]_ ;
  assign \new_[60233]_  = \new_[60232]_  & \new_[60225]_ ;
  assign \new_[60236]_  = ~A234 & A233;
  assign \new_[60239]_  = A265 & ~A235;
  assign \new_[60240]_  = \new_[60239]_  & \new_[60236]_ ;
  assign \new_[60243]_  = ~A267 & A266;
  assign \new_[60246]_  = A301 & ~A268;
  assign \new_[60247]_  = \new_[60246]_  & \new_[60243]_ ;
  assign \new_[60248]_  = \new_[60247]_  & \new_[60240]_ ;
  assign \new_[60251]_  = ~A167 & A170;
  assign \new_[60254]_  = A199 & A166;
  assign \new_[60255]_  = \new_[60254]_  & \new_[60251]_ ;
  assign \new_[60258]_  = ~A201 & A200;
  assign \new_[60261]_  = A232 & ~A202;
  assign \new_[60262]_  = \new_[60261]_  & \new_[60258]_ ;
  assign \new_[60263]_  = \new_[60262]_  & \new_[60255]_ ;
  assign \new_[60266]_  = ~A234 & A233;
  assign \new_[60269]_  = ~A265 & ~A235;
  assign \new_[60270]_  = \new_[60269]_  & \new_[60266]_ ;
  assign \new_[60273]_  = ~A268 & ~A266;
  assign \new_[60276]_  = A300 & A299;
  assign \new_[60277]_  = \new_[60276]_  & \new_[60273]_ ;
  assign \new_[60278]_  = \new_[60277]_  & \new_[60270]_ ;
  assign \new_[60281]_  = ~A167 & A170;
  assign \new_[60284]_  = A199 & A166;
  assign \new_[60285]_  = \new_[60284]_  & \new_[60281]_ ;
  assign \new_[60288]_  = ~A201 & A200;
  assign \new_[60291]_  = A232 & ~A202;
  assign \new_[60292]_  = \new_[60291]_  & \new_[60288]_ ;
  assign \new_[60293]_  = \new_[60292]_  & \new_[60285]_ ;
  assign \new_[60296]_  = ~A234 & A233;
  assign \new_[60299]_  = ~A265 & ~A235;
  assign \new_[60300]_  = \new_[60299]_  & \new_[60296]_ ;
  assign \new_[60303]_  = ~A268 & ~A266;
  assign \new_[60306]_  = A300 & A298;
  assign \new_[60307]_  = \new_[60306]_  & \new_[60303]_ ;
  assign \new_[60308]_  = \new_[60307]_  & \new_[60300]_ ;
  assign \new_[60311]_  = ~A167 & A170;
  assign \new_[60314]_  = A199 & A166;
  assign \new_[60315]_  = \new_[60314]_  & \new_[60311]_ ;
  assign \new_[60318]_  = ~A201 & A200;
  assign \new_[60321]_  = ~A232 & ~A202;
  assign \new_[60322]_  = \new_[60321]_  & \new_[60318]_ ;
  assign \new_[60323]_  = \new_[60322]_  & \new_[60315]_ ;
  assign \new_[60326]_  = ~A235 & ~A233;
  assign \new_[60329]_  = ~A268 & ~A267;
  assign \new_[60330]_  = \new_[60329]_  & \new_[60326]_ ;
  assign \new_[60333]_  = A298 & ~A269;
  assign \new_[60336]_  = A302 & ~A299;
  assign \new_[60337]_  = \new_[60336]_  & \new_[60333]_ ;
  assign \new_[60338]_  = \new_[60337]_  & \new_[60330]_ ;
  assign \new_[60341]_  = ~A167 & A170;
  assign \new_[60344]_  = A199 & A166;
  assign \new_[60345]_  = \new_[60344]_  & \new_[60341]_ ;
  assign \new_[60348]_  = ~A201 & A200;
  assign \new_[60351]_  = ~A232 & ~A202;
  assign \new_[60352]_  = \new_[60351]_  & \new_[60348]_ ;
  assign \new_[60353]_  = \new_[60352]_  & \new_[60345]_ ;
  assign \new_[60356]_  = ~A235 & ~A233;
  assign \new_[60359]_  = ~A268 & ~A267;
  assign \new_[60360]_  = \new_[60359]_  & \new_[60356]_ ;
  assign \new_[60363]_  = ~A298 & ~A269;
  assign \new_[60366]_  = A302 & A299;
  assign \new_[60367]_  = \new_[60366]_  & \new_[60363]_ ;
  assign \new_[60368]_  = \new_[60367]_  & \new_[60360]_ ;
  assign \new_[60371]_  = ~A167 & A170;
  assign \new_[60374]_  = A199 & A166;
  assign \new_[60375]_  = \new_[60374]_  & \new_[60371]_ ;
  assign \new_[60378]_  = ~A201 & A200;
  assign \new_[60381]_  = ~A232 & ~A202;
  assign \new_[60382]_  = \new_[60381]_  & \new_[60378]_ ;
  assign \new_[60383]_  = \new_[60382]_  & \new_[60375]_ ;
  assign \new_[60386]_  = ~A235 & ~A233;
  assign \new_[60389]_  = A266 & A265;
  assign \new_[60390]_  = \new_[60389]_  & \new_[60386]_ ;
  assign \new_[60393]_  = ~A268 & ~A267;
  assign \new_[60396]_  = A300 & A299;
  assign \new_[60397]_  = \new_[60396]_  & \new_[60393]_ ;
  assign \new_[60398]_  = \new_[60397]_  & \new_[60390]_ ;
  assign \new_[60401]_  = ~A167 & A170;
  assign \new_[60404]_  = A199 & A166;
  assign \new_[60405]_  = \new_[60404]_  & \new_[60401]_ ;
  assign \new_[60408]_  = ~A201 & A200;
  assign \new_[60411]_  = ~A232 & ~A202;
  assign \new_[60412]_  = \new_[60411]_  & \new_[60408]_ ;
  assign \new_[60413]_  = \new_[60412]_  & \new_[60405]_ ;
  assign \new_[60416]_  = ~A235 & ~A233;
  assign \new_[60419]_  = A266 & A265;
  assign \new_[60420]_  = \new_[60419]_  & \new_[60416]_ ;
  assign \new_[60423]_  = ~A268 & ~A267;
  assign \new_[60426]_  = A300 & A298;
  assign \new_[60427]_  = \new_[60426]_  & \new_[60423]_ ;
  assign \new_[60428]_  = \new_[60427]_  & \new_[60420]_ ;
  assign \new_[60431]_  = ~A167 & A170;
  assign \new_[60434]_  = A199 & A166;
  assign \new_[60435]_  = \new_[60434]_  & \new_[60431]_ ;
  assign \new_[60438]_  = ~A201 & A200;
  assign \new_[60441]_  = ~A232 & ~A202;
  assign \new_[60442]_  = \new_[60441]_  & \new_[60438]_ ;
  assign \new_[60443]_  = \new_[60442]_  & \new_[60435]_ ;
  assign \new_[60446]_  = ~A235 & ~A233;
  assign \new_[60449]_  = ~A266 & ~A265;
  assign \new_[60450]_  = \new_[60449]_  & \new_[60446]_ ;
  assign \new_[60453]_  = A298 & ~A268;
  assign \new_[60456]_  = A302 & ~A299;
  assign \new_[60457]_  = \new_[60456]_  & \new_[60453]_ ;
  assign \new_[60458]_  = \new_[60457]_  & \new_[60450]_ ;
  assign \new_[60461]_  = ~A167 & A170;
  assign \new_[60464]_  = A199 & A166;
  assign \new_[60465]_  = \new_[60464]_  & \new_[60461]_ ;
  assign \new_[60468]_  = ~A201 & A200;
  assign \new_[60471]_  = ~A232 & ~A202;
  assign \new_[60472]_  = \new_[60471]_  & \new_[60468]_ ;
  assign \new_[60473]_  = \new_[60472]_  & \new_[60465]_ ;
  assign \new_[60476]_  = ~A235 & ~A233;
  assign \new_[60479]_  = ~A266 & ~A265;
  assign \new_[60480]_  = \new_[60479]_  & \new_[60476]_ ;
  assign \new_[60483]_  = ~A298 & ~A268;
  assign \new_[60486]_  = A302 & A299;
  assign \new_[60487]_  = \new_[60486]_  & \new_[60483]_ ;
  assign \new_[60488]_  = \new_[60487]_  & \new_[60480]_ ;
  assign \new_[60491]_  = ~A167 & A170;
  assign \new_[60494]_  = ~A199 & A166;
  assign \new_[60495]_  = \new_[60494]_  & \new_[60491]_ ;
  assign \new_[60498]_  = ~A202 & ~A200;
  assign \new_[60501]_  = ~A235 & ~A234;
  assign \new_[60502]_  = \new_[60501]_  & \new_[60498]_ ;
  assign \new_[60503]_  = \new_[60502]_  & \new_[60495]_ ;
  assign \new_[60506]_  = A265 & ~A236;
  assign \new_[60509]_  = ~A267 & A266;
  assign \new_[60510]_  = \new_[60509]_  & \new_[60506]_ ;
  assign \new_[60513]_  = A298 & ~A268;
  assign \new_[60516]_  = A302 & ~A299;
  assign \new_[60517]_  = \new_[60516]_  & \new_[60513]_ ;
  assign \new_[60518]_  = \new_[60517]_  & \new_[60510]_ ;
  assign \new_[60521]_  = ~A167 & A170;
  assign \new_[60524]_  = ~A199 & A166;
  assign \new_[60525]_  = \new_[60524]_  & \new_[60521]_ ;
  assign \new_[60528]_  = ~A202 & ~A200;
  assign \new_[60531]_  = ~A235 & ~A234;
  assign \new_[60532]_  = \new_[60531]_  & \new_[60528]_ ;
  assign \new_[60533]_  = \new_[60532]_  & \new_[60525]_ ;
  assign \new_[60536]_  = A265 & ~A236;
  assign \new_[60539]_  = ~A267 & A266;
  assign \new_[60540]_  = \new_[60539]_  & \new_[60536]_ ;
  assign \new_[60543]_  = ~A298 & ~A268;
  assign \new_[60546]_  = A302 & A299;
  assign \new_[60547]_  = \new_[60546]_  & \new_[60543]_ ;
  assign \new_[60548]_  = \new_[60547]_  & \new_[60540]_ ;
  assign \new_[60551]_  = ~A167 & A170;
  assign \new_[60554]_  = ~A199 & A166;
  assign \new_[60555]_  = \new_[60554]_  & \new_[60551]_ ;
  assign \new_[60558]_  = ~A202 & ~A200;
  assign \new_[60561]_  = A233 & A232;
  assign \new_[60562]_  = \new_[60561]_  & \new_[60558]_ ;
  assign \new_[60563]_  = \new_[60562]_  & \new_[60555]_ ;
  assign \new_[60566]_  = ~A235 & ~A234;
  assign \new_[60569]_  = ~A268 & ~A267;
  assign \new_[60570]_  = \new_[60569]_  & \new_[60566]_ ;
  assign \new_[60573]_  = A298 & ~A269;
  assign \new_[60576]_  = A302 & ~A299;
  assign \new_[60577]_  = \new_[60576]_  & \new_[60573]_ ;
  assign \new_[60578]_  = \new_[60577]_  & \new_[60570]_ ;
  assign \new_[60581]_  = ~A167 & A170;
  assign \new_[60584]_  = ~A199 & A166;
  assign \new_[60585]_  = \new_[60584]_  & \new_[60581]_ ;
  assign \new_[60588]_  = ~A202 & ~A200;
  assign \new_[60591]_  = A233 & A232;
  assign \new_[60592]_  = \new_[60591]_  & \new_[60588]_ ;
  assign \new_[60593]_  = \new_[60592]_  & \new_[60585]_ ;
  assign \new_[60596]_  = ~A235 & ~A234;
  assign \new_[60599]_  = ~A268 & ~A267;
  assign \new_[60600]_  = \new_[60599]_  & \new_[60596]_ ;
  assign \new_[60603]_  = ~A298 & ~A269;
  assign \new_[60606]_  = A302 & A299;
  assign \new_[60607]_  = \new_[60606]_  & \new_[60603]_ ;
  assign \new_[60608]_  = \new_[60607]_  & \new_[60600]_ ;
  assign \new_[60611]_  = ~A167 & A170;
  assign \new_[60614]_  = ~A199 & A166;
  assign \new_[60615]_  = \new_[60614]_  & \new_[60611]_ ;
  assign \new_[60618]_  = ~A202 & ~A200;
  assign \new_[60621]_  = A233 & A232;
  assign \new_[60622]_  = \new_[60621]_  & \new_[60618]_ ;
  assign \new_[60623]_  = \new_[60622]_  & \new_[60615]_ ;
  assign \new_[60626]_  = ~A235 & ~A234;
  assign \new_[60629]_  = A266 & A265;
  assign \new_[60630]_  = \new_[60629]_  & \new_[60626]_ ;
  assign \new_[60633]_  = ~A268 & ~A267;
  assign \new_[60636]_  = A300 & A299;
  assign \new_[60637]_  = \new_[60636]_  & \new_[60633]_ ;
  assign \new_[60638]_  = \new_[60637]_  & \new_[60630]_ ;
  assign \new_[60641]_  = ~A167 & A170;
  assign \new_[60644]_  = ~A199 & A166;
  assign \new_[60645]_  = \new_[60644]_  & \new_[60641]_ ;
  assign \new_[60648]_  = ~A202 & ~A200;
  assign \new_[60651]_  = A233 & A232;
  assign \new_[60652]_  = \new_[60651]_  & \new_[60648]_ ;
  assign \new_[60653]_  = \new_[60652]_  & \new_[60645]_ ;
  assign \new_[60656]_  = ~A235 & ~A234;
  assign \new_[60659]_  = A266 & A265;
  assign \new_[60660]_  = \new_[60659]_  & \new_[60656]_ ;
  assign \new_[60663]_  = ~A268 & ~A267;
  assign \new_[60666]_  = A300 & A298;
  assign \new_[60667]_  = \new_[60666]_  & \new_[60663]_ ;
  assign \new_[60668]_  = \new_[60667]_  & \new_[60660]_ ;
  assign \new_[60671]_  = ~A167 & A170;
  assign \new_[60674]_  = ~A199 & A166;
  assign \new_[60675]_  = \new_[60674]_  & \new_[60671]_ ;
  assign \new_[60678]_  = ~A202 & ~A200;
  assign \new_[60681]_  = A233 & A232;
  assign \new_[60682]_  = \new_[60681]_  & \new_[60678]_ ;
  assign \new_[60683]_  = \new_[60682]_  & \new_[60675]_ ;
  assign \new_[60686]_  = ~A235 & ~A234;
  assign \new_[60689]_  = ~A266 & ~A265;
  assign \new_[60690]_  = \new_[60689]_  & \new_[60686]_ ;
  assign \new_[60693]_  = A298 & ~A268;
  assign \new_[60696]_  = A302 & ~A299;
  assign \new_[60697]_  = \new_[60696]_  & \new_[60693]_ ;
  assign \new_[60698]_  = \new_[60697]_  & \new_[60690]_ ;
  assign \new_[60701]_  = ~A167 & A170;
  assign \new_[60704]_  = ~A199 & A166;
  assign \new_[60705]_  = \new_[60704]_  & \new_[60701]_ ;
  assign \new_[60708]_  = ~A202 & ~A200;
  assign \new_[60711]_  = A233 & A232;
  assign \new_[60712]_  = \new_[60711]_  & \new_[60708]_ ;
  assign \new_[60713]_  = \new_[60712]_  & \new_[60705]_ ;
  assign \new_[60716]_  = ~A235 & ~A234;
  assign \new_[60719]_  = ~A266 & ~A265;
  assign \new_[60720]_  = \new_[60719]_  & \new_[60716]_ ;
  assign \new_[60723]_  = ~A298 & ~A268;
  assign \new_[60726]_  = A302 & A299;
  assign \new_[60727]_  = \new_[60726]_  & \new_[60723]_ ;
  assign \new_[60728]_  = \new_[60727]_  & \new_[60720]_ ;
  assign \new_[60731]_  = ~A167 & A170;
  assign \new_[60734]_  = ~A199 & A166;
  assign \new_[60735]_  = \new_[60734]_  & \new_[60731]_ ;
  assign \new_[60738]_  = ~A202 & ~A200;
  assign \new_[60741]_  = ~A233 & ~A232;
  assign \new_[60742]_  = \new_[60741]_  & \new_[60738]_ ;
  assign \new_[60743]_  = \new_[60742]_  & \new_[60735]_ ;
  assign \new_[60746]_  = A265 & ~A235;
  assign \new_[60749]_  = ~A267 & A266;
  assign \new_[60750]_  = \new_[60749]_  & \new_[60746]_ ;
  assign \new_[60753]_  = A298 & ~A268;
  assign \new_[60756]_  = A302 & ~A299;
  assign \new_[60757]_  = \new_[60756]_  & \new_[60753]_ ;
  assign \new_[60758]_  = \new_[60757]_  & \new_[60750]_ ;
  assign \new_[60761]_  = ~A167 & A170;
  assign \new_[60764]_  = ~A199 & A166;
  assign \new_[60765]_  = \new_[60764]_  & \new_[60761]_ ;
  assign \new_[60768]_  = ~A202 & ~A200;
  assign \new_[60771]_  = ~A233 & ~A232;
  assign \new_[60772]_  = \new_[60771]_  & \new_[60768]_ ;
  assign \new_[60773]_  = \new_[60772]_  & \new_[60765]_ ;
  assign \new_[60776]_  = A265 & ~A235;
  assign \new_[60779]_  = ~A267 & A266;
  assign \new_[60780]_  = \new_[60779]_  & \new_[60776]_ ;
  assign \new_[60783]_  = ~A298 & ~A268;
  assign \new_[60786]_  = A302 & A299;
  assign \new_[60787]_  = \new_[60786]_  & \new_[60783]_ ;
  assign \new_[60788]_  = \new_[60787]_  & \new_[60780]_ ;
  assign \new_[60791]_  = A199 & A169;
  assign \new_[60794]_  = ~A201 & A200;
  assign \new_[60795]_  = \new_[60794]_  & \new_[60791]_ ;
  assign \new_[60798]_  = A232 & ~A202;
  assign \new_[60801]_  = ~A234 & A233;
  assign \new_[60802]_  = \new_[60801]_  & \new_[60798]_ ;
  assign \new_[60803]_  = \new_[60802]_  & \new_[60795]_ ;
  assign \new_[60806]_  = A265 & ~A235;
  assign \new_[60809]_  = ~A267 & A266;
  assign \new_[60810]_  = \new_[60809]_  & \new_[60806]_ ;
  assign \new_[60813]_  = A298 & ~A268;
  assign \new_[60816]_  = A302 & ~A299;
  assign \new_[60817]_  = \new_[60816]_  & \new_[60813]_ ;
  assign \new_[60818]_  = \new_[60817]_  & \new_[60810]_ ;
  assign \new_[60821]_  = A199 & A169;
  assign \new_[60824]_  = ~A201 & A200;
  assign \new_[60825]_  = \new_[60824]_  & \new_[60821]_ ;
  assign \new_[60828]_  = A232 & ~A202;
  assign \new_[60831]_  = ~A234 & A233;
  assign \new_[60832]_  = \new_[60831]_  & \new_[60828]_ ;
  assign \new_[60833]_  = \new_[60832]_  & \new_[60825]_ ;
  assign \new_[60836]_  = A265 & ~A235;
  assign \new_[60839]_  = ~A267 & A266;
  assign \new_[60840]_  = \new_[60839]_  & \new_[60836]_ ;
  assign \new_[60843]_  = ~A298 & ~A268;
  assign \new_[60846]_  = A302 & A299;
  assign \new_[60847]_  = \new_[60846]_  & \new_[60843]_ ;
  assign \new_[60848]_  = \new_[60847]_  & \new_[60840]_ ;
  assign \new_[60851]_  = ~A167 & ~A169;
  assign \new_[60854]_  = A199 & ~A166;
  assign \new_[60855]_  = \new_[60854]_  & \new_[60851]_ ;
  assign \new_[60858]_  = A232 & A201;
  assign \new_[60861]_  = ~A234 & A233;
  assign \new_[60862]_  = \new_[60861]_  & \new_[60858]_ ;
  assign \new_[60863]_  = \new_[60862]_  & \new_[60855]_ ;
  assign \new_[60866]_  = A265 & ~A235;
  assign \new_[60869]_  = ~A267 & A266;
  assign \new_[60870]_  = \new_[60869]_  & \new_[60866]_ ;
  assign \new_[60873]_  = A298 & ~A268;
  assign \new_[60876]_  = A302 & ~A299;
  assign \new_[60877]_  = \new_[60876]_  & \new_[60873]_ ;
  assign \new_[60878]_  = \new_[60877]_  & \new_[60870]_ ;
  assign \new_[60881]_  = ~A167 & ~A169;
  assign \new_[60884]_  = A199 & ~A166;
  assign \new_[60885]_  = \new_[60884]_  & \new_[60881]_ ;
  assign \new_[60888]_  = A232 & A201;
  assign \new_[60891]_  = ~A234 & A233;
  assign \new_[60892]_  = \new_[60891]_  & \new_[60888]_ ;
  assign \new_[60893]_  = \new_[60892]_  & \new_[60885]_ ;
  assign \new_[60896]_  = A265 & ~A235;
  assign \new_[60899]_  = ~A267 & A266;
  assign \new_[60900]_  = \new_[60899]_  & \new_[60896]_ ;
  assign \new_[60903]_  = ~A298 & ~A268;
  assign \new_[60906]_  = A302 & A299;
  assign \new_[60907]_  = \new_[60906]_  & \new_[60903]_ ;
  assign \new_[60908]_  = \new_[60907]_  & \new_[60900]_ ;
  assign \new_[60911]_  = ~A167 & ~A169;
  assign \new_[60914]_  = A200 & ~A166;
  assign \new_[60915]_  = \new_[60914]_  & \new_[60911]_ ;
  assign \new_[60918]_  = A232 & A201;
  assign \new_[60921]_  = ~A234 & A233;
  assign \new_[60922]_  = \new_[60921]_  & \new_[60918]_ ;
  assign \new_[60923]_  = \new_[60922]_  & \new_[60915]_ ;
  assign \new_[60926]_  = A265 & ~A235;
  assign \new_[60929]_  = ~A267 & A266;
  assign \new_[60930]_  = \new_[60929]_  & \new_[60926]_ ;
  assign \new_[60933]_  = A298 & ~A268;
  assign \new_[60936]_  = A302 & ~A299;
  assign \new_[60937]_  = \new_[60936]_  & \new_[60933]_ ;
  assign \new_[60938]_  = \new_[60937]_  & \new_[60930]_ ;
  assign \new_[60941]_  = ~A167 & ~A169;
  assign \new_[60944]_  = A200 & ~A166;
  assign \new_[60945]_  = \new_[60944]_  & \new_[60941]_ ;
  assign \new_[60948]_  = A232 & A201;
  assign \new_[60951]_  = ~A234 & A233;
  assign \new_[60952]_  = \new_[60951]_  & \new_[60948]_ ;
  assign \new_[60953]_  = \new_[60952]_  & \new_[60945]_ ;
  assign \new_[60956]_  = A265 & ~A235;
  assign \new_[60959]_  = ~A267 & A266;
  assign \new_[60960]_  = \new_[60959]_  & \new_[60956]_ ;
  assign \new_[60963]_  = ~A298 & ~A268;
  assign \new_[60966]_  = A302 & A299;
  assign \new_[60967]_  = \new_[60966]_  & \new_[60963]_ ;
  assign \new_[60968]_  = \new_[60967]_  & \new_[60960]_ ;
  assign \new_[60971]_  = ~A167 & ~A169;
  assign \new_[60974]_  = ~A199 & ~A166;
  assign \new_[60975]_  = \new_[60974]_  & \new_[60971]_ ;
  assign \new_[60978]_  = A203 & A200;
  assign \new_[60981]_  = ~A235 & ~A234;
  assign \new_[60982]_  = \new_[60981]_  & \new_[60978]_ ;
  assign \new_[60983]_  = \new_[60982]_  & \new_[60975]_ ;
  assign \new_[60986]_  = A265 & ~A236;
  assign \new_[60989]_  = ~A267 & A266;
  assign \new_[60990]_  = \new_[60989]_  & \new_[60986]_ ;
  assign \new_[60993]_  = A298 & ~A268;
  assign \new_[60996]_  = A302 & ~A299;
  assign \new_[60997]_  = \new_[60996]_  & \new_[60993]_ ;
  assign \new_[60998]_  = \new_[60997]_  & \new_[60990]_ ;
  assign \new_[61001]_  = ~A167 & ~A169;
  assign \new_[61004]_  = ~A199 & ~A166;
  assign \new_[61005]_  = \new_[61004]_  & \new_[61001]_ ;
  assign \new_[61008]_  = A203 & A200;
  assign \new_[61011]_  = ~A235 & ~A234;
  assign \new_[61012]_  = \new_[61011]_  & \new_[61008]_ ;
  assign \new_[61013]_  = \new_[61012]_  & \new_[61005]_ ;
  assign \new_[61016]_  = A265 & ~A236;
  assign \new_[61019]_  = ~A267 & A266;
  assign \new_[61020]_  = \new_[61019]_  & \new_[61016]_ ;
  assign \new_[61023]_  = ~A298 & ~A268;
  assign \new_[61026]_  = A302 & A299;
  assign \new_[61027]_  = \new_[61026]_  & \new_[61023]_ ;
  assign \new_[61028]_  = \new_[61027]_  & \new_[61020]_ ;
  assign \new_[61031]_  = ~A167 & ~A169;
  assign \new_[61034]_  = ~A199 & ~A166;
  assign \new_[61035]_  = \new_[61034]_  & \new_[61031]_ ;
  assign \new_[61038]_  = A203 & A200;
  assign \new_[61041]_  = A233 & A232;
  assign \new_[61042]_  = \new_[61041]_  & \new_[61038]_ ;
  assign \new_[61043]_  = \new_[61042]_  & \new_[61035]_ ;
  assign \new_[61046]_  = ~A235 & ~A234;
  assign \new_[61049]_  = ~A268 & ~A267;
  assign \new_[61050]_  = \new_[61049]_  & \new_[61046]_ ;
  assign \new_[61053]_  = A298 & ~A269;
  assign \new_[61056]_  = A302 & ~A299;
  assign \new_[61057]_  = \new_[61056]_  & \new_[61053]_ ;
  assign \new_[61058]_  = \new_[61057]_  & \new_[61050]_ ;
  assign \new_[61061]_  = ~A167 & ~A169;
  assign \new_[61064]_  = ~A199 & ~A166;
  assign \new_[61065]_  = \new_[61064]_  & \new_[61061]_ ;
  assign \new_[61068]_  = A203 & A200;
  assign \new_[61071]_  = A233 & A232;
  assign \new_[61072]_  = \new_[61071]_  & \new_[61068]_ ;
  assign \new_[61073]_  = \new_[61072]_  & \new_[61065]_ ;
  assign \new_[61076]_  = ~A235 & ~A234;
  assign \new_[61079]_  = ~A268 & ~A267;
  assign \new_[61080]_  = \new_[61079]_  & \new_[61076]_ ;
  assign \new_[61083]_  = ~A298 & ~A269;
  assign \new_[61086]_  = A302 & A299;
  assign \new_[61087]_  = \new_[61086]_  & \new_[61083]_ ;
  assign \new_[61088]_  = \new_[61087]_  & \new_[61080]_ ;
  assign \new_[61091]_  = ~A167 & ~A169;
  assign \new_[61094]_  = ~A199 & ~A166;
  assign \new_[61095]_  = \new_[61094]_  & \new_[61091]_ ;
  assign \new_[61098]_  = A203 & A200;
  assign \new_[61101]_  = A233 & A232;
  assign \new_[61102]_  = \new_[61101]_  & \new_[61098]_ ;
  assign \new_[61103]_  = \new_[61102]_  & \new_[61095]_ ;
  assign \new_[61106]_  = ~A235 & ~A234;
  assign \new_[61109]_  = A266 & A265;
  assign \new_[61110]_  = \new_[61109]_  & \new_[61106]_ ;
  assign \new_[61113]_  = ~A268 & ~A267;
  assign \new_[61116]_  = A300 & A299;
  assign \new_[61117]_  = \new_[61116]_  & \new_[61113]_ ;
  assign \new_[61118]_  = \new_[61117]_  & \new_[61110]_ ;
  assign \new_[61121]_  = ~A167 & ~A169;
  assign \new_[61124]_  = ~A199 & ~A166;
  assign \new_[61125]_  = \new_[61124]_  & \new_[61121]_ ;
  assign \new_[61128]_  = A203 & A200;
  assign \new_[61131]_  = A233 & A232;
  assign \new_[61132]_  = \new_[61131]_  & \new_[61128]_ ;
  assign \new_[61133]_  = \new_[61132]_  & \new_[61125]_ ;
  assign \new_[61136]_  = ~A235 & ~A234;
  assign \new_[61139]_  = A266 & A265;
  assign \new_[61140]_  = \new_[61139]_  & \new_[61136]_ ;
  assign \new_[61143]_  = ~A268 & ~A267;
  assign \new_[61146]_  = A300 & A298;
  assign \new_[61147]_  = \new_[61146]_  & \new_[61143]_ ;
  assign \new_[61148]_  = \new_[61147]_  & \new_[61140]_ ;
  assign \new_[61151]_  = ~A167 & ~A169;
  assign \new_[61154]_  = ~A199 & ~A166;
  assign \new_[61155]_  = \new_[61154]_  & \new_[61151]_ ;
  assign \new_[61158]_  = A203 & A200;
  assign \new_[61161]_  = A233 & A232;
  assign \new_[61162]_  = \new_[61161]_  & \new_[61158]_ ;
  assign \new_[61163]_  = \new_[61162]_  & \new_[61155]_ ;
  assign \new_[61166]_  = ~A235 & ~A234;
  assign \new_[61169]_  = ~A266 & ~A265;
  assign \new_[61170]_  = \new_[61169]_  & \new_[61166]_ ;
  assign \new_[61173]_  = A298 & ~A268;
  assign \new_[61176]_  = A302 & ~A299;
  assign \new_[61177]_  = \new_[61176]_  & \new_[61173]_ ;
  assign \new_[61178]_  = \new_[61177]_  & \new_[61170]_ ;
  assign \new_[61181]_  = ~A167 & ~A169;
  assign \new_[61184]_  = ~A199 & ~A166;
  assign \new_[61185]_  = \new_[61184]_  & \new_[61181]_ ;
  assign \new_[61188]_  = A203 & A200;
  assign \new_[61191]_  = A233 & A232;
  assign \new_[61192]_  = \new_[61191]_  & \new_[61188]_ ;
  assign \new_[61193]_  = \new_[61192]_  & \new_[61185]_ ;
  assign \new_[61196]_  = ~A235 & ~A234;
  assign \new_[61199]_  = ~A266 & ~A265;
  assign \new_[61200]_  = \new_[61199]_  & \new_[61196]_ ;
  assign \new_[61203]_  = ~A298 & ~A268;
  assign \new_[61206]_  = A302 & A299;
  assign \new_[61207]_  = \new_[61206]_  & \new_[61203]_ ;
  assign \new_[61208]_  = \new_[61207]_  & \new_[61200]_ ;
  assign \new_[61211]_  = ~A167 & ~A169;
  assign \new_[61214]_  = ~A199 & ~A166;
  assign \new_[61215]_  = \new_[61214]_  & \new_[61211]_ ;
  assign \new_[61218]_  = A203 & A200;
  assign \new_[61221]_  = ~A233 & ~A232;
  assign \new_[61222]_  = \new_[61221]_  & \new_[61218]_ ;
  assign \new_[61223]_  = \new_[61222]_  & \new_[61215]_ ;
  assign \new_[61226]_  = A265 & ~A235;
  assign \new_[61229]_  = ~A267 & A266;
  assign \new_[61230]_  = \new_[61229]_  & \new_[61226]_ ;
  assign \new_[61233]_  = A298 & ~A268;
  assign \new_[61236]_  = A302 & ~A299;
  assign \new_[61237]_  = \new_[61236]_  & \new_[61233]_ ;
  assign \new_[61238]_  = \new_[61237]_  & \new_[61230]_ ;
  assign \new_[61241]_  = ~A167 & ~A169;
  assign \new_[61244]_  = ~A199 & ~A166;
  assign \new_[61245]_  = \new_[61244]_  & \new_[61241]_ ;
  assign \new_[61248]_  = A203 & A200;
  assign \new_[61251]_  = ~A233 & ~A232;
  assign \new_[61252]_  = \new_[61251]_  & \new_[61248]_ ;
  assign \new_[61253]_  = \new_[61252]_  & \new_[61245]_ ;
  assign \new_[61256]_  = A265 & ~A235;
  assign \new_[61259]_  = ~A267 & A266;
  assign \new_[61260]_  = \new_[61259]_  & \new_[61256]_ ;
  assign \new_[61263]_  = ~A298 & ~A268;
  assign \new_[61266]_  = A302 & A299;
  assign \new_[61267]_  = \new_[61266]_  & \new_[61263]_ ;
  assign \new_[61268]_  = \new_[61267]_  & \new_[61260]_ ;
  assign \new_[61271]_  = ~A167 & ~A169;
  assign \new_[61274]_  = A199 & ~A166;
  assign \new_[61275]_  = \new_[61274]_  & \new_[61271]_ ;
  assign \new_[61278]_  = A203 & ~A200;
  assign \new_[61281]_  = ~A235 & ~A234;
  assign \new_[61282]_  = \new_[61281]_  & \new_[61278]_ ;
  assign \new_[61283]_  = \new_[61282]_  & \new_[61275]_ ;
  assign \new_[61286]_  = A265 & ~A236;
  assign \new_[61289]_  = ~A267 & A266;
  assign \new_[61290]_  = \new_[61289]_  & \new_[61286]_ ;
  assign \new_[61293]_  = A298 & ~A268;
  assign \new_[61296]_  = A302 & ~A299;
  assign \new_[61297]_  = \new_[61296]_  & \new_[61293]_ ;
  assign \new_[61298]_  = \new_[61297]_  & \new_[61290]_ ;
  assign \new_[61301]_  = ~A167 & ~A169;
  assign \new_[61304]_  = A199 & ~A166;
  assign \new_[61305]_  = \new_[61304]_  & \new_[61301]_ ;
  assign \new_[61308]_  = A203 & ~A200;
  assign \new_[61311]_  = ~A235 & ~A234;
  assign \new_[61312]_  = \new_[61311]_  & \new_[61308]_ ;
  assign \new_[61313]_  = \new_[61312]_  & \new_[61305]_ ;
  assign \new_[61316]_  = A265 & ~A236;
  assign \new_[61319]_  = ~A267 & A266;
  assign \new_[61320]_  = \new_[61319]_  & \new_[61316]_ ;
  assign \new_[61323]_  = ~A298 & ~A268;
  assign \new_[61326]_  = A302 & A299;
  assign \new_[61327]_  = \new_[61326]_  & \new_[61323]_ ;
  assign \new_[61328]_  = \new_[61327]_  & \new_[61320]_ ;
  assign \new_[61331]_  = ~A167 & ~A169;
  assign \new_[61334]_  = A199 & ~A166;
  assign \new_[61335]_  = \new_[61334]_  & \new_[61331]_ ;
  assign \new_[61338]_  = A203 & ~A200;
  assign \new_[61341]_  = A233 & A232;
  assign \new_[61342]_  = \new_[61341]_  & \new_[61338]_ ;
  assign \new_[61343]_  = \new_[61342]_  & \new_[61335]_ ;
  assign \new_[61346]_  = ~A235 & ~A234;
  assign \new_[61349]_  = ~A268 & ~A267;
  assign \new_[61350]_  = \new_[61349]_  & \new_[61346]_ ;
  assign \new_[61353]_  = A298 & ~A269;
  assign \new_[61356]_  = A302 & ~A299;
  assign \new_[61357]_  = \new_[61356]_  & \new_[61353]_ ;
  assign \new_[61358]_  = \new_[61357]_  & \new_[61350]_ ;
  assign \new_[61361]_  = ~A167 & ~A169;
  assign \new_[61364]_  = A199 & ~A166;
  assign \new_[61365]_  = \new_[61364]_  & \new_[61361]_ ;
  assign \new_[61368]_  = A203 & ~A200;
  assign \new_[61371]_  = A233 & A232;
  assign \new_[61372]_  = \new_[61371]_  & \new_[61368]_ ;
  assign \new_[61373]_  = \new_[61372]_  & \new_[61365]_ ;
  assign \new_[61376]_  = ~A235 & ~A234;
  assign \new_[61379]_  = ~A268 & ~A267;
  assign \new_[61380]_  = \new_[61379]_  & \new_[61376]_ ;
  assign \new_[61383]_  = ~A298 & ~A269;
  assign \new_[61386]_  = A302 & A299;
  assign \new_[61387]_  = \new_[61386]_  & \new_[61383]_ ;
  assign \new_[61388]_  = \new_[61387]_  & \new_[61380]_ ;
  assign \new_[61391]_  = ~A167 & ~A169;
  assign \new_[61394]_  = A199 & ~A166;
  assign \new_[61395]_  = \new_[61394]_  & \new_[61391]_ ;
  assign \new_[61398]_  = A203 & ~A200;
  assign \new_[61401]_  = A233 & A232;
  assign \new_[61402]_  = \new_[61401]_  & \new_[61398]_ ;
  assign \new_[61403]_  = \new_[61402]_  & \new_[61395]_ ;
  assign \new_[61406]_  = ~A235 & ~A234;
  assign \new_[61409]_  = A266 & A265;
  assign \new_[61410]_  = \new_[61409]_  & \new_[61406]_ ;
  assign \new_[61413]_  = ~A268 & ~A267;
  assign \new_[61416]_  = A300 & A299;
  assign \new_[61417]_  = \new_[61416]_  & \new_[61413]_ ;
  assign \new_[61418]_  = \new_[61417]_  & \new_[61410]_ ;
  assign \new_[61421]_  = ~A167 & ~A169;
  assign \new_[61424]_  = A199 & ~A166;
  assign \new_[61425]_  = \new_[61424]_  & \new_[61421]_ ;
  assign \new_[61428]_  = A203 & ~A200;
  assign \new_[61431]_  = A233 & A232;
  assign \new_[61432]_  = \new_[61431]_  & \new_[61428]_ ;
  assign \new_[61433]_  = \new_[61432]_  & \new_[61425]_ ;
  assign \new_[61436]_  = ~A235 & ~A234;
  assign \new_[61439]_  = A266 & A265;
  assign \new_[61440]_  = \new_[61439]_  & \new_[61436]_ ;
  assign \new_[61443]_  = ~A268 & ~A267;
  assign \new_[61446]_  = A300 & A298;
  assign \new_[61447]_  = \new_[61446]_  & \new_[61443]_ ;
  assign \new_[61448]_  = \new_[61447]_  & \new_[61440]_ ;
  assign \new_[61451]_  = ~A167 & ~A169;
  assign \new_[61454]_  = A199 & ~A166;
  assign \new_[61455]_  = \new_[61454]_  & \new_[61451]_ ;
  assign \new_[61458]_  = A203 & ~A200;
  assign \new_[61461]_  = A233 & A232;
  assign \new_[61462]_  = \new_[61461]_  & \new_[61458]_ ;
  assign \new_[61463]_  = \new_[61462]_  & \new_[61455]_ ;
  assign \new_[61466]_  = ~A235 & ~A234;
  assign \new_[61469]_  = ~A266 & ~A265;
  assign \new_[61470]_  = \new_[61469]_  & \new_[61466]_ ;
  assign \new_[61473]_  = A298 & ~A268;
  assign \new_[61476]_  = A302 & ~A299;
  assign \new_[61477]_  = \new_[61476]_  & \new_[61473]_ ;
  assign \new_[61478]_  = \new_[61477]_  & \new_[61470]_ ;
  assign \new_[61481]_  = ~A167 & ~A169;
  assign \new_[61484]_  = A199 & ~A166;
  assign \new_[61485]_  = \new_[61484]_  & \new_[61481]_ ;
  assign \new_[61488]_  = A203 & ~A200;
  assign \new_[61491]_  = A233 & A232;
  assign \new_[61492]_  = \new_[61491]_  & \new_[61488]_ ;
  assign \new_[61493]_  = \new_[61492]_  & \new_[61485]_ ;
  assign \new_[61496]_  = ~A235 & ~A234;
  assign \new_[61499]_  = ~A266 & ~A265;
  assign \new_[61500]_  = \new_[61499]_  & \new_[61496]_ ;
  assign \new_[61503]_  = ~A298 & ~A268;
  assign \new_[61506]_  = A302 & A299;
  assign \new_[61507]_  = \new_[61506]_  & \new_[61503]_ ;
  assign \new_[61508]_  = \new_[61507]_  & \new_[61500]_ ;
  assign \new_[61511]_  = ~A167 & ~A169;
  assign \new_[61514]_  = A199 & ~A166;
  assign \new_[61515]_  = \new_[61514]_  & \new_[61511]_ ;
  assign \new_[61518]_  = A203 & ~A200;
  assign \new_[61521]_  = ~A233 & ~A232;
  assign \new_[61522]_  = \new_[61521]_  & \new_[61518]_ ;
  assign \new_[61523]_  = \new_[61522]_  & \new_[61515]_ ;
  assign \new_[61526]_  = A265 & ~A235;
  assign \new_[61529]_  = ~A267 & A266;
  assign \new_[61530]_  = \new_[61529]_  & \new_[61526]_ ;
  assign \new_[61533]_  = A298 & ~A268;
  assign \new_[61536]_  = A302 & ~A299;
  assign \new_[61537]_  = \new_[61536]_  & \new_[61533]_ ;
  assign \new_[61538]_  = \new_[61537]_  & \new_[61530]_ ;
  assign \new_[61541]_  = ~A167 & ~A169;
  assign \new_[61544]_  = A199 & ~A166;
  assign \new_[61545]_  = \new_[61544]_  & \new_[61541]_ ;
  assign \new_[61548]_  = A203 & ~A200;
  assign \new_[61551]_  = ~A233 & ~A232;
  assign \new_[61552]_  = \new_[61551]_  & \new_[61548]_ ;
  assign \new_[61553]_  = \new_[61552]_  & \new_[61545]_ ;
  assign \new_[61556]_  = A265 & ~A235;
  assign \new_[61559]_  = ~A267 & A266;
  assign \new_[61560]_  = \new_[61559]_  & \new_[61556]_ ;
  assign \new_[61563]_  = ~A298 & ~A268;
  assign \new_[61566]_  = A302 & A299;
  assign \new_[61567]_  = \new_[61566]_  & \new_[61563]_ ;
  assign \new_[61568]_  = \new_[61567]_  & \new_[61560]_ ;
  assign \new_[61571]_  = ~A168 & ~A169;
  assign \new_[61574]_  = A166 & A167;
  assign \new_[61575]_  = \new_[61574]_  & \new_[61571]_ ;
  assign \new_[61578]_  = A232 & A202;
  assign \new_[61581]_  = ~A234 & A233;
  assign \new_[61582]_  = \new_[61581]_  & \new_[61578]_ ;
  assign \new_[61583]_  = \new_[61582]_  & \new_[61575]_ ;
  assign \new_[61586]_  = A265 & ~A235;
  assign \new_[61589]_  = ~A267 & A266;
  assign \new_[61590]_  = \new_[61589]_  & \new_[61586]_ ;
  assign \new_[61593]_  = A298 & ~A268;
  assign \new_[61596]_  = A302 & ~A299;
  assign \new_[61597]_  = \new_[61596]_  & \new_[61593]_ ;
  assign \new_[61598]_  = \new_[61597]_  & \new_[61590]_ ;
  assign \new_[61601]_  = ~A168 & ~A169;
  assign \new_[61604]_  = A166 & A167;
  assign \new_[61605]_  = \new_[61604]_  & \new_[61601]_ ;
  assign \new_[61608]_  = A232 & A202;
  assign \new_[61611]_  = ~A234 & A233;
  assign \new_[61612]_  = \new_[61611]_  & \new_[61608]_ ;
  assign \new_[61613]_  = \new_[61612]_  & \new_[61605]_ ;
  assign \new_[61616]_  = A265 & ~A235;
  assign \new_[61619]_  = ~A267 & A266;
  assign \new_[61620]_  = \new_[61619]_  & \new_[61616]_ ;
  assign \new_[61623]_  = ~A298 & ~A268;
  assign \new_[61626]_  = A302 & A299;
  assign \new_[61627]_  = \new_[61626]_  & \new_[61623]_ ;
  assign \new_[61628]_  = \new_[61627]_  & \new_[61620]_ ;
  assign \new_[61631]_  = ~A168 & ~A169;
  assign \new_[61634]_  = A166 & A167;
  assign \new_[61635]_  = \new_[61634]_  & \new_[61631]_ ;
  assign \new_[61638]_  = A201 & A199;
  assign \new_[61641]_  = ~A235 & ~A234;
  assign \new_[61642]_  = \new_[61641]_  & \new_[61638]_ ;
  assign \new_[61643]_  = \new_[61642]_  & \new_[61635]_ ;
  assign \new_[61646]_  = A265 & ~A236;
  assign \new_[61649]_  = ~A267 & A266;
  assign \new_[61650]_  = \new_[61649]_  & \new_[61646]_ ;
  assign \new_[61653]_  = A298 & ~A268;
  assign \new_[61656]_  = A302 & ~A299;
  assign \new_[61657]_  = \new_[61656]_  & \new_[61653]_ ;
  assign \new_[61658]_  = \new_[61657]_  & \new_[61650]_ ;
  assign \new_[61661]_  = ~A168 & ~A169;
  assign \new_[61664]_  = A166 & A167;
  assign \new_[61665]_  = \new_[61664]_  & \new_[61661]_ ;
  assign \new_[61668]_  = A201 & A199;
  assign \new_[61671]_  = ~A235 & ~A234;
  assign \new_[61672]_  = \new_[61671]_  & \new_[61668]_ ;
  assign \new_[61673]_  = \new_[61672]_  & \new_[61665]_ ;
  assign \new_[61676]_  = A265 & ~A236;
  assign \new_[61679]_  = ~A267 & A266;
  assign \new_[61680]_  = \new_[61679]_  & \new_[61676]_ ;
  assign \new_[61683]_  = ~A298 & ~A268;
  assign \new_[61686]_  = A302 & A299;
  assign \new_[61687]_  = \new_[61686]_  & \new_[61683]_ ;
  assign \new_[61688]_  = \new_[61687]_  & \new_[61680]_ ;
  assign \new_[61691]_  = ~A168 & ~A169;
  assign \new_[61694]_  = A166 & A167;
  assign \new_[61695]_  = \new_[61694]_  & \new_[61691]_ ;
  assign \new_[61698]_  = A201 & A199;
  assign \new_[61701]_  = A233 & A232;
  assign \new_[61702]_  = \new_[61701]_  & \new_[61698]_ ;
  assign \new_[61703]_  = \new_[61702]_  & \new_[61695]_ ;
  assign \new_[61706]_  = ~A235 & ~A234;
  assign \new_[61709]_  = ~A268 & ~A267;
  assign \new_[61710]_  = \new_[61709]_  & \new_[61706]_ ;
  assign \new_[61713]_  = A298 & ~A269;
  assign \new_[61716]_  = A302 & ~A299;
  assign \new_[61717]_  = \new_[61716]_  & \new_[61713]_ ;
  assign \new_[61718]_  = \new_[61717]_  & \new_[61710]_ ;
  assign \new_[61721]_  = ~A168 & ~A169;
  assign \new_[61724]_  = A166 & A167;
  assign \new_[61725]_  = \new_[61724]_  & \new_[61721]_ ;
  assign \new_[61728]_  = A201 & A199;
  assign \new_[61731]_  = A233 & A232;
  assign \new_[61732]_  = \new_[61731]_  & \new_[61728]_ ;
  assign \new_[61733]_  = \new_[61732]_  & \new_[61725]_ ;
  assign \new_[61736]_  = ~A235 & ~A234;
  assign \new_[61739]_  = ~A268 & ~A267;
  assign \new_[61740]_  = \new_[61739]_  & \new_[61736]_ ;
  assign \new_[61743]_  = ~A298 & ~A269;
  assign \new_[61746]_  = A302 & A299;
  assign \new_[61747]_  = \new_[61746]_  & \new_[61743]_ ;
  assign \new_[61748]_  = \new_[61747]_  & \new_[61740]_ ;
  assign \new_[61751]_  = ~A168 & ~A169;
  assign \new_[61754]_  = A166 & A167;
  assign \new_[61755]_  = \new_[61754]_  & \new_[61751]_ ;
  assign \new_[61758]_  = A201 & A199;
  assign \new_[61761]_  = A233 & A232;
  assign \new_[61762]_  = \new_[61761]_  & \new_[61758]_ ;
  assign \new_[61763]_  = \new_[61762]_  & \new_[61755]_ ;
  assign \new_[61766]_  = ~A235 & ~A234;
  assign \new_[61769]_  = A266 & A265;
  assign \new_[61770]_  = \new_[61769]_  & \new_[61766]_ ;
  assign \new_[61773]_  = ~A268 & ~A267;
  assign \new_[61776]_  = A300 & A299;
  assign \new_[61777]_  = \new_[61776]_  & \new_[61773]_ ;
  assign \new_[61778]_  = \new_[61777]_  & \new_[61770]_ ;
  assign \new_[61781]_  = ~A168 & ~A169;
  assign \new_[61784]_  = A166 & A167;
  assign \new_[61785]_  = \new_[61784]_  & \new_[61781]_ ;
  assign \new_[61788]_  = A201 & A199;
  assign \new_[61791]_  = A233 & A232;
  assign \new_[61792]_  = \new_[61791]_  & \new_[61788]_ ;
  assign \new_[61793]_  = \new_[61792]_  & \new_[61785]_ ;
  assign \new_[61796]_  = ~A235 & ~A234;
  assign \new_[61799]_  = A266 & A265;
  assign \new_[61800]_  = \new_[61799]_  & \new_[61796]_ ;
  assign \new_[61803]_  = ~A268 & ~A267;
  assign \new_[61806]_  = A300 & A298;
  assign \new_[61807]_  = \new_[61806]_  & \new_[61803]_ ;
  assign \new_[61808]_  = \new_[61807]_  & \new_[61800]_ ;
  assign \new_[61811]_  = ~A168 & ~A169;
  assign \new_[61814]_  = A166 & A167;
  assign \new_[61815]_  = \new_[61814]_  & \new_[61811]_ ;
  assign \new_[61818]_  = A201 & A199;
  assign \new_[61821]_  = A233 & A232;
  assign \new_[61822]_  = \new_[61821]_  & \new_[61818]_ ;
  assign \new_[61823]_  = \new_[61822]_  & \new_[61815]_ ;
  assign \new_[61826]_  = ~A235 & ~A234;
  assign \new_[61829]_  = ~A266 & ~A265;
  assign \new_[61830]_  = \new_[61829]_  & \new_[61826]_ ;
  assign \new_[61833]_  = A298 & ~A268;
  assign \new_[61836]_  = A302 & ~A299;
  assign \new_[61837]_  = \new_[61836]_  & \new_[61833]_ ;
  assign \new_[61838]_  = \new_[61837]_  & \new_[61830]_ ;
  assign \new_[61841]_  = ~A168 & ~A169;
  assign \new_[61844]_  = A166 & A167;
  assign \new_[61845]_  = \new_[61844]_  & \new_[61841]_ ;
  assign \new_[61848]_  = A201 & A199;
  assign \new_[61851]_  = A233 & A232;
  assign \new_[61852]_  = \new_[61851]_  & \new_[61848]_ ;
  assign \new_[61853]_  = \new_[61852]_  & \new_[61845]_ ;
  assign \new_[61856]_  = ~A235 & ~A234;
  assign \new_[61859]_  = ~A266 & ~A265;
  assign \new_[61860]_  = \new_[61859]_  & \new_[61856]_ ;
  assign \new_[61863]_  = ~A298 & ~A268;
  assign \new_[61866]_  = A302 & A299;
  assign \new_[61867]_  = \new_[61866]_  & \new_[61863]_ ;
  assign \new_[61868]_  = \new_[61867]_  & \new_[61860]_ ;
  assign \new_[61871]_  = ~A168 & ~A169;
  assign \new_[61874]_  = A166 & A167;
  assign \new_[61875]_  = \new_[61874]_  & \new_[61871]_ ;
  assign \new_[61878]_  = A201 & A199;
  assign \new_[61881]_  = ~A233 & ~A232;
  assign \new_[61882]_  = \new_[61881]_  & \new_[61878]_ ;
  assign \new_[61883]_  = \new_[61882]_  & \new_[61875]_ ;
  assign \new_[61886]_  = A265 & ~A235;
  assign \new_[61889]_  = ~A267 & A266;
  assign \new_[61890]_  = \new_[61889]_  & \new_[61886]_ ;
  assign \new_[61893]_  = A298 & ~A268;
  assign \new_[61896]_  = A302 & ~A299;
  assign \new_[61897]_  = \new_[61896]_  & \new_[61893]_ ;
  assign \new_[61898]_  = \new_[61897]_  & \new_[61890]_ ;
  assign \new_[61901]_  = ~A168 & ~A169;
  assign \new_[61904]_  = A166 & A167;
  assign \new_[61905]_  = \new_[61904]_  & \new_[61901]_ ;
  assign \new_[61908]_  = A201 & A199;
  assign \new_[61911]_  = ~A233 & ~A232;
  assign \new_[61912]_  = \new_[61911]_  & \new_[61908]_ ;
  assign \new_[61913]_  = \new_[61912]_  & \new_[61905]_ ;
  assign \new_[61916]_  = A265 & ~A235;
  assign \new_[61919]_  = ~A267 & A266;
  assign \new_[61920]_  = \new_[61919]_  & \new_[61916]_ ;
  assign \new_[61923]_  = ~A298 & ~A268;
  assign \new_[61926]_  = A302 & A299;
  assign \new_[61927]_  = \new_[61926]_  & \new_[61923]_ ;
  assign \new_[61928]_  = \new_[61927]_  & \new_[61920]_ ;
  assign \new_[61931]_  = ~A168 & ~A169;
  assign \new_[61934]_  = A166 & A167;
  assign \new_[61935]_  = \new_[61934]_  & \new_[61931]_ ;
  assign \new_[61938]_  = A201 & A200;
  assign \new_[61941]_  = ~A235 & ~A234;
  assign \new_[61942]_  = \new_[61941]_  & \new_[61938]_ ;
  assign \new_[61943]_  = \new_[61942]_  & \new_[61935]_ ;
  assign \new_[61946]_  = A265 & ~A236;
  assign \new_[61949]_  = ~A267 & A266;
  assign \new_[61950]_  = \new_[61949]_  & \new_[61946]_ ;
  assign \new_[61953]_  = A298 & ~A268;
  assign \new_[61956]_  = A302 & ~A299;
  assign \new_[61957]_  = \new_[61956]_  & \new_[61953]_ ;
  assign \new_[61958]_  = \new_[61957]_  & \new_[61950]_ ;
  assign \new_[61961]_  = ~A168 & ~A169;
  assign \new_[61964]_  = A166 & A167;
  assign \new_[61965]_  = \new_[61964]_  & \new_[61961]_ ;
  assign \new_[61968]_  = A201 & A200;
  assign \new_[61971]_  = ~A235 & ~A234;
  assign \new_[61972]_  = \new_[61971]_  & \new_[61968]_ ;
  assign \new_[61973]_  = \new_[61972]_  & \new_[61965]_ ;
  assign \new_[61976]_  = A265 & ~A236;
  assign \new_[61979]_  = ~A267 & A266;
  assign \new_[61980]_  = \new_[61979]_  & \new_[61976]_ ;
  assign \new_[61983]_  = ~A298 & ~A268;
  assign \new_[61986]_  = A302 & A299;
  assign \new_[61987]_  = \new_[61986]_  & \new_[61983]_ ;
  assign \new_[61988]_  = \new_[61987]_  & \new_[61980]_ ;
  assign \new_[61991]_  = ~A168 & ~A169;
  assign \new_[61994]_  = A166 & A167;
  assign \new_[61995]_  = \new_[61994]_  & \new_[61991]_ ;
  assign \new_[61998]_  = A201 & A200;
  assign \new_[62001]_  = A233 & A232;
  assign \new_[62002]_  = \new_[62001]_  & \new_[61998]_ ;
  assign \new_[62003]_  = \new_[62002]_  & \new_[61995]_ ;
  assign \new_[62006]_  = ~A235 & ~A234;
  assign \new_[62009]_  = ~A268 & ~A267;
  assign \new_[62010]_  = \new_[62009]_  & \new_[62006]_ ;
  assign \new_[62013]_  = A298 & ~A269;
  assign \new_[62016]_  = A302 & ~A299;
  assign \new_[62017]_  = \new_[62016]_  & \new_[62013]_ ;
  assign \new_[62018]_  = \new_[62017]_  & \new_[62010]_ ;
  assign \new_[62021]_  = ~A168 & ~A169;
  assign \new_[62024]_  = A166 & A167;
  assign \new_[62025]_  = \new_[62024]_  & \new_[62021]_ ;
  assign \new_[62028]_  = A201 & A200;
  assign \new_[62031]_  = A233 & A232;
  assign \new_[62032]_  = \new_[62031]_  & \new_[62028]_ ;
  assign \new_[62033]_  = \new_[62032]_  & \new_[62025]_ ;
  assign \new_[62036]_  = ~A235 & ~A234;
  assign \new_[62039]_  = ~A268 & ~A267;
  assign \new_[62040]_  = \new_[62039]_  & \new_[62036]_ ;
  assign \new_[62043]_  = ~A298 & ~A269;
  assign \new_[62046]_  = A302 & A299;
  assign \new_[62047]_  = \new_[62046]_  & \new_[62043]_ ;
  assign \new_[62048]_  = \new_[62047]_  & \new_[62040]_ ;
  assign \new_[62051]_  = ~A168 & ~A169;
  assign \new_[62054]_  = A166 & A167;
  assign \new_[62055]_  = \new_[62054]_  & \new_[62051]_ ;
  assign \new_[62058]_  = A201 & A200;
  assign \new_[62061]_  = A233 & A232;
  assign \new_[62062]_  = \new_[62061]_  & \new_[62058]_ ;
  assign \new_[62063]_  = \new_[62062]_  & \new_[62055]_ ;
  assign \new_[62066]_  = ~A235 & ~A234;
  assign \new_[62069]_  = A266 & A265;
  assign \new_[62070]_  = \new_[62069]_  & \new_[62066]_ ;
  assign \new_[62073]_  = ~A268 & ~A267;
  assign \new_[62076]_  = A300 & A299;
  assign \new_[62077]_  = \new_[62076]_  & \new_[62073]_ ;
  assign \new_[62078]_  = \new_[62077]_  & \new_[62070]_ ;
  assign \new_[62081]_  = ~A168 & ~A169;
  assign \new_[62084]_  = A166 & A167;
  assign \new_[62085]_  = \new_[62084]_  & \new_[62081]_ ;
  assign \new_[62088]_  = A201 & A200;
  assign \new_[62091]_  = A233 & A232;
  assign \new_[62092]_  = \new_[62091]_  & \new_[62088]_ ;
  assign \new_[62093]_  = \new_[62092]_  & \new_[62085]_ ;
  assign \new_[62096]_  = ~A235 & ~A234;
  assign \new_[62099]_  = A266 & A265;
  assign \new_[62100]_  = \new_[62099]_  & \new_[62096]_ ;
  assign \new_[62103]_  = ~A268 & ~A267;
  assign \new_[62106]_  = A300 & A298;
  assign \new_[62107]_  = \new_[62106]_  & \new_[62103]_ ;
  assign \new_[62108]_  = \new_[62107]_  & \new_[62100]_ ;
  assign \new_[62111]_  = ~A168 & ~A169;
  assign \new_[62114]_  = A166 & A167;
  assign \new_[62115]_  = \new_[62114]_  & \new_[62111]_ ;
  assign \new_[62118]_  = A201 & A200;
  assign \new_[62121]_  = A233 & A232;
  assign \new_[62122]_  = \new_[62121]_  & \new_[62118]_ ;
  assign \new_[62123]_  = \new_[62122]_  & \new_[62115]_ ;
  assign \new_[62126]_  = ~A235 & ~A234;
  assign \new_[62129]_  = ~A266 & ~A265;
  assign \new_[62130]_  = \new_[62129]_  & \new_[62126]_ ;
  assign \new_[62133]_  = A298 & ~A268;
  assign \new_[62136]_  = A302 & ~A299;
  assign \new_[62137]_  = \new_[62136]_  & \new_[62133]_ ;
  assign \new_[62138]_  = \new_[62137]_  & \new_[62130]_ ;
  assign \new_[62141]_  = ~A168 & ~A169;
  assign \new_[62144]_  = A166 & A167;
  assign \new_[62145]_  = \new_[62144]_  & \new_[62141]_ ;
  assign \new_[62148]_  = A201 & A200;
  assign \new_[62151]_  = A233 & A232;
  assign \new_[62152]_  = \new_[62151]_  & \new_[62148]_ ;
  assign \new_[62153]_  = \new_[62152]_  & \new_[62145]_ ;
  assign \new_[62156]_  = ~A235 & ~A234;
  assign \new_[62159]_  = ~A266 & ~A265;
  assign \new_[62160]_  = \new_[62159]_  & \new_[62156]_ ;
  assign \new_[62163]_  = ~A298 & ~A268;
  assign \new_[62166]_  = A302 & A299;
  assign \new_[62167]_  = \new_[62166]_  & \new_[62163]_ ;
  assign \new_[62168]_  = \new_[62167]_  & \new_[62160]_ ;
  assign \new_[62171]_  = ~A168 & ~A169;
  assign \new_[62174]_  = A166 & A167;
  assign \new_[62175]_  = \new_[62174]_  & \new_[62171]_ ;
  assign \new_[62178]_  = A201 & A200;
  assign \new_[62181]_  = ~A233 & ~A232;
  assign \new_[62182]_  = \new_[62181]_  & \new_[62178]_ ;
  assign \new_[62183]_  = \new_[62182]_  & \new_[62175]_ ;
  assign \new_[62186]_  = A265 & ~A235;
  assign \new_[62189]_  = ~A267 & A266;
  assign \new_[62190]_  = \new_[62189]_  & \new_[62186]_ ;
  assign \new_[62193]_  = A298 & ~A268;
  assign \new_[62196]_  = A302 & ~A299;
  assign \new_[62197]_  = \new_[62196]_  & \new_[62193]_ ;
  assign \new_[62198]_  = \new_[62197]_  & \new_[62190]_ ;
  assign \new_[62201]_  = ~A168 & ~A169;
  assign \new_[62204]_  = A166 & A167;
  assign \new_[62205]_  = \new_[62204]_  & \new_[62201]_ ;
  assign \new_[62208]_  = A201 & A200;
  assign \new_[62211]_  = ~A233 & ~A232;
  assign \new_[62212]_  = \new_[62211]_  & \new_[62208]_ ;
  assign \new_[62213]_  = \new_[62212]_  & \new_[62205]_ ;
  assign \new_[62216]_  = A265 & ~A235;
  assign \new_[62219]_  = ~A267 & A266;
  assign \new_[62220]_  = \new_[62219]_  & \new_[62216]_ ;
  assign \new_[62223]_  = ~A298 & ~A268;
  assign \new_[62226]_  = A302 & A299;
  assign \new_[62227]_  = \new_[62226]_  & \new_[62223]_ ;
  assign \new_[62228]_  = \new_[62227]_  & \new_[62220]_ ;
  assign \new_[62231]_  = ~A168 & ~A169;
  assign \new_[62234]_  = A166 & A167;
  assign \new_[62235]_  = \new_[62234]_  & \new_[62231]_ ;
  assign \new_[62238]_  = A200 & ~A199;
  assign \new_[62241]_  = ~A234 & A203;
  assign \new_[62242]_  = \new_[62241]_  & \new_[62238]_ ;
  assign \new_[62243]_  = \new_[62242]_  & \new_[62235]_ ;
  assign \new_[62246]_  = ~A236 & ~A235;
  assign \new_[62249]_  = ~A268 & ~A267;
  assign \new_[62250]_  = \new_[62249]_  & \new_[62246]_ ;
  assign \new_[62253]_  = A298 & ~A269;
  assign \new_[62256]_  = A302 & ~A299;
  assign \new_[62257]_  = \new_[62256]_  & \new_[62253]_ ;
  assign \new_[62258]_  = \new_[62257]_  & \new_[62250]_ ;
  assign \new_[62261]_  = ~A168 & ~A169;
  assign \new_[62264]_  = A166 & A167;
  assign \new_[62265]_  = \new_[62264]_  & \new_[62261]_ ;
  assign \new_[62268]_  = A200 & ~A199;
  assign \new_[62271]_  = ~A234 & A203;
  assign \new_[62272]_  = \new_[62271]_  & \new_[62268]_ ;
  assign \new_[62273]_  = \new_[62272]_  & \new_[62265]_ ;
  assign \new_[62276]_  = ~A236 & ~A235;
  assign \new_[62279]_  = ~A268 & ~A267;
  assign \new_[62280]_  = \new_[62279]_  & \new_[62276]_ ;
  assign \new_[62283]_  = ~A298 & ~A269;
  assign \new_[62286]_  = A302 & A299;
  assign \new_[62287]_  = \new_[62286]_  & \new_[62283]_ ;
  assign \new_[62288]_  = \new_[62287]_  & \new_[62280]_ ;
  assign \new_[62291]_  = ~A168 & ~A169;
  assign \new_[62294]_  = A166 & A167;
  assign \new_[62295]_  = \new_[62294]_  & \new_[62291]_ ;
  assign \new_[62298]_  = A200 & ~A199;
  assign \new_[62301]_  = ~A234 & A203;
  assign \new_[62302]_  = \new_[62301]_  & \new_[62298]_ ;
  assign \new_[62303]_  = \new_[62302]_  & \new_[62295]_ ;
  assign \new_[62306]_  = ~A236 & ~A235;
  assign \new_[62309]_  = A266 & A265;
  assign \new_[62310]_  = \new_[62309]_  & \new_[62306]_ ;
  assign \new_[62313]_  = ~A268 & ~A267;
  assign \new_[62316]_  = A300 & A299;
  assign \new_[62317]_  = \new_[62316]_  & \new_[62313]_ ;
  assign \new_[62318]_  = \new_[62317]_  & \new_[62310]_ ;
  assign \new_[62321]_  = ~A168 & ~A169;
  assign \new_[62324]_  = A166 & A167;
  assign \new_[62325]_  = \new_[62324]_  & \new_[62321]_ ;
  assign \new_[62328]_  = A200 & ~A199;
  assign \new_[62331]_  = ~A234 & A203;
  assign \new_[62332]_  = \new_[62331]_  & \new_[62328]_ ;
  assign \new_[62333]_  = \new_[62332]_  & \new_[62325]_ ;
  assign \new_[62336]_  = ~A236 & ~A235;
  assign \new_[62339]_  = A266 & A265;
  assign \new_[62340]_  = \new_[62339]_  & \new_[62336]_ ;
  assign \new_[62343]_  = ~A268 & ~A267;
  assign \new_[62346]_  = A300 & A298;
  assign \new_[62347]_  = \new_[62346]_  & \new_[62343]_ ;
  assign \new_[62348]_  = \new_[62347]_  & \new_[62340]_ ;
  assign \new_[62351]_  = ~A168 & ~A169;
  assign \new_[62354]_  = A166 & A167;
  assign \new_[62355]_  = \new_[62354]_  & \new_[62351]_ ;
  assign \new_[62358]_  = A200 & ~A199;
  assign \new_[62361]_  = ~A234 & A203;
  assign \new_[62362]_  = \new_[62361]_  & \new_[62358]_ ;
  assign \new_[62363]_  = \new_[62362]_  & \new_[62355]_ ;
  assign \new_[62366]_  = ~A236 & ~A235;
  assign \new_[62369]_  = ~A266 & ~A265;
  assign \new_[62370]_  = \new_[62369]_  & \new_[62366]_ ;
  assign \new_[62373]_  = A298 & ~A268;
  assign \new_[62376]_  = A302 & ~A299;
  assign \new_[62377]_  = \new_[62376]_  & \new_[62373]_ ;
  assign \new_[62378]_  = \new_[62377]_  & \new_[62370]_ ;
  assign \new_[62381]_  = ~A168 & ~A169;
  assign \new_[62384]_  = A166 & A167;
  assign \new_[62385]_  = \new_[62384]_  & \new_[62381]_ ;
  assign \new_[62388]_  = A200 & ~A199;
  assign \new_[62391]_  = ~A234 & A203;
  assign \new_[62392]_  = \new_[62391]_  & \new_[62388]_ ;
  assign \new_[62393]_  = \new_[62392]_  & \new_[62385]_ ;
  assign \new_[62396]_  = ~A236 & ~A235;
  assign \new_[62399]_  = ~A266 & ~A265;
  assign \new_[62400]_  = \new_[62399]_  & \new_[62396]_ ;
  assign \new_[62403]_  = ~A298 & ~A268;
  assign \new_[62406]_  = A302 & A299;
  assign \new_[62407]_  = \new_[62406]_  & \new_[62403]_ ;
  assign \new_[62408]_  = \new_[62407]_  & \new_[62400]_ ;
  assign \new_[62411]_  = ~A168 & ~A169;
  assign \new_[62414]_  = A166 & A167;
  assign \new_[62415]_  = \new_[62414]_  & \new_[62411]_ ;
  assign \new_[62418]_  = A200 & ~A199;
  assign \new_[62421]_  = A232 & A203;
  assign \new_[62422]_  = \new_[62421]_  & \new_[62418]_ ;
  assign \new_[62423]_  = \new_[62422]_  & \new_[62415]_ ;
  assign \new_[62426]_  = ~A234 & A233;
  assign \new_[62429]_  = ~A267 & ~A235;
  assign \new_[62430]_  = \new_[62429]_  & \new_[62426]_ ;
  assign \new_[62433]_  = ~A269 & ~A268;
  assign \new_[62436]_  = A300 & A299;
  assign \new_[62437]_  = \new_[62436]_  & \new_[62433]_ ;
  assign \new_[62438]_  = \new_[62437]_  & \new_[62430]_ ;
  assign \new_[62441]_  = ~A168 & ~A169;
  assign \new_[62444]_  = A166 & A167;
  assign \new_[62445]_  = \new_[62444]_  & \new_[62441]_ ;
  assign \new_[62448]_  = A200 & ~A199;
  assign \new_[62451]_  = A232 & A203;
  assign \new_[62452]_  = \new_[62451]_  & \new_[62448]_ ;
  assign \new_[62453]_  = \new_[62452]_  & \new_[62445]_ ;
  assign \new_[62456]_  = ~A234 & A233;
  assign \new_[62459]_  = ~A267 & ~A235;
  assign \new_[62460]_  = \new_[62459]_  & \new_[62456]_ ;
  assign \new_[62463]_  = ~A269 & ~A268;
  assign \new_[62466]_  = A300 & A298;
  assign \new_[62467]_  = \new_[62466]_  & \new_[62463]_ ;
  assign \new_[62468]_  = \new_[62467]_  & \new_[62460]_ ;
  assign \new_[62471]_  = ~A168 & ~A169;
  assign \new_[62474]_  = A166 & A167;
  assign \new_[62475]_  = \new_[62474]_  & \new_[62471]_ ;
  assign \new_[62478]_  = A200 & ~A199;
  assign \new_[62481]_  = A232 & A203;
  assign \new_[62482]_  = \new_[62481]_  & \new_[62478]_ ;
  assign \new_[62483]_  = \new_[62482]_  & \new_[62475]_ ;
  assign \new_[62486]_  = ~A234 & A233;
  assign \new_[62489]_  = A265 & ~A235;
  assign \new_[62490]_  = \new_[62489]_  & \new_[62486]_ ;
  assign \new_[62493]_  = ~A267 & A266;
  assign \new_[62496]_  = A301 & ~A268;
  assign \new_[62497]_  = \new_[62496]_  & \new_[62493]_ ;
  assign \new_[62498]_  = \new_[62497]_  & \new_[62490]_ ;
  assign \new_[62501]_  = ~A168 & ~A169;
  assign \new_[62504]_  = A166 & A167;
  assign \new_[62505]_  = \new_[62504]_  & \new_[62501]_ ;
  assign \new_[62508]_  = A200 & ~A199;
  assign \new_[62511]_  = A232 & A203;
  assign \new_[62512]_  = \new_[62511]_  & \new_[62508]_ ;
  assign \new_[62513]_  = \new_[62512]_  & \new_[62505]_ ;
  assign \new_[62516]_  = ~A234 & A233;
  assign \new_[62519]_  = ~A265 & ~A235;
  assign \new_[62520]_  = \new_[62519]_  & \new_[62516]_ ;
  assign \new_[62523]_  = ~A268 & ~A266;
  assign \new_[62526]_  = A300 & A299;
  assign \new_[62527]_  = \new_[62526]_  & \new_[62523]_ ;
  assign \new_[62528]_  = \new_[62527]_  & \new_[62520]_ ;
  assign \new_[62531]_  = ~A168 & ~A169;
  assign \new_[62534]_  = A166 & A167;
  assign \new_[62535]_  = \new_[62534]_  & \new_[62531]_ ;
  assign \new_[62538]_  = A200 & ~A199;
  assign \new_[62541]_  = A232 & A203;
  assign \new_[62542]_  = \new_[62541]_  & \new_[62538]_ ;
  assign \new_[62543]_  = \new_[62542]_  & \new_[62535]_ ;
  assign \new_[62546]_  = ~A234 & A233;
  assign \new_[62549]_  = ~A265 & ~A235;
  assign \new_[62550]_  = \new_[62549]_  & \new_[62546]_ ;
  assign \new_[62553]_  = ~A268 & ~A266;
  assign \new_[62556]_  = A300 & A298;
  assign \new_[62557]_  = \new_[62556]_  & \new_[62553]_ ;
  assign \new_[62558]_  = \new_[62557]_  & \new_[62550]_ ;
  assign \new_[62561]_  = ~A168 & ~A169;
  assign \new_[62564]_  = A166 & A167;
  assign \new_[62565]_  = \new_[62564]_  & \new_[62561]_ ;
  assign \new_[62568]_  = A200 & ~A199;
  assign \new_[62571]_  = ~A232 & A203;
  assign \new_[62572]_  = \new_[62571]_  & \new_[62568]_ ;
  assign \new_[62573]_  = \new_[62572]_  & \new_[62565]_ ;
  assign \new_[62576]_  = ~A235 & ~A233;
  assign \new_[62579]_  = ~A268 & ~A267;
  assign \new_[62580]_  = \new_[62579]_  & \new_[62576]_ ;
  assign \new_[62583]_  = A298 & ~A269;
  assign \new_[62586]_  = A302 & ~A299;
  assign \new_[62587]_  = \new_[62586]_  & \new_[62583]_ ;
  assign \new_[62588]_  = \new_[62587]_  & \new_[62580]_ ;
  assign \new_[62591]_  = ~A168 & ~A169;
  assign \new_[62594]_  = A166 & A167;
  assign \new_[62595]_  = \new_[62594]_  & \new_[62591]_ ;
  assign \new_[62598]_  = A200 & ~A199;
  assign \new_[62601]_  = ~A232 & A203;
  assign \new_[62602]_  = \new_[62601]_  & \new_[62598]_ ;
  assign \new_[62603]_  = \new_[62602]_  & \new_[62595]_ ;
  assign \new_[62606]_  = ~A235 & ~A233;
  assign \new_[62609]_  = ~A268 & ~A267;
  assign \new_[62610]_  = \new_[62609]_  & \new_[62606]_ ;
  assign \new_[62613]_  = ~A298 & ~A269;
  assign \new_[62616]_  = A302 & A299;
  assign \new_[62617]_  = \new_[62616]_  & \new_[62613]_ ;
  assign \new_[62618]_  = \new_[62617]_  & \new_[62610]_ ;
  assign \new_[62621]_  = ~A168 & ~A169;
  assign \new_[62624]_  = A166 & A167;
  assign \new_[62625]_  = \new_[62624]_  & \new_[62621]_ ;
  assign \new_[62628]_  = A200 & ~A199;
  assign \new_[62631]_  = ~A232 & A203;
  assign \new_[62632]_  = \new_[62631]_  & \new_[62628]_ ;
  assign \new_[62633]_  = \new_[62632]_  & \new_[62625]_ ;
  assign \new_[62636]_  = ~A235 & ~A233;
  assign \new_[62639]_  = A266 & A265;
  assign \new_[62640]_  = \new_[62639]_  & \new_[62636]_ ;
  assign \new_[62643]_  = ~A268 & ~A267;
  assign \new_[62646]_  = A300 & A299;
  assign \new_[62647]_  = \new_[62646]_  & \new_[62643]_ ;
  assign \new_[62648]_  = \new_[62647]_  & \new_[62640]_ ;
  assign \new_[62651]_  = ~A168 & ~A169;
  assign \new_[62654]_  = A166 & A167;
  assign \new_[62655]_  = \new_[62654]_  & \new_[62651]_ ;
  assign \new_[62658]_  = A200 & ~A199;
  assign \new_[62661]_  = ~A232 & A203;
  assign \new_[62662]_  = \new_[62661]_  & \new_[62658]_ ;
  assign \new_[62663]_  = \new_[62662]_  & \new_[62655]_ ;
  assign \new_[62666]_  = ~A235 & ~A233;
  assign \new_[62669]_  = A266 & A265;
  assign \new_[62670]_  = \new_[62669]_  & \new_[62666]_ ;
  assign \new_[62673]_  = ~A268 & ~A267;
  assign \new_[62676]_  = A300 & A298;
  assign \new_[62677]_  = \new_[62676]_  & \new_[62673]_ ;
  assign \new_[62678]_  = \new_[62677]_  & \new_[62670]_ ;
  assign \new_[62681]_  = ~A168 & ~A169;
  assign \new_[62684]_  = A166 & A167;
  assign \new_[62685]_  = \new_[62684]_  & \new_[62681]_ ;
  assign \new_[62688]_  = A200 & ~A199;
  assign \new_[62691]_  = ~A232 & A203;
  assign \new_[62692]_  = \new_[62691]_  & \new_[62688]_ ;
  assign \new_[62693]_  = \new_[62692]_  & \new_[62685]_ ;
  assign \new_[62696]_  = ~A235 & ~A233;
  assign \new_[62699]_  = ~A266 & ~A265;
  assign \new_[62700]_  = \new_[62699]_  & \new_[62696]_ ;
  assign \new_[62703]_  = A298 & ~A268;
  assign \new_[62706]_  = A302 & ~A299;
  assign \new_[62707]_  = \new_[62706]_  & \new_[62703]_ ;
  assign \new_[62708]_  = \new_[62707]_  & \new_[62700]_ ;
  assign \new_[62711]_  = ~A168 & ~A169;
  assign \new_[62714]_  = A166 & A167;
  assign \new_[62715]_  = \new_[62714]_  & \new_[62711]_ ;
  assign \new_[62718]_  = A200 & ~A199;
  assign \new_[62721]_  = ~A232 & A203;
  assign \new_[62722]_  = \new_[62721]_  & \new_[62718]_ ;
  assign \new_[62723]_  = \new_[62722]_  & \new_[62715]_ ;
  assign \new_[62726]_  = ~A235 & ~A233;
  assign \new_[62729]_  = ~A266 & ~A265;
  assign \new_[62730]_  = \new_[62729]_  & \new_[62726]_ ;
  assign \new_[62733]_  = ~A298 & ~A268;
  assign \new_[62736]_  = A302 & A299;
  assign \new_[62737]_  = \new_[62736]_  & \new_[62733]_ ;
  assign \new_[62738]_  = \new_[62737]_  & \new_[62730]_ ;
  assign \new_[62741]_  = ~A168 & ~A169;
  assign \new_[62744]_  = A166 & A167;
  assign \new_[62745]_  = \new_[62744]_  & \new_[62741]_ ;
  assign \new_[62748]_  = ~A200 & A199;
  assign \new_[62751]_  = ~A234 & A203;
  assign \new_[62752]_  = \new_[62751]_  & \new_[62748]_ ;
  assign \new_[62753]_  = \new_[62752]_  & \new_[62745]_ ;
  assign \new_[62756]_  = ~A236 & ~A235;
  assign \new_[62759]_  = ~A268 & ~A267;
  assign \new_[62760]_  = \new_[62759]_  & \new_[62756]_ ;
  assign \new_[62763]_  = A298 & ~A269;
  assign \new_[62766]_  = A302 & ~A299;
  assign \new_[62767]_  = \new_[62766]_  & \new_[62763]_ ;
  assign \new_[62768]_  = \new_[62767]_  & \new_[62760]_ ;
  assign \new_[62771]_  = ~A168 & ~A169;
  assign \new_[62774]_  = A166 & A167;
  assign \new_[62775]_  = \new_[62774]_  & \new_[62771]_ ;
  assign \new_[62778]_  = ~A200 & A199;
  assign \new_[62781]_  = ~A234 & A203;
  assign \new_[62782]_  = \new_[62781]_  & \new_[62778]_ ;
  assign \new_[62783]_  = \new_[62782]_  & \new_[62775]_ ;
  assign \new_[62786]_  = ~A236 & ~A235;
  assign \new_[62789]_  = ~A268 & ~A267;
  assign \new_[62790]_  = \new_[62789]_  & \new_[62786]_ ;
  assign \new_[62793]_  = ~A298 & ~A269;
  assign \new_[62796]_  = A302 & A299;
  assign \new_[62797]_  = \new_[62796]_  & \new_[62793]_ ;
  assign \new_[62798]_  = \new_[62797]_  & \new_[62790]_ ;
  assign \new_[62801]_  = ~A168 & ~A169;
  assign \new_[62804]_  = A166 & A167;
  assign \new_[62805]_  = \new_[62804]_  & \new_[62801]_ ;
  assign \new_[62808]_  = ~A200 & A199;
  assign \new_[62811]_  = ~A234 & A203;
  assign \new_[62812]_  = \new_[62811]_  & \new_[62808]_ ;
  assign \new_[62813]_  = \new_[62812]_  & \new_[62805]_ ;
  assign \new_[62816]_  = ~A236 & ~A235;
  assign \new_[62819]_  = A266 & A265;
  assign \new_[62820]_  = \new_[62819]_  & \new_[62816]_ ;
  assign \new_[62823]_  = ~A268 & ~A267;
  assign \new_[62826]_  = A300 & A299;
  assign \new_[62827]_  = \new_[62826]_  & \new_[62823]_ ;
  assign \new_[62828]_  = \new_[62827]_  & \new_[62820]_ ;
  assign \new_[62831]_  = ~A168 & ~A169;
  assign \new_[62834]_  = A166 & A167;
  assign \new_[62835]_  = \new_[62834]_  & \new_[62831]_ ;
  assign \new_[62838]_  = ~A200 & A199;
  assign \new_[62841]_  = ~A234 & A203;
  assign \new_[62842]_  = \new_[62841]_  & \new_[62838]_ ;
  assign \new_[62843]_  = \new_[62842]_  & \new_[62835]_ ;
  assign \new_[62846]_  = ~A236 & ~A235;
  assign \new_[62849]_  = A266 & A265;
  assign \new_[62850]_  = \new_[62849]_  & \new_[62846]_ ;
  assign \new_[62853]_  = ~A268 & ~A267;
  assign \new_[62856]_  = A300 & A298;
  assign \new_[62857]_  = \new_[62856]_  & \new_[62853]_ ;
  assign \new_[62858]_  = \new_[62857]_  & \new_[62850]_ ;
  assign \new_[62861]_  = ~A168 & ~A169;
  assign \new_[62864]_  = A166 & A167;
  assign \new_[62865]_  = \new_[62864]_  & \new_[62861]_ ;
  assign \new_[62868]_  = ~A200 & A199;
  assign \new_[62871]_  = ~A234 & A203;
  assign \new_[62872]_  = \new_[62871]_  & \new_[62868]_ ;
  assign \new_[62873]_  = \new_[62872]_  & \new_[62865]_ ;
  assign \new_[62876]_  = ~A236 & ~A235;
  assign \new_[62879]_  = ~A266 & ~A265;
  assign \new_[62880]_  = \new_[62879]_  & \new_[62876]_ ;
  assign \new_[62883]_  = A298 & ~A268;
  assign \new_[62886]_  = A302 & ~A299;
  assign \new_[62887]_  = \new_[62886]_  & \new_[62883]_ ;
  assign \new_[62888]_  = \new_[62887]_  & \new_[62880]_ ;
  assign \new_[62891]_  = ~A168 & ~A169;
  assign \new_[62894]_  = A166 & A167;
  assign \new_[62895]_  = \new_[62894]_  & \new_[62891]_ ;
  assign \new_[62898]_  = ~A200 & A199;
  assign \new_[62901]_  = ~A234 & A203;
  assign \new_[62902]_  = \new_[62901]_  & \new_[62898]_ ;
  assign \new_[62903]_  = \new_[62902]_  & \new_[62895]_ ;
  assign \new_[62906]_  = ~A236 & ~A235;
  assign \new_[62909]_  = ~A266 & ~A265;
  assign \new_[62910]_  = \new_[62909]_  & \new_[62906]_ ;
  assign \new_[62913]_  = ~A298 & ~A268;
  assign \new_[62916]_  = A302 & A299;
  assign \new_[62917]_  = \new_[62916]_  & \new_[62913]_ ;
  assign \new_[62918]_  = \new_[62917]_  & \new_[62910]_ ;
  assign \new_[62921]_  = ~A168 & ~A169;
  assign \new_[62924]_  = A166 & A167;
  assign \new_[62925]_  = \new_[62924]_  & \new_[62921]_ ;
  assign \new_[62928]_  = ~A200 & A199;
  assign \new_[62931]_  = A232 & A203;
  assign \new_[62932]_  = \new_[62931]_  & \new_[62928]_ ;
  assign \new_[62933]_  = \new_[62932]_  & \new_[62925]_ ;
  assign \new_[62936]_  = ~A234 & A233;
  assign \new_[62939]_  = ~A267 & ~A235;
  assign \new_[62940]_  = \new_[62939]_  & \new_[62936]_ ;
  assign \new_[62943]_  = ~A269 & ~A268;
  assign \new_[62946]_  = A300 & A299;
  assign \new_[62947]_  = \new_[62946]_  & \new_[62943]_ ;
  assign \new_[62948]_  = \new_[62947]_  & \new_[62940]_ ;
  assign \new_[62951]_  = ~A168 & ~A169;
  assign \new_[62954]_  = A166 & A167;
  assign \new_[62955]_  = \new_[62954]_  & \new_[62951]_ ;
  assign \new_[62958]_  = ~A200 & A199;
  assign \new_[62961]_  = A232 & A203;
  assign \new_[62962]_  = \new_[62961]_  & \new_[62958]_ ;
  assign \new_[62963]_  = \new_[62962]_  & \new_[62955]_ ;
  assign \new_[62966]_  = ~A234 & A233;
  assign \new_[62969]_  = ~A267 & ~A235;
  assign \new_[62970]_  = \new_[62969]_  & \new_[62966]_ ;
  assign \new_[62973]_  = ~A269 & ~A268;
  assign \new_[62976]_  = A300 & A298;
  assign \new_[62977]_  = \new_[62976]_  & \new_[62973]_ ;
  assign \new_[62978]_  = \new_[62977]_  & \new_[62970]_ ;
  assign \new_[62981]_  = ~A168 & ~A169;
  assign \new_[62984]_  = A166 & A167;
  assign \new_[62985]_  = \new_[62984]_  & \new_[62981]_ ;
  assign \new_[62988]_  = ~A200 & A199;
  assign \new_[62991]_  = A232 & A203;
  assign \new_[62992]_  = \new_[62991]_  & \new_[62988]_ ;
  assign \new_[62993]_  = \new_[62992]_  & \new_[62985]_ ;
  assign \new_[62996]_  = ~A234 & A233;
  assign \new_[62999]_  = A265 & ~A235;
  assign \new_[63000]_  = \new_[62999]_  & \new_[62996]_ ;
  assign \new_[63003]_  = ~A267 & A266;
  assign \new_[63006]_  = A301 & ~A268;
  assign \new_[63007]_  = \new_[63006]_  & \new_[63003]_ ;
  assign \new_[63008]_  = \new_[63007]_  & \new_[63000]_ ;
  assign \new_[63011]_  = ~A168 & ~A169;
  assign \new_[63014]_  = A166 & A167;
  assign \new_[63015]_  = \new_[63014]_  & \new_[63011]_ ;
  assign \new_[63018]_  = ~A200 & A199;
  assign \new_[63021]_  = A232 & A203;
  assign \new_[63022]_  = \new_[63021]_  & \new_[63018]_ ;
  assign \new_[63023]_  = \new_[63022]_  & \new_[63015]_ ;
  assign \new_[63026]_  = ~A234 & A233;
  assign \new_[63029]_  = ~A265 & ~A235;
  assign \new_[63030]_  = \new_[63029]_  & \new_[63026]_ ;
  assign \new_[63033]_  = ~A268 & ~A266;
  assign \new_[63036]_  = A300 & A299;
  assign \new_[63037]_  = \new_[63036]_  & \new_[63033]_ ;
  assign \new_[63038]_  = \new_[63037]_  & \new_[63030]_ ;
  assign \new_[63041]_  = ~A168 & ~A169;
  assign \new_[63044]_  = A166 & A167;
  assign \new_[63045]_  = \new_[63044]_  & \new_[63041]_ ;
  assign \new_[63048]_  = ~A200 & A199;
  assign \new_[63051]_  = A232 & A203;
  assign \new_[63052]_  = \new_[63051]_  & \new_[63048]_ ;
  assign \new_[63053]_  = \new_[63052]_  & \new_[63045]_ ;
  assign \new_[63056]_  = ~A234 & A233;
  assign \new_[63059]_  = ~A265 & ~A235;
  assign \new_[63060]_  = \new_[63059]_  & \new_[63056]_ ;
  assign \new_[63063]_  = ~A268 & ~A266;
  assign \new_[63066]_  = A300 & A298;
  assign \new_[63067]_  = \new_[63066]_  & \new_[63063]_ ;
  assign \new_[63068]_  = \new_[63067]_  & \new_[63060]_ ;
  assign \new_[63071]_  = ~A168 & ~A169;
  assign \new_[63074]_  = A166 & A167;
  assign \new_[63075]_  = \new_[63074]_  & \new_[63071]_ ;
  assign \new_[63078]_  = ~A200 & A199;
  assign \new_[63081]_  = ~A232 & A203;
  assign \new_[63082]_  = \new_[63081]_  & \new_[63078]_ ;
  assign \new_[63083]_  = \new_[63082]_  & \new_[63075]_ ;
  assign \new_[63086]_  = ~A235 & ~A233;
  assign \new_[63089]_  = ~A268 & ~A267;
  assign \new_[63090]_  = \new_[63089]_  & \new_[63086]_ ;
  assign \new_[63093]_  = A298 & ~A269;
  assign \new_[63096]_  = A302 & ~A299;
  assign \new_[63097]_  = \new_[63096]_  & \new_[63093]_ ;
  assign \new_[63098]_  = \new_[63097]_  & \new_[63090]_ ;
  assign \new_[63101]_  = ~A168 & ~A169;
  assign \new_[63104]_  = A166 & A167;
  assign \new_[63105]_  = \new_[63104]_  & \new_[63101]_ ;
  assign \new_[63108]_  = ~A200 & A199;
  assign \new_[63111]_  = ~A232 & A203;
  assign \new_[63112]_  = \new_[63111]_  & \new_[63108]_ ;
  assign \new_[63113]_  = \new_[63112]_  & \new_[63105]_ ;
  assign \new_[63116]_  = ~A235 & ~A233;
  assign \new_[63119]_  = ~A268 & ~A267;
  assign \new_[63120]_  = \new_[63119]_  & \new_[63116]_ ;
  assign \new_[63123]_  = ~A298 & ~A269;
  assign \new_[63126]_  = A302 & A299;
  assign \new_[63127]_  = \new_[63126]_  & \new_[63123]_ ;
  assign \new_[63128]_  = \new_[63127]_  & \new_[63120]_ ;
  assign \new_[63131]_  = ~A168 & ~A169;
  assign \new_[63134]_  = A166 & A167;
  assign \new_[63135]_  = \new_[63134]_  & \new_[63131]_ ;
  assign \new_[63138]_  = ~A200 & A199;
  assign \new_[63141]_  = ~A232 & A203;
  assign \new_[63142]_  = \new_[63141]_  & \new_[63138]_ ;
  assign \new_[63143]_  = \new_[63142]_  & \new_[63135]_ ;
  assign \new_[63146]_  = ~A235 & ~A233;
  assign \new_[63149]_  = A266 & A265;
  assign \new_[63150]_  = \new_[63149]_  & \new_[63146]_ ;
  assign \new_[63153]_  = ~A268 & ~A267;
  assign \new_[63156]_  = A300 & A299;
  assign \new_[63157]_  = \new_[63156]_  & \new_[63153]_ ;
  assign \new_[63158]_  = \new_[63157]_  & \new_[63150]_ ;
  assign \new_[63161]_  = ~A168 & ~A169;
  assign \new_[63164]_  = A166 & A167;
  assign \new_[63165]_  = \new_[63164]_  & \new_[63161]_ ;
  assign \new_[63168]_  = ~A200 & A199;
  assign \new_[63171]_  = ~A232 & A203;
  assign \new_[63172]_  = \new_[63171]_  & \new_[63168]_ ;
  assign \new_[63173]_  = \new_[63172]_  & \new_[63165]_ ;
  assign \new_[63176]_  = ~A235 & ~A233;
  assign \new_[63179]_  = A266 & A265;
  assign \new_[63180]_  = \new_[63179]_  & \new_[63176]_ ;
  assign \new_[63183]_  = ~A268 & ~A267;
  assign \new_[63186]_  = A300 & A298;
  assign \new_[63187]_  = \new_[63186]_  & \new_[63183]_ ;
  assign \new_[63188]_  = \new_[63187]_  & \new_[63180]_ ;
  assign \new_[63191]_  = ~A168 & ~A169;
  assign \new_[63194]_  = A166 & A167;
  assign \new_[63195]_  = \new_[63194]_  & \new_[63191]_ ;
  assign \new_[63198]_  = ~A200 & A199;
  assign \new_[63201]_  = ~A232 & A203;
  assign \new_[63202]_  = \new_[63201]_  & \new_[63198]_ ;
  assign \new_[63203]_  = \new_[63202]_  & \new_[63195]_ ;
  assign \new_[63206]_  = ~A235 & ~A233;
  assign \new_[63209]_  = ~A266 & ~A265;
  assign \new_[63210]_  = \new_[63209]_  & \new_[63206]_ ;
  assign \new_[63213]_  = A298 & ~A268;
  assign \new_[63216]_  = A302 & ~A299;
  assign \new_[63217]_  = \new_[63216]_  & \new_[63213]_ ;
  assign \new_[63218]_  = \new_[63217]_  & \new_[63210]_ ;
  assign \new_[63221]_  = ~A168 & ~A169;
  assign \new_[63224]_  = A166 & A167;
  assign \new_[63225]_  = \new_[63224]_  & \new_[63221]_ ;
  assign \new_[63228]_  = ~A200 & A199;
  assign \new_[63231]_  = ~A232 & A203;
  assign \new_[63232]_  = \new_[63231]_  & \new_[63228]_ ;
  assign \new_[63233]_  = \new_[63232]_  & \new_[63225]_ ;
  assign \new_[63236]_  = ~A235 & ~A233;
  assign \new_[63239]_  = ~A266 & ~A265;
  assign \new_[63240]_  = \new_[63239]_  & \new_[63236]_ ;
  assign \new_[63243]_  = ~A298 & ~A268;
  assign \new_[63246]_  = A302 & A299;
  assign \new_[63247]_  = \new_[63246]_  & \new_[63243]_ ;
  assign \new_[63248]_  = \new_[63247]_  & \new_[63240]_ ;
  assign \new_[63251]_  = ~A169 & ~A170;
  assign \new_[63254]_  = A199 & ~A168;
  assign \new_[63255]_  = \new_[63254]_  & \new_[63251]_ ;
  assign \new_[63258]_  = A232 & A201;
  assign \new_[63261]_  = ~A234 & A233;
  assign \new_[63262]_  = \new_[63261]_  & \new_[63258]_ ;
  assign \new_[63263]_  = \new_[63262]_  & \new_[63255]_ ;
  assign \new_[63266]_  = A265 & ~A235;
  assign \new_[63269]_  = ~A267 & A266;
  assign \new_[63270]_  = \new_[63269]_  & \new_[63266]_ ;
  assign \new_[63273]_  = A298 & ~A268;
  assign \new_[63276]_  = A302 & ~A299;
  assign \new_[63277]_  = \new_[63276]_  & \new_[63273]_ ;
  assign \new_[63278]_  = \new_[63277]_  & \new_[63270]_ ;
  assign \new_[63281]_  = ~A169 & ~A170;
  assign \new_[63284]_  = A199 & ~A168;
  assign \new_[63285]_  = \new_[63284]_  & \new_[63281]_ ;
  assign \new_[63288]_  = A232 & A201;
  assign \new_[63291]_  = ~A234 & A233;
  assign \new_[63292]_  = \new_[63291]_  & \new_[63288]_ ;
  assign \new_[63293]_  = \new_[63292]_  & \new_[63285]_ ;
  assign \new_[63296]_  = A265 & ~A235;
  assign \new_[63299]_  = ~A267 & A266;
  assign \new_[63300]_  = \new_[63299]_  & \new_[63296]_ ;
  assign \new_[63303]_  = ~A298 & ~A268;
  assign \new_[63306]_  = A302 & A299;
  assign \new_[63307]_  = \new_[63306]_  & \new_[63303]_ ;
  assign \new_[63308]_  = \new_[63307]_  & \new_[63300]_ ;
  assign \new_[63311]_  = ~A169 & ~A170;
  assign \new_[63314]_  = A200 & ~A168;
  assign \new_[63315]_  = \new_[63314]_  & \new_[63311]_ ;
  assign \new_[63318]_  = A232 & A201;
  assign \new_[63321]_  = ~A234 & A233;
  assign \new_[63322]_  = \new_[63321]_  & \new_[63318]_ ;
  assign \new_[63323]_  = \new_[63322]_  & \new_[63315]_ ;
  assign \new_[63326]_  = A265 & ~A235;
  assign \new_[63329]_  = ~A267 & A266;
  assign \new_[63330]_  = \new_[63329]_  & \new_[63326]_ ;
  assign \new_[63333]_  = A298 & ~A268;
  assign \new_[63336]_  = A302 & ~A299;
  assign \new_[63337]_  = \new_[63336]_  & \new_[63333]_ ;
  assign \new_[63338]_  = \new_[63337]_  & \new_[63330]_ ;
  assign \new_[63341]_  = ~A169 & ~A170;
  assign \new_[63344]_  = A200 & ~A168;
  assign \new_[63345]_  = \new_[63344]_  & \new_[63341]_ ;
  assign \new_[63348]_  = A232 & A201;
  assign \new_[63351]_  = ~A234 & A233;
  assign \new_[63352]_  = \new_[63351]_  & \new_[63348]_ ;
  assign \new_[63353]_  = \new_[63352]_  & \new_[63345]_ ;
  assign \new_[63356]_  = A265 & ~A235;
  assign \new_[63359]_  = ~A267 & A266;
  assign \new_[63360]_  = \new_[63359]_  & \new_[63356]_ ;
  assign \new_[63363]_  = ~A298 & ~A268;
  assign \new_[63366]_  = A302 & A299;
  assign \new_[63367]_  = \new_[63366]_  & \new_[63363]_ ;
  assign \new_[63368]_  = \new_[63367]_  & \new_[63360]_ ;
  assign \new_[63371]_  = ~A169 & ~A170;
  assign \new_[63374]_  = ~A199 & ~A168;
  assign \new_[63375]_  = \new_[63374]_  & \new_[63371]_ ;
  assign \new_[63378]_  = A203 & A200;
  assign \new_[63381]_  = ~A235 & ~A234;
  assign \new_[63382]_  = \new_[63381]_  & \new_[63378]_ ;
  assign \new_[63383]_  = \new_[63382]_  & \new_[63375]_ ;
  assign \new_[63386]_  = A265 & ~A236;
  assign \new_[63389]_  = ~A267 & A266;
  assign \new_[63390]_  = \new_[63389]_  & \new_[63386]_ ;
  assign \new_[63393]_  = A298 & ~A268;
  assign \new_[63396]_  = A302 & ~A299;
  assign \new_[63397]_  = \new_[63396]_  & \new_[63393]_ ;
  assign \new_[63398]_  = \new_[63397]_  & \new_[63390]_ ;
  assign \new_[63401]_  = ~A169 & ~A170;
  assign \new_[63404]_  = ~A199 & ~A168;
  assign \new_[63405]_  = \new_[63404]_  & \new_[63401]_ ;
  assign \new_[63408]_  = A203 & A200;
  assign \new_[63411]_  = ~A235 & ~A234;
  assign \new_[63412]_  = \new_[63411]_  & \new_[63408]_ ;
  assign \new_[63413]_  = \new_[63412]_  & \new_[63405]_ ;
  assign \new_[63416]_  = A265 & ~A236;
  assign \new_[63419]_  = ~A267 & A266;
  assign \new_[63420]_  = \new_[63419]_  & \new_[63416]_ ;
  assign \new_[63423]_  = ~A298 & ~A268;
  assign \new_[63426]_  = A302 & A299;
  assign \new_[63427]_  = \new_[63426]_  & \new_[63423]_ ;
  assign \new_[63428]_  = \new_[63427]_  & \new_[63420]_ ;
  assign \new_[63431]_  = ~A169 & ~A170;
  assign \new_[63434]_  = ~A199 & ~A168;
  assign \new_[63435]_  = \new_[63434]_  & \new_[63431]_ ;
  assign \new_[63438]_  = A203 & A200;
  assign \new_[63441]_  = A233 & A232;
  assign \new_[63442]_  = \new_[63441]_  & \new_[63438]_ ;
  assign \new_[63443]_  = \new_[63442]_  & \new_[63435]_ ;
  assign \new_[63446]_  = ~A235 & ~A234;
  assign \new_[63449]_  = ~A268 & ~A267;
  assign \new_[63450]_  = \new_[63449]_  & \new_[63446]_ ;
  assign \new_[63453]_  = A298 & ~A269;
  assign \new_[63456]_  = A302 & ~A299;
  assign \new_[63457]_  = \new_[63456]_  & \new_[63453]_ ;
  assign \new_[63458]_  = \new_[63457]_  & \new_[63450]_ ;
  assign \new_[63461]_  = ~A169 & ~A170;
  assign \new_[63464]_  = ~A199 & ~A168;
  assign \new_[63465]_  = \new_[63464]_  & \new_[63461]_ ;
  assign \new_[63468]_  = A203 & A200;
  assign \new_[63471]_  = A233 & A232;
  assign \new_[63472]_  = \new_[63471]_  & \new_[63468]_ ;
  assign \new_[63473]_  = \new_[63472]_  & \new_[63465]_ ;
  assign \new_[63476]_  = ~A235 & ~A234;
  assign \new_[63479]_  = ~A268 & ~A267;
  assign \new_[63480]_  = \new_[63479]_  & \new_[63476]_ ;
  assign \new_[63483]_  = ~A298 & ~A269;
  assign \new_[63486]_  = A302 & A299;
  assign \new_[63487]_  = \new_[63486]_  & \new_[63483]_ ;
  assign \new_[63488]_  = \new_[63487]_  & \new_[63480]_ ;
  assign \new_[63491]_  = ~A169 & ~A170;
  assign \new_[63494]_  = ~A199 & ~A168;
  assign \new_[63495]_  = \new_[63494]_  & \new_[63491]_ ;
  assign \new_[63498]_  = A203 & A200;
  assign \new_[63501]_  = A233 & A232;
  assign \new_[63502]_  = \new_[63501]_  & \new_[63498]_ ;
  assign \new_[63503]_  = \new_[63502]_  & \new_[63495]_ ;
  assign \new_[63506]_  = ~A235 & ~A234;
  assign \new_[63509]_  = A266 & A265;
  assign \new_[63510]_  = \new_[63509]_  & \new_[63506]_ ;
  assign \new_[63513]_  = ~A268 & ~A267;
  assign \new_[63516]_  = A300 & A299;
  assign \new_[63517]_  = \new_[63516]_  & \new_[63513]_ ;
  assign \new_[63518]_  = \new_[63517]_  & \new_[63510]_ ;
  assign \new_[63521]_  = ~A169 & ~A170;
  assign \new_[63524]_  = ~A199 & ~A168;
  assign \new_[63525]_  = \new_[63524]_  & \new_[63521]_ ;
  assign \new_[63528]_  = A203 & A200;
  assign \new_[63531]_  = A233 & A232;
  assign \new_[63532]_  = \new_[63531]_  & \new_[63528]_ ;
  assign \new_[63533]_  = \new_[63532]_  & \new_[63525]_ ;
  assign \new_[63536]_  = ~A235 & ~A234;
  assign \new_[63539]_  = A266 & A265;
  assign \new_[63540]_  = \new_[63539]_  & \new_[63536]_ ;
  assign \new_[63543]_  = ~A268 & ~A267;
  assign \new_[63546]_  = A300 & A298;
  assign \new_[63547]_  = \new_[63546]_  & \new_[63543]_ ;
  assign \new_[63548]_  = \new_[63547]_  & \new_[63540]_ ;
  assign \new_[63551]_  = ~A169 & ~A170;
  assign \new_[63554]_  = ~A199 & ~A168;
  assign \new_[63555]_  = \new_[63554]_  & \new_[63551]_ ;
  assign \new_[63558]_  = A203 & A200;
  assign \new_[63561]_  = A233 & A232;
  assign \new_[63562]_  = \new_[63561]_  & \new_[63558]_ ;
  assign \new_[63563]_  = \new_[63562]_  & \new_[63555]_ ;
  assign \new_[63566]_  = ~A235 & ~A234;
  assign \new_[63569]_  = ~A266 & ~A265;
  assign \new_[63570]_  = \new_[63569]_  & \new_[63566]_ ;
  assign \new_[63573]_  = A298 & ~A268;
  assign \new_[63576]_  = A302 & ~A299;
  assign \new_[63577]_  = \new_[63576]_  & \new_[63573]_ ;
  assign \new_[63578]_  = \new_[63577]_  & \new_[63570]_ ;
  assign \new_[63581]_  = ~A169 & ~A170;
  assign \new_[63584]_  = ~A199 & ~A168;
  assign \new_[63585]_  = \new_[63584]_  & \new_[63581]_ ;
  assign \new_[63588]_  = A203 & A200;
  assign \new_[63591]_  = A233 & A232;
  assign \new_[63592]_  = \new_[63591]_  & \new_[63588]_ ;
  assign \new_[63593]_  = \new_[63592]_  & \new_[63585]_ ;
  assign \new_[63596]_  = ~A235 & ~A234;
  assign \new_[63599]_  = ~A266 & ~A265;
  assign \new_[63600]_  = \new_[63599]_  & \new_[63596]_ ;
  assign \new_[63603]_  = ~A298 & ~A268;
  assign \new_[63606]_  = A302 & A299;
  assign \new_[63607]_  = \new_[63606]_  & \new_[63603]_ ;
  assign \new_[63608]_  = \new_[63607]_  & \new_[63600]_ ;
  assign \new_[63611]_  = ~A169 & ~A170;
  assign \new_[63614]_  = ~A199 & ~A168;
  assign \new_[63615]_  = \new_[63614]_  & \new_[63611]_ ;
  assign \new_[63618]_  = A203 & A200;
  assign \new_[63621]_  = ~A233 & ~A232;
  assign \new_[63622]_  = \new_[63621]_  & \new_[63618]_ ;
  assign \new_[63623]_  = \new_[63622]_  & \new_[63615]_ ;
  assign \new_[63626]_  = A265 & ~A235;
  assign \new_[63629]_  = ~A267 & A266;
  assign \new_[63630]_  = \new_[63629]_  & \new_[63626]_ ;
  assign \new_[63633]_  = A298 & ~A268;
  assign \new_[63636]_  = A302 & ~A299;
  assign \new_[63637]_  = \new_[63636]_  & \new_[63633]_ ;
  assign \new_[63638]_  = \new_[63637]_  & \new_[63630]_ ;
  assign \new_[63641]_  = ~A169 & ~A170;
  assign \new_[63644]_  = ~A199 & ~A168;
  assign \new_[63645]_  = \new_[63644]_  & \new_[63641]_ ;
  assign \new_[63648]_  = A203 & A200;
  assign \new_[63651]_  = ~A233 & ~A232;
  assign \new_[63652]_  = \new_[63651]_  & \new_[63648]_ ;
  assign \new_[63653]_  = \new_[63652]_  & \new_[63645]_ ;
  assign \new_[63656]_  = A265 & ~A235;
  assign \new_[63659]_  = ~A267 & A266;
  assign \new_[63660]_  = \new_[63659]_  & \new_[63656]_ ;
  assign \new_[63663]_  = ~A298 & ~A268;
  assign \new_[63666]_  = A302 & A299;
  assign \new_[63667]_  = \new_[63666]_  & \new_[63663]_ ;
  assign \new_[63668]_  = \new_[63667]_  & \new_[63660]_ ;
  assign \new_[63671]_  = ~A169 & ~A170;
  assign \new_[63674]_  = A199 & ~A168;
  assign \new_[63675]_  = \new_[63674]_  & \new_[63671]_ ;
  assign \new_[63678]_  = A203 & ~A200;
  assign \new_[63681]_  = ~A235 & ~A234;
  assign \new_[63682]_  = \new_[63681]_  & \new_[63678]_ ;
  assign \new_[63683]_  = \new_[63682]_  & \new_[63675]_ ;
  assign \new_[63686]_  = A265 & ~A236;
  assign \new_[63689]_  = ~A267 & A266;
  assign \new_[63690]_  = \new_[63689]_  & \new_[63686]_ ;
  assign \new_[63693]_  = A298 & ~A268;
  assign \new_[63696]_  = A302 & ~A299;
  assign \new_[63697]_  = \new_[63696]_  & \new_[63693]_ ;
  assign \new_[63698]_  = \new_[63697]_  & \new_[63690]_ ;
  assign \new_[63701]_  = ~A169 & ~A170;
  assign \new_[63704]_  = A199 & ~A168;
  assign \new_[63705]_  = \new_[63704]_  & \new_[63701]_ ;
  assign \new_[63708]_  = A203 & ~A200;
  assign \new_[63711]_  = ~A235 & ~A234;
  assign \new_[63712]_  = \new_[63711]_  & \new_[63708]_ ;
  assign \new_[63713]_  = \new_[63712]_  & \new_[63705]_ ;
  assign \new_[63716]_  = A265 & ~A236;
  assign \new_[63719]_  = ~A267 & A266;
  assign \new_[63720]_  = \new_[63719]_  & \new_[63716]_ ;
  assign \new_[63723]_  = ~A298 & ~A268;
  assign \new_[63726]_  = A302 & A299;
  assign \new_[63727]_  = \new_[63726]_  & \new_[63723]_ ;
  assign \new_[63728]_  = \new_[63727]_  & \new_[63720]_ ;
  assign \new_[63731]_  = ~A169 & ~A170;
  assign \new_[63734]_  = A199 & ~A168;
  assign \new_[63735]_  = \new_[63734]_  & \new_[63731]_ ;
  assign \new_[63738]_  = A203 & ~A200;
  assign \new_[63741]_  = A233 & A232;
  assign \new_[63742]_  = \new_[63741]_  & \new_[63738]_ ;
  assign \new_[63743]_  = \new_[63742]_  & \new_[63735]_ ;
  assign \new_[63746]_  = ~A235 & ~A234;
  assign \new_[63749]_  = ~A268 & ~A267;
  assign \new_[63750]_  = \new_[63749]_  & \new_[63746]_ ;
  assign \new_[63753]_  = A298 & ~A269;
  assign \new_[63756]_  = A302 & ~A299;
  assign \new_[63757]_  = \new_[63756]_  & \new_[63753]_ ;
  assign \new_[63758]_  = \new_[63757]_  & \new_[63750]_ ;
  assign \new_[63761]_  = ~A169 & ~A170;
  assign \new_[63764]_  = A199 & ~A168;
  assign \new_[63765]_  = \new_[63764]_  & \new_[63761]_ ;
  assign \new_[63768]_  = A203 & ~A200;
  assign \new_[63771]_  = A233 & A232;
  assign \new_[63772]_  = \new_[63771]_  & \new_[63768]_ ;
  assign \new_[63773]_  = \new_[63772]_  & \new_[63765]_ ;
  assign \new_[63776]_  = ~A235 & ~A234;
  assign \new_[63779]_  = ~A268 & ~A267;
  assign \new_[63780]_  = \new_[63779]_  & \new_[63776]_ ;
  assign \new_[63783]_  = ~A298 & ~A269;
  assign \new_[63786]_  = A302 & A299;
  assign \new_[63787]_  = \new_[63786]_  & \new_[63783]_ ;
  assign \new_[63788]_  = \new_[63787]_  & \new_[63780]_ ;
  assign \new_[63791]_  = ~A169 & ~A170;
  assign \new_[63794]_  = A199 & ~A168;
  assign \new_[63795]_  = \new_[63794]_  & \new_[63791]_ ;
  assign \new_[63798]_  = A203 & ~A200;
  assign \new_[63801]_  = A233 & A232;
  assign \new_[63802]_  = \new_[63801]_  & \new_[63798]_ ;
  assign \new_[63803]_  = \new_[63802]_  & \new_[63795]_ ;
  assign \new_[63806]_  = ~A235 & ~A234;
  assign \new_[63809]_  = A266 & A265;
  assign \new_[63810]_  = \new_[63809]_  & \new_[63806]_ ;
  assign \new_[63813]_  = ~A268 & ~A267;
  assign \new_[63816]_  = A300 & A299;
  assign \new_[63817]_  = \new_[63816]_  & \new_[63813]_ ;
  assign \new_[63818]_  = \new_[63817]_  & \new_[63810]_ ;
  assign \new_[63821]_  = ~A169 & ~A170;
  assign \new_[63824]_  = A199 & ~A168;
  assign \new_[63825]_  = \new_[63824]_  & \new_[63821]_ ;
  assign \new_[63828]_  = A203 & ~A200;
  assign \new_[63831]_  = A233 & A232;
  assign \new_[63832]_  = \new_[63831]_  & \new_[63828]_ ;
  assign \new_[63833]_  = \new_[63832]_  & \new_[63825]_ ;
  assign \new_[63836]_  = ~A235 & ~A234;
  assign \new_[63839]_  = A266 & A265;
  assign \new_[63840]_  = \new_[63839]_  & \new_[63836]_ ;
  assign \new_[63843]_  = ~A268 & ~A267;
  assign \new_[63846]_  = A300 & A298;
  assign \new_[63847]_  = \new_[63846]_  & \new_[63843]_ ;
  assign \new_[63848]_  = \new_[63847]_  & \new_[63840]_ ;
  assign \new_[63851]_  = ~A169 & ~A170;
  assign \new_[63854]_  = A199 & ~A168;
  assign \new_[63855]_  = \new_[63854]_  & \new_[63851]_ ;
  assign \new_[63858]_  = A203 & ~A200;
  assign \new_[63861]_  = A233 & A232;
  assign \new_[63862]_  = \new_[63861]_  & \new_[63858]_ ;
  assign \new_[63863]_  = \new_[63862]_  & \new_[63855]_ ;
  assign \new_[63866]_  = ~A235 & ~A234;
  assign \new_[63869]_  = ~A266 & ~A265;
  assign \new_[63870]_  = \new_[63869]_  & \new_[63866]_ ;
  assign \new_[63873]_  = A298 & ~A268;
  assign \new_[63876]_  = A302 & ~A299;
  assign \new_[63877]_  = \new_[63876]_  & \new_[63873]_ ;
  assign \new_[63878]_  = \new_[63877]_  & \new_[63870]_ ;
  assign \new_[63881]_  = ~A169 & ~A170;
  assign \new_[63884]_  = A199 & ~A168;
  assign \new_[63885]_  = \new_[63884]_  & \new_[63881]_ ;
  assign \new_[63888]_  = A203 & ~A200;
  assign \new_[63891]_  = A233 & A232;
  assign \new_[63892]_  = \new_[63891]_  & \new_[63888]_ ;
  assign \new_[63893]_  = \new_[63892]_  & \new_[63885]_ ;
  assign \new_[63896]_  = ~A235 & ~A234;
  assign \new_[63899]_  = ~A266 & ~A265;
  assign \new_[63900]_  = \new_[63899]_  & \new_[63896]_ ;
  assign \new_[63903]_  = ~A298 & ~A268;
  assign \new_[63906]_  = A302 & A299;
  assign \new_[63907]_  = \new_[63906]_  & \new_[63903]_ ;
  assign \new_[63908]_  = \new_[63907]_  & \new_[63900]_ ;
  assign \new_[63911]_  = ~A169 & ~A170;
  assign \new_[63914]_  = A199 & ~A168;
  assign \new_[63915]_  = \new_[63914]_  & \new_[63911]_ ;
  assign \new_[63918]_  = A203 & ~A200;
  assign \new_[63921]_  = ~A233 & ~A232;
  assign \new_[63922]_  = \new_[63921]_  & \new_[63918]_ ;
  assign \new_[63923]_  = \new_[63922]_  & \new_[63915]_ ;
  assign \new_[63926]_  = A265 & ~A235;
  assign \new_[63929]_  = ~A267 & A266;
  assign \new_[63930]_  = \new_[63929]_  & \new_[63926]_ ;
  assign \new_[63933]_  = A298 & ~A268;
  assign \new_[63936]_  = A302 & ~A299;
  assign \new_[63937]_  = \new_[63936]_  & \new_[63933]_ ;
  assign \new_[63938]_  = \new_[63937]_  & \new_[63930]_ ;
  assign \new_[63941]_  = ~A169 & ~A170;
  assign \new_[63944]_  = A199 & ~A168;
  assign \new_[63945]_  = \new_[63944]_  & \new_[63941]_ ;
  assign \new_[63948]_  = A203 & ~A200;
  assign \new_[63951]_  = ~A233 & ~A232;
  assign \new_[63952]_  = \new_[63951]_  & \new_[63948]_ ;
  assign \new_[63953]_  = \new_[63952]_  & \new_[63945]_ ;
  assign \new_[63956]_  = A265 & ~A235;
  assign \new_[63959]_  = ~A267 & A266;
  assign \new_[63960]_  = \new_[63959]_  & \new_[63956]_ ;
  assign \new_[63963]_  = ~A298 & ~A268;
  assign \new_[63966]_  = A302 & A299;
  assign \new_[63967]_  = \new_[63966]_  & \new_[63963]_ ;
  assign \new_[63968]_  = \new_[63967]_  & \new_[63960]_ ;
  assign \new_[63971]_  = A166 & A168;
  assign \new_[63974]_  = A200 & A199;
  assign \new_[63975]_  = \new_[63974]_  & \new_[63971]_ ;
  assign \new_[63978]_  = ~A202 & ~A201;
  assign \new_[63981]_  = A233 & A232;
  assign \new_[63982]_  = \new_[63981]_  & \new_[63978]_ ;
  assign \new_[63983]_  = \new_[63982]_  & \new_[63975]_ ;
  assign \new_[63986]_  = ~A235 & ~A234;
  assign \new_[63989]_  = A266 & A265;
  assign \new_[63990]_  = \new_[63989]_  & \new_[63986]_ ;
  assign \new_[63993]_  = ~A268 & ~A267;
  assign \new_[63997]_  = A302 & ~A299;
  assign \new_[63998]_  = A298 & \new_[63997]_ ;
  assign \new_[63999]_  = \new_[63998]_  & \new_[63993]_ ;
  assign \new_[64000]_  = \new_[63999]_  & \new_[63990]_ ;
  assign \new_[64003]_  = A166 & A168;
  assign \new_[64006]_  = A200 & A199;
  assign \new_[64007]_  = \new_[64006]_  & \new_[64003]_ ;
  assign \new_[64010]_  = ~A202 & ~A201;
  assign \new_[64013]_  = A233 & A232;
  assign \new_[64014]_  = \new_[64013]_  & \new_[64010]_ ;
  assign \new_[64015]_  = \new_[64014]_  & \new_[64007]_ ;
  assign \new_[64018]_  = ~A235 & ~A234;
  assign \new_[64021]_  = A266 & A265;
  assign \new_[64022]_  = \new_[64021]_  & \new_[64018]_ ;
  assign \new_[64025]_  = ~A268 & ~A267;
  assign \new_[64029]_  = A302 & A299;
  assign \new_[64030]_  = ~A298 & \new_[64029]_ ;
  assign \new_[64031]_  = \new_[64030]_  & \new_[64025]_ ;
  assign \new_[64032]_  = \new_[64031]_  & \new_[64022]_ ;
  assign \new_[64035]_  = A167 & A168;
  assign \new_[64038]_  = A200 & A199;
  assign \new_[64039]_  = \new_[64038]_  & \new_[64035]_ ;
  assign \new_[64042]_  = ~A202 & ~A201;
  assign \new_[64045]_  = A233 & A232;
  assign \new_[64046]_  = \new_[64045]_  & \new_[64042]_ ;
  assign \new_[64047]_  = \new_[64046]_  & \new_[64039]_ ;
  assign \new_[64050]_  = ~A235 & ~A234;
  assign \new_[64053]_  = A266 & A265;
  assign \new_[64054]_  = \new_[64053]_  & \new_[64050]_ ;
  assign \new_[64057]_  = ~A268 & ~A267;
  assign \new_[64061]_  = A302 & ~A299;
  assign \new_[64062]_  = A298 & \new_[64061]_ ;
  assign \new_[64063]_  = \new_[64062]_  & \new_[64057]_ ;
  assign \new_[64064]_  = \new_[64063]_  & \new_[64054]_ ;
  assign \new_[64067]_  = A167 & A168;
  assign \new_[64070]_  = A200 & A199;
  assign \new_[64071]_  = \new_[64070]_  & \new_[64067]_ ;
  assign \new_[64074]_  = ~A202 & ~A201;
  assign \new_[64077]_  = A233 & A232;
  assign \new_[64078]_  = \new_[64077]_  & \new_[64074]_ ;
  assign \new_[64079]_  = \new_[64078]_  & \new_[64071]_ ;
  assign \new_[64082]_  = ~A235 & ~A234;
  assign \new_[64085]_  = A266 & A265;
  assign \new_[64086]_  = \new_[64085]_  & \new_[64082]_ ;
  assign \new_[64089]_  = ~A268 & ~A267;
  assign \new_[64093]_  = A302 & A299;
  assign \new_[64094]_  = ~A298 & \new_[64093]_ ;
  assign \new_[64095]_  = \new_[64094]_  & \new_[64089]_ ;
  assign \new_[64096]_  = \new_[64095]_  & \new_[64086]_ ;
  assign \new_[64099]_  = A167 & A170;
  assign \new_[64102]_  = ~A201 & ~A166;
  assign \new_[64103]_  = \new_[64102]_  & \new_[64099]_ ;
  assign \new_[64106]_  = ~A203 & ~A202;
  assign \new_[64109]_  = A233 & A232;
  assign \new_[64110]_  = \new_[64109]_  & \new_[64106]_ ;
  assign \new_[64111]_  = \new_[64110]_  & \new_[64103]_ ;
  assign \new_[64114]_  = ~A235 & ~A234;
  assign \new_[64117]_  = A266 & A265;
  assign \new_[64118]_  = \new_[64117]_  & \new_[64114]_ ;
  assign \new_[64121]_  = ~A268 & ~A267;
  assign \new_[64125]_  = A302 & ~A299;
  assign \new_[64126]_  = A298 & \new_[64125]_ ;
  assign \new_[64127]_  = \new_[64126]_  & \new_[64121]_ ;
  assign \new_[64128]_  = \new_[64127]_  & \new_[64118]_ ;
  assign \new_[64131]_  = A167 & A170;
  assign \new_[64134]_  = ~A201 & ~A166;
  assign \new_[64135]_  = \new_[64134]_  & \new_[64131]_ ;
  assign \new_[64138]_  = ~A203 & ~A202;
  assign \new_[64141]_  = A233 & A232;
  assign \new_[64142]_  = \new_[64141]_  & \new_[64138]_ ;
  assign \new_[64143]_  = \new_[64142]_  & \new_[64135]_ ;
  assign \new_[64146]_  = ~A235 & ~A234;
  assign \new_[64149]_  = A266 & A265;
  assign \new_[64150]_  = \new_[64149]_  & \new_[64146]_ ;
  assign \new_[64153]_  = ~A268 & ~A267;
  assign \new_[64157]_  = A302 & A299;
  assign \new_[64158]_  = ~A298 & \new_[64157]_ ;
  assign \new_[64159]_  = \new_[64158]_  & \new_[64153]_ ;
  assign \new_[64160]_  = \new_[64159]_  & \new_[64150]_ ;
  assign \new_[64163]_  = A167 & A170;
  assign \new_[64166]_  = A199 & ~A166;
  assign \new_[64167]_  = \new_[64166]_  & \new_[64163]_ ;
  assign \new_[64170]_  = ~A201 & A200;
  assign \new_[64173]_  = ~A234 & ~A202;
  assign \new_[64174]_  = \new_[64173]_  & \new_[64170]_ ;
  assign \new_[64175]_  = \new_[64174]_  & \new_[64167]_ ;
  assign \new_[64178]_  = ~A236 & ~A235;
  assign \new_[64181]_  = A266 & A265;
  assign \new_[64182]_  = \new_[64181]_  & \new_[64178]_ ;
  assign \new_[64185]_  = ~A268 & ~A267;
  assign \new_[64189]_  = A302 & ~A299;
  assign \new_[64190]_  = A298 & \new_[64189]_ ;
  assign \new_[64191]_  = \new_[64190]_  & \new_[64185]_ ;
  assign \new_[64192]_  = \new_[64191]_  & \new_[64182]_ ;
  assign \new_[64195]_  = A167 & A170;
  assign \new_[64198]_  = A199 & ~A166;
  assign \new_[64199]_  = \new_[64198]_  & \new_[64195]_ ;
  assign \new_[64202]_  = ~A201 & A200;
  assign \new_[64205]_  = ~A234 & ~A202;
  assign \new_[64206]_  = \new_[64205]_  & \new_[64202]_ ;
  assign \new_[64207]_  = \new_[64206]_  & \new_[64199]_ ;
  assign \new_[64210]_  = ~A236 & ~A235;
  assign \new_[64213]_  = A266 & A265;
  assign \new_[64214]_  = \new_[64213]_  & \new_[64210]_ ;
  assign \new_[64217]_  = ~A268 & ~A267;
  assign \new_[64221]_  = A302 & A299;
  assign \new_[64222]_  = ~A298 & \new_[64221]_ ;
  assign \new_[64223]_  = \new_[64222]_  & \new_[64217]_ ;
  assign \new_[64224]_  = \new_[64223]_  & \new_[64214]_ ;
  assign \new_[64227]_  = A167 & A170;
  assign \new_[64230]_  = A199 & ~A166;
  assign \new_[64231]_  = \new_[64230]_  & \new_[64227]_ ;
  assign \new_[64234]_  = ~A201 & A200;
  assign \new_[64237]_  = A232 & ~A202;
  assign \new_[64238]_  = \new_[64237]_  & \new_[64234]_ ;
  assign \new_[64239]_  = \new_[64238]_  & \new_[64231]_ ;
  assign \new_[64242]_  = ~A234 & A233;
  assign \new_[64245]_  = ~A267 & ~A235;
  assign \new_[64246]_  = \new_[64245]_  & \new_[64242]_ ;
  assign \new_[64249]_  = ~A269 & ~A268;
  assign \new_[64253]_  = A302 & ~A299;
  assign \new_[64254]_  = A298 & \new_[64253]_ ;
  assign \new_[64255]_  = \new_[64254]_  & \new_[64249]_ ;
  assign \new_[64256]_  = \new_[64255]_  & \new_[64246]_ ;
  assign \new_[64259]_  = A167 & A170;
  assign \new_[64262]_  = A199 & ~A166;
  assign \new_[64263]_  = \new_[64262]_  & \new_[64259]_ ;
  assign \new_[64266]_  = ~A201 & A200;
  assign \new_[64269]_  = A232 & ~A202;
  assign \new_[64270]_  = \new_[64269]_  & \new_[64266]_ ;
  assign \new_[64271]_  = \new_[64270]_  & \new_[64263]_ ;
  assign \new_[64274]_  = ~A234 & A233;
  assign \new_[64277]_  = ~A267 & ~A235;
  assign \new_[64278]_  = \new_[64277]_  & \new_[64274]_ ;
  assign \new_[64281]_  = ~A269 & ~A268;
  assign \new_[64285]_  = A302 & A299;
  assign \new_[64286]_  = ~A298 & \new_[64285]_ ;
  assign \new_[64287]_  = \new_[64286]_  & \new_[64281]_ ;
  assign \new_[64288]_  = \new_[64287]_  & \new_[64278]_ ;
  assign \new_[64291]_  = A167 & A170;
  assign \new_[64294]_  = A199 & ~A166;
  assign \new_[64295]_  = \new_[64294]_  & \new_[64291]_ ;
  assign \new_[64298]_  = ~A201 & A200;
  assign \new_[64301]_  = A232 & ~A202;
  assign \new_[64302]_  = \new_[64301]_  & \new_[64298]_ ;
  assign \new_[64303]_  = \new_[64302]_  & \new_[64295]_ ;
  assign \new_[64306]_  = ~A234 & A233;
  assign \new_[64309]_  = A265 & ~A235;
  assign \new_[64310]_  = \new_[64309]_  & \new_[64306]_ ;
  assign \new_[64313]_  = ~A267 & A266;
  assign \new_[64317]_  = A300 & A299;
  assign \new_[64318]_  = ~A268 & \new_[64317]_ ;
  assign \new_[64319]_  = \new_[64318]_  & \new_[64313]_ ;
  assign \new_[64320]_  = \new_[64319]_  & \new_[64310]_ ;
  assign \new_[64323]_  = A167 & A170;
  assign \new_[64326]_  = A199 & ~A166;
  assign \new_[64327]_  = \new_[64326]_  & \new_[64323]_ ;
  assign \new_[64330]_  = ~A201 & A200;
  assign \new_[64333]_  = A232 & ~A202;
  assign \new_[64334]_  = \new_[64333]_  & \new_[64330]_ ;
  assign \new_[64335]_  = \new_[64334]_  & \new_[64327]_ ;
  assign \new_[64338]_  = ~A234 & A233;
  assign \new_[64341]_  = A265 & ~A235;
  assign \new_[64342]_  = \new_[64341]_  & \new_[64338]_ ;
  assign \new_[64345]_  = ~A267 & A266;
  assign \new_[64349]_  = A300 & A298;
  assign \new_[64350]_  = ~A268 & \new_[64349]_ ;
  assign \new_[64351]_  = \new_[64350]_  & \new_[64345]_ ;
  assign \new_[64352]_  = \new_[64351]_  & \new_[64342]_ ;
  assign \new_[64355]_  = A167 & A170;
  assign \new_[64358]_  = A199 & ~A166;
  assign \new_[64359]_  = \new_[64358]_  & \new_[64355]_ ;
  assign \new_[64362]_  = ~A201 & A200;
  assign \new_[64365]_  = A232 & ~A202;
  assign \new_[64366]_  = \new_[64365]_  & \new_[64362]_ ;
  assign \new_[64367]_  = \new_[64366]_  & \new_[64359]_ ;
  assign \new_[64370]_  = ~A234 & A233;
  assign \new_[64373]_  = ~A265 & ~A235;
  assign \new_[64374]_  = \new_[64373]_  & \new_[64370]_ ;
  assign \new_[64377]_  = ~A268 & ~A266;
  assign \new_[64381]_  = A302 & ~A299;
  assign \new_[64382]_  = A298 & \new_[64381]_ ;
  assign \new_[64383]_  = \new_[64382]_  & \new_[64377]_ ;
  assign \new_[64384]_  = \new_[64383]_  & \new_[64374]_ ;
  assign \new_[64387]_  = A167 & A170;
  assign \new_[64390]_  = A199 & ~A166;
  assign \new_[64391]_  = \new_[64390]_  & \new_[64387]_ ;
  assign \new_[64394]_  = ~A201 & A200;
  assign \new_[64397]_  = A232 & ~A202;
  assign \new_[64398]_  = \new_[64397]_  & \new_[64394]_ ;
  assign \new_[64399]_  = \new_[64398]_  & \new_[64391]_ ;
  assign \new_[64402]_  = ~A234 & A233;
  assign \new_[64405]_  = ~A265 & ~A235;
  assign \new_[64406]_  = \new_[64405]_  & \new_[64402]_ ;
  assign \new_[64409]_  = ~A268 & ~A266;
  assign \new_[64413]_  = A302 & A299;
  assign \new_[64414]_  = ~A298 & \new_[64413]_ ;
  assign \new_[64415]_  = \new_[64414]_  & \new_[64409]_ ;
  assign \new_[64416]_  = \new_[64415]_  & \new_[64406]_ ;
  assign \new_[64419]_  = A167 & A170;
  assign \new_[64422]_  = A199 & ~A166;
  assign \new_[64423]_  = \new_[64422]_  & \new_[64419]_ ;
  assign \new_[64426]_  = ~A201 & A200;
  assign \new_[64429]_  = ~A232 & ~A202;
  assign \new_[64430]_  = \new_[64429]_  & \new_[64426]_ ;
  assign \new_[64431]_  = \new_[64430]_  & \new_[64423]_ ;
  assign \new_[64434]_  = ~A235 & ~A233;
  assign \new_[64437]_  = A266 & A265;
  assign \new_[64438]_  = \new_[64437]_  & \new_[64434]_ ;
  assign \new_[64441]_  = ~A268 & ~A267;
  assign \new_[64445]_  = A302 & ~A299;
  assign \new_[64446]_  = A298 & \new_[64445]_ ;
  assign \new_[64447]_  = \new_[64446]_  & \new_[64441]_ ;
  assign \new_[64448]_  = \new_[64447]_  & \new_[64438]_ ;
  assign \new_[64451]_  = A167 & A170;
  assign \new_[64454]_  = A199 & ~A166;
  assign \new_[64455]_  = \new_[64454]_  & \new_[64451]_ ;
  assign \new_[64458]_  = ~A201 & A200;
  assign \new_[64461]_  = ~A232 & ~A202;
  assign \new_[64462]_  = \new_[64461]_  & \new_[64458]_ ;
  assign \new_[64463]_  = \new_[64462]_  & \new_[64455]_ ;
  assign \new_[64466]_  = ~A235 & ~A233;
  assign \new_[64469]_  = A266 & A265;
  assign \new_[64470]_  = \new_[64469]_  & \new_[64466]_ ;
  assign \new_[64473]_  = ~A268 & ~A267;
  assign \new_[64477]_  = A302 & A299;
  assign \new_[64478]_  = ~A298 & \new_[64477]_ ;
  assign \new_[64479]_  = \new_[64478]_  & \new_[64473]_ ;
  assign \new_[64480]_  = \new_[64479]_  & \new_[64470]_ ;
  assign \new_[64483]_  = A167 & A170;
  assign \new_[64486]_  = ~A199 & ~A166;
  assign \new_[64487]_  = \new_[64486]_  & \new_[64483]_ ;
  assign \new_[64490]_  = ~A202 & ~A200;
  assign \new_[64493]_  = A233 & A232;
  assign \new_[64494]_  = \new_[64493]_  & \new_[64490]_ ;
  assign \new_[64495]_  = \new_[64494]_  & \new_[64487]_ ;
  assign \new_[64498]_  = ~A235 & ~A234;
  assign \new_[64501]_  = A266 & A265;
  assign \new_[64502]_  = \new_[64501]_  & \new_[64498]_ ;
  assign \new_[64505]_  = ~A268 & ~A267;
  assign \new_[64509]_  = A302 & ~A299;
  assign \new_[64510]_  = A298 & \new_[64509]_ ;
  assign \new_[64511]_  = \new_[64510]_  & \new_[64505]_ ;
  assign \new_[64512]_  = \new_[64511]_  & \new_[64502]_ ;
  assign \new_[64515]_  = A167 & A170;
  assign \new_[64518]_  = ~A199 & ~A166;
  assign \new_[64519]_  = \new_[64518]_  & \new_[64515]_ ;
  assign \new_[64522]_  = ~A202 & ~A200;
  assign \new_[64525]_  = A233 & A232;
  assign \new_[64526]_  = \new_[64525]_  & \new_[64522]_ ;
  assign \new_[64527]_  = \new_[64526]_  & \new_[64519]_ ;
  assign \new_[64530]_  = ~A235 & ~A234;
  assign \new_[64533]_  = A266 & A265;
  assign \new_[64534]_  = \new_[64533]_  & \new_[64530]_ ;
  assign \new_[64537]_  = ~A268 & ~A267;
  assign \new_[64541]_  = A302 & A299;
  assign \new_[64542]_  = ~A298 & \new_[64541]_ ;
  assign \new_[64543]_  = \new_[64542]_  & \new_[64537]_ ;
  assign \new_[64544]_  = \new_[64543]_  & \new_[64534]_ ;
  assign \new_[64547]_  = ~A167 & A170;
  assign \new_[64550]_  = ~A201 & A166;
  assign \new_[64551]_  = \new_[64550]_  & \new_[64547]_ ;
  assign \new_[64554]_  = ~A203 & ~A202;
  assign \new_[64557]_  = A233 & A232;
  assign \new_[64558]_  = \new_[64557]_  & \new_[64554]_ ;
  assign \new_[64559]_  = \new_[64558]_  & \new_[64551]_ ;
  assign \new_[64562]_  = ~A235 & ~A234;
  assign \new_[64565]_  = A266 & A265;
  assign \new_[64566]_  = \new_[64565]_  & \new_[64562]_ ;
  assign \new_[64569]_  = ~A268 & ~A267;
  assign \new_[64573]_  = A302 & ~A299;
  assign \new_[64574]_  = A298 & \new_[64573]_ ;
  assign \new_[64575]_  = \new_[64574]_  & \new_[64569]_ ;
  assign \new_[64576]_  = \new_[64575]_  & \new_[64566]_ ;
  assign \new_[64579]_  = ~A167 & A170;
  assign \new_[64582]_  = ~A201 & A166;
  assign \new_[64583]_  = \new_[64582]_  & \new_[64579]_ ;
  assign \new_[64586]_  = ~A203 & ~A202;
  assign \new_[64589]_  = A233 & A232;
  assign \new_[64590]_  = \new_[64589]_  & \new_[64586]_ ;
  assign \new_[64591]_  = \new_[64590]_  & \new_[64583]_ ;
  assign \new_[64594]_  = ~A235 & ~A234;
  assign \new_[64597]_  = A266 & A265;
  assign \new_[64598]_  = \new_[64597]_  & \new_[64594]_ ;
  assign \new_[64601]_  = ~A268 & ~A267;
  assign \new_[64605]_  = A302 & A299;
  assign \new_[64606]_  = ~A298 & \new_[64605]_ ;
  assign \new_[64607]_  = \new_[64606]_  & \new_[64601]_ ;
  assign \new_[64608]_  = \new_[64607]_  & \new_[64598]_ ;
  assign \new_[64611]_  = ~A167 & A170;
  assign \new_[64614]_  = A199 & A166;
  assign \new_[64615]_  = \new_[64614]_  & \new_[64611]_ ;
  assign \new_[64618]_  = ~A201 & A200;
  assign \new_[64621]_  = ~A234 & ~A202;
  assign \new_[64622]_  = \new_[64621]_  & \new_[64618]_ ;
  assign \new_[64623]_  = \new_[64622]_  & \new_[64615]_ ;
  assign \new_[64626]_  = ~A236 & ~A235;
  assign \new_[64629]_  = A266 & A265;
  assign \new_[64630]_  = \new_[64629]_  & \new_[64626]_ ;
  assign \new_[64633]_  = ~A268 & ~A267;
  assign \new_[64637]_  = A302 & ~A299;
  assign \new_[64638]_  = A298 & \new_[64637]_ ;
  assign \new_[64639]_  = \new_[64638]_  & \new_[64633]_ ;
  assign \new_[64640]_  = \new_[64639]_  & \new_[64630]_ ;
  assign \new_[64643]_  = ~A167 & A170;
  assign \new_[64646]_  = A199 & A166;
  assign \new_[64647]_  = \new_[64646]_  & \new_[64643]_ ;
  assign \new_[64650]_  = ~A201 & A200;
  assign \new_[64653]_  = ~A234 & ~A202;
  assign \new_[64654]_  = \new_[64653]_  & \new_[64650]_ ;
  assign \new_[64655]_  = \new_[64654]_  & \new_[64647]_ ;
  assign \new_[64658]_  = ~A236 & ~A235;
  assign \new_[64661]_  = A266 & A265;
  assign \new_[64662]_  = \new_[64661]_  & \new_[64658]_ ;
  assign \new_[64665]_  = ~A268 & ~A267;
  assign \new_[64669]_  = A302 & A299;
  assign \new_[64670]_  = ~A298 & \new_[64669]_ ;
  assign \new_[64671]_  = \new_[64670]_  & \new_[64665]_ ;
  assign \new_[64672]_  = \new_[64671]_  & \new_[64662]_ ;
  assign \new_[64675]_  = ~A167 & A170;
  assign \new_[64678]_  = A199 & A166;
  assign \new_[64679]_  = \new_[64678]_  & \new_[64675]_ ;
  assign \new_[64682]_  = ~A201 & A200;
  assign \new_[64685]_  = A232 & ~A202;
  assign \new_[64686]_  = \new_[64685]_  & \new_[64682]_ ;
  assign \new_[64687]_  = \new_[64686]_  & \new_[64679]_ ;
  assign \new_[64690]_  = ~A234 & A233;
  assign \new_[64693]_  = ~A267 & ~A235;
  assign \new_[64694]_  = \new_[64693]_  & \new_[64690]_ ;
  assign \new_[64697]_  = ~A269 & ~A268;
  assign \new_[64701]_  = A302 & ~A299;
  assign \new_[64702]_  = A298 & \new_[64701]_ ;
  assign \new_[64703]_  = \new_[64702]_  & \new_[64697]_ ;
  assign \new_[64704]_  = \new_[64703]_  & \new_[64694]_ ;
  assign \new_[64707]_  = ~A167 & A170;
  assign \new_[64710]_  = A199 & A166;
  assign \new_[64711]_  = \new_[64710]_  & \new_[64707]_ ;
  assign \new_[64714]_  = ~A201 & A200;
  assign \new_[64717]_  = A232 & ~A202;
  assign \new_[64718]_  = \new_[64717]_  & \new_[64714]_ ;
  assign \new_[64719]_  = \new_[64718]_  & \new_[64711]_ ;
  assign \new_[64722]_  = ~A234 & A233;
  assign \new_[64725]_  = ~A267 & ~A235;
  assign \new_[64726]_  = \new_[64725]_  & \new_[64722]_ ;
  assign \new_[64729]_  = ~A269 & ~A268;
  assign \new_[64733]_  = A302 & A299;
  assign \new_[64734]_  = ~A298 & \new_[64733]_ ;
  assign \new_[64735]_  = \new_[64734]_  & \new_[64729]_ ;
  assign \new_[64736]_  = \new_[64735]_  & \new_[64726]_ ;
  assign \new_[64739]_  = ~A167 & A170;
  assign \new_[64742]_  = A199 & A166;
  assign \new_[64743]_  = \new_[64742]_  & \new_[64739]_ ;
  assign \new_[64746]_  = ~A201 & A200;
  assign \new_[64749]_  = A232 & ~A202;
  assign \new_[64750]_  = \new_[64749]_  & \new_[64746]_ ;
  assign \new_[64751]_  = \new_[64750]_  & \new_[64743]_ ;
  assign \new_[64754]_  = ~A234 & A233;
  assign \new_[64757]_  = A265 & ~A235;
  assign \new_[64758]_  = \new_[64757]_  & \new_[64754]_ ;
  assign \new_[64761]_  = ~A267 & A266;
  assign \new_[64765]_  = A300 & A299;
  assign \new_[64766]_  = ~A268 & \new_[64765]_ ;
  assign \new_[64767]_  = \new_[64766]_  & \new_[64761]_ ;
  assign \new_[64768]_  = \new_[64767]_  & \new_[64758]_ ;
  assign \new_[64771]_  = ~A167 & A170;
  assign \new_[64774]_  = A199 & A166;
  assign \new_[64775]_  = \new_[64774]_  & \new_[64771]_ ;
  assign \new_[64778]_  = ~A201 & A200;
  assign \new_[64781]_  = A232 & ~A202;
  assign \new_[64782]_  = \new_[64781]_  & \new_[64778]_ ;
  assign \new_[64783]_  = \new_[64782]_  & \new_[64775]_ ;
  assign \new_[64786]_  = ~A234 & A233;
  assign \new_[64789]_  = A265 & ~A235;
  assign \new_[64790]_  = \new_[64789]_  & \new_[64786]_ ;
  assign \new_[64793]_  = ~A267 & A266;
  assign \new_[64797]_  = A300 & A298;
  assign \new_[64798]_  = ~A268 & \new_[64797]_ ;
  assign \new_[64799]_  = \new_[64798]_  & \new_[64793]_ ;
  assign \new_[64800]_  = \new_[64799]_  & \new_[64790]_ ;
  assign \new_[64803]_  = ~A167 & A170;
  assign \new_[64806]_  = A199 & A166;
  assign \new_[64807]_  = \new_[64806]_  & \new_[64803]_ ;
  assign \new_[64810]_  = ~A201 & A200;
  assign \new_[64813]_  = A232 & ~A202;
  assign \new_[64814]_  = \new_[64813]_  & \new_[64810]_ ;
  assign \new_[64815]_  = \new_[64814]_  & \new_[64807]_ ;
  assign \new_[64818]_  = ~A234 & A233;
  assign \new_[64821]_  = ~A265 & ~A235;
  assign \new_[64822]_  = \new_[64821]_  & \new_[64818]_ ;
  assign \new_[64825]_  = ~A268 & ~A266;
  assign \new_[64829]_  = A302 & ~A299;
  assign \new_[64830]_  = A298 & \new_[64829]_ ;
  assign \new_[64831]_  = \new_[64830]_  & \new_[64825]_ ;
  assign \new_[64832]_  = \new_[64831]_  & \new_[64822]_ ;
  assign \new_[64835]_  = ~A167 & A170;
  assign \new_[64838]_  = A199 & A166;
  assign \new_[64839]_  = \new_[64838]_  & \new_[64835]_ ;
  assign \new_[64842]_  = ~A201 & A200;
  assign \new_[64845]_  = A232 & ~A202;
  assign \new_[64846]_  = \new_[64845]_  & \new_[64842]_ ;
  assign \new_[64847]_  = \new_[64846]_  & \new_[64839]_ ;
  assign \new_[64850]_  = ~A234 & A233;
  assign \new_[64853]_  = ~A265 & ~A235;
  assign \new_[64854]_  = \new_[64853]_  & \new_[64850]_ ;
  assign \new_[64857]_  = ~A268 & ~A266;
  assign \new_[64861]_  = A302 & A299;
  assign \new_[64862]_  = ~A298 & \new_[64861]_ ;
  assign \new_[64863]_  = \new_[64862]_  & \new_[64857]_ ;
  assign \new_[64864]_  = \new_[64863]_  & \new_[64854]_ ;
  assign \new_[64867]_  = ~A167 & A170;
  assign \new_[64870]_  = A199 & A166;
  assign \new_[64871]_  = \new_[64870]_  & \new_[64867]_ ;
  assign \new_[64874]_  = ~A201 & A200;
  assign \new_[64877]_  = ~A232 & ~A202;
  assign \new_[64878]_  = \new_[64877]_  & \new_[64874]_ ;
  assign \new_[64879]_  = \new_[64878]_  & \new_[64871]_ ;
  assign \new_[64882]_  = ~A235 & ~A233;
  assign \new_[64885]_  = A266 & A265;
  assign \new_[64886]_  = \new_[64885]_  & \new_[64882]_ ;
  assign \new_[64889]_  = ~A268 & ~A267;
  assign \new_[64893]_  = A302 & ~A299;
  assign \new_[64894]_  = A298 & \new_[64893]_ ;
  assign \new_[64895]_  = \new_[64894]_  & \new_[64889]_ ;
  assign \new_[64896]_  = \new_[64895]_  & \new_[64886]_ ;
  assign \new_[64899]_  = ~A167 & A170;
  assign \new_[64902]_  = A199 & A166;
  assign \new_[64903]_  = \new_[64902]_  & \new_[64899]_ ;
  assign \new_[64906]_  = ~A201 & A200;
  assign \new_[64909]_  = ~A232 & ~A202;
  assign \new_[64910]_  = \new_[64909]_  & \new_[64906]_ ;
  assign \new_[64911]_  = \new_[64910]_  & \new_[64903]_ ;
  assign \new_[64914]_  = ~A235 & ~A233;
  assign \new_[64917]_  = A266 & A265;
  assign \new_[64918]_  = \new_[64917]_  & \new_[64914]_ ;
  assign \new_[64921]_  = ~A268 & ~A267;
  assign \new_[64925]_  = A302 & A299;
  assign \new_[64926]_  = ~A298 & \new_[64925]_ ;
  assign \new_[64927]_  = \new_[64926]_  & \new_[64921]_ ;
  assign \new_[64928]_  = \new_[64927]_  & \new_[64918]_ ;
  assign \new_[64931]_  = ~A167 & A170;
  assign \new_[64934]_  = ~A199 & A166;
  assign \new_[64935]_  = \new_[64934]_  & \new_[64931]_ ;
  assign \new_[64938]_  = ~A202 & ~A200;
  assign \new_[64941]_  = A233 & A232;
  assign \new_[64942]_  = \new_[64941]_  & \new_[64938]_ ;
  assign \new_[64943]_  = \new_[64942]_  & \new_[64935]_ ;
  assign \new_[64946]_  = ~A235 & ~A234;
  assign \new_[64949]_  = A266 & A265;
  assign \new_[64950]_  = \new_[64949]_  & \new_[64946]_ ;
  assign \new_[64953]_  = ~A268 & ~A267;
  assign \new_[64957]_  = A302 & ~A299;
  assign \new_[64958]_  = A298 & \new_[64957]_ ;
  assign \new_[64959]_  = \new_[64958]_  & \new_[64953]_ ;
  assign \new_[64960]_  = \new_[64959]_  & \new_[64950]_ ;
  assign \new_[64963]_  = ~A167 & A170;
  assign \new_[64966]_  = ~A199 & A166;
  assign \new_[64967]_  = \new_[64966]_  & \new_[64963]_ ;
  assign \new_[64970]_  = ~A202 & ~A200;
  assign \new_[64973]_  = A233 & A232;
  assign \new_[64974]_  = \new_[64973]_  & \new_[64970]_ ;
  assign \new_[64975]_  = \new_[64974]_  & \new_[64967]_ ;
  assign \new_[64978]_  = ~A235 & ~A234;
  assign \new_[64981]_  = A266 & A265;
  assign \new_[64982]_  = \new_[64981]_  & \new_[64978]_ ;
  assign \new_[64985]_  = ~A268 & ~A267;
  assign \new_[64989]_  = A302 & A299;
  assign \new_[64990]_  = ~A298 & \new_[64989]_ ;
  assign \new_[64991]_  = \new_[64990]_  & \new_[64985]_ ;
  assign \new_[64992]_  = \new_[64991]_  & \new_[64982]_ ;
  assign \new_[64995]_  = ~A167 & ~A169;
  assign \new_[64998]_  = ~A199 & ~A166;
  assign \new_[64999]_  = \new_[64998]_  & \new_[64995]_ ;
  assign \new_[65002]_  = A203 & A200;
  assign \new_[65005]_  = A233 & A232;
  assign \new_[65006]_  = \new_[65005]_  & \new_[65002]_ ;
  assign \new_[65007]_  = \new_[65006]_  & \new_[64999]_ ;
  assign \new_[65010]_  = ~A235 & ~A234;
  assign \new_[65013]_  = A266 & A265;
  assign \new_[65014]_  = \new_[65013]_  & \new_[65010]_ ;
  assign \new_[65017]_  = ~A268 & ~A267;
  assign \new_[65021]_  = A302 & ~A299;
  assign \new_[65022]_  = A298 & \new_[65021]_ ;
  assign \new_[65023]_  = \new_[65022]_  & \new_[65017]_ ;
  assign \new_[65024]_  = \new_[65023]_  & \new_[65014]_ ;
  assign \new_[65027]_  = ~A167 & ~A169;
  assign \new_[65030]_  = ~A199 & ~A166;
  assign \new_[65031]_  = \new_[65030]_  & \new_[65027]_ ;
  assign \new_[65034]_  = A203 & A200;
  assign \new_[65037]_  = A233 & A232;
  assign \new_[65038]_  = \new_[65037]_  & \new_[65034]_ ;
  assign \new_[65039]_  = \new_[65038]_  & \new_[65031]_ ;
  assign \new_[65042]_  = ~A235 & ~A234;
  assign \new_[65045]_  = A266 & A265;
  assign \new_[65046]_  = \new_[65045]_  & \new_[65042]_ ;
  assign \new_[65049]_  = ~A268 & ~A267;
  assign \new_[65053]_  = A302 & A299;
  assign \new_[65054]_  = ~A298 & \new_[65053]_ ;
  assign \new_[65055]_  = \new_[65054]_  & \new_[65049]_ ;
  assign \new_[65056]_  = \new_[65055]_  & \new_[65046]_ ;
  assign \new_[65059]_  = ~A167 & ~A169;
  assign \new_[65062]_  = A199 & ~A166;
  assign \new_[65063]_  = \new_[65062]_  & \new_[65059]_ ;
  assign \new_[65066]_  = A203 & ~A200;
  assign \new_[65069]_  = A233 & A232;
  assign \new_[65070]_  = \new_[65069]_  & \new_[65066]_ ;
  assign \new_[65071]_  = \new_[65070]_  & \new_[65063]_ ;
  assign \new_[65074]_  = ~A235 & ~A234;
  assign \new_[65077]_  = A266 & A265;
  assign \new_[65078]_  = \new_[65077]_  & \new_[65074]_ ;
  assign \new_[65081]_  = ~A268 & ~A267;
  assign \new_[65085]_  = A302 & ~A299;
  assign \new_[65086]_  = A298 & \new_[65085]_ ;
  assign \new_[65087]_  = \new_[65086]_  & \new_[65081]_ ;
  assign \new_[65088]_  = \new_[65087]_  & \new_[65078]_ ;
  assign \new_[65091]_  = ~A167 & ~A169;
  assign \new_[65094]_  = A199 & ~A166;
  assign \new_[65095]_  = \new_[65094]_  & \new_[65091]_ ;
  assign \new_[65098]_  = A203 & ~A200;
  assign \new_[65101]_  = A233 & A232;
  assign \new_[65102]_  = \new_[65101]_  & \new_[65098]_ ;
  assign \new_[65103]_  = \new_[65102]_  & \new_[65095]_ ;
  assign \new_[65106]_  = ~A235 & ~A234;
  assign \new_[65109]_  = A266 & A265;
  assign \new_[65110]_  = \new_[65109]_  & \new_[65106]_ ;
  assign \new_[65113]_  = ~A268 & ~A267;
  assign \new_[65117]_  = A302 & A299;
  assign \new_[65118]_  = ~A298 & \new_[65117]_ ;
  assign \new_[65119]_  = \new_[65118]_  & \new_[65113]_ ;
  assign \new_[65120]_  = \new_[65119]_  & \new_[65110]_ ;
  assign \new_[65123]_  = ~A168 & ~A169;
  assign \new_[65126]_  = A166 & A167;
  assign \new_[65127]_  = \new_[65126]_  & \new_[65123]_ ;
  assign \new_[65130]_  = A201 & A199;
  assign \new_[65133]_  = A233 & A232;
  assign \new_[65134]_  = \new_[65133]_  & \new_[65130]_ ;
  assign \new_[65135]_  = \new_[65134]_  & \new_[65127]_ ;
  assign \new_[65138]_  = ~A235 & ~A234;
  assign \new_[65141]_  = A266 & A265;
  assign \new_[65142]_  = \new_[65141]_  & \new_[65138]_ ;
  assign \new_[65145]_  = ~A268 & ~A267;
  assign \new_[65149]_  = A302 & ~A299;
  assign \new_[65150]_  = A298 & \new_[65149]_ ;
  assign \new_[65151]_  = \new_[65150]_  & \new_[65145]_ ;
  assign \new_[65152]_  = \new_[65151]_  & \new_[65142]_ ;
  assign \new_[65155]_  = ~A168 & ~A169;
  assign \new_[65158]_  = A166 & A167;
  assign \new_[65159]_  = \new_[65158]_  & \new_[65155]_ ;
  assign \new_[65162]_  = A201 & A199;
  assign \new_[65165]_  = A233 & A232;
  assign \new_[65166]_  = \new_[65165]_  & \new_[65162]_ ;
  assign \new_[65167]_  = \new_[65166]_  & \new_[65159]_ ;
  assign \new_[65170]_  = ~A235 & ~A234;
  assign \new_[65173]_  = A266 & A265;
  assign \new_[65174]_  = \new_[65173]_  & \new_[65170]_ ;
  assign \new_[65177]_  = ~A268 & ~A267;
  assign \new_[65181]_  = A302 & A299;
  assign \new_[65182]_  = ~A298 & \new_[65181]_ ;
  assign \new_[65183]_  = \new_[65182]_  & \new_[65177]_ ;
  assign \new_[65184]_  = \new_[65183]_  & \new_[65174]_ ;
  assign \new_[65187]_  = ~A168 & ~A169;
  assign \new_[65190]_  = A166 & A167;
  assign \new_[65191]_  = \new_[65190]_  & \new_[65187]_ ;
  assign \new_[65194]_  = A201 & A200;
  assign \new_[65197]_  = A233 & A232;
  assign \new_[65198]_  = \new_[65197]_  & \new_[65194]_ ;
  assign \new_[65199]_  = \new_[65198]_  & \new_[65191]_ ;
  assign \new_[65202]_  = ~A235 & ~A234;
  assign \new_[65205]_  = A266 & A265;
  assign \new_[65206]_  = \new_[65205]_  & \new_[65202]_ ;
  assign \new_[65209]_  = ~A268 & ~A267;
  assign \new_[65213]_  = A302 & ~A299;
  assign \new_[65214]_  = A298 & \new_[65213]_ ;
  assign \new_[65215]_  = \new_[65214]_  & \new_[65209]_ ;
  assign \new_[65216]_  = \new_[65215]_  & \new_[65206]_ ;
  assign \new_[65219]_  = ~A168 & ~A169;
  assign \new_[65222]_  = A166 & A167;
  assign \new_[65223]_  = \new_[65222]_  & \new_[65219]_ ;
  assign \new_[65226]_  = A201 & A200;
  assign \new_[65229]_  = A233 & A232;
  assign \new_[65230]_  = \new_[65229]_  & \new_[65226]_ ;
  assign \new_[65231]_  = \new_[65230]_  & \new_[65223]_ ;
  assign \new_[65234]_  = ~A235 & ~A234;
  assign \new_[65237]_  = A266 & A265;
  assign \new_[65238]_  = \new_[65237]_  & \new_[65234]_ ;
  assign \new_[65241]_  = ~A268 & ~A267;
  assign \new_[65245]_  = A302 & A299;
  assign \new_[65246]_  = ~A298 & \new_[65245]_ ;
  assign \new_[65247]_  = \new_[65246]_  & \new_[65241]_ ;
  assign \new_[65248]_  = \new_[65247]_  & \new_[65238]_ ;
  assign \new_[65251]_  = ~A168 & ~A169;
  assign \new_[65254]_  = A166 & A167;
  assign \new_[65255]_  = \new_[65254]_  & \new_[65251]_ ;
  assign \new_[65258]_  = A200 & ~A199;
  assign \new_[65261]_  = ~A234 & A203;
  assign \new_[65262]_  = \new_[65261]_  & \new_[65258]_ ;
  assign \new_[65263]_  = \new_[65262]_  & \new_[65255]_ ;
  assign \new_[65266]_  = ~A236 & ~A235;
  assign \new_[65269]_  = A266 & A265;
  assign \new_[65270]_  = \new_[65269]_  & \new_[65266]_ ;
  assign \new_[65273]_  = ~A268 & ~A267;
  assign \new_[65277]_  = A302 & ~A299;
  assign \new_[65278]_  = A298 & \new_[65277]_ ;
  assign \new_[65279]_  = \new_[65278]_  & \new_[65273]_ ;
  assign \new_[65280]_  = \new_[65279]_  & \new_[65270]_ ;
  assign \new_[65283]_  = ~A168 & ~A169;
  assign \new_[65286]_  = A166 & A167;
  assign \new_[65287]_  = \new_[65286]_  & \new_[65283]_ ;
  assign \new_[65290]_  = A200 & ~A199;
  assign \new_[65293]_  = ~A234 & A203;
  assign \new_[65294]_  = \new_[65293]_  & \new_[65290]_ ;
  assign \new_[65295]_  = \new_[65294]_  & \new_[65287]_ ;
  assign \new_[65298]_  = ~A236 & ~A235;
  assign \new_[65301]_  = A266 & A265;
  assign \new_[65302]_  = \new_[65301]_  & \new_[65298]_ ;
  assign \new_[65305]_  = ~A268 & ~A267;
  assign \new_[65309]_  = A302 & A299;
  assign \new_[65310]_  = ~A298 & \new_[65309]_ ;
  assign \new_[65311]_  = \new_[65310]_  & \new_[65305]_ ;
  assign \new_[65312]_  = \new_[65311]_  & \new_[65302]_ ;
  assign \new_[65315]_  = ~A168 & ~A169;
  assign \new_[65318]_  = A166 & A167;
  assign \new_[65319]_  = \new_[65318]_  & \new_[65315]_ ;
  assign \new_[65322]_  = A200 & ~A199;
  assign \new_[65325]_  = A232 & A203;
  assign \new_[65326]_  = \new_[65325]_  & \new_[65322]_ ;
  assign \new_[65327]_  = \new_[65326]_  & \new_[65319]_ ;
  assign \new_[65330]_  = ~A234 & A233;
  assign \new_[65333]_  = ~A267 & ~A235;
  assign \new_[65334]_  = \new_[65333]_  & \new_[65330]_ ;
  assign \new_[65337]_  = ~A269 & ~A268;
  assign \new_[65341]_  = A302 & ~A299;
  assign \new_[65342]_  = A298 & \new_[65341]_ ;
  assign \new_[65343]_  = \new_[65342]_  & \new_[65337]_ ;
  assign \new_[65344]_  = \new_[65343]_  & \new_[65334]_ ;
  assign \new_[65347]_  = ~A168 & ~A169;
  assign \new_[65350]_  = A166 & A167;
  assign \new_[65351]_  = \new_[65350]_  & \new_[65347]_ ;
  assign \new_[65354]_  = A200 & ~A199;
  assign \new_[65357]_  = A232 & A203;
  assign \new_[65358]_  = \new_[65357]_  & \new_[65354]_ ;
  assign \new_[65359]_  = \new_[65358]_  & \new_[65351]_ ;
  assign \new_[65362]_  = ~A234 & A233;
  assign \new_[65365]_  = ~A267 & ~A235;
  assign \new_[65366]_  = \new_[65365]_  & \new_[65362]_ ;
  assign \new_[65369]_  = ~A269 & ~A268;
  assign \new_[65373]_  = A302 & A299;
  assign \new_[65374]_  = ~A298 & \new_[65373]_ ;
  assign \new_[65375]_  = \new_[65374]_  & \new_[65369]_ ;
  assign \new_[65376]_  = \new_[65375]_  & \new_[65366]_ ;
  assign \new_[65379]_  = ~A168 & ~A169;
  assign \new_[65382]_  = A166 & A167;
  assign \new_[65383]_  = \new_[65382]_  & \new_[65379]_ ;
  assign \new_[65386]_  = A200 & ~A199;
  assign \new_[65389]_  = A232 & A203;
  assign \new_[65390]_  = \new_[65389]_  & \new_[65386]_ ;
  assign \new_[65391]_  = \new_[65390]_  & \new_[65383]_ ;
  assign \new_[65394]_  = ~A234 & A233;
  assign \new_[65397]_  = A265 & ~A235;
  assign \new_[65398]_  = \new_[65397]_  & \new_[65394]_ ;
  assign \new_[65401]_  = ~A267 & A266;
  assign \new_[65405]_  = A300 & A299;
  assign \new_[65406]_  = ~A268 & \new_[65405]_ ;
  assign \new_[65407]_  = \new_[65406]_  & \new_[65401]_ ;
  assign \new_[65408]_  = \new_[65407]_  & \new_[65398]_ ;
  assign \new_[65411]_  = ~A168 & ~A169;
  assign \new_[65414]_  = A166 & A167;
  assign \new_[65415]_  = \new_[65414]_  & \new_[65411]_ ;
  assign \new_[65418]_  = A200 & ~A199;
  assign \new_[65421]_  = A232 & A203;
  assign \new_[65422]_  = \new_[65421]_  & \new_[65418]_ ;
  assign \new_[65423]_  = \new_[65422]_  & \new_[65415]_ ;
  assign \new_[65426]_  = ~A234 & A233;
  assign \new_[65429]_  = A265 & ~A235;
  assign \new_[65430]_  = \new_[65429]_  & \new_[65426]_ ;
  assign \new_[65433]_  = ~A267 & A266;
  assign \new_[65437]_  = A300 & A298;
  assign \new_[65438]_  = ~A268 & \new_[65437]_ ;
  assign \new_[65439]_  = \new_[65438]_  & \new_[65433]_ ;
  assign \new_[65440]_  = \new_[65439]_  & \new_[65430]_ ;
  assign \new_[65443]_  = ~A168 & ~A169;
  assign \new_[65446]_  = A166 & A167;
  assign \new_[65447]_  = \new_[65446]_  & \new_[65443]_ ;
  assign \new_[65450]_  = A200 & ~A199;
  assign \new_[65453]_  = A232 & A203;
  assign \new_[65454]_  = \new_[65453]_  & \new_[65450]_ ;
  assign \new_[65455]_  = \new_[65454]_  & \new_[65447]_ ;
  assign \new_[65458]_  = ~A234 & A233;
  assign \new_[65461]_  = ~A265 & ~A235;
  assign \new_[65462]_  = \new_[65461]_  & \new_[65458]_ ;
  assign \new_[65465]_  = ~A268 & ~A266;
  assign \new_[65469]_  = A302 & ~A299;
  assign \new_[65470]_  = A298 & \new_[65469]_ ;
  assign \new_[65471]_  = \new_[65470]_  & \new_[65465]_ ;
  assign \new_[65472]_  = \new_[65471]_  & \new_[65462]_ ;
  assign \new_[65475]_  = ~A168 & ~A169;
  assign \new_[65478]_  = A166 & A167;
  assign \new_[65479]_  = \new_[65478]_  & \new_[65475]_ ;
  assign \new_[65482]_  = A200 & ~A199;
  assign \new_[65485]_  = A232 & A203;
  assign \new_[65486]_  = \new_[65485]_  & \new_[65482]_ ;
  assign \new_[65487]_  = \new_[65486]_  & \new_[65479]_ ;
  assign \new_[65490]_  = ~A234 & A233;
  assign \new_[65493]_  = ~A265 & ~A235;
  assign \new_[65494]_  = \new_[65493]_  & \new_[65490]_ ;
  assign \new_[65497]_  = ~A268 & ~A266;
  assign \new_[65501]_  = A302 & A299;
  assign \new_[65502]_  = ~A298 & \new_[65501]_ ;
  assign \new_[65503]_  = \new_[65502]_  & \new_[65497]_ ;
  assign \new_[65504]_  = \new_[65503]_  & \new_[65494]_ ;
  assign \new_[65507]_  = ~A168 & ~A169;
  assign \new_[65510]_  = A166 & A167;
  assign \new_[65511]_  = \new_[65510]_  & \new_[65507]_ ;
  assign \new_[65514]_  = A200 & ~A199;
  assign \new_[65517]_  = ~A232 & A203;
  assign \new_[65518]_  = \new_[65517]_  & \new_[65514]_ ;
  assign \new_[65519]_  = \new_[65518]_  & \new_[65511]_ ;
  assign \new_[65522]_  = ~A235 & ~A233;
  assign \new_[65525]_  = A266 & A265;
  assign \new_[65526]_  = \new_[65525]_  & \new_[65522]_ ;
  assign \new_[65529]_  = ~A268 & ~A267;
  assign \new_[65533]_  = A302 & ~A299;
  assign \new_[65534]_  = A298 & \new_[65533]_ ;
  assign \new_[65535]_  = \new_[65534]_  & \new_[65529]_ ;
  assign \new_[65536]_  = \new_[65535]_  & \new_[65526]_ ;
  assign \new_[65539]_  = ~A168 & ~A169;
  assign \new_[65542]_  = A166 & A167;
  assign \new_[65543]_  = \new_[65542]_  & \new_[65539]_ ;
  assign \new_[65546]_  = A200 & ~A199;
  assign \new_[65549]_  = ~A232 & A203;
  assign \new_[65550]_  = \new_[65549]_  & \new_[65546]_ ;
  assign \new_[65551]_  = \new_[65550]_  & \new_[65543]_ ;
  assign \new_[65554]_  = ~A235 & ~A233;
  assign \new_[65557]_  = A266 & A265;
  assign \new_[65558]_  = \new_[65557]_  & \new_[65554]_ ;
  assign \new_[65561]_  = ~A268 & ~A267;
  assign \new_[65565]_  = A302 & A299;
  assign \new_[65566]_  = ~A298 & \new_[65565]_ ;
  assign \new_[65567]_  = \new_[65566]_  & \new_[65561]_ ;
  assign \new_[65568]_  = \new_[65567]_  & \new_[65558]_ ;
  assign \new_[65571]_  = ~A168 & ~A169;
  assign \new_[65574]_  = A166 & A167;
  assign \new_[65575]_  = \new_[65574]_  & \new_[65571]_ ;
  assign \new_[65578]_  = ~A200 & A199;
  assign \new_[65581]_  = ~A234 & A203;
  assign \new_[65582]_  = \new_[65581]_  & \new_[65578]_ ;
  assign \new_[65583]_  = \new_[65582]_  & \new_[65575]_ ;
  assign \new_[65586]_  = ~A236 & ~A235;
  assign \new_[65589]_  = A266 & A265;
  assign \new_[65590]_  = \new_[65589]_  & \new_[65586]_ ;
  assign \new_[65593]_  = ~A268 & ~A267;
  assign \new_[65597]_  = A302 & ~A299;
  assign \new_[65598]_  = A298 & \new_[65597]_ ;
  assign \new_[65599]_  = \new_[65598]_  & \new_[65593]_ ;
  assign \new_[65600]_  = \new_[65599]_  & \new_[65590]_ ;
  assign \new_[65603]_  = ~A168 & ~A169;
  assign \new_[65606]_  = A166 & A167;
  assign \new_[65607]_  = \new_[65606]_  & \new_[65603]_ ;
  assign \new_[65610]_  = ~A200 & A199;
  assign \new_[65613]_  = ~A234 & A203;
  assign \new_[65614]_  = \new_[65613]_  & \new_[65610]_ ;
  assign \new_[65615]_  = \new_[65614]_  & \new_[65607]_ ;
  assign \new_[65618]_  = ~A236 & ~A235;
  assign \new_[65621]_  = A266 & A265;
  assign \new_[65622]_  = \new_[65621]_  & \new_[65618]_ ;
  assign \new_[65625]_  = ~A268 & ~A267;
  assign \new_[65629]_  = A302 & A299;
  assign \new_[65630]_  = ~A298 & \new_[65629]_ ;
  assign \new_[65631]_  = \new_[65630]_  & \new_[65625]_ ;
  assign \new_[65632]_  = \new_[65631]_  & \new_[65622]_ ;
  assign \new_[65635]_  = ~A168 & ~A169;
  assign \new_[65638]_  = A166 & A167;
  assign \new_[65639]_  = \new_[65638]_  & \new_[65635]_ ;
  assign \new_[65642]_  = ~A200 & A199;
  assign \new_[65645]_  = A232 & A203;
  assign \new_[65646]_  = \new_[65645]_  & \new_[65642]_ ;
  assign \new_[65647]_  = \new_[65646]_  & \new_[65639]_ ;
  assign \new_[65650]_  = ~A234 & A233;
  assign \new_[65653]_  = ~A267 & ~A235;
  assign \new_[65654]_  = \new_[65653]_  & \new_[65650]_ ;
  assign \new_[65657]_  = ~A269 & ~A268;
  assign \new_[65661]_  = A302 & ~A299;
  assign \new_[65662]_  = A298 & \new_[65661]_ ;
  assign \new_[65663]_  = \new_[65662]_  & \new_[65657]_ ;
  assign \new_[65664]_  = \new_[65663]_  & \new_[65654]_ ;
  assign \new_[65667]_  = ~A168 & ~A169;
  assign \new_[65670]_  = A166 & A167;
  assign \new_[65671]_  = \new_[65670]_  & \new_[65667]_ ;
  assign \new_[65674]_  = ~A200 & A199;
  assign \new_[65677]_  = A232 & A203;
  assign \new_[65678]_  = \new_[65677]_  & \new_[65674]_ ;
  assign \new_[65679]_  = \new_[65678]_  & \new_[65671]_ ;
  assign \new_[65682]_  = ~A234 & A233;
  assign \new_[65685]_  = ~A267 & ~A235;
  assign \new_[65686]_  = \new_[65685]_  & \new_[65682]_ ;
  assign \new_[65689]_  = ~A269 & ~A268;
  assign \new_[65693]_  = A302 & A299;
  assign \new_[65694]_  = ~A298 & \new_[65693]_ ;
  assign \new_[65695]_  = \new_[65694]_  & \new_[65689]_ ;
  assign \new_[65696]_  = \new_[65695]_  & \new_[65686]_ ;
  assign \new_[65699]_  = ~A168 & ~A169;
  assign \new_[65702]_  = A166 & A167;
  assign \new_[65703]_  = \new_[65702]_  & \new_[65699]_ ;
  assign \new_[65706]_  = ~A200 & A199;
  assign \new_[65709]_  = A232 & A203;
  assign \new_[65710]_  = \new_[65709]_  & \new_[65706]_ ;
  assign \new_[65711]_  = \new_[65710]_  & \new_[65703]_ ;
  assign \new_[65714]_  = ~A234 & A233;
  assign \new_[65717]_  = A265 & ~A235;
  assign \new_[65718]_  = \new_[65717]_  & \new_[65714]_ ;
  assign \new_[65721]_  = ~A267 & A266;
  assign \new_[65725]_  = A300 & A299;
  assign \new_[65726]_  = ~A268 & \new_[65725]_ ;
  assign \new_[65727]_  = \new_[65726]_  & \new_[65721]_ ;
  assign \new_[65728]_  = \new_[65727]_  & \new_[65718]_ ;
  assign \new_[65731]_  = ~A168 & ~A169;
  assign \new_[65734]_  = A166 & A167;
  assign \new_[65735]_  = \new_[65734]_  & \new_[65731]_ ;
  assign \new_[65738]_  = ~A200 & A199;
  assign \new_[65741]_  = A232 & A203;
  assign \new_[65742]_  = \new_[65741]_  & \new_[65738]_ ;
  assign \new_[65743]_  = \new_[65742]_  & \new_[65735]_ ;
  assign \new_[65746]_  = ~A234 & A233;
  assign \new_[65749]_  = A265 & ~A235;
  assign \new_[65750]_  = \new_[65749]_  & \new_[65746]_ ;
  assign \new_[65753]_  = ~A267 & A266;
  assign \new_[65757]_  = A300 & A298;
  assign \new_[65758]_  = ~A268 & \new_[65757]_ ;
  assign \new_[65759]_  = \new_[65758]_  & \new_[65753]_ ;
  assign \new_[65760]_  = \new_[65759]_  & \new_[65750]_ ;
  assign \new_[65763]_  = ~A168 & ~A169;
  assign \new_[65766]_  = A166 & A167;
  assign \new_[65767]_  = \new_[65766]_  & \new_[65763]_ ;
  assign \new_[65770]_  = ~A200 & A199;
  assign \new_[65773]_  = A232 & A203;
  assign \new_[65774]_  = \new_[65773]_  & \new_[65770]_ ;
  assign \new_[65775]_  = \new_[65774]_  & \new_[65767]_ ;
  assign \new_[65778]_  = ~A234 & A233;
  assign \new_[65781]_  = ~A265 & ~A235;
  assign \new_[65782]_  = \new_[65781]_  & \new_[65778]_ ;
  assign \new_[65785]_  = ~A268 & ~A266;
  assign \new_[65789]_  = A302 & ~A299;
  assign \new_[65790]_  = A298 & \new_[65789]_ ;
  assign \new_[65791]_  = \new_[65790]_  & \new_[65785]_ ;
  assign \new_[65792]_  = \new_[65791]_  & \new_[65782]_ ;
  assign \new_[65795]_  = ~A168 & ~A169;
  assign \new_[65798]_  = A166 & A167;
  assign \new_[65799]_  = \new_[65798]_  & \new_[65795]_ ;
  assign \new_[65802]_  = ~A200 & A199;
  assign \new_[65805]_  = A232 & A203;
  assign \new_[65806]_  = \new_[65805]_  & \new_[65802]_ ;
  assign \new_[65807]_  = \new_[65806]_  & \new_[65799]_ ;
  assign \new_[65810]_  = ~A234 & A233;
  assign \new_[65813]_  = ~A265 & ~A235;
  assign \new_[65814]_  = \new_[65813]_  & \new_[65810]_ ;
  assign \new_[65817]_  = ~A268 & ~A266;
  assign \new_[65821]_  = A302 & A299;
  assign \new_[65822]_  = ~A298 & \new_[65821]_ ;
  assign \new_[65823]_  = \new_[65822]_  & \new_[65817]_ ;
  assign \new_[65824]_  = \new_[65823]_  & \new_[65814]_ ;
  assign \new_[65827]_  = ~A168 & ~A169;
  assign \new_[65830]_  = A166 & A167;
  assign \new_[65831]_  = \new_[65830]_  & \new_[65827]_ ;
  assign \new_[65834]_  = ~A200 & A199;
  assign \new_[65837]_  = ~A232 & A203;
  assign \new_[65838]_  = \new_[65837]_  & \new_[65834]_ ;
  assign \new_[65839]_  = \new_[65838]_  & \new_[65831]_ ;
  assign \new_[65842]_  = ~A235 & ~A233;
  assign \new_[65845]_  = A266 & A265;
  assign \new_[65846]_  = \new_[65845]_  & \new_[65842]_ ;
  assign \new_[65849]_  = ~A268 & ~A267;
  assign \new_[65853]_  = A302 & ~A299;
  assign \new_[65854]_  = A298 & \new_[65853]_ ;
  assign \new_[65855]_  = \new_[65854]_  & \new_[65849]_ ;
  assign \new_[65856]_  = \new_[65855]_  & \new_[65846]_ ;
  assign \new_[65859]_  = ~A168 & ~A169;
  assign \new_[65862]_  = A166 & A167;
  assign \new_[65863]_  = \new_[65862]_  & \new_[65859]_ ;
  assign \new_[65866]_  = ~A200 & A199;
  assign \new_[65869]_  = ~A232 & A203;
  assign \new_[65870]_  = \new_[65869]_  & \new_[65866]_ ;
  assign \new_[65871]_  = \new_[65870]_  & \new_[65863]_ ;
  assign \new_[65874]_  = ~A235 & ~A233;
  assign \new_[65877]_  = A266 & A265;
  assign \new_[65878]_  = \new_[65877]_  & \new_[65874]_ ;
  assign \new_[65881]_  = ~A268 & ~A267;
  assign \new_[65885]_  = A302 & A299;
  assign \new_[65886]_  = ~A298 & \new_[65885]_ ;
  assign \new_[65887]_  = \new_[65886]_  & \new_[65881]_ ;
  assign \new_[65888]_  = \new_[65887]_  & \new_[65878]_ ;
  assign \new_[65891]_  = ~A169 & ~A170;
  assign \new_[65894]_  = ~A199 & ~A168;
  assign \new_[65895]_  = \new_[65894]_  & \new_[65891]_ ;
  assign \new_[65898]_  = A203 & A200;
  assign \new_[65901]_  = A233 & A232;
  assign \new_[65902]_  = \new_[65901]_  & \new_[65898]_ ;
  assign \new_[65903]_  = \new_[65902]_  & \new_[65895]_ ;
  assign \new_[65906]_  = ~A235 & ~A234;
  assign \new_[65909]_  = A266 & A265;
  assign \new_[65910]_  = \new_[65909]_  & \new_[65906]_ ;
  assign \new_[65913]_  = ~A268 & ~A267;
  assign \new_[65917]_  = A302 & ~A299;
  assign \new_[65918]_  = A298 & \new_[65917]_ ;
  assign \new_[65919]_  = \new_[65918]_  & \new_[65913]_ ;
  assign \new_[65920]_  = \new_[65919]_  & \new_[65910]_ ;
  assign \new_[65923]_  = ~A169 & ~A170;
  assign \new_[65926]_  = ~A199 & ~A168;
  assign \new_[65927]_  = \new_[65926]_  & \new_[65923]_ ;
  assign \new_[65930]_  = A203 & A200;
  assign \new_[65933]_  = A233 & A232;
  assign \new_[65934]_  = \new_[65933]_  & \new_[65930]_ ;
  assign \new_[65935]_  = \new_[65934]_  & \new_[65927]_ ;
  assign \new_[65938]_  = ~A235 & ~A234;
  assign \new_[65941]_  = A266 & A265;
  assign \new_[65942]_  = \new_[65941]_  & \new_[65938]_ ;
  assign \new_[65945]_  = ~A268 & ~A267;
  assign \new_[65949]_  = A302 & A299;
  assign \new_[65950]_  = ~A298 & \new_[65949]_ ;
  assign \new_[65951]_  = \new_[65950]_  & \new_[65945]_ ;
  assign \new_[65952]_  = \new_[65951]_  & \new_[65942]_ ;
  assign \new_[65955]_  = ~A169 & ~A170;
  assign \new_[65958]_  = A199 & ~A168;
  assign \new_[65959]_  = \new_[65958]_  & \new_[65955]_ ;
  assign \new_[65962]_  = A203 & ~A200;
  assign \new_[65965]_  = A233 & A232;
  assign \new_[65966]_  = \new_[65965]_  & \new_[65962]_ ;
  assign \new_[65967]_  = \new_[65966]_  & \new_[65959]_ ;
  assign \new_[65970]_  = ~A235 & ~A234;
  assign \new_[65973]_  = A266 & A265;
  assign \new_[65974]_  = \new_[65973]_  & \new_[65970]_ ;
  assign \new_[65977]_  = ~A268 & ~A267;
  assign \new_[65981]_  = A302 & ~A299;
  assign \new_[65982]_  = A298 & \new_[65981]_ ;
  assign \new_[65983]_  = \new_[65982]_  & \new_[65977]_ ;
  assign \new_[65984]_  = \new_[65983]_  & \new_[65974]_ ;
  assign \new_[65987]_  = ~A169 & ~A170;
  assign \new_[65990]_  = A199 & ~A168;
  assign \new_[65991]_  = \new_[65990]_  & \new_[65987]_ ;
  assign \new_[65994]_  = A203 & ~A200;
  assign \new_[65997]_  = A233 & A232;
  assign \new_[65998]_  = \new_[65997]_  & \new_[65994]_ ;
  assign \new_[65999]_  = \new_[65998]_  & \new_[65991]_ ;
  assign \new_[66002]_  = ~A235 & ~A234;
  assign \new_[66005]_  = A266 & A265;
  assign \new_[66006]_  = \new_[66005]_  & \new_[66002]_ ;
  assign \new_[66009]_  = ~A268 & ~A267;
  assign \new_[66013]_  = A302 & A299;
  assign \new_[66014]_  = ~A298 & \new_[66013]_ ;
  assign \new_[66015]_  = \new_[66014]_  & \new_[66009]_ ;
  assign \new_[66016]_  = \new_[66015]_  & \new_[66006]_ ;
  assign \new_[66019]_  = A167 & A170;
  assign \new_[66022]_  = A199 & ~A166;
  assign \new_[66023]_  = \new_[66022]_  & \new_[66019]_ ;
  assign \new_[66026]_  = ~A201 & A200;
  assign \new_[66030]_  = A233 & A232;
  assign \new_[66031]_  = ~A202 & \new_[66030]_ ;
  assign \new_[66032]_  = \new_[66031]_  & \new_[66026]_ ;
  assign \new_[66033]_  = \new_[66032]_  & \new_[66023]_ ;
  assign \new_[66036]_  = ~A235 & ~A234;
  assign \new_[66039]_  = A266 & A265;
  assign \new_[66040]_  = \new_[66039]_  & \new_[66036]_ ;
  assign \new_[66043]_  = ~A268 & ~A267;
  assign \new_[66047]_  = A302 & ~A299;
  assign \new_[66048]_  = A298 & \new_[66047]_ ;
  assign \new_[66049]_  = \new_[66048]_  & \new_[66043]_ ;
  assign \new_[66050]_  = \new_[66049]_  & \new_[66040]_ ;
  assign \new_[66053]_  = A167 & A170;
  assign \new_[66056]_  = A199 & ~A166;
  assign \new_[66057]_  = \new_[66056]_  & \new_[66053]_ ;
  assign \new_[66060]_  = ~A201 & A200;
  assign \new_[66064]_  = A233 & A232;
  assign \new_[66065]_  = ~A202 & \new_[66064]_ ;
  assign \new_[66066]_  = \new_[66065]_  & \new_[66060]_ ;
  assign \new_[66067]_  = \new_[66066]_  & \new_[66057]_ ;
  assign \new_[66070]_  = ~A235 & ~A234;
  assign \new_[66073]_  = A266 & A265;
  assign \new_[66074]_  = \new_[66073]_  & \new_[66070]_ ;
  assign \new_[66077]_  = ~A268 & ~A267;
  assign \new_[66081]_  = A302 & A299;
  assign \new_[66082]_  = ~A298 & \new_[66081]_ ;
  assign \new_[66083]_  = \new_[66082]_  & \new_[66077]_ ;
  assign \new_[66084]_  = \new_[66083]_  & \new_[66074]_ ;
  assign \new_[66087]_  = ~A167 & A170;
  assign \new_[66090]_  = A199 & A166;
  assign \new_[66091]_  = \new_[66090]_  & \new_[66087]_ ;
  assign \new_[66094]_  = ~A201 & A200;
  assign \new_[66098]_  = A233 & A232;
  assign \new_[66099]_  = ~A202 & \new_[66098]_ ;
  assign \new_[66100]_  = \new_[66099]_  & \new_[66094]_ ;
  assign \new_[66101]_  = \new_[66100]_  & \new_[66091]_ ;
  assign \new_[66104]_  = ~A235 & ~A234;
  assign \new_[66107]_  = A266 & A265;
  assign \new_[66108]_  = \new_[66107]_  & \new_[66104]_ ;
  assign \new_[66111]_  = ~A268 & ~A267;
  assign \new_[66115]_  = A302 & ~A299;
  assign \new_[66116]_  = A298 & \new_[66115]_ ;
  assign \new_[66117]_  = \new_[66116]_  & \new_[66111]_ ;
  assign \new_[66118]_  = \new_[66117]_  & \new_[66108]_ ;
  assign \new_[66121]_  = ~A167 & A170;
  assign \new_[66124]_  = A199 & A166;
  assign \new_[66125]_  = \new_[66124]_  & \new_[66121]_ ;
  assign \new_[66128]_  = ~A201 & A200;
  assign \new_[66132]_  = A233 & A232;
  assign \new_[66133]_  = ~A202 & \new_[66132]_ ;
  assign \new_[66134]_  = \new_[66133]_  & \new_[66128]_ ;
  assign \new_[66135]_  = \new_[66134]_  & \new_[66125]_ ;
  assign \new_[66138]_  = ~A235 & ~A234;
  assign \new_[66141]_  = A266 & A265;
  assign \new_[66142]_  = \new_[66141]_  & \new_[66138]_ ;
  assign \new_[66145]_  = ~A268 & ~A267;
  assign \new_[66149]_  = A302 & A299;
  assign \new_[66150]_  = ~A298 & \new_[66149]_ ;
  assign \new_[66151]_  = \new_[66150]_  & \new_[66145]_ ;
  assign \new_[66152]_  = \new_[66151]_  & \new_[66142]_ ;
  assign \new_[66155]_  = ~A168 & ~A169;
  assign \new_[66158]_  = A166 & A167;
  assign \new_[66159]_  = \new_[66158]_  & \new_[66155]_ ;
  assign \new_[66162]_  = A200 & ~A199;
  assign \new_[66166]_  = A233 & A232;
  assign \new_[66167]_  = A203 & \new_[66166]_ ;
  assign \new_[66168]_  = \new_[66167]_  & \new_[66162]_ ;
  assign \new_[66169]_  = \new_[66168]_  & \new_[66159]_ ;
  assign \new_[66172]_  = ~A235 & ~A234;
  assign \new_[66175]_  = A266 & A265;
  assign \new_[66176]_  = \new_[66175]_  & \new_[66172]_ ;
  assign \new_[66179]_  = ~A268 & ~A267;
  assign \new_[66183]_  = A302 & ~A299;
  assign \new_[66184]_  = A298 & \new_[66183]_ ;
  assign \new_[66185]_  = \new_[66184]_  & \new_[66179]_ ;
  assign \new_[66186]_  = \new_[66185]_  & \new_[66176]_ ;
  assign \new_[66189]_  = ~A168 & ~A169;
  assign \new_[66192]_  = A166 & A167;
  assign \new_[66193]_  = \new_[66192]_  & \new_[66189]_ ;
  assign \new_[66196]_  = A200 & ~A199;
  assign \new_[66200]_  = A233 & A232;
  assign \new_[66201]_  = A203 & \new_[66200]_ ;
  assign \new_[66202]_  = \new_[66201]_  & \new_[66196]_ ;
  assign \new_[66203]_  = \new_[66202]_  & \new_[66193]_ ;
  assign \new_[66206]_  = ~A235 & ~A234;
  assign \new_[66209]_  = A266 & A265;
  assign \new_[66210]_  = \new_[66209]_  & \new_[66206]_ ;
  assign \new_[66213]_  = ~A268 & ~A267;
  assign \new_[66217]_  = A302 & A299;
  assign \new_[66218]_  = ~A298 & \new_[66217]_ ;
  assign \new_[66219]_  = \new_[66218]_  & \new_[66213]_ ;
  assign \new_[66220]_  = \new_[66219]_  & \new_[66210]_ ;
  assign \new_[66223]_  = ~A168 & ~A169;
  assign \new_[66226]_  = A166 & A167;
  assign \new_[66227]_  = \new_[66226]_  & \new_[66223]_ ;
  assign \new_[66230]_  = ~A200 & A199;
  assign \new_[66234]_  = A233 & A232;
  assign \new_[66235]_  = A203 & \new_[66234]_ ;
  assign \new_[66236]_  = \new_[66235]_  & \new_[66230]_ ;
  assign \new_[66237]_  = \new_[66236]_  & \new_[66227]_ ;
  assign \new_[66240]_  = ~A235 & ~A234;
  assign \new_[66243]_  = A266 & A265;
  assign \new_[66244]_  = \new_[66243]_  & \new_[66240]_ ;
  assign \new_[66247]_  = ~A268 & ~A267;
  assign \new_[66251]_  = A302 & ~A299;
  assign \new_[66252]_  = A298 & \new_[66251]_ ;
  assign \new_[66253]_  = \new_[66252]_  & \new_[66247]_ ;
  assign \new_[66254]_  = \new_[66253]_  & \new_[66244]_ ;
  assign \new_[66257]_  = ~A168 & ~A169;
  assign \new_[66260]_  = A166 & A167;
  assign \new_[66261]_  = \new_[66260]_  & \new_[66257]_ ;
  assign \new_[66264]_  = ~A200 & A199;
  assign \new_[66268]_  = A233 & A232;
  assign \new_[66269]_  = A203 & \new_[66268]_ ;
  assign \new_[66270]_  = \new_[66269]_  & \new_[66264]_ ;
  assign \new_[66271]_  = \new_[66270]_  & \new_[66261]_ ;
  assign \new_[66274]_  = ~A235 & ~A234;
  assign \new_[66277]_  = A266 & A265;
  assign \new_[66278]_  = \new_[66277]_  & \new_[66274]_ ;
  assign \new_[66281]_  = ~A268 & ~A267;
  assign \new_[66285]_  = A302 & A299;
  assign \new_[66286]_  = ~A298 & \new_[66285]_ ;
  assign \new_[66287]_  = \new_[66286]_  & \new_[66281]_ ;
  assign \new_[66288]_  = \new_[66287]_  & \new_[66278]_ ;
endmodule


