module top ( clock, 
    p_10, p_12, p_11, pclk, p_14, p_13, p_16, p_15, p_9, p_18, p_8, p_17,
    p_7, p_6, p_5, p_4, p_3, p_1,
    p_50  );
  input  clock;
  input  p_10, p_12, p_11, pclk, p_14, p_13, p_16, p_15, p_9, p_18, p_8,
    p_17, p_7, p_6, p_5, p_4, p_3, p_1;
  output p_50;
  reg n_28, n_24, n_25, n_26, n_27, n_20, n_21, n_22, n_23, n_2, n_29, n_40,
    n_30, n_39, n_31, n_42, n_32, n_41, n_33, n_44, n_34, n_43, n_35, n_46,
    n_36, n_45, n_37, n_48, n_38, n_47;
  wire new_n110_1_, new_n111_, new_n112_, new_n113_, new_n114_, new_n115_1_,
    new_n117_, new_n118_, new_n119_, new_n120_1_, new_n121_, new_n122_,
    new_n124_, new_n125_1_, new_n126_, new_n127_, new_n128_, new_n129_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_1_, new_n136_,
    new_n138_, new_n139_, new_n140_1_, new_n141_, new_n142_, new_n143_,
    new_n145_1_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_1_,
    new_n152_, new_n153_, new_n154_, new_n155_1_, new_n156_, new_n157_,
    new_n159_, new_n160_1_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n166_, new_n167_, new_n168_, new_n169_, new_n170_1_, new_n171_,
    new_n173_, new_n174_, new_n175_1_, new_n176_, new_n177_, new_n178_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_1_, new_n186_,
    new_n188_, new_n189_, new_n190_, new_n191_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n224_, new_n225_, new_n226_, new_n227_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n286_, new_n287_, new_n288_, new_n289_, n40,
    n45, n50, n55, n60, n65, n70, n75, n80, n85, n90, n95, n100, n105,
    n110, n115, n120, n125, n130, n135, n140, n145, n150, n155, n160, n165,
    n170, n175, n180, n185;
  assign new_n110_1_ = ~n_20 & n_34;
  assign new_n111_ = n_20 & ~n_34;
  assign new_n112_ = ~new_n110_1_ & ~new_n111_;
  assign new_n113_ = p_3 & p_1;
  assign new_n114_ = ~new_n112_ & ~new_n113_;
  assign new_n115_1_ = new_n112_ & new_n113_;
  assign p_50 = new_n114_ | new_n115_1_;
  assign new_n117_ = ~n_29 & n_43;
  assign new_n118_ = n_29 & ~n_43;
  assign new_n119_ = ~new_n117_ & ~new_n118_;
  assign new_n120_1_ = p_12 & p_1;
  assign new_n121_ = ~new_n119_ & ~new_n120_1_;
  assign new_n122_ = new_n119_ & new_n120_1_;
  assign n40 = new_n121_ | new_n122_;
  assign new_n124_ = ~n_25 & n_39;
  assign new_n125_1_ = n_25 & ~n_39;
  assign new_n126_ = ~new_n124_ & ~new_n125_1_;
  assign new_n127_ = p_8 & p_1;
  assign new_n128_ = ~new_n126_ & ~new_n127_;
  assign new_n129_ = new_n126_ & new_n127_;
  assign n45 = new_n128_ | new_n129_;
  assign new_n131_ = ~n_26 & n_40;
  assign new_n132_ = n_26 & ~n_40;
  assign new_n133_ = ~new_n131_ & ~new_n132_;
  assign new_n134_ = p_9 & p_1;
  assign new_n135_1_ = ~new_n133_ & ~new_n134_;
  assign new_n136_ = new_n133_ & new_n134_;
  assign n50 = new_n135_1_ | new_n136_;
  assign new_n138_ = ~n_27 & n_41;
  assign new_n139_ = n_27 & ~n_41;
  assign new_n140_1_ = ~new_n138_ & ~new_n139_;
  assign new_n141_ = p_10 & p_1;
  assign new_n142_ = ~new_n140_1_ & ~new_n141_;
  assign new_n143_ = new_n140_1_ & new_n141_;
  assign n55 = new_n142_ | new_n143_;
  assign new_n145_1_ = ~n_28 & n_42;
  assign new_n146_ = n_28 & ~n_42;
  assign new_n147_ = ~new_n145_1_ & ~new_n146_;
  assign new_n148_ = p_11 & p_1;
  assign new_n149_ = ~new_n147_ & ~new_n148_;
  assign new_n150_1_ = new_n147_ & new_n148_;
  assign n60 = new_n149_ | new_n150_1_;
  assign new_n152_ = ~n_21 & n_35;
  assign new_n153_ = n_21 & ~n_35;
  assign new_n154_ = ~new_n152_ & ~new_n153_;
  assign new_n155_1_ = p_4 & p_1;
  assign new_n156_ = ~new_n154_ & ~new_n155_1_;
  assign new_n157_ = new_n154_ & new_n155_1_;
  assign n65 = new_n156_ | new_n157_;
  assign new_n159_ = ~n_22 & n_36;
  assign new_n160_1_ = n_22 & ~n_36;
  assign new_n161_ = ~new_n159_ & ~new_n160_1_;
  assign new_n162_ = p_5 & p_1;
  assign new_n163_ = ~new_n161_ & ~new_n162_;
  assign new_n164_ = new_n161_ & new_n162_;
  assign n70 = new_n163_ | new_n164_;
  assign new_n166_ = ~n_23 & n_37;
  assign new_n167_ = n_23 & ~n_37;
  assign new_n168_ = ~new_n166_ & ~new_n167_;
  assign new_n169_ = p_6 & p_1;
  assign new_n170_1_ = ~new_n168_ & ~new_n169_;
  assign new_n171_ = new_n168_ & new_n169_;
  assign n75 = new_n170_1_ | new_n171_;
  assign new_n173_ = ~n_24 & n_38;
  assign new_n174_ = n_24 & ~n_38;
  assign new_n175_1_ = ~new_n173_ & ~new_n174_;
  assign new_n176_ = p_7 & p_1;
  assign new_n177_ = ~new_n175_1_ & ~new_n176_;
  assign new_n178_ = new_n175_1_ & new_n176_;
  assign n80 = new_n177_ | new_n178_;
  assign n85 = p_18 & p_1;
  assign new_n181_ = ~n_30 & n_44;
  assign new_n182_ = n_30 & ~n_44;
  assign new_n183_ = ~new_n181_ & ~new_n182_;
  assign new_n184_ = p_13 & p_1;
  assign new_n185_1_ = ~new_n183_ & ~new_n184_;
  assign new_n186_ = new_n183_ & new_n184_;
  assign n90 = new_n185_1_ | new_n186_;
  assign new_n188_ = n_26 & new_n134_;
  assign new_n189_ = n_40 & new_n134_;
  assign new_n190_ = ~new_n188_ & ~new_n189_;
  assign new_n191_ = n_26 & n_40;
  assign n95 = ~new_n190_ | new_n191_;
  assign new_n193_ = ~n_31 & n_45;
  assign new_n194_ = n_31 & ~n_45;
  assign new_n195_ = ~new_n193_ & ~new_n194_;
  assign new_n196_ = p_14 & p_1;
  assign new_n197_ = ~new_n195_ & ~new_n196_;
  assign new_n198_ = new_n195_ & new_n196_;
  assign n100 = new_n197_ | new_n198_;
  assign new_n200_ = n_25 & new_n127_;
  assign new_n201_ = n_39 & new_n127_;
  assign new_n202_ = ~new_n200_ & ~new_n201_;
  assign new_n203_ = n_25 & n_39;
  assign n105 = ~new_n202_ | new_n203_;
  assign new_n205_ = ~n_32 & n_46;
  assign new_n206_ = n_32 & ~n_46;
  assign new_n207_ = ~new_n205_ & ~new_n206_;
  assign new_n208_ = p_15 & p_1;
  assign new_n209_ = ~new_n207_ & ~new_n208_;
  assign new_n210_ = new_n207_ & new_n208_;
  assign n110 = new_n209_ | new_n210_;
  assign new_n212_ = n_28 & new_n148_;
  assign new_n213_ = n_42 & new_n148_;
  assign new_n214_ = ~new_n212_ & ~new_n213_;
  assign new_n215_ = n_28 & n_42;
  assign n115 = ~new_n214_ | new_n215_;
  assign new_n217_ = ~n_33 & n_47;
  assign new_n218_ = n_33 & ~n_47;
  assign new_n219_ = ~new_n217_ & ~new_n218_;
  assign new_n220_ = p_16 & p_1;
  assign new_n221_ = ~new_n219_ & ~new_n220_;
  assign new_n222_ = new_n219_ & new_n220_;
  assign n120 = new_n221_ | new_n222_;
  assign new_n224_ = n_27 & new_n141_;
  assign new_n225_ = n_41 & new_n141_;
  assign new_n226_ = ~new_n224_ & ~new_n225_;
  assign new_n227_ = n_27 & n_41;
  assign n125 = ~new_n226_ | new_n227_;
  assign new_n229_ = ~n_2 & n_48;
  assign new_n230_ = n_2 & ~n_48;
  assign new_n231_ = ~new_n229_ & ~new_n230_;
  assign new_n232_ = p_17 & p_1;
  assign new_n233_ = ~new_n231_ & ~new_n232_;
  assign new_n234_ = new_n231_ & new_n232_;
  assign n130 = new_n233_ | new_n234_;
  assign new_n236_ = n_30 & new_n184_;
  assign new_n237_ = n_44 & new_n184_;
  assign new_n238_ = ~new_n236_ & ~new_n237_;
  assign new_n239_ = n_30 & n_44;
  assign n135 = ~new_n238_ | new_n239_;
  assign new_n241_ = n_20 & new_n113_;
  assign new_n242_ = n_34 & new_n113_;
  assign new_n243_ = ~new_n241_ & ~new_n242_;
  assign new_n244_ = n_20 & n_34;
  assign n140 = ~new_n243_ | new_n244_;
  assign new_n246_ = n_29 & new_n120_1_;
  assign new_n247_ = n_43 & new_n120_1_;
  assign new_n248_ = ~new_n246_ & ~new_n247_;
  assign new_n249_ = n_29 & n_43;
  assign n145 = ~new_n248_ | new_n249_;
  assign new_n251_ = n_21 & new_n155_1_;
  assign new_n252_ = n_35 & new_n155_1_;
  assign new_n253_ = ~new_n251_ & ~new_n252_;
  assign new_n254_ = n_21 & n_35;
  assign n150 = ~new_n253_ | new_n254_;
  assign new_n256_ = n_32 & new_n208_;
  assign new_n257_ = n_46 & new_n208_;
  assign new_n258_ = ~new_n256_ & ~new_n257_;
  assign new_n259_ = n_32 & n_46;
  assign n155 = ~new_n258_ | new_n259_;
  assign new_n261_ = n_22 & new_n162_;
  assign new_n262_ = n_36 & new_n162_;
  assign new_n263_ = ~new_n261_ & ~new_n262_;
  assign new_n264_ = n_22 & n_36;
  assign n160 = ~new_n263_ | new_n264_;
  assign new_n266_ = n_31 & new_n196_;
  assign new_n267_ = n_45 & new_n196_;
  assign new_n268_ = ~new_n266_ & ~new_n267_;
  assign new_n269_ = n_31 & n_45;
  assign n165 = ~new_n268_ | new_n269_;
  assign new_n271_ = n_23 & new_n169_;
  assign new_n272_ = n_37 & new_n169_;
  assign new_n273_ = ~new_n271_ & ~new_n272_;
  assign new_n274_ = n_23 & n_37;
  assign n170 = ~new_n273_ | new_n274_;
  assign new_n276_ = n_2 & new_n232_;
  assign new_n277_ = n_48 & new_n232_;
  assign new_n278_ = ~new_n276_ & ~new_n277_;
  assign new_n279_ = n_2 & n_48;
  assign n175 = ~new_n278_ | new_n279_;
  assign new_n281_ = n_24 & new_n176_;
  assign new_n282_ = n_38 & new_n176_;
  assign new_n283_ = ~new_n281_ & ~new_n282_;
  assign new_n284_ = n_24 & n_38;
  assign n180 = ~new_n283_ | new_n284_;
  assign new_n286_ = n_33 & new_n220_;
  assign new_n287_ = n_47 & new_n220_;
  assign new_n288_ = ~new_n286_ & ~new_n287_;
  assign new_n289_ = n_33 & n_47;
  assign n185 = ~new_n288_ | new_n289_;
  always @ (posedge clock) begin
    n_28 <= n40;
    n_24 <= n45;
    n_25 <= n50;
    n_26 <= n55;
    n_27 <= n60;
    n_20 <= n65;
    n_21 <= n70;
    n_22 <= n75;
    n_23 <= n80;
    n_2 <= n85;
    n_29 <= n90;
    n_40 <= n95;
    n_30 <= n100;
    n_39 <= n105;
    n_31 <= n110;
    n_42 <= n115;
    n_32 <= n120;
    n_41 <= n125;
    n_33 <= n130;
    n_44 <= n135;
    n_34 <= n140;
    n_43 <= n145;
    n_35 <= n150;
    n_46 <= n155;
    n_36 <= n160;
    n_45 <= n165;
    n_37 <= n170;
    n_48 <= n175;
    n_38 <= n180;
    n_47 <= n185;
  end
endmodule

