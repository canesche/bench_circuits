module frg2 ( 
    a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, x,
    y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0,
    q0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1,
    j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2,
    b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2,
    t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3,
    l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4,
    d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4,
    o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5,
    g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, x5,
    y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6,
    q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7,
    i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7,
    a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8, r8,
    s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, j9,
    k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9  );
  input  a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u,
    v, w, x, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0,
    o0, p0, q0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1,
    h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1,
    z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2,
    r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3,
    j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4,
    b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4;
  output o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5,
    f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5,
    x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6,
    p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7,
    h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7,
    z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8,
    r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9,
    j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9;
  wire new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_,
    new_n308_, new_n309_, new_n310_, new_n311_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n356_, new_n357_, new_n358_, new_n359_, new_n361_,
    new_n362_, new_n363_, new_n364_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n371_, new_n372_, new_n373_, new_n374_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n395_, new_n397_, new_n399_, new_n401_, new_n403_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n416_, new_n427_,
    new_n428_, new_n430_, new_n431_, new_n432_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n537_, new_n538_, new_n539_,
    new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_,
    new_n546_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_,
    new_n972_, new_n973_, new_n974_, new_n975_, new_n977_, new_n978_,
    new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_,
    new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_,
    new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_,
    new_n1022_, new_n1023_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_,
    new_n1063_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_,
    new_n1070_, new_n1071_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_,
    new_n1118_, new_n1119_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1227_, new_n1228_, new_n1229_, new_n1230_,
    new_n1231_, new_n1232_, new_n1234_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1311_, new_n1312_, new_n1313_, new_n1314_,
    new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_, new_n1321_,
    new_n1322_, new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_,
    new_n1328_, new_n1329_, new_n1330_, new_n1331_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1395_, new_n1396_, new_n1397_, new_n1398_,
    new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_, new_n1404_,
    new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_, new_n1410_,
    new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_, new_n1416_,
    new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_, new_n1422_,
    new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_, new_n1428_,
    new_n1430_, new_n1431_, new_n1432_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_;
  assign new_n283_ = l0 & l3;
  assign new_n284_ = ~d3 & ~new_n283_;
  assign new_n285_ = l0 & ~l3;
  assign new_n286_ = ~new_n284_ & ~new_n285_;
  assign new_n287_ = ~l0 & l3;
  assign new_n288_ = ~d3 & ~new_n287_;
  assign new_n289_ = ~l0 & ~l3;
  assign new_n290_ = ~new_n288_ & ~new_n289_;
  assign new_n291_ = ~m0 & ~t3;
  assign new_n292_ = k0 & ~new_n290_;
  assign new_n293_ = new_n286_ & ~new_n292_;
  assign new_n294_ = k0 & new_n290_;
  assign new_n295_ = m0 & ~new_n294_;
  assign new_n296_ = ~new_n293_ & new_n295_;
  assign p4 = ~new_n291_ & ~new_n296_;
  assign new_n298_ = l0 & k3;
  assign new_n299_ = ~c3 & ~new_n298_;
  assign new_n300_ = l0 & ~k3;
  assign new_n301_ = ~new_n299_ & ~new_n300_;
  assign new_n302_ = ~l0 & k3;
  assign new_n303_ = ~c3 & ~new_n302_;
  assign new_n304_ = ~l0 & ~k3;
  assign new_n305_ = ~new_n303_ & ~new_n304_;
  assign new_n306_ = ~m0 & ~s3;
  assign new_n307_ = k0 & ~new_n305_;
  assign new_n308_ = new_n301_ & ~new_n307_;
  assign new_n309_ = k0 & new_n305_;
  assign new_n310_ = m0 & ~new_n309_;
  assign new_n311_ = ~new_n308_ & new_n310_;
  assign q4 = ~new_n306_ & ~new_n311_;
  assign new_n313_ = l0 & j3;
  assign new_n314_ = ~b3 & ~new_n313_;
  assign new_n315_ = l0 & ~j3;
  assign new_n316_ = ~new_n314_ & ~new_n315_;
  assign new_n317_ = ~l0 & j3;
  assign new_n318_ = ~b3 & ~new_n317_;
  assign new_n319_ = ~l0 & ~j3;
  assign new_n320_ = ~new_n318_ & ~new_n319_;
  assign new_n321_ = ~m0 & ~r3;
  assign new_n322_ = k0 & ~new_n320_;
  assign new_n323_ = new_n316_ & ~new_n322_;
  assign new_n324_ = k0 & new_n320_;
  assign new_n325_ = m0 & ~new_n324_;
  assign new_n326_ = ~new_n323_ & new_n325_;
  assign r4 = ~new_n321_ & ~new_n326_;
  assign new_n328_ = l0 & i3;
  assign new_n329_ = ~a3 & ~new_n328_;
  assign new_n330_ = l0 & ~i3;
  assign new_n331_ = ~new_n329_ & ~new_n330_;
  assign new_n332_ = ~l0 & i3;
  assign new_n333_ = ~a3 & ~new_n332_;
  assign new_n334_ = ~l0 & ~i3;
  assign new_n335_ = ~new_n333_ & ~new_n334_;
  assign new_n336_ = ~m0 & ~q3;
  assign new_n337_ = k0 & ~new_n335_;
  assign new_n338_ = new_n331_ & ~new_n337_;
  assign new_n339_ = k0 & new_n335_;
  assign new_n340_ = m0 & ~new_n339_;
  assign new_n341_ = ~new_n338_ & new_n340_;
  assign s4 = ~new_n336_ & ~new_n341_;
  assign new_n343_ = k0 & l0;
  assign new_n344_ = ~k0 & ~l0;
  assign new_n345_ = ~new_n343_ & ~new_n344_;
  assign new_n346_ = ~e3 & ~new_n345_;
  assign new_n347_ = m0 & ~new_n346_;
  assign new_n348_ = ~m3 & ~new_n344_;
  assign new_n349_ = ~new_n343_ & new_n348_;
  assign v4 = new_n347_ & ~new_n349_;
  assign new_n351_ = ~f3 & ~new_n345_;
  assign new_n352_ = m0 & ~new_n351_;
  assign new_n353_ = ~n3 & ~new_n344_;
  assign new_n354_ = ~new_n343_ & new_n353_;
  assign w4 = new_n352_ & ~new_n354_;
  assign new_n356_ = ~g3 & ~new_n345_;
  assign new_n357_ = m0 & ~new_n356_;
  assign new_n358_ = ~o3 & ~new_n344_;
  assign new_n359_ = ~new_n343_ & new_n358_;
  assign x4 = new_n357_ & ~new_n359_;
  assign new_n361_ = ~h3 & ~new_n345_;
  assign new_n362_ = m0 & ~new_n361_;
  assign new_n363_ = ~p3 & ~new_n344_;
  assign new_n364_ = ~new_n343_ & new_n363_;
  assign y4 = new_n362_ & ~new_n364_;
  assign new_n366_ = ~i3 & ~new_n345_;
  assign new_n367_ = m0 & ~new_n366_;
  assign new_n368_ = ~q3 & ~new_n344_;
  assign new_n369_ = ~new_n343_ & new_n368_;
  assign z4 = new_n367_ & ~new_n369_;
  assign new_n371_ = ~j3 & ~new_n345_;
  assign new_n372_ = m0 & ~new_n371_;
  assign new_n373_ = ~r3 & ~new_n344_;
  assign new_n374_ = ~new_n343_ & new_n373_;
  assign a5 = new_n372_ & ~new_n374_;
  assign new_n376_ = ~k3 & ~new_n345_;
  assign new_n377_ = m0 & ~new_n376_;
  assign new_n378_ = ~s3 & ~new_n344_;
  assign new_n379_ = ~new_n343_ & new_n378_;
  assign b5 = new_n377_ & ~new_n379_;
  assign new_n381_ = ~l3 & ~new_n345_;
  assign new_n382_ = m0 & ~new_n381_;
  assign new_n383_ = ~t3 & ~new_n344_;
  assign new_n384_ = ~new_n343_ & new_n383_;
  assign c5 = new_n382_ & ~new_n384_;
  assign d5 = m0 & m3;
  assign e5 = m0 & n3;
  assign f5 = m0 & o3;
  assign g5 = m0 & p3;
  assign h5 = m0 & q3;
  assign i5 = m0 & r3;
  assign j5 = m0 & s3;
  assign k5 = m0 & t3;
  assign l5 = g1 & ~j4;
  assign new_n395_ = h1 & ~k4;
  assign n5 = n0 | ~new_n395_;
  assign new_n397_ = i1 & ~k4;
  assign o5 = n0 | ~new_n397_;
  assign new_n399_ = j1 & ~k4;
  assign p5 = n0 | ~new_n399_;
  assign new_n401_ = k1 & ~k4;
  assign q5 = n0 | ~new_n401_;
  assign new_n403_ = l1 & ~k4;
  assign r5 = n0 | ~new_n403_;
  assign new_n405_ = y3 & z3;
  assign new_n406_ = ~b4 & ~c4;
  assign new_n407_ = ~a4 & new_n406_;
  assign new_n408_ = ~f1 & i4;
  assign new_n409_ = f1 & ~i4;
  assign new_n410_ = ~new_n408_ & ~new_n409_;
  assign new_n411_ = new_n405_ & new_n407_;
  assign new_n412_ = ~n1 & ~new_n411_;
  assign new_n413_ = new_n407_ & ~new_n410_;
  assign new_n414_ = new_n405_ & new_n413_;
  assign s5 = ~new_n412_ & ~new_n414_;
  assign new_n416_ = m1 & ~k4;
  assign x5 = ~h1 | ~new_n416_;
  assign y5 = ~i1 | ~new_n416_;
  assign z5 = ~j1 | ~new_n416_;
  assign a6 = ~k1 | ~new_n416_;
  assign b6 = ~l1 | ~new_n416_;
  assign c6 = ~h1 | ~l4;
  assign d6 = ~i1 | ~l4;
  assign e6 = ~j1 | ~l4;
  assign f6 = ~k1 | ~l4;
  assign g6 = ~l1 | ~l4;
  assign new_n427_ = f1 & i4;
  assign new_n428_ = ~f1 & ~i4;
  assign n6 = new_n427_ | new_n428_;
  assign new_n430_ = z3 & ~a4;
  assign new_n431_ = x3 & y3;
  assign new_n432_ = new_n430_ & new_n431_;
  assign o6 = new_n406_ & new_n432_;
  assign new_n434_ = ~g4 & ~h4;
  assign new_n435_ = e4 & f4;
  assign new_n436_ = new_n434_ & new_n435_;
  assign new_n437_ = ~g1 & d4;
  assign new_n438_ = new_n435_ & new_n437_;
  assign new_n439_ = new_n434_ & new_n438_;
  assign new_n440_ = ~b1 & l1;
  assign new_n441_ = ~new_n436_ & ~new_n440_;
  assign new_n442_ = n4 & new_n441_;
  assign new_n443_ = ~new_n439_ & ~new_n442_;
  assign new_n444_ = ~z0 & j1;
  assign new_n445_ = ~a1 & k1;
  assign new_n446_ = ~new_n444_ & ~new_n445_;
  assign new_n447_ = ~new_n436_ & ~new_n446_;
  assign new_n448_ = ~new_n443_ & ~new_n447_;
  assign new_n449_ = ~x0 & h1;
  assign new_n450_ = ~y0 & i1;
  assign new_n451_ = ~new_n449_ & ~new_n450_;
  assign new_n452_ = ~new_n436_ & ~new_n451_;
  assign new_n453_ = new_n448_ & ~new_n452_;
  assign new_n454_ = ~q0 & new_n453_;
  assign p6 = o0 & new_n454_;
  assign new_n456_ = ~q0 & ~c1;
  assign new_n457_ = o0 & new_n456_;
  assign new_n458_ = ~i1 & ~j1;
  assign new_n459_ = ~h1 & new_n458_;
  assign new_n460_ = ~k1 & ~l1;
  assign new_n461_ = new_n459_ & new_n460_;
  assign new_n462_ = ~e1 & new_n461_;
  assign new_n463_ = ~d1 & new_n462_;
  assign new_n464_ = ~g1 & h1;
  assign new_n465_ = ~q0 & new_n464_;
  assign new_n466_ = ~c1 & ~d1;
  assign new_n467_ = e1 & ~new_n466_;
  assign new_n468_ = ~n0 & new_n461_;
  assign new_n469_ = ~new_n467_ & new_n468_;
  assign new_n470_ = new_n465_ & ~new_n469_;
  assign new_n471_ = o0 & new_n470_;
  assign new_n472_ = new_n457_ & new_n463_;
  assign new_n473_ = ~n0 & new_n472_;
  assign q6 = new_n471_ | new_n473_;
  assign new_n475_ = d1 & e1;
  assign new_n476_ = ~c1 & ~new_n475_;
  assign new_n477_ = d1 & ~e1;
  assign new_n478_ = ~new_n476_ & ~new_n477_;
  assign new_n479_ = ~n0 & new_n462_;
  assign new_n480_ = ~i1 & ~new_n479_;
  assign new_n481_ = o0 & ~q0;
  assign new_n482_ = ~new_n480_ & new_n481_;
  assign new_n483_ = g1 & ~new_n479_;
  assign new_n484_ = ~n0 & ~new_n478_;
  assign new_n485_ = new_n461_ & new_n484_;
  assign new_n486_ = ~new_n483_ & ~new_n485_;
  assign r6 = new_n482_ & new_n486_;
  assign new_n488_ = c1 & e1;
  assign new_n489_ = ~d1 & ~new_n488_;
  assign new_n490_ = c1 & ~e1;
  assign new_n491_ = ~new_n489_ & ~new_n490_;
  assign new_n492_ = ~j1 & ~new_n479_;
  assign new_n493_ = new_n481_ & ~new_n492_;
  assign new_n494_ = ~n0 & ~new_n491_;
  assign new_n495_ = new_n461_ & new_n494_;
  assign new_n496_ = ~new_n483_ & ~new_n495_;
  assign s6 = new_n493_ & new_n496_;
  assign new_n498_ = ~d1 & ~e1;
  assign new_n499_ = ~new_n476_ & ~new_n498_;
  assign new_n500_ = ~k1 & ~new_n479_;
  assign new_n501_ = new_n481_ & ~new_n500_;
  assign new_n502_ = ~n0 & ~new_n499_;
  assign new_n503_ = new_n461_ & new_n502_;
  assign new_n504_ = ~new_n483_ & ~new_n503_;
  assign t6 = new_n501_ & new_n504_;
  assign new_n506_ = ~d1 & new_n461_;
  assign new_n507_ = ~n0 & ~c1;
  assign new_n508_ = new_n506_ & new_n507_;
  assign new_n509_ = ~q0 & ~new_n479_;
  assign new_n510_ = o0 & new_n509_;
  assign new_n511_ = ~g1 & l1;
  assign new_n512_ = ~new_n508_ & ~new_n511_;
  assign u6 = new_n510_ & ~new_n512_;
  assign new_n514_ = m1 & new_n453_;
  assign new_n515_ = ~q0 & ~new_n514_;
  assign new_n516_ = o0 & new_n515_;
  assign new_n517_ = ~n0 & p0;
  assign new_n518_ = ~m1 & ~new_n517_;
  assign v6 = new_n516_ & ~new_n518_;
  assign new_n520_ = ~x3 & y3;
  assign new_n521_ = new_n430_ & new_n520_;
  assign new_n522_ = new_n406_ & new_n521_;
  assign new_n523_ = ~o1 & l4;
  assign new_n524_ = l4 & ~new_n522_;
  assign new_n525_ = ~j0 & new_n468_;
  assign new_n526_ = ~q0 & ~new_n525_;
  assign new_n527_ = o0 & new_n526_;
  assign new_n528_ = ~new_n461_ & ~new_n524_;
  assign new_n529_ = ~n1 & new_n528_;
  assign new_n530_ = new_n527_ & ~new_n529_;
  assign new_n531_ = n0 & ~new_n524_;
  assign new_n532_ = ~n1 & new_n531_;
  assign new_n533_ = ~new_n468_ & new_n523_;
  assign new_n534_ = ~new_n522_ & new_n533_;
  assign new_n535_ = ~new_n532_ & ~new_n534_;
  assign w6 = new_n530_ & new_n535_;
  assign new_n537_ = ~p1 & l4;
  assign new_n538_ = ~i0 & new_n468_;
  assign new_n539_ = ~q0 & ~new_n538_;
  assign new_n540_ = o0 & new_n539_;
  assign new_n541_ = ~o1 & new_n528_;
  assign new_n542_ = new_n540_ & ~new_n541_;
  assign new_n543_ = ~o1 & new_n531_;
  assign new_n544_ = ~new_n468_ & new_n537_;
  assign new_n545_ = ~new_n522_ & new_n544_;
  assign new_n546_ = ~new_n543_ & ~new_n545_;
  assign x6 = new_n542_ & new_n546_;
  assign new_n548_ = ~q1 & l4;
  assign new_n549_ = ~h0 & new_n468_;
  assign new_n550_ = ~q0 & ~new_n549_;
  assign new_n551_ = o0 & new_n550_;
  assign new_n552_ = ~p1 & new_n528_;
  assign new_n553_ = new_n551_ & ~new_n552_;
  assign new_n554_ = ~p1 & new_n531_;
  assign new_n555_ = ~new_n468_ & new_n548_;
  assign new_n556_ = ~new_n522_ & new_n555_;
  assign new_n557_ = ~new_n554_ & ~new_n556_;
  assign y6 = new_n553_ & new_n557_;
  assign new_n559_ = ~r1 & l4;
  assign new_n560_ = ~g0 & new_n468_;
  assign new_n561_ = ~q0 & ~new_n560_;
  assign new_n562_ = o0 & new_n561_;
  assign new_n563_ = ~q1 & new_n528_;
  assign new_n564_ = new_n562_ & ~new_n563_;
  assign new_n565_ = ~q1 & new_n531_;
  assign new_n566_ = ~new_n468_ & new_n559_;
  assign new_n567_ = ~new_n522_ & new_n566_;
  assign new_n568_ = ~new_n565_ & ~new_n567_;
  assign z6 = new_n564_ & new_n568_;
  assign new_n570_ = ~s1 & l4;
  assign new_n571_ = ~f0 & new_n468_;
  assign new_n572_ = ~q0 & ~new_n571_;
  assign new_n573_ = o0 & new_n572_;
  assign new_n574_ = ~r1 & new_n528_;
  assign new_n575_ = new_n573_ & ~new_n574_;
  assign new_n576_ = ~r1 & new_n531_;
  assign new_n577_ = ~new_n468_ & new_n570_;
  assign new_n578_ = ~new_n522_ & new_n577_;
  assign new_n579_ = ~new_n576_ & ~new_n578_;
  assign a7 = new_n575_ & new_n579_;
  assign new_n581_ = ~t1 & l4;
  assign new_n582_ = ~e0 & new_n468_;
  assign new_n583_ = ~q0 & ~new_n582_;
  assign new_n584_ = o0 & new_n583_;
  assign new_n585_ = ~s1 & new_n528_;
  assign new_n586_ = new_n584_ & ~new_n585_;
  assign new_n587_ = ~s1 & new_n531_;
  assign new_n588_ = ~new_n468_ & new_n581_;
  assign new_n589_ = ~new_n522_ & new_n588_;
  assign new_n590_ = ~new_n587_ & ~new_n589_;
  assign b7 = new_n586_ & new_n590_;
  assign new_n592_ = ~u1 & l4;
  assign new_n593_ = ~d0 & new_n468_;
  assign new_n594_ = ~q0 & ~new_n593_;
  assign new_n595_ = o0 & new_n594_;
  assign new_n596_ = ~t1 & new_n528_;
  assign new_n597_ = new_n595_ & ~new_n596_;
  assign new_n598_ = ~t1 & new_n531_;
  assign new_n599_ = ~new_n468_ & new_n592_;
  assign new_n600_ = ~new_n522_ & new_n599_;
  assign new_n601_ = ~new_n598_ & ~new_n600_;
  assign c7 = new_n597_ & new_n601_;
  assign new_n603_ = ~v1 & l4;
  assign new_n604_ = ~m0 & new_n468_;
  assign new_n605_ = ~q0 & ~new_n604_;
  assign new_n606_ = o0 & new_n605_;
  assign new_n607_ = ~u1 & new_n528_;
  assign new_n608_ = new_n606_ & ~new_n607_;
  assign new_n609_ = ~u1 & new_n531_;
  assign new_n610_ = ~new_n468_ & new_n603_;
  assign new_n611_ = ~new_n522_ & new_n610_;
  assign new_n612_ = ~new_n609_ & ~new_n611_;
  assign d7 = new_n608_ & new_n612_;
  assign new_n614_ = ~w1 & l4;
  assign new_n615_ = ~k0 & new_n468_;
  assign new_n616_ = ~q0 & ~new_n615_;
  assign new_n617_ = o0 & new_n616_;
  assign new_n618_ = ~v1 & new_n528_;
  assign new_n619_ = new_n617_ & ~new_n618_;
  assign new_n620_ = ~v1 & new_n531_;
  assign new_n621_ = ~new_n468_ & new_n614_;
  assign new_n622_ = ~new_n522_ & new_n621_;
  assign new_n623_ = ~new_n620_ & ~new_n622_;
  assign e7 = new_n619_ & new_n623_;
  assign new_n625_ = ~x1 & l4;
  assign new_n626_ = ~l0 & new_n468_;
  assign new_n627_ = ~q0 & ~new_n626_;
  assign new_n628_ = o0 & new_n627_;
  assign new_n629_ = ~w1 & new_n528_;
  assign new_n630_ = new_n628_ & ~new_n629_;
  assign new_n631_ = ~w1 & new_n531_;
  assign new_n632_ = ~new_n468_ & new_n625_;
  assign new_n633_ = ~new_n522_ & new_n632_;
  assign new_n634_ = ~new_n631_ & ~new_n633_;
  assign f7 = new_n630_ & new_n634_;
  assign new_n636_ = ~y1 & l4;
  assign new_n637_ = ~q & new_n468_;
  assign new_n638_ = ~q0 & ~new_n637_;
  assign new_n639_ = o0 & new_n638_;
  assign new_n640_ = ~x1 & new_n528_;
  assign new_n641_ = new_n639_ & ~new_n640_;
  assign new_n642_ = ~x1 & new_n531_;
  assign new_n643_ = ~new_n468_ & new_n636_;
  assign new_n644_ = ~new_n522_ & new_n643_;
  assign new_n645_ = ~new_n642_ & ~new_n644_;
  assign g7 = new_n641_ & new_n645_;
  assign new_n647_ = ~z1 & l4;
  assign new_n648_ = ~r & new_n468_;
  assign new_n649_ = ~q0 & ~new_n648_;
  assign new_n650_ = o0 & new_n649_;
  assign new_n651_ = ~y1 & new_n528_;
  assign new_n652_ = new_n650_ & ~new_n651_;
  assign new_n653_ = ~y1 & new_n531_;
  assign new_n654_ = ~new_n468_ & new_n647_;
  assign new_n655_ = ~new_n522_ & new_n654_;
  assign new_n656_ = ~new_n653_ & ~new_n655_;
  assign h7 = new_n652_ & new_n656_;
  assign new_n658_ = ~a2 & l4;
  assign new_n659_ = ~s & new_n468_;
  assign new_n660_ = ~q0 & ~new_n659_;
  assign new_n661_ = o0 & new_n660_;
  assign new_n662_ = ~z1 & new_n528_;
  assign new_n663_ = new_n661_ & ~new_n662_;
  assign new_n664_ = ~z1 & new_n531_;
  assign new_n665_ = ~new_n468_ & new_n658_;
  assign new_n666_ = ~new_n522_ & new_n665_;
  assign new_n667_ = ~new_n664_ & ~new_n666_;
  assign i7 = new_n663_ & new_n667_;
  assign new_n669_ = ~b2 & l4;
  assign new_n670_ = ~t & new_n468_;
  assign new_n671_ = ~q0 & ~new_n670_;
  assign new_n672_ = o0 & new_n671_;
  assign new_n673_ = ~a2 & new_n528_;
  assign new_n674_ = new_n672_ & ~new_n673_;
  assign new_n675_ = ~a2 & new_n531_;
  assign new_n676_ = ~new_n468_ & new_n669_;
  assign new_n677_ = ~new_n522_ & new_n676_;
  assign new_n678_ = ~new_n675_ & ~new_n677_;
  assign j7 = new_n674_ & new_n678_;
  assign new_n680_ = ~c2 & l4;
  assign new_n681_ = ~u & new_n468_;
  assign new_n682_ = ~q0 & ~new_n681_;
  assign new_n683_ = o0 & new_n682_;
  assign new_n684_ = ~b2 & new_n528_;
  assign new_n685_ = new_n683_ & ~new_n684_;
  assign new_n686_ = ~b2 & new_n531_;
  assign new_n687_ = ~new_n468_ & new_n680_;
  assign new_n688_ = ~new_n522_ & new_n687_;
  assign new_n689_ = ~new_n686_ & ~new_n688_;
  assign k7 = new_n685_ & new_n689_;
  assign new_n691_ = ~d2 & l4;
  assign new_n692_ = ~v & new_n468_;
  assign new_n693_ = ~q0 & ~new_n692_;
  assign new_n694_ = o0 & new_n693_;
  assign new_n695_ = ~c2 & new_n528_;
  assign new_n696_ = new_n694_ & ~new_n695_;
  assign new_n697_ = ~c2 & new_n531_;
  assign new_n698_ = ~new_n468_ & new_n691_;
  assign new_n699_ = ~new_n522_ & new_n698_;
  assign new_n700_ = ~new_n697_ & ~new_n699_;
  assign l7 = new_n696_ & new_n700_;
  assign new_n702_ = ~e2 & l4;
  assign new_n703_ = ~w & new_n468_;
  assign new_n704_ = ~q0 & ~new_n703_;
  assign new_n705_ = o0 & new_n704_;
  assign new_n706_ = ~d2 & new_n528_;
  assign new_n707_ = new_n705_ & ~new_n706_;
  assign new_n708_ = ~d2 & new_n531_;
  assign new_n709_ = ~new_n468_ & new_n702_;
  assign new_n710_ = ~new_n522_ & new_n709_;
  assign new_n711_ = ~new_n708_ & ~new_n710_;
  assign m7 = new_n707_ & new_n711_;
  assign new_n713_ = ~f2 & l4;
  assign new_n714_ = ~x & new_n468_;
  assign new_n715_ = ~q0 & ~new_n714_;
  assign new_n716_ = o0 & new_n715_;
  assign new_n717_ = ~e2 & new_n528_;
  assign new_n718_ = new_n716_ & ~new_n717_;
  assign new_n719_ = ~e2 & new_n531_;
  assign new_n720_ = ~new_n468_ & new_n713_;
  assign new_n721_ = ~new_n522_ & new_n720_;
  assign new_n722_ = ~new_n719_ & ~new_n721_;
  assign n7 = new_n718_ & new_n722_;
  assign new_n724_ = ~g2 & l4;
  assign new_n725_ = ~y & new_n468_;
  assign new_n726_ = ~q0 & ~new_n725_;
  assign new_n727_ = o0 & new_n726_;
  assign new_n728_ = ~f2 & new_n528_;
  assign new_n729_ = new_n727_ & ~new_n728_;
  assign new_n730_ = ~f2 & new_n531_;
  assign new_n731_ = ~new_n468_ & new_n724_;
  assign new_n732_ = ~new_n522_ & new_n731_;
  assign new_n733_ = ~new_n730_ & ~new_n732_;
  assign o7 = new_n729_ & new_n733_;
  assign new_n735_ = ~h2 & l4;
  assign new_n736_ = ~z & new_n468_;
  assign new_n737_ = ~q0 & ~new_n736_;
  assign new_n738_ = o0 & new_n737_;
  assign new_n739_ = ~g2 & new_n528_;
  assign new_n740_ = new_n738_ & ~new_n739_;
  assign new_n741_ = ~g2 & new_n531_;
  assign new_n742_ = ~new_n468_ & new_n735_;
  assign new_n743_ = ~new_n522_ & new_n742_;
  assign new_n744_ = ~new_n741_ & ~new_n743_;
  assign p7 = new_n740_ & new_n744_;
  assign new_n746_ = ~i2 & l4;
  assign new_n747_ = ~a0 & new_n468_;
  assign new_n748_ = ~q0 & ~new_n747_;
  assign new_n749_ = o0 & new_n748_;
  assign new_n750_ = ~h2 & new_n528_;
  assign new_n751_ = new_n749_ & ~new_n750_;
  assign new_n752_ = ~h2 & new_n531_;
  assign new_n753_ = ~new_n468_ & new_n746_;
  assign new_n754_ = ~new_n522_ & new_n753_;
  assign new_n755_ = ~new_n752_ & ~new_n754_;
  assign q7 = new_n751_ & new_n755_;
  assign new_n757_ = ~j2 & l4;
  assign new_n758_ = ~b0 & new_n468_;
  assign new_n759_ = ~q0 & ~new_n758_;
  assign new_n760_ = o0 & new_n759_;
  assign new_n761_ = ~i2 & new_n528_;
  assign new_n762_ = new_n760_ & ~new_n761_;
  assign new_n763_ = ~i2 & new_n531_;
  assign new_n764_ = ~new_n468_ & new_n757_;
  assign new_n765_ = ~new_n522_ & new_n764_;
  assign new_n766_ = ~new_n763_ & ~new_n765_;
  assign r7 = new_n762_ & new_n766_;
  assign new_n768_ = ~k2 & l4;
  assign new_n769_ = ~c0 & new_n468_;
  assign new_n770_ = ~q0 & ~new_n769_;
  assign new_n771_ = o0 & new_n770_;
  assign new_n772_ = ~j2 & new_n528_;
  assign new_n773_ = new_n771_ & ~new_n772_;
  assign new_n774_ = ~j2 & new_n531_;
  assign new_n775_ = ~new_n468_ & new_n768_;
  assign new_n776_ = ~new_n522_ & new_n775_;
  assign new_n777_ = ~new_n774_ & ~new_n776_;
  assign s7 = new_n773_ & new_n777_;
  assign new_n779_ = i & ~l0;
  assign new_n780_ = k0 & new_n779_;
  assign new_n781_ = k0 & ~l0;
  assign new_n782_ = a & ~new_n781_;
  assign new_n783_ = ~new_n780_ & ~new_n782_;
  assign new_n784_ = ~l2 & l4;
  assign new_n785_ = ~new_n524_ & ~new_n604_;
  assign new_n786_ = ~k2 & new_n785_;
  assign new_n787_ = new_n468_ & new_n783_;
  assign new_n788_ = ~m0 & new_n787_;
  assign new_n789_ = ~new_n604_ & new_n784_;
  assign new_n790_ = ~new_n522_ & new_n789_;
  assign new_n791_ = ~new_n788_ & ~new_n790_;
  assign new_n792_ = ~new_n786_ & new_n791_;
  assign t7 = new_n481_ & new_n792_;
  assign new_n794_ = j & ~l0;
  assign new_n795_ = k0 & new_n794_;
  assign new_n796_ = b & ~new_n781_;
  assign new_n797_ = ~new_n795_ & ~new_n796_;
  assign new_n798_ = ~m2 & l4;
  assign new_n799_ = ~l2 & new_n785_;
  assign new_n800_ = new_n468_ & new_n797_;
  assign new_n801_ = ~m0 & new_n800_;
  assign new_n802_ = ~new_n604_ & new_n798_;
  assign new_n803_ = ~new_n522_ & new_n802_;
  assign new_n804_ = ~new_n801_ & ~new_n803_;
  assign new_n805_ = ~new_n799_ & new_n804_;
  assign u7 = new_n481_ & new_n805_;
  assign new_n807_ = k & ~l0;
  assign new_n808_ = k0 & new_n807_;
  assign new_n809_ = c & ~new_n781_;
  assign new_n810_ = ~new_n808_ & ~new_n809_;
  assign new_n811_ = ~n2 & l4;
  assign new_n812_ = ~m2 & new_n785_;
  assign new_n813_ = new_n468_ & new_n810_;
  assign new_n814_ = ~m0 & new_n813_;
  assign new_n815_ = ~new_n604_ & new_n811_;
  assign new_n816_ = ~new_n522_ & new_n815_;
  assign new_n817_ = ~new_n814_ & ~new_n816_;
  assign new_n818_ = ~new_n812_ & new_n817_;
  assign v7 = new_n481_ & new_n818_;
  assign new_n820_ = l & ~l0;
  assign new_n821_ = k0 & new_n820_;
  assign new_n822_ = d & ~new_n781_;
  assign new_n823_ = ~new_n821_ & ~new_n822_;
  assign new_n824_ = ~o2 & l4;
  assign new_n825_ = ~n2 & new_n785_;
  assign new_n826_ = new_n468_ & new_n823_;
  assign new_n827_ = ~m0 & new_n826_;
  assign new_n828_ = ~new_n604_ & new_n824_;
  assign new_n829_ = ~new_n522_ & new_n828_;
  assign new_n830_ = ~new_n827_ & ~new_n829_;
  assign new_n831_ = ~new_n825_ & new_n830_;
  assign w7 = new_n481_ & new_n831_;
  assign new_n833_ = m & ~l0;
  assign new_n834_ = k0 & new_n833_;
  assign new_n835_ = e & ~new_n781_;
  assign new_n836_ = ~new_n834_ & ~new_n835_;
  assign new_n837_ = ~p2 & l4;
  assign new_n838_ = ~o2 & new_n785_;
  assign new_n839_ = new_n468_ & new_n836_;
  assign new_n840_ = ~m0 & new_n839_;
  assign new_n841_ = ~new_n604_ & new_n837_;
  assign new_n842_ = ~new_n522_ & new_n841_;
  assign new_n843_ = ~new_n840_ & ~new_n842_;
  assign new_n844_ = ~new_n838_ & new_n843_;
  assign x7 = new_n481_ & new_n844_;
  assign new_n846_ = n & ~l0;
  assign new_n847_ = k0 & new_n846_;
  assign new_n848_ = f & ~new_n781_;
  assign new_n849_ = ~new_n847_ & ~new_n848_;
  assign new_n850_ = ~q2 & l4;
  assign new_n851_ = ~p2 & new_n785_;
  assign new_n852_ = new_n468_ & new_n849_;
  assign new_n853_ = ~m0 & new_n852_;
  assign new_n854_ = ~new_n604_ & new_n850_;
  assign new_n855_ = ~new_n522_ & new_n854_;
  assign new_n856_ = ~new_n853_ & ~new_n855_;
  assign new_n857_ = ~new_n851_ & new_n856_;
  assign y7 = new_n481_ & new_n857_;
  assign new_n859_ = o & ~l0;
  assign new_n860_ = k0 & new_n859_;
  assign new_n861_ = g & ~new_n781_;
  assign new_n862_ = ~new_n860_ & ~new_n861_;
  assign new_n863_ = ~r2 & l4;
  assign new_n864_ = ~q2 & new_n785_;
  assign new_n865_ = new_n468_ & new_n862_;
  assign new_n866_ = ~m0 & new_n865_;
  assign new_n867_ = ~new_n604_ & new_n863_;
  assign new_n868_ = ~new_n522_ & new_n867_;
  assign new_n869_ = ~new_n866_ & ~new_n868_;
  assign new_n870_ = ~new_n864_ & new_n869_;
  assign z7 = new_n481_ & new_n870_;
  assign new_n872_ = p & ~l0;
  assign new_n873_ = k0 & new_n872_;
  assign new_n874_ = h & ~new_n781_;
  assign new_n875_ = ~new_n873_ & ~new_n874_;
  assign new_n876_ = ~s2 & l4;
  assign new_n877_ = ~r2 & new_n785_;
  assign new_n878_ = new_n468_ & new_n875_;
  assign new_n879_ = ~m0 & new_n878_;
  assign new_n880_ = ~new_n604_ & new_n876_;
  assign new_n881_ = ~new_n522_ & new_n880_;
  assign new_n882_ = ~new_n879_ & ~new_n881_;
  assign new_n883_ = ~new_n877_ & new_n882_;
  assign a8 = new_n481_ & new_n883_;
  assign new_n885_ = t2 & l4;
  assign new_n886_ = ~new_n345_ & new_n461_;
  assign new_n887_ = ~m0 & ~n0;
  assign new_n888_ = new_n886_ & new_n887_;
  assign new_n889_ = ~k0 & l0;
  assign new_n890_ = ~new_n781_ & ~new_n889_;
  assign new_n891_ = new_n461_ & new_n890_;
  assign new_n892_ = new_n887_ & new_n891_;
  assign new_n893_ = s2 & ~new_n892_;
  assign new_n894_ = ~l4 & new_n893_;
  assign new_n895_ = new_n604_ & new_n890_;
  assign new_n896_ = i & new_n895_;
  assign new_n897_ = ~new_n894_ & ~new_n896_;
  assign new_n898_ = ~new_n522_ & new_n885_;
  assign new_n899_ = ~s2 & ~new_n898_;
  assign new_n900_ = ~new_n522_ & ~new_n885_;
  assign new_n901_ = ~new_n888_ & ~new_n900_;
  assign new_n902_ = ~new_n899_ & new_n901_;
  assign new_n903_ = new_n897_ & ~new_n902_;
  assign b8 = new_n481_ & ~new_n903_;
  assign new_n905_ = u2 & l4;
  assign new_n906_ = t2 & ~new_n892_;
  assign new_n907_ = ~l4 & new_n906_;
  assign new_n908_ = j & new_n895_;
  assign new_n909_ = ~new_n907_ & ~new_n908_;
  assign new_n910_ = ~new_n522_ & new_n905_;
  assign new_n911_ = ~t2 & ~new_n910_;
  assign new_n912_ = ~new_n522_ & ~new_n905_;
  assign new_n913_ = ~new_n888_ & ~new_n912_;
  assign new_n914_ = ~new_n911_ & new_n913_;
  assign new_n915_ = new_n909_ & ~new_n914_;
  assign c8 = new_n481_ & ~new_n915_;
  assign new_n917_ = v2 & l4;
  assign new_n918_ = u2 & ~new_n892_;
  assign new_n919_ = ~l4 & new_n918_;
  assign new_n920_ = k & new_n895_;
  assign new_n921_ = ~new_n919_ & ~new_n920_;
  assign new_n922_ = ~new_n522_ & new_n917_;
  assign new_n923_ = ~u2 & ~new_n922_;
  assign new_n924_ = ~new_n522_ & ~new_n917_;
  assign new_n925_ = ~new_n888_ & ~new_n924_;
  assign new_n926_ = ~new_n923_ & new_n925_;
  assign new_n927_ = new_n921_ & ~new_n926_;
  assign d8 = new_n481_ & ~new_n927_;
  assign new_n929_ = w2 & l4;
  assign new_n930_ = v2 & ~new_n892_;
  assign new_n931_ = ~l4 & new_n930_;
  assign new_n932_ = l & new_n895_;
  assign new_n933_ = ~new_n931_ & ~new_n932_;
  assign new_n934_ = ~new_n522_ & new_n929_;
  assign new_n935_ = ~v2 & ~new_n934_;
  assign new_n936_ = ~new_n522_ & ~new_n929_;
  assign new_n937_ = ~new_n888_ & ~new_n936_;
  assign new_n938_ = ~new_n935_ & new_n937_;
  assign new_n939_ = new_n933_ & ~new_n938_;
  assign e8 = new_n481_ & ~new_n939_;
  assign new_n941_ = x2 & l4;
  assign new_n942_ = w2 & ~new_n892_;
  assign new_n943_ = ~l4 & new_n942_;
  assign new_n944_ = m & new_n895_;
  assign new_n945_ = ~new_n943_ & ~new_n944_;
  assign new_n946_ = ~new_n522_ & new_n941_;
  assign new_n947_ = ~w2 & ~new_n946_;
  assign new_n948_ = ~new_n522_ & ~new_n941_;
  assign new_n949_ = ~new_n888_ & ~new_n948_;
  assign new_n950_ = ~new_n947_ & new_n949_;
  assign new_n951_ = new_n945_ & ~new_n950_;
  assign f8 = new_n481_ & ~new_n951_;
  assign new_n953_ = y2 & l4;
  assign new_n954_ = x2 & ~new_n892_;
  assign new_n955_ = ~l4 & new_n954_;
  assign new_n956_ = n & new_n895_;
  assign new_n957_ = ~new_n955_ & ~new_n956_;
  assign new_n958_ = ~new_n522_ & new_n953_;
  assign new_n959_ = ~x2 & ~new_n958_;
  assign new_n960_ = ~new_n522_ & ~new_n953_;
  assign new_n961_ = ~new_n888_ & ~new_n960_;
  assign new_n962_ = ~new_n959_ & new_n961_;
  assign new_n963_ = new_n957_ & ~new_n962_;
  assign g8 = new_n481_ & ~new_n963_;
  assign new_n965_ = z2 & l4;
  assign new_n966_ = y2 & ~new_n892_;
  assign new_n967_ = ~l4 & new_n966_;
  assign new_n968_ = o & new_n895_;
  assign new_n969_ = ~new_n967_ & ~new_n968_;
  assign new_n970_ = ~new_n522_ & new_n965_;
  assign new_n971_ = ~y2 & ~new_n970_;
  assign new_n972_ = ~new_n522_ & ~new_n965_;
  assign new_n973_ = ~new_n888_ & ~new_n972_;
  assign new_n974_ = ~new_n971_ & new_n973_;
  assign new_n975_ = new_n969_ & ~new_n974_;
  assign h8 = new_n481_ & ~new_n975_;
  assign new_n977_ = p & new_n887_;
  assign new_n978_ = ~q0 & new_n461_;
  assign new_n979_ = o0 & new_n978_;
  assign new_n980_ = ~q0 & z2;
  assign new_n981_ = new_n468_ & new_n890_;
  assign new_n982_ = ~m0 & new_n981_;
  assign new_n983_ = ~new_n524_ & ~new_n982_;
  assign new_n984_ = new_n980_ & new_n983_;
  assign new_n985_ = o0 & new_n984_;
  assign new_n986_ = new_n890_ & new_n979_;
  assign new_n987_ = new_n977_ & new_n986_;
  assign i8 = new_n985_ | new_n987_;
  assign new_n989_ = ~new_n440_ & new_n446_;
  assign new_n990_ = new_n451_ & new_n989_;
  assign new_n991_ = ~q0 & ~new_n990_;
  assign new_n992_ = o0 & new_n991_;
  assign new_n993_ = f4 & ~g4;
  assign new_n994_ = e4 & new_n993_;
  assign new_n995_ = ~h4 & new_n994_;
  assign new_n996_ = b3 & k4;
  assign new_n997_ = ~new_n995_ & new_n996_;
  assign new_n998_ = new_n458_ & new_n460_;
  assign new_n999_ = ~j1 & new_n460_;
  assign new_n1000_ = k1 & l1;
  assign new_n1001_ = j1 & ~new_n460_;
  assign new_n1002_ = ~new_n1000_ & ~new_n1001_;
  assign new_n1003_ = ~h1 & new_n999_;
  assign new_n1004_ = ~i1 & new_n1003_;
  assign new_n1005_ = new_n1002_ & ~new_n1004_;
  assign new_n1006_ = h1 & ~new_n998_;
  assign new_n1007_ = i1 & ~new_n999_;
  assign new_n1008_ = ~new_n1006_ & ~new_n1007_;
  assign new_n1009_ = new_n1005_ & new_n1008_;
  assign new_n1010_ = ~q0 & a3;
  assign new_n1011_ = j1 & k1;
  assign new_n1012_ = ~new_n990_ & ~new_n1011_;
  assign new_n1013_ = ~new_n461_ & new_n1012_;
  assign new_n1014_ = j1 & l1;
  assign new_n1015_ = new_n1013_ & ~new_n1014_;
  assign new_n1016_ = ~new_n995_ & new_n1015_;
  assign new_n1017_ = k4 & ~new_n1000_;
  assign new_n1018_ = new_n1016_ & new_n1017_;
  assign new_n1019_ = new_n1008_ & new_n1018_;
  assign new_n1020_ = new_n1010_ & ~new_n1019_;
  assign new_n1021_ = o0 & new_n1020_;
  assign new_n1022_ = new_n997_ & new_n1009_;
  assign new_n1023_ = new_n992_ & new_n1022_;
  assign j8 = new_n1021_ | new_n1023_;
  assign new_n1025_ = c3 & k4;
  assign new_n1026_ = ~new_n995_ & new_n1025_;
  assign new_n1027_ = ~q0 & b3;
  assign new_n1028_ = ~new_n1019_ & new_n1027_;
  assign new_n1029_ = o0 & new_n1028_;
  assign new_n1030_ = new_n1009_ & new_n1026_;
  assign new_n1031_ = new_n992_ & new_n1030_;
  assign k8 = new_n1029_ | new_n1031_;
  assign new_n1033_ = d3 & k4;
  assign new_n1034_ = ~new_n995_ & new_n1033_;
  assign new_n1035_ = ~q0 & c3;
  assign new_n1036_ = ~new_n1019_ & new_n1035_;
  assign new_n1037_ = o0 & new_n1036_;
  assign new_n1038_ = new_n1009_ & new_n1034_;
  assign new_n1039_ = new_n992_ & new_n1038_;
  assign l8 = new_n1037_ | new_n1039_;
  assign new_n1041_ = e3 & k4;
  assign new_n1042_ = ~new_n995_ & new_n1041_;
  assign new_n1043_ = ~q0 & d3;
  assign new_n1044_ = ~new_n1019_ & new_n1043_;
  assign new_n1045_ = o0 & new_n1044_;
  assign new_n1046_ = new_n1009_ & new_n1042_;
  assign new_n1047_ = new_n992_ & new_n1046_;
  assign m8 = new_n1045_ | new_n1047_;
  assign new_n1049_ = f3 & k4;
  assign new_n1050_ = ~new_n995_ & new_n1049_;
  assign new_n1051_ = ~q0 & e3;
  assign new_n1052_ = ~new_n1019_ & new_n1051_;
  assign new_n1053_ = o0 & new_n1052_;
  assign new_n1054_ = new_n1009_ & new_n1050_;
  assign new_n1055_ = new_n992_ & new_n1054_;
  assign n8 = new_n1053_ | new_n1055_;
  assign new_n1057_ = g3 & k4;
  assign new_n1058_ = ~new_n995_ & new_n1057_;
  assign new_n1059_ = ~q0 & f3;
  assign new_n1060_ = ~new_n1019_ & new_n1059_;
  assign new_n1061_ = o0 & new_n1060_;
  assign new_n1062_ = new_n1009_ & new_n1058_;
  assign new_n1063_ = new_n992_ & new_n1062_;
  assign o8 = new_n1061_ | new_n1063_;
  assign new_n1065_ = h3 & k4;
  assign new_n1066_ = ~new_n995_ & new_n1065_;
  assign new_n1067_ = ~q0 & g3;
  assign new_n1068_ = ~new_n1019_ & new_n1067_;
  assign new_n1069_ = o0 & new_n1068_;
  assign new_n1070_ = new_n1009_ & new_n1066_;
  assign new_n1071_ = new_n992_ & new_n1070_;
  assign p8 = new_n1069_ | new_n1071_;
  assign new_n1073_ = i3 & k4;
  assign new_n1074_ = ~new_n995_ & new_n1073_;
  assign new_n1075_ = ~q0 & h3;
  assign new_n1076_ = ~new_n1019_ & new_n1075_;
  assign new_n1077_ = o0 & new_n1076_;
  assign new_n1078_ = new_n1009_ & new_n1074_;
  assign new_n1079_ = new_n992_ & new_n1078_;
  assign q8 = new_n1077_ | new_n1079_;
  assign new_n1081_ = j3 & k4;
  assign new_n1082_ = ~new_n995_ & new_n1081_;
  assign new_n1083_ = ~q0 & i3;
  assign new_n1084_ = ~new_n1019_ & new_n1083_;
  assign new_n1085_ = o0 & new_n1084_;
  assign new_n1086_ = new_n1009_ & new_n1082_;
  assign new_n1087_ = new_n992_ & new_n1086_;
  assign r8 = new_n1085_ | new_n1087_;
  assign new_n1089_ = k3 & k4;
  assign new_n1090_ = ~new_n995_ & new_n1089_;
  assign new_n1091_ = ~q0 & j3;
  assign new_n1092_ = ~new_n1019_ & new_n1091_;
  assign new_n1093_ = o0 & new_n1092_;
  assign new_n1094_ = new_n1009_ & new_n1090_;
  assign new_n1095_ = new_n992_ & new_n1094_;
  assign s8 = new_n1093_ | new_n1095_;
  assign new_n1097_ = l3 & k4;
  assign new_n1098_ = ~new_n995_ & new_n1097_;
  assign new_n1099_ = ~q0 & k3;
  assign new_n1100_ = ~new_n1019_ & new_n1099_;
  assign new_n1101_ = o0 & new_n1100_;
  assign new_n1102_ = new_n1009_ & new_n1098_;
  assign new_n1103_ = new_n992_ & new_n1102_;
  assign t8 = new_n1101_ | new_n1103_;
  assign new_n1105_ = m3 & k4;
  assign new_n1106_ = ~new_n995_ & new_n1105_;
  assign new_n1107_ = ~q0 & l3;
  assign new_n1108_ = ~new_n1019_ & new_n1107_;
  assign new_n1109_ = o0 & new_n1108_;
  assign new_n1110_ = new_n1009_ & new_n1106_;
  assign new_n1111_ = new_n992_ & new_n1110_;
  assign u8 = new_n1109_ | new_n1111_;
  assign new_n1113_ = n3 & k4;
  assign new_n1114_ = ~new_n995_ & new_n1113_;
  assign new_n1115_ = ~q0 & m3;
  assign new_n1116_ = ~new_n1019_ & new_n1115_;
  assign new_n1117_ = o0 & new_n1116_;
  assign new_n1118_ = new_n1009_ & new_n1114_;
  assign new_n1119_ = new_n992_ & new_n1118_;
  assign v8 = new_n1117_ | new_n1119_;
  assign new_n1121_ = o3 & k4;
  assign new_n1122_ = ~new_n995_ & new_n1121_;
  assign new_n1123_ = ~q0 & n3;
  assign new_n1124_ = ~new_n1019_ & new_n1123_;
  assign new_n1125_ = o0 & new_n1124_;
  assign new_n1126_ = new_n1009_ & new_n1122_;
  assign new_n1127_ = new_n992_ & new_n1126_;
  assign w8 = new_n1125_ | new_n1127_;
  assign new_n1129_ = p3 & k4;
  assign new_n1130_ = ~new_n995_ & new_n1129_;
  assign new_n1131_ = ~q0 & o3;
  assign new_n1132_ = ~new_n1019_ & new_n1131_;
  assign new_n1133_ = o0 & new_n1132_;
  assign new_n1134_ = new_n1009_ & new_n1130_;
  assign new_n1135_ = new_n992_ & new_n1134_;
  assign x8 = new_n1133_ | new_n1135_;
  assign new_n1137_ = q3 & k4;
  assign new_n1138_ = ~new_n995_ & new_n1137_;
  assign new_n1139_ = ~q0 & p3;
  assign new_n1140_ = ~new_n1019_ & new_n1139_;
  assign new_n1141_ = o0 & new_n1140_;
  assign new_n1142_ = new_n1009_ & new_n1138_;
  assign new_n1143_ = new_n992_ & new_n1142_;
  assign y8 = new_n1141_ | new_n1143_;
  assign new_n1145_ = r3 & k4;
  assign new_n1146_ = ~new_n995_ & new_n1145_;
  assign new_n1147_ = ~q0 & q3;
  assign new_n1148_ = ~new_n1019_ & new_n1147_;
  assign new_n1149_ = o0 & new_n1148_;
  assign new_n1150_ = new_n1009_ & new_n1146_;
  assign new_n1151_ = new_n992_ & new_n1150_;
  assign z8 = new_n1149_ | new_n1151_;
  assign new_n1153_ = s3 & k4;
  assign new_n1154_ = ~new_n995_ & new_n1153_;
  assign new_n1155_ = ~q0 & r3;
  assign new_n1156_ = ~new_n1019_ & new_n1155_;
  assign new_n1157_ = o0 & new_n1156_;
  assign new_n1158_ = new_n1009_ & new_n1154_;
  assign new_n1159_ = new_n992_ & new_n1158_;
  assign a9 = new_n1157_ | new_n1159_;
  assign new_n1161_ = t3 & k4;
  assign new_n1162_ = ~new_n995_ & new_n1161_;
  assign new_n1163_ = ~q0 & s3;
  assign new_n1164_ = ~new_n1019_ & new_n1163_;
  assign new_n1165_ = o0 & new_n1164_;
  assign new_n1166_ = new_n1009_ & new_n1162_;
  assign new_n1167_ = new_n992_ & new_n1166_;
  assign b9 = new_n1165_ | new_n1167_;
  assign new_n1169_ = u3 & k4;
  assign new_n1170_ = ~new_n995_ & new_n1169_;
  assign new_n1171_ = ~q0 & t3;
  assign new_n1172_ = ~new_n1019_ & new_n1171_;
  assign new_n1173_ = o0 & new_n1172_;
  assign new_n1174_ = new_n1009_ & new_n1170_;
  assign new_n1175_ = new_n992_ & new_n1174_;
  assign c9 = new_n1173_ | new_n1175_;
  assign new_n1177_ = v3 & k4;
  assign new_n1178_ = ~new_n995_ & new_n1177_;
  assign new_n1179_ = ~q0 & u3;
  assign new_n1180_ = ~new_n1019_ & new_n1179_;
  assign new_n1181_ = o0 & new_n1180_;
  assign new_n1182_ = new_n1009_ & new_n1178_;
  assign new_n1183_ = new_n992_ & new_n1182_;
  assign d9 = new_n1181_ | new_n1183_;
  assign new_n1185_ = w3 & k4;
  assign new_n1186_ = ~new_n995_ & new_n1185_;
  assign new_n1187_ = ~q0 & v3;
  assign new_n1188_ = ~new_n1019_ & new_n1187_;
  assign new_n1189_ = o0 & new_n1188_;
  assign new_n1190_ = new_n1009_ & new_n1186_;
  assign new_n1191_ = new_n992_ & new_n1190_;
  assign e9 = new_n1189_ | new_n1191_;
  assign new_n1193_ = k4 & ~new_n995_;
  assign new_n1194_ = ~new_n990_ & new_n1193_;
  assign new_n1195_ = h1 & ~i1;
  assign new_n1196_ = ~k1 & l1;
  assign new_n1197_ = ~j1 & k1;
  assign new_n1198_ = v0 & new_n1197_;
  assign new_n1199_ = ~l1 & new_n1198_;
  assign new_n1200_ = u0 & new_n460_;
  assign new_n1201_ = ~j1 & new_n1196_;
  assign new_n1202_ = w0 & new_n1201_;
  assign new_n1203_ = ~new_n1200_ & ~new_n1202_;
  assign new_n1204_ = w0 & new_n1196_;
  assign new_n1205_ = ~j1 & ~new_n1204_;
  assign new_n1206_ = ~new_n1203_ & ~new_n1205_;
  assign new_n1207_ = ~new_n1199_ & ~new_n1206_;
  assign new_n1208_ = t0 & new_n999_;
  assign new_n1209_ = i1 & new_n1208_;
  assign new_n1210_ = ~i1 & ~new_n1207_;
  assign new_n1211_ = ~new_n1209_ & ~new_n1210_;
  assign new_n1212_ = ~h1 & ~new_n1211_;
  assign new_n1213_ = new_n999_ & new_n1195_;
  assign new_n1214_ = s0 & new_n1213_;
  assign new_n1215_ = ~new_n1212_ & ~new_n1214_;
  assign new_n1216_ = ~q0 & w3;
  assign new_n1217_ = ~new_n1001_ & ~new_n1004_;
  assign new_n1218_ = ~new_n1000_ & new_n1217_;
  assign new_n1219_ = ~new_n990_ & new_n1218_;
  assign new_n1220_ = new_n1193_ & new_n1219_;
  assign new_n1221_ = new_n1008_ & new_n1220_;
  assign new_n1222_ = new_n1216_ & ~new_n1221_;
  assign new_n1223_ = o0 & new_n1222_;
  assign new_n1224_ = new_n1194_ & ~new_n1215_;
  assign new_n1225_ = new_n481_ & new_n1224_;
  assign f9 = new_n1223_ | new_n1225_;
  assign new_n1227_ = ~q0 & ~new_n468_;
  assign new_n1228_ = o0 & new_n1227_;
  assign new_n1229_ = x3 & ~new_n522_;
  assign new_n1230_ = l4 & new_n1229_;
  assign new_n1231_ = new_n1228_ & ~new_n1230_;
  assign new_n1232_ = ~x3 & ~new_n524_;
  assign g9 = new_n1231_ & ~new_n1232_;
  assign new_n1234_ = ~x3 & l4;
  assign new_n1235_ = ~new_n522_ & new_n1234_;
  assign new_n1236_ = ~x3 & ~y3;
  assign new_n1237_ = ~new_n522_ & new_n1236_;
  assign new_n1238_ = l4 & new_n1237_;
  assign new_n1239_ = ~new_n468_ & ~new_n1238_;
  assign new_n1240_ = ~q0 & new_n1239_;
  assign new_n1241_ = y3 & ~new_n1235_;
  assign new_n1242_ = o0 & ~new_n1241_;
  assign h9 = ~new_n1240_ | ~new_n1242_;
  assign new_n1244_ = y3 & l4;
  assign new_n1245_ = ~x3 & ~new_n522_;
  assign new_n1246_ = new_n1244_ & new_n1245_;
  assign new_n1247_ = new_n520_ & ~new_n522_;
  assign new_n1248_ = ~z3 & l4;
  assign new_n1249_ = new_n1247_ & new_n1248_;
  assign new_n1250_ = ~new_n468_ & ~new_n1249_;
  assign new_n1251_ = ~q0 & new_n1250_;
  assign new_n1252_ = z3 & ~new_n1246_;
  assign new_n1253_ = o0 & ~new_n1252_;
  assign i9 = ~new_n1251_ | ~new_n1253_;
  assign new_n1255_ = ~a4 & l4;
  assign new_n1256_ = z3 & new_n1255_;
  assign new_n1257_ = z3 & l4;
  assign new_n1258_ = y3 & new_n1257_;
  assign new_n1259_ = new_n1245_ & new_n1258_;
  assign new_n1260_ = n0 & new_n461_;
  assign new_n1261_ = ~new_n461_ & new_n1259_;
  assign new_n1262_ = ~new_n1260_ & ~new_n1261_;
  assign new_n1263_ = a4 & ~new_n461_;
  assign new_n1264_ = ~a4 & ~new_n461_;
  assign new_n1265_ = ~m0 & ~new_n890_;
  assign new_n1266_ = ~new_n1264_ & ~new_n1265_;
  assign new_n1267_ = ~new_n1263_ & ~new_n1266_;
  assign new_n1268_ = new_n1262_ & ~new_n1267_;
  assign new_n1269_ = ~new_n468_ & new_n1256_;
  assign new_n1270_ = new_n1247_ & new_n1269_;
  assign new_n1271_ = n0 & ~new_n1259_;
  assign new_n1272_ = a4 & new_n1271_;
  assign new_n1273_ = ~new_n1270_ & ~new_n1272_;
  assign new_n1274_ = ~new_n1268_ & new_n1273_;
  assign j9 = new_n481_ & ~new_n1274_;
  assign new_n1276_ = ~b4 & l4;
  assign new_n1277_ = ~a4 & new_n1276_;
  assign new_n1278_ = o0 & new_n405_;
  assign new_n1279_ = new_n1277_ & new_n1278_;
  assign new_n1280_ = ~q0 & new_n1245_;
  assign new_n1281_ = ~q0 & b4;
  assign new_n1282_ = new_n520_ & new_n1256_;
  assign new_n1283_ = ~new_n522_ & new_n1282_;
  assign new_n1284_ = ~new_n468_ & ~new_n1283_;
  assign new_n1285_ = ~n0 & o0;
  assign new_n1286_ = m0 & new_n1285_;
  assign new_n1287_ = new_n978_ & new_n1286_;
  assign new_n1288_ = new_n1281_ & new_n1284_;
  assign new_n1289_ = o0 & new_n1288_;
  assign new_n1290_ = ~new_n468_ & new_n1280_;
  assign new_n1291_ = new_n1279_ & new_n1290_;
  assign new_n1292_ = ~new_n1289_ & ~new_n1291_;
  assign k9 = new_n1287_ | ~new_n1292_;
  assign new_n1294_ = y3 & new_n430_;
  assign new_n1295_ = ~c4 & l4;
  assign new_n1296_ = ~b4 & new_n1295_;
  assign new_n1297_ = o0 & new_n1294_;
  assign new_n1298_ = new_n1296_ & new_n1297_;
  assign new_n1299_ = ~q0 & c4;
  assign new_n1300_ = ~x3 & new_n405_;
  assign new_n1301_ = new_n1277_ & new_n1300_;
  assign new_n1302_ = ~new_n522_ & new_n1301_;
  assign new_n1303_ = ~new_n468_ & ~new_n1302_;
  assign new_n1304_ = ~m0 & new_n1285_;
  assign new_n1305_ = new_n978_ & new_n1304_;
  assign new_n1306_ = new_n1299_ & new_n1303_;
  assign new_n1307_ = o0 & new_n1306_;
  assign new_n1308_ = new_n1290_ & new_n1298_;
  assign new_n1309_ = ~new_n1307_ & ~new_n1308_;
  assign l9 = new_n1305_ | ~new_n1309_;
  assign new_n1311_ = ~q0 & ~g1;
  assign new_n1312_ = d4 & k4;
  assign new_n1313_ = ~d4 & ~new_n1194_;
  assign new_n1314_ = ~new_n990_ & new_n1312_;
  assign new_n1315_ = ~new_n995_ & new_n1314_;
  assign new_n1316_ = ~new_n1313_ & ~new_n1315_;
  assign new_n1317_ = new_n1311_ & new_n1316_;
  assign new_n1318_ = ~n0 & new_n978_;
  assign new_n1319_ = ~new_n1317_ & ~new_n1318_;
  assign m9 = o0 & ~new_n1319_;
  assign new_n1321_ = ~d4 & k4;
  assign new_n1322_ = ~new_n990_ & ~new_n995_;
  assign new_n1323_ = new_n1321_ & new_n1322_;
  assign new_n1324_ = ~e4 & k4;
  assign new_n1325_ = ~d4 & new_n1324_;
  assign new_n1326_ = ~new_n990_ & new_n1325_;
  assign new_n1327_ = ~new_n995_ & new_n1326_;
  assign new_n1328_ = ~new_n468_ & ~new_n1327_;
  assign new_n1329_ = new_n1311_ & new_n1328_;
  assign new_n1330_ = e4 & ~new_n1323_;
  assign new_n1331_ = o0 & ~new_n1330_;
  assign n9 = ~new_n1329_ | ~new_n1331_;
  assign new_n1333_ = e4 & k4;
  assign new_n1334_ = ~d4 & new_n1333_;
  assign new_n1335_ = new_n1322_ & new_n1334_;
  assign new_n1336_ = ~d4 & ~new_n995_;
  assign new_n1337_ = ~f4 & k4;
  assign new_n1338_ = e4 & new_n1337_;
  assign new_n1339_ = new_n1336_ & new_n1338_;
  assign new_n1340_ = ~new_n990_ & new_n1339_;
  assign new_n1341_ = ~new_n468_ & ~new_n1340_;
  assign new_n1342_ = new_n1311_ & new_n1341_;
  assign new_n1343_ = f4 & ~new_n1335_;
  assign new_n1344_ = o0 & ~new_n1343_;
  assign o9 = ~new_n1342_ | ~new_n1344_;
  assign new_n1346_ = ~d4 & e4;
  assign new_n1347_ = ~g1 & new_n1346_;
  assign new_n1348_ = ~g4 & k4;
  assign new_n1349_ = f4 & new_n1348_;
  assign new_n1350_ = o0 & new_n1347_;
  assign new_n1351_ = new_n1349_ & new_n1350_;
  assign new_n1352_ = ~q0 & new_n1322_;
  assign new_n1353_ = ~g1 & g4;
  assign new_n1354_ = ~q0 & new_n1353_;
  assign new_n1355_ = f4 & k4;
  assign new_n1356_ = e4 & new_n1355_;
  assign new_n1357_ = new_n1336_ & new_n1356_;
  assign new_n1358_ = ~new_n990_ & new_n1357_;
  assign new_n1359_ = ~new_n468_ & ~new_n1358_;
  assign new_n1360_ = m0 & ~new_n890_;
  assign new_n1361_ = ~n0 & ~new_n1360_;
  assign new_n1362_ = o0 & new_n1361_;
  assign new_n1363_ = new_n978_ & new_n1362_;
  assign new_n1364_ = new_n1354_ & new_n1359_;
  assign new_n1365_ = o0 & new_n1364_;
  assign new_n1366_ = ~new_n468_ & new_n1352_;
  assign new_n1367_ = new_n1351_ & new_n1366_;
  assign new_n1368_ = ~new_n1365_ & ~new_n1367_;
  assign p9 = new_n1363_ | ~new_n1368_;
  assign new_n1370_ = ~g1 & ~new_n995_;
  assign new_n1371_ = ~d4 & new_n435_;
  assign new_n1372_ = ~h4 & k4;
  assign new_n1373_ = ~g4 & new_n1372_;
  assign new_n1374_ = new_n1370_ & new_n1371_;
  assign new_n1375_ = new_n1373_ & new_n1374_;
  assign new_n1376_ = ~g1 & h4;
  assign new_n1377_ = ~q0 & new_n1376_;
  assign new_n1378_ = ~new_n995_ & new_n1346_;
  assign new_n1379_ = new_n1349_ & new_n1378_;
  assign new_n1380_ = ~new_n990_ & new_n1379_;
  assign new_n1381_ = ~new_n468_ & ~new_n1380_;
  assign new_n1382_ = new_n1377_ & new_n1381_;
  assign new_n1383_ = o0 & new_n1382_;
  assign new_n1384_ = ~new_n468_ & new_n992_;
  assign new_n1385_ = new_n1375_ & new_n1384_;
  assign new_n1386_ = ~new_n1383_ & ~new_n1385_;
  assign q9 = new_n1287_ | ~new_n1386_;
  assign new_n1388_ = ~q0 & ~new_n522_;
  assign new_n1389_ = o0 & new_n1388_;
  assign new_n1390_ = n1 & i4;
  assign new_n1391_ = new_n1389_ & ~new_n1390_;
  assign new_n1392_ = ~n1 & ~i4;
  assign new_n1393_ = new_n1391_ & ~new_n1392_;
  assign r9 = l4 & new_n1393_;
  assign new_n1395_ = k4 & n4;
  assign new_n1396_ = ~j4 & new_n1395_;
  assign new_n1397_ = new_n481_ & new_n1396_;
  assign new_n1398_ = ~new_n990_ & new_n1370_;
  assign new_n1399_ = ~g1 & j4;
  assign new_n1400_ = ~q0 & new_n1399_;
  assign new_n1401_ = ~v0 & ~l1;
  assign new_n1402_ = w0 & l1;
  assign new_n1403_ = ~k1 & ~new_n1402_;
  assign new_n1404_ = ~new_n1401_ & ~new_n1403_;
  assign new_n1405_ = s0 & ~i1;
  assign new_n1406_ = new_n999_ & new_n1405_;
  assign new_n1407_ = ~i1 & new_n460_;
  assign new_n1408_ = t0 & ~j1;
  assign new_n1409_ = new_n460_ & new_n1408_;
  assign new_n1410_ = ~new_n995_ & ~new_n1001_;
  assign new_n1411_ = ~new_n990_ & ~new_n1000_;
  assign new_n1412_ = new_n1410_ & new_n1411_;
  assign new_n1413_ = new_n1395_ & new_n1412_;
  assign new_n1414_ = ~u0 & new_n1407_;
  assign new_n1415_ = ~h1 & new_n1414_;
  assign new_n1416_ = i1 & ~new_n1409_;
  assign new_n1417_ = ~new_n1415_ & ~new_n1416_;
  assign new_n1418_ = new_n1413_ & new_n1417_;
  assign new_n1419_ = h1 & new_n1406_;
  assign new_n1420_ = h1 & ~new_n1406_;
  assign new_n1421_ = new_n458_ & ~new_n1404_;
  assign new_n1422_ = ~new_n1420_ & ~new_n1421_;
  assign new_n1423_ = ~new_n1419_ & ~new_n1422_;
  assign new_n1424_ = new_n1418_ & ~new_n1423_;
  assign new_n1425_ = new_n1400_ & ~new_n1424_;
  assign new_n1426_ = o0 & new_n1425_;
  assign new_n1427_ = ~new_n1215_ & new_n1398_;
  assign new_n1428_ = new_n1397_ & new_n1427_;
  assign s9 = new_n1426_ | new_n1428_;
  assign new_n1430_ = ~q0 & m1;
  assign new_n1431_ = o0 & new_n1430_;
  assign new_n1432_ = new_n1294_ & new_n1431_;
  assign t9 = new_n406_ & new_n1432_;
  assign u9 = m1 & new_n1389_;
  assign new_n1435_ = ~new_n440_ & ~new_n445_;
  assign new_n1436_ = ~new_n995_ & new_n1435_;
  assign new_n1437_ = ~new_n444_ & ~new_n450_;
  assign new_n1438_ = new_n1436_ & new_n1437_;
  assign new_n1439_ = n4 & ~new_n449_;
  assign new_n1440_ = new_n1438_ & new_n1439_;
  assign new_n1441_ = new_n990_ & ~new_n1440_;
  assign new_n1442_ = ~q0 & ~new_n1441_;
  assign new_n1443_ = o0 & new_n1442_;
  assign new_n1444_ = ~new_n453_ & ~new_n1440_;
  assign v9 = new_n1443_ & ~new_n1444_;
  assign w9 = k4 & new_n992_;
  assign o4 = ~g1;
  assign h6 = ~h1;
  assign i6 = ~i1;
  assign j6 = ~j1;
  assign k6 = ~k1;
  assign l6 = ~l1;
  assign t4 = u3;
  assign u4 = v3;
  assign m5 = m4;
  assign t5 = s5;
  assign u5 = s5;
  assign v5 = s5;
  assign w5 = s5;
  assign m6 = k4;
endmodule

