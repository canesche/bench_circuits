// Benchmark "testing" written by ABC on Thu Oct  8 22:16:59 2020

module testing ( 
    A743, A742, A741, A740, A739, A738, A676, A675, A674, A673, A672, A671,
    A609, A608, A607, A606, A605, A604, A542, A541, A540, A539, A538, A537,
    A475, A474, A473, A472, A471, A470, A403, A404, A405, A406, A407, A408,
    A347, A346, A345, A344, A343, A342, A280, A279, A278, A277, A276, A275,
    A213, A212, A211, A210, A209, A208, A146, A145, A144, A143, A142, A141,
    A79, A78, A77, A76, A75, A74, A7, A8, A9, A10, A11, A12  );
  input  A743, A742, A741, A740, A739, A738, A676, A675, A674, A673,
    A672, A671, A609, A608, A607, A606, A605, A604, A542, A541, A540, A539,
    A538, A537, A475, A474, A473, A472, A471, A470, A403, A404, A405, A406,
    A407, A408;
  output A347, A346, A345, A344, A343, A342, A280, A279, A278, A277, A276,
    A275, A213, A212, A211, A210, A209, A208, A146, A145, A144, A143, A142,
    A141, A79, A78, A77, A76, A75, A74, A7, A8, A9, A10, A11, A12;
  wire new_A469_, new_A468_, new_A467_, new_A466_, new_A465_, new_A464_,
    new_A463_, new_A462_, new_A461_, new_A460_, new_A459_, new_A458_,
    new_A457_, new_A456_, new_A455_, new_A454_, new_A453_, new_A452_,
    new_A451_, new_A450_, new_A449_, new_A448_, new_A447_, new_A446_,
    new_A445_, new_A444_, new_A443_, new_A442_, new_A441_, new_A440_,
    new_A439_, new_A438_, new_A437_, new_A436_, new_A435_, new_A434_,
    new_A433_, new_A432_, new_A431_, new_A430_, new_A429_, new_A428_,
    new_A427_, new_A426_, new_A425_, new_A424_, new_A423_, new_A422_,
    new_A421_, new_A420_, new_A419_, new_A418_, new_A417_, new_A416_,
    new_A415_, new_A414_, new_A413_, new_A412_, new_A411_, new_A410_,
    new_A409_, new_A476_, new_A477_, new_A478_, new_A479_, new_A480_,
    new_A481_, new_A482_, new_A483_, new_A484_, new_A485_, new_A486_,
    new_A487_, new_A488_, new_A489_, new_A490_, new_A491_, new_A492_,
    new_A493_, new_A494_, new_A495_, new_A496_, new_A497_, new_A498_,
    new_A499_, new_A500_, new_A501_, new_A502_, new_A503_, new_A504_,
    new_A505_, new_A506_, new_A507_, new_A508_, new_A509_, new_A510_,
    new_A511_, new_A512_, new_A513_, new_A514_, new_A515_, new_A516_,
    new_A517_, new_A518_, new_A519_, new_A520_, new_A521_, new_A522_,
    new_A523_, new_A524_, new_A525_, new_A526_, new_A527_, new_A528_,
    new_A529_, new_A530_, new_A531_, new_A532_, new_A533_, new_A534_,
    new_A535_, new_A536_, new_A543_, new_A544_, new_A545_, new_A546_,
    new_A547_, new_A548_, new_A549_, new_A550_, new_A551_, new_A552_,
    new_A553_, new_A554_, new_A555_, new_A556_, new_A557_, new_A558_,
    new_A559_, new_A560_, new_A561_, new_A562_, new_A563_, new_A564_,
    new_A565_, new_A566_, new_A567_, new_A568_, new_A569_, new_A570_,
    new_A571_, new_A572_, new_A573_, new_A574_, new_A575_, new_A576_,
    new_A577_, new_A578_, new_A579_, new_A580_, new_A581_, new_A582_,
    new_A583_, new_A584_, new_A585_, new_A586_, new_A587_, new_A588_,
    new_A589_, new_A590_, new_A591_, new_A592_, new_A593_, new_A594_,
    new_A595_, new_A596_, new_A597_, new_A598_, new_A599_, new_A600_,
    new_A601_, new_A602_, new_A603_, new_A610_, new_A611_, new_A612_,
    new_A613_, new_A614_, new_A615_, new_A616_, new_A617_, new_A618_,
    new_A619_, new_A620_, new_A621_, new_A622_, new_A623_, new_A624_,
    new_A625_, new_A626_, new_A627_, new_A628_, new_A629_, new_A630_,
    new_A631_, new_A632_, new_A633_, new_A634_, new_A635_, new_A636_,
    new_A637_, new_A638_, new_A639_, new_A640_, new_A641_, new_A642_,
    new_A643_, new_A644_, new_A645_, new_A646_, new_A647_, new_A648_,
    new_A649_, new_A650_, new_A651_, new_A652_, new_A653_, new_A654_,
    new_A655_, new_A656_, new_A657_, new_A658_, new_A659_, new_A660_,
    new_A661_, new_A662_, new_A663_, new_A664_, new_A665_, new_A666_,
    new_A667_, new_A668_, new_A669_, new_A670_, new_A677_, new_A678_,
    new_A679_, new_A680_, new_A681_, new_A682_, new_A683_, new_A684_,
    new_A685_, new_A686_, new_A687_, new_A688_, new_A689_, new_A690_,
    new_A691_, new_A692_, new_A693_, new_A694_, new_A695_, new_A696_,
    new_A697_, new_A698_, new_A699_, new_A700_, new_A701_, new_A702_,
    new_A703_, new_A704_, new_A705_, new_A706_, new_A707_, new_A708_,
    new_A709_, new_A710_, new_A711_, new_A712_, new_A713_, new_A714_,
    new_A715_, new_A716_, new_A717_, new_A718_, new_A719_, new_A720_,
    new_A721_, new_A722_, new_A723_, new_A724_, new_A725_, new_A726_,
    new_A727_, new_A728_, new_A729_, new_A730_, new_A731_, new_A732_,
    new_A733_, new_A734_, new_A735_, new_A736_, new_A737_, new_A744_,
    new_A745_, new_A746_, new_A747_, new_A748_, new_A749_, new_A750_,
    new_A751_, new_A752_, new_A753_, new_A754_, new_A755_, new_A756_,
    new_A757_, new_A758_, new_A759_, new_A760_, new_A761_, new_A762_,
    new_A763_, new_A764_, new_A765_, new_A766_, new_A767_, new_A768_,
    new_A769_, new_A770_, new_A771_, new_A772_, new_A773_, new_A774_,
    new_A775_, new_A776_, new_A777_, new_A778_, new_A779_, new_A780_,
    new_A781_, new_A782_, new_A783_, new_A784_, new_A785_, new_A786_,
    new_A787_, new_A788_, new_A789_, new_A790_, new_A791_, new_A792_,
    new_A793_, new_A794_, new_A795_, new_A796_, new_A797_, new_A798_,
    new_A799_, new_A800_, new_A801_, new_A802_, new_A803_, new_A804_,
    new_A402_, new_A401_, new_A400_, new_A399_, new_A398_, new_A397_,
    new_A396_, new_A395_, new_A394_, new_A393_, new_A392_, new_A391_,
    new_A390_, new_A389_, new_A388_, new_A387_, new_A386_, new_A385_,
    new_A384_, new_A383_, new_A382_, new_A381_, new_A380_, new_A379_,
    new_A378_, new_A377_, new_A376_, new_A375_, new_A374_, new_A373_,
    new_A372_, new_A371_, new_A370_, new_A369_, new_A368_, new_A367_,
    new_A366_, new_A365_, new_A364_, new_A363_, new_A362_, new_A361_,
    new_A360_, new_A359_, new_A358_, new_A357_, new_A356_, new_A355_,
    new_A354_, new_A353_, new_A352_, new_A351_, new_A350_, new_A349_,
    new_A348_, new_A341_, new_A340_, new_A339_, new_A338_, new_A337_,
    new_A336_, new_A335_, new_A334_, new_A333_, new_A332_, new_A331_,
    new_A330_, new_A329_, new_A328_, new_A327_, new_A326_, new_A325_,
    new_A324_, new_A323_, new_A322_, new_A321_, new_A320_, new_A319_,
    new_A318_, new_A317_, new_A316_, new_A315_, new_A314_, new_A313_,
    new_A312_, new_A311_, new_A310_, new_A309_, new_A308_, new_A307_,
    new_A306_, new_A305_, new_A304_, new_A303_, new_A302_, new_A301_,
    new_A300_, new_A299_, new_A298_, new_A297_, new_A296_, new_A295_,
    new_A294_, new_A293_, new_A292_, new_A291_, new_A290_, new_A289_,
    new_A288_, new_A287_, new_A286_, new_A285_, new_A284_, new_A283_,
    new_A282_, new_A281_, new_A274_, new_A273_, new_A272_, new_A271_,
    new_A270_, new_A269_, new_A268_, new_A267_, new_A266_, new_A265_,
    new_A264_, new_A263_, new_A262_, new_A261_, new_A260_, new_A259_,
    new_A258_, new_A257_, new_A256_, new_A255_, new_A254_, new_A253_,
    new_A252_, new_A251_, new_A250_, new_A249_, new_A248_, new_A247_,
    new_A246_, new_A245_, new_A244_, new_A243_, new_A242_, new_A241_,
    new_A240_, new_A239_, new_A238_, new_A237_, new_A236_, new_A235_,
    new_A234_, new_A233_, new_A232_, new_A231_, new_A230_, new_A229_,
    new_A228_, new_A227_, new_A226_, new_A225_, new_A224_, new_A223_,
    new_A222_, new_A221_, new_A220_, new_A219_, new_A218_, new_A217_,
    new_A216_, new_A215_, new_A214_, new_A207_, new_A206_, new_A205_,
    new_A204_, new_A203_, new_A202_, new_A201_, new_A200_, new_A199_,
    new_A198_, new_A197_, new_A196_, new_A195_, new_A194_, new_A193_,
    new_A192_, new_A191_, new_A190_, new_A189_, new_A188_, new_A187_,
    new_A186_, new_A185_, new_A184_, new_A183_, new_A182_, new_A181_,
    new_A180_, new_A179_, new_A178_, new_A177_, new_A176_, new_A175_,
    new_A174_, new_A173_, new_A172_, new_A171_, new_A170_, new_A169_,
    new_A168_, new_A167_, new_A166_, new_A165_, new_A164_, new_A163_,
    new_A162_, new_A161_, new_A160_, new_A159_, new_A158_, new_A157_,
    new_A156_, new_A155_, new_A154_, new_A153_, new_A152_, new_A151_,
    new_A150_, new_A149_, new_A148_, new_A147_, new_A140_, new_A139_,
    new_A138_, new_A137_, new_A136_, new_A135_, new_A134_, new_A133_,
    new_A132_, new_A131_, new_A130_, new_A129_, new_A128_, new_A127_,
    new_A126_, new_A125_, new_A124_, new_A123_, new_A122_, new_A121_,
    new_A120_, new_A119_, new_A118_, new_A117_, new_A116_, new_A115_,
    new_A114_, new_A113_, new_A112_, new_A111_, new_A110_, new_A109_,
    new_A108_, new_A107_, new_A106_, new_A105_, new_A104_, new_A103_,
    new_A102_, new_A101_, new_A100_, new_A99_, new_A98_, new_A97_,
    new_A96_, new_A95_, new_A94_, new_A93_, new_A92_, new_A91_, new_A90_,
    new_A89_, new_A88_, new_A87_, new_A86_, new_A85_, new_A84_, new_A83_,
    new_A82_, new_A81_, new_A80_, new_A73_, new_A72_, new_A71_, new_A70_,
    new_A69_, new_A68_, new_A1_, new_A2_, new_A3_, new_A4_, new_A5_,
    new_A6_, new_A13_, new_A14_, new_A15_, new_A16_, new_A17_, new_A18_,
    new_A19_, new_A20_, new_A21_, new_A22_, new_A23_, new_A24_, new_A25_,
    new_A26_, new_A27_, new_A28_, new_A29_, new_A30_, new_A31_, new_A32_,
    new_A33_, new_A34_, new_A35_, new_A36_, new_A37_, new_A38_, new_A39_,
    new_A40_, new_A41_, new_A42_, new_A43_, new_A44_, new_A45_, new_A46_,
    new_A47_, new_A48_, new_A49_, new_A50_, new_A51_, new_A52_, new_A53_,
    new_A54_, new_A55_, new_A56_, new_A57_, new_A58_, new_A59_, new_A60_,
    new_A61_, new_A62_, new_A63_, new_A64_, new_A65_, new_A66_, new_A67_;
  assign new_A469_ = ~A408 & new_A422_;
  assign new_A468_ = A408 & ~new_A422_;
  assign new_A467_ = A408 & ~new_A422_;
  assign new_A466_ = ~A408 & ~new_A422_;
  assign new_A465_ = A408 & new_A422_;
  assign new_A464_ = new_A468_ | new_A469_;
  assign new_A463_ = ~A408 & new_A422_;
  assign new_A462_ = new_A466_ | new_A467_;
  assign new_A461_ = ~new_A437_ & ~new_A457_;
  assign new_A460_ = new_A437_ & new_A457_;
  assign new_A459_ = ~A404 | ~new_A429_;
  assign new_A458_ = new_A422_ & new_A459_;
  assign new_A457_ = A405 | A406;
  assign new_A456_ = A405 | new_A422_;
  assign new_A455_ = ~new_A422_ & ~new_A458_;
  assign new_A454_ = new_A422_ | new_A459_;
  assign new_A453_ = A405 & ~A406;
  assign new_A452_ = ~A405 & A406;
  assign new_A451_ = new_A415_ | new_A448_;
  assign new_A450_ = ~new_A415_ & ~new_A449_;
  assign new_A449_ = new_A415_ & new_A448_;
  assign new_A448_ = ~A404 | ~new_A429_;
  assign new_A447_ = ~A405 & new_A415_;
  assign new_A446_ = A405 & ~new_A415_;
  assign new_A445_ = A407 & new_A444_;
  assign new_A444_ = new_A463_ | new_A462_;
  assign new_A443_ = ~A407 & new_A442_;
  assign new_A442_ = new_A465_ | new_A464_;
  assign new_A441_ = A407 | new_A440_;
  assign new_A440_ = new_A461_ | new_A460_;
  assign new_A439_ = ~new_A419_ & ~new_A429_;
  assign new_A438_ = new_A419_ & new_A429_;
  assign new_A437_ = ~new_A419_ | new_A429_;
  assign new_A436_ = A403 & ~A404;
  assign new_A435_ = ~A403 & A404;
  assign new_A434_ = new_A456_ & ~new_A457_;
  assign new_A433_ = ~new_A456_ & new_A457_;
  assign new_A432_ = ~new_A455_ | ~new_A454_;
  assign new_A431_ = new_A447_ | new_A446_;
  assign new_A430_ = new_A453_ | new_A452_;
  assign new_A429_ = new_A443_ | new_A445_;
  assign new_A428_ = ~new_A450_ | ~new_A451_;
  assign new_A427_ = A403 & ~A404;
  assign new_A426_ = new_A417_ & ~new_A429_;
  assign new_A425_ = ~new_A417_ & new_A429_;
  assign new_A424_ = ~new_A415_ & new_A441_;
  assign new_A423_ = new_A439_ | new_A438_;
  assign new_A422_ = new_A436_ | new_A435_;
  assign new_A421_ = A404 | new_A437_;
  assign new_A420_ = new_A429_ & new_A432_;
  assign new_A419_ = new_A434_ | new_A433_;
  assign new_A418_ = new_A429_ & new_A428_;
  assign new_A417_ = new_A431_ & new_A430_;
  assign new_A416_ = new_A426_ | new_A425_;
  assign new_A415_ = A404 | new_A427_;
  assign new_A414_ = new_A415_ | new_A424_;
  assign new_A413_ = new_A422_ & new_A423_;
  assign new_A412_ = new_A422_ & new_A421_;
  assign new_A411_ = new_A420_ | new_A419_;
  assign new_A410_ = new_A418_ | new_A417_;
  assign new_A409_ = new_A416_ & new_A415_;
  assign new_A476_ = new_A483_ & new_A482_;
  assign new_A477_ = new_A485_ | new_A484_;
  assign new_A478_ = new_A487_ | new_A486_;
  assign new_A479_ = new_A489_ & new_A488_;
  assign new_A480_ = new_A489_ & new_A490_;
  assign new_A481_ = new_A482_ | new_A491_;
  assign new_A482_ = A471 | new_A494_;
  assign new_A483_ = new_A493_ | new_A492_;
  assign new_A484_ = new_A498_ & new_A497_;
  assign new_A485_ = new_A496_ & new_A495_;
  assign new_A486_ = new_A501_ | new_A500_;
  assign new_A487_ = new_A496_ & new_A499_;
  assign new_A488_ = A471 | new_A504_;
  assign new_A489_ = new_A503_ | new_A502_;
  assign new_A490_ = new_A506_ | new_A505_;
  assign new_A491_ = ~new_A482_ & new_A508_;
  assign new_A492_ = ~new_A484_ & new_A496_;
  assign new_A493_ = new_A484_ & ~new_A496_;
  assign new_A494_ = A470 & ~A471;
  assign new_A495_ = ~new_A517_ | ~new_A518_;
  assign new_A496_ = new_A510_ | new_A512_;
  assign new_A497_ = new_A520_ | new_A519_;
  assign new_A498_ = new_A514_ | new_A513_;
  assign new_A499_ = ~new_A522_ | ~new_A521_;
  assign new_A500_ = ~new_A523_ & new_A524_;
  assign new_A501_ = new_A523_ & ~new_A524_;
  assign new_A502_ = ~A470 & A471;
  assign new_A503_ = A470 & ~A471;
  assign new_A504_ = ~new_A486_ | new_A496_;
  assign new_A505_ = new_A486_ & new_A496_;
  assign new_A506_ = ~new_A486_ & ~new_A496_;
  assign new_A507_ = new_A528_ | new_A527_;
  assign new_A508_ = A474 | new_A507_;
  assign new_A509_ = new_A532_ | new_A531_;
  assign new_A510_ = ~A474 & new_A509_;
  assign new_A511_ = new_A530_ | new_A529_;
  assign new_A512_ = A474 & new_A511_;
  assign new_A513_ = A472 & ~new_A482_;
  assign new_A514_ = ~A472 & new_A482_;
  assign new_A515_ = ~A471 | ~new_A496_;
  assign new_A516_ = new_A482_ & new_A515_;
  assign new_A517_ = ~new_A482_ & ~new_A516_;
  assign new_A518_ = new_A482_ | new_A515_;
  assign new_A519_ = ~A472 & A473;
  assign new_A520_ = A472 & ~A473;
  assign new_A521_ = new_A489_ | new_A526_;
  assign new_A522_ = ~new_A489_ & ~new_A525_;
  assign new_A523_ = A472 | new_A489_;
  assign new_A524_ = A472 | A473;
  assign new_A525_ = new_A489_ & new_A526_;
  assign new_A526_ = ~A471 | ~new_A496_;
  assign new_A527_ = new_A504_ & new_A524_;
  assign new_A528_ = ~new_A504_ & ~new_A524_;
  assign new_A529_ = new_A533_ | new_A534_;
  assign new_A530_ = ~A475 & new_A489_;
  assign new_A531_ = new_A535_ | new_A536_;
  assign new_A532_ = A475 & new_A489_;
  assign new_A533_ = ~A475 & ~new_A489_;
  assign new_A534_ = A475 & ~new_A489_;
  assign new_A535_ = A475 & ~new_A489_;
  assign new_A536_ = ~A475 & new_A489_;
  assign new_A543_ = new_A550_ & new_A549_;
  assign new_A544_ = new_A552_ | new_A551_;
  assign new_A545_ = new_A554_ | new_A553_;
  assign new_A546_ = new_A556_ & new_A555_;
  assign new_A547_ = new_A556_ & new_A557_;
  assign new_A548_ = new_A549_ | new_A558_;
  assign new_A549_ = A538 | new_A561_;
  assign new_A550_ = new_A560_ | new_A559_;
  assign new_A551_ = new_A565_ & new_A564_;
  assign new_A552_ = new_A563_ & new_A562_;
  assign new_A553_ = new_A568_ | new_A567_;
  assign new_A554_ = new_A563_ & new_A566_;
  assign new_A555_ = A538 | new_A571_;
  assign new_A556_ = new_A570_ | new_A569_;
  assign new_A557_ = new_A573_ | new_A572_;
  assign new_A558_ = ~new_A549_ & new_A575_;
  assign new_A559_ = ~new_A551_ & new_A563_;
  assign new_A560_ = new_A551_ & ~new_A563_;
  assign new_A561_ = A537 & ~A538;
  assign new_A562_ = ~new_A584_ | ~new_A585_;
  assign new_A563_ = new_A577_ | new_A579_;
  assign new_A564_ = new_A587_ | new_A586_;
  assign new_A565_ = new_A581_ | new_A580_;
  assign new_A566_ = ~new_A589_ | ~new_A588_;
  assign new_A567_ = ~new_A590_ & new_A591_;
  assign new_A568_ = new_A590_ & ~new_A591_;
  assign new_A569_ = ~A537 & A538;
  assign new_A570_ = A537 & ~A538;
  assign new_A571_ = ~new_A553_ | new_A563_;
  assign new_A572_ = new_A553_ & new_A563_;
  assign new_A573_ = ~new_A553_ & ~new_A563_;
  assign new_A574_ = new_A595_ | new_A594_;
  assign new_A575_ = A541 | new_A574_;
  assign new_A576_ = new_A599_ | new_A598_;
  assign new_A577_ = ~A541 & new_A576_;
  assign new_A578_ = new_A597_ | new_A596_;
  assign new_A579_ = A541 & new_A578_;
  assign new_A580_ = A539 & ~new_A549_;
  assign new_A581_ = ~A539 & new_A549_;
  assign new_A582_ = ~A538 | ~new_A563_;
  assign new_A583_ = new_A549_ & new_A582_;
  assign new_A584_ = ~new_A549_ & ~new_A583_;
  assign new_A585_ = new_A549_ | new_A582_;
  assign new_A586_ = ~A539 & A540;
  assign new_A587_ = A539 & ~A540;
  assign new_A588_ = new_A556_ | new_A593_;
  assign new_A589_ = ~new_A556_ & ~new_A592_;
  assign new_A590_ = A539 | new_A556_;
  assign new_A591_ = A539 | A540;
  assign new_A592_ = new_A556_ & new_A593_;
  assign new_A593_ = ~A538 | ~new_A563_;
  assign new_A594_ = new_A571_ & new_A591_;
  assign new_A595_ = ~new_A571_ & ~new_A591_;
  assign new_A596_ = new_A600_ | new_A601_;
  assign new_A597_ = ~A542 & new_A556_;
  assign new_A598_ = new_A602_ | new_A603_;
  assign new_A599_ = A542 & new_A556_;
  assign new_A600_ = ~A542 & ~new_A556_;
  assign new_A601_ = A542 & ~new_A556_;
  assign new_A602_ = A542 & ~new_A556_;
  assign new_A603_ = ~A542 & new_A556_;
  assign new_A610_ = new_A617_ & new_A616_;
  assign new_A611_ = new_A619_ | new_A618_;
  assign new_A612_ = new_A621_ | new_A620_;
  assign new_A613_ = new_A623_ & new_A622_;
  assign new_A614_ = new_A623_ & new_A624_;
  assign new_A615_ = new_A616_ | new_A625_;
  assign new_A616_ = A605 | new_A628_;
  assign new_A617_ = new_A627_ | new_A626_;
  assign new_A618_ = new_A632_ & new_A631_;
  assign new_A619_ = new_A630_ & new_A629_;
  assign new_A620_ = new_A635_ | new_A634_;
  assign new_A621_ = new_A630_ & new_A633_;
  assign new_A622_ = A605 | new_A638_;
  assign new_A623_ = new_A637_ | new_A636_;
  assign new_A624_ = new_A640_ | new_A639_;
  assign new_A625_ = ~new_A616_ & new_A642_;
  assign new_A626_ = ~new_A618_ & new_A630_;
  assign new_A627_ = new_A618_ & ~new_A630_;
  assign new_A628_ = A604 & ~A605;
  assign new_A629_ = ~new_A651_ | ~new_A652_;
  assign new_A630_ = new_A644_ | new_A646_;
  assign new_A631_ = new_A654_ | new_A653_;
  assign new_A632_ = new_A648_ | new_A647_;
  assign new_A633_ = ~new_A656_ | ~new_A655_;
  assign new_A634_ = ~new_A657_ & new_A658_;
  assign new_A635_ = new_A657_ & ~new_A658_;
  assign new_A636_ = ~A604 & A605;
  assign new_A637_ = A604 & ~A605;
  assign new_A638_ = ~new_A620_ | new_A630_;
  assign new_A639_ = new_A620_ & new_A630_;
  assign new_A640_ = ~new_A620_ & ~new_A630_;
  assign new_A641_ = new_A662_ | new_A661_;
  assign new_A642_ = A608 | new_A641_;
  assign new_A643_ = new_A666_ | new_A665_;
  assign new_A644_ = ~A608 & new_A643_;
  assign new_A645_ = new_A664_ | new_A663_;
  assign new_A646_ = A608 & new_A645_;
  assign new_A647_ = A606 & ~new_A616_;
  assign new_A648_ = ~A606 & new_A616_;
  assign new_A649_ = ~A605 | ~new_A630_;
  assign new_A650_ = new_A616_ & new_A649_;
  assign new_A651_ = ~new_A616_ & ~new_A650_;
  assign new_A652_ = new_A616_ | new_A649_;
  assign new_A653_ = ~A606 & A607;
  assign new_A654_ = A606 & ~A607;
  assign new_A655_ = new_A623_ | new_A660_;
  assign new_A656_ = ~new_A623_ & ~new_A659_;
  assign new_A657_ = A606 | new_A623_;
  assign new_A658_ = A606 | A607;
  assign new_A659_ = new_A623_ & new_A660_;
  assign new_A660_ = ~A605 | ~new_A630_;
  assign new_A661_ = new_A638_ & new_A658_;
  assign new_A662_ = ~new_A638_ & ~new_A658_;
  assign new_A663_ = new_A667_ | new_A668_;
  assign new_A664_ = ~A609 & new_A623_;
  assign new_A665_ = new_A669_ | new_A670_;
  assign new_A666_ = A609 & new_A623_;
  assign new_A667_ = ~A609 & ~new_A623_;
  assign new_A668_ = A609 & ~new_A623_;
  assign new_A669_ = A609 & ~new_A623_;
  assign new_A670_ = ~A609 & new_A623_;
  assign new_A677_ = new_A684_ & new_A683_;
  assign new_A678_ = new_A686_ | new_A685_;
  assign new_A679_ = new_A688_ | new_A687_;
  assign new_A680_ = new_A690_ & new_A689_;
  assign new_A681_ = new_A690_ & new_A691_;
  assign new_A682_ = new_A683_ | new_A692_;
  assign new_A683_ = A672 | new_A695_;
  assign new_A684_ = new_A694_ | new_A693_;
  assign new_A685_ = new_A699_ & new_A698_;
  assign new_A686_ = new_A697_ & new_A696_;
  assign new_A687_ = new_A702_ | new_A701_;
  assign new_A688_ = new_A697_ & new_A700_;
  assign new_A689_ = A672 | new_A705_;
  assign new_A690_ = new_A704_ | new_A703_;
  assign new_A691_ = new_A707_ | new_A706_;
  assign new_A692_ = ~new_A683_ & new_A709_;
  assign new_A693_ = ~new_A685_ & new_A697_;
  assign new_A694_ = new_A685_ & ~new_A697_;
  assign new_A695_ = A671 & ~A672;
  assign new_A696_ = ~new_A718_ | ~new_A719_;
  assign new_A697_ = new_A711_ | new_A713_;
  assign new_A698_ = new_A721_ | new_A720_;
  assign new_A699_ = new_A715_ | new_A714_;
  assign new_A700_ = ~new_A723_ | ~new_A722_;
  assign new_A701_ = ~new_A724_ & new_A725_;
  assign new_A702_ = new_A724_ & ~new_A725_;
  assign new_A703_ = ~A671 & A672;
  assign new_A704_ = A671 & ~A672;
  assign new_A705_ = ~new_A687_ | new_A697_;
  assign new_A706_ = new_A687_ & new_A697_;
  assign new_A707_ = ~new_A687_ & ~new_A697_;
  assign new_A708_ = new_A729_ | new_A728_;
  assign new_A709_ = A675 | new_A708_;
  assign new_A710_ = new_A733_ | new_A732_;
  assign new_A711_ = ~A675 & new_A710_;
  assign new_A712_ = new_A731_ | new_A730_;
  assign new_A713_ = A675 & new_A712_;
  assign new_A714_ = A673 & ~new_A683_;
  assign new_A715_ = ~A673 & new_A683_;
  assign new_A716_ = ~A672 | ~new_A697_;
  assign new_A717_ = new_A683_ & new_A716_;
  assign new_A718_ = ~new_A683_ & ~new_A717_;
  assign new_A719_ = new_A683_ | new_A716_;
  assign new_A720_ = ~A673 & A674;
  assign new_A721_ = A673 & ~A674;
  assign new_A722_ = new_A690_ | new_A727_;
  assign new_A723_ = ~new_A690_ & ~new_A726_;
  assign new_A724_ = A673 | new_A690_;
  assign new_A725_ = A673 | A674;
  assign new_A726_ = new_A690_ & new_A727_;
  assign new_A727_ = ~A672 | ~new_A697_;
  assign new_A728_ = new_A705_ & new_A725_;
  assign new_A729_ = ~new_A705_ & ~new_A725_;
  assign new_A730_ = new_A734_ | new_A735_;
  assign new_A731_ = ~A676 & new_A690_;
  assign new_A732_ = new_A736_ | new_A737_;
  assign new_A733_ = A676 & new_A690_;
  assign new_A734_ = ~A676 & ~new_A690_;
  assign new_A735_ = A676 & ~new_A690_;
  assign new_A736_ = A676 & ~new_A690_;
  assign new_A737_ = ~A676 & new_A690_;
  assign new_A744_ = new_A751_ & new_A750_;
  assign new_A745_ = new_A753_ | new_A752_;
  assign new_A746_ = new_A755_ | new_A754_;
  assign new_A747_ = new_A757_ & new_A756_;
  assign new_A748_ = new_A757_ & new_A758_;
  assign new_A749_ = new_A750_ | new_A759_;
  assign new_A750_ = A739 | new_A762_;
  assign new_A751_ = new_A761_ | new_A760_;
  assign new_A752_ = new_A766_ & new_A765_;
  assign new_A753_ = new_A764_ & new_A763_;
  assign new_A754_ = new_A769_ | new_A768_;
  assign new_A755_ = new_A764_ & new_A767_;
  assign new_A756_ = A739 | new_A772_;
  assign new_A757_ = new_A771_ | new_A770_;
  assign new_A758_ = new_A774_ | new_A773_;
  assign new_A759_ = ~new_A750_ & new_A776_;
  assign new_A760_ = ~new_A752_ & new_A764_;
  assign new_A761_ = new_A752_ & ~new_A764_;
  assign new_A762_ = A738 & ~A739;
  assign new_A763_ = ~new_A785_ | ~new_A786_;
  assign new_A764_ = new_A778_ | new_A780_;
  assign new_A765_ = new_A788_ | new_A787_;
  assign new_A766_ = new_A782_ | new_A781_;
  assign new_A767_ = ~new_A790_ | ~new_A789_;
  assign new_A768_ = ~new_A791_ & new_A792_;
  assign new_A769_ = new_A791_ & ~new_A792_;
  assign new_A770_ = ~A738 & A739;
  assign new_A771_ = A738 & ~A739;
  assign new_A772_ = ~new_A754_ | new_A764_;
  assign new_A773_ = new_A754_ & new_A764_;
  assign new_A774_ = ~new_A754_ & ~new_A764_;
  assign new_A775_ = new_A796_ | new_A795_;
  assign new_A776_ = A742 | new_A775_;
  assign new_A777_ = new_A800_ | new_A799_;
  assign new_A778_ = ~A742 & new_A777_;
  assign new_A779_ = new_A798_ | new_A797_;
  assign new_A780_ = A742 & new_A779_;
  assign new_A781_ = A740 & ~new_A750_;
  assign new_A782_ = ~A740 & new_A750_;
  assign new_A783_ = ~A739 | ~new_A764_;
  assign new_A784_ = new_A750_ & new_A783_;
  assign new_A785_ = ~new_A750_ & ~new_A784_;
  assign new_A786_ = new_A750_ | new_A783_;
  assign new_A787_ = ~A740 & A741;
  assign new_A788_ = A740 & ~A741;
  assign new_A789_ = new_A757_ | new_A794_;
  assign new_A790_ = ~new_A757_ & ~new_A793_;
  assign new_A791_ = A740 | new_A757_;
  assign new_A792_ = A740 | A741;
  assign new_A793_ = new_A757_ & new_A794_;
  assign new_A794_ = ~A739 | ~new_A764_;
  assign new_A795_ = new_A772_ & new_A792_;
  assign new_A796_ = ~new_A772_ & ~new_A792_;
  assign new_A797_ = new_A801_ | new_A802_;
  assign new_A798_ = ~A743 & new_A757_;
  assign new_A799_ = new_A803_ | new_A804_;
  assign new_A800_ = A743 & new_A757_;
  assign new_A801_ = ~A743 & ~new_A757_;
  assign new_A802_ = A743 & ~new_A757_;
  assign new_A803_ = A743 & ~new_A757_;
  assign new_A804_ = ~A743 & new_A757_;
  assign new_A402_ = ~new_A341_ & new_A355_;
  assign new_A401_ = new_A341_ & ~new_A355_;
  assign new_A400_ = new_A341_ & ~new_A355_;
  assign new_A399_ = ~new_A341_ & ~new_A355_;
  assign new_A398_ = new_A341_ & new_A355_;
  assign new_A397_ = new_A401_ | new_A402_;
  assign new_A396_ = ~new_A341_ & new_A355_;
  assign new_A395_ = new_A399_ | new_A400_;
  assign new_A394_ = ~new_A370_ & ~new_A390_;
  assign new_A393_ = new_A370_ & new_A390_;
  assign new_A392_ = ~new_A337_ | ~new_A362_;
  assign new_A391_ = new_A355_ & new_A392_;
  assign new_A390_ = new_A338_ | new_A339_;
  assign new_A389_ = new_A338_ | new_A355_;
  assign new_A388_ = ~new_A355_ & ~new_A391_;
  assign new_A387_ = new_A355_ | new_A392_;
  assign new_A386_ = new_A338_ & ~new_A339_;
  assign new_A385_ = ~new_A338_ & new_A339_;
  assign new_A384_ = new_A348_ | new_A381_;
  assign new_A383_ = ~new_A348_ & ~new_A382_;
  assign new_A382_ = new_A348_ & new_A381_;
  assign new_A381_ = ~new_A337_ | ~new_A362_;
  assign new_A380_ = ~new_A338_ & new_A348_;
  assign new_A379_ = new_A338_ & ~new_A348_;
  assign new_A378_ = new_A340_ & new_A377_;
  assign new_A377_ = new_A396_ | new_A395_;
  assign new_A376_ = ~new_A340_ & new_A375_;
  assign new_A375_ = new_A398_ | new_A397_;
  assign new_A374_ = new_A340_ | new_A373_;
  assign new_A373_ = new_A394_ | new_A393_;
  assign new_A372_ = ~new_A352_ & ~new_A362_;
  assign new_A371_ = new_A352_ & new_A362_;
  assign new_A370_ = ~new_A352_ | new_A362_;
  assign new_A369_ = new_A336_ & ~new_A337_;
  assign new_A368_ = ~new_A336_ & new_A337_;
  assign new_A367_ = new_A389_ & ~new_A390_;
  assign new_A366_ = ~new_A389_ & new_A390_;
  assign new_A365_ = ~new_A388_ | ~new_A387_;
  assign new_A364_ = new_A380_ | new_A379_;
  assign new_A363_ = new_A386_ | new_A385_;
  assign new_A362_ = new_A376_ | new_A378_;
  assign new_A361_ = ~new_A383_ | ~new_A384_;
  assign new_A360_ = new_A336_ & ~new_A337_;
  assign new_A359_ = new_A350_ & ~new_A362_;
  assign new_A358_ = ~new_A350_ & new_A362_;
  assign new_A357_ = ~new_A348_ & new_A374_;
  assign new_A356_ = new_A372_ | new_A371_;
  assign new_A355_ = new_A369_ | new_A368_;
  assign new_A354_ = new_A337_ | new_A370_;
  assign new_A353_ = new_A362_ & new_A365_;
  assign new_A352_ = new_A367_ | new_A366_;
  assign new_A351_ = new_A362_ & new_A361_;
  assign new_A350_ = new_A364_ & new_A363_;
  assign new_A349_ = new_A359_ | new_A358_;
  assign new_A348_ = new_A337_ | new_A360_;
  assign A347 = new_A348_ | new_A357_;
  assign A346 = new_A355_ & new_A356_;
  assign A345 = new_A355_ & new_A354_;
  assign A344 = new_A353_ | new_A352_;
  assign A343 = new_A351_ | new_A350_;
  assign A342 = new_A349_ & new_A348_;
  assign new_A341_ = new_A749_;
  assign new_A340_ = new_A682_;
  assign new_A339_ = new_A615_;
  assign new_A338_ = new_A548_;
  assign new_A337_ = new_A481_;
  assign new_A336_ = new_A409_;
  assign new_A335_ = ~new_A274_ & new_A288_;
  assign new_A334_ = new_A274_ & ~new_A288_;
  assign new_A333_ = new_A274_ & ~new_A288_;
  assign new_A332_ = ~new_A274_ & ~new_A288_;
  assign new_A331_ = new_A274_ & new_A288_;
  assign new_A330_ = new_A334_ | new_A335_;
  assign new_A329_ = ~new_A274_ & new_A288_;
  assign new_A328_ = new_A332_ | new_A333_;
  assign new_A327_ = ~new_A303_ & ~new_A323_;
  assign new_A326_ = new_A303_ & new_A323_;
  assign new_A325_ = ~new_A270_ | ~new_A295_;
  assign new_A324_ = new_A288_ & new_A325_;
  assign new_A323_ = new_A271_ | new_A272_;
  assign new_A322_ = new_A271_ | new_A288_;
  assign new_A321_ = ~new_A288_ & ~new_A324_;
  assign new_A320_ = new_A288_ | new_A325_;
  assign new_A319_ = new_A271_ & ~new_A272_;
  assign new_A318_ = ~new_A271_ & new_A272_;
  assign new_A317_ = new_A281_ | new_A314_;
  assign new_A316_ = ~new_A281_ & ~new_A315_;
  assign new_A315_ = new_A281_ & new_A314_;
  assign new_A314_ = ~new_A270_ | ~new_A295_;
  assign new_A313_ = ~new_A271_ & new_A281_;
  assign new_A312_ = new_A271_ & ~new_A281_;
  assign new_A311_ = new_A273_ & new_A310_;
  assign new_A310_ = new_A329_ | new_A328_;
  assign new_A309_ = ~new_A273_ & new_A308_;
  assign new_A308_ = new_A331_ | new_A330_;
  assign new_A307_ = new_A273_ | new_A306_;
  assign new_A306_ = new_A327_ | new_A326_;
  assign new_A305_ = ~new_A285_ & ~new_A295_;
  assign new_A304_ = new_A285_ & new_A295_;
  assign new_A303_ = ~new_A285_ | new_A295_;
  assign new_A302_ = new_A269_ & ~new_A270_;
  assign new_A301_ = ~new_A269_ & new_A270_;
  assign new_A300_ = new_A322_ & ~new_A323_;
  assign new_A299_ = ~new_A322_ & new_A323_;
  assign new_A298_ = ~new_A321_ | ~new_A320_;
  assign new_A297_ = new_A313_ | new_A312_;
  assign new_A296_ = new_A319_ | new_A318_;
  assign new_A295_ = new_A309_ | new_A311_;
  assign new_A294_ = ~new_A316_ | ~new_A317_;
  assign new_A293_ = new_A269_ & ~new_A270_;
  assign new_A292_ = new_A283_ & ~new_A295_;
  assign new_A291_ = ~new_A283_ & new_A295_;
  assign new_A290_ = ~new_A281_ & new_A307_;
  assign new_A289_ = new_A305_ | new_A304_;
  assign new_A288_ = new_A302_ | new_A301_;
  assign new_A287_ = new_A270_ | new_A303_;
  assign new_A286_ = new_A295_ & new_A298_;
  assign new_A285_ = new_A300_ | new_A299_;
  assign new_A284_ = new_A295_ & new_A294_;
  assign new_A283_ = new_A297_ & new_A296_;
  assign new_A282_ = new_A292_ | new_A291_;
  assign new_A281_ = new_A270_ | new_A293_;
  assign A280 = new_A281_ | new_A290_;
  assign A279 = new_A288_ & new_A289_;
  assign A278 = new_A288_ & new_A287_;
  assign A277 = new_A286_ | new_A285_;
  assign A276 = new_A284_ | new_A283_;
  assign A275 = new_A282_ & new_A281_;
  assign new_A274_ = new_A748_;
  assign new_A273_ = new_A681_;
  assign new_A272_ = new_A614_;
  assign new_A271_ = new_A547_;
  assign new_A270_ = new_A480_;
  assign new_A269_ = new_A410_;
  assign new_A268_ = ~new_A207_ & new_A221_;
  assign new_A267_ = new_A207_ & ~new_A221_;
  assign new_A266_ = new_A207_ & ~new_A221_;
  assign new_A265_ = ~new_A207_ & ~new_A221_;
  assign new_A264_ = new_A207_ & new_A221_;
  assign new_A263_ = new_A267_ | new_A268_;
  assign new_A262_ = ~new_A207_ & new_A221_;
  assign new_A261_ = new_A265_ | new_A266_;
  assign new_A260_ = ~new_A236_ & ~new_A256_;
  assign new_A259_ = new_A236_ & new_A256_;
  assign new_A258_ = ~new_A203_ | ~new_A228_;
  assign new_A257_ = new_A221_ & new_A258_;
  assign new_A256_ = new_A204_ | new_A205_;
  assign new_A255_ = new_A204_ | new_A221_;
  assign new_A254_ = ~new_A221_ & ~new_A257_;
  assign new_A253_ = new_A221_ | new_A258_;
  assign new_A252_ = new_A204_ & ~new_A205_;
  assign new_A251_ = ~new_A204_ & new_A205_;
  assign new_A250_ = new_A214_ | new_A247_;
  assign new_A249_ = ~new_A214_ & ~new_A248_;
  assign new_A248_ = new_A214_ & new_A247_;
  assign new_A247_ = ~new_A203_ | ~new_A228_;
  assign new_A246_ = ~new_A204_ & new_A214_;
  assign new_A245_ = new_A204_ & ~new_A214_;
  assign new_A244_ = new_A206_ & new_A243_;
  assign new_A243_ = new_A262_ | new_A261_;
  assign new_A242_ = ~new_A206_ & new_A241_;
  assign new_A241_ = new_A264_ | new_A263_;
  assign new_A240_ = new_A206_ | new_A239_;
  assign new_A239_ = new_A260_ | new_A259_;
  assign new_A238_ = ~new_A218_ & ~new_A228_;
  assign new_A237_ = new_A218_ & new_A228_;
  assign new_A236_ = ~new_A218_ | new_A228_;
  assign new_A235_ = new_A202_ & ~new_A203_;
  assign new_A234_ = ~new_A202_ & new_A203_;
  assign new_A233_ = new_A255_ & ~new_A256_;
  assign new_A232_ = ~new_A255_ & new_A256_;
  assign new_A231_ = ~new_A254_ | ~new_A253_;
  assign new_A230_ = new_A246_ | new_A245_;
  assign new_A229_ = new_A252_ | new_A251_;
  assign new_A228_ = new_A242_ | new_A244_;
  assign new_A227_ = ~new_A249_ | ~new_A250_;
  assign new_A226_ = new_A202_ & ~new_A203_;
  assign new_A225_ = new_A216_ & ~new_A228_;
  assign new_A224_ = ~new_A216_ & new_A228_;
  assign new_A223_ = ~new_A214_ & new_A240_;
  assign new_A222_ = new_A238_ | new_A237_;
  assign new_A221_ = new_A235_ | new_A234_;
  assign new_A220_ = new_A203_ | new_A236_;
  assign new_A219_ = new_A228_ & new_A231_;
  assign new_A218_ = new_A233_ | new_A232_;
  assign new_A217_ = new_A228_ & new_A227_;
  assign new_A216_ = new_A230_ & new_A229_;
  assign new_A215_ = new_A225_ | new_A224_;
  assign new_A214_ = new_A203_ | new_A226_;
  assign A213 = new_A214_ | new_A223_;
  assign A212 = new_A221_ & new_A222_;
  assign A211 = new_A221_ & new_A220_;
  assign A210 = new_A219_ | new_A218_;
  assign A209 = new_A217_ | new_A216_;
  assign A208 = new_A215_ & new_A214_;
  assign new_A207_ = new_A747_;
  assign new_A206_ = new_A680_;
  assign new_A205_ = new_A613_;
  assign new_A204_ = new_A546_;
  assign new_A203_ = new_A479_;
  assign new_A202_ = new_A411_;
  assign new_A201_ = ~new_A140_ & new_A154_;
  assign new_A200_ = new_A140_ & ~new_A154_;
  assign new_A199_ = new_A140_ & ~new_A154_;
  assign new_A198_ = ~new_A140_ & ~new_A154_;
  assign new_A197_ = new_A140_ & new_A154_;
  assign new_A196_ = new_A200_ | new_A201_;
  assign new_A195_ = ~new_A140_ & new_A154_;
  assign new_A194_ = new_A198_ | new_A199_;
  assign new_A193_ = ~new_A169_ & ~new_A189_;
  assign new_A192_ = new_A169_ & new_A189_;
  assign new_A191_ = ~new_A136_ | ~new_A161_;
  assign new_A190_ = new_A154_ & new_A191_;
  assign new_A189_ = new_A137_ | new_A138_;
  assign new_A188_ = new_A137_ | new_A154_;
  assign new_A187_ = ~new_A154_ & ~new_A190_;
  assign new_A186_ = new_A154_ | new_A191_;
  assign new_A185_ = new_A137_ & ~new_A138_;
  assign new_A184_ = ~new_A137_ & new_A138_;
  assign new_A183_ = new_A147_ | new_A180_;
  assign new_A182_ = ~new_A147_ & ~new_A181_;
  assign new_A181_ = new_A147_ & new_A180_;
  assign new_A180_ = ~new_A136_ | ~new_A161_;
  assign new_A179_ = ~new_A137_ & new_A147_;
  assign new_A178_ = new_A137_ & ~new_A147_;
  assign new_A177_ = new_A139_ & new_A176_;
  assign new_A176_ = new_A195_ | new_A194_;
  assign new_A175_ = ~new_A139_ & new_A174_;
  assign new_A174_ = new_A197_ | new_A196_;
  assign new_A173_ = new_A139_ | new_A172_;
  assign new_A172_ = new_A193_ | new_A192_;
  assign new_A171_ = ~new_A151_ & ~new_A161_;
  assign new_A170_ = new_A151_ & new_A161_;
  assign new_A169_ = ~new_A151_ | new_A161_;
  assign new_A168_ = new_A135_ & ~new_A136_;
  assign new_A167_ = ~new_A135_ & new_A136_;
  assign new_A166_ = new_A188_ & ~new_A189_;
  assign new_A165_ = ~new_A188_ & new_A189_;
  assign new_A164_ = ~new_A187_ | ~new_A186_;
  assign new_A163_ = new_A179_ | new_A178_;
  assign new_A162_ = new_A185_ | new_A184_;
  assign new_A161_ = new_A175_ | new_A177_;
  assign new_A160_ = ~new_A182_ | ~new_A183_;
  assign new_A159_ = new_A135_ & ~new_A136_;
  assign new_A158_ = new_A149_ & ~new_A161_;
  assign new_A157_ = ~new_A149_ & new_A161_;
  assign new_A156_ = ~new_A147_ & new_A173_;
  assign new_A155_ = new_A171_ | new_A170_;
  assign new_A154_ = new_A168_ | new_A167_;
  assign new_A153_ = new_A136_ | new_A169_;
  assign new_A152_ = new_A161_ & new_A164_;
  assign new_A151_ = new_A166_ | new_A165_;
  assign new_A150_ = new_A161_ & new_A160_;
  assign new_A149_ = new_A163_ & new_A162_;
  assign new_A148_ = new_A158_ | new_A157_;
  assign new_A147_ = new_A136_ | new_A159_;
  assign A146 = new_A147_ | new_A156_;
  assign A145 = new_A154_ & new_A155_;
  assign A144 = new_A154_ & new_A153_;
  assign A143 = new_A152_ | new_A151_;
  assign A142 = new_A150_ | new_A149_;
  assign A141 = new_A148_ & new_A147_;
  assign new_A140_ = new_A746_;
  assign new_A139_ = new_A679_;
  assign new_A138_ = new_A612_;
  assign new_A137_ = new_A545_;
  assign new_A136_ = new_A478_;
  assign new_A135_ = new_A412_;
  assign new_A134_ = ~new_A73_ & new_A87_;
  assign new_A133_ = new_A73_ & ~new_A87_;
  assign new_A132_ = new_A73_ & ~new_A87_;
  assign new_A131_ = ~new_A73_ & ~new_A87_;
  assign new_A130_ = new_A73_ & new_A87_;
  assign new_A129_ = new_A133_ | new_A134_;
  assign new_A128_ = ~new_A73_ & new_A87_;
  assign new_A127_ = new_A131_ | new_A132_;
  assign new_A126_ = ~new_A102_ & ~new_A122_;
  assign new_A125_ = new_A102_ & new_A122_;
  assign new_A124_ = ~new_A69_ | ~new_A94_;
  assign new_A123_ = new_A87_ & new_A124_;
  assign new_A122_ = new_A70_ | new_A71_;
  assign new_A121_ = new_A70_ | new_A87_;
  assign new_A120_ = ~new_A87_ & ~new_A123_;
  assign new_A119_ = new_A87_ | new_A124_;
  assign new_A118_ = new_A70_ & ~new_A71_;
  assign new_A117_ = ~new_A70_ & new_A71_;
  assign new_A116_ = new_A80_ | new_A113_;
  assign new_A115_ = ~new_A80_ & ~new_A114_;
  assign new_A114_ = new_A80_ & new_A113_;
  assign new_A113_ = ~new_A69_ | ~new_A94_;
  assign new_A112_ = ~new_A70_ & new_A80_;
  assign new_A111_ = new_A70_ & ~new_A80_;
  assign new_A110_ = new_A72_ & new_A109_;
  assign new_A109_ = new_A128_ | new_A127_;
  assign new_A108_ = ~new_A72_ & new_A107_;
  assign new_A107_ = new_A130_ | new_A129_;
  assign new_A106_ = new_A72_ | new_A105_;
  assign new_A105_ = new_A126_ | new_A125_;
  assign new_A104_ = ~new_A84_ & ~new_A94_;
  assign new_A103_ = new_A84_ & new_A94_;
  assign new_A102_ = ~new_A84_ | new_A94_;
  assign new_A101_ = new_A68_ & ~new_A69_;
  assign new_A100_ = ~new_A68_ & new_A69_;
  assign new_A99_ = new_A121_ & ~new_A122_;
  assign new_A98_ = ~new_A121_ & new_A122_;
  assign new_A97_ = ~new_A120_ | ~new_A119_;
  assign new_A96_ = new_A112_ | new_A111_;
  assign new_A95_ = new_A118_ | new_A117_;
  assign new_A94_ = new_A108_ | new_A110_;
  assign new_A93_ = ~new_A115_ | ~new_A116_;
  assign new_A92_ = new_A68_ & ~new_A69_;
  assign new_A91_ = new_A82_ & ~new_A94_;
  assign new_A90_ = ~new_A82_ & new_A94_;
  assign new_A89_ = ~new_A80_ & new_A106_;
  assign new_A88_ = new_A104_ | new_A103_;
  assign new_A87_ = new_A101_ | new_A100_;
  assign new_A86_ = new_A69_ | new_A102_;
  assign new_A85_ = new_A94_ & new_A97_;
  assign new_A84_ = new_A99_ | new_A98_;
  assign new_A83_ = new_A94_ & new_A93_;
  assign new_A82_ = new_A96_ & new_A95_;
  assign new_A81_ = new_A91_ | new_A90_;
  assign new_A80_ = new_A69_ | new_A92_;
  assign A79 = new_A80_ | new_A89_;
  assign A78 = new_A87_ & new_A88_;
  assign A77 = new_A87_ & new_A86_;
  assign A76 = new_A85_ | new_A84_;
  assign A75 = new_A83_ | new_A82_;
  assign A74 = new_A81_ & new_A80_;
  assign new_A73_ = new_A745_;
  assign new_A72_ = new_A678_;
  assign new_A71_ = new_A611_;
  assign new_A70_ = new_A544_;
  assign new_A69_ = new_A477_;
  assign new_A68_ = new_A413_;
  assign new_A1_ = new_A744_;
  assign new_A2_ = new_A677_;
  assign new_A3_ = new_A610_;
  assign new_A4_ = new_A543_;
  assign new_A5_ = new_A476_;
  assign new_A6_ = new_A414_;
  assign A7 = new_A14_ & new_A13_;
  assign A8 = new_A16_ | new_A15_;
  assign A9 = new_A18_ | new_A17_;
  assign A10 = new_A20_ & new_A19_;
  assign A11 = new_A20_ & new_A21_;
  assign A12 = new_A13_ | new_A22_;
  assign new_A13_ = new_A2_ | new_A25_;
  assign new_A14_ = new_A24_ | new_A23_;
  assign new_A15_ = new_A29_ & new_A28_;
  assign new_A16_ = new_A27_ & new_A26_;
  assign new_A17_ = new_A32_ | new_A31_;
  assign new_A18_ = new_A27_ & new_A30_;
  assign new_A19_ = new_A2_ | new_A35_;
  assign new_A20_ = new_A34_ | new_A33_;
  assign new_A21_ = new_A37_ | new_A36_;
  assign new_A22_ = ~new_A13_ & new_A39_;
  assign new_A23_ = ~new_A15_ & new_A27_;
  assign new_A24_ = new_A15_ & ~new_A27_;
  assign new_A25_ = new_A1_ & ~new_A2_;
  assign new_A26_ = ~new_A48_ | ~new_A49_;
  assign new_A27_ = new_A41_ | new_A43_;
  assign new_A28_ = new_A51_ | new_A50_;
  assign new_A29_ = new_A45_ | new_A44_;
  assign new_A30_ = ~new_A53_ | ~new_A52_;
  assign new_A31_ = ~new_A54_ & new_A55_;
  assign new_A32_ = new_A54_ & ~new_A55_;
  assign new_A33_ = ~new_A1_ & new_A2_;
  assign new_A34_ = new_A1_ & ~new_A2_;
  assign new_A35_ = ~new_A17_ | new_A27_;
  assign new_A36_ = new_A17_ & new_A27_;
  assign new_A37_ = ~new_A17_ & ~new_A27_;
  assign new_A38_ = new_A59_ | new_A58_;
  assign new_A39_ = new_A5_ | new_A38_;
  assign new_A40_ = new_A63_ | new_A62_;
  assign new_A41_ = ~new_A5_ & new_A40_;
  assign new_A42_ = new_A61_ | new_A60_;
  assign new_A43_ = new_A5_ & new_A42_;
  assign new_A44_ = new_A3_ & ~new_A13_;
  assign new_A45_ = ~new_A3_ & new_A13_;
  assign new_A46_ = ~new_A2_ | ~new_A27_;
  assign new_A47_ = new_A13_ & new_A46_;
  assign new_A48_ = ~new_A13_ & ~new_A47_;
  assign new_A49_ = new_A13_ | new_A46_;
  assign new_A50_ = ~new_A3_ & new_A4_;
  assign new_A51_ = new_A3_ & ~new_A4_;
  assign new_A52_ = new_A20_ | new_A57_;
  assign new_A53_ = ~new_A20_ & ~new_A56_;
  assign new_A54_ = new_A3_ | new_A20_;
  assign new_A55_ = new_A3_ | new_A4_;
  assign new_A56_ = new_A20_ & new_A57_;
  assign new_A57_ = ~new_A2_ | ~new_A27_;
  assign new_A58_ = new_A35_ & new_A55_;
  assign new_A59_ = ~new_A35_ & ~new_A55_;
  assign new_A60_ = new_A64_ | new_A65_;
  assign new_A61_ = ~new_A6_ & new_A20_;
  assign new_A62_ = new_A66_ | new_A67_;
  assign new_A63_ = new_A6_ & new_A20_;
  assign new_A64_ = ~new_A6_ & ~new_A20_;
  assign new_A65_ = new_A6_ & ~new_A20_;
  assign new_A66_ = new_A6_ & ~new_A20_;
  assign new_A67_ = ~new_A6_ & new_A20_;
endmodule


