module top ( clock, 
    p_10, p_12, p_11, pclk, p_9, p_8, p_7, p_6, p_5, p_4, p_3, p_2, p_1,
    p_40, p_45, p_46, p_47, p_41, p_42, p_43, p_44, p_39  );
  input  clock;
  input  p_10, p_12, p_11, pclk, p_9, p_8, p_7, p_6, p_5, p_4, p_3, p_2,
    p_1;
  output p_40, p_45, p_46, p_47, p_41, p_42, p_43, p_44, p_39;
  reg n_22, n_18, n_19, n_20, n_21, n_14, n_15, n_16, n_17, n_13, n_23,
    n_34, n_24, n_33, n_25, n_36, n_26, n_35, n_27, n_38, n_28, n_37, n_29,
    n_30, n_31, n_32;
  wire new_n101_1_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_1_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_1_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_1_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_1_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_1_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_1_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_1_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_1_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_1_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_1_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_1_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_1_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_1_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_1_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n536_,
    new_n537_, new_n539_, new_n540_, new_n542_, new_n543_, new_n545_,
    new_n546_, new_n548_, new_n549_, new_n551_, new_n552_, new_n554_,
    new_n555_, new_n557_, new_n558_, new_n560_, new_n561_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n569_, new_n570_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n578_,
    new_n579_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n587_, new_n588_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n634_, new_n635_, n46, n51, n56, n61, n66, n71, n76,
    n81, n86, n91, n96, n101, n106, n111, n116, n121, n126, n131, n136,
    n141, n146, n151, n156, n161, n166, n171;
  assign new_n101_1_ = ~p_3 & p_2;
  assign new_n102_ = ~p_1 & new_n101_1_;
  assign new_n103_ = ~n_36 & ~n_37;
  assign new_n104_ = ~n_35 & new_n103_;
  assign new_n105_ = ~n_34 & new_n104_;
  assign new_n106_1_ = ~n_33 & new_n105_;
  assign new_n107_ = ~n_32 & new_n106_1_;
  assign new_n108_ = ~n_31 & new_n107_;
  assign new_n109_ = ~n_30 & new_n108_;
  assign new_n110_ = n_29 & new_n109_;
  assign new_n111_1_ = n_28 & new_n110_;
  assign new_n112_ = n_27 & new_n111_1_;
  assign new_n113_ = n_26 & new_n112_;
  assign new_n114_ = n_25 & new_n113_;
  assign new_n115_ = n_24 & new_n114_;
  assign new_n116_1_ = n_23 & new_n115_;
  assign new_n117_ = n_22 & new_n116_1_;
  assign new_n118_ = new_n102_ & new_n117_;
  assign new_n119_ = n_21 & n_38;
  assign new_n120_ = ~n_21 & ~n_38;
  assign new_n121_1_ = ~new_n119_ & ~new_n120_;
  assign new_n122_ = new_n118_ & ~new_n121_1_;
  assign new_n123_ = n_32 & ~new_n122_;
  assign new_n124_ = new_n102_ & new_n123_;
  assign new_n125_ = n_30 & ~new_n122_;
  assign new_n126_1_ = new_n102_ & new_n125_;
  assign new_n127_ = ~p_4 & new_n126_1_;
  assign new_n128_ = p_4 & ~new_n126_1_;
  assign new_n129_ = ~new_n127_ & ~new_n128_;
  assign new_n130_ = p_4 & ~new_n129_;
  assign new_n131_1_ = n_31 & ~new_n122_;
  assign new_n132_ = new_n102_ & new_n131_1_;
  assign new_n133_ = ~p_5 & new_n132_;
  assign new_n134_ = p_5 & ~new_n132_;
  assign new_n135_ = ~new_n133_ & ~new_n134_;
  assign new_n136_1_ = new_n130_ & new_n135_;
  assign new_n137_ = p_5 & ~new_n135_;
  assign new_n138_ = ~new_n136_1_ & ~new_n137_;
  assign new_n139_ = ~p_6 & new_n124_;
  assign new_n140_ = p_6 & ~new_n124_;
  assign new_n141_1_ = ~new_n139_ & ~new_n140_;
  assign new_n142_ = ~new_n138_ & new_n141_1_;
  assign new_n143_ = p_6 & ~new_n141_1_;
  assign new_n144_ = ~new_n142_ & ~new_n143_;
  assign new_n145_ = n_33 & ~new_n122_;
  assign new_n146_1_ = new_n102_ & new_n145_;
  assign new_n147_ = ~p_7 & new_n146_1_;
  assign new_n148_ = p_7 & ~new_n146_1_;
  assign new_n149_ = ~new_n147_ & ~new_n148_;
  assign new_n150_ = ~new_n144_ & new_n149_;
  assign new_n151_1_ = p_7 & ~new_n149_;
  assign new_n152_ = ~new_n150_ & ~new_n151_1_;
  assign new_n153_ = n_34 & ~new_n122_;
  assign new_n154_ = new_n102_ & new_n153_;
  assign new_n155_ = ~p_8 & new_n154_;
  assign new_n156_1_ = p_8 & ~new_n154_;
  assign new_n157_ = ~new_n155_ & ~new_n156_1_;
  assign new_n158_ = ~new_n152_ & new_n157_;
  assign new_n159_ = p_8 & ~new_n157_;
  assign new_n160_ = ~new_n158_ & ~new_n159_;
  assign new_n161_1_ = n_35 & ~new_n122_;
  assign new_n162_ = new_n102_ & new_n161_1_;
  assign new_n163_ = ~p_9 & new_n162_;
  assign new_n164_ = p_9 & ~new_n162_;
  assign new_n165_ = ~new_n163_ & ~new_n164_;
  assign new_n166_1_ = ~new_n160_ & new_n165_;
  assign new_n167_ = p_9 & ~new_n165_;
  assign new_n168_ = ~new_n166_1_ & ~new_n167_;
  assign new_n169_ = n_36 & ~new_n122_;
  assign new_n170_ = new_n102_ & new_n169_;
  assign new_n171_1_ = ~p_10 & new_n170_;
  assign new_n172_ = p_10 & ~new_n170_;
  assign new_n173_ = ~new_n171_1_ & ~new_n172_;
  assign new_n174_ = ~new_n168_ & new_n173_;
  assign new_n175_ = p_10 & ~new_n173_;
  assign new_n176_ = ~new_n174_ & ~new_n175_;
  assign new_n177_ = n_37 & ~new_n122_;
  assign new_n178_ = new_n102_ & new_n177_;
  assign new_n179_ = ~p_11 & new_n178_;
  assign new_n180_ = p_11 & ~new_n178_;
  assign new_n181_ = ~new_n179_ & ~new_n180_;
  assign new_n182_ = ~new_n176_ & new_n181_;
  assign new_n183_ = p_11 & ~new_n181_;
  assign new_n184_ = ~new_n182_ & ~new_n183_;
  assign new_n185_ = ~new_n120_ & ~new_n122_;
  assign new_n186_ = new_n102_ & new_n185_;
  assign new_n187_ = ~p_12 & new_n186_;
  assign new_n188_ = p_12 & ~new_n186_;
  assign new_n189_ = ~new_n187_ & ~new_n188_;
  assign new_n190_ = ~new_n184_ & new_n189_;
  assign new_n191_ = p_12 & ~new_n189_;
  assign new_n192_ = ~new_n190_ & ~new_n191_;
  assign new_n193_ = new_n102_ & ~new_n192_;
  assign new_n194_ = new_n124_ & ~new_n193_;
  assign new_n195_ = p_6 & new_n193_;
  assign new_n196_ = ~new_n194_ & ~new_n195_;
  assign new_n197_ = new_n102_ & ~new_n196_;
  assign new_n198_ = n_22 & ~new_n122_;
  assign new_n199_ = ~new_n122_ & ~new_n198_;
  assign new_n200_ = new_n102_ & ~new_n199_;
  assign new_n201_ = ~p_4 & new_n200_;
  assign new_n202_ = p_4 & ~new_n200_;
  assign new_n203_ = ~new_n201_ & ~new_n202_;
  assign new_n204_ = p_4 & ~new_n203_;
  assign new_n205_ = n_23 & ~new_n122_;
  assign new_n206_ = ~new_n122_ & ~new_n205_;
  assign new_n207_ = new_n102_ & ~new_n206_;
  assign new_n208_ = ~p_5 & new_n207_;
  assign new_n209_ = p_5 & ~new_n207_;
  assign new_n210_ = ~new_n208_ & ~new_n209_;
  assign new_n211_ = new_n204_ & new_n210_;
  assign new_n212_ = p_5 & ~new_n210_;
  assign new_n213_ = ~new_n211_ & ~new_n212_;
  assign new_n214_ = n_24 & ~new_n122_;
  assign new_n215_ = ~new_n122_ & ~new_n214_;
  assign new_n216_ = new_n102_ & ~new_n215_;
  assign new_n217_ = ~p_6 & new_n216_;
  assign new_n218_ = p_6 & ~new_n216_;
  assign new_n219_ = ~new_n217_ & ~new_n218_;
  assign new_n220_ = ~new_n213_ & new_n219_;
  assign new_n221_ = p_6 & ~new_n219_;
  assign new_n222_ = ~new_n220_ & ~new_n221_;
  assign new_n223_ = n_25 & ~new_n122_;
  assign new_n224_ = ~new_n122_ & ~new_n223_;
  assign new_n225_ = new_n102_ & ~new_n224_;
  assign new_n226_ = ~p_7 & new_n225_;
  assign new_n227_ = p_7 & ~new_n225_;
  assign new_n228_ = ~new_n226_ & ~new_n227_;
  assign new_n229_ = ~new_n222_ & new_n228_;
  assign new_n230_ = p_7 & ~new_n228_;
  assign new_n231_ = ~new_n229_ & ~new_n230_;
  assign new_n232_ = n_26 & ~new_n122_;
  assign new_n233_ = ~new_n122_ & ~new_n232_;
  assign new_n234_ = new_n102_ & ~new_n233_;
  assign new_n235_ = ~p_8 & new_n234_;
  assign new_n236_ = p_8 & ~new_n234_;
  assign new_n237_ = ~new_n235_ & ~new_n236_;
  assign new_n238_ = ~new_n231_ & new_n237_;
  assign new_n239_ = p_8 & ~new_n237_;
  assign new_n240_ = ~new_n238_ & ~new_n239_;
  assign new_n241_ = n_27 & ~new_n122_;
  assign new_n242_ = ~new_n122_ & ~new_n241_;
  assign new_n243_ = new_n102_ & ~new_n242_;
  assign new_n244_ = ~p_9 & new_n243_;
  assign new_n245_ = p_9 & ~new_n243_;
  assign new_n246_ = ~new_n244_ & ~new_n245_;
  assign new_n247_ = ~new_n240_ & new_n246_;
  assign new_n248_ = p_9 & ~new_n246_;
  assign new_n249_ = ~new_n247_ & ~new_n248_;
  assign new_n250_ = n_28 & ~new_n122_;
  assign new_n251_ = ~new_n122_ & ~new_n250_;
  assign new_n252_ = new_n102_ & ~new_n251_;
  assign new_n253_ = ~p_10 & new_n252_;
  assign new_n254_ = p_10 & ~new_n252_;
  assign new_n255_ = ~new_n253_ & ~new_n254_;
  assign new_n256_ = ~new_n249_ & new_n255_;
  assign new_n257_ = p_10 & ~new_n255_;
  assign new_n258_ = ~new_n256_ & ~new_n257_;
  assign new_n259_ = n_29 & ~new_n122_;
  assign new_n260_ = ~new_n122_ & ~new_n259_;
  assign new_n261_ = new_n102_ & ~new_n260_;
  assign new_n262_ = ~p_11 & new_n261_;
  assign new_n263_ = p_11 & ~new_n261_;
  assign new_n264_ = ~new_n262_ & ~new_n263_;
  assign new_n265_ = ~new_n258_ & new_n264_;
  assign new_n266_ = p_11 & ~new_n264_;
  assign new_n267_ = ~new_n265_ & ~new_n266_;
  assign new_n268_ = new_n119_ & ~new_n122_;
  assign new_n269_ = ~new_n122_ & ~new_n268_;
  assign new_n270_ = new_n102_ & ~new_n269_;
  assign new_n271_ = ~p_12 & new_n270_;
  assign new_n272_ = p_12 & ~new_n270_;
  assign new_n273_ = ~new_n271_ & ~new_n272_;
  assign new_n274_ = ~new_n267_ & new_n273_;
  assign new_n275_ = p_12 & ~new_n273_;
  assign new_n276_ = ~new_n274_ & ~new_n275_;
  assign new_n277_ = new_n102_ & ~new_n276_;
  assign new_n278_ = p_6 & ~new_n277_;
  assign new_n279_ = new_n216_ & new_n277_;
  assign new_n280_ = ~new_n278_ & ~new_n279_;
  assign new_n281_ = new_n102_ & ~new_n280_;
  assign new_n282_ = p_5 & ~new_n277_;
  assign new_n283_ = new_n207_ & new_n277_;
  assign new_n284_ = ~new_n282_ & ~new_n283_;
  assign new_n285_ = new_n102_ & ~new_n284_;
  assign new_n286_ = new_n132_ & ~new_n193_;
  assign new_n287_ = p_5 & new_n193_;
  assign new_n288_ = ~new_n286_ & ~new_n287_;
  assign new_n289_ = new_n102_ & ~new_n288_;
  assign new_n290_ = new_n285_ & new_n289_;
  assign new_n291_ = p_4 & ~new_n277_;
  assign new_n292_ = new_n200_ & new_n277_;
  assign new_n293_ = ~new_n291_ & ~new_n292_;
  assign new_n294_ = new_n102_ & ~new_n293_;
  assign new_n295_ = new_n126_1_ & ~new_n193_;
  assign new_n296_ = p_4 & new_n193_;
  assign new_n297_ = ~new_n295_ & ~new_n296_;
  assign new_n298_ = new_n102_ & ~new_n297_;
  assign new_n299_ = new_n294_ & new_n298_;
  assign new_n300_ = new_n289_ & new_n299_;
  assign new_n301_ = new_n285_ & new_n299_;
  assign new_n302_ = ~new_n290_ & ~new_n300_;
  assign new_n303_ = ~new_n301_ & new_n302_;
  assign new_n304_ = new_n197_ & new_n281_;
  assign new_n305_ = ~new_n303_ & new_n304_;
  assign new_n306_ = ~new_n197_ & new_n281_;
  assign new_n307_ = new_n303_ & new_n306_;
  assign new_n308_ = new_n197_ & ~new_n281_;
  assign new_n309_ = new_n303_ & new_n308_;
  assign new_n310_ = ~new_n197_ & ~new_n281_;
  assign new_n311_ = ~new_n303_ & new_n310_;
  assign new_n312_ = ~new_n305_ & ~new_n307_;
  assign new_n313_ = ~new_n309_ & ~new_n311_;
  assign new_n314_ = new_n312_ & new_n313_;
  assign new_n315_ = ~p_3 & ~new_n314_;
  assign new_n316_ = p_5 & p_3;
  assign new_n317_ = ~new_n315_ & ~new_n316_;
  assign new_n318_ = p_2 & ~new_n317_;
  assign new_n319_ = ~p_2 & n_14;
  assign new_n320_ = ~new_n318_ & ~new_n319_;
  assign p_40 = ~p_1 & ~new_n320_;
  assign new_n322_ = new_n178_ & ~new_n193_;
  assign new_n323_ = p_11 & new_n193_;
  assign new_n324_ = ~new_n322_ & ~new_n323_;
  assign new_n325_ = new_n102_ & ~new_n324_;
  assign new_n326_ = p_11 & ~new_n277_;
  assign new_n327_ = new_n261_ & new_n277_;
  assign new_n328_ = ~new_n326_ & ~new_n327_;
  assign new_n329_ = new_n102_ & ~new_n328_;
  assign new_n330_ = p_10 & ~new_n277_;
  assign new_n331_ = new_n252_ & new_n277_;
  assign new_n332_ = ~new_n330_ & ~new_n331_;
  assign new_n333_ = new_n102_ & ~new_n332_;
  assign new_n334_ = new_n170_ & ~new_n193_;
  assign new_n335_ = p_10 & new_n193_;
  assign new_n336_ = ~new_n334_ & ~new_n335_;
  assign new_n337_ = new_n102_ & ~new_n336_;
  assign new_n338_ = new_n333_ & new_n337_;
  assign new_n339_ = p_9 & ~new_n277_;
  assign new_n340_ = new_n243_ & new_n277_;
  assign new_n341_ = ~new_n339_ & ~new_n340_;
  assign new_n342_ = new_n102_ & ~new_n341_;
  assign new_n343_ = new_n162_ & ~new_n193_;
  assign new_n344_ = p_9 & new_n193_;
  assign new_n345_ = ~new_n343_ & ~new_n344_;
  assign new_n346_ = new_n102_ & ~new_n345_;
  assign new_n347_ = new_n342_ & new_n346_;
  assign new_n348_ = p_8 & ~new_n277_;
  assign new_n349_ = new_n234_ & new_n277_;
  assign new_n350_ = ~new_n348_ & ~new_n349_;
  assign new_n351_ = new_n102_ & ~new_n350_;
  assign new_n352_ = new_n154_ & ~new_n193_;
  assign new_n353_ = p_8 & new_n193_;
  assign new_n354_ = ~new_n352_ & ~new_n353_;
  assign new_n355_ = new_n102_ & ~new_n354_;
  assign new_n356_ = new_n351_ & new_n355_;
  assign new_n357_ = p_7 & ~new_n277_;
  assign new_n358_ = new_n225_ & new_n277_;
  assign new_n359_ = ~new_n357_ & ~new_n358_;
  assign new_n360_ = new_n102_ & ~new_n359_;
  assign new_n361_ = new_n146_1_ & ~new_n193_;
  assign new_n362_ = p_7 & new_n193_;
  assign new_n363_ = ~new_n361_ & ~new_n362_;
  assign new_n364_ = new_n102_ & ~new_n363_;
  assign new_n365_ = new_n360_ & new_n364_;
  assign new_n366_ = new_n197_ & ~new_n303_;
  assign new_n367_ = new_n281_ & ~new_n303_;
  assign new_n368_ = ~new_n304_ & ~new_n366_;
  assign new_n369_ = ~new_n367_ & new_n368_;
  assign new_n370_ = new_n364_ & ~new_n369_;
  assign new_n371_ = new_n360_ & ~new_n369_;
  assign new_n372_ = ~new_n365_ & ~new_n370_;
  assign new_n373_ = ~new_n371_ & new_n372_;
  assign new_n374_ = new_n355_ & ~new_n373_;
  assign new_n375_ = new_n351_ & ~new_n373_;
  assign new_n376_ = ~new_n356_ & ~new_n374_;
  assign new_n377_ = ~new_n375_ & new_n376_;
  assign new_n378_ = new_n346_ & ~new_n377_;
  assign new_n379_ = new_n342_ & ~new_n377_;
  assign new_n380_ = ~new_n347_ & ~new_n378_;
  assign new_n381_ = ~new_n379_ & new_n380_;
  assign new_n382_ = new_n337_ & ~new_n381_;
  assign new_n383_ = new_n333_ & ~new_n381_;
  assign new_n384_ = ~new_n338_ & ~new_n382_;
  assign new_n385_ = ~new_n383_ & new_n384_;
  assign new_n386_ = new_n325_ & new_n329_;
  assign new_n387_ = ~new_n385_ & new_n386_;
  assign new_n388_ = ~new_n325_ & new_n329_;
  assign new_n389_ = new_n385_ & new_n388_;
  assign new_n390_ = new_n325_ & ~new_n329_;
  assign new_n391_ = new_n385_ & new_n390_;
  assign new_n392_ = ~new_n325_ & ~new_n329_;
  assign new_n393_ = ~new_n385_ & new_n392_;
  assign new_n394_ = ~new_n387_ & ~new_n389_;
  assign new_n395_ = ~new_n391_ & ~new_n393_;
  assign new_n396_ = new_n394_ & new_n395_;
  assign new_n397_ = ~p_3 & ~new_n396_;
  assign new_n398_ = p_10 & p_3;
  assign new_n399_ = ~new_n397_ & ~new_n398_;
  assign new_n400_ = p_2 & ~new_n399_;
  assign new_n401_ = ~p_2 & n_19;
  assign new_n402_ = ~new_n400_ & ~new_n401_;
  assign p_45 = ~p_1 & ~new_n402_;
  assign new_n404_ = new_n186_ & ~new_n193_;
  assign new_n405_ = p_12 & new_n193_;
  assign new_n406_ = ~new_n404_ & ~new_n405_;
  assign new_n407_ = new_n102_ & ~new_n406_;
  assign new_n408_ = p_12 & ~new_n277_;
  assign new_n409_ = new_n270_ & new_n277_;
  assign new_n410_ = ~new_n408_ & ~new_n409_;
  assign new_n411_ = new_n102_ & ~new_n410_;
  assign new_n412_ = new_n325_ & ~new_n385_;
  assign new_n413_ = new_n329_ & ~new_n385_;
  assign new_n414_ = ~new_n386_ & ~new_n412_;
  assign new_n415_ = ~new_n413_ & new_n414_;
  assign new_n416_ = new_n407_ & new_n411_;
  assign new_n417_ = ~new_n415_ & new_n416_;
  assign new_n418_ = ~new_n407_ & new_n411_;
  assign new_n419_ = new_n415_ & new_n418_;
  assign new_n420_ = new_n407_ & ~new_n411_;
  assign new_n421_ = new_n415_ & new_n420_;
  assign new_n422_ = ~new_n407_ & ~new_n411_;
  assign new_n423_ = ~new_n415_ & new_n422_;
  assign new_n424_ = ~new_n417_ & ~new_n419_;
  assign new_n425_ = ~new_n421_ & ~new_n423_;
  assign new_n426_ = new_n424_ & new_n425_;
  assign new_n427_ = ~p_3 & ~new_n426_;
  assign new_n428_ = p_11 & p_3;
  assign new_n429_ = ~new_n427_ & ~new_n428_;
  assign new_n430_ = p_2 & ~new_n429_;
  assign new_n431_ = ~p_2 & n_20;
  assign new_n432_ = ~new_n430_ & ~new_n431_;
  assign p_46 = ~p_1 & ~new_n432_;
  assign new_n434_ = new_n407_ & ~new_n415_;
  assign new_n435_ = new_n411_ & ~new_n415_;
  assign new_n436_ = ~new_n416_ & ~new_n434_;
  assign new_n437_ = ~new_n435_ & new_n436_;
  assign new_n438_ = ~p_3 & ~new_n437_;
  assign new_n439_ = p_12 & p_3;
  assign new_n440_ = ~new_n438_ & ~new_n439_;
  assign new_n441_ = p_2 & ~new_n440_;
  assign new_n442_ = ~p_2 & n_21;
  assign new_n443_ = ~new_n441_ & ~new_n442_;
  assign p_47 = ~p_1 & ~new_n443_;
  assign new_n445_ = new_n365_ & ~new_n369_;
  assign new_n446_ = new_n360_ & ~new_n364_;
  assign new_n447_ = new_n369_ & new_n446_;
  assign new_n448_ = ~new_n360_ & new_n364_;
  assign new_n449_ = new_n369_ & new_n448_;
  assign new_n450_ = ~new_n360_ & ~new_n364_;
  assign new_n451_ = ~new_n369_ & new_n450_;
  assign new_n452_ = ~new_n445_ & ~new_n447_;
  assign new_n453_ = ~new_n449_ & ~new_n451_;
  assign new_n454_ = new_n452_ & new_n453_;
  assign new_n455_ = ~p_3 & ~new_n454_;
  assign new_n456_ = p_6 & p_3;
  assign new_n457_ = ~new_n455_ & ~new_n456_;
  assign new_n458_ = p_2 & ~new_n457_;
  assign new_n459_ = ~p_2 & n_15;
  assign new_n460_ = ~new_n458_ & ~new_n459_;
  assign p_41 = ~p_1 & ~new_n460_;
  assign new_n462_ = new_n356_ & ~new_n373_;
  assign new_n463_ = new_n351_ & ~new_n355_;
  assign new_n464_ = new_n373_ & new_n463_;
  assign new_n465_ = ~new_n351_ & new_n355_;
  assign new_n466_ = new_n373_ & new_n465_;
  assign new_n467_ = ~new_n351_ & ~new_n355_;
  assign new_n468_ = ~new_n373_ & new_n467_;
  assign new_n469_ = ~new_n462_ & ~new_n464_;
  assign new_n470_ = ~new_n466_ & ~new_n468_;
  assign new_n471_ = new_n469_ & new_n470_;
  assign new_n472_ = ~p_3 & ~new_n471_;
  assign new_n473_ = p_7 & p_3;
  assign new_n474_ = ~new_n472_ & ~new_n473_;
  assign new_n475_ = p_2 & ~new_n474_;
  assign new_n476_ = ~p_2 & n_16;
  assign new_n477_ = ~new_n475_ & ~new_n476_;
  assign p_42 = ~p_1 & ~new_n477_;
  assign new_n479_ = new_n347_ & ~new_n377_;
  assign new_n480_ = new_n342_ & ~new_n346_;
  assign new_n481_ = new_n377_ & new_n480_;
  assign new_n482_ = ~new_n342_ & new_n346_;
  assign new_n483_ = new_n377_ & new_n482_;
  assign new_n484_ = ~new_n342_ & ~new_n346_;
  assign new_n485_ = ~new_n377_ & new_n484_;
  assign new_n486_ = ~new_n479_ & ~new_n481_;
  assign new_n487_ = ~new_n483_ & ~new_n485_;
  assign new_n488_ = new_n486_ & new_n487_;
  assign new_n489_ = ~p_3 & ~new_n488_;
  assign new_n490_ = p_8 & p_3;
  assign new_n491_ = ~new_n489_ & ~new_n490_;
  assign new_n492_ = p_2 & ~new_n491_;
  assign new_n493_ = ~p_2 & n_17;
  assign new_n494_ = ~new_n492_ & ~new_n493_;
  assign p_43 = ~p_1 & ~new_n494_;
  assign new_n496_ = new_n338_ & ~new_n381_;
  assign new_n497_ = new_n333_ & ~new_n337_;
  assign new_n498_ = new_n381_ & new_n497_;
  assign new_n499_ = ~new_n333_ & new_n337_;
  assign new_n500_ = new_n381_ & new_n499_;
  assign new_n501_ = ~new_n333_ & ~new_n337_;
  assign new_n502_ = ~new_n381_ & new_n501_;
  assign new_n503_ = ~new_n496_ & ~new_n498_;
  assign new_n504_ = ~new_n500_ & ~new_n502_;
  assign new_n505_ = new_n503_ & new_n504_;
  assign new_n506_ = ~p_3 & ~new_n505_;
  assign new_n507_ = p_9 & p_3;
  assign new_n508_ = ~new_n506_ & ~new_n507_;
  assign new_n509_ = p_2 & ~new_n508_;
  assign new_n510_ = ~p_2 & n_18;
  assign new_n511_ = ~new_n509_ & ~new_n510_;
  assign p_44 = ~p_1 & ~new_n511_;
  assign new_n513_ = new_n290_ & new_n299_;
  assign new_n514_ = new_n285_ & ~new_n289_;
  assign new_n515_ = ~new_n299_ & new_n514_;
  assign new_n516_ = ~new_n285_ & new_n289_;
  assign new_n517_ = ~new_n299_ & new_n516_;
  assign new_n518_ = ~new_n285_ & ~new_n289_;
  assign new_n519_ = new_n299_ & new_n518_;
  assign new_n520_ = ~new_n513_ & ~new_n515_;
  assign new_n521_ = ~new_n517_ & ~new_n519_;
  assign new_n522_ = new_n520_ & new_n521_;
  assign new_n523_ = ~p_3 & ~new_n522_;
  assign new_n524_ = p_4 & p_3;
  assign new_n525_ = ~new_n523_ & ~new_n524_;
  assign new_n526_ = p_2 & ~new_n525_;
  assign new_n527_ = ~p_2 & n_13;
  assign new_n528_ = ~new_n526_ & ~new_n527_;
  assign p_39 = ~p_1 & ~new_n528_;
  assign new_n530_ = ~p_3 & new_n294_;
  assign new_n531_ = ~p_3 & ~new_n530_;
  assign new_n532_ = p_2 & ~new_n531_;
  assign new_n533_ = p_2 & ~new_n532_;
  assign new_n534_ = ~p_1 & ~new_n533_;
  assign n46 = p_1 | new_n534_;
  assign new_n536_ = p_9 & p_2;
  assign new_n537_ = ~new_n510_ & ~new_n536_;
  assign n51 = ~p_1 & ~new_n537_;
  assign new_n539_ = p_10 & p_2;
  assign new_n540_ = ~new_n401_ & ~new_n539_;
  assign n56 = ~p_1 & ~new_n540_;
  assign new_n542_ = p_11 & p_2;
  assign new_n543_ = ~new_n431_ & ~new_n542_;
  assign n61 = ~p_1 & ~new_n543_;
  assign new_n545_ = p_12 & p_2;
  assign new_n546_ = ~new_n442_ & ~new_n545_;
  assign n66 = ~p_1 & ~new_n546_;
  assign new_n548_ = p_5 & p_2;
  assign new_n549_ = ~new_n319_ & ~new_n548_;
  assign n71 = ~p_1 & ~new_n549_;
  assign new_n551_ = p_6 & p_2;
  assign new_n552_ = ~new_n459_ & ~new_n551_;
  assign n76 = ~p_1 & ~new_n552_;
  assign new_n554_ = p_7 & p_2;
  assign new_n555_ = ~new_n476_ & ~new_n554_;
  assign n81 = ~p_1 & ~new_n555_;
  assign new_n557_ = p_8 & p_2;
  assign new_n558_ = ~new_n493_ & ~new_n557_;
  assign n86 = ~p_1 & ~new_n558_;
  assign new_n560_ = p_4 & p_2;
  assign new_n561_ = ~new_n527_ & ~new_n560_;
  assign n91 = ~p_1 & ~new_n561_;
  assign new_n563_ = ~p_3 & new_n285_;
  assign new_n564_ = ~p_3 & ~new_n563_;
  assign new_n565_ = p_2 & ~new_n564_;
  assign new_n566_ = p_2 & ~new_n565_;
  assign new_n567_ = ~p_1 & ~new_n566_;
  assign n96 = p_1 | new_n567_;
  assign new_n569_ = ~p_3 & new_n355_;
  assign new_n570_ = p_2 & new_n569_;
  assign n101 = ~p_1 & new_n570_;
  assign new_n572_ = ~p_3 & new_n281_;
  assign new_n573_ = ~p_3 & ~new_n572_;
  assign new_n574_ = p_2 & ~new_n573_;
  assign new_n575_ = p_2 & ~new_n574_;
  assign new_n576_ = ~p_1 & ~new_n575_;
  assign n106 = p_1 | new_n576_;
  assign new_n578_ = ~p_3 & new_n364_;
  assign new_n579_ = p_2 & new_n578_;
  assign n111 = ~p_1 & new_n579_;
  assign new_n581_ = ~p_3 & new_n360_;
  assign new_n582_ = ~p_3 & ~new_n581_;
  assign new_n583_ = p_2 & ~new_n582_;
  assign new_n584_ = p_2 & ~new_n583_;
  assign new_n585_ = ~p_1 & ~new_n584_;
  assign n116 = p_1 | new_n585_;
  assign new_n587_ = ~p_3 & new_n337_;
  assign new_n588_ = p_2 & new_n587_;
  assign n121 = ~p_1 & new_n588_;
  assign new_n590_ = ~p_3 & new_n351_;
  assign new_n591_ = ~p_3 & ~new_n590_;
  assign new_n592_ = p_2 & ~new_n591_;
  assign new_n593_ = p_2 & ~new_n592_;
  assign new_n594_ = ~p_1 & ~new_n593_;
  assign n126 = p_1 | new_n594_;
  assign new_n596_ = ~p_3 & new_n346_;
  assign new_n597_ = p_2 & new_n596_;
  assign n131 = ~p_1 & new_n597_;
  assign new_n599_ = ~p_3 & new_n342_;
  assign new_n600_ = ~p_3 & ~new_n599_;
  assign new_n601_ = p_2 & ~new_n600_;
  assign new_n602_ = p_2 & ~new_n601_;
  assign new_n603_ = ~p_1 & ~new_n602_;
  assign n136 = p_1 | new_n603_;
  assign new_n605_ = p_12 & new_n411_;
  assign new_n606_ = ~p_12 & new_n407_;
  assign new_n607_ = ~new_n605_ & ~new_n606_;
  assign new_n608_ = ~p_3 & ~new_n607_;
  assign new_n609_ = ~new_n439_ & ~new_n608_;
  assign new_n610_ = p_2 & ~new_n609_;
  assign new_n611_ = ~new_n442_ & ~new_n610_;
  assign n141 = ~p_1 & ~new_n611_;
  assign new_n613_ = ~p_3 & new_n333_;
  assign new_n614_ = ~p_3 & ~new_n613_;
  assign new_n615_ = p_2 & ~new_n614_;
  assign new_n616_ = p_2 & ~new_n615_;
  assign new_n617_ = ~p_1 & ~new_n616_;
  assign n146 = p_1 | new_n617_;
  assign new_n619_ = ~p_3 & new_n325_;
  assign new_n620_ = p_2 & new_n619_;
  assign n151 = ~p_1 & new_n620_;
  assign new_n622_ = ~p_3 & new_n329_;
  assign new_n623_ = ~p_3 & ~new_n622_;
  assign new_n624_ = p_2 & ~new_n623_;
  assign new_n625_ = p_2 & ~new_n624_;
  assign new_n626_ = ~p_1 & ~new_n625_;
  assign n156 = p_1 | new_n626_;
  assign new_n628_ = ~p_3 & new_n298_;
  assign new_n629_ = p_2 & new_n628_;
  assign n161 = ~p_1 & new_n629_;
  assign new_n631_ = ~p_3 & new_n289_;
  assign new_n632_ = p_2 & new_n631_;
  assign n166 = ~p_1 & new_n632_;
  assign new_n634_ = ~p_3 & new_n197_;
  assign new_n635_ = p_2 & new_n634_;
  assign n171 = ~p_1 & new_n635_;
  always @ (posedge clock) begin
    n_22 <= n46;
    n_18 <= n51;
    n_19 <= n56;
    n_20 <= n61;
    n_21 <= n66;
    n_14 <= n71;
    n_15 <= n76;
    n_16 <= n81;
    n_17 <= n86;
    n_13 <= n91;
    n_23 <= n96;
    n_34 <= n101;
    n_24 <= n106;
    n_33 <= n111;
    n_25 <= n116;
    n_36 <= n121;
    n_26 <= n126;
    n_35 <= n131;
    n_27 <= n136;
    n_38 <= n141;
    n_28 <= n146;
    n_37 <= n151;
    n_29 <= n156;
    n_30 <= n161;
    n_31 <= n166;
    n_32 <= n171;
  end
endmodule

